# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_ls__a311oi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_ls__a311oi_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.760000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.300000 1.350000 3.235000 1.550000 ;
        RECT 2.870000 1.550000 3.235000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.180000 1.315000 1.220000 ;
        RECT 1.085000 1.220000 2.090000 1.550000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.470000 1.220000 0.835000 1.550000 ;
        RECT 0.605000 1.180000 0.835000 1.220000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.447000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485000 1.350000 4.675000 1.780000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.447000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.845000 1.350000 5.175000 1.780000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  0.935400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.555000 0.850000 3.745000 1.010000 ;
        RECT 2.555000 1.010000 5.635000 1.180000 ;
        RECT 3.495000 0.350000 3.745000 0.850000 ;
        RECT 4.685000 0.350000 5.635000 1.010000 ;
        RECT 4.850000 1.950000 5.635000 2.120000 ;
        RECT 4.850000 2.120000 5.020000 2.735000 ;
        RECT 5.405000 1.180000 5.635000 1.950000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.760000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000000 0.000000 5.760000 0.245000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.660000 5.950000 3.520000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.760000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.760000 0.085000 ;
      RECT 0.000000  3.245000 5.760000 3.415000 ;
      RECT 0.170000  1.820000 0.420000 3.245000 ;
      RECT 0.185000  0.350000 0.435000 0.840000 ;
      RECT 0.185000  0.840000 2.235000 1.010000 ;
      RECT 0.185000  1.010000 0.435000 1.050000 ;
      RECT 0.615000  0.085000 0.945000 0.670000 ;
      RECT 0.620000  1.720000 2.700000 1.890000 ;
      RECT 0.620000  1.890000 0.950000 2.980000 ;
      RECT 1.125000  0.330000 1.295000 0.770000 ;
      RECT 1.125000  0.770000 2.235000 0.840000 ;
      RECT 1.150000  2.060000 1.320000 3.245000 ;
      RECT 1.475000  0.350000 3.315000 0.600000 ;
      RECT 1.520000  1.890000 1.850000 2.980000 ;
      RECT 1.905000  1.010000 2.235000 1.050000 ;
      RECT 2.050000  2.060000 2.330000 3.245000 ;
      RECT 2.530000  1.890000 2.700000 1.950000 ;
      RECT 2.530000  1.950000 4.120000 2.120000 ;
      RECT 2.530000  2.120000 2.700000 2.980000 ;
      RECT 2.900000  2.290000 3.230000 3.245000 ;
      RECT 2.985000  0.600000 3.315000 0.680000 ;
      RECT 3.420000  2.290000 3.755000 2.905000 ;
      RECT 3.420000  2.905000 5.550000 3.075000 ;
      RECT 3.915000  0.085000 4.515000 0.840000 ;
      RECT 3.925000  2.120000 4.120000 2.735000 ;
      RECT 4.320000  1.950000 4.650000 2.905000 ;
      RECT 5.220000  2.290000 5.550000 2.905000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
  END
END sky130_fd_sc_ls__a311oi_2
END LIBRARY
