* File: sky130_fd_sc_ls__decaphe_3.spice
* Created: Wed Sep  2 10:59:47 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__decaphe_3.pex.spice"
.subckt sky130_fd_sc_ls__decaphe_3  VNB VPB VGND VPWR
* 
* VPWR	VPWR
* VGND	VGND
* VPB	VPB
* VNB	VNB
MM1000 N_VGND_M1000_s N_VPWR_M1000_g N_VGND_M1000_s VNB NSHORT L=0.65 W=0.775
+ AD=0.2015 AS=0.2015 PD=2.07 PS=2.07 NRD=0 NRS=0 M=1 R=1.19231 SA=325000
+ SB=325000 A=0.50375 P=2.85 MULT=1
MM1001 N_VPWR_M1001_s N_VGND_M1001_g N_VPWR_M1001_s VPB PSHORT L=0.65 W=1.255
+ AD=0.3263 AS=0.3263 PD=3.03 PS=3.03 NRD=0 NRS=0 M=1 R=1.93077 SA=325000
+ SB=325000 A=0.81575 P=3.81 MULT=1
DX2_noxref VNB VPB NWDIODE A=3.3852 P=7.36
*
.include "sky130_fd_sc_ls__decaphe_3.pxi.spice"
*
.ends
*
*
