* File: sky130_fd_sc_ls__dfxbp_1.pex.spice
* Created: Fri Aug 28 13:16:04 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__DFXBP_1%CLK 1 3 4 6 7 11
c29 11 0 2.6712e-20 $X=0.335 $Y=1.385
c30 4 0 1.73501e-19 $X=0.5 $Y=1.765
r31 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.335
+ $Y=1.385 $X2=0.335 $Y2=1.385
r32 7 11 2.95898 $w=3.68e-07 $l=9.5e-08 $layer=LI1_cond $X=0.24 $Y=1.365
+ $X2=0.335 $Y2=1.365
r33 4 10 70.4572 $w=3.25e-07 $l=4.3589e-07 $layer=POLY_cond $X=0.5 $Y=1.765
+ $X2=0.38 $Y2=1.385
r34 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.5 $Y=1.765 $X2=0.5
+ $Y2=2.4
r35 1 10 38.571 $w=3.25e-07 $l=2.14942e-07 $layer=POLY_cond $X=0.495 $Y=1.22
+ $X2=0.38 $Y2=1.385
r36 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.495 $Y=1.22 $X2=0.495
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__DFXBP_1%A_27_74# 1 2 7 9 10 12 15 18 19 21 22 24 26
+ 30 33 37 41 45 48 49 50 51 53 55 56 59 60 61 62 65 68 70 75 76 78 80 83 84 85
c243 80 0 4.89519e-20 $X=0.965 $Y=1.385
c244 75 0 6.57199e-20 $X=5.55 $Y=0.455
c245 65 0 2.11133e-19 $X=3.285 $Y=1.91
c246 37 0 6.7972e-20 $X=5.64 $Y=1.3
c247 33 0 5.93116e-20 $X=5.34 $Y=1.97
c248 30 0 1.76992e-19 $X=5.64 $Y=0.94
c249 26 0 3.57825e-20 $X=5.34 $Y=1.895
c250 18 0 1.34618e-19 $X=3.175 $Y=2.375
c251 15 0 4.57052e-20 $X=3.015 $Y=0.805
c252 10 0 2.6712e-20 $X=1.135 $Y=1.22
c253 7 0 8.80023e-20 $X=0.95 $Y=1.765
r254 87 89 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=3.015 $Y=1.91
+ $X2=3.175 $Y2=1.91
r255 84 85 8.63679 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=4.48 $Y=0.52
+ $X2=4.65 $Y2=0.52
r256 80 82 8.7366 $w=4.18e-07 $l=1.65e-07 $layer=LI1_cond $X=0.88 $Y=1.385
+ $X2=0.88 $Y2=1.55
r257 80 81 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.965
+ $Y=1.385 $X2=0.965 $Y2=1.385
r258 76 94 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.55 $Y=0.455
+ $X2=5.55 $Y2=0.62
r259 75 85 31.4303 $w=3.28e-07 $l=9e-07 $layer=LI1_cond $X=5.55 $Y=0.455
+ $X2=4.65 $Y2=0.455
r260 75 76 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.55
+ $Y=0.455 $X2=5.55 $Y2=0.455
r261 72 83 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.655 $Y=0.665
+ $X2=3.57 $Y2=0.665
r262 72 84 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=3.655 $Y=0.665
+ $X2=4.48 $Y2=0.665
r263 69 83 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.57 $Y=0.75
+ $X2=3.57 $Y2=0.665
r264 69 70 65.2406 $w=1.68e-07 $l=1e-06 $layer=LI1_cond $X=3.57 $Y=0.75 $X2=3.57
+ $Y2=1.75
r265 68 83 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.57 $Y=0.58
+ $X2=3.57 $Y2=0.665
r266 67 68 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=3.57 $Y=0.425
+ $X2=3.57 $Y2=0.58
r267 65 89 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=3.285 $Y=1.91
+ $X2=3.175 $Y2=1.91
r268 64 65 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.285
+ $Y=1.91 $X2=3.285 $Y2=1.91
r269 62 70 7.72402 $w=3.25e-07 $l=2.00035e-07 $layer=LI1_cond $X=3.485 $Y=1.912
+ $X2=3.57 $Y2=1.75
r270 62 64 7.09196 $w=3.23e-07 $l=2e-07 $layer=LI1_cond $X=3.485 $Y=1.912
+ $X2=3.285 $Y2=1.912
r271 60 67 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.485 $Y=0.34
+ $X2=3.57 $Y2=0.425
r272 60 61 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=3.485 $Y=0.34
+ $X2=2.545 $Y2=0.34
r273 58 61 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.46 $Y=0.425
+ $X2=2.545 $Y2=0.34
r274 58 59 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.46 $Y=0.425
+ $X2=2.46 $Y2=0.73
r275 57 78 10.1275 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=1.09 $Y=0.815
+ $X2=0.88 $Y2=0.815
r276 56 59 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.375 $Y=0.815
+ $X2=2.46 $Y2=0.73
r277 56 57 83.8342 $w=1.68e-07 $l=1.285e-06 $layer=LI1_cond $X=2.375 $Y=0.815
+ $X2=1.09 $Y2=0.815
r278 55 82 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.755 $Y=1.72
+ $X2=0.755 $Y2=1.55
r279 53 80 1.23476 $w=4.18e-07 $l=4.5e-08 $layer=LI1_cond $X=0.88 $Y=1.34
+ $X2=0.88 $Y2=1.385
r280 52 78 1.60615 $w=4.2e-07 $l=8.5e-08 $layer=LI1_cond $X=0.88 $Y=0.9 $X2=0.88
+ $Y2=0.815
r281 52 53 12.0732 $w=4.18e-07 $l=4.4e-07 $layer=LI1_cond $X=0.88 $Y=0.9
+ $X2=0.88 $Y2=1.34
r282 50 78 10.1275 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=0.67 $Y=0.815
+ $X2=0.88 $Y2=0.815
r283 50 51 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.67 $Y=0.815
+ $X2=0.445 $Y2=0.815
r284 48 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.67 $Y=1.805
+ $X2=0.755 $Y2=1.72
r285 48 49 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.67 $Y=1.805
+ $X2=0.36 $Y2=1.805
r286 45 51 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=0.73
+ $X2=0.445 $Y2=0.815
r287 45 47 1.84848 $w=3.3e-07 $l=5e-08 $layer=LI1_cond $X=0.28 $Y=0.73 $X2=0.28
+ $Y2=0.68
r288 41 43 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=0.235 $Y=1.985
+ $X2=0.235 $Y2=2.815
r289 39 49 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.235 $Y=1.89
+ $X2=0.36 $Y2=1.805
r290 39 41 4.37928 $w=2.48e-07 $l=9.5e-08 $layer=LI1_cond $X=0.235 $Y=1.89
+ $X2=0.235 $Y2=1.985
r291 35 37 153.83 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=5.34 $Y=1.3 $X2=5.64
+ $Y2=1.3
r292 31 33 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=5.18 $Y=1.97
+ $X2=5.34 $Y2=1.97
r293 30 94 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=5.64 $Y=0.94
+ $X2=5.64 $Y2=0.62
r294 28 37 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.64 $Y=1.225
+ $X2=5.64 $Y2=1.3
r295 28 30 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=5.64 $Y=1.225
+ $X2=5.64 $Y2=0.94
r296 26 33 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.34 $Y=1.895
+ $X2=5.34 $Y2=1.97
r297 25 35 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.34 $Y=1.375
+ $X2=5.34 $Y2=1.3
r298 25 26 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=5.34 $Y=1.375
+ $X2=5.34 $Y2=1.895
r299 22 31 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.18 $Y=2.045
+ $X2=5.18 $Y2=1.97
r300 22 24 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=5.18 $Y=2.045
+ $X2=5.18 $Y2=2.54
r301 19 21 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.175 $Y=2.465
+ $X2=3.175 $Y2=2.75
r302 18 19 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.175 $Y=2.375
+ $X2=3.175 $Y2=2.465
r303 17 89 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.175 $Y=2.075
+ $X2=3.175 $Y2=1.91
r304 17 18 116.613 $w=1.8e-07 $l=3e-07 $layer=POLY_cond $X=3.175 $Y=2.075
+ $X2=3.175 $Y2=2.375
r305 13 87 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.015 $Y=1.745
+ $X2=3.015 $Y2=1.91
r306 13 15 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=3.015 $Y=1.745
+ $X2=3.015 $Y2=0.805
r307 10 81 38.5462 $w=3.19e-07 $l=2.20624e-07 $layer=POLY_cond $X=1.135 $Y=1.22
+ $X2=1.005 $Y2=1.385
r308 10 12 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.135 $Y=1.22
+ $X2=1.135 $Y2=0.74
r309 7 81 71.0321 $w=3.19e-07 $l=4.06571e-07 $layer=POLY_cond $X=0.95 $Y=1.765
+ $X2=1.005 $Y2=1.385
r310 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.95 $Y=1.765
+ $X2=0.95 $Y2=2.4
r311 2 43 400 $w=1.7e-07 $l=1.04265e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.275 $Y2=2.815
r312 2 41 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.275 $Y2=1.985
r313 1 47 182 $w=1.7e-07 $l=3.75566e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_LS__DFXBP_1%D 1 3 4 6 8 10 15 17 18 23 35
c59 35 0 8.5492e-20 $X=2.16 $Y=1.665
c60 17 0 4.57052e-20 $X=2.16 $Y=1.295
c61 15 0 4.61005e-19 $X=1.995 $Y=2.19
c62 4 0 1.35673e-19 $X=2.51 $Y=1.2
c63 1 0 3.08123e-19 $X=2.025 $Y=2.44
r64 29 35 2.0808 $w=3.58e-07 $l=6.5e-08 $layer=LI1_cond $X=2.09 $Y=1.6 $X2=2.09
+ $Y2=1.665
r65 23 26 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.175 $Y=1.2 $X2=2.175
+ $Y2=1.29
r66 18 37 6.59029 $w=3.58e-07 $l=1.05e-07 $layer=LI1_cond $X=2.09 $Y=1.675
+ $X2=2.09 $Y2=1.78
r67 18 35 0.320123 $w=3.58e-07 $l=1e-08 $layer=LI1_cond $X=2.09 $Y=1.675
+ $X2=2.09 $Y2=1.665
r68 18 29 0.320123 $w=3.58e-07 $l=1e-08 $layer=LI1_cond $X=2.09 $Y=1.59 $X2=2.09
+ $Y2=1.6
r69 17 18 9.60369 $w=3.58e-07 $l=3e-07 $layer=LI1_cond $X=2.09 $Y=1.29 $X2=2.09
+ $Y2=1.59
r70 17 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.175
+ $Y=1.29 $X2=2.175 $Y2=1.29
r71 12 15 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=1.865 $Y=2.19
+ $X2=1.995 $Y2=2.19
r72 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.865
+ $Y=2.19 $X2=1.865 $Y2=2.19
r73 10 15 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.995 $Y=2.025
+ $X2=1.995 $Y2=2.19
r74 10 37 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.995 $Y=2.025
+ $X2=1.995 $Y2=1.78
r75 6 8 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.585 $Y=1.125
+ $X2=2.585 $Y2=0.805
r76 5 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.34 $Y=1.2
+ $X2=2.175 $Y2=1.2
r77 4 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.51 $Y=1.2
+ $X2=2.585 $Y2=1.125
r78 4 5 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=2.51 $Y=1.2 $X2=2.34
+ $Y2=1.2
r79 1 13 50.1894 $w=3.66e-07 $l=3.03315e-07 $layer=POLY_cond $X=2.025 $Y=2.44
+ $X2=1.907 $Y2=2.19
r80 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.025 $Y=2.44 $X2=2.025
+ $Y2=2.725
.ends

.subckt PM_SKY130_FD_SC_LS__DFXBP_1%A_205_368# 1 2 9 10 11 14 15 17 20 24 27 28
+ 30 32 35 37 39 41 43 46 47 50 53 56 57 60 64 68 74 76 78 80 81 85
c235 80 0 1.10354e-19 $X=5.825 $Y=1.78
c236 74 0 1.49219e-19 $X=4.89 $Y=1.52
c237 57 0 1.73501e-19 $X=1.222 $Y=2.63
c238 56 0 4.89519e-20 $X=1.635 $Y=1.65
c239 53 0 1.3952e-19 $X=1.43 $Y=1.756
c240 39 0 1.89237e-19 $X=3.12 $Y=2.8
c241 20 0 4.21193e-20 $X=3.49 $Y=0.72
c242 15 0 1.53541e-19 $X=2.64 $Y=2.16
c243 14 0 1.10948e-19 $X=2.64 $Y=2.07
c244 11 0 1.08514e-19 $X=2.55 $Y=1.74
r245 81 91 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=5.825 $Y=1.78
+ $X2=5.715 $Y2=1.78
r246 80 83 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=5.825 $Y=1.78
+ $X2=5.825 $Y2=1.945
r247 80 81 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.825
+ $Y=1.78 $X2=5.825 $Y2=1.78
r248 74 89 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.89 $Y=1.52
+ $X2=4.89 $Y2=1.355
r249 73 76 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=4.89 $Y=1.52
+ $X2=5.065 $Y2=1.52
r250 73 74 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.89
+ $Y=1.52 $X2=4.89 $Y2=1.52
r251 64 66 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=3.205 $Y=2.67
+ $X2=3.205 $Y2=2.8
r252 60 62 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.14 $Y=2.63
+ $X2=2.14 $Y2=2.8
r253 57 59 6.14986 $w=3.67e-07 $l=1.85e-07 $layer=LI1_cond $X=1.222 $Y=2.63
+ $X2=1.222 $Y2=2.815
r254 56 86 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.635 $Y=1.65
+ $X2=1.635 $Y2=1.74
r255 56 85 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.635 $Y=1.65
+ $X2=1.635 $Y2=1.485
r256 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.635
+ $Y=1.65 $X2=1.635 $Y2=1.65
r257 53 55 7.39941 $w=3.38e-07 $l=2.05e-07 $layer=LI1_cond $X=1.43 $Y=1.756
+ $X2=1.635 $Y2=1.756
r258 52 53 9.20414 $w=3.38e-07 $l=3.51312e-07 $layer=LI1_cond $X=1.175 $Y=1.985
+ $X2=1.43 $Y2=1.756
r259 50 83 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=5.905 $Y=2.905
+ $X2=5.905 $Y2=1.945
r260 48 78 4.10697 $w=2.22e-07 $l=1.08305e-07 $layer=LI1_cond $X=5.15 $Y=2.99
+ $X2=5.065 $Y2=2.937
r261 47 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.82 $Y=2.99
+ $X2=5.905 $Y2=2.905
r262 47 48 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.82 $Y=2.99
+ $X2=5.15 $Y2=2.99
r263 46 78 2.32734 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=5.065 $Y=2.8
+ $X2=5.065 $Y2=2.937
r264 45 76 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.065 $Y=1.685
+ $X2=5.065 $Y2=1.52
r265 45 46 72.7433 $w=1.68e-07 $l=1.115e-06 $layer=LI1_cond $X=5.065 $Y=1.685
+ $X2=5.065 $Y2=2.8
r266 44 68 17.4193 $w=1.68e-07 $l=2.67e-07 $layer=LI1_cond $X=4.385 $Y=2.937
+ $X2=4.385 $Y2=2.67
r267 43 78 4.10697 $w=2.22e-07 $l=8.5e-08 $layer=LI1_cond $X=4.98 $Y=2.937
+ $X2=5.065 $Y2=2.937
r268 43 44 21.3726 $w=2.73e-07 $l=5.1e-07 $layer=LI1_cond $X=4.98 $Y=2.937
+ $X2=4.47 $Y2=2.937
r269 42 64 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.29 $Y=2.67
+ $X2=3.205 $Y2=2.67
r270 41 68 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.3 $Y=2.67
+ $X2=4.385 $Y2=2.67
r271 41 42 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=4.3 $Y=2.67
+ $X2=3.29 $Y2=2.67
r272 40 62 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.225 $Y=2.8
+ $X2=2.14 $Y2=2.8
r273 39 66 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.12 $Y=2.8
+ $X2=3.205 $Y2=2.8
r274 39 40 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=3.12 $Y=2.8
+ $X2=2.225 $Y2=2.8
r275 38 57 5.25812 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=1.435 $Y=2.63
+ $X2=1.222 $Y2=2.63
r276 37 60 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.055 $Y=2.63
+ $X2=2.14 $Y2=2.63
r277 37 38 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=2.055 $Y=2.63
+ $X2=1.435 $Y2=2.63
r278 33 53 0.862142 $w=3.3e-07 $l=2.71e-07 $layer=LI1_cond $X=1.43 $Y=1.485
+ $X2=1.43 $Y2=1.756
r279 33 35 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=1.43 $Y=1.485
+ $X2=1.43 $Y2=1.155
r280 32 57 2.70071 $w=4.25e-07 $l=8.5e-08 $layer=LI1_cond $X=1.222 $Y=2.545
+ $X2=1.222 $Y2=2.63
r281 32 52 14.0462 $w=4.23e-07 $l=5.18e-07 $layer=LI1_cond $X=1.222 $Y=2.545
+ $X2=1.222 $Y2=2.027
r282 28 30 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=5.715 $Y=2.335
+ $X2=5.715 $Y2=2.62
r283 27 28 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.715 $Y=2.245
+ $X2=5.715 $Y2=2.335
r284 26 91 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.715 $Y=1.945
+ $X2=5.715 $Y2=1.78
r285 26 27 116.613 $w=1.8e-07 $l=3e-07 $layer=POLY_cond $X=5.715 $Y=1.945
+ $X2=5.715 $Y2=2.245
r286 24 89 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.95 $Y=0.875
+ $X2=4.95 $Y2=1.355
r287 18 20 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.49 $Y=0.255
+ $X2=3.49 $Y2=0.72
r288 15 17 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.64 $Y=2.16
+ $X2=2.64 $Y2=2.445
r289 14 15 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.64 $Y=2.07 $X2=2.64
+ $Y2=2.16
r290 13 14 99.121 $w=1.8e-07 $l=2.55e-07 $layer=POLY_cond $X=2.64 $Y=1.815
+ $X2=2.64 $Y2=2.07
r291 12 86 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.8 $Y=1.74
+ $X2=1.635 $Y2=1.74
r292 11 13 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=2.55 $Y=1.74
+ $X2=2.64 $Y2=1.815
r293 11 12 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=2.55 $Y=1.74
+ $X2=1.8 $Y2=1.74
r294 9 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.415 $Y=0.18
+ $X2=3.49 $Y2=0.255
r295 9 10 828.117 $w=1.5e-07 $l=1.615e-06 $layer=POLY_cond $X=3.415 $Y=0.18
+ $X2=1.8 $Y2=0.18
r296 7 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.725 $Y=0.255
+ $X2=1.8 $Y2=0.18
r297 7 85 630.702 $w=1.5e-07 $l=1.23e-06 $layer=POLY_cond $X=1.725 $Y=0.255
+ $X2=1.725 $Y2=1.485
r298 2 59 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.025
+ $Y=1.84 $X2=1.175 $Y2=2.815
r299 2 52 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.025
+ $Y=1.84 $X2=1.175 $Y2=1.985
r300 1 35 182 $w=1.7e-07 $l=8.88214e-07 $layer=licon1_NDIFF $count=1 $X=1.21
+ $Y=0.37 $X2=1.43 $Y2=1.155
.ends

.subckt PM_SKY130_FD_SC_LS__DFXBP_1%A_701_463# 1 2 7 9 11 12 14 17 19 25 28 32
+ 34 37 40
c89 34 0 1.27123e-19 $X=4.45 $Y=1.015
c90 32 0 5.93116e-20 $X=4.725 $Y=2.42
c91 28 0 1.76992e-19 $X=4.735 $Y=1.005
c92 19 0 4.21193e-20 $X=4.45 $Y=1.192
r93 35 37 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=4.535 $Y=1.94
+ $X2=4.725 $Y2=1.94
r94 30 37 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.725 $Y=2.025
+ $X2=4.725 $Y2=1.94
r95 30 32 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=4.725 $Y=2.025
+ $X2=4.725 $Y2=2.42
r96 26 34 3.05675 $w=3.1e-07 $l=1.8759e-07 $layer=LI1_cond $X=4.62 $Y=1.052
+ $X2=4.45 $Y2=1.015
r97 26 28 5.00117 $w=2.63e-07 $l=1.15e-07 $layer=LI1_cond $X=4.62 $Y=1.052
+ $X2=4.735 $Y2=1.052
r98 25 35 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.535 $Y=1.855
+ $X2=4.535 $Y2=1.94
r99 24 34 3.57226 $w=1.7e-07 $l=3.95221e-07 $layer=LI1_cond $X=4.535 $Y=1.37
+ $X2=4.45 $Y2=1.015
r100 24 25 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=4.535 $Y=1.37
+ $X2=4.535 $Y2=1.855
r101 22 40 20.6994 $w=3.26e-07 $l=1.4e-07 $layer=POLY_cond $X=3.99 $Y=1.23
+ $X2=3.85 $Y2=1.23
r102 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.99
+ $Y=1.205 $X2=3.99 $Y2=1.205
r103 19 34 3.05675 $w=3.1e-07 $l=1.77e-07 $layer=LI1_cond $X=4.45 $Y=1.192
+ $X2=4.45 $Y2=1.015
r104 19 21 14.9331 $w=3.53e-07 $l=4.6e-07 $layer=LI1_cond $X=4.45 $Y=1.192
+ $X2=3.99 $Y2=1.192
r105 15 17 71.7872 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=3.595 $Y=2.39
+ $X2=3.735 $Y2=2.39
r106 12 40 20.933 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=3.85 $Y=1.04
+ $X2=3.85 $Y2=1.23
r107 12 14 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.85 $Y=1.04
+ $X2=3.85 $Y2=0.72
r108 11 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.735 $Y=2.315
+ $X2=3.735 $Y2=2.39
r109 10 40 17.0031 $w=3.26e-07 $l=2.40728e-07 $layer=POLY_cond $X=3.735 $Y=1.42
+ $X2=3.85 $Y2=1.23
r110 10 11 458.926 $w=1.5e-07 $l=8.95e-07 $layer=POLY_cond $X=3.735 $Y=1.42
+ $X2=3.735 $Y2=2.315
r111 7 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.595 $Y=2.465
+ $X2=3.595 $Y2=2.39
r112 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.595 $Y=2.465
+ $X2=3.595 $Y2=2.75
r113 2 32 600 $w=1.7e-07 $l=3.96863e-07 $layer=licon1_PDIFF $count=1 $X=4.5
+ $Y=2.12 $X2=4.725 $Y2=2.42
r114 1 28 182 $w=1.7e-07 $l=7.26722e-07 $layer=licon1_NDIFF $count=1 $X=4.515
+ $Y=0.38 $X2=4.735 $Y2=1.005
.ends

.subckt PM_SKY130_FD_SC_LS__DFXBP_1%A_543_447# 1 2 7 9 12 15 16 18 20 24
c88 20 0 1.35673e-19 $X=3.23 $Y=0.77
r89 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.185
+ $Y=1.795 $X2=4.185 $Y2=1.795
r90 22 24 19.9461 $w=2.58e-07 $l=4.5e-07 $layer=LI1_cond $X=4.15 $Y=2.245
+ $X2=4.15 $Y2=1.795
r91 18 27 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=3.19 $Y=1.495
+ $X2=2.865 $Y2=1.495
r92 18 20 29.5025 $w=2.48e-07 $l=6.4e-07 $layer=LI1_cond $X=3.19 $Y=1.41
+ $X2=3.19 $Y2=0.77
r93 17 32 3.40825 $w=1.7e-07 $l=1.12916e-07 $layer=LI1_cond $X=2.95 $Y=2.33
+ $X2=2.865 $Y2=2.395
r94 16 22 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=4.02 $Y=2.33
+ $X2=4.15 $Y2=2.245
r95 16 17 69.8075 $w=1.68e-07 $l=1.07e-06 $layer=LI1_cond $X=4.02 $Y=2.33
+ $X2=2.95 $Y2=2.33
r96 15 32 3.40825 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=2.865 $Y=2.245
+ $X2=2.865 $Y2=2.395
r97 14 27 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.865 $Y=1.58
+ $X2=2.865 $Y2=1.495
r98 14 15 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=2.865 $Y=1.58
+ $X2=2.865 $Y2=2.245
r99 10 25 40.2182 $w=4.3e-07 $l=2.41814e-07 $layer=POLY_cond $X=4.44 $Y=1.63
+ $X2=4.267 $Y2=1.795
r100 10 12 499.947 $w=1.5e-07 $l=9.75e-07 $layer=POLY_cond $X=4.44 $Y=1.63
+ $X2=4.44 $Y2=0.655
r101 7 25 49.7461 $w=4.3e-07 $l=3.19374e-07 $layer=POLY_cond $X=4.425 $Y=2.045
+ $X2=4.267 $Y2=1.795
r102 7 9 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=4.425 $Y=2.045
+ $X2=4.425 $Y2=2.54
r103 2 32 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.715
+ $Y=2.235 $X2=2.865 $Y2=2.38
r104 1 20 182 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=1 $X=3.09
+ $Y=0.595 $X2=3.23 $Y2=0.77
.ends

.subckt PM_SKY130_FD_SC_LS__DFXBP_1%A_1191_120# 1 2 7 9 10 12 17 19 21 22 23 26
+ 28 30 33 38 41 42 45 49 51 52 53 54 59 63 65
c146 33 0 4.23824e-20 $X=6.305 $Y=1.3
c147 23 0 3.58297e-19 $X=7.695 $Y=1.515
c148 7 0 1.54211e-19 $X=6.03 $Y=1.225
r149 70 71 1.89764 $w=3.81e-07 $l=1.5e-08 $layer=POLY_cond $X=7.59 $Y=1.557
+ $X2=7.605 $Y2=1.557
r150 64 70 3.16273 $w=3.81e-07 $l=2.5e-08 $layer=POLY_cond $X=7.565 $Y=1.557
+ $X2=7.59 $Y2=1.557
r151 63 66 6.96826 $w=4.28e-07 $l=2.6e-07 $layer=LI1_cond $X=7.515 $Y=1.515
+ $X2=7.515 $Y2=1.775
r152 63 65 8.78489 $w=4.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.515 $Y=1.515
+ $X2=7.515 $Y2=1.35
r153 63 64 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.565
+ $Y=1.515 $X2=7.565 $Y2=1.515
r154 58 61 9.97615 $w=5.87e-07 $l=4.8e-07 $layer=LI1_cond $X=6.395 $Y=1.885
+ $X2=6.875 $Y2=1.885
r155 58 59 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.395
+ $Y=1.715 $X2=6.395 $Y2=1.715
r156 55 65 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=7.385 $Y=1.02
+ $X2=7.385 $Y2=1.35
r157 54 61 10.2728 $w=5.87e-07 $l=2.13014e-07 $layer=LI1_cond $X=7.04 $Y=1.775
+ $X2=6.875 $Y2=1.885
r158 53 66 6.22023 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=7.3 $Y=1.775
+ $X2=7.515 $Y2=1.775
r159 53 54 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=7.3 $Y=1.775
+ $X2=7.04 $Y2=1.775
r160 51 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.3 $Y=0.935
+ $X2=7.385 $Y2=1.02
r161 51 52 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=7.3 $Y=0.935
+ $X2=6.97 $Y2=0.935
r162 47 61 4.10774 $w=3.3e-07 $l=3.35e-07 $layer=LI1_cond $X=6.875 $Y=2.22
+ $X2=6.875 $Y2=1.885
r163 47 49 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=6.875 $Y=2.22
+ $X2=6.875 $Y2=2.695
r164 43 52 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.805 $Y=0.85
+ $X2=6.97 $Y2=0.935
r165 43 45 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=6.805 $Y=0.85
+ $X2=6.805 $Y2=0.645
r166 41 59 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.395 $Y=1.55
+ $X2=6.395 $Y2=1.715
r167 38 59 82.1848 $w=3.3e-07 $l=4.7e-07 $layer=POLY_cond $X=6.395 $Y=2.185
+ $X2=6.395 $Y2=1.715
r168 35 38 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=6.105 $Y=2.26
+ $X2=6.395 $Y2=2.26
r169 31 33 141.011 $w=1.5e-07 $l=2.75e-07 $layer=POLY_cond $X=6.03 $Y=1.3
+ $X2=6.305 $Y2=1.3
r170 28 42 37.0704 $w=1.5e-07 $l=4.57794e-07 $layer=POLY_cond $X=8.595 $Y=1.765
+ $X2=8.505 $Y2=1.35
r171 28 30 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=8.595 $Y=1.765
+ $X2=8.595 $Y2=2.26
r172 24 42 37.0704 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.58 $Y=1.35
+ $X2=8.505 $Y2=1.35
r173 24 26 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=8.58 $Y=1.35
+ $X2=8.58 $Y2=0.835
r174 23 71 12.3804 $w=3.81e-07 $l=1.08995e-07 $layer=POLY_cond $X=7.695 $Y=1.515
+ $X2=7.605 $Y2=1.557
r175 22 42 5.03009 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.505 $Y=1.515
+ $X2=8.505 $Y2=1.35
r176 22 23 141.638 $w=3.3e-07 $l=8.1e-07 $layer=POLY_cond $X=8.505 $Y=1.515
+ $X2=7.695 $Y2=1.515
r177 19 71 24.6764 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=7.605 $Y=1.765
+ $X2=7.605 $Y2=1.557
r178 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.605 $Y=1.765
+ $X2=7.605 $Y2=2.4
r179 15 70 24.6764 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.59 $Y=1.35
+ $X2=7.59 $Y2=1.557
r180 15 17 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.59 $Y=1.35
+ $X2=7.59 $Y2=0.74
r181 13 33 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.305 $Y=1.375
+ $X2=6.305 $Y2=1.3
r182 13 41 89.734 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=6.305 $Y=1.375
+ $X2=6.305 $Y2=1.55
r183 10 35 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.105 $Y=2.335
+ $X2=6.105 $Y2=2.26
r184 10 12 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.105 $Y=2.335
+ $X2=6.105 $Y2=2.62
r185 7 31 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.03 $Y=1.225
+ $X2=6.03 $Y2=1.3
r186 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.03 $Y=1.225 $X2=6.03
+ $Y2=0.94
r187 2 61 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=6.735
+ $Y=1.84 $X2=6.875 $Y2=1.985
r188 2 49 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=6.735
+ $Y=1.84 $X2=6.875 $Y2=2.695
r189 1 45 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=6.66
+ $Y=0.37 $X2=6.805 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_LS__DFXBP_1%A_1005_120# 1 2 9 11 13 14 16 18 25 27 29
c81 27 0 2.55347e-19 $X=6.965 $Y=1.355
c82 14 0 5.7879e-20 $X=5.405 $Y=1.38
c83 9 0 2.43826e-20 $X=7.02 $Y=0.645
r84 27 29 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=6.965 $Y=1.355
+ $X2=6.8 $Y2=1.355
r85 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.965
+ $Y=1.355 $X2=6.965 $Y2=1.355
r86 23 24 10.9446 $w=3.79e-07 $l=3.4e-07 $layer=LI1_cond $X=5.357 $Y=0.955
+ $X2=5.357 $Y2=1.295
r87 21 24 5.45184 $w=1.7e-07 $l=2.33e-07 $layer=LI1_cond $X=5.59 $Y=1.295
+ $X2=5.357 $Y2=1.295
r88 21 29 78.9412 $w=1.68e-07 $l=1.21e-06 $layer=LI1_cond $X=5.59 $Y=1.295
+ $X2=6.8 $Y2=1.295
r89 16 25 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=5.445 $Y=2.24
+ $X2=5.445 $Y2=2.115
r90 16 18 14.0598 $w=2.48e-07 $l=3.05e-07 $layer=LI1_cond $X=5.445 $Y=2.24
+ $X2=5.445 $Y2=2.545
r91 14 24 6.49482 $w=3.79e-07 $l=1.06325e-07 $layer=LI1_cond $X=5.405 $Y=1.38
+ $X2=5.357 $Y2=1.295
r92 14 25 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=5.405 $Y=1.38
+ $X2=5.405 $Y2=2.115
r93 11 28 80.4178 $w=2.83e-07 $l=4.59511e-07 $layer=POLY_cond $X=7.1 $Y=1.765
+ $X2=6.995 $Y2=1.355
r94 11 13 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=7.1 $Y=1.765
+ $X2=7.1 $Y2=2.34
r95 7 28 38.6899 $w=2.83e-07 $l=1.77059e-07 $layer=POLY_cond $X=7.02 $Y=1.19
+ $X2=6.995 $Y2=1.355
r96 7 9 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=7.02 $Y=1.19 $X2=7.02
+ $Y2=0.645
r97 2 18 600 $w=1.7e-07 $l=4.94343e-07 $layer=licon1_PDIFF $count=1 $X=5.255
+ $Y=2.12 $X2=5.405 $Y2=2.545
r98 1 23 182 $w=1.7e-07 $l=4.69148e-07 $layer=licon1_NDIFF $count=1 $X=5.025
+ $Y=0.6 $X2=5.29 $Y2=0.955
.ends

.subckt PM_SKY130_FD_SC_LS__DFXBP_1%A_1644_112# 1 2 9 11 13 16 20 24 27
r50 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.06
+ $Y=1.465 $X2=9.06 $Y2=1.465
r51 22 27 0.182887 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=8.53 $Y=1.465
+ $X2=8.405 $Y2=1.465
r52 22 24 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=8.53 $Y=1.465
+ $X2=9.06 $Y2=1.465
r53 18 27 7.32358 $w=2.12e-07 $l=1.83016e-07 $layer=LI1_cond $X=8.367 $Y=1.63
+ $X2=8.405 $Y2=1.465
r54 18 20 22.4987 $w=1.73e-07 $l=3.55e-07 $layer=LI1_cond $X=8.367 $Y=1.63
+ $X2=8.367 $Y2=1.985
r55 14 27 7.32358 $w=2.12e-07 $l=1.65e-07 $layer=LI1_cond $X=8.405 $Y=1.3
+ $X2=8.405 $Y2=1.465
r56 14 16 21.4354 $w=2.48e-07 $l=4.65e-07 $layer=LI1_cond $X=8.405 $Y=1.3
+ $X2=8.405 $Y2=0.835
r57 11 25 61.4066 $w=2.86e-07 $l=3.19374e-07 $layer=POLY_cond $X=9.1 $Y=1.765
+ $X2=9.06 $Y2=1.465
r58 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=9.1 $Y=1.765
+ $X2=9.1 $Y2=2.4
r59 7 25 38.6549 $w=2.86e-07 $l=1.79374e-07 $layer=POLY_cond $X=9.09 $Y=1.3
+ $X2=9.06 $Y2=1.465
r60 7 9 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=9.09 $Y=1.3 $X2=9.09
+ $Y2=0.74
r61 2 20 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=8.235
+ $Y=1.84 $X2=8.37 $Y2=1.985
r62 1 16 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=8.22
+ $Y=0.56 $X2=8.365 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_LS__DFXBP_1%VPWR 1 2 3 4 5 6 21 25 29 33 37 40 41 42 44
+ 49 54 66 70 77 78 81 84 87 94 97
r122 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r123 94 95 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r124 90 91 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r125 87 90 9.45594 $w=3.88e-07 $l=3.2e-07 $layer=LI1_cond $X=3.935 $Y=3.01
+ $X2=3.935 $Y2=3.33
r126 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r127 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r128 78 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=8.88 $Y2=3.33
r129 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r130 75 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.985 $Y=3.33
+ $X2=8.82 $Y2=3.33
r131 75 77 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=8.985 $Y=3.33
+ $X2=9.36 $Y2=3.33
r132 74 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=8.88 $Y2=3.33
r133 74 95 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=7.44 $Y2=3.33
r134 73 74 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r135 71 94 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.49 $Y=3.33
+ $X2=7.365 $Y2=3.33
r136 71 73 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=7.49 $Y=3.33 $X2=8.4
+ $Y2=3.33
r137 70 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.655 $Y=3.33
+ $X2=8.82 $Y2=3.33
r138 70 73 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=8.655 $Y=3.33
+ $X2=8.4 $Y2=3.33
r139 69 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.44 $Y2=3.33
r140 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r141 66 94 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.24 $Y=3.33
+ $X2=7.365 $Y2=3.33
r142 66 68 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=7.24 $Y=3.33
+ $X2=6.96 $Y2=3.33
r143 65 69 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.96
+ $Y2=3.33
r144 64 65 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r145 62 90 5.6248 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=4.13 $Y=3.33
+ $X2=3.935 $Y2=3.33
r146 62 64 122 $w=1.68e-07 $l=1.87e-06 $layer=LI1_cond $X=4.13 $Y=3.33 $X2=6
+ $Y2=3.33
r147 61 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r148 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r149 58 61 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.6 $Y2=3.33
r150 58 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r151 57 60 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=3.6 $Y2=3.33
r152 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r153 55 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.885 $Y=3.33
+ $X2=1.72 $Y2=3.33
r154 55 57 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.885 $Y=3.33
+ $X2=2.16 $Y2=3.33
r155 54 90 5.6248 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=3.74 $Y=3.33
+ $X2=3.935 $Y2=3.33
r156 54 60 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=3.74 $Y=3.33
+ $X2=3.6 $Y2=3.33
r157 53 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r158 53 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r159 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r160 50 81 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.81 $Y=3.33
+ $X2=0.685 $Y2=3.33
r161 50 52 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=0.81 $Y=3.33
+ $X2=1.2 $Y2=3.33
r162 49 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.555 $Y=3.33
+ $X2=1.72 $Y2=3.33
r163 49 52 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=1.555 $Y=3.33
+ $X2=1.2 $Y2=3.33
r164 47 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r165 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r166 44 81 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.56 $Y=3.33
+ $X2=0.685 $Y2=3.33
r167 44 46 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.56 $Y=3.33
+ $X2=0.24 $Y2=3.33
r168 42 65 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=4.8 $Y=3.33 $X2=6
+ $Y2=3.33
r169 42 91 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=4.8 $Y=3.33
+ $X2=4.08 $Y2=3.33
r170 40 64 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=6.165 $Y=3.33
+ $X2=6 $Y2=3.33
r171 40 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.165 $Y=3.33
+ $X2=6.33 $Y2=3.33
r172 39 68 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=6.495 $Y=3.33
+ $X2=6.96 $Y2=3.33
r173 39 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.495 $Y=3.33
+ $X2=6.33 $Y2=3.33
r174 35 97 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.82 $Y=3.245
+ $X2=8.82 $Y2=3.33
r175 35 37 44.0024 $w=3.28e-07 $l=1.26e-06 $layer=LI1_cond $X=8.82 $Y=3.245
+ $X2=8.82 $Y2=1.985
r176 31 94 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.365 $Y=3.245
+ $X2=7.365 $Y2=3.33
r177 31 33 48.4026 $w=2.48e-07 $l=1.05e-06 $layer=LI1_cond $X=7.365 $Y=3.245
+ $X2=7.365 $Y2=2.195
r178 27 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.33 $Y=3.245
+ $X2=6.33 $Y2=3.33
r179 27 29 21.8266 $w=3.28e-07 $l=6.25e-07 $layer=LI1_cond $X=6.33 $Y=3.245
+ $X2=6.33 $Y2=2.62
r180 23 84 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.72 $Y=3.245
+ $X2=1.72 $Y2=3.33
r181 23 25 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=1.72 $Y=3.245
+ $X2=1.72 $Y2=3.05
r182 19 81 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.685 $Y=3.245
+ $X2=0.685 $Y2=3.33
r183 19 21 47.0197 $w=2.48e-07 $l=1.02e-06 $layer=LI1_cond $X=0.685 $Y=3.245
+ $X2=0.685 $Y2=2.225
r184 6 37 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=8.67
+ $Y=1.84 $X2=8.82 $Y2=1.985
r185 5 33 300 $w=1.7e-07 $l=4.23409e-07 $layer=licon1_PDIFF $count=2 $X=7.175
+ $Y=1.84 $X2=7.325 $Y2=2.195
r186 4 29 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=6.18
+ $Y=2.41 $X2=6.33 $Y2=2.62
r187 3 87 600 $w=1.7e-07 $l=5.8775e-07 $layer=licon1_PDIFF $count=1 $X=3.67
+ $Y=2.54 $X2=3.935 $Y2=3.01
r188 2 25 600 $w=1.7e-07 $l=6.00937e-07 $layer=licon1_PDIFF $count=1 $X=1.58
+ $Y=2.515 $X2=1.72 $Y2=3.05
r189 1 21 300 $w=1.7e-07 $l=4.53845e-07 $layer=licon1_PDIFF $count=2 $X=0.575
+ $Y=1.84 $X2=0.725 $Y2=2.225
.ends

.subckt PM_SKY130_FD_SC_LS__DFXBP_1%A_420_503# 1 2 8 11 16 20
c40 16 0 1.56514e-19 $X=2.525 $Y=2.21
c41 8 0 1.68603e-19 $X=2.525 $Y=2.045
r42 18 20 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.525 $Y=1.155
+ $X2=2.8 $Y2=1.155
r43 14 16 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=2.335 $Y=2.21
+ $X2=2.525 $Y2=2.21
r44 9 20 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.8 $Y=1.07 $X2=2.8
+ $Y2=1.155
r45 9 11 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.8 $Y=1.07 $X2=2.8
+ $Y2=0.815
r46 8 16 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.525 $Y=2.045
+ $X2=2.525 $Y2=2.21
r47 7 18 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.525 $Y=1.24
+ $X2=2.525 $Y2=1.155
r48 7 8 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=2.525 $Y=1.24
+ $X2=2.525 $Y2=2.045
r49 2 14 600 $w=1.7e-07 $l=4.05832e-07 $layer=licon1_PDIFF $count=1 $X=2.1
+ $Y=2.515 $X2=2.335 $Y2=2.21
r50 1 11 182 $w=1.7e-07 $l=2.81425e-07 $layer=licon1_NDIFF $count=1 $X=2.66
+ $Y=0.595 $X2=2.8 $Y2=0.815
.ends

.subckt PM_SKY130_FD_SC_LS__DFXBP_1%Q 1 2 9 13 16 17 18 19
c36 13 0 2.43826e-20 $X=7.855 $Y=1.13
r37 18 19 10.5285 $w=4.03e-07 $l=3.7e-07 $layer=LI1_cond $X=7.867 $Y=2.405
+ $X2=7.867 $Y2=2.775
r38 16 17 8.6688 $w=4.03e-07 $l=1.65e-07 $layer=LI1_cond $X=7.867 $Y=2.195
+ $X2=7.867 $Y2=2.03
r39 14 18 4.92278 $w=4.03e-07 $l=1.73e-07 $layer=LI1_cond $X=7.867 $Y=2.232
+ $X2=7.867 $Y2=2.405
r40 14 16 1.05285 $w=4.03e-07 $l=3.7e-08 $layer=LI1_cond $X=7.867 $Y=2.232
+ $X2=7.867 $Y2=2.195
r41 13 17 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=7.985 $Y=1.13
+ $X2=7.985 $Y2=2.03
r42 7 13 10.1249 $w=4.28e-07 $l=2.15e-07 $layer=LI1_cond $X=7.855 $Y=0.915
+ $X2=7.855 $Y2=1.13
r43 7 9 10.7204 $w=4.28e-07 $l=4e-07 $layer=LI1_cond $X=7.855 $Y=0.915 $X2=7.855
+ $Y2=0.515
r44 2 16 300 $w=1.7e-07 $l=4.23409e-07 $layer=licon1_PDIFF $count=2 $X=7.68
+ $Y=1.84 $X2=7.83 $Y2=2.195
r45 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.665
+ $Y=0.37 $X2=7.805 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__DFXBP_1%Q_N 1 2 9 13 14 15 16 23 32
r23 21 23 1.2336 $w=3.53e-07 $l=3.8e-08 $layer=LI1_cond $X=9.337 $Y=1.997
+ $X2=9.337 $Y2=2.035
r24 15 16 12.0114 $w=3.53e-07 $l=3.7e-07 $layer=LI1_cond $X=9.337 $Y=2.405
+ $X2=9.337 $Y2=2.775
r25 14 21 0.779116 $w=3.53e-07 $l=2.4e-08 $layer=LI1_cond $X=9.337 $Y=1.973
+ $X2=9.337 $Y2=1.997
r26 14 32 8.1095 $w=3.53e-07 $l=1.53e-07 $layer=LI1_cond $X=9.337 $Y=1.973
+ $X2=9.337 $Y2=1.82
r27 14 15 11.2647 $w=3.53e-07 $l=3.47e-07 $layer=LI1_cond $X=9.337 $Y=2.058
+ $X2=9.337 $Y2=2.405
r28 14 23 0.746653 $w=3.53e-07 $l=2.3e-08 $layer=LI1_cond $X=9.337 $Y=2.058
+ $X2=9.337 $Y2=2.035
r29 13 32 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=9.43 $Y=1.13 $X2=9.43
+ $Y2=1.82
r30 7 13 9.23056 $w=3.73e-07 $l=1.87e-07 $layer=LI1_cond $X=9.327 $Y=0.943
+ $X2=9.327 $Y2=1.13
r31 7 9 13.1532 $w=3.73e-07 $l=4.28e-07 $layer=LI1_cond $X=9.327 $Y=0.943
+ $X2=9.327 $Y2=0.515
r32 2 14 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=9.175
+ $Y=1.84 $X2=9.325 $Y2=1.985
r33 2 16 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=9.175
+ $Y=1.84 $X2=9.325 $Y2=2.815
r34 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.165
+ $Y=0.37 $X2=9.305 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__DFXBP_1%VGND 1 2 3 4 5 6 21 25 29 33 37 42 43 45 46
+ 47 49 54 59 71 80 81 84 87 91 97
c120 33 0 1.91441e-19 $X=7.305 $Y=0.515
r121 97 98 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r122 91 94 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=4.145 $Y=0
+ $X2=4.145 $Y2=0.325
r123 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r124 87 88 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r125 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r126 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r127 78 81 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=9.36
+ $Y2=0
r128 78 98 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=7.44
+ $Y2=0
r129 77 78 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r130 75 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.47 $Y=0 $X2=7.305
+ $Y2=0
r131 75 77 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=7.47 $Y=0 $X2=8.4
+ $Y2=0
r132 74 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r133 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r134 71 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.14 $Y=0 $X2=7.305
+ $Y2=0
r135 71 73 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=7.14 $Y=0 $X2=6.96
+ $Y2=0
r136 70 74 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.96
+ $Y2=0
r137 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6 $Y2=0
r138 67 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r139 66 69 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=4.56 $Y=0 $X2=6
+ $Y2=0
r140 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r141 64 91 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.31 $Y=0 $X2=4.145
+ $Y2=0
r142 64 66 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=4.31 $Y=0 $X2=4.56
+ $Y2=0
r143 63 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r144 63 88 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=3.6 $Y=0 $X2=2.16
+ $Y2=0
r145 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r146 60 87 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=2.205 $Y=0 $X2=2.03
+ $Y2=0
r147 60 62 91.0107 $w=1.68e-07 $l=1.395e-06 $layer=LI1_cond $X=2.205 $Y=0
+ $X2=3.6 $Y2=0
r148 59 91 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.98 $Y=0 $X2=4.145
+ $Y2=0
r149 59 62 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=3.98 $Y=0 $X2=3.6
+ $Y2=0
r150 58 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r151 58 85 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r152 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r153 55 84 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.005 $Y=0 $X2=0.815
+ $Y2=0
r154 55 57 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=1.005 $Y=0
+ $X2=1.68 $Y2=0
r155 54 87 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=1.855 $Y=0 $X2=2.03
+ $Y2=0
r156 54 57 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.855 $Y=0
+ $X2=1.68 $Y2=0
r157 52 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r158 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r159 49 84 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.625 $Y=0 $X2=0.815
+ $Y2=0
r160 49 51 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.625 $Y=0
+ $X2=0.24 $Y2=0
r161 47 70 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=4.8 $Y=0 $X2=6
+ $Y2=0
r162 47 67 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.8 $Y=0 $X2=4.56
+ $Y2=0
r163 45 77 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=8.71 $Y=0 $X2=8.4
+ $Y2=0
r164 45 46 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.71 $Y=0 $X2=8.835
+ $Y2=0
r165 44 80 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=8.96 $Y=0 $X2=9.36
+ $Y2=0
r166 44 46 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.96 $Y=0 $X2=8.835
+ $Y2=0
r167 42 69 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=6.08 $Y=0 $X2=6 $Y2=0
r168 42 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.08 $Y=0 $X2=6.245
+ $Y2=0
r169 41 73 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=6.41 $Y=0 $X2=6.96
+ $Y2=0
r170 41 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.41 $Y=0 $X2=6.245
+ $Y2=0
r171 37 39 20.744 $w=2.48e-07 $l=4.5e-07 $layer=LI1_cond $X=8.835 $Y=0.515
+ $X2=8.835 $Y2=0.965
r172 35 46 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.835 $Y=0.085
+ $X2=8.835 $Y2=0
r173 35 37 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=8.835 $Y=0.085
+ $X2=8.835 $Y2=0.515
r174 31 97 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.305 $Y=0.085
+ $X2=7.305 $Y2=0
r175 31 33 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=7.305 $Y=0.085
+ $X2=7.305 $Y2=0.515
r176 27 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.245 $Y=0.085
+ $X2=6.245 $Y2=0
r177 27 29 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=6.245 $Y=0.085
+ $X2=6.245 $Y2=0.875
r178 23 87 1.07557 $w=3.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.03 $Y=0.085
+ $X2=2.03 $Y2=0
r179 23 25 12.8415 $w=3.48e-07 $l=3.9e-07 $layer=LI1_cond $X=2.03 $Y=0.085
+ $X2=2.03 $Y2=0.475
r180 19 84 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=0.085
+ $X2=0.815 $Y2=0
r181 19 21 9.40151 $w=3.78e-07 $l=3.1e-07 $layer=LI1_cond $X=0.815 $Y=0.085
+ $X2=0.815 $Y2=0.395
r182 6 39 182 $w=1.7e-07 $l=5.03115e-07 $layer=licon1_NDIFF $count=1 $X=8.655
+ $Y=0.56 $X2=8.875 $Y2=0.965
r183 6 37 182 $w=1.7e-07 $l=2.41454e-07 $layer=licon1_NDIFF $count=1 $X=8.655
+ $Y=0.56 $X2=8.875 $Y2=0.515
r184 5 33 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=7.095
+ $Y=0.37 $X2=7.305 $Y2=0.515
r185 4 29 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=6.105
+ $Y=0.73 $X2=6.245 $Y2=0.875
r186 3 94 182 $w=1.7e-07 $l=2.98496e-07 $layer=licon1_NDIFF $count=1 $X=3.925
+ $Y=0.51 $X2=4.145 $Y2=0.325
r187 2 25 182 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=1 $X=1.875
+ $Y=0.33 $X2=2.03 $Y2=0.475
r188 1 21 182 $w=1.7e-07 $l=2.57196e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.815 $Y2=0.395
.ends

