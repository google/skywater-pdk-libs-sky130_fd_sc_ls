* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
M1000 a_509_392# B2 a_310_392# VPB phighvt w=1e+06u l=150000u
+  ad=6.05e+11p pd=5.21e+06u as=6e+11p ps=5.2e+06u
M1001 a_148_260# C1 VGND VNB nshort w=640000u l=150000u
+  ad=4.192e+11p pd=3.87e+06u as=8.64875e+11p ps=5.71e+06u
M1002 a_417_79# A2 VGND VNB nshort w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1003 a_148_260# A1 a_417_79# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND a_148_260# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=1.961e+11p ps=2.01e+06u
M1005 a_597_79# B1 a_148_260# VNB nshort w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1006 VGND B2 a_597_79# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR a_148_260# X VPB phighvt w=1.12e+06u l=150000u
+  ad=6.73e+11p pd=5.52e+06u as=3.08e+11p ps=2.79e+06u
M1008 a_310_392# A2 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_148_260# C1 a_509_392# VPB phighvt w=1e+06u l=150000u
+  ad=2.75e+11p pd=2.55e+06u as=0p ps=0u
M1010 VPWR A1 a_310_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_310_392# B1 a_509_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
