* File: sky130_fd_sc_ls__dlclkp_4.pex.spice
* Created: Fri Aug 28 13:17:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__DLCLKP_4%A_84_48# 1 2 7 9 10 12 14 15 17 18 20 22 23
+ 25 27 29 31
c86 10 0 6.50014e-20 $X=0.6 $Y=1.765
r87 34 36 8.4794 $w=3.43e-07 $l=1.65e-07 $layer=LI1_cond $X=0.707 $Y=1.385
+ $X2=0.707 $Y2=1.55
r88 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.695
+ $Y=1.385 $X2=0.695 $Y2=1.385
r89 31 34 3.67446 $w=3.43e-07 $l=1.1e-07 $layer=LI1_cond $X=0.707 $Y=1.275
+ $X2=0.707 $Y2=1.385
r90 27 29 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=1.605 $Y=2.685
+ $X2=2.15 $Y2=2.685
r91 23 25 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=1.605 $Y=0.815
+ $X2=2.06 $Y2=0.815
r92 22 27 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.52 $Y=2.52
+ $X2=1.605 $Y2=2.685
r93 21 22 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=1.52 $Y=2.14
+ $X2=1.52 $Y2=2.52
r94 19 23 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.52 $Y=0.98
+ $X2=1.605 $Y2=0.815
r95 19 20 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=1.52 $Y=0.98
+ $X2=1.52 $Y2=1.19
r96 17 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.435 $Y=2.055
+ $X2=1.52 $Y2=2.14
r97 17 18 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=1.435 $Y=2.055
+ $X2=0.88 $Y2=2.055
r98 16 31 4.88813 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.88 $Y=1.275
+ $X2=0.707 $Y2=1.275
r99 15 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.435 $Y=1.275
+ $X2=1.52 $Y2=1.19
r100 15 16 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=1.435 $Y=1.275
+ $X2=0.88 $Y2=1.275
r101 14 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.795 $Y=1.97
+ $X2=0.88 $Y2=2.055
r102 14 36 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=0.795 $Y=1.97
+ $X2=0.795 $Y2=1.55
r103 10 35 69.4037 $w=3.37e-07 $l=3.995e-07 $layer=POLY_cond $X=0.6 $Y=1.765
+ $X2=0.64 $Y2=1.385
r104 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.6 $Y=1.765
+ $X2=0.6 $Y2=2.4
r105 7 35 38.6529 $w=3.37e-07 $l=2.26164e-07 $layer=POLY_cond $X=0.495 $Y=1.22
+ $X2=0.64 $Y2=1.385
r106 7 9 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.495 $Y=1.22
+ $X2=0.495 $Y2=0.74
r107 2 29 600 $w=1.7e-07 $l=8.68332e-07 $layer=licon1_PDIFF $count=1 $X=1.835
+ $Y=1.96 $X2=2.15 $Y2=2.685
r108 1 25 182 $w=1.7e-07 $l=5.21368e-07 $layer=licon1_NDIFF $count=1 $X=1.82
+ $Y=0.4 $X2=2.06 $Y2=0.815
.ends

.subckt PM_SKY130_FD_SC_LS__DLCLKP_4%GATE 1 3 6 8
c32 8 0 6.50014e-20 $X=1.2 $Y=1.665
c33 1 0 1.40564e-19 $X=1.34 $Y=1.885
r34 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.265
+ $Y=1.635 $X2=1.265 $Y2=1.635
r35 4 11 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=1.355 $Y=1.47
+ $X2=1.265 $Y2=1.635
r36 4 6 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=1.355 $Y=1.47
+ $X2=1.355 $Y2=0.72
r37 1 11 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=1.34 $Y=1.885
+ $X2=1.265 $Y2=1.635
r38 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.34 $Y=1.885
+ $X2=1.34 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_LS__DLCLKP_4%A_334_54# 1 2 7 9 10 12 13 15 19 22 23 25
+ 26 30 31 32 33 34 37 41 45
c122 37 0 2.3821e-19 $X=3.98 $Y=0.35
c123 26 0 1.40564e-19 $X=2.065 $Y=2.2
c124 19 0 1.80208e-19 $X=3.695 $Y=0.995
r125 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.49
+ $Y=1.795 $X2=3.49 $Y2=1.795
r126 43 45 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=4.445 $Y=0.515
+ $X2=4.445 $Y2=0.685
r127 39 41 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=4.37 $Y=2.52
+ $X2=4.37 $Y2=2.255
r128 37 57 49.8355 $w=3.3e-07 $l=2.85e-07 $layer=POLY_cond $X=3.98 $Y=0.35
+ $X2=3.695 $Y2=0.35
r129 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.98
+ $Y=0.35 $X2=3.98 $Y2=0.35
r130 34 43 6.94204 $w=2.6e-07 $l=2.20624e-07 $layer=LI1_cond $X=4.28 $Y=0.385
+ $X2=4.445 $Y2=0.515
r131 34 36 13.2974 $w=2.58e-07 $l=3e-07 $layer=LI1_cond $X=4.28 $Y=0.385
+ $X2=3.98 $Y2=0.385
r132 32 39 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.205 $Y=2.605
+ $X2=4.37 $Y2=2.52
r133 32 33 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=4.205 $Y=2.605
+ $X2=3.475 $Y2=2.605
r134 31 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.39 $Y=2.52
+ $X2=3.475 $Y2=2.605
r135 30 31 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.39 $Y=2.35
+ $X2=3.39 $Y2=2.52
r136 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.47
+ $Y=2.215 $X2=2.47 $Y2=2.215
r137 26 28 15.558 $w=2.98e-07 $l=4.05e-07 $layer=LI1_cond $X=2.065 $Y=2.2
+ $X2=2.47 $Y2=2.2
r138 25 30 8.65646 $w=2.42e-07 $l=1.8775e-07 $layer=LI1_cond $X=3.475 $Y=2.2
+ $X2=3.39 $Y2=2.35
r139 25 48 20.4174 $w=2.42e-07 $l=4.05e-07 $layer=LI1_cond $X=3.475 $Y=2.2
+ $X2=3.475 $Y2=1.795
r140 25 28 32.0763 $w=2.98e-07 $l=8.35e-07 $layer=LI1_cond $X=3.305 $Y=2.2
+ $X2=2.47 $Y2=2.2
r141 23 51 27.1035 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=1.9 $Y=1.315
+ $X2=1.745 $Y2=1.315
r142 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.9
+ $Y=1.315 $X2=1.9 $Y2=1.315
r143 20 26 6.81904 $w=3e-07 $l=2.10357e-07 $layer=LI1_cond $X=1.92 $Y=2.05
+ $X2=2.065 $Y2=2.2
r144 20 22 29.2085 $w=2.88e-07 $l=7.35e-07 $layer=LI1_cond $X=1.92 $Y=2.05
+ $X2=1.92 $Y2=1.315
r145 17 49 39.3952 $w=3.9e-07 $l=2.27255e-07 $layer=POLY_cond $X=3.695 $Y=1.63
+ $X2=3.547 $Y2=1.795
r146 17 19 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.695 $Y=1.63
+ $X2=3.695 $Y2=0.995
r147 16 57 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.695 $Y=0.515
+ $X2=3.695 $Y2=0.35
r148 16 19 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.695 $Y=0.515
+ $X2=3.695 $Y2=0.995
r149 13 49 49.9004 $w=3.9e-07 $l=2.68328e-07 $layer=POLY_cond $X=3.585 $Y=2.045
+ $X2=3.547 $Y2=1.795
r150 13 15 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=3.585 $Y=2.045
+ $X2=3.585 $Y2=2.54
r151 10 29 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=2.545 $Y=2.465
+ $X2=2.47 $Y2=2.215
r152 10 12 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.545 $Y=2.465
+ $X2=2.545 $Y2=2.75
r153 7 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.745 $Y=1.15
+ $X2=1.745 $Y2=1.315
r154 7 9 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.745 $Y=1.15
+ $X2=1.745 $Y2=0.72
r155 2 41 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=4.225
+ $Y=2.11 $X2=4.37 $Y2=2.255
r156 1 45 182 $w=1.7e-07 $l=3.80657e-07 $layer=licon1_NDIFF $count=1 $X=4.3
+ $Y=0.37 $X2=4.445 $Y2=0.685
.ends

.subckt PM_SKY130_FD_SC_LS__DLCLKP_4%A_334_338# 1 2 7 9 10 11 14 19 20 24 29 32
+ 34
c78 29 0 1.04843e-19 $X=3.91 $Y=2.265
c79 20 0 8.09841e-20 $X=2.47 $Y=1.445
r80 31 34 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=3.91 $Y=1.485 $X2=3.99
+ $Y2=1.485
r81 31 32 5.10546 $w=2.48e-07 $l=8.5e-08 $layer=LI1_cond $X=3.91 $Y=1.485
+ $X2=3.825 $Y2=1.485
r82 27 29 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=3.81 $Y=2.265 $X2=3.91
+ $Y2=2.265
r83 24 38 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=2.47 $Y=1.64
+ $X2=2.47 $Y2=1.765
r84 24 37 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.47 $Y=1.64
+ $X2=2.47 $Y2=1.475
r85 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.47
+ $Y=1.64 $X2=2.47 $Y2=1.64
r86 20 23 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=2.47 $Y=1.445
+ $X2=2.47 $Y2=1.64
r87 19 29 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.91 $Y=2.18
+ $X2=3.91 $Y2=2.265
r88 18 31 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.91 $Y=1.61
+ $X2=3.91 $Y2=1.485
r89 18 19 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=3.91 $Y=1.61
+ $X2=3.91 $Y2=2.18
r90 17 20 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.635 $Y=1.445
+ $X2=2.47 $Y2=1.445
r91 17 32 77.6364 $w=1.68e-07 $l=1.19e-06 $layer=LI1_cond $X=2.635 $Y=1.445
+ $X2=3.825 $Y2=1.445
r92 14 37 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=2.38 $Y=0.83
+ $X2=2.38 $Y2=1.475
r93 10 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.305 $Y=1.765
+ $X2=2.47 $Y2=1.765
r94 10 11 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=2.305 $Y=1.765
+ $X2=1.85 $Y2=1.765
r95 7 11 26.9307 $w=1.5e-07 $l=1.58745e-07 $layer=POLY_cond $X=1.76 $Y=1.885
+ $X2=1.85 $Y2=1.765
r96 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.76 $Y=1.885
+ $X2=1.76 $Y2=2.46
r97 2 27 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=3.66
+ $Y=2.12 $X2=3.81 $Y2=2.265
r98 1 34 182 $w=1.7e-07 $l=9.23472e-07 $layer=licon1_NDIFF $count=1 $X=3.77
+ $Y=0.625 $X2=3.99 $Y2=1.445
.ends

.subckt PM_SKY130_FD_SC_LS__DLCLKP_4%A_27_74# 1 2 7 8 9 11 15 18 20 22 26 32 34
+ 37 38 39 40 41 42 43 45 47 48 51
c139 41 0 9.8676e-20 $X=2.98 $Y=1.02
c140 40 0 1.39534e-19 $X=2.98 $Y=0.425
c141 15 0 8.09841e-20 $X=2.98 $Y=1.155
c142 8 0 1.04843e-19 $X=2.965 $Y=2.375
r143 54 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.64
+ $Y=1.465 $X2=5.64 $Y2=1.465
r144 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.98
+ $Y=0.38 $X2=2.98 $Y2=0.38
r145 47 48 6.41202 $w=4.23e-07 $l=1.65e-07 $layer=LI1_cond $X=0.327 $Y=1.985
+ $X2=0.327 $Y2=1.82
r146 42 54 11.8065 $w=3.72e-07 $l=4.76991e-07 $layer=LI1_cond $X=5.26 $Y=1.105
+ $X2=5.532 $Y2=1.465
r147 42 43 137.984 $w=1.68e-07 $l=2.115e-06 $layer=LI1_cond $X=5.26 $Y=1.105
+ $X2=3.145 $Y2=1.105
r148 41 43 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.98 $Y=1.02
+ $X2=3.145 $Y2=1.105
r149 40 50 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.98 $Y=0.425
+ $X2=2.98 $Y2=0.34
r150 40 41 20.7789 $w=3.28e-07 $l=5.95e-07 $layer=LI1_cond $X=2.98 $Y=0.425
+ $X2=2.98 $Y2=1.02
r151 38 50 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.815 $Y=0.34
+ $X2=2.98 $Y2=0.34
r152 38 39 101.123 $w=1.68e-07 $l=1.55e-06 $layer=LI1_cond $X=2.815 $Y=0.34
+ $X2=1.265 $Y2=0.34
r153 36 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.18 $Y=0.425
+ $X2=1.265 $Y2=0.34
r154 36 37 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=1.18 $Y=0.425
+ $X2=1.18 $Y2=0.85
r155 35 45 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.365 $Y=0.935
+ $X2=0.24 $Y2=0.935
r156 34 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.095 $Y=0.935
+ $X2=1.18 $Y2=0.85
r157 34 35 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.095 $Y=0.935
+ $X2=0.365 $Y2=0.935
r158 30 47 1.27447 $w=4.23e-07 $l=4.7e-08 $layer=LI1_cond $X=0.327 $Y=2.032
+ $X2=0.327 $Y2=1.985
r159 30 32 21.2321 $w=4.23e-07 $l=7.83e-07 $layer=LI1_cond $X=0.327 $Y=2.032
+ $X2=0.327 $Y2=2.815
r160 28 45 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.24 $Y=1.02
+ $X2=0.24 $Y2=0.935
r161 28 48 36.8782 $w=2.48e-07 $l=8e-07 $layer=LI1_cond $X=0.24 $Y=1.02 $X2=0.24
+ $Y2=1.82
r162 24 45 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.24 $Y=0.85
+ $X2=0.24 $Y2=0.935
r163 24 26 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=0.24 $Y=0.85
+ $X2=0.24 $Y2=0.515
r164 20 55 61.4066 $w=2.86e-07 $l=3.04959e-07 $layer=POLY_cond $X=5.63 $Y=1.765
+ $X2=5.64 $Y2=1.465
r165 20 22 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.63 $Y=1.765
+ $X2=5.63 $Y2=2.4
r166 16 55 38.6549 $w=2.86e-07 $l=2.05122e-07 $layer=POLY_cond $X=5.55 $Y=1.3
+ $X2=5.64 $Y2=1.465
r167 16 18 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=5.55 $Y=1.3
+ $X2=5.55 $Y2=0.74
r168 15 23 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.98 $Y=1.155
+ $X2=2.98 $Y2=1.44
r169 12 51 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.98 $Y=0.545
+ $X2=2.98 $Y2=0.38
r170 12 15 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.98 $Y=0.545
+ $X2=2.98 $Y2=1.155
r171 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.965 $Y=2.465
+ $X2=2.965 $Y2=2.75
r172 8 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.965 $Y=2.375
+ $X2=2.965 $Y2=2.465
r173 7 23 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.965 $Y=1.53
+ $X2=2.965 $Y2=1.44
r174 7 8 328.46 $w=1.8e-07 $l=8.45e-07 $layer=POLY_cond $X=2.965 $Y=1.53
+ $X2=2.965 $Y2=2.375
r175 2 47 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.23
+ $Y=1.84 $X2=0.375 $Y2=1.985
r176 2 32 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.23
+ $Y=1.84 $X2=0.375 $Y2=2.815
r177 1 45 182 $w=1.7e-07 $l=6.63551e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.965
r178 1 26 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__DLCLKP_4%CLK 2 3 5 8 10 12 15 17 26 27
c47 26 0 1.80208e-19 $X=4.905 $Y=1.515
r48 27 28 2.07759 $w=3.48e-07 $l=1.5e-08 $layer=POLY_cond $X=5.145 $Y=1.557
+ $X2=5.16 $Y2=1.557
r49 25 27 33.2414 $w=3.48e-07 $l=2.4e-07 $layer=POLY_cond $X=4.905 $Y=1.557
+ $X2=5.145 $Y2=1.557
r50 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.905
+ $Y=1.515 $X2=4.905 $Y2=1.515
r51 23 25 24.2385 $w=3.48e-07 $l=1.75e-07 $layer=POLY_cond $X=4.73 $Y=1.557
+ $X2=4.905 $Y2=1.557
r52 21 26 9.3293 $w=4.18e-07 $l=3.4e-07 $layer=LI1_cond $X=4.565 $Y=1.57
+ $X2=4.905 $Y2=1.57
r53 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.565
+ $Y=1.515 $X2=4.565 $Y2=1.515
r54 17 21 0.137196 $w=4.18e-07 $l=5e-09 $layer=LI1_cond $X=4.56 $Y=1.57
+ $X2=4.565 $Y2=1.57
r55 13 28 22.4912 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.16 $Y=1.35
+ $X2=5.16 $Y2=1.557
r56 13 15 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.16 $Y=1.35
+ $X2=5.16 $Y2=0.74
r57 10 27 22.4912 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=5.145 $Y=1.765
+ $X2=5.145 $Y2=1.557
r58 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.145 $Y=1.765
+ $X2=5.145 $Y2=2.4
r59 6 23 22.4912 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.73 $Y=1.35
+ $X2=4.73 $Y2=1.557
r60 6 8 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.73 $Y=1.35 $X2=4.73
+ $Y2=0.74
r61 3 5 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=4.595 $Y=2.035
+ $X2=4.595 $Y2=2.53
r62 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=4.595 $Y=1.945 $X2=4.595
+ $Y2=2.035
r63 1 23 18.6983 $w=3.48e-07 $l=1.35e-07 $layer=POLY_cond $X=4.595 $Y=1.557
+ $X2=4.73 $Y2=1.557
r64 1 20 4.15517 $w=3.48e-07 $l=3e-08 $layer=POLY_cond $X=4.595 $Y=1.557
+ $X2=4.565 $Y2=1.557
r65 1 2 103.008 $w=1.8e-07 $l=2.65e-07 $layer=POLY_cond $X=4.595 $Y=1.68
+ $X2=4.595 $Y2=1.945
.ends

.subckt PM_SKY130_FD_SC_LS__DLCLKP_4%A_1044_368# 1 2 7 9 11 14 16 18 21 23 24 25
+ 27 30 32 34 37 45 47 49 51 53 56 64 65
c120 45 0 1.31164e-19 $X=8.135 $Y=1.582
c121 24 0 1.35311e-19 $X=7.29 $Y=1.54
c122 16 0 4.22657e-20 $X=7.2 $Y=1.765
r123 64 65 98.7966 $w=3.3e-07 $l=5.65e-07 $layer=POLY_cond $X=6.185 $Y=0.835
+ $X2=6.185 $Y2=1.4
r124 63 64 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=6.185
+ $Y=0.835 $X2=6.185 $Y2=0.835
r125 61 63 6.55034 $w=5.96e-07 $l=3.2e-07 $layer=LI1_cond $X=5.975 $Y=0.515
+ $X2=5.975 $Y2=0.835
r126 57 65 12.47 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=6.185 $Y=1.54
+ $X2=6.185 $Y2=1.4
r127 56 57 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=6.185
+ $Y=1.515 $X2=6.185 $Y2=1.515
r128 54 56 9.3732 $w=3.73e-07 $l=3.05e-07 $layer=LI1_cond $X=6.162 $Y=1.82
+ $X2=6.162 $Y2=1.515
r129 53 63 7.70783 $w=5.96e-07 $l=3.77081e-07 $layer=LI1_cond $X=6.162 $Y=1.13
+ $X2=5.975 $Y2=0.835
r130 53 56 11.8317 $w=3.73e-07 $l=3.85e-07 $layer=LI1_cond $X=6.162 $Y=1.13
+ $X2=6.162 $Y2=1.515
r131 52 59 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.57 $Y=1.905
+ $X2=5.405 $Y2=1.905
r132 51 54 8.1532 $w=1.7e-07 $l=2.2553e-07 $layer=LI1_cond $X=5.975 $Y=1.905
+ $X2=6.162 $Y2=1.82
r133 51 52 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=5.975 $Y=1.905
+ $X2=5.57 $Y2=1.905
r134 47 59 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.405 $Y=1.99
+ $X2=5.405 $Y2=1.905
r135 47 49 28.8111 $w=3.28e-07 $l=8.25e-07 $layer=LI1_cond $X=5.405 $Y=1.99
+ $X2=5.405 $Y2=2.815
r136 45 46 1.47401 $w=3.27e-07 $l=1e-08 $layer=POLY_cond $X=8.135 $Y=1.582
+ $X2=8.145 $Y2=1.582
r137 44 45 61.9083 $w=3.27e-07 $l=4.2e-07 $layer=POLY_cond $X=7.715 $Y=1.582
+ $X2=8.135 $Y2=1.582
r138 43 44 4.42202 $w=3.27e-07 $l=3e-08 $layer=POLY_cond $X=7.685 $Y=1.582
+ $X2=7.715 $Y2=1.582
r139 41 42 2.21101 $w=3.27e-07 $l=1.5e-08 $layer=POLY_cond $X=7.2 $Y=1.582
+ $X2=7.215 $Y2=1.582
r140 40 41 61.1713 $w=3.27e-07 $l=4.15e-07 $layer=POLY_cond $X=6.785 $Y=1.582
+ $X2=7.2 $Y2=1.582
r141 39 40 7.37003 $w=3.27e-07 $l=5e-08 $layer=POLY_cond $X=6.735 $Y=1.582
+ $X2=6.785 $Y2=1.582
r142 35 46 21.0057 $w=1.5e-07 $l=1.82e-07 $layer=POLY_cond $X=8.145 $Y=1.4
+ $X2=8.145 $Y2=1.582
r143 35 37 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.145 $Y=1.4
+ $X2=8.145 $Y2=0.74
r144 32 45 21.0057 $w=1.5e-07 $l=1.83e-07 $layer=POLY_cond $X=8.135 $Y=1.765
+ $X2=8.135 $Y2=1.582
r145 32 34 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.135 $Y=1.765
+ $X2=8.135 $Y2=2.4
r146 28 44 21.0057 $w=1.5e-07 $l=1.82e-07 $layer=POLY_cond $X=7.715 $Y=1.4
+ $X2=7.715 $Y2=1.582
r147 28 30 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.715 $Y=1.4
+ $X2=7.715 $Y2=0.74
r148 25 43 21.0057 $w=1.5e-07 $l=1.83e-07 $layer=POLY_cond $X=7.685 $Y=1.765
+ $X2=7.685 $Y2=1.582
r149 25 27 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.685 $Y=1.765
+ $X2=7.685 $Y2=2.4
r150 24 42 12.1866 $w=3.27e-07 $l=9.3675e-08 $layer=POLY_cond $X=7.29 $Y=1.54
+ $X2=7.215 $Y2=1.582
r151 23 43 14.3976 $w=3.27e-07 $l=1.08995e-07 $layer=POLY_cond $X=7.595 $Y=1.54
+ $X2=7.685 $Y2=1.582
r152 23 24 65.3429 $w=2.8e-07 $l=3.05e-07 $layer=POLY_cond $X=7.595 $Y=1.54
+ $X2=7.29 $Y2=1.54
r153 19 42 21.0057 $w=1.5e-07 $l=1.82e-07 $layer=POLY_cond $X=7.215 $Y=1.4
+ $X2=7.215 $Y2=1.582
r154 19 21 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.215 $Y=1.4
+ $X2=7.215 $Y2=0.74
r155 16 41 21.0057 $w=1.5e-07 $l=1.83e-07 $layer=POLY_cond $X=7.2 $Y=1.765
+ $X2=7.2 $Y2=1.582
r156 16 18 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.2 $Y=1.765
+ $X2=7.2 $Y2=2.4
r157 12 40 21.0057 $w=1.5e-07 $l=1.82e-07 $layer=POLY_cond $X=6.785 $Y=1.4
+ $X2=6.785 $Y2=1.582
r158 12 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.785 $Y=1.4
+ $X2=6.785 $Y2=0.74
r159 9 39 21.0057 $w=1.5e-07 $l=1.83e-07 $layer=POLY_cond $X=6.735 $Y=1.765
+ $X2=6.735 $Y2=1.582
r160 9 11 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.735 $Y=1.765
+ $X2=6.735 $Y2=2.4
r161 8 57 14.6968 $w=2.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.35 $Y=1.54
+ $X2=6.185 $Y2=1.54
r162 7 39 14.3976 $w=3.27e-07 $l=1.08995e-07 $layer=POLY_cond $X=6.645 $Y=1.54
+ $X2=6.735 $Y2=1.582
r163 7 8 63.2005 $w=2.8e-07 $l=2.95e-07 $layer=POLY_cond $X=6.645 $Y=1.54
+ $X2=6.35 $Y2=1.54
r164 2 59 400 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=1 $X=5.22
+ $Y=1.84 $X2=5.405 $Y2=1.985
r165 2 49 400 $w=1.7e-07 $l=1.06348e-06 $layer=licon1_PDIFF $count=1 $X=5.22
+ $Y=1.84 $X2=5.405 $Y2=2.815
r166 1 61 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.625
+ $Y=0.37 $X2=5.765 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__DLCLKP_4%VPWR 1 2 3 4 5 6 21 25 29 33 37 41 43 48 49
+ 51 52 53 59 70 74 79 85 88 91 95
r102 94 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33 $X2=8.4
+ $Y2=3.33
r103 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r104 88 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r105 85 86 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r106 83 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r107 83 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=7.44 $Y2=3.33
r108 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r109 80 91 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.545 $Y=3.33
+ $X2=7.42 $Y2=3.33
r110 80 82 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=7.545 $Y=3.33
+ $X2=7.92 $Y2=3.33
r111 79 94 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=8.195 $Y=3.33
+ $X2=8.417 $Y2=3.33
r112 79 82 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=8.195 $Y=3.33
+ $X2=7.92 $Y2=3.33
r113 78 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.44 $Y2=3.33
r114 78 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6.48 $Y2=3.33
r115 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r116 75 88 15.3799 $w=1.7e-07 $l=4.43e-07 $layer=LI1_cond $X=6.625 $Y=3.33
+ $X2=6.182 $Y2=3.33
r117 75 77 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=6.625 $Y=3.33
+ $X2=6.96 $Y2=3.33
r118 74 91 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.295 $Y=3.33
+ $X2=7.42 $Y2=3.33
r119 74 77 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=7.295 $Y=3.33
+ $X2=6.96 $Y2=3.33
r120 73 89 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6.48 $Y2=3.33
r121 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r122 70 88 15.3799 $w=1.7e-07 $l=4.42e-07 $layer=LI1_cond $X=5.74 $Y=3.33
+ $X2=6.182 $Y2=3.33
r123 70 72 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=5.74 $Y=3.33
+ $X2=5.52 $Y2=3.33
r124 69 73 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r125 68 69 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r126 66 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r127 65 68 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.6 $Y=3.33 $X2=4.56
+ $Y2=3.33
r128 65 66 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r129 63 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.44 $Y=3.33
+ $X2=3.275 $Y2=3.33
r130 63 65 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=3.44 $Y=3.33
+ $X2=3.6 $Y2=3.33
r131 62 86 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=3.12 $Y2=3.33
r132 61 62 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r133 59 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.11 $Y=3.33
+ $X2=3.275 $Y2=3.33
r134 59 61 124.61 $w=1.68e-07 $l=1.91e-06 $layer=LI1_cond $X=3.11 $Y=3.33
+ $X2=1.2 $Y2=3.33
r135 57 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r136 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r137 53 69 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=3.33
+ $X2=4.56 $Y2=3.33
r138 53 66 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=4.32 $Y=3.33
+ $X2=3.6 $Y2=3.33
r139 51 68 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=4.74 $Y=3.33
+ $X2=4.56 $Y2=3.33
r140 51 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.74 $Y=3.33
+ $X2=4.905 $Y2=3.33
r141 50 72 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=5.07 $Y=3.33
+ $X2=5.52 $Y2=3.33
r142 50 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.07 $Y=3.33
+ $X2=4.905 $Y2=3.33
r143 48 56 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=0.785 $Y=3.33
+ $X2=0.72 $Y2=3.33
r144 48 49 9.39981 $w=1.7e-07 $l=1.87e-07 $layer=LI1_cond $X=0.785 $Y=3.33
+ $X2=0.972 $Y2=3.33
r145 47 61 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=1.16 $Y=3.33 $X2=1.2
+ $Y2=3.33
r146 47 49 9.39981 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=1.16 $Y=3.33
+ $X2=0.972 $Y2=3.33
r147 43 46 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=8.36 $Y=2.035
+ $X2=8.36 $Y2=2.815
r148 41 94 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=8.36 $Y=3.245
+ $X2=8.417 $Y2=3.33
r149 41 46 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=8.36 $Y=3.245
+ $X2=8.36 $Y2=2.815
r150 37 40 35.0343 $w=2.48e-07 $l=7.6e-07 $layer=LI1_cond $X=7.42 $Y=2.055
+ $X2=7.42 $Y2=2.815
r151 35 91 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.42 $Y=3.245
+ $X2=7.42 $Y2=3.33
r152 35 40 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=7.42 $Y=3.245
+ $X2=7.42 $Y2=2.815
r153 31 88 3.31993 $w=8.85e-07 $l=8.5e-08 $layer=LI1_cond $X=6.182 $Y=3.245
+ $X2=6.182 $Y2=3.33
r154 31 33 13.5785 $w=8.83e-07 $l=9.85e-07 $layer=LI1_cond $X=6.182 $Y=3.245
+ $X2=6.182 $Y2=2.26
r155 27 52 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.905 $Y=3.245
+ $X2=4.905 $Y2=3.33
r156 27 29 34.5733 $w=3.28e-07 $l=9.9e-07 $layer=LI1_cond $X=4.905 $Y=3.245
+ $X2=4.905 $Y2=2.255
r157 23 85 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.275 $Y=3.245
+ $X2=3.275 $Y2=3.33
r158 23 25 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=3.275 $Y=3.245
+ $X2=3.275 $Y2=3.025
r159 19 49 1.28102 $w=3.75e-07 $l=8.5e-08 $layer=LI1_cond $X=0.972 $Y=3.245
+ $X2=0.972 $Y2=3.33
r160 19 21 25.6611 $w=3.73e-07 $l=8.35e-07 $layer=LI1_cond $X=0.972 $Y=3.245
+ $X2=0.972 $Y2=2.41
r161 6 46 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=8.21
+ $Y=1.84 $X2=8.36 $Y2=2.815
r162 6 43 400 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=8.21
+ $Y=1.84 $X2=8.36 $Y2=2.035
r163 5 40 400 $w=1.7e-07 $l=1.06348e-06 $layer=licon1_PDIFF $count=1 $X=7.275
+ $Y=1.84 $X2=7.46 $Y2=2.815
r164 5 37 400 $w=1.7e-07 $l=2.93258e-07 $layer=licon1_PDIFF $count=1 $X=7.275
+ $Y=1.84 $X2=7.46 $Y2=2.055
r165 4 33 150 $w=1.7e-07 $l=9.41873e-07 $layer=licon1_PDIFF $count=4 $X=5.705
+ $Y=1.84 $X2=6.46 $Y2=2.26
r166 3 29 300 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=2 $X=4.67
+ $Y=2.11 $X2=4.905 $Y2=2.255
r167 2 25 600 $w=1.7e-07 $l=5.90931e-07 $layer=licon1_PDIFF $count=1 $X=3.04
+ $Y=2.54 $X2=3.275 $Y2=3.025
r168 1 21 300 $w=1.7e-07 $l=7.00143e-07 $layer=licon1_PDIFF $count=2 $X=0.675
+ $Y=1.84 $X2=0.965 $Y2=2.41
.ends

.subckt PM_SKY130_FD_SC_LS__DLCLKP_4%GCLK 1 2 3 4 15 21 23 24 25 26 29 35 38 39
+ 40 41
c71 40 0 1.77576e-19 $X=7.92 $Y=1.665
c72 15 0 1.31164e-19 $X=6.96 $Y=1.985
r73 41 44 19.2909 $w=2.28e-07 $l=3.85e-07 $layer=LI1_cond $X=8.4 $Y=1.665
+ $X2=8.015 $Y2=1.665
r74 40 44 3.48671 $w=2.3e-07 $l=1.35e-07 $layer=LI1_cond $X=7.88 $Y=1.665
+ $X2=8.015 $Y2=1.665
r75 38 40 2.63492 $w=2.1e-07 $l=1.29132e-07 $layer=LI1_cond $X=7.91 $Y=1.55
+ $X2=7.88 $Y2=1.665
r76 37 39 3.98977 $w=2.3e-07 $l=9.44722e-08 $layer=LI1_cond $X=7.91 $Y=1.38
+ $X2=7.89 $Y2=1.295
r77 37 38 8.97835 $w=2.08e-07 $l=1.7e-07 $layer=LI1_cond $X=7.91 $Y=1.38
+ $X2=7.91 $Y2=1.55
r78 33 39 3.98977 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.89 $Y=1.21 $X2=7.89
+ $Y2=1.295
r79 33 35 32.0379 $w=2.48e-07 $l=6.95e-07 $layer=LI1_cond $X=7.89 $Y=1.21
+ $X2=7.89 $Y2=0.515
r80 29 31 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=7.87 $Y=1.985
+ $X2=7.87 $Y2=2.815
r81 27 40 2.63492 $w=2.5e-07 $l=1.19896e-07 $layer=LI1_cond $X=7.87 $Y=1.78
+ $X2=7.88 $Y2=1.665
r82 27 29 9.45003 $w=2.48e-07 $l=2.05e-07 $layer=LI1_cond $X=7.87 $Y=1.78
+ $X2=7.87 $Y2=1.985
r83 25 39 2.45049 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.765 $Y=1.295
+ $X2=7.89 $Y2=1.295
r84 25 26 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=7.765 $Y=1.295
+ $X2=7.165 $Y2=1.295
r85 23 40 3.48671 $w=1.7e-07 $l=1.49248e-07 $layer=LI1_cond $X=7.745 $Y=1.635
+ $X2=7.88 $Y2=1.665
r86 23 24 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=7.745 $Y=1.635
+ $X2=7.125 $Y2=1.635
r87 19 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7 $Y=1.21
+ $X2=7.165 $Y2=1.295
r88 19 21 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=7 $Y=1.21 $X2=7
+ $Y2=0.515
r89 15 17 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=6.96 $Y=1.985
+ $X2=6.96 $Y2=2.815
r90 13 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.96 $Y=1.72
+ $X2=7.125 $Y2=1.635
r91 13 15 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=6.96 $Y=1.72
+ $X2=6.96 $Y2=1.985
r92 4 31 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=7.76
+ $Y=1.84 $X2=7.91 $Y2=2.815
r93 4 29 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=7.76
+ $Y=1.84 $X2=7.91 $Y2=1.985
r94 3 17 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=6.81
+ $Y=1.84 $X2=6.96 $Y2=2.815
r95 3 15 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=6.81
+ $Y=1.84 $X2=6.96 $Y2=1.985
r96 2 35 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.79
+ $Y=0.37 $X2=7.93 $Y2=0.515
r97 1 21 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.86
+ $Y=0.37 $X2=7 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__DLCLKP_4%VGND 1 2 3 4 5 6 21 25 29 33 35 37 39 41 46
+ 54 59 64 69 75 78 81 91 95
r98 94 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r99 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r100 81 82 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r101 78 79 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r102 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r103 73 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.4
+ $Y2=0
r104 73 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=7.44
+ $Y2=0
r105 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r106 70 91 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.585 $Y=0 $X2=7.46
+ $Y2=0
r107 70 72 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=7.585 $Y=0
+ $X2=7.92 $Y2=0
r108 69 94 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=8.195 $Y=0
+ $X2=8.417 $Y2=0
r109 69 72 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=8.195 $Y=0
+ $X2=7.92 $Y2=0
r110 68 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r111 68 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=6.48
+ $Y2=0
r112 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r113 65 67 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=6.655 $Y=0
+ $X2=6.96 $Y2=0
r114 64 91 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.335 $Y=0 $X2=7.46
+ $Y2=0
r115 64 67 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=7.335 $Y=0
+ $X2=6.96 $Y2=0
r116 63 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r117 63 82 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.04
+ $Y2=0
r118 62 63 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r119 60 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.11 $Y=0 $X2=4.945
+ $Y2=0
r120 60 62 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=5.11 $Y=0 $X2=6
+ $Y2=0
r121 59 88 8.09467 $w=4.93e-07 $l=3.35e-07 $layer=LI1_cond $X=6.407 $Y=0
+ $X2=6.407 $Y2=0.335
r122 59 65 7.09362 $w=1.7e-07 $l=2.48e-07 $layer=LI1_cond $X=6.407 $Y=0
+ $X2=6.655 $Y2=0
r123 59 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r124 59 62 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=6.16 $Y=0 $X2=6
+ $Y2=0
r125 58 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r126 57 58 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r127 55 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.645 $Y=0 $X2=3.48
+ $Y2=0
r128 55 57 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=3.645 $Y=0
+ $X2=4.56 $Y2=0
r129 54 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.78 $Y=0 $X2=4.945
+ $Y2=0
r130 54 57 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=4.78 $Y=0 $X2=4.56
+ $Y2=0
r131 53 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r132 52 53 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r133 50 53 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r134 50 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r135 49 52 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r136 49 50 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r137 47 75 9.39981 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=0.925 $Y=0
+ $X2=0.737 $Y2=0
r138 47 49 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.925 $Y=0 $X2=1.2
+ $Y2=0
r139 46 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.315 $Y=0 $X2=3.48
+ $Y2=0
r140 46 52 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=3.315 $Y=0
+ $X2=3.12 $Y2=0
r141 44 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r142 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r143 41 75 9.39981 $w=1.7e-07 $l=1.87e-07 $layer=LI1_cond $X=0.55 $Y=0 $X2=0.737
+ $Y2=0
r144 41 43 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.55 $Y=0 $X2=0.24
+ $Y2=0
r145 39 58 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=0
+ $X2=4.56 $Y2=0
r146 39 79 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=4.32 $Y=0 $X2=3.6
+ $Y2=0
r147 35 94 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=8.36 $Y=0.085
+ $X2=8.417 $Y2=0
r148 35 37 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=8.36 $Y=0.085
+ $X2=8.36 $Y2=0.515
r149 31 91 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.46 $Y=0.085
+ $X2=7.46 $Y2=0
r150 31 33 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=7.46 $Y=0.085
+ $X2=7.46 $Y2=0.515
r151 27 81 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.945 $Y=0.085
+ $X2=4.945 $Y2=0
r152 27 29 20.9535 $w=3.28e-07 $l=6e-07 $layer=LI1_cond $X=4.945 $Y=0.085
+ $X2=4.945 $Y2=0.685
r153 23 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.48 $Y=0.085
+ $X2=3.48 $Y2=0
r154 23 25 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=3.48 $Y=0.085
+ $X2=3.48 $Y2=0.765
r155 19 75 1.28102 $w=3.75e-07 $l=8.5e-08 $layer=LI1_cond $X=0.737 $Y=0.085
+ $X2=0.737 $Y2=0
r156 19 21 13.2147 $w=3.73e-07 $l=4.3e-07 $layer=LI1_cond $X=0.737 $Y=0.085
+ $X2=0.737 $Y2=0.515
r157 6 37 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.22
+ $Y=0.37 $X2=8.36 $Y2=0.515
r158 5 33 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=7.29
+ $Y=0.37 $X2=7.5 $Y2=0.515
r159 4 88 182 $w=1.7e-07 $l=2.88531e-07 $layer=licon1_NDIFF $count=1 $X=6.18
+ $Y=0.19 $X2=6.405 $Y2=0.335
r160 3 29 182 $w=1.7e-07 $l=3.78583e-07 $layer=licon1_NDIFF $count=1 $X=4.805
+ $Y=0.37 $X2=4.945 $Y2=0.685
r161 2 25 182 $w=1.7e-07 $l=5.07075e-07 $layer=licon1_NDIFF $count=1 $X=3.055
+ $Y=0.945 $X2=3.48 $Y2=0.765
r162 1 21 182 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.735 $Y2=0.515
.ends

