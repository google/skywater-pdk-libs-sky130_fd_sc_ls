# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ls__o22a_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ls__o22a_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.720000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.845000 1.450000 2.275000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.845000 1.450000 1.515000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 0.255000 2.610000 0.570000 ;
        RECT 2.045000 0.570000 2.275000 0.670000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525000 1.450000 3.505000 1.780000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  1.125600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.600000 1.850000 6.105000 2.020000 ;
        RECT 4.600000 2.020000 4.930000 2.980000 ;
        RECT 4.980000 0.350000 5.230000 1.010000 ;
        RECT 4.980000 1.010000 6.105000 1.180000 ;
        RECT 5.775000 2.020000 6.105000 2.980000 ;
        RECT 5.920000 0.350000 6.105000 1.010000 ;
        RECT 5.935000 1.180000 6.595000 1.410000 ;
        RECT 5.935000 1.410000 6.105000 1.850000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.720000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 6.720000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.720000 0.085000 ;
      RECT 0.000000  3.245000 6.720000 3.415000 ;
      RECT 0.115000  0.660000 0.445000 1.110000 ;
      RECT 0.115000  1.110000 4.240000 1.280000 ;
      RECT 0.115000  1.280000 0.445000 1.340000 ;
      RECT 0.115000  1.940000 0.365000 3.245000 ;
      RECT 0.565000  1.950000 0.895000 2.905000 ;
      RECT 0.565000  2.905000 1.895000 3.075000 ;
      RECT 0.615000  0.085000 0.945000 0.940000 ;
      RECT 1.065000  1.950000 3.845000 2.120000 ;
      RECT 1.065000  2.120000 1.395000 2.735000 ;
      RECT 1.125000  0.660000 1.375000 1.110000 ;
      RECT 1.545000  0.085000 1.875000 0.940000 ;
      RECT 1.565000  2.290000 1.895000 2.905000 ;
      RECT 2.045000  0.840000 2.375000 1.090000 ;
      RECT 2.045000  1.090000 4.240000 1.110000 ;
      RECT 2.065000  2.290000 2.395000 3.245000 ;
      RECT 2.545000  0.740000 3.810000 0.750000 ;
      RECT 2.545000  0.750000 4.585000 0.920000 ;
      RECT 2.565000  2.290000 2.895000 2.905000 ;
      RECT 2.565000  2.905000 3.895000 3.075000 ;
      RECT 3.065000  2.120000 3.395000 2.735000 ;
      RECT 3.480000  0.660000 3.810000 0.740000 ;
      RECT 3.565000  2.290000 3.895000 2.905000 ;
      RECT 3.675000  1.510000 5.765000 1.680000 ;
      RECT 3.675000  1.680000 3.845000 1.950000 ;
      RECT 3.910000  1.280000 4.240000 1.340000 ;
      RECT 4.100000  1.850000 4.430000 3.245000 ;
      RECT 4.415000  0.920000 4.585000 1.350000 ;
      RECT 4.415000  1.350000 5.765000 1.510000 ;
      RECT 4.470000  0.085000 4.800000 0.580000 ;
      RECT 5.200000  2.190000 5.530000 3.245000 ;
      RECT 5.410000  0.085000 5.740000 0.790000 ;
      RECT 6.275000  0.085000 6.605000 1.010000 ;
      RECT 6.275000  1.820000 6.605000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
  END
END sky130_fd_sc_ls__o22a_4
