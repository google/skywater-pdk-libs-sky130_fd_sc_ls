* File: sky130_fd_sc_ls__clkinv_16.pxi.spice
* Created: Wed Sep  2 10:58:36 2020
* 
x_PM_SKY130_FD_SC_LS__CLKINV_16%A N_A_M1002_g N_A_c_182_n N_A_M1000_g
+ N_A_M1003_g N_A_c_183_n N_A_M1001_g N_A_M1004_g N_A_c_184_n N_A_M1005_g
+ N_A_M1008_g N_A_c_185_n N_A_M1006_g N_A_M1011_g N_A_c_186_n N_A_M1007_g
+ N_A_M1012_g N_A_c_187_n N_A_M1009_g N_A_c_188_n N_A_M1010_g N_A_M1016_g
+ N_A_M1017_g N_A_c_189_n N_A_M1013_g N_A_c_190_n N_A_M1014_g N_A_M1021_g
+ N_A_c_191_n N_A_M1015_g N_A_M1022_g N_A_c_192_n N_A_M1018_g N_A_M1026_g
+ N_A_c_193_n N_A_M1019_g N_A_M1029_g N_A_c_194_n N_A_M1020_g N_A_M1030_g
+ N_A_c_195_n N_A_M1023_g N_A_M1034_g N_A_c_196_n N_A_M1024_g N_A_M1036_g
+ N_A_M1039_g N_A_c_197_n N_A_M1025_g N_A_c_198_n N_A_M1027_g N_A_c_199_n
+ N_A_M1028_g N_A_c_200_n N_A_M1031_g N_A_c_201_n N_A_M1032_g N_A_c_202_n
+ N_A_M1033_g N_A_c_203_n N_A_M1035_g N_A_c_204_n N_A_M1037_g N_A_c_205_n
+ N_A_M1038_g A N_A_c_172_n N_A_c_173_n N_A_c_174_n N_A_c_175_n N_A_c_176_n
+ N_A_c_177_n N_A_c_178_n N_A_c_179_n N_A_c_180_n N_A_c_181_n
+ PM_SKY130_FD_SC_LS__CLKINV_16%A
x_PM_SKY130_FD_SC_LS__CLKINV_16%VPWR N_VPWR_M1000_d N_VPWR_M1001_d
+ N_VPWR_M1006_d N_VPWR_M1009_d N_VPWR_M1013_d N_VPWR_M1015_d N_VPWR_M1019_d
+ N_VPWR_M1023_d N_VPWR_M1025_d N_VPWR_M1028_d N_VPWR_M1032_d N_VPWR_M1035_d
+ N_VPWR_M1038_d N_VPWR_c_574_n N_VPWR_c_575_n N_VPWR_c_576_n N_VPWR_c_577_n
+ N_VPWR_c_578_n N_VPWR_c_579_n N_VPWR_c_580_n N_VPWR_c_581_n N_VPWR_c_582_n
+ N_VPWR_c_583_n N_VPWR_c_584_n N_VPWR_c_585_n N_VPWR_c_586_n N_VPWR_c_587_n
+ N_VPWR_c_588_n N_VPWR_c_589_n N_VPWR_c_590_n N_VPWR_c_591_n N_VPWR_c_592_n
+ N_VPWR_c_593_n N_VPWR_c_594_n N_VPWR_c_595_n N_VPWR_c_596_n N_VPWR_c_597_n
+ N_VPWR_c_598_n N_VPWR_c_599_n N_VPWR_c_600_n N_VPWR_c_601_n N_VPWR_c_602_n
+ N_VPWR_c_603_n N_VPWR_c_604_n N_VPWR_c_605_n VPWR N_VPWR_c_606_n
+ N_VPWR_c_607_n N_VPWR_c_608_n N_VPWR_c_609_n N_VPWR_c_610_n N_VPWR_c_611_n
+ N_VPWR_c_573_n PM_SKY130_FD_SC_LS__CLKINV_16%VPWR
x_PM_SKY130_FD_SC_LS__CLKINV_16%Y N_Y_M1002_s N_Y_M1004_s N_Y_M1011_s
+ N_Y_M1016_s N_Y_M1021_s N_Y_M1026_s N_Y_M1030_s N_Y_M1036_s N_Y_M1000_s
+ N_Y_M1005_s N_Y_M1007_s N_Y_M1010_s N_Y_M1014_s N_Y_M1018_s N_Y_M1020_s
+ N_Y_M1024_s N_Y_M1027_s N_Y_M1031_s N_Y_M1033_s N_Y_M1037_s N_Y_c_806_n
+ N_Y_c_822_n N_Y_c_823_n N_Y_c_807_n N_Y_c_808_n N_Y_c_809_n N_Y_c_810_n
+ N_Y_c_826_n N_Y_c_811_n N_Y_c_812_n N_Y_c_813_n N_Y_c_814_n N_Y_c_888_n
+ N_Y_c_892_n N_Y_c_815_n N_Y_c_816_n N_Y_c_817_n N_Y_c_912_n Y N_Y_c_829_n
+ N_Y_c_818_n N_Y_c_831_n N_Y_c_832_n N_Y_c_833_n N_Y_c_819_n N_Y_c_835_n
+ N_Y_c_836_n N_Y_c_837_n N_Y_c_838_n N_Y_c_956_n N_Y_c_989_n N_Y_c_820_n
+ N_Y_c_1002_n N_Y_c_821_n PM_SKY130_FD_SC_LS__CLKINV_16%Y
x_PM_SKY130_FD_SC_LS__CLKINV_16%VGND N_VGND_M1002_d N_VGND_M1003_d
+ N_VGND_M1008_d N_VGND_M1012_d N_VGND_M1017_d N_VGND_M1022_d N_VGND_M1029_d
+ N_VGND_M1034_d N_VGND_M1039_d N_VGND_c_1131_n N_VGND_c_1132_n N_VGND_c_1133_n
+ N_VGND_c_1134_n N_VGND_c_1135_n N_VGND_c_1136_n N_VGND_c_1137_n
+ N_VGND_c_1138_n N_VGND_c_1139_n N_VGND_c_1140_n N_VGND_c_1141_n
+ N_VGND_c_1142_n N_VGND_c_1143_n N_VGND_c_1144_n N_VGND_c_1145_n
+ N_VGND_c_1146_n N_VGND_c_1147_n N_VGND_c_1148_n N_VGND_c_1149_n
+ N_VGND_c_1150_n N_VGND_c_1151_n N_VGND_c_1152_n N_VGND_c_1153_n
+ N_VGND_c_1154_n N_VGND_c_1155_n VGND N_VGND_c_1156_n N_VGND_c_1157_n
+ N_VGND_c_1158_n N_VGND_c_1159_n PM_SKY130_FD_SC_LS__CLKINV_16%VGND
cc_1 VNB N_A_M1002_g 0.0516017f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.61
cc_2 VNB N_A_M1003_g 0.034419f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.61
cc_3 VNB N_A_M1004_g 0.0344887f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=0.61
cc_4 VNB N_A_M1008_g 0.0363131f $X=-0.19 $Y=-0.245 $X2=1.785 $Y2=0.61
cc_5 VNB N_A_M1011_g 0.0362251f $X=-0.19 $Y=-0.245 $X2=2.285 $Y2=0.61
cc_6 VNB N_A_M1012_g 0.0348055f $X=-0.19 $Y=-0.245 $X2=2.715 $Y2=0.61
cc_7 VNB N_A_M1016_g 0.0361753f $X=-0.19 $Y=-0.245 $X2=3.215 $Y2=0.61
cc_8 VNB N_A_M1017_g 0.0363124f $X=-0.19 $Y=-0.245 $X2=3.645 $Y2=0.61
cc_9 VNB N_A_M1021_g 0.0363124f $X=-0.19 $Y=-0.245 $X2=4.215 $Y2=0.61
cc_10 VNB N_A_M1022_g 0.0378286f $X=-0.19 $Y=-0.245 $X2=4.645 $Y2=0.61
cc_11 VNB N_A_M1026_g 0.0363229f $X=-0.19 $Y=-0.245 $X2=5.215 $Y2=0.61
cc_12 VNB N_A_M1029_g 0.0339185f $X=-0.19 $Y=-0.245 $X2=5.645 $Y2=0.61
cc_13 VNB N_A_M1030_g 0.0339399f $X=-0.19 $Y=-0.245 $X2=6.075 $Y2=0.61
cc_14 VNB N_A_M1034_g 0.0339103f $X=-0.19 $Y=-0.245 $X2=6.505 $Y2=0.61
cc_15 VNB N_A_M1036_g 0.0338885f $X=-0.19 $Y=-0.245 $X2=6.935 $Y2=0.61
cc_16 VNB N_A_M1039_g 0.0478711f $X=-0.19 $Y=-0.245 $X2=7.365 $Y2=0.61
cc_17 VNB N_A_c_172_n 0.588305f $X=-0.19 $Y=-0.245 $X2=10.75 $Y2=1.485
cc_18 VNB N_A_c_173_n 0.00387801f $X=-0.19 $Y=-0.245 $X2=1.13 $Y2=1.295
cc_19 VNB N_A_c_174_n 0.00654828f $X=-0.19 $Y=-0.245 $X2=2.03 $Y2=1.295
cc_20 VNB N_A_c_175_n 0.00577619f $X=-0.19 $Y=-0.245 $X2=3 $Y2=1.295
cc_21 VNB N_A_c_176_n 0.00517742f $X=-0.19 $Y=-0.245 $X2=3.93 $Y2=1.295
cc_22 VNB N_A_c_177_n 0.00561549f $X=-0.19 $Y=-0.245 $X2=4.92 $Y2=1.295
cc_23 VNB N_A_c_178_n 0.00306139f $X=-0.19 $Y=-0.245 $X2=5.76 $Y2=1.295
cc_24 VNB N_A_c_179_n 0.00330179f $X=-0.19 $Y=-0.245 $X2=6.71 $Y2=1.295
cc_25 VNB N_A_c_180_n 0.0785738f $X=-0.19 $Y=-0.245 $X2=7.83 $Y2=1.295
cc_26 VNB N_A_c_181_n 0.0290559f $X=-0.19 $Y=-0.245 $X2=10.71 $Y2=1.295
cc_27 VNB N_VPWR_c_573_n 0.48212f $X=-0.19 $Y=-0.245 $X2=9.665 $Y2=1.542
cc_28 VNB N_Y_c_806_n 0.00204288f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_Y_c_807_n 0.0068134f $X=-0.19 $Y=-0.245 $X2=5.645 $Y2=1.32
cc_30 VNB N_Y_c_808_n 0.00162022f $X=-0.19 $Y=-0.245 $X2=5.955 $Y2=1.765
cc_31 VNB N_Y_c_809_n 9.15856e-19 $X=-0.19 $Y=-0.245 $X2=5.955 $Y2=2.4
cc_32 VNB N_Y_c_810_n 0.00238225f $X=-0.19 $Y=-0.245 $X2=6.075 $Y2=0.61
cc_33 VNB N_Y_c_811_n 0.0100998f $X=-0.19 $Y=-0.245 $X2=6.505 $Y2=1.32
cc_34 VNB N_Y_c_812_n 0.00273892f $X=-0.19 $Y=-0.245 $X2=6.505 $Y2=0.61
cc_35 VNB N_Y_c_813_n 0.00252649f $X=-0.19 $Y=-0.245 $X2=6.905 $Y2=2.4
cc_36 VNB N_Y_c_814_n 0.00260578f $X=-0.19 $Y=-0.245 $X2=7.365 $Y2=1.32
cc_37 VNB N_Y_c_815_n 0.00364049f $X=-0.19 $Y=-0.245 $X2=7.865 $Y2=2.4
cc_38 VNB N_Y_c_816_n 0.00223955f $X=-0.19 $Y=-0.245 $X2=8.765 $Y2=2.4
cc_39 VNB N_Y_c_817_n 0.00345942f $X=-0.19 $Y=-0.245 $X2=9.215 $Y2=2.4
cc_40 VNB N_Y_c_818_n 0.00402748f $X=-0.19 $Y=-0.245 $X2=11.015 $Y2=2.4
cc_41 VNB N_Y_c_819_n 0.0129955f $X=-0.19 $Y=-0.245 $X2=3.645 $Y2=1.542
cc_42 VNB N_Y_c_820_n 0.00947359f $X=-0.19 $Y=-0.245 $X2=11.015 $Y2=1.542
cc_43 VNB N_Y_c_821_n 0.00406555f $X=-0.19 $Y=-0.245 $X2=1.135 $Y2=1.485
cc_44 VNB N_VGND_c_1131_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=2.4
cc_45 VNB N_VGND_c_1132_n 0.0399637f $X=-0.19 $Y=-0.245 $X2=2.285 $Y2=0.61
cc_46 VNB N_VGND_c_1133_n 0.00793748f $X=-0.19 $Y=-0.245 $X2=2.305 $Y2=2.4
cc_47 VNB N_VGND_c_1134_n 0.0130085f $X=-0.19 $Y=-0.245 $X2=2.715 $Y2=0.61
cc_48 VNB N_VGND_c_1135_n 0.0124212f $X=-0.19 $Y=-0.245 $X2=2.755 $Y2=2.4
cc_49 VNB N_VGND_c_1136_n 0.01271f $X=-0.19 $Y=-0.245 $X2=3.215 $Y2=1.32
cc_50 VNB N_VGND_c_1137_n 0.0124326f $X=-0.19 $Y=-0.245 $X2=3.645 $Y2=1.32
cc_51 VNB N_VGND_c_1138_n 0.00823433f $X=-0.19 $Y=-0.245 $X2=3.655 $Y2=1.765
cc_52 VNB N_VGND_c_1139_n 0.0061123f $X=-0.19 $Y=-0.245 $X2=4.105 $Y2=2.4
cc_53 VNB N_VGND_c_1140_n 0.0154173f $X=-0.19 $Y=-0.245 $X2=4.215 $Y2=0.61
cc_54 VNB N_VGND_c_1141_n 0.00548191f $X=-0.19 $Y=-0.245 $X2=4.215 $Y2=0.61
cc_55 VNB N_VGND_c_1142_n 0.0179248f $X=-0.19 $Y=-0.245 $X2=4.555 $Y2=1.765
cc_56 VNB N_VGND_c_1143_n 0.00538573f $X=-0.19 $Y=-0.245 $X2=4.555 $Y2=2.4
cc_57 VNB N_VGND_c_1144_n 0.0192699f $X=-0.19 $Y=-0.245 $X2=4.645 $Y2=1.32
cc_58 VNB N_VGND_c_1145_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=4.645 $Y2=0.61
cc_59 VNB N_VGND_c_1146_n 0.019099f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_1147_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=5.005 $Y2=1.765
cc_61 VNB N_VGND_c_1148_n 0.0193568f $X=-0.19 $Y=-0.245 $X2=5.005 $Y2=2.4
cc_62 VNB N_VGND_c_1149_n 0.00615512f $X=-0.19 $Y=-0.245 $X2=5.215 $Y2=1.32
cc_63 VNB N_VGND_c_1150_n 0.017363f $X=-0.19 $Y=-0.245 $X2=5.215 $Y2=0.61
cc_64 VNB N_VGND_c_1151_n 0.00548191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_1152_n 0.0165915f $X=-0.19 $Y=-0.245 $X2=5.455 $Y2=2.4
cc_66 VNB N_VGND_c_1153_n 0.00615512f $X=-0.19 $Y=-0.245 $X2=5.455 $Y2=2.4
cc_67 VNB N_VGND_c_1154_n 0.0474172f $X=-0.19 $Y=-0.245 $X2=5.645 $Y2=0.61
cc_68 VNB N_VGND_c_1155_n 0.03761f $X=-0.19 $Y=-0.245 $X2=5.955 $Y2=1.765
cc_69 VNB N_VGND_c_1156_n 0.0335227f $X=-0.19 $Y=-0.245 $X2=7.865 $Y2=2.4
cc_70 VNB N_VGND_c_1157_n 0.0560816f $X=-0.19 $Y=-0.245 $X2=9.215 $Y2=1.765
cc_71 VNB N_VGND_c_1158_n 0.679149f $X=-0.19 $Y=-0.245 $X2=9.215 $Y2=2.4
cc_72 VNB N_VGND_c_1159_n 0.0175452f $X=-0.19 $Y=-0.245 $X2=10.115 $Y2=2.4
cc_73 VPB N_A_c_182_n 0.0190846f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_74 VPB N_A_c_183_n 0.0149759f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.765
cc_75 VPB N_A_c_184_n 0.0152869f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=1.765
cc_76 VPB N_A_c_185_n 0.0155846f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=1.765
cc_77 VPB N_A_c_186_n 0.0152871f $X=-0.19 $Y=1.66 $X2=2.305 $Y2=1.765
cc_78 VPB N_A_c_187_n 0.0155841f $X=-0.19 $Y=1.66 $X2=2.755 $Y2=1.765
cc_79 VPB N_A_c_188_n 0.0156763f $X=-0.19 $Y=1.66 $X2=3.205 $Y2=1.765
cc_80 VPB N_A_c_189_n 0.0152871f $X=-0.19 $Y=1.66 $X2=3.655 $Y2=1.765
cc_81 VPB N_A_c_190_n 0.0155846f $X=-0.19 $Y=1.66 $X2=4.105 $Y2=1.765
cc_82 VPB N_A_c_191_n 0.0152848f $X=-0.19 $Y=1.66 $X2=4.555 $Y2=1.765
cc_83 VPB N_A_c_192_n 0.0155892f $X=-0.19 $Y=1.66 $X2=5.005 $Y2=1.765
cc_84 VPB N_A_c_193_n 0.0156611f $X=-0.19 $Y=1.66 $X2=5.455 $Y2=1.765
cc_85 VPB N_A_c_194_n 0.0158646f $X=-0.19 $Y=1.66 $X2=5.955 $Y2=1.765
cc_86 VPB N_A_c_195_n 0.0157363f $X=-0.19 $Y=1.66 $X2=6.405 $Y2=1.765
cc_87 VPB N_A_c_196_n 0.0165056f $X=-0.19 $Y=1.66 $X2=6.905 $Y2=1.765
cc_88 VPB N_A_c_197_n 0.0154383f $X=-0.19 $Y=1.66 $X2=7.415 $Y2=1.765
cc_89 VPB N_A_c_198_n 0.0149964f $X=-0.19 $Y=1.66 $X2=7.865 $Y2=1.765
cc_90 VPB N_A_c_199_n 0.0149989f $X=-0.19 $Y=1.66 $X2=8.315 $Y2=1.765
cc_91 VPB N_A_c_200_n 0.0156962f $X=-0.19 $Y=1.66 $X2=8.765 $Y2=1.765
cc_92 VPB N_A_c_201_n 0.0150021f $X=-0.19 $Y=1.66 $X2=9.215 $Y2=1.765
cc_93 VPB N_A_c_202_n 0.0149989f $X=-0.19 $Y=1.66 $X2=9.665 $Y2=1.765
cc_94 VPB N_A_c_203_n 0.0149989f $X=-0.19 $Y=1.66 $X2=10.115 $Y2=1.765
cc_95 VPB N_A_c_204_n 0.0149989f $X=-0.19 $Y=1.66 $X2=10.565 $Y2=1.765
cc_96 VPB N_A_c_205_n 0.0187055f $X=-0.19 $Y=1.66 $X2=11.015 $Y2=1.765
cc_97 VPB N_A_c_172_n 0.340562f $X=-0.19 $Y=1.66 $X2=10.75 $Y2=1.485
cc_98 VPB N_VPWR_c_574_n 0.0120106f $X=-0.19 $Y=1.66 $X2=2.755 $Y2=1.765
cc_99 VPB N_VPWR_c_575_n 0.0504452f $X=-0.19 $Y=1.66 $X2=2.755 $Y2=2.4
cc_100 VPB N_VPWR_c_576_n 0.00646409f $X=-0.19 $Y=1.66 $X2=3.215 $Y2=0.61
cc_101 VPB N_VPWR_c_577_n 0.00923549f $X=-0.19 $Y=1.66 $X2=3.655 $Y2=1.765
cc_102 VPB N_VPWR_c_578_n 0.00924893f $X=-0.19 $Y=1.66 $X2=4.215 $Y2=1.32
cc_103 VPB N_VPWR_c_579_n 0.00923549f $X=-0.19 $Y=1.66 $X2=4.555 $Y2=2.4
cc_104 VPB N_VPWR_c_580_n 0.00919269f $X=-0.19 $Y=1.66 $X2=5.005 $Y2=2.4
cc_105 VPB N_VPWR_c_581_n 0.00986066f $X=-0.19 $Y=1.66 $X2=5.455 $Y2=1.765
cc_106 VPB N_VPWR_c_582_n 0.0104904f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB N_VPWR_c_583_n 0.00489832f $X=-0.19 $Y=1.66 $X2=6.075 $Y2=0.61
cc_108 VPB N_VPWR_c_584_n 0.0164465f $X=-0.19 $Y=1.66 $X2=6.405 $Y2=2.4
cc_109 VPB N_VPWR_c_585_n 0.00579511f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_110 VPB N_VPWR_c_586_n 0.00435442f $X=-0.19 $Y=1.66 $X2=6.935 $Y2=0.61
cc_111 VPB N_VPWR_c_587_n 0.00425453f $X=-0.19 $Y=1.66 $X2=7.415 $Y2=1.765
cc_112 VPB N_VPWR_c_588_n 0.0120106f $X=-0.19 $Y=1.66 $X2=7.865 $Y2=2.4
cc_113 VPB N_VPWR_c_589_n 0.0651331f $X=-0.19 $Y=1.66 $X2=8.315 $Y2=1.765
cc_114 VPB N_VPWR_c_590_n 0.0162902f $X=-0.19 $Y=1.66 $X2=8.765 $Y2=2.4
cc_115 VPB N_VPWR_c_591_n 0.00460249f $X=-0.19 $Y=1.66 $X2=9.215 $Y2=1.765
cc_116 VPB N_VPWR_c_592_n 0.0206041f $X=-0.19 $Y=1.66 $X2=9.215 $Y2=2.4
cc_117 VPB N_VPWR_c_593_n 0.00324402f $X=-0.19 $Y=1.66 $X2=9.665 $Y2=1.765
cc_118 VPB N_VPWR_c_594_n 0.0206041f $X=-0.19 $Y=1.66 $X2=9.665 $Y2=2.4
cc_119 VPB N_VPWR_c_595_n 0.00324402f $X=-0.19 $Y=1.66 $X2=10.115 $Y2=1.765
cc_120 VPB N_VPWR_c_596_n 0.0211509f $X=-0.19 $Y=1.66 $X2=10.115 $Y2=2.4
cc_121 VPB N_VPWR_c_597_n 0.00324402f $X=-0.19 $Y=1.66 $X2=10.565 $Y2=1.765
cc_122 VPB N_VPWR_c_598_n 0.0206041f $X=-0.19 $Y=1.66 $X2=10.565 $Y2=2.4
cc_123 VPB N_VPWR_c_599_n 0.00324402f $X=-0.19 $Y=1.66 $X2=11.015 $Y2=1.765
cc_124 VPB N_VPWR_c_600_n 0.0206041f $X=-0.19 $Y=1.66 $X2=11.015 $Y2=2.4
cc_125 VPB N_VPWR_c_601_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0.985 $Y2=1.18
cc_126 VPB N_VPWR_c_602_n 0.0186401f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.542
cc_127 VPB N_VPWR_c_603_n 0.00545601f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.542
cc_128 VPB N_VPWR_c_604_n 0.019519f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.542
cc_129 VPB N_VPWR_c_605_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.542
cc_130 VPB N_VPWR_c_606_n 0.0191503f $X=-0.19 $Y=1.66 $X2=4.645 $Y2=1.542
cc_131 VPB N_VPWR_c_607_n 0.0164465f $X=-0.19 $Y=1.66 $X2=5.215 $Y2=1.542
cc_132 VPB N_VPWR_c_608_n 0.0164465f $X=-0.19 $Y=1.66 $X2=5.76 $Y2=1.485
cc_133 VPB N_VPWR_c_609_n 0.00460249f $X=-0.19 $Y=1.66 $X2=6.935 $Y2=1.542
cc_134 VPB N_VPWR_c_610_n 0.00601644f $X=-0.19 $Y=1.66 $X2=7.69 $Y2=1.542
cc_135 VPB N_VPWR_c_611_n 0.00601644f $X=-0.19 $Y=1.66 $X2=7.865 $Y2=1.542
cc_136 VPB N_VPWR_c_573_n 0.132762f $X=-0.19 $Y=1.66 $X2=9.665 $Y2=1.542
cc_137 VPB N_Y_c_822_n 0.00257348f $X=-0.19 $Y=1.66 $X2=5.005 $Y2=1.765
cc_138 VPB N_Y_c_823_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_Y_c_807_n 0.00135194f $X=-0.19 $Y=1.66 $X2=5.645 $Y2=1.32
cc_140 VPB N_Y_c_809_n 0.00150393f $X=-0.19 $Y=1.66 $X2=5.955 $Y2=2.4
cc_141 VPB N_Y_c_826_n 3.97087e-19 $X=-0.19 $Y=1.66 $X2=6.405 $Y2=2.4
cc_142 VPB N_Y_c_811_n 0.0024558f $X=-0.19 $Y=1.66 $X2=6.505 $Y2=1.32
cc_143 VPB N_Y_c_815_n 0.00150097f $X=-0.19 $Y=1.66 $X2=7.865 $Y2=2.4
cc_144 VPB N_Y_c_829_n 0.00198541f $X=-0.19 $Y=1.66 $X2=10.115 $Y2=1.765
cc_145 VPB N_Y_c_818_n 0.00360064f $X=-0.19 $Y=1.66 $X2=11.015 $Y2=2.4
cc_146 VPB N_Y_c_831_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.542
cc_147 VPB N_Y_c_832_n 0.00257348f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=1.542
cc_148 VPB N_Y_c_833_n 0.00276337f $X=-0.19 $Y=1.66 $X2=2.715 $Y2=1.542
cc_149 VPB N_Y_c_819_n 0.00541142f $X=-0.19 $Y=1.66 $X2=3.645 $Y2=1.542
cc_150 VPB N_Y_c_835_n 0.00303384f $X=-0.19 $Y=1.66 $X2=4.92 $Y2=1.485
cc_151 VPB N_Y_c_836_n 0.00306331f $X=-0.19 $Y=1.66 $X2=5.76 $Y2=1.485
cc_152 VPB N_Y_c_837_n 0.00303384f $X=-0.19 $Y=1.66 $X2=6.905 $Y2=1.542
cc_153 VPB N_Y_c_838_n 0.00303384f $X=-0.19 $Y=1.66 $X2=8.315 $Y2=1.542
cc_154 VPB N_Y_c_820_n 0.00135161f $X=-0.19 $Y=1.66 $X2=11.015 $Y2=1.542
cc_155 VPB N_Y_c_821_n 0.00131968f $X=-0.19 $Y=1.66 $X2=1.135 $Y2=1.485
cc_156 N_A_c_182_n N_VPWR_c_575_n 0.0168926f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_157 N_A_c_183_n N_VPWR_c_575_n 6.23847e-19 $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_158 N_A_c_182_n N_VPWR_c_576_n 7.68816e-19 $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_159 N_A_c_183_n N_VPWR_c_576_n 0.01532f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_160 N_A_c_184_n N_VPWR_c_576_n 0.00703885f $X=1.405 $Y=1.765 $X2=0 $Y2=0
cc_161 N_A_c_172_n N_VPWR_c_576_n 0.00628163f $X=10.75 $Y=1.485 $X2=0 $Y2=0
cc_162 N_A_c_173_n N_VPWR_c_576_n 0.019006f $X=1.13 $Y=1.295 $X2=0 $Y2=0
cc_163 N_A_c_181_n N_VPWR_c_576_n 7.83582e-19 $X=10.71 $Y=1.295 $X2=0 $Y2=0
cc_164 N_A_c_185_n N_VPWR_c_577_n 0.00663139f $X=1.855 $Y=1.765 $X2=0 $Y2=0
cc_165 N_A_c_186_n N_VPWR_c_577_n 0.00654256f $X=2.305 $Y=1.765 $X2=0 $Y2=0
cc_166 N_A_c_172_n N_VPWR_c_577_n 0.00428618f $X=10.75 $Y=1.485 $X2=0 $Y2=0
cc_167 N_A_c_174_n N_VPWR_c_577_n 0.0129137f $X=2.03 $Y=1.295 $X2=0 $Y2=0
cc_168 N_A_c_181_n N_VPWR_c_577_n 5.34739e-19 $X=10.71 $Y=1.295 $X2=0 $Y2=0
cc_169 N_A_c_187_n N_VPWR_c_578_n 0.00657003f $X=2.755 $Y=1.765 $X2=0 $Y2=0
cc_170 N_A_c_188_n N_VPWR_c_578_n 0.00763212f $X=3.205 $Y=1.765 $X2=0 $Y2=0
cc_171 N_A_c_172_n N_VPWR_c_578_n 0.00417652f $X=10.75 $Y=1.485 $X2=0 $Y2=0
cc_172 N_A_c_175_n N_VPWR_c_578_n 0.0129137f $X=3 $Y=1.295 $X2=0 $Y2=0
cc_173 N_A_c_181_n N_VPWR_c_578_n 5.34739e-19 $X=10.71 $Y=1.295 $X2=0 $Y2=0
cc_174 N_A_c_189_n N_VPWR_c_579_n 0.00654256f $X=3.655 $Y=1.765 $X2=0 $Y2=0
cc_175 N_A_c_190_n N_VPWR_c_579_n 0.00658356f $X=4.105 $Y=1.765 $X2=0 $Y2=0
cc_176 N_A_c_172_n N_VPWR_c_579_n 0.00417652f $X=10.75 $Y=1.485 $X2=0 $Y2=0
cc_177 N_A_c_176_n N_VPWR_c_579_n 0.0129137f $X=3.93 $Y=1.295 $X2=0 $Y2=0
cc_178 N_A_c_181_n N_VPWR_c_579_n 5.34739e-19 $X=10.71 $Y=1.295 $X2=0 $Y2=0
cc_179 N_A_c_191_n N_VPWR_c_580_n 0.00650785f $X=4.555 $Y=1.765 $X2=0 $Y2=0
cc_180 N_A_c_192_n N_VPWR_c_580_n 0.00661751f $X=5.005 $Y=1.765 $X2=0 $Y2=0
cc_181 N_A_c_172_n N_VPWR_c_580_n 0.00584842f $X=10.75 $Y=1.485 $X2=0 $Y2=0
cc_182 N_A_c_177_n N_VPWR_c_580_n 0.00830167f $X=4.92 $Y=1.295 $X2=0 $Y2=0
cc_183 N_A_c_181_n N_VPWR_c_580_n 0.00205008f $X=10.71 $Y=1.295 $X2=0 $Y2=0
cc_184 N_A_c_193_n N_VPWR_c_581_n 0.00708127f $X=5.455 $Y=1.765 $X2=0 $Y2=0
cc_185 N_A_c_194_n N_VPWR_c_581_n 0.00810561f $X=5.955 $Y=1.765 $X2=0 $Y2=0
cc_186 N_A_c_172_n N_VPWR_c_581_n 0.006872f $X=10.75 $Y=1.485 $X2=0 $Y2=0
cc_187 N_A_c_178_n N_VPWR_c_581_n 0.0190631f $X=5.76 $Y=1.295 $X2=0 $Y2=0
cc_188 N_A_c_181_n N_VPWR_c_581_n 7.89376e-19 $X=10.71 $Y=1.295 $X2=0 $Y2=0
cc_189 N_A_c_195_n N_VPWR_c_582_n 0.00266116f $X=6.405 $Y=1.765 $X2=0 $Y2=0
cc_190 N_A_c_196_n N_VPWR_c_582_n 0.00967509f $X=6.905 $Y=1.765 $X2=0 $Y2=0
cc_191 N_A_c_172_n N_VPWR_c_582_n 0.0083802f $X=10.75 $Y=1.485 $X2=0 $Y2=0
cc_192 N_A_c_179_n N_VPWR_c_582_n 0.0190631f $X=6.71 $Y=1.295 $X2=0 $Y2=0
cc_193 N_A_c_181_n N_VPWR_c_582_n 0.00178473f $X=10.71 $Y=1.295 $X2=0 $Y2=0
cc_194 N_A_c_196_n N_VPWR_c_583_n 8.74621e-19 $X=6.905 $Y=1.765 $X2=0 $Y2=0
cc_195 N_A_c_197_n N_VPWR_c_583_n 0.015894f $X=7.415 $Y=1.765 $X2=0 $Y2=0
cc_196 N_A_c_198_n N_VPWR_c_583_n 0.0159037f $X=7.865 $Y=1.765 $X2=0 $Y2=0
cc_197 N_A_c_199_n N_VPWR_c_583_n 7.70516e-19 $X=8.315 $Y=1.765 $X2=0 $Y2=0
cc_198 N_A_c_172_n N_VPWR_c_583_n 0.00829349f $X=10.75 $Y=1.485 $X2=0 $Y2=0
cc_199 N_A_c_180_n N_VPWR_c_583_n 0.021312f $X=7.83 $Y=1.295 $X2=0 $Y2=0
cc_200 N_A_c_181_n N_VPWR_c_583_n 0.00224459f $X=10.71 $Y=1.295 $X2=0 $Y2=0
cc_201 N_A_c_198_n N_VPWR_c_584_n 0.00413917f $X=7.865 $Y=1.765 $X2=0 $Y2=0
cc_202 N_A_c_199_n N_VPWR_c_584_n 0.00413917f $X=8.315 $Y=1.765 $X2=0 $Y2=0
cc_203 N_A_c_198_n N_VPWR_c_585_n 7.68816e-19 $X=7.865 $Y=1.765 $X2=0 $Y2=0
cc_204 N_A_c_199_n N_VPWR_c_585_n 0.01532f $X=8.315 $Y=1.765 $X2=0 $Y2=0
cc_205 N_A_c_200_n N_VPWR_c_585_n 0.00707592f $X=8.765 $Y=1.765 $X2=0 $Y2=0
cc_206 N_A_c_172_n N_VPWR_c_585_n 0.0058039f $X=10.75 $Y=1.485 $X2=0 $Y2=0
cc_207 N_A_c_180_n N_VPWR_c_585_n 0.019006f $X=7.83 $Y=1.295 $X2=0 $Y2=0
cc_208 N_A_c_181_n N_VPWR_c_585_n 7.83582e-19 $X=10.71 $Y=1.295 $X2=0 $Y2=0
cc_209 N_A_c_200_n N_VPWR_c_586_n 7.80707e-19 $X=8.765 $Y=1.765 $X2=0 $Y2=0
cc_210 N_A_c_201_n N_VPWR_c_586_n 0.0160348f $X=9.215 $Y=1.765 $X2=0 $Y2=0
cc_211 N_A_c_202_n N_VPWR_c_586_n 0.0159037f $X=9.665 $Y=1.765 $X2=0 $Y2=0
cc_212 N_A_c_203_n N_VPWR_c_586_n 7.70516e-19 $X=10.115 $Y=1.765 $X2=0 $Y2=0
cc_213 N_A_c_172_n N_VPWR_c_586_n 0.00748245f $X=10.75 $Y=1.485 $X2=0 $Y2=0
cc_214 N_A_c_180_n N_VPWR_c_586_n 0.0250982f $X=7.83 $Y=1.295 $X2=0 $Y2=0
cc_215 N_A_c_181_n N_VPWR_c_586_n 0.00103243f $X=10.71 $Y=1.295 $X2=0 $Y2=0
cc_216 N_A_c_202_n N_VPWR_c_587_n 7.70516e-19 $X=9.665 $Y=1.765 $X2=0 $Y2=0
cc_217 N_A_c_203_n N_VPWR_c_587_n 0.0159037f $X=10.115 $Y=1.765 $X2=0 $Y2=0
cc_218 N_A_c_204_n N_VPWR_c_587_n 0.0159037f $X=10.565 $Y=1.765 $X2=0 $Y2=0
cc_219 N_A_c_205_n N_VPWR_c_587_n 7.70516e-19 $X=11.015 $Y=1.765 $X2=0 $Y2=0
cc_220 N_A_c_172_n N_VPWR_c_587_n 0.00748245f $X=10.75 $Y=1.485 $X2=0 $Y2=0
cc_221 N_A_c_180_n N_VPWR_c_587_n 0.0250982f $X=7.83 $Y=1.295 $X2=0 $Y2=0
cc_222 N_A_c_181_n N_VPWR_c_587_n 0.00103243f $X=10.71 $Y=1.295 $X2=0 $Y2=0
cc_223 N_A_c_204_n N_VPWR_c_589_n 6.78853e-19 $X=10.565 $Y=1.765 $X2=0 $Y2=0
cc_224 N_A_c_205_n N_VPWR_c_589_n 0.0185947f $X=11.015 $Y=1.765 $X2=0 $Y2=0
cc_225 N_A_c_172_n N_VPWR_c_589_n 7.80018e-19 $X=10.75 $Y=1.485 $X2=0 $Y2=0
cc_226 N_A_c_182_n N_VPWR_c_590_n 0.00413917f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_227 N_A_c_183_n N_VPWR_c_590_n 0.00413917f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_228 N_A_c_184_n N_VPWR_c_592_n 0.00445602f $X=1.405 $Y=1.765 $X2=0 $Y2=0
cc_229 N_A_c_185_n N_VPWR_c_592_n 0.00445602f $X=1.855 $Y=1.765 $X2=0 $Y2=0
cc_230 N_A_c_186_n N_VPWR_c_594_n 0.00445602f $X=2.305 $Y=1.765 $X2=0 $Y2=0
cc_231 N_A_c_187_n N_VPWR_c_594_n 0.00445602f $X=2.755 $Y=1.765 $X2=0 $Y2=0
cc_232 N_A_c_188_n N_VPWR_c_596_n 0.00461464f $X=3.205 $Y=1.765 $X2=0 $Y2=0
cc_233 N_A_c_189_n N_VPWR_c_596_n 0.00445602f $X=3.655 $Y=1.765 $X2=0 $Y2=0
cc_234 N_A_c_190_n N_VPWR_c_598_n 0.00445602f $X=4.105 $Y=1.765 $X2=0 $Y2=0
cc_235 N_A_c_191_n N_VPWR_c_598_n 0.00445602f $X=4.555 $Y=1.765 $X2=0 $Y2=0
cc_236 N_A_c_192_n N_VPWR_c_600_n 0.00445602f $X=5.005 $Y=1.765 $X2=0 $Y2=0
cc_237 N_A_c_193_n N_VPWR_c_600_n 0.00445602f $X=5.455 $Y=1.765 $X2=0 $Y2=0
cc_238 N_A_c_194_n N_VPWR_c_602_n 0.00445602f $X=5.955 $Y=1.765 $X2=0 $Y2=0
cc_239 N_A_c_195_n N_VPWR_c_602_n 0.00461464f $X=6.405 $Y=1.765 $X2=0 $Y2=0
cc_240 N_A_c_196_n N_VPWR_c_604_n 0.00461464f $X=6.905 $Y=1.765 $X2=0 $Y2=0
cc_241 N_A_c_197_n N_VPWR_c_604_n 0.00413917f $X=7.415 $Y=1.765 $X2=0 $Y2=0
cc_242 N_A_c_200_n N_VPWR_c_606_n 0.00461464f $X=8.765 $Y=1.765 $X2=0 $Y2=0
cc_243 N_A_c_201_n N_VPWR_c_606_n 0.00413917f $X=9.215 $Y=1.765 $X2=0 $Y2=0
cc_244 N_A_c_202_n N_VPWR_c_607_n 0.00413917f $X=9.665 $Y=1.765 $X2=0 $Y2=0
cc_245 N_A_c_203_n N_VPWR_c_607_n 0.00413917f $X=10.115 $Y=1.765 $X2=0 $Y2=0
cc_246 N_A_c_204_n N_VPWR_c_608_n 0.00413917f $X=10.565 $Y=1.765 $X2=0 $Y2=0
cc_247 N_A_c_205_n N_VPWR_c_608_n 0.00413917f $X=11.015 $Y=1.765 $X2=0 $Y2=0
cc_248 N_A_c_182_n N_VPWR_c_573_n 0.00817726f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_249 N_A_c_183_n N_VPWR_c_573_n 0.00817726f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_250 N_A_c_184_n N_VPWR_c_573_n 0.00857589f $X=1.405 $Y=1.765 $X2=0 $Y2=0
cc_251 N_A_c_185_n N_VPWR_c_573_n 0.00857589f $X=1.855 $Y=1.765 $X2=0 $Y2=0
cc_252 N_A_c_186_n N_VPWR_c_573_n 0.00857589f $X=2.305 $Y=1.765 $X2=0 $Y2=0
cc_253 N_A_c_187_n N_VPWR_c_573_n 0.00857589f $X=2.755 $Y=1.765 $X2=0 $Y2=0
cc_254 N_A_c_188_n N_VPWR_c_573_n 0.00908951f $X=3.205 $Y=1.765 $X2=0 $Y2=0
cc_255 N_A_c_189_n N_VPWR_c_573_n 0.00857589f $X=3.655 $Y=1.765 $X2=0 $Y2=0
cc_256 N_A_c_190_n N_VPWR_c_573_n 0.00857589f $X=4.105 $Y=1.765 $X2=0 $Y2=0
cc_257 N_A_c_191_n N_VPWR_c_573_n 0.00857589f $X=4.555 $Y=1.765 $X2=0 $Y2=0
cc_258 N_A_c_192_n N_VPWR_c_573_n 0.00857589f $X=5.005 $Y=1.765 $X2=0 $Y2=0
cc_259 N_A_c_193_n N_VPWR_c_573_n 0.0085805f $X=5.455 $Y=1.765 $X2=0 $Y2=0
cc_260 N_A_c_194_n N_VPWR_c_573_n 0.00857378f $X=5.955 $Y=1.765 $X2=0 $Y2=0
cc_261 N_A_c_195_n N_VPWR_c_573_n 0.00908628f $X=6.405 $Y=1.765 $X2=0 $Y2=0
cc_262 N_A_c_196_n N_VPWR_c_573_n 0.00909288f $X=6.905 $Y=1.765 $X2=0 $Y2=0
cc_263 N_A_c_197_n N_VPWR_c_573_n 0.00818274f $X=7.415 $Y=1.765 $X2=0 $Y2=0
cc_264 N_A_c_198_n N_VPWR_c_573_n 0.00817726f $X=7.865 $Y=1.765 $X2=0 $Y2=0
cc_265 N_A_c_199_n N_VPWR_c_573_n 0.00817726f $X=8.315 $Y=1.765 $X2=0 $Y2=0
cc_266 N_A_c_200_n N_VPWR_c_573_n 0.00908951f $X=8.765 $Y=1.765 $X2=0 $Y2=0
cc_267 N_A_c_201_n N_VPWR_c_573_n 0.00817726f $X=9.215 $Y=1.765 $X2=0 $Y2=0
cc_268 N_A_c_202_n N_VPWR_c_573_n 0.00817726f $X=9.665 $Y=1.765 $X2=0 $Y2=0
cc_269 N_A_c_203_n N_VPWR_c_573_n 0.00817726f $X=10.115 $Y=1.765 $X2=0 $Y2=0
cc_270 N_A_c_204_n N_VPWR_c_573_n 0.00817726f $X=10.565 $Y=1.765 $X2=0 $Y2=0
cc_271 N_A_c_205_n N_VPWR_c_573_n 0.00817726f $X=11.015 $Y=1.765 $X2=0 $Y2=0
cc_272 N_A_M1002_g N_Y_c_806_n 2.05722e-19 $X=0.495 $Y=0.61 $X2=0 $Y2=0
cc_273 N_A_M1003_g N_Y_c_806_n 0.00575088f $X=0.925 $Y=0.61 $X2=0 $Y2=0
cc_274 N_A_c_184_n N_Y_c_822_n 0.0101078f $X=1.405 $Y=1.765 $X2=0 $Y2=0
cc_275 N_A_c_185_n N_Y_c_822_n 0.0101078f $X=1.855 $Y=1.765 $X2=0 $Y2=0
cc_276 N_A_c_186_n N_Y_c_823_n 0.0101078f $X=2.305 $Y=1.765 $X2=0 $Y2=0
cc_277 N_A_c_187_n N_Y_c_823_n 0.0101078f $X=2.755 $Y=1.765 $X2=0 $Y2=0
cc_278 N_A_M1017_g N_Y_c_807_n 0.00113286f $X=3.645 $Y=0.61 $X2=0 $Y2=0
cc_279 N_A_c_190_n N_Y_c_807_n 9.55363e-19 $X=4.105 $Y=1.765 $X2=0 $Y2=0
cc_280 N_A_M1021_g N_Y_c_807_n 0.0177058f $X=4.215 $Y=0.61 $X2=0 $Y2=0
cc_281 N_A_c_191_n N_Y_c_807_n 0.00207923f $X=4.555 $Y=1.765 $X2=0 $Y2=0
cc_282 N_A_M1022_g N_Y_c_807_n 0.00983021f $X=4.645 $Y=0.61 $X2=0 $Y2=0
cc_283 N_A_c_192_n N_Y_c_807_n 2.94132e-19 $X=5.005 $Y=1.765 $X2=0 $Y2=0
cc_284 N_A_c_172_n N_Y_c_807_n 0.0317354f $X=10.75 $Y=1.485 $X2=0 $Y2=0
cc_285 N_A_c_176_n N_Y_c_807_n 0.035492f $X=3.93 $Y=1.295 $X2=0 $Y2=0
cc_286 N_A_c_177_n N_Y_c_807_n 0.0275344f $X=4.92 $Y=1.295 $X2=0 $Y2=0
cc_287 N_A_c_181_n N_Y_c_807_n 0.0332159f $X=10.71 $Y=1.295 $X2=0 $Y2=0
cc_288 N_A_M1029_g N_Y_c_808_n 4.62803e-19 $X=5.645 $Y=0.61 $X2=0 $Y2=0
cc_289 N_A_M1030_g N_Y_c_808_n 0.00646016f $X=6.075 $Y=0.61 $X2=0 $Y2=0
cc_290 N_A_c_194_n N_Y_c_809_n 0.00266055f $X=5.955 $Y=1.765 $X2=0 $Y2=0
cc_291 N_A_M1030_g N_Y_c_809_n 0.0035086f $X=6.075 $Y=0.61 $X2=0 $Y2=0
cc_292 N_A_c_195_n N_Y_c_809_n 0.00166693f $X=6.405 $Y=1.765 $X2=0 $Y2=0
cc_293 N_A_c_196_n N_Y_c_809_n 2.50506e-19 $X=6.905 $Y=1.765 $X2=0 $Y2=0
cc_294 N_A_c_172_n N_Y_c_809_n 0.0346951f $X=10.75 $Y=1.485 $X2=0 $Y2=0
cc_295 N_A_c_178_n N_Y_c_809_n 0.0353686f $X=5.76 $Y=1.295 $X2=0 $Y2=0
cc_296 N_A_c_179_n N_Y_c_809_n 0.0297797f $X=6.71 $Y=1.295 $X2=0 $Y2=0
cc_297 N_A_c_181_n N_Y_c_809_n 0.0329404f $X=10.71 $Y=1.295 $X2=0 $Y2=0
cc_298 N_A_M1030_g N_Y_c_810_n 0.00477496f $X=6.075 $Y=0.61 $X2=0 $Y2=0
cc_299 N_A_M1034_g N_Y_c_810_n 2.07919e-19 $X=6.505 $Y=0.61 $X2=0 $Y2=0
cc_300 N_A_c_183_n N_Y_c_826_n 0.00402199f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_301 N_A_c_172_n N_Y_c_826_n 4.49855e-19 $X=10.75 $Y=1.485 $X2=0 $Y2=0
cc_302 N_A_M1002_g N_Y_c_811_n 0.0117801f $X=0.495 $Y=0.61 $X2=0 $Y2=0
cc_303 N_A_c_182_n N_Y_c_811_n 0.00248883f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_304 N_A_c_183_n N_Y_c_811_n 6.91217e-19 $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_305 N_A_c_172_n N_Y_c_811_n 0.0356393f $X=10.75 $Y=1.485 $X2=0 $Y2=0
cc_306 N_A_c_173_n N_Y_c_811_n 0.0348136f $X=1.13 $Y=1.295 $X2=0 $Y2=0
cc_307 N_A_c_181_n N_Y_c_811_n 0.00159972f $X=10.71 $Y=1.295 $X2=0 $Y2=0
cc_308 N_A_M1004_g N_Y_c_812_n 2.29421e-19 $X=1.355 $Y=0.61 $X2=0 $Y2=0
cc_309 N_A_M1008_g N_Y_c_812_n 2.3112e-19 $X=1.785 $Y=0.61 $X2=0 $Y2=0
cc_310 N_A_c_181_n N_Y_c_812_n 9.91373e-19 $X=10.71 $Y=1.295 $X2=0 $Y2=0
cc_311 N_A_M1011_g N_Y_c_813_n 0.00446178f $X=2.285 $Y=0.61 $X2=0 $Y2=0
cc_312 N_A_M1012_g N_Y_c_813_n 0.00480415f $X=2.715 $Y=0.61 $X2=0 $Y2=0
cc_313 N_A_M1016_g N_Y_c_813_n 0.00108834f $X=3.215 $Y=0.61 $X2=0 $Y2=0
cc_314 N_A_c_181_n N_Y_c_813_n 4.71012e-19 $X=10.71 $Y=1.295 $X2=0 $Y2=0
cc_315 N_A_M1016_g N_Y_c_814_n 2.40073e-19 $X=3.215 $Y=0.61 $X2=0 $Y2=0
cc_316 N_A_M1017_g N_Y_c_814_n 0.00467704f $X=3.645 $Y=0.61 $X2=0 $Y2=0
cc_317 N_A_M1021_g N_Y_c_814_n 0.00113241f $X=4.215 $Y=0.61 $X2=0 $Y2=0
cc_318 N_A_c_181_n N_Y_c_814_n 0.00140445f $X=10.71 $Y=1.295 $X2=0 $Y2=0
cc_319 N_A_c_190_n N_Y_c_888_n 8.25115e-19 $X=4.105 $Y=1.765 $X2=0 $Y2=0
cc_320 N_A_c_191_n N_Y_c_888_n 0.00106087f $X=4.555 $Y=1.765 $X2=0 $Y2=0
cc_321 N_A_c_172_n N_Y_c_888_n 0.00237089f $X=10.75 $Y=1.485 $X2=0 $Y2=0
cc_322 N_A_c_181_n N_Y_c_888_n 0.00262869f $X=10.71 $Y=1.295 $X2=0 $Y2=0
cc_323 N_A_c_192_n N_Y_c_892_n 0.00151945f $X=5.005 $Y=1.765 $X2=0 $Y2=0
cc_324 N_A_c_193_n N_Y_c_892_n 0.00223127f $X=5.455 $Y=1.765 $X2=0 $Y2=0
cc_325 N_A_c_172_n N_Y_c_892_n 0.00672558f $X=10.75 $Y=1.485 $X2=0 $Y2=0
cc_326 N_A_c_177_n N_Y_c_892_n 9.35725e-19 $X=4.92 $Y=1.295 $X2=0 $Y2=0
cc_327 N_A_c_181_n N_Y_c_892_n 0.00476102f $X=10.71 $Y=1.295 $X2=0 $Y2=0
cc_328 N_A_M1022_g N_Y_c_815_n 0.00153159f $X=4.645 $Y=0.61 $X2=0 $Y2=0
cc_329 N_A_c_192_n N_Y_c_815_n 0.00134094f $X=5.005 $Y=1.765 $X2=0 $Y2=0
cc_330 N_A_M1026_g N_Y_c_815_n 0.0120682f $X=5.215 $Y=0.61 $X2=0 $Y2=0
cc_331 N_A_c_193_n N_Y_c_815_n 0.0020199f $X=5.455 $Y=1.765 $X2=0 $Y2=0
cc_332 N_A_M1029_g N_Y_c_815_n 0.00633798f $X=5.645 $Y=0.61 $X2=0 $Y2=0
cc_333 N_A_c_194_n N_Y_c_815_n 2.53518e-19 $X=5.955 $Y=1.765 $X2=0 $Y2=0
cc_334 N_A_c_172_n N_Y_c_815_n 0.0244673f $X=10.75 $Y=1.485 $X2=0 $Y2=0
cc_335 N_A_c_177_n N_Y_c_815_n 0.034848f $X=4.92 $Y=1.295 $X2=0 $Y2=0
cc_336 N_A_c_178_n N_Y_c_815_n 0.0347592f $X=5.76 $Y=1.295 $X2=0 $Y2=0
cc_337 N_A_c_181_n N_Y_c_815_n 0.016141f $X=10.71 $Y=1.295 $X2=0 $Y2=0
cc_338 N_A_M1026_g N_Y_c_816_n 0.00513212f $X=5.215 $Y=0.61 $X2=0 $Y2=0
cc_339 N_A_M1029_g N_Y_c_816_n 2.03144e-19 $X=5.645 $Y=0.61 $X2=0 $Y2=0
cc_340 N_A_c_172_n N_Y_c_816_n 0.00136026f $X=10.75 $Y=1.485 $X2=0 $Y2=0
cc_341 N_A_c_181_n N_Y_c_816_n 0.00460277f $X=10.71 $Y=1.295 $X2=0 $Y2=0
cc_342 N_A_M1034_g N_Y_c_817_n 0.00867347f $X=6.505 $Y=0.61 $X2=0 $Y2=0
cc_343 N_A_c_181_n N_Y_c_912_n 0.00183934f $X=10.71 $Y=1.295 $X2=0 $Y2=0
cc_344 N_A_c_188_n N_Y_c_818_n 0.00178902f $X=3.205 $Y=1.765 $X2=0 $Y2=0
cc_345 N_A_M1016_g N_Y_c_818_n 0.00573532f $X=3.215 $Y=0.61 $X2=0 $Y2=0
cc_346 N_A_M1017_g N_Y_c_818_n 0.0130408f $X=3.645 $Y=0.61 $X2=0 $Y2=0
cc_347 N_A_c_189_n N_Y_c_818_n 0.0135702f $X=3.655 $Y=1.765 $X2=0 $Y2=0
cc_348 N_A_c_190_n N_Y_c_818_n 6.08154e-19 $X=4.105 $Y=1.765 $X2=0 $Y2=0
cc_349 N_A_c_172_n N_Y_c_818_n 0.0310549f $X=10.75 $Y=1.485 $X2=0 $Y2=0
cc_350 N_A_c_175_n N_Y_c_818_n 0.0354598f $X=3 $Y=1.295 $X2=0 $Y2=0
cc_351 N_A_c_176_n N_Y_c_818_n 0.035492f $X=3.93 $Y=1.295 $X2=0 $Y2=0
cc_352 N_A_c_181_n N_Y_c_818_n 0.0325837f $X=10.71 $Y=1.295 $X2=0 $Y2=0
cc_353 N_A_c_190_n N_Y_c_831_n 0.0111833f $X=4.105 $Y=1.765 $X2=0 $Y2=0
cc_354 N_A_c_191_n N_Y_c_831_n 0.0111833f $X=4.555 $Y=1.765 $X2=0 $Y2=0
cc_355 N_A_c_192_n N_Y_c_832_n 0.0103773f $X=5.005 $Y=1.765 $X2=0 $Y2=0
cc_356 N_A_c_193_n N_Y_c_832_n 0.0104526f $X=5.455 $Y=1.765 $X2=0 $Y2=0
cc_357 N_A_c_194_n N_Y_c_833_n 0.00988118f $X=5.955 $Y=1.765 $X2=0 $Y2=0
cc_358 N_A_c_195_n N_Y_c_833_n 4.18282e-19 $X=6.405 $Y=1.765 $X2=0 $Y2=0
cc_359 N_A_c_196_n N_Y_c_819_n 0.00658218f $X=6.905 $Y=1.765 $X2=0 $Y2=0
cc_360 N_A_M1036_g N_Y_c_819_n 0.00968751f $X=6.935 $Y=0.61 $X2=0 $Y2=0
cc_361 N_A_M1039_g N_Y_c_819_n 0.0107483f $X=7.365 $Y=0.61 $X2=0 $Y2=0
cc_362 N_A_c_197_n N_Y_c_819_n 0.00238034f $X=7.415 $Y=1.765 $X2=0 $Y2=0
cc_363 N_A_c_172_n N_Y_c_819_n 0.0330156f $X=10.75 $Y=1.485 $X2=0 $Y2=0
cc_364 N_A_c_179_n N_Y_c_819_n 0.0353594f $X=6.71 $Y=1.295 $X2=0 $Y2=0
cc_365 N_A_c_180_n N_Y_c_819_n 0.0279635f $X=7.83 $Y=1.295 $X2=0 $Y2=0
cc_366 N_A_c_181_n N_Y_c_819_n 0.0317748f $X=10.71 $Y=1.295 $X2=0 $Y2=0
cc_367 N_A_c_198_n N_Y_c_835_n 0.00394046f $X=7.865 $Y=1.765 $X2=0 $Y2=0
cc_368 N_A_c_199_n N_Y_c_835_n 0.00394046f $X=8.315 $Y=1.765 $X2=0 $Y2=0
cc_369 N_A_c_172_n N_Y_c_835_n 0.00412535f $X=10.75 $Y=1.485 $X2=0 $Y2=0
cc_370 N_A_c_180_n N_Y_c_835_n 0.0129137f $X=7.83 $Y=1.295 $X2=0 $Y2=0
cc_371 N_A_c_181_n N_Y_c_835_n 5.34739e-19 $X=10.71 $Y=1.295 $X2=0 $Y2=0
cc_372 N_A_c_200_n N_Y_c_836_n 0.00518028f $X=8.765 $Y=1.765 $X2=0 $Y2=0
cc_373 N_A_c_201_n N_Y_c_836_n 0.00394046f $X=9.215 $Y=1.765 $X2=0 $Y2=0
cc_374 N_A_c_172_n N_Y_c_836_n 0.00412535f $X=10.75 $Y=1.485 $X2=0 $Y2=0
cc_375 N_A_c_180_n N_Y_c_836_n 0.0129137f $X=7.83 $Y=1.295 $X2=0 $Y2=0
cc_376 N_A_c_181_n N_Y_c_836_n 5.34739e-19 $X=10.71 $Y=1.295 $X2=0 $Y2=0
cc_377 N_A_c_202_n N_Y_c_837_n 0.00394046f $X=9.665 $Y=1.765 $X2=0 $Y2=0
cc_378 N_A_c_203_n N_Y_c_837_n 0.00394046f $X=10.115 $Y=1.765 $X2=0 $Y2=0
cc_379 N_A_c_172_n N_Y_c_837_n 0.00412535f $X=10.75 $Y=1.485 $X2=0 $Y2=0
cc_380 N_A_c_180_n N_Y_c_837_n 0.0129137f $X=7.83 $Y=1.295 $X2=0 $Y2=0
cc_381 N_A_c_181_n N_Y_c_837_n 5.34739e-19 $X=10.71 $Y=1.295 $X2=0 $Y2=0
cc_382 N_A_c_204_n N_Y_c_838_n 0.00394046f $X=10.565 $Y=1.765 $X2=0 $Y2=0
cc_383 N_A_c_205_n N_Y_c_838_n 0.00394046f $X=11.015 $Y=1.765 $X2=0 $Y2=0
cc_384 N_A_c_172_n N_Y_c_838_n 0.00412535f $X=10.75 $Y=1.485 $X2=0 $Y2=0
cc_385 N_A_c_180_n N_Y_c_838_n 0.0129137f $X=7.83 $Y=1.295 $X2=0 $Y2=0
cc_386 N_A_c_181_n N_Y_c_838_n 5.34739e-19 $X=10.71 $Y=1.295 $X2=0 $Y2=0
cc_387 N_A_c_182_n N_Y_c_956_n 0.00192824f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_388 N_A_c_183_n N_Y_c_956_n 0.0103148f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_389 N_A_c_184_n N_Y_c_956_n 0.00800853f $X=1.405 $Y=1.765 $X2=0 $Y2=0
cc_390 N_A_c_185_n N_Y_c_956_n 0.00760965f $X=1.855 $Y=1.765 $X2=0 $Y2=0
cc_391 N_A_c_186_n N_Y_c_956_n 0.00800853f $X=2.305 $Y=1.765 $X2=0 $Y2=0
cc_392 N_A_c_187_n N_Y_c_956_n 0.00800853f $X=2.755 $Y=1.765 $X2=0 $Y2=0
cc_393 N_A_c_188_n N_Y_c_956_n 0.00929017f $X=3.205 $Y=1.765 $X2=0 $Y2=0
cc_394 N_A_c_189_n N_Y_c_956_n 0.00800853f $X=3.655 $Y=1.765 $X2=0 $Y2=0
cc_395 N_A_c_190_n N_Y_c_956_n 0.00760965f $X=4.105 $Y=1.765 $X2=0 $Y2=0
cc_396 N_A_c_191_n N_Y_c_956_n 0.00776772f $X=4.555 $Y=1.765 $X2=0 $Y2=0
cc_397 N_A_c_192_n N_Y_c_956_n 0.00715379f $X=5.005 $Y=1.765 $X2=0 $Y2=0
cc_398 N_A_c_193_n N_Y_c_956_n 0.00750353f $X=5.455 $Y=1.765 $X2=0 $Y2=0
cc_399 N_A_c_194_n N_Y_c_956_n 0.00946261f $X=5.955 $Y=1.765 $X2=0 $Y2=0
cc_400 N_A_c_195_n N_Y_c_956_n 0.00869249f $X=6.405 $Y=1.765 $X2=0 $Y2=0
cc_401 N_A_c_196_n N_Y_c_956_n 0.0107838f $X=6.905 $Y=1.765 $X2=0 $Y2=0
cc_402 N_A_c_197_n N_Y_c_956_n 0.00798792f $X=7.415 $Y=1.765 $X2=0 $Y2=0
cc_403 N_A_c_198_n N_Y_c_956_n 0.00715379f $X=7.865 $Y=1.765 $X2=0 $Y2=0
cc_404 N_A_c_199_n N_Y_c_956_n 0.00715379f $X=8.315 $Y=1.765 $X2=0 $Y2=0
cc_405 N_A_c_200_n N_Y_c_956_n 0.00866511f $X=8.765 $Y=1.765 $X2=0 $Y2=0
cc_406 N_A_c_201_n N_Y_c_956_n 0.00715379f $X=9.215 $Y=1.765 $X2=0 $Y2=0
cc_407 N_A_c_202_n N_Y_c_956_n 0.00715379f $X=9.665 $Y=1.765 $X2=0 $Y2=0
cc_408 N_A_c_203_n N_Y_c_956_n 0.00715379f $X=10.115 $Y=1.765 $X2=0 $Y2=0
cc_409 N_A_c_204_n N_Y_c_956_n 0.00715379f $X=10.565 $Y=1.765 $X2=0 $Y2=0
cc_410 N_A_c_172_n N_Y_c_956_n 0.0320851f $X=10.75 $Y=1.485 $X2=0 $Y2=0
cc_411 N_A_c_173_n N_Y_c_956_n 0.00296806f $X=1.13 $Y=1.295 $X2=0 $Y2=0
cc_412 N_A_c_174_n N_Y_c_956_n 0.00511094f $X=2.03 $Y=1.295 $X2=0 $Y2=0
cc_413 N_A_c_175_n N_Y_c_956_n 0.00514555f $X=3 $Y=1.295 $X2=0 $Y2=0
cc_414 N_A_c_176_n N_Y_c_956_n 0.00511094f $X=3.93 $Y=1.295 $X2=0 $Y2=0
cc_415 N_A_c_177_n N_Y_c_956_n 0.00609124f $X=4.92 $Y=1.295 $X2=0 $Y2=0
cc_416 N_A_c_178_n N_Y_c_956_n 0.00312154f $X=5.76 $Y=1.295 $X2=0 $Y2=0
cc_417 N_A_c_179_n N_Y_c_956_n 0.00312154f $X=6.71 $Y=1.295 $X2=0 $Y2=0
cc_418 N_A_c_180_n N_Y_c_956_n 0.0494857f $X=7.83 $Y=1.295 $X2=0 $Y2=0
cc_419 N_A_c_181_n N_Y_c_956_n 0.450235f $X=10.71 $Y=1.295 $X2=0 $Y2=0
cc_420 N_A_c_184_n N_Y_c_989_n 0.00123111f $X=1.405 $Y=1.765 $X2=0 $Y2=0
cc_421 N_A_c_185_n N_Y_c_989_n 0.00156012f $X=1.855 $Y=1.765 $X2=0 $Y2=0
cc_422 N_A_c_172_n N_Y_c_989_n 0.00228314f $X=10.75 $Y=1.485 $X2=0 $Y2=0
cc_423 N_A_c_181_n N_Y_c_989_n 0.00253287f $X=10.71 $Y=1.295 $X2=0 $Y2=0
cc_424 N_A_c_183_n N_Y_c_820_n 6.48882e-19 $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_425 N_A_M1004_g N_Y_c_820_n 0.00571583f $X=1.355 $Y=0.61 $X2=0 $Y2=0
cc_426 N_A_c_184_n N_Y_c_820_n 0.00235453f $X=1.405 $Y=1.765 $X2=0 $Y2=0
cc_427 N_A_M1008_g N_Y_c_820_n 0.00599297f $X=1.785 $Y=0.61 $X2=0 $Y2=0
cc_428 N_A_c_185_n N_Y_c_820_n 0.00110032f $X=1.855 $Y=1.765 $X2=0 $Y2=0
cc_429 N_A_c_172_n N_Y_c_820_n 0.0290857f $X=10.75 $Y=1.485 $X2=0 $Y2=0
cc_430 N_A_c_173_n N_Y_c_820_n 0.035204f $X=1.13 $Y=1.295 $X2=0 $Y2=0
cc_431 N_A_c_174_n N_Y_c_820_n 0.0358472f $X=2.03 $Y=1.295 $X2=0 $Y2=0
cc_432 N_A_c_181_n N_Y_c_820_n 0.029424f $X=10.71 $Y=1.295 $X2=0 $Y2=0
cc_433 N_A_c_186_n N_Y_c_1002_n 0.00123111f $X=2.305 $Y=1.765 $X2=0 $Y2=0
cc_434 N_A_c_187_n N_Y_c_1002_n 0.00156012f $X=2.755 $Y=1.765 $X2=0 $Y2=0
cc_435 N_A_c_181_n N_Y_c_1002_n 6.73203e-19 $X=10.71 $Y=1.295 $X2=0 $Y2=0
cc_436 N_A_c_185_n N_Y_c_821_n 6.08789e-19 $X=1.855 $Y=1.765 $X2=0 $Y2=0
cc_437 N_A_M1011_g N_Y_c_821_n 0.00635294f $X=2.285 $Y=0.61 $X2=0 $Y2=0
cc_438 N_A_c_186_n N_Y_c_821_n 0.00245617f $X=2.305 $Y=1.765 $X2=0 $Y2=0
cc_439 N_A_M1012_g N_Y_c_821_n 0.0132982f $X=2.715 $Y=0.61 $X2=0 $Y2=0
cc_440 N_A_c_187_n N_Y_c_821_n 0.00104269f $X=2.755 $Y=1.765 $X2=0 $Y2=0
cc_441 N_A_c_172_n N_Y_c_821_n 0.0336513f $X=10.75 $Y=1.485 $X2=0 $Y2=0
cc_442 N_A_c_174_n N_Y_c_821_n 0.0362983f $X=2.03 $Y=1.295 $X2=0 $Y2=0
cc_443 N_A_c_175_n N_Y_c_821_n 0.0357176f $X=3 $Y=1.295 $X2=0 $Y2=0
cc_444 N_A_c_181_n N_Y_c_821_n 0.0369752f $X=10.71 $Y=1.295 $X2=0 $Y2=0
cc_445 N_A_M1002_g N_VGND_c_1132_n 0.0119813f $X=0.495 $Y=0.61 $X2=0 $Y2=0
cc_446 N_A_M1003_g N_VGND_c_1132_n 4.54967e-19 $X=0.925 $Y=0.61 $X2=0 $Y2=0
cc_447 N_A_M1002_g N_VGND_c_1133_n 4.54759e-19 $X=0.495 $Y=0.61 $X2=0 $Y2=0
cc_448 N_A_M1003_g N_VGND_c_1133_n 0.00930829f $X=0.925 $Y=0.61 $X2=0 $Y2=0
cc_449 N_A_M1004_g N_VGND_c_1133_n 0.00206942f $X=1.355 $Y=0.61 $X2=0 $Y2=0
cc_450 N_A_c_172_n N_VGND_c_1133_n 5.34284e-19 $X=10.75 $Y=1.485 $X2=0 $Y2=0
cc_451 N_A_c_173_n N_VGND_c_1133_n 0.0142005f $X=1.13 $Y=1.295 $X2=0 $Y2=0
cc_452 N_A_c_181_n N_VGND_c_1133_n 0.00212703f $X=10.71 $Y=1.295 $X2=0 $Y2=0
cc_453 N_A_M1008_g N_VGND_c_1134_n 0.00221156f $X=1.785 $Y=0.61 $X2=0 $Y2=0
cc_454 N_A_M1011_g N_VGND_c_1134_n 0.00555924f $X=2.285 $Y=0.61 $X2=0 $Y2=0
cc_455 N_A_c_172_n N_VGND_c_1134_n 9.08282e-19 $X=10.75 $Y=1.485 $X2=0 $Y2=0
cc_456 N_A_c_174_n N_VGND_c_1134_n 0.0140607f $X=2.03 $Y=1.295 $X2=0 $Y2=0
cc_457 N_A_c_181_n N_VGND_c_1134_n 0.00216974f $X=10.71 $Y=1.295 $X2=0 $Y2=0
cc_458 N_A_M1012_g N_VGND_c_1135_n 0.00340406f $X=2.715 $Y=0.61 $X2=0 $Y2=0
cc_459 N_A_M1016_g N_VGND_c_1135_n 0.00420244f $X=3.215 $Y=0.61 $X2=0 $Y2=0
cc_460 N_A_c_172_n N_VGND_c_1135_n 9.08282e-19 $X=10.75 $Y=1.485 $X2=0 $Y2=0
cc_461 N_A_c_175_n N_VGND_c_1135_n 0.0125433f $X=3 $Y=1.295 $X2=0 $Y2=0
cc_462 N_A_c_181_n N_VGND_c_1135_n 0.00193559f $X=10.71 $Y=1.295 $X2=0 $Y2=0
cc_463 N_A_M1017_g N_VGND_c_1136_n 0.00473938f $X=3.645 $Y=0.61 $X2=0 $Y2=0
cc_464 N_A_M1021_g N_VGND_c_1136_n 0.00473938f $X=4.215 $Y=0.61 $X2=0 $Y2=0
cc_465 N_A_c_172_n N_VGND_c_1136_n 0.00128128f $X=10.75 $Y=1.485 $X2=0 $Y2=0
cc_466 N_A_c_176_n N_VGND_c_1136_n 0.0165894f $X=3.93 $Y=1.295 $X2=0 $Y2=0
cc_467 N_A_c_181_n N_VGND_c_1136_n 0.00255998f $X=10.71 $Y=1.295 $X2=0 $Y2=0
cc_468 N_A_M1022_g N_VGND_c_1137_n 0.00477591f $X=4.645 $Y=0.61 $X2=0 $Y2=0
cc_469 N_A_M1026_g N_VGND_c_1137_n 0.0045678f $X=5.215 $Y=0.61 $X2=0 $Y2=0
cc_470 N_A_c_172_n N_VGND_c_1137_n 0.00127722f $X=10.75 $Y=1.485 $X2=0 $Y2=0
cc_471 N_A_c_177_n N_VGND_c_1137_n 0.0160836f $X=4.92 $Y=1.295 $X2=0 $Y2=0
cc_472 N_A_c_181_n N_VGND_c_1137_n 0.00248193f $X=10.71 $Y=1.295 $X2=0 $Y2=0
cc_473 N_A_M1026_g N_VGND_c_1138_n 5.08429e-19 $X=5.215 $Y=0.61 $X2=0 $Y2=0
cc_474 N_A_M1029_g N_VGND_c_1138_n 0.00958043f $X=5.645 $Y=0.61 $X2=0 $Y2=0
cc_475 N_A_M1030_g N_VGND_c_1138_n 0.00199403f $X=6.075 $Y=0.61 $X2=0 $Y2=0
cc_476 N_A_c_172_n N_VGND_c_1138_n 5.32878e-19 $X=10.75 $Y=1.485 $X2=0 $Y2=0
cc_477 N_A_c_178_n N_VGND_c_1138_n 0.0113456f $X=5.76 $Y=1.295 $X2=0 $Y2=0
cc_478 N_A_c_181_n N_VGND_c_1138_n 0.00431872f $X=10.71 $Y=1.295 $X2=0 $Y2=0
cc_479 N_A_M1030_g N_VGND_c_1139_n 4.63961e-19 $X=6.075 $Y=0.61 $X2=0 $Y2=0
cc_480 N_A_M1034_g N_VGND_c_1139_n 0.0098413f $X=6.505 $Y=0.61 $X2=0 $Y2=0
cc_481 N_A_M1036_g N_VGND_c_1139_n 0.00904542f $X=6.935 $Y=0.61 $X2=0 $Y2=0
cc_482 N_A_M1039_g N_VGND_c_1139_n 4.54543e-19 $X=7.365 $Y=0.61 $X2=0 $Y2=0
cc_483 N_A_c_172_n N_VGND_c_1139_n 5.34284e-19 $X=10.75 $Y=1.485 $X2=0 $Y2=0
cc_484 N_A_c_179_n N_VGND_c_1139_n 0.0157891f $X=6.71 $Y=1.295 $X2=0 $Y2=0
cc_485 N_A_c_181_n N_VGND_c_1139_n 0.00245282f $X=10.71 $Y=1.295 $X2=0 $Y2=0
cc_486 N_A_M1002_g N_VGND_c_1140_n 0.00462012f $X=0.495 $Y=0.61 $X2=0 $Y2=0
cc_487 N_A_M1003_g N_VGND_c_1140_n 0.00462012f $X=0.925 $Y=0.61 $X2=0 $Y2=0
cc_488 N_A_M1004_g N_VGND_c_1142_n 0.0055601f $X=1.355 $Y=0.61 $X2=0 $Y2=0
cc_489 N_A_M1008_g N_VGND_c_1142_n 0.0055601f $X=1.785 $Y=0.61 $X2=0 $Y2=0
cc_490 N_A_M1011_g N_VGND_c_1144_n 0.00546502f $X=2.285 $Y=0.61 $X2=0 $Y2=0
cc_491 N_A_M1012_g N_VGND_c_1144_n 0.00530655f $X=2.715 $Y=0.61 $X2=0 $Y2=0
cc_492 N_A_M1016_g N_VGND_c_1146_n 0.0055601f $X=3.215 $Y=0.61 $X2=0 $Y2=0
cc_493 N_A_M1017_g N_VGND_c_1146_n 0.00530655f $X=3.645 $Y=0.61 $X2=0 $Y2=0
cc_494 N_A_M1021_g N_VGND_c_1148_n 0.00530655f $X=4.215 $Y=0.61 $X2=0 $Y2=0
cc_495 N_A_M1022_g N_VGND_c_1148_n 0.0055601f $X=4.645 $Y=0.61 $X2=0 $Y2=0
cc_496 N_A_M1026_g N_VGND_c_1150_n 0.00519063f $X=5.215 $Y=0.61 $X2=0 $Y2=0
cc_497 N_A_M1029_g N_VGND_c_1150_n 0.00462012f $X=5.645 $Y=0.61 $X2=0 $Y2=0
cc_498 N_A_M1030_g N_VGND_c_1152_n 0.0055601f $X=6.075 $Y=0.61 $X2=0 $Y2=0
cc_499 N_A_M1034_g N_VGND_c_1152_n 0.00462012f $X=6.505 $Y=0.61 $X2=0 $Y2=0
cc_500 N_A_M1039_g N_VGND_c_1156_n 0.00988344f $X=7.365 $Y=0.61 $X2=0 $Y2=0
cc_501 N_A_c_172_n N_VGND_c_1156_n 0.0126349f $X=10.75 $Y=1.485 $X2=0 $Y2=0
cc_502 N_A_c_180_n N_VGND_c_1156_n 0.0875864f $X=7.83 $Y=1.295 $X2=0 $Y2=0
cc_503 N_A_c_181_n N_VGND_c_1156_n 0.0192684f $X=10.71 $Y=1.295 $X2=0 $Y2=0
cc_504 N_A_M1002_g N_VGND_c_1158_n 0.00450456f $X=0.495 $Y=0.61 $X2=0 $Y2=0
cc_505 N_A_M1003_g N_VGND_c_1158_n 0.00450456f $X=0.925 $Y=0.61 $X2=0 $Y2=0
cc_506 N_A_M1004_g N_VGND_c_1158_n 0.00536257f $X=1.355 $Y=0.61 $X2=0 $Y2=0
cc_507 N_A_M1008_g N_VGND_c_1158_n 0.00536257f $X=1.785 $Y=0.61 $X2=0 $Y2=0
cc_508 N_A_M1011_g N_VGND_c_1158_n 0.00536257f $X=2.285 $Y=0.61 $X2=0 $Y2=0
cc_509 N_A_M1012_g N_VGND_c_1158_n 0.00536257f $X=2.715 $Y=0.61 $X2=0 $Y2=0
cc_510 N_A_M1016_g N_VGND_c_1158_n 0.00536257f $X=3.215 $Y=0.61 $X2=0 $Y2=0
cc_511 N_A_M1017_g N_VGND_c_1158_n 0.00536257f $X=3.645 $Y=0.61 $X2=0 $Y2=0
cc_512 N_A_M1021_g N_VGND_c_1158_n 0.00536257f $X=4.215 $Y=0.61 $X2=0 $Y2=0
cc_513 N_A_M1022_g N_VGND_c_1158_n 0.00536257f $X=4.645 $Y=0.61 $X2=0 $Y2=0
cc_514 N_A_M1026_g N_VGND_c_1158_n 0.00536257f $X=5.215 $Y=0.61 $X2=0 $Y2=0
cc_515 N_A_M1029_g N_VGND_c_1158_n 0.00450456f $X=5.645 $Y=0.61 $X2=0 $Y2=0
cc_516 N_A_M1030_g N_VGND_c_1158_n 0.00536257f $X=6.075 $Y=0.61 $X2=0 $Y2=0
cc_517 N_A_M1034_g N_VGND_c_1158_n 0.00450456f $X=6.505 $Y=0.61 $X2=0 $Y2=0
cc_518 N_A_M1036_g N_VGND_c_1158_n 0.00486206f $X=6.935 $Y=0.61 $X2=0 $Y2=0
cc_519 N_A_M1039_g N_VGND_c_1158_n 0.00536257f $X=7.365 $Y=0.61 $X2=0 $Y2=0
cc_520 N_A_M1036_g N_VGND_c_1159_n 0.0049908f $X=6.935 $Y=0.61 $X2=0 $Y2=0
cc_521 N_A_M1039_g N_VGND_c_1159_n 0.0055601f $X=7.365 $Y=0.61 $X2=0 $Y2=0
cc_522 N_VPWR_c_592_n N_Y_c_822_n 0.014552f $X=1.995 $Y=3.33 $X2=0 $Y2=0
cc_523 N_VPWR_c_573_n N_Y_c_822_n 0.0119791f $X=11.28 $Y=3.33 $X2=0 $Y2=0
cc_524 N_VPWR_c_594_n N_Y_c_823_n 0.014552f $X=2.895 $Y=3.33 $X2=0 $Y2=0
cc_525 N_VPWR_c_573_n N_Y_c_823_n 0.0119791f $X=11.28 $Y=3.33 $X2=0 $Y2=0
cc_526 N_VPWR_c_579_n N_Y_c_807_n 0.00151517f $X=3.88 $Y=1.985 $X2=0 $Y2=0
cc_527 N_VPWR_c_580_n N_Y_c_807_n 0.00588171f $X=4.78 $Y=1.985 $X2=0 $Y2=0
cc_528 N_VPWR_c_581_n N_Y_c_809_n 0.00740298f $X=5.68 $Y=1.985 $X2=0 $Y2=0
cc_529 N_VPWR_c_582_n N_Y_c_809_n 0.0075713f $X=6.63 $Y=1.985 $X2=0 $Y2=0
cc_530 N_VPWR_c_576_n N_Y_c_826_n 0.0727885f $X=1.18 $Y=1.985 $X2=0 $Y2=0
cc_531 N_VPWR_c_579_n N_Y_c_888_n 0.0716012f $X=3.88 $Y=1.985 $X2=0 $Y2=0
cc_532 N_VPWR_c_580_n N_Y_c_892_n 0.0716175f $X=4.78 $Y=1.985 $X2=0 $Y2=0
cc_533 N_VPWR_c_580_n N_Y_c_815_n 0.00121873f $X=4.78 $Y=1.985 $X2=0 $Y2=0
cc_534 N_VPWR_c_581_n N_Y_c_815_n 0.0135808f $X=5.68 $Y=1.985 $X2=0 $Y2=0
cc_535 N_VPWR_c_575_n N_Y_c_829_n 0.0414236f $X=0.28 $Y=1.985 $X2=0 $Y2=0
cc_536 N_VPWR_c_590_n N_Y_c_829_n 0.00838873f $X=1.015 $Y=3.33 $X2=0 $Y2=0
cc_537 N_VPWR_c_573_n N_Y_c_829_n 0.00694347f $X=11.28 $Y=3.33 $X2=0 $Y2=0
cc_538 N_VPWR_c_578_n N_Y_c_818_n 0.0326929f $X=2.98 $Y=1.985 $X2=0 $Y2=0
cc_539 N_VPWR_c_579_n N_Y_c_818_n 0.0724821f $X=3.88 $Y=1.985 $X2=0 $Y2=0
cc_540 N_VPWR_c_596_n N_Y_c_818_n 0.0114703f $X=3.795 $Y=3.33 $X2=0 $Y2=0
cc_541 N_VPWR_c_573_n N_Y_c_818_n 0.00946127f $X=11.28 $Y=3.33 $X2=0 $Y2=0
cc_542 N_VPWR_c_580_n N_Y_c_831_n 0.0683223f $X=4.78 $Y=1.985 $X2=0 $Y2=0
cc_543 N_VPWR_c_598_n N_Y_c_831_n 0.014552f $X=4.695 $Y=3.33 $X2=0 $Y2=0
cc_544 N_VPWR_c_573_n N_Y_c_831_n 0.0119791f $X=11.28 $Y=3.33 $X2=0 $Y2=0
cc_545 N_VPWR_c_581_n N_Y_c_832_n 0.0635728f $X=5.68 $Y=1.985 $X2=0 $Y2=0
cc_546 N_VPWR_c_600_n N_Y_c_832_n 0.014552f $X=5.595 $Y=3.33 $X2=0 $Y2=0
cc_547 N_VPWR_c_573_n N_Y_c_832_n 0.0119791f $X=11.28 $Y=3.33 $X2=0 $Y2=0
cc_548 N_VPWR_c_581_n N_Y_c_833_n 0.0403783f $X=5.68 $Y=1.985 $X2=0 $Y2=0
cc_549 N_VPWR_c_582_n N_Y_c_833_n 0.0404231f $X=6.63 $Y=1.985 $X2=0 $Y2=0
cc_550 N_VPWR_c_602_n N_Y_c_833_n 0.0139245f $X=6.51 $Y=3.33 $X2=0 $Y2=0
cc_551 N_VPWR_c_573_n N_Y_c_833_n 0.0114926f $X=11.28 $Y=3.33 $X2=0 $Y2=0
cc_552 N_VPWR_c_582_n N_Y_c_819_n 0.0362611f $X=6.63 $Y=1.985 $X2=0 $Y2=0
cc_553 N_VPWR_c_583_n N_Y_c_819_n 0.0446363f $X=7.64 $Y=1.985 $X2=0 $Y2=0
cc_554 N_VPWR_c_604_n N_Y_c_819_n 0.0108429f $X=7.475 $Y=3.33 $X2=0 $Y2=0
cc_555 N_VPWR_c_573_n N_Y_c_819_n 0.0089748f $X=11.28 $Y=3.33 $X2=0 $Y2=0
cc_556 N_VPWR_c_583_n N_Y_c_835_n 0.0735935f $X=7.64 $Y=1.985 $X2=0 $Y2=0
cc_557 N_VPWR_c_584_n N_Y_c_835_n 0.00749631f $X=8.375 $Y=3.33 $X2=0 $Y2=0
cc_558 N_VPWR_c_585_n N_Y_c_835_n 0.0723029f $X=8.54 $Y=1.985 $X2=0 $Y2=0
cc_559 N_VPWR_c_573_n N_Y_c_835_n 0.0062048f $X=11.28 $Y=3.33 $X2=0 $Y2=0
cc_560 N_VPWR_c_585_n N_Y_c_836_n 0.0577412f $X=8.54 $Y=1.985 $X2=0 $Y2=0
cc_561 N_VPWR_c_586_n N_Y_c_836_n 0.0735935f $X=9.44 $Y=1.985 $X2=0 $Y2=0
cc_562 N_VPWR_c_606_n N_Y_c_836_n 0.00749631f $X=9.275 $Y=3.33 $X2=0 $Y2=0
cc_563 N_VPWR_c_573_n N_Y_c_836_n 0.0062048f $X=11.28 $Y=3.33 $X2=0 $Y2=0
cc_564 N_VPWR_c_586_n N_Y_c_837_n 0.0735935f $X=9.44 $Y=1.985 $X2=0 $Y2=0
cc_565 N_VPWR_c_587_n N_Y_c_837_n 0.0735935f $X=10.34 $Y=1.985 $X2=0 $Y2=0
cc_566 N_VPWR_c_607_n N_Y_c_837_n 0.00749631f $X=10.175 $Y=3.33 $X2=0 $Y2=0
cc_567 N_VPWR_c_573_n N_Y_c_837_n 0.0062048f $X=11.28 $Y=3.33 $X2=0 $Y2=0
cc_568 N_VPWR_c_587_n N_Y_c_838_n 0.0735935f $X=10.34 $Y=1.985 $X2=0 $Y2=0
cc_569 N_VPWR_c_589_n N_Y_c_838_n 0.072981f $X=11.24 $Y=1.985 $X2=0 $Y2=0
cc_570 N_VPWR_c_608_n N_Y_c_838_n 0.00749631f $X=11.075 $Y=3.33 $X2=0 $Y2=0
cc_571 N_VPWR_c_573_n N_Y_c_838_n 0.0062048f $X=11.28 $Y=3.33 $X2=0 $Y2=0
cc_572 N_VPWR_M1001_d N_Y_c_956_n 0.00320842f $X=1.03 $Y=1.84 $X2=0 $Y2=0
cc_573 N_VPWR_M1006_d N_Y_c_956_n 0.00629202f $X=1.93 $Y=1.84 $X2=0 $Y2=0
cc_574 N_VPWR_M1009_d N_Y_c_956_n 0.00618475f $X=2.83 $Y=1.84 $X2=0 $Y2=0
cc_575 N_VPWR_M1013_d N_Y_c_956_n 0.00629202f $X=3.73 $Y=1.84 $X2=0 $Y2=0
cc_576 N_VPWR_M1015_d N_Y_c_956_n 0.00640013f $X=4.63 $Y=1.84 $X2=0 $Y2=0
cc_577 N_VPWR_M1019_d N_Y_c_956_n 0.00492949f $X=5.53 $Y=1.84 $X2=0 $Y2=0
cc_578 N_VPWR_M1023_d N_Y_c_956_n 0.00304088f $X=6.48 $Y=1.84 $X2=0 $Y2=0
cc_579 N_VPWR_M1028_d N_Y_c_956_n 0.0030836f $X=8.39 $Y=1.84 $X2=0 $Y2=0
cc_580 N_VPWR_c_575_n N_Y_c_956_n 0.00707614f $X=0.28 $Y=1.985 $X2=0 $Y2=0
cc_581 N_VPWR_c_576_n N_Y_c_956_n 0.0290346f $X=1.18 $Y=1.985 $X2=0 $Y2=0
cc_582 N_VPWR_c_577_n N_Y_c_956_n 0.0213209f $X=2.08 $Y=1.985 $X2=0 $Y2=0
cc_583 N_VPWR_c_578_n N_Y_c_956_n 0.0220331f $X=2.98 $Y=1.985 $X2=0 $Y2=0
cc_584 N_VPWR_c_579_n N_Y_c_956_n 0.0213209f $X=3.88 $Y=1.985 $X2=0 $Y2=0
cc_585 N_VPWR_c_580_n N_Y_c_956_n 0.0214674f $X=4.78 $Y=1.985 $X2=0 $Y2=0
cc_586 N_VPWR_c_581_n N_Y_c_956_n 0.0287563f $X=5.68 $Y=1.985 $X2=0 $Y2=0
cc_587 N_VPWR_c_582_n N_Y_c_956_n 0.033123f $X=6.63 $Y=1.985 $X2=0 $Y2=0
cc_588 N_VPWR_c_583_n N_Y_c_956_n 0.0366973f $X=7.64 $Y=1.985 $X2=0 $Y2=0
cc_589 N_VPWR_c_585_n N_Y_c_956_n 0.0298424f $X=8.54 $Y=1.985 $X2=0 $Y2=0
cc_590 N_VPWR_c_586_n N_Y_c_956_n 0.0367409f $X=9.44 $Y=1.985 $X2=0 $Y2=0
cc_591 N_VPWR_c_587_n N_Y_c_956_n 0.0367409f $X=10.34 $Y=1.985 $X2=0 $Y2=0
cc_592 N_VPWR_c_589_n N_Y_c_956_n 0.0079968f $X=11.24 $Y=1.985 $X2=0 $Y2=0
cc_593 N_VPWR_c_577_n N_Y_c_989_n 0.069305f $X=2.08 $Y=1.985 $X2=0 $Y2=0
cc_594 N_VPWR_c_576_n N_Y_c_820_n 0.0752512f $X=1.18 $Y=1.985 $X2=0 $Y2=0
cc_595 N_VPWR_c_577_n N_Y_c_820_n 0.00321305f $X=2.08 $Y=1.985 $X2=0 $Y2=0
cc_596 N_VPWR_c_578_n N_Y_c_1002_n 0.069305f $X=2.98 $Y=1.985 $X2=0 $Y2=0
cc_597 N_VPWR_c_577_n N_Y_c_821_n 0.0735027f $X=2.08 $Y=1.985 $X2=0 $Y2=0
cc_598 N_VPWR_c_578_n N_Y_c_821_n 0.00254626f $X=2.98 $Y=1.985 $X2=0 $Y2=0
cc_599 N_Y_c_806_n N_VGND_c_1132_n 0.0155484f $X=0.71 $Y=0.61 $X2=0 $Y2=0
cc_600 N_Y_c_811_n N_VGND_c_1132_n 0.00302225f $X=0.72 $Y=1.82 $X2=0 $Y2=0
cc_601 N_Y_c_806_n N_VGND_c_1133_n 0.0183251f $X=0.71 $Y=0.61 $X2=0 $Y2=0
cc_602 N_Y_c_812_n N_VGND_c_1133_n 0.00147481f $X=1.57 $Y=0.61 $X2=0 $Y2=0
cc_603 N_Y_c_820_n N_VGND_c_1133_n 0.00133383f $X=1.63 $Y=1.885 $X2=0 $Y2=0
cc_604 N_Y_c_812_n N_VGND_c_1134_n 0.00144467f $X=1.57 $Y=0.61 $X2=0 $Y2=0
cc_605 N_Y_c_813_n N_VGND_c_1134_n 0.0144782f $X=2.5 $Y=0.61 $X2=0 $Y2=0
cc_606 N_Y_c_820_n N_VGND_c_1134_n 0.00140486f $X=1.63 $Y=1.885 $X2=0 $Y2=0
cc_607 N_Y_c_821_n N_VGND_c_1134_n 0.00138266f $X=2.53 $Y=1.885 $X2=0 $Y2=0
cc_608 N_Y_c_813_n N_VGND_c_1135_n 0.0177734f $X=2.5 $Y=0.61 $X2=0 $Y2=0
cc_609 N_Y_c_814_n N_VGND_c_1135_n 0.00134573f $X=3.43 $Y=0.61 $X2=0 $Y2=0
cc_610 N_Y_c_818_n N_VGND_c_1135_n 0.00119432f $X=3.43 $Y=1.985 $X2=0 $Y2=0
cc_611 N_Y_c_807_n N_VGND_c_1136_n 0.0182221f $X=4.43 $Y=0.61 $X2=0 $Y2=0
cc_612 N_Y_c_814_n N_VGND_c_1136_n 0.0184653f $X=3.43 $Y=0.61 $X2=0 $Y2=0
cc_613 N_Y_c_807_n N_VGND_c_1137_n 0.002434f $X=4.43 $Y=0.61 $X2=0 $Y2=0
cc_614 N_Y_c_815_n N_VGND_c_1137_n 0.0029897f $X=5.245 $Y=1.85 $X2=0 $Y2=0
cc_615 N_Y_c_816_n N_VGND_c_1137_n 0.0151326f $X=5.43 $Y=0.61 $X2=0 $Y2=0
cc_616 N_Y_c_810_n N_VGND_c_1138_n 0.002894f $X=6.29 $Y=0.61 $X2=0 $Y2=0
cc_617 N_Y_c_815_n N_VGND_c_1138_n 0.00335516f $X=5.245 $Y=1.85 $X2=0 $Y2=0
cc_618 N_Y_c_816_n N_VGND_c_1138_n 0.0152177f $X=5.43 $Y=0.61 $X2=0 $Y2=0
cc_619 N_Y_c_810_n N_VGND_c_1139_n 0.0158711f $X=6.29 $Y=0.61 $X2=0 $Y2=0
cc_620 N_Y_c_817_n N_VGND_c_1139_n 0.00339272f $X=6.217 $Y=1.01 $X2=0 $Y2=0
cc_621 N_Y_c_819_n N_VGND_c_1139_n 0.0186904f $X=7.15 $Y=0.61 $X2=0 $Y2=0
cc_622 N_Y_c_806_n N_VGND_c_1140_n 0.00747177f $X=0.71 $Y=0.61 $X2=0 $Y2=0
cc_623 N_Y_c_812_n N_VGND_c_1142_n 0.0102362f $X=1.57 $Y=0.61 $X2=0 $Y2=0
cc_624 N_Y_c_813_n N_VGND_c_1144_n 0.0123489f $X=2.5 $Y=0.61 $X2=0 $Y2=0
cc_625 N_Y_c_814_n N_VGND_c_1146_n 0.0115462f $X=3.43 $Y=0.61 $X2=0 $Y2=0
cc_626 N_Y_c_807_n N_VGND_c_1148_n 0.0102039f $X=4.43 $Y=0.61 $X2=0 $Y2=0
cc_627 N_Y_c_816_n N_VGND_c_1150_n 0.0102099f $X=5.43 $Y=0.61 $X2=0 $Y2=0
cc_628 N_Y_c_810_n N_VGND_c_1152_n 0.00881546f $X=6.29 $Y=0.61 $X2=0 $Y2=0
cc_629 N_Y_c_819_n N_VGND_c_1156_n 0.0121454f $X=7.15 $Y=0.61 $X2=0 $Y2=0
cc_630 N_Y_c_806_n N_VGND_c_1158_n 0.0068104f $X=0.71 $Y=0.61 $X2=0 $Y2=0
cc_631 N_Y_c_807_n N_VGND_c_1158_n 0.0093336f $X=4.43 $Y=0.61 $X2=0 $Y2=0
cc_632 N_Y_c_810_n N_VGND_c_1158_n 0.00805707f $X=6.29 $Y=0.61 $X2=0 $Y2=0
cc_633 N_Y_c_812_n N_VGND_c_1158_n 0.00933832f $X=1.57 $Y=0.61 $X2=0 $Y2=0
cc_634 N_Y_c_813_n N_VGND_c_1158_n 0.0113107f $X=2.5 $Y=0.61 $X2=0 $Y2=0
cc_635 N_Y_c_814_n N_VGND_c_1158_n 0.0105796f $X=3.43 $Y=0.61 $X2=0 $Y2=0
cc_636 N_Y_c_816_n N_VGND_c_1158_n 0.00956929f $X=5.43 $Y=0.61 $X2=0 $Y2=0
cc_637 N_Y_c_819_n N_VGND_c_1158_n 0.00881068f $X=7.15 $Y=0.61 $X2=0 $Y2=0
cc_638 N_Y_c_819_n N_VGND_c_1159_n 0.0096752f $X=7.15 $Y=0.61 $X2=0 $Y2=0
