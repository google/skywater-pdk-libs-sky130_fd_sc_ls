# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_ls__buf_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_ls__buf_16 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.56000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  1.674000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.775000 1.350000 10.435000 1.780000 ;
    END
  END A
  PIN VNB
    PORT
      LAYER pwell ;
        RECT 0.000000 0.000000 10.560000 0.245000 ;
    END
  END VNB
  PIN VPB
    PORT
      LAYER nwell ;
        RECT -0.190000 1.660000 10.750000 3.520000 ;
    END
  END VPB
  PIN X
    ANTENNADIFFAREA  4.345600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.575000 1.920000 7.255000 2.150000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.560000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 10.560000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 10.560000 0.085000 ;
      RECT  0.000000  3.245000 10.560000 3.415000 ;
      RECT  0.115000  1.820000  0.365000 3.245000 ;
      RECT  0.130000  0.085000  0.380000 1.130000 ;
      RECT  0.560000  0.350000  0.815000 2.980000 ;
      RECT  0.985000  1.300000  1.295000 1.780000 ;
      RECT  0.990000  0.085000  1.285000 1.130000 ;
      RECT  1.095000  1.965000  1.265000 3.245000 ;
      RECT  1.465000  0.350000  1.720000 2.980000 ;
      RECT  1.890000  1.300000  2.175000 1.780000 ;
      RECT  1.895000  0.085000  2.100000 1.130000 ;
      RECT  1.965000  1.965000  2.215000 3.245000 ;
      RECT  2.345000  0.350000  2.610000 1.185000 ;
      RECT  2.345000  1.185000  2.675000 1.355000 ;
      RECT  2.415000  1.355000  2.675000 2.980000 ;
      RECT  2.790000  0.085000  2.960000 1.015000 ;
      RECT  2.845000  1.300000  3.140000 1.780000 ;
      RECT  2.945000  1.965000  3.115000 3.245000 ;
      RECT  3.220000  0.350000  3.480000 1.130000 ;
      RECT  3.310000  1.130000  3.480000 1.820000 ;
      RECT  3.310000  1.820000  3.565000 2.980000 ;
      RECT  3.650000  0.085000  3.820000 1.130000 ;
      RECT  3.655000  1.300000  4.045000 1.655000 ;
      RECT  3.735000  1.655000  4.045000 1.780000 ;
      RECT  3.845000  1.965000  4.015000 3.245000 ;
      RECT  4.000000  0.350000  4.385000 1.130000 ;
      RECT  4.215000  1.130000  4.385000 1.900000 ;
      RECT  4.215000  1.900000  4.545000 2.980000 ;
      RECT  4.555000  0.085000  4.830000 1.130000 ;
      RECT  4.555000  1.300000  4.865000 1.730000 ;
      RECT  4.675000  1.730000  4.865000 1.780000 ;
      RECT  4.745000  1.965000  4.915000 3.245000 ;
      RECT  5.035000  0.350000  5.330000 1.205000 ;
      RECT  5.035000  1.205000  5.410000 1.375000 ;
      RECT  5.115000  1.375000  5.410000 2.980000 ;
      RECT  5.500000  0.085000  5.830000 1.035000 ;
      RECT  5.580000  1.300000  5.890000 1.780000 ;
      RECT  5.645000  1.965000  5.815000 3.245000 ;
      RECT  6.000000  0.350000  6.330000 1.130000 ;
      RECT  6.060000  1.130000  6.330000 2.980000 ;
      RECT  6.500000  0.085000  6.830000 1.130000 ;
      RECT  6.500000  1.300000  6.810000 1.780000 ;
      RECT  6.545000  1.965000  6.715000 3.245000 ;
      RECT  6.980000  1.250000  7.245000 2.980000 ;
      RECT  7.000000  0.350000  7.250000 1.250000 ;
      RECT  7.420000  1.010000  9.945000 1.180000 ;
      RECT  7.420000  1.180000  7.590000 1.950000 ;
      RECT  7.420000  1.950000  9.995000 2.120000 ;
      RECT  7.430000  0.085000  7.760000 0.840000 ;
      RECT  7.445000  2.290000  7.695000 3.245000 ;
      RECT  7.865000  2.120000  8.195000 2.980000 ;
      RECT  7.940000  0.350000  8.110000 1.010000 ;
      RECT  8.290000  0.085000  8.620000 0.840000 ;
      RECT  8.395000  2.290000  8.565000 3.245000 ;
      RECT  8.765000  2.120000  9.095000 2.980000 ;
      RECT  8.800000  0.350000  8.970000 1.010000 ;
      RECT  9.150000  0.085000  9.480000 0.840000 ;
      RECT  9.295000  2.290000  9.465000 3.245000 ;
      RECT  9.665000  2.120000  9.995000 2.980000 ;
      RECT  9.695000  0.350000  9.945000 1.010000 ;
      RECT 10.115000  0.085000 10.445000 1.130000 ;
      RECT 10.195000  1.950000 10.445000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  1.950000  0.805000 2.120000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.055000  1.580000  1.225000 1.750000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.515000  1.950000  1.685000 2.120000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  1.950000  1.580000  2.120000 1.750000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.470000  1.950000  2.640000 2.120000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  2.910000  1.580000  3.080000 1.750000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.360000  1.950000  3.530000 2.120000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.800000  1.580000  3.970000 1.750000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.300000  1.950000  4.470000 2.120000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.680000  1.580000  4.850000 1.750000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.195000  1.950000  5.365000 2.120000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.650000  1.580000  5.820000 1.750000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.095000  1.950000  6.265000 2.120000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.565000  1.580000  6.735000 1.750000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.025000  1.950000  7.195000 2.120000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.420000  1.580000  7.590000 1.750000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
    LAYER met1 ;
      RECT 0.985000 1.550000 7.650000 1.780000 ;
  END
END sky130_fd_sc_ls__buf_16
END LIBRARY
