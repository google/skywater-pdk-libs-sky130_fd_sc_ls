* File: sky130_fd_sc_ls__nand4_2.spice
* Created: Fri Aug 28 13:34:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__nand4_2.pex.spice"
.subckt sky130_fd_sc_ls__nand4_2  VNB VPB D C B A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* B	B
* C	C
* D	D
* VPB	VPB
* VNB	VNB
MM1001 N_A_27_74#_M1001_d N_D_M1001_g N_VGND_M1001_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.1369 PD=2.05 PS=1.11 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75000.2
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1011 N_A_27_74#_M1011_d N_D_M1011_g N_VGND_M1001_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1369 PD=1.02 PS=1.11 NRD=0 NRS=3.24 M=1 R=4.93333 SA=75000.7
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1007 N_A_304_74#_M1007_d N_C_M1007_g N_A_27_74#_M1011_d VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.2 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1013 N_A_304_74#_M1007_d N_C_M1013_g N_A_27_74#_M1013_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.23225 PD=1.02 PS=2.19 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75001.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1004 N_A_515_74#_M1004_d N_B_M1004_g N_A_304_74#_M1004_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1983 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001.5 A=0.111 P=1.78 MULT=1
MM1012 N_A_515_74#_M1012_d N_B_M1012_g N_A_304_74#_M1004_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1010 N_Y_M1010_d N_A_M1010_g N_A_515_74#_M1012_d VNB NSHORT L=0.15 W=0.74
+ AD=0.111 AS=0.1036 PD=1.04 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1015 N_Y_M1010_d N_A_M1015_g N_A_515_74#_M1015_s VNB NSHORT L=0.15 W=0.74
+ AD=0.111 AS=0.22325 PD=1.04 PS=2.15 NRD=3.24 NRS=8.1 M=1 R=4.93333 SA=75001.5
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1006 N_Y_M1006_d N_D_M1006_g N_VPWR_M1006_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.1904 AS=0.336 PD=1.46 PS=2.84 NRD=1.7533 NRS=2.6201 M=1 R=7.46667
+ SA=75000.2 SB=75004 A=0.168 P=2.54 MULT=1
MM1009 N_Y_M1006_d N_D_M1009_g N_VPWR_M1009_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.1904 AS=0.1904 PD=1.46 PS=1.46 NRD=8.7862 NRS=3.5066 M=1 R=7.46667
+ SA=75000.7 SB=75003.5 A=0.168 P=2.54 MULT=1
MM1000 N_Y_M1000_d N_C_M1000_g N_VPWR_M1009_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.1792 AS=0.1904 PD=1.44 PS=1.46 NRD=5.2599 NRS=7.0329 M=1 R=7.46667
+ SA=75001.2 SB=75003 A=0.168 P=2.54 MULT=1
MM1014 N_Y_M1000_d N_C_M1014_g N_VPWR_M1014_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.1792 AS=0.3696 PD=1.44 PS=1.78 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.7 SB=75002.5 A=0.168 P=2.54 MULT=1
MM1002 N_Y_M1002_d N_B_M1002_g N_VPWR_M1014_s VPB PHIGHVT L=0.15 W=1.12 AD=0.168
+ AS=0.3696 PD=1.42 PS=1.78 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75002.5
+ SB=75001.7 A=0.168 P=2.54 MULT=1
MM1005 N_Y_M1002_d N_B_M1005_g N_VPWR_M1005_s VPB PHIGHVT L=0.15 W=1.12 AD=0.168
+ AS=0.2296 PD=1.42 PS=1.53 NRD=1.7533 NRS=10.5395 M=1 R=7.46667 SA=75002.9
+ SB=75001.2 A=0.168 P=2.54 MULT=1
MM1003 N_Y_M1003_d N_A_M1003_g N_VPWR_M1005_s VPB PHIGHVT L=0.15 W=1.12 AD=0.168
+ AS=0.2296 PD=1.42 PS=1.53 NRD=1.7533 NRS=12.2928 M=1 R=7.46667 SA=75003.5
+ SB=75000.7 A=0.168 P=2.54 MULT=1
MM1008 N_Y_M1003_d N_A_M1008_g N_VPWR_M1008_s VPB PHIGHVT L=0.15 W=1.12 AD=0.168
+ AS=0.3528 PD=1.42 PS=2.87 NRD=1.7533 NRS=2.6201 M=1 R=7.46667 SA=75003.9
+ SB=75000.2 A=0.168 P=2.54 MULT=1
DX16_noxref VNB VPB NWDIODE A=9.6348 P=14.08
*
.include "sky130_fd_sc_ls__nand4_2.pxi.spice"
*
.ends
*
*
