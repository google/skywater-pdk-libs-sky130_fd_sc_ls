* NGSPICE file created from sky130_fd_sc_ls__nand2_8.ext - technology: sky130A

.subckt sky130_fd_sc_ls__nand2_8 A B VGND VNB VPB VPWR Y
M1000 VGND B a_27_74# VNB nshort w=740000u l=150000u
+  ad=1.0656e+12p pd=8.8e+06u as=2.14795e+12p ps=1.918e+07u
M1001 a_27_74# A Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=8.288e+11p ps=8.16e+06u
M1002 a_27_74# A Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPWR B Y VPB phighvt w=1.12e+06u l=150000u
+  ad=5.1352e+12p pd=2.261e+07u as=1.456e+12p ps=1.156e+07u
M1004 VPWR B Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y A a_27_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y A VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR A Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y A a_27_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR A Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_27_74# B VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND B a_27_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND B a_27_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_27_74# A Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Y A a_27_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_27_74# B VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_27_74# B VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 Y A a_27_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 Y B VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 Y B VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_27_74# A Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND B a_27_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_27_74# B VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 Y A VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

