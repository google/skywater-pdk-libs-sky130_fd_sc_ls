* File: sky130_fd_sc_ls__o21ai_1.pxi.spice
* Created: Wed Sep  2 11:18:12 2020
* 
x_PM_SKY130_FD_SC_LS__O21AI_1%A1 N_A1_c_36_n N_A1_M1003_g N_A1_c_37_n
+ N_A1_M1000_g A1 N_A1_c_38_n PM_SKY130_FD_SC_LS__O21AI_1%A1
x_PM_SKY130_FD_SC_LS__O21AI_1%A2 N_A2_c_62_n N_A2_M1004_g N_A2_M1001_g A2
+ N_A2_c_64_n PM_SKY130_FD_SC_LS__O21AI_1%A2
x_PM_SKY130_FD_SC_LS__O21AI_1%B1 N_B1_c_91_n N_B1_M1005_g N_B1_M1002_g B1 B1
+ PM_SKY130_FD_SC_LS__O21AI_1%B1
x_PM_SKY130_FD_SC_LS__O21AI_1%VPWR N_VPWR_M1000_s N_VPWR_M1005_d N_VPWR_c_115_n
+ N_VPWR_c_116_n N_VPWR_c_117_n N_VPWR_c_118_n N_VPWR_c_119_n VPWR
+ N_VPWR_c_120_n N_VPWR_c_114_n PM_SKY130_FD_SC_LS__O21AI_1%VPWR
x_PM_SKY130_FD_SC_LS__O21AI_1%Y N_Y_M1002_d N_Y_M1004_d N_Y_c_139_n N_Y_c_140_n
+ N_Y_c_141_n Y Y N_Y_c_143_n N_Y_c_142_n PM_SKY130_FD_SC_LS__O21AI_1%Y
x_PM_SKY130_FD_SC_LS__O21AI_1%A_27_74# N_A_27_74#_M1003_s N_A_27_74#_M1001_d
+ N_A_27_74#_c_177_n N_A_27_74#_c_181_n N_A_27_74#_c_178_n N_A_27_74#_c_179_n
+ PM_SKY130_FD_SC_LS__O21AI_1%A_27_74#
x_PM_SKY130_FD_SC_LS__O21AI_1%VGND N_VGND_M1003_d VGND N_VGND_c_208_n
+ N_VGND_c_209_n N_VGND_c_210_n N_VGND_c_211_n PM_SKY130_FD_SC_LS__O21AI_1%VGND
cc_1 VNB N_A1_c_36_n 0.0240813f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.22
cc_2 VNB N_A1_c_37_n 0.0724919f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=1.765
cc_3 VNB N_A1_c_38_n 0.0206951f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.385
cc_4 VNB N_A2_c_62_n 0.0322642f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.22
cc_5 VNB N_A2_M1001_g 0.0268063f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=2.4
cc_6 VNB N_A2_c_64_n 0.00245973f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.365
cc_7 VNB N_B1_c_91_n 0.0276824f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.22
cc_8 VNB N_B1_M1002_g 0.0329453f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=2.4
cc_9 VNB B1 0.01855f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.385
cc_10 VNB N_VPWR_c_114_n 0.103974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_Y_c_139_n 0.0231532f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.385
cc_12 VNB N_Y_c_140_n 7.88229e-19 $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.385
cc_13 VNB N_Y_c_141_n 0.0281704f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_Y_c_142_n 0.00413149f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_74#_c_177_n 0.0149177f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.385
cc_16 VNB N_A_27_74#_c_178_n 0.0139746f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.365
cc_17 VNB N_A_27_74#_c_179_n 0.00256335f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_VGND_c_208_n 0.031602f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_VGND_c_209_n 0.159013f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_210_n 0.0182531f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_211_n 0.023075f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VPB N_A1_c_37_n 0.0269034f $X=-0.19 $Y=1.66 $X2=0.735 $Y2=1.765
cc_23 VPB N_A2_c_62_n 0.0309127f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.22
cc_24 VPB N_A2_c_64_n 0.00240305f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.365
cc_25 VPB N_B1_c_91_n 0.0328561f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.22
cc_26 VPB B1 0.0182438f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=1.385
cc_27 VPB N_VPWR_c_115_n 0.015156f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=1.385
cc_28 VPB N_VPWR_c_116_n 0.0147219f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_29 VPB N_VPWR_c_117_n 0.0486246f $X=-0.19 $Y=1.66 $X2=0.39 $Y2=1.365
cc_30 VPB N_VPWR_c_118_n 0.011849f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_31 VPB N_VPWR_c_119_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_32 VPB N_VPWR_c_120_n 0.0352341f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_33 VPB N_VPWR_c_114_n 0.0727985f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_34 VPB N_Y_c_143_n 0.00526404f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_35 VPB N_Y_c_142_n 0.00129742f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_36 N_A1_c_37_n N_A2_c_62_n 0.0837915f $X=0.735 $Y=1.765 $X2=-0.19 $Y2=-0.245
cc_37 N_A1_c_37_n N_A2_M1001_g 0.00239f $X=0.735 $Y=1.765 $X2=0 $Y2=0
cc_38 N_A1_c_37_n N_A2_c_64_n 5.01684e-19 $X=0.735 $Y=1.765 $X2=0 $Y2=0
cc_39 N_A1_c_37_n N_VPWR_c_115_n 0.0149384f $X=0.735 $Y=1.765 $X2=0 $Y2=0
cc_40 N_A1_c_38_n N_VPWR_c_115_n 0.0149317f $X=0.39 $Y=1.385 $X2=0 $Y2=0
cc_41 N_A1_c_37_n N_VPWR_c_120_n 0.00366292f $X=0.735 $Y=1.765 $X2=0 $Y2=0
cc_42 N_A1_c_37_n N_VPWR_c_114_n 0.00605395f $X=0.735 $Y=1.765 $X2=0 $Y2=0
cc_43 N_A1_c_36_n N_Y_c_140_n 0.00710272f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_44 N_A1_c_37_n N_Y_c_143_n 0.0276669f $X=0.735 $Y=1.765 $X2=0 $Y2=0
cc_45 N_A1_c_36_n N_Y_c_142_n 7.57456e-19 $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_46 N_A1_c_37_n N_Y_c_142_n 0.0281574f $X=0.735 $Y=1.765 $X2=0 $Y2=0
cc_47 N_A1_c_38_n N_Y_c_142_n 0.0270948f $X=0.39 $Y=1.385 $X2=0 $Y2=0
cc_48 N_A1_c_36_n N_A_27_74#_c_177_n 4.59808e-19 $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_49 N_A1_c_36_n N_A_27_74#_c_181_n 0.0116592f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_50 N_A1_c_37_n N_A_27_74#_c_181_n 0.00454671f $X=0.735 $Y=1.765 $X2=0 $Y2=0
cc_51 N_A1_c_38_n N_A_27_74#_c_181_n 0.00452942f $X=0.39 $Y=1.385 $X2=0 $Y2=0
cc_52 N_A1_c_36_n N_A_27_74#_c_178_n 0.00905744f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_53 N_A1_c_37_n N_A_27_74#_c_178_n 0.0012195f $X=0.735 $Y=1.765 $X2=0 $Y2=0
cc_54 N_A1_c_38_n N_A_27_74#_c_178_n 0.0250699f $X=0.39 $Y=1.385 $X2=0 $Y2=0
cc_55 N_A1_c_36_n N_VGND_c_209_n 0.00429381f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_56 N_A1_c_36_n N_VGND_c_210_n 0.00329909f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_57 N_A1_c_36_n N_VGND_c_211_n 0.00816535f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_58 N_A2_c_62_n N_B1_c_91_n 0.0347773f $X=1.155 $Y=1.765 $X2=-0.19 $Y2=-0.245
cc_59 N_A2_c_64_n N_B1_c_91_n 5.50397e-19 $X=1.23 $Y=1.515 $X2=-0.19 $Y2=-0.245
cc_60 N_A2_M1001_g N_B1_M1002_g 0.0331423f $X=1.405 $Y=0.74 $X2=0 $Y2=0
cc_61 N_A2_c_62_n B1 0.00293689f $X=1.155 $Y=1.765 $X2=0 $Y2=0
cc_62 N_A2_c_64_n B1 0.036629f $X=1.23 $Y=1.515 $X2=0 $Y2=0
cc_63 N_A2_c_62_n N_VPWR_c_117_n 7.87841e-19 $X=1.155 $Y=1.765 $X2=0 $Y2=0
cc_64 N_A2_c_62_n N_VPWR_c_120_n 0.00291513f $X=1.155 $Y=1.765 $X2=0 $Y2=0
cc_65 N_A2_c_62_n N_VPWR_c_114_n 0.00360842f $X=1.155 $Y=1.765 $X2=0 $Y2=0
cc_66 N_A2_c_62_n N_Y_c_139_n 0.00184613f $X=1.155 $Y=1.765 $X2=0 $Y2=0
cc_67 N_A2_M1001_g N_Y_c_139_n 0.0147665f $X=1.405 $Y=0.74 $X2=0 $Y2=0
cc_68 N_A2_c_64_n N_Y_c_139_n 0.0250422f $X=1.23 $Y=1.515 $X2=0 $Y2=0
cc_69 N_A2_c_62_n N_Y_c_143_n 0.0345605f $X=1.155 $Y=1.765 $X2=0 $Y2=0
cc_70 N_A2_c_64_n N_Y_c_143_n 0.024835f $X=1.23 $Y=1.515 $X2=0 $Y2=0
cc_71 N_A2_c_62_n N_Y_c_142_n 0.00583924f $X=1.155 $Y=1.765 $X2=0 $Y2=0
cc_72 N_A2_M1001_g N_Y_c_142_n 0.00317248f $X=1.405 $Y=0.74 $X2=0 $Y2=0
cc_73 N_A2_c_64_n N_Y_c_142_n 0.0323789f $X=1.23 $Y=1.515 $X2=0 $Y2=0
cc_74 N_A2_M1001_g N_A_27_74#_c_181_n 0.01182f $X=1.405 $Y=0.74 $X2=0 $Y2=0
cc_75 N_A2_M1001_g N_A_27_74#_c_179_n 5.92733e-19 $X=1.405 $Y=0.74 $X2=0 $Y2=0
cc_76 N_A2_M1001_g N_VGND_c_208_n 0.00329926f $X=1.405 $Y=0.74 $X2=0 $Y2=0
cc_77 N_A2_M1001_g N_VGND_c_209_n 0.00425862f $X=1.405 $Y=0.74 $X2=0 $Y2=0
cc_78 N_A2_M1001_g N_VGND_c_211_n 0.00816535f $X=1.405 $Y=0.74 $X2=0 $Y2=0
cc_79 N_B1_c_91_n N_VPWR_c_117_n 0.0200806f $X=1.81 $Y=1.765 $X2=0 $Y2=0
cc_80 B1 N_VPWR_c_117_n 0.0263294f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_81 N_B1_c_91_n N_VPWR_c_120_n 0.00413917f $X=1.81 $Y=1.765 $X2=0 $Y2=0
cc_82 N_B1_c_91_n N_VPWR_c_114_n 0.00819352f $X=1.81 $Y=1.765 $X2=0 $Y2=0
cc_83 N_B1_c_91_n N_Y_c_139_n 0.00423142f $X=1.81 $Y=1.765 $X2=0 $Y2=0
cc_84 N_B1_M1002_g N_Y_c_139_n 0.0158149f $X=1.835 $Y=0.74 $X2=0 $Y2=0
cc_85 B1 N_Y_c_139_n 0.0584272f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_86 N_B1_M1002_g N_Y_c_141_n 0.0128452f $X=1.835 $Y=0.74 $X2=0 $Y2=0
cc_87 N_B1_c_91_n N_Y_c_143_n 0.0109265f $X=1.81 $Y=1.765 $X2=0 $Y2=0
cc_88 N_B1_M1002_g N_A_27_74#_c_181_n 0.00214696f $X=1.835 $Y=0.74 $X2=0 $Y2=0
cc_89 N_B1_M1002_g N_A_27_74#_c_179_n 0.00475124f $X=1.835 $Y=0.74 $X2=0 $Y2=0
cc_90 N_B1_M1002_g N_VGND_c_208_n 0.00434272f $X=1.835 $Y=0.74 $X2=0 $Y2=0
cc_91 N_B1_M1002_g N_VGND_c_209_n 0.00825242f $X=1.835 $Y=0.74 $X2=0 $Y2=0
cc_92 N_VPWR_c_117_n N_Y_c_143_n 0.0516113f $X=2.035 $Y=2.115 $X2=0 $Y2=0
cc_93 N_VPWR_c_120_n N_Y_c_143_n 0.0358004f $X=1.87 $Y=3.33 $X2=0 $Y2=0
cc_94 N_VPWR_c_114_n N_Y_c_143_n 0.0290828f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_95 N_VPWR_c_115_n N_Y_c_142_n 0.0922411f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_96 A_162_368# N_Y_c_143_n 0.00577415f $X=0.81 $Y=1.84 $X2=1.38 $Y2=2.115
cc_97 A_162_368# N_Y_c_142_n 0.00127723f $X=0.81 $Y=1.84 $X2=1.135 $Y2=1.95
cc_98 N_Y_c_139_n N_A_27_74#_M1001_d 0.00176461f $X=1.955 $Y=1.095 $X2=0 $Y2=0
cc_99 N_Y_c_139_n N_A_27_74#_c_181_n 0.0525194f $X=1.955 $Y=1.095 $X2=0 $Y2=0
cc_100 N_Y_c_140_n N_A_27_74#_c_181_n 0.0138309f $X=0.895 $Y=1.095 $X2=0 $Y2=0
cc_101 N_Y_c_141_n N_A_27_74#_c_179_n 0.0126166f $X=2.12 $Y=0.515 $X2=0 $Y2=0
cc_102 N_Y_c_139_n N_VGND_M1003_d 0.00498687f $X=1.955 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_103 N_Y_c_140_n N_VGND_M1003_d 0.00350137f $X=0.895 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_104 N_Y_c_141_n N_VGND_c_208_n 0.0146357f $X=2.12 $Y=0.515 $X2=0 $Y2=0
cc_105 N_Y_c_141_n N_VGND_c_209_n 0.0121141f $X=2.12 $Y=0.515 $X2=0 $Y2=0
cc_106 N_A_27_74#_c_181_n N_VGND_M1003_d 0.0171612f $X=1.48 $Y=0.755 $X2=-0.19
+ $Y2=-0.245
cc_107 N_A_27_74#_c_181_n N_VGND_c_208_n 0.00255882f $X=1.48 $Y=0.755 $X2=0
+ $Y2=0
cc_108 N_A_27_74#_c_179_n N_VGND_c_208_n 0.0131355f $X=1.632 $Y=0.67 $X2=0 $Y2=0
cc_109 N_A_27_74#_c_177_n N_VGND_c_209_n 0.0111794f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_110 N_A_27_74#_c_181_n N_VGND_c_209_n 0.0111174f $X=1.48 $Y=0.755 $X2=0 $Y2=0
cc_111 N_A_27_74#_c_178_n N_VGND_c_209_n 5.83956e-19 $X=0.445 $Y=0.755 $X2=0
+ $Y2=0
cc_112 N_A_27_74#_c_179_n N_VGND_c_209_n 0.0109537f $X=1.632 $Y=0.67 $X2=0 $Y2=0
cc_113 N_A_27_74#_c_177_n N_VGND_c_210_n 0.0134907f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_114 N_A_27_74#_c_181_n N_VGND_c_210_n 0.00218193f $X=1.48 $Y=0.755 $X2=0
+ $Y2=0
cc_115 N_A_27_74#_c_178_n N_VGND_c_210_n 3.88305e-19 $X=0.445 $Y=0.755 $X2=0
+ $Y2=0
cc_116 N_A_27_74#_c_177_n N_VGND_c_211_n 0.00658978f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_117 N_A_27_74#_c_181_n N_VGND_c_211_n 0.0495128f $X=1.48 $Y=0.755 $X2=0 $Y2=0
cc_118 N_A_27_74#_c_179_n N_VGND_c_211_n 0.00309085f $X=1.632 $Y=0.67 $X2=0
+ $Y2=0
