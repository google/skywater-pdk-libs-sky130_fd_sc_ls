* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__xor2_2 A B VGND VNB VPB VPWR X
X0 a_313_368# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X1 VGND A a_399_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X2 a_399_74# A VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X3 X B a_399_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X4 X a_183_74# a_313_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X5 VPWR A a_313_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X6 VPWR A a_116_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 a_116_392# B a_183_74# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 a_313_368# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X9 VGND A a_183_74# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X10 a_399_74# B X VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X11 a_313_368# a_183_74# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X12 VGND a_183_74# X VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X13 VPWR B a_313_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X14 a_183_74# B VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
.ends
