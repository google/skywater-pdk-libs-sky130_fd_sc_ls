* File: sky130_fd_sc_ls__nand4bb_2.pex.spice
* Created: Wed Sep  2 11:13:36 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__NAND4BB_2%A_N 1 3 6 8 12
c36 12 0 1.87042e-19 $X=0.6 $Y=1.465
r37 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.6
+ $Y=1.465 $X2=0.6 $Y2=1.465
r38 8 12 5.76222 $w=3.98e-07 $l=2e-07 $layer=LI1_cond $X=0.635 $Y=1.665
+ $X2=0.635 $Y2=1.465
r39 4 11 38.5519 $w=3e-07 $l=2.0106e-07 $layer=POLY_cond $X=0.51 $Y=1.3 $X2=0.59
+ $Y2=1.465
r40 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.51 $Y=1.3 $X2=0.51
+ $Y2=0.69
r41 1 11 60.2419 $w=3e-07 $l=3.39853e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.59 $Y2=1.465
r42 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_LS__NAND4BB_2%B_N 3 6 7 9 10 13
c39 7 0 1.87042e-19 $X=1.125 $Y=1.765
r40 13 16 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.17 $Y=1.345
+ $X2=1.17 $Y2=1.51
r41 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.17 $Y=1.345
+ $X2=1.17 $Y2=1.18
r42 10 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.17
+ $Y=1.345 $X2=1.17 $Y2=1.345
r43 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.125 $Y=1.765
+ $X2=1.125 $Y2=2.34
r44 6 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.125 $Y=1.675 $X2=1.125
+ $Y2=1.765
r45 6 16 64.1371 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.125 $Y=1.675
+ $X2=1.125 $Y2=1.51
r46 3 15 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=1.08 $Y=0.69 $X2=1.08
+ $Y2=1.18
.ends

.subckt PM_SKY130_FD_SC_LS__NAND4BB_2%A_27_368# 1 2 7 9 10 12 13 15 16 18 19 22
+ 26 32 34 38 41 43 44
c97 13 0 2.48037e-20 $X=2.725 $Y=1.185
c98 7 0 1.41504e-19 $X=2.27 $Y=1.185
r99 43 45 9.54881 $w=3.48e-07 $l=2.9e-07 $layer=LI1_cond $X=0.27 $Y=2.035
+ $X2=0.27 $Y2=2.325
r100 43 44 5.85433 $w=3.48e-07 $l=8.5e-08 $layer=LI1_cond $X=0.27 $Y=2.035
+ $X2=0.27 $Y2=1.95
r101 41 44 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=0.18 $Y=1.03
+ $X2=0.18 $Y2=1.95
r102 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.01
+ $Y=1.515 $X2=2.01 $Y2=1.515
r103 36 38 25.3188 $w=3.28e-07 $l=7.25e-07 $layer=LI1_cond $X=2.01 $Y=2.24
+ $X2=2.01 $Y2=1.515
r104 35 45 4.974 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=0.445 $Y=2.325
+ $X2=0.27 $Y2=2.325
r105 34 36 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.845 $Y=2.325
+ $X2=2.01 $Y2=2.24
r106 34 35 91.3369 $w=1.68e-07 $l=1.4e-06 $layer=LI1_cond $X=1.845 $Y=2.325
+ $X2=0.445 $Y2=2.325
r107 30 45 2.79879 $w=3.48e-07 $l=8.5e-08 $layer=LI1_cond $X=0.27 $Y=2.41
+ $X2=0.27 $Y2=2.325
r108 30 32 10.0427 $w=3.48e-07 $l=3.05e-07 $layer=LI1_cond $X=0.27 $Y=2.41
+ $X2=0.27 $Y2=2.715
r109 24 41 9.06106 $w=3.63e-07 $l=1.82e-07 $layer=LI1_cond $X=0.277 $Y=0.848
+ $X2=0.277 $Y2=1.03
r110 24 26 10.5141 $w=3.63e-07 $l=3.33e-07 $layer=LI1_cond $X=0.277 $Y=0.848
+ $X2=0.277 $Y2=0.515
r111 22 23 0.932302 $w=5.17e-07 $l=1e-08 $layer=POLY_cond $X=2.725 $Y=1.475
+ $X2=2.735 $Y2=1.475
r112 21 22 41.0213 $w=5.17e-07 $l=4.4e-07 $layer=POLY_cond $X=2.285 $Y=1.475
+ $X2=2.725 $Y2=1.475
r113 20 21 1.39845 $w=5.17e-07 $l=1.5e-08 $layer=POLY_cond $X=2.27 $Y=1.475
+ $X2=2.285 $Y2=1.475
r114 19 39 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=2.195 $Y=1.515
+ $X2=2.01 $Y2=1.515
r115 19 20 13.276 $w=5.17e-07 $l=9.28709e-08 $layer=POLY_cond $X=2.195 $Y=1.515
+ $X2=2.27 $Y2=1.475
r116 16 23 32.2548 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.735 $Y=1.765
+ $X2=2.735 $Y2=1.475
r117 16 18 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.735 $Y=1.765
+ $X2=2.735 $Y2=2.4
r118 13 22 32.2548 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.725 $Y=1.185
+ $X2=2.725 $Y2=1.475
r119 13 15 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.725 $Y=1.185
+ $X2=2.725 $Y2=0.74
r120 10 21 32.2548 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.285 $Y=1.765
+ $X2=2.285 $Y2=1.475
r121 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.285 $Y=1.765
+ $X2=2.285 $Y2=2.4
r122 7 20 32.2548 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.27 $Y=1.185
+ $X2=2.27 $Y2=1.475
r123 7 9 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.27 $Y=1.185
+ $X2=2.27 $Y2=0.74
r124 2 43 400 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.035
r125 2 32 400 $w=1.7e-07 $l=9.44722e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.715
r126 1 26 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.15
+ $Y=0.37 $X2=0.295 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__NAND4BB_2%A_231_74# 1 2 7 9 12 14 16 19 21 25 26 27
+ 30 32 33 35 41 45
c103 30 0 8.4381e-20 $X=2.43 $Y=1.43
c104 12 0 6.95413e-20 $X=3.315 $Y=0.74
c105 7 0 1.36243e-19 $X=3.285 $Y=1.765
r106 45 46 1.29223 $w=3.73e-07 $l=1e-08 $layer=POLY_cond $X=3.735 $Y=1.557
+ $X2=3.745 $Y2=1.557
r107 42 43 3.87668 $w=3.73e-07 $l=3e-08 $layer=POLY_cond $X=3.285 $Y=1.557
+ $X2=3.315 $Y2=1.557
r108 36 45 13.5684 $w=3.73e-07 $l=1.05e-07 $layer=POLY_cond $X=3.63 $Y=1.557
+ $X2=3.735 $Y2=1.557
r109 36 43 40.7051 $w=3.73e-07 $l=3.15e-07 $layer=POLY_cond $X=3.63 $Y=1.557
+ $X2=3.315 $Y2=1.557
r110 35 36 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.63
+ $Y=1.515 $X2=3.63 $Y2=1.515
r111 33 41 12.7116 $w=2.48e-07 $l=2.5e-07 $layer=LI1_cond $X=3.375 $Y=1.555
+ $X2=3.125 $Y2=1.555
r112 33 35 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=3.375 $Y=1.555
+ $X2=3.63 $Y2=1.555
r113 32 41 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=2.515 $Y=1.515
+ $X2=3.125 $Y2=1.515
r114 30 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.43 $Y=1.43
+ $X2=2.515 $Y2=1.515
r115 29 30 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.43 $Y=1.18
+ $X2=2.43 $Y2=1.43
r116 28 39 15.1197 $w=4.68e-07 $l=7.03378e-07 $layer=LI1_cond $X=1.675 $Y=1.095
+ $X2=1.402 $Y2=0.515
r117 27 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.345 $Y=1.095
+ $X2=2.43 $Y2=1.18
r118 27 28 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.345 $Y=1.095
+ $X2=1.675 $Y2=1.095
r119 25 28 7.42701 $w=4.68e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.59 $Y=1.18
+ $X2=1.675 $Y2=1.095
r120 25 26 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=1.59 $Y=1.18
+ $X2=1.59 $Y2=1.82
r121 21 26 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.505 $Y=1.945
+ $X2=1.59 $Y2=1.82
r122 21 23 4.84026 $w=2.48e-07 $l=1.05e-07 $layer=LI1_cond $X=1.505 $Y=1.945
+ $X2=1.4 $Y2=1.945
r123 17 46 24.162 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.745 $Y=1.35
+ $X2=3.745 $Y2=1.557
r124 17 19 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.745 $Y=1.35
+ $X2=3.745 $Y2=0.74
r125 14 45 24.162 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.735 $Y=1.765
+ $X2=3.735 $Y2=1.557
r126 14 16 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.735 $Y=1.765
+ $X2=3.735 $Y2=2.4
r127 10 43 24.162 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.315 $Y=1.35
+ $X2=3.315 $Y2=1.557
r128 10 12 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.315 $Y=1.35
+ $X2=3.315 $Y2=0.74
r129 7 42 24.162 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.285 $Y=1.765
+ $X2=3.285 $Y2=1.557
r130 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.285 $Y=1.765
+ $X2=3.285 $Y2=2.4
r131 2 23 600 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=1 $X=1.2
+ $Y=1.84 $X2=1.4 $Y2=1.985
r132 1 39 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.155
+ $Y=0.37 $X2=1.295 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__NAND4BB_2%C 1 3 6 8 10 13 15 16 23 24
r57 23 25 9.11892 $w=3.7e-07 $l=7e-08 $layer=POLY_cond $X=5.22 $Y=1.557 $X2=5.29
+ $Y2=1.557
r58 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.22
+ $Y=1.515 $X2=5.22 $Y2=1.515
r59 21 23 7.16487 $w=3.7e-07 $l=5.5e-08 $layer=POLY_cond $X=5.165 $Y=1.557
+ $X2=5.22 $Y2=1.557
r60 20 21 48.8514 $w=3.7e-07 $l=3.75e-07 $layer=POLY_cond $X=4.79 $Y=1.557
+ $X2=5.165 $Y2=1.557
r61 19 20 9.77027 $w=3.7e-07 $l=7.5e-08 $layer=POLY_cond $X=4.715 $Y=1.557
+ $X2=4.79 $Y2=1.557
r62 16 24 4.82418 $w=4.28e-07 $l=1.8e-07 $layer=LI1_cond $X=5.04 $Y=1.565
+ $X2=5.22 $Y2=1.565
r63 15 16 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=4.56 $Y=1.565
+ $X2=5.04 $Y2=1.565
r64 11 25 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.29 $Y=1.35
+ $X2=5.29 $Y2=1.557
r65 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.29 $Y=1.35
+ $X2=5.29 $Y2=0.74
r66 8 21 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=5.165 $Y=1.765
+ $X2=5.165 $Y2=1.557
r67 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.165 $Y=1.765
+ $X2=5.165 $Y2=2.4
r68 4 20 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.79 $Y=1.35
+ $X2=4.79 $Y2=1.557
r69 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.79 $Y=1.35 $X2=4.79
+ $Y2=0.74
r70 1 19 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=4.715 $Y=1.765
+ $X2=4.715 $Y2=1.557
r71 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.715 $Y=1.765
+ $X2=4.715 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__NAND4BB_2%D 1 3 6 8 10 13 20 25 28
c51 6 0 1.4333e-19 $X=5.72 $Y=0.74
r52 25 26 1.928 $w=3.75e-07 $l=1.5e-08 $layer=POLY_cond $X=6.205 $Y=1.557
+ $X2=6.22 $Y2=1.557
r53 22 23 0.642667 $w=3.75e-07 $l=5e-09 $layer=POLY_cond $X=5.715 $Y=1.557
+ $X2=5.72 $Y2=1.557
r54 20 28 3.73456 $w=4.28e-07 $l=1.15e-07 $layer=LI1_cond $X=6.48 $Y=1.565
+ $X2=6.365 $Y2=1.565
r55 18 25 9.64 $w=3.75e-07 $l=7.5e-08 $layer=POLY_cond $X=6.13 $Y=1.557
+ $X2=6.205 $Y2=1.557
r56 18 23 52.6987 $w=3.75e-07 $l=4.1e-07 $layer=POLY_cond $X=6.13 $Y=1.557
+ $X2=5.72 $Y2=1.557
r57 17 28 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=6.13 $Y=1.515
+ $X2=6.365 $Y2=1.515
r58 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.13
+ $Y=1.515 $X2=6.13 $Y2=1.515
r59 11 26 24.2915 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.22 $Y=1.35
+ $X2=6.22 $Y2=1.557
r60 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.22 $Y=1.35
+ $X2=6.22 $Y2=0.74
r61 8 25 24.2915 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=6.205 $Y=1.765
+ $X2=6.205 $Y2=1.557
r62 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.205 $Y=1.765
+ $X2=6.205 $Y2=2.4
r63 4 23 24.2915 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.72 $Y=1.35
+ $X2=5.72 $Y2=1.557
r64 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.72 $Y=1.35 $X2=5.72
+ $Y2=0.74
r65 1 22 24.2915 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=5.715 $Y=1.765
+ $X2=5.715 $Y2=1.557
r66 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.715 $Y=1.765
+ $X2=5.715 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__NAND4BB_2%VPWR 1 2 3 4 5 6 23 27 31 35 39 41 43 48
+ 49 51 52 53 62 66 71 77 80 83 87
r88 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r89 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r90 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r91 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r92 75 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r93 75 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=5.52
+ $Y2=3.33
r94 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r95 72 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.605 $Y=3.33
+ $X2=5.44 $Y2=3.33
r96 72 74 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=5.605 $Y=3.33 $X2=6
+ $Y2=3.33
r97 71 86 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=6.275 $Y=3.33
+ $X2=6.497 $Y2=3.33
r98 71 74 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.275 $Y=3.33 $X2=6
+ $Y2=3.33
r99 70 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r100 70 81 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.08 $Y2=3.33
r101 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r102 67 80 14.259 $w=1.7e-07 $l=3.8e-07 $layer=LI1_cond $X=4.605 $Y=3.33
+ $X2=4.225 $Y2=3.33
r103 67 69 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=4.605 $Y=3.33
+ $X2=5.04 $Y2=3.33
r104 66 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.275 $Y=3.33
+ $X2=5.44 $Y2=3.33
r105 66 69 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=5.275 $Y=3.33
+ $X2=5.04 $Y2=3.33
r106 65 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r107 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r108 62 80 14.259 $w=1.7e-07 $l=3.8e-07 $layer=LI1_cond $X=3.845 $Y=3.33
+ $X2=4.225 $Y2=3.33
r109 62 64 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=3.845 $Y=3.33
+ $X2=3.6 $Y2=3.33
r110 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r111 58 61 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r112 58 78 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r113 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r114 55 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.98 $Y=3.33
+ $X2=0.815 $Y2=3.33
r115 55 57 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=0.98 $Y=3.33 $X2=1.68
+ $Y2=3.33
r116 53 65 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=3.6 $Y2=3.33
r117 53 61 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=2.64 $Y2=3.33
r118 51 60 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=2.845 $Y=3.33
+ $X2=2.64 $Y2=3.33
r119 51 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.845 $Y=3.33
+ $X2=3.01 $Y2=3.33
r120 50 64 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=3.175 $Y=3.33
+ $X2=3.6 $Y2=3.33
r121 50 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.175 $Y=3.33
+ $X2=3.01 $Y2=3.33
r122 48 57 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.845 $Y=3.33
+ $X2=1.68 $Y2=3.33
r123 48 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.845 $Y=3.33
+ $X2=2.01 $Y2=3.33
r124 47 60 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=2.175 $Y=3.33
+ $X2=2.64 $Y2=3.33
r125 47 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.175 $Y=3.33
+ $X2=2.01 $Y2=3.33
r126 43 46 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=6.44 $Y=2.115
+ $X2=6.44 $Y2=2.815
r127 41 86 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=6.44 $Y=3.245
+ $X2=6.497 $Y2=3.33
r128 41 46 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=6.44 $Y=3.245
+ $X2=6.44 $Y2=2.815
r129 37 83 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.44 $Y=3.245
+ $X2=5.44 $Y2=3.33
r130 37 39 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=5.44 $Y=3.245
+ $X2=5.44 $Y2=2.455
r131 33 80 3.03114 $w=7.6e-07 $l=8.5e-08 $layer=LI1_cond $X=4.225 $Y=3.245
+ $X2=4.225 $Y2=3.33
r132 33 35 12.4329 $w=7.58e-07 $l=7.9e-07 $layer=LI1_cond $X=4.225 $Y=3.245
+ $X2=4.225 $Y2=2.455
r133 29 52 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.01 $Y=3.245
+ $X2=3.01 $Y2=3.33
r134 29 31 31.081 $w=3.28e-07 $l=8.9e-07 $layer=LI1_cond $X=3.01 $Y=3.245
+ $X2=3.01 $Y2=2.355
r135 25 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.01 $Y=3.245
+ $X2=2.01 $Y2=3.33
r136 25 27 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=2.01 $Y=3.245
+ $X2=2.01 $Y2=2.78
r137 21 77 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=3.245
+ $X2=0.815 $Y2=3.33
r138 21 23 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=0.815 $Y=3.245
+ $X2=0.815 $Y2=2.745
r139 6 46 400 $w=1.7e-07 $l=1.05196e-06 $layer=licon1_PDIFF $count=1 $X=6.28
+ $Y=1.84 $X2=6.44 $Y2=2.815
r140 6 43 400 $w=1.7e-07 $l=3.45868e-07 $layer=licon1_PDIFF $count=1 $X=6.28
+ $Y=1.84 $X2=6.44 $Y2=2.115
r141 5 39 300 $w=1.7e-07 $l=7.07972e-07 $layer=licon1_PDIFF $count=2 $X=5.24
+ $Y=1.84 $X2=5.44 $Y2=2.455
r142 4 35 150 $w=1.7e-07 $l=9.38403e-07 $layer=licon1_PDIFF $count=4 $X=3.81
+ $Y=1.84 $X2=4.49 $Y2=2.455
r143 3 31 300 $w=1.7e-07 $l=6.06815e-07 $layer=licon1_PDIFF $count=2 $X=2.81
+ $Y=1.84 $X2=3.01 $Y2=2.355
r144 2 27 600 $w=1.7e-07 $l=1.0099e-06 $layer=licon1_PDIFF $count=1 $X=1.865
+ $Y=1.84 $X2=2.01 $Y2=2.78
r145 1 23 600 $w=1.7e-07 $l=1.01573e-06 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.84 $X2=0.815 $Y2=2.745
.ends

.subckt PM_SKY130_FD_SC_LS__NAND4BB_2%Y 1 2 3 4 5 16 20 22 24 27 28 29 32 34 36
+ 40 42 44 46 51 53 55 58 61 63
c121 29 0 8.19262e-20 $X=2.855 $Y=1.175
c122 20 0 1.36243e-19 $X=2.51 $Y=2.02
r123 61 63 1.75372 $w=2.28e-07 $l=3.5e-08 $layer=LI1_cond $X=4.08 $Y=1.26
+ $X2=4.08 $Y2=1.295
r124 58 61 2.9826 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.08 $Y=1.175
+ $X2=4.08 $Y2=1.26
r125 58 63 1.25266 $w=2.28e-07 $l=2.5e-08 $layer=LI1_cond $X=4.08 $Y=1.32
+ $X2=4.08 $Y2=1.295
r126 52 58 26.5563 $w=2.28e-07 $l=5.3e-07 $layer=LI1_cond $X=4.08 $Y=1.85
+ $X2=4.08 $Y2=1.32
r127 52 53 1.18299 $w=2.3e-07 $l=1.35e-07 $layer=LI1_cond $X=4.08 $Y=1.85
+ $X2=4.08 $Y2=1.985
r128 44 57 2.99552 $w=3.3e-07 $l=1.35e-07 $layer=LI1_cond $X=5.94 $Y=2.12
+ $X2=5.94 $Y2=1.985
r129 44 46 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=5.94 $Y=2.12
+ $X2=5.94 $Y2=2.815
r130 43 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.105 $Y=2.035
+ $X2=4.94 $Y2=2.035
r131 42 57 4.77065 $w=1.7e-07 $l=1.88348e-07 $layer=LI1_cond $X=5.775 $Y=2.035
+ $X2=5.94 $Y2=1.985
r132 42 43 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.775 $Y=2.035
+ $X2=5.105 $Y2=2.035
r133 38 55 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.94 $Y=2.12
+ $X2=4.94 $Y2=2.035
r134 38 40 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=4.94 $Y=2.12
+ $X2=4.94 $Y2=2.815
r135 37 53 5.35987 $w=2.2e-07 $l=1.3775e-07 $layer=LI1_cond $X=4.195 $Y=2.035
+ $X2=4.08 $Y2=1.985
r136 36 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.775 $Y=2.035
+ $X2=4.94 $Y2=2.035
r137 36 37 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=4.775 $Y=2.035
+ $X2=4.195 $Y2=2.035
r138 35 51 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=3.675 $Y=1.985
+ $X2=3.51 $Y2=1.985
r139 34 53 5.35987 $w=2.2e-07 $l=1.15e-07 $layer=LI1_cond $X=3.965 $Y=1.985
+ $X2=4.08 $Y2=1.985
r140 34 35 12.3781 $w=2.68e-07 $l=2.9e-07 $layer=LI1_cond $X=3.965 $Y=1.985
+ $X2=3.675 $Y2=1.985
r141 30 51 0.067832 $w=3.3e-07 $l=1.35e-07 $layer=LI1_cond $X=3.51 $Y=2.12
+ $X2=3.51 $Y2=1.985
r142 30 32 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=3.51 $Y=2.12
+ $X2=3.51 $Y2=2.815
r143 28 58 4.03528 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=3.965 $Y=1.175
+ $X2=4.08 $Y2=1.175
r144 28 29 72.4171 $w=1.68e-07 $l=1.11e-06 $layer=LI1_cond $X=3.965 $Y=1.175
+ $X2=2.855 $Y2=1.175
r145 27 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.77 $Y=1.09
+ $X2=2.855 $Y2=1.175
r146 26 27 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.77 $Y=0.84
+ $X2=2.77 $Y2=1.09
r147 25 49 4.99254 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=2.675 $Y=1.935
+ $X2=2.51 $Y2=1.92
r148 24 51 7.13466 $w=2.2e-07 $l=1.88348e-07 $layer=LI1_cond $X=3.345 $Y=1.935
+ $X2=3.51 $Y2=1.985
r149 24 25 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.345 $Y=1.935
+ $X2=2.675 $Y2=1.935
r150 20 49 2.77363 $w=3.3e-07 $l=1e-07 $layer=LI1_cond $X=2.51 $Y=2.02 $X2=2.51
+ $Y2=1.92
r151 20 22 27.7634 $w=3.28e-07 $l=7.95e-07 $layer=LI1_cond $X=2.51 $Y=2.02
+ $X2=2.51 $Y2=2.815
r152 16 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.685 $Y=0.755
+ $X2=2.77 $Y2=0.84
r153 16 18 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.685 $Y=0.755
+ $X2=2.51 $Y2=0.755
r154 5 57 400 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=1 $X=5.79
+ $Y=1.84 $X2=5.94 $Y2=2.015
r155 5 46 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=5.79
+ $Y=1.84 $X2=5.94 $Y2=2.815
r156 4 55 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=4.79
+ $Y=1.84 $X2=4.94 $Y2=2.115
r157 4 40 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=4.79
+ $Y=1.84 $X2=4.94 $Y2=2.815
r158 3 51 400 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=1 $X=3.36
+ $Y=1.84 $X2=3.51 $Y2=2.015
r159 3 32 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=3.36
+ $Y=1.84 $X2=3.51 $Y2=2.815
r160 2 49 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.36
+ $Y=1.84 $X2=2.51 $Y2=1.985
r161 2 22 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.36
+ $Y=1.84 $X2=2.51 $Y2=2.815
r162 1 18 182 $w=1.7e-07 $l=4.60163e-07 $layer=licon1_NDIFF $count=1 $X=2.345
+ $Y=0.37 $X2=2.51 $Y2=0.755
.ends

.subckt PM_SKY130_FD_SC_LS__NAND4BB_2%VGND 1 2 9 13 15 17 22 32 33 36 39
r59 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r60 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r61 33 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r62 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r63 30 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.17 $Y=0 $X2=6.005
+ $Y2=0
r64 30 32 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=6.17 $Y=0 $X2=6.48
+ $Y2=0
r65 29 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r66 28 29 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r67 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r68 25 28 281.84 $w=1.68e-07 $l=4.32e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=5.52
+ $Y2=0
r69 25 26 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r70 23 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.96 $Y=0 $X2=0.795
+ $Y2=0
r71 23 25 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=0.96 $Y=0 $X2=1.2
+ $Y2=0
r72 22 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.84 $Y=0 $X2=6.005
+ $Y2=0
r73 22 28 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=5.84 $Y=0 $X2=5.52
+ $Y2=0
r74 20 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r75 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r76 17 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.63 $Y=0 $X2=0.795
+ $Y2=0
r77 17 19 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=0.63 $Y=0 $X2=0.24
+ $Y2=0
r78 15 29 0.602067 $w=4.9e-07 $l=2.16e-06 $layer=MET1_cond $X=3.36 $Y=0 $X2=5.52
+ $Y2=0
r79 15 26 0.602067 $w=4.9e-07 $l=2.16e-06 $layer=MET1_cond $X=3.36 $Y=0 $X2=1.2
+ $Y2=0
r80 11 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.005 $Y=0.085
+ $X2=6.005 $Y2=0
r81 11 13 19.7312 $w=3.28e-07 $l=5.65e-07 $layer=LI1_cond $X=6.005 $Y=0.085
+ $X2=6.005 $Y2=0.65
r82 7 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.795 $Y=0.085
+ $X2=0.795 $Y2=0
r83 7 9 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.795 $Y=0.085
+ $X2=0.795 $Y2=0.515
r84 2 13 182 $w=1.7e-07 $l=3.70405e-07 $layer=licon1_NDIFF $count=1 $X=5.795
+ $Y=0.37 $X2=6.005 $Y2=0.65
r85 1 9 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=0.585
+ $Y=0.37 $X2=0.795 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__NAND4BB_2%A_373_74# 1 2 3 12 14 15 19 20 22
r38 20 22 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=3.195 $Y=0.835
+ $X2=3.985 $Y2=0.835
r39 19 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.11 $Y=0.75
+ $X2=3.195 $Y2=0.835
r40 18 19 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.11 $Y=0.5 $X2=3.11
+ $Y2=0.75
r41 15 17 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=2.175 $Y=0.415
+ $X2=3.02 $Y2=0.415
r42 14 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.025 $Y=0.415
+ $X2=3.11 $Y2=0.5
r43 14 17 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=3.025 $Y=0.415
+ $X2=3.02 $Y2=0.415
r44 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.01 $Y=0.5
+ $X2=2.175 $Y2=0.415
r45 10 12 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=2.01 $Y=0.5 $X2=2.01
+ $Y2=0.595
r46 3 22 182 $w=1.7e-07 $l=5.41249e-07 $layer=licon1_NDIFF $count=1 $X=3.82
+ $Y=0.37 $X2=3.985 $Y2=0.835
r47 2 17 182 $w=1.7e-07 $l=2.41454e-07 $layer=licon1_NDIFF $count=1 $X=2.8
+ $Y=0.37 $X2=3.02 $Y2=0.415
r48 1 12 182 $w=1.7e-07 $l=2.88531e-07 $layer=licon1_NDIFF $count=1 $X=1.865
+ $Y=0.37 $X2=2.01 $Y2=0.595
.ends

.subckt PM_SKY130_FD_SC_LS__NAND4BB_2%A_678_74# 1 2 7 11 13
c28 11 0 1.4333e-19 $X=5.075 $Y=0.65
c29 7 0 6.95413e-20 $X=4.91 $Y=0.34
r30 13 16 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=3.53 $Y=0.34
+ $X2=3.53 $Y2=0.495
r31 9 11 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=5.075 $Y=0.425
+ $X2=5.075 $Y2=0.65
r32 8 13 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.695 $Y=0.34
+ $X2=3.53 $Y2=0.34
r33 7 9 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.91 $Y=0.34
+ $X2=5.075 $Y2=0.425
r34 7 8 79.2674 $w=1.68e-07 $l=1.215e-06 $layer=LI1_cond $X=4.91 $Y=0.34
+ $X2=3.695 $Y2=0.34
r35 2 11 182 $w=1.7e-07 $l=3.70405e-07 $layer=licon1_NDIFF $count=1 $X=4.865
+ $Y=0.37 $X2=5.075 $Y2=0.65
r36 1 16 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=3.39
+ $Y=0.37 $X2=3.53 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LS__NAND4BB_2%A_886_74# 1 2 3 12 14 15 18 20 24 26
r45 22 24 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=6.475 $Y=1.01
+ $X2=6.475 $Y2=0.515
r46 21 26 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.67 $Y=1.095
+ $X2=5.545 $Y2=1.095
r47 20 22 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.35 $Y=1.095
+ $X2=6.475 $Y2=1.01
r48 20 21 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=6.35 $Y=1.095
+ $X2=5.67 $Y2=1.095
r49 16 26 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.545 $Y=1.01
+ $X2=5.545 $Y2=1.095
r50 16 18 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=5.545 $Y=1.01
+ $X2=5.545 $Y2=0.515
r51 14 26 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.42 $Y=1.095
+ $X2=5.545 $Y2=1.095
r52 14 15 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=5.42 $Y=1.095
+ $X2=4.74 $Y2=1.095
r53 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.575 $Y=1.01
+ $X2=4.74 $Y2=1.095
r54 10 12 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=4.575 $Y=1.01
+ $X2=4.575 $Y2=0.785
r55 3 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.295
+ $Y=0.37 $X2=6.435 $Y2=0.515
r56 2 18 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.365
+ $Y=0.37 $X2=5.505 $Y2=0.515
r57 1 12 182 $w=1.7e-07 $l=4.82079e-07 $layer=licon1_NDIFF $count=1 $X=4.43
+ $Y=0.37 $X2=4.575 $Y2=0.785
.ends

