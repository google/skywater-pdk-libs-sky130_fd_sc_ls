* NGSPICE file created from sky130_fd_sc_ls__or3b_2.ext - technology: sky130A

.subckt sky130_fd_sc_ls__or3b_2 A B C_N VGND VNB VPB VPWR X
M1000 VPWR a_190_260# X VPB phighvt w=1.12e+06u l=150000u
+  ad=1.04315e+12p pd=6.42e+06u as=3.36e+11p ps=2.84e+06u
M1001 a_458_368# A VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1002 a_190_260# a_27_368# a_542_368# VPB phighvt w=1e+06u l=150000u
+  ad=2.95e+11p pd=2.59e+06u as=3.9e+11p ps=2.78e+06u
M1003 X a_190_260# VGND VNB nshort w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=9.1395e+11p ps=6.95e+06u
M1004 VGND C_N a_27_368# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1005 VGND B a_190_260# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=4.064e+11p ps=3.83e+06u
M1006 a_190_260# A VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR C_N a_27_368# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=2.478e+11p ps=2.27e+06u
M1008 VGND a_190_260# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 X a_190_260# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_542_368# B a_458_368# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_190_260# a_27_368# VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

