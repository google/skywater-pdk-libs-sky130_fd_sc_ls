* File: sky130_fd_sc_ls__a211oi_1.pex.spice
* Created: Fri Aug 28 12:49:29 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__A211OI_1%A2 1 3 6 8 12
r26 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.63
+ $Y=1.515 $X2=0.63 $Y2=1.515
r27 8 12 4.67207 $w=3.68e-07 $l=1.5e-07 $layer=LI1_cond $X=0.65 $Y=1.665
+ $X2=0.65 $Y2=1.515
r28 4 11 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=0.72 $Y=1.35
+ $X2=0.63 $Y2=1.515
r29 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.72 $Y=1.35 $X2=0.72
+ $Y2=0.74
r30 1 11 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=0.705 $Y=1.765
+ $X2=0.63 $Y2=1.515
r31 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.705 $Y=1.765
+ $X2=0.705 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__A211OI_1%A1 3 5 7 8 12
r32 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.17
+ $Y=1.515 $X2=1.17 $Y2=1.515
r33 8 12 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.17 $Y=1.665
+ $X2=1.17 $Y2=1.515
r34 5 11 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=1.245 $Y=1.765
+ $X2=1.17 $Y2=1.515
r35 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.245 $Y=1.765
+ $X2=1.245 $Y2=2.4
r36 1 11 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=1.08 $Y=1.35
+ $X2=1.17 $Y2=1.515
r37 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.08 $Y=1.35 $X2=1.08
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__A211OI_1%B1 3 5 7 8 12
c30 12 0 4.72069e-20 $X=1.71 $Y=1.515
r31 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.71
+ $Y=1.515 $X2=1.71 $Y2=1.515
r32 8 12 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.71 $Y=1.665
+ $X2=1.71 $Y2=1.515
r33 5 11 52.2586 $w=2.99e-07 $l=2.57391e-07 $layer=POLY_cond $X=1.695 $Y=1.765
+ $X2=1.71 $Y2=1.515
r34 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.695 $Y=1.765
+ $X2=1.695 $Y2=2.4
r35 1 11 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=1.62 $Y=1.35
+ $X2=1.71 $Y2=1.515
r36 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.62 $Y=1.35 $X2=1.62
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__A211OI_1%C1 3 4 6 8 9 10 13
c29 4 0 2.15901e-19 $X=2.175 $Y=1.765
r30 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.61
+ $Y=1.385 $X2=2.61 $Y2=1.385
r31 10 14 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=2.61 $Y=1.295 $X2=2.61
+ $Y2=1.385
r32 8 13 60.3271 $w=3.3e-07 $l=3.45e-07 $layer=POLY_cond $X=2.265 $Y=1.385
+ $X2=2.61 $Y2=1.385
r33 8 9 66.2869 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.175 $Y=1.385
+ $X2=2.175 $Y2=1.22
r34 4 8 149.859 $w=1.8e-07 $l=3.8e-07 $layer=POLY_cond $X=2.175 $Y=1.765
+ $X2=2.175 $Y2=1.385
r35 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.175 $Y=1.765
+ $X2=2.175 $Y2=2.4
r36 3 9 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.16 $Y=0.74 $X2=2.16
+ $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_LS__A211OI_1%A_71_368# 1 2 7 9 11 13 15
c28 13 0 1.68694e-19 $X=1.47 $Y=2.12
r29 13 20 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.47 $Y=2.12 $X2=1.47
+ $Y2=2.035
r30 13 15 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=1.47 $Y=2.12
+ $X2=1.47 $Y2=2.815
r31 12 18 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.645 $Y=2.035
+ $X2=0.48 $Y2=2.035
r32 11 20 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.305 $Y=2.035
+ $X2=1.47 $Y2=2.035
r33 11 12 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=1.305 $Y=2.035
+ $X2=0.645 $Y2=2.035
r34 7 18 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.48 $Y=2.12 $X2=0.48
+ $Y2=2.035
r35 7 9 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=0.48 $Y=2.12 $X2=0.48
+ $Y2=2.815
r36 2 20 400 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=1.32
+ $Y=1.84 $X2=1.47 $Y2=2.035
r37 2 15 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.32
+ $Y=1.84 $X2=1.47 $Y2=2.815
r38 1 18 400 $w=1.7e-07 $l=2.498e-07 $layer=licon1_PDIFF $count=1 $X=0.355
+ $Y=1.84 $X2=0.48 $Y2=2.035
r39 1 9 400 $w=1.7e-07 $l=1.03562e-06 $layer=licon1_PDIFF $count=1 $X=0.355
+ $Y=1.84 $X2=0.48 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_LS__A211OI_1%VPWR 1 6 9 10 11 21 22
r26 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r27 18 21 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r28 18 19 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r29 15 19 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r30 14 15 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r31 11 22 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=2.64 $Y2=3.33
r32 11 19 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.2 $Y2=3.33
r33 9 14 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=0.815 $Y=3.33
+ $X2=0.72 $Y2=3.33
r34 9 10 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=0.815 $Y=3.33
+ $X2=0.975 $Y2=3.33
r35 8 18 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=1.135 $Y=3.33 $X2=1.2
+ $Y2=3.33
r36 8 10 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=1.135 $Y=3.33
+ $X2=0.975 $Y2=3.33
r37 4 10 0.800721 $w=3.2e-07 $l=8.5e-08 $layer=LI1_cond $X=0.975 $Y=3.245
+ $X2=0.975 $Y2=3.33
r38 4 6 28.4509 $w=3.18e-07 $l=7.9e-07 $layer=LI1_cond $X=0.975 $Y=3.245
+ $X2=0.975 $Y2=2.455
r39 1 6 300 $w=1.7e-07 $l=6.9482e-07 $layer=licon1_PDIFF $count=2 $X=0.78
+ $Y=1.84 $X2=0.95 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_LS__A211OI_1%Y 1 2 3 10 12 18 22 25 26 27 28 29 33
r51 29 33 0.0230313 $w=3.7e-07 $l=1.85e-07 $layer=LI1_cond $X=2.045 $Y=0.81
+ $X2=2.045 $Y2=0.995
r52 28 33 11.3687 $w=3.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.68 $Y=0.995
+ $X2=2.045 $Y2=0.995
r53 28 34 5.60648 $w=3.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.68 $Y=0.995
+ $X2=1.5 $Y2=0.995
r54 27 34 3.62315 $w=3.7e-07 $l=2.08e-07 $layer=LI1_cond $X=1.292 $Y=0.995
+ $X2=1.5 $Y2=0.995
r55 25 26 9.6413 $w=5.18e-07 $l=1.65e-07 $layer=LI1_cond $X=2.305 $Y=1.985
+ $X2=2.305 $Y2=1.82
r56 20 29 7.06239 $w=2.5e-07 $l=3.3e-07 $layer=LI1_cond $X=2.375 $Y=0.81
+ $X2=2.045 $Y2=0.81
r57 20 22 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.375 $Y=0.81
+ $X2=2.375 $Y2=0.515
r58 16 25 2.18514 $w=5.18e-07 $l=9.5e-08 $layer=LI1_cond $X=2.305 $Y=2.08
+ $X2=2.305 $Y2=1.985
r59 16 18 16.9061 $w=5.18e-07 $l=7.35e-07 $layer=LI1_cond $X=2.305 $Y=2.08
+ $X2=2.305 $Y2=2.815
r60 14 29 7.06239 $w=2.5e-07 $l=4.10305e-07 $layer=LI1_cond $X=2.13 $Y=1.18
+ $X2=2.045 $Y2=0.81
r61 14 26 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=2.13 $Y=1.18 $X2=2.13
+ $Y2=1.82
r62 10 27 3.22252 $w=4.15e-07 $l=1.85e-07 $layer=LI1_cond $X=1.292 $Y=0.81
+ $X2=1.292 $Y2=0.995
r63 10 12 8.19206 $w=4.13e-07 $l=2.95e-07 $layer=LI1_cond $X=1.292 $Y=0.81
+ $X2=1.292 $Y2=0.515
r64 3 25 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.25
+ $Y=1.84 $X2=2.4 $Y2=1.985
r65 3 18 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.25
+ $Y=1.84 $X2=2.4 $Y2=2.815
r66 2 22 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.235
+ $Y=0.37 $X2=2.375 $Y2=0.515
r67 1 27 182 $w=1.7e-07 $l=6.70242e-07 $layer=licon1_NDIFF $count=1 $X=1.155
+ $Y=0.37 $X2=1.315 $Y2=0.965
r68 1 12 182 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=1 $X=1.155
+ $Y=0.37 $X2=1.315 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__A211OI_1%VGND 1 2 9 13 16 17 18 24 30 31 34
r35 34 35 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r36 31 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=1.68
+ $Y2=0
r37 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r38 28 34 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=2.04 $Y=0 $X2=1.855
+ $Y2=0
r39 28 30 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=2.04 $Y=0 $X2=2.64
+ $Y2=0
r40 26 27 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r41 24 34 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=1.67 $Y=0 $X2=1.855
+ $Y2=0
r42 24 26 61.9786 $w=1.68e-07 $l=9.5e-07 $layer=LI1_cond $X=1.67 $Y=0 $X2=0.72
+ $Y2=0
r43 22 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r44 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r45 18 35 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.68
+ $Y2=0
r46 18 27 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=0.72
+ $Y2=0
r47 16 21 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=0.34 $Y=0 $X2=0.24
+ $Y2=0
r48 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.34 $Y=0 $X2=0.505
+ $Y2=0
r49 15 26 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=0.67 $Y=0 $X2=0.72
+ $Y2=0
r50 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.67 $Y=0 $X2=0.505
+ $Y2=0
r51 11 34 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.855 $Y=0.085
+ $X2=1.855 $Y2=0
r52 11 13 14.0162 $w=3.68e-07 $l=4.5e-07 $layer=LI1_cond $X=1.855 $Y=0.085
+ $X2=1.855 $Y2=0.535
r53 7 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.505 $Y=0.085
+ $X2=0.505 $Y2=0
r54 7 9 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.505 $Y=0.085
+ $X2=0.505 $Y2=0.515
r55 2 13 182 $w=1.7e-07 $l=2.31571e-07 $layer=licon1_NDIFF $count=1 $X=1.695
+ $Y=0.37 $X2=1.855 $Y2=0.535
r56 1 9 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.38
+ $Y=0.37 $X2=0.505 $Y2=0.515
.ends

