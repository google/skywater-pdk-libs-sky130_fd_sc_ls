* File: sky130_fd_sc_ls__nor4b_2.spice
* Created: Wed Sep  2 11:15:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__nor4b_2.pex.spice"
.subckt sky130_fd_sc_ls__nor4b_2  VNB VPB D_N C B A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* B	B
* C	C
* D_N	D_N
* VPB	VPB
* VNB	VNB
MM1017 N_VGND_M1017_d N_D_N_M1017_g N_A_27_392#_M1017_s VNB NSHORT L=0.15 W=0.64
+ AD=0.136255 AS=0.1824 PD=1.07594 PS=1.85 NRD=13.116 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75004.8 A=0.096 P=1.58 MULT=1
MM1004 N_VGND_M1017_d N_A_27_392#_M1004_g N_Y_M1004_s VNB NSHORT L=0.15 W=0.74
+ AD=0.157545 AS=0.1295 PD=1.24406 PS=1.09 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75000.7 SB=75004.3 A=0.111 P=1.78 MULT=1
MM1006 N_VGND_M1006_d N_A_27_392#_M1006_g N_Y_M1004_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1998 AS=0.1295 PD=1.28 PS=1.09 NRD=15.396 NRS=11.34 M=1 R=4.93333
+ SA=75001.2 SB=75003.8 A=0.111 P=1.78 MULT=1
MM1007 N_VGND_M1006_d N_C_M1007_g N_Y_M1007_s VNB NSHORT L=0.15 W=0.74 AD=0.1998
+ AS=0.1036 PD=1.28 PS=1.02 NRD=26.748 NRS=0 M=1 R=4.93333 SA=75001.9 SB=75003.1
+ A=0.111 P=1.78 MULT=1
MM1016 N_VGND_M1016_d N_C_M1016_g N_Y_M1007_s VNB NSHORT L=0.15 W=0.74 AD=0.148
+ AS=0.1036 PD=1.14 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75002.3 SB=75002.7
+ A=0.111 P=1.78 MULT=1
MM1001 N_Y_M1001_d N_B_M1001_g N_VGND_M1016_d VNB NSHORT L=0.15 W=0.74 AD=0.1369
+ AS=0.148 PD=1.11 PS=1.14 NRD=3.24 NRS=8.1 M=1 R=4.93333 SA=75002.9 SB=75002.1
+ A=0.111 P=1.78 MULT=1
MM1009 N_Y_M1001_d N_B_M1009_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.74 AD=0.1369
+ AS=0.26825 PD=1.11 PS=1.465 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75003.4
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1003 N_VGND_M1009_s N_A_M1003_g N_Y_M1003_s VNB NSHORT L=0.15 W=0.74
+ AD=0.26825 AS=0.12395 PD=1.465 PS=1.075 NRD=0 NRS=0 M=1 R=4.93333 SA=75004.3
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1011 N_VGND_M1011_d N_A_M1011_g N_Y_M1003_s VNB NSHORT L=0.15 W=0.74 AD=0.222
+ AS=0.12395 PD=2.08 PS=1.075 NRD=2.424 NRS=8.916 M=1 R=4.93333 SA=75004.7
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1013 N_VPWR_M1013_d N_D_N_M1013_g N_A_27_392#_M1013_s VPB PHIGHVT L=0.15 W=1
+ AD=0.295 AS=0.295 PD=2.59 PS=2.59 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1008 N_Y_M1008_d N_A_27_392#_M1008_g N_A_229_368#_M1008_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1014 N_Y_M1008_d N_A_27_392#_M1014_g N_A_229_368#_M1014_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1000 N_A_498_368#_M1000_d N_C_M1000_g N_A_229_368#_M1014_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1002 N_A_498_368#_M1000_d N_C_M1002_g N_A_229_368#_M1002_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.6 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1005 N_A_498_368#_M1005_d N_B_M1005_g N_A_701_368#_M1005_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1010 N_A_498_368#_M1005_d N_B_M1010_g N_A_701_368#_M1010_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1012 N_A_701_368#_M1010_s N_A_M1012_g N_VPWR_M1012_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.1736 PD=1.42 PS=1.43 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1015 N_A_701_368#_M1015_d N_A_M1015_g N_VPWR_M1012_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.1736 PD=2.83 PS=1.43 NRD=1.7533 NRS=3.5066 M=1 R=7.46667
+ SA=75001.6 SB=75000.2 A=0.168 P=2.54 MULT=1
DX18_noxref VNB VPB NWDIODE A=11.4204 P=16
*
.include "sky130_fd_sc_ls__nor4b_2.pxi.spice"
*
.ends
*
*
