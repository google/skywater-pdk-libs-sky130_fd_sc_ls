# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ls__ebufn_8
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ls__ebufn_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.56000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.645000 1.180000 9.975000 1.550000 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  1.623000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.265000 1.180000 9.475000 1.550000 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  2.360500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545000 0.595000 0.875000 0.980000 ;
        RECT 0.545000 0.980000 3.760000 1.150000 ;
        RECT 0.545000 1.150000 0.835000 1.820000 ;
        RECT 0.545000 1.820000 3.700000 1.990000 ;
        RECT 0.545000 1.990000 0.900000 2.735000 ;
        RECT 1.430000 0.595000 1.760000 0.980000 ;
        RECT 1.520000 1.990000 1.850000 2.735000 ;
        RECT 2.420000 1.990000 2.750000 2.735000 ;
        RECT 2.430000 0.595000 2.760000 0.980000 ;
        RECT 3.370000 1.990000 3.700000 2.735000 ;
        RECT 3.430000 0.595000 3.760000 0.980000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 10.560000 0.085000 ;
        RECT  4.290000  0.085000  4.620000 0.970000 ;
        RECT  5.230000  0.085000  5.400000 1.130000 ;
        RECT  6.010000  0.085000  6.260000 1.130000 ;
        RECT  6.870000  0.085000  7.120000 1.130000 ;
        RECT  9.330000  0.085000  9.500000 1.010000 ;
        RECT 10.110000  0.085000 10.445000 0.600000 ;
      LAYER mcon ;
        RECT  0.155000 -0.085000  0.325000 0.085000 ;
        RECT  0.635000 -0.085000  0.805000 0.085000 ;
        RECT  1.115000 -0.085000  1.285000 0.085000 ;
        RECT  1.595000 -0.085000  1.765000 0.085000 ;
        RECT  2.075000 -0.085000  2.245000 0.085000 ;
        RECT  2.555000 -0.085000  2.725000 0.085000 ;
        RECT  3.035000 -0.085000  3.205000 0.085000 ;
        RECT  3.515000 -0.085000  3.685000 0.085000 ;
        RECT  3.995000 -0.085000  4.165000 0.085000 ;
        RECT  4.475000 -0.085000  4.645000 0.085000 ;
        RECT  4.955000 -0.085000  5.125000 0.085000 ;
        RECT  5.435000 -0.085000  5.605000 0.085000 ;
        RECT  5.915000 -0.085000  6.085000 0.085000 ;
        RECT  6.395000 -0.085000  6.565000 0.085000 ;
        RECT  6.875000 -0.085000  7.045000 0.085000 ;
        RECT  7.355000 -0.085000  7.525000 0.085000 ;
        RECT  7.835000 -0.085000  8.005000 0.085000 ;
        RECT  8.315000 -0.085000  8.485000 0.085000 ;
        RECT  8.795000 -0.085000  8.965000 0.085000 ;
        RECT  9.275000 -0.085000  9.445000 0.085000 ;
        RECT  9.755000 -0.085000  9.925000 0.085000 ;
        RECT 10.235000 -0.085000 10.405000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.560000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 3.245000 10.560000 3.415000 ;
        RECT  4.370000 2.730000  4.700000 3.245000 ;
        RECT  5.370000 2.730000  5.700000 3.245000 ;
        RECT  6.370000 2.730000  6.700000 3.245000 ;
        RECT  7.405000 2.900000  7.735000 3.245000 ;
        RECT  9.165000 2.560000  9.495000 3.245000 ;
        RECT 10.115000 2.060000 10.445000 3.245000 ;
      LAYER mcon ;
        RECT  0.155000 3.245000  0.325000 3.415000 ;
        RECT  0.635000 3.245000  0.805000 3.415000 ;
        RECT  1.115000 3.245000  1.285000 3.415000 ;
        RECT  1.595000 3.245000  1.765000 3.415000 ;
        RECT  2.075000 3.245000  2.245000 3.415000 ;
        RECT  2.555000 3.245000  2.725000 3.415000 ;
        RECT  3.035000 3.245000  3.205000 3.415000 ;
        RECT  3.515000 3.245000  3.685000 3.415000 ;
        RECT  3.995000 3.245000  4.165000 3.415000 ;
        RECT  4.475000 3.245000  4.645000 3.415000 ;
        RECT  4.955000 3.245000  5.125000 3.415000 ;
        RECT  5.435000 3.245000  5.605000 3.415000 ;
        RECT  5.915000 3.245000  6.085000 3.415000 ;
        RECT  6.395000 3.245000  6.565000 3.415000 ;
        RECT  6.875000 3.245000  7.045000 3.415000 ;
        RECT  7.355000 3.245000  7.525000 3.415000 ;
        RECT  7.835000 3.245000  8.005000 3.415000 ;
        RECT  8.315000 3.245000  8.485000 3.415000 ;
        RECT  8.795000 3.245000  8.965000 3.415000 ;
        RECT  9.275000 3.245000  9.445000 3.415000 ;
        RECT  9.755000 3.245000  9.925000 3.415000 ;
        RECT 10.235000 3.245000 10.405000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 10.560000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.115000 0.255000  4.110000 0.425000 ;
      RECT  0.115000 0.425000  0.365000 1.130000 ;
      RECT  0.120000 1.820000  0.370000 2.905000 ;
      RECT  0.120000 2.905000  4.200000 3.075000 ;
      RECT  1.035000 1.320000  3.655000 1.480000 ;
      RECT  1.035000 1.480000  4.040000 1.650000 ;
      RECT  1.055000 0.425000  1.225000 0.810000 ;
      RECT  1.085000 2.160000  1.350000 2.905000 ;
      RECT  1.930000 0.425000  2.260000 0.810000 ;
      RECT  2.050000 2.160000  2.220000 2.905000 ;
      RECT  2.920000 2.160000  3.190000 2.905000 ;
      RECT  2.930000 0.425000  3.260000 0.810000 ;
      RECT  3.870000 1.650000  4.040000 2.050000 ;
      RECT  3.870000 2.050000  7.755000 2.220000 ;
      RECT  3.870000 2.390000  7.200000 2.560000 ;
      RECT  3.870000 2.560000  4.200000 2.905000 ;
      RECT  3.940000 0.425000  4.110000 1.140000 ;
      RECT  3.940000 1.140000  5.050000 1.300000 ;
      RECT  3.940000 1.300000  7.550000 1.310000 ;
      RECT  4.720000 1.310000  7.550000 1.470000 ;
      RECT  4.800000 0.350000  5.050000 1.140000 ;
      RECT  4.870000 2.560000  5.200000 2.980000 ;
      RECT  5.580000 0.350000  5.830000 1.300000 ;
      RECT  5.870000 2.560000  6.200000 2.980000 ;
      RECT  6.440000 0.350000  6.690000 1.300000 ;
      RECT  6.870000 2.560000  8.270000 2.730000 ;
      RECT  6.870000 2.730000  7.200000 2.980000 ;
      RECT  7.300000 0.350000  7.550000 1.300000 ;
      RECT  7.585000 2.220000  9.945000 2.390000 ;
      RECT  7.720000 0.340000  9.150000 0.670000 ;
      RECT  7.925000 0.670000  9.150000 1.010000 ;
      RECT  7.925000 1.010000  8.095000 1.800000 ;
      RECT  7.925000 1.800000  9.045000 2.050000 ;
      RECT  7.940000 2.730000  8.270000 2.980000 ;
      RECT  9.665000 1.720000 10.315000 1.890000 ;
      RECT  9.665000 1.890000  9.945000 2.220000 ;
      RECT  9.665000 2.390000  9.945000 2.980000 ;
      RECT  9.680000 0.340000  9.930000 0.840000 ;
      RECT  9.680000 0.840000 10.315000 1.010000 ;
      RECT 10.145000 1.010000 10.315000 1.720000 ;
  END
END sky130_fd_sc_ls__ebufn_8
