* NGSPICE file created from sky130_fd_sc_ls__sdfrbp_2.ext - technology: sky130A

.subckt sky130_fd_sc_ls__sdfrbp_2 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q Q_N
M1000 VGND RESET_B a_223_79# VNB nshort w=420000u l=150000u
+  ad=2.20027e+12p pd=1.854e+07u as=2.751e+11p ps=2.99e+06u
M1001 VPWR a_2006_373# a_1955_471# VPB phighvt w=420000u l=150000u
+  ad=3.4219e+12p pd=2.674e+07u as=1.134e+11p ps=1.38e+06u
M1002 a_1370_290# a_1223_119# VGND VNB nshort w=640000u l=150000u
+  ad=1.792e+11p pd=1.84e+06u as=0p ps=0u
M1003 VPWR a_1790_75# Q_N VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.36e+11p ps=2.84e+06u
M1004 a_1790_75# a_852_119# a_1370_290# VPB phighvt w=1e+06u l=150000u
+  ad=4.029e+11p pd=3.28e+06u as=3e+11p ps=2.6e+06u
M1005 a_2604_392# a_1790_75# VGND VNB nshort w=640000u l=150000u
+  ad=1.696e+11p pd=1.81e+06u as=0p ps=0u
M1006 VGND RESET_B a_1401_119# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1007 a_310_79# a_27_79# a_223_79# VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1008 a_223_79# SCD a_547_79# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1009 a_2006_373# RESET_B VPWR VPB phighvt w=420000u l=150000u
+  ad=1.26e+11p pd=1.44e+06u as=0p ps=0u
M1010 a_1223_119# a_852_119# a_388_79# VNB nshort w=420000u l=150000u
+  ad=1.47e+11p pd=1.54e+06u as=3.906e+11p ps=3.54e+06u
M1011 a_1323_119# a_1025_119# a_1223_119# VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1012 a_2604_392# a_1790_75# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.75e+11p pd=2.55e+06u as=0p ps=0u
M1013 a_2006_373# a_1790_75# a_2158_74# VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=8.82e+10p ps=1.26e+06u
M1014 a_538_464# a_27_79# a_388_79# VPB phighvt w=640000u l=150000u
+  ad=1.728e+11p pd=1.82e+06u as=6.808e+11p ps=5.72e+06u
M1015 a_1223_119# RESET_B VPWR VPB phighvt w=420000u l=150000u
+  ad=2.436e+11p pd=2.84e+06u as=0p ps=0u
M1016 a_1790_75# a_1025_119# a_1370_290# VNB nshort w=640000u l=150000u
+  ad=4.3185e+11p pd=3.09e+06u as=0p ps=0u
M1017 Q a_2604_392# VGND VNB nshort w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1018 a_388_79# D a_307_464# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1019 VGND CLK a_852_119# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.018e+11p ps=2.05e+06u
M1020 a_2158_74# RESET_B VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 Q_N a_1790_75# VGND VNB nshort w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1022 a_1325_457# a_852_119# a_1223_119# VPB phighvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1023 a_388_79# D a_310_79# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_1955_471# a_1025_119# a_1790_75# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPWR a_1790_75# a_2006_373# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VPWR SCE a_27_79# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.888e+11p ps=1.87e+06u
M1027 VGND SCE a_27_79# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1028 a_547_79# SCE a_388_79# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_1025_119# a_852_119# VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1030 a_307_464# SCE VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VPWR SCD a_538_464# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 VPWR CLK a_852_119# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.95e+11p ps=2.59e+06u
M1033 a_1223_119# a_1025_119# a_388_79# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 Q a_2604_392# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=0p ps=0u
M1035 a_1025_119# a_852_119# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.75e+11p pd=2.55e+06u as=0p ps=0u
M1036 Q_N a_1790_75# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 VGND a_1790_75# Q_N VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 VGND a_2604_392# Q VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_1370_290# a_1223_119# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1040 a_1401_119# a_1370_290# a_1323_119# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1041 VGND a_2006_373# a_2000_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1042 VPWR a_1370_290# a_1325_457# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1043 VPWR a_2604_392# Q VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1044 a_388_79# RESET_B VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1045 a_2000_74# a_852_119# a_1790_75# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

