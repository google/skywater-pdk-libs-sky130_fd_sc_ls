* File: sky130_fd_sc_ls__o21a_1.pex.spice
* Created: Fri Aug 28 13:44:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__O21A_1%A_83_244# 1 2 7 9 10 12 14 15 17 18 21 25 32
c59 25 0 1.80225e-19 $X=0.7 $Y=1.19
c60 21 0 1.20151e-20 $X=1.31 $Y=0.515
r61 28 30 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.7 $Y=1.385
+ $X2=0.7 $Y2=1.55
r62 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.7
+ $Y=1.385 $X2=0.7 $Y2=1.385
r63 25 28 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=0.7 $Y=1.19 $X2=0.7
+ $Y2=1.385
r64 19 21 27.1977 $w=2.48e-07 $l=5.9e-07 $layer=LI1_cond $X=1.27 $Y=1.105
+ $X2=1.27 $Y2=0.515
r65 17 32 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.36 $Y=2.035
+ $X2=1.525 $Y2=2.035
r66 17 18 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=1.36 $Y=2.035
+ $X2=0.865 $Y2=2.035
r67 16 25 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.865 $Y=1.19
+ $X2=0.7 $Y2=1.19
r68 15 19 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.145 $Y=1.19
+ $X2=1.27 $Y2=1.105
r69 15 16 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1.145 $Y=1.19
+ $X2=0.865 $Y2=1.19
r70 14 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.78 $Y=1.95
+ $X2=0.865 $Y2=2.035
r71 14 30 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=0.78 $Y=1.95 $X2=0.78
+ $Y2=1.55
r72 10 29 68.9212 $w=3.43e-07 $l=4.4238e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.64 $Y2=1.385
r73 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.4
r74 7 29 38.7084 $w=3.43e-07 $l=2.26164e-07 $layer=POLY_cond $X=0.495 $Y=1.22
+ $X2=0.64 $Y2=1.385
r75 7 9 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.495 $Y=1.22 $X2=0.495
+ $Y2=0.74
r76 2 32 300 $w=1.7e-07 $l=2.43721e-07 $layer=licon1_PDIFF $count=2 $X=1.375
+ $Y=1.935 $X2=1.525 $Y2=2.115
r77 1 21 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=1.165
+ $Y=0.37 $X2=1.31 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__O21A_1%B1 2 3 5 8 9 10 11
c42 10 0 1.80225e-19 $X=1.352 $Y=1.235
r43 11 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.27
+ $Y=1.61 $X2=1.27 $Y2=1.61
r44 9 10 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=1.352 $Y=1.085
+ $X2=1.352 $Y2=1.235
r45 8 9 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.525 $Y=0.69
+ $X2=1.525 $Y2=1.085
r46 3 14 53.429 $w=2.79e-07 $l=2.64575e-07 $layer=POLY_cond $X=1.3 $Y=1.86
+ $X2=1.27 $Y2=1.61
r47 3 5 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.3 $Y=1.86 $X2=1.3
+ $Y2=2.355
r48 2 14 1.29086 $w=3.3e-07 $l=8.75758e-08 $layer=POLY_cond $X=1.27 $Y=1.61
+ $X2=1.27 $Y2=1.61
r49 2 10 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=1.27 $Y=1.61 $X2=1.27
+ $Y2=1.235
.ends

.subckt PM_SKY130_FD_SC_LS__O21A_1%A2 1 3 6 8
c31 6 0 1.56978e-19 $X=1.955 $Y=0.69
r32 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.88
+ $Y=1.61 $X2=1.88 $Y2=1.61
r33 8 12 9.63236 $w=3.33e-07 $l=2.8e-07 $layer=LI1_cond $X=2.16 $Y=1.612
+ $X2=1.88 $Y2=1.612
r34 4 11 38.5562 $w=2.99e-07 $l=1.98997e-07 $layer=POLY_cond $X=1.955 $Y=1.445
+ $X2=1.88 $Y2=1.61
r35 4 6 387.138 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=1.955 $Y=1.445
+ $X2=1.955 $Y2=0.69
r36 1 11 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=1.805 $Y=1.86
+ $X2=1.88 $Y2=1.61
r37 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.805 $Y=1.86
+ $X2=1.805 $Y2=2.435
.ends

.subckt PM_SKY130_FD_SC_LS__O21A_1%A1 1 3 6 8 12
r22 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.61
+ $Y=1.465 $X2=2.61 $Y2=1.465
r23 8 12 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=2.61 $Y=1.665 $X2=2.61
+ $Y2=1.465
r24 4 11 38.7502 $w=3.47e-07 $l=2.26164e-07 $layer=POLY_cond $X=2.385 $Y=1.3
+ $X2=2.53 $Y2=1.465
r25 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.385 $Y=1.3 $X2=2.385
+ $Y2=0.69
r26 1 11 70.6983 $w=3.47e-07 $l=4.66101e-07 $layer=POLY_cond $X=2.375 $Y=1.86
+ $X2=2.53 $Y2=1.465
r27 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.375 $Y=1.86
+ $X2=2.375 $Y2=2.435
.ends

.subckt PM_SKY130_FD_SC_LS__O21A_1%X 1 2 7 8 9 10 11 12 13 36
r16 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.28 $Y=2.405
+ $X2=0.28 $Y2=2.775
r17 11 36 0.628605 $w=3.28e-07 $l=1.8e-08 $layer=LI1_cond $X=0.28 $Y=1.967
+ $X2=0.28 $Y2=1.985
r18 11 45 5.83828 $w=3.28e-07 $l=1.47e-07 $layer=LI1_cond $X=0.28 $Y=1.967
+ $X2=0.28 $Y2=1.82
r19 11 12 12.3276 $w=3.28e-07 $l=3.53e-07 $layer=LI1_cond $X=0.28 $Y=2.052
+ $X2=0.28 $Y2=2.405
r20 11 36 2.33981 $w=3.28e-07 $l=6.7e-08 $layer=LI1_cond $X=0.28 $Y=2.052
+ $X2=0.28 $Y2=1.985
r21 10 45 7.14515 $w=2.48e-07 $l=1.55e-07 $layer=LI1_cond $X=0.24 $Y=1.665
+ $X2=0.24 $Y2=1.82
r22 9 10 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=1.295
+ $X2=0.24 $Y2=1.665
r23 8 9 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=0.925 $X2=0.24
+ $Y2=1.295
r24 7 8 18.9001 $w=2.48e-07 $l=4.1e-07 $layer=LI1_cond $X=0.24 $Y=0.515 $X2=0.24
+ $Y2=0.925
r25 2 13 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r26 2 36 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
r27 1 7 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__O21A_1%VPWR 1 2 9 11 13 17 19 24 33 37
r33 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r34 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r35 31 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r36 30 31 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r37 28 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r38 27 30 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r39 27 28 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r40 25 33 12.1365 $w=1.7e-07 $l=2.83e-07 $layer=LI1_cond $X=1.18 $Y=3.33
+ $X2=0.897 $Y2=3.33
r41 25 27 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=1.18 $Y=3.33 $X2=1.2
+ $Y2=3.33
r42 24 36 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=2.435 $Y=3.33
+ $X2=2.657 $Y2=3.33
r43 24 30 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.435 $Y=3.33
+ $X2=2.16 $Y2=3.33
r44 22 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r45 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r46 19 33 12.1365 $w=1.7e-07 $l=2.82e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.897 $Y2=3.33
r47 19 21 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.24 $Y2=3.33
r48 17 31 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=2.16 $Y2=3.33
r49 17 28 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.2 $Y2=3.33
r50 13 16 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=2.6 $Y=2.11 $X2=2.6
+ $Y2=2.79
r51 11 36 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=2.6 $Y=3.245
+ $X2=2.657 $Y2=3.33
r52 11 16 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=2.6 $Y=3.245
+ $X2=2.6 $Y2=2.79
r53 7 33 2.37858 $w=5.65e-07 $l=8.5e-08 $layer=LI1_cond $X=0.897 $Y=3.245
+ $X2=0.897 $Y2=3.33
r54 7 9 16.7239 $w=5.63e-07 $l=7.9e-07 $layer=LI1_cond $X=0.897 $Y=3.245
+ $X2=0.897 $Y2=2.455
r55 2 16 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=2.45
+ $Y=1.935 $X2=2.6 $Y2=2.79
r56 2 13 400 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=1 $X=2.45
+ $Y=1.935 $X2=2.6 $Y2=2.11
r57 1 9 200 $w=1.7e-07 $l=8.26226e-07 $layer=licon1_PDIFF $count=3 $X=0.58
+ $Y=1.84 $X2=1.075 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_LS__O21A_1%VGND 1 2 9 13 15 17 22 29 30 33 36
r39 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r40 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r41 30 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r42 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r43 27 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.335 $Y=0 $X2=2.17
+ $Y2=0
r44 27 29 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.335 $Y=0 $X2=2.64
+ $Y2=0
r45 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r46 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r47 23 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=0.71
+ $Y2=0
r48 23 25 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=1.68
+ $Y2=0
r49 22 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.005 $Y=0 $X2=2.17
+ $Y2=0
r50 22 25 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.005 $Y=0 $X2=1.68
+ $Y2=0
r51 20 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r52 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r53 17 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.71
+ $Y2=0
r54 17 19 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.24
+ $Y2=0
r55 15 26 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.68
+ $Y2=0
r56 15 34 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=0.72
+ $Y2=0
r57 11 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.17 $Y=0.085
+ $X2=2.17 $Y2=0
r58 11 13 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=2.17 $Y=0.085
+ $X2=2.17 $Y2=0.57
r59 7 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=0.085 $X2=0.71
+ $Y2=0
r60 7 9 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0.51
r61 2 13 182 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=1 $X=2.03
+ $Y=0.37 $X2=2.17 $Y2=0.57
r62 1 9 91 $w=1.7e-07 $l=1.9799e-07 $layer=licon1_NDIFF $count=2 $X=0.57 $Y=0.37
+ $X2=0.71 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_LS__O21A_1%A_320_74# 1 2 9 11 12 15
c27 9 0 1.44963e-19 $X=1.74 $Y=0.515
r28 13 15 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=2.64 $Y=0.96
+ $X2=2.64 $Y2=0.515
r29 11 13 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.515 $Y=1.045
+ $X2=2.64 $Y2=0.96
r30 11 12 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.515 $Y=1.045
+ $X2=1.825 $Y2=1.045
r31 7 12 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.7 $Y=0.96
+ $X2=1.825 $Y2=1.045
r32 7 9 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=1.7 $Y=0.96 $X2=1.7
+ $Y2=0.515
r33 2 15 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.46
+ $Y=0.37 $X2=2.6 $Y2=0.515
r34 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.6 $Y=0.37
+ $X2=1.74 $Y2=0.515
.ends

