* File: sky130_fd_sc_ls__o221ai_1.pxi.spice
* Created: Wed Sep  2 11:19:32 2020
* 
x_PM_SKY130_FD_SC_LS__O221AI_1%C1 N_C1_M1008_g N_C1_c_61_n N_C1_M1000_g C1
+ N_C1_c_59_n N_C1_c_60_n PM_SKY130_FD_SC_LS__O221AI_1%C1
x_PM_SKY130_FD_SC_LS__O221AI_1%B1 N_B1_c_88_n N_B1_M1009_g N_B1_M1003_g B1
+ N_B1_c_86_n N_B1_c_87_n PM_SKY130_FD_SC_LS__O221AI_1%B1
x_PM_SKY130_FD_SC_LS__O221AI_1%B2 N_B2_c_119_n N_B2_M1007_g N_B2_M1002_g B2
+ N_B2_c_121_n PM_SKY130_FD_SC_LS__O221AI_1%B2
x_PM_SKY130_FD_SC_LS__O221AI_1%A2 N_A2_c_155_n N_A2_M1004_g N_A2_M1001_g A2 A2
+ A2 A2 N_A2_c_157_n A2 PM_SKY130_FD_SC_LS__O221AI_1%A2
x_PM_SKY130_FD_SC_LS__O221AI_1%A1 N_A1_c_201_n N_A1_M1006_g N_A1_M1005_g A1 A1
+ N_A1_c_200_n PM_SKY130_FD_SC_LS__O221AI_1%A1
x_PM_SKY130_FD_SC_LS__O221AI_1%Y N_Y_M1008_s N_Y_M1000_s N_Y_M1007_d N_Y_c_229_n
+ N_Y_c_226_n N_Y_c_247_n N_Y_c_237_n N_Y_c_253_n N_Y_c_231_n Y Y Y N_Y_c_228_n
+ PM_SKY130_FD_SC_LS__O221AI_1%Y
x_PM_SKY130_FD_SC_LS__O221AI_1%VPWR N_VPWR_M1000_d N_VPWR_M1006_d N_VPWR_c_278_n
+ N_VPWR_c_279_n N_VPWR_c_280_n N_VPWR_c_281_n VPWR N_VPWR_c_282_n
+ N_VPWR_c_283_n N_VPWR_c_277_n N_VPWR_c_285_n PM_SKY130_FD_SC_LS__O221AI_1%VPWR
x_PM_SKY130_FD_SC_LS__O221AI_1%A_114_74# N_A_114_74#_M1008_d N_A_114_74#_M1003_d
+ N_A_114_74#_c_317_n N_A_114_74#_c_318_n N_A_114_74#_c_319_n
+ PM_SKY130_FD_SC_LS__O221AI_1%A_114_74#
x_PM_SKY130_FD_SC_LS__O221AI_1%A_239_74# N_A_239_74#_M1003_s N_A_239_74#_M1002_d
+ N_A_239_74#_M1005_d N_A_239_74#_c_340_n N_A_239_74#_c_341_n
+ N_A_239_74#_c_342_n N_A_239_74#_c_343_n N_A_239_74#_c_344_n
+ N_A_239_74#_c_345_n PM_SKY130_FD_SC_LS__O221AI_1%A_239_74#
x_PM_SKY130_FD_SC_LS__O221AI_1%VGND N_VGND_M1001_d N_VGND_c_386_n VGND
+ N_VGND_c_387_n N_VGND_c_388_n N_VGND_c_389_n N_VGND_c_390_n
+ PM_SKY130_FD_SC_LS__O221AI_1%VGND
cc_1 VNB N_C1_M1008_g 0.0339542f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_C1_c_59_n 0.00448523f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_3 VNB N_C1_c_60_n 0.0699552f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.532
cc_4 VNB N_B1_M1003_g 0.0340087f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_5 VNB N_B1_c_86_n 0.0486827f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.532
cc_6 VNB N_B1_c_87_n 0.0109062f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.532
cc_7 VNB N_B2_c_119_n 0.025098f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.3
cc_8 VNB N_B2_M1002_g 0.0259532f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=2.4
cc_9 VNB N_B2_c_121_n 0.00419897f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_10 VNB N_A2_c_155_n 0.0269917f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.3
cc_11 VNB N_A2_M1001_g 0.0287203f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=2.4
cc_12 VNB N_A2_c_157_n 0.00179855f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A1_M1005_g 0.0335202f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=2.4
cc_14 VNB A1 0.0179013f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A1_c_200_n 0.0656045f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.532
cc_16 VNB N_Y_c_226_n 0.0116419f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_17 VNB Y 0.0258829f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_Y_c_228_n 0.00992326f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_VPWR_c_277_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_114_74#_c_317_n 0.0150295f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=2.4
cc_21 VNB N_A_114_74#_c_318_n 0.00814237f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_114_74#_c_319_n 0.00262119f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.532
cc_23 VNB N_A_239_74#_c_340_n 0.00920118f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.532
cc_24 VNB N_A_239_74#_c_341_n 0.00279871f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.532
cc_25 VNB N_A_239_74#_c_342_n 0.0200423f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_239_74#_c_343_n 0.02581f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_239_74#_c_344_n 0.00726397f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_239_74#_c_345_n 0.00804404f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_386_n 0.0121692f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=2.4
cc_30 VNB N_VGND_c_387_n 0.0713008f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.532
cc_31 VNB N_VGND_c_388_n 0.0191515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_389_n 0.233314f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_390_n 0.0105791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VPB N_C1_c_61_n 0.0220341f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.765
cc_35 VPB N_C1_c_59_n 0.0147422f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_36 VPB N_C1_c_60_n 0.00781219f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.532
cc_37 VPB N_B1_c_88_n 0.0175528f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_38 VPB N_B1_c_86_n 0.0223613f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.532
cc_39 VPB N_B1_c_87_n 0.00559402f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.532
cc_40 VPB N_B2_c_119_n 0.0276986f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.3
cc_41 VPB N_B2_c_121_n 0.00322696f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_42 VPB N_A2_c_155_n 0.0295057f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.3
cc_43 VPB A2 0.00133136f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_44 VPB N_A1_c_201_n 0.0199541f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.3
cc_45 VPB A1 0.0182935f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_A1_c_200_n 0.00756982f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.532
cc_47 VPB N_Y_c_229_n 0.00276769f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_48 VPB N_Y_c_226_n 0.0018342f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_49 VPB N_Y_c_231_n 0.0029874f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_278_n 0.0109451f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_279_n 0.0485725f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.532
cc_52 VPB N_VPWR_c_280_n 0.0465089f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_281_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_282_n 0.0239133f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_283_n 0.0131219f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_277_n 0.0960602f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_285_n 0.0154008f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 N_C1_c_60_n N_B1_c_86_n 0.0145689f $X=0.495 $Y=1.532 $X2=0 $Y2=0
cc_59 N_C1_c_60_n N_B1_c_87_n 8.15661e-19 $X=0.495 $Y=1.532 $X2=0 $Y2=0
cc_60 N_C1_c_61_n N_Y_c_229_n 0.0144227f $X=0.635 $Y=1.765 $X2=0 $Y2=0
cc_61 N_C1_M1008_g N_Y_c_226_n 0.00950615f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_62 N_C1_c_61_n N_Y_c_226_n 0.0113471f $X=0.635 $Y=1.765 $X2=0 $Y2=0
cc_63 N_C1_c_59_n N_Y_c_226_n 0.0355293f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_64 N_C1_c_60_n N_Y_c_226_n 0.010892f $X=0.495 $Y=1.532 $X2=0 $Y2=0
cc_65 N_C1_c_61_n N_Y_c_237_n 0.0146819f $X=0.635 $Y=1.765 $X2=0 $Y2=0
cc_66 N_C1_c_59_n N_Y_c_237_n 0.00880161f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_67 N_C1_c_60_n N_Y_c_237_n 0.00383619f $X=0.495 $Y=1.532 $X2=0 $Y2=0
cc_68 N_C1_M1008_g Y 0.0146416f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_69 N_C1_M1008_g N_Y_c_228_n 0.0173829f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_70 N_C1_c_59_n N_Y_c_228_n 0.0247471f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_71 N_C1_c_60_n N_Y_c_228_n 0.00374051f $X=0.495 $Y=1.532 $X2=0 $Y2=0
cc_72 N_C1_c_61_n N_VPWR_c_278_n 0.00565407f $X=0.635 $Y=1.765 $X2=0 $Y2=0
cc_73 N_C1_c_61_n N_VPWR_c_282_n 0.00445602f $X=0.635 $Y=1.765 $X2=0 $Y2=0
cc_74 N_C1_c_61_n N_VPWR_c_277_n 0.00865571f $X=0.635 $Y=1.765 $X2=0 $Y2=0
cc_75 N_C1_M1008_g N_A_114_74#_c_318_n 0.00122485f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_76 N_C1_M1008_g N_A_239_74#_c_344_n 0.00471147f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_77 N_C1_M1008_g N_VGND_c_387_n 0.00434272f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_78 N_C1_M1008_g N_VGND_c_389_n 0.00829926f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_79 N_B1_c_88_n N_B2_c_119_n 0.0595838f $X=1.545 $Y=1.765 $X2=-0.19 $Y2=-0.245
cc_80 N_B1_c_86_n N_B2_c_119_n 0.0220632f $X=1.47 $Y=1.515 $X2=-0.19 $Y2=-0.245
cc_81 N_B1_c_87_n N_B2_c_119_n 0.00155181f $X=1.47 $Y=1.515 $X2=-0.19 $Y2=-0.245
cc_82 N_B1_M1003_g N_B2_M1002_g 0.0313505f $X=1.555 $Y=0.74 $X2=0 $Y2=0
cc_83 N_B1_c_86_n N_B2_c_121_n 0.00166897f $X=1.47 $Y=1.515 $X2=0 $Y2=0
cc_84 N_B1_c_87_n N_B2_c_121_n 0.0263986f $X=1.47 $Y=1.515 $X2=0 $Y2=0
cc_85 N_B1_c_88_n N_Y_c_226_n 0.00343144f $X=1.545 $Y=1.765 $X2=0 $Y2=0
cc_86 N_B1_c_86_n N_Y_c_226_n 0.00258218f $X=1.47 $Y=1.515 $X2=0 $Y2=0
cc_87 N_B1_c_87_n N_Y_c_226_n 0.0318707f $X=1.47 $Y=1.515 $X2=0 $Y2=0
cc_88 N_B1_c_88_n N_Y_c_247_n 0.0142797f $X=1.545 $Y=1.765 $X2=0 $Y2=0
cc_89 N_B1_c_86_n N_Y_c_247_n 0.00258259f $X=1.47 $Y=1.515 $X2=0 $Y2=0
cc_90 N_B1_c_87_n N_Y_c_247_n 0.0498623f $X=1.47 $Y=1.515 $X2=0 $Y2=0
cc_91 N_B1_c_88_n N_Y_c_231_n 0.0027401f $X=1.545 $Y=1.765 $X2=0 $Y2=0
cc_92 N_B1_c_88_n N_VPWR_c_278_n 0.0243302f $X=1.545 $Y=1.765 $X2=0 $Y2=0
cc_93 N_B1_c_88_n N_VPWR_c_280_n 0.00183185f $X=1.545 $Y=1.765 $X2=0 $Y2=0
cc_94 N_B1_c_88_n N_VPWR_c_277_n 0.00367613f $X=1.545 $Y=1.765 $X2=0 $Y2=0
cc_95 N_B1_M1003_g N_A_114_74#_c_317_n 0.0121776f $X=1.555 $Y=0.74 $X2=0 $Y2=0
cc_96 N_B1_M1003_g N_A_114_74#_c_318_n 0.00672761f $X=1.555 $Y=0.74 $X2=0 $Y2=0
cc_97 N_B1_M1003_g N_A_114_74#_c_319_n 4.44647e-19 $X=1.555 $Y=0.74 $X2=0 $Y2=0
cc_98 N_B1_M1003_g N_A_239_74#_c_340_n 0.00961368f $X=1.555 $Y=0.74 $X2=0 $Y2=0
cc_99 N_B1_c_87_n N_A_239_74#_c_340_n 0.00947557f $X=1.47 $Y=1.515 $X2=0 $Y2=0
cc_100 N_B1_M1003_g N_A_239_74#_c_344_n 0.00723558f $X=1.555 $Y=0.74 $X2=0 $Y2=0
cc_101 N_B1_c_86_n N_A_239_74#_c_344_n 0.00227486f $X=1.47 $Y=1.515 $X2=0 $Y2=0
cc_102 N_B1_c_87_n N_A_239_74#_c_344_n 0.0268812f $X=1.47 $Y=1.515 $X2=0 $Y2=0
cc_103 N_B1_M1003_g N_VGND_c_387_n 0.00291649f $X=1.555 $Y=0.74 $X2=0 $Y2=0
cc_104 N_B1_M1003_g N_VGND_c_389_n 0.00364831f $X=1.555 $Y=0.74 $X2=0 $Y2=0
cc_105 N_B2_c_119_n N_A2_c_155_n 0.03861f $X=1.965 $Y=1.765 $X2=-0.19 $Y2=-0.245
cc_106 N_B2_c_121_n N_A2_c_155_n 0.00286759f $X=2.04 $Y=1.515 $X2=-0.19
+ $Y2=-0.245
cc_107 N_B2_M1002_g N_A2_M1001_g 0.0247498f $X=2.055 $Y=0.74 $X2=0 $Y2=0
cc_108 N_B2_c_119_n A2 8.64739e-19 $X=1.965 $Y=1.765 $X2=0 $Y2=0
cc_109 N_B2_c_121_n A2 0.0058624f $X=2.04 $Y=1.515 $X2=0 $Y2=0
cc_110 N_B2_c_119_n N_A2_c_157_n 3.65288e-19 $X=1.965 $Y=1.765 $X2=0 $Y2=0
cc_111 N_B2_c_121_n N_A2_c_157_n 0.0265213f $X=2.04 $Y=1.515 $X2=0 $Y2=0
cc_112 N_B2_c_119_n N_Y_c_247_n 0.0117753f $X=1.965 $Y=1.765 $X2=0 $Y2=0
cc_113 N_B2_c_121_n N_Y_c_247_n 0.0104762f $X=2.04 $Y=1.515 $X2=0 $Y2=0
cc_114 N_B2_c_119_n N_Y_c_253_n 0.00123893f $X=1.965 $Y=1.765 $X2=0 $Y2=0
cc_115 N_B2_c_121_n N_Y_c_253_n 0.0193965f $X=2.04 $Y=1.515 $X2=0 $Y2=0
cc_116 N_B2_c_119_n N_Y_c_231_n 0.0140982f $X=1.965 $Y=1.765 $X2=0 $Y2=0
cc_117 N_B2_c_119_n N_VPWR_c_278_n 0.00285765f $X=1.965 $Y=1.765 $X2=0 $Y2=0
cc_118 N_B2_c_119_n N_VPWR_c_280_n 0.00445602f $X=1.965 $Y=1.765 $X2=0 $Y2=0
cc_119 N_B2_c_119_n N_VPWR_c_277_n 0.00859212f $X=1.965 $Y=1.765 $X2=0 $Y2=0
cc_120 N_B2_M1002_g N_A_114_74#_c_319_n 0.00617064f $X=2.055 $Y=0.74 $X2=0 $Y2=0
cc_121 N_B2_c_119_n N_A_239_74#_c_340_n 0.00103933f $X=1.965 $Y=1.765 $X2=0
+ $Y2=0
cc_122 N_B2_M1002_g N_A_239_74#_c_340_n 0.015042f $X=2.055 $Y=0.74 $X2=0 $Y2=0
cc_123 N_B2_c_121_n N_A_239_74#_c_340_n 0.0224475f $X=2.04 $Y=1.515 $X2=0 $Y2=0
cc_124 N_B2_M1002_g N_A_239_74#_c_341_n 0.00324276f $X=2.055 $Y=0.74 $X2=0 $Y2=0
cc_125 N_B2_M1002_g N_A_239_74#_c_344_n 6.83744e-19 $X=2.055 $Y=0.74 $X2=0 $Y2=0
cc_126 N_B2_c_119_n N_A_239_74#_c_345_n 2.37442e-19 $X=1.965 $Y=1.765 $X2=0
+ $Y2=0
cc_127 N_B2_c_121_n N_A_239_74#_c_345_n 0.00883898f $X=2.04 $Y=1.515 $X2=0 $Y2=0
cc_128 N_B2_M1002_g N_VGND_c_387_n 0.00434272f $X=2.055 $Y=0.74 $X2=0 $Y2=0
cc_129 N_B2_M1002_g N_VGND_c_389_n 0.00822693f $X=2.055 $Y=0.74 $X2=0 $Y2=0
cc_130 N_A2_c_155_n N_A1_c_201_n 0.0318252f $X=2.535 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_131 A2 N_A1_c_201_n 0.0115418f $X=2.555 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_132 N_A2_M1001_g N_A1_M1005_g 0.0111967f $X=2.555 $Y=0.74 $X2=0 $Y2=0
cc_133 N_A2_c_155_n A1 0.00253478f $X=2.535 $Y=1.765 $X2=0 $Y2=0
cc_134 N_A2_M1001_g A1 0.00109635f $X=2.555 $Y=0.74 $X2=0 $Y2=0
cc_135 N_A2_c_157_n A1 0.0292169f $X=2.61 $Y=1.515 $X2=0 $Y2=0
cc_136 N_A2_c_155_n N_A1_c_200_n 0.0200708f $X=2.535 $Y=1.765 $X2=0 $Y2=0
cc_137 N_A2_M1001_g N_A1_c_200_n 0.00138545f $X=2.555 $Y=0.74 $X2=0 $Y2=0
cc_138 A2 N_A1_c_200_n 3.15765e-19 $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_139 N_A2_c_157_n N_A1_c_200_n 4.11342e-19 $X=2.61 $Y=1.515 $X2=0 $Y2=0
cc_140 N_A2_c_155_n N_Y_c_253_n 0.00150908f $X=2.535 $Y=1.765 $X2=0 $Y2=0
cc_141 A2 N_Y_c_253_n 0.0137716f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_142 N_A2_c_155_n N_Y_c_231_n 0.00882811f $X=2.535 $Y=1.765 $X2=0 $Y2=0
cc_143 A2 N_Y_c_231_n 0.0585277f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_144 N_A2_c_155_n N_VPWR_c_279_n 0.00172253f $X=2.535 $Y=1.765 $X2=0 $Y2=0
cc_145 A2 N_VPWR_c_279_n 0.0376974f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_146 N_A2_c_155_n N_VPWR_c_280_n 0.00372889f $X=2.535 $Y=1.765 $X2=0 $Y2=0
cc_147 A2 N_VPWR_c_280_n 0.00687333f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_148 N_A2_c_155_n N_VPWR_c_277_n 0.00610745f $X=2.535 $Y=1.765 $X2=0 $Y2=0
cc_149 A2 N_VPWR_c_277_n 0.00822835f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_150 A2 A_522_368# 0.0145626f $X=2.555 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_151 N_A2_M1001_g N_A_239_74#_c_341_n 0.013204f $X=2.555 $Y=0.74 $X2=0 $Y2=0
cc_152 N_A2_c_155_n N_A_239_74#_c_342_n 9.61123e-19 $X=2.535 $Y=1.765 $X2=0
+ $Y2=0
cc_153 N_A2_M1001_g N_A_239_74#_c_342_n 0.0127283f $X=2.555 $Y=0.74 $X2=0 $Y2=0
cc_154 N_A2_c_157_n N_A_239_74#_c_342_n 0.0171097f $X=2.61 $Y=1.515 $X2=0 $Y2=0
cc_155 N_A2_c_155_n N_A_239_74#_c_345_n 2.6682e-19 $X=2.535 $Y=1.765 $X2=0 $Y2=0
cc_156 N_A2_M1001_g N_A_239_74#_c_345_n 0.00406658f $X=2.555 $Y=0.74 $X2=0 $Y2=0
cc_157 N_A2_c_157_n N_A_239_74#_c_345_n 0.00488735f $X=2.61 $Y=1.515 $X2=0 $Y2=0
cc_158 N_A2_M1001_g N_VGND_c_386_n 0.00450194f $X=2.555 $Y=0.74 $X2=0 $Y2=0
cc_159 N_A2_M1001_g N_VGND_c_387_n 0.00434272f $X=2.555 $Y=0.74 $X2=0 $Y2=0
cc_160 N_A2_M1001_g N_VGND_c_389_n 0.00823337f $X=2.555 $Y=0.74 $X2=0 $Y2=0
cc_161 N_A1_c_201_n N_VPWR_c_279_n 0.0208463f $X=3.105 $Y=1.765 $X2=0 $Y2=0
cc_162 A1 N_VPWR_c_279_n 0.0265674f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_163 N_A1_c_200_n N_VPWR_c_279_n 0.00154884f $X=3.345 $Y=1.532 $X2=0 $Y2=0
cc_164 N_A1_c_201_n N_VPWR_c_280_n 0.00413917f $X=3.105 $Y=1.765 $X2=0 $Y2=0
cc_165 N_A1_c_201_n N_VPWR_c_277_n 0.00818781f $X=3.105 $Y=1.765 $X2=0 $Y2=0
cc_166 N_A1_M1005_g N_A_239_74#_c_342_n 0.0136182f $X=3.345 $Y=0.74 $X2=0 $Y2=0
cc_167 A1 N_A_239_74#_c_342_n 0.0574315f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_168 N_A1_c_200_n N_A_239_74#_c_342_n 0.012531f $X=3.345 $Y=1.532 $X2=0 $Y2=0
cc_169 N_A1_M1005_g N_A_239_74#_c_343_n 0.0138506f $X=3.345 $Y=0.74 $X2=0 $Y2=0
cc_170 N_A1_M1005_g N_VGND_c_386_n 0.00450194f $X=3.345 $Y=0.74 $X2=0 $Y2=0
cc_171 N_A1_M1005_g N_VGND_c_388_n 0.00434272f $X=3.345 $Y=0.74 $X2=0 $Y2=0
cc_172 N_A1_M1005_g N_VGND_c_389_n 0.00826283f $X=3.345 $Y=0.74 $X2=0 $Y2=0
cc_173 N_Y_c_226_n N_VPWR_M1000_d 0.00200633f $X=0.69 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_174 N_Y_c_247_n N_VPWR_M1000_d 0.0216166f $X=2.025 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_175 N_Y_c_229_n N_VPWR_c_278_n 0.0256941f $X=0.41 $Y=2.815 $X2=0 $Y2=0
cc_176 N_Y_c_237_n N_VPWR_c_278_n 0.0592221f $X=0.775 $Y=2.035 $X2=0 $Y2=0
cc_177 N_Y_c_231_n N_VPWR_c_278_n 0.0242156f $X=2.19 $Y=2.815 $X2=0 $Y2=0
cc_178 N_Y_c_231_n N_VPWR_c_280_n 0.0145938f $X=2.19 $Y=2.815 $X2=0 $Y2=0
cc_179 N_Y_c_229_n N_VPWR_c_282_n 0.0110241f $X=0.41 $Y=2.815 $X2=0 $Y2=0
cc_180 N_Y_c_229_n N_VPWR_c_277_n 0.00909194f $X=0.41 $Y=2.815 $X2=0 $Y2=0
cc_181 N_Y_c_231_n N_VPWR_c_277_n 0.0120466f $X=2.19 $Y=2.815 $X2=0 $Y2=0
cc_182 N_Y_c_247_n A_324_368# 0.0119045f $X=2.025 $Y=2.035 $X2=-0.19 $Y2=-0.245
cc_183 N_Y_c_228_n N_A_114_74#_M1008_d 0.00435283f $X=0.69 $Y=1.045 $X2=-0.19
+ $Y2=-0.245
cc_184 Y N_A_114_74#_c_318_n 0.0165499f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_185 N_Y_c_228_n N_A_114_74#_c_318_n 0.01066f $X=0.69 $Y=1.045 $X2=0 $Y2=0
cc_186 N_Y_c_226_n N_A_239_74#_c_344_n 0.00219497f $X=0.69 $Y=1.95 $X2=0 $Y2=0
cc_187 N_Y_c_228_n N_A_239_74#_c_344_n 0.00790447f $X=0.69 $Y=1.045 $X2=0 $Y2=0
cc_188 Y N_VGND_c_387_n 0.0144497f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_189 Y N_VGND_c_389_n 0.0119539f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_190 N_A_114_74#_c_317_n N_A_239_74#_M1003_s 0.00390908f $X=1.675 $Y=0.435
+ $X2=-0.19 $Y2=-0.245
cc_191 N_A_114_74#_M1003_d N_A_239_74#_c_340_n 0.00277863f $X=1.63 $Y=0.37 $X2=0
+ $Y2=0
cc_192 N_A_114_74#_c_317_n N_A_239_74#_c_340_n 0.00357806f $X=1.675 $Y=0.435
+ $X2=0 $Y2=0
cc_193 N_A_114_74#_c_319_n N_A_239_74#_c_340_n 0.0170103f $X=1.84 $Y=0.435 $X2=0
+ $Y2=0
cc_194 N_A_114_74#_c_319_n N_A_239_74#_c_341_n 0.017488f $X=1.84 $Y=0.435 $X2=0
+ $Y2=0
cc_195 N_A_114_74#_c_317_n N_A_239_74#_c_344_n 0.013123f $X=1.675 $Y=0.435 $X2=0
+ $Y2=0
cc_196 N_A_114_74#_c_317_n N_VGND_c_387_n 0.0290838f $X=1.675 $Y=0.435 $X2=0
+ $Y2=0
cc_197 N_A_114_74#_c_318_n N_VGND_c_387_n 0.0141382f $X=0.78 $Y=0.435 $X2=0
+ $Y2=0
cc_198 N_A_114_74#_c_319_n N_VGND_c_387_n 0.0141284f $X=1.84 $Y=0.435 $X2=0
+ $Y2=0
cc_199 N_A_114_74#_c_317_n N_VGND_c_389_n 0.0250986f $X=1.675 $Y=0.435 $X2=0
+ $Y2=0
cc_200 N_A_114_74#_c_318_n N_VGND_c_389_n 0.0119234f $X=0.78 $Y=0.435 $X2=0
+ $Y2=0
cc_201 N_A_114_74#_c_319_n N_VGND_c_389_n 0.0118299f $X=1.84 $Y=0.435 $X2=0
+ $Y2=0
cc_202 N_A_239_74#_c_342_n N_VGND_M1001_d 0.0079007f $X=3.395 $Y=1.045 $X2=-0.19
+ $Y2=-0.245
cc_203 N_A_239_74#_c_341_n N_VGND_c_386_n 0.0173638f $X=2.34 $Y=0.515 $X2=0
+ $Y2=0
cc_204 N_A_239_74#_c_342_n N_VGND_c_386_n 0.0427946f $X=3.395 $Y=1.045 $X2=0
+ $Y2=0
cc_205 N_A_239_74#_c_343_n N_VGND_c_386_n 0.0173638f $X=3.56 $Y=0.515 $X2=0
+ $Y2=0
cc_206 N_A_239_74#_c_341_n N_VGND_c_387_n 0.0145639f $X=2.34 $Y=0.515 $X2=0
+ $Y2=0
cc_207 N_A_239_74#_c_343_n N_VGND_c_388_n 0.0145639f $X=3.56 $Y=0.515 $X2=0
+ $Y2=0
cc_208 N_A_239_74#_c_341_n N_VGND_c_389_n 0.0119984f $X=2.34 $Y=0.515 $X2=0
+ $Y2=0
cc_209 N_A_239_74#_c_343_n N_VGND_c_389_n 0.0119984f $X=3.56 $Y=0.515 $X2=0
+ $Y2=0
