* NGSPICE file created from sky130_fd_sc_ls__o2111ai_1.ext - technology: sky130A

.subckt sky130_fd_sc_ls__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
M1000 Y B1 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=7e+11p pd=5.73e+06u as=1.2544e+12p ps=8.96e+06u
M1001 a_368_74# B1 a_260_74# VNB nshort w=740000u l=150000u
+  ad=4.773e+11p pd=4.25e+06u as=2.886e+11p ps=2.26e+06u
M1002 VGND A2 a_368_74# VNB nshort w=740000u l=150000u
+  ad=3.256e+11p pd=2.36e+06u as=0p ps=0u
M1003 Y D1 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_368_74# A1 VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR C1 Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_182_74# D1 Y VNB nshort w=740000u l=150000u
+  ad=1.776e+11p pd=1.96e+06u as=4.625e+11p ps=2.73e+06u
M1007 a_260_74# C1 a_182_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_490_368# A2 Y VPB phighvt w=1.12e+06u l=150000u
+  ad=3.416e+11p pd=2.85e+06u as=0p ps=0u
M1009 VPWR A1 a_490_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

