# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_ls__einvp_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_ls__einvp_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.120000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  2.232000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.410000 1.180000 3.460000 1.550000 ;
    END
  END A
  PIN TE
    ANTENNAGATEAREA  1.167000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.435000 1.180000 8.995000 1.410000 ;
        RECT 8.435000 1.410000 8.765000 1.550000 ;
    END
  END TE
  PIN Z
    ANTENNADIFFAREA  2.328200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.560000 1.720000 4.195000 1.890000 ;
        RECT 0.560000 1.890000 0.890000 2.735000 ;
        RECT 0.625000 0.615000 0.875000 0.840000 ;
        RECT 0.625000 0.840000 3.875000 1.010000 ;
        RECT 1.460000 1.890000 1.790000 2.735000 ;
        RECT 1.545000 0.615000 1.875000 0.840000 ;
        RECT 2.360000 1.890000 2.690000 2.735000 ;
        RECT 2.545000 0.615000 2.875000 0.840000 ;
        RECT 3.260000 1.890000 3.590000 2.735000 ;
        RECT 3.545000 0.595000 3.875000 0.840000 ;
        RECT 3.705000 1.010000 3.875000 1.550000 ;
        RECT 3.705000 1.550000 4.195000 1.720000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 9.120000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000000 0.000000 9.120000 0.245000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.660000 9.310000 3.520000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 9.120000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.120000 0.085000 ;
      RECT 0.000000  3.245000 9.120000 3.415000 ;
      RECT 0.110000  1.820000 0.375000 2.905000 ;
      RECT 0.110000  2.905000 3.960000 3.075000 ;
      RECT 0.115000  0.255000 4.225000 0.425000 ;
      RECT 0.115000  0.425000 0.445000 1.010000 ;
      RECT 1.045000  0.425000 1.375000 0.670000 ;
      RECT 1.070000  2.060000 1.275000 2.905000 ;
      RECT 1.970000  2.060000 2.190000 2.905000 ;
      RECT 2.045000  0.425000 2.375000 0.670000 ;
      RECT 2.875000  2.060000 3.075000 2.905000 ;
      RECT 3.045000  0.425000 3.375000 0.670000 ;
      RECT 3.790000  2.060000 4.940000 2.230000 ;
      RECT 3.790000  2.230000 3.960000 2.905000 ;
      RECT 4.055000  0.425000 4.225000 1.210000 ;
      RECT 4.055000  1.210000 7.885000 1.380000 ;
      RECT 4.160000  2.400000 4.490000 3.245000 ;
      RECT 4.405000  0.085000 4.735000 1.040000 ;
      RECT 4.690000  1.550000 7.560000 1.720000 ;
      RECT 4.690000  1.720000 4.940000 2.060000 ;
      RECT 4.690000  2.230000 4.940000 2.980000 ;
      RECT 4.905000  0.350000 5.155000 1.210000 ;
      RECT 5.140000  1.890000 5.310000 3.245000 ;
      RECT 5.335000  0.085000 5.665000 1.040000 ;
      RECT 5.510000  1.720000 5.760000 2.980000 ;
      RECT 5.845000  0.350000 6.015000 1.210000 ;
      RECT 5.960000  1.890000 6.210000 3.245000 ;
      RECT 6.195000  0.085000 6.525000 1.040000 ;
      RECT 6.410000  1.720000 6.660000 2.980000 ;
      RECT 6.705000  0.350000 6.955000 1.210000 ;
      RECT 6.860000  1.890000 7.110000 3.245000 ;
      RECT 7.125000  0.085000 7.455000 1.040000 ;
      RECT 7.310000  1.720000 7.560000 2.980000 ;
      RECT 7.635000  0.350000 7.885000 1.210000 ;
      RECT 7.775000  1.615000 8.225000 1.820000 ;
      RECT 7.775000  1.820000 8.565000 2.965000 ;
      RECT 8.055000  0.350000 8.505000 1.010000 ;
      RECT 8.055000  1.010000 8.225000 1.615000 ;
      RECT 8.235000  2.965000 8.565000 2.980000 ;
      RECT 8.675000  0.085000 8.935000 1.010000 ;
      RECT 8.765000  1.820000 9.015000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
  END
END sky130_fd_sc_ls__einvp_8
END LIBRARY
