* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
M1000 a_231_74# A2 a_159_74# VNB nshort w=740000u l=150000u
+  ad=2.886e+11p pd=2.26e+06u as=1.554e+11p ps=1.9e+06u
M1001 Y C1 VGND VNB nshort w=740000u l=150000u
+  ad=4.847e+11p pd=4.27e+06u as=4.847e+11p ps=4.27e+06u
M1002 a_159_74# A3 VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 Y C1 a_462_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=3.08e+11p pd=2.79e+06u as=3.696e+11p ps=2.9e+06u
M1004 a_156_368# A1 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=6.72e+11p pd=5.68e+06u as=8.456e+11p ps=5.99e+06u
M1005 Y A1 a_231_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_462_368# B1 a_156_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_156_368# A3 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND B1 Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR A2 a_156_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
