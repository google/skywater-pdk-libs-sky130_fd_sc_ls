* File: sky130_fd_sc_ls__o221ai_4.pex.spice
* Created: Wed Sep  2 11:19:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__O221AI_4%C1 3 5 7 10 12 14 17 19 21 24 26 28 29 30
+ 31 44 47
c81 26 0 1.05417e-19 $X=1.965 $Y=1.765
r82 47 48 25.1478 $w=3.45e-07 $l=1.8e-07 $layer=POLY_cond $X=1.785 $Y=1.557
+ $X2=1.965 $Y2=1.557
r83 46 47 41.2145 $w=3.45e-07 $l=2.95e-07 $layer=POLY_cond $X=1.49 $Y=1.557
+ $X2=1.785 $Y2=1.557
r84 45 46 18.8609 $w=3.45e-07 $l=1.35e-07 $layer=POLY_cond $X=1.355 $Y=1.557
+ $X2=1.49 $Y2=1.557
r85 43 45 16.0667 $w=3.45e-07 $l=1.15e-07 $layer=POLY_cond $X=1.24 $Y=1.557
+ $X2=1.355 $Y2=1.557
r86 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.24
+ $Y=1.515 $X2=1.24 $Y2=1.515
r87 41 43 39.8174 $w=3.45e-07 $l=2.85e-07 $layer=POLY_cond $X=0.955 $Y=1.557
+ $X2=1.24 $Y2=1.557
r88 40 41 4.1913 $w=3.45e-07 $l=3e-08 $layer=POLY_cond $X=0.925 $Y=1.557
+ $X2=0.955 $Y2=1.557
r89 38 40 3.49275 $w=3.45e-07 $l=2.5e-08 $layer=POLY_cond $X=0.9 $Y=1.557
+ $X2=0.925 $Y2=1.557
r90 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.9
+ $Y=1.515 $X2=0.9 $Y2=1.515
r91 36 38 55.1855 $w=3.45e-07 $l=3.95e-07 $layer=POLY_cond $X=0.505 $Y=1.557
+ $X2=0.9 $Y2=1.557
r92 35 36 1.3971 $w=3.45e-07 $l=1e-08 $layer=POLY_cond $X=0.495 $Y=1.557
+ $X2=0.505 $Y2=1.557
r93 31 44 1.07204 $w=4.28e-07 $l=4e-08 $layer=LI1_cond $X=1.2 $Y=1.565 $X2=1.24
+ $Y2=1.565
r94 31 39 8.0403 $w=4.28e-07 $l=3e-07 $layer=LI1_cond $X=1.2 $Y=1.565 $X2=0.9
+ $Y2=1.565
r95 30 39 4.82418 $w=4.28e-07 $l=1.8e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=0.9 $Y2=1.565
r96 29 30 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.24 $Y=1.565
+ $X2=0.72 $Y2=1.565
r97 26 48 22.2839 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.965 $Y=1.765
+ $X2=1.965 $Y2=1.557
r98 26 28 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.965 $Y=1.765
+ $X2=1.965 $Y2=2.4
r99 22 47 22.2839 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.785 $Y=1.35
+ $X2=1.785 $Y2=1.557
r100 22 24 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.785 $Y=1.35
+ $X2=1.785 $Y2=0.79
r101 19 46 22.2839 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.49 $Y=1.765
+ $X2=1.49 $Y2=1.557
r102 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.49 $Y=1.765
+ $X2=1.49 $Y2=2.4
r103 15 45 22.2839 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.355 $Y=1.35
+ $X2=1.355 $Y2=1.557
r104 15 17 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.355 $Y=1.35
+ $X2=1.355 $Y2=0.79
r105 12 41 22.2839 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.955 $Y=1.765
+ $X2=0.955 $Y2=1.557
r106 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.955 $Y=1.765
+ $X2=0.955 $Y2=2.4
r107 8 40 22.2839 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.925 $Y=1.35
+ $X2=0.925 $Y2=1.557
r108 8 10 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.925 $Y=1.35
+ $X2=0.925 $Y2=0.79
r109 5 36 22.2839 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=1.557
r110 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.4
r111 1 35 22.2839 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=1.557
r112 1 3 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=0.79
.ends

.subckt PM_SKY130_FD_SC_LS__O221AI_4%B1 1 3 6 8 10 11 13 14 16 17 19 22 24 26 27
+ 32 37 38 46 50
c122 24 0 1.14201e-19 $X=5.815 $Y=1.765
c123 17 0 9.65396e-20 $X=3.635 $Y=1.185
c124 11 0 9.65396e-20 $X=3.205 $Y=1.185
r125 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.835
+ $Y=1.515 $X2=5.835 $Y2=1.515
r126 43 44 35.298 $w=3.96e-07 $l=2.9e-07 $layer=POLY_cond $X=2.915 $Y=1.475
+ $X2=3.205 $Y2=1.475
r127 38 50 3.01532 $w=5.93e-07 $l=1.5e-07 $layer=LI1_cond $X=5.702 $Y=1.665
+ $X2=5.702 $Y2=1.515
r128 36 46 9.12879 $w=3.96e-07 $l=7.5e-08 $layer=POLY_cond $X=3.39 $Y=1.475
+ $X2=3.465 $Y2=1.475
r129 36 44 22.5177 $w=3.96e-07 $l=1.85e-07 $layer=POLY_cond $X=3.39 $Y=1.475
+ $X2=3.205 $Y2=1.475
r130 35 37 9.70437 $w=5.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.39 $Y=1.615
+ $X2=3.555 $Y2=1.615
r131 35 36 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.39
+ $Y=1.515 $X2=3.39 $Y2=1.515
r132 32 38 2.61328 $w=5.93e-07 $l=1.3e-07 $layer=LI1_cond $X=5.702 $Y=1.795
+ $X2=5.702 $Y2=1.665
r133 32 37 120.695 $w=1.68e-07 $l=1.85e-06 $layer=LI1_cond $X=5.405 $Y=1.795
+ $X2=3.555 $Y2=1.795
r134 30 40 29.8207 $w=3.96e-07 $l=2.45e-07 $layer=POLY_cond $X=2.71 $Y=1.475
+ $X2=2.465 $Y2=1.475
r135 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.71
+ $Y=1.515 $X2=2.71 $Y2=1.515
r136 27 35 2.25675 $w=5.28e-07 $l=1e-07 $layer=LI1_cond $X=3.29 $Y=1.615
+ $X2=3.39 $Y2=1.615
r137 27 29 13.0892 $w=5.28e-07 $l=5.8e-07 $layer=LI1_cond $X=3.29 $Y=1.615
+ $X2=2.71 $Y2=1.615
r138 24 49 52.2586 $w=2.99e-07 $l=2.59808e-07 $layer=POLY_cond $X=5.815 $Y=1.765
+ $X2=5.835 $Y2=1.515
r139 24 26 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.815 $Y=1.765
+ $X2=5.815 $Y2=2.4
r140 20 49 38.5562 $w=2.99e-07 $l=1.88348e-07 $layer=POLY_cond $X=5.785 $Y=1.35
+ $X2=5.835 $Y2=1.515
r141 20 22 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.785 $Y=1.35
+ $X2=5.785 $Y2=0.74
r142 17 46 20.6919 $w=3.96e-07 $l=3.6524e-07 $layer=POLY_cond $X=3.635 $Y=1.185
+ $X2=3.465 $Y2=1.475
r143 17 19 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=3.635 $Y=1.185
+ $X2=3.635 $Y2=0.74
r144 14 46 25.6164 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=3.465 $Y=1.765
+ $X2=3.465 $Y2=1.475
r145 14 16 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.465 $Y=1.765
+ $X2=3.465 $Y2=2.4
r146 11 44 25.6164 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=3.205 $Y=1.185
+ $X2=3.205 $Y2=1.475
r147 11 13 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=3.205 $Y=1.185
+ $X2=3.205 $Y2=0.74
r148 8 43 25.6164 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.915 $Y=1.765
+ $X2=2.915 $Y2=1.475
r149 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.915 $Y=1.765
+ $X2=2.915 $Y2=2.4
r150 4 43 17.0404 $w=3.96e-07 $l=1.4e-07 $layer=POLY_cond $X=2.775 $Y=1.475
+ $X2=2.915 $Y2=1.475
r151 4 30 7.91162 $w=3.96e-07 $l=6.5e-08 $layer=POLY_cond $X=2.775 $Y=1.475
+ $X2=2.71 $Y2=1.475
r152 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.775 $Y=1.35
+ $X2=2.775 $Y2=0.74
r153 1 40 25.6164 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.465 $Y=1.765
+ $X2=2.465 $Y2=1.475
r154 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.465 $Y=1.765
+ $X2=2.465 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__O221AI_4%B2 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 26 41
c83 41 0 3.38438e-19 $X=5.315 $Y=1.492
c84 26 0 1.14201e-19 $X=5.04 $Y=1.295
c85 16 0 1.90514e-19 $X=4.925 $Y=1.22
c86 4 0 4.22428e-20 $X=4.065 $Y=1.22
r87 41 42 4.60143 $w=4.19e-07 $l=4e-08 $layer=POLY_cond $X=5.315 $Y=1.492
+ $X2=5.355 $Y2=1.492
r88 39 41 32.7852 $w=4.19e-07 $l=2.85e-07 $layer=POLY_cond $X=5.03 $Y=1.492
+ $X2=5.315 $Y2=1.492
r89 39 40 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=5.03
+ $Y=1.385 $X2=5.03 $Y2=1.385
r90 37 39 12.0788 $w=4.19e-07 $l=1.05e-07 $layer=POLY_cond $X=4.925 $Y=1.492
+ $X2=5.03 $Y2=1.492
r91 36 37 12.6539 $w=4.19e-07 $l=1.1e-07 $layer=POLY_cond $X=4.815 $Y=1.492
+ $X2=4.925 $Y2=1.492
r92 35 36 36.8115 $w=4.19e-07 $l=3.2e-07 $layer=POLY_cond $X=4.495 $Y=1.492
+ $X2=4.815 $Y2=1.492
r93 34 35 14.9547 $w=4.19e-07 $l=1.3e-07 $layer=POLY_cond $X=4.365 $Y=1.492
+ $X2=4.495 $Y2=1.492
r94 32 34 1.72554 $w=4.19e-07 $l=1.5e-08 $layer=POLY_cond $X=4.35 $Y=1.492
+ $X2=4.365 $Y2=1.492
r95 32 33 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=4.35
+ $Y=1.385 $X2=4.35 $Y2=1.385
r96 30 32 32.7852 $w=4.19e-07 $l=2.85e-07 $layer=POLY_cond $X=4.065 $Y=1.492
+ $X2=4.35 $Y2=1.492
r97 26 40 0.320123 $w=3.58e-07 $l=1e-08 $layer=LI1_cond $X=5.04 $Y=1.36 $X2=5.03
+ $Y2=1.36
r98 25 40 15.0458 $w=3.58e-07 $l=4.7e-07 $layer=LI1_cond $X=4.56 $Y=1.36
+ $X2=5.03 $Y2=1.36
r99 25 33 6.72258 $w=3.58e-07 $l=2.1e-07 $layer=LI1_cond $X=4.56 $Y=1.36
+ $X2=4.35 $Y2=1.36
r100 22 42 27.0004 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=5.355 $Y=1.22
+ $X2=5.355 $Y2=1.492
r101 22 24 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.355 $Y=1.22
+ $X2=5.355 $Y2=0.74
r102 19 41 27.0004 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=5.315 $Y=1.765
+ $X2=5.315 $Y2=1.492
r103 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.315 $Y=1.765
+ $X2=5.315 $Y2=2.4
r104 16 37 27.0004 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=4.925 $Y=1.22
+ $X2=4.925 $Y2=1.492
r105 16 18 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.925 $Y=1.22
+ $X2=4.925 $Y2=0.74
r106 13 36 27.0004 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=4.815 $Y=1.765
+ $X2=4.815 $Y2=1.492
r107 13 15 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.815 $Y=1.765
+ $X2=4.815 $Y2=2.4
r108 10 35 27.0004 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=4.495 $Y=1.22
+ $X2=4.495 $Y2=1.492
r109 10 12 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.495 $Y=1.22
+ $X2=4.495 $Y2=0.74
r110 7 34 27.0004 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=4.365 $Y=1.765
+ $X2=4.365 $Y2=1.492
r111 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.365 $Y=1.765
+ $X2=4.365 $Y2=2.4
r112 4 30 27.0004 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=4.065 $Y=1.22
+ $X2=4.065 $Y2=1.492
r113 4 6 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.065 $Y=1.22
+ $X2=4.065 $Y2=0.74
r114 1 30 17.2554 $w=4.19e-07 $l=3.39822e-07 $layer=POLY_cond $X=3.915 $Y=1.765
+ $X2=4.065 $Y2=1.492
r115 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.915 $Y=1.765
+ $X2=3.915 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__O221AI_4%A1 3 5 7 10 12 14 15 17 20 22 24 27 30 35
+ 36 37 38 55 69 71 72
c116 72 0 1.04264e-20 $X=8.455 $Y=1.435
c117 55 0 1.46492e-19 $X=9.57 $Y=1.512
c118 3 0 1.43357e-20 $X=6.285 $Y=0.74
r119 71 72 1.70704 $w=6.88e-07 $l=5.5e-08 $layer=LI1_cond $X=8.4 $Y=1.435
+ $X2=8.455 $Y2=1.435
r120 55 56 1.73381 $w=4.17e-07 $l=1.5e-08 $layer=POLY_cond $X=9.57 $Y=1.512
+ $X2=9.585 $Y2=1.512
r121 53 55 16.7602 $w=4.17e-07 $l=1.45e-07 $layer=POLY_cond $X=9.425 $Y=1.512
+ $X2=9.57 $Y2=1.512
r122 53 54 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=9.425
+ $Y=1.425 $X2=9.425 $Y2=1.425
r123 51 53 31.2086 $w=4.17e-07 $l=2.7e-07 $layer=POLY_cond $X=9.155 $Y=1.512
+ $X2=9.425 $Y2=1.512
r124 50 51 4.04556 $w=4.17e-07 $l=3.5e-08 $layer=POLY_cond $X=9.12 $Y=1.512
+ $X2=9.155 $Y2=1.512
r125 48 50 43.3453 $w=4.17e-07 $l=3.75e-07 $layer=POLY_cond $X=8.745 $Y=1.512
+ $X2=9.12 $Y2=1.512
r126 48 49 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=8.745
+ $Y=1.425 $X2=8.745 $Y2=1.425
r127 46 48 8.66906 $w=4.17e-07 $l=7.5e-08 $layer=POLY_cond $X=8.67 $Y=1.512
+ $X2=8.745 $Y2=1.512
r128 45 46 1.73381 $w=4.17e-07 $l=1.5e-08 $layer=POLY_cond $X=8.655 $Y=1.512
+ $X2=8.67 $Y2=1.512
r129 38 54 9.54563 $w=5.18e-07 $l=4.15e-07 $layer=LI1_cond $X=9.84 $Y=1.52
+ $X2=9.425 $Y2=1.52
r130 37 54 1.4951 $w=5.18e-07 $l=6.5e-08 $layer=LI1_cond $X=9.36 $Y=1.52
+ $X2=9.425 $Y2=1.52
r131 36 37 11.0407 $w=5.18e-07 $l=4.8e-07 $layer=LI1_cond $X=8.88 $Y=1.52
+ $X2=9.36 $Y2=1.52
r132 36 49 3.1052 $w=5.18e-07 $l=1.35e-07 $layer=LI1_cond $X=8.88 $Y=1.52
+ $X2=8.745 $Y2=1.52
r133 35 71 0.260017 $w=6.88e-07 $l=1.5e-08 $layer=LI1_cond $X=8.385 $Y=1.435
+ $X2=8.4 $Y2=1.435
r134 35 69 9.6141 $w=6.88e-07 $l=1e-07 $layer=LI1_cond $X=8.385 $Y=1.435
+ $X2=8.285 $Y2=1.435
r135 35 49 6.32541 $w=5.18e-07 $l=2.75e-07 $layer=LI1_cond $X=8.47 $Y=1.52
+ $X2=8.745 $Y2=1.52
r136 35 72 0.345023 $w=5.18e-07 $l=1.5e-08 $layer=LI1_cond $X=8.47 $Y=1.52
+ $X2=8.455 $Y2=1.52
r137 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.375
+ $Y=1.425 $X2=6.375 $Y2=1.425
r138 30 33 10.2349 $w=2.98e-07 $l=3.29014e-07 $layer=LI1_cond $X=6.575 $Y=1.175
+ $X2=6.392 $Y2=1.425
r139 30 69 111.561 $w=1.68e-07 $l=1.71e-06 $layer=LI1_cond $X=6.575 $Y=1.175
+ $X2=8.285 $Y2=1.175
r140 25 56 26.8826 $w=1.5e-07 $l=2.52e-07 $layer=POLY_cond $X=9.585 $Y=1.26
+ $X2=9.585 $Y2=1.512
r141 25 27 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=9.585 $Y=1.26
+ $X2=9.585 $Y2=0.74
r142 22 55 26.8826 $w=1.5e-07 $l=2.53e-07 $layer=POLY_cond $X=9.57 $Y=1.765
+ $X2=9.57 $Y2=1.512
r143 22 24 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=9.57 $Y=1.765
+ $X2=9.57 $Y2=2.4
r144 18 51 26.8826 $w=1.5e-07 $l=2.52e-07 $layer=POLY_cond $X=9.155 $Y=1.26
+ $X2=9.155 $Y2=1.512
r145 18 20 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=9.155 $Y=1.26
+ $X2=9.155 $Y2=0.74
r146 15 50 26.8826 $w=1.5e-07 $l=2.53e-07 $layer=POLY_cond $X=9.12 $Y=1.765
+ $X2=9.12 $Y2=1.512
r147 15 17 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=9.12 $Y=1.765
+ $X2=9.12 $Y2=2.4
r148 12 46 26.8826 $w=1.5e-07 $l=2.53e-07 $layer=POLY_cond $X=8.67 $Y=1.765
+ $X2=8.67 $Y2=1.512
r149 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.67 $Y=1.765
+ $X2=8.67 $Y2=2.4
r150 8 45 26.8826 $w=1.5e-07 $l=2.52e-07 $layer=POLY_cond $X=8.655 $Y=1.26
+ $X2=8.655 $Y2=1.512
r151 8 10 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=8.655 $Y=1.26
+ $X2=8.655 $Y2=0.74
r152 5 34 69.1012 $w=2.78e-07 $l=3.44964e-07 $layer=POLY_cond $X=6.365 $Y=1.765
+ $X2=6.375 $Y2=1.425
r153 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.365 $Y=1.765
+ $X2=6.365 $Y2=2.4
r154 1 34 38.7595 $w=2.78e-07 $l=2.05122e-07 $layer=POLY_cond $X=6.285 $Y=1.26
+ $X2=6.375 $Y2=1.425
r155 1 3 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=6.285 $Y=1.26
+ $X2=6.285 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__O221AI_4%A2 3 5 7 10 12 14 15 17 20 24 26 28 29 30
+ 31 47
c86 31 0 1.46492e-19 $X=7.92 $Y=1.665
c87 26 0 1.88367e-19 $X=8.22 $Y=1.765
c88 15 0 1.04264e-20 $X=7.77 $Y=1.765
r89 47 48 0.656676 $w=3.67e-07 $l=5e-09 $layer=POLY_cond $X=8.215 $Y=1.557
+ $X2=8.22 $Y2=1.557
r90 46 47 56.4741 $w=3.67e-07 $l=4.3e-07 $layer=POLY_cond $X=7.785 $Y=1.557
+ $X2=8.215 $Y2=1.557
r91 45 46 1.97003 $w=3.67e-07 $l=1.5e-08 $layer=POLY_cond $X=7.77 $Y=1.557
+ $X2=7.785 $Y2=1.557
r92 43 45 10.5068 $w=3.67e-07 $l=8e-08 $layer=POLY_cond $X=7.69 $Y=1.557
+ $X2=7.77 $Y2=1.557
r93 43 44 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.69
+ $Y=1.515 $X2=7.69 $Y2=1.515
r94 41 43 48.594 $w=3.67e-07 $l=3.7e-07 $layer=POLY_cond $X=7.32 $Y=1.557
+ $X2=7.69 $Y2=1.557
r95 40 41 4.59673 $w=3.67e-07 $l=3.5e-08 $layer=POLY_cond $X=7.285 $Y=1.557
+ $X2=7.32 $Y2=1.557
r96 38 40 36.1172 $w=3.67e-07 $l=2.75e-07 $layer=POLY_cond $X=7.01 $Y=1.557
+ $X2=7.285 $Y2=1.557
r97 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.01
+ $Y=1.515 $X2=7.01 $Y2=1.515
r98 36 38 18.3869 $w=3.67e-07 $l=1.4e-07 $layer=POLY_cond $X=6.87 $Y=1.557
+ $X2=7.01 $Y2=1.557
r99 35 36 1.97003 $w=3.67e-07 $l=1.5e-08 $layer=POLY_cond $X=6.855 $Y=1.557
+ $X2=6.87 $Y2=1.557
r100 31 44 7.5732 $w=3.48e-07 $l=2.3e-07 $layer=LI1_cond $X=7.92 $Y=1.605
+ $X2=7.69 $Y2=1.605
r101 30 44 8.23174 $w=3.48e-07 $l=2.5e-07 $layer=LI1_cond $X=7.44 $Y=1.605
+ $X2=7.69 $Y2=1.605
r102 30 39 14.1586 $w=3.48e-07 $l=4.3e-07 $layer=LI1_cond $X=7.44 $Y=1.605
+ $X2=7.01 $Y2=1.605
r103 29 39 1.64635 $w=3.48e-07 $l=5e-08 $layer=LI1_cond $X=6.96 $Y=1.605
+ $X2=7.01 $Y2=1.605
r104 26 48 23.77 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=8.22 $Y=1.765
+ $X2=8.22 $Y2=1.557
r105 26 28 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.22 $Y=1.765
+ $X2=8.22 $Y2=2.4
r106 22 47 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=8.215 $Y=1.35
+ $X2=8.215 $Y2=1.557
r107 22 24 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=8.215 $Y=1.35
+ $X2=8.215 $Y2=0.74
r108 18 46 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.785 $Y=1.35
+ $X2=7.785 $Y2=1.557
r109 18 20 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.785 $Y=1.35
+ $X2=7.785 $Y2=0.74
r110 15 45 23.77 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=7.77 $Y=1.765
+ $X2=7.77 $Y2=1.557
r111 15 17 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.77 $Y=1.765
+ $X2=7.77 $Y2=2.4
r112 12 41 23.77 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=7.32 $Y=1.765
+ $X2=7.32 $Y2=1.557
r113 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.32 $Y=1.765
+ $X2=7.32 $Y2=2.4
r114 8 40 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.285 $Y=1.35
+ $X2=7.285 $Y2=1.557
r115 8 10 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.285 $Y=1.35
+ $X2=7.285 $Y2=0.74
r116 5 36 23.77 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=6.87 $Y=1.765
+ $X2=6.87 $Y2=1.557
r117 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.87 $Y=1.765
+ $X2=6.87 $Y2=2.4
r118 1 35 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.855 $Y=1.35
+ $X2=6.855 $Y2=1.557
r119 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.855 $Y=1.35
+ $X2=6.855 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__O221AI_4%VPWR 1 2 3 4 5 6 7 22 24 30 34 38 42 46 48
+ 50 54 56 61 66 71 76 84 93 96 99 102 105 109
c131 46 0 1.88367e-19 $X=8.895 $Y=2.455
r132 108 109 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r133 105 106 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r134 102 103 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r135 99 100 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r136 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r137 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r138 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r139 88 109 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=9.84 $Y2=3.33
r140 88 106 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=8.88 $Y2=3.33
r141 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r142 85 105 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.98 $Y=3.33
+ $X2=8.855 $Y2=3.33
r143 85 87 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=8.98 $Y=3.33
+ $X2=9.36 $Y2=3.33
r144 84 108 4.0045 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=9.71 $Y=3.33
+ $X2=9.895 $Y2=3.33
r145 84 87 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=9.71 $Y=3.33
+ $X2=9.36 $Y2=3.33
r146 83 106 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=8.88 $Y2=3.33
r147 82 83 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r148 80 83 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=8.4 $Y2=3.33
r149 80 103 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6 $Y2=3.33
r150 79 82 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=6.48 $Y=3.33
+ $X2=8.4 $Y2=3.33
r151 79 80 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r152 77 102 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.255 $Y=3.33
+ $X2=6.09 $Y2=3.33
r153 77 79 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=6.255 $Y=3.33
+ $X2=6.48 $Y2=3.33
r154 76 105 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.73 $Y=3.33
+ $X2=8.855 $Y2=3.33
r155 76 82 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=8.73 $Y=3.33
+ $X2=8.4 $Y2=3.33
r156 75 100 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r157 74 75 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r158 72 99 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.355 $Y=3.33
+ $X2=3.19 $Y2=3.33
r159 72 74 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=3.355 $Y=3.33
+ $X2=3.6 $Y2=3.33
r160 71 102 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.925 $Y=3.33
+ $X2=6.09 $Y2=3.33
r161 71 74 151.684 $w=1.68e-07 $l=2.325e-06 $layer=LI1_cond $X=5.925 $Y=3.33
+ $X2=3.6 $Y2=3.33
r162 70 100 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r163 70 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r164 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r165 67 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.355 $Y=3.33
+ $X2=2.19 $Y2=3.33
r166 67 69 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.355 $Y=3.33
+ $X2=2.64 $Y2=3.33
r167 66 99 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.025 $Y=3.33
+ $X2=3.19 $Y2=3.33
r168 66 69 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=3.025 $Y=3.33
+ $X2=2.64 $Y2=3.33
r169 65 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r170 65 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r171 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r172 62 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.395 $Y=3.33
+ $X2=1.23 $Y2=3.33
r173 62 64 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.395 $Y=3.33
+ $X2=1.68 $Y2=3.33
r174 61 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.025 $Y=3.33
+ $X2=2.19 $Y2=3.33
r175 61 64 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.025 $Y=3.33
+ $X2=1.68 $Y2=3.33
r176 60 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r177 60 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r178 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r179 57 90 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.182 $Y2=3.33
r180 57 59 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.72 $Y2=3.33
r181 56 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.065 $Y=3.33
+ $X2=1.23 $Y2=3.33
r182 56 59 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.065 $Y=3.33
+ $X2=0.72 $Y2=3.33
r183 54 103 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=6 $Y2=3.33
r184 54 75 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=3.6 $Y2=3.33
r185 50 53 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=9.835 $Y=2.115
+ $X2=9.835 $Y2=2.815
r186 48 108 3.13866 $w=2.5e-07 $l=1.11018e-07 $layer=LI1_cond $X=9.835 $Y=3.245
+ $X2=9.895 $Y2=3.33
r187 48 53 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=9.835 $Y=3.245
+ $X2=9.835 $Y2=2.815
r188 44 105 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.855 $Y=3.245
+ $X2=8.855 $Y2=3.33
r189 44 46 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=8.855 $Y=3.245
+ $X2=8.855 $Y2=2.455
r190 40 102 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.09 $Y=3.245
+ $X2=6.09 $Y2=3.33
r191 40 42 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=6.09 $Y=3.245
+ $X2=6.09 $Y2=2.475
r192 36 99 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.19 $Y=3.245
+ $X2=3.19 $Y2=3.33
r193 36 38 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.19 $Y=3.245
+ $X2=3.19 $Y2=2.815
r194 32 96 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.19 $Y=3.245
+ $X2=2.19 $Y2=3.33
r195 32 34 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=2.19 $Y=3.245
+ $X2=2.19 $Y2=2.475
r196 28 93 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.23 $Y=3.245
+ $X2=1.23 $Y2=3.33
r197 28 30 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=1.23 $Y=3.245
+ $X2=1.23 $Y2=2.455
r198 24 27 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=0.24 $Y=2.115
+ $X2=0.24 $Y2=2.815
r199 22 90 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.182 $Y2=3.33
r200 22 27 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.24 $Y2=2.815
r201 7 53 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=9.645
+ $Y=1.84 $X2=9.795 $Y2=2.815
r202 7 50 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=9.645
+ $Y=1.84 $X2=9.795 $Y2=2.115
r203 6 46 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=8.745
+ $Y=1.84 $X2=8.895 $Y2=2.455
r204 5 42 300 $w=1.7e-07 $l=7.28166e-07 $layer=licon1_PDIFF $count=2 $X=5.89
+ $Y=1.84 $X2=6.09 $Y2=2.475
r205 4 38 600 $w=1.7e-07 $l=1.07034e-06 $layer=licon1_PDIFF $count=1 $X=2.99
+ $Y=1.84 $X2=3.19 $Y2=2.815
r206 3 34 300 $w=1.7e-07 $l=7.06028e-07 $layer=licon1_PDIFF $count=2 $X=2.04
+ $Y=1.84 $X2=2.19 $Y2=2.475
r207 2 30 300 $w=1.7e-07 $l=7.07972e-07 $layer=licon1_PDIFF $count=2 $X=1.03
+ $Y=1.84 $X2=1.23 $Y2=2.455
r208 1 27 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r209 1 24 400 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_LS__O221AI_4%Y 1 2 3 4 5 6 7 8 27 29 31 33 34 35 39 45
+ 47 51 53 57 59 61 67 69 70 74 76 78 79
c144 53 0 1.6985e-19 $X=4.925 $Y=2.135
c145 47 0 1.68588e-19 $X=4.055 $Y=2.135
r146 83 84 0.624041 $w=3.91e-07 $l=2e-08 $layer=LI1_cond $X=7.052 $Y=2.115
+ $X2=7.052 $Y2=2.135
r147 81 83 2.49616 $w=3.91e-07 $l=8e-08 $layer=LI1_cond $X=7.052 $Y=2.035
+ $X2=7.052 $Y2=2.115
r148 79 84 8.42455 $w=3.91e-07 $l=2.7e-07 $layer=LI1_cond $X=7.052 $Y=2.405
+ $X2=7.052 $Y2=2.135
r149 71 72 4.60977 $w=2.48e-07 $l=1e-07 $layer=LI1_cond $X=1.7 $Y=2.035 $X2=1.7
+ $Y2=2.135
r150 69 71 2.30489 $w=2.48e-07 $l=5e-08 $layer=LI1_cond $X=1.7 $Y=1.985 $X2=1.7
+ $Y2=2.035
r151 69 70 8.79328 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=1.7 $Y=1.985
+ $X2=1.7 $Y2=1.82
r152 62 81 5.64031 $w=1.7e-07 $l=2.08e-07 $layer=LI1_cond $X=7.26 $Y=2.035
+ $X2=7.052 $Y2=2.035
r153 61 78 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.83 $Y=2.035
+ $X2=7.995 $Y2=2.035
r154 61 62 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=7.83 $Y=2.035
+ $X2=7.26 $Y2=2.035
r155 60 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.255 $Y=2.135
+ $X2=5.09 $Y2=2.135
r156 59 84 5.64031 $w=1.7e-07 $l=2.07e-07 $layer=LI1_cond $X=6.845 $Y=2.135
+ $X2=7.052 $Y2=2.135
r157 59 60 103.733 $w=1.68e-07 $l=1.59e-06 $layer=LI1_cond $X=6.845 $Y=2.135
+ $X2=5.255 $Y2=2.135
r158 55 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.09 $Y=2.22
+ $X2=5.09 $Y2=2.135
r159 55 57 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=5.09 $Y=2.22
+ $X2=5.09 $Y2=2.57
r160 54 74 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.225 $Y=2.135
+ $X2=4.14 $Y2=2.135
r161 53 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.925 $Y=2.135
+ $X2=5.09 $Y2=2.135
r162 53 54 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=4.925 $Y=2.135
+ $X2=4.225 $Y2=2.135
r163 49 74 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.14 $Y=2.22
+ $X2=4.14 $Y2=2.135
r164 49 51 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=4.14 $Y=2.22
+ $X2=4.14 $Y2=2.57
r165 48 72 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.825 $Y=2.135
+ $X2=1.7 $Y2=2.135
r166 47 74 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.055 $Y=2.135
+ $X2=4.14 $Y2=2.135
r167 47 48 145.487 $w=1.68e-07 $l=2.23e-06 $layer=LI1_cond $X=4.055 $Y=2.135
+ $X2=1.825 $Y2=2.135
r168 43 72 3.91831 $w=2.48e-07 $l=8.5e-08 $layer=LI1_cond $X=1.7 $Y=2.22 $X2=1.7
+ $Y2=2.135
r169 43 45 8.29759 $w=2.48e-07 $l=1.8e-07 $layer=LI1_cond $X=1.7 $Y=2.22 $X2=1.7
+ $Y2=2.4
r170 41 67 3.64284 $w=2.55e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.66 $Y=1.18
+ $X2=1.575 $Y2=1.095
r171 41 70 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=1.66 $Y=1.18
+ $X2=1.66 $Y2=1.82
r172 37 67 3.64284 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=1.575 $Y=1.01
+ $X2=1.575 $Y2=1.095
r173 37 39 11.1855 $w=3.38e-07 $l=3.3e-07 $layer=LI1_cond $X=1.575 $Y=1.01
+ $X2=1.575 $Y2=0.68
r174 36 66 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=2.035
+ $X2=0.73 $Y2=2.035
r175 35 71 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.575 $Y=2.035
+ $X2=1.7 $Y2=2.035
r176 35 36 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.575 $Y=2.035
+ $X2=0.895 $Y2=2.035
r177 33 67 2.83584 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=1.405 $Y=1.095
+ $X2=1.575 $Y2=1.095
r178 33 34 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.405 $Y=1.095
+ $X2=0.875 $Y2=1.095
r179 29 66 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=2.12 $X2=0.73
+ $Y2=2.035
r180 29 31 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=0.73 $Y=2.12
+ $X2=0.73 $Y2=2.815
r181 25 34 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.71 $Y=1.01
+ $X2=0.875 $Y2=1.095
r182 25 27 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=0.71 $Y=1.01
+ $X2=0.71 $Y2=0.68
r183 8 78 300 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=2 $X=7.845
+ $Y=1.84 $X2=7.995 $Y2=2.115
r184 7 83 300 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=2 $X=6.945
+ $Y=1.84 $X2=7.095 $Y2=2.115
r185 6 76 600 $w=1.7e-07 $l=3.82132e-07 $layer=licon1_PDIFF $count=1 $X=4.89
+ $Y=1.84 $X2=5.09 $Y2=2.135
r186 6 57 600 $w=1.7e-07 $l=8.23954e-07 $layer=licon1_PDIFF $count=1 $X=4.89
+ $Y=1.84 $X2=5.09 $Y2=2.57
r187 5 74 600 $w=1.7e-07 $l=3.62319e-07 $layer=licon1_PDIFF $count=1 $X=3.99
+ $Y=1.84 $X2=4.14 $Y2=2.135
r188 5 51 600 $w=1.7e-07 $l=8.01499e-07 $layer=licon1_PDIFF $count=1 $X=3.99
+ $Y=1.84 $X2=4.14 $Y2=2.57
r189 4 69 600 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=1.565
+ $Y=1.84 $X2=1.74 $Y2=1.985
r190 4 45 300 $w=1.7e-07 $l=6.41561e-07 $layer=licon1_PDIFF $count=2 $X=1.565
+ $Y=1.84 $X2=1.74 $Y2=2.4
r191 3 66 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.84 $X2=0.73 $Y2=2.115
r192 3 31 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.84 $X2=0.73 $Y2=2.815
r193 2 39 91 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_NDIFF $count=2 $X=1.43
+ $Y=0.42 $X2=1.57 $Y2=0.68
r194 1 27 91 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_NDIFF $count=2 $X=0.57
+ $Y=0.42 $X2=0.71 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_LS__O221AI_4%A_508_368# 1 2 3 4 15 17 18 19 20 23 25 29
+ 32 35
c67 32 0 1.05417e-19 $X=2.69 $Y=2.475
r68 27 29 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=5.59 $Y=2.905
+ $X2=5.59 $Y2=2.475
r69 26 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.755 $Y=2.99
+ $X2=4.59 $Y2=2.99
r70 25 27 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.425 $Y=2.99
+ $X2=5.59 $Y2=2.905
r71 25 26 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.425 $Y=2.99
+ $X2=4.755 $Y2=2.99
r72 21 35 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.59 $Y=2.905
+ $X2=4.59 $Y2=2.99
r73 21 23 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=4.59 $Y=2.905
+ $X2=4.59 $Y2=2.475
r74 19 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.425 $Y=2.99
+ $X2=4.59 $Y2=2.99
r75 19 20 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=4.425 $Y=2.99
+ $X2=3.855 $Y2=2.99
r76 18 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.69 $Y=2.905
+ $X2=3.855 $Y2=2.99
r77 17 34 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.69 $Y=2.56 $X2=3.69
+ $Y2=2.475
r78 17 18 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=3.69 $Y=2.56
+ $X2=3.69 $Y2=2.905
r79 16 32 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.855 $Y=2.475
+ $X2=2.69 $Y2=2.475
r80 15 34 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.525 $Y=2.475
+ $X2=3.69 $Y2=2.475
r81 15 16 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.525 $Y=2.475
+ $X2=2.855 $Y2=2.475
r82 4 29 300 $w=1.7e-07 $l=7.28166e-07 $layer=licon1_PDIFF $count=2 $X=5.39
+ $Y=1.84 $X2=5.59 $Y2=2.475
r83 3 23 300 $w=1.7e-07 $l=7.06028e-07 $layer=licon1_PDIFF $count=2 $X=4.44
+ $Y=1.84 $X2=4.59 $Y2=2.475
r84 2 34 300 $w=1.7e-07 $l=7.06028e-07 $layer=licon1_PDIFF $count=2 $X=3.54
+ $Y=1.84 $X2=3.69 $Y2=2.475
r85 1 32 300 $w=1.7e-07 $l=7.06028e-07 $layer=licon1_PDIFF $count=2 $X=2.54
+ $Y=1.84 $X2=2.69 $Y2=2.475
.ends

.subckt PM_SKY130_FD_SC_LS__O221AI_4%A_1288_368# 1 2 3 4 13 17 19 21 24 25 27 29
+ 32 34
r55 32 33 6.69279 $w=3.19e-07 $l=1.75e-07 $layer=LI1_cond $X=6.592 $Y=2.815
+ $X2=6.592 $Y2=2.99
r56 27 38 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.345 $Y=2.12
+ $X2=9.345 $Y2=2.035
r57 27 29 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=9.345 $Y=2.12
+ $X2=9.345 $Y2=2.815
r58 26 36 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.53 $Y=2.035
+ $X2=8.445 $Y2=2.035
r59 25 38 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.18 $Y=2.035
+ $X2=9.345 $Y2=2.035
r60 25 26 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=9.18 $Y=2.035
+ $X2=8.53 $Y2=2.035
r61 22 24 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=8.445 $Y=2.905
+ $X2=8.445 $Y2=2.815
r62 21 36 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.445 $Y=2.12
+ $X2=8.445 $Y2=2.035
r63 21 24 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=8.445 $Y=2.12
+ $X2=8.445 $Y2=2.815
r64 20 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.63 $Y=2.99
+ $X2=7.545 $Y2=2.99
r65 19 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.36 $Y=2.99
+ $X2=8.445 $Y2=2.905
r66 19 20 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=8.36 $Y=2.99
+ $X2=7.63 $Y2=2.99
r67 15 34 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.545 $Y=2.905
+ $X2=7.545 $Y2=2.99
r68 15 17 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=7.545 $Y=2.905
+ $X2=7.545 $Y2=2.455
r69 14 33 4.42298 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=6.76 $Y=2.99
+ $X2=6.592 $Y2=2.99
r70 13 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.46 $Y=2.99
+ $X2=7.545 $Y2=2.99
r71 13 14 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=7.46 $Y=2.99 $X2=6.76
+ $Y2=2.99
r72 4 38 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=9.195
+ $Y=1.84 $X2=9.345 $Y2=2.115
r73 4 29 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=9.195
+ $Y=1.84 $X2=9.345 $Y2=2.815
r74 3 36 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=8.295
+ $Y=1.84 $X2=8.445 $Y2=2.115
r75 3 24 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=8.295
+ $Y=1.84 $X2=8.445 $Y2=2.815
r76 2 17 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=7.395
+ $Y=1.84 $X2=7.545 $Y2=2.455
r77 1 32 600 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=6.44
+ $Y=1.84 $X2=6.59 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_LS__O221AI_4%A_27_84# 1 2 3 4 5 6 7 24 26 27 30 32 37 38
+ 39 40 46 49 50 57 58
c80 57 0 1.90514e-19 $X=5.57 $Y=0.91
c81 40 0 4.22428e-20 $X=3.685 $Y=1.095
r82 57 58 7.05875 $w=2.78e-07 $l=1.65e-07 $layer=LI1_cond $X=5.57 $Y=0.91
+ $X2=5.405 $Y2=0.91
r83 53 54 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=3.85 $Y=0.95
+ $X2=3.85 $Y2=1.095
r84 50 53 2.09535 $w=3.28e-07 $l=6e-08 $layer=LI1_cond $X=3.85 $Y=0.89 $X2=3.85
+ $Y2=0.95
r85 48 49 8.69073 $w=4.08e-07 $l=1.65e-07 $layer=LI1_cond $X=2.99 $Y=0.975
+ $X2=3.155 $Y2=0.975
r86 45 58 33.3728 $w=2.38e-07 $l=6.95e-07 $layer=LI1_cond $X=4.71 $Y=0.89
+ $X2=5.405 $Y2=0.89
r87 43 50 2.60351 $w=2.4e-07 $l=1.65e-07 $layer=LI1_cond $X=4.015 $Y=0.89
+ $X2=3.85 $Y2=0.89
r88 43 45 33.3728 $w=2.38e-07 $l=6.95e-07 $layer=LI1_cond $X=4.015 $Y=0.89
+ $X2=4.71 $Y2=0.89
r89 40 54 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.685 $Y=1.095
+ $X2=3.85 $Y2=1.095
r90 40 49 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.685 $Y=1.095
+ $X2=3.155 $Y2=1.095
r91 38 48 1.12433 $w=4.08e-07 $l=4e-08 $layer=LI1_cond $X=2.95 $Y=0.975 $X2=2.99
+ $Y2=0.975
r92 38 39 22.0651 $w=4.08e-07 $l=7.85e-07 $layer=LI1_cond $X=2.95 $Y=0.975
+ $X2=2.165 $Y2=0.975
r93 35 39 7.35087 $w=4.1e-07 $l=2.60096e-07 $layer=LI1_cond $X=2.04 $Y=0.77
+ $X2=2.165 $Y2=0.975
r94 35 37 9.45003 $w=2.48e-07 $l=2.05e-07 $layer=LI1_cond $X=2.04 $Y=0.77
+ $X2=2.04 $Y2=0.565
r95 34 37 6.45368 $w=2.48e-07 $l=1.4e-07 $layer=LI1_cond $X=2.04 $Y=0.425
+ $X2=2.04 $Y2=0.565
r96 33 46 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.235 $Y=0.34
+ $X2=1.14 $Y2=0.34
r97 32 34 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.915 $Y=0.34
+ $X2=2.04 $Y2=0.425
r98 32 33 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.915 $Y=0.34
+ $X2=1.235 $Y2=0.34
r99 28 46 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=0.425
+ $X2=1.14 $Y2=0.34
r100 28 30 13.7177 $w=1.88e-07 $l=2.35e-07 $layer=LI1_cond $X=1.14 $Y=0.425
+ $X2=1.14 $Y2=0.66
r101 26 46 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.045 $Y=0.34
+ $X2=1.14 $Y2=0.34
r102 26 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.045 $Y=0.34
+ $X2=0.375 $Y2=0.34
r103 22 27 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.245 $Y=0.425
+ $X2=0.375 $Y2=0.34
r104 22 24 6.20546 $w=2.58e-07 $l=1.4e-07 $layer=LI1_cond $X=0.245 $Y=0.425
+ $X2=0.245 $Y2=0.565
r105 7 57 182 $w=1.7e-07 $l=6.0597e-07 $layer=licon1_NDIFF $count=1 $X=5.43
+ $Y=0.37 $X2=5.57 $Y2=0.91
r106 6 45 182 $w=1.7e-07 $l=5.85833e-07 $layer=licon1_NDIFF $count=1 $X=4.57
+ $Y=0.37 $X2=4.71 $Y2=0.89
r107 5 53 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=3.71
+ $Y=0.37 $X2=3.85 $Y2=0.95
r108 4 48 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=2.85
+ $Y=0.37 $X2=2.99 $Y2=0.95
r109 3 37 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.86
+ $Y=0.42 $X2=2 $Y2=0.565
r110 2 30 182 $w=1.7e-07 $l=3.01993e-07 $layer=licon1_NDIFF $count=1 $X=1
+ $Y=0.42 $X2=1.14 $Y2=0.66
r111 1 24 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.42 $X2=0.28 $Y2=0.565
.ends

.subckt PM_SKY130_FD_SC_LS__O221AI_4%A_483_74# 1 2 3 4 5 6 7 8 9 28 32 38 42 44
+ 48 50 54 56 60 67 75 76 77
c110 32 0 1.43357e-20 $X=5.905 $Y=0.475
c111 28 0 1.93079e-19 $X=3.335 $Y=0.475
r112 77 79 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=8.9 $Y=0.835 $X2=8.9
+ $Y2=0.925
r113 71 73 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=6.07 $Y=0.835
+ $X2=6.07 $Y2=0.925
r114 70 71 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=6.07 $Y=0.515
+ $X2=6.07 $Y2=0.835
r115 67 70 1.3969 $w=3.28e-07 $l=4e-08 $layer=LI1_cond $X=6.07 $Y=0.475 $X2=6.07
+ $Y2=0.515
r116 58 60 18.6696 $w=2.48e-07 $l=4.05e-07 $layer=LI1_cond $X=9.84 $Y=0.92
+ $X2=9.84 $Y2=0.515
r117 57 79 2.99516 $w=1.7e-07 $l=1.60078e-07 $layer=LI1_cond $X=9.025 $Y=1.005
+ $X2=8.9 $Y2=0.925
r118 56 58 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=9.715 $Y=1.005
+ $X2=9.84 $Y2=0.92
r119 56 57 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=9.715 $Y=1.005
+ $X2=9.025 $Y2=1.005
r120 52 77 3.91831 $w=2.48e-07 $l=8.5e-08 $layer=LI1_cond $X=8.9 $Y=0.75 $X2=8.9
+ $Y2=0.835
r121 52 54 10.833 $w=2.48e-07 $l=2.35e-07 $layer=LI1_cond $X=8.9 $Y=0.75 $X2=8.9
+ $Y2=0.515
r122 51 76 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.085 $Y=0.835
+ $X2=7.96 $Y2=0.835
r123 50 77 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.775 $Y=0.835
+ $X2=8.9 $Y2=0.835
r124 50 51 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=8.775 $Y=0.835
+ $X2=8.085 $Y2=0.835
r125 46 76 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.96 $Y=0.75
+ $X2=7.96 $Y2=0.835
r126 46 48 5.30124 $w=2.48e-07 $l=1.15e-07 $layer=LI1_cond $X=7.96 $Y=0.75
+ $X2=7.96 $Y2=0.635
r127 45 75 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.155 $Y=0.835
+ $X2=7.03 $Y2=0.835
r128 44 76 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.835 $Y=0.835
+ $X2=7.96 $Y2=0.835
r129 44 45 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=7.835 $Y=0.835
+ $X2=7.155 $Y2=0.835
r130 40 75 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.03 $Y=0.75
+ $X2=7.03 $Y2=0.835
r131 40 42 5.30124 $w=2.48e-07 $l=1.15e-07 $layer=LI1_cond $X=7.03 $Y=0.75
+ $X2=7.03 $Y2=0.635
r132 39 71 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.235 $Y=0.835
+ $X2=6.07 $Y2=0.835
r133 38 75 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.905 $Y=0.835
+ $X2=7.03 $Y2=0.835
r134 38 39 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.905 $Y=0.835
+ $X2=6.235 $Y2=0.835
r135 35 37 39.644 $w=2.48e-07 $l=8.6e-07 $layer=LI1_cond $X=4.28 $Y=0.475
+ $X2=5.14 $Y2=0.475
r136 32 67 2.36532 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=5.905 $Y=0.475
+ $X2=6.07 $Y2=0.475
r137 32 37 35.2648 $w=2.48e-07 $l=7.65e-07 $layer=LI1_cond $X=5.905 $Y=0.475
+ $X2=5.14 $Y2=0.475
r138 28 65 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=3.42 $Y=0.475
+ $X2=3.42 $Y2=0.595
r139 28 35 35.7257 $w=2.48e-07 $l=7.75e-07 $layer=LI1_cond $X=3.505 $Y=0.475
+ $X2=4.28 $Y2=0.475
r140 28 30 35.7257 $w=2.48e-07 $l=7.75e-07 $layer=LI1_cond $X=3.335 $Y=0.475
+ $X2=2.56 $Y2=0.475
r141 9 60 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.66
+ $Y=0.37 $X2=9.8 $Y2=0.515
r142 8 79 182 $w=1.7e-07 $l=6.51594e-07 $layer=licon1_NDIFF $count=1 $X=8.73
+ $Y=0.37 $X2=8.94 $Y2=0.925
r143 8 54 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=8.73
+ $Y=0.37 $X2=8.94 $Y2=0.515
r144 7 48 182 $w=1.7e-07 $l=3.27605e-07 $layer=licon1_NDIFF $count=1 $X=7.86
+ $Y=0.37 $X2=8 $Y2=0.635
r145 6 42 182 $w=1.7e-07 $l=3.27605e-07 $layer=licon1_NDIFF $count=1 $X=6.93
+ $Y=0.37 $X2=7.07 $Y2=0.635
r146 5 73 182 $w=1.7e-07 $l=6.51594e-07 $layer=licon1_NDIFF $count=1 $X=5.86
+ $Y=0.37 $X2=6.07 $Y2=0.925
r147 5 70 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=5.86
+ $Y=0.37 $X2=6.07 $Y2=0.515
r148 4 37 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=5
+ $Y=0.37 $X2=5.14 $Y2=0.515
r149 3 35 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=4.14
+ $Y=0.37 $X2=4.28 $Y2=0.515
r150 2 65 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=3.28
+ $Y=0.37 $X2=3.42 $Y2=0.595
r151 1 30 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=2.415
+ $Y=0.37 $X2=2.56 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__O221AI_4%VGND 1 2 3 4 15 19 23 27 29 31 36 41 46 53
+ 54 57 60 63 66
r114 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r115 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r116 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r117 57 58 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r118 54 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0 $X2=9.36
+ $Y2=0
r119 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r120 51 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.535 $Y=0 $X2=9.37
+ $Y2=0
r121 51 53 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=9.535 $Y=0
+ $X2=9.84 $Y2=0
r122 50 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=9.36
+ $Y2=0
r123 50 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=8.4
+ $Y2=0
r124 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r125 47 63 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=8.605 $Y=0 $X2=8.435
+ $Y2=0
r126 47 49 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=8.605 $Y=0
+ $X2=8.88 $Y2=0
r127 46 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.205 $Y=0 $X2=9.37
+ $Y2=0
r128 46 49 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=9.205 $Y=0
+ $X2=8.88 $Y2=0
r129 45 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.4
+ $Y2=0
r130 45 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=7.44
+ $Y2=0
r131 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r132 42 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.665 $Y=0 $X2=7.5
+ $Y2=0
r133 42 44 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=7.665 $Y=0
+ $X2=7.92 $Y2=0
r134 41 63 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=8.265 $Y=0 $X2=8.435
+ $Y2=0
r135 41 44 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=8.265 $Y=0 $X2=7.92
+ $Y2=0
r136 40 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r137 40 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=6.48
+ $Y2=0
r138 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r139 37 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.735 $Y=0 $X2=6.57
+ $Y2=0
r140 37 39 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=6.735 $Y=0
+ $X2=6.96 $Y2=0
r141 36 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.335 $Y=0 $X2=7.5
+ $Y2=0
r142 36 39 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=7.335 $Y=0
+ $X2=6.96 $Y2=0
r143 33 34 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r144 31 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.405 $Y=0 $X2=6.57
+ $Y2=0
r145 31 33 402.209 $w=1.68e-07 $l=6.165e-06 $layer=LI1_cond $X=6.405 $Y=0
+ $X2=0.24 $Y2=0
r146 29 58 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=6.48 $Y2=0
r147 29 34 1.33793 $w=4.9e-07 $l=4.8e-06 $layer=MET1_cond $X=5.04 $Y=0 $X2=0.24
+ $Y2=0
r148 25 66 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.37 $Y=0.085
+ $X2=9.37 $Y2=0
r149 25 27 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=9.37 $Y=0.085
+ $X2=9.37 $Y2=0.55
r150 21 63 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=8.435 $Y=0.085
+ $X2=8.435 $Y2=0
r151 21 23 13.8971 $w=3.38e-07 $l=4.1e-07 $layer=LI1_cond $X=8.435 $Y=0.085
+ $X2=8.435 $Y2=0.495
r152 17 60 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.5 $Y=0.085 $X2=7.5
+ $Y2=0
r153 17 19 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=7.5 $Y=0.085
+ $X2=7.5 $Y2=0.495
r154 13 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.57 $Y=0.085
+ $X2=6.57 $Y2=0
r155 13 15 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=6.57 $Y=0.085
+ $X2=6.57 $Y2=0.495
r156 4 27 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=9.23 $Y=0.37
+ $X2=9.37 $Y2=0.55
r157 3 23 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=8.29
+ $Y=0.37 $X2=8.435 $Y2=0.495
r158 2 19 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=7.36
+ $Y=0.37 $X2=7.5 $Y2=0.495
r159 1 15 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=6.36
+ $Y=0.37 $X2=6.57 $Y2=0.495
.ends

