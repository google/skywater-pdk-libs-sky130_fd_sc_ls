* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__einvp_2 A TE VGND VNB VPB VPWR Z
X0 a_263_323# TE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_263_323# TE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X2 a_27_368# a_263_323# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X3 a_27_368# A Z VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X4 Z A a_36_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X5 a_36_74# TE VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X6 VGND TE a_36_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X7 VPWR a_263_323# a_27_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X8 Z A a_27_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X9 a_36_74# A Z VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
.ends
