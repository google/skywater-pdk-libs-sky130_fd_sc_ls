# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ls__or3b_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ls__or3b_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.760000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.411000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.800000 1.150000 3.545000 1.320000 ;
        RECT 0.800000 1.320000 1.130000 1.760000 ;
        RECT 3.005000 1.320000 3.545000 1.380000 ;
        RECT 3.285000 1.380000 3.545000 1.550000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.411000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.340000 1.490000 1.670000 1.550000 ;
        RECT 1.340000 1.550000 3.075000 1.800000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 0.255000 0.775000 0.640000 ;
    END
  END C_N
  PIN X
    ANTENNADIFFAREA  1.104900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.055000 0.350000 4.225000 0.960000 ;
        RECT 4.055000 0.960000 5.635000 1.130000 ;
        RECT 4.055000 1.800000 5.635000 1.970000 ;
        RECT 4.055000 1.970000 4.225000 2.980000 ;
        RECT 4.875000 1.970000 5.205000 2.980000 ;
        RECT 4.885000 0.350000 5.135000 0.960000 ;
        RECT 5.405000 1.130000 5.635000 1.800000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 5.760000 0.085000 ;
        RECT 0.945000  0.085000 1.410000 0.640000 ;
        RECT 2.580000  0.085000 2.910000 0.640000 ;
        RECT 3.510000  0.085000 3.850000 0.600000 ;
        RECT 4.405000  0.085000 4.655000 0.790000 ;
        RECT 5.315000  0.085000 5.645000 0.790000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.760000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 5.760000 3.415000 ;
        RECT 0.560000 1.940000 0.890000 3.245000 ;
        RECT 3.505000 2.310000 3.835000 3.245000 ;
        RECT 4.425000 2.140000 4.675000 3.245000 ;
        RECT 5.405000 2.140000 5.655000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 5.760000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.110000 0.810000 1.910000 0.980000 ;
      RECT 0.110000 0.980000 0.465000 1.340000 ;
      RECT 0.110000 1.340000 0.360000 2.980000 ;
      RECT 1.070000 1.970000 1.400000 2.360000 ;
      RECT 1.070000 2.360000 3.335000 2.530000 ;
      RECT 1.070000 2.530000 1.400000 2.980000 ;
      RECT 1.580000 0.310000 1.910000 0.810000 ;
      RECT 1.580000 2.700000 2.835000 2.980000 ;
      RECT 2.030000 1.970000 3.885000 2.140000 ;
      RECT 2.030000 2.140000 2.385000 2.190000 ;
      RECT 2.080000 0.350000 2.410000 0.810000 ;
      RECT 2.080000 0.810000 3.885000 0.980000 ;
      RECT 3.005000 2.310000 3.335000 2.360000 ;
      RECT 3.005000 2.530000 3.335000 2.980000 ;
      RECT 3.090000 0.350000 3.340000 0.810000 ;
      RECT 3.715000 0.980000 3.885000 1.300000 ;
      RECT 3.715000 1.300000 5.175000 1.630000 ;
      RECT 3.715000 1.630000 3.885000 1.970000 ;
  END
END sky130_fd_sc_ls__or3b_4
