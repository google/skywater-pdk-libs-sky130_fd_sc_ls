* File: sky130_fd_sc_ls__a222o_1.spice
* Created: Wed Sep  2 10:49:46 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__a222o_1.pex.spice"
.subckt sky130_fd_sc_ls__a222o_1  VNB VPB C1 C2 B2 B1 A1 A2 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A2	A2
* A1	A1
* B1	B1
* B2	B2
* C2	C2
* C1	C1
* VPB	VPB
* VNB	VNB
MM1006 A_119_74# N_C1_M1006_g N_A_32_74#_M1006_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0768 AS=0.1824 PD=0.88 PS=1.85 NRD=12.18 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75004 A=0.096 P=1.58 MULT=1
MM1013 N_VGND_M1013_d N_C2_M1013_g A_119_74# VNB NSHORT L=0.15 W=0.64 AD=0.2544
+ AS=0.0768 PD=1.435 PS=0.88 NRD=0 NRS=12.18 M=1 R=4.26667 SA=75000.6 SB=75003.6
+ A=0.096 P=1.58 MULT=1
MM1007 A_386_74# N_B2_M1007_g N_VGND_M1013_d VNB NSHORT L=0.15 W=0.64 AD=0.0768
+ AS=0.2544 PD=0.88 PS=1.435 NRD=12.18 NRS=0 M=1 R=4.26667 SA=75001.5 SB=75002.7
+ A=0.096 P=1.58 MULT=1
MM1008 N_A_32_74#_M1008_d N_B1_M1008_g A_386_74# VNB NSHORT L=0.15 W=0.64
+ AD=0.2512 AS=0.0768 PD=1.425 PS=0.88 NRD=0 NRS=12.18 M=1 R=4.26667 SA=75001.9
+ SB=75002.3 A=0.096 P=1.58 MULT=1
MM1004 A_651_74# N_A1_M1004_g N_A_32_74#_M1008_d VNB NSHORT L=0.15 W=0.64
+ AD=0.0768 AS=0.2512 PD=0.88 PS=1.425 NRD=12.18 NRS=0 M=1 R=4.26667 SA=75002.9
+ SB=75001.3 A=0.096 P=1.58 MULT=1
MM1001 N_VGND_M1001_d N_A2_M1001_g A_651_74# VNB NSHORT L=0.15 W=0.64
+ AD=0.185229 AS=0.0768 PD=1.22899 PS=0.88 NRD=21.552 NRS=12.18 M=1 R=4.26667
+ SA=75003.3 SB=75000.9 A=0.096 P=1.58 MULT=1
MM1000 N_X_M1000_d N_A_32_74#_M1000_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.214171 PD=2.05 PS=1.42101 NRD=0 NRS=30.804 M=1 R=4.93333
+ SA=75003.5 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1009 N_A_32_74#_M1009_d N_C1_M1009_g N_A_27_390#_M1009_s VPB PHIGHVT L=0.15
+ W=1 AD=0.2275 AS=0.295 PD=1.455 PS=2.59 NRD=32.4853 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75001.9 A=0.15 P=2.3 MULT=1
MM1011 N_A_27_390#_M1011_d N_C2_M1011_g N_A_32_74#_M1009_d VPB PHIGHVT L=0.15
+ W=1 AD=0.175 AS=0.2275 PD=1.35 PS=1.455 NRD=11.8003 NRS=1.9503 M=1 R=6.66667
+ SA=75000.8 SB=75001.3 A=0.15 P=2.3 MULT=1
MM1012 N_A_337_390#_M1012_d N_B2_M1012_g N_A_27_390#_M1011_d VPB PHIGHVT L=0.15
+ W=1 AD=0.22 AS=0.175 PD=1.44 PS=1.35 NRD=11.8003 NRS=1.9503 M=1 R=6.66667
+ SA=75001.3 SB=75000.8 A=0.15 P=2.3 MULT=1
MM1002 N_A_27_390#_M1002_d N_B1_M1002_g N_A_337_390#_M1012_d VPB PHIGHVT L=0.15
+ W=1 AD=0.295 AS=0.22 PD=2.59 PS=1.44 NRD=1.9503 NRS=19.7 M=1 R=6.66667
+ SA=75001.9 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1003 N_A_337_390#_M1003_d N_A1_M1003_g N_VPWR_M1003_s VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.345 PD=1.3 PS=2.69 NRD=1.9503 NRS=11.8003 M=1 R=6.66667
+ SA=75000.3 SB=75001.3 A=0.15 P=2.3 MULT=1
MM1010 N_VPWR_M1010_d N_A2_M1010_g N_A_337_390#_M1003_d VPB PHIGHVT L=0.15 W=1
+ AD=0.221887 AS=0.15 PD=1.46698 PS=1.3 NRD=18.715 NRS=1.9503 M=1 R=6.66667
+ SA=75000.7 SB=75000.8 A=0.15 P=2.3 MULT=1
MM1005 N_X_M1005_d N_A_32_74#_M1005_g N_VPWR_M1010_d VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.248513 PD=2.83 PS=1.64302 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75001.2 SB=75000.2 A=0.168 P=2.54 MULT=1
DX14_noxref VNB VPB NWDIODE A=9.6348 P=14.08
*
.include "sky130_fd_sc_ls__a222o_1.pxi.spice"
*
.ends
*
*
