* File: sky130_fd_sc_ls__dfrtn_1.pex.spice
* Created: Fri Aug 28 13:14:06 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__DFRTN_1%D 2 3 4 5 7 10 14 16 21 22 23 28 29
c38 5 0 4.35267e-20 $X=0.5 $Y=2.465
r39 28 29 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.27
+ $Y=1.125 $X2=0.27 $Y2=1.125
r40 22 23 16.0907 $w=2.63e-07 $l=3.7e-07 $layer=LI1_cond $X=0.237 $Y=1.665
+ $X2=0.237 $Y2=2.035
r41 21 22 16.0907 $w=2.63e-07 $l=3.7e-07 $layer=LI1_cond $X=0.237 $Y=1.295
+ $X2=0.237 $Y2=1.665
r42 21 29 7.39303 $w=2.63e-07 $l=1.7e-07 $layer=LI1_cond $X=0.237 $Y=1.295
+ $X2=0.237 $Y2=1.125
r43 15 28 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.27 $Y=1.465
+ $X2=0.27 $Y2=1.125
r44 15 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.27 $Y=1.465
+ $X2=0.27 $Y2=1.63
r45 14 28 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.27 $Y=1.11
+ $X2=0.27 $Y2=1.125
r46 13 14 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=0.352 $Y=0.96
+ $X2=0.352 $Y2=1.11
r47 10 13 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=0.525 $Y=0.58
+ $X2=0.525 $Y2=0.96
r48 5 7 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.5 $Y=2.465 $X2=0.5
+ $Y2=2.75
r49 4 5 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.5 $Y=2.375 $X2=0.5
+ $Y2=2.465
r50 3 17 71.7872 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=0.5 $Y=1.995 $X2=0.36
+ $Y2=1.995
r51 3 4 118.556 $w=1.8e-07 $l=3.05e-07 $layer=POLY_cond $X=0.5 $Y=2.07 $X2=0.5
+ $Y2=2.375
r52 2 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.36 $Y=1.92 $X2=0.36
+ $Y2=1.995
r53 2 16 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=0.36 $Y=1.92 $X2=0.36
+ $Y2=1.63
.ends

.subckt PM_SKY130_FD_SC_LS__DFRTN_1%CLK_N 3 6 7 10 12 13
r43 10 13 60.3205 $w=3.55e-07 $l=2.5e-07 $layer=POLY_cond $X=1.527 $Y=1.41
+ $X2=1.527 $Y2=1.66
r44 10 12 56.2568 $w=3.55e-07 $l=2.25e-07 $layer=POLY_cond $X=1.527 $Y=1.41
+ $X2=1.527 $Y2=1.185
r45 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.54
+ $Y=1.41 $X2=1.54 $Y2=1.41
r46 7 11 3.56279 $w=4.68e-07 $l=1.4e-07 $layer=LI1_cond $X=1.68 $Y=1.415
+ $X2=1.54 $Y2=1.415
r47 6 13 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.455 $Y=2.235
+ $X2=1.455 $Y2=1.66
r48 3 12 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.425 $Y=0.74
+ $X2=1.425 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LS__DFRTN_1%A_507_347# 1 2 7 9 11 13 14 16 18 19 21 23
+ 24 26 28 31 35 39 42 43 44 46 47 48 50 51 52 54 56 57 59 60 71 75 78
c178 78 0 1.01786e-19 $X=7.42 $Y=1.29
c179 75 0 1.68346e-20 $X=3.92 $Y=1.715
c180 59 0 2.79847e-19 $X=7.255 $Y=1.29
c181 57 0 2.84298e-19 $X=7.08 $Y=1.29
c182 56 0 2.21313e-20 $X=6.535 $Y=1.21
c183 42 0 1.36584e-19 $X=3.62 $Y=1.245
c184 35 0 6.28401e-20 $X=4.01 $Y=2.165
c185 31 0 7.26587e-20 $X=3.795 $Y=1.215
c186 23 0 1.07929e-19 $X=6.9 $Y=1.29
r187 74 75 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=3.795 $Y=1.715
+ $X2=3.92 $Y2=1.715
r188 68 74 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=3.565 $Y=1.715
+ $X2=3.795 $Y2=1.715
r189 67 68 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.565
+ $Y=1.715 $X2=3.565 $Y2=1.715
r190 65 67 11.3354 $w=7.63e-07 $l=7.25e-07 $layer=LI1_cond $X=2.84 $Y=1.627
+ $X2=3.565 $Y2=1.627
r191 60 78 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.255 $Y=1.29
+ $X2=7.42 $Y2=1.29
r192 59 60 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.255
+ $Y=1.29 $X2=7.255 $Y2=1.29
r193 57 71 14.2244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=7.08 $Y=1.29
+ $X2=6.75 $Y2=1.29
r194 57 59 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=7.08 $Y=1.29
+ $X2=7.255 $Y2=1.29
r195 56 71 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=6.535 $Y=1.21
+ $X2=6.75 $Y2=1.21
r196 54 56 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.45 $Y=1.125
+ $X2=6.535 $Y2=1.21
r197 53 54 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=6.45 $Y=0.425
+ $X2=6.45 $Y2=1.125
r198 51 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.365 $Y=0.34
+ $X2=6.45 $Y2=0.425
r199 51 52 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.365 $Y=0.34
+ $X2=5.695 $Y2=0.34
r200 49 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.61 $Y=0.425
+ $X2=5.695 $Y2=0.34
r201 49 50 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=5.61 $Y=0.425
+ $X2=5.61 $Y2=0.79
r202 47 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.525 $Y=0.875
+ $X2=5.61 $Y2=0.79
r203 47 48 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.525 $Y=0.875
+ $X2=4.855 $Y2=0.875
r204 46 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.77 $Y=0.79
+ $X2=4.855 $Y2=0.875
r205 45 46 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=4.77 $Y=0.465
+ $X2=4.77 $Y2=0.79
r206 43 45 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=4.685 $Y=0.36
+ $X2=4.77 $Y2=0.465
r207 43 44 51.7576 $w=2.08e-07 $l=9.8e-07 $layer=LI1_cond $X=4.685 $Y=0.36
+ $X2=3.705 $Y2=0.36
r208 42 67 0.859926 $w=7.63e-07 $l=5.5e-08 $layer=LI1_cond $X=3.62 $Y=1.627
+ $X2=3.565 $Y2=1.627
r209 41 44 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=3.62 $Y=0.465
+ $X2=3.705 $Y2=0.36
r210 41 42 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=3.62 $Y=0.465
+ $X2=3.62 $Y2=1.245
r211 37 65 0.515955 $w=7.63e-07 $l=3.3e-08 $layer=LI1_cond $X=2.807 $Y=1.627
+ $X2=2.84 $Y2=1.627
r212 37 39 11.0895 $w=2.63e-07 $l=2.55e-07 $layer=LI1_cond $X=2.807 $Y=1.245
+ $X2=2.807 $Y2=0.99
r213 33 35 46.1489 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.92 $Y=2.165
+ $X2=4.01 $Y2=2.165
r214 29 31 153.83 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=3.495 $Y=1.215
+ $X2=3.795 $Y2=1.215
r215 26 28 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=7.675 $Y=1.125
+ $X2=7.675 $Y2=0.805
r216 24 26 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.6 $Y=1.2
+ $X2=7.675 $Y2=1.125
r217 24 78 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=7.6 $Y=1.2 $X2=7.42
+ $Y2=1.2
r218 23 60 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=6.9 $Y=1.29
+ $X2=7.255 $Y2=1.29
r219 19 21 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.81 $Y=1.885
+ $X2=6.81 $Y2=2.46
r220 18 19 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.81 $Y=1.795
+ $X2=6.81 $Y2=1.885
r221 17 23 18.0464 $w=4.25e-07 $l=2.05122e-07 $layer=POLY_cond $X=6.81 $Y=1.455
+ $X2=6.9 $Y2=1.29
r222 17 18 132.161 $w=1.8e-07 $l=3.4e-07 $layer=POLY_cond $X=6.81 $Y=1.455
+ $X2=6.81 $Y2=1.795
r223 14 35 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.01 $Y=2.24
+ $X2=4.01 $Y2=2.165
r224 14 16 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.01 $Y=2.24
+ $X2=4.01 $Y2=2.525
r225 13 33 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.92 $Y=2.09
+ $X2=3.92 $Y2=2.165
r226 12 75 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.92 $Y=1.88
+ $X2=3.92 $Y2=1.715
r227 12 13 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=3.92 $Y=1.88
+ $X2=3.92 $Y2=2.09
r228 11 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.795 $Y=1.55
+ $X2=3.795 $Y2=1.715
r229 10 31 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.795 $Y=1.29
+ $X2=3.795 $Y2=1.215
r230 10 11 133.319 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=3.795 $Y=1.29
+ $X2=3.795 $Y2=1.55
r231 7 29 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.495 $Y=1.14
+ $X2=3.495 $Y2=1.215
r232 7 9 94.7933 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=3.495 $Y=1.14
+ $X2=3.495 $Y2=0.845
r233 2 65 600 $w=1.7e-07 $l=3.80624e-07 $layer=licon1_PDIFF $count=1 $X=2.535
+ $Y=1.735 $X2=2.84 $Y2=1.905
r234 1 39 182 $w=1.7e-07 $l=6.9208e-07 $layer=licon1_NDIFF $count=1 $X=2.55
+ $Y=0.395 $X2=2.76 $Y2=0.99
.ends

.subckt PM_SKY130_FD_SC_LS__DFRTN_1%A_841_288# 1 2 8 11 14 16 19 20 22 23 26 32
+ 34 36 37
c92 36 0 2.21313e-20 $X=6.11 $Y=2.135
c93 34 0 2.66816e-19 $X=6.03 $Y=1.215
r94 36 38 0.373936 $w=8.33e-07 $l=5e-09 $layer=LI1_cond $X=6.282 $Y=2.135
+ $X2=6.282 $Y2=2.14
r95 36 37 11.6472 $w=8.33e-07 $l=1.65e-07 $layer=LI1_cond $X=6.282 $Y=2.135
+ $X2=6.282 $Y2=1.97
r96 32 38 11.3712 $w=7.08e-07 $l=6.75e-07 $layer=LI1_cond $X=6.345 $Y=2.815
+ $X2=6.345 $Y2=2.14
r97 28 34 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=5.95 $Y=1.3
+ $X2=6.03 $Y2=1.215
r98 28 37 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.95 $Y=1.3 $X2=5.95
+ $Y2=1.97
r99 24 34 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.03 $Y=1.13 $X2=6.03
+ $Y2=1.215
r100 24 26 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=6.03 $Y=1.13
+ $X2=6.03 $Y2=0.76
r101 22 34 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.865 $Y=1.215
+ $X2=6.03 $Y2=1.215
r102 22 23 78.9412 $w=1.68e-07 $l=1.21e-06 $layer=LI1_cond $X=5.865 $Y=1.215
+ $X2=4.655 $Y2=1.215
r103 20 41 42.0275 $w=4.05e-07 $l=2.7e-07 $layer=POLY_cond $X=4.407 $Y=1.61
+ $X2=4.407 $Y2=1.88
r104 20 40 46.4766 $w=4.05e-07 $l=1.7e-07 $layer=POLY_cond $X=4.407 $Y=1.61
+ $X2=4.407 $Y2=1.44
r105 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.37
+ $Y=1.61 $X2=4.37 $Y2=1.61
r106 17 23 8.19669 $w=1.7e-07 $l=2.28583e-07 $layer=LI1_cond $X=4.465 $Y=1.3
+ $X2=4.655 $Y2=1.215
r107 17 19 9.40151 $w=3.78e-07 $l=3.1e-07 $layer=LI1_cond $X=4.465 $Y=1.3
+ $X2=4.465 $Y2=1.61
r108 14 40 305.096 $w=1.5e-07 $l=5.95e-07 $layer=POLY_cond $X=4.535 $Y=0.845
+ $X2=4.535 $Y2=1.44
r109 11 16 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.4 $Y=2.525 $X2=4.4
+ $Y2=2.24
r110 8 16 43.2804 $w=2.85e-07 $l=1.42e-07 $layer=POLY_cond $X=4.467 $Y=2.098
+ $X2=4.467 $Y2=2.24
r111 8 41 45.8847 $w=2.85e-07 $l=2.18e-07 $layer=POLY_cond $X=4.467 $Y=2.098
+ $X2=4.467 $Y2=1.88
r112 2 36 200 $w=1.7e-07 $l=2.40312e-07 $layer=licon1_PDIFF $count=3 $X=5.955
+ $Y=1.96 $X2=6.11 $Y2=2.135
r113 2 32 200 $w=1.7e-07 $l=9.29274e-07 $layer=licon1_PDIFF $count=3 $X=5.955
+ $Y=1.96 $X2=6.11 $Y2=2.815
r114 1 26 91 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=2 $X=5.89
+ $Y=0.595 $X2=6.03 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_LS__DFRTN_1%RESET_B 3 6 7 10 11 12 15 16 19 23 26 29 30
+ 32 33 34 35 36 37 38 43 44 46 49 50 54 55 56 59
c231 35 0 9.76428e-20 $X=4.895 $Y=1.665
r232 59 62 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.545 $Y=1.63
+ $X2=8.545 $Y2=1.795
r233 59 61 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.545 $Y=1.63
+ $X2=8.545 $Y2=1.465
r234 54 57 33.5009 $w=3.45e-07 $l=1.65e-07 $layer=POLY_cond $X=4.992 $Y=1.635
+ $X2=4.992 $Y2=1.8
r235 54 56 33.5009 $w=3.45e-07 $l=1.65e-07 $layer=POLY_cond $X=4.992 $Y=1.635
+ $X2=4.992 $Y2=1.47
r236 54 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5
+ $Y=1.635 $X2=5 $Y2=1.635
r237 50 66 7.25612 $w=4.03e-07 $l=2.55e-07 $layer=LI1_cond $X=1.082 $Y=1.41
+ $X2=1.082 $Y2=1.665
r238 49 52 55.5535 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=0.975 $Y=1.41
+ $X2=0.975 $Y2=1.66
r239 49 51 56.7032 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=0.975 $Y=1.41
+ $X2=0.975 $Y2=1.185
r240 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.975
+ $Y=1.41 $X2=0.975 $Y2=1.41
r241 46 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=1.665
+ $X2=1.2 $Y2=1.665
r242 44 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.545
+ $Y=1.63 $X2=8.545 $Y2=1.63
r243 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=1.665
+ $X2=8.4 $Y2=1.665
r244 40 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=1.665
+ $X2=5.04 $Y2=1.665
r245 38 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.185 $Y=1.665
+ $X2=5.04 $Y2=1.665
r246 37 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.255 $Y=1.665
+ $X2=8.4 $Y2=1.665
r247 37 38 3.7995 $w=1.4e-07 $l=3.07e-06 $layer=MET1_cond $X=8.255 $Y=1.665
+ $X2=5.185 $Y2=1.665
r248 36 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.345 $Y=1.665
+ $X2=1.2 $Y2=1.665
r249 35 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.895 $Y=1.665
+ $X2=5.04 $Y2=1.665
r250 35 36 4.39356 $w=1.4e-07 $l=3.55e-06 $layer=MET1_cond $X=4.895 $Y=1.665
+ $X2=1.345 $Y2=1.665
r251 30 32 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=8.62 $Y=2.465
+ $X2=8.62 $Y2=2.75
r252 29 30 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=8.62 $Y=2.375
+ $X2=8.62 $Y2=2.465
r253 29 62 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=8.62 $Y=2.375
+ $X2=8.62 $Y2=1.795
r254 26 61 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.605 $Y=0.805
+ $X2=8.605 $Y2=1.465
r255 23 34 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.895 $Y=2.525
+ $X2=4.895 $Y2=2.24
r256 21 23 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=4.895 $Y=3.075
+ $X2=4.895 $Y2=2.525
r257 19 34 39.0221 $w=2.35e-07 $l=1.17e-07 $layer=POLY_cond $X=4.937 $Y=2.123
+ $X2=4.937 $Y2=2.24
r258 19 57 85.3729 $w=2.35e-07 $l=3.23e-07 $layer=POLY_cond $X=4.937 $Y=2.123
+ $X2=4.937 $Y2=1.8
r259 16 33 39.0221 $w=2.35e-07 $l=1.17e-07 $layer=POLY_cond $X=4.937 $Y=1.247
+ $X2=4.937 $Y2=1.13
r260 16 56 58.9417 $w=2.35e-07 $l=2.23e-07 $layer=POLY_cond $X=4.937 $Y=1.247
+ $X2=4.937 $Y2=1.47
r261 15 33 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.895 $Y=0.845
+ $X2=4.895 $Y2=1.13
r262 11 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.82 $Y=3.15
+ $X2=4.895 $Y2=3.075
r263 11 12 1945.95 $w=1.5e-07 $l=3.795e-06 $layer=POLY_cond $X=4.82 $Y=3.15
+ $X2=1.025 $Y2=3.15
r264 8 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.95 $Y=3.075
+ $X2=1.025 $Y2=3.15
r265 8 10 166.649 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=0.95 $Y=3.075
+ $X2=0.95 $Y2=2.75
r266 7 10 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=0.95 $Y=2.24
+ $X2=0.95 $Y2=2.75
r267 6 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.95 $Y=2.15 $X2=0.95
+ $Y2=2.24
r268 6 52 190.468 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=0.95 $Y=2.15
+ $X2=0.95 $Y2=1.66
r269 3 51 310.223 $w=1.5e-07 $l=6.05e-07 $layer=POLY_cond $X=0.915 $Y=0.58
+ $X2=0.915 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LS__DFRTN_1%A_714_127# 1 2 3 12 14 16 18 21 23 24 27 29
+ 31
c101 21 0 1.87783e-19 $X=3.96 $Y=0.855
r102 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.54
+ $Y=1.635 $X2=5.54 $Y2=1.635
r103 29 31 10.7241 $w=3.58e-07 $l=3.35e-07 $layer=LI1_cond $X=5.515 $Y=1.97
+ $X2=5.515 $Y2=1.635
r104 25 29 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=5.135 $Y=2.055
+ $X2=5.515 $Y2=2.055
r105 25 27 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=5.135 $Y=2.14
+ $X2=5.135 $Y2=2.55
r106 24 36 15.6857 $w=3.85e-07 $l=5.98235e-07 $layer=LI1_cond $X=4.075 $Y=2.055
+ $X2=3.847 $Y2=2.55
r107 23 25 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=4.97 $Y=2.055
+ $X2=5.135 $Y2=2.055
r108 23 24 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=4.97 $Y=2.055
+ $X2=4.075 $Y2=2.055
r109 19 24 5.49905 $w=3.85e-07 $l=1.36015e-07 $layer=LI1_cond $X=3.975 $Y=1.97
+ $X2=4.075 $Y2=2.055
r110 19 21 61.8318 $w=1.98e-07 $l=1.115e-06 $layer=LI1_cond $X=3.975 $Y=1.97
+ $X2=3.975 $Y2=0.855
r111 18 32 34.9723 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=5.74 $Y=1.635
+ $X2=5.54 $Y2=1.635
r112 14 18 59.8433 $w=2.19e-07 $l=2.62202e-07 $layer=POLY_cond $X=5.88 $Y=1.885
+ $X2=5.855 $Y2=1.635
r113 14 16 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.88 $Y=1.885
+ $X2=5.88 $Y2=2.46
r114 10 18 41.1355 $w=2.19e-07 $l=1.83916e-07 $layer=POLY_cond $X=5.815 $Y=1.47
+ $X2=5.855 $Y2=1.635
r115 10 12 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=5.815 $Y=1.47
+ $X2=5.815 $Y2=0.965
r116 3 27 600 $w=1.7e-07 $l=3.06594e-07 $layer=licon1_PDIFF $count=1 $X=4.97
+ $Y=2.315 $X2=5.135 $Y2=2.55
r117 2 36 600 $w=1.7e-07 $l=3.00791e-07 $layer=licon1_PDIFF $count=1 $X=3.635
+ $Y=2.315 $X2=3.785 $Y2=2.55
r118 1 21 182 $w=1.7e-07 $l=4.8775e-07 $layer=licon1_NDIFF $count=1 $X=3.57
+ $Y=0.635 $X2=3.96 $Y2=0.855
.ends

.subckt PM_SKY130_FD_SC_LS__DFRTN_1%A_300_74# 1 2 7 9 13 14 15 16 19 20 21 22 24
+ 27 29 34 35 37 38 39 40 41 42 49 51 55 56 59 62 63
c195 56 0 1.21652e-19 $X=7.475 $Y=1.86
c196 16 0 3.24367e-19 $X=3.04 $Y=1.435
r197 63 72 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.345 $Y=1.635
+ $X2=6.345 $Y2=1.47
r198 62 65 3.0228 $w=3.03e-07 $l=8e-08 $layer=LI1_cond $X=6.357 $Y=1.635
+ $X2=6.357 $Y2=1.715
r199 62 63 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.345
+ $Y=1.635 $X2=6.345 $Y2=1.635
r200 59 60 10.1051 $w=4.95e-07 $l=4.1e-07 $layer=LI1_cond $X=1.64 $Y=0.68
+ $X2=2.05 $Y2=0.68
r201 55 56 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.475
+ $Y=1.86 $X2=7.475 $Y2=1.86
r202 53 55 2.76586 $w=2.48e-07 $l=6e-08 $layer=LI1_cond $X=7.435 $Y=1.8
+ $X2=7.435 $Y2=1.86
r203 52 65 4.15824 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=6.51 $Y=1.715
+ $X2=6.357 $Y2=1.715
r204 51 53 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=7.31 $Y=1.715
+ $X2=7.435 $Y2=1.8
r205 51 52 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=7.31 $Y=1.715
+ $X2=6.51 $Y2=1.715
r206 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.08
+ $Y=1.41 $X2=2.08 $Y2=1.41
r207 47 49 20.5435 $w=2.28e-07 $l=4.1e-07 $layer=LI1_cond $X=2.05 $Y=1.82
+ $X2=2.05 $Y2=1.41
r208 46 60 5.23959 $w=2.3e-07 $l=3.3e-07 $layer=LI1_cond $X=2.05 $Y=1.01
+ $X2=2.05 $Y2=0.68
r209 46 49 20.0425 $w=2.28e-07 $l=4e-07 $layer=LI1_cond $X=2.05 $Y=1.01 $X2=2.05
+ $Y2=1.41
r210 42 47 6.89722 $w=1.9e-07 $l=1.55403e-07 $layer=LI1_cond $X=1.935 $Y=1.915
+ $X2=2.05 $Y2=1.82
r211 42 44 14.8852 $w=1.88e-07 $l=2.55e-07 $layer=LI1_cond $X=1.935 $Y=1.915
+ $X2=1.68 $Y2=1.915
r212 41 56 40.6942 $w=4.1e-07 $l=3e-07 $layer=POLY_cond $X=7.515 $Y=2.16
+ $X2=7.515 $Y2=1.86
r213 38 50 37.6949 $w=4.5e-07 $l=3.05e-07 $layer=POLY_cond $X=2.385 $Y=1.435
+ $X2=2.08 $Y2=1.435
r214 38 39 1.87879 $w=4.5e-07 $l=8.2e-08 $layer=POLY_cond $X=2.385 $Y=1.435
+ $X2=2.467 $Y2=1.435
r215 35 41 44.6839 $w=3.29e-07 $l=3.70473e-07 $layer=POLY_cond $X=7.66 $Y=2.465
+ $X2=7.515 $Y2=2.16
r216 35 37 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.66 $Y=2.465
+ $X2=7.66 $Y2=2.75
r217 34 72 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=6.255 $Y=0.965
+ $X2=6.255 $Y2=1.47
r218 31 34 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=6.255 $Y=0.255
+ $X2=6.255 $Y2=0.965
r219 30 40 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.25 $Y=0.18
+ $X2=4.175 $Y2=0.18
r220 29 31 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.18 $Y=0.18
+ $X2=6.255 $Y2=0.255
r221 29 30 989.638 $w=1.5e-07 $l=1.93e-06 $layer=POLY_cond $X=6.18 $Y=0.18
+ $X2=4.25 $Y2=0.18
r222 25 40 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.175 $Y=0.255
+ $X2=4.175 $Y2=0.18
r223 25 27 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=4.175 $Y=0.255
+ $X2=4.175 $Y2=0.845
r224 22 24 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.56 $Y=2.24
+ $X2=3.56 $Y2=2.525
r225 20 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.485 $Y=2.165
+ $X2=3.56 $Y2=2.24
r226 20 21 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=3.485 $Y=2.165
+ $X2=3.19 $Y2=2.165
r227 19 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.115 $Y=2.09
+ $X2=3.19 $Y2=2.165
r228 18 19 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.115 $Y=1.66
+ $X2=3.115 $Y2=2.09
r229 17 39 1.87879 $w=4.5e-07 $l=8.3e-08 $layer=POLY_cond $X=2.55 $Y=1.435
+ $X2=2.467 $Y2=1.435
r230 16 18 36.8 $w=4.5e-07 $l=2.59808e-07 $layer=POLY_cond $X=3.04 $Y=1.435
+ $X2=3.115 $Y2=1.66
r231 16 17 60.559 $w=4.5e-07 $l=4.9e-07 $layer=POLY_cond $X=3.04 $Y=1.435
+ $X2=2.55 $Y2=1.435
r232 14 40 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.1 $Y=0.18
+ $X2=4.175 $Y2=0.18
r233 14 15 794.787 $w=1.5e-07 $l=1.55e-06 $layer=POLY_cond $X=4.1 $Y=0.18
+ $X2=2.55 $Y2=0.18
r234 11 39 27.1559 $w=1.5e-07 $l=2.28965e-07 $layer=POLY_cond $X=2.475 $Y=1.21
+ $X2=2.467 $Y2=1.435
r235 11 13 228.181 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.475 $Y=1.21
+ $X2=2.475 $Y2=0.765
r236 10 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.475 $Y=0.255
+ $X2=2.55 $Y2=0.18
r237 10 13 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=2.475 $Y=0.255
+ $X2=2.475 $Y2=0.765
r238 7 39 27.1559 $w=1.5e-07 $l=2.28473e-07 $layer=POLY_cond $X=2.46 $Y=1.66
+ $X2=2.467 $Y2=1.435
r239 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.46 $Y=1.66
+ $X2=2.46 $Y2=2.235
r240 2 44 600 $w=1.7e-07 $l=2.33238e-07 $layer=licon1_PDIFF $count=1 $X=1.53
+ $Y=1.735 $X2=1.68 $Y2=1.905
r241 1 59 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.5
+ $Y=0.37 $X2=1.64 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__DFRTN_1%A_1598_93# 1 2 9 11 13 14 21 23 26 27 31
c89 9 0 1.58195e-19 $X=8.065 $Y=0.805
r90 29 31 8.03677 $w=3.78e-07 $l=2.65e-07 $layer=LI1_cond $X=9.21 $Y=0.765
+ $X2=9.475 $Y2=0.765
r91 25 31 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=9.475 $Y=0.955
+ $X2=9.475 $Y2=0.765
r92 25 26 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=9.475 $Y=0.955
+ $X2=9.475 $Y2=1.965
r93 24 27 6.08426 $w=2.7e-07 $l=2.29619e-07 $layer=LI1_cond $X=9.05 $Y=2.05
+ $X2=8.865 $Y2=2.15
r94 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.39 $Y=2.05
+ $X2=9.475 $Y2=1.965
r95 23 24 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=9.39 $Y=2.05
+ $X2=9.05 $Y2=2.05
r96 19 27 0.630948 $w=3.3e-07 $l=1.94743e-07 $layer=LI1_cond $X=8.845 $Y=2.335
+ $X2=8.865 $Y2=2.15
r97 19 21 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=8.845 $Y=2.335
+ $X2=8.845 $Y2=2.75
r98 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.155
+ $Y=2.17 $X2=8.155 $Y2=2.17
r99 14 27 6.08426 $w=2.7e-07 $l=1.85e-07 $layer=LI1_cond $X=8.68 $Y=2.15
+ $X2=8.865 $Y2=2.15
r100 14 16 16.3522 $w=3.68e-07 $l=5.25e-07 $layer=LI1_cond $X=8.68 $Y=2.15
+ $X2=8.155 $Y2=2.15
r101 11 17 60.4771 $w=2.87e-07 $l=3.30379e-07 $layer=POLY_cond $X=8.08 $Y=2.465
+ $X2=8.155 $Y2=2.17
r102 11 13 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=8.08 $Y=2.465
+ $X2=8.08 $Y2=2.75
r103 7 17 38.6443 $w=2.87e-07 $l=2.05122e-07 $layer=POLY_cond $X=8.065 $Y=2.005
+ $X2=8.155 $Y2=2.17
r104 7 9 615.319 $w=1.5e-07 $l=1.2e-06 $layer=POLY_cond $X=8.065 $Y=2.005
+ $X2=8.065 $Y2=0.805
r105 2 21 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=8.695
+ $Y=2.54 $X2=8.845 $Y2=2.75
r106 1 29 182 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_NDIFF $count=1 $X=9.07
+ $Y=0.595 $X2=9.21 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LS__DFRTN_1%A_1266_119# 1 2 7 9 10 11 12 14 15 17 19 21
+ 22 24 26 29 33 38 40 41 46 48 50 51
c138 48 0 2.64234e-19 $X=7.815 $Y=1.21
r139 50 51 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.085
+ $Y=1.29 $X2=9.085 $Y2=1.29
r140 46 47 20.5133 $w=2.26e-07 $l=3.8e-07 $layer=LI1_cond $X=7.435 $Y=2.7
+ $X2=7.815 $Y2=2.7
r141 42 48 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.9 $Y=1.21
+ $X2=7.815 $Y2=1.21
r142 41 50 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=8.92 $Y=1.21
+ $X2=9.07 $Y2=1.21
r143 41 42 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=8.92 $Y=1.21
+ $X2=7.9 $Y2=1.21
r144 40 47 2.4068 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.815 $Y=2.535
+ $X2=7.815 $Y2=2.7
r145 39 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.815 $Y=1.295
+ $X2=7.815 $Y2=1.21
r146 39 40 80.8984 $w=1.68e-07 $l=1.24e-06 $layer=LI1_cond $X=7.815 $Y=1.295
+ $X2=7.815 $Y2=2.535
r147 38 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.815 $Y=1.125
+ $X2=7.815 $Y2=1.21
r148 37 38 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=7.815 $Y=0.955
+ $X2=7.815 $Y2=1.125
r149 33 46 1.22073 $w=3.3e-07 $l=1.75152e-07 $layer=LI1_cond $X=7.435 $Y=2.7
+ $X2=7.435 $Y2=2.7
r150 33 35 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=7.435 $Y=2.7 $X2=7.035
+ $Y2=2.7
r151 29 37 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.73 $Y=0.79
+ $X2=7.815 $Y2=0.955
r152 29 31 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=7.73 $Y=0.79
+ $X2=7.46 $Y2=0.79
r153 27 51 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=9.085 $Y=1.63
+ $X2=9.085 $Y2=1.29
r154 27 28 50.3824 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=9.085 $Y=1.63
+ $X2=9.085 $Y2=1.97
r155 25 51 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=9.085 $Y=1.275
+ $X2=9.085 $Y2=1.29
r156 25 26 13.5877 $w=2.4e-07 $l=7.5e-08 $layer=POLY_cond $X=9.085 $Y=1.275
+ $X2=9.085 $Y2=1.2
r157 22 24 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=10.04 $Y=2.045
+ $X2=10.04 $Y2=2.54
r158 19 21 122.107 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=10.03 $Y=1.125
+ $X2=10.03 $Y2=0.745
r159 18 28 18.414 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.25 $Y=1.97
+ $X2=9.085 $Y2=1.97
r160 17 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.965 $Y=1.97
+ $X2=10.04 $Y2=2.045
r161 17 18 366.628 $w=1.5e-07 $l=7.15e-07 $layer=POLY_cond $X=9.965 $Y=1.97
+ $X2=9.25 $Y2=1.97
r162 16 26 12.1617 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.25 $Y=1.2
+ $X2=9.085 $Y2=1.2
r163 15 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.955 $Y=1.2
+ $X2=10.03 $Y2=1.125
r164 15 16 361.5 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=9.955 $Y=1.2
+ $X2=9.25 $Y2=1.2
r165 12 14 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=9.07 $Y=2.465
+ $X2=9.07 $Y2=2.75
r166 11 12 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=9.07 $Y=2.375
+ $X2=9.07 $Y2=2.465
r167 10 28 19.4594 $w=2.93e-07 $l=8.21584e-08 $layer=POLY_cond $X=9.07 $Y=2.045
+ $X2=9.085 $Y2=1.97
r168 10 11 128.274 $w=1.8e-07 $l=3.3e-07 $layer=POLY_cond $X=9.07 $Y=2.045
+ $X2=9.07 $Y2=2.375
r169 7 26 13.5877 $w=2.4e-07 $l=1.21861e-07 $layer=POLY_cond $X=8.995 $Y=1.125
+ $X2=9.085 $Y2=1.2
r170 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=8.995 $Y=1.125
+ $X2=8.995 $Y2=0.805
r171 2 46 600 $w=1.7e-07 $l=9.77036e-07 $layer=licon1_PDIFF $count=1 $X=6.885
+ $Y=1.96 $X2=7.435 $Y2=2.7
r172 2 35 600 $w=1.7e-07 $l=8.11542e-07 $layer=licon1_PDIFF $count=1 $X=6.885
+ $Y=1.96 $X2=7.035 $Y2=2.7
r173 1 31 91 $w=1.7e-07 $l=1.22362e-06 $layer=licon1_NDIFF $count=2 $X=6.33
+ $Y=0.595 $X2=7.46 $Y2=0.79
.ends

.subckt PM_SKY130_FD_SC_LS__DFRTN_1%A_1934_94# 1 2 7 9 10 12 13 15 19 24 27 31
r60 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.48
+ $Y=1.485 $X2=10.48 $Y2=1.485
r61 25 31 0.364692 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=9.98 $Y=1.485
+ $X2=9.855 $Y2=1.485
r62 25 27 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=9.98 $Y=1.485
+ $X2=10.48 $Y2=1.485
r63 24 30 1.61342 $w=2.48e-07 $l=3.5e-08 $layer=LI1_cond $X=9.855 $Y=2.27
+ $X2=9.855 $Y2=2.305
r64 21 31 6.46576 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=9.855 $Y=1.65
+ $X2=9.855 $Y2=1.485
r65 21 24 28.5806 $w=2.48e-07 $l=6.2e-07 $layer=LI1_cond $X=9.855 $Y=1.65
+ $X2=9.855 $Y2=2.27
r66 17 31 6.46576 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=9.855 $Y=1.32
+ $X2=9.855 $Y2=1.485
r67 17 19 26.5062 $w=2.48e-07 $l=5.75e-07 $layer=LI1_cond $X=9.855 $Y=1.32
+ $X2=9.855 $Y2=0.745
r68 13 30 6.46688 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=9.815 $Y=2.47
+ $X2=9.815 $Y2=2.305
r69 13 15 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=9.815 $Y=2.47
+ $X2=9.815 $Y2=2.815
r70 10 28 57.6553 $w=2.91e-07 $l=3.10805e-07 $layer=POLY_cond $X=10.545 $Y=1.765
+ $X2=10.48 $Y2=1.485
r71 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=10.545 $Y=1.765
+ $X2=10.545 $Y2=2.4
r72 7 28 38.6072 $w=2.91e-07 $l=1.92678e-07 $layer=POLY_cond $X=10.54 $Y=1.32
+ $X2=10.48 $Y2=1.485
r73 7 9 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=10.54 $Y=1.32 $X2=10.54
+ $Y2=0.84
r74 2 24 600 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_PDIFF $count=1 $X=9.69
+ $Y=2.12 $X2=9.815 $Y2=2.27
r75 2 15 600 $w=1.7e-07 $l=7.54917e-07 $layer=licon1_PDIFF $count=1 $X=9.69
+ $Y=2.12 $X2=9.815 $Y2=2.815
r76 1 19 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=9.67
+ $Y=0.47 $X2=9.815 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_LS__DFRTN_1%VPWR 1 2 3 4 5 6 7 8 25 27 31 35 39 41 45 49
+ 53 57 60 61 63 64 65 67 72 77 92 101 102 108 111 114 117 120
c132 31 0 4.35267e-20 $X=1.18 $Y=2.685
r133 120 121 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r134 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r135 111 112 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r136 108 109 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r137 105 106 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r138 101 102 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r139 99 102 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=10.8 $Y2=3.33
r140 99 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=9.36 $Y2=3.33
r141 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r142 96 120 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.46 $Y=3.33
+ $X2=9.335 $Y2=3.33
r143 96 98 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=9.46 $Y=3.33
+ $X2=9.84 $Y2=3.33
r144 95 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=9.36 $Y2=3.33
r145 94 95 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r146 92 120 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.21 $Y=3.33
+ $X2=9.335 $Y2=3.33
r147 92 94 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=9.21 $Y=3.33
+ $X2=8.88 $Y2=3.33
r148 91 95 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.88 $Y2=3.33
r149 90 91 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r150 88 91 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=7.92 $Y2=3.33
r151 87 90 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=6 $Y=3.33 $X2=7.92
+ $Y2=3.33
r152 87 88 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r153 85 117 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.82 $Y=3.33
+ $X2=5.655 $Y2=3.33
r154 85 87 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=5.82 $Y=3.33 $X2=6
+ $Y2=3.33
r155 84 115 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r156 83 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r157 81 84 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=4.08 $Y2=3.33
r158 81 112 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r159 80 83 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.64 $Y=3.33
+ $X2=4.08 $Y2=3.33
r160 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r161 78 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.4 $Y=3.33
+ $X2=2.235 $Y2=3.33
r162 78 80 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=2.4 $Y=3.33
+ $X2=2.64 $Y2=3.33
r163 77 114 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.46 $Y=3.33
+ $X2=4.625 $Y2=3.33
r164 77 83 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=4.46 $Y=3.33
+ $X2=4.08 $Y2=3.33
r165 76 112 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r166 76 109 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r167 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r168 73 108 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.37 $Y=3.33
+ $X2=1.205 $Y2=3.33
r169 73 75 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1.37 $Y=3.33
+ $X2=1.68 $Y2=3.33
r170 72 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.07 $Y=3.33
+ $X2=2.235 $Y2=3.33
r171 72 75 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=2.07 $Y=3.33
+ $X2=1.68 $Y2=3.33
r172 71 109 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r173 71 106 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r174 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r175 68 105 4.746 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=0.44 $Y=3.33 $X2=0.22
+ $Y2=3.33
r176 68 70 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.44 $Y=3.33
+ $X2=0.72 $Y2=3.33
r177 67 108 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.04 $Y=3.33
+ $X2=1.205 $Y2=3.33
r178 67 70 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.04 $Y=3.33
+ $X2=0.72 $Y2=3.33
r179 65 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33 $X2=6
+ $Y2=3.33
r180 65 115 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=4.56 $Y2=3.33
r181 65 117 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r182 63 98 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=10.15 $Y=3.33
+ $X2=9.84 $Y2=3.33
r183 63 64 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.15 $Y=3.33
+ $X2=10.275 $Y2=3.33
r184 62 101 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=10.4 $Y=3.33
+ $X2=10.8 $Y2=3.33
r185 62 64 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.4 $Y=3.33
+ $X2=10.275 $Y2=3.33
r186 60 90 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=8.14 $Y=3.33
+ $X2=7.92 $Y2=3.33
r187 60 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.14 $Y=3.33
+ $X2=8.305 $Y2=3.33
r188 59 94 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=8.47 $Y=3.33
+ $X2=8.88 $Y2=3.33
r189 59 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.47 $Y=3.33
+ $X2=8.305 $Y2=3.33
r190 55 64 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=10.275 $Y=3.245
+ $X2=10.275 $Y2=3.33
r191 55 57 45.1758 $w=2.48e-07 $l=9.8e-07 $layer=LI1_cond $X=10.275 $Y=3.245
+ $X2=10.275 $Y2=2.265
r192 51 120 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.335 $Y=3.245
+ $X2=9.335 $Y2=3.33
r193 51 53 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=9.335 $Y=3.245
+ $X2=9.335 $Y2=2.75
r194 47 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.305 $Y=3.245
+ $X2=8.305 $Y2=3.33
r195 47 49 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=8.305 $Y=3.245
+ $X2=8.305 $Y2=2.75
r196 43 117 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.655 $Y=3.245
+ $X2=5.655 $Y2=3.33
r197 43 45 27.938 $w=3.28e-07 $l=8e-07 $layer=LI1_cond $X=5.655 $Y=3.245
+ $X2=5.655 $Y2=2.445
r198 42 114 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.79 $Y=3.33
+ $X2=4.625 $Y2=3.33
r199 41 117 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.49 $Y=3.33
+ $X2=5.655 $Y2=3.33
r200 41 42 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=5.49 $Y=3.33 $X2=4.79
+ $Y2=3.33
r201 37 114 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.625 $Y=3.245
+ $X2=4.625 $Y2=3.33
r202 37 39 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=4.625 $Y=3.245
+ $X2=4.625 $Y2=2.55
r203 33 111 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.235 $Y=3.245
+ $X2=2.235 $Y2=3.33
r204 33 35 22.3504 $w=3.28e-07 $l=6.4e-07 $layer=LI1_cond $X=2.235 $Y=3.245
+ $X2=2.235 $Y2=2.605
r205 29 108 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=3.245
+ $X2=1.205 $Y2=3.33
r206 29 31 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=1.205 $Y=3.245
+ $X2=1.205 $Y2=2.685
r207 25 105 3.02018 $w=3.3e-07 $l=1.09087e-07 $layer=LI1_cond $X=0.275 $Y=3.245
+ $X2=0.22 $Y2=3.33
r208 25 27 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=0.275 $Y=3.245
+ $X2=0.275 $Y2=2.75
r209 8 57 300 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=2 $X=10.115
+ $Y=2.12 $X2=10.315 $Y2=2.265
r210 7 53 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=9.145
+ $Y=2.54 $X2=9.295 $Y2=2.75
r211 6 49 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=8.155
+ $Y=2.54 $X2=8.305 $Y2=2.75
r212 5 45 300 $w=1.7e-07 $l=5.43921e-07 $layer=licon1_PDIFF $count=2 $X=5.53
+ $Y=1.96 $X2=5.655 $Y2=2.445
r213 4 39 600 $w=1.7e-07 $l=3.00791e-07 $layer=licon1_PDIFF $count=1 $X=4.475
+ $Y=2.315 $X2=4.625 $Y2=2.55
r214 3 35 600 $w=1.7e-07 $l=9.39707e-07 $layer=licon1_PDIFF $count=1 $X=2.09
+ $Y=1.735 $X2=2.235 $Y2=2.605
r215 2 31 600 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=1 $X=1.025
+ $Y=2.54 $X2=1.18 $Y2=2.685
r216 1 27 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.54 $X2=0.275 $Y2=2.75
.ends

.subckt PM_SKY130_FD_SC_LS__DFRTN_1%A_33_74# 1 2 3 4 14 17 19 21 22 23 25 29 33
+ 38 40 42
c104 23 0 5.46906e-20 $X=3.17 $Y=2.265
c105 14 0 1.52323e-19 $X=0.625 $Y=2.18
r106 36 38 8.25044 $w=4.38e-07 $l=3.15e-07 $layer=LI1_cond $X=0.31 $Y=0.57
+ $X2=0.625 $Y2=0.57
r107 31 33 9.21954 $w=2.48e-07 $l=2e-07 $layer=LI1_cond $X=3.295 $Y=2.35
+ $X2=3.295 $Y2=2.55
r108 27 29 9.21954 $w=2.48e-07 $l=2e-07 $layer=LI1_cond $X=3.24 $Y=0.655
+ $X2=3.24 $Y2=0.855
r109 26 41 1.47909 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=2.575 $Y=0.57
+ $X2=2.455 $Y2=0.57
r110 25 27 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.115 $Y=0.57
+ $X2=3.24 $Y2=0.655
r111 25 26 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=3.115 $Y=0.57
+ $X2=2.575 $Y2=0.57
r112 24 42 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.505 $Y=2.265
+ $X2=2.42 $Y2=2.265
r113 23 31 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.17 $Y=2.265
+ $X2=3.295 $Y2=2.35
r114 23 24 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=3.17 $Y=2.265
+ $X2=2.505 $Y2=2.265
r115 22 42 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.42 $Y=2.18
+ $X2=2.42 $Y2=2.265
r116 21 41 10.0019 $w=1.93e-07 $l=1.7161e-07 $layer=LI1_cond $X=2.42 $Y=0.725
+ $X2=2.455 $Y2=0.57
r117 21 22 94.9251 $w=1.68e-07 $l=1.455e-06 $layer=LI1_cond $X=2.42 $Y=0.725
+ $X2=2.42 $Y2=2.18
r118 20 40 1.93381 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.87 $Y=2.265
+ $X2=0.705 $Y2=2.265
r119 19 42 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.335 $Y=2.265
+ $X2=2.42 $Y2=2.265
r120 19 20 95.5775 $w=1.68e-07 $l=1.465e-06 $layer=LI1_cond $X=2.335 $Y=2.265
+ $X2=0.87 $Y2=2.265
r121 15 40 4.50329 $w=2e-07 $l=1.07121e-07 $layer=LI1_cond $X=0.755 $Y=2.35
+ $X2=0.705 $Y2=2.265
r122 15 17 20.0425 $w=2.28e-07 $l=4e-07 $layer=LI1_cond $X=0.755 $Y=2.35
+ $X2=0.755 $Y2=2.75
r123 14 40 4.50329 $w=2e-07 $l=1.18427e-07 $layer=LI1_cond $X=0.625 $Y=2.18
+ $X2=0.705 $Y2=2.265
r124 13 38 6.36164 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=0.625 $Y=0.79
+ $X2=0.625 $Y2=0.57
r125 13 14 90.6845 $w=1.68e-07 $l=1.39e-06 $layer=LI1_cond $X=0.625 $Y=0.79
+ $X2=0.625 $Y2=2.18
r126 4 33 600 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=1 $X=3.19
+ $Y=2.315 $X2=3.335 $Y2=2.55
r127 3 17 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=0.575
+ $Y=2.54 $X2=0.725 $Y2=2.75
r128 2 29 182 $w=1.7e-07 $l=2.755e-07 $layer=licon1_NDIFF $count=1 $X=3.155
+ $Y=0.635 $X2=3.28 $Y2=0.855
r129 1 36 182 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_NDIFF $count=1 $X=0.165
+ $Y=0.37 $X2=0.31 $Y2=0.57
.ends

.subckt PM_SKY130_FD_SC_LS__DFRTN_1%Q 1 2 9 13 14 15 16 23 32
r26 21 23 1.31708 $w=3.48e-07 $l=4e-08 $layer=LI1_cond $X=10.78 $Y=1.995
+ $X2=10.78 $Y2=2.035
r27 15 16 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=10.78 $Y=2.405
+ $X2=10.78 $Y2=2.775
r28 14 21 0.75732 $w=3.48e-07 $l=2.3e-08 $layer=LI1_cond $X=10.78 $Y=1.972
+ $X2=10.78 $Y2=1.995
r29 14 32 8.06043 $w=3.48e-07 $l=1.52e-07 $layer=LI1_cond $X=10.78 $Y=1.972
+ $X2=10.78 $Y2=1.82
r30 14 15 11.4586 $w=3.48e-07 $l=3.48e-07 $layer=LI1_cond $X=10.78 $Y=2.057
+ $X2=10.78 $Y2=2.405
r31 14 23 0.724393 $w=3.48e-07 $l=2.2e-08 $layer=LI1_cond $X=10.78 $Y=2.057
+ $X2=10.78 $Y2=2.035
r32 13 32 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=10.87 $Y=1.15
+ $X2=10.87 $Y2=1.82
r33 7 13 9.06106 $w=3.63e-07 $l=1.82e-07 $layer=LI1_cond $X=10.772 $Y=0.968
+ $X2=10.772 $Y2=1.15
r34 7 9 11.4613 $w=3.63e-07 $l=3.63e-07 $layer=LI1_cond $X=10.772 $Y=0.968
+ $X2=10.772 $Y2=0.605
r35 2 14 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=10.62
+ $Y=1.84 $X2=10.77 $Y2=1.985
r36 2 16 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=10.62
+ $Y=1.84 $X2=10.77 $Y2=2.815
r37 1 9 91 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=2 $X=10.615
+ $Y=0.47 $X2=10.755 $Y2=0.605
.ends

.subckt PM_SKY130_FD_SC_LS__DFRTN_1%VGND 1 2 3 4 5 18 22 26 30 34 36 38 43 48 53
+ 61 71 72 75 78 81 84 87
r105 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r106 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r107 81 82 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r108 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r109 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r110 72 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=10.32 $Y2=0
r111 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=0 $X2=10.8
+ $Y2=0
r112 69 87 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.41 $Y=0
+ $X2=10.285 $Y2=0
r113 69 71 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=10.41 $Y=0 $X2=10.8
+ $Y2=0
r114 68 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=10.32 $Y2=0
r115 67 68 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r116 65 68 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=9.84
+ $Y2=0
r117 65 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=8.4
+ $Y2=0
r118 64 67 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=8.88 $Y=0 $X2=9.84
+ $Y2=0
r119 64 65 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r120 62 84 10.4332 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=8.555 $Y=0 $X2=8.335
+ $Y2=0
r121 62 64 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=8.555 $Y=0
+ $X2=8.88 $Y2=0
r122 61 87 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.16 $Y=0
+ $X2=10.285 $Y2=0
r123 61 67 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=10.16 $Y=0 $X2=9.84
+ $Y2=0
r124 60 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.4
+ $Y2=0
r125 59 60 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r126 56 59 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=5.52 $Y=0 $X2=7.92
+ $Y2=0
r127 54 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.355 $Y=0 $X2=5.19
+ $Y2=0
r128 54 56 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=5.355 $Y=0
+ $X2=5.52 $Y2=0
r129 53 84 10.4332 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=8.115 $Y=0 $X2=8.335
+ $Y2=0
r130 53 59 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=8.115 $Y=0
+ $X2=7.92 $Y2=0
r131 52 82 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=2.64 $Y=0 $X2=5.04
+ $Y2=0
r132 52 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r133 51 52 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r134 49 78 6.70225 $w=1.7e-07 $l=1.18e-07 $layer=LI1_cond $X=2.255 $Y=0
+ $X2=2.137 $Y2=0
r135 49 51 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=2.255 $Y=0
+ $X2=2.64 $Y2=0
r136 48 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.025 $Y=0 $X2=5.19
+ $Y2=0
r137 48 51 155.599 $w=1.68e-07 $l=2.385e-06 $layer=LI1_cond $X=5.025 $Y=0
+ $X2=2.64 $Y2=0
r138 47 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r139 47 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r140 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r141 44 75 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.295 $Y=0 $X2=1.17
+ $Y2=0
r142 44 46 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=1.295 $Y=0
+ $X2=1.68 $Y2=0
r143 43 78 6.70225 $w=1.7e-07 $l=1.17e-07 $layer=LI1_cond $X=2.02 $Y=0 $X2=2.137
+ $Y2=0
r144 43 46 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.02 $Y=0 $X2=1.68
+ $Y2=0
r145 41 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r146 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r147 38 75 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.045 $Y=0 $X2=1.17
+ $Y2=0
r148 38 40 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.045 $Y=0
+ $X2=0.72 $Y2=0
r149 36 60 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=5.52 $Y=0 $X2=7.92
+ $Y2=0
r150 36 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r151 36 56 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r152 32 87 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=10.285 $Y=0.085
+ $X2=10.285 $Y2=0
r153 32 34 23.9708 $w=2.48e-07 $l=5.2e-07 $layer=LI1_cond $X=10.285 $Y=0.085
+ $X2=10.285 $Y2=0.605
r154 28 84 1.73497 $w=4.4e-07 $l=8.5e-08 $layer=LI1_cond $X=8.335 $Y=0.085
+ $X2=8.335 $Y2=0
r155 28 30 17.1557 $w=4.38e-07 $l=6.55e-07 $layer=LI1_cond $X=8.335 $Y=0.085
+ $X2=8.335 $Y2=0.74
r156 24 81 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.19 $Y=0.085
+ $X2=5.19 $Y2=0
r157 24 26 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=5.19 $Y=0.085
+ $X2=5.19 $Y2=0.535
r158 20 78 0.207053 $w=2.35e-07 $l=8.5e-08 $layer=LI1_cond $X=2.137 $Y=0.085
+ $X2=2.137 $Y2=0
r159 20 22 10.5436 $w=2.33e-07 $l=2.15e-07 $layer=LI1_cond $X=2.137 $Y=0.085
+ $X2=2.137 $Y2=0.3
r160 16 75 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.17 $Y=0.085
+ $X2=1.17 $Y2=0
r161 16 18 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=1.17 $Y=0.085
+ $X2=1.17 $Y2=0.58
r162 5 34 91 $w=1.7e-07 $l=2.79464e-07 $layer=licon1_NDIFF $count=2 $X=10.105
+ $Y=0.47 $X2=10.325 $Y2=0.605
r163 4 30 182 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_NDIFF $count=1 $X=8.14
+ $Y=0.595 $X2=8.335 $Y2=0.74
r164 3 26 182 $w=1.7e-07 $l=2.6533e-07 $layer=licon1_NDIFF $count=1 $X=4.97
+ $Y=0.635 $X2=5.19 $Y2=0.535
r165 2 22 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=2.045
+ $Y=0.155 $X2=2.17 $Y2=0.3
r166 1 18 182 $w=1.7e-07 $l=3.07571e-07 $layer=licon1_NDIFF $count=1 $X=0.99
+ $Y=0.37 $X2=1.21 $Y2=0.58
.ends

