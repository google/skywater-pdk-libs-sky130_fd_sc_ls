* NGSPICE file created from sky130_fd_sc_ls__and3_4.ext - technology: sky130A

.subckt sky130_fd_sc_ls__and3_4 A B C VGND VNB VPB VPWR X
M1000 VPWR a_83_260# X VPB phighvt w=1.12e+06u l=150000u
+  ad=2.3268e+12p pd=1.666e+07u as=6.72e+11p ps=5.68e+06u
M1001 a_686_74# B a_489_74# VNB nshort w=640000u l=150000u
+  ad=5.76e+11p pd=5.64e+06u as=3.84e+11p ps=3.76e+06u
M1002 a_489_74# B a_686_74# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_83_260# C VPWR VPB phighvt w=840000u l=150000u
+  ad=7.896e+11p pd=6.92e+06u as=0p ps=0u
M1004 VPWR B a_83_260# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_83_260# A VPWR VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_489_74# C VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=9.013e+11p ps=8.26e+06u
M1007 a_83_260# A a_686_74# VNB nshort w=640000u l=150000u
+  ad=2.368e+11p pd=2.02e+06u as=0p ps=0u
M1008 VPWR A a_83_260# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND a_83_260# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=4.144e+11p ps=4.08e+06u
M1010 VPWR C a_83_260# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 X a_83_260# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR a_83_260# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND C a_489_74# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 X a_83_260# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 X a_83_260# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_83_260# B VPWR VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 X a_83_260# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND a_83_260# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_686_74# A a_83_260# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

