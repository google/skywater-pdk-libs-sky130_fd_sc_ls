* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__and4_4 A B C D VGND VNB VPB VPWR X
X0 a_116_392# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_116_392# A a_119_119# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X2 VPWR a_116_392# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X3 a_32_119# C a_463_119# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X4 VPWR C a_116_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_32_119# B a_119_119# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X6 VGND a_116_392# X VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X7 VPWR A a_116_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 X a_116_392# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X9 VPWR D a_116_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 X a_116_392# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X11 X a_116_392# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X12 VPWR B a_116_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 VPWR a_116_392# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X14 a_116_392# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 a_116_392# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 VGND D a_463_119# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X17 X a_116_392# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X18 a_119_119# A a_116_392# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X19 a_119_119# B a_32_119# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X20 a_463_119# D VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X21 VGND a_116_392# X VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X22 a_116_392# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X23 a_463_119# C a_32_119# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
.ends
