* File: sky130_fd_sc_ls__dlxtp_1.pxi.spice
* Created: Wed Sep  2 11:05:02 2020
* 
x_PM_SKY130_FD_SC_LS__DLXTP_1%D N_D_c_150_n N_D_M1009_g N_D_M1006_g N_D_c_147_n
+ D D N_D_c_149_n PM_SKY130_FD_SC_LS__DLXTP_1%D
x_PM_SKY130_FD_SC_LS__DLXTP_1%A_116_424# N_A_116_424#_M1006_d
+ N_A_116_424#_M1009_d N_A_116_424#_c_175_n N_A_116_424#_c_176_n
+ N_A_116_424#_c_185_n N_A_116_424#_M1011_g N_A_116_424#_c_177_n
+ N_A_116_424#_M1017_g N_A_116_424#_c_178_n N_A_116_424#_c_179_n
+ N_A_116_424#_c_186_n N_A_116_424#_c_187_n N_A_116_424#_c_180_n
+ N_A_116_424#_c_181_n N_A_116_424#_c_182_n N_A_116_424#_c_189_n
+ N_A_116_424#_c_183_n PM_SKY130_FD_SC_LS__DLXTP_1%A_116_424#
x_PM_SKY130_FD_SC_LS__DLXTP_1%A_386_326# N_A_386_326#_M1008_s
+ N_A_386_326#_M1001_s N_A_386_326#_c_258_n N_A_386_326#_M1015_g
+ N_A_386_326#_c_246_n N_A_386_326#_M1010_g N_A_386_326#_c_248_n
+ N_A_386_326#_M1016_g N_A_386_326#_M1004_g N_A_386_326#_c_250_n
+ N_A_386_326#_c_251_n N_A_386_326#_c_273_p N_A_386_326#_c_252_n
+ N_A_386_326#_c_253_n N_A_386_326#_c_254_n N_A_386_326#_c_255_n
+ N_A_386_326#_c_263_n N_A_386_326#_c_305_p N_A_386_326#_c_256_n
+ N_A_386_326#_c_257_n PM_SKY130_FD_SC_LS__DLXTP_1%A_386_326#
x_PM_SKY130_FD_SC_LS__DLXTP_1%A_562_123# N_A_562_123#_M1014_s
+ N_A_562_123#_M1007_s N_A_562_123#_M1003_g N_A_562_123#_c_388_n
+ N_A_562_123#_M1000_g N_A_562_123#_c_398_n N_A_562_123#_M1012_g
+ N_A_562_123#_M1002_g N_A_562_123#_c_390_n N_A_562_123#_c_391_n
+ N_A_562_123#_c_400_n N_A_562_123#_c_392_n N_A_562_123#_c_402_n
+ N_A_562_123#_c_403_n N_A_562_123#_c_431_p N_A_562_123#_c_404_n
+ N_A_562_123#_c_393_n N_A_562_123#_c_405_n N_A_562_123#_c_394_n
+ N_A_562_123#_c_395_n N_A_562_123#_c_396_n
+ PM_SKY130_FD_SC_LS__DLXTP_1%A_562_123#
x_PM_SKY130_FD_SC_LS__DLXTP_1%A_685_59# N_A_685_59#_M1002_d N_A_685_59#_M1012_d
+ N_A_685_59#_M1013_g N_A_685_59#_c_529_n N_A_685_59#_c_530_n
+ N_A_685_59#_M1005_g N_A_685_59#_c_521_n N_A_685_59#_c_522_n
+ N_A_685_59#_c_523_n N_A_685_59#_c_524_n N_A_685_59#_c_525_n
+ N_A_685_59#_c_526_n N_A_685_59#_c_533_n N_A_685_59#_c_534_n
+ N_A_685_59#_c_527_n N_A_685_59#_c_528_n PM_SKY130_FD_SC_LS__DLXTP_1%A_685_59#
x_PM_SKY130_FD_SC_LS__DLXTP_1%A_592_149# N_A_592_149#_M1003_d
+ N_A_592_149#_M1000_d N_A_592_149#_c_612_n N_A_592_149#_c_613_n
+ N_A_592_149#_c_614_n N_A_592_149#_c_624_n N_A_592_149#_M1001_g
+ N_A_592_149#_c_615_n N_A_592_149#_M1008_g N_A_592_149#_c_616_n
+ N_A_592_149#_c_617_n N_A_592_149#_c_643_n N_A_592_149#_c_626_n
+ N_A_592_149#_c_627_n N_A_592_149#_c_618_n N_A_592_149#_c_619_n
+ N_A_592_149#_c_620_n N_A_592_149#_c_621_n N_A_592_149#_c_622_n
+ PM_SKY130_FD_SC_LS__DLXTP_1%A_592_149#
x_PM_SKY130_FD_SC_LS__DLXTP_1%GATE N_GATE_M1014_g N_GATE_c_719_n N_GATE_M1007_g
+ GATE N_GATE_c_720_n PM_SKY130_FD_SC_LS__DLXTP_1%GATE
x_PM_SKY130_FD_SC_LS__DLXTP_1%VPWR N_VPWR_M1009_s N_VPWR_M1011_d N_VPWR_M1001_d
+ N_VPWR_M1007_d N_VPWR_c_752_n N_VPWR_c_753_n N_VPWR_c_754_n N_VPWR_c_755_n
+ VPWR N_VPWR_c_756_n N_VPWR_c_757_n N_VPWR_c_758_n N_VPWR_c_759_n
+ N_VPWR_c_751_n N_VPWR_c_761_n N_VPWR_c_762_n N_VPWR_c_763_n
+ PM_SKY130_FD_SC_LS__DLXTP_1%VPWR
x_PM_SKY130_FD_SC_LS__DLXTP_1%A_229_392# N_A_229_392#_M1011_s
+ N_A_229_392#_M1000_s N_A_229_392#_c_818_n N_A_229_392#_c_819_n
+ N_A_229_392#_c_820_n N_A_229_392#_c_821_n N_A_229_392#_c_822_n
+ PM_SKY130_FD_SC_LS__DLXTP_1%A_229_392#
x_PM_SKY130_FD_SC_LS__DLXTP_1%A_419_392# N_A_419_392#_M1015_d
+ N_A_419_392#_M1005_d N_A_419_392#_c_859_n N_A_419_392#_c_860_n
+ N_A_419_392#_c_861_n N_A_419_392#_c_877_n N_A_419_392#_c_880_n
+ N_A_419_392#_c_862_n N_A_419_392#_c_863_n N_A_419_392#_c_864_n
+ PM_SKY130_FD_SC_LS__DLXTP_1%A_419_392#
x_PM_SKY130_FD_SC_LS__DLXTP_1%Q N_Q_M1004_d N_Q_M1016_d N_Q_c_914_n N_Q_c_915_n
+ Q Q Q Q N_Q_c_916_n PM_SKY130_FD_SC_LS__DLXTP_1%Q
x_PM_SKY130_FD_SC_LS__DLXTP_1%VGND N_VGND_M1006_s N_VGND_M1017_d N_VGND_M1008_d
+ N_VGND_M1014_d N_VGND_c_936_n N_VGND_c_937_n N_VGND_c_938_n VGND
+ N_VGND_c_939_n N_VGND_c_940_n N_VGND_c_941_n N_VGND_c_942_n N_VGND_c_943_n
+ N_VGND_c_944_n N_VGND_c_945_n PM_SKY130_FD_SC_LS__DLXTP_1%VGND
x_PM_SKY130_FD_SC_LS__DLXTP_1%A_239_85# N_A_239_85#_M1017_s N_A_239_85#_M1013_d
+ N_A_239_85#_c_1002_n N_A_239_85#_c_1003_n N_A_239_85#_c_1004_n
+ N_A_239_85#_c_1005_n N_A_239_85#_c_1006_n N_A_239_85#_c_1032_n
+ N_A_239_85#_c_1036_n N_A_239_85#_c_1007_n N_A_239_85#_c_1008_n
+ N_A_239_85#_c_1009_n PM_SKY130_FD_SC_LS__DLXTP_1%A_239_85#
cc_1 VNB N_D_M1006_g 0.0293871f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.715
cc_2 VNB N_D_c_147_n 0.0255643f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.685
cc_3 VNB D 0.0216595f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_D_c_149_n 0.0185426f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.345
cc_5 VNB N_A_116_424#_c_175_n 0.0137405f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.18
cc_6 VNB N_A_116_424#_c_176_n 0.0185508f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_7 VNB N_A_116_424#_c_177_n 0.0195539f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.345
cc_8 VNB N_A_116_424#_c_178_n 0.0141747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_116_424#_c_179_n 0.0073213f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=1.665
cc_10 VNB N_A_116_424#_c_180_n 0.0212568f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_116_424#_c_181_n 0.00173165f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_116_424#_c_182_n 0.0421531f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_116_424#_c_183_n 5.29461e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_386_326#_c_246_n 0.0103436f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.685
cc_15 VNB N_A_386_326#_M1010_g 0.0288227f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.345
cc_16 VNB N_A_386_326#_c_248_n 0.0348926f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.345
cc_17 VNB N_A_386_326#_M1004_g 0.027505f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=1.345
cc_18 VNB N_A_386_326#_c_250_n 0.00571323f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_386_326#_c_251_n 0.0442704f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_386_326#_c_252_n 0.00398307f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_386_326#_c_253_n 0.00773815f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_386_326#_c_254_n 0.00331008f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_386_326#_c_255_n 0.00461843f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_386_326#_c_256_n 0.00264351f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_386_326#_c_257_n 0.0537079f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_562_123#_M1003_g 0.0249529f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.18
cc_27 VNB N_A_562_123#_c_388_n 0.0227058f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_28 VNB N_A_562_123#_M1002_g 0.0277582f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_562_123#_c_390_n 0.0256723f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=1.345
cc_30 VNB N_A_562_123#_c_391_n 0.0177402f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=1.665
cc_31 VNB N_A_562_123#_c_392_n 0.00541649f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_562_123#_c_393_n 0.00260442f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_562_123#_c_394_n 0.00393894f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_562_123#_c_395_n 0.0107544f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_562_123#_c_396_n 0.0251887f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_685_59#_c_521_n 0.0186701f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.345
cc_37 VNB N_A_685_59#_c_522_n 0.0217776f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.345
cc_38 VNB N_A_685_59#_c_523_n 0.0029799f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_685_59#_c_524_n 0.0064491f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=1.345
cc_40 VNB N_A_685_59#_c_525_n 0.0204596f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_685_59#_c_526_n 0.00246741f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_685_59#_c_527_n 0.00456952f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_685_59#_c_528_n 0.00480596f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_592_149#_c_612_n 0.0137834f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_592_149#_c_613_n 0.0209814f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.345
cc_46 VNB N_A_592_149#_c_614_n 0.00857213f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.685
cc_47 VNB N_A_592_149#_c_615_n 0.0171293f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_592_149#_c_616_n 0.0195486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_592_149#_c_617_n 0.00290329f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=1.665
cc_50 VNB N_A_592_149#_c_618_n 0.00448004f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_592_149#_c_619_n 0.00220735f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_592_149#_c_620_n 0.00402759f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_592_149#_c_621_n 0.00372743f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_592_149#_c_622_n 0.045578f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_GATE_M1014_g 0.0288503f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.54
cc_56 VNB N_GATE_c_719_n 0.0243079f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.715
cc_57 VNB N_GATE_c_720_n 0.00505132f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_58 VNB N_VPWR_c_751_n 0.322901f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_Q_c_914_n 0.0260019f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.18
cc_60 VNB N_Q_c_915_n 0.00874531f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_Q_c_916_n 0.0237646f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_936_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_937_n 0.0439288f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.345
cc_64 VNB N_VGND_c_938_n 0.0202602f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_939_n 0.0345439f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_940_n 0.0691667f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_941_n 0.0542831f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_942_n 0.0194271f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_943_n 0.442226f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_944_n 0.00634414f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_945_n 0.0158736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_239_85#_c_1002_n 0.00675372f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.18
cc_73 VNB N_A_239_85#_c_1003_n 0.00103024f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_74 VNB N_A_239_85#_c_1004_n 0.0275945f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_239_85#_c_1005_n 0.00205182f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_239_85#_c_1006_n 0.00419449f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.345
cc_77 VNB N_A_239_85#_c_1007_n 0.00623433f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=1.345
cc_78 VNB N_A_239_85#_c_1008_n 0.0027321f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_239_85#_c_1009_n 0.00286487f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VPB N_D_c_150_n 0.0222056f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.045
cc_81 VPB N_D_c_147_n 0.0389278f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.685
cc_82 VPB D 0.0105206f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_83 VPB N_A_116_424#_c_176_n 0.00786178f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_84 VPB N_A_116_424#_c_185_n 0.0278815f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_A_116_424#_c_186_n 0.00703133f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_A_116_424#_c_187_n 0.0100658f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_A_116_424#_c_182_n 0.0163485f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_A_116_424#_c_189_n 0.00711835f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_A_116_424#_c_183_n 0.00839962f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB N_A_386_326#_c_258_n 0.0170091f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB N_A_386_326#_c_246_n 0.0193107f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.685
cc_92 VPB N_A_386_326#_c_248_n 0.0295185f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.345
cc_93 VPB N_A_386_326#_c_250_n 0.0130076f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB N_A_386_326#_c_252_n 0.00426023f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_95 VPB N_A_386_326#_c_263_n 0.00657379f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB N_A_562_123#_c_388_n 0.0417724f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_97 VPB N_A_562_123#_c_398_n 0.0168624f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_A_562_123#_c_391_n 0.00744684f $X=-0.19 $Y=1.66 $X2=0.36 $Y2=1.665
cc_99 VPB N_A_562_123#_c_400_n 0.00508842f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 VPB N_A_562_123#_c_392_n 0.00467423f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB N_A_562_123#_c_402_n 0.00992746f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_102 VPB N_A_562_123#_c_403_n 0.0168443f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 VPB N_A_562_123#_c_404_n 0.00585209f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB N_A_562_123#_c_405_n 0.040563f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_105 VPB N_A_562_123#_c_396_n 0.0147743f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_A_685_59#_c_529_n 0.0408224f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_107 VPB N_A_685_59#_c_530_n 0.0268779f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_108 VPB N_A_685_59#_c_523_n 0.0177586f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_109 VPB N_A_685_59#_c_526_n 0.0107548f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_110 VPB N_A_685_59#_c_533_n 0.00890014f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_A_685_59#_c_534_n 0.00374796f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_A_685_59#_c_527_n 0.00122718f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_A_592_149#_c_614_n 9.30309e-19 $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.685
cc_114 VPB N_A_592_149#_c_624_n 0.02624f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_115 VPB N_A_592_149#_c_617_n 0.00405557f $X=-0.19 $Y=1.66 $X2=0.36 $Y2=1.665
cc_116 VPB N_A_592_149#_c_626_n 0.0063065f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_A_592_149#_c_627_n 0.00156376f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_GATE_c_719_n 0.0324622f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=0.715
cc_119 VPB N_GATE_c_720_n 0.00575224f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_120 VPB N_VPWR_c_752_n 0.0120106f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_753_n 0.0459344f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.345
cc_122 VPB N_VPWR_c_754_n 0.0213835f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_755_n 0.0202785f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_756_n 0.0324821f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_757_n 0.0723317f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_758_n 0.043529f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_759_n 0.0190372f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_751_n 0.109586f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_761_n 0.016933f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_762_n 0.00631563f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_VPWR_c_763_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_A_229_392#_c_818_n 0.0121389f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.18
cc_133 VPB N_A_229_392#_c_819_n 0.0115889f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.345
cc_134 VPB N_A_229_392#_c_820_n 0.00578657f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.345
cc_135 VPB N_A_229_392#_c_821_n 0.00991886f $X=-0.19 $Y=1.66 $X2=0.36 $Y2=1.345
cc_136 VPB N_A_229_392#_c_822_n 0.0102748f $X=-0.19 $Y=1.66 $X2=0.36 $Y2=1.665
cc_137 VPB N_A_419_392#_c_859_n 0.00214599f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.18
cc_138 VPB N_A_419_392#_c_860_n 0.00461189f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_139 VPB N_A_419_392#_c_861_n 0.00231845f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_140 VPB N_A_419_392#_c_862_n 0.00216417f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.345
cc_141 VPB N_A_419_392#_c_863_n 0.00725767f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_142 VPB N_A_419_392#_c_864_n 0.00735108f $X=-0.19 $Y=1.66 $X2=0.36 $Y2=1.345
cc_143 VPB Q 0.00991834f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_144 VPB Q 0.0418938f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_145 VPB N_Q_c_916_n 0.00776232f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_146 N_D_M1006_g N_A_116_424#_c_179_n 0.00205721f $X=0.52 $Y=0.715 $X2=0 $Y2=0
cc_147 N_D_c_150_n N_A_116_424#_c_186_n 0.00694909f $X=0.505 $Y=2.045 $X2=0
+ $Y2=0
cc_148 N_D_M1006_g N_A_116_424#_c_180_n 0.00771334f $X=0.52 $Y=0.715 $X2=0 $Y2=0
cc_149 D N_A_116_424#_c_180_n 0.0091069f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_150 D N_A_116_424#_c_181_n 0.0431681f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_151 N_D_c_149_n N_A_116_424#_c_181_n 0.00571717f $X=0.43 $Y=1.345 $X2=0 $Y2=0
cc_152 N_D_M1006_g N_A_116_424#_c_182_n 0.017533f $X=0.52 $Y=0.715 $X2=0 $Y2=0
cc_153 D N_A_116_424#_c_182_n 6.6718e-19 $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_154 N_D_c_149_n N_A_116_424#_c_182_n 0.017533f $X=0.43 $Y=1.345 $X2=0 $Y2=0
cc_155 N_D_c_150_n N_A_116_424#_c_189_n 0.00179961f $X=0.505 $Y=2.045 $X2=0
+ $Y2=0
cc_156 N_D_c_147_n N_A_116_424#_c_183_n 0.00571717f $X=0.43 $Y=1.685 $X2=0 $Y2=0
cc_157 N_D_c_150_n N_VPWR_c_753_n 0.0208523f $X=0.505 $Y=2.045 $X2=0 $Y2=0
cc_158 N_D_c_147_n N_VPWR_c_753_n 0.00161586f $X=0.43 $Y=1.685 $X2=0 $Y2=0
cc_159 D N_VPWR_c_753_n 0.0217756f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_160 N_D_c_150_n N_VPWR_c_756_n 0.00413917f $X=0.505 $Y=2.045 $X2=0 $Y2=0
cc_161 N_D_c_150_n N_VPWR_c_751_n 0.00822528f $X=0.505 $Y=2.045 $X2=0 $Y2=0
cc_162 N_D_M1006_g N_VGND_c_937_n 0.00912487f $X=0.52 $Y=0.715 $X2=0 $Y2=0
cc_163 D N_VGND_c_937_n 0.0289511f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_164 N_D_c_149_n N_VGND_c_937_n 0.00140112f $X=0.43 $Y=1.345 $X2=0 $Y2=0
cc_165 N_D_M1006_g N_VGND_c_939_n 0.00526206f $X=0.52 $Y=0.715 $X2=0 $Y2=0
cc_166 N_D_M1006_g N_VGND_c_943_n 0.00523671f $X=0.52 $Y=0.715 $X2=0 $Y2=0
cc_167 N_D_M1006_g N_A_239_85#_c_1002_n 0.00118246f $X=0.52 $Y=0.715 $X2=0 $Y2=0
cc_168 N_A_116_424#_c_185_n N_A_386_326#_c_258_n 0.020051f $X=1.515 $Y=1.885
+ $X2=0 $Y2=0
cc_169 N_A_116_424#_c_176_n N_A_386_326#_c_250_n 0.0123399f $X=1.515 $Y=1.795
+ $X2=0 $Y2=0
cc_170 N_A_116_424#_c_177_n N_A_386_326#_c_257_n 0.00458971f $X=1.6 $Y=1.24
+ $X2=0 $Y2=0
cc_171 N_A_116_424#_c_186_n N_VPWR_c_753_n 0.05986f $X=0.795 $Y=2.25 $X2=0 $Y2=0
cc_172 N_A_116_424#_c_185_n N_VPWR_c_756_n 0.00314797f $X=1.515 $Y=1.885 $X2=0
+ $Y2=0
cc_173 N_A_116_424#_c_187_n N_VPWR_c_756_n 0.013297f $X=0.73 $Y=2.265 $X2=0
+ $Y2=0
cc_174 N_A_116_424#_c_185_n N_VPWR_c_751_n 0.00397822f $X=1.515 $Y=1.885 $X2=0
+ $Y2=0
cc_175 N_A_116_424#_c_187_n N_VPWR_c_751_n 0.0110061f $X=0.73 $Y=2.265 $X2=0
+ $Y2=0
cc_176 N_A_116_424#_c_185_n N_VPWR_c_761_n 0.00508459f $X=1.515 $Y=1.885 $X2=0
+ $Y2=0
cc_177 N_A_116_424#_c_175_n N_A_229_392#_c_818_n 0.00221207f $X=1.425 $Y=1.315
+ $X2=0 $Y2=0
cc_178 N_A_116_424#_c_185_n N_A_229_392#_c_818_n 0.016306f $X=1.515 $Y=1.885
+ $X2=0 $Y2=0
cc_179 N_A_116_424#_c_182_n N_A_229_392#_c_818_n 2.97498e-19 $X=1 $Y=1.265 $X2=0
+ $Y2=0
cc_180 N_A_116_424#_c_189_n N_A_229_392#_c_818_n 0.0409741f $X=0.795 $Y=2.1
+ $X2=0 $Y2=0
cc_181 N_A_116_424#_c_183_n N_A_229_392#_c_818_n 0.00338425f $X=0.97 $Y=1.77
+ $X2=0 $Y2=0
cc_182 N_A_116_424#_c_185_n N_A_229_392#_c_820_n 0.00880689f $X=1.515 $Y=1.885
+ $X2=0 $Y2=0
cc_183 N_A_116_424#_c_186_n N_A_229_392#_c_820_n 0.0409741f $X=0.795 $Y=2.25
+ $X2=0 $Y2=0
cc_184 N_A_116_424#_c_185_n N_A_229_392#_c_821_n 0.0151578f $X=1.515 $Y=1.885
+ $X2=0 $Y2=0
cc_185 N_A_116_424#_c_185_n N_A_229_392#_c_822_n 0.00462681f $X=1.515 $Y=1.885
+ $X2=0 $Y2=0
cc_186 N_A_116_424#_c_185_n N_A_419_392#_c_859_n 0.00101945f $X=1.515 $Y=1.885
+ $X2=0 $Y2=0
cc_187 N_A_116_424#_c_185_n N_A_419_392#_c_861_n 5.16815e-19 $X=1.515 $Y=1.885
+ $X2=0 $Y2=0
cc_188 N_A_116_424#_c_179_n N_VGND_c_937_n 0.0151023f $X=0.78 $Y=0.715 $X2=0
+ $Y2=0
cc_189 N_A_116_424#_c_180_n N_VGND_c_937_n 0.00430388f $X=0.97 $Y=1.295 $X2=0
+ $Y2=0
cc_190 N_A_116_424#_c_177_n N_VGND_c_938_n 0.00930917f $X=1.6 $Y=1.24 $X2=0
+ $Y2=0
cc_191 N_A_116_424#_c_177_n N_VGND_c_939_n 0.00536686f $X=1.6 $Y=1.24 $X2=0
+ $Y2=0
cc_192 N_A_116_424#_c_179_n N_VGND_c_939_n 0.0113526f $X=0.78 $Y=0.715 $X2=0
+ $Y2=0
cc_193 N_A_116_424#_c_177_n N_VGND_c_943_n 0.00528353f $X=1.6 $Y=1.24 $X2=0
+ $Y2=0
cc_194 N_A_116_424#_c_179_n N_VGND_c_943_n 0.0115594f $X=0.78 $Y=0.715 $X2=0
+ $Y2=0
cc_195 N_A_116_424#_c_177_n N_A_239_85#_c_1002_n 0.00749565f $X=1.6 $Y=1.24
+ $X2=0 $Y2=0
cc_196 N_A_116_424#_c_179_n N_A_239_85#_c_1002_n 0.0285858f $X=0.78 $Y=0.715
+ $X2=0 $Y2=0
cc_197 N_A_116_424#_c_175_n N_A_239_85#_c_1003_n 0.00471495f $X=1.425 $Y=1.315
+ $X2=0 $Y2=0
cc_198 N_A_116_424#_c_178_n N_A_239_85#_c_1003_n 0.00524714f $X=1.55 $Y=1.315
+ $X2=0 $Y2=0
cc_199 N_A_116_424#_c_180_n N_A_239_85#_c_1003_n 0.0217614f $X=0.97 $Y=1.295
+ $X2=0 $Y2=0
cc_200 N_A_116_424#_c_181_n N_A_239_85#_c_1003_n 0.00427066f $X=0.97 $Y=1.575
+ $X2=0 $Y2=0
cc_201 N_A_116_424#_c_182_n N_A_239_85#_c_1003_n 4.73506e-19 $X=1 $Y=1.265 $X2=0
+ $Y2=0
cc_202 N_A_116_424#_c_176_n N_A_239_85#_c_1004_n 0.00878425f $X=1.515 $Y=1.795
+ $X2=0 $Y2=0
cc_203 N_A_116_424#_c_178_n N_A_239_85#_c_1004_n 0.0098925f $X=1.55 $Y=1.315
+ $X2=0 $Y2=0
cc_204 N_A_116_424#_c_175_n N_A_239_85#_c_1005_n 8.00681e-19 $X=1.425 $Y=1.315
+ $X2=0 $Y2=0
cc_205 N_A_116_424#_c_176_n N_A_239_85#_c_1005_n 0.00499084f $X=1.515 $Y=1.795
+ $X2=0 $Y2=0
cc_206 N_A_116_424#_c_178_n N_A_239_85#_c_1005_n 2.6366e-19 $X=1.55 $Y=1.315
+ $X2=0 $Y2=0
cc_207 N_A_116_424#_c_181_n N_A_239_85#_c_1005_n 0.0143061f $X=0.97 $Y=1.575
+ $X2=0 $Y2=0
cc_208 N_A_116_424#_c_182_n N_A_239_85#_c_1005_n 9.1358e-19 $X=1 $Y=1.265 $X2=0
+ $Y2=0
cc_209 N_A_116_424#_c_177_n N_A_239_85#_c_1006_n 0.00360374f $X=1.6 $Y=1.24
+ $X2=0 $Y2=0
cc_210 N_A_116_424#_c_175_n N_A_239_85#_c_1008_n 0.00589353f $X=1.425 $Y=1.315
+ $X2=0 $Y2=0
cc_211 N_A_116_424#_c_180_n N_A_239_85#_c_1008_n 0.00575056f $X=0.97 $Y=1.295
+ $X2=0 $Y2=0
cc_212 N_A_386_326#_c_253_n N_A_562_123#_M1014_s 0.00758073f $X=6.895 $Y=0.665
+ $X2=-0.19 $Y2=-0.245
cc_213 N_A_386_326#_M1010_g N_A_562_123#_M1003_g 0.0300741f $X=2.495 $Y=0.955
+ $X2=0 $Y2=0
cc_214 N_A_386_326#_c_251_n N_A_562_123#_M1003_g 9.7971e-19 $X=4.565 $Y=0.34
+ $X2=0 $Y2=0
cc_215 N_A_386_326#_c_246_n N_A_562_123#_c_388_n 0.0305045f $X=2.42 $Y=1.705
+ $X2=0 $Y2=0
cc_216 N_A_386_326#_c_252_n N_A_562_123#_c_398_n 4.15804e-19 $X=4.69 $Y=1.665
+ $X2=0 $Y2=0
cc_217 N_A_386_326#_c_263_n N_A_562_123#_c_398_n 0.00117923f $X=4.69 $Y=1.83
+ $X2=0 $Y2=0
cc_218 N_A_386_326#_c_273_p N_A_562_123#_M1002_g 6.97948e-19 $X=4.65 $Y=0.555
+ $X2=0 $Y2=0
cc_219 N_A_386_326#_c_252_n N_A_562_123#_M1002_g 0.0012083f $X=4.69 $Y=1.665
+ $X2=0 $Y2=0
cc_220 N_A_386_326#_c_253_n N_A_562_123#_M1002_g 0.0140652f $X=6.895 $Y=0.665
+ $X2=0 $Y2=0
cc_221 N_A_386_326#_c_253_n N_A_562_123#_c_390_n 4.45051e-19 $X=6.895 $Y=0.665
+ $X2=0 $Y2=0
cc_222 N_A_386_326#_c_252_n N_A_562_123#_c_391_n 0.00207833f $X=4.69 $Y=1.665
+ $X2=0 $Y2=0
cc_223 N_A_386_326#_c_253_n N_A_562_123#_c_391_n 0.00337467f $X=6.895 $Y=0.665
+ $X2=0 $Y2=0
cc_224 N_A_386_326#_M1010_g N_A_562_123#_c_392_n 3.11059e-19 $X=2.495 $Y=0.955
+ $X2=0 $Y2=0
cc_225 N_A_386_326#_M1001_s N_A_562_123#_c_403_n 0.00916709f $X=4.29 $Y=1.685
+ $X2=0 $Y2=0
cc_226 N_A_386_326#_c_253_n N_A_562_123#_c_393_n 0.00484455f $X=6.895 $Y=0.665
+ $X2=0 $Y2=0
cc_227 N_A_386_326#_c_253_n N_A_562_123#_c_395_n 0.0260907f $X=6.895 $Y=0.665
+ $X2=0 $Y2=0
cc_228 N_A_386_326#_c_254_n N_A_562_123#_c_395_n 0.00828008f $X=6.98 $Y=1.32
+ $X2=0 $Y2=0
cc_229 N_A_386_326#_c_253_n N_A_562_123#_c_396_n 8.08962e-19 $X=6.895 $Y=0.665
+ $X2=0 $Y2=0
cc_230 N_A_386_326#_c_253_n N_A_685_59#_M1002_d 0.00691035f $X=6.895 $Y=0.665
+ $X2=-0.19 $Y2=-0.245
cc_231 N_A_386_326#_c_251_n N_A_685_59#_c_521_n 0.0123027f $X=4.565 $Y=0.34
+ $X2=0 $Y2=0
cc_232 N_A_386_326#_c_252_n N_A_685_59#_c_524_n 0.0106374f $X=4.69 $Y=1.665
+ $X2=0 $Y2=0
cc_233 N_A_386_326#_c_252_n N_A_685_59#_c_526_n 0.00462326f $X=4.69 $Y=1.665
+ $X2=0 $Y2=0
cc_234 N_A_386_326#_c_263_n N_A_685_59#_c_526_n 0.0272018f $X=4.69 $Y=1.83 $X2=0
+ $Y2=0
cc_235 N_A_386_326#_M1001_s N_A_685_59#_c_533_n 0.00721306f $X=4.29 $Y=1.685
+ $X2=0 $Y2=0
cc_236 N_A_386_326#_c_263_n N_A_685_59#_c_533_n 0.0331232f $X=4.69 $Y=1.83 $X2=0
+ $Y2=0
cc_237 N_A_386_326#_c_252_n N_A_685_59#_c_527_n 0.015174f $X=4.69 $Y=1.665 $X2=0
+ $Y2=0
cc_238 N_A_386_326#_c_263_n N_A_685_59#_c_527_n 0.00478602f $X=4.69 $Y=1.83
+ $X2=0 $Y2=0
cc_239 N_A_386_326#_c_252_n N_A_685_59#_c_528_n 0.00369591f $X=4.69 $Y=1.665
+ $X2=0 $Y2=0
cc_240 N_A_386_326#_c_253_n N_A_685_59#_c_528_n 0.0290457f $X=6.895 $Y=0.665
+ $X2=0 $Y2=0
cc_241 N_A_386_326#_c_252_n N_A_592_149#_c_612_n 0.00681063f $X=4.69 $Y=1.665
+ $X2=0 $Y2=0
cc_242 N_A_386_326#_c_263_n N_A_592_149#_c_613_n 0.00941891f $X=4.69 $Y=1.83
+ $X2=0 $Y2=0
cc_243 N_A_386_326#_c_252_n N_A_592_149#_c_614_n 0.00554298f $X=4.69 $Y=1.665
+ $X2=0 $Y2=0
cc_244 N_A_386_326#_c_252_n N_A_592_149#_c_624_n 0.00643165f $X=4.69 $Y=1.665
+ $X2=0 $Y2=0
cc_245 N_A_386_326#_c_263_n N_A_592_149#_c_624_n 0.0104706f $X=4.69 $Y=1.83
+ $X2=0 $Y2=0
cc_246 N_A_386_326#_c_251_n N_A_592_149#_c_615_n 0.005196f $X=4.565 $Y=0.34
+ $X2=0 $Y2=0
cc_247 N_A_386_326#_c_273_p N_A_592_149#_c_615_n 0.00307059f $X=4.65 $Y=0.555
+ $X2=0 $Y2=0
cc_248 N_A_386_326#_c_252_n N_A_592_149#_c_615_n 0.0107557f $X=4.69 $Y=1.665
+ $X2=0 $Y2=0
cc_249 N_A_386_326#_c_253_n N_A_592_149#_c_615_n 0.0123434f $X=6.895 $Y=0.665
+ $X2=0 $Y2=0
cc_250 N_A_386_326#_c_305_p N_A_592_149#_c_615_n 3.84191e-19 $X=4.69 $Y=0.665
+ $X2=0 $Y2=0
cc_251 N_A_386_326#_c_252_n N_A_592_149#_c_616_n 0.00837347f $X=4.69 $Y=1.665
+ $X2=0 $Y2=0
cc_252 N_A_386_326#_c_258_n N_A_592_149#_c_617_n 0.00128813f $X=2.02 $Y=1.885
+ $X2=0 $Y2=0
cc_253 N_A_386_326#_c_246_n N_A_592_149#_c_617_n 0.00909586f $X=2.42 $Y=1.705
+ $X2=0 $Y2=0
cc_254 N_A_386_326#_M1010_g N_A_592_149#_c_617_n 0.0103388f $X=2.495 $Y=0.955
+ $X2=0 $Y2=0
cc_255 N_A_386_326#_c_250_n N_A_592_149#_c_617_n 0.00286215f $X=2.02 $Y=1.705
+ $X2=0 $Y2=0
cc_256 N_A_386_326#_M1010_g N_A_592_149#_c_643_n 0.00470683f $X=2.495 $Y=0.955
+ $X2=0 $Y2=0
cc_257 N_A_386_326#_c_258_n N_A_592_149#_c_626_n 5.66015e-19 $X=2.02 $Y=1.885
+ $X2=0 $Y2=0
cc_258 N_A_386_326#_c_251_n N_A_592_149#_c_618_n 0.00598461f $X=4.565 $Y=0.34
+ $X2=0 $Y2=0
cc_259 N_A_386_326#_c_251_n N_A_592_149#_c_621_n 0.0126277f $X=4.565 $Y=0.34
+ $X2=0 $Y2=0
cc_260 N_A_386_326#_c_252_n N_A_592_149#_c_621_n 0.025079f $X=4.69 $Y=1.665
+ $X2=0 $Y2=0
cc_261 N_A_386_326#_c_263_n N_A_592_149#_c_621_n 0.00399806f $X=4.69 $Y=1.83
+ $X2=0 $Y2=0
cc_262 N_A_386_326#_c_251_n N_A_592_149#_c_622_n 0.00196387f $X=4.565 $Y=0.34
+ $X2=0 $Y2=0
cc_263 N_A_386_326#_c_252_n N_A_592_149#_c_622_n 0.00549048f $X=4.69 $Y=1.665
+ $X2=0 $Y2=0
cc_264 N_A_386_326#_c_248_n N_GATE_M1014_g 8.08286e-19 $X=7.17 $Y=1.765 $X2=0
+ $Y2=0
cc_265 N_A_386_326#_M1004_g N_GATE_M1014_g 0.0152937f $X=7.185 $Y=0.78 $X2=0
+ $Y2=0
cc_266 N_A_386_326#_c_253_n N_GATE_M1014_g 0.016091f $X=6.895 $Y=0.665 $X2=0
+ $Y2=0
cc_267 N_A_386_326#_c_254_n N_GATE_M1014_g 0.00801253f $X=6.98 $Y=1.32 $X2=0
+ $Y2=0
cc_268 N_A_386_326#_c_256_n N_GATE_M1014_g 5.77738e-19 $X=7.09 $Y=1.485 $X2=0
+ $Y2=0
cc_269 N_A_386_326#_c_248_n N_GATE_c_719_n 0.0430027f $X=7.17 $Y=1.765 $X2=0
+ $Y2=0
cc_270 N_A_386_326#_c_253_n N_GATE_c_719_n 7.23523e-19 $X=6.895 $Y=0.665 $X2=0
+ $Y2=0
cc_271 N_A_386_326#_c_256_n N_GATE_c_719_n 0.00170854f $X=7.09 $Y=1.485 $X2=0
+ $Y2=0
cc_272 N_A_386_326#_c_248_n N_GATE_c_720_n 0.0025254f $X=7.17 $Y=1.765 $X2=0
+ $Y2=0
cc_273 N_A_386_326#_c_253_n N_GATE_c_720_n 0.0074181f $X=6.895 $Y=0.665 $X2=0
+ $Y2=0
cc_274 N_A_386_326#_c_256_n N_GATE_c_720_n 0.0230297f $X=7.09 $Y=1.485 $X2=0
+ $Y2=0
cc_275 N_A_386_326#_c_248_n N_VPWR_c_755_n 0.0163842f $X=7.17 $Y=1.765 $X2=0
+ $Y2=0
cc_276 N_A_386_326#_c_256_n N_VPWR_c_755_n 0.00826396f $X=7.09 $Y=1.485 $X2=0
+ $Y2=0
cc_277 N_A_386_326#_c_248_n N_VPWR_c_759_n 0.00445602f $X=7.17 $Y=1.765 $X2=0
+ $Y2=0
cc_278 N_A_386_326#_c_248_n N_VPWR_c_751_n 0.0086523f $X=7.17 $Y=1.765 $X2=0
+ $Y2=0
cc_279 N_A_386_326#_c_258_n N_A_229_392#_c_818_n 0.00183633f $X=2.02 $Y=1.885
+ $X2=0 $Y2=0
cc_280 N_A_386_326#_c_258_n N_A_229_392#_c_821_n 0.00643965f $X=2.02 $Y=1.885
+ $X2=0 $Y2=0
cc_281 N_A_386_326#_c_258_n N_A_419_392#_c_859_n 0.00716039f $X=2.02 $Y=1.885
+ $X2=0 $Y2=0
cc_282 N_A_386_326#_c_246_n N_A_419_392#_c_859_n 0.00511664f $X=2.42 $Y=1.705
+ $X2=0 $Y2=0
cc_283 N_A_386_326#_c_250_n N_A_419_392#_c_859_n 4.41735e-19 $X=2.02 $Y=1.705
+ $X2=0 $Y2=0
cc_284 N_A_386_326#_c_246_n N_A_419_392#_c_860_n 0.00467553f $X=2.42 $Y=1.705
+ $X2=0 $Y2=0
cc_285 N_A_386_326#_c_258_n N_A_419_392#_c_861_n 0.00495686f $X=2.02 $Y=1.885
+ $X2=0 $Y2=0
cc_286 N_A_386_326#_c_258_n N_A_419_392#_c_864_n 0.00197423f $X=2.02 $Y=1.885
+ $X2=0 $Y2=0
cc_287 N_A_386_326#_c_246_n N_A_419_392#_c_864_n 4.94042e-19 $X=2.42 $Y=1.705
+ $X2=0 $Y2=0
cc_288 N_A_386_326#_M1004_g N_Q_c_914_n 0.0132797f $X=7.185 $Y=0.78 $X2=0 $Y2=0
cc_289 N_A_386_326#_M1004_g N_Q_c_915_n 0.0021929f $X=7.185 $Y=0.78 $X2=0 $Y2=0
cc_290 N_A_386_326#_c_256_n N_Q_c_915_n 0.00151667f $X=7.09 $Y=1.485 $X2=0 $Y2=0
cc_291 N_A_386_326#_c_248_n Q 0.00422325f $X=7.17 $Y=1.765 $X2=0 $Y2=0
cc_292 N_A_386_326#_c_256_n Q 0.00196075f $X=7.09 $Y=1.485 $X2=0 $Y2=0
cc_293 N_A_386_326#_c_248_n Q 0.0110598f $X=7.17 $Y=1.765 $X2=0 $Y2=0
cc_294 N_A_386_326#_M1004_g N_Q_c_916_n 0.0140755f $X=7.185 $Y=0.78 $X2=0 $Y2=0
cc_295 N_A_386_326#_c_254_n N_Q_c_916_n 0.00535893f $X=6.98 $Y=1.32 $X2=0 $Y2=0
cc_296 N_A_386_326#_c_256_n N_Q_c_916_n 0.0249377f $X=7.09 $Y=1.485 $X2=0 $Y2=0
cc_297 N_A_386_326#_c_253_n N_VGND_M1008_d 0.0143787f $X=6.895 $Y=0.665 $X2=0
+ $Y2=0
cc_298 N_A_386_326#_c_253_n N_VGND_M1014_d 0.0168228f $X=6.895 $Y=0.665 $X2=0
+ $Y2=0
cc_299 N_A_386_326#_c_254_n N_VGND_M1014_d 0.00893215f $X=6.98 $Y=1.32 $X2=0
+ $Y2=0
cc_300 N_A_386_326#_M1010_g N_VGND_c_938_n 0.0026503f $X=2.495 $Y=0.955 $X2=0
+ $Y2=0
cc_301 N_A_386_326#_c_255_n N_VGND_c_938_n 0.026116f $X=2.34 $Y=0.34 $X2=0 $Y2=0
cc_302 N_A_386_326#_c_257_n N_VGND_c_938_n 0.00367328f $X=2.495 $Y=0.42 $X2=0
+ $Y2=0
cc_303 N_A_386_326#_c_251_n N_VGND_c_940_n 0.150405f $X=4.565 $Y=0.34 $X2=0
+ $Y2=0
cc_304 N_A_386_326#_c_253_n N_VGND_c_940_n 0.00294479f $X=6.895 $Y=0.665 $X2=0
+ $Y2=0
cc_305 N_A_386_326#_c_255_n N_VGND_c_940_n 0.0212434f $X=2.34 $Y=0.34 $X2=0
+ $Y2=0
cc_306 N_A_386_326#_c_257_n N_VGND_c_940_n 0.00386462f $X=2.495 $Y=0.42 $X2=0
+ $Y2=0
cc_307 N_A_386_326#_M1004_g N_VGND_c_941_n 0.00379265f $X=7.185 $Y=0.78 $X2=0
+ $Y2=0
cc_308 N_A_386_326#_c_253_n N_VGND_c_941_n 0.0587995f $X=6.895 $Y=0.665 $X2=0
+ $Y2=0
cc_309 N_A_386_326#_M1004_g N_VGND_c_942_n 0.00523933f $X=7.185 $Y=0.78 $X2=0
+ $Y2=0
cc_310 N_A_386_326#_M1004_g N_VGND_c_943_n 0.00533081f $X=7.185 $Y=0.78 $X2=0
+ $Y2=0
cc_311 N_A_386_326#_c_251_n N_VGND_c_943_n 0.0871302f $X=4.565 $Y=0.34 $X2=0
+ $Y2=0
cc_312 N_A_386_326#_c_253_n N_VGND_c_943_n 0.0471749f $X=6.895 $Y=0.665 $X2=0
+ $Y2=0
cc_313 N_A_386_326#_c_255_n N_VGND_c_943_n 0.0123341f $X=2.34 $Y=0.34 $X2=0
+ $Y2=0
cc_314 N_A_386_326#_c_257_n N_VGND_c_943_n 0.00241264f $X=2.495 $Y=0.42 $X2=0
+ $Y2=0
cc_315 N_A_386_326#_c_251_n N_VGND_c_945_n 0.0125682f $X=4.565 $Y=0.34 $X2=0
+ $Y2=0
cc_316 N_A_386_326#_c_253_n N_VGND_c_945_n 0.0244835f $X=6.895 $Y=0.665 $X2=0
+ $Y2=0
cc_317 N_A_386_326#_c_246_n N_A_239_85#_c_1004_n 0.00467906f $X=2.42 $Y=1.705
+ $X2=0 $Y2=0
cc_318 N_A_386_326#_M1010_g N_A_239_85#_c_1004_n 0.00381815f $X=2.495 $Y=0.955
+ $X2=0 $Y2=0
cc_319 N_A_386_326#_c_250_n N_A_239_85#_c_1004_n 0.00898486f $X=2.02 $Y=1.705
+ $X2=0 $Y2=0
cc_320 N_A_386_326#_M1010_g N_A_239_85#_c_1006_n 0.010286f $X=2.495 $Y=0.955
+ $X2=0 $Y2=0
cc_321 N_A_386_326#_M1010_g N_A_239_85#_c_1032_n 0.0138414f $X=2.495 $Y=0.955
+ $X2=0 $Y2=0
cc_322 N_A_386_326#_c_251_n N_A_239_85#_c_1032_n 0.00556984f $X=4.565 $Y=0.34
+ $X2=0 $Y2=0
cc_323 N_A_386_326#_c_255_n N_A_239_85#_c_1032_n 0.00924645f $X=2.34 $Y=0.34
+ $X2=0 $Y2=0
cc_324 N_A_386_326#_c_257_n N_A_239_85#_c_1032_n 4.02158e-19 $X=2.495 $Y=0.42
+ $X2=0 $Y2=0
cc_325 N_A_386_326#_c_255_n N_A_239_85#_c_1036_n 0.0135204f $X=2.34 $Y=0.34
+ $X2=0 $Y2=0
cc_326 N_A_386_326#_c_257_n N_A_239_85#_c_1036_n 0.00133759f $X=2.495 $Y=0.42
+ $X2=0 $Y2=0
cc_327 N_A_386_326#_c_251_n N_A_239_85#_c_1007_n 0.0690104f $X=4.565 $Y=0.34
+ $X2=0 $Y2=0
cc_328 N_A_386_326#_c_252_n N_A_239_85#_c_1007_n 4.28062e-19 $X=4.69 $Y=1.665
+ $X2=0 $Y2=0
cc_329 N_A_386_326#_c_305_p N_A_239_85#_c_1007_n 0.00520638f $X=4.69 $Y=0.665
+ $X2=0 $Y2=0
cc_330 N_A_386_326#_M1010_g N_A_239_85#_c_1009_n 0.00256415f $X=2.495 $Y=0.955
+ $X2=0 $Y2=0
cc_331 N_A_386_326#_c_251_n N_A_239_85#_c_1009_n 0.0125599f $X=4.565 $Y=0.34
+ $X2=0 $Y2=0
cc_332 N_A_562_123#_c_405_n N_A_685_59#_M1012_d 0.00434337f $X=6.01 $Y=2.325
+ $X2=0 $Y2=0
cc_333 N_A_562_123#_c_388_n N_A_685_59#_c_529_n 0.0121258f $X=3.03 $Y=1.885
+ $X2=0 $Y2=0
cc_334 N_A_562_123#_c_400_n N_A_685_59#_c_529_n 0.0096809f $X=3.59 $Y=1.8 $X2=0
+ $Y2=0
cc_335 N_A_562_123#_c_402_n N_A_685_59#_c_529_n 0.017338f $X=3.675 $Y=2.505
+ $X2=0 $Y2=0
cc_336 N_A_562_123#_c_388_n N_A_685_59#_c_530_n 0.0159914f $X=3.03 $Y=1.885
+ $X2=0 $Y2=0
cc_337 N_A_562_123#_c_402_n N_A_685_59#_c_530_n 0.00451529f $X=3.675 $Y=2.505
+ $X2=0 $Y2=0
cc_338 N_A_562_123#_c_431_p N_A_685_59#_c_530_n 0.00728303f $X=3.76 $Y=2.59
+ $X2=0 $Y2=0
cc_339 N_A_562_123#_M1003_g N_A_685_59#_c_521_n 0.0180485f $X=2.885 $Y=0.955
+ $X2=0 $Y2=0
cc_340 N_A_562_123#_c_400_n N_A_685_59#_c_522_n 0.00140172f $X=3.59 $Y=1.8 $X2=0
+ $Y2=0
cc_341 N_A_562_123#_c_388_n N_A_685_59#_c_523_n 0.00916653f $X=3.03 $Y=1.885
+ $X2=0 $Y2=0
cc_342 N_A_562_123#_c_400_n N_A_685_59#_c_523_n 0.00996571f $X=3.59 $Y=1.8 $X2=0
+ $Y2=0
cc_343 N_A_562_123#_c_392_n N_A_685_59#_c_523_n 0.00115804f $X=3.355 $Y=1.8
+ $X2=0 $Y2=0
cc_344 N_A_562_123#_M1003_g N_A_685_59#_c_524_n 7.46303e-19 $X=2.885 $Y=0.955
+ $X2=0 $Y2=0
cc_345 N_A_562_123#_c_400_n N_A_685_59#_c_524_n 0.0179102f $X=3.59 $Y=1.8 $X2=0
+ $Y2=0
cc_346 N_A_562_123#_c_392_n N_A_685_59#_c_524_n 0.00937071f $X=3.355 $Y=1.8
+ $X2=0 $Y2=0
cc_347 N_A_562_123#_M1003_g N_A_685_59#_c_525_n 0.00107053f $X=2.885 $Y=0.955
+ $X2=0 $Y2=0
cc_348 N_A_562_123#_c_388_n N_A_685_59#_c_525_n 0.0069901f $X=3.03 $Y=1.885
+ $X2=0 $Y2=0
cc_349 N_A_562_123#_c_392_n N_A_685_59#_c_525_n 0.00197703f $X=3.355 $Y=1.8
+ $X2=0 $Y2=0
cc_350 N_A_562_123#_c_400_n N_A_685_59#_c_526_n 0.0139236f $X=3.59 $Y=1.8 $X2=0
+ $Y2=0
cc_351 N_A_562_123#_c_392_n N_A_685_59#_c_526_n 0.00589522f $X=3.355 $Y=1.8
+ $X2=0 $Y2=0
cc_352 N_A_562_123#_c_402_n N_A_685_59#_c_526_n 0.021007f $X=3.675 $Y=2.505
+ $X2=0 $Y2=0
cc_353 N_A_562_123#_c_398_n N_A_685_59#_c_533_n 0.013139f $X=5.315 $Y=1.61 $X2=0
+ $Y2=0
cc_354 N_A_562_123#_c_403_n N_A_685_59#_c_533_n 0.0768671f $X=5.34 $Y=2.59 $X2=0
+ $Y2=0
cc_355 N_A_562_123#_c_405_n N_A_685_59#_c_533_n 0.0310555f $X=6.01 $Y=2.325
+ $X2=0 $Y2=0
cc_356 N_A_562_123#_c_402_n N_A_685_59#_c_534_n 0.0143568f $X=3.675 $Y=2.505
+ $X2=0 $Y2=0
cc_357 N_A_562_123#_c_403_n N_A_685_59#_c_534_n 0.014265f $X=5.34 $Y=2.59 $X2=0
+ $Y2=0
cc_358 N_A_562_123#_c_398_n N_A_685_59#_c_527_n 0.0111628f $X=5.315 $Y=1.61
+ $X2=0 $Y2=0
cc_359 N_A_562_123#_M1002_g N_A_685_59#_c_527_n 0.00698684f $X=5.455 $Y=0.78
+ $X2=0 $Y2=0
cc_360 N_A_562_123#_c_390_n N_A_685_59#_c_527_n 0.00761918f $X=5.845 $Y=1.425
+ $X2=0 $Y2=0
cc_361 N_A_562_123#_c_391_n N_A_685_59#_c_527_n 0.0117749f $X=5.53 $Y=1.425
+ $X2=0 $Y2=0
cc_362 N_A_562_123#_c_393_n N_A_685_59#_c_527_n 0.0383754f $X=6.01 $Y=1.515
+ $X2=0 $Y2=0
cc_363 N_A_562_123#_c_405_n N_A_685_59#_c_527_n 0.0151941f $X=6.01 $Y=2.325
+ $X2=0 $Y2=0
cc_364 N_A_562_123#_c_394_n N_A_685_59#_c_527_n 0.00798634f $X=6.01 $Y=1.35
+ $X2=0 $Y2=0
cc_365 N_A_562_123#_c_396_n N_A_685_59#_c_527_n 0.00147605f $X=6.01 $Y=1.425
+ $X2=0 $Y2=0
cc_366 N_A_562_123#_M1002_g N_A_685_59#_c_528_n 0.00792994f $X=5.455 $Y=0.78
+ $X2=0 $Y2=0
cc_367 N_A_562_123#_c_390_n N_A_685_59#_c_528_n 0.00793048f $X=5.845 $Y=1.425
+ $X2=0 $Y2=0
cc_368 N_A_562_123#_c_395_n N_A_685_59#_c_528_n 0.0217027f $X=6.235 $Y=1.005
+ $X2=0 $Y2=0
cc_369 N_A_562_123#_c_391_n N_A_592_149#_c_614_n 0.00570465f $X=5.53 $Y=1.425
+ $X2=0 $Y2=0
cc_370 N_A_562_123#_c_398_n N_A_592_149#_c_624_n 0.0247415f $X=5.315 $Y=1.61
+ $X2=0 $Y2=0
cc_371 N_A_562_123#_c_403_n N_A_592_149#_c_624_n 0.0144641f $X=5.34 $Y=2.59
+ $X2=0 $Y2=0
cc_372 N_A_562_123#_c_405_n N_A_592_149#_c_624_n 6.77567e-19 $X=6.01 $Y=2.325
+ $X2=0 $Y2=0
cc_373 N_A_562_123#_M1002_g N_A_592_149#_c_615_n 0.0263176f $X=5.455 $Y=0.78
+ $X2=0 $Y2=0
cc_374 N_A_562_123#_c_391_n N_A_592_149#_c_616_n 0.00126227f $X=5.53 $Y=1.425
+ $X2=0 $Y2=0
cc_375 N_A_562_123#_M1003_g N_A_592_149#_c_617_n 0.00569551f $X=2.885 $Y=0.955
+ $X2=0 $Y2=0
cc_376 N_A_562_123#_c_388_n N_A_592_149#_c_617_n 0.00383164f $X=3.03 $Y=1.885
+ $X2=0 $Y2=0
cc_377 N_A_562_123#_c_392_n N_A_592_149#_c_617_n 0.0305203f $X=3.355 $Y=1.8
+ $X2=0 $Y2=0
cc_378 N_A_562_123#_c_388_n N_A_592_149#_c_626_n 0.0133727f $X=3.03 $Y=1.885
+ $X2=0 $Y2=0
cc_379 N_A_562_123#_c_392_n N_A_592_149#_c_626_n 0.0124167f $X=3.355 $Y=1.8
+ $X2=0 $Y2=0
cc_380 N_A_562_123#_c_402_n N_A_592_149#_c_626_n 0.00325293f $X=3.675 $Y=2.505
+ $X2=0 $Y2=0
cc_381 N_A_562_123#_c_388_n N_A_592_149#_c_627_n 0.00449176f $X=3.03 $Y=1.885
+ $X2=0 $Y2=0
cc_382 N_A_562_123#_c_400_n N_A_592_149#_c_627_n 0.00479689f $X=3.59 $Y=1.8
+ $X2=0 $Y2=0
cc_383 N_A_562_123#_c_392_n N_A_592_149#_c_627_n 0.020349f $X=3.355 $Y=1.8 $X2=0
+ $Y2=0
cc_384 N_A_562_123#_c_402_n N_A_592_149#_c_627_n 0.0134146f $X=3.675 $Y=2.505
+ $X2=0 $Y2=0
cc_385 N_A_562_123#_c_400_n N_A_592_149#_c_618_n 0.0037683f $X=3.59 $Y=1.8 $X2=0
+ $Y2=0
cc_386 N_A_562_123#_M1003_g N_A_592_149#_c_619_n 0.011968f $X=2.885 $Y=0.955
+ $X2=0 $Y2=0
cc_387 N_A_562_123#_c_388_n N_A_592_149#_c_619_n 0.0016309f $X=3.03 $Y=1.885
+ $X2=0 $Y2=0
cc_388 N_A_562_123#_c_392_n N_A_592_149#_c_619_n 0.0397344f $X=3.355 $Y=1.8
+ $X2=0 $Y2=0
cc_389 N_A_562_123#_c_394_n N_GATE_M1014_g 0.00586999f $X=6.01 $Y=1.35 $X2=0
+ $Y2=0
cc_390 N_A_562_123#_c_395_n N_GATE_M1014_g 0.00548315f $X=6.235 $Y=1.005 $X2=0
+ $Y2=0
cc_391 N_A_562_123#_c_404_n N_GATE_c_719_n 0.00538385f $X=6.01 $Y=1.95 $X2=0
+ $Y2=0
cc_392 N_A_562_123#_c_393_n N_GATE_c_719_n 3.98767e-19 $X=6.01 $Y=1.515 $X2=0
+ $Y2=0
cc_393 N_A_562_123#_c_405_n N_GATE_c_719_n 0.0100851f $X=6.01 $Y=2.325 $X2=0
+ $Y2=0
cc_394 N_A_562_123#_c_396_n N_GATE_c_719_n 0.0212619f $X=6.01 $Y=1.425 $X2=0
+ $Y2=0
cc_395 N_A_562_123#_c_393_n N_GATE_c_720_n 0.0318395f $X=6.01 $Y=1.515 $X2=0
+ $Y2=0
cc_396 N_A_562_123#_c_405_n N_GATE_c_720_n 0.0114037f $X=6.01 $Y=2.325 $X2=0
+ $Y2=0
cc_397 N_A_562_123#_c_395_n N_GATE_c_720_n 0.00332637f $X=6.235 $Y=1.005 $X2=0
+ $Y2=0
cc_398 N_A_562_123#_c_396_n N_GATE_c_720_n 0.00197366f $X=6.01 $Y=1.425 $X2=0
+ $Y2=0
cc_399 N_A_562_123#_c_403_n N_VPWR_M1001_d 0.00821677f $X=5.34 $Y=2.59 $X2=0
+ $Y2=0
cc_400 N_A_562_123#_c_403_n N_VPWR_c_754_n 0.0252482f $X=5.34 $Y=2.59 $X2=0
+ $Y2=0
cc_401 N_A_562_123#_c_405_n N_VPWR_c_755_n 0.0534822f $X=6.01 $Y=2.325 $X2=0
+ $Y2=0
cc_402 N_A_562_123#_c_388_n N_VPWR_c_757_n 0.00444415f $X=3.03 $Y=1.885 $X2=0
+ $Y2=0
cc_403 N_A_562_123#_c_403_n N_VPWR_c_757_n 0.012541f $X=5.34 $Y=2.59 $X2=0 $Y2=0
cc_404 N_A_562_123#_c_398_n N_VPWR_c_758_n 5.65108e-19 $X=5.315 $Y=1.61 $X2=0
+ $Y2=0
cc_405 N_A_562_123#_c_403_n N_VPWR_c_758_n 0.00295476f $X=5.34 $Y=2.59 $X2=0
+ $Y2=0
cc_406 N_A_562_123#_c_405_n N_VPWR_c_758_n 0.0233045f $X=6.01 $Y=2.325 $X2=0
+ $Y2=0
cc_407 N_A_562_123#_c_388_n N_VPWR_c_751_n 0.00443106f $X=3.03 $Y=1.885 $X2=0
+ $Y2=0
cc_408 N_A_562_123#_c_403_n N_VPWR_c_751_n 0.0291491f $X=5.34 $Y=2.59 $X2=0
+ $Y2=0
cc_409 N_A_562_123#_c_405_n N_VPWR_c_751_n 0.0352734f $X=6.01 $Y=2.325 $X2=0
+ $Y2=0
cc_410 N_A_562_123#_c_388_n N_A_229_392#_c_819_n 0.00327191f $X=3.03 $Y=1.885
+ $X2=0 $Y2=0
cc_411 N_A_562_123#_c_388_n N_A_229_392#_c_822_n 0.00190162f $X=3.03 $Y=1.885
+ $X2=0 $Y2=0
cc_412 N_A_562_123#_c_403_n N_A_419_392#_M1005_d 0.00405842f $X=5.34 $Y=2.59
+ $X2=0 $Y2=0
cc_413 N_A_562_123#_c_431_p N_A_419_392#_M1005_d 6.7409e-19 $X=3.76 $Y=2.59
+ $X2=0 $Y2=0
cc_414 N_A_562_123#_c_388_n N_A_419_392#_c_859_n 0.00218148f $X=3.03 $Y=1.885
+ $X2=0 $Y2=0
cc_415 N_A_562_123#_c_388_n N_A_419_392#_c_877_n 0.0126481f $X=3.03 $Y=1.885
+ $X2=0 $Y2=0
cc_416 N_A_562_123#_c_402_n N_A_419_392#_c_877_n 0.0058422f $X=3.675 $Y=2.505
+ $X2=0 $Y2=0
cc_417 N_A_562_123#_c_431_p N_A_419_392#_c_877_n 0.00354594f $X=3.76 $Y=2.59
+ $X2=0 $Y2=0
cc_418 N_A_562_123#_c_431_p N_A_419_392#_c_880_n 0.00585258f $X=3.76 $Y=2.59
+ $X2=0 $Y2=0
cc_419 N_A_562_123#_c_388_n N_A_419_392#_c_862_n 0.0019436f $X=3.03 $Y=1.885
+ $X2=0 $Y2=0
cc_420 N_A_562_123#_c_403_n N_A_419_392#_c_863_n 0.0193689f $X=5.34 $Y=2.59
+ $X2=0 $Y2=0
cc_421 N_A_562_123#_c_431_p N_A_419_392#_c_863_n 0.00842254f $X=3.76 $Y=2.59
+ $X2=0 $Y2=0
cc_422 N_A_562_123#_c_388_n N_A_419_392#_c_864_n 0.00429406f $X=3.03 $Y=1.885
+ $X2=0 $Y2=0
cc_423 N_A_562_123#_M1002_g N_VGND_c_941_n 0.00414982f $X=5.455 $Y=0.78 $X2=0
+ $Y2=0
cc_424 N_A_562_123#_M1002_g N_VGND_c_943_n 0.00533081f $X=5.455 $Y=0.78 $X2=0
+ $Y2=0
cc_425 N_A_562_123#_M1002_g N_VGND_c_945_n 0.00378066f $X=5.455 $Y=0.78 $X2=0
+ $Y2=0
cc_426 N_A_562_123#_M1003_g N_A_239_85#_c_1007_n 0.00845704f $X=2.885 $Y=0.955
+ $X2=0 $Y2=0
cc_427 N_A_562_123#_M1003_g N_A_239_85#_c_1009_n 0.00706284f $X=2.885 $Y=0.955
+ $X2=0 $Y2=0
cc_428 N_A_685_59#_c_522_n N_A_592_149#_c_613_n 0.00934639f $X=3.64 $Y=1.39
+ $X2=0 $Y2=0
cc_429 N_A_685_59#_c_524_n N_A_592_149#_c_613_n 0.00510189f $X=3.93 $Y=1.41
+ $X2=0 $Y2=0
cc_430 N_A_685_59#_c_524_n N_A_592_149#_c_614_n 0.00105015f $X=3.93 $Y=1.41
+ $X2=0 $Y2=0
cc_431 N_A_685_59#_c_527_n N_A_592_149#_c_614_n 2.2559e-19 $X=5.54 $Y=1.83 $X2=0
+ $Y2=0
cc_432 N_A_685_59#_c_526_n N_A_592_149#_c_624_n 0.00471994f $X=4.015 $Y=2.165
+ $X2=0 $Y2=0
cc_433 N_A_685_59#_c_533_n N_A_592_149#_c_624_n 0.0133171f $X=5.375 $Y=2.25
+ $X2=0 $Y2=0
cc_434 N_A_685_59#_c_527_n N_A_592_149#_c_624_n 0.00111405f $X=5.54 $Y=1.83
+ $X2=0 $Y2=0
cc_435 N_A_685_59#_c_527_n N_A_592_149#_c_615_n 0.00147828f $X=5.54 $Y=1.83
+ $X2=0 $Y2=0
cc_436 N_A_685_59#_c_528_n N_A_592_149#_c_615_n 8.50659e-19 $X=5.67 $Y=1.005
+ $X2=0 $Y2=0
cc_437 N_A_685_59#_c_529_n N_A_592_149#_c_626_n 4.03212e-19 $X=3.565 $Y=2.375
+ $X2=0 $Y2=0
cc_438 N_A_685_59#_c_529_n N_A_592_149#_c_627_n 0.00156512f $X=3.565 $Y=2.375
+ $X2=0 $Y2=0
cc_439 N_A_685_59#_c_521_n N_A_592_149#_c_618_n 0.0129061f $X=3.64 $Y=1.24 $X2=0
+ $Y2=0
cc_440 N_A_685_59#_c_522_n N_A_592_149#_c_618_n 0.00723426f $X=3.64 $Y=1.39
+ $X2=0 $Y2=0
cc_441 N_A_685_59#_c_524_n N_A_592_149#_c_618_n 0.0389883f $X=3.93 $Y=1.41 $X2=0
+ $Y2=0
cc_442 N_A_685_59#_c_521_n N_A_592_149#_c_620_n 0.00532445f $X=3.64 $Y=1.24
+ $X2=0 $Y2=0
cc_443 N_A_685_59#_c_521_n N_A_592_149#_c_621_n 6.62218e-19 $X=3.64 $Y=1.24
+ $X2=0 $Y2=0
cc_444 N_A_685_59#_c_524_n N_A_592_149#_c_621_n 0.0027282f $X=3.93 $Y=1.41 $X2=0
+ $Y2=0
cc_445 N_A_685_59#_c_521_n N_A_592_149#_c_622_n 0.0111292f $X=3.64 $Y=1.24 $X2=0
+ $Y2=0
cc_446 N_A_685_59#_c_528_n N_GATE_M1014_g 3.79315e-19 $X=5.67 $Y=1.005 $X2=0
+ $Y2=0
cc_447 N_A_685_59#_c_533_n N_VPWR_M1001_d 0.0183998f $X=5.375 $Y=2.25 $X2=0
+ $Y2=0
cc_448 N_A_685_59#_c_530_n N_VPWR_c_757_n 0.00286838f $X=3.565 $Y=2.465 $X2=0
+ $Y2=0
cc_449 N_A_685_59#_c_530_n N_VPWR_c_751_n 0.00361977f $X=3.565 $Y=2.465 $X2=0
+ $Y2=0
cc_450 N_A_685_59#_c_530_n N_A_419_392#_c_877_n 0.00153124f $X=3.565 $Y=2.465
+ $X2=0 $Y2=0
cc_451 N_A_685_59#_c_530_n N_A_419_392#_c_880_n 0.00447905f $X=3.565 $Y=2.465
+ $X2=0 $Y2=0
cc_452 N_A_685_59#_c_530_n N_A_419_392#_c_863_n 0.0145454f $X=3.565 $Y=2.465
+ $X2=0 $Y2=0
cc_453 N_A_685_59#_c_521_n N_VGND_c_940_n 8.63546e-19 $X=3.64 $Y=1.24 $X2=0
+ $Y2=0
cc_454 N_A_685_59#_c_521_n N_A_239_85#_c_1007_n 0.00935421f $X=3.64 $Y=1.24
+ $X2=0 $Y2=0
cc_455 N_A_685_59#_c_521_n N_A_239_85#_c_1009_n 8.42574e-19 $X=3.64 $Y=1.24
+ $X2=0 $Y2=0
cc_456 N_A_592_149#_c_624_n N_VPWR_c_754_n 0.00372286f $X=4.695 $Y=1.61 $X2=0
+ $Y2=0
cc_457 N_A_592_149#_c_624_n N_VPWR_c_757_n 0.00364445f $X=4.695 $Y=1.61 $X2=0
+ $Y2=0
cc_458 N_A_592_149#_c_624_n N_VPWR_c_751_n 0.0049796f $X=4.695 $Y=1.61 $X2=0
+ $Y2=0
cc_459 N_A_592_149#_c_626_n N_A_229_392#_M1000_s 0.00624139f $X=3.015 $Y=2.14
+ $X2=0 $Y2=0
cc_460 N_A_592_149#_c_626_n N_A_419_392#_c_859_n 0.017373f $X=3.015 $Y=2.14
+ $X2=0 $Y2=0
cc_461 N_A_592_149#_M1000_d N_A_419_392#_c_877_n 0.00364382f $X=3.105 $Y=1.96
+ $X2=0 $Y2=0
cc_462 N_A_592_149#_c_626_n N_A_419_392#_c_877_n 0.0167142f $X=3.015 $Y=2.14
+ $X2=0 $Y2=0
cc_463 N_A_592_149#_c_627_n N_A_419_392#_c_877_n 0.0179831f $X=3.255 $Y=2.14
+ $X2=0 $Y2=0
cc_464 N_A_592_149#_M1000_d N_A_419_392#_c_880_n 0.00414139f $X=3.105 $Y=1.96
+ $X2=0 $Y2=0
cc_465 N_A_592_149#_M1000_d N_A_419_392#_c_862_n 9.42062e-19 $X=3.105 $Y=1.96
+ $X2=0 $Y2=0
cc_466 N_A_592_149#_M1000_d N_A_419_392#_c_863_n 0.00270409f $X=3.105 $Y=1.96
+ $X2=0 $Y2=0
cc_467 N_A_592_149#_c_624_n N_A_419_392#_c_863_n 0.00238819f $X=4.695 $Y=1.61
+ $X2=0 $Y2=0
cc_468 N_A_592_149#_c_627_n N_A_419_392#_c_863_n 0.00304765f $X=3.255 $Y=2.14
+ $X2=0 $Y2=0
cc_469 N_A_592_149#_c_626_n N_A_419_392#_c_864_n 0.0139565f $X=3.015 $Y=2.14
+ $X2=0 $Y2=0
cc_470 N_A_592_149#_c_615_n N_VGND_c_940_n 0.00360834f $X=4.865 $Y=1.225 $X2=0
+ $Y2=0
cc_471 N_A_592_149#_c_615_n N_VGND_c_943_n 0.00444234f $X=4.865 $Y=1.225 $X2=0
+ $Y2=0
cc_472 N_A_592_149#_c_615_n N_VGND_c_945_n 0.00124503f $X=4.865 $Y=1.225 $X2=0
+ $Y2=0
cc_473 N_A_592_149#_c_618_n N_A_239_85#_M1013_d 0.00571125f $X=4.065 $Y=1.02
+ $X2=0 $Y2=0
cc_474 N_A_592_149#_c_617_n N_A_239_85#_c_1004_n 0.0137144f $X=2.6 $Y=1.935
+ $X2=0 $Y2=0
cc_475 N_A_592_149#_c_617_n N_A_239_85#_c_1006_n 0.00636489f $X=2.6 $Y=1.935
+ $X2=0 $Y2=0
cc_476 N_A_592_149#_c_643_n N_A_239_85#_c_1006_n 0.0134926f $X=2.685 $Y=1.18
+ $X2=0 $Y2=0
cc_477 N_A_592_149#_c_643_n N_A_239_85#_c_1032_n 0.00809485f $X=2.685 $Y=1.18
+ $X2=0 $Y2=0
cc_478 N_A_592_149#_M1003_d N_A_239_85#_c_1007_n 0.00626188f $X=2.96 $Y=0.745
+ $X2=0 $Y2=0
cc_479 N_A_592_149#_c_619_n N_A_239_85#_c_1007_n 0.00458218f $X=3.015 $Y=1.1
+ $X2=0 $Y2=0
cc_480 N_A_592_149#_c_620_n N_A_239_85#_c_1007_n 0.0560276f $X=3.355 $Y=1.1
+ $X2=0 $Y2=0
cc_481 N_A_592_149#_c_643_n N_A_239_85#_c_1009_n 7.702e-19 $X=2.685 $Y=1.18
+ $X2=0 $Y2=0
cc_482 N_A_592_149#_c_619_n N_A_239_85#_c_1009_n 0.00762632f $X=3.015 $Y=1.1
+ $X2=0 $Y2=0
cc_483 N_A_592_149#_c_643_n A_514_149# 6.32083e-19 $X=2.685 $Y=1.18 $X2=-0.19
+ $Y2=-0.245
cc_484 N_A_592_149#_c_619_n A_514_149# 7.12223e-19 $X=3.015 $Y=1.1 $X2=-0.19
+ $Y2=-0.245
cc_485 N_GATE_c_719_n N_VPWR_c_755_n 0.0103676f $X=6.585 $Y=1.765 $X2=0 $Y2=0
cc_486 N_GATE_c_719_n N_VPWR_c_758_n 0.00393265f $X=6.585 $Y=1.765 $X2=0 $Y2=0
cc_487 N_GATE_c_719_n N_VPWR_c_751_n 0.00462577f $X=6.585 $Y=1.765 $X2=0 $Y2=0
cc_488 N_GATE_c_719_n Q 7.39082e-19 $X=6.585 $Y=1.765 $X2=0 $Y2=0
cc_489 N_GATE_M1014_g N_VGND_c_941_n 0.00836411f $X=6.46 $Y=0.78 $X2=0 $Y2=0
cc_490 N_GATE_M1014_g N_VGND_c_943_n 0.00533081f $X=6.46 $Y=0.78 $X2=0 $Y2=0
cc_491 N_VPWR_c_756_n N_A_229_392#_c_820_n 0.0145938f $X=1.66 $Y=3.33 $X2=0
+ $Y2=0
cc_492 N_VPWR_c_751_n N_A_229_392#_c_820_n 0.0120466f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_493 N_VPWR_c_761_n N_A_229_392#_c_820_n 0.00171364f $X=1.825 $Y=3.04 $X2=0
+ $Y2=0
cc_494 N_VPWR_M1011_d N_A_229_392#_c_821_n 0.0108714f $X=1.59 $Y=1.96 $X2=0
+ $Y2=0
cc_495 N_VPWR_c_756_n N_A_229_392#_c_821_n 0.00373946f $X=1.66 $Y=3.33 $X2=0
+ $Y2=0
cc_496 N_VPWR_c_757_n N_A_229_392#_c_821_n 0.00378997f $X=4.84 $Y=3.33 $X2=0
+ $Y2=0
cc_497 N_VPWR_c_751_n N_A_229_392#_c_821_n 0.0126785f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_498 N_VPWR_c_761_n N_A_229_392#_c_821_n 0.0247939f $X=1.825 $Y=3.04 $X2=0
+ $Y2=0
cc_499 N_VPWR_c_757_n N_A_229_392#_c_822_n 0.0341429f $X=4.84 $Y=3.33 $X2=0
+ $Y2=0
cc_500 N_VPWR_c_751_n N_A_229_392#_c_822_n 0.0288709f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_501 N_VPWR_c_761_n N_A_229_392#_c_822_n 0.00256814f $X=1.825 $Y=3.04 $X2=0
+ $Y2=0
cc_502 N_VPWR_c_751_n N_A_419_392#_c_877_n 0.00574011f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_503 N_VPWR_c_757_n N_A_419_392#_c_862_n 0.00876015f $X=4.84 $Y=3.33 $X2=0
+ $Y2=0
cc_504 N_VPWR_c_751_n N_A_419_392#_c_862_n 0.00638906f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_505 N_VPWR_c_757_n N_A_419_392#_c_863_n 0.0334884f $X=4.84 $Y=3.33 $X2=0
+ $Y2=0
cc_506 N_VPWR_c_751_n N_A_419_392#_c_863_n 0.0257212f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_507 N_VPWR_c_755_n Q 0.0400013f $X=6.895 $Y=2.115 $X2=0 $Y2=0
cc_508 N_VPWR_c_759_n Q 0.0161555f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_509 N_VPWR_c_751_n Q 0.0133393f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_510 N_A_229_392#_c_818_n N_A_419_392#_c_859_n 0.00833623f $X=1.29 $Y=2.105
+ $X2=0 $Y2=0
cc_511 N_A_229_392#_c_819_n N_A_419_392#_c_860_n 0.00907605f $X=2.805 $Y=2.82
+ $X2=0 $Y2=0
cc_512 N_A_229_392#_c_822_n N_A_419_392#_c_860_n 3.6241e-19 $X=2.335 $Y=2.8
+ $X2=0 $Y2=0
cc_513 N_A_229_392#_c_818_n N_A_419_392#_c_861_n 0.00442219f $X=1.29 $Y=2.105
+ $X2=0 $Y2=0
cc_514 N_A_229_392#_c_821_n N_A_419_392#_c_861_n 0.0212859f $X=2.165 $Y=2.8
+ $X2=0 $Y2=0
cc_515 N_A_229_392#_M1000_s N_A_419_392#_c_877_n 0.00651211f $X=2.66 $Y=1.96
+ $X2=0 $Y2=0
cc_516 N_A_229_392#_c_819_n N_A_419_392#_c_877_n 0.0171242f $X=2.805 $Y=2.82
+ $X2=0 $Y2=0
cc_517 N_A_229_392#_c_819_n N_A_419_392#_c_862_n 0.00695999f $X=2.805 $Y=2.82
+ $X2=0 $Y2=0
cc_518 N_A_229_392#_M1000_s N_A_419_392#_c_864_n 0.00247455f $X=2.66 $Y=1.96
+ $X2=0 $Y2=0
cc_519 N_A_229_392#_c_819_n N_A_419_392#_c_864_n 0.0131419f $X=2.805 $Y=2.82
+ $X2=0 $Y2=0
cc_520 N_A_229_392#_c_818_n N_A_239_85#_c_1005_n 0.00578551f $X=1.29 $Y=2.105
+ $X2=0 $Y2=0
cc_521 N_A_419_392#_c_859_n N_A_239_85#_c_1004_n 0.01161f $X=2.245 $Y=2.17 $X2=0
+ $Y2=0
cc_522 N_Q_c_914_n N_VGND_c_941_n 0.00156813f $X=7.4 $Y=0.555 $X2=0 $Y2=0
cc_523 N_Q_c_914_n N_VGND_c_942_n 0.0136906f $X=7.4 $Y=0.555 $X2=0 $Y2=0
cc_524 N_Q_c_914_n N_VGND_c_943_n 0.012877f $X=7.4 $Y=0.555 $X2=0 $Y2=0
cc_525 N_VGND_c_938_n N_A_239_85#_c_1002_n 0.0193118f $X=1.84 $Y=0.955 $X2=0
+ $Y2=0
cc_526 N_VGND_c_939_n N_A_239_85#_c_1002_n 0.0118717f $X=1.675 $Y=0 $X2=0 $Y2=0
cc_527 N_VGND_c_943_n N_A_239_85#_c_1002_n 0.0116501f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_528 N_VGND_c_938_n N_A_239_85#_c_1004_n 0.0277029f $X=1.84 $Y=0.955 $X2=0
+ $Y2=0
cc_529 N_VGND_M1017_d N_A_239_85#_c_1006_n 0.00637985f $X=1.675 $Y=0.425 $X2=0
+ $Y2=0
cc_530 N_VGND_c_938_n N_A_239_85#_c_1006_n 0.0198906f $X=1.84 $Y=0.955 $X2=0
+ $Y2=0
cc_531 N_VGND_M1017_d N_A_239_85#_c_1032_n 7.87578e-19 $X=1.675 $Y=0.425 $X2=0
+ $Y2=0
cc_532 N_VGND_c_943_n N_A_239_85#_c_1032_n 7.15647e-19 $X=7.44 $Y=0 $X2=0 $Y2=0
cc_533 N_VGND_M1017_d N_A_239_85#_c_1036_n 0.00365385f $X=1.675 $Y=0.425 $X2=0
+ $Y2=0
cc_534 N_VGND_c_938_n N_A_239_85#_c_1036_n 0.0141417f $X=1.84 $Y=0.955 $X2=0
+ $Y2=0
cc_535 N_VGND_c_943_n N_A_239_85#_c_1036_n 3.82042e-19 $X=7.44 $Y=0 $X2=0 $Y2=0
cc_536 N_VGND_c_938_n N_A_239_85#_c_1009_n 0.00480999f $X=1.84 $Y=0.955 $X2=0
+ $Y2=0
cc_537 N_A_239_85#_c_1032_n A_514_149# 0.00158593f $X=2.675 $Y=0.84 $X2=-0.19
+ $Y2=-0.245
cc_538 N_A_239_85#_c_1009_n A_514_149# 0.00139332f $X=2.76 $Y=0.68 $X2=-0.19
+ $Y2=-0.245
