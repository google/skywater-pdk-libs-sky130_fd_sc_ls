* File: sky130_fd_sc_ls__einvn_4.pxi.spice
* Created: Fri Aug 28 13:23:45 2020
* 
x_PM_SKY130_FD_SC_LS__EINVN_4%A_114_74# N_A_114_74#_M1013_d N_A_114_74#_M1006_d
+ N_A_114_74#_c_98_n N_A_114_74#_c_99_n N_A_114_74#_c_100_n N_A_114_74#_M1002_g
+ N_A_114_74#_c_101_n N_A_114_74#_c_102_n N_A_114_74#_M1003_g
+ N_A_114_74#_c_103_n N_A_114_74#_c_104_n N_A_114_74#_M1009_g
+ N_A_114_74#_c_105_n N_A_114_74#_c_106_n N_A_114_74#_M1016_g
+ N_A_114_74#_c_107_n N_A_114_74#_c_108_n N_A_114_74#_c_109_n
+ N_A_114_74#_c_110_n N_A_114_74#_c_111_n N_A_114_74#_c_112_n
+ PM_SKY130_FD_SC_LS__EINVN_4%A_114_74#
x_PM_SKY130_FD_SC_LS__EINVN_4%TE_B N_TE_B_M1013_g N_TE_B_c_187_n N_TE_B_M1006_g
+ N_TE_B_c_188_n N_TE_B_c_198_n N_TE_B_M1007_g N_TE_B_c_189_n N_TE_B_c_200_n
+ N_TE_B_M1011_g N_TE_B_c_190_n N_TE_B_c_202_n N_TE_B_M1012_g N_TE_B_c_191_n
+ N_TE_B_c_204_n N_TE_B_M1017_g N_TE_B_c_192_n N_TE_B_c_193_n N_TE_B_c_194_n
+ TE_B N_TE_B_c_195_n PM_SKY130_FD_SC_LS__EINVN_4%TE_B
x_PM_SKY130_FD_SC_LS__EINVN_4%A N_A_c_287_n N_A_M1001_g N_A_c_281_n N_A_M1000_g
+ N_A_c_288_n N_A_M1005_g N_A_c_282_n N_A_M1004_g N_A_c_289_n N_A_M1010_g
+ N_A_c_283_n N_A_M1008_g N_A_c_290_n N_A_M1014_g N_A_c_284_n N_A_M1015_g A A
+ N_A_c_286_n PM_SKY130_FD_SC_LS__EINVN_4%A
x_PM_SKY130_FD_SC_LS__EINVN_4%VPWR N_VPWR_M1006_s N_VPWR_M1007_s N_VPWR_M1012_s
+ N_VPWR_c_369_n N_VPWR_c_370_n N_VPWR_c_371_n N_VPWR_c_372_n VPWR
+ N_VPWR_c_373_n N_VPWR_c_374_n N_VPWR_c_375_n N_VPWR_c_368_n N_VPWR_c_377_n
+ N_VPWR_c_378_n PM_SKY130_FD_SC_LS__EINVN_4%VPWR
x_PM_SKY130_FD_SC_LS__EINVN_4%A_241_368# N_A_241_368#_M1007_d
+ N_A_241_368#_M1011_d N_A_241_368#_M1017_d N_A_241_368#_M1005_s
+ N_A_241_368#_M1014_s N_A_241_368#_c_434_n N_A_241_368#_c_430_n
+ N_A_241_368#_c_431_n N_A_241_368#_c_435_n N_A_241_368#_c_432_n
+ N_A_241_368#_c_436_n N_A_241_368#_c_437_n N_A_241_368#_c_438_n
+ N_A_241_368#_c_480_n N_A_241_368#_c_439_n N_A_241_368#_c_440_n
+ N_A_241_368#_c_433_n N_A_241_368#_c_441_n
+ PM_SKY130_FD_SC_LS__EINVN_4%A_241_368#
x_PM_SKY130_FD_SC_LS__EINVN_4%Z N_Z_M1000_s N_Z_M1008_s N_Z_M1001_d N_Z_M1010_d
+ N_Z_c_529_n N_Z_c_531_n N_Z_c_536_n N_Z_c_540_n N_Z_c_526_n N_Z_c_546_n Z
+ N_Z_c_527_n PM_SKY130_FD_SC_LS__EINVN_4%Z
x_PM_SKY130_FD_SC_LS__EINVN_4%VGND N_VGND_M1013_s N_VGND_M1002_s N_VGND_M1009_s
+ N_VGND_c_577_n N_VGND_c_578_n N_VGND_c_579_n N_VGND_c_580_n N_VGND_c_581_n
+ N_VGND_c_582_n N_VGND_c_583_n N_VGND_c_584_n VGND N_VGND_c_585_n
+ N_VGND_c_586_n PM_SKY130_FD_SC_LS__EINVN_4%VGND
x_PM_SKY130_FD_SC_LS__EINVN_4%A_281_74# N_A_281_74#_M1002_d N_A_281_74#_M1003_d
+ N_A_281_74#_M1016_d N_A_281_74#_M1004_d N_A_281_74#_M1015_d
+ N_A_281_74#_c_638_n N_A_281_74#_c_639_n N_A_281_74#_c_640_n
+ N_A_281_74#_c_641_n N_A_281_74#_c_642_n N_A_281_74#_c_643_n
+ N_A_281_74#_c_644_n N_A_281_74#_c_645_n N_A_281_74#_c_646_n
+ N_A_281_74#_c_647_n N_A_281_74#_c_670_n N_A_281_74#_c_648_n
+ PM_SKY130_FD_SC_LS__EINVN_4%A_281_74#
cc_1 VNB N_A_114_74#_c_98_n 0.0208628f $X=-0.19 $Y=-0.245 $X2=1.69 $Y2=1.26
cc_2 VNB N_A_114_74#_c_99_n 0.0139628f $X=-0.19 $Y=-0.245 $X2=1.295 $Y2=1.26
cc_3 VNB N_A_114_74#_c_100_n 0.0166447f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=1.185
cc_4 VNB N_A_114_74#_c_101_n 0.0122635f $X=-0.19 $Y=-0.245 $X2=2.12 $Y2=1.26
cc_5 VNB N_A_114_74#_c_102_n 0.0143129f $X=-0.19 $Y=-0.245 $X2=2.195 $Y2=1.185
cc_6 VNB N_A_114_74#_c_103_n 0.0122635f $X=-0.19 $Y=-0.245 $X2=2.55 $Y2=1.26
cc_7 VNB N_A_114_74#_c_104_n 0.0143129f $X=-0.19 $Y=-0.245 $X2=2.625 $Y2=1.185
cc_8 VNB N_A_114_74#_c_105_n 0.0200435f $X=-0.19 $Y=-0.245 $X2=2.98 $Y2=1.26
cc_9 VNB N_A_114_74#_c_106_n 0.0145547f $X=-0.19 $Y=-0.245 $X2=3.055 $Y2=1.185
cc_10 VNB N_A_114_74#_c_107_n 0.00511446f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=1.26
cc_11 VNB N_A_114_74#_c_108_n 0.00511435f $X=-0.19 $Y=-0.245 $X2=2.195 $Y2=1.26
cc_12 VNB N_A_114_74#_c_109_n 0.00511446f $X=-0.19 $Y=-0.245 $X2=2.625 $Y2=1.26
cc_13 VNB N_A_114_74#_c_110_n 0.0146868f $X=-0.19 $Y=-0.245 $X2=0.79 $Y2=1.31
cc_14 VNB N_A_114_74#_c_111_n 0.0066218f $X=-0.19 $Y=-0.245 $X2=0.79 $Y2=1.985
cc_15 VNB N_A_114_74#_c_112_n 0.0711714f $X=-0.19 $Y=-0.245 $X2=1.13 $Y2=0.465
cc_16 VNB N_TE_B_M1013_g 0.0294944f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_TE_B_c_187_n 0.0577213f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_TE_B_c_188_n 0.0235484f $X=-0.19 $Y=-0.245 $X2=1.295 $Y2=1.26
cc_19 VNB N_TE_B_c_189_n 0.00553319f $X=-0.19 $Y=-0.245 $X2=1.84 $Y2=1.26
cc_20 VNB N_TE_B_c_190_n 0.00547506f $X=-0.19 $Y=-0.245 $X2=2.27 $Y2=1.26
cc_21 VNB N_TE_B_c_191_n 0.0113445f $X=-0.19 $Y=-0.245 $X2=2.7 $Y2=1.26
cc_22 VNB N_TE_B_c_192_n 0.00370817f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=1.26
cc_23 VNB N_TE_B_c_193_n 0.0036966f $X=-0.19 $Y=-0.245 $X2=2.195 $Y2=1.26
cc_24 VNB N_TE_B_c_194_n 0.00370817f $X=-0.19 $Y=-0.245 $X2=2.625 $Y2=1.26
cc_25 VNB N_TE_B_c_195_n 0.00440334f $X=-0.19 $Y=-0.245 $X2=0.79 $Y2=2.815
cc_26 VNB N_A_c_281_n 0.0157318f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_c_282_n 0.0161778f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=0.74
cc_28 VNB N_A_c_283_n 0.0159974f $X=-0.19 $Y=-0.245 $X2=2.195 $Y2=0.74
cc_29 VNB N_A_c_284_n 0.0207336f $X=-0.19 $Y=-0.245 $X2=2.98 $Y2=1.26
cc_30 VNB A 0.0256668f $X=-0.19 $Y=-0.245 $X2=3.055 $Y2=0.74
cc_31 VNB N_A_c_286_n 0.122505f $X=-0.19 $Y=-0.245 $X2=1.13 $Y2=0.465
cc_32 VNB N_VPWR_c_368_n 0.223389f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_241_368#_c_430_n 0.00395162f $X=-0.19 $Y=-0.245 $X2=2.98 $Y2=1.26
cc_34 VNB N_A_241_368#_c_431_n 0.00301433f $X=-0.19 $Y=-0.245 $X2=2.7 $Y2=1.26
cc_35 VNB N_A_241_368#_c_432_n 0.00757f $X=-0.19 $Y=-0.245 $X2=2.625 $Y2=1.26
cc_36 VNB N_A_241_368#_c_433_n 0.00151865f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_Z_c_526_n 4.62656e-19 $X=-0.19 $Y=-0.245 $X2=0.79 $Y2=1.31
cc_38 VNB N_Z_c_527_n 0.00122353f $X=-0.19 $Y=-0.245 $X2=1.13 $Y2=1.145
cc_39 VNB N_VGND_c_577_n 0.010678f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=0.74
cc_40 VNB N_VGND_c_578_n 0.0420905f $X=-0.19 $Y=-0.245 $X2=2.12 $Y2=1.26
cc_41 VNB N_VGND_c_579_n 0.00323505f $X=-0.19 $Y=-0.245 $X2=2.195 $Y2=0.74
cc_42 VNB N_VGND_c_580_n 0.00323505f $X=-0.19 $Y=-0.245 $X2=2.625 $Y2=0.74
cc_43 VNB N_VGND_c_581_n 0.0381462f $X=-0.19 $Y=-0.245 $X2=2.7 $Y2=1.26
cc_44 VNB N_VGND_c_582_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=3.055 $Y2=1.185
cc_45 VNB N_VGND_c_583_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=3.055 $Y2=0.74
cc_46 VNB N_VGND_c_584_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=1.13 $Y2=1.185
cc_47 VNB N_VGND_c_585_n 0.0552148f $X=-0.19 $Y=-0.245 $X2=1.13 $Y2=1.145
cc_48 VNB N_VGND_c_586_n 0.305559f $X=-0.19 $Y=-0.245 $X2=1.13 $Y2=0.465
cc_49 VNB N_A_281_74#_c_638_n 0.00221876f $X=-0.19 $Y=-0.245 $X2=2.27 $Y2=1.26
cc_50 VNB N_A_281_74#_c_639_n 0.00627739f $X=-0.19 $Y=-0.245 $X2=2.625 $Y2=0.74
cc_51 VNB N_A_281_74#_c_640_n 2.75804e-19 $X=-0.19 $Y=-0.245 $X2=2.625 $Y2=0.74
cc_52 VNB N_A_281_74#_c_641_n 0.00229766f $X=-0.19 $Y=-0.245 $X2=3.055 $Y2=1.185
cc_53 VNB N_A_281_74#_c_642_n 0.0106645f $X=-0.19 $Y=-0.245 $X2=3.055 $Y2=0.74
cc_54 VNB N_A_281_74#_c_643_n 0.00251555f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=1.26
cc_55 VNB N_A_281_74#_c_644_n 2.66637e-19 $X=-0.19 $Y=-0.245 $X2=2.195 $Y2=1.26
cc_56 VNB N_A_281_74#_c_645_n 0.00304162f $X=-0.19 $Y=-0.245 $X2=2.625 $Y2=1.26
cc_57 VNB N_A_281_74#_c_646_n 0.01171f $X=-0.19 $Y=-0.245 $X2=0.79 $Y2=1.985
cc_58 VNB N_A_281_74#_c_647_n 0.0226357f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_281_74#_c_648_n 0.00105952f $X=-0.19 $Y=-0.245 $X2=1.13 $Y2=1.145
cc_60 VPB N_A_114_74#_c_111_n 0.0138015f $X=-0.19 $Y=1.66 $X2=0.79 $Y2=1.985
cc_61 VPB N_TE_B_c_187_n 0.0437465f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_TE_B_c_188_n 0.0346273f $X=-0.19 $Y=1.66 $X2=1.295 $Y2=1.26
cc_63 VPB N_TE_B_c_198_n 0.0184246f $X=-0.19 $Y=1.66 $X2=1.765 $Y2=0.74
cc_64 VPB N_TE_B_c_189_n 0.00889325f $X=-0.19 $Y=1.66 $X2=1.84 $Y2=1.26
cc_65 VPB N_TE_B_c_200_n 0.0152836f $X=-0.19 $Y=1.66 $X2=2.195 $Y2=0.74
cc_66 VPB N_TE_B_c_190_n 0.0104465f $X=-0.19 $Y=1.66 $X2=2.27 $Y2=1.26
cc_67 VPB N_TE_B_c_202_n 0.0153585f $X=-0.19 $Y=1.66 $X2=2.625 $Y2=0.74
cc_68 VPB N_TE_B_c_191_n 0.0148222f $X=-0.19 $Y=1.66 $X2=2.7 $Y2=1.26
cc_69 VPB N_TE_B_c_204_n 0.0152983f $X=-0.19 $Y=1.66 $X2=3.055 $Y2=0.74
cc_70 VPB N_TE_B_c_192_n 0.00460198f $X=-0.19 $Y=1.66 $X2=1.765 $Y2=1.26
cc_71 VPB N_TE_B_c_193_n 0.00435393f $X=-0.19 $Y=1.66 $X2=2.195 $Y2=1.26
cc_72 VPB N_TE_B_c_194_n 0.00448698f $X=-0.19 $Y=1.66 $X2=2.625 $Y2=1.26
cc_73 VPB N_TE_B_c_195_n 0.00780393f $X=-0.19 $Y=1.66 $X2=0.79 $Y2=2.815
cc_74 VPB N_A_c_287_n 0.0145656f $X=-0.19 $Y=1.66 $X2=0.57 $Y2=0.37
cc_75 VPB N_A_c_288_n 0.0141098f $X=-0.19 $Y=1.66 $X2=1.69 $Y2=1.26
cc_76 VPB N_A_c_289_n 0.0141098f $X=-0.19 $Y=1.66 $X2=1.84 $Y2=1.26
cc_77 VPB N_A_c_290_n 0.0181207f $X=-0.19 $Y=1.66 $X2=2.625 $Y2=1.185
cc_78 VPB N_A_c_286_n 0.0585457f $X=-0.19 $Y=1.66 $X2=1.13 $Y2=0.465
cc_79 VPB N_VPWR_c_369_n 0.012566f $X=-0.19 $Y=1.66 $X2=1.765 $Y2=0.74
cc_80 VPB N_VPWR_c_370_n 0.0495285f $X=-0.19 $Y=1.66 $X2=2.12 $Y2=1.26
cc_81 VPB N_VPWR_c_371_n 0.00655511f $X=-0.19 $Y=1.66 $X2=2.27 $Y2=1.26
cc_82 VPB N_VPWR_c_372_n 0.00756064f $X=-0.19 $Y=1.66 $X2=3.055 $Y2=1.185
cc_83 VPB N_VPWR_c_373_n 0.0337833f $X=-0.19 $Y=1.66 $X2=2.625 $Y2=1.26
cc_84 VPB N_VPWR_c_374_n 0.0185253f $X=-0.19 $Y=1.66 $X2=0.79 $Y2=2.815
cc_85 VPB N_VPWR_c_375_n 0.0583247f $X=-0.19 $Y=1.66 $X2=1.13 $Y2=0.465
cc_86 VPB N_VPWR_c_368_n 0.0867306f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_377_n 0.00460249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_378_n 0.00613757f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_A_241_368#_c_434_n 0.0143194f $X=-0.19 $Y=1.66 $X2=2.27 $Y2=1.26
cc_90 VPB N_A_241_368#_c_435_n 0.00319836f $X=-0.19 $Y=1.66 $X2=3.055 $Y2=0.74
cc_91 VPB N_A_241_368#_c_436_n 0.00133794f $X=-0.19 $Y=1.66 $X2=0.79 $Y2=2.815
cc_92 VPB N_A_241_368#_c_437_n 0.0030474f $X=-0.19 $Y=1.66 $X2=1.13 $Y2=0.465
cc_93 VPB N_A_241_368#_c_438_n 0.00170344f $X=-0.19 $Y=1.66 $X2=1.13 $Y2=0.465
cc_94 VPB N_A_241_368#_c_439_n 0.0124059f $X=-0.19 $Y=1.66 $X2=1.13 $Y2=1.145
cc_95 VPB N_A_241_368#_c_440_n 0.0425963f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB N_A_241_368#_c_441_n 0.00123754f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 N_A_114_74#_c_110_n N_TE_B_M1013_g 0.0183768f $X=0.79 $Y=1.31 $X2=0 $Y2=0
cc_98 N_A_114_74#_c_112_n N_TE_B_M1013_g 0.0180863f $X=1.13 $Y=0.465 $X2=0 $Y2=0
cc_99 N_A_114_74#_c_99_n N_TE_B_c_187_n 0.00138455f $X=1.295 $Y=1.26 $X2=0 $Y2=0
cc_100 N_A_114_74#_c_110_n N_TE_B_c_187_n 0.0037134f $X=0.79 $Y=1.31 $X2=0 $Y2=0
cc_101 N_A_114_74#_c_111_n N_TE_B_c_187_n 0.0351803f $X=0.79 $Y=1.985 $X2=0
+ $Y2=0
cc_102 N_A_114_74#_c_99_n N_TE_B_c_188_n 0.0163096f $X=1.295 $Y=1.26 $X2=0 $Y2=0
cc_103 N_A_114_74#_c_110_n N_TE_B_c_188_n 0.00181554f $X=0.79 $Y=1.31 $X2=0
+ $Y2=0
cc_104 N_A_114_74#_c_111_n N_TE_B_c_188_n 0.0210449f $X=0.79 $Y=1.985 $X2=0
+ $Y2=0
cc_105 N_A_114_74#_c_107_n N_TE_B_c_189_n 0.0163096f $X=1.765 $Y=1.26 $X2=0
+ $Y2=0
cc_106 N_A_114_74#_c_108_n N_TE_B_c_190_n 0.0163096f $X=2.195 $Y=1.26 $X2=0
+ $Y2=0
cc_107 N_A_114_74#_c_109_n N_TE_B_c_191_n 0.0163096f $X=2.625 $Y=1.26 $X2=0
+ $Y2=0
cc_108 N_A_114_74#_c_98_n N_TE_B_c_192_n 0.0163096f $X=1.69 $Y=1.26 $X2=0 $Y2=0
cc_109 N_A_114_74#_c_101_n N_TE_B_c_193_n 0.0163096f $X=2.12 $Y=1.26 $X2=0 $Y2=0
cc_110 N_A_114_74#_c_103_n N_TE_B_c_194_n 0.0163096f $X=2.55 $Y=1.26 $X2=0 $Y2=0
cc_111 N_A_114_74#_c_110_n N_TE_B_c_195_n 7.97299e-19 $X=0.79 $Y=1.31 $X2=0
+ $Y2=0
cc_112 N_A_114_74#_c_111_n N_TE_B_c_195_n 0.0354205f $X=0.79 $Y=1.985 $X2=0
+ $Y2=0
cc_113 N_A_114_74#_c_106_n N_A_c_281_n 0.00903267f $X=3.055 $Y=1.185 $X2=0 $Y2=0
cc_114 N_A_114_74#_c_105_n N_A_c_286_n 0.00903267f $X=2.98 $Y=1.26 $X2=0 $Y2=0
cc_115 N_A_114_74#_c_111_n N_VPWR_c_370_n 0.0690922f $X=0.79 $Y=1.985 $X2=0
+ $Y2=0
cc_116 N_A_114_74#_c_111_n N_VPWR_c_373_n 0.0145938f $X=0.79 $Y=1.985 $X2=0
+ $Y2=0
cc_117 N_A_114_74#_c_111_n N_VPWR_c_368_n 0.0120466f $X=0.79 $Y=1.985 $X2=0
+ $Y2=0
cc_118 N_A_114_74#_c_111_n N_A_241_368#_c_434_n 0.087169f $X=0.79 $Y=1.985 $X2=0
+ $Y2=0
cc_119 N_A_114_74#_c_98_n N_A_241_368#_c_430_n 0.00442459f $X=1.69 $Y=1.26 $X2=0
+ $Y2=0
cc_120 N_A_114_74#_c_99_n N_A_241_368#_c_431_n 0.0048544f $X=1.295 $Y=1.26 $X2=0
+ $Y2=0
cc_121 N_A_114_74#_c_110_n N_A_241_368#_c_431_n 0.00980665f $X=0.79 $Y=1.31
+ $X2=0 $Y2=0
cc_122 N_A_114_74#_c_111_n N_A_241_368#_c_431_n 0.0114923f $X=0.79 $Y=1.985
+ $X2=0 $Y2=0
cc_123 N_A_114_74#_c_103_n N_A_241_368#_c_432_n 0.00438974f $X=2.55 $Y=1.26
+ $X2=0 $Y2=0
cc_124 N_A_114_74#_c_105_n N_A_241_368#_c_432_n 0.00205135f $X=2.98 $Y=1.26
+ $X2=0 $Y2=0
cc_125 N_A_114_74#_c_101_n N_A_241_368#_c_433_n 0.00188621f $X=2.12 $Y=1.26
+ $X2=0 $Y2=0
cc_126 N_A_114_74#_c_110_n N_VGND_c_578_n 0.0367724f $X=0.79 $Y=1.31 $X2=0 $Y2=0
cc_127 N_A_114_74#_c_100_n N_VGND_c_579_n 0.0122703f $X=1.765 $Y=1.185 $X2=0
+ $Y2=0
cc_128 N_A_114_74#_c_101_n N_VGND_c_579_n 7.11061e-19 $X=2.12 $Y=1.26 $X2=0
+ $Y2=0
cc_129 N_A_114_74#_c_102_n N_VGND_c_579_n 0.0106722f $X=2.195 $Y=1.185 $X2=0
+ $Y2=0
cc_130 N_A_114_74#_c_104_n N_VGND_c_579_n 5.10431e-19 $X=2.625 $Y=1.185 $X2=0
+ $Y2=0
cc_131 N_A_114_74#_c_110_n N_VGND_c_579_n 0.00159476f $X=0.79 $Y=1.31 $X2=0
+ $Y2=0
cc_132 N_A_114_74#_c_102_n N_VGND_c_580_n 5.10431e-19 $X=2.195 $Y=1.185 $X2=0
+ $Y2=0
cc_133 N_A_114_74#_c_104_n N_VGND_c_580_n 0.0106722f $X=2.625 $Y=1.185 $X2=0
+ $Y2=0
cc_134 N_A_114_74#_c_105_n N_VGND_c_580_n 7.11061e-19 $X=2.98 $Y=1.26 $X2=0
+ $Y2=0
cc_135 N_A_114_74#_c_106_n N_VGND_c_580_n 0.010039f $X=3.055 $Y=1.185 $X2=0
+ $Y2=0
cc_136 N_A_114_74#_c_100_n N_VGND_c_581_n 0.00383152f $X=1.765 $Y=1.185 $X2=0
+ $Y2=0
cc_137 N_A_114_74#_c_110_n N_VGND_c_581_n 0.0406574f $X=0.79 $Y=1.31 $X2=0 $Y2=0
cc_138 N_A_114_74#_c_112_n N_VGND_c_581_n 0.00199209f $X=1.13 $Y=0.465 $X2=0
+ $Y2=0
cc_139 N_A_114_74#_c_102_n N_VGND_c_583_n 0.00383152f $X=2.195 $Y=1.185 $X2=0
+ $Y2=0
cc_140 N_A_114_74#_c_104_n N_VGND_c_583_n 0.00383152f $X=2.625 $Y=1.185 $X2=0
+ $Y2=0
cc_141 N_A_114_74#_c_106_n N_VGND_c_585_n 0.00383152f $X=3.055 $Y=1.185 $X2=0
+ $Y2=0
cc_142 N_A_114_74#_c_100_n N_VGND_c_586_n 0.00762539f $X=1.765 $Y=1.185 $X2=0
+ $Y2=0
cc_143 N_A_114_74#_c_102_n N_VGND_c_586_n 0.0075754f $X=2.195 $Y=1.185 $X2=0
+ $Y2=0
cc_144 N_A_114_74#_c_104_n N_VGND_c_586_n 0.0075754f $X=2.625 $Y=1.185 $X2=0
+ $Y2=0
cc_145 N_A_114_74#_c_106_n N_VGND_c_586_n 0.00757637f $X=3.055 $Y=1.185 $X2=0
+ $Y2=0
cc_146 N_A_114_74#_c_110_n N_VGND_c_586_n 0.0281533f $X=0.79 $Y=1.31 $X2=0 $Y2=0
cc_147 N_A_114_74#_c_100_n N_A_281_74#_c_638_n 0.00122824f $X=1.765 $Y=1.185
+ $X2=0 $Y2=0
cc_148 N_A_114_74#_c_110_n N_A_281_74#_c_638_n 0.0621205f $X=0.79 $Y=1.31 $X2=0
+ $Y2=0
cc_149 N_A_114_74#_c_112_n N_A_281_74#_c_638_n 0.00274841f $X=1.13 $Y=0.465
+ $X2=0 $Y2=0
cc_150 N_A_114_74#_c_98_n N_A_281_74#_c_639_n 8.87202e-19 $X=1.69 $Y=1.26 $X2=0
+ $Y2=0
cc_151 N_A_114_74#_c_100_n N_A_281_74#_c_639_n 0.0075146f $X=1.765 $Y=1.185
+ $X2=0 $Y2=0
cc_152 N_A_114_74#_c_101_n N_A_281_74#_c_639_n 0.00614039f $X=2.12 $Y=1.26 $X2=0
+ $Y2=0
cc_153 N_A_114_74#_c_102_n N_A_281_74#_c_639_n 0.00752307f $X=2.195 $Y=1.185
+ $X2=0 $Y2=0
cc_154 N_A_114_74#_c_103_n N_A_281_74#_c_639_n 8.86022e-19 $X=2.55 $Y=1.26 $X2=0
+ $Y2=0
cc_155 N_A_114_74#_c_107_n N_A_281_74#_c_639_n 0.00251095f $X=1.765 $Y=1.26
+ $X2=0 $Y2=0
cc_156 N_A_114_74#_c_108_n N_A_281_74#_c_639_n 0.00250761f $X=2.195 $Y=1.26
+ $X2=0 $Y2=0
cc_157 N_A_114_74#_c_98_n N_A_281_74#_c_640_n 0.00791143f $X=1.69 $Y=1.26 $X2=0
+ $Y2=0
cc_158 N_A_114_74#_c_110_n N_A_281_74#_c_640_n 0.0145349f $X=0.79 $Y=1.31 $X2=0
+ $Y2=0
cc_159 N_A_114_74#_c_102_n N_A_281_74#_c_641_n 0.00106896f $X=2.195 $Y=1.185
+ $X2=0 $Y2=0
cc_160 N_A_114_74#_c_104_n N_A_281_74#_c_641_n 0.00106896f $X=2.625 $Y=1.185
+ $X2=0 $Y2=0
cc_161 N_A_114_74#_c_103_n N_A_281_74#_c_642_n 8.87202e-19 $X=2.55 $Y=1.26 $X2=0
+ $Y2=0
cc_162 N_A_114_74#_c_104_n N_A_281_74#_c_642_n 0.00753499f $X=2.625 $Y=1.185
+ $X2=0 $Y2=0
cc_163 N_A_114_74#_c_105_n N_A_281_74#_c_642_n 0.0101675f $X=2.98 $Y=1.26 $X2=0
+ $Y2=0
cc_164 N_A_114_74#_c_106_n N_A_281_74#_c_642_n 0.00752307f $X=3.055 $Y=1.185
+ $X2=0 $Y2=0
cc_165 N_A_114_74#_c_109_n N_A_281_74#_c_642_n 0.00251095f $X=2.625 $Y=1.26
+ $X2=0 $Y2=0
cc_166 N_A_114_74#_c_106_n N_A_281_74#_c_643_n 9.48753e-19 $X=3.055 $Y=1.185
+ $X2=0 $Y2=0
cc_167 N_A_114_74#_c_106_n N_A_281_74#_c_644_n 9.80302e-19 $X=3.055 $Y=1.185
+ $X2=0 $Y2=0
cc_168 N_A_114_74#_c_103_n N_A_281_74#_c_670_n 0.00526155f $X=2.55 $Y=1.26 $X2=0
+ $Y2=0
cc_169 N_TE_B_c_204_n N_A_c_287_n 0.00992225f $X=2.975 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_170 N_TE_B_c_191_n N_A_c_286_n 0.00879305f $X=2.885 $Y=1.65 $X2=0 $Y2=0
cc_171 N_TE_B_c_187_n N_VPWR_c_370_n 0.0100063f $X=0.565 $Y=1.765 $X2=0 $Y2=0
cc_172 N_TE_B_c_195_n N_VPWR_c_370_n 0.0222388f $X=0.29 $Y=1.465 $X2=0 $Y2=0
cc_173 N_TE_B_c_198_n N_VPWR_c_371_n 0.0193133f $X=1.575 $Y=1.765 $X2=0 $Y2=0
cc_174 N_TE_B_c_189_n N_VPWR_c_371_n 0.00477816f $X=1.935 $Y=1.65 $X2=0 $Y2=0
cc_175 N_TE_B_c_200_n N_VPWR_c_371_n 0.00588051f $X=2.025 $Y=1.765 $X2=0 $Y2=0
cc_176 N_TE_B_c_192_n N_VPWR_c_371_n 3.61478e-19 $X=1.575 $Y=1.67 $X2=0 $Y2=0
cc_177 N_TE_B_c_200_n N_VPWR_c_372_n 7.29261e-19 $X=2.025 $Y=1.765 $X2=0 $Y2=0
cc_178 N_TE_B_c_202_n N_VPWR_c_372_n 0.016713f $X=2.475 $Y=1.765 $X2=0 $Y2=0
cc_179 N_TE_B_c_191_n N_VPWR_c_372_n 0.00653031f $X=2.885 $Y=1.65 $X2=0 $Y2=0
cc_180 N_TE_B_c_204_n N_VPWR_c_372_n 0.00752981f $X=2.975 $Y=1.765 $X2=0 $Y2=0
cc_181 N_TE_B_c_194_n N_VPWR_c_372_n 3.61478e-19 $X=2.475 $Y=1.67 $X2=0 $Y2=0
cc_182 N_TE_B_c_187_n N_VPWR_c_373_n 0.00445602f $X=0.565 $Y=1.765 $X2=0 $Y2=0
cc_183 N_TE_B_c_198_n N_VPWR_c_373_n 0.00413917f $X=1.575 $Y=1.765 $X2=0 $Y2=0
cc_184 N_TE_B_c_200_n N_VPWR_c_374_n 0.00445602f $X=2.025 $Y=1.765 $X2=0 $Y2=0
cc_185 N_TE_B_c_202_n N_VPWR_c_374_n 0.00413917f $X=2.475 $Y=1.765 $X2=0 $Y2=0
cc_186 N_TE_B_c_204_n N_VPWR_c_375_n 0.0044313f $X=2.975 $Y=1.765 $X2=0 $Y2=0
cc_187 N_TE_B_c_187_n N_VPWR_c_368_n 0.00866068f $X=0.565 $Y=1.765 $X2=0 $Y2=0
cc_188 N_TE_B_c_198_n N_VPWR_c_368_n 0.00822528f $X=1.575 $Y=1.765 $X2=0 $Y2=0
cc_189 N_TE_B_c_200_n N_VPWR_c_368_n 0.00857589f $X=2.025 $Y=1.765 $X2=0 $Y2=0
cc_190 N_TE_B_c_202_n N_VPWR_c_368_n 0.00817726f $X=2.475 $Y=1.765 $X2=0 $Y2=0
cc_191 N_TE_B_c_204_n N_VPWR_c_368_n 0.00853234f $X=2.975 $Y=1.765 $X2=0 $Y2=0
cc_192 N_TE_B_c_187_n N_A_241_368#_c_434_n 0.00240926f $X=0.565 $Y=1.765 $X2=0
+ $Y2=0
cc_193 N_TE_B_c_188_n N_A_241_368#_c_434_n 0.0109801f $X=1.485 $Y=1.65 $X2=0
+ $Y2=0
cc_194 N_TE_B_c_198_n N_A_241_368#_c_434_n 0.0072359f $X=1.575 $Y=1.765 $X2=0
+ $Y2=0
cc_195 N_TE_B_c_192_n N_A_241_368#_c_434_n 0.00118386f $X=1.575 $Y=1.67 $X2=0
+ $Y2=0
cc_196 N_TE_B_c_188_n N_A_241_368#_c_430_n 0.00237072f $X=1.485 $Y=1.65 $X2=0
+ $Y2=0
cc_197 N_TE_B_c_189_n N_A_241_368#_c_430_n 0.00661792f $X=1.935 $Y=1.65 $X2=0
+ $Y2=0
cc_198 N_TE_B_c_192_n N_A_241_368#_c_430_n 0.00904558f $X=1.575 $Y=1.67 $X2=0
+ $Y2=0
cc_199 N_TE_B_c_193_n N_A_241_368#_c_430_n 0.00827334f $X=2.025 $Y=1.67 $X2=0
+ $Y2=0
cc_200 N_TE_B_c_187_n N_A_241_368#_c_431_n 4.01997e-19 $X=0.565 $Y=1.765 $X2=0
+ $Y2=0
cc_201 N_TE_B_c_188_n N_A_241_368#_c_431_n 0.00428963f $X=1.485 $Y=1.65 $X2=0
+ $Y2=0
cc_202 N_TE_B_c_198_n N_A_241_368#_c_435_n 5.59846e-19 $X=1.575 $Y=1.765 $X2=0
+ $Y2=0
cc_203 N_TE_B_c_200_n N_A_241_368#_c_435_n 0.0143126f $X=2.025 $Y=1.765 $X2=0
+ $Y2=0
cc_204 N_TE_B_c_190_n N_A_241_368#_c_435_n 0.0101931f $X=2.385 $Y=1.65 $X2=0
+ $Y2=0
cc_205 N_TE_B_c_202_n N_A_241_368#_c_435_n 0.00579845f $X=2.475 $Y=1.765 $X2=0
+ $Y2=0
cc_206 N_TE_B_c_193_n N_A_241_368#_c_435_n 0.00379988f $X=2.025 $Y=1.67 $X2=0
+ $Y2=0
cc_207 N_TE_B_c_194_n N_A_241_368#_c_435_n 0.00103579f $X=2.475 $Y=1.67 $X2=0
+ $Y2=0
cc_208 N_TE_B_c_190_n N_A_241_368#_c_432_n 0.00237072f $X=2.385 $Y=1.65 $X2=0
+ $Y2=0
cc_209 N_TE_B_c_191_n N_A_241_368#_c_432_n 0.0159486f $X=2.885 $Y=1.65 $X2=0
+ $Y2=0
cc_210 N_TE_B_c_194_n N_A_241_368#_c_432_n 0.00904558f $X=2.475 $Y=1.67 $X2=0
+ $Y2=0
cc_211 N_TE_B_c_202_n N_A_241_368#_c_436_n 5.34422e-19 $X=2.475 $Y=1.765 $X2=0
+ $Y2=0
cc_212 N_TE_B_c_191_n N_A_241_368#_c_436_n 0.00575686f $X=2.885 $Y=1.65 $X2=0
+ $Y2=0
cc_213 N_TE_B_c_204_n N_A_241_368#_c_436_n 0.0125105f $X=2.975 $Y=1.765 $X2=0
+ $Y2=0
cc_214 N_TE_B_c_204_n N_A_241_368#_c_438_n 0.00311631f $X=2.975 $Y=1.765 $X2=0
+ $Y2=0
cc_215 N_TE_B_c_190_n N_A_241_368#_c_433_n 0.00261868f $X=2.385 $Y=1.65 $X2=0
+ $Y2=0
cc_216 N_TE_B_c_193_n N_A_241_368#_c_433_n 3.61456e-19 $X=2.025 $Y=1.67 $X2=0
+ $Y2=0
cc_217 N_TE_B_c_204_n Z 3.49656e-19 $X=2.975 $Y=1.765 $X2=0 $Y2=0
cc_218 N_TE_B_M1013_g N_VGND_c_578_n 0.00555851f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_219 N_TE_B_c_187_n N_VGND_c_578_n 0.00187637f $X=0.565 $Y=1.765 $X2=0 $Y2=0
cc_220 N_TE_B_c_195_n N_VGND_c_578_n 0.0206988f $X=0.29 $Y=1.465 $X2=0 $Y2=0
cc_221 N_TE_B_M1013_g N_VGND_c_581_n 0.00431986f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_222 N_TE_B_M1013_g N_VGND_c_586_n 0.00824594f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_223 N_TE_B_c_192_n N_A_281_74#_c_639_n 7.07907e-19 $X=1.575 $Y=1.67 $X2=0
+ $Y2=0
cc_224 N_TE_B_c_194_n N_A_281_74#_c_642_n 5.84787e-19 $X=2.475 $Y=1.67 $X2=0
+ $Y2=0
cc_225 N_A_c_287_n N_VPWR_c_375_n 0.00278271f $X=3.425 $Y=1.765 $X2=0 $Y2=0
cc_226 N_A_c_288_n N_VPWR_c_375_n 0.00278271f $X=3.875 $Y=1.765 $X2=0 $Y2=0
cc_227 N_A_c_289_n N_VPWR_c_375_n 0.00278271f $X=4.325 $Y=1.765 $X2=0 $Y2=0
cc_228 N_A_c_290_n N_VPWR_c_375_n 0.00278271f $X=4.775 $Y=1.765 $X2=0 $Y2=0
cc_229 N_A_c_287_n N_VPWR_c_368_n 0.00353907f $X=3.425 $Y=1.765 $X2=0 $Y2=0
cc_230 N_A_c_288_n N_VPWR_c_368_n 0.00353823f $X=3.875 $Y=1.765 $X2=0 $Y2=0
cc_231 N_A_c_289_n N_VPWR_c_368_n 0.00353823f $X=4.325 $Y=1.765 $X2=0 $Y2=0
cc_232 N_A_c_290_n N_VPWR_c_368_n 0.00357317f $X=4.775 $Y=1.765 $X2=0 $Y2=0
cc_233 N_A_c_286_n N_A_241_368#_c_432_n 0.00371655f $X=4.785 $Y=1.492 $X2=0
+ $Y2=0
cc_234 N_A_c_287_n N_A_241_368#_c_436_n 0.0074781f $X=3.425 $Y=1.765 $X2=0 $Y2=0
cc_235 N_A_c_286_n N_A_241_368#_c_436_n 0.00101907f $X=4.785 $Y=1.492 $X2=0
+ $Y2=0
cc_236 N_A_c_287_n N_A_241_368#_c_437_n 0.0128006f $X=3.425 $Y=1.765 $X2=0 $Y2=0
cc_237 N_A_c_288_n N_A_241_368#_c_437_n 0.0127857f $X=3.875 $Y=1.765 $X2=0 $Y2=0
cc_238 N_A_c_288_n N_A_241_368#_c_480_n 0.0062909f $X=3.875 $Y=1.765 $X2=0 $Y2=0
cc_239 N_A_c_289_n N_A_241_368#_c_480_n 0.0062909f $X=4.325 $Y=1.765 $X2=0 $Y2=0
cc_240 N_A_c_286_n N_A_241_368#_c_480_n 8.93776e-19 $X=4.785 $Y=1.492 $X2=0
+ $Y2=0
cc_241 N_A_c_289_n N_A_241_368#_c_439_n 0.0128349f $X=4.325 $Y=1.765 $X2=0 $Y2=0
cc_242 N_A_c_290_n N_A_241_368#_c_439_n 0.0136604f $X=4.775 $Y=1.765 $X2=0 $Y2=0
cc_243 N_A_c_290_n N_A_241_368#_c_440_n 0.00807045f $X=4.775 $Y=1.765 $X2=0
+ $Y2=0
cc_244 A N_A_241_368#_c_440_n 0.0148634f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_245 N_A_c_286_n N_A_241_368#_c_440_n 0.00381921f $X=4.785 $Y=1.492 $X2=0
+ $Y2=0
cc_246 N_A_c_287_n N_Z_c_529_n 0.00875043f $X=3.425 $Y=1.765 $X2=0 $Y2=0
cc_247 N_A_c_288_n N_Z_c_529_n 0.00999614f $X=3.875 $Y=1.765 $X2=0 $Y2=0
cc_248 N_A_c_288_n N_Z_c_531_n 0.00980715f $X=3.875 $Y=1.765 $X2=0 $Y2=0
cc_249 N_A_c_289_n N_Z_c_531_n 0.0101302f $X=4.325 $Y=1.765 $X2=0 $Y2=0
cc_250 N_A_c_290_n N_Z_c_531_n 0.00418463f $X=4.775 $Y=1.765 $X2=0 $Y2=0
cc_251 A N_Z_c_531_n 0.0517544f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_252 N_A_c_286_n N_Z_c_531_n 0.0370793f $X=4.785 $Y=1.492 $X2=0 $Y2=0
cc_253 N_A_c_282_n N_Z_c_536_n 0.013849f $X=3.915 $Y=1.22 $X2=0 $Y2=0
cc_254 N_A_c_283_n N_Z_c_536_n 0.0112736f $X=4.355 $Y=1.22 $X2=0 $Y2=0
cc_255 A N_Z_c_536_n 0.030527f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_256 N_A_c_286_n N_Z_c_536_n 7.08101e-19 $X=4.785 $Y=1.492 $X2=0 $Y2=0
cc_257 N_A_c_288_n N_Z_c_540_n 6.41034e-19 $X=3.875 $Y=1.765 $X2=0 $Y2=0
cc_258 N_A_c_289_n N_Z_c_540_n 0.00999614f $X=4.325 $Y=1.765 $X2=0 $Y2=0
cc_259 N_A_c_290_n N_Z_c_540_n 0.00925235f $X=4.775 $Y=1.765 $X2=0 $Y2=0
cc_260 N_A_c_281_n N_Z_c_526_n 7.88797e-19 $X=3.485 $Y=1.22 $X2=0 $Y2=0
cc_261 N_A_c_282_n N_Z_c_526_n 0.0045177f $X=3.915 $Y=1.22 $X2=0 $Y2=0
cc_262 N_A_c_283_n N_Z_c_526_n 6.97036e-19 $X=4.355 $Y=1.22 $X2=0 $Y2=0
cc_263 A N_Z_c_546_n 0.0140706f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_264 N_A_c_286_n N_Z_c_546_n 6.73793e-19 $X=4.785 $Y=1.492 $X2=0 $Y2=0
cc_265 N_A_c_287_n Z 0.00218937f $X=3.425 $Y=1.765 $X2=0 $Y2=0
cc_266 N_A_c_288_n Z 0.00145587f $X=3.875 $Y=1.765 $X2=0 $Y2=0
cc_267 N_A_c_289_n Z 7.00941e-19 $X=4.325 $Y=1.765 $X2=0 $Y2=0
cc_268 N_A_c_286_n Z 0.031018f $X=4.785 $Y=1.492 $X2=0 $Y2=0
cc_269 N_A_c_282_n N_Z_c_527_n 0.00160429f $X=3.915 $Y=1.22 $X2=0 $Y2=0
cc_270 A N_Z_c_527_n 0.023376f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_271 N_A_c_286_n N_Z_c_527_n 0.0219011f $X=4.785 $Y=1.492 $X2=0 $Y2=0
cc_272 N_A_c_281_n N_VGND_c_580_n 3.79623e-19 $X=3.485 $Y=1.22 $X2=0 $Y2=0
cc_273 N_A_c_281_n N_VGND_c_585_n 0.00278247f $X=3.485 $Y=1.22 $X2=0 $Y2=0
cc_274 N_A_c_282_n N_VGND_c_585_n 0.00278271f $X=3.915 $Y=1.22 $X2=0 $Y2=0
cc_275 N_A_c_283_n N_VGND_c_585_n 0.00278271f $X=4.355 $Y=1.22 $X2=0 $Y2=0
cc_276 N_A_c_284_n N_VGND_c_585_n 0.00278247f $X=4.785 $Y=1.22 $X2=0 $Y2=0
cc_277 N_A_c_281_n N_VGND_c_586_n 0.00353524f $X=3.485 $Y=1.22 $X2=0 $Y2=0
cc_278 N_A_c_282_n N_VGND_c_586_n 0.00352619f $X=3.915 $Y=1.22 $X2=0 $Y2=0
cc_279 N_A_c_283_n N_VGND_c_586_n 0.00353528f $X=4.355 $Y=1.22 $X2=0 $Y2=0
cc_280 N_A_c_284_n N_VGND_c_586_n 0.00357084f $X=4.785 $Y=1.22 $X2=0 $Y2=0
cc_281 N_A_c_281_n N_A_281_74#_c_642_n 0.00174914f $X=3.485 $Y=1.22 $X2=0 $Y2=0
cc_282 N_A_c_286_n N_A_281_74#_c_642_n 0.00712155f $X=4.785 $Y=1.492 $X2=0 $Y2=0
cc_283 N_A_c_281_n N_A_281_74#_c_643_n 0.00194824f $X=3.485 $Y=1.22 $X2=0 $Y2=0
cc_284 N_A_c_281_n N_A_281_74#_c_644_n 0.00761102f $X=3.485 $Y=1.22 $X2=0 $Y2=0
cc_285 N_A_c_282_n N_A_281_74#_c_644_n 9.14331e-19 $X=3.915 $Y=1.22 $X2=0 $Y2=0
cc_286 N_A_c_281_n N_A_281_74#_c_645_n 0.0146721f $X=3.485 $Y=1.22 $X2=0 $Y2=0
cc_287 N_A_c_282_n N_A_281_74#_c_645_n 0.0130518f $X=3.915 $Y=1.22 $X2=0 $Y2=0
cc_288 N_A_c_286_n N_A_281_74#_c_645_n 2.98942e-19 $X=4.785 $Y=1.492 $X2=0 $Y2=0
cc_289 N_A_c_283_n N_A_281_74#_c_646_n 0.00708406f $X=4.355 $Y=1.22 $X2=0 $Y2=0
cc_290 N_A_c_284_n N_A_281_74#_c_646_n 0.0140292f $X=4.785 $Y=1.22 $X2=0 $Y2=0
cc_291 N_A_c_283_n N_A_281_74#_c_647_n 5.5198e-19 $X=4.355 $Y=1.22 $X2=0 $Y2=0
cc_292 N_A_c_284_n N_A_281_74#_c_647_n 0.0114766f $X=4.785 $Y=1.22 $X2=0 $Y2=0
cc_293 A N_A_281_74#_c_647_n 0.0251801f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_294 N_A_c_286_n N_A_281_74#_c_647_n 0.00114751f $X=4.785 $Y=1.492 $X2=0 $Y2=0
cc_295 N_A_c_283_n N_A_281_74#_c_648_n 0.00529157f $X=4.355 $Y=1.22 $X2=0 $Y2=0
cc_296 N_A_c_284_n N_A_281_74#_c_648_n 5.01714e-19 $X=4.785 $Y=1.22 $X2=0 $Y2=0
cc_297 N_VPWR_c_371_n N_A_241_368#_c_434_n 0.0762465f $X=1.8 $Y=1.985 $X2=0
+ $Y2=0
cc_298 N_VPWR_c_373_n N_A_241_368#_c_434_n 0.011066f $X=1.635 $Y=3.33 $X2=0
+ $Y2=0
cc_299 N_VPWR_c_368_n N_A_241_368#_c_434_n 0.00915947f $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_300 N_VPWR_c_371_n N_A_241_368#_c_430_n 0.0199103f $X=1.8 $Y=1.985 $X2=0
+ $Y2=0
cc_301 N_VPWR_c_371_n N_A_241_368#_c_435_n 0.0762465f $X=1.8 $Y=1.985 $X2=0
+ $Y2=0
cc_302 N_VPWR_c_372_n N_A_241_368#_c_435_n 0.0778383f $X=2.7 $Y=1.985 $X2=0
+ $Y2=0
cc_303 N_VPWR_c_374_n N_A_241_368#_c_435_n 0.0110241f $X=2.535 $Y=3.33 $X2=0
+ $Y2=0
cc_304 N_VPWR_c_368_n N_A_241_368#_c_435_n 0.00909194f $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_305 N_VPWR_c_372_n N_A_241_368#_c_432_n 0.0263643f $X=2.7 $Y=1.985 $X2=0
+ $Y2=0
cc_306 N_VPWR_c_372_n N_A_241_368#_c_436_n 0.0397705f $X=2.7 $Y=1.985 $X2=0
+ $Y2=0
cc_307 N_VPWR_c_375_n N_A_241_368#_c_437_n 0.0460675f $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_308 N_VPWR_c_368_n N_A_241_368#_c_437_n 0.0260697f $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_309 N_VPWR_c_372_n N_A_241_368#_c_438_n 0.0119239f $X=2.7 $Y=1.985 $X2=0
+ $Y2=0
cc_310 N_VPWR_c_375_n N_A_241_368#_c_438_n 0.0178001f $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_311 N_VPWR_c_368_n N_A_241_368#_c_438_n 0.00964081f $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_312 N_VPWR_c_375_n N_A_241_368#_c_439_n 0.0640155f $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_313 N_VPWR_c_368_n N_A_241_368#_c_439_n 0.0357926f $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_314 N_VPWR_c_375_n N_A_241_368#_c_441_n 0.0121867f $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_315 N_VPWR_c_368_n N_A_241_368#_c_441_n 0.00660921f $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_316 N_A_241_368#_c_437_n N_Z_M1001_d 0.00197722f $X=4.015 $Y=2.99 $X2=0 $Y2=0
cc_317 N_A_241_368#_c_439_n N_Z_M1010_d 0.00197722f $X=4.915 $Y=2.99 $X2=0 $Y2=0
cc_318 N_A_241_368#_c_437_n N_Z_c_529_n 0.0160777f $X=4.015 $Y=2.99 $X2=0 $Y2=0
cc_319 N_A_241_368#_c_480_n N_Z_c_529_n 0.0439674f $X=4.1 $Y=2.225 $X2=0 $Y2=0
cc_320 N_A_241_368#_M1005_s N_Z_c_531_n 0.00247267f $X=3.95 $Y=1.84 $X2=0 $Y2=0
cc_321 N_A_241_368#_c_480_n N_Z_c_531_n 0.0136682f $X=4.1 $Y=2.225 $X2=0 $Y2=0
cc_322 N_A_241_368#_c_440_n N_Z_c_531_n 0.00501285f $X=5 $Y=1.985 $X2=0 $Y2=0
cc_323 N_A_241_368#_c_480_n N_Z_c_540_n 0.0439674f $X=4.1 $Y=2.225 $X2=0 $Y2=0
cc_324 N_A_241_368#_c_439_n N_Z_c_540_n 0.0160777f $X=4.915 $Y=2.99 $X2=0 $Y2=0
cc_325 N_A_241_368#_c_440_n N_Z_c_540_n 0.0566253f $X=5 $Y=1.985 $X2=0 $Y2=0
cc_326 N_A_241_368#_c_432_n Z 0.00746325f $X=3.035 $Y=1.565 $X2=0 $Y2=0
cc_327 N_A_241_368#_c_436_n Z 0.0729293f $X=3.2 $Y=1.985 $X2=0 $Y2=0
cc_328 N_A_241_368#_c_432_n N_Z_c_527_n 0.00346621f $X=3.035 $Y=1.565 $X2=0
+ $Y2=0
cc_329 N_A_241_368#_c_430_n N_A_281_74#_c_639_n 0.0320456f $X=2.085 $Y=1.565
+ $X2=0 $Y2=0
cc_330 N_A_241_368#_c_433_n N_A_281_74#_c_639_n 0.0192612f $X=2.21 $Y=1.565
+ $X2=0 $Y2=0
cc_331 N_A_241_368#_c_430_n N_A_281_74#_c_640_n 0.0135853f $X=2.085 $Y=1.565
+ $X2=0 $Y2=0
cc_332 N_A_241_368#_c_432_n N_A_281_74#_c_642_n 0.0600906f $X=3.035 $Y=1.565
+ $X2=0 $Y2=0
cc_333 N_A_241_368#_c_432_n N_A_281_74#_c_670_n 0.0127483f $X=3.035 $Y=1.565
+ $X2=0 $Y2=0
cc_334 N_A_241_368#_c_433_n N_A_281_74#_c_670_n 8.91514e-19 $X=2.21 $Y=1.565
+ $X2=0 $Y2=0
cc_335 N_Z_c_536_n N_A_281_74#_M1004_d 0.00351264f $X=4.485 $Y=0.89 $X2=0 $Y2=0
cc_336 N_Z_c_527_n N_A_281_74#_c_642_n 0.0127735f $X=3.65 $Y=1.55 $X2=0 $Y2=0
cc_337 N_Z_c_526_n N_A_281_74#_c_644_n 0.0137359f $X=3.74 $Y=0.89 $X2=0 $Y2=0
cc_338 N_Z_M1000_s N_A_281_74#_c_645_n 0.00171549f $X=3.56 $Y=0.37 $X2=0 $Y2=0
cc_339 N_Z_c_536_n N_A_281_74#_c_645_n 0.023966f $X=4.485 $Y=0.89 $X2=0 $Y2=0
cc_340 N_Z_c_526_n N_A_281_74#_c_645_n 0.0154405f $X=3.74 $Y=0.89 $X2=0 $Y2=0
cc_341 N_Z_M1008_s N_A_281_74#_c_646_n 0.00176461f $X=4.43 $Y=0.37 $X2=0 $Y2=0
cc_342 N_Z_c_536_n N_A_281_74#_c_646_n 0.00424866f $X=4.485 $Y=0.89 $X2=0 $Y2=0
cc_343 N_Z_c_546_n N_A_281_74#_c_646_n 0.0121701f $X=4.57 $Y=0.8 $X2=0 $Y2=0
cc_344 N_VGND_c_579_n N_A_281_74#_c_638_n 0.0229082f $X=1.98 $Y=0.515 $X2=0
+ $Y2=0
cc_345 N_VGND_c_581_n N_A_281_74#_c_638_n 0.00749631f $X=1.815 $Y=0 $X2=0 $Y2=0
cc_346 N_VGND_c_586_n N_A_281_74#_c_638_n 0.0062048f $X=5.04 $Y=0 $X2=0 $Y2=0
cc_347 N_VGND_c_579_n N_A_281_74#_c_639_n 0.0216086f $X=1.98 $Y=0.515 $X2=0
+ $Y2=0
cc_348 N_VGND_c_579_n N_A_281_74#_c_641_n 0.0229082f $X=1.98 $Y=0.515 $X2=0
+ $Y2=0
cc_349 N_VGND_c_580_n N_A_281_74#_c_641_n 0.0229082f $X=2.84 $Y=0.515 $X2=0
+ $Y2=0
cc_350 N_VGND_c_583_n N_A_281_74#_c_641_n 0.00749631f $X=2.675 $Y=0 $X2=0 $Y2=0
cc_351 N_VGND_c_586_n N_A_281_74#_c_641_n 0.0062048f $X=5.04 $Y=0 $X2=0 $Y2=0
cc_352 N_VGND_c_580_n N_A_281_74#_c_642_n 0.0216086f $X=2.84 $Y=0.515 $X2=0
+ $Y2=0
cc_353 N_VGND_c_580_n N_A_281_74#_c_643_n 0.0175237f $X=2.84 $Y=0.515 $X2=0
+ $Y2=0
cc_354 N_VGND_c_585_n N_A_281_74#_c_643_n 0.0178338f $X=5.04 $Y=0 $X2=0 $Y2=0
cc_355 N_VGND_c_586_n N_A_281_74#_c_643_n 0.00960503f $X=5.04 $Y=0 $X2=0 $Y2=0
cc_356 N_VGND_c_585_n N_A_281_74#_c_645_n 0.0912556f $X=5.04 $Y=0 $X2=0 $Y2=0
cc_357 N_VGND_c_586_n N_A_281_74#_c_645_n 0.0506361f $X=5.04 $Y=0 $X2=0 $Y2=0
cc_358 N_VGND_c_585_n N_A_281_74#_c_646_n 0.0235688f $X=5.04 $Y=0 $X2=0 $Y2=0
cc_359 N_VGND_c_586_n N_A_281_74#_c_646_n 0.0127152f $X=5.04 $Y=0 $X2=0 $Y2=0
