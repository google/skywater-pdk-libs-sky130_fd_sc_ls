* File: sky130_fd_sc_ls__o21bai_2.pxi.spice
* Created: Fri Aug 28 13:46:47 2020
* 
x_PM_SKY130_FD_SC_LS__O21BAI_2%B1_N N_B1_N_M1012_g N_B1_N_c_79_n N_B1_N_M1011_g
+ B1_N N_B1_N_c_80_n PM_SKY130_FD_SC_LS__O21BAI_2%B1_N
x_PM_SKY130_FD_SC_LS__O21BAI_2%A_27_74# N_A_27_74#_M1012_s N_A_27_74#_M1011_s
+ N_A_27_74#_c_121_n N_A_27_74#_M1006_g N_A_27_74#_c_111_n N_A_27_74#_M1005_g
+ N_A_27_74#_c_112_n N_A_27_74#_c_113_n N_A_27_74#_M1013_g N_A_27_74#_c_123_n
+ N_A_27_74#_M1010_g N_A_27_74#_c_114_n N_A_27_74#_c_115_n N_A_27_74#_c_116_n
+ N_A_27_74#_c_125_n N_A_27_74#_c_117_n N_A_27_74#_c_118_n N_A_27_74#_c_119_n
+ N_A_27_74#_c_126_n N_A_27_74#_c_120_n PM_SKY130_FD_SC_LS__O21BAI_2%A_27_74#
x_PM_SKY130_FD_SC_LS__O21BAI_2%A1 N_A1_M1001_g N_A1_c_199_n N_A1_M1000_g
+ N_A1_M1004_g N_A1_c_201_n N_A1_M1009_g N_A1_c_202_n N_A1_c_217_p N_A1_c_214_n
+ A1 N_A1_c_203_n A1 PM_SKY130_FD_SC_LS__O21BAI_2%A1
x_PM_SKY130_FD_SC_LS__O21BAI_2%A2 N_A2_c_283_n N_A2_M1003_g N_A2_M1002_g
+ N_A2_c_284_n N_A2_M1007_g N_A2_M1008_g A2 N_A2_c_281_n N_A2_c_282_n
+ PM_SKY130_FD_SC_LS__O21BAI_2%A2
x_PM_SKY130_FD_SC_LS__O21BAI_2%VPWR N_VPWR_M1011_d N_VPWR_M1010_s N_VPWR_M1009_s
+ N_VPWR_c_339_n N_VPWR_c_340_n N_VPWR_c_341_n N_VPWR_c_342_n VPWR
+ N_VPWR_c_343_n N_VPWR_c_344_n N_VPWR_c_345_n N_VPWR_c_346_n N_VPWR_c_347_n
+ N_VPWR_c_338_n PM_SKY130_FD_SC_LS__O21BAI_2%VPWR
x_PM_SKY130_FD_SC_LS__O21BAI_2%Y N_Y_M1005_s N_Y_M1006_d N_Y_M1003_d N_Y_c_394_n
+ N_Y_c_400_n N_Y_c_420_n N_Y_c_396_n Y Y Y Y PM_SKY130_FD_SC_LS__O21BAI_2%Y
x_PM_SKY130_FD_SC_LS__O21BAI_2%A_507_368# N_A_507_368#_M1000_d
+ N_A_507_368#_M1007_s N_A_507_368#_c_440_n N_A_507_368#_c_446_n
+ N_A_507_368#_c_441_n PM_SKY130_FD_SC_LS__O21BAI_2%A_507_368#
x_PM_SKY130_FD_SC_LS__O21BAI_2%VGND N_VGND_M1012_d N_VGND_M1001_s N_VGND_M1008_s
+ N_VGND_c_471_n N_VGND_c_472_n N_VGND_c_473_n VGND N_VGND_c_474_n
+ N_VGND_c_475_n N_VGND_c_476_n N_VGND_c_477_n N_VGND_c_478_n N_VGND_c_479_n
+ N_VGND_c_480_n N_VGND_c_481_n PM_SKY130_FD_SC_LS__O21BAI_2%VGND
x_PM_SKY130_FD_SC_LS__O21BAI_2%A_225_74# N_A_225_74#_M1005_d N_A_225_74#_M1013_d
+ N_A_225_74#_M1002_d N_A_225_74#_M1004_d N_A_225_74#_c_525_n
+ N_A_225_74#_c_526_n N_A_225_74#_c_527_n N_A_225_74#_c_546_n
+ N_A_225_74#_c_528_n N_A_225_74#_c_529_n N_A_225_74#_c_530_n
+ N_A_225_74#_c_531_n N_A_225_74#_c_532_n N_A_225_74#_c_533_n
+ PM_SKY130_FD_SC_LS__O21BAI_2%A_225_74#
cc_1 VNB N_B1_N_M1012_g 0.0392908f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.69
cc_2 VNB N_B1_N_c_79_n 0.0306379f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.765
cc_3 VNB N_B1_N_c_80_n 0.00536388f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.515
cc_4 VNB N_A_27_74#_c_111_n 0.0184105f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.515
cc_5 VNB N_A_27_74#_c_112_n 0.00663413f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_A_27_74#_c_113_n 0.016529f $X=-0.19 $Y=-0.245 $X2=0.647 $Y2=1.665
cc_7 VNB N_A_27_74#_c_114_n 0.0396459f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_27_74#_c_115_n 0.0411124f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_27_74#_c_116_n 0.0266107f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_27_74#_c_117_n 0.0243345f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_27_74#_c_118_n 0.00511234f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_74#_c_119_n 0.0109678f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_74#_c_120_n 0.022547f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A1_M1001_g 0.025715f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.69
cc_15 VNB N_A1_c_199_n 0.0270222f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.765
cc_16 VNB N_A1_M1004_g 0.030416f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.515
cc_17 VNB N_A1_c_201_n 0.0354747f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.515
cc_18 VNB N_A1_c_202_n 0.00166985f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A1_c_203_n 0.0191473f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB A1 8.32086e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A2_M1002_g 0.024925f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=2.34
cc_22 VNB N_A2_M1008_g 0.0230333f $X=-0.19 $Y=-0.245 $X2=0.647 $Y2=1.515
cc_23 VNB N_A2_c_281_n 0.00138642f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A2_c_282_n 0.03662f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VPWR_c_338_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_Y_c_394_n 4.51115e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB Y 0.00224001f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_471_n 0.0107462f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.515
cc_29 VNB N_VGND_c_472_n 0.00842841f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_473_n 0.00327765f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_474_n 0.0173909f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_475_n 0.0405043f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_476_n 0.0162351f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_477_n 0.0180274f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_478_n 0.262471f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_479_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_480_n 0.00634377f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_481_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_225_74#_c_525_n 0.00379275f $X=-0.19 $Y=-0.245 $X2=0.647 $Y2=1.665
cc_40 VNB N_A_225_74#_c_526_n 0.00452721f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_225_74#_c_527_n 0.00417961f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_225_74#_c_528_n 0.00968069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_225_74#_c_529_n 0.0100176f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_225_74#_c_530_n 0.00179461f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_225_74#_c_531_n 0.015761f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_225_74#_c_532_n 0.0255089f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_225_74#_c_533_n 0.00193677f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VPB N_B1_N_c_79_n 0.0347524f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.765
cc_49 VPB N_B1_N_c_80_n 0.00650654f $X=-0.19 $Y=1.66 $X2=0.625 $Y2=1.515
cc_50 VPB N_A_27_74#_c_121_n 0.0166835f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=2.34
cc_51 VPB N_A_27_74#_c_112_n 6.93118e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_A_27_74#_c_123_n 0.0212458f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_A_27_74#_c_115_n 0.00761635f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_A_27_74#_c_125_n 0.0358186f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_A_27_74#_c_126_n 0.0137373f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_A_27_74#_c_120_n 0.0143493f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_A1_c_199_n 0.0260039f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.765
cc_58 VPB N_A1_c_201_n 0.0278171f $X=-0.19 $Y=1.66 $X2=0.625 $Y2=1.515
cc_59 VPB N_A1_c_202_n 0.00270844f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB A1 0.00324651f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_A2_c_283_n 0.0147591f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.35
cc_62 VPB N_A2_c_284_n 0.0149173f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_63 VPB N_A2_c_281_n 0.00322323f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_A2_c_282_n 0.020345f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_339_n 0.015617f $X=-0.19 $Y=1.66 $X2=0.625 $Y2=1.515
cc_66 VPB N_VPWR_c_340_n 0.00595534f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_341_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_342_n 0.0577101f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_343_n 0.030897f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_344_n 0.0183662f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_345_n 0.0388892f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_346_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_347_n 0.00690733f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_338_n 0.079556f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_Y_c_396_n 0.00216998f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_A_507_368#_c_440_n 0.00435633f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=2.34
cc_77 VPB N_A_507_368#_c_441_n 0.00216812f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 N_B1_N_c_79_n N_A_27_74#_c_121_n 0.0131934f $X=0.7 $Y=1.765 $X2=0 $Y2=0
cc_79 N_B1_N_c_80_n N_A_27_74#_c_121_n 2.54649e-19 $X=0.625 $Y=1.515 $X2=0 $Y2=0
cc_80 N_B1_N_M1012_g N_A_27_74#_c_114_n 0.0040089f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_81 N_B1_N_c_79_n N_A_27_74#_c_114_n 0.0111951f $X=0.7 $Y=1.765 $X2=0 $Y2=0
cc_82 N_B1_N_c_80_n N_A_27_74#_c_114_n 0.00135338f $X=0.625 $Y=1.515 $X2=0 $Y2=0
cc_83 N_B1_N_c_79_n N_A_27_74#_c_115_n 0.00318173f $X=0.7 $Y=1.765 $X2=0 $Y2=0
cc_84 N_B1_N_c_80_n N_A_27_74#_c_115_n 0.00376061f $X=0.625 $Y=1.515 $X2=0 $Y2=0
cc_85 N_B1_N_M1012_g N_A_27_74#_c_116_n 4.43891e-19 $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_86 N_B1_N_c_79_n N_A_27_74#_c_125_n 0.0102926f $X=0.7 $Y=1.765 $X2=0 $Y2=0
cc_87 N_B1_N_M1012_g N_A_27_74#_c_117_n 0.0189149f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_88 N_B1_N_c_79_n N_A_27_74#_c_117_n 0.00153593f $X=0.7 $Y=1.765 $X2=0 $Y2=0
cc_89 N_B1_N_c_80_n N_A_27_74#_c_117_n 0.0285306f $X=0.625 $Y=1.515 $X2=0 $Y2=0
cc_90 N_B1_N_M1012_g N_A_27_74#_c_118_n 0.00179141f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_91 N_B1_N_c_79_n N_A_27_74#_c_118_n 2.33686e-19 $X=0.7 $Y=1.765 $X2=0 $Y2=0
cc_92 N_B1_N_c_80_n N_A_27_74#_c_118_n 0.014429f $X=0.625 $Y=1.515 $X2=0 $Y2=0
cc_93 N_B1_N_c_79_n N_A_27_74#_c_126_n 0.0066951f $X=0.7 $Y=1.765 $X2=0 $Y2=0
cc_94 N_B1_N_c_80_n N_A_27_74#_c_126_n 0.013098f $X=0.625 $Y=1.515 $X2=0 $Y2=0
cc_95 N_B1_N_M1012_g N_A_27_74#_c_120_n 0.0139236f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_96 N_B1_N_c_79_n N_A_27_74#_c_120_n 0.00377891f $X=0.7 $Y=1.765 $X2=0 $Y2=0
cc_97 N_B1_N_c_80_n N_A_27_74#_c_120_n 0.0323502f $X=0.625 $Y=1.515 $X2=0 $Y2=0
cc_98 N_B1_N_c_79_n N_VPWR_c_339_n 0.0153815f $X=0.7 $Y=1.765 $X2=0 $Y2=0
cc_99 N_B1_N_c_79_n N_VPWR_c_343_n 0.00481995f $X=0.7 $Y=1.765 $X2=0 $Y2=0
cc_100 N_B1_N_c_79_n N_VPWR_c_338_n 0.00508379f $X=0.7 $Y=1.765 $X2=0 $Y2=0
cc_101 N_B1_N_M1012_g N_VGND_c_471_n 0.0156976f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_102 N_B1_N_M1012_g N_VGND_c_474_n 0.00383152f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_103 N_B1_N_M1012_g N_VGND_c_478_n 0.00761198f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_104 N_B1_N_M1012_g N_A_225_74#_c_525_n 8.38994e-19 $X=0.495 $Y=0.69 $X2=0
+ $Y2=0
cc_105 N_B1_N_M1012_g N_A_225_74#_c_527_n 7.24903e-19 $X=0.495 $Y=0.69 $X2=0
+ $Y2=0
cc_106 N_A_27_74#_c_113_n N_A1_M1001_g 0.0238637f $X=1.915 $Y=1.22 $X2=0 $Y2=0
cc_107 N_A_27_74#_c_123_n N_A1_c_199_n 0.0344574f $X=1.92 $Y=1.765 $X2=0 $Y2=0
cc_108 N_A_27_74#_c_115_n N_A1_c_199_n 0.0176849f $X=1.915 $Y=1.492 $X2=0 $Y2=0
cc_109 N_A_27_74#_c_123_n N_A1_c_202_n 0.00224923f $X=1.92 $Y=1.765 $X2=0 $Y2=0
cc_110 N_A_27_74#_c_115_n N_A1_c_202_n 0.00136385f $X=1.915 $Y=1.492 $X2=0 $Y2=0
cc_111 N_A_27_74#_c_123_n N_A1_c_214_n 0.00156633f $X=1.92 $Y=1.765 $X2=0 $Y2=0
cc_112 N_A_27_74#_c_121_n N_VPWR_c_339_n 0.0167791f $X=1.47 $Y=1.765 $X2=0 $Y2=0
cc_113 N_A_27_74#_c_114_n N_VPWR_c_339_n 0.00226699f $X=1.38 $Y=1.385 $X2=0
+ $Y2=0
cc_114 N_A_27_74#_c_117_n N_VPWR_c_339_n 7.87179e-19 $X=1.03 $Y=1.095 $X2=0
+ $Y2=0
cc_115 N_A_27_74#_c_118_n N_VPWR_c_339_n 0.0187766f $X=1.195 $Y=1.385 $X2=0
+ $Y2=0
cc_116 N_A_27_74#_c_126_n N_VPWR_c_339_n 0.0406203f $X=0.475 $Y=2.035 $X2=0
+ $Y2=0
cc_117 N_A_27_74#_c_121_n N_VPWR_c_340_n 4.44619e-19 $X=1.47 $Y=1.765 $X2=0
+ $Y2=0
cc_118 N_A_27_74#_c_123_n N_VPWR_c_340_n 0.00761915f $X=1.92 $Y=1.765 $X2=0
+ $Y2=0
cc_119 N_A_27_74#_c_125_n N_VPWR_c_343_n 0.0156448f $X=0.475 $Y=2.715 $X2=0
+ $Y2=0
cc_120 N_A_27_74#_c_121_n N_VPWR_c_344_n 0.00445602f $X=1.47 $Y=1.765 $X2=0
+ $Y2=0
cc_121 N_A_27_74#_c_123_n N_VPWR_c_344_n 0.00413917f $X=1.92 $Y=1.765 $X2=0
+ $Y2=0
cc_122 N_A_27_74#_c_121_n N_VPWR_c_338_n 0.00862279f $X=1.47 $Y=1.765 $X2=0
+ $Y2=0
cc_123 N_A_27_74#_c_123_n N_VPWR_c_338_n 0.00817726f $X=1.92 $Y=1.765 $X2=0
+ $Y2=0
cc_124 N_A_27_74#_c_125_n N_VPWR_c_338_n 0.0178521f $X=0.475 $Y=2.715 $X2=0
+ $Y2=0
cc_125 N_A_27_74#_c_111_n N_Y_c_394_n 0.00107507f $X=1.485 $Y=1.22 $X2=0 $Y2=0
cc_126 N_A_27_74#_c_113_n N_Y_c_394_n 0.00779056f $X=1.915 $Y=1.22 $X2=0 $Y2=0
cc_127 N_A_27_74#_c_117_n N_Y_c_394_n 0.00446815f $X=1.03 $Y=1.095 $X2=0 $Y2=0
cc_128 N_A_27_74#_c_123_n N_Y_c_400_n 0.0153804f $X=1.92 $Y=1.765 $X2=0 $Y2=0
cc_129 N_A_27_74#_c_121_n N_Y_c_396_n 0.00788856f $X=1.47 $Y=1.765 $X2=0 $Y2=0
cc_130 N_A_27_74#_c_123_n N_Y_c_396_n 0.00655006f $X=1.92 $Y=1.765 $X2=0 $Y2=0
cc_131 N_A_27_74#_c_121_n Y 0.00852736f $X=1.47 $Y=1.765 $X2=0 $Y2=0
cc_132 N_A_27_74#_c_111_n Y 0.00240384f $X=1.485 $Y=1.22 $X2=0 $Y2=0
cc_133 N_A_27_74#_c_112_n Y 0.00411229f $X=1.92 $Y=1.675 $X2=0 $Y2=0
cc_134 N_A_27_74#_c_113_n Y 0.0012234f $X=1.915 $Y=1.22 $X2=0 $Y2=0
cc_135 N_A_27_74#_c_123_n Y 0.0126986f $X=1.92 $Y=1.765 $X2=0 $Y2=0
cc_136 N_A_27_74#_c_115_n Y 0.0359062f $X=1.915 $Y=1.492 $X2=0 $Y2=0
cc_137 N_A_27_74#_c_118_n Y 0.0278451f $X=1.195 $Y=1.385 $X2=0 $Y2=0
cc_138 N_A_27_74#_c_111_n N_VGND_c_471_n 0.00184366f $X=1.485 $Y=1.22 $X2=0
+ $Y2=0
cc_139 N_A_27_74#_c_116_n N_VGND_c_471_n 0.0182902f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_140 N_A_27_74#_c_117_n N_VGND_c_471_n 0.0243991f $X=1.03 $Y=1.095 $X2=0 $Y2=0
cc_141 N_A_27_74#_c_116_n N_VGND_c_474_n 0.011066f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_142 N_A_27_74#_c_111_n N_VGND_c_475_n 0.00278247f $X=1.485 $Y=1.22 $X2=0
+ $Y2=0
cc_143 N_A_27_74#_c_113_n N_VGND_c_475_n 0.00278271f $X=1.915 $Y=1.22 $X2=0
+ $Y2=0
cc_144 N_A_27_74#_c_111_n N_VGND_c_478_n 0.00358425f $X=1.485 $Y=1.22 $X2=0
+ $Y2=0
cc_145 N_A_27_74#_c_113_n N_VGND_c_478_n 0.0035414f $X=1.915 $Y=1.22 $X2=0 $Y2=0
cc_146 N_A_27_74#_c_116_n N_VGND_c_478_n 0.00915947f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_147 N_A_27_74#_c_117_n N_A_225_74#_M1005_d 0.00281428f $X=1.03 $Y=1.095
+ $X2=-0.19 $Y2=-0.245
cc_148 N_A_27_74#_c_111_n N_A_225_74#_c_525_n 0.00809982f $X=1.485 $Y=1.22 $X2=0
+ $Y2=0
cc_149 N_A_27_74#_c_113_n N_A_225_74#_c_525_n 5.5293e-19 $X=1.915 $Y=1.22 $X2=0
+ $Y2=0
cc_150 N_A_27_74#_c_114_n N_A_225_74#_c_525_n 0.00120271f $X=1.38 $Y=1.385 $X2=0
+ $Y2=0
cc_151 N_A_27_74#_c_117_n N_A_225_74#_c_525_n 0.0217145f $X=1.03 $Y=1.095 $X2=0
+ $Y2=0
cc_152 N_A_27_74#_c_111_n N_A_225_74#_c_526_n 0.0100711f $X=1.485 $Y=1.22 $X2=0
+ $Y2=0
cc_153 N_A_27_74#_c_113_n N_A_225_74#_c_526_n 0.0133867f $X=1.915 $Y=1.22 $X2=0
+ $Y2=0
cc_154 N_A_27_74#_c_111_n N_A_225_74#_c_527_n 0.00395315f $X=1.485 $Y=1.22 $X2=0
+ $Y2=0
cc_155 N_A_27_74#_c_113_n N_A_225_74#_c_529_n 0.00116009f $X=1.915 $Y=1.22 $X2=0
+ $Y2=0
cc_156 N_A1_c_199_n N_A2_c_283_n 0.0410296f $X=2.46 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_157 N_A1_c_202_n N_A2_c_283_n 0.00165633f $X=2.415 $Y=1.515 $X2=-0.19
+ $Y2=-0.245
cc_158 N_A1_c_217_p N_A2_c_283_n 0.0106753f $X=3.485 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_159 N_A1_M1001_g N_A2_M1002_g 0.0254412f $X=2.415 $Y=0.74 $X2=0 $Y2=0
cc_160 N_A1_c_201_n N_A2_c_284_n 0.0215775f $X=3.815 $Y=1.765 $X2=0 $Y2=0
cc_161 N_A1_c_217_p N_A2_c_284_n 0.0191296f $X=3.485 $Y=2.035 $X2=0 $Y2=0
cc_162 A1 N_A2_c_284_n 0.00215749f $X=3.6 $Y=1.665 $X2=0 $Y2=0
cc_163 N_A1_M1004_g N_A2_M1008_g 0.0314638f $X=3.805 $Y=0.74 $X2=0 $Y2=0
cc_164 N_A1_c_201_n N_A2_M1008_g 0.0192099f $X=3.815 $Y=1.765 $X2=0 $Y2=0
cc_165 N_A1_c_203_n N_A2_M1008_g 0.0043055f $X=3.89 $Y=1.485 $X2=0 $Y2=0
cc_166 N_A1_c_199_n N_A2_c_281_n 0.00137209f $X=2.46 $Y=1.765 $X2=0 $Y2=0
cc_167 N_A1_c_201_n N_A2_c_281_n 2.15819e-19 $X=3.815 $Y=1.765 $X2=0 $Y2=0
cc_168 N_A1_c_202_n N_A2_c_281_n 0.0254228f $X=2.415 $Y=1.515 $X2=0 $Y2=0
cc_169 N_A1_c_217_p N_A2_c_281_n 0.0292378f $X=3.485 $Y=2.035 $X2=0 $Y2=0
cc_170 N_A1_c_203_n N_A2_c_281_n 0.0189163f $X=3.89 $Y=1.485 $X2=0 $Y2=0
cc_171 A1 N_A2_c_281_n 0.00805578f $X=3.6 $Y=1.665 $X2=0 $Y2=0
cc_172 N_A1_c_199_n N_A2_c_282_n 0.0216797f $X=2.46 $Y=1.765 $X2=0 $Y2=0
cc_173 N_A1_c_202_n N_A2_c_282_n 0.00188444f $X=2.415 $Y=1.515 $X2=0 $Y2=0
cc_174 N_A1_c_217_p N_A2_c_282_n 0.00117801f $X=3.485 $Y=2.035 $X2=0 $Y2=0
cc_175 A1 N_A2_c_282_n 0.00106815f $X=3.6 $Y=1.665 $X2=0 $Y2=0
cc_176 N_A1_c_202_n N_VPWR_M1010_s 0.00135567f $X=2.415 $Y=1.515 $X2=0 $Y2=0
cc_177 N_A1_c_214_n N_VPWR_M1010_s 0.00301618f $X=2.58 $Y=2.035 $X2=0 $Y2=0
cc_178 N_A1_c_199_n N_VPWR_c_340_n 0.00329185f $X=2.46 $Y=1.765 $X2=0 $Y2=0
cc_179 N_A1_c_201_n N_VPWR_c_342_n 0.0139116f $X=3.815 $Y=1.765 $X2=0 $Y2=0
cc_180 N_A1_c_203_n N_VPWR_c_342_n 0.008349f $X=3.89 $Y=1.485 $X2=0 $Y2=0
cc_181 A1 N_VPWR_c_342_n 0.00449553f $X=3.6 $Y=1.665 $X2=0 $Y2=0
cc_182 N_A1_c_199_n N_VPWR_c_345_n 0.00444353f $X=2.46 $Y=1.765 $X2=0 $Y2=0
cc_183 N_A1_c_201_n N_VPWR_c_345_n 0.0044313f $X=3.815 $Y=1.765 $X2=0 $Y2=0
cc_184 N_A1_c_199_n N_VPWR_c_338_n 0.0085731f $X=2.46 $Y=1.765 $X2=0 $Y2=0
cc_185 N_A1_c_201_n N_VPWR_c_338_n 0.00856984f $X=3.815 $Y=1.765 $X2=0 $Y2=0
cc_186 N_A1_c_217_p N_Y_M1003_d 0.00381047f $X=3.485 $Y=2.035 $X2=0 $Y2=0
cc_187 N_A1_c_199_n N_Y_c_400_n 0.0153145f $X=2.46 $Y=1.765 $X2=0 $Y2=0
cc_188 N_A1_c_217_p N_Y_c_400_n 0.037593f $X=3.485 $Y=2.035 $X2=0 $Y2=0
cc_189 N_A1_c_214_n N_Y_c_400_n 0.0177274f $X=2.58 $Y=2.035 $X2=0 $Y2=0
cc_190 N_A1_M1001_g Y 7.96105e-19 $X=2.415 $Y=0.74 $X2=0 $Y2=0
cc_191 N_A1_c_199_n Y 0.00215496f $X=2.46 $Y=1.765 $X2=0 $Y2=0
cc_192 N_A1_c_202_n Y 0.0242167f $X=2.415 $Y=1.515 $X2=0 $Y2=0
cc_193 N_A1_c_214_n Y 0.00748808f $X=2.58 $Y=2.035 $X2=0 $Y2=0
cc_194 N_A1_c_217_p N_A_507_368#_M1000_d 0.00907897f $X=3.485 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_195 N_A1_c_217_p N_A_507_368#_M1007_s 0.00269219f $X=3.485 $Y=2.035 $X2=0
+ $Y2=0
cc_196 A1 N_A_507_368#_M1007_s 4.10256e-19 $X=3.6 $Y=1.665 $X2=0 $Y2=0
cc_197 N_A1_c_201_n N_A_507_368#_c_440_n 0.0033408f $X=3.815 $Y=1.765 $X2=0
+ $Y2=0
cc_198 N_A1_c_201_n N_A_507_368#_c_446_n 0.00761772f $X=3.815 $Y=1.765 $X2=0
+ $Y2=0
cc_199 N_A1_c_217_p N_A_507_368#_c_446_n 0.0177862f $X=3.485 $Y=2.035 $X2=0
+ $Y2=0
cc_200 N_A1_c_203_n N_A_507_368#_c_446_n 7.41312e-19 $X=3.89 $Y=1.485 $X2=0
+ $Y2=0
cc_201 N_A1_c_199_n N_A_507_368#_c_441_n 0.00611929f $X=2.46 $Y=1.765 $X2=0
+ $Y2=0
cc_202 N_A1_M1001_g N_VGND_c_472_n 0.00404801f $X=2.415 $Y=0.74 $X2=0 $Y2=0
cc_203 N_A1_M1004_g N_VGND_c_473_n 0.0129724f $X=3.805 $Y=0.74 $X2=0 $Y2=0
cc_204 N_A1_M1001_g N_VGND_c_475_n 0.00430908f $X=2.415 $Y=0.74 $X2=0 $Y2=0
cc_205 N_A1_M1004_g N_VGND_c_477_n 0.00383152f $X=3.805 $Y=0.74 $X2=0 $Y2=0
cc_206 N_A1_M1001_g N_VGND_c_478_n 0.00817122f $X=2.415 $Y=0.74 $X2=0 $Y2=0
cc_207 N_A1_M1004_g N_VGND_c_478_n 0.00761264f $X=3.805 $Y=0.74 $X2=0 $Y2=0
cc_208 N_A1_M1001_g N_A_225_74#_c_526_n 0.00347348f $X=2.415 $Y=0.74 $X2=0 $Y2=0
cc_209 N_A1_M1001_g N_A_225_74#_c_546_n 0.00831216f $X=2.415 $Y=0.74 $X2=0 $Y2=0
cc_210 N_A1_M1001_g N_A_225_74#_c_528_n 0.0116199f $X=2.415 $Y=0.74 $X2=0 $Y2=0
cc_211 N_A1_c_199_n N_A_225_74#_c_528_n 6.22749e-19 $X=2.46 $Y=1.765 $X2=0 $Y2=0
cc_212 N_A1_c_202_n N_A_225_74#_c_528_n 0.0166004f $X=2.415 $Y=1.515 $X2=0 $Y2=0
cc_213 N_A1_M1001_g N_A_225_74#_c_529_n 0.00158144f $X=2.415 $Y=0.74 $X2=0 $Y2=0
cc_214 N_A1_c_199_n N_A_225_74#_c_529_n 7.04412e-19 $X=2.46 $Y=1.765 $X2=0 $Y2=0
cc_215 N_A1_c_202_n N_A_225_74#_c_529_n 0.010051f $X=2.415 $Y=1.515 $X2=0 $Y2=0
cc_216 N_A1_M1004_g N_A_225_74#_c_531_n 0.012998f $X=3.805 $Y=0.74 $X2=0 $Y2=0
cc_217 N_A1_c_201_n N_A_225_74#_c_531_n 0.00420647f $X=3.815 $Y=1.765 $X2=0
+ $Y2=0
cc_218 N_A1_c_203_n N_A_225_74#_c_531_n 0.0443322f $X=3.89 $Y=1.485 $X2=0 $Y2=0
cc_219 N_A1_M1004_g N_A_225_74#_c_532_n 0.00159319f $X=3.805 $Y=0.74 $X2=0 $Y2=0
cc_220 N_A2_c_283_n N_VPWR_c_345_n 0.00279479f $X=2.91 $Y=1.765 $X2=0 $Y2=0
cc_221 N_A2_c_284_n N_VPWR_c_345_n 0.00278257f $X=3.36 $Y=1.765 $X2=0 $Y2=0
cc_222 N_A2_c_283_n N_VPWR_c_338_n 0.00352997f $X=2.91 $Y=1.765 $X2=0 $Y2=0
cc_223 N_A2_c_284_n N_VPWR_c_338_n 0.0035395f $X=3.36 $Y=1.765 $X2=0 $Y2=0
cc_224 N_A2_c_283_n N_Y_c_400_n 0.0100252f $X=2.91 $Y=1.765 $X2=0 $Y2=0
cc_225 N_A2_c_284_n N_Y_c_400_n 8.55285e-19 $X=3.36 $Y=1.765 $X2=0 $Y2=0
cc_226 N_A2_c_283_n N_Y_c_420_n 0.00374827f $X=2.91 $Y=1.765 $X2=0 $Y2=0
cc_227 N_A2_c_284_n N_Y_c_420_n 9.95708e-19 $X=3.36 $Y=1.765 $X2=0 $Y2=0
cc_228 N_A2_c_283_n N_A_507_368#_c_440_n 0.00857014f $X=2.91 $Y=1.765 $X2=0
+ $Y2=0
cc_229 N_A2_c_284_n N_A_507_368#_c_440_n 0.0125777f $X=3.36 $Y=1.765 $X2=0 $Y2=0
cc_230 N_A2_c_283_n N_A_507_368#_c_446_n 6.467e-19 $X=2.91 $Y=1.765 $X2=0 $Y2=0
cc_231 N_A2_c_284_n N_A_507_368#_c_446_n 0.00827398f $X=3.36 $Y=1.765 $X2=0
+ $Y2=0
cc_232 N_A2_c_283_n N_A_507_368#_c_441_n 0.0064347f $X=2.91 $Y=1.765 $X2=0 $Y2=0
cc_233 N_A2_c_284_n N_A_507_368#_c_441_n 6.14126e-19 $X=3.36 $Y=1.765 $X2=0
+ $Y2=0
cc_234 N_A2_M1002_g N_VGND_c_472_n 0.00261709f $X=2.945 $Y=0.74 $X2=0 $Y2=0
cc_235 N_A2_M1002_g N_VGND_c_473_n 4.66963e-19 $X=2.945 $Y=0.74 $X2=0 $Y2=0
cc_236 N_A2_M1008_g N_VGND_c_473_n 0.00999938f $X=3.375 $Y=0.74 $X2=0 $Y2=0
cc_237 N_A2_M1002_g N_VGND_c_476_n 0.00461464f $X=2.945 $Y=0.74 $X2=0 $Y2=0
cc_238 N_A2_M1008_g N_VGND_c_476_n 0.00383152f $X=3.375 $Y=0.74 $X2=0 $Y2=0
cc_239 N_A2_M1002_g N_VGND_c_478_n 0.00908164f $X=2.945 $Y=0.74 $X2=0 $Y2=0
cc_240 N_A2_M1008_g N_VGND_c_478_n 0.0075754f $X=3.375 $Y=0.74 $X2=0 $Y2=0
cc_241 N_A2_M1002_g N_A_225_74#_c_546_n 8.0819e-19 $X=2.945 $Y=0.74 $X2=0 $Y2=0
cc_242 N_A2_M1002_g N_A_225_74#_c_528_n 0.0142114f $X=2.945 $Y=0.74 $X2=0 $Y2=0
cc_243 N_A2_c_281_n N_A_225_74#_c_528_n 0.0189798f $X=3.03 $Y=1.515 $X2=0 $Y2=0
cc_244 N_A2_c_282_n N_A_225_74#_c_528_n 3.41739e-19 $X=3.36 $Y=1.557 $X2=0 $Y2=0
cc_245 N_A2_M1002_g N_A_225_74#_c_530_n 4.00651e-19 $X=2.945 $Y=0.74 $X2=0 $Y2=0
cc_246 N_A2_M1008_g N_A_225_74#_c_530_n 3.92313e-19 $X=3.375 $Y=0.74 $X2=0 $Y2=0
cc_247 N_A2_M1008_g N_A_225_74#_c_531_n 0.0172403f $X=3.375 $Y=0.74 $X2=0 $Y2=0
cc_248 N_A2_M1008_g N_A_225_74#_c_533_n 9.49306e-19 $X=3.375 $Y=0.74 $X2=0 $Y2=0
cc_249 N_A2_c_281_n N_A_225_74#_c_533_n 0.0137234f $X=3.03 $Y=1.515 $X2=0 $Y2=0
cc_250 N_A2_c_282_n N_A_225_74#_c_533_n 7.91474e-19 $X=3.36 $Y=1.557 $X2=0 $Y2=0
cc_251 N_VPWR_M1010_s N_Y_c_400_n 0.01166f $X=1.995 $Y=1.84 $X2=0 $Y2=0
cc_252 N_VPWR_c_340_n N_Y_c_400_n 0.0216022f $X=2.165 $Y=2.815 $X2=0 $Y2=0
cc_253 N_VPWR_c_339_n N_Y_c_396_n 0.0481799f $X=1.17 $Y=1.985 $X2=0 $Y2=0
cc_254 N_VPWR_c_340_n N_Y_c_396_n 0.0223484f $X=2.165 $Y=2.815 $X2=0 $Y2=0
cc_255 N_VPWR_c_344_n N_Y_c_396_n 0.0110241f $X=1.98 $Y=3.33 $X2=0 $Y2=0
cc_256 N_VPWR_c_338_n N_Y_c_396_n 0.00909194f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_257 N_VPWR_c_339_n Y 0.0328581f $X=1.17 $Y=1.985 $X2=0 $Y2=0
cc_258 N_VPWR_c_342_n N_A_507_368#_c_440_n 0.012272f $X=4.04 $Y=1.985 $X2=0
+ $Y2=0
cc_259 N_VPWR_c_345_n N_A_507_368#_c_440_n 0.0597832f $X=3.955 $Y=3.33 $X2=0
+ $Y2=0
cc_260 N_VPWR_c_338_n N_A_507_368#_c_440_n 0.0330807f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_261 N_VPWR_c_342_n N_A_507_368#_c_446_n 0.0412501f $X=4.04 $Y=1.985 $X2=0
+ $Y2=0
cc_262 N_VPWR_c_340_n N_A_507_368#_c_441_n 0.0207727f $X=2.165 $Y=2.815 $X2=0
+ $Y2=0
cc_263 N_VPWR_c_345_n N_A_507_368#_c_441_n 0.0226868f $X=3.955 $Y=3.33 $X2=0
+ $Y2=0
cc_264 N_VPWR_c_338_n N_A_507_368#_c_441_n 0.0124868f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_265 N_VPWR_c_342_n N_A_225_74#_c_531_n 0.00464454f $X=4.04 $Y=1.985 $X2=0
+ $Y2=0
cc_266 N_Y_c_400_n N_A_507_368#_M1000_d 0.00395925f $X=3.05 $Y=2.375 $X2=-0.19
+ $Y2=-0.245
cc_267 N_Y_M1003_d N_A_507_368#_c_440_n 0.00226507f $X=2.985 $Y=1.84 $X2=0 $Y2=0
cc_268 N_Y_c_400_n N_A_507_368#_c_440_n 0.00445035f $X=3.05 $Y=2.375 $X2=0 $Y2=0
cc_269 N_Y_c_420_n N_A_507_368#_c_440_n 0.0123811f $X=3.135 $Y=2.46 $X2=0 $Y2=0
cc_270 N_Y_c_400_n N_A_507_368#_c_446_n 0.0123947f $X=3.05 $Y=2.375 $X2=0 $Y2=0
cc_271 N_Y_c_420_n N_A_507_368#_c_446_n 0.0179013f $X=3.135 $Y=2.46 $X2=0 $Y2=0
cc_272 N_Y_c_400_n N_A_507_368#_c_441_n 0.0166041f $X=3.05 $Y=2.375 $X2=0 $Y2=0
cc_273 N_Y_c_420_n N_A_507_368#_c_441_n 0.00683937f $X=3.135 $Y=2.46 $X2=0 $Y2=0
cc_274 N_Y_M1005_s N_A_225_74#_c_526_n 0.00184993f $X=1.56 $Y=0.37 $X2=0 $Y2=0
cc_275 N_Y_c_394_n N_A_225_74#_c_526_n 0.0129924f $X=1.7 $Y=0.8 $X2=0 $Y2=0
cc_276 N_Y_c_394_n N_A_225_74#_c_529_n 0.00932276f $X=1.7 $Y=0.8 $X2=0 $Y2=0
cc_277 N_VGND_c_471_n N_A_225_74#_c_525_n 0.027945f $X=0.71 $Y=0.675 $X2=0 $Y2=0
cc_278 N_VGND_c_472_n N_A_225_74#_c_526_n 0.011924f $X=2.7 $Y=0.675 $X2=0 $Y2=0
cc_279 N_VGND_c_475_n N_A_225_74#_c_526_n 0.0613638f $X=2.535 $Y=0 $X2=0 $Y2=0
cc_280 N_VGND_c_478_n N_A_225_74#_c_526_n 0.034015f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_281 N_VGND_c_471_n N_A_225_74#_c_527_n 0.0121616f $X=0.71 $Y=0.675 $X2=0
+ $Y2=0
cc_282 N_VGND_c_475_n N_A_225_74#_c_527_n 0.0233048f $X=2.535 $Y=0 $X2=0 $Y2=0
cc_283 N_VGND_c_478_n N_A_225_74#_c_527_n 0.0126653f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_284 N_VGND_M1001_s N_A_225_74#_c_528_n 0.00293722f $X=2.49 $Y=0.37 $X2=0
+ $Y2=0
cc_285 N_VGND_c_472_n N_A_225_74#_c_528_n 0.0216414f $X=2.7 $Y=0.675 $X2=0 $Y2=0
cc_286 N_VGND_c_472_n N_A_225_74#_c_530_n 0.00129758f $X=2.7 $Y=0.675 $X2=0
+ $Y2=0
cc_287 N_VGND_c_473_n N_A_225_74#_c_530_n 0.0171736f $X=3.59 $Y=0.645 $X2=0
+ $Y2=0
cc_288 N_VGND_c_476_n N_A_225_74#_c_530_n 0.00749631f $X=3.425 $Y=0 $X2=0 $Y2=0
cc_289 N_VGND_c_478_n N_A_225_74#_c_530_n 0.0062048f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_290 N_VGND_M1008_s N_A_225_74#_c_531_n 0.00176461f $X=3.45 $Y=0.37 $X2=0
+ $Y2=0
cc_291 N_VGND_c_473_n N_A_225_74#_c_531_n 0.0170777f $X=3.59 $Y=0.645 $X2=0
+ $Y2=0
cc_292 N_VGND_c_473_n N_A_225_74#_c_532_n 0.017215f $X=3.59 $Y=0.645 $X2=0 $Y2=0
cc_293 N_VGND_c_477_n N_A_225_74#_c_532_n 0.011066f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_294 N_VGND_c_478_n N_A_225_74#_c_532_n 0.00915947f $X=4.08 $Y=0 $X2=0 $Y2=0
