* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__dfbbp_1 CLK D RESET_B SET_B VGND VNB VPB VPWR Q Q_N
X0 a_422_125# a_214_74# a_520_87# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_422_125# a_27_74# a_520_87# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 VPWR SET_B a_671_93# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X3 a_671_93# a_1062_93# a_872_119# VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X4 a_520_87# a_27_74# a_713_379# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 a_1318_119# a_214_74# a_1311_424# VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X6 a_2320_410# a_1474_446# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 VPWR a_671_93# a_1203_379# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X8 a_1708_74# a_1311_424# a_1474_446# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X9 VGND a_1474_446# Q_N VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X10 a_872_119# a_520_87# a_671_93# VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X11 VGND a_2320_410# Q VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X12 a_520_87# a_214_74# a_606_87# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 a_27_74# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X14 a_1311_424# a_27_74# a_1498_74# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 VPWR a_1474_446# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X16 a_1498_74# a_1474_446# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 a_1062_93# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 a_1311_424# a_214_74# a_1418_508# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X19 a_606_87# a_671_93# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 VGND SET_B a_1708_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X21 VPWR D a_422_125# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X22 VPWR SET_B a_1474_446# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X23 a_713_379# a_671_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X24 a_2320_410# a_1474_446# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X25 VPWR a_2320_410# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X26 VGND a_671_93# a_1318_119# VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X27 VGND SET_B a_872_119# VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X28 a_1062_93# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X29 a_1017_379# a_1062_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X30 a_1814_392# a_1062_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X31 a_27_74# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X32 VGND a_27_74# a_214_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X33 a_1203_379# a_27_74# a_1311_424# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X34 VGND D a_422_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X35 VPWR a_27_74# a_214_74# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X36 a_1418_508# a_1474_446# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X37 a_1474_446# a_1062_93# a_1708_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X38 a_671_93# a_520_87# a_1017_379# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X39 a_1474_446# a_1311_424# a_1814_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends
