* File: sky130_fd_sc_ls__nor2_8.pxi.spice
* Created: Wed Sep  2 11:14:13 2020
* 
x_PM_SKY130_FD_SC_LS__NOR2_8%A N_A_c_142_n N_A_M1000_g N_A_c_130_n N_A_c_131_n
+ N_A_c_145_n N_A_M1005_g N_A_c_132_n N_A_c_147_n N_A_M1013_g N_A_c_133_n
+ N_A_M1004_g N_A_c_149_n N_A_M1016_g N_A_M1007_g N_A_c_150_n N_A_M1017_g
+ N_A_c_151_n N_A_M1019_g N_A_M1012_g N_A_c_152_n N_A_M1021_g N_A_M1015_g
+ N_A_c_153_n N_A_M1023_g N_A_c_138_n N_A_c_139_n A A A A A N_A_c_141_n
+ PM_SKY130_FD_SC_LS__NOR2_8%A
x_PM_SKY130_FD_SC_LS__NOR2_8%B N_B_c_269_n N_B_M1003_g N_B_c_270_n N_B_c_295_n
+ N_B_M1001_g N_B_c_271_n N_B_c_272_n N_B_c_297_n N_B_M1002_g N_B_c_273_n
+ N_B_c_274_n N_B_c_299_n N_B_M1006_g N_B_c_275_n N_B_M1009_g N_B_c_276_n
+ N_B_c_277_n N_B_c_301_n N_B_M1008_g N_B_c_278_n N_B_M1010_g N_B_c_279_n
+ N_B_c_303_n N_B_M1011_g N_B_c_280_n N_B_M1020_g N_B_c_281_n N_B_c_282_n
+ N_B_c_283_n N_B_c_305_n N_B_M1014_g N_B_c_284_n N_B_c_285_n N_B_c_307_n
+ N_B_M1018_g N_B_c_286_n N_B_c_309_n N_B_M1022_g N_B_c_287_n N_B_c_288_n
+ N_B_c_289_n N_B_c_290_n N_B_c_291_n B B N_B_c_292_n N_B_c_293_n
+ PM_SKY130_FD_SC_LS__NOR2_8%B
x_PM_SKY130_FD_SC_LS__NOR2_8%A_27_368# N_A_27_368#_M1000_d N_A_27_368#_M1005_d
+ N_A_27_368#_M1016_d N_A_27_368#_M1019_d N_A_27_368#_M1023_d
+ N_A_27_368#_M1002_d N_A_27_368#_M1008_d N_A_27_368#_M1014_d
+ N_A_27_368#_M1022_d N_A_27_368#_c_423_n N_A_27_368#_c_424_n
+ N_A_27_368#_c_425_n N_A_27_368#_c_426_n N_A_27_368#_c_451_n
+ N_A_27_368#_c_427_n N_A_27_368#_c_460_n N_A_27_368#_c_428_n
+ N_A_27_368#_c_467_n N_A_27_368#_c_471_n N_A_27_368#_c_472_n
+ N_A_27_368#_c_429_n N_A_27_368#_c_430_n N_A_27_368#_c_491_n
+ N_A_27_368#_c_431_n N_A_27_368#_c_432_n N_A_27_368#_c_433_n
+ N_A_27_368#_c_434_n N_A_27_368#_c_435_n N_A_27_368#_c_436_n
+ N_A_27_368#_c_437_n N_A_27_368#_c_478_n N_A_27_368#_c_481_n
+ N_A_27_368#_c_438_n N_A_27_368#_c_439_n N_A_27_368#_c_440_n
+ PM_SKY130_FD_SC_LS__NOR2_8%A_27_368#
x_PM_SKY130_FD_SC_LS__NOR2_8%VPWR N_VPWR_M1000_s N_VPWR_M1013_s N_VPWR_M1017_s
+ N_VPWR_M1021_s N_VPWR_c_563_n N_VPWR_c_564_n N_VPWR_c_565_n N_VPWR_c_566_n
+ VPWR N_VPWR_c_567_n N_VPWR_c_568_n N_VPWR_c_569_n N_VPWR_c_570_n
+ N_VPWR_c_571_n N_VPWR_c_562_n N_VPWR_c_573_n N_VPWR_c_574_n N_VPWR_c_575_n
+ N_VPWR_c_576_n PM_SKY130_FD_SC_LS__NOR2_8%VPWR
x_PM_SKY130_FD_SC_LS__NOR2_8%Y N_Y_M1004_s N_Y_M1012_s N_Y_M1003_s N_Y_M1010_s
+ N_Y_M1001_s N_Y_M1006_s N_Y_M1011_s N_Y_M1018_s N_Y_c_661_n N_Y_c_662_n
+ N_Y_c_663_n N_Y_c_664_n N_Y_c_665_n N_Y_c_670_n N_Y_c_694_n N_Y_c_666_n
+ N_Y_c_701_n N_Y_c_667_n N_Y_c_668_n N_Y_c_736_n N_Y_c_669_n Y Y
+ PM_SKY130_FD_SC_LS__NOR2_8%Y
x_PM_SKY130_FD_SC_LS__NOR2_8%VGND N_VGND_M1004_d N_VGND_M1007_d N_VGND_M1015_d
+ N_VGND_M1009_d N_VGND_M1020_d N_VGND_c_781_n N_VGND_c_782_n N_VGND_c_783_n
+ N_VGND_c_784_n N_VGND_c_785_n N_VGND_c_786_n N_VGND_c_787_n VGND
+ N_VGND_c_788_n N_VGND_c_789_n N_VGND_c_790_n N_VGND_c_791_n N_VGND_c_792_n
+ N_VGND_c_793_n N_VGND_c_794_n N_VGND_c_795_n N_VGND_c_796_n
+ PM_SKY130_FD_SC_LS__NOR2_8%VGND
cc_1 VNB N_A_c_130_n 0.0125911f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=1.65
cc_2 VNB N_A_c_131_n 0.0160597f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.65
cc_3 VNB N_A_c_132_n 0.00968592f $X=-0.19 $Y=-0.245 $X2=1.365 $Y2=1.65
cc_4 VNB N_A_c_133_n 0.00705127f $X=-0.19 $Y=-0.245 $X2=1.735 $Y2=1.65
cc_5 VNB N_A_M1004_g 0.0315514f $X=-0.19 $Y=-0.245 $X2=1.81 $Y2=0.74
cc_6 VNB N_A_M1007_g 0.0315587f $X=-0.19 $Y=-0.245 $X2=2.31 $Y2=0.74
cc_7 VNB N_A_M1012_g 0.0307539f $X=-0.19 $Y=-0.245 $X2=3.21 $Y2=0.74
cc_8 VNB N_A_M1015_g 0.0247574f $X=-0.19 $Y=-0.245 $X2=3.71 $Y2=0.74
cc_9 VNB N_A_c_138_n 0.00723254f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.67
cc_10 VNB N_A_c_139_n 0.00723254f $X=-0.19 $Y=-0.245 $X2=1.455 $Y2=1.67
cc_11 VNB A 0.012161f $X=-0.19 $Y=-0.245 $X2=3.515 $Y2=1.58
cc_12 VNB N_A_c_141_n 0.110096f $X=-0.19 $Y=-0.245 $X2=3.71 $Y2=1.557
cc_13 VNB N_B_c_269_n 0.0200058f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_14 VNB N_B_c_270_n 0.0196625f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.65
cc_15 VNB N_B_c_271_n 0.0181613f $X=-0.19 $Y=-0.245 $X2=1.365 $Y2=1.65
cc_16 VNB N_B_c_272_n 0.0158298f $X=-0.19 $Y=-0.245 $X2=1.455 $Y2=2.4
cc_17 VNB N_B_c_273_n 0.0166202f $X=-0.19 $Y=-0.245 $X2=1.81 $Y2=1.35
cc_18 VNB N_B_c_274_n 0.015177f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_B_c_275_n 0.020416f $X=-0.19 $Y=-0.245 $X2=2.31 $Y2=1.35
cc_20 VNB N_B_c_276_n 0.0117381f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_B_c_277_n 0.0145655f $X=-0.19 $Y=-0.245 $X2=2.355 $Y2=2.4
cc_22 VNB N_B_c_278_n 0.0157738f $X=-0.19 $Y=-0.245 $X2=3.21 $Y2=1.35
cc_23 VNB N_B_c_279_n 0.015156f $X=-0.19 $Y=-0.245 $X2=3.305 $Y2=1.765
cc_24 VNB N_B_c_280_n 0.0169231f $X=-0.19 $Y=-0.245 $X2=3.71 $Y2=0.74
cc_25 VNB N_B_c_281_n 0.00635223f $X=-0.19 $Y=-0.245 $X2=3.855 $Y2=1.765
cc_26 VNB N_B_c_282_n 0.0193657f $X=-0.19 $Y=-0.245 $X2=3.855 $Y2=2.4
cc_27 VNB N_B_c_283_n 0.0163843f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.67
cc_28 VNB N_B_c_284_n 0.0188047f $X=-0.19 $Y=-0.245 $X2=2.555 $Y2=1.58
cc_29 VNB N_B_c_285_n 0.0164034f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_B_c_286_n 0.0264902f $X=-0.19 $Y=-0.245 $X2=1.81 $Y2=1.557
cc_31 VNB N_B_c_287_n 0.0109819f $X=-0.19 $Y=-0.245 $X2=2.06 $Y2=1.515
cc_32 VNB N_B_c_288_n 0.00800291f $X=-0.19 $Y=-0.245 $X2=2.31 $Y2=1.557
cc_33 VNB N_B_c_289_n 0.00294508f $X=-0.19 $Y=-0.245 $X2=2.355 $Y2=1.557
cc_34 VNB N_B_c_290_n 0.00734323f $X=-0.19 $Y=-0.245 $X2=3.42 $Y2=1.515
cc_35 VNB N_B_c_291_n 0.0206427f $X=-0.19 $Y=-0.245 $X2=3.71 $Y2=1.557
cc_36 VNB N_B_c_292_n 0.150322f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_B_c_293_n 0.00258269f $X=-0.19 $Y=-0.245 $X2=2.64 $Y2=1.565
cc_38 VNB N_VPWR_c_562_n 0.342803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_Y_c_661_n 0.00280455f $X=-0.19 $Y=-0.245 $X2=2.355 $Y2=1.765
cc_40 VNB N_Y_c_662_n 0.00636217f $X=-0.19 $Y=-0.245 $X2=2.355 $Y2=2.4
cc_41 VNB N_Y_c_663_n 0.00231148f $X=-0.19 $Y=-0.245 $X2=2.855 $Y2=1.765
cc_42 VNB N_Y_c_664_n 0.00280455f $X=-0.19 $Y=-0.245 $X2=3.21 $Y2=1.35
cc_43 VNB N_Y_c_665_n 0.00879444f $X=-0.19 $Y=-0.245 $X2=3.21 $Y2=0.74
cc_44 VNB N_Y_c_666_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=2.555 $Y2=1.58
cc_45 VNB N_Y_c_667_n 0.0135921f $X=-0.19 $Y=-0.245 $X2=1.81 $Y2=1.557
cc_46 VNB N_Y_c_668_n 0.0298908f $X=-0.19 $Y=-0.245 $X2=1.905 $Y2=1.557
cc_47 VNB N_Y_c_669_n 0.00231148f $X=-0.19 $Y=-0.245 $X2=3.21 $Y2=1.557
cc_48 VNB N_VGND_c_781_n 0.065313f $X=-0.19 $Y=-0.245 $X2=1.905 $Y2=1.765
cc_49 VNB N_VGND_c_782_n 0.00936836f $X=-0.19 $Y=-0.245 $X2=2.31 $Y2=0.74
cc_50 VNB N_VGND_c_783_n 0.00585698f $X=-0.19 $Y=-0.245 $X2=2.355 $Y2=2.4
cc_51 VNB N_VGND_c_784_n 0.0351261f $X=-0.19 $Y=-0.245 $X2=2.855 $Y2=2.4
cc_52 VNB N_VGND_c_785_n 0.00899973f $X=-0.19 $Y=-0.245 $X2=3.21 $Y2=0.74
cc_53 VNB N_VGND_c_786_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=3.305 $Y2=1.765
cc_54 VNB N_VGND_c_787_n 0.0211799f $X=-0.19 $Y=-0.245 $X2=3.71 $Y2=0.74
cc_55 VNB N_VGND_c_788_n 0.0185368f $X=-0.19 $Y=-0.245 $X2=3.855 $Y2=2.4
cc_56 VNB N_VGND_c_789_n 0.0185368f $X=-0.19 $Y=-0.245 $X2=2.075 $Y2=1.58
cc_57 VNB N_VGND_c_790_n 0.0433909f $X=-0.19 $Y=-0.245 $X2=1.905 $Y2=1.557
cc_58 VNB N_VGND_c_791_n 0.474712f $X=-0.19 $Y=-0.245 $X2=2.06 $Y2=1.557
cc_59 VNB N_VGND_c_792_n 0.0428317f $X=-0.19 $Y=-0.245 $X2=2.31 $Y2=1.557
cc_60 VNB N_VGND_c_793_n 0.0138518f $X=-0.19 $Y=-0.245 $X2=3.42 $Y2=1.557
cc_61 VNB N_VGND_c_794_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=3.71 $Y2=1.557
cc_62 VNB N_VGND_c_795_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_796_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=2.16 $Y2=1.565
cc_64 VPB N_A_c_142_n 0.0201143f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_65 VPB N_A_c_130_n 0.00895896f $X=-0.19 $Y=1.66 $X2=0.915 $Y2=1.65
cc_66 VPB N_A_c_131_n 0.00893071f $X=-0.19 $Y=1.66 $X2=0.595 $Y2=1.65
cc_67 VPB N_A_c_145_n 0.0149072f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.765
cc_68 VPB N_A_c_132_n 0.00759523f $X=-0.19 $Y=1.66 $X2=1.365 $Y2=1.65
cc_69 VPB N_A_c_147_n 0.0150613f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=1.765
cc_70 VPB N_A_c_133_n 0.00657536f $X=-0.19 $Y=1.66 $X2=1.735 $Y2=1.65
cc_71 VPB N_A_c_149_n 0.0149599f $X=-0.19 $Y=1.66 $X2=1.905 $Y2=1.765
cc_72 VPB N_A_c_150_n 0.0158869f $X=-0.19 $Y=1.66 $X2=2.355 $Y2=1.765
cc_73 VPB N_A_c_151_n 0.0153815f $X=-0.19 $Y=1.66 $X2=2.855 $Y2=1.765
cc_74 VPB N_A_c_152_n 0.0162352f $X=-0.19 $Y=1.66 $X2=3.305 $Y2=1.765
cc_75 VPB N_A_c_153_n 0.0160915f $X=-0.19 $Y=1.66 $X2=3.855 $Y2=1.765
cc_76 VPB N_A_c_138_n 0.00409953f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.67
cc_77 VPB N_A_c_139_n 0.00404919f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=1.67
cc_78 VPB A 0.0156195f $X=-0.19 $Y=1.66 $X2=3.515 $Y2=1.58
cc_79 VPB N_A_c_141_n 0.0678482f $X=-0.19 $Y=1.66 $X2=3.71 $Y2=1.557
cc_80 VPB N_B_c_270_n 7.92394e-19 $X=-0.19 $Y=1.66 $X2=0.595 $Y2=1.65
cc_81 VPB N_B_c_295_n 0.0215615f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.765
cc_82 VPB N_B_c_272_n 6.84003e-19 $X=-0.19 $Y=1.66 $X2=1.455 $Y2=2.4
cc_83 VPB N_B_c_297_n 0.020382f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=2.4
cc_84 VPB N_B_c_274_n 6.55797e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_B_c_299_n 0.0198258f $X=-0.19 $Y=1.66 $X2=1.905 $Y2=1.765
cc_86 VPB N_B_c_277_n 6.85396e-19 $X=-0.19 $Y=1.66 $X2=2.355 $Y2=2.4
cc_87 VPB N_B_c_301_n 0.0200857f $X=-0.19 $Y=1.66 $X2=2.855 $Y2=1.765
cc_88 VPB N_B_c_279_n 6.8539e-19 $X=-0.19 $Y=1.66 $X2=3.305 $Y2=1.765
cc_89 VPB N_B_c_303_n 0.0200814f $X=-0.19 $Y=1.66 $X2=3.305 $Y2=2.4
cc_90 VPB N_B_c_283_n 7.13681e-19 $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.67
cc_91 VPB N_B_c_305_n 0.0206453f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=1.67
cc_92 VPB N_B_c_285_n 7.13681e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_B_c_307_n 0.0206632f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB N_B_c_286_n 0.00111912f $X=-0.19 $Y=1.66 $X2=1.81 $Y2=1.557
cc_95 VPB N_B_c_309_n 0.0265697f $X=-0.19 $Y=1.66 $X2=1.905 $Y2=1.557
cc_96 VPB N_A_27_368#_c_423_n 0.0418511f $X=-0.19 $Y=1.66 $X2=2.855 $Y2=1.765
cc_97 VPB N_A_27_368#_c_424_n 0.00399078f $X=-0.19 $Y=1.66 $X2=3.21 $Y2=0.74
cc_98 VPB N_A_27_368#_c_425_n 0.0196833f $X=-0.19 $Y=1.66 $X2=3.21 $Y2=0.74
cc_99 VPB N_A_27_368#_c_426_n 0.00180921f $X=-0.19 $Y=1.66 $X2=3.305 $Y2=2.4
cc_100 VPB N_A_27_368#_c_427_n 0.00216998f $X=-0.19 $Y=1.66 $X2=3.855 $Y2=1.765
cc_101 VPB N_A_27_368#_c_428_n 0.00216998f $X=-0.19 $Y=1.66 $X2=2.075 $Y2=1.58
cc_102 VPB N_A_27_368#_c_429_n 0.00280532f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 VPB N_A_27_368#_c_430_n 0.0021839f $X=-0.19 $Y=1.66 $X2=1.81 $Y2=1.557
cc_104 VPB N_A_27_368#_c_431_n 0.0027626f $X=-0.19 $Y=1.66 $X2=2.855 $Y2=1.557
cc_105 VPB N_A_27_368#_c_432_n 0.00201157f $X=-0.19 $Y=1.66 $X2=3.42 $Y2=1.515
cc_106 VPB N_A_27_368#_c_433_n 0.0027982f $X=-0.19 $Y=1.66 $X2=1.68 $Y2=1.565
cc_107 VPB N_A_27_368#_c_434_n 0.00245482f $X=-0.19 $Y=1.66 $X2=2.16 $Y2=1.565
cc_108 VPB N_A_27_368#_c_435_n 0.0128449f $X=-0.19 $Y=1.66 $X2=3.12 $Y2=1.565
cc_109 VPB N_A_27_368#_c_436_n 0.0548523f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_110 VPB N_A_27_368#_c_437_n 0.00228583f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_A_27_368#_c_438_n 0.00189272f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_A_27_368#_c_439_n 0.00149233f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_A_27_368#_c_440_n 0.00189272f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_VPWR_c_563_n 0.00584464f $X=-0.19 $Y=1.66 $X2=1.545 $Y2=1.65
cc_115 VPB N_VPWR_c_564_n 0.0026822f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_VPWR_c_565_n 0.00511574f $X=-0.19 $Y=1.66 $X2=2.31 $Y2=1.35
cc_117 VPB N_VPWR_c_566_n 0.00849451f $X=-0.19 $Y=1.66 $X2=2.355 $Y2=1.765
cc_118 VPB N_VPWR_c_567_n 0.0191515f $X=-0.19 $Y=1.66 $X2=2.855 $Y2=2.4
cc_119 VPB N_VPWR_c_568_n 0.0164465f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_569_n 0.0175706f $X=-0.19 $Y=1.66 $X2=3.71 $Y2=0.74
cc_121 VPB N_VPWR_c_570_n 0.0175706f $X=-0.19 $Y=1.66 $X2=3.855 $Y2=2.4
cc_122 VPB N_VPWR_c_571_n 0.102588f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_562_n 0.0902801f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_573_n 0.00614127f $X=-0.19 $Y=1.66 $X2=1.905 $Y2=1.557
cc_125 VPB N_VPWR_c_574_n 0.00601644f $X=-0.19 $Y=1.66 $X2=2.06 $Y2=1.515
cc_126 VPB N_VPWR_c_575_n 0.00614127f $X=-0.19 $Y=1.66 $X2=2.855 $Y2=1.557
cc_127 VPB N_VPWR_c_576_n 0.00631788f $X=-0.19 $Y=1.66 $X2=3.42 $Y2=1.557
cc_128 VPB N_Y_c_670_n 8.08642e-19 $X=-0.19 $Y=1.66 $X2=3.305 $Y2=2.4
cc_129 VPB N_Y_c_668_n 0.00797804f $X=-0.19 $Y=1.66 $X2=1.905 $Y2=1.557
cc_130 N_A_M1015_g N_B_c_269_n 0.0286926f $X=3.71 $Y=0.74 $X2=-0.19 $Y2=-0.245
cc_131 N_A_M1015_g N_B_c_270_n 0.00677313f $X=3.71 $Y=0.74 $X2=0 $Y2=0
cc_132 A N_B_c_270_n 0.00174415f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_133 N_A_c_141_n N_B_c_270_n 0.00932947f $X=3.71 $Y=1.557 $X2=0 $Y2=0
cc_134 N_A_c_153_n N_B_c_295_n 0.00894277f $X=3.855 $Y=1.765 $X2=0 $Y2=0
cc_135 N_A_c_142_n N_A_27_368#_c_423_n 0.0128821f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_136 N_A_c_145_n N_A_27_368#_c_423_n 9.88307e-19 $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_137 N_A_c_142_n N_A_27_368#_c_424_n 0.0156179f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_138 N_A_c_130_n N_A_27_368#_c_424_n 0.00946668f $X=0.915 $Y=1.65 $X2=0 $Y2=0
cc_139 N_A_c_131_n N_A_27_368#_c_424_n 6.25096e-19 $X=0.595 $Y=1.65 $X2=0 $Y2=0
cc_140 N_A_c_145_n N_A_27_368#_c_424_n 0.014467f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_141 N_A_c_132_n N_A_27_368#_c_424_n 0.00136939f $X=1.365 $Y=1.65 $X2=0 $Y2=0
cc_142 N_A_c_138_n N_A_27_368#_c_424_n 9.13093e-19 $X=1.005 $Y=1.67 $X2=0 $Y2=0
cc_143 N_A_c_142_n N_A_27_368#_c_425_n 0.00211856f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_144 N_A_c_131_n N_A_27_368#_c_425_n 7.47253e-19 $X=0.595 $Y=1.65 $X2=0 $Y2=0
cc_145 N_A_c_132_n N_A_27_368#_c_451_n 9.11152e-19 $X=1.365 $Y=1.65 $X2=0 $Y2=0
cc_146 N_A_c_147_n N_A_27_368#_c_451_n 0.0167176f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_147 N_A_c_133_n N_A_27_368#_c_451_n 0.00139628f $X=1.735 $Y=1.65 $X2=0 $Y2=0
cc_148 N_A_c_149_n N_A_27_368#_c_451_n 0.0125795f $X=1.905 $Y=1.765 $X2=0 $Y2=0
cc_149 A N_A_27_368#_c_451_n 0.0322199f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_150 N_A_c_141_n N_A_27_368#_c_451_n 2.1846e-19 $X=3.71 $Y=1.557 $X2=0 $Y2=0
cc_151 N_A_c_149_n N_A_27_368#_c_427_n 0.00610108f $X=1.905 $Y=1.765 $X2=0 $Y2=0
cc_152 N_A_c_150_n N_A_27_368#_c_427_n 0.0100427f $X=2.355 $Y=1.765 $X2=0 $Y2=0
cc_153 N_A_c_151_n N_A_27_368#_c_427_n 8.89687e-19 $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_154 N_A_c_150_n N_A_27_368#_c_460_n 0.0122806f $X=2.355 $Y=1.765 $X2=0 $Y2=0
cc_155 N_A_c_151_n N_A_27_368#_c_460_n 0.0129585f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_156 A N_A_27_368#_c_460_n 0.0475353f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_157 N_A_c_141_n N_A_27_368#_c_460_n 0.00199109f $X=3.71 $Y=1.557 $X2=0 $Y2=0
cc_158 N_A_c_151_n N_A_27_368#_c_428_n 0.00610108f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_159 N_A_c_152_n N_A_27_368#_c_428_n 0.0103558f $X=3.305 $Y=1.765 $X2=0 $Y2=0
cc_160 N_A_c_153_n N_A_27_368#_c_428_n 6.65337e-19 $X=3.855 $Y=1.765 $X2=0 $Y2=0
cc_161 N_A_c_152_n N_A_27_368#_c_467_n 0.0125195f $X=3.305 $Y=1.765 $X2=0 $Y2=0
cc_162 N_A_c_153_n N_A_27_368#_c_467_n 0.0161633f $X=3.855 $Y=1.765 $X2=0 $Y2=0
cc_163 A N_A_27_368#_c_467_n 0.034429f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_164 N_A_c_141_n N_A_27_368#_c_467_n 0.00311572f $X=3.71 $Y=1.557 $X2=0 $Y2=0
cc_165 N_A_c_153_n N_A_27_368#_c_471_n 8.9215e-19 $X=3.855 $Y=1.765 $X2=0 $Y2=0
cc_166 N_A_c_152_n N_A_27_368#_c_472_n 6.4805e-19 $X=3.305 $Y=1.765 $X2=0 $Y2=0
cc_167 N_A_c_153_n N_A_27_368#_c_472_n 0.00932822f $X=3.855 $Y=1.765 $X2=0 $Y2=0
cc_168 N_A_c_153_n N_A_27_368#_c_430_n 0.00313312f $X=3.855 $Y=1.765 $X2=0 $Y2=0
cc_169 N_A_c_145_n N_A_27_368#_c_437_n 0.00628092f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_170 N_A_c_132_n N_A_27_368#_c_437_n 0.00524054f $X=1.365 $Y=1.65 $X2=0 $Y2=0
cc_171 N_A_c_147_n N_A_27_368#_c_437_n 0.00920037f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_172 N_A_c_150_n N_A_27_368#_c_478_n 4.27055e-19 $X=2.355 $Y=1.765 $X2=0 $Y2=0
cc_173 A N_A_27_368#_c_478_n 0.0193936f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_174 N_A_c_141_n N_A_27_368#_c_478_n 0.0013819f $X=3.71 $Y=1.557 $X2=0 $Y2=0
cc_175 N_A_c_152_n N_A_27_368#_c_481_n 4.27055e-19 $X=3.305 $Y=1.765 $X2=0 $Y2=0
cc_176 A N_A_27_368#_c_481_n 0.0193936f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_177 N_A_c_141_n N_A_27_368#_c_481_n 0.00137857f $X=3.71 $Y=1.557 $X2=0 $Y2=0
cc_178 N_A_c_142_n N_VPWR_c_563_n 0.00777421f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_179 N_A_c_145_n N_VPWR_c_563_n 0.014403f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_180 N_A_c_147_n N_VPWR_c_563_n 5.87661e-19 $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_181 N_A_c_145_n N_VPWR_c_564_n 5.35985e-19 $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_182 N_A_c_147_n N_VPWR_c_564_n 0.0110266f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_183 N_A_c_149_n N_VPWR_c_564_n 0.0111104f $X=1.905 $Y=1.765 $X2=0 $Y2=0
cc_184 N_A_c_150_n N_VPWR_c_564_n 5.51351e-19 $X=2.355 $Y=1.765 $X2=0 $Y2=0
cc_185 N_A_c_150_n N_VPWR_c_565_n 0.00541712f $X=2.355 $Y=1.765 $X2=0 $Y2=0
cc_186 N_A_c_151_n N_VPWR_c_565_n 0.011046f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_187 N_A_c_152_n N_VPWR_c_565_n 5.51351e-19 $X=3.305 $Y=1.765 $X2=0 $Y2=0
cc_188 N_A_c_152_n N_VPWR_c_566_n 0.00592199f $X=3.305 $Y=1.765 $X2=0 $Y2=0
cc_189 N_A_c_153_n N_VPWR_c_566_n 0.00546951f $X=3.855 $Y=1.765 $X2=0 $Y2=0
cc_190 N_A_c_142_n N_VPWR_c_567_n 0.00445602f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_191 N_A_c_145_n N_VPWR_c_568_n 0.00413917f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_192 N_A_c_147_n N_VPWR_c_568_n 0.00413917f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_193 N_A_c_149_n N_VPWR_c_569_n 0.00413917f $X=1.905 $Y=1.765 $X2=0 $Y2=0
cc_194 N_A_c_150_n N_VPWR_c_569_n 0.00445602f $X=2.355 $Y=1.765 $X2=0 $Y2=0
cc_195 N_A_c_151_n N_VPWR_c_570_n 0.00413917f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_196 N_A_c_152_n N_VPWR_c_570_n 0.00445602f $X=3.305 $Y=1.765 $X2=0 $Y2=0
cc_197 N_A_c_153_n N_VPWR_c_571_n 0.0044313f $X=3.855 $Y=1.765 $X2=0 $Y2=0
cc_198 N_A_c_142_n N_VPWR_c_562_n 0.00860873f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_199 N_A_c_145_n N_VPWR_c_562_n 0.00817726f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_200 N_A_c_147_n N_VPWR_c_562_n 0.00817726f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_201 N_A_c_149_n N_VPWR_c_562_n 0.00817726f $X=1.905 $Y=1.765 $X2=0 $Y2=0
cc_202 N_A_c_150_n N_VPWR_c_562_n 0.00857378f $X=2.355 $Y=1.765 $X2=0 $Y2=0
cc_203 N_A_c_151_n N_VPWR_c_562_n 0.00817726f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_204 N_A_c_152_n N_VPWR_c_562_n 0.00857797f $X=3.305 $Y=1.765 $X2=0 $Y2=0
cc_205 N_A_c_153_n N_VPWR_c_562_n 0.00853652f $X=3.855 $Y=1.765 $X2=0 $Y2=0
cc_206 N_A_M1004_g N_Y_c_661_n 0.00821243f $X=1.81 $Y=0.74 $X2=0 $Y2=0
cc_207 N_A_M1007_g N_Y_c_661_n 0.00350341f $X=2.31 $Y=0.74 $X2=0 $Y2=0
cc_208 N_A_M1007_g N_Y_c_662_n 0.0167736f $X=2.31 $Y=0.74 $X2=0 $Y2=0
cc_209 N_A_M1012_g N_Y_c_662_n 0.0131906f $X=3.21 $Y=0.74 $X2=0 $Y2=0
cc_210 A N_Y_c_662_n 0.0809793f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_211 N_A_c_141_n N_Y_c_662_n 0.0136367f $X=3.71 $Y=1.557 $X2=0 $Y2=0
cc_212 N_A_M1004_g N_Y_c_663_n 0.00499186f $X=1.81 $Y=0.74 $X2=0 $Y2=0
cc_213 A N_Y_c_663_n 0.0282341f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_214 N_A_c_141_n N_Y_c_663_n 0.00408616f $X=3.71 $Y=1.557 $X2=0 $Y2=0
cc_215 N_A_M1012_g N_Y_c_664_n 0.0137366f $X=3.21 $Y=0.74 $X2=0 $Y2=0
cc_216 N_A_M1015_g N_Y_c_664_n 0.00350341f $X=3.71 $Y=0.74 $X2=0 $Y2=0
cc_217 N_A_M1015_g N_Y_c_665_n 0.0169005f $X=3.71 $Y=0.74 $X2=0 $Y2=0
cc_218 A N_Y_c_665_n 0.00925196f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_219 N_A_c_141_n N_Y_c_665_n 0.00515795f $X=3.71 $Y=1.557 $X2=0 $Y2=0
cc_220 N_A_M1015_g N_Y_c_668_n 0.00133266f $X=3.71 $Y=0.74 $X2=0 $Y2=0
cc_221 N_A_M1012_g N_Y_c_669_n 0.00173883f $X=3.21 $Y=0.74 $X2=0 $Y2=0
cc_222 A N_Y_c_669_n 0.0282341f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_223 N_A_c_141_n N_Y_c_669_n 0.00408616f $X=3.71 $Y=1.557 $X2=0 $Y2=0
cc_224 N_A_c_130_n N_VGND_c_781_n 0.0217371f $X=0.915 $Y=1.65 $X2=0 $Y2=0
cc_225 N_A_c_133_n N_VGND_c_781_n 6.06424e-19 $X=1.735 $Y=1.65 $X2=0 $Y2=0
cc_226 N_A_M1004_g N_VGND_c_781_n 0.00556557f $X=1.81 $Y=0.74 $X2=0 $Y2=0
cc_227 A N_VGND_c_781_n 0.00932589f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_228 N_A_M1004_g N_VGND_c_782_n 4.95933e-19 $X=1.81 $Y=0.74 $X2=0 $Y2=0
cc_229 N_A_M1007_g N_VGND_c_782_n 0.0137423f $X=2.31 $Y=0.74 $X2=0 $Y2=0
cc_230 N_A_M1012_g N_VGND_c_782_n 0.00607183f $X=3.21 $Y=0.74 $X2=0 $Y2=0
cc_231 N_A_M1012_g N_VGND_c_783_n 4.99121e-19 $X=3.21 $Y=0.74 $X2=0 $Y2=0
cc_232 N_A_M1015_g N_VGND_c_783_n 0.0109084f $X=3.71 $Y=0.74 $X2=0 $Y2=0
cc_233 N_A_M1004_g N_VGND_c_788_n 0.00434272f $X=1.81 $Y=0.74 $X2=0 $Y2=0
cc_234 N_A_M1007_g N_VGND_c_788_n 0.00383152f $X=2.31 $Y=0.74 $X2=0 $Y2=0
cc_235 N_A_M1012_g N_VGND_c_789_n 0.00434272f $X=3.21 $Y=0.74 $X2=0 $Y2=0
cc_236 N_A_M1015_g N_VGND_c_789_n 0.00383152f $X=3.71 $Y=0.74 $X2=0 $Y2=0
cc_237 N_A_M1004_g N_VGND_c_791_n 0.00825717f $X=1.81 $Y=0.74 $X2=0 $Y2=0
cc_238 N_A_M1007_g N_VGND_c_791_n 0.00758198f $X=2.31 $Y=0.74 $X2=0 $Y2=0
cc_239 N_A_M1012_g N_VGND_c_791_n 0.00825717f $X=3.21 $Y=0.74 $X2=0 $Y2=0
cc_240 N_A_M1015_g N_VGND_c_791_n 0.00758198f $X=3.71 $Y=0.74 $X2=0 $Y2=0
cc_241 N_B_c_295_n N_A_27_368#_c_471_n 0.00235486f $X=4.305 $Y=1.765 $X2=0 $Y2=0
cc_242 N_B_c_287_n N_A_27_368#_c_471_n 0.00179981f $X=4.265 $Y=1.26 $X2=0 $Y2=0
cc_243 N_B_c_295_n N_A_27_368#_c_472_n 0.0091139f $X=4.305 $Y=1.765 $X2=0 $Y2=0
cc_244 N_B_c_297_n N_A_27_368#_c_472_n 5.33746e-19 $X=4.805 $Y=1.765 $X2=0 $Y2=0
cc_245 N_B_c_295_n N_A_27_368#_c_429_n 0.0111147f $X=4.305 $Y=1.765 $X2=0 $Y2=0
cc_246 N_B_c_297_n N_A_27_368#_c_429_n 0.014127f $X=4.805 $Y=1.765 $X2=0 $Y2=0
cc_247 N_B_c_295_n N_A_27_368#_c_430_n 0.00171731f $X=4.305 $Y=1.765 $X2=0 $Y2=0
cc_248 N_B_c_273_n N_A_27_368#_c_491_n 4.59311e-19 $X=5.215 $Y=1.26 $X2=0 $Y2=0
cc_249 N_B_c_299_n N_A_27_368#_c_431_n 0.0130187f $X=5.305 $Y=1.765 $X2=0 $Y2=0
cc_250 N_B_c_301_n N_A_27_368#_c_431_n 0.0127907f $X=5.755 $Y=1.765 $X2=0 $Y2=0
cc_251 N_B_c_301_n N_A_27_368#_c_432_n 3.7884e-19 $X=5.755 $Y=1.765 $X2=0 $Y2=0
cc_252 N_B_c_303_n N_A_27_368#_c_432_n 3.76405e-19 $X=6.205 $Y=1.765 $X2=0 $Y2=0
cc_253 N_B_c_282_n N_A_27_368#_c_432_n 3.5899e-19 $X=6.4 $Y=1.26 $X2=0 $Y2=0
cc_254 N_B_c_303_n N_A_27_368#_c_433_n 0.0128349f $X=6.205 $Y=1.765 $X2=0 $Y2=0
cc_255 N_B_c_305_n N_A_27_368#_c_433_n 0.0138537f $X=6.655 $Y=1.765 $X2=0 $Y2=0
cc_256 N_B_c_305_n N_A_27_368#_c_434_n 0.00571878f $X=6.655 $Y=1.765 $X2=0 $Y2=0
cc_257 N_B_c_307_n N_A_27_368#_c_434_n 4.27567e-19 $X=7.155 $Y=1.765 $X2=0 $Y2=0
cc_258 N_B_c_307_n N_A_27_368#_c_435_n 0.0130187f $X=7.155 $Y=1.765 $X2=0 $Y2=0
cc_259 N_B_c_309_n N_A_27_368#_c_435_n 0.014991f $X=7.605 $Y=1.765 $X2=0 $Y2=0
cc_260 N_B_c_309_n N_A_27_368#_c_436_n 0.0213106f $X=7.605 $Y=1.765 $X2=0 $Y2=0
cc_261 N_B_c_295_n N_VPWR_c_571_n 0.00278257f $X=4.305 $Y=1.765 $X2=0 $Y2=0
cc_262 N_B_c_297_n N_VPWR_c_571_n 0.00278271f $X=4.805 $Y=1.765 $X2=0 $Y2=0
cc_263 N_B_c_299_n N_VPWR_c_571_n 0.00278271f $X=5.305 $Y=1.765 $X2=0 $Y2=0
cc_264 N_B_c_301_n N_VPWR_c_571_n 0.00278271f $X=5.755 $Y=1.765 $X2=0 $Y2=0
cc_265 N_B_c_303_n N_VPWR_c_571_n 0.00278271f $X=6.205 $Y=1.765 $X2=0 $Y2=0
cc_266 N_B_c_305_n N_VPWR_c_571_n 0.00278271f $X=6.655 $Y=1.765 $X2=0 $Y2=0
cc_267 N_B_c_307_n N_VPWR_c_571_n 0.00278271f $X=7.155 $Y=1.765 $X2=0 $Y2=0
cc_268 N_B_c_309_n N_VPWR_c_571_n 0.00278271f $X=7.605 $Y=1.765 $X2=0 $Y2=0
cc_269 N_B_c_295_n N_VPWR_c_562_n 0.00354366f $X=4.305 $Y=1.765 $X2=0 $Y2=0
cc_270 N_B_c_297_n N_VPWR_c_562_n 0.00354745f $X=4.805 $Y=1.765 $X2=0 $Y2=0
cc_271 N_B_c_299_n N_VPWR_c_562_n 0.00354284f $X=5.305 $Y=1.765 $X2=0 $Y2=0
cc_272 N_B_c_301_n N_VPWR_c_562_n 0.00353823f $X=5.755 $Y=1.765 $X2=0 $Y2=0
cc_273 N_B_c_303_n N_VPWR_c_562_n 0.00353823f $X=6.205 $Y=1.765 $X2=0 $Y2=0
cc_274 N_B_c_305_n N_VPWR_c_562_n 0.00354284f $X=6.655 $Y=1.765 $X2=0 $Y2=0
cc_275 N_B_c_307_n N_VPWR_c_562_n 0.00354284f $X=7.155 $Y=1.765 $X2=0 $Y2=0
cc_276 N_B_c_309_n N_VPWR_c_562_n 0.00357472f $X=7.605 $Y=1.765 $X2=0 $Y2=0
cc_277 N_B_c_269_n N_Y_c_665_n 0.0147808f $X=4.21 $Y=1.185 $X2=0 $Y2=0
cc_278 N_B_c_295_n N_Y_c_670_n 0.00643948f $X=4.305 $Y=1.765 $X2=0 $Y2=0
cc_279 N_B_c_297_n N_Y_c_670_n 0.0117002f $X=4.805 $Y=1.765 $X2=0 $Y2=0
cc_280 N_B_c_299_n N_Y_c_670_n 6.36423e-19 $X=5.305 $Y=1.765 $X2=0 $Y2=0
cc_281 N_B_c_297_n N_Y_c_694_n 7.05539e-19 $X=4.805 $Y=1.765 $X2=0 $Y2=0
cc_282 N_B_c_299_n N_Y_c_694_n 0.0117292f $X=5.305 $Y=1.765 $X2=0 $Y2=0
cc_283 N_B_c_301_n N_Y_c_694_n 0.0104688f $X=5.755 $Y=1.765 $X2=0 $Y2=0
cc_284 N_B_c_303_n N_Y_c_694_n 3.69512e-19 $X=6.205 $Y=1.765 $X2=0 $Y2=0
cc_285 N_B_c_275_n N_Y_c_666_n 6.54586e-19 $X=5.325 $Y=1.185 $X2=0 $Y2=0
cc_286 N_B_c_278_n N_Y_c_666_n 0.0113581f $X=5.895 $Y=1.185 $X2=0 $Y2=0
cc_287 N_B_c_280_n N_Y_c_666_n 0.0102239f $X=6.325 $Y=1.185 $X2=0 $Y2=0
cc_288 N_B_c_277_n N_Y_c_701_n 3.32215e-19 $X=5.755 $Y=1.675 $X2=0 $Y2=0
cc_289 N_B_c_301_n N_Y_c_701_n 4.18148e-19 $X=5.755 $Y=1.765 $X2=0 $Y2=0
cc_290 N_B_c_279_n N_Y_c_701_n 7.08536e-19 $X=6.205 $Y=1.675 $X2=0 $Y2=0
cc_291 N_B_c_303_n N_Y_c_701_n 0.0141785f $X=6.205 $Y=1.765 $X2=0 $Y2=0
cc_292 N_B_c_283_n N_Y_c_701_n 7.32832e-19 $X=6.655 $Y=1.675 $X2=0 $Y2=0
cc_293 N_B_c_305_n N_Y_c_701_n 0.0142979f $X=6.655 $Y=1.765 $X2=0 $Y2=0
cc_294 N_B_c_285_n N_Y_c_701_n 3.44604e-19 $X=7.155 $Y=1.675 $X2=0 $Y2=0
cc_295 N_B_c_307_n N_Y_c_701_n 3.85846e-19 $X=7.155 $Y=1.765 $X2=0 $Y2=0
cc_296 N_B_c_283_n N_Y_c_667_n 0.0135684f $X=6.655 $Y=1.675 $X2=0 $Y2=0
cc_297 N_B_c_284_n N_Y_c_667_n 0.00492465f $X=7.065 $Y=1.26 $X2=0 $Y2=0
cc_298 N_B_c_285_n N_Y_c_667_n 0.0209772f $X=7.155 $Y=1.675 $X2=0 $Y2=0
cc_299 N_B_c_286_n N_Y_c_667_n 0.0105573f $X=7.605 $Y=1.675 $X2=0 $Y2=0
cc_300 N_B_c_291_n N_Y_c_667_n 0.00252388f $X=7.38 $Y=1.26 $X2=0 $Y2=0
cc_301 N_B_c_293_n N_Y_c_667_n 0.0282229f $X=7.39 $Y=0.465 $X2=0 $Y2=0
cc_302 N_B_c_269_n N_Y_c_668_n 0.0127495f $X=4.21 $Y=1.185 $X2=0 $Y2=0
cc_303 N_B_c_270_n N_Y_c_668_n 0.0145311f $X=4.305 $Y=1.675 $X2=0 $Y2=0
cc_304 N_B_c_295_n N_Y_c_668_n 4.95215e-19 $X=4.305 $Y=1.765 $X2=0 $Y2=0
cc_305 N_B_c_271_n N_Y_c_668_n 0.0172053f $X=4.715 $Y=1.26 $X2=0 $Y2=0
cc_306 N_B_c_272_n N_Y_c_668_n 0.0140589f $X=4.805 $Y=1.675 $X2=0 $Y2=0
cc_307 N_B_c_297_n N_Y_c_668_n 0.00936307f $X=4.805 $Y=1.765 $X2=0 $Y2=0
cc_308 N_B_c_273_n N_Y_c_668_n 0.0140604f $X=5.215 $Y=1.26 $X2=0 $Y2=0
cc_309 N_B_c_274_n N_Y_c_668_n 0.0141477f $X=5.305 $Y=1.675 $X2=0 $Y2=0
cc_310 N_B_c_299_n N_Y_c_668_n 0.00939569f $X=5.305 $Y=1.765 $X2=0 $Y2=0
cc_311 N_B_c_275_n N_Y_c_668_n 0.0190402f $X=5.325 $Y=1.185 $X2=0 $Y2=0
cc_312 N_B_c_276_n N_Y_c_668_n 0.00848084f $X=5.665 $Y=1.26 $X2=0 $Y2=0
cc_313 N_B_c_277_n N_Y_c_668_n 0.0182482f $X=5.755 $Y=1.675 $X2=0 $Y2=0
cc_314 N_B_c_301_n N_Y_c_668_n 0.00355833f $X=5.755 $Y=1.765 $X2=0 $Y2=0
cc_315 N_B_c_278_n N_Y_c_668_n 0.00632967f $X=5.895 $Y=1.185 $X2=0 $Y2=0
cc_316 N_B_c_279_n N_Y_c_668_n 0.0193546f $X=6.205 $Y=1.675 $X2=0 $Y2=0
cc_317 N_B_c_280_n N_Y_c_668_n 0.00260099f $X=6.325 $Y=1.185 $X2=0 $Y2=0
cc_318 N_B_c_282_n N_Y_c_668_n 0.0256212f $X=6.4 $Y=1.26 $X2=0 $Y2=0
cc_319 N_B_c_283_n N_Y_c_668_n 0.00382311f $X=6.655 $Y=1.675 $X2=0 $Y2=0
cc_320 N_B_c_287_n N_Y_c_668_n 0.0113753f $X=4.265 $Y=1.26 $X2=0 $Y2=0
cc_321 N_B_c_288_n N_Y_c_668_n 0.0070628f $X=4.805 $Y=1.26 $X2=0 $Y2=0
cc_322 N_B_c_289_n N_Y_c_668_n 0.00261306f $X=5.307 $Y=1.26 $X2=0 $Y2=0
cc_323 N_B_c_283_n N_Y_c_736_n 3.44604e-19 $X=6.655 $Y=1.675 $X2=0 $Y2=0
cc_324 N_B_c_305_n N_Y_c_736_n 3.85846e-19 $X=6.655 $Y=1.765 $X2=0 $Y2=0
cc_325 N_B_c_285_n N_Y_c_736_n 7.32832e-19 $X=7.155 $Y=1.675 $X2=0 $Y2=0
cc_326 N_B_c_307_n N_Y_c_736_n 0.0143001f $X=7.155 $Y=1.765 $X2=0 $Y2=0
cc_327 N_B_c_286_n N_Y_c_736_n 0.00128334f $X=7.605 $Y=1.675 $X2=0 $Y2=0
cc_328 N_B_c_309_n N_Y_c_736_n 0.0179284f $X=7.605 $Y=1.765 $X2=0 $Y2=0
cc_329 N_B_c_269_n N_VGND_c_783_n 0.00571001f $X=4.21 $Y=1.185 $X2=0 $Y2=0
cc_330 N_B_c_269_n N_VGND_c_784_n 0.00433139f $X=4.21 $Y=1.185 $X2=0 $Y2=0
cc_331 N_B_c_275_n N_VGND_c_784_n 0.00433139f $X=5.325 $Y=1.185 $X2=0 $Y2=0
cc_332 N_B_c_275_n N_VGND_c_785_n 0.00701523f $X=5.325 $Y=1.185 $X2=0 $Y2=0
cc_333 N_B_c_276_n N_VGND_c_785_n 0.00167326f $X=5.665 $Y=1.26 $X2=0 $Y2=0
cc_334 N_B_c_278_n N_VGND_c_785_n 0.00563364f $X=5.895 $Y=1.185 $X2=0 $Y2=0
cc_335 N_B_c_278_n N_VGND_c_786_n 0.00434272f $X=5.895 $Y=1.185 $X2=0 $Y2=0
cc_336 N_B_c_280_n N_VGND_c_786_n 0.00434272f $X=6.325 $Y=1.185 $X2=0 $Y2=0
cc_337 N_B_c_280_n N_VGND_c_787_n 0.00963146f $X=6.325 $Y=1.185 $X2=0 $Y2=0
cc_338 N_B_c_281_n N_VGND_c_787_n 0.00977659f $X=6.565 $Y=1.26 $X2=0 $Y2=0
cc_339 N_B_c_292_n N_VGND_c_787_n 0.0104159f $X=7.39 $Y=0.465 $X2=0 $Y2=0
cc_340 N_B_c_293_n N_VGND_c_787_n 0.0317365f $X=7.39 $Y=0.465 $X2=0 $Y2=0
cc_341 N_B_c_292_n N_VGND_c_790_n 0.0127398f $X=7.39 $Y=0.465 $X2=0 $Y2=0
cc_342 N_B_c_293_n N_VGND_c_790_n 0.0172176f $X=7.39 $Y=0.465 $X2=0 $Y2=0
cc_343 N_B_c_269_n N_VGND_c_791_n 0.00822102f $X=4.21 $Y=1.185 $X2=0 $Y2=0
cc_344 N_B_c_275_n N_VGND_c_791_n 0.00822624f $X=5.325 $Y=1.185 $X2=0 $Y2=0
cc_345 N_B_c_278_n N_VGND_c_791_n 0.00821294f $X=5.895 $Y=1.185 $X2=0 $Y2=0
cc_346 N_B_c_280_n N_VGND_c_791_n 0.00825059f $X=6.325 $Y=1.185 $X2=0 $Y2=0
cc_347 N_B_c_292_n N_VGND_c_791_n 0.010606f $X=7.39 $Y=0.465 $X2=0 $Y2=0
cc_348 N_B_c_293_n N_VGND_c_791_n 0.0122345f $X=7.39 $Y=0.465 $X2=0 $Y2=0
cc_349 N_A_27_368#_c_424_n N_VPWR_M1000_s 0.00250873f $X=1.145 $Y=1.865
+ $X2=-0.19 $Y2=1.66
cc_350 N_A_27_368#_c_451_n N_VPWR_M1013_s 0.00356523f $X=2.045 $Y=2.035 $X2=0
+ $Y2=0
cc_351 N_A_27_368#_c_460_n N_VPWR_M1017_s 0.00452363f $X=2.995 $Y=2.035 $X2=0
+ $Y2=0
cc_352 N_A_27_368#_c_467_n N_VPWR_M1021_s 0.00588226f $X=3.915 $Y=2.035 $X2=0
+ $Y2=0
cc_353 N_A_27_368#_c_423_n N_VPWR_c_563_n 0.0330597f $X=0.28 $Y=1.985 $X2=0
+ $Y2=0
cc_354 N_A_27_368#_c_424_n N_VPWR_c_563_n 0.0202249f $X=1.145 $Y=1.865 $X2=0
+ $Y2=0
cc_355 N_A_27_368#_c_426_n N_VPWR_c_563_n 0.0560128f $X=1.23 $Y=2.435 $X2=0
+ $Y2=0
cc_356 N_A_27_368#_c_426_n N_VPWR_c_564_n 0.0449718f $X=1.23 $Y=2.435 $X2=0
+ $Y2=0
cc_357 N_A_27_368#_c_451_n N_VPWR_c_564_n 0.0171813f $X=2.045 $Y=2.035 $X2=0
+ $Y2=0
cc_358 N_A_27_368#_c_427_n N_VPWR_c_564_n 0.0462948f $X=2.13 $Y=2.435 $X2=0
+ $Y2=0
cc_359 N_A_27_368#_c_427_n N_VPWR_c_565_n 0.0256025f $X=2.13 $Y=2.435 $X2=0
+ $Y2=0
cc_360 N_A_27_368#_c_460_n N_VPWR_c_565_n 0.0202249f $X=2.995 $Y=2.035 $X2=0
+ $Y2=0
cc_361 N_A_27_368#_c_428_n N_VPWR_c_565_n 0.0462948f $X=3.08 $Y=2.435 $X2=0
+ $Y2=0
cc_362 N_A_27_368#_c_428_n N_VPWR_c_566_n 0.0256025f $X=3.08 $Y=2.435 $X2=0
+ $Y2=0
cc_363 N_A_27_368#_c_467_n N_VPWR_c_566_n 0.0232685f $X=3.915 $Y=2.035 $X2=0
+ $Y2=0
cc_364 N_A_27_368#_c_430_n N_VPWR_c_566_n 0.0119239f $X=4.245 $Y=2.99 $X2=0
+ $Y2=0
cc_365 N_A_27_368#_c_423_n N_VPWR_c_567_n 0.0145938f $X=0.28 $Y=1.985 $X2=0
+ $Y2=0
cc_366 N_A_27_368#_c_426_n N_VPWR_c_568_n 0.00749631f $X=1.23 $Y=2.435 $X2=0
+ $Y2=0
cc_367 N_A_27_368#_c_427_n N_VPWR_c_569_n 0.0110241f $X=2.13 $Y=2.435 $X2=0
+ $Y2=0
cc_368 N_A_27_368#_c_428_n N_VPWR_c_570_n 0.0110241f $X=3.08 $Y=2.435 $X2=0
+ $Y2=0
cc_369 N_A_27_368#_c_429_n N_VPWR_c_571_n 0.0429194f $X=4.925 $Y=2.99 $X2=0
+ $Y2=0
cc_370 N_A_27_368#_c_430_n N_VPWR_c_571_n 0.0235512f $X=4.245 $Y=2.99 $X2=0
+ $Y2=0
cc_371 N_A_27_368#_c_431_n N_VPWR_c_571_n 0.043517f $X=5.875 $Y=2.99 $X2=0 $Y2=0
cc_372 N_A_27_368#_c_433_n N_VPWR_c_571_n 0.0438391f $X=6.775 $Y=2.99 $X2=0
+ $Y2=0
cc_373 N_A_27_368#_c_435_n N_VPWR_c_571_n 0.0665295f $X=7.715 $Y=2.99 $X2=0
+ $Y2=0
cc_374 N_A_27_368#_c_438_n N_VPWR_c_571_n 0.0186386f $X=5.055 $Y=2.99 $X2=0
+ $Y2=0
cc_375 N_A_27_368#_c_439_n N_VPWR_c_571_n 0.0146958f $X=5.977 $Y=2.99 $X2=0
+ $Y2=0
cc_376 N_A_27_368#_c_440_n N_VPWR_c_571_n 0.0186386f $X=6.905 $Y=2.99 $X2=0
+ $Y2=0
cc_377 N_A_27_368#_c_423_n N_VPWR_c_562_n 0.0120466f $X=0.28 $Y=1.985 $X2=0
+ $Y2=0
cc_378 N_A_27_368#_c_426_n N_VPWR_c_562_n 0.0062048f $X=1.23 $Y=2.435 $X2=0
+ $Y2=0
cc_379 N_A_27_368#_c_427_n N_VPWR_c_562_n 0.00909194f $X=2.13 $Y=2.435 $X2=0
+ $Y2=0
cc_380 N_A_27_368#_c_428_n N_VPWR_c_562_n 0.00909194f $X=3.08 $Y=2.435 $X2=0
+ $Y2=0
cc_381 N_A_27_368#_c_429_n N_VPWR_c_562_n 0.0242621f $X=4.925 $Y=2.99 $X2=0
+ $Y2=0
cc_382 N_A_27_368#_c_430_n N_VPWR_c_562_n 0.0126924f $X=4.245 $Y=2.99 $X2=0
+ $Y2=0
cc_383 N_A_27_368#_c_431_n N_VPWR_c_562_n 0.0245693f $X=5.875 $Y=2.99 $X2=0
+ $Y2=0
cc_384 N_A_27_368#_c_433_n N_VPWR_c_562_n 0.0247572f $X=6.775 $Y=2.99 $X2=0
+ $Y2=0
cc_385 N_A_27_368#_c_435_n N_VPWR_c_562_n 0.0370229f $X=7.715 $Y=2.99 $X2=0
+ $Y2=0
cc_386 N_A_27_368#_c_438_n N_VPWR_c_562_n 0.0101082f $X=5.055 $Y=2.99 $X2=0
+ $Y2=0
cc_387 N_A_27_368#_c_439_n N_VPWR_c_562_n 0.00796993f $X=5.977 $Y=2.99 $X2=0
+ $Y2=0
cc_388 N_A_27_368#_c_440_n N_VPWR_c_562_n 0.0101082f $X=6.905 $Y=2.99 $X2=0
+ $Y2=0
cc_389 N_A_27_368#_c_429_n N_Y_M1001_s 0.00250873f $X=4.925 $Y=2.99 $X2=0 $Y2=0
cc_390 N_A_27_368#_c_431_n N_Y_M1006_s 0.00197722f $X=5.875 $Y=2.99 $X2=0 $Y2=0
cc_391 N_A_27_368#_c_433_n N_Y_M1011_s 0.00197722f $X=6.775 $Y=2.99 $X2=0 $Y2=0
cc_392 N_A_27_368#_c_435_n N_Y_M1018_s 0.00197722f $X=7.715 $Y=2.99 $X2=0 $Y2=0
cc_393 N_A_27_368#_c_429_n N_Y_c_670_n 0.018923f $X=4.925 $Y=2.99 $X2=0 $Y2=0
cc_394 N_A_27_368#_c_431_n N_Y_c_694_n 0.0160777f $X=5.875 $Y=2.99 $X2=0 $Y2=0
cc_395 N_A_27_368#_c_432_n N_Y_c_694_n 0.0335012f $X=5.98 $Y=1.985 $X2=0 $Y2=0
cc_396 N_A_27_368#_c_432_n N_Y_c_701_n 0.0327761f $X=5.98 $Y=1.985 $X2=0 $Y2=0
cc_397 N_A_27_368#_c_433_n N_Y_c_701_n 0.0160777f $X=6.775 $Y=2.99 $X2=0 $Y2=0
cc_398 N_A_27_368#_c_434_n N_Y_c_701_n 0.0335271f $X=6.93 $Y=1.985 $X2=0 $Y2=0
cc_399 N_A_27_368#_c_434_n N_Y_c_667_n 0.0217907f $X=6.93 $Y=1.985 $X2=0 $Y2=0
cc_400 N_A_27_368#_c_491_n N_Y_c_668_n 0.0227261f $X=5.08 $Y=2.115 $X2=0 $Y2=0
cc_401 N_A_27_368#_c_432_n N_Y_c_668_n 0.0189809f $X=5.98 $Y=1.985 $X2=0 $Y2=0
cc_402 N_A_27_368#_c_434_n N_Y_c_736_n 0.0335271f $X=6.93 $Y=1.985 $X2=0 $Y2=0
cc_403 N_A_27_368#_c_435_n N_Y_c_736_n 0.0160777f $X=7.715 $Y=2.99 $X2=0 $Y2=0
cc_404 N_A_27_368#_c_436_n N_Y_c_736_n 0.0351235f $X=7.88 $Y=1.985 $X2=0 $Y2=0
cc_405 N_A_27_368#_c_424_n N_VGND_c_781_n 0.0156334f $X=1.145 $Y=1.865 $X2=0
+ $Y2=0
cc_406 N_A_27_368#_c_437_n N_VGND_c_781_n 0.00606686f $X=1.23 $Y=1.865 $X2=0
+ $Y2=0
cc_407 N_Y_c_662_n N_VGND_M1007_d 0.00889788f $X=3.26 $Y=1.095 $X2=0 $Y2=0
cc_408 N_Y_c_665_n N_VGND_M1015_d 0.00250873f $X=4.26 $Y=1.095 $X2=0 $Y2=0
cc_409 N_Y_c_661_n N_VGND_c_781_n 0.0256093f $X=2.025 $Y=0.515 $X2=0 $Y2=0
cc_410 N_Y_c_663_n N_VGND_c_781_n 0.00594067f $X=2.19 $Y=1.095 $X2=0 $Y2=0
cc_411 N_Y_c_661_n N_VGND_c_782_n 0.0213338f $X=2.025 $Y=0.515 $X2=0 $Y2=0
cc_412 N_Y_c_662_n N_VGND_c_782_n 0.0535301f $X=3.26 $Y=1.095 $X2=0 $Y2=0
cc_413 N_Y_c_664_n N_VGND_c_782_n 0.019268f $X=3.425 $Y=0.515 $X2=0 $Y2=0
cc_414 N_Y_c_664_n N_VGND_c_783_n 0.0191765f $X=3.425 $Y=0.515 $X2=0 $Y2=0
cc_415 N_Y_c_665_n N_VGND_c_783_n 0.0209867f $X=4.26 $Y=1.095 $X2=0 $Y2=0
cc_416 N_Y_c_668_n N_VGND_c_783_n 0.0214346f $X=6.595 $Y=1.565 $X2=0 $Y2=0
cc_417 N_Y_c_668_n N_VGND_c_784_n 0.0451408f $X=6.595 $Y=1.565 $X2=0 $Y2=0
cc_418 N_Y_c_666_n N_VGND_c_785_n 0.0240544f $X=6.11 $Y=0.515 $X2=0 $Y2=0
cc_419 N_Y_c_668_n N_VGND_c_785_n 0.0560141f $X=6.595 $Y=1.565 $X2=0 $Y2=0
cc_420 N_Y_c_666_n N_VGND_c_786_n 0.0144922f $X=6.11 $Y=0.515 $X2=0 $Y2=0
cc_421 N_Y_c_666_n N_VGND_c_787_n 0.0308485f $X=6.11 $Y=0.515 $X2=0 $Y2=0
cc_422 N_Y_c_667_n N_VGND_c_787_n 0.0085367f $X=7.215 $Y=1.565 $X2=0 $Y2=0
cc_423 N_Y_c_668_n N_VGND_c_787_n 0.00828005f $X=6.595 $Y=1.565 $X2=0 $Y2=0
cc_424 N_Y_c_661_n N_VGND_c_788_n 0.0145639f $X=2.025 $Y=0.515 $X2=0 $Y2=0
cc_425 N_Y_c_664_n N_VGND_c_789_n 0.0145639f $X=3.425 $Y=0.515 $X2=0 $Y2=0
cc_426 N_Y_c_661_n N_VGND_c_791_n 0.0119984f $X=2.025 $Y=0.515 $X2=0 $Y2=0
cc_427 N_Y_c_664_n N_VGND_c_791_n 0.0119984f $X=3.425 $Y=0.515 $X2=0 $Y2=0
cc_428 N_Y_c_666_n N_VGND_c_791_n 0.0118826f $X=6.11 $Y=0.515 $X2=0 $Y2=0
cc_429 N_Y_c_668_n N_VGND_c_791_n 0.0372462f $X=6.595 $Y=1.565 $X2=0 $Y2=0
