* File: sky130_fd_sc_ls__sdfbbp_1.spice
* Created: Wed Sep  2 11:26:46 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__sdfbbp_1.pex.spice"
.subckt sky130_fd_sc_ls__sdfbbp_1  VNB VPB SCD D SCE CLK SET_B RESET_B VPWR Q_N
+ Q VGND
* 
* VGND	VGND
* Q	Q
* Q_N	Q_N
* VPWR	VPWR
* RESET_B	RESET_B
* SET_B	SET_B
* CLK	CLK
* SCE	SCE
* D	D
* SCD	SCD
* VPB	VPB
* VNB	VNB
MM1006 A_119_119# N_SCD_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.2 A=0.063 P=1.14 MULT=1
MM1029 N_A_197_119#_M1029_d N_SCE_M1029_g A_119_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.0756 AS=0.0504 PD=0.78 PS=0.66 NRD=22.848 NRS=18.564 M=1 R=2.8 SA=75000.6
+ SB=75001.8 A=0.063 P=1.14 MULT=1
MM1009 A_299_119# N_D_M1009_g N_A_197_119#_M1029_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0756 PD=0.63 PS=0.78 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001.1
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1012 N_VGND_M1012_d N_A_341_93#_M1012_g A_299_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.1155 AS=0.0441 PD=0.97 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.5
+ SB=75000.9 A=0.063 P=1.14 MULT=1
MM1041 N_A_341_93#_M1041_d N_SCE_M1041_g N_VGND_M1012_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.1155 PD=1.41 PS=0.97 NRD=0 NRS=77.136 M=1 R=2.8 SA=75002.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1042 N_VGND_M1042_d N_CLK_M1042_g N_A_622_98#_M1042_s VNB NSHORT L=0.15 W=0.74
+ AD=0.30025 AS=0.2109 PD=1.74 PS=2.05 NRD=56.868 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1000 N_A_877_98#_M1000_d N_A_622_98#_M1000_g N_VGND_M1042_d VNB NSHORT L=0.15
+ W=0.74 AD=0.2516 AS=0.30025 PD=2.16 PS=1.74 NRD=4.044 NRS=56.868 M=1 R=4.93333
+ SA=75001.1 SB=75000.3 A=0.111 P=1.78 MULT=1
MM1035 N_A_1092_96#_M1035_d N_A_622_98#_M1035_g N_A_197_119#_M1035_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0735 AS=0.1197 PD=0.77 PS=1.41 NRD=19.992 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002.3 A=0.063 P=1.14 MULT=1
MM1030 A_1192_96# N_A_877_98#_M1030_g N_A_1092_96#_M1035_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0809375 AS=0.0735 PD=0.89 PS=0.77 NRD=39.336 NRS=0 M=1 R=2.8
+ SA=75000.7 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1046 N_VGND_M1046_d N_A_1250_231#_M1046_g A_1192_96# VNB NSHORT L=0.15 W=0.42
+ AD=0.151254 AS=0.0809375 PD=1.16907 PS=0.89 NRD=87.168 NRS=39.336 M=1 R=2.8
+ SA=75000.8 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1022 N_A_1418_125#_M1022_d N_SET_B_M1022_g N_VGND_M1046_d VNB NSHORT L=0.15
+ W=0.55 AD=0.229287 AS=0.198071 PD=1.45 PS=1.53093 NRD=78.948 NRS=66.564 M=1
+ R=3.66667 SA=75001.2 SB=75001.5 A=0.0825 P=1.4 MULT=1
MM1015 N_A_1250_231#_M1015_d N_A_1092_96#_M1015_g N_A_1418_125#_M1022_d VNB
+ NSHORT L=0.15 W=0.55 AD=0.077 AS=0.229287 PD=0.83 PS=1.45 NRD=0 NRS=78.948 M=1
+ R=3.66667 SA=75001.9 SB=75000.8 A=0.0825 P=1.4 MULT=1
MM1016 N_A_1418_125#_M1016_d N_A_1625_93#_M1016_g N_A_1250_231#_M1015_d VNB
+ NSHORT L=0.15 W=0.55 AD=0.322425 AS=0.077 PD=2.47 PS=0.83 NRD=115.896 NRS=0
+ M=1 R=3.66667 SA=75002.3 SB=75000.3 A=0.0825 P=1.4 MULT=1
MM1013 A_1880_119# N_A_1250_231#_M1013_g N_VGND_M1013_s VNB NSHORT L=0.15 W=0.55
+ AD=0.05775 AS=0.15675 PD=0.76 PS=1.67 NRD=10.908 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75001.5 A=0.0825 P=1.4 MULT=1
MM1001 N_A_1878_420#_M1001_d N_A_877_98#_M1001_g A_1880_119# VNB NSHORT L=0.15
+ W=0.55 AD=0.132936 AS=0.05775 PD=1.3268 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667
+ SA=75000.6 SB=75001.1 A=0.0825 P=1.4 MULT=1
MM1023 A_2061_74# N_A_622_98#_M1023_g N_A_1878_420#_M1001_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0819 AS=0.101514 PD=0.81 PS=1.0132 NRD=39.996 NRS=53.34 M=1 R=2.8
+ SA=75000.6 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1047 N_VGND_M1047_d N_A_2037_442#_M1047_g A_2061_74# VNB NSHORT L=0.15 W=0.42
+ AD=0.0877655 AS=0.0819 PD=0.796552 PS=0.81 NRD=23.568 NRS=39.996 M=1 R=2.8
+ SA=75001.2 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1002 N_A_2271_74#_M1002_d N_SET_B_M1002_g N_VGND_M1047_d VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.154634 PD=1.02 PS=1.40345 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001 SB=75001.2 A=0.111 P=1.78 MULT=1
MM1031 N_A_2037_442#_M1031_d N_A_1878_420#_M1031_g N_A_2271_74#_M1002_d VNB
+ NSHORT L=0.15 W=0.74 AD=0.1443 AS=0.1036 PD=1.13 PS=1.02 NRD=17.832 NRS=0 M=1
+ R=4.93333 SA=75001.5 SB=75000.8 A=0.111 P=1.78 MULT=1
MM1043 N_A_2271_74#_M1043_d N_A_1625_93#_M1043_g N_A_2037_442#_M1031_d VNB
+ NSHORT L=0.15 W=0.74 AD=0.2146 AS=0.1443 PD=2.06 PS=1.13 NRD=0.804 NRS=0 M=1
+ R=4.93333 SA=75002 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1007 N_VGND_M1007_d N_RESET_B_M1007_g N_A_1625_93#_M1007_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0783879 AS=0.1197 PD=0.771207 PS=1.41 NRD=5.712 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1032 N_Q_N_M1032_d N_A_2037_442#_M1032_g N_VGND_M1007_d VNB NSHORT L=0.15
+ W=0.74 AD=0.2109 AS=0.138112 PD=2.05 PS=1.35879 NRD=0 NRS=4.044 M=1 R=4.93333
+ SA=75000.5 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1025 N_VGND_M1025_d N_A_2037_442#_M1025_g N_A_2881_74#_M1025_s VNB NSHORT
+ L=0.15 W=0.55 AD=0.129591 AS=0.15675 PD=0.997674 PS=1.67 NRD=18 NRS=0 M=1
+ R=3.66667 SA=75000.2 SB=75000.8 A=0.0825 P=1.4 MULT=1
MM1003 N_Q_M1003_d N_A_2881_74#_M1003_g N_VGND_M1025_d VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.174359 PD=2.05 PS=1.34233 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75000.7 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1026 N_VPWR_M1026_d N_SCD_M1026_g N_A_27_464#_M1026_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1152 AS=0.1888 PD=1 PS=1.87 NRD=18.4589 NRS=3.0732 M=1 R=4.26667
+ SA=75000.2 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1018 A_218_464# N_SCE_M1018_g N_VPWR_M1026_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0864 AS=0.1152 PD=0.91 PS=1 NRD=24.625 NRS=6.1464 M=1 R=4.26667
+ SA=75000.7 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1010 N_A_197_119#_M1010_d N_D_M1010_g A_218_464# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.096 AS=0.0864 PD=0.94 PS=0.91 NRD=3.0732 NRS=24.625 M=1 R=4.26667
+ SA=75001.1 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1019 N_A_27_464#_M1019_d N_A_341_93#_M1019_g N_A_197_119#_M1010_d VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.1888 AS=0.096 PD=1.87 PS=0.94 NRD=3.0732 NRS=3.0732 M=1
+ R=4.26667 SA=75001.6 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1027 N_A_341_93#_M1027_d N_SCE_M1027_g N_VPWR_M1027_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1888 AS=0.1888 PD=1.87 PS=1.87 NRD=3.0732 NRS=3.0732 M=1 R=4.26667
+ SA=75000.2 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1040 N_VPWR_M1040_d N_CLK_M1040_g N_A_622_98#_M1040_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1004 N_A_877_98#_M1004_d N_A_622_98#_M1004_g N_VPWR_M1040_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1014 N_A_1092_96#_M1014_d N_A_877_98#_M1014_g N_A_197_119#_M1014_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.140438 AS=0.1888 PD=1.27396 PS=1.87 NRD=27.6982 NRS=3.0732
+ M=1 R=4.26667 SA=75000.2 SB=75002.7 A=0.096 P=1.58 MULT=1
MM1005 A_1221_419# N_A_622_98#_M1005_g N_A_1092_96#_M1014_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0567 AS=0.0921623 PD=0.69 PS=0.836038 NRD=37.5088 NRS=21.0987 M=1
+ R=2.8 SA=75000.8 SB=75003.5 A=0.063 P=1.14 MULT=1
MM1045 N_VPWR_M1045_d N_A_1250_231#_M1045_g A_1221_419# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1572 AS=0.0567 PD=1.01667 PS=0.69 NRD=45.7237 NRS=37.5088 M=1
+ R=2.8 SA=75001.2 SB=75003.1 A=0.063 P=1.14 MULT=1
MM1024 N_A_1250_231#_M1024_d N_SET_B_M1024_g N_VPWR_M1045_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.1638 AS=0.3144 PD=1.23 PS=2.03333 NRD=23.443 NRS=72.693 M=1 R=5.6
+ SA=75001.2 SB=75002.9 A=0.126 P=1.98 MULT=1
MM1039 A_1580_379# N_A_1092_96#_M1039_g N_A_1250_231#_M1024_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.1134 AS=0.1638 PD=1.11 PS=1.23 NRD=18.7544 NRS=2.3443 M=1 R=5.6
+ SA=75001.7 SB=75002.3 A=0.126 P=1.98 MULT=1
MM1033 N_VPWR_M1033_d N_A_1625_93#_M1033_g A_1580_379# VPB PHIGHVT L=0.15 W=0.84
+ AD=0.1512 AS=0.1134 PD=1.2 PS=1.11 NRD=9.3772 NRS=18.7544 M=1 R=5.6 SA=75002.2
+ SB=75001.9 A=0.126 P=1.98 MULT=1
MM1034 A_1766_379# N_A_1250_231#_M1034_g N_VPWR_M1033_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.1845 AS=0.1512 PD=1.455 PS=1.2 NRD=38.612 NRS=9.3772 M=1 R=5.6
+ SA=75002.7 SB=75001.4 A=0.126 P=1.98 MULT=1
MM1008 N_A_1878_420#_M1008_d N_A_622_98#_M1008_g A_1766_379# VPB PHIGHVT L=0.15
+ W=0.84 AD=0.1932 AS=0.1845 PD=1.64 PS=1.455 NRD=2.3443 NRS=38.612 M=1 R=5.6
+ SA=75002.7 SB=75001.7 A=0.126 P=1.98 MULT=1
MM1020 A_1986_504# N_A_877_98#_M1020_g N_A_1878_420#_M1008_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0567 AS=0.0966 PD=0.69 PS=0.82 NRD=37.5088 NRS=46.886 M=1 R=2.8
+ SA=75001.9 SB=75002.6 A=0.063 P=1.14 MULT=1
MM1036 N_VPWR_M1036_d N_A_2037_442#_M1036_g A_1986_504# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.158491 AS=0.0567 PD=1.11211 PS=0.69 NRD=51.5943 NRS=37.5088 M=1
+ R=2.8 SA=75002.4 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1037 N_A_2037_442#_M1037_d N_SET_B_M1037_g N_VPWR_M1036_d VPB PHIGHVT L=0.15
+ W=1 AD=0.2 AS=0.377359 PD=1.4 PS=2.64789 NRD=21.67 NRS=18.715 M=1 R=6.66667
+ SA=75001.5 SB=75001.1 A=0.15 P=2.3 MULT=1
MM1044 A_2384_392# N_A_1878_420#_M1044_g N_A_2037_442#_M1037_d VPB PHIGHVT
+ L=0.15 W=1 AD=0.12 AS=0.2 PD=1.24 PS=1.4 NRD=12.7853 NRS=1.9503 M=1 R=6.66667
+ SA=75002.1 SB=75000.6 A=0.15 P=2.3 MULT=1
MM1017 N_VPWR_M1017_d N_A_1625_93#_M1017_g A_2384_392# VPB PHIGHVT L=0.15 W=1
+ AD=0.28 AS=0.12 PD=2.56 PS=1.24 NRD=1.9503 NRS=12.7853 M=1 R=6.66667
+ SA=75002.5 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1028 N_VPWR_M1028_d N_RESET_B_M1028_g N_A_1625_93#_M1028_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.132945 AS=0.1792 PD=1.08 PS=1.84 NRD=47.0042 NRS=3.0732 M=1
+ R=4.26667 SA=75000.2 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1021 N_Q_N_M1021_d N_A_2037_442#_M1021_g N_VPWR_M1028_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.308 AS=0.232655 PD=2.79 PS=1.89 NRD=1.7533 NRS=1.7533 M=1
+ R=7.46667 SA=75000.5 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1011 N_VPWR_M1011_d N_A_2037_442#_M1011_g N_A_2881_74#_M1011_s VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.1614 AS=0.2478 PD=1.26857 PS=2.27 NRD=15.2281 NRS=2.3443
+ M=1 R=5.6 SA=75000.2 SB=75000.7 A=0.126 P=1.98 MULT=1
MM1038 N_Q_M1038_d N_A_2881_74#_M1038_g N_VPWR_M1011_d VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3192 AS=0.2152 PD=2.81 PS=1.69143 NRD=1.7533 NRS=2.6201 M=1 R=7.46667
+ SA=75000.6 SB=75000.2 A=0.168 P=2.54 MULT=1
DX48_noxref VNB VPB NWDIODE A=30.3272 P=36.36
c_177 VNB 0 3.53193e-20 $X=0 $Y=0
c_2191 A_218_464# 0 1.00461e-19 $X=1.09 $Y=2.32
c_2372 A_1766_379# 0 9.6863e-20 $X=8.83 $Y=1.895
*
.include "sky130_fd_sc_ls__sdfbbp_1.pxi.spice"
*
.ends
*
*
