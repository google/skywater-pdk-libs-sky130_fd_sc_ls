* NGSPICE file created from sky130_fd_sc_ls__nor3_2.ext - technology: sky130A

.subckt sky130_fd_sc_ls__nor3_2 A B C VGND VNB VPB VPWR Y
M1000 a_306_368# A VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=7.056e+11p pd=5.74e+06u as=3.584e+11p ps=2.88e+06u
M1001 VPWR A a_306_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_27_368# B a_306_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=9.968e+11p pd=8.5e+06u as=0p ps=0u
M1003 a_27_368# C Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.92e+11p ps=2.94e+06u
M1004 Y C a_27_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_306_368# B a_27_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND C Y VNB nshort w=740000u l=150000u
+  ad=9.176e+11p pd=5.44e+06u as=4.699e+11p ps=4.23e+06u
M1007 VGND A Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y B VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

