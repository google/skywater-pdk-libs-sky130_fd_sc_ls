# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ls__nor2_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_ls__nor2_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.160000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  1.788000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 1.350000 3.715000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.788000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.225000 0.300000 7.555000 1.310000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  2.839300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.860000 0.350000 2.190000 1.010000 ;
        RECT 1.860000 1.010000 5.275000 1.140000 ;
        RECT 1.860000 1.140000 6.275000 1.180000 ;
        RECT 3.260000 0.350000 3.590000 1.010000 ;
        RECT 4.260000 0.350000 5.275000 1.010000 ;
        RECT 4.260000 1.180000 6.275000 1.310000 ;
        RECT 4.415000 1.310000 6.275000 1.480000 ;
        RECT 4.415000 1.480000 7.545000 1.650000 ;
        RECT 4.415000 1.650000 5.695000 1.780000 ;
        RECT 4.415000 1.780000 4.745000 2.735000 ;
        RECT 5.365000 1.780000 5.695000 2.735000 ;
        RECT 5.945000 0.350000 6.275000 1.140000 ;
        RECT 6.265000 1.650000 6.595000 2.735000 ;
        RECT 7.215000 1.650000 7.545000 2.735000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.160000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.160000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.160000 0.085000 ;
      RECT 0.000000  3.245000 8.160000 3.415000 ;
      RECT 0.115000  1.780000 1.315000 1.950000 ;
      RECT 0.115000  1.950000 0.445000 2.980000 ;
      RECT 0.615000  2.120000 0.945000 3.245000 ;
      RECT 0.650000  0.085000 1.690000 1.130000 ;
      RECT 1.145000  1.950000 4.245000 2.120000 ;
      RECT 1.145000  2.120000 1.315000 2.980000 ;
      RECT 1.515000  2.290000 1.845000 3.245000 ;
      RECT 2.045000  2.120000 2.295000 2.980000 ;
      RECT 2.360000  0.085000 3.090000 0.840000 ;
      RECT 2.465000  2.290000 2.795000 3.245000 ;
      RECT 2.995000  2.120000 3.245000 2.980000 ;
      RECT 3.415000  2.290000 3.745000 3.245000 ;
      RECT 3.760000  0.085000 4.090000 0.840000 ;
      RECT 3.915000  2.120000 4.245000 2.905000 ;
      RECT 3.915000  2.905000 8.045000 3.075000 ;
      RECT 4.925000  1.950000 5.185000 2.905000 ;
      RECT 5.445000  0.085000 5.775000 0.970000 ;
      RECT 5.875000  1.820000 6.080000 2.905000 ;
      RECT 6.445000  0.085000 6.775000 1.130000 ;
      RECT 6.775000  1.820000 7.035000 2.905000 ;
      RECT 7.715000  1.820000 8.045000 2.905000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
  END
END sky130_fd_sc_ls__nor2_8
END LIBRARY
