* File: sky130_fd_sc_ls__a222oi_2.spice
* Created: Fri Aug 28 12:54:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__a222oi_2.pex.spice"
.subckt sky130_fd_sc_ls__a222oi_2  VNB VPB C2 C1 B1 B2 A1 A2 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A2	A2
* A1	A1
* B2	B2
* B1	B1
* C1	C1
* C2	C2
* VPB	VPB
* VNB	VNB
MM1006 N_VGND_M1006_d N_C2_M1006_g N_A_137_74#_M1006_s VNB NSHORT L=0.15 W=0.64
+ AD=0.264125 AS=0.0896 PD=2.13 PS=0.92 NRD=18.744 NRS=0 M=1 R=4.26667
+ SA=75000.3 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1000 N_A_137_74#_M1006_s N_C1_M1000_g N_Y_M1000_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.8
+ SB=75001.1 A=0.096 P=1.58 MULT=1
MM1009 N_A_137_74#_M1009_d N_C1_M1009_g N_Y_M1000_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75001.2
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1008 N_VGND_M1008_d N_C2_M1008_g N_A_137_74#_M1009_d VNB NSHORT L=0.15 W=0.64
+ AD=0.1824 AS=0.0896 PD=1.85 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75001.6
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1018 N_A_593_74#_M1018_d N_B1_M1018_g N_Y_M1018_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.1824 PD=0.92 PS=1.85 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75003.5 A=0.096 P=1.58 MULT=1
MM1007 N_VGND_M1007_d N_B2_M1007_g N_A_593_74#_M1018_d VNB NSHORT L=0.15 W=0.64
+ AD=0.19325 AS=0.0896 PD=1.33 PS=0.92 NRD=46.296 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75003.1 A=0.096 P=1.58 MULT=1
MM1013 N_VGND_M1007_d N_B2_M1013_g N_A_593_74#_M1013_s VNB NSHORT L=0.15 W=0.64
+ AD=0.19325 AS=0.0896 PD=1.33 PS=0.92 NRD=46.296 NRS=0 M=1 R=4.26667 SA=75001.3
+ SB=75002.4 A=0.096 P=1.58 MULT=1
MM1020 N_A_593_74#_M1013_s N_B1_M1020_g N_Y_M1020_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75001.7
+ SB=75002 A=0.096 P=1.58 MULT=1
MM1002 N_A_981_74#_M1002_d N_A1_M1002_g N_Y_M1020_s VNB NSHORT L=0.15 W=0.64
+ AD=0.112 AS=0.0896 PD=0.99 PS=0.92 NRD=0.936 NRS=0 M=1 R=4.26667 SA=75002.1
+ SB=75001.6 A=0.096 P=1.58 MULT=1
MM1022 N_VGND_M1022_d N_A2_M1022_g N_A_981_74#_M1002_d VNB NSHORT L=0.15 W=0.64
+ AD=0.0928 AS=0.112 PD=0.93 PS=0.99 NRD=0.936 NRS=12.18 M=1 R=4.26667
+ SA=75002.6 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1023 N_VGND_M1022_d N_A2_M1023_g N_A_981_74#_M1023_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0928 AS=0.0896 PD=0.93 PS=0.92 NRD=0.936 NRS=0 M=1 R=4.26667 SA=75003.1
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1005 N_A_981_74#_M1023_s N_A1_M1005_g N_Y_M1005_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.1824 PD=0.92 PS=1.85 NRD=0 NRS=0 M=1 R=4.26667 SA=75003.5
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1010 N_Y_M1010_d N_C2_M1010_g N_A_116_392#_M1010_s VPB PHIGHVT L=0.15 W=1
+ AD=0.295 AS=0.15 PD=2.59 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75000.2
+ SB=75001.6 A=0.15 P=2.3 MULT=1
MM1003 N_A_116_392#_M1010_s N_C1_M1003_g N_Y_M1003_s VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.165 PD=1.3 PS=1.33 NRD=1.9503 NRS=4.9053 M=1 R=6.66667 SA=75000.7
+ SB=75001.2 A=0.15 P=2.3 MULT=1
MM1014 N_A_116_392#_M1014_d N_C1_M1014_g N_Y_M1003_s VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.165 PD=1.3 PS=1.33 NRD=1.9503 NRS=4.9053 M=1 R=6.66667 SA=75001.1
+ SB=75000.7 A=0.15 P=2.3 MULT=1
MM1016 N_Y_M1016_d N_C2_M1016_g N_A_116_392#_M1014_d VPB PHIGHVT L=0.15 W=1
+ AD=0.345 AS=0.15 PD=2.69 PS=1.3 NRD=11.8003 NRS=1.9503 M=1 R=6.66667
+ SA=75001.6 SB=75000.3 A=0.15 P=2.3 MULT=1
MM1011 N_A_515_392#_M1011_d N_B1_M1011_g N_A_116_392#_M1011_s VPB PHIGHVT L=0.15
+ W=1 AD=0.295 AS=0.15 PD=2.59 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75003.5 A=0.15 P=2.3 MULT=1
MM1001 N_A_116_392#_M1011_s N_B2_M1001_g N_A_515_392#_M1001_s VPB PHIGHVT L=0.15
+ W=1 AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75000.7 SB=75003 A=0.15 P=2.3 MULT=1
MM1021 N_A_116_392#_M1021_d N_B2_M1021_g N_A_515_392#_M1001_s VPB PHIGHVT L=0.15
+ W=1 AD=0.195 AS=0.15 PD=1.39 PS=1.3 NRD=10.8153 NRS=1.9503 M=1 R=6.66667
+ SA=75001.1 SB=75002.6 A=0.15 P=2.3 MULT=1
MM1015 N_A_515_392#_M1015_d N_B1_M1015_g N_A_116_392#_M1021_d VPB PHIGHVT L=0.15
+ W=1 AD=0.15 AS=0.195 PD=1.3 PS=1.39 NRD=1.9503 NRS=10.8153 M=1 R=6.66667
+ SA=75001.7 SB=75002 A=0.15 P=2.3 MULT=1
MM1017 N_A_515_392#_M1015_d N_A1_M1017_g N_VPWR_M1017_s VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.165 PD=1.3 PS=1.33 NRD=1.9503 NRS=4.9053 M=1 R=6.66667 SA=75002.1
+ SB=75001.6 A=0.15 P=2.3 MULT=1
MM1004 N_A_515_392#_M1004_d N_A2_M1004_g N_VPWR_M1017_s VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.165 PD=1.3 PS=1.33 NRD=1.9503 NRS=4.9053 M=1 R=6.66667 SA=75002.6
+ SB=75001.1 A=0.15 P=2.3 MULT=1
MM1012 N_A_515_392#_M1004_d N_A2_M1012_g N_VPWR_M1012_s VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75003
+ SB=75000.7 A=0.15 P=2.3 MULT=1
MM1019 N_A_515_392#_M1019_d N_A1_M1019_g N_VPWR_M1012_s VPB PHIGHVT L=0.15 W=1
+ AD=0.295 AS=0.15 PD=2.59 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75003.5
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX24_noxref VNB VPB NWDIODE A=13.206 P=17.92
c_125 VPB 0 1.3759e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_ls__a222oi_2.pxi.spice"
*
.ends
*
*
