* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__or2_2 A B VGND VNB VPB VPWR X
M1000 VPWR A a_114_368# VPB phighvt w=1e+06u l=150000u
+  ad=7.558e+11p pd=5.85e+06u as=2.4e+11p ps=2.48e+06u
M1001 VPWR a_27_368# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.584e+11p ps=2.88e+06u
M1002 VGND a_27_368# X VNB nshort w=740000u l=150000u
+  ad=6.823e+11p pd=6.18e+06u as=2.072e+11p ps=2.04e+06u
M1003 X a_27_368# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_27_368# B VGND VNB nshort w=640000u l=150000u
+  ad=1.792e+11p pd=1.84e+06u as=0p ps=0u
M1005 VGND A a_27_368# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 X a_27_368# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_114_368# B a_27_368# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.85e+11p ps=2.57e+06u
.ends
