* File: sky130_fd_sc_ls__inv_8.pex.spice
* Created: Fri Aug 28 13:28:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__INV_8%A 1 3 4 6 7 9 10 12 15 17 19 22 24 26 29 31 33
+ 36 38 40 43 45 47 48 50 52 54 55 56 57 74
r144 73 74 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=2.085
+ $Y=1.515 $X2=2.085 $Y2=1.515
r145 71 73 22.1893 $w=3.91e-07 $l=1.8e-07 $layer=POLY_cond $X=1.905 $Y=1.482
+ $X2=2.085 $Y2=1.482
r146 66 67 1.8491 $w=3.91e-07 $l=1.5e-08 $layer=POLY_cond $X=0.94 $Y=1.482
+ $X2=0.955 $Y2=1.482
r147 64 66 26.5038 $w=3.91e-07 $l=2.15e-07 $layer=POLY_cond $X=0.725 $Y=1.482
+ $X2=0.94 $Y2=1.482
r148 64 65 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=0.725
+ $Y=1.515 $X2=0.725 $Y2=1.515
r149 62 64 26.5038 $w=3.91e-07 $l=2.15e-07 $layer=POLY_cond $X=0.51 $Y=1.482
+ $X2=0.725 $Y2=1.482
r150 61 62 0.616368 $w=3.91e-07 $l=5e-09 $layer=POLY_cond $X=0.505 $Y=1.482
+ $X2=0.51 $Y2=1.482
r151 57 74 10.8544 $w=4.28e-07 $l=4.05e-07 $layer=LI1_cond $X=1.68 $Y=1.565
+ $X2=2.085 $Y2=1.565
r152 56 57 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.565
+ $X2=1.68 $Y2=1.565
r153 56 65 12.7305 $w=4.28e-07 $l=4.75e-07 $layer=LI1_cond $X=1.2 $Y=1.565
+ $X2=0.725 $Y2=1.565
r154 55 65 0.134005 $w=4.28e-07 $l=5e-09 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=0.725 $Y2=1.565
r155 52 82 25.3065 $w=1.5e-07 $l=2.83e-07 $layer=POLY_cond $X=3.755 $Y=1.765
+ $X2=3.755 $Y2=1.482
r156 52 54 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.755 $Y=1.765
+ $X2=3.755 $Y2=2.4
r157 48 82 3.08184 $w=3.91e-07 $l=2.5e-08 $layer=POLY_cond $X=3.73 $Y=1.482
+ $X2=3.755 $Y2=1.482
r158 48 80 52.3913 $w=3.91e-07 $l=4.25e-07 $layer=POLY_cond $X=3.73 $Y=1.482
+ $X2=3.305 $Y2=1.482
r159 48 50 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.73 $Y=1.35
+ $X2=3.73 $Y2=0.74
r160 45 80 25.3065 $w=1.5e-07 $l=2.83e-07 $layer=POLY_cond $X=3.305 $Y=1.765
+ $X2=3.305 $Y2=1.482
r161 45 47 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.305 $Y=1.765
+ $X2=3.305 $Y2=2.4
r162 41 80 0.616368 $w=3.91e-07 $l=5e-09 $layer=POLY_cond $X=3.3 $Y=1.482
+ $X2=3.305 $Y2=1.482
r163 41 78 61.0205 $w=3.91e-07 $l=4.95e-07 $layer=POLY_cond $X=3.3 $Y=1.482
+ $X2=2.805 $Y2=1.482
r164 41 43 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.3 $Y=1.35 $X2=3.3
+ $Y2=0.74
r165 38 78 25.3065 $w=1.5e-07 $l=2.83e-07 $layer=POLY_cond $X=2.805 $Y=1.765
+ $X2=2.805 $Y2=1.482
r166 38 40 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.805 $Y=1.765
+ $X2=2.805 $Y2=2.4
r167 34 78 9.24552 $w=3.91e-07 $l=7.5e-08 $layer=POLY_cond $X=2.73 $Y=1.482
+ $X2=2.805 $Y2=1.482
r168 34 76 46.2276 $w=3.91e-07 $l=3.75e-07 $layer=POLY_cond $X=2.73 $Y=1.482
+ $X2=2.355 $Y2=1.482
r169 34 36 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.73 $Y=1.35
+ $X2=2.73 $Y2=0.74
r170 31 76 25.3065 $w=1.5e-07 $l=2.83e-07 $layer=POLY_cond $X=2.355 $Y=1.765
+ $X2=2.355 $Y2=1.482
r171 31 33 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.355 $Y=1.765
+ $X2=2.355 $Y2=2.4
r172 27 76 6.78005 $w=3.91e-07 $l=5.5e-08 $layer=POLY_cond $X=2.3 $Y=1.482
+ $X2=2.355 $Y2=1.482
r173 27 73 26.5038 $w=3.91e-07 $l=2.15e-07 $layer=POLY_cond $X=2.3 $Y=1.482
+ $X2=2.085 $Y2=1.482
r174 27 29 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.3 $Y=1.35 $X2=2.3
+ $Y2=0.74
r175 24 71 25.3065 $w=1.5e-07 $l=2.83e-07 $layer=POLY_cond $X=1.905 $Y=1.765
+ $X2=1.905 $Y2=1.482
r176 24 26 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.905 $Y=1.765
+ $X2=1.905 $Y2=2.4
r177 20 71 12.9437 $w=3.91e-07 $l=1.05e-07 $layer=POLY_cond $X=1.8 $Y=1.482
+ $X2=1.905 $Y2=1.482
r178 20 69 42.5294 $w=3.91e-07 $l=3.45e-07 $layer=POLY_cond $X=1.8 $Y=1.482
+ $X2=1.455 $Y2=1.482
r179 20 22 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.8 $Y=1.35 $X2=1.8
+ $Y2=0.74
r180 17 69 25.3065 $w=1.5e-07 $l=2.83e-07 $layer=POLY_cond $X=1.455 $Y=1.765
+ $X2=1.455 $Y2=1.482
r181 17 19 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.455 $Y=1.765
+ $X2=1.455 $Y2=2.4
r182 13 69 10.4783 $w=3.91e-07 $l=8.5e-08 $layer=POLY_cond $X=1.37 $Y=1.482
+ $X2=1.455 $Y2=1.482
r183 13 67 51.1586 $w=3.91e-07 $l=4.15e-07 $layer=POLY_cond $X=1.37 $Y=1.482
+ $X2=0.955 $Y2=1.482
r184 13 15 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.37 $Y=1.35
+ $X2=1.37 $Y2=0.74
r185 10 67 25.3065 $w=1.5e-07 $l=2.83e-07 $layer=POLY_cond $X=0.955 $Y=1.765
+ $X2=0.955 $Y2=1.482
r186 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.955 $Y=1.765
+ $X2=0.955 $Y2=2.4
r187 7 66 25.3065 $w=1.5e-07 $l=2.82e-07 $layer=POLY_cond $X=0.94 $Y=1.2
+ $X2=0.94 $Y2=1.482
r188 7 9 147.813 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=0.94 $Y=1.2 $X2=0.94
+ $Y2=0.74
r189 4 62 25.3065 $w=1.5e-07 $l=2.82e-07 $layer=POLY_cond $X=0.51 $Y=1.2
+ $X2=0.51 $Y2=1.482
r190 4 6 147.813 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=0.51 $Y=1.2 $X2=0.51
+ $Y2=0.74
r191 1 61 25.3065 $w=1.5e-07 $l=2.83e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=1.482
r192 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__INV_8%VPWR 1 2 3 4 5 16 18 24 28 32 36 38 43 44 45
+ 47 52 61 69 72 76
r69 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r70 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r71 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r72 64 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r73 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r74 61 75 4.71369 $w=1.7e-07 $l=2.27e-07 $layer=LI1_cond $X=3.865 $Y=3.33
+ $X2=4.092 $Y2=3.33
r75 61 63 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.865 $Y=3.33
+ $X2=3.6 $Y2=3.33
r76 60 64 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r77 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r78 57 72 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.295 $Y=3.33
+ $X2=2.17 $Y2=3.33
r79 57 59 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.295 $Y=3.33
+ $X2=2.64 $Y2=3.33
r80 56 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r81 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r82 53 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.345 $Y=3.33
+ $X2=1.18 $Y2=3.33
r83 53 55 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.345 $Y=3.33
+ $X2=1.68 $Y2=3.33
r84 52 72 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.045 $Y=3.33
+ $X2=2.17 $Y2=3.33
r85 52 55 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.045 $Y=3.33
+ $X2=1.68 $Y2=3.33
r86 51 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r87 51 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r88 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r89 48 66 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.182 $Y2=3.33
r90 48 50 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.72 $Y2=3.33
r91 47 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.015 $Y=3.33
+ $X2=1.18 $Y2=3.33
r92 47 50 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.015 $Y=3.33
+ $X2=0.72 $Y2=3.33
r93 45 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r94 45 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r95 45 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r96 43 59 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.865 $Y=3.33
+ $X2=2.64 $Y2=3.33
r97 43 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.865 $Y=3.33
+ $X2=3.03 $Y2=3.33
r98 42 63 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=3.195 $Y=3.33
+ $X2=3.6 $Y2=3.33
r99 42 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.195 $Y=3.33
+ $X2=3.03 $Y2=3.33
r100 38 41 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=4.03 $Y=1.985
+ $X2=4.03 $Y2=2.815
r101 36 75 3.05248 $w=3.3e-07 $l=1.11781e-07 $layer=LI1_cond $X=4.03 $Y=3.245
+ $X2=4.092 $Y2=3.33
r102 36 41 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=4.03 $Y=3.245
+ $X2=4.03 $Y2=2.815
r103 32 35 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=3.03 $Y=1.985
+ $X2=3.03 $Y2=2.815
r104 30 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.03 $Y=3.245
+ $X2=3.03 $Y2=3.33
r105 30 35 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.03 $Y=3.245
+ $X2=3.03 $Y2=2.815
r106 26 72 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.17 $Y=3.245
+ $X2=2.17 $Y2=3.33
r107 26 28 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=2.17 $Y=3.245
+ $X2=2.17 $Y2=2.455
r108 22 69 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.18 $Y=3.245
+ $X2=1.18 $Y2=3.33
r109 22 24 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=1.18 $Y=3.245
+ $X2=1.18 $Y2=2.455
r110 18 21 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=0.24 $Y=1.985
+ $X2=0.24 $Y2=2.815
r111 16 66 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.182 $Y2=3.33
r112 16 21 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.24 $Y2=2.815
r113 5 41 400 $w=1.7e-07 $l=1.07034e-06 $layer=licon1_PDIFF $count=1 $X=3.83
+ $Y=1.84 $X2=4.03 $Y2=2.815
r114 5 38 400 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=1 $X=3.83
+ $Y=1.84 $X2=4.03 $Y2=1.985
r115 4 35 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.88
+ $Y=1.84 $X2=3.03 $Y2=2.815
r116 4 32 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.88
+ $Y=1.84 $X2=3.03 $Y2=1.985
r117 3 28 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=1.98
+ $Y=1.84 $X2=2.13 $Y2=2.455
r118 2 24 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=1.03
+ $Y=1.84 $X2=1.18 $Y2=2.455
r119 1 21 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r120 1 18 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_LS__INV_8%Y 1 2 3 4 5 6 7 8 27 29 31 33 34 35 39 43 45
+ 47 51 54 57 59 63 67 73 75 76 78 80 81
r133 79 81 9.59355 $w=4.78e-07 $l=3.85e-07 $layer=LI1_cond $X=3.695 $Y=1.38
+ $X2=4.08 $Y2=1.38
r134 79 80 1.71002 $w=4.8e-07 $l=1.73e-07 $layer=LI1_cond $X=3.695 $Y=1.38
+ $X2=3.522 $Y2=1.38
r135 67 69 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=3.53 $Y=1.985
+ $X2=3.53 $Y2=2.815
r136 65 80 4.64884 $w=3.3e-07 $l=2.43967e-07 $layer=LI1_cond $X=3.53 $Y=1.62
+ $X2=3.522 $Y2=1.38
r137 65 67 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=3.53 $Y=1.62
+ $X2=3.53 $Y2=1.985
r138 61 80 4.64884 $w=2.6e-07 $l=2.60154e-07 $layer=LI1_cond $X=3.48 $Y=1.14
+ $X2=3.522 $Y2=1.38
r139 61 63 27.703 $w=2.58e-07 $l=6.25e-07 $layer=LI1_cond $X=3.48 $Y=1.14
+ $X2=3.48 $Y2=0.515
r140 60 76 2.29025 $w=4.8e-07 $l=5.0892e-07 $layer=LI1_cond $X=2.68 $Y=1.38
+ $X2=2.35 $Y2=1.01
r141 59 80 1.71002 $w=4.8e-07 $l=1.72e-07 $layer=LI1_cond $X=3.35 $Y=1.38
+ $X2=3.522 $Y2=1.38
r142 59 60 16.6953 $w=4.78e-07 $l=6.7e-07 $layer=LI1_cond $X=3.35 $Y=1.38
+ $X2=2.68 $Y2=1.38
r143 55 78 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.58 $Y=2.12
+ $X2=2.58 $Y2=2.035
r144 55 57 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=2.58 $Y=2.12
+ $X2=2.58 $Y2=2.4
r145 54 78 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.58 $Y=1.95
+ $X2=2.58 $Y2=2.035
r146 53 76 3.88572 $w=1.7e-07 $l=7.15821e-07 $layer=LI1_cond $X=2.58 $Y=1.62
+ $X2=2.35 $Y2=1.01
r147 53 54 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.58 $Y=1.62
+ $X2=2.58 $Y2=1.95
r148 49 76 3.88572 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=2.515 $Y=1.01
+ $X2=2.35 $Y2=1.01
r149 49 51 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=2.515 $Y=1.01
+ $X2=2.515 $Y2=0.515
r150 48 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.845 $Y=2.035
+ $X2=1.68 $Y2=2.035
r151 47 78 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.495 $Y=2.035
+ $X2=2.58 $Y2=2.035
r152 47 48 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=2.495 $Y=2.035
+ $X2=1.845 $Y2=2.035
r153 46 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.67 $Y=1.095
+ $X2=1.585 $Y2=1.095
r154 45 76 2.29025 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.35 $Y=1.095
+ $X2=2.35 $Y2=1.01
r155 45 46 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.35 $Y=1.095
+ $X2=1.67 $Y2=1.095
r156 41 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.68 $Y=2.12
+ $X2=1.68 $Y2=2.035
r157 41 43 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=1.68 $Y=2.12
+ $X2=1.68 $Y2=2.815
r158 37 73 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.585 $Y=1.01
+ $X2=1.585 $Y2=1.095
r159 37 39 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=1.585 $Y=1.01
+ $X2=1.585 $Y2=0.515
r160 36 72 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.815 $Y=2.035
+ $X2=0.69 $Y2=2.035
r161 35 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.515 $Y=2.035
+ $X2=1.68 $Y2=2.035
r162 35 36 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.515 $Y=2.035
+ $X2=0.815 $Y2=2.035
r163 33 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.5 $Y=1.095
+ $X2=1.585 $Y2=1.095
r164 33 34 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.5 $Y=1.095
+ $X2=0.81 $Y2=1.095
r165 29 72 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=2.12
+ $X2=0.69 $Y2=2.035
r166 29 31 32.0379 $w=2.48e-07 $l=6.95e-07 $layer=LI1_cond $X=0.69 $Y=2.12
+ $X2=0.69 $Y2=2.815
r167 25 34 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.685 $Y=1.01
+ $X2=0.81 $Y2=1.095
r168 25 27 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=0.685 $Y=1.01
+ $X2=0.685 $Y2=0.515
r169 8 69 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=3.38
+ $Y=1.84 $X2=3.53 $Y2=2.815
r170 8 67 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=3.38
+ $Y=1.84 $X2=3.53 $Y2=1.985
r171 7 78 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.43
+ $Y=1.84 $X2=2.58 $Y2=1.985
r172 7 57 300 $w=1.7e-07 $l=6.30555e-07 $layer=licon1_PDIFF $count=2 $X=2.43
+ $Y=1.84 $X2=2.58 $Y2=2.4
r173 6 75 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=1.53
+ $Y=1.84 $X2=1.68 $Y2=2.115
r174 6 43 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.53
+ $Y=1.84 $X2=1.68 $Y2=2.815
r175 5 72 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.84 $X2=0.73 $Y2=2.115
r176 5 31 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.84 $X2=0.73 $Y2=2.815
r177 4 63 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.375
+ $Y=0.37 $X2=3.515 $Y2=0.515
r178 3 51 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.375
+ $Y=0.37 $X2=2.515 $Y2=0.515
r179 2 39 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.445
+ $Y=0.37 $X2=1.585 $Y2=0.515
r180 1 27 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.585
+ $Y=0.37 $X2=0.725 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__INV_8%VGND 1 2 3 4 5 16 18 22 26 30 32 34 37 38 40
+ 41 42 44 56 64 68
r67 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r68 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r69 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r70 59 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r71 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r72 56 67 4.55841 $w=1.7e-07 $l=2.7e-07 $layer=LI1_cond $X=3.78 $Y=0 $X2=4.05
+ $Y2=0
r73 56 58 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=3.78 $Y=0 $X2=3.6
+ $Y2=0
r74 55 59 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r75 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r76 52 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r77 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r78 49 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.32 $Y=0 $X2=1.155
+ $Y2=0
r79 49 51 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=1.32 $Y=0 $X2=1.68
+ $Y2=0
r80 48 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r81 48 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r82 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r83 45 61 3.99177 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.38 $Y=0 $X2=0.19
+ $Y2=0
r84 45 47 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.38 $Y=0 $X2=0.72
+ $Y2=0
r85 44 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.99 $Y=0 $X2=1.155
+ $Y2=0
r86 44 47 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.99 $Y=0 $X2=0.72
+ $Y2=0
r87 42 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r88 42 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r89 40 54 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=2.85 $Y=0 $X2=2.64
+ $Y2=0
r90 40 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.85 $Y=0 $X2=3.015
+ $Y2=0
r91 39 58 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=3.18 $Y=0 $X2=3.6
+ $Y2=0
r92 39 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.18 $Y=0 $X2=3.015
+ $Y2=0
r93 37 51 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.85 $Y=0 $X2=1.68
+ $Y2=0
r94 37 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.85 $Y=0 $X2=2.015
+ $Y2=0
r95 36 54 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=2.18 $Y=0 $X2=2.64
+ $Y2=0
r96 36 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.18 $Y=0 $X2=2.015
+ $Y2=0
r97 32 67 3.20777 $w=3.3e-07 $l=1.41244e-07 $layer=LI1_cond $X=3.945 $Y=0.085
+ $X2=4.05 $Y2=0
r98 32 34 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.945 $Y=0.085
+ $X2=3.945 $Y2=0.515
r99 28 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.015 $Y=0.085
+ $X2=3.015 $Y2=0
r100 28 30 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=3.015 $Y=0.085
+ $X2=3.015 $Y2=0.495
r101 24 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.015 $Y=0.085
+ $X2=2.015 $Y2=0
r102 24 26 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=2.015 $Y=0.085
+ $X2=2.015 $Y2=0.675
r103 20 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.155 $Y=0.085
+ $X2=1.155 $Y2=0
r104 20 22 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=1.155 $Y=0.085
+ $X2=1.155 $Y2=0.675
r105 16 61 3.1514 $w=2.5e-07 $l=1.12916e-07 $layer=LI1_cond $X=0.255 $Y=0.085
+ $X2=0.19 $Y2=0
r106 16 18 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.255 $Y=0.085
+ $X2=0.255 $Y2=0.515
r107 5 34 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.805
+ $Y=0.37 $X2=3.945 $Y2=0.515
r108 4 30 91 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=2 $X=2.805
+ $Y=0.37 $X2=3.015 $Y2=0.495
r109 3 26 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=1.875
+ $Y=0.37 $X2=2.015 $Y2=0.675
r110 2 22 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=1.015
+ $Y=0.37 $X2=1.155 $Y2=0.675
r111 1 18 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.15
+ $Y=0.37 $X2=0.295 $Y2=0.515
.ends

