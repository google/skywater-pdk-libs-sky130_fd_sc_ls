* File: sky130_fd_sc_ls__o211a_2.pxi.spice
* Created: Fri Aug 28 13:43:21 2020
* 
x_PM_SKY130_FD_SC_LS__O211A_2%C1 N_C1_c_63_n N_C1_M1004_g N_C1_c_64_n
+ N_C1_M1009_g C1 PM_SKY130_FD_SC_LS__O211A_2%C1
x_PM_SKY130_FD_SC_LS__O211A_2%B1 N_B1_M1002_g N_B1_c_86_n N_B1_M1008_g B1
+ N_B1_c_87_n PM_SKY130_FD_SC_LS__O211A_2%B1
x_PM_SKY130_FD_SC_LS__O211A_2%A2 N_A2_M1007_g N_A2_c_118_n N_A2_M1011_g A2
+ PM_SKY130_FD_SC_LS__O211A_2%A2
x_PM_SKY130_FD_SC_LS__O211A_2%A1 N_A1_c_149_n N_A1_M1005_g N_A1_M1010_g A1
+ N_A1_c_151_n PM_SKY130_FD_SC_LS__O211A_2%A1
x_PM_SKY130_FD_SC_LS__O211A_2%A_27_368# N_A_27_368#_M1009_s N_A_27_368#_M1004_s
+ N_A_27_368#_M1008_d N_A_27_368#_c_190_n N_A_27_368#_M1000_g
+ N_A_27_368#_c_184_n N_A_27_368#_M1001_g N_A_27_368#_c_191_n
+ N_A_27_368#_M1006_g N_A_27_368#_c_185_n N_A_27_368#_M1003_g
+ N_A_27_368#_c_192_n N_A_27_368#_c_193_n N_A_27_368#_c_200_n
+ N_A_27_368#_c_186_n N_A_27_368#_c_194_n N_A_27_368#_c_220_n
+ N_A_27_368#_c_187_n N_A_27_368#_c_195_n N_A_27_368#_c_188_n
+ N_A_27_368#_c_215_n N_A_27_368#_c_189_n PM_SKY130_FD_SC_LS__O211A_2%A_27_368#
x_PM_SKY130_FD_SC_LS__O211A_2%VPWR N_VPWR_M1004_d N_VPWR_M1005_d N_VPWR_M1006_d
+ N_VPWR_c_299_n N_VPWR_c_300_n N_VPWR_c_301_n N_VPWR_c_302_n VPWR
+ N_VPWR_c_303_n N_VPWR_c_304_n N_VPWR_c_305_n N_VPWR_c_306_n N_VPWR_c_307_n
+ N_VPWR_c_298_n PM_SKY130_FD_SC_LS__O211A_2%VPWR
x_PM_SKY130_FD_SC_LS__O211A_2%X N_X_M1001_d N_X_M1000_s N_X_c_350_n N_X_c_351_n
+ N_X_c_347_n X X X X X PM_SKY130_FD_SC_LS__O211A_2%X
x_PM_SKY130_FD_SC_LS__O211A_2%A_195_74# N_A_195_74#_M1002_d N_A_195_74#_M1010_d
+ N_A_195_74#_c_383_n N_A_195_74#_c_380_n N_A_195_74#_c_381_n
+ PM_SKY130_FD_SC_LS__O211A_2%A_195_74#
x_PM_SKY130_FD_SC_LS__O211A_2%VGND N_VGND_M1007_d N_VGND_M1001_s N_VGND_M1003_s
+ N_VGND_c_407_n N_VGND_c_408_n N_VGND_c_409_n N_VGND_c_410_n VGND
+ N_VGND_c_411_n N_VGND_c_412_n N_VGND_c_413_n N_VGND_c_414_n N_VGND_c_415_n
+ N_VGND_c_416_n PM_SKY130_FD_SC_LS__O211A_2%VGND
cc_1 VNB N_C1_c_63_n 0.0670849f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.765
cc_2 VNB N_C1_c_64_n 0.0226984f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.22
cc_3 VNB C1 0.00891253f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_B1_M1002_g 0.0246592f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.34
cc_5 VNB N_B1_c_86_n 0.0217744f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.74
cc_6 VNB N_B1_c_87_n 0.00613118f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.295
cc_7 VNB N_A2_M1007_g 0.0267529f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.34
cc_8 VNB N_A2_c_118_n 0.0216741f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.74
cc_9 VNB A2 0.00508898f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A1_c_149_n 0.0317625f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.765
cc_11 VNB N_A1_M1010_g 0.0290764f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.74
cc_12 VNB N_A1_c_151_n 0.00231998f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.295
cc_13 VNB N_A_27_368#_c_184_n 0.0161558f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_368#_c_185_n 0.0184695f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_368#_c_186_n 0.0284016f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_27_368#_c_187_n 0.00677368f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_27_368#_c_188_n 0.0341051f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_27_368#_c_189_n 0.096444f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_VPWR_c_298_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_X_c_347_n 5.40438e-19 $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_21 VNB X 0.00210995f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB X 8.99291e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_195_74#_c_380_n 0.0028557f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_24 VNB N_A_195_74#_c_381_n 0.00734199f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_25 VNB N_VGND_c_407_n 0.00560579f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.295
cc_26 VNB N_VGND_c_408_n 0.0129885f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_409_n 0.0115487f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_410_n 0.0510963f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_411_n 0.0423577f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_412_n 0.0210122f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_413_n 0.0172134f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_414_n 0.00477896f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_415_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_416_n 0.236934f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VPB N_C1_c_63_n 0.0308401f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.765
cc_36 VPB N_B1_c_86_n 0.0263273f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=0.74
cc_37 VPB N_B1_c_87_n 0.00549423f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.295
cc_38 VPB N_A2_c_118_n 0.0256896f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=0.74
cc_39 VPB A2 0.00438576f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_40 VPB N_A1_c_149_n 0.0312161f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.765
cc_41 VPB N_A1_c_151_n 0.0030812f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.295
cc_42 VPB N_A_27_368#_c_190_n 0.0169399f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_43 VPB N_A_27_368#_c_191_n 0.0174014f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_44 VPB N_A_27_368#_c_192_n 0.014539f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_45 VPB N_A_27_368#_c_193_n 0.0316952f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_A_27_368#_c_194_n 0.00324157f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB N_A_27_368#_c_195_n 0.00197537f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 VPB N_A_27_368#_c_189_n 0.0265046f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_299_n 0.0198253f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.295
cc_50 VPB N_VPWR_c_300_n 0.0163777f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_301_n 0.0121909f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_302_n 0.0685555f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_303_n 0.0193716f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_304_n 0.0325718f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_305_n 0.0186948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_306_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_307_n 0.0134384f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_298_n 0.0813545f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_X_c_350_n 0.00341966f $X=-0.19 $Y=1.66 $X2=0.345 $Y2=1.385
cc_60 VPB N_X_c_351_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_61 VPB N_X_c_347_n 0.00116518f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_62 N_C1_c_64_n N_B1_M1002_g 0.0568681f $X=0.51 $Y=1.22 $X2=0 $Y2=0
cc_63 C1 N_B1_M1002_g 6.12064e-19 $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_64 N_C1_c_63_n N_B1_c_86_n 0.0455697f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_65 N_C1_c_63_n N_B1_c_87_n 0.00878524f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_66 C1 N_B1_c_87_n 0.0164128f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_67 N_C1_c_63_n N_A_27_368#_c_192_n 0.00608673f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_68 C1 N_A_27_368#_c_192_n 0.0197435f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_69 N_C1_c_63_n N_A_27_368#_c_193_n 0.00933129f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_70 N_C1_c_63_n N_A_27_368#_c_200_n 0.0165f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_71 N_C1_c_63_n N_A_27_368#_c_194_n 6.30044e-19 $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_72 N_C1_c_63_n N_A_27_368#_c_188_n 0.00198616f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_73 N_C1_c_64_n N_A_27_368#_c_188_n 0.0264367f $X=0.51 $Y=1.22 $X2=0 $Y2=0
cc_74 C1 N_A_27_368#_c_188_n 0.0241619f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_75 N_C1_c_63_n N_VPWR_c_299_n 0.00660268f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_76 N_C1_c_63_n N_VPWR_c_303_n 0.00481995f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_77 N_C1_c_63_n N_VPWR_c_298_n 0.00508379f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_78 N_C1_c_64_n N_VGND_c_411_n 0.00291513f $X=0.51 $Y=1.22 $X2=0 $Y2=0
cc_79 N_C1_c_64_n N_VGND_c_416_n 0.00362434f $X=0.51 $Y=1.22 $X2=0 $Y2=0
cc_80 N_B1_M1002_g N_A2_M1007_g 0.0298942f $X=0.9 $Y=0.74 $X2=0 $Y2=0
cc_81 N_B1_c_86_n N_A2_c_118_n 0.033955f $X=1.035 $Y=1.765 $X2=0 $Y2=0
cc_82 N_B1_c_87_n N_A2_c_118_n 5.5756e-19 $X=0.96 $Y=1.515 $X2=0 $Y2=0
cc_83 N_B1_c_86_n A2 8.00115e-19 $X=1.035 $Y=1.765 $X2=0 $Y2=0
cc_84 N_B1_c_87_n A2 0.0295439f $X=0.96 $Y=1.515 $X2=0 $Y2=0
cc_85 N_B1_c_86_n N_A_27_368#_c_192_n 5.93323e-19 $X=1.035 $Y=1.765 $X2=0 $Y2=0
cc_86 N_B1_c_86_n N_A_27_368#_c_193_n 3.81051e-19 $X=1.035 $Y=1.765 $X2=0 $Y2=0
cc_87 N_B1_c_86_n N_A_27_368#_c_200_n 0.0138784f $X=1.035 $Y=1.765 $X2=0 $Y2=0
cc_88 N_B1_c_87_n N_A_27_368#_c_200_n 0.0359529f $X=0.96 $Y=1.515 $X2=0 $Y2=0
cc_89 N_B1_M1002_g N_A_27_368#_c_186_n 0.0147907f $X=0.9 $Y=0.74 $X2=0 $Y2=0
cc_90 N_B1_c_86_n N_A_27_368#_c_186_n 0.00458387f $X=1.035 $Y=1.765 $X2=0 $Y2=0
cc_91 N_B1_c_87_n N_A_27_368#_c_186_n 0.0263338f $X=0.96 $Y=1.515 $X2=0 $Y2=0
cc_92 N_B1_c_86_n N_A_27_368#_c_194_n 0.00849717f $X=1.035 $Y=1.765 $X2=0 $Y2=0
cc_93 N_B1_M1002_g N_A_27_368#_c_188_n 0.00255489f $X=0.9 $Y=0.74 $X2=0 $Y2=0
cc_94 N_B1_c_87_n N_A_27_368#_c_188_n 0.0153286f $X=0.96 $Y=1.515 $X2=0 $Y2=0
cc_95 N_B1_c_87_n N_A_27_368#_c_215_n 0.00101752f $X=0.96 $Y=1.515 $X2=0 $Y2=0
cc_96 N_B1_c_86_n N_VPWR_c_299_n 0.0034425f $X=1.035 $Y=1.765 $X2=0 $Y2=0
cc_97 N_B1_c_86_n N_VPWR_c_304_n 0.00490606f $X=1.035 $Y=1.765 $X2=0 $Y2=0
cc_98 N_B1_c_86_n N_VPWR_c_298_n 0.00508379f $X=1.035 $Y=1.765 $X2=0 $Y2=0
cc_99 N_B1_M1002_g N_A_195_74#_c_380_n 0.00267731f $X=0.9 $Y=0.74 $X2=0 $Y2=0
cc_100 N_B1_M1002_g N_VGND_c_411_n 0.00461464f $X=0.9 $Y=0.74 $X2=0 $Y2=0
cc_101 N_B1_M1002_g N_VGND_c_416_n 0.00909821f $X=0.9 $Y=0.74 $X2=0 $Y2=0
cc_102 N_A2_c_118_n N_A1_c_149_n 0.0696068f $X=1.495 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_103 A2 N_A1_c_149_n 0.00312363f $X=1.595 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_104 N_A2_M1007_g N_A1_M1010_g 0.0308987f $X=1.41 $Y=0.74 $X2=0 $Y2=0
cc_105 N_A2_c_118_n N_A1_c_151_n 3.56421e-19 $X=1.495 $Y=1.765 $X2=0 $Y2=0
cc_106 A2 N_A1_c_151_n 0.0349136f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_107 N_A2_M1007_g N_A_27_368#_c_186_n 0.0114661f $X=1.41 $Y=0.74 $X2=0 $Y2=0
cc_108 N_A2_c_118_n N_A_27_368#_c_186_n 0.00438688f $X=1.495 $Y=1.765 $X2=0
+ $Y2=0
cc_109 A2 N_A_27_368#_c_186_n 0.0352799f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_110 N_A2_c_118_n N_A_27_368#_c_194_n 0.0137081f $X=1.495 $Y=1.765 $X2=0 $Y2=0
cc_111 N_A2_c_118_n N_A_27_368#_c_220_n 0.0124263f $X=1.495 $Y=1.765 $X2=0 $Y2=0
cc_112 A2 N_A_27_368#_c_220_n 0.0256676f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_113 N_A2_c_118_n N_A_27_368#_c_215_n 7.48251e-19 $X=1.495 $Y=1.765 $X2=0
+ $Y2=0
cc_114 A2 N_A_27_368#_c_215_n 0.00613412f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_115 N_A2_c_118_n N_VPWR_c_300_n 0.00220919f $X=1.495 $Y=1.765 $X2=0 $Y2=0
cc_116 N_A2_c_118_n N_VPWR_c_304_n 0.00481995f $X=1.495 $Y=1.765 $X2=0 $Y2=0
cc_117 N_A2_c_118_n N_VPWR_c_298_n 0.00508379f $X=1.495 $Y=1.765 $X2=0 $Y2=0
cc_118 N_A2_M1007_g N_A_195_74#_c_383_n 0.00989989f $X=1.41 $Y=0.74 $X2=0 $Y2=0
cc_119 N_A2_M1007_g N_A_195_74#_c_380_n 0.00739554f $X=1.41 $Y=0.74 $X2=0 $Y2=0
cc_120 N_A2_M1007_g N_A_195_74#_c_381_n 6.56032e-19 $X=1.41 $Y=0.74 $X2=0 $Y2=0
cc_121 N_A2_M1007_g N_VGND_c_407_n 0.00400267f $X=1.41 $Y=0.74 $X2=0 $Y2=0
cc_122 N_A2_M1007_g N_VGND_c_411_n 0.00325937f $X=1.41 $Y=0.74 $X2=0 $Y2=0
cc_123 N_A2_M1007_g N_VGND_c_416_n 0.00413498f $X=1.41 $Y=0.74 $X2=0 $Y2=0
cc_124 N_A1_c_149_n N_A_27_368#_c_190_n 0.00869429f $X=1.965 $Y=1.765 $X2=0
+ $Y2=0
cc_125 N_A1_c_149_n N_A_27_368#_c_186_n 0.00254235f $X=1.965 $Y=1.765 $X2=0
+ $Y2=0
cc_126 N_A1_M1010_g N_A_27_368#_c_186_n 0.0151825f $X=1.97 $Y=0.74 $X2=0 $Y2=0
cc_127 N_A1_c_151_n N_A_27_368#_c_186_n 0.0249861f $X=2.13 $Y=1.515 $X2=0 $Y2=0
cc_128 N_A1_c_149_n N_A_27_368#_c_194_n 0.00250227f $X=1.965 $Y=1.765 $X2=0
+ $Y2=0
cc_129 N_A1_c_149_n N_A_27_368#_c_220_n 0.019788f $X=1.965 $Y=1.765 $X2=0 $Y2=0
cc_130 N_A1_c_151_n N_A_27_368#_c_220_n 0.0236735f $X=2.13 $Y=1.515 $X2=0 $Y2=0
cc_131 N_A1_c_149_n N_A_27_368#_c_187_n 0.00102181f $X=1.965 $Y=1.765 $X2=0
+ $Y2=0
cc_132 N_A1_M1010_g N_A_27_368#_c_187_n 0.00103826f $X=1.97 $Y=0.74 $X2=0 $Y2=0
cc_133 N_A1_c_151_n N_A_27_368#_c_187_n 0.0178205f $X=2.13 $Y=1.515 $X2=0 $Y2=0
cc_134 N_A1_c_149_n N_A_27_368#_c_195_n 0.00325521f $X=1.965 $Y=1.765 $X2=0
+ $Y2=0
cc_135 N_A1_c_151_n N_A_27_368#_c_195_n 0.00964976f $X=2.13 $Y=1.515 $X2=0 $Y2=0
cc_136 N_A1_c_149_n N_A_27_368#_c_189_n 0.0225204f $X=1.965 $Y=1.765 $X2=0 $Y2=0
cc_137 N_A1_M1010_g N_A_27_368#_c_189_n 0.00356504f $X=1.97 $Y=0.74 $X2=0 $Y2=0
cc_138 N_A1_c_151_n N_A_27_368#_c_189_n 9.27871e-19 $X=2.13 $Y=1.515 $X2=0 $Y2=0
cc_139 N_A1_c_149_n N_VPWR_c_300_n 0.0155728f $X=1.965 $Y=1.765 $X2=0 $Y2=0
cc_140 N_A1_c_149_n N_VPWR_c_304_n 0.00443511f $X=1.965 $Y=1.765 $X2=0 $Y2=0
cc_141 N_A1_c_149_n N_VPWR_c_298_n 0.00460931f $X=1.965 $Y=1.765 $X2=0 $Y2=0
cc_142 N_A1_M1010_g N_A_195_74#_c_383_n 0.00966375f $X=1.97 $Y=0.74 $X2=0 $Y2=0
cc_143 N_A1_M1010_g N_A_195_74#_c_380_n 6.37625e-19 $X=1.97 $Y=0.74 $X2=0 $Y2=0
cc_144 N_A1_M1010_g N_A_195_74#_c_381_n 0.00876423f $X=1.97 $Y=0.74 $X2=0 $Y2=0
cc_145 N_A1_M1010_g N_VGND_c_407_n 0.0040624f $X=1.97 $Y=0.74 $X2=0 $Y2=0
cc_146 N_A1_M1010_g N_VGND_c_408_n 0.00369425f $X=1.97 $Y=0.74 $X2=0 $Y2=0
cc_147 N_A1_M1010_g N_VGND_c_412_n 0.00324657f $X=1.97 $Y=0.74 $X2=0 $Y2=0
cc_148 N_A1_M1010_g N_VGND_c_416_n 0.00416919f $X=1.97 $Y=0.74 $X2=0 $Y2=0
cc_149 N_A_27_368#_c_200_n N_VPWR_M1004_d 0.0059417f $X=1.105 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_150 N_A_27_368#_c_220_n N_VPWR_M1005_d 0.0217482f $X=2.505 $Y=2.035 $X2=0
+ $Y2=0
cc_151 N_A_27_368#_c_195_n N_VPWR_M1005_d 0.00302199f $X=2.59 $Y=1.95 $X2=0
+ $Y2=0
cc_152 N_A_27_368#_c_193_n N_VPWR_c_299_n 0.0221782f $X=0.27 $Y=2.695 $X2=0
+ $Y2=0
cc_153 N_A_27_368#_c_200_n N_VPWR_c_299_n 0.022455f $X=1.105 $Y=2.035 $X2=0
+ $Y2=0
cc_154 N_A_27_368#_c_194_n N_VPWR_c_299_n 0.0221782f $X=1.27 $Y=2.715 $X2=0
+ $Y2=0
cc_155 N_A_27_368#_c_190_n N_VPWR_c_300_n 0.0101725f $X=2.835 $Y=1.765 $X2=0
+ $Y2=0
cc_156 N_A_27_368#_c_194_n N_VPWR_c_300_n 0.0162323f $X=1.27 $Y=2.715 $X2=0
+ $Y2=0
cc_157 N_A_27_368#_c_220_n N_VPWR_c_300_n 0.0494195f $X=2.505 $Y=2.035 $X2=0
+ $Y2=0
cc_158 N_A_27_368#_c_187_n N_VPWR_c_300_n 0.00104666f $X=2.59 $Y=1.63 $X2=0
+ $Y2=0
cc_159 N_A_27_368#_c_189_n N_VPWR_c_300_n 0.0014794f $X=3.285 $Y=1.475 $X2=0
+ $Y2=0
cc_160 N_A_27_368#_c_191_n N_VPWR_c_302_n 0.0261486f $X=3.285 $Y=1.765 $X2=0
+ $Y2=0
cc_161 N_A_27_368#_c_189_n N_VPWR_c_302_n 0.00135549f $X=3.285 $Y=1.475 $X2=0
+ $Y2=0
cc_162 N_A_27_368#_c_193_n N_VPWR_c_303_n 0.0097982f $X=0.27 $Y=2.695 $X2=0
+ $Y2=0
cc_163 N_A_27_368#_c_194_n N_VPWR_c_304_n 0.00978791f $X=1.27 $Y=2.715 $X2=0
+ $Y2=0
cc_164 N_A_27_368#_c_190_n N_VPWR_c_305_n 0.00445602f $X=2.835 $Y=1.765 $X2=0
+ $Y2=0
cc_165 N_A_27_368#_c_191_n N_VPWR_c_305_n 0.00445602f $X=3.285 $Y=1.765 $X2=0
+ $Y2=0
cc_166 N_A_27_368#_c_190_n N_VPWR_c_298_n 0.00861719f $X=2.835 $Y=1.765 $X2=0
+ $Y2=0
cc_167 N_A_27_368#_c_191_n N_VPWR_c_298_n 0.00860566f $X=3.285 $Y=1.765 $X2=0
+ $Y2=0
cc_168 N_A_27_368#_c_193_n N_VPWR_c_298_n 0.0111907f $X=0.27 $Y=2.695 $X2=0
+ $Y2=0
cc_169 N_A_27_368#_c_194_n N_VPWR_c_298_n 0.0111866f $X=1.27 $Y=2.715 $X2=0
+ $Y2=0
cc_170 N_A_27_368#_c_220_n A_314_368# 0.0110255f $X=2.505 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_171 N_A_27_368#_c_190_n N_X_c_350_n 0.00282707f $X=2.835 $Y=1.765 $X2=0 $Y2=0
cc_172 N_A_27_368#_c_191_n N_X_c_350_n 0.00188635f $X=3.285 $Y=1.765 $X2=0 $Y2=0
cc_173 N_A_27_368#_c_220_n N_X_c_350_n 0.0114771f $X=2.505 $Y=2.035 $X2=0 $Y2=0
cc_174 N_A_27_368#_c_195_n N_X_c_350_n 0.00786832f $X=2.59 $Y=1.95 $X2=0 $Y2=0
cc_175 N_A_27_368#_c_189_n N_X_c_350_n 8.22785e-19 $X=3.285 $Y=1.475 $X2=0 $Y2=0
cc_176 N_A_27_368#_c_190_n N_X_c_351_n 0.0166285f $X=2.835 $Y=1.765 $X2=0 $Y2=0
cc_177 N_A_27_368#_c_191_n N_X_c_351_n 0.0109216f $X=3.285 $Y=1.765 $X2=0 $Y2=0
cc_178 N_A_27_368#_c_190_n N_X_c_347_n 4.87241e-19 $X=2.835 $Y=1.765 $X2=0 $Y2=0
cc_179 N_A_27_368#_c_191_n N_X_c_347_n 0.00264043f $X=3.285 $Y=1.765 $X2=0 $Y2=0
cc_180 N_A_27_368#_c_195_n N_X_c_347_n 0.00878595f $X=2.59 $Y=1.95 $X2=0 $Y2=0
cc_181 N_A_27_368#_c_189_n N_X_c_347_n 0.0260629f $X=3.285 $Y=1.475 $X2=0 $Y2=0
cc_182 N_A_27_368#_c_184_n X 0.0131366f $X=2.93 $Y=1.185 $X2=0 $Y2=0
cc_183 N_A_27_368#_c_185_n X 0.00191951f $X=3.36 $Y=1.185 $X2=0 $Y2=0
cc_184 N_A_27_368#_c_184_n X 0.00341227f $X=2.93 $Y=1.185 $X2=0 $Y2=0
cc_185 N_A_27_368#_c_187_n X 0.00625242f $X=2.59 $Y=1.63 $X2=0 $Y2=0
cc_186 N_A_27_368#_c_184_n X 5.79411e-19 $X=2.93 $Y=1.185 $X2=0 $Y2=0
cc_187 N_A_27_368#_c_187_n X 0.0319634f $X=2.59 $Y=1.63 $X2=0 $Y2=0
cc_188 N_A_27_368#_c_189_n X 0.0205638f $X=3.285 $Y=1.475 $X2=0 $Y2=0
cc_189 N_A_27_368#_c_186_n N_A_195_74#_M1002_d 0.00261503f $X=2.505 $Y=1.095
+ $X2=-0.19 $Y2=-0.245
cc_190 N_A_27_368#_c_186_n N_A_195_74#_M1010_d 0.0027574f $X=2.505 $Y=1.095
+ $X2=0 $Y2=0
cc_191 N_A_27_368#_c_186_n N_A_195_74#_c_383_n 0.0387834f $X=2.505 $Y=1.095
+ $X2=0 $Y2=0
cc_192 N_A_27_368#_c_186_n N_A_195_74#_c_380_n 0.0208988f $X=2.505 $Y=1.095
+ $X2=0 $Y2=0
cc_193 N_A_27_368#_c_188_n N_A_195_74#_c_380_n 0.0012754f $X=0.295 $Y=0.515
+ $X2=0 $Y2=0
cc_194 N_A_27_368#_c_186_n N_A_195_74#_c_381_n 0.0214503f $X=2.505 $Y=1.095
+ $X2=0 $Y2=0
cc_195 N_A_27_368#_c_186_n N_VGND_M1007_d 0.00342819f $X=2.505 $Y=1.095
+ $X2=-0.19 $Y2=-0.245
cc_196 N_A_27_368#_c_187_n N_VGND_M1001_s 0.00210817f $X=2.59 $Y=1.63 $X2=0
+ $Y2=0
cc_197 N_A_27_368#_c_184_n N_VGND_c_408_n 0.00505083f $X=2.93 $Y=1.185 $X2=0
+ $Y2=0
cc_198 N_A_27_368#_c_187_n N_VGND_c_408_n 0.016027f $X=2.59 $Y=1.63 $X2=0 $Y2=0
cc_199 N_A_27_368#_c_189_n N_VGND_c_408_n 0.00368888f $X=3.285 $Y=1.475 $X2=0
+ $Y2=0
cc_200 N_A_27_368#_c_184_n N_VGND_c_410_n 6.08778e-19 $X=2.93 $Y=1.185 $X2=0
+ $Y2=0
cc_201 N_A_27_368#_c_185_n N_VGND_c_410_n 0.015817f $X=3.36 $Y=1.185 $X2=0 $Y2=0
cc_202 N_A_27_368#_c_188_n N_VGND_c_411_n 0.0282878f $X=0.295 $Y=0.515 $X2=0
+ $Y2=0
cc_203 N_A_27_368#_c_184_n N_VGND_c_413_n 0.00434272f $X=2.93 $Y=1.185 $X2=0
+ $Y2=0
cc_204 N_A_27_368#_c_185_n N_VGND_c_413_n 0.00383152f $X=3.36 $Y=1.185 $X2=0
+ $Y2=0
cc_205 N_A_27_368#_c_184_n N_VGND_c_416_n 0.00825283f $X=2.93 $Y=1.185 $X2=0
+ $Y2=0
cc_206 N_A_27_368#_c_185_n N_VGND_c_416_n 0.0075754f $X=3.36 $Y=1.185 $X2=0
+ $Y2=0
cc_207 N_A_27_368#_c_188_n N_VGND_c_416_n 0.0230808f $X=0.295 $Y=0.515 $X2=0
+ $Y2=0
cc_208 N_VPWR_c_302_n N_X_c_350_n 0.0450694f $X=3.56 $Y=1.985 $X2=0 $Y2=0
cc_209 N_VPWR_c_300_n N_X_c_351_n 0.026776f $X=2.56 $Y=2.375 $X2=0 $Y2=0
cc_210 N_VPWR_c_305_n N_X_c_351_n 0.014552f $X=3.395 $Y=3.33 $X2=0 $Y2=0
cc_211 N_VPWR_c_298_n N_X_c_351_n 0.0119791f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_212 X N_VGND_c_408_n 0.0176099f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_213 X N_VGND_c_410_n 0.0300842f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_214 X N_VGND_c_413_n 0.0112174f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_215 X N_VGND_c_416_n 0.00922837f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_216 N_A_195_74#_c_383_n N_VGND_M1007_d 0.0070032f $X=2.02 $Y=0.755 $X2=-0.19
+ $Y2=-0.245
cc_217 N_A_195_74#_c_383_n N_VGND_c_407_n 0.017876f $X=2.02 $Y=0.755 $X2=0 $Y2=0
cc_218 N_A_195_74#_c_380_n N_VGND_c_407_n 0.00638631f $X=1.19 $Y=0.595 $X2=0
+ $Y2=0
cc_219 N_A_195_74#_c_381_n N_VGND_c_407_n 0.00861021f $X=2.185 $Y=0.595 $X2=0
+ $Y2=0
cc_220 N_A_195_74#_c_381_n N_VGND_c_408_n 0.035653f $X=2.185 $Y=0.595 $X2=0
+ $Y2=0
cc_221 N_A_195_74#_c_383_n N_VGND_c_411_n 0.00230811f $X=2.02 $Y=0.755 $X2=0
+ $Y2=0
cc_222 N_A_195_74#_c_380_n N_VGND_c_411_n 0.0142392f $X=1.19 $Y=0.595 $X2=0
+ $Y2=0
cc_223 N_A_195_74#_c_383_n N_VGND_c_412_n 0.00340448f $X=2.02 $Y=0.755 $X2=0
+ $Y2=0
cc_224 N_A_195_74#_c_381_n N_VGND_c_412_n 0.0142249f $X=2.185 $Y=0.595 $X2=0
+ $Y2=0
cc_225 N_A_195_74#_c_383_n N_VGND_c_416_n 0.0113875f $X=2.02 $Y=0.755 $X2=0
+ $Y2=0
cc_226 N_A_195_74#_c_380_n N_VGND_c_416_n 0.0118911f $X=1.19 $Y=0.595 $X2=0
+ $Y2=0
cc_227 N_A_195_74#_c_381_n N_VGND_c_416_n 0.011867f $X=2.185 $Y=0.595 $X2=0
+ $Y2=0
