# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ls__sdfrtp_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ls__sdfrtp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  14.40000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 0.810000 2.100000 1.265000 ;
        RECT 1.605000 0.595000 2.100000 0.810000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.525000 0.350000 13.855000 1.410000 ;
        RECT 13.525000 1.410000 13.785000 2.980000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.411000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  3.785000 1.830000  4.165000 2.160000 ;
        RECT  3.920000 2.160000  4.165000 2.190000 ;
        RECT  7.775000 1.795000  8.570000 2.150000 ;
        RECT 11.110000 1.920000 11.440000 2.220000 ;
      LAYER mcon ;
        RECT  3.995000 1.950000  4.165000 2.120000 ;
        RECT  8.315000 1.950000  8.485000 2.120000 ;
        RECT 11.195000 1.950000 11.365000 2.120000 ;
      LAYER met1 ;
        RECT  3.935000 1.920000  4.225000 1.965000 ;
        RECT  3.935000 1.965000 11.425000 2.105000 ;
        RECT  3.935000 2.105000  4.225000 2.150000 ;
        RECT  8.255000 1.920000  8.545000 1.965000 ;
        RECT  8.255000 2.105000  8.545000 2.150000 ;
        RECT 11.135000 1.920000 11.425000 1.965000 ;
        RECT 11.135000 2.105000 11.425000 2.150000 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.875000 2.000000 3.275000 2.175000 ;
        RECT 2.945000 1.440000 3.275000 2.000000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.455000 1.490000 2.705000 1.660000 ;
        RECT 0.455000 1.660000 2.205000 1.835000 ;
        RECT 2.375000 1.260000 2.705000 1.490000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.785000 0.920000 4.060000 1.180000 ;
        RECT 3.785000 1.180000 4.195000 1.260000 ;
        RECT 3.785000 1.260000 4.645000 1.630000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 14.400000 0.085000 ;
        RECT  0.545000  0.085000  0.875000 0.765000 ;
        RECT  3.610000  0.085000  3.880000 0.730000 ;
        RECT  4.705000  0.085000  5.035000 0.710000 ;
        RECT  7.430000  0.085000  7.760000 0.410000 ;
        RECT 10.755000  0.085000 11.085000 0.810000 ;
        RECT 12.105000  0.085000 12.435000 0.600000 ;
        RECT 13.095000  0.085000 13.345000 1.130000 ;
        RECT 14.035000  0.085000 14.285000 1.130000 ;
      LAYER mcon ;
        RECT  0.155000 -0.085000  0.325000 0.085000 ;
        RECT  0.635000 -0.085000  0.805000 0.085000 ;
        RECT  1.115000 -0.085000  1.285000 0.085000 ;
        RECT  1.595000 -0.085000  1.765000 0.085000 ;
        RECT  2.075000 -0.085000  2.245000 0.085000 ;
        RECT  2.555000 -0.085000  2.725000 0.085000 ;
        RECT  3.035000 -0.085000  3.205000 0.085000 ;
        RECT  3.515000 -0.085000  3.685000 0.085000 ;
        RECT  3.995000 -0.085000  4.165000 0.085000 ;
        RECT  4.475000 -0.085000  4.645000 0.085000 ;
        RECT  4.955000 -0.085000  5.125000 0.085000 ;
        RECT  5.435000 -0.085000  5.605000 0.085000 ;
        RECT  5.915000 -0.085000  6.085000 0.085000 ;
        RECT  6.395000 -0.085000  6.565000 0.085000 ;
        RECT  6.875000 -0.085000  7.045000 0.085000 ;
        RECT  7.355000 -0.085000  7.525000 0.085000 ;
        RECT  7.835000 -0.085000  8.005000 0.085000 ;
        RECT  8.315000 -0.085000  8.485000 0.085000 ;
        RECT  8.795000 -0.085000  8.965000 0.085000 ;
        RECT  9.275000 -0.085000  9.445000 0.085000 ;
        RECT  9.755000 -0.085000  9.925000 0.085000 ;
        RECT 10.235000 -0.085000 10.405000 0.085000 ;
        RECT 10.715000 -0.085000 10.885000 0.085000 ;
        RECT 11.195000 -0.085000 11.365000 0.085000 ;
        RECT 11.675000 -0.085000 11.845000 0.085000 ;
        RECT 12.155000 -0.085000 12.325000 0.085000 ;
        RECT 12.635000 -0.085000 12.805000 0.085000 ;
        RECT 13.115000 -0.085000 13.285000 0.085000 ;
        RECT 13.595000 -0.085000 13.765000 0.085000 ;
        RECT 14.075000 -0.085000 14.245000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 14.400000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 3.245000 14.400000 3.415000 ;
        RECT  0.615000 2.345000  1.565000 3.245000 ;
        RECT  3.095000 2.685000  3.425000 3.245000 ;
        RECT  4.705000 2.750000  5.035000 3.245000 ;
        RECT  7.025000 2.345000  7.265000 3.245000 ;
        RECT  8.245000 2.330000  8.580000 3.245000 ;
        RECT 10.560000 2.730000 11.240000 3.245000 ;
        RECT 11.945000 1.940000 12.275000 3.245000 ;
        RECT 13.005000 1.820000 13.335000 3.245000 ;
        RECT 13.955000 1.820000 14.285000 3.245000 ;
      LAYER mcon ;
        RECT  0.155000 3.245000  0.325000 3.415000 ;
        RECT  0.635000 3.245000  0.805000 3.415000 ;
        RECT  1.115000 3.245000  1.285000 3.415000 ;
        RECT  1.595000 3.245000  1.765000 3.415000 ;
        RECT  2.075000 3.245000  2.245000 3.415000 ;
        RECT  2.555000 3.245000  2.725000 3.415000 ;
        RECT  3.035000 3.245000  3.205000 3.415000 ;
        RECT  3.515000 3.245000  3.685000 3.415000 ;
        RECT  3.995000 3.245000  4.165000 3.415000 ;
        RECT  4.475000 3.245000  4.645000 3.415000 ;
        RECT  4.955000 3.245000  5.125000 3.415000 ;
        RECT  5.435000 3.245000  5.605000 3.415000 ;
        RECT  5.915000 3.245000  6.085000 3.415000 ;
        RECT  6.395000 3.245000  6.565000 3.415000 ;
        RECT  6.875000 3.245000  7.045000 3.415000 ;
        RECT  7.355000 3.245000  7.525000 3.415000 ;
        RECT  7.835000 3.245000  8.005000 3.415000 ;
        RECT  8.315000 3.245000  8.485000 3.415000 ;
        RECT  8.795000 3.245000  8.965000 3.415000 ;
        RECT  9.275000 3.245000  9.445000 3.415000 ;
        RECT  9.755000 3.245000  9.925000 3.415000 ;
        RECT 10.235000 3.245000 10.405000 3.415000 ;
        RECT 10.715000 3.245000 10.885000 3.415000 ;
        RECT 11.195000 3.245000 11.365000 3.415000 ;
        RECT 11.675000 3.245000 11.845000 3.415000 ;
        RECT 12.155000 3.245000 12.325000 3.415000 ;
        RECT 12.635000 3.245000 12.805000 3.415000 ;
        RECT 13.115000 3.245000 13.285000 3.415000 ;
        RECT 13.595000 3.245000 13.765000 3.415000 ;
        RECT 14.075000 3.245000 14.245000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 14.400000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.115000 0.350000  0.365000 0.935000 ;
      RECT  0.115000 0.935000  1.140000 1.265000 ;
      RECT  0.115000 1.265000  0.285000 2.005000 ;
      RECT  0.115000 2.005000  2.705000 2.175000 ;
      RECT  0.115000 2.175000  0.445000 2.980000 ;
      RECT  1.105000 0.255000  3.430000 0.425000 ;
      RECT  1.105000 0.425000  1.435000 0.640000 ;
      RECT  2.095000 2.345000  3.785000 2.385000 ;
      RECT  2.095000 2.385000  4.230000 2.400000 ;
      RECT  2.095000 2.400000  4.250000 2.420000 ;
      RECT  2.095000 2.420000  6.075000 2.515000 ;
      RECT  2.095000 2.515000  2.425000 2.980000 ;
      RECT  2.270000 0.595000  3.020000 0.810000 ;
      RECT  2.270000 0.810000  3.040000 0.835000 ;
      RECT  2.270000 0.835000  3.055000 0.845000 ;
      RECT  2.375000 1.830000  2.705000 2.005000 ;
      RECT  2.785000 0.845000  3.055000 0.855000 ;
      RECT  2.785000 0.855000  3.065000 0.865000 ;
      RECT  2.810000 0.865000  3.085000 0.880000 ;
      RECT  2.830000 0.880000  3.110000 0.890000 ;
      RECT  2.840000 0.890000  3.110000 0.900000 ;
      RECT  2.840000 0.900000  3.615000 0.910000 ;
      RECT  2.855000 0.910000  3.615000 0.935000 ;
      RECT  2.875000 0.935000  3.615000 1.270000 ;
      RECT  3.190000 0.425000  3.430000 0.730000 ;
      RECT  3.445000 1.270000  3.615000 2.330000 ;
      RECT  3.445000 2.330000  3.785000 2.345000 ;
      RECT  3.615000 2.515000  6.075000 2.580000 ;
      RECT  3.615000 2.580000  4.645000 2.585000 ;
      RECT  3.615000 2.585000  4.630000 2.590000 ;
      RECT  3.615000 2.590000  4.610000 2.600000 ;
      RECT  3.615000 2.600000  4.580000 2.620000 ;
      RECT  3.615000 2.620000  3.995000 2.980000 ;
      RECT  4.135000 0.500000  4.535000 0.750000 ;
      RECT  4.230000 0.750000  4.535000 0.790000 ;
      RECT  4.230000 0.790000  4.555000 0.815000 ;
      RECT  4.230000 0.815000  4.570000 0.835000 ;
      RECT  4.230000 0.835000  4.580000 0.845000 ;
      RECT  4.300000 0.845000  4.600000 0.860000 ;
      RECT  4.300000 0.860000  4.625000 0.865000 ;
      RECT  4.325000 0.865000  4.625000 0.880000 ;
      RECT  4.335000 1.820000  4.985000 2.195000 ;
      RECT  4.335000 2.195000  4.505000 2.250000 ;
      RECT  4.345000 0.880000  5.045000 0.890000 ;
      RECT  4.355000 0.890000  5.045000 0.910000 ;
      RECT  4.370000 0.910000  5.045000 0.935000 ;
      RECT  4.390000 0.935000  5.045000 1.080000 ;
      RECT  4.555000 2.415000  6.075000 2.420000 ;
      RECT  4.570000 2.410000  6.075000 2.415000 ;
      RECT  4.590000 2.400000  6.075000 2.410000 ;
      RECT  4.615000 2.385000  6.075000 2.400000 ;
      RECT  4.815000 1.080000  5.045000 1.455000 ;
      RECT  4.815000 1.455000  5.280000 1.775000 ;
      RECT  4.815000 1.775000  4.985000 1.820000 ;
      RECT  5.155000 1.955000  5.630000 2.215000 ;
      RECT  5.215000 0.255000  7.220000 0.425000 ;
      RECT  5.215000 0.425000  5.620000 1.070000 ;
      RECT  5.215000 1.070000  5.630000 1.285000 ;
      RECT  5.450000 1.285000  5.630000 1.545000 ;
      RECT  5.450000 1.545000  6.175000 1.875000 ;
      RECT  5.450000 1.875000  5.630000 1.955000 ;
      RECT  5.795000 0.595000  5.975000 0.995000 ;
      RECT  5.800000 0.995000  5.975000 1.200000 ;
      RECT  5.800000 1.200000  6.515000 1.370000 ;
      RECT  5.825000 2.045000  6.515000 2.215000 ;
      RECT  5.825000 2.215000  6.075000 2.385000 ;
      RECT  5.825000 2.580000  6.075000 2.725000 ;
      RECT  6.145000 0.595000  6.470000 0.860000 ;
      RECT  6.145000 0.860000  6.855000 1.030000 ;
      RECT  6.250000 2.385000  6.855000 2.725000 ;
      RECT  6.345000 1.370000  6.515000 2.045000 ;
      RECT  6.685000 1.030000  6.855000 1.985000 ;
      RECT  6.685000 1.985000  7.605000 2.165000 ;
      RECT  6.685000 2.165000  6.855000 2.385000 ;
      RECT  7.025000 0.920000  8.920000 1.090000 ;
      RECT  7.025000 1.090000  7.265000 1.805000 ;
      RECT  7.050000 0.425000  7.220000 0.580000 ;
      RECT  7.050000 0.580000  8.100000 0.750000 ;
      RECT  7.435000 1.260000  8.485000 1.545000 ;
      RECT  7.435000 1.545000  7.605000 1.985000 ;
      RECT  7.435000 2.165000  7.605000 2.320000 ;
      RECT  7.435000 2.320000  7.765000 2.745000 ;
      RECT  7.930000 0.255000  9.260000 0.425000 ;
      RECT  7.930000 0.425000  8.100000 0.580000 ;
      RECT  8.270000 0.595000  8.920000 0.920000 ;
      RECT  8.750000 1.090000  8.920000 1.715000 ;
      RECT  8.750000 1.715000  9.115000 2.755000 ;
      RECT  9.090000 0.425000  9.260000 1.005000 ;
      RECT  9.090000 1.005000 10.050000 1.335000 ;
      RECT  9.320000 1.840000  9.600000 2.520000 ;
      RECT  9.320000 2.520000 10.390000 2.850000 ;
      RECT  9.430000 0.480000 10.390000 0.810000 ;
      RECT  9.785000 1.335000 10.050000 2.330000 ;
      RECT 10.220000 0.810000 10.390000 1.030000 ;
      RECT 10.220000 1.030000 11.190000 1.110000 ;
      RECT 10.220000 1.110000 11.890000 1.200000 ;
      RECT 10.220000 1.200000 10.390000 2.520000 ;
      RECT 10.560000 1.370000 10.850000 1.580000 ;
      RECT 10.560000 1.580000 12.230000 1.750000 ;
      RECT 10.560000 1.750000 10.850000 2.390000 ;
      RECT 10.560000 2.390000 11.740000 2.560000 ;
      RECT 11.020000 1.200000 11.890000 1.410000 ;
      RECT 11.410000 2.560000 11.740000 2.980000 ;
      RECT 11.545000 0.350000 11.875000 0.770000 ;
      RECT 11.545000 0.770000 12.230000 0.940000 ;
      RECT 12.060000 0.940000 12.230000 1.580000 ;
      RECT 12.445000 1.940000 12.775000 2.980000 ;
      RECT 12.605000 0.350000 12.865000 1.300000 ;
      RECT 12.605000 1.300000 13.355000 1.630000 ;
      RECT 12.605000 1.630000 12.775000 1.940000 ;
  END
END sky130_fd_sc_ls__sdfrtp_2
