# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ls__o2111a_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ls__o2111a_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.160000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.522000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.325000 1.450000 5.655000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.522000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485000 1.450000 5.155000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.474000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.985000 1.450000 3.315000 1.780000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.474000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.450000 1.795000 1.780000 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.474000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.450000 0.550000 1.780000 ;
    END
  END D1
  PIN X
    ANTENNADIFFAREA  1.142400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.185000 0.350000 6.515000 1.010000 ;
        RECT 6.185000 1.010000 8.035000 1.180000 ;
        RECT 6.315000 1.850000 7.545000 2.180000 ;
        RECT 6.315000 2.180000 6.590000 2.980000 ;
        RECT 7.185000 0.350000 7.515000 1.010000 ;
        RECT 7.295000 1.480000 8.035000 1.650000 ;
        RECT 7.295000 1.650000 7.545000 1.850000 ;
        RECT 7.295000 2.180000 7.545000 2.980000 ;
        RECT 7.805000 1.180000 8.035000 1.480000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.160000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.160000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.160000 0.085000 ;
      RECT 0.000000  3.245000 8.160000 3.415000 ;
      RECT 0.115000  0.255000 2.250000 0.425000 ;
      RECT 0.115000  0.425000 1.230000 0.600000 ;
      RECT 0.115000  0.600000 0.380000 1.115000 ;
      RECT 0.115000  1.950000 6.145000 2.120000 ;
      RECT 0.115000  2.120000 0.445000 2.820000 ;
      RECT 0.550000  0.770000 0.890000 1.130000 ;
      RECT 0.615000  2.315000 0.945000 3.245000 ;
      RECT 0.720000  1.130000 0.890000 1.950000 ;
      RECT 1.060000  0.600000 1.230000 1.130000 ;
      RECT 1.115000  2.120000 1.445000 2.820000 ;
      RECT 1.410000  0.595000 1.740000 0.710000 ;
      RECT 1.410000  0.710000 3.125000 0.880000 ;
      RECT 1.410000  0.880000 1.740000 1.130000 ;
      RECT 1.615000  2.315000 1.945000 3.245000 ;
      RECT 1.920000  0.425000 2.250000 0.540000 ;
      RECT 2.150000  1.940000 2.480000 1.950000 ;
      RECT 2.150000  2.120000 2.480000 2.820000 ;
      RECT 2.365000  1.050000 3.555000 1.110000 ;
      RECT 2.365000  1.110000 5.505000 1.280000 ;
      RECT 2.365000  1.280000 2.775000 1.300000 ;
      RECT 2.685000  2.315000 3.015000 3.245000 ;
      RECT 2.875000  0.520000 3.125000 0.710000 ;
      RECT 3.220000  2.120000 3.550000 2.905000 ;
      RECT 3.220000  2.905000 4.550000 3.075000 ;
      RECT 3.305000  0.520000 3.555000 1.050000 ;
      RECT 3.720000  2.290000 5.610000 2.460000 ;
      RECT 3.720000  2.460000 4.050000 2.735000 ;
      RECT 3.735000  0.085000 4.065000 0.940000 ;
      RECT 4.220000  2.630000 4.550000 2.905000 ;
      RECT 4.235000  0.520000 4.565000 1.110000 ;
      RECT 4.780000  2.630000 5.110000 3.245000 ;
      RECT 4.825000  0.085000 5.155000 0.940000 ;
      RECT 5.280000  2.460000 5.610000 2.980000 ;
      RECT 5.335000  0.350000 5.505000 1.110000 ;
      RECT 5.685000  0.085000 6.015000 1.130000 ;
      RECT 5.815000  2.290000 6.145000 3.245000 ;
      RECT 5.975000  1.350000 7.125000 1.680000 ;
      RECT 5.975000  1.680000 6.145000 1.950000 ;
      RECT 6.685000  0.085000 7.015000 0.815000 ;
      RECT 6.765000  2.350000 7.095000 3.245000 ;
      RECT 7.685000  0.085000 8.015000 0.815000 ;
      RECT 7.715000  1.820000 8.045000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
  END
END sky130_fd_sc_ls__o2111a_4
END LIBRARY
