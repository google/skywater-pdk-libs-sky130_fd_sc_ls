* File: sky130_fd_sc_ls__or4bb_2.pxi.spice
* Created: Wed Sep  2 11:26:17 2020
* 
x_PM_SKY130_FD_SC_LS__OR4BB_2%D_N N_D_N_c_96_n N_D_N_c_100_n N_D_N_c_101_n
+ N_D_N_M1010_g N_D_N_c_97_n N_D_N_M1004_g D_N N_D_N_c_98_n
+ PM_SKY130_FD_SC_LS__OR4BB_2%D_N
x_PM_SKY130_FD_SC_LS__OR4BB_2%A_182_270# N_A_182_270#_M1011_d
+ N_A_182_270#_M1000_d N_A_182_270#_M1009_s N_A_182_270#_c_138_n
+ N_A_182_270#_M1008_g N_A_182_270#_M1002_g N_A_182_270#_c_128_n
+ N_A_182_270#_c_129_n N_A_182_270#_c_130_n N_A_182_270#_M1003_g
+ N_A_182_270#_c_131_n N_A_182_270#_M1013_g N_A_182_270#_c_132_n
+ N_A_182_270#_c_133_n N_A_182_270#_c_134_n N_A_182_270#_c_135_n
+ N_A_182_270#_c_180_p N_A_182_270#_c_136_n N_A_182_270#_c_143_n
+ N_A_182_270#_c_137_n N_A_182_270#_c_181_p
+ PM_SKY130_FD_SC_LS__OR4BB_2%A_182_270#
x_PM_SKY130_FD_SC_LS__OR4BB_2%A_27_424# N_A_27_424#_M1004_s N_A_27_424#_M1010_s
+ N_A_27_424#_M1011_g N_A_27_424#_c_253_n N_A_27_424#_M1009_g
+ N_A_27_424#_c_248_n N_A_27_424#_c_261_n N_A_27_424#_c_249_n
+ N_A_27_424#_c_250_n N_A_27_424#_c_255_n N_A_27_424#_c_251_n
+ N_A_27_424#_c_257_n N_A_27_424#_c_258_n N_A_27_424#_c_252_n
+ PM_SKY130_FD_SC_LS__OR4BB_2%A_27_424#
x_PM_SKY130_FD_SC_LS__OR4BB_2%A_548_110# N_A_548_110#_M1007_d
+ N_A_548_110#_M1001_d N_A_548_110#_M1014_g N_A_548_110#_c_336_n
+ N_A_548_110#_M1005_g N_A_548_110#_c_337_n N_A_548_110#_c_398_p
+ N_A_548_110#_c_338_n N_A_548_110#_c_339_n N_A_548_110#_c_340_n
+ N_A_548_110#_c_356_n N_A_548_110#_c_344_n
+ PM_SKY130_FD_SC_LS__OR4BB_2%A_548_110#
x_PM_SKY130_FD_SC_LS__OR4BB_2%B N_B_M1000_g N_B_c_412_n N_B_c_413_n N_B_c_418_n
+ N_B_M1006_g N_B_c_414_n B N_B_c_416_n PM_SKY130_FD_SC_LS__OR4BB_2%B
x_PM_SKY130_FD_SC_LS__OR4BB_2%A N_A_c_456_n N_A_M1015_g N_A_M1012_g A
+ N_A_c_458_n PM_SKY130_FD_SC_LS__OR4BB_2%A
x_PM_SKY130_FD_SC_LS__OR4BB_2%C_N N_C_N_c_490_n N_C_N_c_495_n N_C_N_M1001_g
+ N_C_N_M1007_g C_N N_C_N_c_492_n N_C_N_c_493_n PM_SKY130_FD_SC_LS__OR4BB_2%C_N
x_PM_SKY130_FD_SC_LS__OR4BB_2%VPWR N_VPWR_M1010_d N_VPWR_M1013_s N_VPWR_M1015_d
+ N_VPWR_c_523_n N_VPWR_c_524_n N_VPWR_c_525_n N_VPWR_c_526_n N_VPWR_c_527_n
+ VPWR N_VPWR_c_528_n N_VPWR_c_529_n N_VPWR_c_530_n N_VPWR_c_522_n
+ N_VPWR_c_532_n N_VPWR_c_533_n PM_SKY130_FD_SC_LS__OR4BB_2%VPWR
x_PM_SKY130_FD_SC_LS__OR4BB_2%X N_X_M1002_d N_X_M1008_d N_X_c_580_n N_X_c_582_n
+ N_X_c_576_n X X PM_SKY130_FD_SC_LS__OR4BB_2%X
x_PM_SKY130_FD_SC_LS__OR4BB_2%VGND N_VGND_M1004_d N_VGND_M1003_s N_VGND_M1014_d
+ N_VGND_M1012_d N_VGND_c_609_n N_VGND_c_610_n N_VGND_c_611_n N_VGND_c_612_n
+ N_VGND_c_613_n N_VGND_c_614_n N_VGND_c_637_n VGND N_VGND_c_615_n
+ N_VGND_c_616_n N_VGND_c_617_n N_VGND_c_618_n N_VGND_c_619_n N_VGND_c_620_n
+ N_VGND_c_621_n N_VGND_c_622_n PM_SKY130_FD_SC_LS__OR4BB_2%VGND
cc_1 VNB N_D_N_c_96_n 0.0330083f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.77
cc_2 VNB N_D_N_c_97_n 0.0247296f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.35
cc_3 VNB N_D_N_c_98_n 0.0146969f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.515
cc_4 VNB N_A_182_270#_c_128_n 0.0166342f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.665
cc_5 VNB N_A_182_270#_c_129_n 0.0151503f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_A_182_270#_c_130_n 0.0180833f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_182_270#_c_131_n 0.0236464f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_182_270#_c_132_n 0.0166056f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_182_270#_c_133_n 0.00956212f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_182_270#_c_134_n 0.0050273f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_182_270#_c_135_n 0.00374555f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_182_270#_c_136_n 0.00568326f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_182_270#_c_137_n 2.17555e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_424#_M1011_g 0.0282719f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_15 VNB N_A_27_424#_c_248_n 0.0171251f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_27_424#_c_249_n 0.00736922f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_27_424#_c_250_n 0.00754568f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_27_424#_c_251_n 0.00134284f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_27_424#_c_252_n 0.0277155f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_548_110#_M1014_g 0.0215462f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_21 VNB N_A_548_110#_c_336_n 0.0180701f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1.515
cc_22 VNB N_A_548_110#_c_337_n 0.00168047f $X=-0.19 $Y=-0.245 $X2=0.337
+ $Y2=1.665
cc_23 VNB N_A_548_110#_c_338_n 0.00291601f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_548_110#_c_339_n 0.00967002f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_548_110#_c_340_n 0.0220417f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_B_M1000_g 0.0106411f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.54
cc_27 VNB N_B_c_412_n 0.00605878f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.54
cc_28 VNB N_B_c_413_n 0.008989f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.35
cc_29 VNB N_B_c_414_n 0.0460464f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.515
cc_30 VNB B 0.00867424f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.665
cc_31 VNB N_B_c_416_n 0.00287377f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_c_456_n 0.0184029f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.77
cc_33 VNB N_A_M1012_g 0.0205097f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.35
cc_34 VNB N_A_c_458_n 0.00326462f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.515
cc_35 VNB N_C_N_c_490_n 0.00147691f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.955
cc_36 VNB N_C_N_M1007_g 0.0364307f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.965
cc_37 VNB N_C_N_c_492_n 0.056522f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.665
cc_38 VNB N_C_N_c_493_n 0.00392685f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VPWR_c_522_n 0.203486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_X_c_576_n 0.00125868f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.515
cc_41 VNB X 0.00272487f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_609_n 0.0260483f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_610_n 0.0280682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_611_n 0.0175939f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_612_n 0.012565f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_613_n 0.0229698f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_614_n 0.00326658f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_615_n 0.0208292f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_616_n 0.0203964f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_617_n 0.0238907f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_618_n 0.0178467f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_619_n 0.303661f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_620_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_621_n 0.00884799f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_622_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VPB N_D_N_c_96_n 0.0134976f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.77
cc_57 VPB N_D_N_c_100_n 0.0159532f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.955
cc_58 VPB N_D_N_c_101_n 0.0299571f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.045
cc_59 VPB N_D_N_c_98_n 0.00794482f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.515
cc_60 VPB N_A_182_270#_c_138_n 0.0152697f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_A_182_270#_c_129_n 0.00641233f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_A_182_270#_c_131_n 0.0302866f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_A_182_270#_c_135_n 0.00179111f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_A_182_270#_c_136_n 0.00320718f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_A_182_270#_c_143_n 0.00635123f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_A_27_424#_c_253_n 0.0170253f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=1.515
cc_67 VPB N_A_27_424#_c_250_n 0.00331819f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_A_27_424#_c_255_n 0.0154131f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_A_27_424#_c_251_n 0.00776083f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_A_27_424#_c_257_n 0.0235469f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_A_27_424#_c_258_n 0.020866f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_A_27_424#_c_252_n 0.0316049f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_A_548_110#_c_336_n 0.0357559f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=1.515
cc_74 VPB N_A_548_110#_c_337_n 0.00217087f $X=-0.19 $Y=1.66 $X2=0.337 $Y2=1.665
cc_75 VPB N_A_548_110#_c_338_n 0.00271194f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_A_548_110#_c_344_n 0.0402575f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_B_c_413_n 0.00692257f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=1.35
cc_78 VPB N_B_c_418_n 0.0220608f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=0.965
cc_79 VPB N_A_c_456_n 0.0350637f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.77
cc_80 VPB N_A_c_458_n 0.00285797f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.515
cc_81 VPB N_C_N_c_490_n 0.00719311f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.955
cc_82 VPB N_C_N_c_495_n 0.0289617f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.045
cc_83 VPB N_C_N_c_493_n 0.00740371f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_523_n 0.00590389f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.515
cc_85 VPB N_VPWR_c_524_n 0.00981352f $X=-0.19 $Y=1.66 $X2=0.337 $Y2=1.665
cc_86 VPB N_VPWR_c_525_n 0.0125415f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_526_n 0.0590149f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_527_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_528_n 0.0188333f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_529_n 0.017918f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_530_n 0.0209571f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_522_n 0.112881f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_532_n 0.00614589f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_533_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_95 VPB N_X_c_576_n 0.0016224f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.515
cc_96 N_D_N_c_96_n N_A_182_270#_c_138_n 0.00750183f $X=0.495 $Y=1.77 $X2=0 $Y2=0
cc_97 N_D_N_c_101_n N_A_182_270#_c_138_n 0.0258655f $X=0.495 $Y=2.045 $X2=0
+ $Y2=0
cc_98 N_D_N_c_96_n N_A_182_270#_c_129_n 0.012965f $X=0.495 $Y=1.77 $X2=0 $Y2=0
cc_99 N_D_N_c_97_n N_A_182_270#_c_132_n 0.0168398f $X=0.5 $Y=1.35 $X2=0 $Y2=0
cc_100 N_D_N_c_97_n N_A_27_424#_c_248_n 0.00665298f $X=0.5 $Y=1.35 $X2=0 $Y2=0
cc_101 N_D_N_c_97_n N_A_27_424#_c_261_n 0.0116766f $X=0.5 $Y=1.35 $X2=0 $Y2=0
cc_102 N_D_N_c_98_n N_A_27_424#_c_261_n 0.00722636f $X=0.385 $Y=1.515 $X2=0
+ $Y2=0
cc_103 N_D_N_c_96_n N_A_27_424#_c_249_n 0.00141403f $X=0.495 $Y=1.77 $X2=0 $Y2=0
cc_104 N_D_N_c_97_n N_A_27_424#_c_249_n 0.00194462f $X=0.5 $Y=1.35 $X2=0 $Y2=0
cc_105 N_D_N_c_98_n N_A_27_424#_c_249_n 0.0246812f $X=0.385 $Y=1.515 $X2=0 $Y2=0
cc_106 N_D_N_c_96_n N_A_27_424#_c_250_n 0.0065997f $X=0.495 $Y=1.77 $X2=0 $Y2=0
cc_107 N_D_N_c_101_n N_A_27_424#_c_250_n 0.00120561f $X=0.495 $Y=2.045 $X2=0
+ $Y2=0
cc_108 N_D_N_c_97_n N_A_27_424#_c_250_n 0.00617026f $X=0.5 $Y=1.35 $X2=0 $Y2=0
cc_109 N_D_N_c_98_n N_A_27_424#_c_250_n 0.0329139f $X=0.385 $Y=1.515 $X2=0 $Y2=0
cc_110 N_D_N_c_101_n N_A_27_424#_c_257_n 0.0105346f $X=0.495 $Y=2.045 $X2=0
+ $Y2=0
cc_111 N_D_N_c_96_n N_A_27_424#_c_258_n 0.00101847f $X=0.495 $Y=1.77 $X2=0 $Y2=0
cc_112 N_D_N_c_101_n N_A_27_424#_c_258_n 0.0207121f $X=0.495 $Y=2.045 $X2=0
+ $Y2=0
cc_113 N_D_N_c_98_n N_A_27_424#_c_258_n 0.0221141f $X=0.385 $Y=1.515 $X2=0 $Y2=0
cc_114 N_D_N_c_101_n N_VPWR_c_523_n 0.00519769f $X=0.495 $Y=2.045 $X2=0 $Y2=0
cc_115 N_D_N_c_101_n N_VPWR_c_528_n 0.00445602f $X=0.495 $Y=2.045 $X2=0 $Y2=0
cc_116 N_D_N_c_101_n N_VPWR_c_522_n 0.00860933f $X=0.495 $Y=2.045 $X2=0 $Y2=0
cc_117 N_D_N_c_97_n X 7.18431e-19 $X=0.5 $Y=1.35 $X2=0 $Y2=0
cc_118 N_D_N_c_97_n N_VGND_c_609_n 0.00390595f $X=0.5 $Y=1.35 $X2=0 $Y2=0
cc_119 N_D_N_c_97_n N_VGND_c_615_n 0.0036924f $X=0.5 $Y=1.35 $X2=0 $Y2=0
cc_120 N_D_N_c_97_n N_VGND_c_619_n 0.00451834f $X=0.5 $Y=1.35 $X2=0 $Y2=0
cc_121 N_A_182_270#_c_130_n N_A_27_424#_M1011_g 0.0133144f $X=1.445 $Y=1.35
+ $X2=0 $Y2=0
cc_122 N_A_182_270#_c_131_n N_A_27_424#_M1011_g 0.00343657f $X=1.45 $Y=1.765
+ $X2=0 $Y2=0
cc_123 N_A_182_270#_c_133_n N_A_27_424#_M1011_g 0.0168494f $X=2.31 $Y=1.215
+ $X2=0 $Y2=0
cc_124 N_A_182_270#_c_134_n N_A_27_424#_M1011_g 0.00377486f $X=2.475 $Y=0.745
+ $X2=0 $Y2=0
cc_125 N_A_182_270#_c_135_n N_A_27_424#_M1011_g 0.0026842f $X=2.52 $Y=2.61 $X2=0
+ $Y2=0
cc_126 N_A_182_270#_c_136_n N_A_27_424#_M1011_g 0.00161653f $X=1.565 $Y=1.215
+ $X2=0 $Y2=0
cc_127 N_A_182_270#_c_135_n N_A_27_424#_c_253_n 0.0177427f $X=2.52 $Y=2.61 $X2=0
+ $Y2=0
cc_128 N_A_182_270#_c_143_n N_A_27_424#_c_253_n 0.0129527f $X=2.215 $Y=2.795
+ $X2=0 $Y2=0
cc_129 N_A_182_270#_c_132_n N_A_27_424#_c_248_n 5.28751e-19 $X=1 $Y=1.35 $X2=0
+ $Y2=0
cc_130 N_A_182_270#_c_138_n N_A_27_424#_c_250_n 0.00195921f $X=1 $Y=1.765 $X2=0
+ $Y2=0
cc_131 N_A_182_270#_c_129_n N_A_27_424#_c_250_n 0.00400056f $X=1.09 $Y=1.467
+ $X2=0 $Y2=0
cc_132 N_A_182_270#_c_132_n N_A_27_424#_c_250_n 0.00120976f $X=1 $Y=1.35 $X2=0
+ $Y2=0
cc_133 N_A_182_270#_M1009_s N_A_27_424#_c_255_n 0.00510534f $X=2.08 $Y=1.96
+ $X2=0 $Y2=0
cc_134 N_A_182_270#_c_138_n N_A_27_424#_c_255_n 0.0192233f $X=1 $Y=1.765 $X2=0
+ $Y2=0
cc_135 N_A_182_270#_c_128_n N_A_27_424#_c_255_n 4.0436e-19 $X=1.36 $Y=1.467
+ $X2=0 $Y2=0
cc_136 N_A_182_270#_c_131_n N_A_27_424#_c_255_n 0.0194491f $X=1.45 $Y=1.765
+ $X2=0 $Y2=0
cc_137 N_A_182_270#_c_135_n N_A_27_424#_c_255_n 0.0134181f $X=2.52 $Y=2.61 $X2=0
+ $Y2=0
cc_138 N_A_182_270#_c_136_n N_A_27_424#_c_255_n 0.00827027f $X=1.565 $Y=1.215
+ $X2=0 $Y2=0
cc_139 N_A_182_270#_c_143_n N_A_27_424#_c_255_n 0.0186031f $X=2.215 $Y=2.795
+ $X2=0 $Y2=0
cc_140 N_A_182_270#_M1009_s N_A_27_424#_c_251_n 0.00539353f $X=2.08 $Y=1.96
+ $X2=0 $Y2=0
cc_141 N_A_182_270#_c_131_n N_A_27_424#_c_251_n 0.0112335f $X=1.45 $Y=1.765
+ $X2=0 $Y2=0
cc_142 N_A_182_270#_c_133_n N_A_27_424#_c_251_n 0.0228543f $X=2.31 $Y=1.215
+ $X2=0 $Y2=0
cc_143 N_A_182_270#_c_135_n N_A_27_424#_c_251_n 0.0579813f $X=2.52 $Y=2.61 $X2=0
+ $Y2=0
cc_144 N_A_182_270#_c_136_n N_A_27_424#_c_251_n 0.0119071f $X=1.565 $Y=1.215
+ $X2=0 $Y2=0
cc_145 N_A_182_270#_c_138_n N_A_27_424#_c_257_n 8.57658e-19 $X=1 $Y=1.765 $X2=0
+ $Y2=0
cc_146 N_A_182_270#_c_131_n N_A_27_424#_c_252_n 0.0155414f $X=1.45 $Y=1.765
+ $X2=0 $Y2=0
cc_147 N_A_182_270#_c_133_n N_A_27_424#_c_252_n 0.00271878f $X=2.31 $Y=1.215
+ $X2=0 $Y2=0
cc_148 N_A_182_270#_c_135_n N_A_27_424#_c_252_n 0.0131024f $X=2.52 $Y=2.61 $X2=0
+ $Y2=0
cc_149 N_A_182_270#_c_136_n N_A_27_424#_c_252_n 8.56237e-19 $X=1.565 $Y=1.215
+ $X2=0 $Y2=0
cc_150 N_A_182_270#_c_137_n N_A_27_424#_c_252_n 0.00584755f $X=2.475 $Y=1.215
+ $X2=0 $Y2=0
cc_151 N_A_182_270#_c_134_n N_A_548_110#_M1014_g 0.00820624f $X=2.475 $Y=0.745
+ $X2=0 $Y2=0
cc_152 N_A_182_270#_c_135_n N_A_548_110#_M1014_g 0.00622541f $X=2.52 $Y=2.61
+ $X2=0 $Y2=0
cc_153 N_A_182_270#_c_180_p N_A_548_110#_M1014_g 0.0149081f $X=3.405 $Y=1.215
+ $X2=0 $Y2=0
cc_154 N_A_182_270#_c_181_p N_A_548_110#_M1014_g 6.67717e-19 $X=3.57 $Y=1.07
+ $X2=0 $Y2=0
cc_155 N_A_182_270#_c_135_n N_A_548_110#_c_336_n 0.0110943f $X=2.52 $Y=2.61
+ $X2=0 $Y2=0
cc_156 N_A_182_270#_c_180_p N_A_548_110#_c_336_n 0.00113283f $X=3.405 $Y=1.215
+ $X2=0 $Y2=0
cc_157 N_A_182_270#_c_143_n N_A_548_110#_c_336_n 0.00533687f $X=2.215 $Y=2.795
+ $X2=0 $Y2=0
cc_158 N_A_182_270#_c_135_n N_A_548_110#_c_337_n 0.037138f $X=2.52 $Y=2.61 $X2=0
+ $Y2=0
cc_159 N_A_182_270#_c_180_p N_A_548_110#_c_337_n 0.0206464f $X=3.405 $Y=1.215
+ $X2=0 $Y2=0
cc_160 N_A_182_270#_c_181_p N_A_548_110#_c_338_n 0.0070468f $X=3.57 $Y=1.07
+ $X2=0 $Y2=0
cc_161 N_A_182_270#_c_181_p N_A_548_110#_c_339_n 0.00769979f $X=3.57 $Y=1.07
+ $X2=0 $Y2=0
cc_162 N_A_182_270#_c_180_p N_A_548_110#_c_356_n 0.00666702f $X=3.405 $Y=1.215
+ $X2=0 $Y2=0
cc_163 N_A_182_270#_c_181_p N_A_548_110#_c_356_n 7.22293e-19 $X=3.57 $Y=1.07
+ $X2=0 $Y2=0
cc_164 N_A_182_270#_c_180_p N_B_M1000_g 0.0118685f $X=3.405 $Y=1.215 $X2=0 $Y2=0
cc_165 N_A_182_270#_c_181_p N_B_M1000_g 0.00764803f $X=3.57 $Y=1.07 $X2=0 $Y2=0
cc_166 N_A_182_270#_c_180_p N_B_c_414_n 0.00128204f $X=3.405 $Y=1.215 $X2=0
+ $Y2=0
cc_167 N_A_182_270#_c_181_p B 0.0170437f $X=3.57 $Y=1.07 $X2=0 $Y2=0
cc_168 N_A_182_270#_c_180_p N_B_c_416_n 0.00494392f $X=3.405 $Y=1.215 $X2=0
+ $Y2=0
cc_169 N_A_182_270#_c_181_p N_B_c_416_n 0.00258991f $X=3.57 $Y=1.07 $X2=0 $Y2=0
cc_170 N_A_182_270#_c_181_p N_A_M1012_g 0.00833003f $X=3.57 $Y=1.07 $X2=0 $Y2=0
cc_171 N_A_182_270#_c_181_p N_A_c_458_n 0.0181575f $X=3.57 $Y=1.07 $X2=0 $Y2=0
cc_172 N_A_182_270#_c_181_p N_C_N_M1007_g 8.62984e-19 $X=3.57 $Y=1.07 $X2=0
+ $Y2=0
cc_173 N_A_182_270#_c_138_n N_VPWR_c_523_n 0.0101642f $X=1 $Y=1.765 $X2=0 $Y2=0
cc_174 N_A_182_270#_c_131_n N_VPWR_c_523_n 0.00140807f $X=1.45 $Y=1.765 $X2=0
+ $Y2=0
cc_175 N_A_182_270#_c_138_n N_VPWR_c_524_n 0.00142182f $X=1 $Y=1.765 $X2=0 $Y2=0
cc_176 N_A_182_270#_c_131_n N_VPWR_c_524_n 0.0115353f $X=1.45 $Y=1.765 $X2=0
+ $Y2=0
cc_177 N_A_182_270#_c_143_n N_VPWR_c_524_n 0.027168f $X=2.215 $Y=2.795 $X2=0
+ $Y2=0
cc_178 N_A_182_270#_c_143_n N_VPWR_c_526_n 0.0183917f $X=2.215 $Y=2.795 $X2=0
+ $Y2=0
cc_179 N_A_182_270#_c_138_n N_VPWR_c_529_n 0.00429299f $X=1 $Y=1.765 $X2=0 $Y2=0
cc_180 N_A_182_270#_c_131_n N_VPWR_c_529_n 0.00413917f $X=1.45 $Y=1.765 $X2=0
+ $Y2=0
cc_181 N_A_182_270#_c_138_n N_VPWR_c_522_n 0.00847721f $X=1 $Y=1.765 $X2=0 $Y2=0
cc_182 N_A_182_270#_c_131_n N_VPWR_c_522_n 0.00817726f $X=1.45 $Y=1.765 $X2=0
+ $Y2=0
cc_183 N_A_182_270#_c_143_n N_VPWR_c_522_n 0.0183559f $X=2.215 $Y=2.795 $X2=0
+ $Y2=0
cc_184 N_A_182_270#_c_128_n N_X_c_580_n 0.0014328f $X=1.36 $Y=1.467 $X2=0 $Y2=0
cc_185 N_A_182_270#_c_132_n N_X_c_580_n 0.00133297f $X=1 $Y=1.35 $X2=0 $Y2=0
cc_186 N_A_182_270#_c_138_n N_X_c_582_n 0.00256871f $X=1 $Y=1.765 $X2=0 $Y2=0
cc_187 N_A_182_270#_c_128_n N_X_c_582_n 0.00319311f $X=1.36 $Y=1.467 $X2=0 $Y2=0
cc_188 N_A_182_270#_c_131_n N_X_c_582_n 0.00574199f $X=1.45 $Y=1.765 $X2=0 $Y2=0
cc_189 N_A_182_270#_c_138_n N_X_c_576_n 0.00137915f $X=1 $Y=1.765 $X2=0 $Y2=0
cc_190 N_A_182_270#_c_128_n N_X_c_576_n 0.0105814f $X=1.36 $Y=1.467 $X2=0 $Y2=0
cc_191 N_A_182_270#_c_129_n N_X_c_576_n 0.00627796f $X=1.09 $Y=1.467 $X2=0 $Y2=0
cc_192 N_A_182_270#_c_130_n N_X_c_576_n 0.00120456f $X=1.445 $Y=1.35 $X2=0 $Y2=0
cc_193 N_A_182_270#_c_131_n N_X_c_576_n 0.00425475f $X=1.45 $Y=1.765 $X2=0 $Y2=0
cc_194 N_A_182_270#_c_132_n N_X_c_576_n 0.00278431f $X=1 $Y=1.35 $X2=0 $Y2=0
cc_195 N_A_182_270#_c_136_n N_X_c_576_n 0.0308971f $X=1.565 $Y=1.215 $X2=0 $Y2=0
cc_196 N_A_182_270#_c_130_n X 5.16304e-19 $X=1.445 $Y=1.35 $X2=0 $Y2=0
cc_197 N_A_182_270#_c_132_n X 0.00898935f $X=1 $Y=1.35 $X2=0 $Y2=0
cc_198 N_A_182_270#_c_135_n A_503_392# 0.00707252f $X=2.52 $Y=2.61 $X2=-0.19
+ $Y2=-0.245
cc_199 N_A_182_270#_c_143_n A_503_392# 0.0028132f $X=2.215 $Y=2.795 $X2=-0.19
+ $Y2=-0.245
cc_200 N_A_182_270#_c_133_n N_VGND_M1003_s 0.00461621f $X=2.31 $Y=1.215 $X2=0
+ $Y2=0
cc_201 N_A_182_270#_c_136_n N_VGND_M1003_s 0.00222344f $X=1.565 $Y=1.215 $X2=0
+ $Y2=0
cc_202 N_A_182_270#_c_180_p N_VGND_M1014_d 0.00756824f $X=3.405 $Y=1.215 $X2=0
+ $Y2=0
cc_203 N_A_182_270#_c_132_n N_VGND_c_609_n 0.00523841f $X=1 $Y=1.35 $X2=0 $Y2=0
cc_204 N_A_182_270#_c_130_n N_VGND_c_610_n 0.00735637f $X=1.445 $Y=1.35 $X2=0
+ $Y2=0
cc_205 N_A_182_270#_c_131_n N_VGND_c_610_n 7.4832e-19 $X=1.45 $Y=1.765 $X2=0
+ $Y2=0
cc_206 N_A_182_270#_c_133_n N_VGND_c_610_n 0.0203901f $X=2.31 $Y=1.215 $X2=0
+ $Y2=0
cc_207 N_A_182_270#_c_134_n N_VGND_c_610_n 0.0103558f $X=2.475 $Y=0.745 $X2=0
+ $Y2=0
cc_208 N_A_182_270#_c_136_n N_VGND_c_610_n 0.011201f $X=1.565 $Y=1.215 $X2=0
+ $Y2=0
cc_209 N_A_182_270#_c_134_n N_VGND_c_611_n 0.0119895f $X=2.475 $Y=0.745 $X2=0
+ $Y2=0
cc_210 N_A_182_270#_c_134_n N_VGND_c_613_n 0.00749442f $X=2.475 $Y=0.745 $X2=0
+ $Y2=0
cc_211 N_A_182_270#_c_134_n N_VGND_c_637_n 0.0172025f $X=2.475 $Y=0.745 $X2=0
+ $Y2=0
cc_212 N_A_182_270#_c_180_p N_VGND_c_637_n 0.0238294f $X=3.405 $Y=1.215 $X2=0
+ $Y2=0
cc_213 N_A_182_270#_c_181_p N_VGND_c_637_n 0.00797901f $X=3.57 $Y=1.07 $X2=0
+ $Y2=0
cc_214 N_A_182_270#_c_130_n N_VGND_c_616_n 0.00487664f $X=1.445 $Y=1.35 $X2=0
+ $Y2=0
cc_215 N_A_182_270#_c_132_n N_VGND_c_616_n 0.00462542f $X=1 $Y=1.35 $X2=0 $Y2=0
cc_216 N_A_182_270#_c_130_n N_VGND_c_619_n 0.00505379f $X=1.445 $Y=1.35 $X2=0
+ $Y2=0
cc_217 N_A_182_270#_c_132_n N_VGND_c_619_n 0.00505379f $X=1 $Y=1.35 $X2=0 $Y2=0
cc_218 N_A_182_270#_c_134_n N_VGND_c_619_n 0.0103757f $X=2.475 $Y=0.745 $X2=0
+ $Y2=0
cc_219 N_A_182_270#_c_181_p N_VGND_c_619_n 0.00125724f $X=3.57 $Y=1.07 $X2=0
+ $Y2=0
cc_220 N_A_27_424#_M1011_g N_A_548_110#_M1014_g 0.0156102f $X=2.18 $Y=0.92 $X2=0
+ $Y2=0
cc_221 N_A_27_424#_c_253_n N_A_548_110#_c_336_n 0.0545306f $X=2.44 $Y=1.885
+ $X2=0 $Y2=0
cc_222 N_A_27_424#_c_252_n N_A_548_110#_c_336_n 0.0248603f $X=2.18 $Y=1.677
+ $X2=0 $Y2=0
cc_223 N_A_27_424#_c_253_n N_A_548_110#_c_337_n 2.11464e-19 $X=2.44 $Y=1.885
+ $X2=0 $Y2=0
cc_224 N_A_27_424#_c_252_n N_A_548_110#_c_337_n 4.26403e-19 $X=2.18 $Y=1.677
+ $X2=0 $Y2=0
cc_225 N_A_27_424#_c_250_n N_VPWR_M1010_d 0.00512532f $X=0.805 $Y=2.1 $X2=-0.19
+ $Y2=-0.245
cc_226 N_A_27_424#_c_258_n N_VPWR_M1010_d 0.00558252f $X=0.89 $Y=2.27 $X2=-0.19
+ $Y2=-0.245
cc_227 N_A_27_424#_c_255_n N_VPWR_M1013_s 0.00896348f $X=1.97 $Y=2.355 $X2=0
+ $Y2=0
cc_228 N_A_27_424#_c_257_n N_VPWR_c_523_n 0.0146738f $X=0.27 $Y=2.265 $X2=0
+ $Y2=0
cc_229 N_A_27_424#_c_258_n N_VPWR_c_523_n 0.0212113f $X=0.89 $Y=2.27 $X2=0 $Y2=0
cc_230 N_A_27_424#_c_253_n N_VPWR_c_524_n 0.00340466f $X=2.44 $Y=1.885 $X2=0
+ $Y2=0
cc_231 N_A_27_424#_c_255_n N_VPWR_c_524_n 0.0220234f $X=1.97 $Y=2.355 $X2=0
+ $Y2=0
cc_232 N_A_27_424#_c_253_n N_VPWR_c_526_n 0.00314081f $X=2.44 $Y=1.885 $X2=0
+ $Y2=0
cc_233 N_A_27_424#_c_257_n N_VPWR_c_528_n 0.0143526f $X=0.27 $Y=2.265 $X2=0
+ $Y2=0
cc_234 N_A_27_424#_c_253_n N_VPWR_c_522_n 0.0039522f $X=2.44 $Y=1.885 $X2=0
+ $Y2=0
cc_235 N_A_27_424#_c_257_n N_VPWR_c_522_n 0.0119532f $X=0.27 $Y=2.265 $X2=0
+ $Y2=0
cc_236 N_A_27_424#_c_255_n N_X_M1008_d 0.00894051f $X=1.97 $Y=2.355 $X2=0 $Y2=0
cc_237 N_A_27_424#_c_255_n N_X_c_582_n 0.0165593f $X=1.97 $Y=2.355 $X2=0 $Y2=0
cc_238 N_A_27_424#_c_251_n N_X_c_582_n 0.00776338f $X=2.135 $Y=1.635 $X2=0 $Y2=0
cc_239 N_A_27_424#_c_250_n N_X_c_576_n 0.05445f $X=0.805 $Y=2.1 $X2=0 $Y2=0
cc_240 N_A_27_424#_c_248_n X 0.00432689f $X=0.285 $Y=0.925 $X2=0 $Y2=0
cc_241 N_A_27_424#_c_261_n N_VGND_M1004_d 0.0071895f $X=0.72 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_242 N_A_27_424#_c_250_n N_VGND_M1004_d 0.00108513f $X=0.805 $Y=2.1 $X2=-0.19
+ $Y2=-0.245
cc_243 N_A_27_424#_c_248_n N_VGND_c_609_n 0.006821f $X=0.285 $Y=0.925 $X2=0
+ $Y2=0
cc_244 N_A_27_424#_c_261_n N_VGND_c_609_n 0.0214588f $X=0.72 $Y=1.095 $X2=0
+ $Y2=0
cc_245 N_A_27_424#_M1011_g N_VGND_c_610_n 0.00770585f $X=2.18 $Y=0.92 $X2=0
+ $Y2=0
cc_246 N_A_27_424#_M1011_g N_VGND_c_611_n 0.00201029f $X=2.18 $Y=0.92 $X2=0
+ $Y2=0
cc_247 N_A_27_424#_M1011_g N_VGND_c_613_n 0.00428744f $X=2.18 $Y=0.92 $X2=0
+ $Y2=0
cc_248 N_A_27_424#_c_248_n N_VGND_c_615_n 0.00599771f $X=0.285 $Y=0.925 $X2=0
+ $Y2=0
cc_249 N_A_27_424#_M1011_g N_VGND_c_619_n 0.00476395f $X=2.18 $Y=0.92 $X2=0
+ $Y2=0
cc_250 N_A_27_424#_c_248_n N_VGND_c_619_n 0.0095399f $X=0.285 $Y=0.925 $X2=0
+ $Y2=0
cc_251 N_A_548_110#_M1014_g N_B_M1000_g 0.0202228f $X=2.815 $Y=1 $X2=0 $Y2=0
cc_252 N_A_548_110#_c_336_n N_B_c_412_n 0.0199464f $X=2.86 $Y=1.885 $X2=0 $Y2=0
cc_253 N_A_548_110#_c_337_n N_B_c_412_n 0.00120288f $X=2.905 $Y=1.635 $X2=0
+ $Y2=0
cc_254 N_A_548_110#_c_336_n N_B_c_418_n 0.0468166f $X=2.86 $Y=1.885 $X2=0 $Y2=0
cc_255 N_A_548_110#_c_337_n N_B_c_418_n 0.0037935f $X=2.905 $Y=1.635 $X2=0 $Y2=0
cc_256 N_A_548_110#_c_356_n N_B_c_418_n 0.0173721f $X=4.095 $Y=2.045 $X2=0 $Y2=0
cc_257 N_A_548_110#_M1014_g N_B_c_414_n 9.97833e-19 $X=2.815 $Y=1 $X2=0 $Y2=0
cc_258 N_A_548_110#_c_338_n N_A_c_456_n 0.00499815f $X=4.18 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_259 N_A_548_110#_c_356_n N_A_c_456_n 0.0193549f $X=4.095 $Y=2.045 $X2=-0.19
+ $Y2=-0.245
cc_260 N_A_548_110#_c_344_n N_A_c_456_n 0.00111902f $X=4.525 $Y=2.115 $X2=-0.19
+ $Y2=-0.245
cc_261 N_A_548_110#_c_338_n N_A_M1012_g 0.00467745f $X=4.18 $Y=1.95 $X2=0 $Y2=0
cc_262 N_A_548_110#_c_339_n N_A_M1012_g 0.00149697f $X=4.56 $Y=0.96 $X2=0 $Y2=0
cc_263 N_A_548_110#_c_337_n N_A_c_458_n 0.0135637f $X=2.905 $Y=1.635 $X2=0 $Y2=0
cc_264 N_A_548_110#_c_338_n N_A_c_458_n 0.0253244f $X=4.18 $Y=1.95 $X2=0 $Y2=0
cc_265 N_A_548_110#_c_356_n N_A_c_458_n 0.0281285f $X=4.095 $Y=2.045 $X2=0 $Y2=0
cc_266 N_A_548_110#_c_338_n N_C_N_c_490_n 0.00339822f $X=4.18 $Y=1.95 $X2=0
+ $Y2=0
cc_267 N_A_548_110#_c_338_n N_C_N_c_495_n 0.00818867f $X=4.18 $Y=1.95 $X2=0
+ $Y2=0
cc_268 N_A_548_110#_c_344_n N_C_N_c_495_n 0.0298828f $X=4.525 $Y=2.115 $X2=0
+ $Y2=0
cc_269 N_A_548_110#_c_338_n N_C_N_M1007_g 0.008544f $X=4.18 $Y=1.95 $X2=0 $Y2=0
cc_270 N_A_548_110#_c_339_n N_C_N_M1007_g 0.0181834f $X=4.56 $Y=0.96 $X2=0 $Y2=0
cc_271 N_A_548_110#_c_340_n N_C_N_M1007_g 0.00264672f $X=4.52 $Y=0.73 $X2=0
+ $Y2=0
cc_272 N_A_548_110#_c_338_n N_C_N_c_492_n 0.00863054f $X=4.18 $Y=1.95 $X2=0
+ $Y2=0
cc_273 N_A_548_110#_c_339_n N_C_N_c_492_n 0.00398336f $X=4.56 $Y=0.96 $X2=0
+ $Y2=0
cc_274 N_A_548_110#_c_344_n N_C_N_c_492_n 0.00273979f $X=4.525 $Y=2.115 $X2=0
+ $Y2=0
cc_275 N_A_548_110#_c_338_n N_C_N_c_493_n 0.0341912f $X=4.18 $Y=1.95 $X2=0 $Y2=0
cc_276 N_A_548_110#_c_339_n N_C_N_c_493_n 0.0193576f $X=4.56 $Y=0.96 $X2=0 $Y2=0
cc_277 N_A_548_110#_c_344_n N_C_N_c_493_n 0.0210109f $X=4.525 $Y=2.115 $X2=0
+ $Y2=0
cc_278 N_A_548_110#_c_356_n N_VPWR_M1015_d 0.00707426f $X=4.095 $Y=2.045 $X2=0
+ $Y2=0
cc_279 N_A_548_110#_c_344_n N_VPWR_M1015_d 0.00145521f $X=4.525 $Y=2.115 $X2=0
+ $Y2=0
cc_280 N_A_548_110#_c_356_n N_VPWR_c_525_n 0.0219301f $X=4.095 $Y=2.045 $X2=0
+ $Y2=0
cc_281 N_A_548_110#_c_344_n N_VPWR_c_525_n 0.0336818f $X=4.525 $Y=2.115 $X2=0
+ $Y2=0
cc_282 N_A_548_110#_c_336_n N_VPWR_c_526_n 0.00461464f $X=2.86 $Y=1.885 $X2=0
+ $Y2=0
cc_283 N_A_548_110#_c_344_n N_VPWR_c_530_n 0.00880551f $X=4.525 $Y=2.115 $X2=0
+ $Y2=0
cc_284 N_A_548_110#_c_336_n N_VPWR_c_522_n 0.00910115f $X=2.86 $Y=1.885 $X2=0
+ $Y2=0
cc_285 N_A_548_110#_c_344_n N_VPWR_c_522_n 0.0108814f $X=4.525 $Y=2.115 $X2=0
+ $Y2=0
cc_286 N_A_548_110#_c_398_p A_587_392# 0.00346735f $X=3.07 $Y=2.055 $X2=-0.19
+ $Y2=-0.245
cc_287 N_A_548_110#_c_356_n A_587_392# 0.00989643f $X=4.095 $Y=2.045 $X2=-0.19
+ $Y2=-0.245
cc_288 N_A_548_110#_c_356_n A_689_392# 0.00615027f $X=4.095 $Y=2.045 $X2=-0.19
+ $Y2=-0.245
cc_289 N_A_548_110#_c_338_n N_VGND_M1012_d 0.00229478f $X=4.18 $Y=1.95 $X2=0
+ $Y2=0
cc_290 N_A_548_110#_c_339_n N_VGND_M1012_d 0.00293742f $X=4.56 $Y=0.96 $X2=0
+ $Y2=0
cc_291 N_A_548_110#_M1014_g N_VGND_c_611_n 0.00606464f $X=2.815 $Y=1 $X2=0 $Y2=0
cc_292 N_A_548_110#_c_339_n N_VGND_c_612_n 0.00813205f $X=4.56 $Y=0.96 $X2=0
+ $Y2=0
cc_293 N_A_548_110#_c_340_n N_VGND_c_612_n 0.0134516f $X=4.52 $Y=0.73 $X2=0
+ $Y2=0
cc_294 N_A_548_110#_M1014_g N_VGND_c_613_n 0.00180013f $X=2.815 $Y=1 $X2=0 $Y2=0
cc_295 N_A_548_110#_M1014_g N_VGND_c_637_n 0.0043994f $X=2.815 $Y=1 $X2=0 $Y2=0
cc_296 N_A_548_110#_c_340_n N_VGND_c_618_n 0.00808175f $X=4.52 $Y=0.73 $X2=0
+ $Y2=0
cc_297 N_A_548_110#_M1014_g N_VGND_c_619_n 0.00215127f $X=2.815 $Y=1 $X2=0 $Y2=0
cc_298 N_A_548_110#_c_340_n N_VGND_c_619_n 0.00859001f $X=4.52 $Y=0.73 $X2=0
+ $Y2=0
cc_299 N_B_c_412_n N_A_c_456_n 0.0248418f $X=3.37 $Y=1.485 $X2=-0.19 $Y2=-0.245
cc_300 N_B_c_418_n N_A_c_456_n 0.0654639f $X=3.37 $Y=1.885 $X2=-0.19 $Y2=-0.245
cc_301 N_B_M1000_g N_A_M1012_g 0.0180889f $X=3.355 $Y=1 $X2=0 $Y2=0
cc_302 N_B_c_412_n N_A_M1012_g 0.00387691f $X=3.37 $Y=1.485 $X2=0 $Y2=0
cc_303 N_B_c_414_n N_A_M1012_g 9.87758e-19 $X=3.315 $Y=0.405 $X2=0 $Y2=0
cc_304 B N_A_M1012_g 0.00105619f $X=3.515 $Y=0.47 $X2=0 $Y2=0
cc_305 N_B_c_412_n N_A_c_458_n 0.00381682f $X=3.37 $Y=1.485 $X2=0 $Y2=0
cc_306 B N_C_N_M1007_g 7.14048e-19 $X=3.515 $Y=0.47 $X2=0 $Y2=0
cc_307 N_B_c_418_n N_VPWR_c_525_n 0.00380728f $X=3.37 $Y=1.885 $X2=0 $Y2=0
cc_308 N_B_c_418_n N_VPWR_c_526_n 0.00461464f $X=3.37 $Y=1.885 $X2=0 $Y2=0
cc_309 N_B_c_418_n N_VPWR_c_522_n 0.00909821f $X=3.37 $Y=1.885 $X2=0 $Y2=0
cc_310 N_B_M1000_g N_VGND_c_611_n 0.00210807f $X=3.355 $Y=1 $X2=0 $Y2=0
cc_311 N_B_c_414_n N_VGND_c_611_n 0.00268668f $X=3.315 $Y=0.405 $X2=0 $Y2=0
cc_312 B N_VGND_c_611_n 0.0035728f $X=3.515 $Y=0.47 $X2=0 $Y2=0
cc_313 N_B_c_416_n N_VGND_c_611_n 0.0246471f $X=3.485 $Y=0.462 $X2=0 $Y2=0
cc_314 N_B_c_414_n N_VGND_c_612_n 0.00171528f $X=3.315 $Y=0.405 $X2=0 $Y2=0
cc_315 B N_VGND_c_612_n 0.030525f $X=3.515 $Y=0.47 $X2=0 $Y2=0
cc_316 N_B_M1000_g N_VGND_c_637_n 0.00388229f $X=3.355 $Y=1 $X2=0 $Y2=0
cc_317 N_B_c_414_n N_VGND_c_637_n 0.00101497f $X=3.315 $Y=0.405 $X2=0 $Y2=0
cc_318 N_B_c_416_n N_VGND_c_637_n 0.00325267f $X=3.485 $Y=0.462 $X2=0 $Y2=0
cc_319 N_B_c_414_n N_VGND_c_617_n 0.00584621f $X=3.315 $Y=0.405 $X2=0 $Y2=0
cc_320 N_B_c_416_n N_VGND_c_617_n 0.0372487f $X=3.485 $Y=0.462 $X2=0 $Y2=0
cc_321 N_B_c_414_n N_VGND_c_619_n 0.00760356f $X=3.315 $Y=0.405 $X2=0 $Y2=0
cc_322 N_B_c_416_n N_VGND_c_619_n 0.0200827f $X=3.485 $Y=0.462 $X2=0 $Y2=0
cc_323 N_A_c_456_n N_C_N_c_495_n 0.0204175f $X=3.76 $Y=1.885 $X2=0 $Y2=0
cc_324 N_A_M1012_g N_C_N_M1007_g 0.0179449f $X=3.795 $Y=1 $X2=0 $Y2=0
cc_325 N_A_c_456_n N_C_N_c_492_n 0.0203581f $X=3.76 $Y=1.885 $X2=0 $Y2=0
cc_326 N_A_M1012_g N_C_N_c_492_n 0.00537499f $X=3.795 $Y=1 $X2=0 $Y2=0
cc_327 N_A_c_458_n N_C_N_c_492_n 2.8993e-19 $X=3.835 $Y=1.635 $X2=0 $Y2=0
cc_328 N_A_c_456_n N_VPWR_c_525_n 0.0164805f $X=3.76 $Y=1.885 $X2=0 $Y2=0
cc_329 N_A_c_456_n N_VPWR_c_526_n 0.00413917f $X=3.76 $Y=1.885 $X2=0 $Y2=0
cc_330 N_A_c_456_n N_VPWR_c_522_n 0.00817239f $X=3.76 $Y=1.885 $X2=0 $Y2=0
cc_331 N_A_c_456_n N_VGND_c_612_n 0.00193096f $X=3.76 $Y=1.885 $X2=0 $Y2=0
cc_332 N_A_M1012_g N_VGND_c_612_n 0.00194916f $X=3.795 $Y=1 $X2=0 $Y2=0
cc_333 N_A_M1012_g N_VGND_c_617_n 0.0038748f $X=3.795 $Y=1 $X2=0 $Y2=0
cc_334 N_A_M1012_g N_VGND_c_619_n 0.00454494f $X=3.795 $Y=1 $X2=0 $Y2=0
cc_335 N_C_N_c_495_n N_VPWR_c_525_n 0.00771509f $X=4.3 $Y=1.885 $X2=0 $Y2=0
cc_336 N_C_N_c_495_n N_VPWR_c_530_n 0.00458031f $X=4.3 $Y=1.885 $X2=0 $Y2=0
cc_337 N_C_N_c_495_n N_VPWR_c_522_n 0.0049649f $X=4.3 $Y=1.885 $X2=0 $Y2=0
cc_338 N_C_N_M1007_g N_VGND_c_612_n 0.0121094f $X=4.305 $Y=0.73 $X2=0 $Y2=0
cc_339 N_C_N_M1007_g N_VGND_c_618_n 0.00429764f $X=4.305 $Y=0.73 $X2=0 $Y2=0
cc_340 N_C_N_M1007_g N_VGND_c_619_n 0.00435987f $X=4.305 $Y=0.73 $X2=0 $Y2=0
cc_341 X N_VGND_c_609_n 0.0286165f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_342 X N_VGND_c_610_n 0.00367254f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_343 X N_VGND_c_616_n 0.00819614f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_344 X N_VGND_c_619_n 0.00879294f $X=1.115 $Y=0.47 $X2=0 $Y2=0
