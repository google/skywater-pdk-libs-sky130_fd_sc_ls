* File: sky130_fd_sc_ls__o211a_4.spice
* Created: Fri Aug 28 13:43:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__o211a_4.pex.spice"
.subckt sky130_fd_sc_ls__o211a_4  VNB VPB C1 B1 A2 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A2	A2
* B1	B1
* C1	C1
* VPB	VPB
* VNB	VNB
MM1007 N_X_M1007_d N_A_91_48#_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1015 N_X_M1007_d N_A_91_48#_M1015_g N_VGND_M1015_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1016 N_X_M1016_d N_A_91_48#_M1016_g N_VGND_M1015_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.1
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1023 N_X_M1016_d N_A_91_48#_M1023_g N_VGND_M1023_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1011 N_A_510_125#_M1011_d N_B1_M1011_g N_A_597_125#_M1011_s VNB NSHORT L=0.15
+ W=0.64 AD=0.1817 AS=0.0896 PD=1.85 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75003.5 A=0.096 P=1.58 MULT=1
MM1013 N_A_597_125#_M1011_s N_C1_M1013_g N_A_91_48#_M1013_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75003.1 A=0.096 P=1.58 MULT=1
MM1021 N_A_597_125#_M1021_d N_C1_M1021_g N_A_91_48#_M1013_s VNB NSHORT L=0.15
+ W=0.64 AD=0.112 AS=0.0896 PD=0.99 PS=0.92 NRD=13.116 NRS=0 M=1 R=4.26667
+ SA=75001.1 SB=75002.7 A=0.096 P=1.58 MULT=1
MM1018 N_A_510_125#_M1018_d N_B1_M1018_g N_A_597_125#_M1021_d VNB NSHORT L=0.15
+ W=0.64 AD=0.1152 AS=0.112 PD=1 PS=0.99 NRD=0 NRS=0 M=1 R=4.26667 SA=75001.6
+ SB=75002.2 A=0.096 P=1.58 MULT=1
MM1006 N_VGND_M1006_d N_A1_M1006_g N_A_510_125#_M1018_d VNB NSHORT L=0.15 W=0.64
+ AD=0.0992 AS=0.1152 PD=0.95 PS=1 NRD=0.936 NRS=14.988 M=1 R=4.26667 SA=75002.1
+ SB=75001.7 A=0.096 P=1.58 MULT=1
MM1002 N_A_510_125#_M1002_d N_A2_M1002_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.64
+ AD=0.1072 AS=0.0992 PD=0.975 PS=0.95 NRD=10.308 NRS=4.68 M=1 R=4.26667
+ SA=75002.5 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1019 N_A_510_125#_M1002_d N_A2_M1019_g N_VGND_M1019_s VNB NSHORT L=0.15 W=0.64
+ AD=0.1072 AS=0.112 PD=0.975 PS=0.99 NRD=0 NRS=0 M=1 R=4.26667 SA=75003
+ SB=75000.7 A=0.096 P=1.58 MULT=1
MM1020 N_VGND_M1019_s N_A1_M1020_g N_A_510_125#_M1020_s VNB NSHORT L=0.15 W=0.64
+ AD=0.112 AS=0.1824 PD=0.99 PS=1.85 NRD=13.116 NRS=0 M=1 R=4.26667 SA=75003.5
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1008 N_VPWR_M1008_d N_A_91_48#_M1008_g N_X_M1008_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3864 AS=0.168 PD=2.93 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75000.3 SB=75004.8 A=0.168 P=2.54 MULT=1
MM1012 N_VPWR_M1012_d N_A_91_48#_M1012_g N_X_M1008_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.224 AS=0.168 PD=1.52 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75004.4 A=0.168 P=2.54 MULT=1
MM1017 N_VPWR_M1012_d N_A_91_48#_M1017_g N_X_M1017_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.224 AS=0.168 PD=1.52 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75001.3 SB=75003.8 A=0.168 P=2.54 MULT=1
MM1022 N_VPWR_M1022_d N_A_91_48#_M1022_g N_X_M1017_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.318743 AS=0.168 PD=1.92 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75001.7 SB=75003.4 A=0.168 P=2.54 MULT=1
MM1003 N_A_91_48#_M1003_d N_B1_M1003_g N_VPWR_M1022_d VPB PHIGHVT L=0.15 W=0.84
+ AD=0.126 AS=0.239057 PD=1.14 PS=1.44 NRD=2.3443 NRS=52.1656 M=1 R=5.6
+ SA=75002.4 SB=75003.7 A=0.126 P=1.98 MULT=1
MM1004 N_A_91_48#_M1003_d N_C1_M1004_g N_VPWR_M1004_s VPB PHIGHVT L=0.15 W=0.84
+ AD=0.126 AS=0.1743 PD=1.14 PS=1.255 NRD=2.3443 NRS=14.0658 M=1 R=5.6
+ SA=75002.9 SB=75003.3 A=0.126 P=1.98 MULT=1
MM1009 N_A_91_48#_M1009_d N_C1_M1009_g N_VPWR_M1004_s VPB PHIGHVT L=0.15 W=0.84
+ AD=0.126 AS=0.1743 PD=1.14 PS=1.255 NRD=2.3443 NRS=17.5724 M=1 R=5.6
+ SA=75003.4 SB=75002.7 A=0.126 P=1.98 MULT=1
MM1010 N_A_91_48#_M1009_d N_B1_M1010_g N_VPWR_M1010_s VPB PHIGHVT L=0.15 W=0.84
+ AD=0.126 AS=0.192013 PD=1.14 PS=1.31022 NRD=2.3443 NRS=22.852 M=1 R=5.6
+ SA=75003.9 SB=75002.3 A=0.126 P=1.98 MULT=1
MM1000 N_A_968_391#_M1000_d N_A1_M1000_g N_VPWR_M1010_s VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.228587 PD=1.3 PS=1.55978 NRD=1.9503 NRS=11.8003 M=1 R=6.66667
+ SA=75003.8 SB=75001.7 A=0.15 P=2.3 MULT=1
MM1001 N_A_91_48#_M1001_d N_A2_M1001_g N_A_968_391#_M1000_d VPB PHIGHVT L=0.15
+ W=1 AD=0.175 AS=0.15 PD=1.35 PS=1.3 NRD=11.8003 NRS=1.9503 M=1 R=6.66667
+ SA=75004.3 SB=75001.2 A=0.15 P=2.3 MULT=1
MM1005 N_A_91_48#_M1001_d N_A2_M1005_g N_A_968_391#_M1005_s VPB PHIGHVT L=0.15
+ W=1 AD=0.175 AS=0.15 PD=1.35 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75004.8 SB=75000.7 A=0.15 P=2.3 MULT=1
MM1014 N_A_968_391#_M1005_s N_A1_M1014_g N_VPWR_M1014_s VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.345 PD=1.3 PS=2.69 NRD=1.9503 NRS=11.8003 M=1 R=6.66667
+ SA=75005.2 SB=75000.3 A=0.15 P=2.3 MULT=1
DX24_noxref VNB VPB NWDIODE A=13.206 P=17.92
*
.include "sky130_fd_sc_ls__o211a_4.pxi.spice"
*
.ends
*
*
