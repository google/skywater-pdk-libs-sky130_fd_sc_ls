* File: sky130_fd_sc_ls__decap_8.pex.spice
* Created: Wed Sep  2 10:59:26 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__DECAP_8%VGND 1 12 17 21 24 25 29 32 35 36 39 42 43
+ 45 47 53 62 68 69 72 75
r46 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r47 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r48 69 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r49 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r50 66 75 12.7913 $w=1.7e-07 $l=3.1e-07 $layer=LI1_cond $X=3.29 $Y=0 $X2=2.98
+ $Y2=0
r51 66 68 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=3.29 $Y=0 $X2=3.6
+ $Y2=0
r52 65 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r53 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r54 62 75 12.7913 $w=1.7e-07 $l=3.1e-07 $layer=LI1_cond $X=2.67 $Y=0 $X2=2.98
+ $Y2=0
r55 62 64 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=2.67 $Y=0 $X2=2.64
+ $Y2=0
r56 61 73 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r57 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r58 58 72 12.1365 $w=1.7e-07 $l=2.83e-07 $layer=LI1_cond $X=1.13 $Y=0 $X2=0.847
+ $Y2=0
r59 58 60 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=1.13 $Y=0 $X2=1.68
+ $Y2=0
r60 56 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r61 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r62 53 72 12.1365 $w=1.7e-07 $l=2.82e-07 $layer=LI1_cond $X=0.565 $Y=0 $X2=0.847
+ $Y2=0
r63 53 55 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.565 $Y=0 $X2=0.24
+ $Y2=0
r64 47 65 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.64
+ $Y2=0
r65 47 61 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r66 45 46 4.71681 $w=6.18e-07 $l=1.7e-07 $layer=LI1_cond $X=2.98 $Y=0.64
+ $X2=2.98 $Y2=0.81
r67 42 60 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.765 $Y=0 $X2=1.68
+ $Y2=0
r68 42 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.765 $Y=0 $X2=1.93
+ $Y2=0
r69 41 64 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=2.095 $Y=0 $X2=2.64
+ $Y2=0
r70 41 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.095 $Y=0 $X2=1.93
+ $Y2=0
r71 39 40 5.65072 $w=5.63e-07 $l=1.7e-07 $layer=LI1_cond $X=0.847 $Y=0.64
+ $X2=0.847 $Y2=0.81
r72 35 46 17.3578 $w=4.03e-07 $l=6.1e-07 $layer=LI1_cond $X=2.872 $Y=1.42
+ $X2=2.872 $Y2=0.81
r73 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.91
+ $Y=1.42 $X2=2.91 $Y2=1.42
r74 32 45 2.70082 $w=6.18e-07 $l=1.4e-07 $layer=LI1_cond $X=2.98 $Y=0.5 $X2=2.98
+ $Y2=0.64
r75 31 75 2.59604 $w=6.2e-07 $l=8.5e-08 $layer=LI1_cond $X=2.98 $Y=0.085
+ $X2=2.98 $Y2=0
r76 31 32 8.00601 $w=6.18e-07 $l=4.15e-07 $layer=LI1_cond $X=2.98 $Y=0.085
+ $X2=2.98 $Y2=0.5
r77 27 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.93 $Y=0.085
+ $X2=1.93 $Y2=0
r78 27 29 19.382 $w=3.28e-07 $l=5.55e-07 $layer=LI1_cond $X=1.93 $Y=0.085
+ $X2=1.93 $Y2=0.64
r79 24 40 21.3027 $w=3.28e-07 $l=6.1e-07 $layer=LI1_cond $X=0.965 $Y=1.42
+ $X2=0.965 $Y2=0.81
r80 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.965
+ $Y=1.42 $X2=0.965 $Y2=1.42
r81 21 39 2.37099 $w=5.63e-07 $l=1.12e-07 $layer=LI1_cond $X=0.847 $Y=0.528
+ $X2=0.847 $Y2=0.64
r82 20 72 2.37858 $w=5.65e-07 $l=8.5e-08 $layer=LI1_cond $X=0.847 $Y=0.085
+ $X2=0.847 $Y2=0
r83 20 21 9.3781 $w=5.63e-07 $l=4.43e-07 $layer=LI1_cond $X=0.847 $Y=0.085
+ $X2=0.847 $Y2=0.528
r84 18 36 71.6931 $w=3.3e-07 $l=4.1e-07 $layer=POLY_cond $X=2.91 $Y=1.83
+ $X2=2.91 $Y2=1.42
r85 17 18 57.2398 $w=1e-06 $l=6.3e-07 $layer=POLY_cond $X=2.575 $Y=2.46
+ $X2=2.575 $Y2=1.83
r86 13 25 71.6931 $w=3.3e-07 $l=4.1e-07 $layer=POLY_cond $X=0.965 $Y=1.83
+ $X2=0.965 $Y2=1.42
r87 12 13 57.2398 $w=1e-06 $l=6.3e-07 $layer=POLY_cond $X=1.3 $Y=2.46 $X2=1.3
+ $Y2=1.83
r88 1 45 182 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=1 $X=3.065
+ $Y=0.425 $X2=3.205 $Y2=0.64
r89 1 39 182 $w=1.7e-07 $l=5.36843e-07 $layer=licon1_NDIFF $count=1 $X=1.79
+ $Y=0.425 $X2=0.65 $Y2=0.64
r90 1 29 182 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=1 $X=1.79
+ $Y=0.425 $X2=1.93 $Y2=0.64
.ends

.subckt PM_SKY130_FD_SC_LS__DECAP_8%VPWR 1 12 16 17 23 27 29 32 35 36 41 48 49
+ 52 55 58
r41 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r42 56 59 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r43 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r44 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r45 49 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r46 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r47 46 58 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.3 $Y=3.33
+ $X2=3.175 $Y2=3.33
r48 46 48 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=3.3 $Y=3.33 $X2=3.6
+ $Y2=3.33
r49 45 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r50 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r51 42 52 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.815 $Y=3.33
+ $X2=0.69 $Y2=3.33
r52 42 44 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.815 $Y=3.33
+ $X2=1.2 $Y2=3.33
r53 41 55 15.7884 $w=1.7e-07 $l=4.67e-07 $layer=LI1_cond $X=1.46 $Y=3.33
+ $X2=1.927 $Y2=3.33
r54 41 44 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=1.46 $Y=3.33 $X2=1.2
+ $Y2=3.33
r55 39 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r56 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r57 36 52 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.69 $Y2=3.33
r58 36 38 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.24 $Y2=3.33
r59 29 56 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.16 $Y2=3.33
r60 29 45 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.2 $Y2=3.33
r61 25 58 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.175 $Y=3.245
+ $X2=3.175 $Y2=3.33
r62 25 27 36.1867 $w=2.48e-07 $l=7.85e-07 $layer=LI1_cond $X=3.175 $Y=3.245
+ $X2=3.175 $Y2=2.46
r63 24 55 15.7884 $w=1.7e-07 $l=4.68e-07 $layer=LI1_cond $X=2.395 $Y=3.33
+ $X2=1.927 $Y2=3.33
r64 23 58 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.05 $Y=3.33
+ $X2=3.175 $Y2=3.33
r65 23 24 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=3.05 $Y=3.33
+ $X2=2.395 $Y2=3.33
r66 20 22 9.26417 $w=9.33e-07 $l=7.1e-07 $layer=LI1_cond $X=1.927 $Y=2.105
+ $X2=1.927 $Y2=2.815
r67 17 35 17.6663 $w=9.14e-07 $l=3.35e-07 $layer=POLY_cond $X=2.23 $Y=0.712
+ $X2=2.565 $Y2=0.712
r68 17 32 49.5711 $w=9.14e-07 $l=9.4e-07 $layer=POLY_cond $X=2.23 $Y=0.712
+ $X2=1.29 $Y2=0.712
r69 16 20 9.00321 $w=9.33e-07 $l=6.9e-07 $layer=LI1_cond $X=1.927 $Y=1.415
+ $X2=1.927 $Y2=2.105
r70 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.23
+ $Y=1.415 $X2=2.23 $Y2=1.415
r71 14 55 3.4167 $w=9.35e-07 $l=8.5e-08 $layer=LI1_cond $X=1.927 $Y=3.245
+ $X2=1.927 $Y2=3.33
r72 14 22 5.6107 $w=9.33e-07 $l=4.3e-07 $layer=LI1_cond $X=1.927 $Y=3.245
+ $X2=1.927 $Y2=2.815
r73 10 52 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=3.245
+ $X2=0.69 $Y2=3.33
r74 10 12 36.1867 $w=2.48e-07 $l=7.85e-07 $layer=LI1_cond $X=0.69 $Y=3.245
+ $X2=0.69 $Y2=2.46
r75 1 27 300 $w=1.7e-07 $l=5.65685e-07 $layer=licon1_PDIFF $count=2 $X=3.075
+ $Y=1.96 $X2=3.215 $Y2=2.46
r76 1 22 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.8
+ $Y=1.96 $X2=1.94 $Y2=2.815
r77 1 20 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.8
+ $Y=1.96 $X2=1.94 $Y2=2.105
r78 1 12 300 $w=1.7e-07 $l=7.22997e-07 $layer=licon1_PDIFF $count=2 $X=1.8
+ $Y=1.96 $X2=0.65 $Y2=2.46
.ends

