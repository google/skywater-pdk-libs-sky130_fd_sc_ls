# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ls__sdfstp_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ls__sdfstp_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  15.84000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.105000 1.820000 1.575000 2.150000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  1.201100 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.895000 0.350000 14.225000 0.980000 ;
        RECT 13.895000 0.980000 15.225000 1.150000 ;
        RECT 14.045000 1.820000 15.195000 2.150000 ;
        RECT 14.045000 2.150000 14.325000 2.980000 ;
        RECT 14.895000 0.350000 15.225000 0.980000 ;
        RECT 14.895000 1.150000 15.225000 1.270000 ;
        RECT 14.895000 1.270000 15.715000 1.440000 ;
        RECT 15.025000 1.610000 15.715000 1.780000 ;
        RECT 15.025000 1.780000 15.195000 1.820000 ;
        RECT 15.025000 2.150000 15.195000 2.980000 ;
        RECT 15.485000 1.440000 15.715000 1.610000 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.555000 1.100000 2.835000 2.150000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.525000 1.410000 2.045000 1.580000 ;
        RECT 0.525000 1.580000 0.855000 2.150000 ;
        RECT 1.715000 1.250000 2.045000 1.410000 ;
    END
  END SCE
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  7.195000 1.450000  7.555000 1.780000 ;
        RECT 11.470000 1.470000 11.870000 2.140000 ;
      LAYER mcon ;
        RECT  7.355000 1.580000  7.525000 1.750000 ;
        RECT 11.675000 1.580000 11.845000 1.750000 ;
      LAYER met1 ;
        RECT  7.295000 1.550000  7.585000 1.595000 ;
        RECT  7.295000 1.595000 11.905000 1.735000 ;
        RECT  7.295000 1.735000  7.585000 1.780000 ;
        RECT 11.615000 1.550000 11.905000 1.595000 ;
        RECT 11.615000 1.735000 11.905000 1.780000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.345000 1.180000 3.715000 1.550000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 15.840000 0.085000 ;
        RECT  0.615000  0.085000  0.945000 0.740000 ;
        RECT  2.450000  0.085000  2.780000 0.740000 ;
        RECT  3.560000  0.085000  3.890000 1.010000 ;
        RECT  6.210000  0.085000  6.540000 0.600000 ;
        RECT  7.590000  0.085000  8.260000 0.930000 ;
        RECT  8.790000  0.085000  9.120000 0.940000 ;
        RECT 11.650000  0.085000 12.150000 0.680000 ;
        RECT 13.380000  0.085000 13.710000 1.130000 ;
        RECT 14.395000  0.085000 14.725000 0.810000 ;
        RECT 15.395000  0.085000 15.725000 1.100000 ;
      LAYER mcon ;
        RECT  0.155000 -0.085000  0.325000 0.085000 ;
        RECT  0.635000 -0.085000  0.805000 0.085000 ;
        RECT  1.115000 -0.085000  1.285000 0.085000 ;
        RECT  1.595000 -0.085000  1.765000 0.085000 ;
        RECT  2.075000 -0.085000  2.245000 0.085000 ;
        RECT  2.555000 -0.085000  2.725000 0.085000 ;
        RECT  3.035000 -0.085000  3.205000 0.085000 ;
        RECT  3.515000 -0.085000  3.685000 0.085000 ;
        RECT  3.995000 -0.085000  4.165000 0.085000 ;
        RECT  4.475000 -0.085000  4.645000 0.085000 ;
        RECT  4.955000 -0.085000  5.125000 0.085000 ;
        RECT  5.435000 -0.085000  5.605000 0.085000 ;
        RECT  5.915000 -0.085000  6.085000 0.085000 ;
        RECT  6.395000 -0.085000  6.565000 0.085000 ;
        RECT  6.875000 -0.085000  7.045000 0.085000 ;
        RECT  7.355000 -0.085000  7.525000 0.085000 ;
        RECT  7.835000 -0.085000  8.005000 0.085000 ;
        RECT  8.315000 -0.085000  8.485000 0.085000 ;
        RECT  8.795000 -0.085000  8.965000 0.085000 ;
        RECT  9.275000 -0.085000  9.445000 0.085000 ;
        RECT  9.755000 -0.085000  9.925000 0.085000 ;
        RECT 10.235000 -0.085000 10.405000 0.085000 ;
        RECT 10.715000 -0.085000 10.885000 0.085000 ;
        RECT 11.195000 -0.085000 11.365000 0.085000 ;
        RECT 11.675000 -0.085000 11.845000 0.085000 ;
        RECT 12.155000 -0.085000 12.325000 0.085000 ;
        RECT 12.635000 -0.085000 12.805000 0.085000 ;
        RECT 13.115000 -0.085000 13.285000 0.085000 ;
        RECT 13.595000 -0.085000 13.765000 0.085000 ;
        RECT 14.075000 -0.085000 14.245000 0.085000 ;
        RECT 14.555000 -0.085000 14.725000 0.085000 ;
        RECT 15.035000 -0.085000 15.205000 0.085000 ;
        RECT 15.515000 -0.085000 15.685000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 15.840000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 3.245000 15.840000 3.415000 ;
        RECT  0.555000 2.660000  0.885000 3.245000 ;
        RECT  2.560000 2.830000  2.890000 3.245000 ;
        RECT  3.570000 2.580000  3.900000 3.245000 ;
        RECT  6.275000 2.630000  6.525000 3.245000 ;
        RECT  7.715000 2.290000  7.885000 3.245000 ;
        RECT  8.535000 2.460000  8.865000 3.245000 ;
        RECT 11.125000 2.650000 11.375000 3.245000 ;
        RECT 12.720000 2.520000 12.970000 3.245000 ;
        RECT 13.540000 2.100000 13.870000 3.245000 ;
        RECT 14.495000 2.320000 14.825000 3.245000 ;
        RECT 15.395000 1.950000 15.725000 3.245000 ;
      LAYER mcon ;
        RECT  0.155000 3.245000  0.325000 3.415000 ;
        RECT  0.635000 3.245000  0.805000 3.415000 ;
        RECT  1.115000 3.245000  1.285000 3.415000 ;
        RECT  1.595000 3.245000  1.765000 3.415000 ;
        RECT  2.075000 3.245000  2.245000 3.415000 ;
        RECT  2.555000 3.245000  2.725000 3.415000 ;
        RECT  3.035000 3.245000  3.205000 3.415000 ;
        RECT  3.515000 3.245000  3.685000 3.415000 ;
        RECT  3.995000 3.245000  4.165000 3.415000 ;
        RECT  4.475000 3.245000  4.645000 3.415000 ;
        RECT  4.955000 3.245000  5.125000 3.415000 ;
        RECT  5.435000 3.245000  5.605000 3.415000 ;
        RECT  5.915000 3.245000  6.085000 3.415000 ;
        RECT  6.395000 3.245000  6.565000 3.415000 ;
        RECT  6.875000 3.245000  7.045000 3.415000 ;
        RECT  7.355000 3.245000  7.525000 3.415000 ;
        RECT  7.835000 3.245000  8.005000 3.415000 ;
        RECT  8.315000 3.245000  8.485000 3.415000 ;
        RECT  8.795000 3.245000  8.965000 3.415000 ;
        RECT  9.275000 3.245000  9.445000 3.415000 ;
        RECT  9.755000 3.245000  9.925000 3.415000 ;
        RECT 10.235000 3.245000 10.405000 3.415000 ;
        RECT 10.715000 3.245000 10.885000 3.415000 ;
        RECT 11.195000 3.245000 11.365000 3.415000 ;
        RECT 11.675000 3.245000 11.845000 3.415000 ;
        RECT 12.155000 3.245000 12.325000 3.415000 ;
        RECT 12.635000 3.245000 12.805000 3.415000 ;
        RECT 13.115000 3.245000 13.285000 3.415000 ;
        RECT 13.595000 3.245000 13.765000 3.415000 ;
        RECT 14.075000 3.245000 14.245000 3.415000 ;
        RECT 14.555000 3.245000 14.725000 3.415000 ;
        RECT 15.035000 3.245000 15.205000 3.415000 ;
        RECT 15.515000 3.245000 15.685000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 15.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.105000 0.350000  0.445000 0.910000 ;
      RECT  0.105000 0.910000  1.140000 1.240000 ;
      RECT  0.105000 1.240000  0.355000 2.320000 ;
      RECT  0.105000 2.320000  2.045000 2.490000 ;
      RECT  0.105000 2.490000  0.355000 2.980000 ;
      RECT  1.425000 2.660000  2.385000 2.910000 ;
      RECT  1.475000 0.410000  1.960000 0.740000 ;
      RECT  1.785000 1.830000  2.045000 2.320000 ;
      RECT  1.790000 0.740000  1.960000 0.910000 ;
      RECT  1.790000 0.910000  2.385000 1.080000 ;
      RECT  2.215000 1.080000  2.385000 2.490000 ;
      RECT  2.215000 2.490000  3.175000 2.660000 ;
      RECT  3.005000 0.350000  3.390000 1.010000 ;
      RECT  3.005000 1.010000  3.175000 1.820000 ;
      RECT  3.005000 1.820000  4.215000 2.070000 ;
      RECT  3.005000 2.240000  5.030000 2.410000 ;
      RECT  3.005000 2.410000  3.175000 2.490000 ;
      RECT  3.885000 1.350000  4.215000 1.820000 ;
      RECT  4.070000 0.255000  5.140000 0.425000 ;
      RECT  4.070000 0.425000  4.240000 1.130000 ;
      RECT  4.070000 2.580000  4.400000 2.895000 ;
      RECT  4.070000 2.895000  5.830000 3.065000 ;
      RECT  4.410000 0.595000  4.800000 0.925000 ;
      RECT  4.410000 0.925000  4.580000 1.900000 ;
      RECT  4.410000 1.900000  5.030000 2.240000 ;
      RECT  4.700000 2.410000  5.030000 2.725000 ;
      RECT  4.750000 1.095000  5.140000 1.265000 ;
      RECT  4.750000 1.265000  5.030000 1.730000 ;
      RECT  4.970000 0.425000  5.140000 1.095000 ;
      RECT  5.200000 1.435000  6.955000 1.605000 ;
      RECT  5.200000 1.605000  5.370000 2.275000 ;
      RECT  5.200000 2.275000  5.480000 2.725000 ;
      RECT  5.310000 0.385000  5.640000 1.435000 ;
      RECT  5.540000 1.775000  5.830000 2.105000 ;
      RECT  5.660000 2.105000  5.830000 2.290000 ;
      RECT  5.660000 2.290000  6.865000 2.460000 ;
      RECT  5.660000 2.460000  5.830000 2.895000 ;
      RECT  6.005000 0.770000  7.100000 0.940000 ;
      RECT  6.005000 0.940000  6.335000 1.265000 ;
      RECT  6.040000 1.780000  6.370000 1.950000 ;
      RECT  6.040000 1.950000  7.205000 2.120000 ;
      RECT  6.625000 1.110000  8.265000 1.280000 ;
      RECT  6.625000 1.280000  6.955000 1.435000 ;
      RECT  6.625000 1.605000  6.955000 1.780000 ;
      RECT  6.695000 2.460000  6.865000 2.895000 ;
      RECT  6.695000 2.895000  7.545000 3.065000 ;
      RECT  6.770000 0.350000  7.100000 0.770000 ;
      RECT  7.035000 2.120000  7.205000 2.725000 ;
      RECT  7.375000 1.950000  7.895000 2.120000 ;
      RECT  7.375000 2.120000  7.545000 2.895000 ;
      RECT  7.725000 1.780000 10.765000 1.930000 ;
      RECT  7.725000 1.930000  9.375000 1.950000 ;
      RECT  7.935000 1.280000  8.265000 1.450000 ;
      RECT  8.085000 2.120000  9.875000 2.290000 ;
      RECT  8.085000 2.290000  8.365000 2.715000 ;
      RECT  8.440000 0.350000  8.610000 1.110000 ;
      RECT  8.440000 1.110000 10.030000 1.280000 ;
      RECT  9.045000 1.450000  9.375000 1.760000 ;
      RECT  9.045000 1.760000 10.765000 1.780000 ;
      RECT  9.095000 2.600000  9.375000 2.860000 ;
      RECT  9.095000 2.860000 10.375000 3.075000 ;
      RECT  9.350000 0.255000 10.540000 0.425000 ;
      RECT  9.350000 0.425000  9.680000 0.940000 ;
      RECT  9.545000 2.100000  9.875000 2.120000 ;
      RECT  9.545000 2.290000  9.875000 2.690000 ;
      RECT  9.860000 0.595000 10.030000 1.110000 ;
      RECT 10.045000 2.310000 12.210000 2.480000 ;
      RECT 10.045000 2.480000 10.375000 2.860000 ;
      RECT 10.210000 0.425000 10.540000 1.400000 ;
      RECT 10.210000 1.400000 11.105000 1.570000 ;
      RECT 10.435000 1.930000 10.765000 2.135000 ;
      RECT 10.545000 2.650000 10.955000 2.980000 ;
      RECT 10.935000 1.570000 11.105000 2.310000 ;
      RECT 10.955000 0.900000 12.710000 1.070000 ;
      RECT 10.955000 1.070000 11.285000 1.230000 ;
      RECT 11.575000 2.480000 11.905000 2.980000 ;
      RECT 12.040000 1.340000 12.370000 2.010000 ;
      RECT 12.040000 2.010000 12.210000 2.310000 ;
      RECT 12.135000 2.650000 12.550000 2.980000 ;
      RECT 12.320000 0.350000 12.710000 0.900000 ;
      RECT 12.380000 2.180000 12.710000 2.350000 ;
      RECT 12.380000 2.350000 12.550000 2.650000 ;
      RECT 12.540000 1.070000 12.710000 2.180000 ;
      RECT 12.880000 0.350000 13.210000 1.320000 ;
      RECT 12.880000 1.320000 14.695000 1.490000 ;
      RECT 13.170000 1.490000 14.695000 1.650000 ;
      RECT 13.170000 1.650000 13.340000 2.980000 ;
  END
END sky130_fd_sc_ls__sdfstp_4
