* File: sky130_fd_sc_ls__o311a_2.pex.spice
* Created: Wed Sep  2 11:21:20 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__O311A_2%C1 3 4 6 8 9 10
c27 4 0 4.75566e-20 $X=0.615 $Y=1.765
r28 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.385 $X2=0.27 $Y2=1.385
r29 10 14 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.27 $Y=1.295 $X2=0.27
+ $Y2=1.385
r30 8 13 44.5896 $w=3.3e-07 $l=2.55e-07 $layer=POLY_cond $X=0.525 $Y=1.385
+ $X2=0.27 $Y2=1.385
r31 8 9 66.2869 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.615 $Y=1.385
+ $X2=0.615 $Y2=1.22
r32 4 8 149.859 $w=1.8e-07 $l=3.8e-07 $layer=POLY_cond $X=0.615 $Y=1.765
+ $X2=0.615 $Y2=1.385
r33 4 6 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.615 $Y=1.765
+ $X2=0.615 $Y2=2.34
r34 3 9 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.6 $Y=0.74 $X2=0.6
+ $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_LS__O311A_2%B1 3 5 7 8 12
c32 12 0 4.75566e-20 $X=1.11 $Y=1.515
c33 5 0 1.35203e-19 $X=1.185 $Y=1.765
r34 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.11
+ $Y=1.515 $X2=1.11 $Y2=1.515
r35 8 12 4.67207 $w=3.68e-07 $l=1.5e-07 $layer=LI1_cond $X=1.13 $Y=1.665
+ $X2=1.13 $Y2=1.515
r36 5 11 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=1.185 $Y=1.765
+ $X2=1.11 $Y2=1.515
r37 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.185 $Y=1.765
+ $X2=1.185 $Y2=2.34
r38 1 11 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=1.02 $Y=1.35
+ $X2=1.11 $Y2=1.515
r39 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.02 $Y=1.35 $X2=1.02
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__O311A_2%A3 3 5 7 8 12
r30 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.65
+ $Y=1.515 $X2=1.65 $Y2=1.515
r31 8 12 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.65 $Y=1.665
+ $X2=1.65 $Y2=1.515
r32 5 11 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=1.725 $Y=1.765
+ $X2=1.65 $Y2=1.515
r33 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.725 $Y=1.765
+ $X2=1.725 $Y2=2.4
r34 1 11 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=1.56 $Y=1.35
+ $X2=1.65 $Y2=1.515
r35 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.56 $Y=1.35 $X2=1.56
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__O311A_2%A2 1 3 6 8 9 10 11 18
c32 1 0 1.68448e-19 $X=2.145 $Y=1.765
r33 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.19
+ $Y=1.515 $X2=2.19 $Y2=1.515
r34 10 11 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.19 $Y=2.405
+ $X2=2.19 $Y2=2.775
r35 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.19 $Y=2.035
+ $X2=2.19 $Y2=2.405
r36 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.19 $Y=1.665 $X2=2.19
+ $Y2=2.035
r37 8 18 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=2.19 $Y=1.665
+ $X2=2.19 $Y2=1.515
r38 4 17 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=2.28 $Y=1.35
+ $X2=2.19 $Y2=1.515
r39 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.28 $Y=1.35 $X2=2.28
+ $Y2=0.74
r40 1 17 52.2586 $w=2.99e-07 $l=2.7157e-07 $layer=POLY_cond $X=2.145 $Y=1.765
+ $X2=2.19 $Y2=1.515
r41 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.145 $Y=1.765
+ $X2=2.145 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__O311A_2%A1 1 3 6 8 12
c29 12 0 1.28711e-19 $X=2.76 $Y=1.515
c30 6 0 3.01101e-20 $X=2.71 $Y=0.74
r31 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.76
+ $Y=1.515 $X2=2.76 $Y2=1.515
r32 8 12 4.32166 $w=3.98e-07 $l=1.5e-07 $layer=LI1_cond $X=2.725 $Y=1.665
+ $X2=2.725 $Y2=1.515
r33 4 11 38.5562 $w=2.99e-07 $l=1.88348e-07 $layer=POLY_cond $X=2.71 $Y=1.35
+ $X2=2.76 $Y2=1.515
r34 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.71 $Y=1.35 $X2=2.71
+ $Y2=0.74
r35 1 11 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=2.685 $Y=1.765
+ $X2=2.76 $Y2=1.515
r36 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.685 $Y=1.765
+ $X2=2.685 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__O311A_2%A_32_74# 1 2 3 10 12 13 15 16 18 19 21 24 26
+ 28 30 32 34 40 41 53
c103 40 0 1.35203e-19 $X=0.39 $Y=1.985
c104 32 0 1.68448e-19 $X=1.5 $Y=2.12
c105 13 0 1.73007e-19 $X=3.305 $Y=1.22
c106 10 0 1.28711e-19 $X=3.27 $Y=1.765
r107 53 54 1.59956 $w=4.52e-07 $l=1.5e-08 $layer=POLY_cond $X=3.72 $Y=1.492
+ $X2=3.735 $Y2=1.492
r108 50 51 3.7323 $w=4.52e-07 $l=3.5e-08 $layer=POLY_cond $X=3.27 $Y=1.492
+ $X2=3.305 $Y2=1.492
r109 49 53 39.9889 $w=4.52e-07 $l=3.75e-07 $layer=POLY_cond $X=3.345 $Y=1.492
+ $X2=3.72 $Y2=1.492
r110 49 51 4.26549 $w=4.52e-07 $l=4e-08 $layer=POLY_cond $X=3.345 $Y=1.492
+ $X2=3.305 $Y2=1.492
r111 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.345
+ $Y=1.385 $X2=3.345 $Y2=1.385
r112 42 43 3.00192 $w=5.48e-07 $l=8.5e-08 $layer=LI1_cond $X=0.5 $Y=2.035
+ $X2=0.5 $Y2=2.12
r113 40 42 1.08734 $w=5.48e-07 $l=5e-08 $layer=LI1_cond $X=0.5 $Y=1.985 $X2=0.5
+ $Y2=2.035
r114 40 41 9.83198 $w=5.48e-07 $l=1.65e-07 $layer=LI1_cond $X=0.5 $Y=1.985
+ $X2=0.5 $Y2=1.82
r115 32 45 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.5 $Y=2.12 $X2=1.5
+ $Y2=2.035
r116 32 34 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=1.5 $Y=2.12
+ $X2=1.5 $Y2=2.815
r117 31 42 7.75927 $w=1.7e-07 $l=2.75e-07 $layer=LI1_cond $X=0.775 $Y=2.035
+ $X2=0.5 $Y2=2.035
r118 30 45 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.335 $Y=2.035
+ $X2=1.5 $Y2=2.035
r119 30 31 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.335 $Y=2.035
+ $X2=0.775 $Y2=2.035
r120 29 37 14.5 $w=4.88e-07 $l=7.08308e-07 $layer=LI1_cond $X=0.775 $Y=1.095
+ $X2=0.49 $Y2=0.515
r121 28 48 11.0909 $w=3.19e-07 $l=3.79645e-07 $layer=LI1_cond $X=3.095 $Y=1.095
+ $X2=3.302 $Y2=1.385
r122 28 29 151.358 $w=1.68e-07 $l=2.32e-06 $layer=LI1_cond $X=3.095 $Y=1.095
+ $X2=0.775 $Y2=1.095
r123 26 29 7.63306 $w=4.88e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.69 $Y=1.18
+ $X2=0.775 $Y2=1.095
r124 26 41 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=0.69 $Y=1.18
+ $X2=0.69 $Y2=1.82
r125 24 43 17.4383 $w=3.78e-07 $l=5.75e-07 $layer=LI1_cond $X=0.415 $Y=2.695
+ $X2=0.415 $Y2=2.12
r126 19 54 28.877 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=3.735 $Y=1.22
+ $X2=3.735 $Y2=1.492
r127 19 21 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.735 $Y=1.22
+ $X2=3.735 $Y2=0.74
r128 16 53 28.877 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=3.72 $Y=1.765
+ $X2=3.72 $Y2=1.492
r129 16 18 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.72 $Y=1.765
+ $X2=3.72 $Y2=2.4
r130 13 51 28.877 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=3.305 $Y=1.22
+ $X2=3.305 $Y2=1.492
r131 13 15 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.305 $Y=1.22
+ $X2=3.305 $Y2=0.74
r132 10 50 28.877 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=3.27 $Y=1.765
+ $X2=3.27 $Y2=1.492
r133 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.27 $Y=1.765
+ $X2=3.27 $Y2=2.4
r134 3 45 300 $w=1.7e-07 $l=3.76331e-07 $layer=licon1_PDIFF $count=2 $X=1.26
+ $Y=1.84 $X2=1.5 $Y2=2.115
r135 3 34 600 $w=1.7e-07 $l=1.0884e-06 $layer=licon1_PDIFF $count=1 $X=1.26
+ $Y=1.84 $X2=1.5 $Y2=2.815
r136 2 40 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.245
+ $Y=1.84 $X2=0.39 $Y2=1.985
r137 2 24 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.245
+ $Y=1.84 $X2=0.39 $Y2=2.695
r138 1 37 91 $w=1.7e-07 $l=2.88531e-07 $layer=licon1_NDIFF $count=2 $X=0.16
+ $Y=0.37 $X2=0.385 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__O311A_2%VPWR 1 2 3 12 16 20 22 27 28 30 31 32 44 50
r53 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r54 47 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r55 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r56 44 49 4.64076 $w=1.7e-07 $l=2.45e-07 $layer=LI1_cond $X=3.83 $Y=3.33
+ $X2=4.075 $Y2=3.33
r57 44 46 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=3.83 $Y=3.33 $X2=3.6
+ $Y2=3.33
r58 43 47 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r59 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r60 39 42 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r61 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r62 36 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r63 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r64 32 43 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r65 32 40 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.2 $Y2=3.33
r66 30 42 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=2.745 $Y=3.33
+ $X2=2.64 $Y2=3.33
r67 30 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.745 $Y=3.33
+ $X2=2.91 $Y2=3.33
r68 29 46 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=3.075 $Y=3.33
+ $X2=3.6 $Y2=3.33
r69 29 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.075 $Y=3.33
+ $X2=2.91 $Y2=3.33
r70 27 35 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=0.775 $Y=3.33
+ $X2=0.72 $Y2=3.33
r71 27 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.775 $Y=3.33
+ $X2=0.94 $Y2=3.33
r72 26 39 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=1.105 $Y=3.33
+ $X2=1.2 $Y2=3.33
r73 26 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.105 $Y=3.33
+ $X2=0.94 $Y2=3.33
r74 22 25 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=3.995 $Y=2.145
+ $X2=3.995 $Y2=2.825
r75 20 49 3.12541 $w=3.3e-07 $l=1.18427e-07 $layer=LI1_cond $X=3.995 $Y=3.245
+ $X2=4.075 $Y2=3.33
r76 20 25 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=3.995 $Y=3.245
+ $X2=3.995 $Y2=2.825
r77 16 19 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=2.91 $Y=2.115 $X2=2.91
+ $Y2=2.815
r78 14 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.91 $Y=3.245
+ $X2=2.91 $Y2=3.33
r79 14 19 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.91 $Y=3.245
+ $X2=2.91 $Y2=2.815
r80 10 28 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.94 $Y=3.245
+ $X2=0.94 $Y2=3.33
r81 10 12 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=0.94 $Y=3.245
+ $X2=0.94 $Y2=2.375
r82 3 25 400 $w=1.7e-07 $l=1.08038e-06 $layer=licon1_PDIFF $count=1 $X=3.795
+ $Y=1.84 $X2=3.995 $Y2=2.825
r83 3 22 400 $w=1.7e-07 $l=3.9246e-07 $layer=licon1_PDIFF $count=1 $X=3.795
+ $Y=1.84 $X2=3.995 $Y2=2.145
r84 2 19 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.76
+ $Y=1.84 $X2=2.91 $Y2=2.815
r85 2 16 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=2.76
+ $Y=1.84 $X2=2.91 $Y2=2.115
r86 1 12 300 $w=1.7e-07 $l=6.48055e-07 $layer=licon1_PDIFF $count=2 $X=0.69
+ $Y=1.84 $X2=0.94 $Y2=2.375
.ends

.subckt PM_SKY130_FD_SC_LS__O311A_2%X 1 2 9 15 17 18 19 20 21 22 23 28 29 34
c45 15 0 1.73007e-19 $X=3.52 $Y=0.515
r46 29 34 2.75584 $w=2.28e-07 $l=5.5e-08 $layer=LI1_cond $X=4.08 $Y=1.72
+ $X2=4.08 $Y2=1.665
r47 23 29 2.9826 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.08 $Y=1.805 $X2=4.08
+ $Y2=1.72
r48 23 34 0.751593 $w=2.28e-07 $l=1.5e-08 $layer=LI1_cond $X=4.08 $Y=1.65
+ $X2=4.08 $Y2=1.665
r49 22 23 17.7877 $w=2.28e-07 $l=3.55e-07 $layer=LI1_cond $X=4.08 $Y=1.295
+ $X2=4.08 $Y2=1.65
r50 22 28 12.276 $w=2.28e-07 $l=2.45e-07 $layer=LI1_cond $X=4.08 $Y=1.295
+ $X2=4.08 $Y2=1.05
r51 21 28 3.48281 $w=2.3e-07 $l=1.2e-07 $layer=LI1_cond $X=4.08 $Y=0.93 $X2=4.08
+ $Y2=1.05
r52 19 21 3.33769 $w=2.4e-07 $l=1.15e-07 $layer=LI1_cond $X=3.965 $Y=0.93
+ $X2=4.08 $Y2=0.93
r53 19 20 13.4452 $w=2.38e-07 $l=2.8e-07 $layer=LI1_cond $X=3.965 $Y=0.93
+ $X2=3.685 $Y2=0.93
r54 17 23 4.03528 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=3.965 $Y=1.805
+ $X2=4.08 $Y2=1.805
r55 17 18 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.965 $Y=1.805
+ $X2=3.66 $Y2=1.805
r56 13 20 6.82018 $w=2.4e-07 $l=1.75e-07 $layer=LI1_cond $X=3.56 $Y=0.81
+ $X2=3.685 $Y2=0.93
r57 13 15 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=3.56 $Y=0.81
+ $X2=3.56 $Y2=0.515
r58 9 11 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=3.495 $Y=1.985
+ $X2=3.495 $Y2=2.815
r59 7 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.495 $Y=1.89
+ $X2=3.66 $Y2=1.805
r60 7 9 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=3.495 $Y=1.89
+ $X2=3.495 $Y2=1.985
r61 2 11 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=3.345
+ $Y=1.84 $X2=3.495 $Y2=2.815
r62 2 9 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=3.345
+ $Y=1.84 $X2=3.495 $Y2=1.985
r63 1 15 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.38
+ $Y=0.37 $X2=3.52 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__O311A_2%A_219_74# 1 2 7 10 15
c28 7 0 3.01101e-20 $X=2.33 $Y=0.755
r29 15 17 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=2.495 $Y=0.595
+ $X2=2.495 $Y2=0.755
r30 10 12 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=1.345 $Y=0.595
+ $X2=1.345 $Y2=0.755
r31 8 12 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.51 $Y=0.755
+ $X2=1.345 $Y2=0.755
r32 7 17 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.33 $Y=0.755
+ $X2=2.495 $Y2=0.755
r33 7 8 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=2.33 $Y=0.755 $X2=1.51
+ $Y2=0.755
r34 2 15 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=2.355
+ $Y=0.37 $X2=2.495 $Y2=0.595
r35 1 10 182 $w=1.7e-07 $l=3.44601e-07 $layer=licon1_NDIFF $count=1 $X=1.095
+ $Y=0.37 $X2=1.345 $Y2=0.595
.ends

.subckt PM_SKY130_FD_SC_LS__O311A_2%VGND 1 2 3 12 14 16 18 19 26 27 28 40 46
r56 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r57 43 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r58 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r59 40 45 4.9234 $w=1.7e-07 $l=2.32e-07 $layer=LI1_cond $X=3.855 $Y=0 $X2=4.087
+ $Y2=0
r60 40 42 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=3.855 $Y=0 $X2=3.6
+ $Y2=0
r61 39 43 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r62 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r63 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r64 32 36 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.68
+ $Y2=0
r65 31 35 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=1.68
+ $Y2=0
r66 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r67 28 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r68 28 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r69 26 38 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=2.83 $Y=0 $X2=2.64
+ $Y2=0
r70 26 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.83 $Y=0 $X2=2.995
+ $Y2=0
r71 25 42 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=3.16 $Y=0 $X2=3.6
+ $Y2=0
r72 25 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.16 $Y=0 $X2=2.995
+ $Y2=0
r73 21 38 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=2.15 $Y=0 $X2=2.64
+ $Y2=0
r74 19 35 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=1.69 $Y=0 $X2=1.68
+ $Y2=0
r75 18 23 8.71057 $w=4.58e-07 $l=3.35e-07 $layer=LI1_cond $X=1.92 $Y=0 $X2=1.92
+ $Y2=0.335
r76 18 21 6.6364 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=1.92 $Y=0 $X2=2.15
+ $Y2=0
r77 18 19 6.6364 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=1.92 $Y=0 $X2=1.69
+ $Y2=0
r78 14 45 3.01346 $w=3.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=4.03 $Y=0.085
+ $X2=4.087 $Y2=0
r79 14 16 14.1586 $w=3.48e-07 $l=4.3e-07 $layer=LI1_cond $X=4.03 $Y=0.085
+ $X2=4.03 $Y2=0.515
r80 10 27 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.995 $Y=0.085
+ $X2=2.995 $Y2=0
r81 10 12 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=2.995 $Y=0.085
+ $X2=2.995 $Y2=0.595
r82 3 16 182 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_NDIFF $count=1 $X=3.81
+ $Y=0.37 $X2=4.03 $Y2=0.515
r83 2 12 182 $w=1.7e-07 $l=3.1285e-07 $layer=licon1_NDIFF $count=1 $X=2.785
+ $Y=0.37 $X2=2.995 $Y2=0.595
r84 1 23 182 $w=1.7e-07 $l=3.01993e-07 $layer=licon1_NDIFF $count=1 $X=1.635
+ $Y=0.37 $X2=1.92 $Y2=0.335
.ends

