* File: sky130_fd_sc_ls__nand4_1.pxi.spice
* Created: Fri Aug 28 13:34:35 2020
* 
x_PM_SKY130_FD_SC_LS__NAND4_1%D N_D_c_43_n N_D_M1003_g N_D_c_44_n N_D_M1000_g D
+ PM_SKY130_FD_SC_LS__NAND4_1%D
x_PM_SKY130_FD_SC_LS__NAND4_1%C N_C_c_69_n N_C_M1001_g N_C_c_70_n N_C_M1005_g C
+ N_C_c_71_n PM_SKY130_FD_SC_LS__NAND4_1%C
x_PM_SKY130_FD_SC_LS__NAND4_1%B N_B_c_98_n N_B_M1002_g N_B_c_99_n N_B_M1004_g B
+ PM_SKY130_FD_SC_LS__NAND4_1%B
x_PM_SKY130_FD_SC_LS__NAND4_1%A N_A_c_129_n N_A_M1007_g N_A_c_130_n N_A_M1006_g
+ A PM_SKY130_FD_SC_LS__NAND4_1%A
x_PM_SKY130_FD_SC_LS__NAND4_1%VPWR N_VPWR_M1003_s N_VPWR_M1005_d N_VPWR_M1006_d
+ N_VPWR_c_151_n N_VPWR_c_152_n N_VPWR_c_153_n N_VPWR_c_154_n N_VPWR_c_155_n
+ N_VPWR_c_156_n N_VPWR_c_157_n N_VPWR_c_158_n VPWR N_VPWR_c_159_n
+ N_VPWR_c_150_n PM_SKY130_FD_SC_LS__NAND4_1%VPWR
x_PM_SKY130_FD_SC_LS__NAND4_1%Y N_Y_M1007_d N_Y_M1003_d N_Y_M1004_d N_Y_c_189_n
+ N_Y_c_190_n N_Y_c_191_n N_Y_c_194_n N_Y_c_195_n N_Y_c_196_n N_Y_c_197_n
+ N_Y_c_198_n N_Y_c_192_n N_Y_c_199_n N_Y_c_200_n Y
+ PM_SKY130_FD_SC_LS__NAND4_1%Y
x_PM_SKY130_FD_SC_LS__NAND4_1%VGND N_VGND_M1000_s VGND N_VGND_c_262_n
+ N_VGND_c_263_n N_VGND_c_264_n PM_SKY130_FD_SC_LS__NAND4_1%VGND
cc_1 VNB N_D_c_43_n 0.0417131f $X=-0.19 $Y=-0.245 $X2=0.815 $Y2=1.765
cc_2 VNB N_D_c_44_n 0.0194922f $X=-0.19 $Y=-0.245 $X2=0.83 $Y2=1.22
cc_3 VNB D 0.00341988f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_4 VNB N_C_c_69_n 0.0183508f $X=-0.19 $Y=-0.245 $X2=0.815 $Y2=1.765
cc_5 VNB N_C_c_70_n 0.0350896f $X=-0.19 $Y=-0.245 $X2=0.83 $Y2=1.22
cc_6 VNB N_C_c_71_n 0.00766751f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=1.385
cc_7 VNB N_B_c_98_n 0.0199072f $X=-0.19 $Y=-0.245 $X2=0.815 $Y2=1.765
cc_8 VNB N_B_c_99_n 0.0354333f $X=-0.19 $Y=-0.245 $X2=0.83 $Y2=1.22
cc_9 VNB B 0.0119609f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_10 VNB N_A_c_129_n 0.0243771f $X=-0.19 $Y=-0.245 $X2=0.815 $Y2=1.765
cc_11 VNB N_A_c_130_n 0.0686476f $X=-0.19 $Y=-0.245 $X2=0.83 $Y2=1.22
cc_12 VNB A 0.00941175f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_13 VNB N_VPWR_c_150_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_Y_c_189_n 0.0314733f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=1.385
cc_15 VNB N_Y_c_190_n 0.0122962f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=1.295
cc_16 VNB N_Y_c_191_n 0.00970183f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_Y_c_192_n 0.021252f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_VGND_c_262_n 0.0660892f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_VGND_c_263_n 0.186373f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=1.385
cc_20 VNB N_VGND_c_264_n 0.0431564f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=1.295
cc_21 VPB N_D_c_43_n 0.0240524f $X=-0.19 $Y=1.66 $X2=0.815 $Y2=1.765
cc_22 VPB N_C_c_70_n 0.0237667f $X=-0.19 $Y=1.66 $X2=0.83 $Y2=1.22
cc_23 VPB N_B_c_99_n 0.0248195f $X=-0.19 $Y=1.66 $X2=0.83 $Y2=1.22
cc_24 VPB N_A_c_130_n 0.0298134f $X=-0.19 $Y=1.66 $X2=0.83 $Y2=1.22
cc_25 VPB N_VPWR_c_151_n 0.047631f $X=-0.19 $Y=1.66 $X2=0.74 $Y2=1.295
cc_26 VPB N_VPWR_c_152_n 0.00986028f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_27 VPB N_VPWR_c_153_n 0.0120106f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_28 VPB N_VPWR_c_154_n 0.0558238f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_29 VPB N_VPWR_c_155_n 0.0140765f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_30 VPB N_VPWR_c_156_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_31 VPB N_VPWR_c_157_n 0.0194903f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_32 VPB N_VPWR_c_158_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_33 VPB N_VPWR_c_159_n 0.0196506f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_34 VPB N_VPWR_c_150_n 0.0685036f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_35 VPB N_Y_c_189_n 0.00301672f $X=-0.19 $Y=1.66 $X2=0.74 $Y2=1.385
cc_36 VPB N_Y_c_194_n 0.00729924f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_37 VPB N_Y_c_195_n 0.0138507f $X=-0.19 $Y=1.66 $X2=0.74 $Y2=1.385
cc_38 VPB N_Y_c_196_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_39 VPB N_Y_c_197_n 0.00337359f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_40 VPB N_Y_c_198_n 0.00289722f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_41 VPB N_Y_c_199_n 0.00807857f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_42 VPB N_Y_c_200_n 0.0106363f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_43 N_D_c_44_n N_C_c_69_n 0.0359258f $X=0.83 $Y=1.22 $X2=-0.19 $Y2=-0.245
cc_44 D N_C_c_69_n 4.15144e-19 $X=0.635 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_45 N_D_c_43_n N_C_c_70_n 0.0574431f $X=0.815 $Y=1.765 $X2=0 $Y2=0
cc_46 N_D_c_44_n N_C_c_71_n 0.00224093f $X=0.83 $Y=1.22 $X2=0 $Y2=0
cc_47 D N_C_c_71_n 0.0283697f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_48 N_D_c_43_n N_VPWR_c_151_n 0.0227729f $X=0.815 $Y=1.765 $X2=0 $Y2=0
cc_49 N_D_c_43_n N_VPWR_c_157_n 0.00445602f $X=0.815 $Y=1.765 $X2=0 $Y2=0
cc_50 N_D_c_43_n N_VPWR_c_150_n 0.00861803f $X=0.815 $Y=1.765 $X2=0 $Y2=0
cc_51 N_D_c_43_n N_Y_c_189_n 0.0124478f $X=0.815 $Y=1.765 $X2=0 $Y2=0
cc_52 N_D_c_44_n N_Y_c_189_n 0.00497484f $X=0.83 $Y=1.22 $X2=0 $Y2=0
cc_53 D N_Y_c_189_n 0.027973f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_54 N_D_c_43_n N_Y_c_190_n 0.00101144f $X=0.815 $Y=1.765 $X2=0 $Y2=0
cc_55 N_D_c_44_n N_Y_c_190_n 0.0131907f $X=0.83 $Y=1.22 $X2=0 $Y2=0
cc_56 D N_Y_c_190_n 0.0228656f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_57 N_D_c_43_n N_Y_c_194_n 0.0151942f $X=0.815 $Y=1.765 $X2=0 $Y2=0
cc_58 D N_Y_c_194_n 0.0221856f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_59 N_D_c_43_n N_Y_c_196_n 0.00925663f $X=0.815 $Y=1.765 $X2=0 $Y2=0
cc_60 N_D_c_43_n N_Y_c_199_n 0.0112726f $X=0.815 $Y=1.765 $X2=0 $Y2=0
cc_61 D N_Y_c_199_n 0.00234631f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_62 N_D_c_44_n N_VGND_c_262_n 0.0036777f $X=0.83 $Y=1.22 $X2=0 $Y2=0
cc_63 N_D_c_44_n N_VGND_c_263_n 0.00366857f $X=0.83 $Y=1.22 $X2=0 $Y2=0
cc_64 N_D_c_44_n N_VGND_c_264_n 0.0112037f $X=0.83 $Y=1.22 $X2=0 $Y2=0
cc_65 N_C_c_69_n N_B_c_98_n 0.032462f $X=1.22 $Y=1.22 $X2=-0.19 $Y2=-0.245
cc_66 N_C_c_70_n N_B_c_99_n 0.050956f $X=1.265 $Y=1.765 $X2=0 $Y2=0
cc_67 N_C_c_71_n N_B_c_99_n 4.20537e-19 $X=1.31 $Y=1.385 $X2=0 $Y2=0
cc_68 N_C_c_70_n B 4.18645e-19 $X=1.265 $Y=1.765 $X2=0 $Y2=0
cc_69 N_C_c_71_n B 0.02242f $X=1.31 $Y=1.385 $X2=0 $Y2=0
cc_70 N_C_c_70_n N_VPWR_c_152_n 0.00976006f $X=1.265 $Y=1.765 $X2=0 $Y2=0
cc_71 N_C_c_70_n N_VPWR_c_157_n 0.00445602f $X=1.265 $Y=1.765 $X2=0 $Y2=0
cc_72 N_C_c_70_n N_VPWR_c_150_n 0.00858896f $X=1.265 $Y=1.765 $X2=0 $Y2=0
cc_73 N_C_c_69_n N_Y_c_190_n 0.0122562f $X=1.22 $Y=1.22 $X2=0 $Y2=0
cc_74 N_C_c_70_n N_Y_c_190_n 0.00101661f $X=1.265 $Y=1.765 $X2=0 $Y2=0
cc_75 N_C_c_71_n N_Y_c_190_n 0.0255539f $X=1.31 $Y=1.385 $X2=0 $Y2=0
cc_76 N_C_c_70_n N_Y_c_196_n 0.0112008f $X=1.265 $Y=1.765 $X2=0 $Y2=0
cc_77 N_C_c_70_n N_Y_c_198_n 8.84595e-19 $X=1.265 $Y=1.765 $X2=0 $Y2=0
cc_78 N_C_c_70_n N_Y_c_199_n 0.00572103f $X=1.265 $Y=1.765 $X2=0 $Y2=0
cc_79 N_C_c_71_n N_Y_c_199_n 0.0103162f $X=1.31 $Y=1.385 $X2=0 $Y2=0
cc_80 N_C_c_70_n N_Y_c_200_n 0.0214733f $X=1.265 $Y=1.765 $X2=0 $Y2=0
cc_81 N_C_c_71_n N_Y_c_200_n 0.0146699f $X=1.31 $Y=1.385 $X2=0 $Y2=0
cc_82 N_C_c_69_n N_VGND_c_262_n 0.00461464f $X=1.22 $Y=1.22 $X2=0 $Y2=0
cc_83 N_C_c_69_n N_VGND_c_263_n 0.00465551f $X=1.22 $Y=1.22 $X2=0 $Y2=0
cc_84 N_C_c_69_n N_VGND_c_264_n 0.00180509f $X=1.22 $Y=1.22 $X2=0 $Y2=0
cc_85 N_B_c_98_n N_A_c_129_n 0.029851f $X=1.79 $Y=1.22 $X2=-0.19 $Y2=-0.245
cc_86 B N_A_c_129_n 0.00346899f $X=2.075 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_87 N_B_c_99_n N_A_c_130_n 0.0494262f $X=1.875 $Y=1.765 $X2=0 $Y2=0
cc_88 N_B_c_99_n A 2.22676e-19 $X=1.875 $Y=1.765 $X2=0 $Y2=0
cc_89 B A 0.0306948f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_90 N_B_c_99_n N_VPWR_c_152_n 0.00969525f $X=1.875 $Y=1.765 $X2=0 $Y2=0
cc_91 N_B_c_99_n N_VPWR_c_154_n 8.29197e-19 $X=1.875 $Y=1.765 $X2=0 $Y2=0
cc_92 N_B_c_99_n N_VPWR_c_159_n 0.00445602f $X=1.875 $Y=1.765 $X2=0 $Y2=0
cc_93 N_B_c_99_n N_VPWR_c_150_n 0.0085955f $X=1.875 $Y=1.765 $X2=0 $Y2=0
cc_94 N_B_c_98_n N_Y_c_190_n 0.013201f $X=1.79 $Y=1.22 $X2=0 $Y2=0
cc_95 N_B_c_99_n N_Y_c_190_n 0.0010133f $X=1.875 $Y=1.765 $X2=0 $Y2=0
cc_96 B N_Y_c_190_n 0.0392923f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_97 N_B_c_99_n N_Y_c_196_n 8.78223e-19 $X=1.875 $Y=1.765 $X2=0 $Y2=0
cc_98 N_B_c_99_n N_Y_c_197_n 0.00318394f $X=1.875 $Y=1.765 $X2=0 $Y2=0
cc_99 B N_Y_c_197_n 0.020755f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_100 N_B_c_99_n N_Y_c_198_n 0.0113478f $X=1.875 $Y=1.765 $X2=0 $Y2=0
cc_101 N_B_c_98_n N_Y_c_192_n 0.00223389f $X=1.79 $Y=1.22 $X2=0 $Y2=0
cc_102 N_B_c_99_n N_Y_c_199_n 4.34855e-19 $X=1.875 $Y=1.765 $X2=0 $Y2=0
cc_103 N_B_c_99_n N_Y_c_200_n 0.0206771f $X=1.875 $Y=1.765 $X2=0 $Y2=0
cc_104 B N_Y_c_200_n 0.0118424f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_105 N_B_c_98_n N_VGND_c_262_n 0.00461464f $X=1.79 $Y=1.22 $X2=0 $Y2=0
cc_106 N_B_c_98_n N_VGND_c_263_n 0.00467093f $X=1.79 $Y=1.22 $X2=0 $Y2=0
cc_107 N_A_c_130_n N_VPWR_c_154_n 0.0206403f $X=2.375 $Y=1.765 $X2=0 $Y2=0
cc_108 A N_VPWR_c_154_n 0.0191865f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_109 N_A_c_130_n N_VPWR_c_159_n 0.00413917f $X=2.375 $Y=1.765 $X2=0 $Y2=0
cc_110 N_A_c_130_n N_VPWR_c_150_n 0.00818241f $X=2.375 $Y=1.765 $X2=0 $Y2=0
cc_111 N_A_c_129_n N_Y_c_190_n 0.0145395f $X=2.36 $Y=1.22 $X2=0 $Y2=0
cc_112 N_A_c_130_n N_Y_c_190_n 0.00194404f $X=2.375 $Y=1.765 $X2=0 $Y2=0
cc_113 A N_Y_c_190_n 0.0237695f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_114 N_A_c_130_n N_Y_c_197_n 0.00183618f $X=2.375 $Y=1.765 $X2=0 $Y2=0
cc_115 N_A_c_130_n N_Y_c_198_n 0.00448083f $X=2.375 $Y=1.765 $X2=0 $Y2=0
cc_116 N_A_c_129_n N_Y_c_192_n 0.0109821f $X=2.36 $Y=1.22 $X2=0 $Y2=0
cc_117 N_A_c_129_n N_VGND_c_262_n 0.00434272f $X=2.36 $Y=1.22 $X2=0 $Y2=0
cc_118 N_A_c_129_n N_VGND_c_263_n 0.0045104f $X=2.36 $Y=1.22 $X2=0 $Y2=0
cc_119 N_VPWR_M1003_s N_Y_c_194_n 0.00332155f $X=0.395 $Y=1.84 $X2=0 $Y2=0
cc_120 N_VPWR_c_151_n N_Y_c_194_n 0.0225812f $X=0.54 $Y=2.145 $X2=0 $Y2=0
cc_121 N_VPWR_c_151_n N_Y_c_195_n 0.00268187f $X=0.54 $Y=2.145 $X2=0 $Y2=0
cc_122 N_VPWR_c_151_n N_Y_c_196_n 0.0318965f $X=0.54 $Y=2.145 $X2=0 $Y2=0
cc_123 N_VPWR_c_152_n N_Y_c_196_n 0.0461248f $X=1.565 $Y=2.405 $X2=0 $Y2=0
cc_124 N_VPWR_c_157_n N_Y_c_196_n 0.014552f $X=1.4 $Y=3.33 $X2=0 $Y2=0
cc_125 N_VPWR_c_150_n N_Y_c_196_n 0.0119791f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_126 N_VPWR_c_154_n N_Y_c_197_n 0.0133269f $X=2.6 $Y=1.985 $X2=0 $Y2=0
cc_127 N_VPWR_c_152_n N_Y_c_198_n 0.0443902f $X=1.565 $Y=2.405 $X2=0 $Y2=0
cc_128 N_VPWR_c_154_n N_Y_c_198_n 0.0319341f $X=2.6 $Y=1.985 $X2=0 $Y2=0
cc_129 N_VPWR_c_159_n N_Y_c_198_n 0.0145938f $X=2.435 $Y=3.33 $X2=0 $Y2=0
cc_130 N_VPWR_c_150_n N_Y_c_198_n 0.0120466f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_131 N_VPWR_M1005_d N_Y_c_200_n 0.00584768f $X=1.34 $Y=1.84 $X2=0 $Y2=0
cc_132 N_VPWR_c_152_n N_Y_c_200_n 0.0279337f $X=1.565 $Y=2.405 $X2=0 $Y2=0
cc_133 N_Y_c_190_n N_VGND_M1000_s 0.00674372f $X=2.41 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_134 N_Y_c_192_n N_VGND_c_262_n 0.0145323f $X=2.575 $Y=0.515 $X2=0 $Y2=0
cc_135 N_Y_c_190_n N_VGND_c_263_n 0.0536444f $X=2.41 $Y=0.925 $X2=0 $Y2=0
cc_136 N_Y_c_191_n N_VGND_c_263_n 7.38843e-19 $X=0.405 $Y=0.925 $X2=0 $Y2=0
cc_137 N_Y_c_192_n N_VGND_c_263_n 0.0119861f $X=2.575 $Y=0.515 $X2=0 $Y2=0
cc_138 N_Y_c_190_n N_VGND_c_264_n 0.0192102f $X=2.41 $Y=0.925 $X2=0 $Y2=0
cc_139 N_Y_c_191_n N_VGND_c_264_n 0.0114495f $X=0.405 $Y=0.925 $X2=0 $Y2=0
cc_140 N_Y_c_190_n A_181_74# 0.00722635f $X=2.41 $Y=0.925 $X2=-0.19 $Y2=-0.245
cc_141 N_Y_c_190_n A_259_74# 0.0147367f $X=2.41 $Y=0.925 $X2=-0.19 $Y2=-0.245
cc_142 N_Y_c_190_n A_373_74# 0.00970428f $X=2.41 $Y=0.925 $X2=-0.19 $Y2=-0.245
