* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__clkinv_4 A VGND VNB VPB VPWR Y
M1000 VPWR A Y VPB phighvt w=1.12e+06u l=150000u
+  ad=1.4448e+12p pd=1.154e+07u as=1.008e+12p ps=8.52e+06u
M1001 Y A VGND VNB nshort w=420000u l=150000u
+  ad=4.242e+11p pd=3.7e+06u as=6.216e+11p ps=5.48e+06u
M1002 Y A VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPWR A Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND A Y VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y A VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR A Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND A Y VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y A VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y A VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
