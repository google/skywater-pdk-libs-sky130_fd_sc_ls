# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_ls__o22ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_ls__o22ai_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.160000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.540000 1.320000 1.550000 1.650000 ;
        RECT 1.380000 1.650000 1.550000 1.720000 ;
        RECT 1.380000 1.720000 3.810000 1.890000 ;
        RECT 2.525000 1.890000 3.235000 2.150000 ;
        RECT 3.640000 1.350000 3.970000 1.680000 ;
        RECT 3.640000 1.680000 3.810000 1.720000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.885000 1.180000 3.235000 1.550000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.290000 1.300000 5.635000 1.630000 ;
        RECT 5.405000 1.090000 7.730000 1.260000 ;
        RECT 5.405000 1.260000 5.635000 1.300000 ;
        RECT 7.400000 1.260000 7.730000 1.550000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.805000 1.430000 7.155000 1.680000 ;
        RECT 6.365000 1.680000 7.155000 1.780000 ;
    END
  END B2
  PIN VNB
    PORT
      LAYER pwell ;
        RECT 0.000000 0.000000 8.160000 0.245000 ;
    END
  END VNB
  PIN VPB
    PORT
      LAYER nwell ;
        RECT -0.190000 1.660000 8.350000 3.520000 ;
    END
  END VPB
  PIN Y
    ANTENNADIFFAREA  2.388000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.020000 2.060000 2.350000 2.320000 ;
        RECT 2.020000 2.320000 4.150000 2.490000 ;
        RECT 3.980000 1.850000 6.100000 1.950000 ;
        RECT 3.980000 1.950000 8.070000 2.020000 ;
        RECT 3.980000 2.020000 4.150000 2.320000 ;
        RECT 4.405000 0.750000 8.070000 0.920000 ;
        RECT 4.405000 0.920000 5.155000 1.130000 ;
        RECT 5.770000 2.020000 8.070000 2.120000 ;
        RECT 5.770000 2.120000 6.100000 2.735000 ;
        RECT 6.205000 0.595000 6.535000 0.750000 ;
        RECT 6.670000 2.120000 7.000000 2.735000 ;
        RECT 7.205000 0.595000 7.535000 0.750000 ;
        RECT 7.900000 0.920000 8.070000 1.950000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.160000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.160000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.160000 0.085000 ;
      RECT 0.000000  3.245000 8.160000 3.415000 ;
      RECT 0.115000  0.350000 0.445000 0.980000 ;
      RECT 0.115000  0.980000 4.235000 1.010000 ;
      RECT 0.115000  1.010000 1.375000 1.150000 ;
      RECT 0.120000  1.820000 0.370000 3.245000 ;
      RECT 0.570000  1.820000 0.900000 2.060000 ;
      RECT 0.570000  2.060000 1.850000 2.230000 ;
      RECT 0.570000  2.230000 0.850000 2.980000 ;
      RECT 0.615000  0.085000 0.945000 0.810000 ;
      RECT 1.020000  2.400000 1.350000 3.245000 ;
      RECT 1.125000  0.350000 1.375000 0.840000 ;
      RECT 1.125000  0.840000 4.235000 0.980000 ;
      RECT 1.520000  2.230000 1.850000 2.660000 ;
      RECT 1.520000  2.660000 3.700000 2.980000 ;
      RECT 1.545000  0.085000 1.875000 0.670000 ;
      RECT 2.055000  0.350000 2.305000 0.840000 ;
      RECT 2.475000  0.085000 2.805000 0.670000 ;
      RECT 2.985000  0.350000 3.235000 0.840000 ;
      RECT 3.405000  0.085000 3.735000 0.670000 ;
      RECT 3.870000  2.660000 4.200000 3.245000 ;
      RECT 3.905000  0.255000 8.045000 0.425000 ;
      RECT 3.905000  0.425000 6.035000 0.580000 ;
      RECT 3.905000  0.580000 4.235000 0.840000 ;
      RECT 3.905000  1.010000 4.235000 1.130000 ;
      RECT 4.370000  2.190000 5.570000 2.360000 ;
      RECT 4.370000  2.360000 4.700000 2.980000 ;
      RECT 4.900000  2.530000 5.150000 3.245000 ;
      RECT 5.320000  2.360000 5.570000 2.905000 ;
      RECT 5.320000  2.905000 7.500000 3.075000 ;
      RECT 6.300000  2.290000 6.470000 2.905000 ;
      RECT 6.705000  0.425000 7.035000 0.580000 ;
      RECT 7.170000  2.290000 7.500000 2.905000 ;
      RECT 7.670000  2.290000 8.000000 3.245000 ;
      RECT 7.715000  0.425000 8.045000 0.580000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
  END
END sky130_fd_sc_ls__o22ai_4
END LIBRARY
