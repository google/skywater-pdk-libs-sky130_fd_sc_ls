* File: sky130_fd_sc_ls__a311oi_4.pex.spice
* Created: Wed Sep  2 10:52:02 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__A311OI_4%A3 1 3 6 8 10 13 17 19 21 24 26 28 29 30 31
+ 46 47
c76 47 0 1.91457e-19 $X=1.82 $Y=1.557
c77 46 0 1.16815e-20 $X=1.71 $Y=1.515
c78 26 0 9.70031e-20 $X=1.845 $Y=1.765
r79 47 48 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=1.82 $Y=1.557
+ $X2=1.845 $Y2=1.557
r80 45 47 14.3297 $w=3.7e-07 $l=1.1e-07 $layer=POLY_cond $X=1.71 $Y=1.557
+ $X2=1.82 $Y2=1.557
r81 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.71
+ $Y=1.515 $X2=1.71 $Y2=1.515
r82 43 45 41.0351 $w=3.7e-07 $l=3.15e-07 $layer=POLY_cond $X=1.395 $Y=1.557
+ $X2=1.71 $Y2=1.557
r83 42 43 0.651351 $w=3.7e-07 $l=5e-09 $layer=POLY_cond $X=1.39 $Y=1.557
+ $X2=1.395 $Y2=1.557
r84 41 42 56.0162 $w=3.7e-07 $l=4.3e-07 $layer=POLY_cond $X=0.96 $Y=1.557
+ $X2=1.39 $Y2=1.557
r85 40 41 1.95405 $w=3.7e-07 $l=1.5e-08 $layer=POLY_cond $X=0.945 $Y=1.557
+ $X2=0.96 $Y2=1.557
r86 38 40 33.2189 $w=3.7e-07 $l=2.55e-07 $layer=POLY_cond $X=0.69 $Y=1.557
+ $X2=0.945 $Y2=1.557
r87 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.69
+ $Y=1.515 $X2=0.69 $Y2=1.515
r88 36 38 20.8432 $w=3.7e-07 $l=1.6e-07 $layer=POLY_cond $X=0.53 $Y=1.557
+ $X2=0.69 $Y2=1.557
r89 35 36 4.55946 $w=3.7e-07 $l=3.5e-08 $layer=POLY_cond $X=0.495 $Y=1.557
+ $X2=0.53 $Y2=1.557
r90 31 46 0.80403 $w=4.28e-07 $l=3e-08 $layer=LI1_cond $X=1.68 $Y=1.565 $X2=1.71
+ $Y2=1.565
r91 30 31 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.565
+ $X2=1.68 $Y2=1.565
r92 29 30 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=1.2 $Y2=1.565
r93 29 39 0.80403 $w=4.28e-07 $l=3e-08 $layer=LI1_cond $X=0.72 $Y=1.565 $X2=0.69
+ $Y2=1.565
r94 26 48 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.845 $Y=1.765
+ $X2=1.845 $Y2=1.557
r95 26 28 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.845 $Y=1.765
+ $X2=1.845 $Y2=2.4
r96 22 47 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.82 $Y=1.35
+ $X2=1.82 $Y2=1.557
r97 22 24 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.82 $Y=1.35
+ $X2=1.82 $Y2=0.74
r98 19 43 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.395 $Y=1.765
+ $X2=1.395 $Y2=1.557
r99 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.395 $Y=1.765
+ $X2=1.395 $Y2=2.4
r100 15 42 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.39 $Y=1.35
+ $X2=1.39 $Y2=1.557
r101 15 17 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.39 $Y=1.35
+ $X2=1.39 $Y2=0.74
r102 11 41 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.96 $Y=1.35
+ $X2=0.96 $Y2=1.557
r103 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.96 $Y=1.35
+ $X2=0.96 $Y2=0.74
r104 8 40 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.945 $Y=1.765
+ $X2=0.945 $Y2=1.557
r105 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.945 $Y=1.765
+ $X2=0.945 $Y2=2.4
r106 4 36 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.53 $Y=1.35
+ $X2=0.53 $Y2=1.557
r107 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.53 $Y=1.35 $X2=0.53
+ $Y2=0.74
r108 1 35 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.495 $Y=1.765
+ $X2=0.495 $Y2=1.557
r109 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.495 $Y=1.765
+ $X2=0.495 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__A311OI_4%A2 3 5 7 10 12 14 17 19 21 24 26 28 29 30
+ 31 32 49
c84 49 0 3.84326e-19 $X=3.54 $Y=1.557
c85 32 0 1.75706e-19 $X=3.6 $Y=1.665
c86 5 0 1.16815e-20 $X=2.295 $Y=1.765
r87 49 50 13.8658 $w=3.65e-07 $l=1.05e-07 $layer=POLY_cond $X=3.54 $Y=1.557
+ $X2=3.645 $Y2=1.557
r88 47 49 19.8082 $w=3.65e-07 $l=1.5e-07 $layer=POLY_cond $X=3.39 $Y=1.557
+ $X2=3.54 $Y2=1.557
r89 47 48 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.39
+ $Y=1.515 $X2=3.39 $Y2=1.515
r90 45 47 25.7507 $w=3.65e-07 $l=1.95e-07 $layer=POLY_cond $X=3.195 $Y=1.557
+ $X2=3.39 $Y2=1.557
r91 44 45 11.2247 $w=3.65e-07 $l=8.5e-08 $layer=POLY_cond $X=3.11 $Y=1.557
+ $X2=3.195 $Y2=1.557
r92 43 44 48.2 $w=3.65e-07 $l=3.65e-07 $layer=POLY_cond $X=2.745 $Y=1.557
+ $X2=3.11 $Y2=1.557
r93 42 43 8.58356 $w=3.65e-07 $l=6.5e-08 $layer=POLY_cond $X=2.68 $Y=1.557
+ $X2=2.745 $Y2=1.557
r94 40 42 40.937 $w=3.65e-07 $l=3.1e-07 $layer=POLY_cond $X=2.37 $Y=1.557
+ $X2=2.68 $Y2=1.557
r95 40 41 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.37
+ $Y=1.515 $X2=2.37 $Y2=1.515
r96 38 40 9.90411 $w=3.65e-07 $l=7.5e-08 $layer=POLY_cond $X=2.295 $Y=1.557
+ $X2=2.37 $Y2=1.557
r97 37 38 5.94247 $w=3.65e-07 $l=4.5e-08 $layer=POLY_cond $X=2.25 $Y=1.557
+ $X2=2.295 $Y2=1.557
r98 32 48 5.62821 $w=4.28e-07 $l=2.1e-07 $layer=LI1_cond $X=3.6 $Y=1.565
+ $X2=3.39 $Y2=1.565
r99 31 48 7.23627 $w=4.28e-07 $l=2.7e-07 $layer=LI1_cond $X=3.12 $Y=1.565
+ $X2=3.39 $Y2=1.565
r100 30 31 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=2.64 $Y=1.565
+ $X2=3.12 $Y2=1.565
r101 30 41 7.23627 $w=4.28e-07 $l=2.7e-07 $layer=LI1_cond $X=2.64 $Y=1.565
+ $X2=2.37 $Y2=1.565
r102 29 41 5.62821 $w=4.28e-07 $l=2.1e-07 $layer=LI1_cond $X=2.16 $Y=1.565
+ $X2=2.37 $Y2=1.565
r103 26 50 23.6381 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.645 $Y=1.765
+ $X2=3.645 $Y2=1.557
r104 26 28 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.645 $Y=1.765
+ $X2=3.645 $Y2=2.4
r105 22 49 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.54 $Y=1.35
+ $X2=3.54 $Y2=1.557
r106 22 24 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.54 $Y=1.35
+ $X2=3.54 $Y2=0.74
r107 19 45 23.6381 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.195 $Y=1.765
+ $X2=3.195 $Y2=1.557
r108 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.195 $Y=1.765
+ $X2=3.195 $Y2=2.4
r109 15 44 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.11 $Y=1.35
+ $X2=3.11 $Y2=1.557
r110 15 17 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.11 $Y=1.35
+ $X2=3.11 $Y2=0.74
r111 12 43 23.6381 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.745 $Y=1.765
+ $X2=2.745 $Y2=1.557
r112 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.745 $Y=1.765
+ $X2=2.745 $Y2=2.4
r113 8 42 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.68 $Y=1.35
+ $X2=2.68 $Y2=1.557
r114 8 10 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.68 $Y=1.35
+ $X2=2.68 $Y2=0.74
r115 5 38 23.6381 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.295 $Y=1.765
+ $X2=2.295 $Y2=1.557
r116 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.295 $Y=1.765
+ $X2=2.295 $Y2=2.4
r117 1 37 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.25 $Y=1.35
+ $X2=2.25 $Y2=1.557
r118 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.25 $Y=1.35 $X2=2.25
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__A311OI_4%A1 1 3 4 6 8 11 13 15 18 20 22 25 29 31 33
+ 34 47
c85 47 0 1.98771e-19 $X=5.91 $Y=1.515
c86 29 0 8.65694e-20 $X=6 $Y=0.74
c87 1 0 7.87025e-20 $X=4.095 $Y=1.765
r88 47 49 12.8343 $w=3.38e-07 $l=9e-08 $layer=POLY_cond $X=5.91 $Y=1.557 $X2=6
+ $Y2=1.557
r89 47 48 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.91
+ $Y=1.515 $X2=5.91 $Y2=1.515
r90 45 47 48.4852 $w=3.38e-07 $l=3.4e-07 $layer=POLY_cond $X=5.57 $Y=1.557
+ $X2=5.91 $Y2=1.557
r91 44 45 17.8254 $w=3.38e-07 $l=1.25e-07 $layer=POLY_cond $X=5.445 $Y=1.557
+ $X2=5.57 $Y2=1.557
r92 42 44 34.9379 $w=3.38e-07 $l=2.45e-07 $layer=POLY_cond $X=5.2 $Y=1.557
+ $X2=5.445 $Y2=1.557
r93 42 43 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.2
+ $Y=1.515 $X2=5.2 $Y2=1.515
r94 40 42 8.55621 $w=3.38e-07 $l=6e-08 $layer=POLY_cond $X=5.14 $Y=1.557 $X2=5.2
+ $Y2=1.557
r95 39 40 20.6775 $w=3.38e-07 $l=1.45e-07 $layer=POLY_cond $X=4.995 $Y=1.557
+ $X2=5.14 $Y2=1.557
r96 38 39 40.642 $w=3.38e-07 $l=2.85e-07 $layer=POLY_cond $X=4.71 $Y=1.557
+ $X2=4.995 $Y2=1.557
r97 37 38 23.5296 $w=3.38e-07 $l=1.65e-07 $layer=POLY_cond $X=4.545 $Y=1.557
+ $X2=4.71 $Y2=1.557
r98 34 48 2.41209 $w=4.28e-07 $l=9e-08 $layer=LI1_cond $X=6 $Y=1.565 $X2=5.91
+ $Y2=1.565
r99 33 48 10.4524 $w=4.28e-07 $l=3.9e-07 $layer=LI1_cond $X=5.52 $Y=1.565
+ $X2=5.91 $Y2=1.565
r100 33 43 8.57632 $w=4.28e-07 $l=3.2e-07 $layer=LI1_cond $X=5.52 $Y=1.565
+ $X2=5.2 $Y2=1.565
r101 27 49 21.7938 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6 $Y=1.35 $X2=6
+ $Y2=1.557
r102 27 29 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6 $Y=1.35 $X2=6
+ $Y2=0.74
r103 23 45 21.7938 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.57 $Y=1.35
+ $X2=5.57 $Y2=1.557
r104 23 25 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.57 $Y=1.35
+ $X2=5.57 $Y2=0.74
r105 20 44 21.7938 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=5.445 $Y=1.765
+ $X2=5.445 $Y2=1.557
r106 20 22 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.445 $Y=1.765
+ $X2=5.445 $Y2=2.4
r107 16 40 21.7938 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.14 $Y=1.35
+ $X2=5.14 $Y2=1.557
r108 16 18 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.14 $Y=1.35
+ $X2=5.14 $Y2=0.74
r109 13 39 21.7938 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=4.995 $Y=1.765
+ $X2=4.995 $Y2=1.557
r110 13 15 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.995 $Y=1.765
+ $X2=4.995 $Y2=2.4
r111 9 38 21.7938 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.71 $Y=1.35
+ $X2=4.71 $Y2=1.557
r112 9 11 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.71 $Y=1.35
+ $X2=4.71 $Y2=0.74
r113 6 37 21.7938 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=4.545 $Y=1.765
+ $X2=4.545 $Y2=1.557
r114 6 8 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.545 $Y=1.765
+ $X2=4.545 $Y2=2.4
r115 5 31 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.185 $Y=1.605
+ $X2=4.095 $Y2=1.605
r116 4 37 27.9663 $w=3.38e-07 $l=1.11445e-07 $layer=POLY_cond $X=4.455 $Y=1.605
+ $X2=4.545 $Y2=1.557
r117 4 5 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=4.455 $Y=1.605
+ $X2=4.185 $Y2=1.605
r118 1 31 64.3434 $w=1.8e-07 $l=1.6e-07 $layer=POLY_cond $X=4.095 $Y=1.765
+ $X2=4.095 $Y2=1.605
r119 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.095 $Y=1.765
+ $X2=4.095 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__A311OI_4%B1 1 3 6 8 10 11 13 16 18 20 21 22 35 37
c77 37 0 2.85341e-19 $X=7.32 $Y=1.415
c78 18 0 1.69938e-19 $X=7.765 $Y=1.765
c79 6 0 1.0484e-19 $X=6.43 $Y=0.74
r80 35 36 7.06933 $w=3.75e-07 $l=5.5e-08 $layer=POLY_cond $X=7.71 $Y=1.542
+ $X2=7.765 $Y2=1.542
r81 33 35 11.568 $w=3.75e-07 $l=9e-08 $layer=POLY_cond $X=7.62 $Y=1.542 $X2=7.71
+ $Y2=1.542
r82 33 34 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=7.62
+ $Y=1.485 $X2=7.62 $Y2=1.485
r83 31 33 39.2027 $w=3.75e-07 $l=3.05e-07 $layer=POLY_cond $X=7.315 $Y=1.542
+ $X2=7.62 $Y2=1.542
r84 29 31 48.2 $w=3.75e-07 $l=3.75e-07 $layer=POLY_cond $X=6.94 $Y=1.542
+ $X2=7.315 $Y2=1.542
r85 29 30 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=6.94
+ $Y=1.485 $X2=6.94 $Y2=1.485
r86 27 29 9.64 $w=3.75e-07 $l=7.5e-08 $layer=POLY_cond $X=6.865 $Y=1.542
+ $X2=6.94 $Y2=1.542
r87 26 27 55.912 $w=3.75e-07 $l=4.35e-07 $layer=POLY_cond $X=6.43 $Y=1.542
+ $X2=6.865 $Y2=1.542
r88 25 26 1.928 $w=3.75e-07 $l=1.5e-08 $layer=POLY_cond $X=6.415 $Y=1.542
+ $X2=6.43 $Y2=1.542
r89 22 34 5.49 $w=4e-07 $l=1.8e-07 $layer=LI1_cond $X=7.44 $Y=1.415 $X2=7.62
+ $Y2=1.415
r90 22 37 3.4204 $w=4.7e-07 $l=1.2e-07 $layer=LI1_cond $X=7.44 $Y=1.415 $X2=7.32
+ $Y2=1.415
r91 21 37 9.16145 $w=4.68e-07 $l=3.6e-07 $layer=LI1_cond $X=6.96 $Y=1.415
+ $X2=7.32 $Y2=1.415
r92 21 30 0.50897 $w=4.68e-07 $l=2e-08 $layer=LI1_cond $X=6.96 $Y=1.415 $X2=6.94
+ $Y2=1.415
r93 18 36 24.2915 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=7.765 $Y=1.765
+ $X2=7.765 $Y2=1.542
r94 18 20 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.765 $Y=1.765
+ $X2=7.765 $Y2=2.4
r95 14 35 24.2915 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=7.71 $Y=1.32
+ $X2=7.71 $Y2=1.542
r96 14 16 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=7.71 $Y=1.32
+ $X2=7.71 $Y2=0.74
r97 11 31 24.2915 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=7.315 $Y=1.765
+ $X2=7.315 $Y2=1.542
r98 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.315 $Y=1.765
+ $X2=7.315 $Y2=2.4
r99 8 27 24.2915 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=6.865 $Y=1.765
+ $X2=6.865 $Y2=1.542
r100 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.865 $Y=1.765
+ $X2=6.865 $Y2=2.4
r101 4 26 24.2915 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=6.43 $Y=1.32
+ $X2=6.43 $Y2=1.542
r102 4 6 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.43 $Y=1.32 $X2=6.43
+ $Y2=0.74
r103 1 25 24.2915 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=6.415 $Y=1.765
+ $X2=6.415 $Y2=1.542
r104 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.415 $Y=1.765
+ $X2=6.415 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__A311OI_4%C1 1 3 4 6 7 9 10 12 13 15 16 17 19 20 22
+ 23 24 36 38 47
c78 1 0 1.44963e-19 $X=8.14 $Y=1.22
r79 38 47 2.36628 $w=3.7e-07 $l=7e-08 $layer=LI1_cond $X=8.47 $Y=1.365 $X2=8.4
+ $Y2=1.365
r80 35 37 22.9258 $w=4.31e-07 $l=2.05e-07 $layer=POLY_cond $X=8.91 $Y=1.492
+ $X2=9.115 $Y2=1.492
r81 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.91
+ $Y=1.385 $X2=8.91 $Y2=1.385
r82 33 35 27.3991 $w=4.31e-07 $l=2.45e-07 $layer=POLY_cond $X=8.665 $Y=1.492
+ $X2=8.91 $Y2=1.492
r83 31 33 10.6241 $w=4.31e-07 $l=9.5e-08 $layer=POLY_cond $X=8.57 $Y=1.492
+ $X2=8.665 $Y2=1.492
r84 31 32 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.57
+ $Y=1.385 $X2=8.57 $Y2=1.385
r85 29 31 39.7007 $w=4.31e-07 $l=3.55e-07 $layer=POLY_cond $X=8.215 $Y=1.492
+ $X2=8.57 $Y2=1.492
r86 28 29 8.38747 $w=4.31e-07 $l=7.5e-08 $layer=POLY_cond $X=8.14 $Y=1.492
+ $X2=8.215 $Y2=1.492
r87 24 36 0.934413 $w=3.68e-07 $l=3e-08 $layer=LI1_cond $X=8.88 $Y=1.365
+ $X2=8.91 $Y2=1.365
r88 24 32 9.6556 $w=3.68e-07 $l=3.1e-07 $layer=LI1_cond $X=8.88 $Y=1.365
+ $X2=8.57 $Y2=1.365
r89 23 47 0.28046 $w=3.48e-07 $l=8e-09 $layer=LI1_cond $X=8.392 $Y=1.365 $X2=8.4
+ $Y2=1.365
r90 23 32 2.89668 $w=3.68e-07 $l=9.3e-08 $layer=LI1_cond $X=8.477 $Y=1.365
+ $X2=8.57 $Y2=1.365
r91 23 38 0.21803 $w=3.68e-07 $l=7e-09 $layer=LI1_cond $X=8.477 $Y=1.365
+ $X2=8.47 $Y2=1.365
r92 20 22 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=9.565 $Y=1.765
+ $X2=9.565 $Y2=2.4
r93 19 20 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=9.565 $Y=1.675
+ $X2=9.565 $Y2=1.765
r94 18 19 79.6855 $w=1.8e-07 $l=2.05e-07 $layer=POLY_cond $X=9.565 $Y=1.47
+ $X2=9.565 $Y2=1.675
r95 17 37 18.4942 $w=4.31e-07 $l=1.86652e-07 $layer=POLY_cond $X=9.205 $Y=1.345
+ $X2=9.115 $Y2=1.492
r96 16 18 27.8695 $w=2.5e-07 $l=1.63936e-07 $layer=POLY_cond $X=9.475 $Y=1.345
+ $X2=9.565 $Y2=1.47
r97 16 17 67.0825 $w=2.5e-07 $l=2.7e-07 $layer=POLY_cond $X=9.475 $Y=1.345
+ $X2=9.205 $Y2=1.345
r98 13 37 27.6969 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=9.115 $Y=1.765
+ $X2=9.115 $Y2=1.492
r99 13 15 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=9.115 $Y=1.765
+ $X2=9.115 $Y2=2.4
r100 10 33 27.6969 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=8.665 $Y=1.765
+ $X2=8.665 $Y2=1.492
r101 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.665 $Y=1.765
+ $X2=8.665 $Y2=2.4
r102 7 31 27.6969 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=8.57 $Y=1.22
+ $X2=8.57 $Y2=1.492
r103 7 9 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=8.57 $Y=1.22 $X2=8.57
+ $Y2=0.74
r104 4 29 27.6969 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=8.215 $Y=1.765
+ $X2=8.215 $Y2=1.492
r105 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.215 $Y=1.765
+ $X2=8.215 $Y2=2.4
r106 1 28 27.6969 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=8.14 $Y=1.22
+ $X2=8.14 $Y2=1.492
r107 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=8.14 $Y=1.22 $X2=8.14
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__A311OI_4%VPWR 1 2 3 4 5 6 7 22 24 30 34 38 42 46 48
+ 52 55 56 58 59 61 62 63 64 65 67 90 91 97 100
r142 100 101 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r143 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r144 94 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r145 90 91 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r146 88 91 1.07034 $w=4.9e-07 $l=3.84e-06 $layer=MET1_cond $X=6 $Y=3.33 $X2=9.84
+ $Y2=3.33
r147 88 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=5.52 $Y2=3.33
r148 87 90 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=6 $Y=3.33 $X2=9.84
+ $Y2=3.33
r149 87 88 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=6 $Y=3.33
+ $X2=6 $Y2=3.33
r150 85 100 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.835 $Y=3.33
+ $X2=5.67 $Y2=3.33
r151 85 87 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=5.835 $Y=3.33
+ $X2=6 $Y2=3.33
r152 83 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r153 81 84 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r154 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r155 78 81 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r156 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r157 75 78 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r158 75 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r159 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r160 72 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.335 $Y=3.33
+ $X2=1.17 $Y2=3.33
r161 72 74 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.335 $Y=3.33
+ $X2=1.68 $Y2=3.33
r162 71 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r163 71 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r164 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r165 68 94 4.02368 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=0.355 $Y=3.33
+ $X2=0.177 $Y2=3.33
r166 68 70 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.355 $Y=3.33
+ $X2=0.72 $Y2=3.33
r167 67 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.005 $Y=3.33
+ $X2=1.17 $Y2=3.33
r168 67 70 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.005 $Y=3.33
+ $X2=0.72 $Y2=3.33
r169 65 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r170 65 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r171 63 83 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=4.605 $Y=3.33
+ $X2=4.56 $Y2=3.33
r172 63 64 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.605 $Y=3.33
+ $X2=4.73 $Y2=3.33
r173 61 80 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=3.705 $Y=3.33
+ $X2=3.6 $Y2=3.33
r174 61 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.705 $Y=3.33
+ $X2=3.87 $Y2=3.33
r175 60 83 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=4.035 $Y=3.33
+ $X2=4.56 $Y2=3.33
r176 60 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.035 $Y=3.33
+ $X2=3.87 $Y2=3.33
r177 58 77 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.805 $Y=3.33
+ $X2=2.64 $Y2=3.33
r178 58 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.805 $Y=3.33
+ $X2=2.97 $Y2=3.33
r179 57 80 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=3.135 $Y=3.33
+ $X2=3.6 $Y2=3.33
r180 57 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.135 $Y=3.33
+ $X2=2.97 $Y2=3.33
r181 55 74 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=1.905 $Y=3.33
+ $X2=1.68 $Y2=3.33
r182 55 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.905 $Y=3.33
+ $X2=2.07 $Y2=3.33
r183 54 77 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=2.235 $Y=3.33
+ $X2=2.64 $Y2=3.33
r184 54 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.235 $Y=3.33
+ $X2=2.07 $Y2=3.33
r185 50 100 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.67 $Y=3.245
+ $X2=5.67 $Y2=3.33
r186 50 52 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=5.67 $Y=3.245
+ $X2=5.67 $Y2=2.455
r187 49 64 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.855 $Y=3.33
+ $X2=4.73 $Y2=3.33
r188 48 100 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.505 $Y=3.33
+ $X2=5.67 $Y2=3.33
r189 48 49 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=5.505 $Y=3.33
+ $X2=4.855 $Y2=3.33
r190 44 64 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.73 $Y=3.245
+ $X2=4.73 $Y2=3.33
r191 44 46 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=4.73 $Y=3.245
+ $X2=4.73 $Y2=2.455
r192 40 62 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.87 $Y=3.245
+ $X2=3.87 $Y2=3.33
r193 40 42 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=3.87 $Y=3.245
+ $X2=3.87 $Y2=2.455
r194 36 59 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.97 $Y=3.245
+ $X2=2.97 $Y2=3.33
r195 36 38 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=2.97 $Y=3.245
+ $X2=2.97 $Y2=2.455
r196 32 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.07 $Y=3.245
+ $X2=2.07 $Y2=3.33
r197 32 34 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=2.07 $Y=3.245
+ $X2=2.07 $Y2=2.455
r198 28 97 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.17 $Y=3.245
+ $X2=1.17 $Y2=3.33
r199 28 30 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=1.17 $Y=3.245
+ $X2=1.17 $Y2=2.455
r200 24 27 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=0.23 $Y=1.985
+ $X2=0.23 $Y2=2.815
r201 22 94 3.11948 $w=2.5e-07 $l=1.08305e-07 $layer=LI1_cond $X=0.23 $Y=3.245
+ $X2=0.177 $Y2=3.33
r202 22 27 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.23 $Y=3.245
+ $X2=0.23 $Y2=2.815
r203 7 52 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=5.52
+ $Y=1.84 $X2=5.67 $Y2=2.455
r204 6 46 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=4.62
+ $Y=1.84 $X2=4.77 $Y2=2.455
r205 5 42 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=3.72
+ $Y=1.84 $X2=3.87 $Y2=2.455
r206 4 38 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=2.82
+ $Y=1.84 $X2=2.97 $Y2=2.455
r207 3 34 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=1.92
+ $Y=1.84 $X2=2.07 $Y2=2.455
r208 2 30 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=1.02
+ $Y=1.84 $X2=1.17 $Y2=2.455
r209 1 27 400 $w=1.7e-07 $l=1.03562e-06 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.84 $X2=0.27 $Y2=2.815
r210 1 24 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.84 $X2=0.27 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_LS__A311OI_4%A_114_368# 1 2 3 4 5 6 7 8 25 27 29 33 35
+ 39 41 45 47 51 53 57 59 63 65 67 69 74 76 78 80 82 84
c119 67 0 1.69938e-19 $X=7.54 $Y=2.15
c120 47 0 1.91457e-19 $X=4.235 $Y=2.035
c121 35 0 3.84326e-19 $X=2.435 $Y=2.035
r122 67 86 4.18573 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=7.54 $Y=2.15
+ $X2=7.54 $Y2=1.985
r123 67 69 21.0446 $w=2.28e-07 $l=4.2e-07 $layer=LI1_cond $X=7.54 $Y=2.15
+ $X2=7.54 $Y2=2.57
r124 66 84 4.81705 $w=2.5e-07 $l=1.4e-07 $layer=LI1_cond $X=6.755 $Y=1.985
+ $X2=6.615 $Y2=1.985
r125 65 86 2.91733 $w=3.3e-07 $l=1.15e-07 $layer=LI1_cond $X=7.425 $Y=1.985
+ $X2=7.54 $Y2=1.985
r126 65 66 23.3981 $w=3.28e-07 $l=6.7e-07 $layer=LI1_cond $X=7.425 $Y=1.985
+ $X2=6.755 $Y2=1.985
r127 61 84 1.64447 $w=2.3e-07 $l=1.77059e-07 $layer=LI1_cond $X=6.64 $Y=2.15
+ $X2=6.615 $Y2=1.985
r128 61 63 21.0446 $w=2.28e-07 $l=4.2e-07 $layer=LI1_cond $X=6.64 $Y=2.15
+ $X2=6.64 $Y2=2.57
r129 60 82 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.305 $Y=2.035
+ $X2=5.18 $Y2=2.035
r130 59 84 4.81705 $w=2.5e-07 $l=1.63095e-07 $layer=LI1_cond $X=6.475 $Y=2.035
+ $X2=6.615 $Y2=1.985
r131 59 60 76.3316 $w=1.68e-07 $l=1.17e-06 $layer=LI1_cond $X=6.475 $Y=2.035
+ $X2=5.305 $Y2=2.035
r132 55 82 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.18 $Y=2.12
+ $X2=5.18 $Y2=2.035
r133 55 57 32.0379 $w=2.48e-07 $l=6.95e-07 $layer=LI1_cond $X=5.18 $Y=2.12
+ $X2=5.18 $Y2=2.815
r134 54 80 5.16603 $w=1.7e-07 $l=1.12916e-07 $layer=LI1_cond $X=4.405 $Y=2.035
+ $X2=4.32 $Y2=1.97
r135 53 82 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.055 $Y=2.035
+ $X2=5.18 $Y2=2.035
r136 53 54 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=5.055 $Y=2.035
+ $X2=4.405 $Y2=2.035
r137 49 80 1.34256 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=4.32 $Y=2.12
+ $X2=4.32 $Y2=1.97
r138 49 51 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=4.32 $Y=2.12
+ $X2=4.32 $Y2=2.4
r139 48 78 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.505 $Y=2.035
+ $X2=3.42 $Y2=2.035
r140 47 80 5.16603 $w=1.7e-07 $l=1.12916e-07 $layer=LI1_cond $X=4.235 $Y=2.035
+ $X2=4.32 $Y2=1.97
r141 47 48 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=4.235 $Y=2.035
+ $X2=3.505 $Y2=2.035
r142 43 78 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.42 $Y=2.12
+ $X2=3.42 $Y2=2.035
r143 43 45 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=3.42 $Y=2.12
+ $X2=3.42 $Y2=2.815
r144 42 76 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.605 $Y=2.035
+ $X2=2.52 $Y2=2.035
r145 41 78 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.335 $Y=2.035
+ $X2=3.42 $Y2=2.035
r146 41 42 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=3.335 $Y=2.035
+ $X2=2.605 $Y2=2.035
r147 37 76 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.52 $Y=2.12
+ $X2=2.52 $Y2=2.035
r148 37 39 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=2.52 $Y=2.12
+ $X2=2.52 $Y2=2.815
r149 36 74 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.705 $Y=2.035
+ $X2=1.62 $Y2=2.035
r150 35 76 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.435 $Y=2.035
+ $X2=2.52 $Y2=2.035
r151 35 36 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=2.435 $Y=2.035
+ $X2=1.705 $Y2=2.035
r152 31 74 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.62 $Y=2.12
+ $X2=1.62 $Y2=2.035
r153 31 33 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=1.62 $Y=2.12
+ $X2=1.62 $Y2=2.815
r154 30 72 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.805 $Y=2.035
+ $X2=0.68 $Y2=2.035
r155 29 74 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.535 $Y=2.035
+ $X2=1.62 $Y2=2.035
r156 29 30 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.535 $Y=2.035
+ $X2=0.805 $Y2=2.035
r157 25 72 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.12
+ $X2=0.68 $Y2=2.035
r158 25 27 32.0379 $w=2.48e-07 $l=6.95e-07 $layer=LI1_cond $X=0.68 $Y=2.12
+ $X2=0.68 $Y2=2.815
r159 8 86 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=7.39
+ $Y=1.84 $X2=7.54 $Y2=1.985
r160 8 69 600 $w=1.7e-07 $l=8.01499e-07 $layer=licon1_PDIFF $count=1 $X=7.39
+ $Y=1.84 $X2=7.54 $Y2=2.57
r161 7 84 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=6.49
+ $Y=1.84 $X2=6.64 $Y2=1.985
r162 7 63 600 $w=1.7e-07 $l=8.01499e-07 $layer=licon1_PDIFF $count=1 $X=6.49
+ $Y=1.84 $X2=6.64 $Y2=2.57
r163 6 82 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=5.07
+ $Y=1.84 $X2=5.22 $Y2=2.115
r164 6 57 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=5.07
+ $Y=1.84 $X2=5.22 $Y2=2.815
r165 5 80 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=4.17
+ $Y=1.84 $X2=4.32 $Y2=1.985
r166 5 51 300 $w=1.7e-07 $l=6.30555e-07 $layer=licon1_PDIFF $count=2 $X=4.17
+ $Y=1.84 $X2=4.32 $Y2=2.4
r167 4 78 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=3.27
+ $Y=1.84 $X2=3.42 $Y2=2.115
r168 4 45 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=3.27
+ $Y=1.84 $X2=3.42 $Y2=2.815
r169 3 76 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=2.37
+ $Y=1.84 $X2=2.52 $Y2=2.115
r170 3 39 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.37
+ $Y=1.84 $X2=2.52 $Y2=2.815
r171 2 74 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=1.47
+ $Y=1.84 $X2=1.62 $Y2=2.115
r172 2 33 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.47
+ $Y=1.84 $X2=1.62 $Y2=2.815
r173 1 72 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=0.57
+ $Y=1.84 $X2=0.72 $Y2=2.115
r174 1 27 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=0.57
+ $Y=1.84 $X2=0.72 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_LS__A311OI_4%A_1213_368# 1 2 3 4 5 18 20 21 24 26 30 34
+ 38 40 44 48 49 50
r85 44 47 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=9.79 $Y=1.985
+ $X2=9.79 $Y2=2.815
r86 42 47 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=9.79 $Y=2.905 $X2=9.79
+ $Y2=2.815
r87 41 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.055 $Y=2.99
+ $X2=8.89 $Y2=2.99
r88 40 42 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.625 $Y=2.99
+ $X2=9.79 $Y2=2.905
r89 40 41 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=9.625 $Y=2.99
+ $X2=9.055 $Y2=2.99
r90 36 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.89 $Y=2.905
+ $X2=8.89 $Y2=2.99
r91 36 38 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=8.89 $Y=2.905
+ $X2=8.89 $Y2=2.225
r92 35 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.155 $Y=2.99
+ $X2=7.99 $Y2=2.99
r93 34 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.725 $Y=2.99
+ $X2=8.89 $Y2=2.99
r94 34 35 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=8.725 $Y=2.99
+ $X2=8.155 $Y2=2.99
r95 30 33 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=7.99 $Y=1.985
+ $X2=7.99 $Y2=2.815
r96 28 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.99 $Y=2.905
+ $X2=7.99 $Y2=2.99
r97 28 33 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=7.99 $Y=2.905 $X2=7.99
+ $Y2=2.815
r98 27 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.255 $Y=2.99
+ $X2=7.09 $Y2=2.99
r99 26 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.825 $Y=2.99
+ $X2=7.99 $Y2=2.99
r100 26 27 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=7.825 $Y=2.99
+ $X2=7.255 $Y2=2.99
r101 22 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.09 $Y=2.905
+ $X2=7.09 $Y2=2.99
r102 22 24 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=7.09 $Y=2.905
+ $X2=7.09 $Y2=2.405
r103 20 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.925 $Y=2.99
+ $X2=7.09 $Y2=2.99
r104 20 21 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=6.925 $Y=2.99
+ $X2=6.355 $Y2=2.99
r105 16 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.19 $Y=2.905
+ $X2=6.355 $Y2=2.99
r106 16 18 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=6.19 $Y=2.905
+ $X2=6.19 $Y2=2.405
r107 5 47 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=9.64
+ $Y=1.84 $X2=9.79 $Y2=2.815
r108 5 44 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=9.64
+ $Y=1.84 $X2=9.79 $Y2=1.985
r109 4 38 300 $w=1.7e-07 $l=4.53845e-07 $layer=licon1_PDIFF $count=2 $X=8.74
+ $Y=1.84 $X2=8.89 $Y2=2.225
r110 3 33 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=7.84
+ $Y=1.84 $X2=7.99 $Y2=2.815
r111 3 30 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=7.84
+ $Y=1.84 $X2=7.99 $Y2=1.985
r112 2 24 300 $w=1.7e-07 $l=6.3559e-07 $layer=licon1_PDIFF $count=2 $X=6.94
+ $Y=1.84 $X2=7.09 $Y2=2.405
r113 1 18 300 $w=1.7e-07 $l=6.2438e-07 $layer=licon1_PDIFF $count=2 $X=6.065
+ $Y=1.84 $X2=6.19 $Y2=2.405
.ends

.subckt PM_SKY130_FD_SC_LS__A311OI_4%Y 1 2 3 4 5 6 7 22 28 30 34 40 42 43 45 48
+ 53 55 56 57 58 59 60 72 79 80
c99 34 0 1.44963e-19 $X=7.925 $Y=0.515
r100 79 80 4.36053 $w=6.58e-07 $l=6.5e-08 $layer=LI1_cond $X=9.36 $Y=0.68
+ $X2=9.425 $Y2=0.68
r101 71 72 9.09709 $w=6.58e-07 $l=8.5e-08 $layer=LI1_cond $X=8.785 $Y=0.68
+ $X2=8.7 $Y2=0.68
r102 59 79 0.181224 $w=6.58e-07 $l=1e-08 $layer=LI1_cond $X=9.35 $Y=0.68
+ $X2=9.36 $Y2=0.68
r103 59 76 0.181224 $w=6.58e-07 $l=1e-08 $layer=LI1_cond $X=9.35 $Y=0.68
+ $X2=9.34 $Y2=0.68
r104 59 60 14.5856 $w=3.18e-07 $l=4.05e-07 $layer=LI1_cond $X=9.435 $Y=0.51
+ $X2=9.84 $Y2=0.51
r105 59 80 0.360138 $w=3.18e-07 $l=1e-08 $layer=LI1_cond $X=9.435 $Y=0.51
+ $X2=9.425 $Y2=0.51
r106 58 76 8.3363 $w=6.58e-07 $l=4.6e-07 $layer=LI1_cond $X=8.88 $Y=0.68
+ $X2=9.34 $Y2=0.68
r107 58 71 1.72163 $w=6.58e-07 $l=9.5e-08 $layer=LI1_cond $X=8.88 $Y=0.68
+ $X2=8.785 $Y2=0.68
r108 51 53 5.88189 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=4.495 $Y=0.95
+ $X2=4.66 $Y2=0.95
r109 46 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.34 $Y=1.89
+ $X2=9.34 $Y2=1.805
r110 46 48 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=9.34 $Y=1.89
+ $X2=9.34 $Y2=1.985
r111 45 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.34 $Y=1.72
+ $X2=9.34 $Y2=1.805
r112 44 76 8.93547 $w=1.7e-07 $l=3.3e-07 $layer=LI1_cond $X=9.34 $Y=1.01
+ $X2=9.34 $Y2=0.68
r113 44 45 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=9.34 $Y=1.01
+ $X2=9.34 $Y2=1.72
r114 42 57 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.255 $Y=1.805
+ $X2=9.34 $Y2=1.805
r115 42 43 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=9.255 $Y=1.805
+ $X2=8.525 $Y2=1.805
r116 38 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.44 $Y=1.89
+ $X2=8.525 $Y2=1.805
r117 38 40 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=8.44 $Y=1.89
+ $X2=8.44 $Y2=1.985
r118 37 56 7.02821 $w=1.7e-07 $l=1.34629e-07 $layer=LI1_cond $X=8.01 $Y=0.925
+ $X2=7.885 $Y2=0.945
r119 37 72 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=8.01 $Y=0.925
+ $X2=8.7 $Y2=0.925
r120 32 56 0.00168595 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=7.885 $Y=0.84
+ $X2=7.885 $Y2=0.945
r121 32 34 14.9818 $w=2.48e-07 $l=3.25e-07 $layer=LI1_cond $X=7.885 $Y=0.84
+ $X2=7.885 $Y2=0.515
r122 31 55 5.63431 $w=2.25e-07 $l=1.52069e-07 $layer=LI1_cond $X=6.38 $Y=0.925
+ $X2=6.255 $Y2=0.985
r123 30 56 7.02821 $w=1.7e-07 $l=1.34629e-07 $layer=LI1_cond $X=7.76 $Y=0.925
+ $X2=7.885 $Y2=0.945
r124 30 31 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=7.76 $Y=0.925
+ $X2=6.38 $Y2=0.925
r125 26 55 0.966048 $w=2.5e-07 $l=1.45e-07 $layer=LI1_cond $X=6.255 $Y=0.84
+ $X2=6.255 $Y2=0.985
r126 26 28 14.9818 $w=2.48e-07 $l=3.25e-07 $layer=LI1_cond $X=6.255 $Y=0.84
+ $X2=6.255 $Y2=0.515
r127 25 53 28.6053 $w=2.78e-07 $l=6.95e-07 $layer=LI1_cond $X=5.355 $Y=0.99
+ $X2=4.66 $Y2=0.99
r128 22 55 5.63431 $w=2.25e-07 $l=1.27475e-07 $layer=LI1_cond $X=6.13 $Y=0.99
+ $X2=6.255 $Y2=0.985
r129 22 25 31.898 $w=2.78e-07 $l=7.75e-07 $layer=LI1_cond $X=6.13 $Y=0.99
+ $X2=5.355 $Y2=0.99
r130 7 48 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=9.19
+ $Y=1.84 $X2=9.34 $Y2=1.985
r131 6 40 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=8.29
+ $Y=1.84 $X2=8.44 $Y2=1.985
r132 5 71 182 $w=1.7e-07 $l=6.21068e-07 $layer=licon1_NDIFF $count=1 $X=8.645
+ $Y=0.37 $X2=8.785 $Y2=0.925
r133 5 71 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=8.645
+ $Y=0.37 $X2=8.785 $Y2=0.515
r134 4 34 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.785
+ $Y=0.37 $X2=7.925 $Y2=0.515
r135 3 55 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=6.075
+ $Y=0.37 $X2=6.215 $Y2=0.965
r136 3 28 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=6.075
+ $Y=0.37 $X2=6.215 $Y2=0.515
r137 2 25 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=5.215
+ $Y=0.37 $X2=5.355 $Y2=0.95
r138 1 51 182 $w=1.7e-07 $l=6.39453e-07 $layer=licon1_NDIFF $count=1 $X=4.37
+ $Y=0.37 $X2=4.495 $Y2=0.95
.ends

.subckt PM_SKY130_FD_SC_LS__A311OI_4%A_34_74# 1 2 3 4 5 18 20 21 24 26 30 34 36
+ 37 40 41 43
r74 43 45 4.43516 $w=3.28e-07 $l=1.27e-07 $layer=LI1_cond $X=3.755 $Y=0.95
+ $X2=3.755 $Y2=1.077
r75 39 41 7.51706 $w=4.08e-07 $l=1.65e-07 $layer=LI1_cond $X=2.895 $Y=0.975
+ $X2=3.06 $Y2=0.975
r76 39 40 7.51706 $w=4.08e-07 $l=1.65e-07 $layer=LI1_cond $X=2.895 $Y=0.975
+ $X2=2.73 $Y2=0.975
r77 34 45 3.54104 $w=2.05e-07 $l=1.65e-07 $layer=LI1_cond $X=3.59 $Y=1.077
+ $X2=3.755 $Y2=1.077
r78 34 41 28.6741 $w=2.03e-07 $l=5.3e-07 $layer=LI1_cond $X=3.59 $Y=1.077
+ $X2=3.06 $Y2=1.077
r79 33 37 4.7579 $w=1.87e-07 $l=8.5e-08 $layer=LI1_cond $X=2.12 $Y=1.077
+ $X2=2.035 $Y2=1.077
r80 33 40 33.0022 $w=2.03e-07 $l=6.1e-07 $layer=LI1_cond $X=2.12 $Y=1.077
+ $X2=2.73 $Y2=1.077
r81 28 37 1.69765 $w=1.7e-07 $l=1.02e-07 $layer=LI1_cond $X=2.035 $Y=0.975
+ $X2=2.035 $Y2=1.077
r82 28 30 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=2.035 $Y=0.975
+ $X2=2.035 $Y2=0.515
r83 27 36 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.26 $Y=1.095
+ $X2=1.135 $Y2=1.095
r84 26 37 4.7579 $w=1.87e-07 $l=9.35682e-08 $layer=LI1_cond $X=1.95 $Y=1.095
+ $X2=2.035 $Y2=1.077
r85 26 27 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.95 $Y=1.095
+ $X2=1.26 $Y2=1.095
r86 22 36 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.135 $Y=1.01
+ $X2=1.135 $Y2=1.095
r87 22 24 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=1.135 $Y=1.01
+ $X2=1.135 $Y2=0.515
r88 20 36 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.01 $Y=1.095
+ $X2=1.135 $Y2=1.095
r89 20 21 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=1.01 $Y=1.095
+ $X2=0.4 $Y2=1.095
r90 16 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.275 $Y=1.01
+ $X2=0.4 $Y2=1.095
r91 16 18 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=0.275 $Y=1.01
+ $X2=0.275 $Y2=0.515
r92 5 43 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=3.615
+ $Y=0.37 $X2=3.755 $Y2=0.95
r93 4 39 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=2.755
+ $Y=0.37 $X2=2.895 $Y2=0.95
r94 3 30 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.895
+ $Y=0.37 $X2=2.035 $Y2=0.515
r95 2 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.035
+ $Y=0.37 $X2=1.175 $Y2=0.515
r96 1 18 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.17
+ $Y=0.37 $X2=0.315 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__A311OI_4%VGND 1 2 3 4 15 19 23 25 27 32 45 55 56 59
+ 62 66 72 74
r89 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r90 70 72 10.9168 $w=7.53e-07 $l=1.5e-07 $layer=LI1_cond $X=7.44 $Y=0.292
+ $X2=7.59 $Y2=0.292
r91 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r92 68 70 0.237631 $w=7.53e-07 $l=1.5e-08 $layer=LI1_cond $X=7.425 $Y=0.292
+ $X2=7.44 $Y2=0.292
r93 65 68 11.2479 $w=7.53e-07 $l=7.1e-07 $layer=LI1_cond $X=6.715 $Y=0.292
+ $X2=7.425 $Y2=0.292
r94 65 66 11.1544 $w=7.53e-07 $l=1.65e-07 $layer=LI1_cond $X=6.715 $Y=0.292
+ $X2=6.55 $Y2=0.292
r95 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r96 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r97 55 56 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r98 53 56 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=9.84
+ $Y2=0
r99 53 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=8.4
+ $Y2=0
r100 52 55 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=8.88 $Y=0 $X2=9.84
+ $Y2=0
r101 52 53 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r102 50 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.52 $Y=0 $X2=8.355
+ $Y2=0
r103 50 52 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=8.52 $Y=0 $X2=8.88
+ $Y2=0
r104 49 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.4
+ $Y2=0
r105 49 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=7.44
+ $Y2=0
r106 48 72 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=7.92 $Y=0 $X2=7.59
+ $Y2=0
r107 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r108 45 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.19 $Y=0 $X2=8.355
+ $Y2=0
r109 45 48 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=8.19 $Y=0 $X2=7.92
+ $Y2=0
r110 44 71 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=7.44
+ $Y2=0
r111 43 66 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=6.48 $Y=0 $X2=6.55
+ $Y2=0
r112 43 44 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r113 41 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r114 40 43 281.84 $w=1.68e-07 $l=4.32e-06 $layer=LI1_cond $X=2.16 $Y=0 $X2=6.48
+ $Y2=0
r115 40 41 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r116 38 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.77 $Y=0 $X2=1.605
+ $Y2=0
r117 38 40 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=1.77 $Y=0 $X2=2.16
+ $Y2=0
r118 36 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r119 36 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r120 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r121 33 59 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.83 $Y=0 $X2=0.705
+ $Y2=0
r122 33 35 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.83 $Y=0 $X2=1.2
+ $Y2=0
r123 32 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.44 $Y=0 $X2=1.605
+ $Y2=0
r124 32 35 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=1.44 $Y=0 $X2=1.2
+ $Y2=0
r125 30 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r126 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r127 27 59 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.58 $Y=0 $X2=0.705
+ $Y2=0
r128 27 29 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.58 $Y=0 $X2=0.24
+ $Y2=0
r129 25 44 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=6.48 $Y2=0
r130 25 41 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=2.16 $Y2=0
r131 21 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.355 $Y=0.085
+ $X2=8.355 $Y2=0
r132 21 23 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=8.355 $Y=0.085
+ $X2=8.355 $Y2=0.55
r133 17 62 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.605 $Y=0.085
+ $X2=1.605 $Y2=0
r134 17 19 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=1.605 $Y=0.085
+ $X2=1.605 $Y2=0.675
r135 13 59 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=0.085
+ $X2=0.705 $Y2=0
r136 13 15 27.1977 $w=2.48e-07 $l=5.9e-07 $layer=LI1_cond $X=0.705 $Y=0.085
+ $X2=0.705 $Y2=0.675
r137 4 23 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=8.215
+ $Y=0.37 $X2=8.355 $Y2=0.55
r138 3 68 121.333 $w=1.7e-07 $l=1.00598e-06 $layer=licon1_NDIFF $count=1
+ $X=6.505 $Y=0.37 $X2=7.425 $Y2=0.55
r139 3 65 121.333 $w=1.7e-07 $l=2.86182e-07 $layer=licon1_NDIFF $count=1
+ $X=6.505 $Y=0.37 $X2=6.715 $Y2=0.55
r140 2 19 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=1.465
+ $Y=0.37 $X2=1.605 $Y2=0.675
r141 1 15 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=0.605
+ $Y=0.37 $X2=0.745 $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_LS__A311OI_4%A_465_74# 1 2 3 4 22 25 26 28 29
c37 28 0 1.0484e-19 $X=5.785 $Y=0.515
r38 28 29 6.46688 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=5.785 $Y=0.515
+ $X2=5.62 $Y2=0.515
r39 24 26 4.02231 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=3.325 $Y=0.515
+ $X2=3.42 $Y2=0.515
r40 24 25 4.02231 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=3.325 $Y=0.515
+ $X2=3.23 $Y2=0.515
r41 22 25 30.8855 $w=2.48e-07 $l=6.7e-07 $layer=LI1_cond $X=2.56 $Y=0.475
+ $X2=3.23 $Y2=0.475
r42 20 22 4.02231 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=2.465 $Y=0.515
+ $X2=2.56 $Y2=0.515
r43 18 29 32.0379 $w=2.48e-07 $l=6.95e-07 $layer=LI1_cond $X=4.925 $Y=0.475
+ $X2=5.62 $Y2=0.475
r44 18 26 69.3771 $w=2.48e-07 $l=1.505e-06 $layer=LI1_cond $X=4.925 $Y=0.475
+ $X2=3.42 $Y2=0.475
r45 4 28 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=5.645
+ $Y=0.37 $X2=5.785 $Y2=0.515
r46 3 18 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=4.785
+ $Y=0.37 $X2=4.925 $Y2=0.515
r47 2 24 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.185
+ $Y=0.37 $X2=3.325 $Y2=0.515
r48 1 20 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.325
+ $Y=0.37 $X2=2.465 $Y2=0.515
.ends

