* File: sky130_fd_sc_ls__o32a_2.pxi.spice
* Created: Fri Aug 28 13:54:08 2020
* 
x_PM_SKY130_FD_SC_LS__O32A_2%A_83_264# N_A_83_264#_M1002_d N_A_83_264#_M1004_d
+ N_A_83_264#_c_80_n N_A_83_264#_c_88_n N_A_83_264#_M1008_g N_A_83_264#_M1007_g
+ N_A_83_264#_c_89_n N_A_83_264#_M1009_g N_A_83_264#_M1013_g N_A_83_264#_c_83_n
+ N_A_83_264#_c_97_p N_A_83_264#_c_137_p N_A_83_264#_c_91_n N_A_83_264#_c_92_n
+ N_A_83_264#_c_128_p N_A_83_264#_c_84_n N_A_83_264#_c_85_n N_A_83_264#_c_86_n
+ N_A_83_264#_c_112_p N_A_83_264#_c_115_p PM_SKY130_FD_SC_LS__O32A_2%A_83_264#
x_PM_SKY130_FD_SC_LS__O32A_2%A1 N_A1_c_189_n N_A1_M1001_g N_A1_M1005_g A1
+ N_A1_c_191_n PM_SKY130_FD_SC_LS__O32A_2%A1
x_PM_SKY130_FD_SC_LS__O32A_2%A2 N_A2_c_223_n N_A2_M1011_g N_A2_M1010_g A2
+ N_A2_c_225_n PM_SKY130_FD_SC_LS__O32A_2%A2
x_PM_SKY130_FD_SC_LS__O32A_2%A3 N_A3_c_255_n N_A3_M1004_g N_A3_M1003_g A3
+ N_A3_c_257_n PM_SKY130_FD_SC_LS__O32A_2%A3
x_PM_SKY130_FD_SC_LS__O32A_2%B2 N_B2_M1002_g N_B2_c_287_n N_B2_M1000_g B2
+ PM_SKY130_FD_SC_LS__O32A_2%B2
x_PM_SKY130_FD_SC_LS__O32A_2%B1 N_B1_c_323_n N_B1_M1012_g N_B1_c_317_n
+ N_B1_c_318_n N_B1_M1006_g N_B1_c_319_n N_B1_c_320_n B1 B1 B1 B1 B1
+ N_B1_c_322_n PM_SKY130_FD_SC_LS__O32A_2%B1
x_PM_SKY130_FD_SC_LS__O32A_2%VPWR N_VPWR_M1008_s N_VPWR_M1009_s N_VPWR_M1012_d
+ N_VPWR_c_354_n N_VPWR_c_355_n N_VPWR_c_356_n N_VPWR_c_357_n N_VPWR_c_358_n
+ N_VPWR_c_359_n VPWR N_VPWR_c_360_n N_VPWR_c_361_n N_VPWR_c_353_n
+ N_VPWR_c_363_n PM_SKY130_FD_SC_LS__O32A_2%VPWR
x_PM_SKY130_FD_SC_LS__O32A_2%X N_X_M1007_d N_X_M1008_d N_X_c_403_n N_X_c_404_n X
+ X X X N_X_c_405_n PM_SKY130_FD_SC_LS__O32A_2%X
x_PM_SKY130_FD_SC_LS__O32A_2%VGND N_VGND_M1007_s N_VGND_M1013_s N_VGND_M1010_d
+ N_VGND_c_447_n N_VGND_c_448_n N_VGND_c_449_n N_VGND_c_450_n N_VGND_c_451_n
+ N_VGND_c_452_n N_VGND_c_453_n N_VGND_c_454_n N_VGND_c_455_n N_VGND_c_456_n
+ VGND N_VGND_c_457_n N_VGND_c_458_n PM_SKY130_FD_SC_LS__O32A_2%VGND
x_PM_SKY130_FD_SC_LS__O32A_2%A_349_74# N_A_349_74#_M1005_d N_A_349_74#_M1003_d
+ N_A_349_74#_M1006_d N_A_349_74#_c_507_n N_A_349_74#_c_508_n
+ N_A_349_74#_c_509_n N_A_349_74#_c_510_n N_A_349_74#_c_527_n
+ N_A_349_74#_c_511_n N_A_349_74#_c_512_n PM_SKY130_FD_SC_LS__O32A_2%A_349_74#
cc_1 VNB N_A_83_264#_c_80_n 0.0150953f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.675
cc_2 VNB N_A_83_264#_M1007_g 0.0249445f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=0.74
cc_3 VNB N_A_83_264#_M1013_g 0.0241735f $X=-0.19 $Y=-0.245 $X2=1.1 $Y2=0.74
cc_4 VNB N_A_83_264#_c_83_n 2.18704e-19 $X=-0.19 $Y=-0.245 $X2=1.15 $Y2=1.95
cc_5 VNB N_A_83_264#_c_84_n 0.0105334f $X=-0.19 $Y=-0.245 $X2=4.1 $Y2=1.95
cc_6 VNB N_A_83_264#_c_85_n 0.0521656f $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=1.485
cc_7 VNB N_A_83_264#_c_86_n 0.00302828f $X=-0.19 $Y=-0.245 $X2=1.15 $Y2=1.485
cc_8 VNB N_A1_c_189_n 0.0247507f $X=-0.19 $Y=-0.245 $X2=3.245 $Y2=0.37
cc_9 VNB N_A1_M1005_g 0.0261215f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A1_c_191_n 0.00555649f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.32
cc_11 VNB N_A2_c_223_n 0.0266119f $X=-0.19 $Y=-0.245 $X2=3.245 $Y2=0.37
cc_12 VNB N_A2_M1010_g 0.0257807f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A2_c_225_n 0.00165774f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.32
cc_14 VNB N_A3_c_255_n 0.0266037f $X=-0.19 $Y=-0.245 $X2=3.245 $Y2=0.37
cc_15 VNB N_A3_M1003_g 0.0267316f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A3_c_257_n 0.00165645f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.32
cc_17 VNB N_B2_M1002_g 0.0357125f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_B2_c_287_n 0.0236669f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB B2 0.00601402f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.675
cc_20 VNB N_B1_c_317_n 0.0218972f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_B1_c_318_n 0.0274572f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_B1_c_319_n 0.0157488f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_23 VNB N_B1_c_320_n 0.0180432f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.32
cc_24 VNB B1 0.0118942f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=0.74
cc_25 VNB N_B1_c_322_n 0.0543697f $X=-0.19 $Y=-0.245 $X2=1.15 $Y2=1.95
cc_26 VNB N_VPWR_c_353_n 0.203486f $X=-0.19 $Y=-0.245 $X2=2.892 $Y2=2.035
cc_27 VNB N_X_c_403_n 0.00500933f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_28 VNB N_X_c_404_n 0.00239713f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_29 VNB N_X_c_405_n 0.00759022f $X=-0.19 $Y=-0.245 $X2=4.1 $Y2=1.045
cc_30 VNB N_VGND_c_447_n 0.0140441f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_31 VNB N_VGND_c_448_n 0.0226334f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=0.74
cc_32 VNB N_VGND_c_449_n 0.0175838f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.765
cc_33 VNB N_VGND_c_450_n 0.0178579f $X=-0.19 $Y=-0.245 $X2=1.1 $Y2=0.74
cc_34 VNB N_VGND_c_451_n 0.00899389f $X=-0.19 $Y=-0.245 $X2=1.15 $Y2=1.95
cc_35 VNB N_VGND_c_452_n 0.00829839f $X=-0.19 $Y=-0.245 $X2=1.235 $Y2=2.035
cc_36 VNB N_VGND_c_453_n 0.019013f $X=-0.19 $Y=-0.245 $X2=2.892 $Y2=2.715
cc_37 VNB N_VGND_c_454_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=2.9 $Y2=2.715
cc_38 VNB N_VGND_c_455_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=4.015 $Y2=2.035
cc_39 VNB N_VGND_c_456_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=3.11 $Y2=2.035
cc_40 VNB N_VGND_c_457_n 0.0589592f $X=-0.19 $Y=-0.245 $X2=4.02 $Y2=0.88
cc_41 VNB N_VGND_c_458_n 0.27806f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.47
cc_42 VNB N_A_349_74#_c_507_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.32
cc_43 VNB N_A_349_74#_c_508_n 0.0183106f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=0.74
cc_44 VNB N_A_349_74#_c_509_n 0.00851793f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_349_74#_c_510_n 0.00261637f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.765
cc_46 VNB N_A_349_74#_c_511_n 0.00879016f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_47 VNB N_A_349_74#_c_512_n 0.00311899f $X=-0.19 $Y=-0.245 $X2=2.675 $Y2=2.035
cc_48 VPB N_A_83_264#_c_80_n 0.00111912f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.675
cc_49 VPB N_A_83_264#_c_88_n 0.0258256f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_50 VPB N_A_83_264#_c_89_n 0.0166755f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.765
cc_51 VPB N_A_83_264#_c_83_n 0.00279969f $X=-0.19 $Y=1.66 $X2=1.15 $Y2=1.95
cc_52 VPB N_A_83_264#_c_91_n 0.00499005f $X=-0.19 $Y=1.66 $X2=2.9 $Y2=2.715
cc_53 VPB N_A_83_264#_c_92_n 0.00378081f $X=-0.19 $Y=1.66 $X2=4.015 $Y2=2.035
cc_54 VPB N_A_83_264#_c_84_n 0.00503195f $X=-0.19 $Y=1.66 $X2=4.1 $Y2=1.95
cc_55 VPB N_A_83_264#_c_85_n 0.0074211f $X=-0.19 $Y=1.66 $X2=1.04 $Y2=1.485
cc_56 VPB N_A1_c_189_n 0.02753f $X=-0.19 $Y=1.66 $X2=3.245 $Y2=0.37
cc_57 VPB N_A1_c_191_n 0.00326892f $X=-0.19 $Y=1.66 $X2=0.67 $Y2=1.32
cc_58 VPB N_A2_c_223_n 0.0267962f $X=-0.19 $Y=1.66 $X2=3.245 $Y2=0.37
cc_59 VPB N_A2_c_225_n 0.00241954f $X=-0.19 $Y=1.66 $X2=0.67 $Y2=1.32
cc_60 VPB N_A3_c_255_n 0.0280587f $X=-0.19 $Y=1.66 $X2=3.245 $Y2=0.37
cc_61 VPB N_A3_c_257_n 0.00246053f $X=-0.19 $Y=1.66 $X2=0.67 $Y2=1.32
cc_62 VPB N_B2_c_287_n 0.0279241f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB B2 0.00496903f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.675
cc_64 VPB N_B1_c_323_n 0.0176208f $X=-0.19 $Y=1.66 $X2=3.245 $Y2=0.37
cc_65 VPB N_B1_c_319_n 0.00689027f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_66 VPB B1 0.0736665f $X=-0.19 $Y=1.66 $X2=0.67 $Y2=0.74
cc_67 VPB N_VPWR_c_354_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_68 VPB N_VPWR_c_355_n 0.0587306f $X=-0.19 $Y=1.66 $X2=0.67 $Y2=1.32
cc_69 VPB N_VPWR_c_356_n 0.0144674f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_70 VPB N_VPWR_c_357_n 0.0248954f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_358_n 0.06763f $X=-0.19 $Y=1.66 $X2=2.675 $Y2=2.035
cc_72 VPB N_VPWR_c_359_n 0.00632158f $X=-0.19 $Y=1.66 $X2=1.235 $Y2=2.035
cc_73 VPB N_VPWR_c_360_n 0.0194151f $X=-0.19 $Y=1.66 $X2=2.9 $Y2=2.715
cc_74 VPB N_VPWR_c_361_n 0.0208395f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_353_n 0.124453f $X=-0.19 $Y=1.66 $X2=2.892 $Y2=2.035
cc_76 VPB N_VPWR_c_363_n 0.0102647f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.617
cc_77 VPB X 0.00472837f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_78 VPB X 0.00257348f $X=-0.19 $Y=1.66 $X2=1.235 $Y2=2.035
cc_79 VPB N_X_c_405_n 0.00123421f $X=-0.19 $Y=1.66 $X2=4.1 $Y2=1.045
cc_80 N_A_83_264#_c_89_n N_A1_c_189_n 0.0127624f $X=0.955 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_81 N_A_83_264#_c_83_n N_A1_c_189_n 0.00385953f $X=1.15 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_82 N_A_83_264#_c_97_p N_A1_c_189_n 0.0161824f $X=2.675 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_83 N_A_83_264#_c_85_n N_A1_c_189_n 0.0213682f $X=1.04 $Y=1.485 $X2=-0.19
+ $Y2=-0.245
cc_84 N_A_83_264#_c_86_n N_A1_c_189_n 0.00170854f $X=1.15 $Y=1.485 $X2=-0.19
+ $Y2=-0.245
cc_85 N_A_83_264#_M1013_g N_A1_M1005_g 0.0233513f $X=1.1 $Y=0.74 $X2=0 $Y2=0
cc_86 N_A_83_264#_c_85_n N_A1_M1005_g 8.1421e-19 $X=1.04 $Y=1.485 $X2=0 $Y2=0
cc_87 N_A_83_264#_c_86_n N_A1_M1005_g 5.77738e-19 $X=1.15 $Y=1.485 $X2=0 $Y2=0
cc_88 N_A_83_264#_c_83_n N_A1_c_191_n 0.0096933f $X=1.15 $Y=1.95 $X2=0 $Y2=0
cc_89 N_A_83_264#_c_97_p N_A1_c_191_n 0.0250874f $X=2.675 $Y=2.035 $X2=0 $Y2=0
cc_90 N_A_83_264#_c_85_n N_A1_c_191_n 3.50433e-19 $X=1.04 $Y=1.485 $X2=0 $Y2=0
cc_91 N_A_83_264#_c_86_n N_A1_c_191_n 0.0231673f $X=1.15 $Y=1.485 $X2=0 $Y2=0
cc_92 N_A_83_264#_c_97_p N_A2_c_223_n 0.0162159f $X=2.675 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_93 N_A_83_264#_c_91_n N_A2_c_223_n 0.00344942f $X=2.9 $Y=2.715 $X2=-0.19
+ $Y2=-0.245
cc_94 N_A_83_264#_c_97_p N_A2_c_225_n 0.0226548f $X=2.675 $Y=2.035 $X2=0 $Y2=0
cc_95 N_A_83_264#_c_97_p N_A3_c_255_n 0.0124019f $X=2.675 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_96 N_A_83_264#_c_91_n N_A3_c_255_n 0.0265233f $X=2.9 $Y=2.715 $X2=-0.19
+ $Y2=-0.245
cc_97 N_A_83_264#_c_112_p N_A3_c_255_n 0.00395226f $X=2.9 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_98 N_A_83_264#_c_97_p N_A3_c_257_n 0.0104762f $X=2.675 $Y=2.035 $X2=0 $Y2=0
cc_99 N_A_83_264#_c_112_p N_A3_c_257_n 0.0132222f $X=2.9 $Y=2.035 $X2=0 $Y2=0
cc_100 N_A_83_264#_c_115_p N_B2_M1002_g 0.00419034f $X=4.02 $Y=0.88 $X2=0 $Y2=0
cc_101 N_A_83_264#_c_91_n N_B2_c_287_n 0.00607101f $X=2.9 $Y=2.715 $X2=0 $Y2=0
cc_102 N_A_83_264#_c_92_n N_B2_c_287_n 0.0143839f $X=4.015 $Y=2.035 $X2=0 $Y2=0
cc_103 N_A_83_264#_c_84_n N_B2_c_287_n 2.63846e-19 $X=4.1 $Y=1.95 $X2=0 $Y2=0
cc_104 N_A_83_264#_c_112_p N_B2_c_287_n 0.00268655f $X=2.9 $Y=2.035 $X2=0 $Y2=0
cc_105 N_A_83_264#_c_115_p N_B2_c_287_n 0.00363041f $X=4.02 $Y=0.88 $X2=0 $Y2=0
cc_106 N_A_83_264#_c_92_n B2 0.0427777f $X=4.015 $Y=2.035 $X2=0 $Y2=0
cc_107 N_A_83_264#_c_84_n B2 0.0217679f $X=4.1 $Y=1.95 $X2=0 $Y2=0
cc_108 N_A_83_264#_c_115_p B2 0.0247412f $X=4.02 $Y=0.88 $X2=0 $Y2=0
cc_109 N_A_83_264#_c_92_n N_B1_c_323_n 0.0200732f $X=4.015 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_110 N_A_83_264#_c_84_n N_B1_c_323_n 0.00600924f $X=4.1 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_111 N_A_83_264#_c_92_n N_B1_c_317_n 0.00396467f $X=4.015 $Y=2.035 $X2=0 $Y2=0
cc_112 N_A_83_264#_c_84_n N_B1_c_317_n 0.0113712f $X=4.1 $Y=1.95 $X2=0 $Y2=0
cc_113 N_A_83_264#_c_128_p N_B1_c_318_n 0.00517368f $X=4.1 $Y=1.045 $X2=0 $Y2=0
cc_114 N_A_83_264#_c_84_n N_B1_c_318_n 0.00830667f $X=4.1 $Y=1.95 $X2=0 $Y2=0
cc_115 N_A_83_264#_c_84_n N_B1_c_319_n 0.004573f $X=4.1 $Y=1.95 $X2=0 $Y2=0
cc_116 N_A_83_264#_c_115_p N_B1_c_319_n 0.0101464f $X=4.02 $Y=0.88 $X2=0 $Y2=0
cc_117 N_A_83_264#_c_84_n N_B1_c_320_n 0.00891863f $X=4.1 $Y=1.95 $X2=0 $Y2=0
cc_118 N_A_83_264#_c_92_n B1 0.0150384f $X=4.015 $Y=2.035 $X2=0 $Y2=0
cc_119 N_A_83_264#_c_84_n B1 0.0582284f $X=4.1 $Y=1.95 $X2=0 $Y2=0
cc_120 N_A_83_264#_c_83_n N_VPWR_M1009_s 0.00234639f $X=1.15 $Y=1.95 $X2=0 $Y2=0
cc_121 N_A_83_264#_c_97_p N_VPWR_M1009_s 0.0123554f $X=2.675 $Y=2.035 $X2=0
+ $Y2=0
cc_122 N_A_83_264#_c_137_p N_VPWR_M1009_s 0.00300113f $X=1.235 $Y=2.035 $X2=0
+ $Y2=0
cc_123 N_A_83_264#_c_92_n N_VPWR_M1012_d 0.0054166f $X=4.015 $Y=2.035 $X2=0
+ $Y2=0
cc_124 N_A_83_264#_c_84_n N_VPWR_M1012_d 0.00193485f $X=4.1 $Y=1.95 $X2=0 $Y2=0
cc_125 N_A_83_264#_c_88_n N_VPWR_c_355_n 0.00954146f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_126 N_A_83_264#_c_89_n N_VPWR_c_356_n 0.007483f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_127 N_A_83_264#_c_97_p N_VPWR_c_356_n 0.0248f $X=2.675 $Y=2.035 $X2=0 $Y2=0
cc_128 N_A_83_264#_c_137_p N_VPWR_c_356_n 0.0129456f $X=1.235 $Y=2.035 $X2=0
+ $Y2=0
cc_129 N_A_83_264#_c_85_n N_VPWR_c_356_n 4.01954e-19 $X=1.04 $Y=1.485 $X2=0
+ $Y2=0
cc_130 N_A_83_264#_c_92_n N_VPWR_c_357_n 0.0230547f $X=4.015 $Y=2.035 $X2=0
+ $Y2=0
cc_131 N_A_83_264#_c_91_n N_VPWR_c_358_n 0.0137085f $X=2.9 $Y=2.715 $X2=0 $Y2=0
cc_132 N_A_83_264#_c_88_n N_VPWR_c_360_n 0.00411612f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_133 N_A_83_264#_c_89_n N_VPWR_c_360_n 0.00445602f $X=0.955 $Y=1.765 $X2=0
+ $Y2=0
cc_134 N_A_83_264#_c_88_n N_VPWR_c_353_n 0.00751023f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_135 N_A_83_264#_c_89_n N_VPWR_c_353_n 0.00861719f $X=0.955 $Y=1.765 $X2=0
+ $Y2=0
cc_136 N_A_83_264#_c_91_n N_VPWR_c_353_n 0.0149817f $X=2.9 $Y=2.715 $X2=0 $Y2=0
cc_137 N_A_83_264#_M1007_g N_X_c_403_n 0.0127873f $X=0.67 $Y=0.74 $X2=0 $Y2=0
cc_138 N_A_83_264#_M1013_g N_X_c_403_n 0.002387f $X=1.1 $Y=0.74 $X2=0 $Y2=0
cc_139 N_A_83_264#_c_85_n N_X_c_403_n 0.00341242f $X=1.04 $Y=1.485 $X2=0 $Y2=0
cc_140 N_A_83_264#_c_86_n N_X_c_403_n 0.0120032f $X=1.15 $Y=1.485 $X2=0 $Y2=0
cc_141 N_A_83_264#_M1007_g N_X_c_404_n 0.00875007f $X=0.67 $Y=0.74 $X2=0 $Y2=0
cc_142 N_A_83_264#_M1013_g N_X_c_404_n 0.00755147f $X=1.1 $Y=0.74 $X2=0 $Y2=0
cc_143 N_A_83_264#_c_88_n X 0.00240464f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_144 N_A_83_264#_c_89_n X 0.00219207f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_145 N_A_83_264#_c_83_n X 0.00565815f $X=1.15 $Y=1.95 $X2=0 $Y2=0
cc_146 N_A_83_264#_c_85_n X 0.00345893f $X=1.04 $Y=1.485 $X2=0 $Y2=0
cc_147 N_A_83_264#_c_86_n X 0.00153915f $X=1.15 $Y=1.485 $X2=0 $Y2=0
cc_148 N_A_83_264#_c_88_n X 0.0130738f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_149 N_A_83_264#_c_89_n X 0.012608f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_150 N_A_83_264#_c_80_n N_X_c_405_n 0.0100858f $X=0.505 $Y=1.675 $X2=0 $Y2=0
cc_151 N_A_83_264#_c_88_n N_X_c_405_n 0.00745465f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_152 N_A_83_264#_M1007_g N_X_c_405_n 0.00770058f $X=0.67 $Y=0.74 $X2=0 $Y2=0
cc_153 N_A_83_264#_c_89_n N_X_c_405_n 4.19687e-19 $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_154 N_A_83_264#_M1013_g N_X_c_405_n 0.00109865f $X=1.1 $Y=0.74 $X2=0 $Y2=0
cc_155 N_A_83_264#_c_83_n N_X_c_405_n 0.00756912f $X=1.15 $Y=1.95 $X2=0 $Y2=0
cc_156 N_A_83_264#_c_85_n N_X_c_405_n 0.0136932f $X=1.04 $Y=1.485 $X2=0 $Y2=0
cc_157 N_A_83_264#_c_86_n N_X_c_405_n 0.0243803f $X=1.15 $Y=1.485 $X2=0 $Y2=0
cc_158 N_A_83_264#_c_97_p A_346_368# 0.0117119f $X=2.675 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_159 N_A_83_264#_c_97_p A_430_368# 0.018186f $X=2.675 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_160 N_A_83_264#_c_92_n A_652_368# 0.015282f $X=4.015 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_161 N_A_83_264#_M1007_g N_VGND_c_448_n 0.00671933f $X=0.67 $Y=0.74 $X2=0
+ $Y2=0
cc_162 N_A_83_264#_M1007_g N_VGND_c_449_n 0.00453882f $X=0.67 $Y=0.74 $X2=0
+ $Y2=0
cc_163 N_A_83_264#_M1013_g N_VGND_c_450_n 0.00806966f $X=1.1 $Y=0.74 $X2=0 $Y2=0
cc_164 N_A_83_264#_c_86_n N_VGND_c_450_n 0.00114473f $X=1.15 $Y=1.485 $X2=0
+ $Y2=0
cc_165 N_A_83_264#_c_85_n N_VGND_c_452_n 0.0039922f $X=1.04 $Y=1.485 $X2=0 $Y2=0
cc_166 N_A_83_264#_M1007_g N_VGND_c_453_n 0.00434272f $X=0.67 $Y=0.74 $X2=0
+ $Y2=0
cc_167 N_A_83_264#_M1013_g N_VGND_c_453_n 0.00434272f $X=1.1 $Y=0.74 $X2=0 $Y2=0
cc_168 N_A_83_264#_M1007_g N_VGND_c_458_n 0.00824408f $X=0.67 $Y=0.74 $X2=0
+ $Y2=0
cc_169 N_A_83_264#_M1013_g N_VGND_c_458_n 0.00821312f $X=1.1 $Y=0.74 $X2=0 $Y2=0
cc_170 N_A_83_264#_M1013_g N_A_349_74#_c_509_n 2.49809e-19 $X=1.1 $Y=0.74 $X2=0
+ $Y2=0
cc_171 N_A_83_264#_M1002_d N_A_349_74#_c_511_n 0.0136122f $X=3.245 $Y=0.37 $X2=0
+ $Y2=0
cc_172 N_A_83_264#_c_128_p N_A_349_74#_c_511_n 0.0076481f $X=4.1 $Y=1.045 $X2=0
+ $Y2=0
cc_173 N_A_83_264#_c_115_p N_A_349_74#_c_511_n 0.0478533f $X=4.02 $Y=0.88 $X2=0
+ $Y2=0
cc_174 N_A1_c_189_n N_A2_c_223_n 0.0805105f $X=1.655 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_175 N_A1_c_191_n N_A2_c_223_n 0.00257062f $X=1.58 $Y=1.515 $X2=-0.19
+ $Y2=-0.245
cc_176 N_A1_M1005_g N_A2_M1010_g 0.019972f $X=1.67 $Y=0.74 $X2=0 $Y2=0
cc_177 N_A1_c_189_n N_A2_c_225_n 5.26454e-19 $X=1.655 $Y=1.765 $X2=0 $Y2=0
cc_178 N_A1_c_191_n N_A2_c_225_n 0.0317261f $X=1.58 $Y=1.515 $X2=0 $Y2=0
cc_179 N_A1_c_189_n N_VPWR_c_356_n 0.0203583f $X=1.655 $Y=1.765 $X2=0 $Y2=0
cc_180 N_A1_c_189_n N_VPWR_c_358_n 0.00427043f $X=1.655 $Y=1.765 $X2=0 $Y2=0
cc_181 N_A1_c_189_n N_VPWR_c_353_n 0.00443985f $X=1.655 $Y=1.765 $X2=0 $Y2=0
cc_182 N_A1_c_189_n X 7.29858e-19 $X=1.655 $Y=1.765 $X2=0 $Y2=0
cc_183 N_A1_c_189_n N_VGND_c_450_n 0.00101787f $X=1.655 $Y=1.765 $X2=0 $Y2=0
cc_184 N_A1_M1005_g N_VGND_c_450_n 0.00666787f $X=1.67 $Y=0.74 $X2=0 $Y2=0
cc_185 N_A1_c_191_n N_VGND_c_450_n 0.00945165f $X=1.58 $Y=1.515 $X2=0 $Y2=0
cc_186 N_A1_M1005_g N_VGND_c_455_n 0.00434272f $X=1.67 $Y=0.74 $X2=0 $Y2=0
cc_187 N_A1_M1005_g N_VGND_c_458_n 0.0082141f $X=1.67 $Y=0.74 $X2=0 $Y2=0
cc_188 N_A1_M1005_g N_A_349_74#_c_507_n 0.00795429f $X=1.67 $Y=0.74 $X2=0 $Y2=0
cc_189 N_A1_M1005_g N_A_349_74#_c_509_n 0.00350994f $X=1.67 $Y=0.74 $X2=0 $Y2=0
cc_190 N_A1_c_191_n N_A_349_74#_c_509_n 0.00648331f $X=1.58 $Y=1.515 $X2=0 $Y2=0
cc_191 N_A2_c_223_n N_A3_c_255_n 0.0624378f $X=2.075 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_192 N_A2_c_225_n N_A3_c_255_n 0.00179181f $X=2.15 $Y=1.515 $X2=-0.19
+ $Y2=-0.245
cc_193 N_A2_M1010_g N_A3_M1003_g 0.0260254f $X=2.1 $Y=0.74 $X2=0 $Y2=0
cc_194 N_A2_c_223_n N_A3_c_257_n 0.00127792f $X=2.075 $Y=1.765 $X2=0 $Y2=0
cc_195 N_A2_c_225_n N_A3_c_257_n 0.0277337f $X=2.15 $Y=1.515 $X2=0 $Y2=0
cc_196 N_A2_c_223_n N_VPWR_c_356_n 0.00327604f $X=2.075 $Y=1.765 $X2=0 $Y2=0
cc_197 N_A2_c_223_n N_VPWR_c_358_n 0.0049405f $X=2.075 $Y=1.765 $X2=0 $Y2=0
cc_198 N_A2_c_223_n N_VPWR_c_353_n 0.00508379f $X=2.075 $Y=1.765 $X2=0 $Y2=0
cc_199 N_A2_M1010_g N_VGND_c_451_n 0.00484409f $X=2.1 $Y=0.74 $X2=0 $Y2=0
cc_200 N_A2_M1010_g N_VGND_c_455_n 0.00434272f $X=2.1 $Y=0.74 $X2=0 $Y2=0
cc_201 N_A2_M1010_g N_VGND_c_458_n 0.0082141f $X=2.1 $Y=0.74 $X2=0 $Y2=0
cc_202 N_A2_M1010_g N_A_349_74#_c_507_n 0.00966073f $X=2.1 $Y=0.74 $X2=0 $Y2=0
cc_203 N_A2_c_223_n N_A_349_74#_c_508_n 9.79877e-19 $X=2.075 $Y=1.765 $X2=0
+ $Y2=0
cc_204 N_A2_M1010_g N_A_349_74#_c_508_n 0.0117933f $X=2.1 $Y=0.74 $X2=0 $Y2=0
cc_205 N_A2_c_225_n N_A_349_74#_c_508_n 0.019847f $X=2.15 $Y=1.515 $X2=0 $Y2=0
cc_206 N_A2_c_223_n N_A_349_74#_c_509_n 3.05922e-19 $X=2.075 $Y=1.765 $X2=0
+ $Y2=0
cc_207 N_A2_M1010_g N_A_349_74#_c_509_n 0.0015571f $X=2.1 $Y=0.74 $X2=0 $Y2=0
cc_208 N_A2_c_225_n N_A_349_74#_c_509_n 0.00541082f $X=2.15 $Y=1.515 $X2=0 $Y2=0
cc_209 N_A2_M1010_g N_A_349_74#_c_527_n 5.94859e-19 $X=2.1 $Y=0.74 $X2=0 $Y2=0
cc_210 N_A3_M1003_g N_B2_M1002_g 0.0247403f $X=2.67 $Y=0.74 $X2=0 $Y2=0
cc_211 N_A3_c_255_n N_B2_c_287_n 0.0508832f $X=2.615 $Y=1.765 $X2=0 $Y2=0
cc_212 N_A3_c_257_n N_B2_c_287_n 8.19164e-19 $X=2.69 $Y=1.515 $X2=0 $Y2=0
cc_213 N_A3_c_255_n B2 0.0013426f $X=2.615 $Y=1.765 $X2=0 $Y2=0
cc_214 N_A3_c_257_n B2 0.0261927f $X=2.69 $Y=1.515 $X2=0 $Y2=0
cc_215 N_A3_c_255_n N_VPWR_c_358_n 0.00481822f $X=2.615 $Y=1.765 $X2=0 $Y2=0
cc_216 N_A3_c_255_n N_VPWR_c_353_n 0.00508379f $X=2.615 $Y=1.765 $X2=0 $Y2=0
cc_217 N_A3_M1003_g N_VGND_c_451_n 0.00622568f $X=2.67 $Y=0.74 $X2=0 $Y2=0
cc_218 N_A3_M1003_g N_VGND_c_457_n 0.00433139f $X=2.67 $Y=0.74 $X2=0 $Y2=0
cc_219 N_A3_M1003_g N_VGND_c_458_n 0.00818355f $X=2.67 $Y=0.74 $X2=0 $Y2=0
cc_220 N_A3_M1003_g N_A_349_74#_c_507_n 6.28869e-19 $X=2.67 $Y=0.74 $X2=0 $Y2=0
cc_221 N_A3_c_255_n N_A_349_74#_c_508_n 0.00134355f $X=2.615 $Y=1.765 $X2=0
+ $Y2=0
cc_222 N_A3_M1003_g N_A_349_74#_c_508_n 0.0133747f $X=2.67 $Y=0.74 $X2=0 $Y2=0
cc_223 N_A3_c_257_n N_A_349_74#_c_508_n 0.0259036f $X=2.69 $Y=1.515 $X2=0 $Y2=0
cc_224 N_A3_M1003_g N_A_349_74#_c_510_n 0.00227367f $X=2.67 $Y=0.74 $X2=0 $Y2=0
cc_225 N_A3_M1003_g N_A_349_74#_c_527_n 0.00745726f $X=2.67 $Y=0.74 $X2=0 $Y2=0
cc_226 N_B2_c_287_n N_B1_c_323_n 0.0335204f $X=3.185 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_227 B2 N_B1_c_323_n 8.97324e-19 $X=3.515 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_228 N_B2_c_287_n N_B1_c_319_n 0.0178581f $X=3.185 $Y=1.765 $X2=0 $Y2=0
cc_229 B2 N_B1_c_319_n 0.012373f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_230 B2 N_B1_c_320_n 2.68126e-19 $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_231 N_B2_c_287_n N_VPWR_c_357_n 0.00305222f $X=3.185 $Y=1.765 $X2=0 $Y2=0
cc_232 N_B2_c_287_n N_VPWR_c_358_n 0.0049405f $X=3.185 $Y=1.765 $X2=0 $Y2=0
cc_233 N_B2_c_287_n N_VPWR_c_353_n 0.00508379f $X=3.185 $Y=1.765 $X2=0 $Y2=0
cc_234 N_B2_M1002_g N_VGND_c_457_n 0.00291649f $X=3.17 $Y=0.74 $X2=0 $Y2=0
cc_235 N_B2_M1002_g N_VGND_c_458_n 0.00364831f $X=3.17 $Y=0.74 $X2=0 $Y2=0
cc_236 N_B2_M1002_g N_A_349_74#_c_508_n 0.0028014f $X=3.17 $Y=0.74 $X2=0 $Y2=0
cc_237 N_B2_M1002_g N_A_349_74#_c_511_n 0.0161408f $X=3.17 $Y=0.74 $X2=0 $Y2=0
cc_238 N_B1_c_323_n N_VPWR_c_357_n 0.0164769f $X=3.755 $Y=1.765 $X2=0 $Y2=0
cc_239 B1 N_VPWR_c_357_n 0.0430855f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_240 N_B1_c_323_n N_VPWR_c_358_n 0.00443511f $X=3.755 $Y=1.765 $X2=0 $Y2=0
cc_241 B1 N_VPWR_c_361_n 0.0107254f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_242 N_B1_c_323_n N_VPWR_c_353_n 0.00460931f $X=3.755 $Y=1.765 $X2=0 $Y2=0
cc_243 B1 N_VPWR_c_353_n 0.0114362f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_244 N_B1_c_318_n N_VGND_c_457_n 0.00291649f $X=4.235 $Y=1.22 $X2=0 $Y2=0
cc_245 N_B1_c_318_n N_VGND_c_458_n 0.00367994f $X=4.235 $Y=1.22 $X2=0 $Y2=0
cc_246 N_B1_c_318_n N_A_349_74#_c_511_n 0.0141061f $X=4.235 $Y=1.22 $X2=0 $Y2=0
cc_247 B1 N_A_349_74#_c_512_n 0.0231725f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_248 N_B1_c_322_n N_A_349_74#_c_512_n 0.00178757f $X=4.52 $Y=1.385 $X2=0 $Y2=0
cc_249 N_VPWR_c_355_n X 0.0887573f $X=0.28 $Y=1.985 $X2=0 $Y2=0
cc_250 N_VPWR_c_356_n X 0.0270879f $X=1.425 $Y=2.385 $X2=0 $Y2=0
cc_251 N_VPWR_c_360_n X 0.0158009f $X=1.065 $Y=3.33 $X2=0 $Y2=0
cc_252 N_VPWR_c_353_n X 0.0129424f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_253 N_VPWR_c_355_n N_VGND_c_449_n 0.00876255f $X=0.28 $Y=1.985 $X2=0 $Y2=0
cc_254 N_X_c_403_n N_VGND_M1007_s 0.00163897f $X=0.885 $Y=0.96 $X2=-0.19
+ $Y2=-0.245
cc_255 N_X_c_404_n N_VGND_c_448_n 0.016559f $X=0.885 $Y=0.515 $X2=0 $Y2=0
cc_256 N_X_c_403_n N_VGND_c_449_n 0.013787f $X=0.885 $Y=0.96 $X2=0 $Y2=0
cc_257 N_X_c_404_n N_VGND_c_449_n 0.0073154f $X=0.885 $Y=0.515 $X2=0 $Y2=0
cc_258 N_X_c_405_n N_VGND_c_449_n 7.75603e-19 $X=0.715 $Y=1.82 $X2=0 $Y2=0
cc_259 N_X_c_403_n N_VGND_c_450_n 0.00753583f $X=0.885 $Y=0.96 $X2=0 $Y2=0
cc_260 N_X_c_404_n N_VGND_c_450_n 0.0236791f $X=0.885 $Y=0.515 $X2=0 $Y2=0
cc_261 N_X_c_404_n N_VGND_c_453_n 0.014379f $X=0.885 $Y=0.515 $X2=0 $Y2=0
cc_262 N_X_c_404_n N_VGND_c_458_n 0.0118382f $X=0.885 $Y=0.515 $X2=0 $Y2=0
cc_263 N_VGND_c_450_n N_A_349_74#_c_507_n 0.0255177f $X=1.385 $Y=0.515 $X2=0
+ $Y2=0
cc_264 N_VGND_c_451_n N_A_349_74#_c_507_n 0.0191765f $X=2.385 $Y=0.675 $X2=0
+ $Y2=0
cc_265 N_VGND_c_455_n N_A_349_74#_c_507_n 0.0144922f $X=2.22 $Y=0 $X2=0 $Y2=0
cc_266 N_VGND_c_458_n N_A_349_74#_c_507_n 0.0118826f $X=4.56 $Y=0 $X2=0 $Y2=0
cc_267 N_VGND_M1010_d N_A_349_74#_c_508_n 0.00358162f $X=2.175 $Y=0.37 $X2=0
+ $Y2=0
cc_268 N_VGND_c_451_n N_A_349_74#_c_508_n 0.0248957f $X=2.385 $Y=0.675 $X2=0
+ $Y2=0
cc_269 N_VGND_c_450_n N_A_349_74#_c_509_n 0.00584871f $X=1.385 $Y=0.515 $X2=0
+ $Y2=0
cc_270 N_VGND_c_451_n N_A_349_74#_c_510_n 0.00795492f $X=2.385 $Y=0.675 $X2=0
+ $Y2=0
cc_271 N_VGND_c_457_n N_A_349_74#_c_510_n 0.0146502f $X=4.56 $Y=0 $X2=0 $Y2=0
cc_272 N_VGND_c_458_n N_A_349_74#_c_510_n 0.0120674f $X=4.56 $Y=0 $X2=0 $Y2=0
cc_273 N_VGND_c_457_n N_A_349_74#_c_511_n 0.0518789f $X=4.56 $Y=0 $X2=0 $Y2=0
cc_274 N_VGND_c_458_n N_A_349_74#_c_511_n 0.0447063f $X=4.56 $Y=0 $X2=0 $Y2=0
cc_275 N_VGND_c_457_n N_A_349_74#_c_512_n 0.0115764f $X=4.56 $Y=0 $X2=0 $Y2=0
cc_276 N_VGND_c_458_n N_A_349_74#_c_512_n 0.00959296f $X=4.56 $Y=0 $X2=0 $Y2=0
