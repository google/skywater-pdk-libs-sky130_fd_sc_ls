* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
M1000 Y C1 a_834_74# VNB nshort w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=1.0434e+12p ps=1.022e+07u
M1001 VPWR B1 Y VPB phighvt w=1.12e+06u l=150000u
+  ad=2.3744e+12p pd=1.544e+07u as=1.5008e+12p ps=1.164e+07u
M1002 VGND A2 a_27_74# VNB nshort w=740000u l=150000u
+  ad=9.472e+11p pd=8.48e+06u as=1.4578e+12p ps=1.43e+07u
M1003 VPWR C1 Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_30_368# A2 Y VPB phighvt w=1.12e+06u l=150000u
+  ad=1.7808e+12p pd=1.438e+07u as=0p ps=0u
M1005 VGND A2 a_27_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_834_74# B1 a_27_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_30_368# A1 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_27_74# A2 VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR A1 a_30_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_27_74# A1 VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Y A2 a_30_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_27_74# B1 a_834_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR A1 a_30_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_27_74# A2 VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_834_74# C1 Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_30_368# A2 Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_27_74# A1 VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_834_74# C1 Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_834_74# B1 a_27_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_27_74# B1 a_834_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 Y B1 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND A1 a_27_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_30_368# A1 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND A1 a_27_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 Y A2 a_30_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 Y C1 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 Y C1 a_834_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
