* File: sky130_fd_sc_ls__decap_8.spice
* Created: Fri Aug 28 13:11:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__decap_8.pex.spice"
.subckt sky130_fd_sc_ls__decap_8  VNB VPB VGND VPWR
* 
* VPWR	VPWR
* VGND	VGND
* VPB	VPB
* VNB	VNB
MM1000 N_VGND_M1000_s N_VPWR_M1000_g N_VGND_M1000_s VNB NSHORT L=1 W=0.42
+ AD=0.05775 AS=0.2436 PD=0.695 PS=2 NRD=0 NRS=0 M=1 R=0.42 SA=500000 SB=500001
+ A=0.42 P=2.84 MULT=1
MM1001 N_VGND_M1000_s N_VPWR_M1001_g N_VGND_M1000_s VNB NSHORT L=1 W=0.42
+ AD=0.2688 AS=0.05775 PD=2.12 PS=0.695 NRD=0 NRS=0 M=1 R=0.42 SA=500001
+ SB=500000 A=0.42 P=2.84 MULT=1
MM1002 N_VPWR_M1002_s N_VGND_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=1 W=1
+ AD=0.1375 AS=0.665 PD=1.275 PS=3.33 NRD=0 NRS=1.9503 M=1 R=1 SA=500000
+ SB=500001 A=1 P=4 MULT=1
MM1003 N_VPWR_M1002_s N_VGND_M1003_g N_VPWR_M1002_s VPB PHIGHVT L=1 W=1 AD=0.63
+ AS=0.1375 PD=3.26 PS=1.275 NRD=0 NRS=0 M=1 R=1 SA=500001 SB=500000 A=1 P=4
+ MULT=1
DX4_noxref VNB VPB NWDIODE A=7.8492 P=12.16
*
.include "sky130_fd_sc_ls__decap_8.pxi.spice"
*
.ends
*
*
