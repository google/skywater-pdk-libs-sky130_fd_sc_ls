* File: sky130_fd_sc_ls__nor2b_1.pex.spice
* Created: Fri Aug 28 13:37:39 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__NOR2B_1%B_N 1 3 4 6 8 9
r27 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.275
+ $Y=1.385 $X2=0.275 $Y2=1.385
r28 9 13 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.275 $Y=1.295
+ $X2=0.275 $Y2=1.385
r29 8 12 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.615 $Y=1.385
+ $X2=0.275 $Y2=1.385
r30 4 8 48.459 $w=1.66e-07 $l=1.72337e-07 $layer=POLY_cond $X=0.72 $Y=1.22
+ $X2=0.705 $Y2=1.385
r31 4 6 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=0.72 $Y=1.22 $X2=0.72
+ $Y2=0.835
r32 1 8 110.887 $w=1.66e-07 $l=3.8e-07 $layer=POLY_cond $X=0.705 $Y=1.765
+ $X2=0.705 $Y2=1.385
r33 1 3 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.705 $Y=1.765
+ $X2=0.705 $Y2=2.26
.ends

.subckt PM_SKY130_FD_SC_LS__NOR2B_1%A 1 3 4 6 7
c30 4 0 8.85114e-20 $X=1.33 $Y=1.22
r31 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.2
+ $Y=1.385 $X2=1.2 $Y2=1.385
r32 7 11 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=1.2 $Y=1.295 $X2=1.2
+ $Y2=1.385
r33 4 10 38.578 $w=2.95e-07 $l=2.13014e-07 $layer=POLY_cond $X=1.33 $Y=1.22
+ $X2=1.22 $Y2=1.385
r34 4 6 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.33 $Y=1.22 $X2=1.33
+ $Y2=0.74
r35 1 10 73.7068 $w=2.95e-07 $l=4.24853e-07 $layer=POLY_cond $X=1.315 $Y=1.765
+ $X2=1.22 $Y2=1.385
r36 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.315 $Y=1.765
+ $X2=1.315 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__NOR2B_1%A_27_112# 1 2 7 9 12 14 20 23 24 26 28
c63 14 0 8.85114e-20 $X=0.61 $Y=0.845
r64 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.81
+ $Y=1.485 $X2=1.81 $Y2=1.485
r65 25 26 2.76166 $w=1.7e-07 $l=2.33e-07 $layer=LI1_cond $X=0.78 $Y=1.805
+ $X2=0.547 $Y2=1.805
r66 24 28 11.9755 $w=3.26e-07 $l=4.15692e-07 $layer=LI1_cond $X=1.535 $Y=1.805
+ $X2=1.755 $Y2=1.485
r67 24 25 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=1.535 $Y=1.805
+ $X2=0.78 $Y2=1.805
r68 23 26 3.70735 $w=2.5e-07 $l=1.85699e-07 $layer=LI1_cond $X=0.695 $Y=1.72
+ $X2=0.547 $Y2=1.805
r69 22 23 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=0.695 $Y=1.01
+ $X2=0.695 $Y2=1.72
r70 18 26 3.70735 $w=2.5e-07 $l=1.13666e-07 $layer=LI1_cond $X=0.48 $Y=1.89
+ $X2=0.547 $Y2=1.805
r71 18 20 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=0.48 $Y=1.89
+ $X2=0.48 $Y2=1.985
r72 14 22 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.61 $Y=0.845
+ $X2=0.695 $Y2=1.01
r73 14 16 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=0.61 $Y=0.845
+ $X2=0.505 $Y2=0.845
r74 10 29 38.6072 $w=2.91e-07 $l=1.77059e-07 $layer=POLY_cond $X=1.835 $Y=1.32
+ $X2=1.81 $Y2=1.485
r75 10 12 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.835 $Y=1.32
+ $X2=1.835 $Y2=0.74
r76 7 29 57.6553 $w=2.91e-07 $l=3.15278e-07 $layer=POLY_cond $X=1.735 $Y=1.765
+ $X2=1.81 $Y2=1.485
r77 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.735 $Y=1.765
+ $X2=1.735 $Y2=2.4
r78 2 20 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.335
+ $Y=1.84 $X2=0.48 $Y2=1.985
r79 1 16 182 $w=1.7e-07 $l=4.92291e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.56 $X2=0.505 $Y2=0.845
.ends

.subckt PM_SKY130_FD_SC_LS__NOR2B_1%VPWR 1 6 10 12 19 20 23
r23 19 20 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r24 17 23 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.255 $Y=3.33
+ $X2=1.09 $Y2=3.33
r25 17 19 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=1.255 $Y=3.33
+ $X2=2.16 $Y2=3.33
r26 14 15 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r27 12 23 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.925 $Y=3.33
+ $X2=1.09 $Y2=3.33
r28 12 14 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=0.925 $Y=3.33
+ $X2=0.72 $Y2=3.33
r29 10 20 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r30 10 15 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r31 10 23 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r32 6 9 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.09 $Y=2.145 $X2=1.09
+ $Y2=2.825
r33 4 23 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.09 $Y=3.245 $X2=1.09
+ $Y2=3.33
r34 4 9 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=1.09 $Y=3.245 $X2=1.09
+ $Y2=2.825
r35 1 9 600 $w=1.7e-07 $l=1.12941e-06 $layer=licon1_PDIFF $count=1 $X=0.78
+ $Y=1.84 $X2=1.09 $Y2=2.825
r36 1 6 300 $w=1.7e-07 $l=4.36635e-07 $layer=licon1_PDIFF $count=2 $X=0.78
+ $Y=1.84 $X2=1.09 $Y2=2.145
.ends

.subckt PM_SKY130_FD_SC_LS__NOR2B_1%Y 1 2 9 11 12 15 16 17 32 33 36
r31 32 33 8.83531 $w=4.38e-07 $l=1.65e-07 $layer=LI1_cond $X=2.095 $Y=1.985
+ $X2=2.095 $Y2=1.82
r32 22 36 0.130959 $w=4.38e-07 $l=5e-09 $layer=LI1_cond $X=2.095 $Y=2.04
+ $X2=2.095 $Y2=2.035
r33 17 29 1.04768 $w=4.38e-07 $l=4e-08 $layer=LI1_cond $X=2.095 $Y=2.775
+ $X2=2.095 $Y2=2.815
r34 16 17 9.691 $w=4.38e-07 $l=3.7e-07 $layer=LI1_cond $X=2.095 $Y=2.405
+ $X2=2.095 $Y2=2.775
r35 15 36 1.04768 $w=4.38e-07 $l=4e-08 $layer=LI1_cond $X=2.095 $Y=1.995
+ $X2=2.095 $Y2=2.035
r36 15 32 0.261919 $w=4.38e-07 $l=1e-08 $layer=LI1_cond $X=2.095 $Y=1.995
+ $X2=2.095 $Y2=1.985
r37 15 16 8.51236 $w=4.38e-07 $l=3.25e-07 $layer=LI1_cond $X=2.095 $Y=2.08
+ $X2=2.095 $Y2=2.405
r38 15 22 1.04768 $w=4.38e-07 $l=4e-08 $layer=LI1_cond $X=2.095 $Y=2.08
+ $X2=2.095 $Y2=2.04
r39 13 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.23 $Y=1.15
+ $X2=2.23 $Y2=1.82
r40 11 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.145 $Y=1.065
+ $X2=2.23 $Y2=1.15
r41 11 12 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=2.145 $Y=1.065
+ $X2=1.785 $Y2=1.065
r42 7 12 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.66 $Y=0.98
+ $X2=1.785 $Y2=1.065
r43 7 9 21.4354 $w=2.48e-07 $l=4.65e-07 $layer=LI1_cond $X=1.66 $Y=0.98 $X2=1.66
+ $Y2=0.515
r44 2 32 400 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=1 $X=1.81
+ $Y=1.84 $X2=1.965 $Y2=1.985
r45 2 29 400 $w=1.7e-07 $l=1.04964e-06 $layer=licon1_PDIFF $count=1 $X=1.81
+ $Y=1.84 $X2=1.965 $Y2=2.815
r46 1 9 91 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_NDIFF $count=2 $X=1.405
+ $Y=0.37 $X2=1.62 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__NOR2B_1%VGND 1 2 9 11 13 16 17 18 24 30
r29 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r30 27 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r31 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r32 24 29 4.14667 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=1.955 $Y=0 $X2=2.177
+ $Y2=0
r33 24 26 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.955 $Y=0 $X2=1.68
+ $Y2=0
r34 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r35 18 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r36 18 22 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r37 16 21 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=0.95 $Y=0 $X2=0.72
+ $Y2=0
r38 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.95 $Y=0 $X2=1.115
+ $Y2=0
r39 15 26 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=1.28 $Y=0 $X2=1.68
+ $Y2=0
r40 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.28 $Y=0 $X2=1.115
+ $Y2=0
r41 11 29 3.17537 $w=2.75e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.092 $Y=0.085
+ $X2=2.177 $Y2=0
r42 11 13 23.4679 $w=2.73e-07 $l=5.6e-07 $layer=LI1_cond $X=2.092 $Y=0.085
+ $X2=2.092 $Y2=0.645
r43 7 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.115 $Y=0.085
+ $X2=1.115 $Y2=0
r44 7 9 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=1.115 $Y=0.085
+ $X2=1.115 $Y2=0.515
r45 2 13 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=1.91
+ $Y=0.37 $X2=2.05 $Y2=0.645
r46 1 9 91 $w=1.7e-07 $l=3.4176e-07 $layer=licon1_NDIFF $count=2 $X=0.795
+ $Y=0.56 $X2=1.115 $Y2=0.515
.ends

