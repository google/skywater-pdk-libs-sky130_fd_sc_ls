* File: sky130_fd_sc_ls__and3_2.spice
* Created: Wed Sep  2 10:54:51 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__and3_2.pex.spice"
.subckt sky130_fd_sc_ls__and3_2  VNB VPB A B C VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* C	C
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1006 A_133_136# N_A_M1006_g N_A_41_384#_M1006_s VNB NSHORT L=0.15 W=0.64
+ AD=0.1344 AS=0.1824 PD=1.06 PS=1.85 NRD=29.052 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75002.1 A=0.096 P=1.58 MULT=1
MM1005 A_247_136# N_B_M1005_g A_133_136# VNB NSHORT L=0.15 W=0.64 AD=0.0768
+ AS=0.1344 PD=0.88 PS=1.06 NRD=12.18 NRS=29.052 M=1 R=4.26667 SA=75000.8
+ SB=75001.5 A=0.096 P=1.58 MULT=1
MM1003 N_VGND_M1003_d N_C_M1003_g A_247_136# VNB NSHORT L=0.15 W=0.64 AD=0.15789
+ AS=0.0768 PD=1.2429 PS=0.88 NRD=14.988 NRS=12.18 M=1 R=4.26667 SA=75001.2
+ SB=75001.1 A=0.096 P=1.58 MULT=1
MM1007 N_VGND_M1003_d N_A_41_384#_M1007_g N_X_M1007_s VNB NSHORT L=0.15 W=0.74
+ AD=0.18256 AS=0.1184 PD=1.4371 PS=1.06 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75001.2 SB=75000.9 A=0.111 P=1.78 MULT=1
MM1009 N_VGND_M1009_d N_A_41_384#_M1009_g N_X_M1007_s VNB NSHORT L=0.15 W=0.74
+ AD=0.3552 AS=0.1184 PD=2.44 PS=1.06 NRD=27.564 NRS=6.48 M=1 R=4.93333
+ SA=75001.7 SB=75000.4 A=0.111 P=1.78 MULT=1
MM1000 N_VPWR_M1000_d N_A_M1000_g N_A_41_384#_M1000_s VPB PHIGHVT L=0.15 W=0.84
+ AD=0.1764 AS=0.2478 PD=1.26 PS=2.27 NRD=14.0658 NRS=2.3443 M=1 R=5.6
+ SA=75000.2 SB=75002.5 A=0.126 P=1.98 MULT=1
MM1008 N_A_41_384#_M1008_d N_B_M1008_g N_VPWR_M1000_d VPB PHIGHVT L=0.15 W=0.84
+ AD=0.126 AS=0.1764 PD=1.14 PS=1.26 NRD=2.3443 NRS=18.7544 M=1 R=5.6 SA=75000.8
+ SB=75001.9 A=0.126 P=1.98 MULT=1
MM1002 N_VPWR_M1002_d N_C_M1002_g N_A_41_384#_M1008_d VPB PHIGHVT L=0.15 W=0.84
+ AD=0.243857 AS=0.126 PD=1.44857 PS=1.14 NRD=121.943 NRS=0 M=1 R=5.6 SA=75001.2
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1001 N_X_M1001_d N_A_41_384#_M1001_g N_VPWR_M1002_d VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.325143 PD=1.42 PS=1.93143 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75001.5 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1004 N_X_M1001_d N_A_41_384#_M1004_g N_VPWR_M1004_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.4088 PD=1.42 PS=2.97 NRD=1.7533 NRS=14.0658 M=1 R=7.46667
+ SA=75002 SB=75000.3 A=0.168 P=2.54 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9564 P=11.2
c_55 VPB 0 1.15e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_ls__and3_2.pxi.spice"
*
.ends
*
*
