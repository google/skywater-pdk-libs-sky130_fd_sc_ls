* File: sky130_fd_sc_ls__sdfstp_4.pxi.spice
* Created: Fri Aug 28 14:04:53 2020
* 
x_PM_SKY130_FD_SC_LS__SDFSTP_4%SCE N_SCE_M1045_g N_SCE_c_346_n N_SCE_M1043_g
+ N_SCE_c_347_n N_SCE_M1044_g N_SCE_M1017_g N_SCE_c_341_n N_SCE_c_342_n
+ N_SCE_c_343_n SCE N_SCE_c_344_n N_SCE_c_345_n PM_SKY130_FD_SC_LS__SDFSTP_4%SCE
x_PM_SKY130_FD_SC_LS__SDFSTP_4%A_27_74# N_A_27_74#_M1045_s N_A_27_74#_M1043_s
+ N_A_27_74#_M1041_g N_A_27_74#_c_423_n N_A_27_74#_M1012_g N_A_27_74#_c_417_n
+ N_A_27_74#_c_418_n N_A_27_74#_c_435_n N_A_27_74#_c_419_n N_A_27_74#_c_420_n
+ N_A_27_74#_c_425_n N_A_27_74#_c_421_n N_A_27_74#_c_426_n N_A_27_74#_c_422_n
+ PM_SKY130_FD_SC_LS__SDFSTP_4%A_27_74#
x_PM_SKY130_FD_SC_LS__SDFSTP_4%D N_D_c_492_n N_D_M1034_g N_D_M1042_g D
+ N_D_c_494_n PM_SKY130_FD_SC_LS__SDFSTP_4%D
x_PM_SKY130_FD_SC_LS__SDFSTP_4%SCD N_SCD_M1018_g N_SCD_c_528_n N_SCD_c_532_n
+ N_SCD_M1001_g SCD SCD SCD N_SCD_c_530_n PM_SKY130_FD_SC_LS__SDFSTP_4%SCD
x_PM_SKY130_FD_SC_LS__SDFSTP_4%CLK N_CLK_c_569_n N_CLK_M1025_g N_CLK_c_570_n
+ N_CLK_M1028_g CLK PM_SKY130_FD_SC_LS__SDFSTP_4%CLK
x_PM_SKY130_FD_SC_LS__SDFSTP_4%A_803_74# N_A_803_74#_M1021_d N_A_803_74#_M1040_d
+ N_A_803_74#_c_622_n N_A_803_74#_c_623_n N_A_803_74#_M1029_g
+ N_A_803_74#_c_603_n N_A_803_74#_M1020_g N_A_803_74#_c_605_n
+ N_A_803_74#_c_606_n N_A_803_74#_c_607_n N_A_803_74#_M1010_g
+ N_A_803_74#_c_608_n N_A_803_74#_c_609_n N_A_803_74#_M1036_g
+ N_A_803_74#_c_625_n N_A_803_74#_c_626_n N_A_803_74#_M1009_g
+ N_A_803_74#_c_610_n N_A_803_74#_c_611_n N_A_803_74#_c_612_n
+ N_A_803_74#_c_613_n N_A_803_74#_c_614_n N_A_803_74#_c_628_n
+ N_A_803_74#_c_615_n N_A_803_74#_c_630_n N_A_803_74#_c_650_p
+ N_A_803_74#_c_651_p N_A_803_74#_c_631_n N_A_803_74#_c_632_n
+ N_A_803_74#_c_633_n N_A_803_74#_c_634_n N_A_803_74#_c_635_n
+ N_A_803_74#_c_636_n N_A_803_74#_c_637_n N_A_803_74#_c_638_n
+ N_A_803_74#_c_639_n N_A_803_74#_c_616_n N_A_803_74#_c_617_n
+ N_A_803_74#_c_640_n N_A_803_74#_c_641_n N_A_803_74#_c_642_n
+ N_A_803_74#_c_643_n N_A_803_74#_c_618_n N_A_803_74#_c_619_n
+ N_A_803_74#_c_646_n N_A_803_74#_c_647_n N_A_803_74#_c_620_n
+ N_A_803_74#_c_621_n PM_SKY130_FD_SC_LS__SDFSTP_4%A_803_74#
x_PM_SKY130_FD_SC_LS__SDFSTP_4%A_1201_55# N_A_1201_55#_M1024_s
+ N_A_1201_55#_M1031_d N_A_1201_55#_M1019_g N_A_1201_55#_c_907_n
+ N_A_1201_55#_M1004_g N_A_1201_55#_c_901_n N_A_1201_55#_c_902_n
+ N_A_1201_55#_c_909_n N_A_1201_55#_c_903_n N_A_1201_55#_c_910_n
+ N_A_1201_55#_c_904_n N_A_1201_55#_c_905_n N_A_1201_55#_c_911_n
+ N_A_1201_55#_c_906_n PM_SKY130_FD_SC_LS__SDFSTP_4%A_1201_55#
x_PM_SKY130_FD_SC_LS__SDFSTP_4%A_1017_81# N_A_1017_81#_M1002_d
+ N_A_1017_81#_M1029_d N_A_1017_81#_c_1002_n N_A_1017_81#_c_1003_n
+ N_A_1017_81#_M1031_g N_A_1017_81#_c_987_n N_A_1017_81#_M1024_g
+ N_A_1017_81#_c_988_n N_A_1017_81#_c_1005_n N_A_1017_81#_M1035_g
+ N_A_1017_81#_c_989_n N_A_1017_81#_M1014_g N_A_1017_81#_c_990_n
+ N_A_1017_81#_c_1007_n N_A_1017_81#_M1047_g N_A_1017_81#_c_991_n
+ N_A_1017_81#_M1048_g N_A_1017_81#_c_992_n N_A_1017_81#_c_993_n
+ N_A_1017_81#_c_1009_n N_A_1017_81#_c_1010_n N_A_1017_81#_c_994_n
+ N_A_1017_81#_c_995_n N_A_1017_81#_c_996_n N_A_1017_81#_c_997_n
+ N_A_1017_81#_c_1011_n N_A_1017_81#_c_998_n N_A_1017_81#_c_999_n
+ N_A_1017_81#_c_1000_n N_A_1017_81#_c_1001_n
+ PM_SKY130_FD_SC_LS__SDFSTP_4%A_1017_81#
x_PM_SKY130_FD_SC_LS__SDFSTP_4%SET_B N_SET_B_c_1169_n N_SET_B_c_1170_n
+ N_SET_B_M1006_g N_SET_B_M1003_g N_SET_B_c_1171_n N_SET_B_c_1172_n
+ N_SET_B_c_1173_n N_SET_B_M1005_g N_SET_B_M1038_g N_SET_B_c_1174_n
+ N_SET_B_c_1163_n N_SET_B_c_1176_n SET_B N_SET_B_c_1165_n N_SET_B_c_1166_n
+ N_SET_B_c_1167_n N_SET_B_c_1168_n PM_SKY130_FD_SC_LS__SDFSTP_4%SET_B
x_PM_SKY130_FD_SC_LS__SDFSTP_4%A_616_74# N_A_616_74#_M1025_s N_A_616_74#_M1028_s
+ N_A_616_74#_M1021_g N_A_616_74#_c_1317_n N_A_616_74#_M1040_g
+ N_A_616_74#_c_1305_n N_A_616_74#_c_1306_n N_A_616_74#_c_1319_n
+ N_A_616_74#_c_1320_n N_A_616_74#_c_1307_n N_A_616_74#_c_1308_n
+ N_A_616_74#_c_1321_n N_A_616_74#_c_1322_n N_A_616_74#_M1002_g
+ N_A_616_74#_c_1323_n N_A_616_74#_M1032_g N_A_616_74#_c_1324_n
+ N_A_616_74#_c_1325_n N_A_616_74#_M1016_g N_A_616_74#_c_1326_n
+ N_A_616_74#_c_1327_n N_A_616_74#_c_1328_n N_A_616_74#_M1030_g
+ N_A_616_74#_c_1310_n N_A_616_74#_c_1311_n N_A_616_74#_M1026_g
+ N_A_616_74#_c_1331_n N_A_616_74#_c_1332_n N_A_616_74#_c_1333_n
+ N_A_616_74#_c_1313_n N_A_616_74#_c_1314_n N_A_616_74#_c_1335_n
+ N_A_616_74#_c_1336_n N_A_616_74#_c_1315_n N_A_616_74#_c_1316_n
+ PM_SKY130_FD_SC_LS__SDFSTP_4%A_616_74#
x_PM_SKY130_FD_SC_LS__SDFSTP_4%A_2191_180# N_A_2191_180#_M1039_d
+ N_A_2191_180#_M1013_s N_A_2191_180#_c_1504_n N_A_2191_180#_M1007_g
+ N_A_2191_180#_c_1513_n N_A_2191_180#_M1046_g N_A_2191_180#_c_1505_n
+ N_A_2191_180#_c_1506_n N_A_2191_180#_c_1514_n N_A_2191_180#_c_1507_n
+ N_A_2191_180#_c_1508_n N_A_2191_180#_c_1509_n N_A_2191_180#_c_1516_n
+ N_A_2191_180#_c_1510_n N_A_2191_180#_c_1517_n N_A_2191_180#_c_1511_n
+ PM_SKY130_FD_SC_LS__SDFSTP_4%A_2191_180#
x_PM_SKY130_FD_SC_LS__SDFSTP_4%A_1823_524# N_A_1823_524#_M1010_d
+ N_A_1823_524#_M1036_d N_A_1823_524#_M1016_s N_A_1823_524#_M1030_s
+ N_A_1823_524#_M1005_d N_A_1823_524#_M1039_g N_A_1823_524#_c_1621_n
+ N_A_1823_524#_c_1622_n N_A_1823_524#_M1013_g N_A_1823_524#_c_1623_n
+ N_A_1823_524#_c_1624_n N_A_1823_524#_M1022_g N_A_1823_524#_M1008_g
+ N_A_1823_524#_c_1626_n N_A_1823_524#_M1033_g N_A_1823_524#_c_1627_n
+ N_A_1823_524#_c_1612_n N_A_1823_524#_c_1628_n N_A_1823_524#_c_1613_n
+ N_A_1823_524#_c_1614_n N_A_1823_524#_c_1647_n N_A_1823_524#_c_1615_n
+ N_A_1823_524#_c_1629_n N_A_1823_524#_c_1630_n N_A_1823_524#_c_1616_n
+ N_A_1823_524#_c_1617_n N_A_1823_524#_c_1618_n N_A_1823_524#_c_1632_n
+ N_A_1823_524#_c_1633_n N_A_1823_524#_c_1619_n N_A_1823_524#_c_1620_n
+ N_A_1823_524#_c_1635_n N_A_1823_524#_c_1636_n N_A_1823_524#_c_1637_n
+ N_A_1823_524#_c_1638_n N_A_1823_524#_c_1700_n
+ PM_SKY130_FD_SC_LS__SDFSTP_4%A_1823_524#
x_PM_SKY130_FD_SC_LS__SDFSTP_4%A_2580_74# N_A_2580_74#_M1008_s
+ N_A_2580_74#_M1022_d N_A_2580_74#_M1000_g N_A_2580_74#_c_1838_n
+ N_A_2580_74#_M1011_g N_A_2580_74#_M1015_g N_A_2580_74#_c_1839_n
+ N_A_2580_74#_M1037_g N_A_2580_74#_M1023_g N_A_2580_74#_c_1840_n
+ N_A_2580_74#_M1049_g N_A_2580_74#_c_1829_n N_A_2580_74#_c_1830_n
+ N_A_2580_74#_M1027_g N_A_2580_74#_c_1832_n N_A_2580_74#_c_1843_n
+ N_A_2580_74#_M1050_g N_A_2580_74#_c_1833_n N_A_2580_74#_c_1834_n
+ N_A_2580_74#_c_1835_n N_A_2580_74#_c_1836_n N_A_2580_74#_c_1837_n
+ PM_SKY130_FD_SC_LS__SDFSTP_4%A_2580_74#
x_PM_SKY130_FD_SC_LS__SDFSTP_4%VPWR N_VPWR_M1043_d N_VPWR_M1001_d N_VPWR_M1028_d
+ N_VPWR_M1004_d N_VPWR_M1006_d N_VPWR_M1047_s N_VPWR_M1046_d N_VPWR_M1013_d
+ N_VPWR_M1033_s N_VPWR_M1037_s N_VPWR_M1050_s N_VPWR_c_1948_n N_VPWR_c_1949_n
+ N_VPWR_c_1950_n N_VPWR_c_1951_n N_VPWR_c_1952_n N_VPWR_c_1953_n
+ N_VPWR_c_1954_n N_VPWR_c_1955_n N_VPWR_c_1956_n N_VPWR_c_1957_n
+ N_VPWR_c_1958_n N_VPWR_c_1959_n N_VPWR_c_1960_n N_VPWR_c_1961_n
+ N_VPWR_c_1962_n N_VPWR_c_1963_n N_VPWR_c_1964_n VPWR N_VPWR_c_1965_n
+ N_VPWR_c_1966_n N_VPWR_c_1967_n N_VPWR_c_1968_n N_VPWR_c_1969_n
+ N_VPWR_c_1970_n N_VPWR_c_1971_n N_VPWR_c_1972_n N_VPWR_c_1973_n
+ N_VPWR_c_1974_n N_VPWR_c_1975_n N_VPWR_c_1976_n N_VPWR_c_1977_n
+ N_VPWR_c_1978_n N_VPWR_c_1979_n N_VPWR_c_1980_n N_VPWR_c_1947_n
+ PM_SKY130_FD_SC_LS__SDFSTP_4%VPWR
x_PM_SKY130_FD_SC_LS__SDFSTP_4%A_288_464# N_A_288_464#_M1042_d
+ N_A_288_464#_M1002_s N_A_288_464#_M1034_d N_A_288_464#_M1029_s
+ N_A_288_464#_c_2173_n N_A_288_464#_c_2161_n N_A_288_464#_c_2162_n
+ N_A_288_464#_c_2163_n N_A_288_464#_c_2164_n N_A_288_464#_c_2168_n
+ N_A_288_464#_c_2169_n N_A_288_464#_c_2165_n N_A_288_464#_c_2182_n
+ N_A_288_464#_c_2194_n N_A_288_464#_c_2171_n N_A_288_464#_c_2166_n
+ N_A_288_464#_c_2172_n PM_SKY130_FD_SC_LS__SDFSTP_4%A_288_464#
x_PM_SKY130_FD_SC_LS__SDFSTP_4%A_1620_373# N_A_1620_373#_M1035_d
+ N_A_1620_373#_M1016_d N_A_1620_373#_c_2293_n N_A_1620_373#_c_2289_n
+ N_A_1620_373#_c_2290_n N_A_1620_373#_c_2291_n
+ PM_SKY130_FD_SC_LS__SDFSTP_4%A_1620_373#
x_PM_SKY130_FD_SC_LS__SDFSTP_4%Q N_Q_M1000_d N_Q_M1023_d N_Q_M1011_d N_Q_M1049_d
+ N_Q_c_2330_n N_Q_c_2339_n N_Q_c_2340_n N_Q_c_2331_n N_Q_c_2332_n N_Q_c_2341_n
+ N_Q_c_2333_n N_Q_c_2342_n N_Q_c_2334_n N_Q_c_2335_n N_Q_c_2376_n N_Q_c_2336_n
+ Q N_Q_c_2338_n PM_SKY130_FD_SC_LS__SDFSTP_4%Q
x_PM_SKY130_FD_SC_LS__SDFSTP_4%VGND N_VGND_M1045_d N_VGND_M1018_d N_VGND_M1025_d
+ N_VGND_M1019_d N_VGND_M1003_d N_VGND_M1048_d N_VGND_M1038_d N_VGND_M1008_d
+ N_VGND_M1015_s N_VGND_M1027_s N_VGND_c_2414_n N_VGND_c_2415_n N_VGND_c_2416_n
+ N_VGND_c_2417_n N_VGND_c_2418_n N_VGND_c_2419_n N_VGND_c_2420_n
+ N_VGND_c_2421_n N_VGND_c_2422_n N_VGND_c_2423_n N_VGND_c_2424_n
+ N_VGND_c_2425_n N_VGND_c_2426_n N_VGND_c_2427_n VGND N_VGND_c_2428_n
+ N_VGND_c_2429_n N_VGND_c_2430_n N_VGND_c_2431_n N_VGND_c_2432_n
+ N_VGND_c_2433_n N_VGND_c_2434_n N_VGND_c_2435_n N_VGND_c_2436_n
+ N_VGND_c_2437_n N_VGND_c_2438_n N_VGND_c_2439_n N_VGND_c_2440_n
+ N_VGND_c_2441_n N_VGND_c_2442_n N_VGND_c_2443_n N_VGND_c_2444_n
+ PM_SKY130_FD_SC_LS__SDFSTP_4%VGND
x_PM_SKY130_FD_SC_LS__SDFSTP_4%A_1677_74# N_A_1677_74#_M1014_s
+ N_A_1677_74#_M1010_s N_A_1677_74#_c_2590_n N_A_1677_74#_c_2591_n
+ N_A_1677_74#_c_2592_n N_A_1677_74#_c_2593_n
+ PM_SKY130_FD_SC_LS__SDFSTP_4%A_1677_74#
cc_1 VNB N_SCE_M1045_g 0.0611748f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.58
cc_2 VNB N_SCE_M1017_g 0.0364115f $X=-0.19 $Y=-0.245 $X2=2.01 $Y2=0.58
cc_3 VNB N_SCE_c_341_n 0.0228124f $X=-0.19 $Y=-0.245 $X2=1.715 $Y2=1.495
cc_4 VNB N_SCE_c_342_n 0.00253001f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=1.495
cc_5 VNB N_SCE_c_343_n 0.00689606f $X=-0.19 $Y=-0.245 $X2=1.88 $Y2=1.415
cc_6 VNB N_SCE_c_344_n 0.0287309f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.645
cc_7 VNB N_SCE_c_345_n 0.0354393f $X=-0.19 $Y=-0.245 $X2=2.01 $Y2=1.415
cc_8 VNB N_A_27_74#_c_417_n 0.0247424f $X=-0.19 $Y=-0.245 $X2=1.715 $Y2=1.495
cc_9 VNB N_A_27_74#_c_418_n 0.0211704f $X=-0.19 $Y=-0.245 $X2=1.88 $Y2=1.415
cc_10 VNB N_A_27_74#_c_419_n 0.0086247f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.58
cc_11 VNB N_A_27_74#_c_420_n 0.0312447f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.645
cc_12 VNB N_A_27_74#_c_421_n 0.017304f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_74#_c_422_n 0.0190463f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_D_M1042_g 0.0665196f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.64
cc_15 VNB N_SCD_M1018_g 0.0310746f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.58
cc_16 VNB N_SCD_c_528_n 0.0290233f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.64
cc_17 VNB SCD 0.00507163f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=2.64
cc_18 VNB N_SCD_c_530_n 0.037007f $X=-0.19 $Y=-0.245 $X2=1.88 $Y2=1.415
cc_19 VNB N_CLK_c_569_n 0.0202389f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.48
cc_20 VNB N_CLK_c_570_n 0.0394431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB CLK 0.00726127f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.64
cc_22 VNB N_A_803_74#_c_603_n 0.0122973f $X=-0.19 $Y=-0.245 $X2=2.01 $Y2=0.58
cc_23 VNB N_A_803_74#_M1020_g 0.0550132f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=1.495
cc_24 VNB N_A_803_74#_c_605_n 0.0184994f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_803_74#_c_606_n 0.012774f $X=-0.19 $Y=-0.245 $X2=1.88 $Y2=1.495
cc_26 VNB N_A_803_74#_c_607_n 0.0185719f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_803_74#_c_608_n 0.0185984f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.58
cc_28 VNB N_A_803_74#_c_609_n 0.0147194f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.645
cc_29 VNB N_A_803_74#_c_610_n 0.0096129f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_803_74#_c_611_n 0.00666874f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_803_74#_c_612_n 0.0017973f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_803_74#_c_613_n 0.0162254f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_803_74#_c_614_n 0.00264685f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_803_74#_c_615_n 0.00203104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_803_74#_c_616_n 0.00189663f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_803_74#_c_617_n 0.0029028f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_803_74#_c_618_n 0.00167208f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_803_74#_c_619_n 0.0228906f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_803_74#_c_620_n 0.0283661f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_803_74#_c_621_n 0.0186444f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_1201_55#_c_901_n 0.0212464f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_1201_55#_c_902_n 0.00998322f $X=-0.19 $Y=-0.245 $X2=1.715
+ $Y2=1.495
cc_43 VNB N_A_1201_55#_c_903_n 0.00762292f $X=-0.19 $Y=-0.245 $X2=1.88 $Y2=1.495
cc_44 VNB N_A_1201_55#_c_904_n 0.0016556f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.645
cc_45 VNB N_A_1201_55#_c_905_n 0.0340515f $X=-0.19 $Y=-0.245 $X2=2.01 $Y2=1.415
cc_46 VNB N_A_1201_55#_c_906_n 0.0174151f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_1017_81#_c_987_n 0.0177343f $X=-0.19 $Y=-0.245 $X2=2.01 $Y2=0.58
cc_48 VNB N_A_1017_81#_c_988_n 0.0112637f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=1.495
cc_49 VNB N_A_1017_81#_c_989_n 0.0167979f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_1017_81#_c_990_n 0.0123419f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_1017_81#_c_991_n 0.0188668f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.645
cc_52 VNB N_A_1017_81#_c_992_n 0.0251433f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_1017_81#_c_993_n 0.00327901f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_1017_81#_c_994_n 0.0103511f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_1017_81#_c_995_n 0.0249608f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_1017_81#_c_996_n 0.0235339f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_1017_81#_c_997_n 0.00533446f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_1017_81#_c_998_n 0.00167982f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_1017_81#_c_999_n 0.0511294f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_1017_81#_c_1000_n 0.00339281f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_1017_81#_c_1001_n 0.064725f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_SET_B_M1003_g 0.0517031f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=2.245
cc_63 VNB N_SET_B_M1038_g 0.0527186f $X=-0.19 $Y=-0.245 $X2=1.88 $Y2=1.415
cc_64 VNB N_SET_B_c_1163_n 0.021194f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB SET_B 0.0011916f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.645
cc_66 VNB N_SET_B_c_1165_n 0.00146978f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_SET_B_c_1166_n 0.0227613f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_SET_B_c_1167_n 0.0193627f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_SET_B_c_1168_n 0.00417821f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_616_74#_M1021_g 0.0253006f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=2.64
cc_71 VNB N_A_616_74#_c_1305_n 0.0102921f $X=-0.19 $Y=-0.245 $X2=1.715 $Y2=1.495
cc_72 VNB N_A_616_74#_c_1306_n 0.0373616f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=1.495
cc_73 VNB N_A_616_74#_c_1307_n 0.0348939f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_616_74#_c_1308_n 0.00997874f $X=-0.19 $Y=-0.245 $X2=1.88 $Y2=1.495
cc_75 VNB N_A_616_74#_M1002_g 0.0255966f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.645
cc_76 VNB N_A_616_74#_c_1310_n 0.0419085f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_616_74#_c_1311_n 0.0143162f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_616_74#_M1026_g 0.0476321f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_616_74#_c_1313_n 0.00870938f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_616_74#_c_1314_n 0.0117023f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_616_74#_c_1315_n 0.00112234f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_616_74#_c_1316_n 0.00305136f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_2191_180#_c_1504_n 0.0237375f $X=-0.19 $Y=-0.245 $X2=0.945
+ $Y2=2.245
cc_84 VNB N_A_2191_180#_c_1505_n 0.026758f $X=-0.19 $Y=-0.245 $X2=1.715
+ $Y2=1.495
cc_85 VNB N_A_2191_180#_c_1506_n 0.0091707f $X=-0.19 $Y=-0.245 $X2=1.88
+ $Y2=1.415
cc_86 VNB N_A_2191_180#_c_1507_n 0.0078782f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_2191_180#_c_1508_n 0.00870653f $X=-0.19 $Y=-0.245 $X2=0.72
+ $Y2=1.58
cc_88 VNB N_A_2191_180#_c_1509_n 0.0312307f $X=-0.19 $Y=-0.245 $X2=1.88
+ $Y2=1.415
cc_89 VNB N_A_2191_180#_c_1510_n 0.00469145f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_2191_180#_c_1511_n 0.0185566f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_1823_524#_M1039_g 0.0527305f $X=-0.19 $Y=-0.245 $X2=1.88 $Y2=1.415
cc_92 VNB N_A_1823_524#_M1008_g 0.0477828f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_1823_524#_c_1612_n 0.00465656f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_1823_524#_c_1613_n 0.00597265f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_1823_524#_c_1614_n 0.00418558f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_1823_524#_c_1615_n 0.0113657f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_1823_524#_c_1616_n 0.0111225f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_A_1823_524#_c_1617_n 0.00183274f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_A_1823_524#_c_1618_n 0.00106587f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_A_1823_524#_c_1619_n 0.00199125f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_A_1823_524#_c_1620_n 0.0448785f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_A_2580_74#_M1000_g 0.0245919f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=2.64
cc_103 VNB N_A_2580_74#_M1015_g 0.0240442f $X=-0.19 $Y=-0.245 $X2=0.855
+ $Y2=1.495
cc_104 VNB N_A_2580_74#_M1023_g 0.0219865f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_105 VNB N_A_2580_74#_c_1829_n 0.0085538f $X=-0.19 $Y=-0.245 $X2=0.69
+ $Y2=1.645
cc_106 VNB N_A_2580_74#_c_1830_n 0.0866428f $X=-0.19 $Y=-0.245 $X2=1.88
+ $Y2=1.415
cc_107 VNB N_A_2580_74#_M1027_g 0.0271852f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_A_2580_74#_c_1832_n 0.0110307f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_A_2580_74#_c_1833_n 0.0098689f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_A_2580_74#_c_1834_n 0.0113182f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_A_2580_74#_c_1835_n 2.17078e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_A_2580_74#_c_1836_n 0.00847829f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_A_2580_74#_c_1837_n 0.00989086f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_VPWR_c_1947_n 0.661241f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_A_288_464#_c_2161_n 0.00125762f $X=-0.19 $Y=-0.245 $X2=1.88
+ $Y2=1.415
cc_116 VNB N_A_288_464#_c_2162_n 0.0133432f $X=-0.19 $Y=-0.245 $X2=1.88
+ $Y2=1.415
cc_117 VNB N_A_288_464#_c_2163_n 0.00269445f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_A_288_464#_c_2164_n 0.00627521f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_A_288_464#_c_2165_n 0.00576506f $X=-0.19 $Y=-0.245 $X2=0.69
+ $Y2=1.645
cc_120 VNB N_A_288_464#_c_2166_n 0.00759569f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_Q_c_2330_n 0.00328157f $X=-0.19 $Y=-0.245 $X2=1.715 $Y2=1.495
cc_122 VNB N_Q_c_2331_n 0.00353042f $X=-0.19 $Y=-0.245 $X2=1.88 $Y2=1.495
cc_123 VNB N_Q_c_2332_n 0.00283061f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_Q_c_2333_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.645
cc_125 VNB N_Q_c_2334_n 7.02455e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_Q_c_2335_n 0.012186f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_Q_c_2336_n 0.00132987f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB Q 0.00825292f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_Q_c_2338_n 0.00224342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_2414_n 0.0098348f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_2415_n 0.0105594f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_VGND_c_2416_n 0.0217656f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_VGND_c_2417_n 0.00641543f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_VGND_c_2418_n 0.0121589f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_VGND_c_2419_n 0.00858618f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_VGND_c_2420_n 0.0108564f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_VGND_c_2421_n 0.00826914f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB N_VGND_c_2422_n 0.00957908f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VNB N_VGND_c_2423_n 0.00571618f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_VGND_c_2424_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_141 VNB N_VGND_c_2425_n 0.041823f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_142 VNB N_VGND_c_2426_n 0.0334841f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_143 VNB N_VGND_c_2427_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_144 VNB N_VGND_c_2428_n 0.0190734f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_145 VNB N_VGND_c_2429_n 0.0443033f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_146 VNB N_VGND_c_2430_n 0.0611603f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_147 VNB N_VGND_c_2431_n 0.0306291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_148 VNB N_VGND_c_2432_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_149 VNB N_VGND_c_2433_n 0.068796f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_150 VNB N_VGND_c_2434_n 0.0188561f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_151 VNB N_VGND_c_2435_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_152 VNB N_VGND_c_2436_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_153 VNB N_VGND_c_2437_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_154 VNB N_VGND_c_2438_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_155 VNB N_VGND_c_2439_n 0.00632182f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_156 VNB N_VGND_c_2440_n 0.0125082f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_157 VNB N_VGND_c_2441_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_158 VNB N_VGND_c_2442_n 0.00942782f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_159 VNB N_VGND_c_2443_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_160 VNB N_VGND_c_2444_n 0.878417f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_161 VNB N_A_1677_74#_c_2590_n 0.00313319f $X=-0.19 $Y=-0.245 $X2=0.945
+ $Y2=2.64
cc_162 VNB N_A_1677_74#_c_2591_n 0.0200036f $X=-0.19 $Y=-0.245 $X2=2.01 $Y2=1.25
cc_163 VNB N_A_1677_74#_c_2592_n 5.50194e-19 $X=-0.19 $Y=-0.245 $X2=2.01
+ $Y2=0.58
cc_164 VNB N_A_1677_74#_c_2593_n 0.00110774f $X=-0.19 $Y=-0.245 $X2=1.715
+ $Y2=1.495
cc_165 VPB N_SCE_c_346_n 0.0184724f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.245
cc_166 VPB N_SCE_c_347_n 0.0151594f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=2.245
cc_167 VPB SCE 0.00252604f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_168 VPB N_SCE_c_344_n 0.0736647f $X=-0.19 $Y=1.66 $X2=0.69 $Y2=1.645
cc_169 VPB N_A_27_74#_c_423_n 0.0547416f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=2.64
cc_170 VPB N_A_27_74#_c_418_n 0.033356f $X=-0.19 $Y=1.66 $X2=1.88 $Y2=1.415
cc_171 VPB N_A_27_74#_c_425_n 0.00371646f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_172 VPB N_A_27_74#_c_426_n 0.0276635f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_173 VPB N_D_c_492_n 0.0509057f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.48
cc_174 VPB N_D_M1042_g 0.0134326f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.64
cc_175 VPB N_D_c_494_n 0.00717623f $X=-0.19 $Y=1.66 $X2=2.01 $Y2=0.58
cc_176 VPB N_SCD_c_528_n 0.0204346f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.64
cc_177 VPB N_SCD_c_532_n 0.0626646f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.64
cc_178 VPB SCD 0.00427107f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=2.64
cc_179 VPB N_CLK_c_570_n 0.024646f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_180 VPB N_A_803_74#_c_622_n 0.0229899f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=2.245
cc_181 VPB N_A_803_74#_c_623_n 0.0209544f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=2.64
cc_182 VPB N_A_803_74#_c_603_n 0.00636183f $X=-0.19 $Y=1.66 $X2=2.01 $Y2=0.58
cc_183 VPB N_A_803_74#_c_625_n 0.0147617f $X=-0.19 $Y=1.66 $X2=2.01 $Y2=1.415
cc_184 VPB N_A_803_74#_c_626_n 0.0224245f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_185 VPB N_A_803_74#_c_610_n 0.00405686f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_186 VPB N_A_803_74#_c_628_n 0.0235721f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_187 VPB N_A_803_74#_c_615_n 0.00233121f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_188 VPB N_A_803_74#_c_630_n 0.00342798f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_189 VPB N_A_803_74#_c_631_n 0.0022219f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_190 VPB N_A_803_74#_c_632_n 0.0147183f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_191 VPB N_A_803_74#_c_633_n 0.00268235f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_192 VPB N_A_803_74#_c_634_n 0.00389685f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_193 VPB N_A_803_74#_c_635_n 0.00654961f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_194 VPB N_A_803_74#_c_636_n 5.47995e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_195 VPB N_A_803_74#_c_637_n 0.0102665f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_196 VPB N_A_803_74#_c_638_n 0.0147919f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_197 VPB N_A_803_74#_c_639_n 0.00779773f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_198 VPB N_A_803_74#_c_640_n 0.00154337f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_199 VPB N_A_803_74#_c_641_n 0.0344636f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_200 VPB N_A_803_74#_c_642_n 4.0899e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_201 VPB N_A_803_74#_c_643_n 0.00289013f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_202 VPB N_A_803_74#_c_618_n 0.00406864f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_203 VPB N_A_803_74#_c_619_n 0.018862f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_204 VPB N_A_803_74#_c_646_n 0.00420976f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_205 VPB N_A_803_74#_c_647_n 0.0376148f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_206 VPB N_A_803_74#_c_620_n 0.0119965f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_207 VPB N_A_1201_55#_c_907_n 0.0560942f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=2.64
cc_208 VPB N_A_1201_55#_c_901_n 0.00671929f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_209 VPB N_A_1201_55#_c_909_n 0.0162369f $X=-0.19 $Y=1.66 $X2=1.88 $Y2=1.415
cc_210 VPB N_A_1201_55#_c_910_n 0.00417007f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.58
cc_211 VPB N_A_1201_55#_c_911_n 0.00278009f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_212 VPB N_A_1017_81#_c_1002_n 0.0192476f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=2.245
cc_213 VPB N_A_1017_81#_c_1003_n 0.0216148f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=2.64
cc_214 VPB N_A_1017_81#_c_988_n 0.00185123f $X=-0.19 $Y=1.66 $X2=0.855 $Y2=1.495
cc_215 VPB N_A_1017_81#_c_1005_n 0.0197751f $X=-0.19 $Y=1.66 $X2=1.88 $Y2=1.415
cc_216 VPB N_A_1017_81#_c_990_n 0.00204908f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_217 VPB N_A_1017_81#_c_1007_n 0.0211174f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.58
cc_218 VPB N_A_1017_81#_c_993_n 0.0129792f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_219 VPB N_A_1017_81#_c_1009_n 0.00263488f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_220 VPB N_A_1017_81#_c_1010_n 0.00105507f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_221 VPB N_A_1017_81#_c_1011_n 0.00924191f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_222 VPB N_A_1017_81#_c_998_n 0.00139883f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_223 VPB N_SET_B_c_1169_n 0.0210478f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.58
cc_224 VPB N_SET_B_c_1170_n 0.0204031f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.58
cc_225 VPB N_SET_B_c_1171_n 0.0201693f $X=-0.19 $Y=1.66 $X2=2.01 $Y2=1.25
cc_226 VPB N_SET_B_c_1172_n 0.0148784f $X=-0.19 $Y=1.66 $X2=2.01 $Y2=0.58
cc_227 VPB N_SET_B_c_1173_n 0.0262679f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_228 VPB N_SET_B_c_1174_n 0.0198787f $X=-0.19 $Y=1.66 $X2=1.88 $Y2=1.495
cc_229 VPB N_SET_B_c_1163_n 0.021685f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_230 VPB N_SET_B_c_1176_n 0.0010787f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_231 VPB SET_B 0.00128963f $X=-0.19 $Y=1.66 $X2=0.69 $Y2=1.645
cc_232 VPB N_SET_B_c_1165_n 8.36861e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_233 VPB N_SET_B_c_1166_n 0.0175149f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_234 VPB N_SET_B_c_1168_n 0.00522473f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_235 VPB N_A_616_74#_c_1317_n 0.0153539f $X=-0.19 $Y=1.66 $X2=2.01 $Y2=1.25
cc_236 VPB N_A_616_74#_c_1306_n 0.0174886f $X=-0.19 $Y=1.66 $X2=0.855 $Y2=1.495
cc_237 VPB N_A_616_74#_c_1319_n 0.0153198f $X=-0.19 $Y=1.66 $X2=1.88 $Y2=1.415
cc_238 VPB N_A_616_74#_c_1320_n 0.0576823f $X=-0.19 $Y=1.66 $X2=1.88 $Y2=1.415
cc_239 VPB N_A_616_74#_c_1321_n 0.0651825f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_240 VPB N_A_616_74#_c_1322_n 0.0124023f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_241 VPB N_A_616_74#_c_1323_n 0.0148554f $X=-0.19 $Y=1.66 $X2=0.69 $Y2=1.645
cc_242 VPB N_A_616_74#_c_1324_n 0.279863f $X=-0.19 $Y=1.66 $X2=2.01 $Y2=1.415
cc_243 VPB N_A_616_74#_c_1325_n 0.018406f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_244 VPB N_A_616_74#_c_1326_n 0.0356022f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_245 VPB N_A_616_74#_c_1327_n 0.0185558f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_246 VPB N_A_616_74#_c_1328_n 0.00741659f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_247 VPB N_A_616_74#_M1030_g 0.00737632f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_248 VPB N_A_616_74#_c_1311_n 0.00182704f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_249 VPB N_A_616_74#_c_1331_n 0.0136753f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_250 VPB N_A_616_74#_c_1332_n 0.0180862f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_251 VPB N_A_616_74#_c_1333_n 0.0122239f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_252 VPB N_A_616_74#_c_1314_n 0.00348613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_253 VPB N_A_616_74#_c_1335_n 0.013182f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_254 VPB N_A_616_74#_c_1336_n 0.00396556f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_255 VPB N_A_616_74#_c_1315_n 8.77165e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_256 VPB N_A_2191_180#_c_1504_n 0.0382593f $X=-0.19 $Y=1.66 $X2=0.945
+ $Y2=2.245
cc_257 VPB N_A_2191_180#_c_1513_n 0.0219836f $X=-0.19 $Y=1.66 $X2=2.01 $Y2=0.58
cc_258 VPB N_A_2191_180#_c_1514_n 0.00214288f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_259 VPB N_A_2191_180#_c_1507_n 0.00327448f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_260 VPB N_A_2191_180#_c_1516_n 0.00583651f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_261 VPB N_A_2191_180#_c_1517_n 0.00494054f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_262 VPB N_A_1823_524#_c_1621_n 0.0207651f $X=-0.19 $Y=1.66 $X2=1.88 $Y2=1.495
cc_263 VPB N_A_1823_524#_c_1622_n 0.0272898f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_264 VPB N_A_1823_524#_c_1623_n 0.0239104f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.58
cc_265 VPB N_A_1823_524#_c_1624_n 0.0154364f $X=-0.19 $Y=1.66 $X2=0.69 $Y2=1.645
cc_266 VPB N_A_1823_524#_M1008_g 0.0135742f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_267 VPB N_A_1823_524#_c_1626_n 0.0154743f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_268 VPB N_A_1823_524#_c_1627_n 0.036786f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_269 VPB N_A_1823_524#_c_1628_n 0.00408783f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_270 VPB N_A_1823_524#_c_1629_n 0.00866228f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_271 VPB N_A_1823_524#_c_1630_n 9.06755e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_272 VPB N_A_1823_524#_c_1618_n 0.00625106f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_273 VPB N_A_1823_524#_c_1632_n 0.00776284f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_274 VPB N_A_1823_524#_c_1633_n 0.00860505f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_275 VPB N_A_1823_524#_c_1620_n 0.0473428f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_276 VPB N_A_1823_524#_c_1635_n 0.00559393f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_277 VPB N_A_1823_524#_c_1636_n 0.00596772f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_278 VPB N_A_1823_524#_c_1637_n 8.90709e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_279 VPB N_A_1823_524#_c_1638_n 0.0164557f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_280 VPB N_A_2580_74#_c_1838_n 0.0167004f $X=-0.19 $Y=1.66 $X2=2.01 $Y2=1.25
cc_281 VPB N_A_2580_74#_c_1839_n 0.014884f $X=-0.19 $Y=1.66 $X2=1.88 $Y2=1.415
cc_282 VPB N_A_2580_74#_c_1840_n 0.0148648f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.58
cc_283 VPB N_A_2580_74#_c_1830_n 0.0205499f $X=-0.19 $Y=1.66 $X2=1.88 $Y2=1.415
cc_284 VPB N_A_2580_74#_c_1832_n 8.48304e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_285 VPB N_A_2580_74#_c_1843_n 0.0250879f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_286 VPB N_A_2580_74#_c_1835_n 0.00870003f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_287 VPB N_VPWR_c_1948_n 0.00396467f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_288 VPB N_VPWR_c_1949_n 0.0107937f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_289 VPB N_VPWR_c_1950_n 0.0202345f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_290 VPB N_VPWR_c_1951_n 0.00396467f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_291 VPB N_VPWR_c_1952_n 0.00579541f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_292 VPB N_VPWR_c_1953_n 0.0095436f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_293 VPB N_VPWR_c_1954_n 0.0111943f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_294 VPB N_VPWR_c_1955_n 0.00571271f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_295 VPB N_VPWR_c_1956_n 0.00499983f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_296 VPB N_VPWR_c_1957_n 0.00628728f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_297 VPB N_VPWR_c_1958_n 0.00268828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_298 VPB N_VPWR_c_1959_n 0.0120106f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_299 VPB N_VPWR_c_1960_n 0.0482331f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_300 VPB N_VPWR_c_1961_n 0.0278712f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_301 VPB N_VPWR_c_1962_n 0.00223798f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_302 VPB N_VPWR_c_1963_n 0.0172393f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_303 VPB N_VPWR_c_1964_n 0.00436868f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_304 VPB N_VPWR_c_1965_n 0.0177091f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_305 VPB N_VPWR_c_1966_n 0.0458211f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_306 VPB N_VPWR_c_1967_n 0.0581f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_307 VPB N_VPWR_c_1968_n 0.055019f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_308 VPB N_VPWR_c_1969_n 0.036934f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_309 VPB N_VPWR_c_1970_n 0.0164465f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_310 VPB N_VPWR_c_1971_n 0.0174954f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_311 VPB N_VPWR_c_1972_n 0.0164337f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_312 VPB N_VPWR_c_1973_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_313 VPB N_VPWR_c_1974_n 0.00631651f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_314 VPB N_VPWR_c_1975_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_315 VPB N_VPWR_c_1976_n 0.00330333f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_316 VPB N_VPWR_c_1977_n 0.00460249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_317 VPB N_VPWR_c_1978_n 0.00460249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_318 VPB N_VPWR_c_1979_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_319 VPB N_VPWR_c_1980_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_320 VPB N_VPWR_c_1947_n 0.116047f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_321 VPB N_A_288_464#_c_2164_n 0.00852439f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_322 VPB N_A_288_464#_c_2168_n 0.00754889f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_323 VPB N_A_288_464#_c_2169_n 0.00236749f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.58
cc_324 VPB N_A_288_464#_c_2165_n 0.00230536f $X=-0.19 $Y=1.66 $X2=0.69 $Y2=1.645
cc_325 VPB N_A_288_464#_c_2171_n 0.00818704f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_326 VPB N_A_288_464#_c_2172_n 0.0164949f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_327 VPB N_A_1620_373#_c_2289_n 0.0023794f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=2.64
cc_328 VPB N_A_1620_373#_c_2290_n 0.0135101f $X=-0.19 $Y=1.66 $X2=2.01 $Y2=1.25
cc_329 VPB N_A_1620_373#_c_2291_n 0.0024493f $X=-0.19 $Y=1.66 $X2=1.88 $Y2=1.415
cc_330 VPB A_2103_508# 0.00396022f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.48
cc_331 VPB N_Q_c_2339_n 0.0016237f $X=-0.19 $Y=1.66 $X2=1.88 $Y2=1.415
cc_332 VPB N_Q_c_2340_n 0.00243101f $X=-0.19 $Y=1.66 $X2=1.88 $Y2=1.415
cc_333 VPB N_Q_c_2341_n 0.00296149f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_334 VPB N_Q_c_2342_n 0.00180921f $X=-0.19 $Y=1.66 $X2=2.01 $Y2=1.415
cc_335 VPB N_Q_c_2334_n 0.0028771f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_336 VPB N_Q_c_2336_n 0.00223834f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_337 VPB N_Q_c_2338_n 0.00752918f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_338 N_SCE_c_343_n N_A_27_74#_c_423_n 3.29655e-19 $X=1.88 $Y=1.415 $X2=0 $Y2=0
cc_339 N_SCE_c_345_n N_A_27_74#_c_423_n 0.0164827f $X=2.01 $Y=1.415 $X2=0 $Y2=0
cc_340 N_SCE_M1045_g N_A_27_74#_c_417_n 0.0110711f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_341 N_SCE_M1045_g N_A_27_74#_c_418_n 0.00832591f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_342 N_SCE_c_346_n N_A_27_74#_c_418_n 0.00295538f $X=0.495 $Y=2.245 $X2=0
+ $Y2=0
cc_343 N_SCE_c_342_n N_A_27_74#_c_418_n 0.0139292f $X=0.855 $Y=1.495 $X2=0 $Y2=0
cc_344 SCE N_A_27_74#_c_418_n 0.0440891f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_345 N_SCE_c_344_n N_A_27_74#_c_418_n 0.0237634f $X=0.69 $Y=1.645 $X2=0 $Y2=0
cc_346 N_SCE_c_346_n N_A_27_74#_c_435_n 0.0130372f $X=0.495 $Y=2.245 $X2=0 $Y2=0
cc_347 N_SCE_c_347_n N_A_27_74#_c_435_n 0.0163062f $X=0.945 $Y=2.245 $X2=0 $Y2=0
cc_348 SCE N_A_27_74#_c_435_n 0.0220993f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_349 N_SCE_c_344_n N_A_27_74#_c_435_n 0.0016922f $X=0.69 $Y=1.645 $X2=0 $Y2=0
cc_350 N_SCE_M1045_g N_A_27_74#_c_419_n 0.0172929f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_351 N_SCE_c_341_n N_A_27_74#_c_419_n 0.021382f $X=1.715 $Y=1.495 $X2=0 $Y2=0
cc_352 N_SCE_c_342_n N_A_27_74#_c_419_n 0.0286153f $X=0.855 $Y=1.495 $X2=0 $Y2=0
cc_353 N_SCE_c_344_n N_A_27_74#_c_419_n 0.0016773f $X=0.69 $Y=1.645 $X2=0 $Y2=0
cc_354 N_SCE_M1045_g N_A_27_74#_c_420_n 0.0180926f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_355 N_SCE_c_341_n N_A_27_74#_c_420_n 0.00431973f $X=1.715 $Y=1.495 $X2=0
+ $Y2=0
cc_356 N_SCE_c_342_n N_A_27_74#_c_420_n 2.93992e-19 $X=0.855 $Y=1.495 $X2=0
+ $Y2=0
cc_357 N_SCE_c_344_n N_A_27_74#_c_420_n 0.0104595f $X=0.69 $Y=1.645 $X2=0 $Y2=0
cc_358 N_SCE_c_343_n N_A_27_74#_c_425_n 0.0151292f $X=1.88 $Y=1.415 $X2=0 $Y2=0
cc_359 N_SCE_c_345_n N_A_27_74#_c_425_n 3.27047e-19 $X=2.01 $Y=1.415 $X2=0 $Y2=0
cc_360 N_SCE_M1045_g N_A_27_74#_c_421_n 0.00879173f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_361 N_SCE_c_344_n N_A_27_74#_c_421_n 6.73206e-19 $X=0.69 $Y=1.645 $X2=0 $Y2=0
cc_362 N_SCE_c_346_n N_A_27_74#_c_426_n 0.00507302f $X=0.495 $Y=2.245 $X2=0
+ $Y2=0
cc_363 N_SCE_M1045_g N_A_27_74#_c_422_n 0.0122777f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_364 N_SCE_c_347_n N_D_c_492_n 0.0400037f $X=0.945 $Y=2.245 $X2=-0.19
+ $Y2=-0.245
cc_365 N_SCE_c_341_n N_D_c_492_n 0.0040855f $X=1.715 $Y=1.495 $X2=-0.19
+ $Y2=-0.245
cc_366 SCE N_D_c_492_n 2.62595e-19 $X=0.635 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_367 N_SCE_c_344_n N_D_c_492_n 0.0252607f $X=0.69 $Y=1.645 $X2=-0.19
+ $Y2=-0.245
cc_368 N_SCE_M1017_g N_D_M1042_g 0.0271445f $X=2.01 $Y=0.58 $X2=0 $Y2=0
cc_369 N_SCE_c_341_n N_D_M1042_g 0.0156564f $X=1.715 $Y=1.495 $X2=0 $Y2=0
cc_370 N_SCE_c_343_n N_D_M1042_g 0.00117677f $X=1.88 $Y=1.415 $X2=0 $Y2=0
cc_371 SCE N_D_M1042_g 0.00108399f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_372 N_SCE_c_344_n N_D_M1042_g 0.013509f $X=0.69 $Y=1.645 $X2=0 $Y2=0
cc_373 N_SCE_c_345_n N_D_M1042_g 0.0208078f $X=2.01 $Y=1.415 $X2=0 $Y2=0
cc_374 N_SCE_c_341_n N_D_c_494_n 0.0273112f $X=1.715 $Y=1.495 $X2=0 $Y2=0
cc_375 SCE N_D_c_494_n 0.0201046f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_376 N_SCE_c_344_n N_D_c_494_n 0.00300344f $X=0.69 $Y=1.645 $X2=0 $Y2=0
cc_377 N_SCE_M1017_g N_SCD_M1018_g 0.0346554f $X=2.01 $Y=0.58 $X2=0 $Y2=0
cc_378 N_SCE_c_343_n N_SCD_c_530_n 3.16269e-19 $X=1.88 $Y=1.415 $X2=0 $Y2=0
cc_379 N_SCE_c_345_n N_SCD_c_530_n 0.0346554f $X=2.01 $Y=1.415 $X2=0 $Y2=0
cc_380 N_SCE_c_346_n N_VPWR_c_1948_n 0.0101271f $X=0.495 $Y=2.245 $X2=0 $Y2=0
cc_381 N_SCE_c_347_n N_VPWR_c_1948_n 0.00946621f $X=0.945 $Y=2.245 $X2=0 $Y2=0
cc_382 N_SCE_c_346_n N_VPWR_c_1965_n 0.00413917f $X=0.495 $Y=2.245 $X2=0 $Y2=0
cc_383 N_SCE_c_347_n N_VPWR_c_1966_n 0.00413917f $X=0.945 $Y=2.245 $X2=0 $Y2=0
cc_384 N_SCE_c_346_n N_VPWR_c_1947_n 0.00417966f $X=0.495 $Y=2.245 $X2=0 $Y2=0
cc_385 N_SCE_c_347_n N_VPWR_c_1947_n 0.00414311f $X=0.945 $Y=2.245 $X2=0 $Y2=0
cc_386 N_SCE_c_347_n N_A_288_464#_c_2173_n 7.12872e-19 $X=0.945 $Y=2.245 $X2=0
+ $Y2=0
cc_387 N_SCE_M1017_g N_A_288_464#_c_2161_n 0.00470829f $X=2.01 $Y=0.58 $X2=0
+ $Y2=0
cc_388 N_SCE_M1017_g N_A_288_464#_c_2162_n 0.0118354f $X=2.01 $Y=0.58 $X2=0
+ $Y2=0
cc_389 N_SCE_c_343_n N_A_288_464#_c_2162_n 0.00599602f $X=1.88 $Y=1.415 $X2=0
+ $Y2=0
cc_390 N_SCE_M1017_g N_A_288_464#_c_2163_n 0.00250448f $X=2.01 $Y=0.58 $X2=0
+ $Y2=0
cc_391 N_SCE_c_343_n N_A_288_464#_c_2163_n 0.0135249f $X=1.88 $Y=1.415 $X2=0
+ $Y2=0
cc_392 N_SCE_c_345_n N_A_288_464#_c_2163_n 0.00107899f $X=2.01 $Y=1.415 $X2=0
+ $Y2=0
cc_393 N_SCE_M1017_g N_A_288_464#_c_2164_n 0.00565285f $X=2.01 $Y=0.58 $X2=0
+ $Y2=0
cc_394 N_SCE_c_343_n N_A_288_464#_c_2164_n 0.0248004f $X=1.88 $Y=1.415 $X2=0
+ $Y2=0
cc_395 N_SCE_M1017_g N_A_288_464#_c_2182_n 0.0111806f $X=2.01 $Y=0.58 $X2=0
+ $Y2=0
cc_396 N_SCE_c_341_n N_A_288_464#_c_2182_n 0.00592824f $X=1.715 $Y=1.495 $X2=0
+ $Y2=0
cc_397 N_SCE_c_343_n N_A_288_464#_c_2182_n 0.00248464f $X=1.88 $Y=1.415 $X2=0
+ $Y2=0
cc_398 N_SCE_c_345_n N_A_288_464#_c_2182_n 4.42746e-19 $X=2.01 $Y=1.415 $X2=0
+ $Y2=0
cc_399 N_SCE_M1045_g N_VGND_c_2414_n 0.00543785f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_400 N_SCE_M1017_g N_VGND_c_2415_n 0.00179638f $X=2.01 $Y=0.58 $X2=0 $Y2=0
cc_401 N_SCE_M1045_g N_VGND_c_2428_n 0.00434272f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_402 N_SCE_M1017_g N_VGND_c_2429_n 0.00434485f $X=2.01 $Y=0.58 $X2=0 $Y2=0
cc_403 N_SCE_M1045_g N_VGND_c_2444_n 0.00824747f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_404 N_SCE_M1017_g N_VGND_c_2444_n 0.00818993f $X=2.01 $Y=0.58 $X2=0 $Y2=0
cc_405 N_A_27_74#_c_423_n N_D_c_492_n 0.0433856f $X=1.995 $Y=2.245 $X2=-0.19
+ $Y2=-0.245
cc_406 N_A_27_74#_c_435_n N_D_c_492_n 0.0153081f $X=1.785 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_407 N_A_27_74#_c_425_n N_D_c_492_n 0.00363007f $X=1.95 $Y=1.995 $X2=-0.19
+ $Y2=-0.245
cc_408 N_A_27_74#_c_419_n N_D_M1042_g 0.00172934f $X=0.975 $Y=1.075 $X2=0 $Y2=0
cc_409 N_A_27_74#_c_420_n N_D_M1042_g 0.0196496f $X=0.975 $Y=1.075 $X2=0 $Y2=0
cc_410 N_A_27_74#_c_422_n N_D_M1042_g 0.0348158f $X=0.975 $Y=0.91 $X2=0 $Y2=0
cc_411 N_A_27_74#_c_423_n N_D_c_494_n 0.00111089f $X=1.995 $Y=2.245 $X2=0 $Y2=0
cc_412 N_A_27_74#_c_435_n N_D_c_494_n 0.0307759f $X=1.785 $Y=2.405 $X2=0 $Y2=0
cc_413 N_A_27_74#_c_425_n N_D_c_494_n 0.0205002f $X=1.95 $Y=1.995 $X2=0 $Y2=0
cc_414 N_A_27_74#_c_423_n N_SCD_c_528_n 0.0204489f $X=1.995 $Y=2.245 $X2=0 $Y2=0
cc_415 N_A_27_74#_c_425_n N_SCD_c_528_n 3.79863e-19 $X=1.95 $Y=1.995 $X2=0 $Y2=0
cc_416 N_A_27_74#_c_423_n N_SCD_c_532_n 0.0422835f $X=1.995 $Y=2.245 $X2=0 $Y2=0
cc_417 N_A_27_74#_c_435_n N_VPWR_M1043_d 0.00350365f $X=1.785 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_418 N_A_27_74#_c_435_n N_VPWR_c_1948_n 0.0168032f $X=1.785 $Y=2.405 $X2=0
+ $Y2=0
cc_419 N_A_27_74#_c_426_n N_VPWR_c_1948_n 0.0214859f $X=0.27 $Y=2.465 $X2=0
+ $Y2=0
cc_420 N_A_27_74#_c_426_n N_VPWR_c_1965_n 0.011066f $X=0.27 $Y=2.465 $X2=0 $Y2=0
cc_421 N_A_27_74#_c_423_n N_VPWR_c_1966_n 0.00300876f $X=1.995 $Y=2.245 $X2=0
+ $Y2=0
cc_422 N_A_27_74#_c_423_n N_VPWR_c_1947_n 0.00370184f $X=1.995 $Y=2.245 $X2=0
+ $Y2=0
cc_423 N_A_27_74#_c_435_n N_VPWR_c_1947_n 0.0242263f $X=1.785 $Y=2.405 $X2=0
+ $Y2=0
cc_424 N_A_27_74#_c_426_n N_VPWR_c_1947_n 0.00915947f $X=0.27 $Y=2.465 $X2=0
+ $Y2=0
cc_425 N_A_27_74#_c_435_n A_204_464# 0.0055687f $X=1.785 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_426 N_A_27_74#_c_435_n N_A_288_464#_M1034_d 0.0134049f $X=1.785 $Y=2.405
+ $X2=0 $Y2=0
cc_427 N_A_27_74#_c_423_n N_A_288_464#_c_2173_n 0.0147338f $X=1.995 $Y=2.245
+ $X2=0 $Y2=0
cc_428 N_A_27_74#_c_435_n N_A_288_464#_c_2173_n 0.0377979f $X=1.785 $Y=2.405
+ $X2=0 $Y2=0
cc_429 N_A_27_74#_c_419_n N_A_288_464#_c_2163_n 0.00531239f $X=0.975 $Y=1.075
+ $X2=0 $Y2=0
cc_430 N_A_27_74#_c_423_n N_A_288_464#_c_2164_n 0.00750203f $X=1.995 $Y=2.245
+ $X2=0 $Y2=0
cc_431 N_A_27_74#_c_435_n N_A_288_464#_c_2164_n 0.0133253f $X=1.785 $Y=2.405
+ $X2=0 $Y2=0
cc_432 N_A_27_74#_c_425_n N_A_288_464#_c_2164_n 0.0360921f $X=1.95 $Y=1.995
+ $X2=0 $Y2=0
cc_433 N_A_27_74#_c_422_n N_A_288_464#_c_2182_n 9.45341e-19 $X=0.975 $Y=0.91
+ $X2=0 $Y2=0
cc_434 N_A_27_74#_c_423_n N_A_288_464#_c_2194_n 2.67314e-19 $X=1.995 $Y=2.245
+ $X2=0 $Y2=0
cc_435 N_A_27_74#_c_417_n N_VGND_c_2414_n 0.0154913f $X=0.28 $Y=0.58 $X2=0 $Y2=0
cc_436 N_A_27_74#_c_419_n N_VGND_c_2414_n 0.02555f $X=0.975 $Y=1.075 $X2=0 $Y2=0
cc_437 N_A_27_74#_c_420_n N_VGND_c_2414_n 0.00299669f $X=0.975 $Y=1.075 $X2=0
+ $Y2=0
cc_438 N_A_27_74#_c_422_n N_VGND_c_2414_n 0.0038508f $X=0.975 $Y=0.91 $X2=0
+ $Y2=0
cc_439 N_A_27_74#_c_417_n N_VGND_c_2428_n 0.0150101f $X=0.28 $Y=0.58 $X2=0 $Y2=0
cc_440 N_A_27_74#_c_422_n N_VGND_c_2429_n 0.00461464f $X=0.975 $Y=0.91 $X2=0
+ $Y2=0
cc_441 N_A_27_74#_c_417_n N_VGND_c_2444_n 0.0123677f $X=0.28 $Y=0.58 $X2=0 $Y2=0
cc_442 N_A_27_74#_c_422_n N_VGND_c_2444_n 0.00908175f $X=0.975 $Y=0.91 $X2=0
+ $Y2=0
cc_443 N_D_c_492_n N_VPWR_c_1948_n 0.0016042f $X=1.365 $Y=2.245 $X2=0 $Y2=0
cc_444 N_D_c_492_n N_VPWR_c_1966_n 0.00445405f $X=1.365 $Y=2.245 $X2=0 $Y2=0
cc_445 N_D_c_492_n N_VPWR_c_1947_n 0.00456649f $X=1.365 $Y=2.245 $X2=0 $Y2=0
cc_446 N_D_c_492_n N_A_288_464#_c_2173_n 0.00888514f $X=1.365 $Y=2.245 $X2=0
+ $Y2=0
cc_447 N_D_M1042_g N_A_288_464#_c_2161_n 0.0032439f $X=1.425 $Y=0.58 $X2=0 $Y2=0
cc_448 N_D_M1042_g N_A_288_464#_c_2163_n 0.00195305f $X=1.425 $Y=0.58 $X2=0
+ $Y2=0
cc_449 N_D_c_494_n N_A_288_464#_c_2164_n 2.53081e-19 $X=1.41 $Y=1.985 $X2=0
+ $Y2=0
cc_450 N_D_M1042_g N_A_288_464#_c_2182_n 0.0120673f $X=1.425 $Y=0.58 $X2=0 $Y2=0
cc_451 N_D_M1042_g N_VGND_c_2429_n 0.00434485f $X=1.425 $Y=0.58 $X2=0 $Y2=0
cc_452 N_D_M1042_g N_VGND_c_2444_n 0.00819992f $X=1.425 $Y=0.58 $X2=0 $Y2=0
cc_453 N_SCD_c_530_n N_CLK_c_569_n 0.00195011f $X=2.695 $Y=1.265 $X2=-0.19
+ $Y2=-0.245
cc_454 N_SCD_c_528_n N_CLK_c_570_n 0.00634023f $X=2.592 $Y=1.843 $X2=0 $Y2=0
cc_455 N_SCD_c_530_n N_CLK_c_570_n 0.00642894f $X=2.695 $Y=1.265 $X2=0 $Y2=0
cc_456 N_SCD_M1018_g N_A_616_74#_c_1313_n 0.00807309f $X=2.4 $Y=0.58 $X2=0 $Y2=0
cc_457 SCD N_A_616_74#_c_1314_n 0.0533653f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_458 N_SCD_c_530_n N_A_616_74#_c_1314_n 0.00726202f $X=2.695 $Y=1.265 $X2=0
+ $Y2=0
cc_459 N_SCD_c_528_n N_A_616_74#_c_1336_n 0.00294822f $X=2.592 $Y=1.843 $X2=0
+ $Y2=0
cc_460 SCD N_A_616_74#_c_1336_n 0.0208115f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_461 N_SCD_c_532_n N_VPWR_c_1949_n 0.00917244f $X=2.415 $Y=2.245 $X2=0 $Y2=0
cc_462 N_SCD_c_532_n N_VPWR_c_1966_n 0.00322244f $X=2.415 $Y=2.245 $X2=0 $Y2=0
cc_463 N_SCD_c_532_n N_VPWR_c_1947_n 0.00409406f $X=2.415 $Y=2.245 $X2=0 $Y2=0
cc_464 N_SCD_c_532_n N_A_288_464#_c_2173_n 2.98199e-19 $X=2.415 $Y=2.245 $X2=0
+ $Y2=0
cc_465 N_SCD_M1018_g N_A_288_464#_c_2161_n 8.48135e-19 $X=2.4 $Y=0.58 $X2=0
+ $Y2=0
cc_466 N_SCD_M1018_g N_A_288_464#_c_2162_n 0.00879847f $X=2.4 $Y=0.58 $X2=0
+ $Y2=0
cc_467 N_SCD_M1018_g N_A_288_464#_c_2164_n 5.26815e-19 $X=2.4 $Y=0.58 $X2=0
+ $Y2=0
cc_468 N_SCD_c_528_n N_A_288_464#_c_2164_n 0.014425f $X=2.592 $Y=1.843 $X2=0
+ $Y2=0
cc_469 N_SCD_c_532_n N_A_288_464#_c_2164_n 0.0191424f $X=2.415 $Y=2.245 $X2=0
+ $Y2=0
cc_470 SCD N_A_288_464#_c_2164_n 0.0740228f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_471 N_SCD_c_530_n N_A_288_464#_c_2164_n 0.00657468f $X=2.695 $Y=1.265 $X2=0
+ $Y2=0
cc_472 N_SCD_c_532_n N_A_288_464#_c_2168_n 0.016511f $X=2.415 $Y=2.245 $X2=0
+ $Y2=0
cc_473 SCD N_A_288_464#_c_2168_n 0.0140907f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_474 N_SCD_M1018_g N_A_288_464#_c_2182_n 9.27271e-19 $X=2.4 $Y=0.58 $X2=0
+ $Y2=0
cc_475 N_SCD_c_532_n N_A_288_464#_c_2194_n 0.0126627f $X=2.415 $Y=2.245 $X2=0
+ $Y2=0
cc_476 N_SCD_c_532_n N_A_288_464#_c_2171_n 0.00425835f $X=2.415 $Y=2.245 $X2=0
+ $Y2=0
cc_477 N_SCD_M1018_g N_VGND_c_2415_n 0.0127827f $X=2.4 $Y=0.58 $X2=0 $Y2=0
cc_478 SCD N_VGND_c_2415_n 0.0109414f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_479 N_SCD_c_530_n N_VGND_c_2415_n 0.00366449f $X=2.695 $Y=1.265 $X2=0 $Y2=0
cc_480 N_SCD_M1018_g N_VGND_c_2429_n 0.00383152f $X=2.4 $Y=0.58 $X2=0 $Y2=0
cc_481 N_SCD_M1018_g N_VGND_c_2444_n 0.0075725f $X=2.4 $Y=0.58 $X2=0 $Y2=0
cc_482 N_CLK_c_569_n N_A_616_74#_M1021_g 0.0175852f $X=3.44 $Y=1.22 $X2=0 $Y2=0
cc_483 N_CLK_c_570_n N_A_616_74#_M1021_g 0.020775f $X=3.51 $Y=1.765 $X2=0 $Y2=0
cc_484 CLK N_A_616_74#_M1021_g 0.00539117f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_485 N_CLK_c_570_n N_A_616_74#_c_1317_n 0.0413548f $X=3.51 $Y=1.765 $X2=0
+ $Y2=0
cc_486 N_CLK_c_570_n N_A_616_74#_c_1306_n 0.0104637f $X=3.51 $Y=1.765 $X2=0
+ $Y2=0
cc_487 N_CLK_c_569_n N_A_616_74#_c_1313_n 0.00583023f $X=3.44 $Y=1.22 $X2=0
+ $Y2=0
cc_488 N_CLK_c_569_n N_A_616_74#_c_1314_n 0.00340241f $X=3.44 $Y=1.22 $X2=0
+ $Y2=0
cc_489 N_CLK_c_570_n N_A_616_74#_c_1314_n 0.00863617f $X=3.51 $Y=1.765 $X2=0
+ $Y2=0
cc_490 CLK N_A_616_74#_c_1314_n 0.0282001f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_491 N_CLK_c_570_n N_A_616_74#_c_1335_n 0.0161956f $X=3.51 $Y=1.765 $X2=0
+ $Y2=0
cc_492 CLK N_A_616_74#_c_1335_n 0.0201123f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_493 N_CLK_c_570_n N_A_616_74#_c_1315_n 0.00187439f $X=3.51 $Y=1.765 $X2=0
+ $Y2=0
cc_494 CLK N_A_616_74#_c_1315_n 0.0159704f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_495 N_CLK_c_569_n N_A_616_74#_c_1316_n 0.00229489f $X=3.44 $Y=1.22 $X2=0
+ $Y2=0
cc_496 CLK N_A_616_74#_c_1316_n 0.00273603f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_497 N_CLK_c_570_n N_VPWR_c_1949_n 0.00646829f $X=3.51 $Y=1.765 $X2=0 $Y2=0
cc_498 N_CLK_c_570_n N_VPWR_c_1950_n 0.00413917f $X=3.51 $Y=1.765 $X2=0 $Y2=0
cc_499 N_CLK_c_570_n N_VPWR_c_1951_n 0.021577f $X=3.51 $Y=1.765 $X2=0 $Y2=0
cc_500 N_CLK_c_570_n N_VPWR_c_1947_n 0.00822528f $X=3.51 $Y=1.765 $X2=0 $Y2=0
cc_501 N_CLK_c_570_n N_A_288_464#_c_2169_n 0.01598f $X=3.51 $Y=1.765 $X2=0 $Y2=0
cc_502 N_CLK_c_570_n N_A_288_464#_c_2171_n 0.00750031f $X=3.51 $Y=1.765 $X2=0
+ $Y2=0
cc_503 N_CLK_c_569_n N_VGND_c_2415_n 0.00328908f $X=3.44 $Y=1.22 $X2=0 $Y2=0
cc_504 N_CLK_c_569_n N_VGND_c_2416_n 0.00434272f $X=3.44 $Y=1.22 $X2=0 $Y2=0
cc_505 N_CLK_c_569_n N_VGND_c_2417_n 0.00659657f $X=3.44 $Y=1.22 $X2=0 $Y2=0
cc_506 N_CLK_c_570_n N_VGND_c_2417_n 6.35135e-19 $X=3.51 $Y=1.765 $X2=0 $Y2=0
cc_507 CLK N_VGND_c_2417_n 0.0129689f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_508 N_CLK_c_569_n N_VGND_c_2444_n 0.00825771f $X=3.44 $Y=1.22 $X2=0 $Y2=0
cc_509 N_A_803_74#_c_630_n N_A_1201_55#_c_907_n 0.00586266f $X=5.745 $Y=2.29
+ $X2=0 $Y2=0
cc_510 N_A_803_74#_c_650_p N_A_1201_55#_c_907_n 0.00510269f $X=5.745 $Y=2.895
+ $X2=0 $Y2=0
cc_511 N_A_803_74#_c_651_p N_A_1201_55#_c_907_n 0.0141646f $X=6.695 $Y=2.375
+ $X2=0 $Y2=0
cc_512 N_A_803_74#_c_631_n N_A_1201_55#_c_907_n 0.00295016f $X=6.78 $Y=2.895
+ $X2=0 $Y2=0
cc_513 N_A_803_74#_c_640_n N_A_1201_55#_c_907_n 0.00113262f $X=5.665 $Y=1.94
+ $X2=0 $Y2=0
cc_514 N_A_803_74#_c_641_n N_A_1201_55#_c_907_n 0.0198057f $X=5.665 $Y=1.94
+ $X2=0 $Y2=0
cc_515 N_A_803_74#_M1020_g N_A_1201_55#_c_901_n 0.00882513f $X=5.69 $Y=0.615
+ $X2=0 $Y2=0
cc_516 N_A_803_74#_c_610_n N_A_1201_55#_c_901_n 0.0087626f $X=5.665 $Y=1.655
+ $X2=0 $Y2=0
cc_517 N_A_803_74#_c_651_p N_A_1201_55#_c_909_n 0.034957f $X=6.695 $Y=2.375
+ $X2=0 $Y2=0
cc_518 N_A_803_74#_c_636_n N_A_1201_55#_c_909_n 0.0144283f $X=7.545 $Y=2.035
+ $X2=0 $Y2=0
cc_519 N_A_803_74#_c_651_p N_A_1201_55#_c_910_n 0.0133617f $X=6.695 $Y=2.375
+ $X2=0 $Y2=0
cc_520 N_A_803_74#_c_631_n N_A_1201_55#_c_910_n 0.0185965f $X=6.78 $Y=2.895
+ $X2=0 $Y2=0
cc_521 N_A_803_74#_c_632_n N_A_1201_55#_c_910_n 0.0133013f $X=7.375 $Y=2.98
+ $X2=0 $Y2=0
cc_522 N_A_803_74#_c_634_n N_A_1201_55#_c_910_n 0.0426105f $X=7.46 $Y=2.895
+ $X2=0 $Y2=0
cc_523 N_A_803_74#_M1020_g N_A_1201_55#_c_904_n 0.00171735f $X=5.69 $Y=0.615
+ $X2=0 $Y2=0
cc_524 N_A_803_74#_c_651_p N_A_1201_55#_c_911_n 0.0220592f $X=6.695 $Y=2.375
+ $X2=0 $Y2=0
cc_525 N_A_803_74#_c_640_n N_A_1201_55#_c_911_n 0.0213242f $X=5.665 $Y=1.94
+ $X2=0 $Y2=0
cc_526 N_A_803_74#_c_641_n N_A_1201_55#_c_911_n 0.00113194f $X=5.665 $Y=1.94
+ $X2=0 $Y2=0
cc_527 N_A_803_74#_M1020_g N_A_1201_55#_c_906_n 0.0499897f $X=5.69 $Y=0.615
+ $X2=0 $Y2=0
cc_528 N_A_803_74#_c_651_p N_A_1017_81#_c_1003_n 0.00665677f $X=6.695 $Y=2.375
+ $X2=0 $Y2=0
cc_529 N_A_803_74#_c_631_n N_A_1017_81#_c_1003_n 0.0107045f $X=6.78 $Y=2.895
+ $X2=0 $Y2=0
cc_530 N_A_803_74#_c_632_n N_A_1017_81#_c_1003_n 0.00220266f $X=7.375 $Y=2.98
+ $X2=0 $Y2=0
cc_531 N_A_803_74#_c_634_n N_A_1017_81#_c_1003_n 4.76836e-19 $X=7.46 $Y=2.895
+ $X2=0 $Y2=0
cc_532 N_A_803_74#_c_634_n N_A_1017_81#_c_1005_n 0.00207205f $X=7.46 $Y=2.895
+ $X2=0 $Y2=0
cc_533 N_A_803_74#_c_637_n N_A_1017_81#_c_1005_n 0.0159292f $X=9.045 $Y=1.865
+ $X2=0 $Y2=0
cc_534 N_A_803_74#_c_643_n N_A_1017_81#_c_1005_n 5.52576e-19 $X=7.81 $Y=1.865
+ $X2=0 $Y2=0
cc_535 N_A_803_74#_c_618_n N_A_1017_81#_c_990_n 0.00209777f $X=9.21 $Y=1.615
+ $X2=0 $Y2=0
cc_536 N_A_803_74#_c_619_n N_A_1017_81#_c_990_n 0.00901343f $X=9.21 $Y=1.615
+ $X2=0 $Y2=0
cc_537 N_A_803_74#_c_637_n N_A_1017_81#_c_1007_n 0.0142926f $X=9.045 $Y=1.865
+ $X2=0 $Y2=0
cc_538 N_A_803_74#_c_618_n N_A_1017_81#_c_1007_n 3.93494e-19 $X=9.21 $Y=1.615
+ $X2=0 $Y2=0
cc_539 N_A_803_74#_c_603_n N_A_1017_81#_c_1009_n 6.45562e-19 $X=5.5 $Y=1.655
+ $X2=0 $Y2=0
cc_540 N_A_803_74#_c_630_n N_A_1017_81#_c_1009_n 0.00109141f $X=5.745 $Y=2.29
+ $X2=0 $Y2=0
cc_541 N_A_803_74#_c_642_n N_A_1017_81#_c_1009_n 0.0137049f $X=5.745 $Y=2.375
+ $X2=0 $Y2=0
cc_542 N_A_803_74#_c_628_n N_A_1017_81#_c_1010_n 0.0214489f $X=5.66 $Y=2.98
+ $X2=0 $Y2=0
cc_543 N_A_803_74#_c_650_p N_A_1017_81#_c_1010_n 0.0185063f $X=5.745 $Y=2.895
+ $X2=0 $Y2=0
cc_544 N_A_803_74#_M1020_g N_A_1017_81#_c_994_n 0.0286052f $X=5.69 $Y=0.615
+ $X2=0 $Y2=0
cc_545 N_A_803_74#_c_613_n N_A_1017_81#_c_994_n 0.00252794f $X=4.97 $Y=0.34
+ $X2=0 $Y2=0
cc_546 N_A_803_74#_c_615_n N_A_1017_81#_c_994_n 0.00968151f $X=4.9 $Y=1.565
+ $X2=0 $Y2=0
cc_547 N_A_803_74#_c_616_n N_A_1017_81#_c_994_n 0.0517056f $X=4.945 $Y=1.095
+ $X2=0 $Y2=0
cc_548 N_A_803_74#_c_620_n N_A_1017_81#_c_994_n 3.84912e-19 $X=5.18 $Y=1.565
+ $X2=0 $Y2=0
cc_549 N_A_803_74#_M1020_g N_A_1017_81#_c_995_n 0.00941404f $X=5.69 $Y=0.615
+ $X2=0 $Y2=0
cc_550 N_A_803_74#_c_610_n N_A_1017_81#_c_995_n 0.00445914f $X=5.665 $Y=1.655
+ $X2=0 $Y2=0
cc_551 N_A_803_74#_c_640_n N_A_1017_81#_c_995_n 0.0142753f $X=5.665 $Y=1.94
+ $X2=0 $Y2=0
cc_552 N_A_803_74#_c_635_n N_A_1017_81#_c_996_n 0.00175651f $X=7.725 $Y=2.035
+ $X2=0 $Y2=0
cc_553 N_A_803_74#_c_637_n N_A_1017_81#_c_996_n 6.44876e-19 $X=9.045 $Y=1.865
+ $X2=0 $Y2=0
cc_554 N_A_803_74#_c_643_n N_A_1017_81#_c_996_n 0.00285102f $X=7.81 $Y=1.865
+ $X2=0 $Y2=0
cc_555 N_A_803_74#_c_603_n N_A_1017_81#_c_997_n 0.0114032f $X=5.5 $Y=1.655 $X2=0
+ $Y2=0
cc_556 N_A_803_74#_M1020_g N_A_1017_81#_c_997_n 0.0025116f $X=5.69 $Y=0.615
+ $X2=0 $Y2=0
cc_557 N_A_803_74#_c_610_n N_A_1017_81#_c_997_n 0.00662768f $X=5.665 $Y=1.655
+ $X2=0 $Y2=0
cc_558 N_A_803_74#_c_615_n N_A_1017_81#_c_997_n 0.0140626f $X=4.9 $Y=1.565 $X2=0
+ $Y2=0
cc_559 N_A_803_74#_c_640_n N_A_1017_81#_c_997_n 0.00794388f $X=5.665 $Y=1.94
+ $X2=0 $Y2=0
cc_560 N_A_803_74#_c_620_n N_A_1017_81#_c_997_n 0.00182765f $X=5.18 $Y=1.565
+ $X2=0 $Y2=0
cc_561 N_A_803_74#_c_622_n N_A_1017_81#_c_1011_n 0.00657969f $X=5.09 $Y=2.12
+ $X2=0 $Y2=0
cc_562 N_A_803_74#_c_623_n N_A_1017_81#_c_1011_n 0.0023445f $X=5.09 $Y=2.21
+ $X2=0 $Y2=0
cc_563 N_A_803_74#_c_603_n N_A_1017_81#_c_1011_n 0.00915303f $X=5.5 $Y=1.655
+ $X2=0 $Y2=0
cc_564 N_A_803_74#_c_615_n N_A_1017_81#_c_1011_n 0.00916981f $X=4.9 $Y=1.565
+ $X2=0 $Y2=0
cc_565 N_A_803_74#_c_630_n N_A_1017_81#_c_1011_n 0.00621153f $X=5.745 $Y=2.29
+ $X2=0 $Y2=0
cc_566 N_A_803_74#_c_640_n N_A_1017_81#_c_1011_n 0.0245577f $X=5.665 $Y=1.94
+ $X2=0 $Y2=0
cc_567 N_A_803_74#_c_641_n N_A_1017_81#_c_1011_n 0.0034199f $X=5.665 $Y=1.94
+ $X2=0 $Y2=0
cc_568 N_A_803_74#_c_637_n N_A_1017_81#_c_1000_n 0.00800314f $X=9.045 $Y=1.865
+ $X2=0 $Y2=0
cc_569 N_A_803_74#_c_606_n N_A_1017_81#_c_1001_n 0.00437955f $X=9.375 $Y=1.16
+ $X2=0 $Y2=0
cc_570 N_A_803_74#_c_637_n N_A_1017_81#_c_1001_n 0.00271175f $X=9.045 $Y=1.865
+ $X2=0 $Y2=0
cc_571 N_A_803_74#_c_621_n N_A_1017_81#_c_1001_n 0.00487076f $X=9.21 $Y=1.45
+ $X2=0 $Y2=0
cc_572 N_A_803_74#_c_636_n N_SET_B_c_1169_n 0.00554667f $X=7.545 $Y=2.035 $X2=0
+ $Y2=0
cc_573 N_A_803_74#_c_643_n N_SET_B_c_1169_n 0.00358031f $X=7.81 $Y=1.865 $X2=0
+ $Y2=0
cc_574 N_A_803_74#_c_631_n N_SET_B_c_1170_n 4.36583e-19 $X=6.78 $Y=2.895 $X2=0
+ $Y2=0
cc_575 N_A_803_74#_c_632_n N_SET_B_c_1170_n 0.00294494f $X=7.375 $Y=2.98 $X2=0
+ $Y2=0
cc_576 N_A_803_74#_c_634_n N_SET_B_c_1170_n 0.0180094f $X=7.46 $Y=2.895 $X2=0
+ $Y2=0
cc_577 N_A_803_74#_c_608_n N_SET_B_c_1163_n 9.08689e-19 $X=10.085 $Y=1.16 $X2=0
+ $Y2=0
cc_578 N_A_803_74#_c_635_n N_SET_B_c_1163_n 0.00408641f $X=7.725 $Y=2.035 $X2=0
+ $Y2=0
cc_579 N_A_803_74#_c_637_n N_SET_B_c_1163_n 0.0402396f $X=9.045 $Y=1.865 $X2=0
+ $Y2=0
cc_580 N_A_803_74#_c_638_n N_SET_B_c_1163_n 0.0385897f $X=10.435 $Y=1.845 $X2=0
+ $Y2=0
cc_581 N_A_803_74#_c_643_n N_SET_B_c_1163_n 0.00609828f $X=7.81 $Y=1.865 $X2=0
+ $Y2=0
cc_582 N_A_803_74#_c_618_n N_SET_B_c_1163_n 0.0218675f $X=9.21 $Y=1.615 $X2=0
+ $Y2=0
cc_583 N_A_803_74#_c_619_n N_SET_B_c_1163_n 0.00265151f $X=9.21 $Y=1.615 $X2=0
+ $Y2=0
cc_584 N_A_803_74#_c_646_n N_SET_B_c_1163_n 0.0101538f $X=10.6 $Y=1.845 $X2=0
+ $Y2=0
cc_585 N_A_803_74#_c_635_n N_SET_B_c_1176_n 0.00114052f $X=7.725 $Y=2.035 $X2=0
+ $Y2=0
cc_586 N_A_803_74#_c_636_n N_SET_B_c_1176_n 0.00414922f $X=7.545 $Y=2.035 $X2=0
+ $Y2=0
cc_587 N_A_803_74#_c_635_n N_SET_B_c_1165_n 6.00858e-19 $X=7.725 $Y=2.035 $X2=0
+ $Y2=0
cc_588 N_A_803_74#_c_636_n N_SET_B_c_1165_n 0.011802f $X=7.545 $Y=2.035 $X2=0
+ $Y2=0
cc_589 N_A_803_74#_c_635_n N_SET_B_c_1166_n 0.00182453f $X=7.725 $Y=2.035 $X2=0
+ $Y2=0
cc_590 N_A_803_74#_c_636_n N_SET_B_c_1166_n 0.0020884f $X=7.545 $Y=2.035 $X2=0
+ $Y2=0
cc_591 N_A_803_74#_c_612_n N_A_616_74#_M1021_g 0.00162741f $X=4.155 $Y=0.515
+ $X2=0 $Y2=0
cc_592 N_A_803_74#_c_614_n N_A_616_74#_M1021_g 0.00266901f $X=4.24 $Y=0.34 $X2=0
+ $Y2=0
cc_593 N_A_803_74#_c_639_n N_A_616_74#_c_1317_n 0.00335712f $X=4.235 $Y=2.78
+ $X2=0 $Y2=0
cc_594 N_A_803_74#_c_617_n N_A_616_74#_c_1305_n 6.69154e-19 $X=4.945 $Y=1.265
+ $X2=0 $Y2=0
cc_595 N_A_803_74#_c_612_n N_A_616_74#_c_1306_n 0.00188848f $X=4.155 $Y=0.515
+ $X2=0 $Y2=0
cc_596 N_A_803_74#_c_615_n N_A_616_74#_c_1306_n 0.00102684f $X=4.9 $Y=1.565
+ $X2=0 $Y2=0
cc_597 N_A_803_74#_c_620_n N_A_616_74#_c_1306_n 0.0214155f $X=5.18 $Y=1.565
+ $X2=0 $Y2=0
cc_598 N_A_803_74#_c_622_n N_A_616_74#_c_1319_n 0.00492463f $X=5.09 $Y=2.12
+ $X2=0 $Y2=0
cc_599 N_A_803_74#_c_623_n N_A_616_74#_c_1320_n 0.0142877f $X=5.09 $Y=2.21 $X2=0
+ $Y2=0
cc_600 N_A_803_74#_c_628_n N_A_616_74#_c_1320_n 0.0127037f $X=5.66 $Y=2.98 $X2=0
+ $Y2=0
cc_601 N_A_803_74#_c_639_n N_A_616_74#_c_1320_n 0.00704372f $X=4.235 $Y=2.78
+ $X2=0 $Y2=0
cc_602 N_A_803_74#_c_613_n N_A_616_74#_c_1307_n 0.00190744f $X=4.97 $Y=0.34
+ $X2=0 $Y2=0
cc_603 N_A_803_74#_c_616_n N_A_616_74#_c_1307_n 0.00224787f $X=4.945 $Y=1.095
+ $X2=0 $Y2=0
cc_604 N_A_803_74#_c_617_n N_A_616_74#_c_1307_n 0.0116925f $X=4.945 $Y=1.265
+ $X2=0 $Y2=0
cc_605 N_A_803_74#_c_620_n N_A_616_74#_c_1307_n 0.0227674f $X=5.18 $Y=1.565
+ $X2=0 $Y2=0
cc_606 N_A_803_74#_c_612_n N_A_616_74#_c_1308_n 7.84041e-19 $X=4.155 $Y=0.515
+ $X2=0 $Y2=0
cc_607 N_A_803_74#_c_613_n N_A_616_74#_c_1308_n 9.3219e-19 $X=4.97 $Y=0.34 $X2=0
+ $Y2=0
cc_608 N_A_803_74#_c_623_n N_A_616_74#_c_1321_n 0.00737233f $X=5.09 $Y=2.21
+ $X2=0 $Y2=0
cc_609 N_A_803_74#_c_628_n N_A_616_74#_c_1321_n 0.0192654f $X=5.66 $Y=2.98 $X2=0
+ $Y2=0
cc_610 N_A_803_74#_M1020_g N_A_616_74#_M1002_g 0.012438f $X=5.69 $Y=0.615 $X2=0
+ $Y2=0
cc_611 N_A_803_74#_c_612_n N_A_616_74#_M1002_g 0.00380453f $X=4.155 $Y=0.515
+ $X2=0 $Y2=0
cc_612 N_A_803_74#_c_613_n N_A_616_74#_M1002_g 0.0101814f $X=4.97 $Y=0.34 $X2=0
+ $Y2=0
cc_613 N_A_803_74#_c_616_n N_A_616_74#_M1002_g 0.0218233f $X=4.945 $Y=1.095
+ $X2=0 $Y2=0
cc_614 N_A_803_74#_c_623_n N_A_616_74#_c_1323_n 0.00808094f $X=5.09 $Y=2.21
+ $X2=0 $Y2=0
cc_615 N_A_803_74#_c_628_n N_A_616_74#_c_1323_n 0.00861452f $X=5.66 $Y=2.98
+ $X2=0 $Y2=0
cc_616 N_A_803_74#_c_650_p N_A_616_74#_c_1323_n 0.0118724f $X=5.745 $Y=2.895
+ $X2=0 $Y2=0
cc_617 N_A_803_74#_c_640_n N_A_616_74#_c_1323_n 8.34741e-19 $X=5.665 $Y=1.94
+ $X2=0 $Y2=0
cc_618 N_A_803_74#_c_641_n N_A_616_74#_c_1323_n 0.00846394f $X=5.665 $Y=1.94
+ $X2=0 $Y2=0
cc_619 N_A_803_74#_c_642_n N_A_616_74#_c_1323_n 0.00337651f $X=5.745 $Y=2.375
+ $X2=0 $Y2=0
cc_620 N_A_803_74#_c_628_n N_A_616_74#_c_1324_n 0.00281269f $X=5.66 $Y=2.98
+ $X2=0 $Y2=0
cc_621 N_A_803_74#_c_651_p N_A_616_74#_c_1324_n 0.0100157f $X=6.695 $Y=2.375
+ $X2=0 $Y2=0
cc_622 N_A_803_74#_c_632_n N_A_616_74#_c_1324_n 0.0124701f $X=7.375 $Y=2.98
+ $X2=0 $Y2=0
cc_623 N_A_803_74#_c_633_n N_A_616_74#_c_1324_n 0.00297952f $X=6.865 $Y=2.98
+ $X2=0 $Y2=0
cc_624 N_A_803_74#_c_638_n N_A_616_74#_c_1325_n 0.00453866f $X=10.435 $Y=1.845
+ $X2=0 $Y2=0
cc_625 N_A_803_74#_c_626_n N_A_616_74#_c_1326_n 0.00209279f $X=10.44 $Y=2.465
+ $X2=0 $Y2=0
cc_626 N_A_803_74#_c_638_n N_A_616_74#_c_1327_n 0.0188003f $X=10.435 $Y=1.845
+ $X2=0 $Y2=0
cc_627 N_A_803_74#_c_618_n N_A_616_74#_c_1327_n 9.5574e-19 $X=9.21 $Y=1.615
+ $X2=0 $Y2=0
cc_628 N_A_803_74#_c_646_n N_A_616_74#_c_1327_n 7.89963e-19 $X=10.6 $Y=1.845
+ $X2=0 $Y2=0
cc_629 N_A_803_74#_c_647_n N_A_616_74#_c_1327_n 0.0095945f $X=10.6 $Y=1.97 $X2=0
+ $Y2=0
cc_630 N_A_803_74#_c_626_n N_A_616_74#_M1030_g 0.0106525f $X=10.44 $Y=2.465
+ $X2=0 $Y2=0
cc_631 N_A_803_74#_c_646_n N_A_616_74#_M1030_g 3.92296e-19 $X=10.6 $Y=1.845
+ $X2=0 $Y2=0
cc_632 N_A_803_74#_c_647_n N_A_616_74#_M1030_g 0.0147687f $X=10.6 $Y=1.97 $X2=0
+ $Y2=0
cc_633 N_A_803_74#_c_638_n N_A_616_74#_c_1310_n 0.00828996f $X=10.435 $Y=1.845
+ $X2=0 $Y2=0
cc_634 N_A_803_74#_c_646_n N_A_616_74#_c_1310_n 0.00161435f $X=10.6 $Y=1.845
+ $X2=0 $Y2=0
cc_635 N_A_803_74#_c_647_n N_A_616_74#_c_1310_n 0.0267607f $X=10.6 $Y=1.97 $X2=0
+ $Y2=0
cc_636 N_A_803_74#_c_608_n N_A_616_74#_c_1311_n 0.0256532f $X=10.085 $Y=1.16
+ $X2=0 $Y2=0
cc_637 N_A_803_74#_c_618_n N_A_616_74#_c_1311_n 0.00217356f $X=9.21 $Y=1.615
+ $X2=0 $Y2=0
cc_638 N_A_803_74#_c_619_n N_A_616_74#_c_1311_n 0.0050123f $X=9.21 $Y=1.615
+ $X2=0 $Y2=0
cc_639 N_A_803_74#_c_621_n N_A_616_74#_c_1311_n 0.00433442f $X=9.21 $Y=1.45
+ $X2=0 $Y2=0
cc_640 N_A_803_74#_c_609_n N_A_616_74#_M1026_g 0.0179159f $X=10.16 $Y=1.085
+ $X2=0 $Y2=0
cc_641 N_A_803_74#_c_622_n N_A_616_74#_c_1331_n 0.00337584f $X=5.09 $Y=2.12
+ $X2=0 $Y2=0
cc_642 N_A_803_74#_c_628_n N_A_616_74#_c_1332_n 0.00766255f $X=5.66 $Y=2.98
+ $X2=0 $Y2=0
cc_643 N_A_803_74#_M1040_d N_A_616_74#_c_1335_n 0.00345847f $X=4.035 $Y=1.84
+ $X2=0 $Y2=0
cc_644 N_A_803_74#_c_612_n N_A_616_74#_c_1315_n 0.010537f $X=4.155 $Y=0.515
+ $X2=0 $Y2=0
cc_645 N_A_803_74#_c_625_n N_A_2191_180#_c_1504_n 0.00378106f $X=10.44 $Y=2.375
+ $X2=0 $Y2=0
cc_646 N_A_803_74#_c_646_n N_A_2191_180#_c_1504_n 6.86031e-19 $X=10.6 $Y=1.845
+ $X2=0 $Y2=0
cc_647 N_A_803_74#_c_647_n N_A_2191_180#_c_1504_n 0.0209128f $X=10.6 $Y=1.97
+ $X2=0 $Y2=0
cc_648 N_A_803_74#_c_626_n N_A_2191_180#_c_1513_n 0.0162229f $X=10.44 $Y=2.465
+ $X2=0 $Y2=0
cc_649 N_A_803_74#_c_606_n N_A_1823_524#_c_1612_n 0.00620571f $X=9.375 $Y=1.16
+ $X2=0 $Y2=0
cc_650 N_A_803_74#_c_607_n N_A_1823_524#_c_1612_n 0.00684765f $X=9.73 $Y=1.085
+ $X2=0 $Y2=0
cc_651 N_A_803_74#_c_609_n N_A_1823_524#_c_1612_n 6.02622e-19 $X=10.16 $Y=1.085
+ $X2=0 $Y2=0
cc_652 N_A_803_74#_c_626_n N_A_1823_524#_c_1628_n 0.00515847f $X=10.44 $Y=2.465
+ $X2=0 $Y2=0
cc_653 N_A_803_74#_c_607_n N_A_1823_524#_c_1613_n 0.0100711f $X=9.73 $Y=1.085
+ $X2=0 $Y2=0
cc_654 N_A_803_74#_c_608_n N_A_1823_524#_c_1613_n 2.69874e-19 $X=10.085 $Y=1.16
+ $X2=0 $Y2=0
cc_655 N_A_803_74#_c_609_n N_A_1823_524#_c_1613_n 0.0119826f $X=10.16 $Y=1.085
+ $X2=0 $Y2=0
cc_656 N_A_803_74#_c_607_n N_A_1823_524#_c_1614_n 0.00281658f $X=9.73 $Y=1.085
+ $X2=0 $Y2=0
cc_657 N_A_803_74#_c_626_n N_A_1823_524#_c_1647_n 0.00621217f $X=10.44 $Y=2.465
+ $X2=0 $Y2=0
cc_658 N_A_803_74#_c_607_n N_A_1823_524#_c_1615_n 6.45594e-19 $X=9.73 $Y=1.085
+ $X2=0 $Y2=0
cc_659 N_A_803_74#_c_608_n N_A_1823_524#_c_1615_n 0.00456139f $X=10.085 $Y=1.16
+ $X2=0 $Y2=0
cc_660 N_A_803_74#_c_609_n N_A_1823_524#_c_1615_n 0.00890023f $X=10.16 $Y=1.085
+ $X2=0 $Y2=0
cc_661 N_A_803_74#_c_625_n N_A_1823_524#_c_1629_n 0.00448992f $X=10.44 $Y=2.375
+ $X2=0 $Y2=0
cc_662 N_A_803_74#_c_626_n N_A_1823_524#_c_1629_n 0.00663072f $X=10.44 $Y=2.465
+ $X2=0 $Y2=0
cc_663 N_A_803_74#_c_638_n N_A_1823_524#_c_1629_n 0.00183155f $X=10.435 $Y=1.845
+ $X2=0 $Y2=0
cc_664 N_A_803_74#_c_646_n N_A_1823_524#_c_1629_n 0.0234423f $X=10.6 $Y=1.845
+ $X2=0 $Y2=0
cc_665 N_A_803_74#_c_647_n N_A_1823_524#_c_1629_n 0.00163915f $X=10.6 $Y=1.97
+ $X2=0 $Y2=0
cc_666 N_A_803_74#_c_625_n N_A_1823_524#_c_1630_n 0.0014663f $X=10.44 $Y=2.375
+ $X2=0 $Y2=0
cc_667 N_A_803_74#_c_626_n N_A_1823_524#_c_1630_n 0.00179803f $X=10.44 $Y=2.465
+ $X2=0 $Y2=0
cc_668 N_A_803_74#_c_638_n N_A_1823_524#_c_1630_n 0.0126895f $X=10.435 $Y=1.845
+ $X2=0 $Y2=0
cc_669 N_A_803_74#_c_646_n N_A_1823_524#_c_1616_n 0.0116831f $X=10.6 $Y=1.845
+ $X2=0 $Y2=0
cc_670 N_A_803_74#_c_647_n N_A_1823_524#_c_1616_n 3.42788e-19 $X=10.6 $Y=1.97
+ $X2=0 $Y2=0
cc_671 N_A_803_74#_c_638_n N_A_1823_524#_c_1617_n 0.0122097f $X=10.435 $Y=1.845
+ $X2=0 $Y2=0
cc_672 N_A_803_74#_c_646_n N_A_1823_524#_c_1617_n 0.00602652f $X=10.6 $Y=1.845
+ $X2=0 $Y2=0
cc_673 N_A_803_74#_c_647_n N_A_1823_524#_c_1617_n 2.04636e-19 $X=10.6 $Y=1.97
+ $X2=0 $Y2=0
cc_674 N_A_803_74#_c_625_n N_A_1823_524#_c_1618_n 0.00294488f $X=10.44 $Y=2.375
+ $X2=0 $Y2=0
cc_675 N_A_803_74#_c_646_n N_A_1823_524#_c_1618_n 0.0283689f $X=10.6 $Y=1.845
+ $X2=0 $Y2=0
cc_676 N_A_803_74#_c_647_n N_A_1823_524#_c_1618_n 0.0017947f $X=10.6 $Y=1.97
+ $X2=0 $Y2=0
cc_677 N_A_803_74#_c_651_p N_VPWR_M1004_d 0.0122668f $X=6.695 $Y=2.375 $X2=0
+ $Y2=0
cc_678 N_A_803_74#_c_631_n N_VPWR_M1004_d 0.00328856f $X=6.78 $Y=2.895 $X2=0
+ $Y2=0
cc_679 N_A_803_74#_c_634_n N_VPWR_M1006_d 0.00387922f $X=7.46 $Y=2.895 $X2=0
+ $Y2=0
cc_680 N_A_803_74#_c_635_n N_VPWR_M1006_d 0.00274975f $X=7.725 $Y=2.035 $X2=0
+ $Y2=0
cc_681 N_A_803_74#_c_643_n N_VPWR_M1006_d 0.00407918f $X=7.81 $Y=1.865 $X2=0
+ $Y2=0
cc_682 N_A_803_74#_c_637_n N_VPWR_M1047_s 0.00254193f $X=9.045 $Y=1.865 $X2=0
+ $Y2=0
cc_683 N_A_803_74#_c_639_n N_VPWR_c_1951_n 0.0225252f $X=4.235 $Y=2.78 $X2=0
+ $Y2=0
cc_684 N_A_803_74#_c_628_n N_VPWR_c_1952_n 0.00756371f $X=5.66 $Y=2.98 $X2=0
+ $Y2=0
cc_685 N_A_803_74#_c_650_p N_VPWR_c_1952_n 0.0100041f $X=5.745 $Y=2.895 $X2=0
+ $Y2=0
cc_686 N_A_803_74#_c_651_p N_VPWR_c_1952_n 0.0201769f $X=6.695 $Y=2.375 $X2=0
+ $Y2=0
cc_687 N_A_803_74#_c_631_n N_VPWR_c_1952_n 0.0200357f $X=6.78 $Y=2.895 $X2=0
+ $Y2=0
cc_688 N_A_803_74#_c_633_n N_VPWR_c_1952_n 0.014681f $X=6.865 $Y=2.98 $X2=0
+ $Y2=0
cc_689 N_A_803_74#_c_632_n N_VPWR_c_1953_n 0.0143583f $X=7.375 $Y=2.98 $X2=0
+ $Y2=0
cc_690 N_A_803_74#_c_634_n N_VPWR_c_1953_n 0.0444111f $X=7.46 $Y=2.895 $X2=0
+ $Y2=0
cc_691 N_A_803_74#_c_635_n N_VPWR_c_1953_n 7.09171e-19 $X=7.725 $Y=2.035 $X2=0
+ $Y2=0
cc_692 N_A_803_74#_c_643_n N_VPWR_c_1953_n 0.0131499f $X=7.81 $Y=1.865 $X2=0
+ $Y2=0
cc_693 N_A_803_74#_c_626_n N_VPWR_c_1955_n 5.52504e-19 $X=10.44 $Y=2.465 $X2=0
+ $Y2=0
cc_694 N_A_803_74#_c_632_n N_VPWR_c_1961_n 0.0423147f $X=7.375 $Y=2.98 $X2=0
+ $Y2=0
cc_695 N_A_803_74#_c_633_n N_VPWR_c_1961_n 0.0114574f $X=6.865 $Y=2.98 $X2=0
+ $Y2=0
cc_696 N_A_803_74#_c_628_n N_VPWR_c_1967_n 0.0868345f $X=5.66 $Y=2.98 $X2=0
+ $Y2=0
cc_697 N_A_803_74#_c_639_n N_VPWR_c_1967_n 0.021564f $X=4.235 $Y=2.78 $X2=0
+ $Y2=0
cc_698 N_A_803_74#_c_626_n N_VPWR_c_1968_n 0.00449242f $X=10.44 $Y=2.465 $X2=0
+ $Y2=0
cc_699 N_A_803_74#_c_626_n N_VPWR_c_1947_n 0.0046176f $X=10.44 $Y=2.465 $X2=0
+ $Y2=0
cc_700 N_A_803_74#_c_628_n N_VPWR_c_1947_n 0.0478959f $X=5.66 $Y=2.98 $X2=0
+ $Y2=0
cc_701 N_A_803_74#_c_632_n N_VPWR_c_1947_n 0.0229174f $X=7.375 $Y=2.98 $X2=0
+ $Y2=0
cc_702 N_A_803_74#_c_633_n N_VPWR_c_1947_n 0.00589978f $X=6.865 $Y=2.98 $X2=0
+ $Y2=0
cc_703 N_A_803_74#_c_639_n N_VPWR_c_1947_n 0.0125777f $X=4.235 $Y=2.78 $X2=0
+ $Y2=0
cc_704 N_A_803_74#_c_613_n N_A_288_464#_M1002_s 0.00378448f $X=4.97 $Y=0.34
+ $X2=0 $Y2=0
cc_705 N_A_803_74#_M1040_d N_A_288_464#_c_2169_n 0.00517424f $X=4.035 $Y=1.84
+ $X2=0 $Y2=0
cc_706 N_A_803_74#_c_628_n N_A_288_464#_c_2169_n 3.46483e-19 $X=5.66 $Y=2.98
+ $X2=0 $Y2=0
cc_707 N_A_803_74#_c_639_n N_A_288_464#_c_2169_n 0.0245989f $X=4.235 $Y=2.78
+ $X2=0 $Y2=0
cc_708 N_A_803_74#_c_622_n N_A_288_464#_c_2165_n 0.00132424f $X=5.09 $Y=2.12
+ $X2=0 $Y2=0
cc_709 N_A_803_74#_c_612_n N_A_288_464#_c_2165_n 0.0148507f $X=4.155 $Y=0.515
+ $X2=0 $Y2=0
cc_710 N_A_803_74#_c_616_n N_A_288_464#_c_2165_n 0.0063104f $X=4.945 $Y=1.095
+ $X2=0 $Y2=0
cc_711 N_A_803_74#_c_617_n N_A_288_464#_c_2165_n 0.0479185f $X=4.945 $Y=1.265
+ $X2=0 $Y2=0
cc_712 N_A_803_74#_c_620_n N_A_288_464#_c_2165_n 0.00192596f $X=5.18 $Y=1.565
+ $X2=0 $Y2=0
cc_713 N_A_803_74#_c_612_n N_A_288_464#_c_2166_n 0.0260385f $X=4.155 $Y=0.515
+ $X2=0 $Y2=0
cc_714 N_A_803_74#_c_613_n N_A_288_464#_c_2166_n 0.0283886f $X=4.97 $Y=0.34
+ $X2=0 $Y2=0
cc_715 N_A_803_74#_c_616_n N_A_288_464#_c_2166_n 0.0247538f $X=4.945 $Y=1.095
+ $X2=0 $Y2=0
cc_716 N_A_803_74#_c_617_n N_A_288_464#_c_2166_n 0.00409016f $X=4.945 $Y=1.265
+ $X2=0 $Y2=0
cc_717 N_A_803_74#_c_622_n N_A_288_464#_c_2172_n 0.00638897f $X=5.09 $Y=2.12
+ $X2=0 $Y2=0
cc_718 N_A_803_74#_c_623_n N_A_288_464#_c_2172_n 0.00974949f $X=5.09 $Y=2.21
+ $X2=0 $Y2=0
cc_719 N_A_803_74#_c_628_n N_A_288_464#_c_2172_n 0.0365228f $X=5.66 $Y=2.98
+ $X2=0 $Y2=0
cc_720 N_A_803_74#_c_615_n N_A_288_464#_c_2172_n 0.0245583f $X=4.9 $Y=1.565
+ $X2=0 $Y2=0
cc_721 N_A_803_74#_c_639_n N_A_288_464#_c_2172_n 0.00814501f $X=4.235 $Y=2.78
+ $X2=0 $Y2=0
cc_722 N_A_803_74#_c_620_n N_A_288_464#_c_2172_n 0.00268183f $X=5.18 $Y=1.565
+ $X2=0 $Y2=0
cc_723 N_A_803_74#_c_650_p A_1140_495# 0.00566423f $X=5.745 $Y=2.895 $X2=-0.19
+ $Y2=-0.245
cc_724 N_A_803_74#_c_651_p A_1140_495# 0.00920595f $X=6.695 $Y=2.375 $X2=-0.19
+ $Y2=-0.245
cc_725 N_A_803_74#_c_637_n N_A_1620_373#_M1035_d 0.00197722f $X=9.045 $Y=1.865
+ $X2=-0.19 $Y2=-0.245
cc_726 N_A_803_74#_c_634_n N_A_1620_373#_c_2293_n 0.00561307f $X=7.46 $Y=2.895
+ $X2=0 $Y2=0
cc_727 N_A_803_74#_c_637_n N_A_1620_373#_c_2293_n 0.0151437f $X=9.045 $Y=1.865
+ $X2=0 $Y2=0
cc_728 N_A_803_74#_c_637_n N_A_1620_373#_c_2290_n 0.0403185f $X=9.045 $Y=1.865
+ $X2=0 $Y2=0
cc_729 N_A_803_74#_c_638_n N_A_1620_373#_c_2290_n 0.00951534f $X=10.435 $Y=1.845
+ $X2=0 $Y2=0
cc_730 N_A_803_74#_c_618_n N_A_1620_373#_c_2290_n 0.0247616f $X=9.21 $Y=1.615
+ $X2=0 $Y2=0
cc_731 N_A_803_74#_c_619_n N_A_1620_373#_c_2290_n 0.00149284f $X=9.21 $Y=1.615
+ $X2=0 $Y2=0
cc_732 N_A_803_74#_c_638_n N_A_1620_373#_c_2291_n 0.0256373f $X=10.435 $Y=1.845
+ $X2=0 $Y2=0
cc_733 N_A_803_74#_c_646_n N_A_1620_373#_c_2291_n 0.00101189f $X=10.6 $Y=1.845
+ $X2=0 $Y2=0
cc_734 N_A_803_74#_c_647_n N_A_1620_373#_c_2291_n 8.54694e-19 $X=10.6 $Y=1.97
+ $X2=0 $Y2=0
cc_735 N_A_803_74#_c_626_n A_2103_508# 0.00233754f $X=10.44 $Y=2.465 $X2=-0.19
+ $Y2=-0.245
cc_736 N_A_803_74#_c_614_n N_VGND_c_2417_n 0.0112234f $X=4.24 $Y=0.34 $X2=0
+ $Y2=0
cc_737 N_A_803_74#_c_607_n N_VGND_c_2420_n 0.00176715f $X=9.73 $Y=1.085 $X2=0
+ $Y2=0
cc_738 N_A_803_74#_M1020_g N_VGND_c_2430_n 0.00527282f $X=5.69 $Y=0.615 $X2=0
+ $Y2=0
cc_739 N_A_803_74#_c_613_n N_VGND_c_2430_n 0.0591538f $X=4.97 $Y=0.34 $X2=0
+ $Y2=0
cc_740 N_A_803_74#_c_614_n N_VGND_c_2430_n 0.0121867f $X=4.24 $Y=0.34 $X2=0
+ $Y2=0
cc_741 N_A_803_74#_c_607_n N_VGND_c_2433_n 0.00278247f $X=9.73 $Y=1.085 $X2=0
+ $Y2=0
cc_742 N_A_803_74#_c_609_n N_VGND_c_2433_n 0.00278247f $X=10.16 $Y=1.085 $X2=0
+ $Y2=0
cc_743 N_A_803_74#_M1020_g N_VGND_c_2444_n 0.00534666f $X=5.69 $Y=0.615 $X2=0
+ $Y2=0
cc_744 N_A_803_74#_c_607_n N_VGND_c_2444_n 0.00358425f $X=9.73 $Y=1.085 $X2=0
+ $Y2=0
cc_745 N_A_803_74#_c_609_n N_VGND_c_2444_n 0.0035422f $X=10.16 $Y=1.085 $X2=0
+ $Y2=0
cc_746 N_A_803_74#_c_613_n N_VGND_c_2444_n 0.0340476f $X=4.97 $Y=0.34 $X2=0
+ $Y2=0
cc_747 N_A_803_74#_c_614_n N_VGND_c_2444_n 0.00660921f $X=4.24 $Y=0.34 $X2=0
+ $Y2=0
cc_748 N_A_803_74#_c_605_n N_A_1677_74#_c_2591_n 0.00893137f $X=9.655 $Y=1.16
+ $X2=0 $Y2=0
cc_749 N_A_803_74#_c_606_n N_A_1677_74#_c_2591_n 0.00849831f $X=9.375 $Y=1.16
+ $X2=0 $Y2=0
cc_750 N_A_803_74#_c_608_n N_A_1677_74#_c_2591_n 0.00792883f $X=10.085 $Y=1.16
+ $X2=0 $Y2=0
cc_751 N_A_803_74#_c_611_n N_A_1677_74#_c_2591_n 0.00988318f $X=9.73 $Y=1.16
+ $X2=0 $Y2=0
cc_752 N_A_803_74#_c_637_n N_A_1677_74#_c_2591_n 0.00700312f $X=9.045 $Y=1.865
+ $X2=0 $Y2=0
cc_753 N_A_803_74#_c_638_n N_A_1677_74#_c_2591_n 0.0112447f $X=10.435 $Y=1.845
+ $X2=0 $Y2=0
cc_754 N_A_803_74#_c_618_n N_A_1677_74#_c_2591_n 0.0234872f $X=9.21 $Y=1.615
+ $X2=0 $Y2=0
cc_755 N_A_803_74#_c_619_n N_A_1677_74#_c_2591_n 0.00126186f $X=9.21 $Y=1.615
+ $X2=0 $Y2=0
cc_756 N_A_803_74#_c_621_n N_A_1677_74#_c_2591_n 0.00448379f $X=9.21 $Y=1.45
+ $X2=0 $Y2=0
cc_757 N_A_803_74#_c_637_n N_A_1677_74#_c_2592_n 0.00261373f $X=9.045 $Y=1.865
+ $X2=0 $Y2=0
cc_758 N_A_803_74#_c_607_n N_A_1677_74#_c_2593_n 0.00187125f $X=9.73 $Y=1.085
+ $X2=0 $Y2=0
cc_759 N_A_803_74#_c_608_n N_A_1677_74#_c_2593_n 0.00397268f $X=10.085 $Y=1.16
+ $X2=0 $Y2=0
cc_760 N_A_803_74#_c_609_n N_A_1677_74#_c_2593_n 6.33289e-19 $X=10.16 $Y=1.085
+ $X2=0 $Y2=0
cc_761 N_A_1201_55#_c_907_n N_A_1017_81#_c_1002_n 0.0126216f $X=6.13 $Y=2.21
+ $X2=0 $Y2=0
cc_762 N_A_1201_55#_c_909_n N_A_1017_81#_c_1002_n 0.0146017f $X=7.035 $Y=2.035
+ $X2=0 $Y2=0
cc_763 N_A_1201_55#_c_911_n N_A_1017_81#_c_1002_n 0.0011051f $X=6.205 $Y=1.945
+ $X2=0 $Y2=0
cc_764 N_A_1201_55#_c_907_n N_A_1017_81#_c_1003_n 0.00954336f $X=6.13 $Y=2.21
+ $X2=0 $Y2=0
cc_765 N_A_1201_55#_c_910_n N_A_1017_81#_c_1003_n 0.00527003f $X=7.12 $Y=2.495
+ $X2=0 $Y2=0
cc_766 N_A_1201_55#_c_902_n N_A_1017_81#_c_987_n 0.00371558f $X=6.77 $Y=0.855
+ $X2=0 $Y2=0
cc_767 N_A_1201_55#_c_903_n N_A_1017_81#_c_987_n 0.00789289f $X=6.935 $Y=0.58
+ $X2=0 $Y2=0
cc_768 N_A_1201_55#_c_901_n N_A_1017_81#_c_992_n 0.0147338f $X=6.26 $Y=1.78
+ $X2=0 $Y2=0
cc_769 N_A_1201_55#_c_909_n N_A_1017_81#_c_993_n 0.00103763f $X=7.035 $Y=2.035
+ $X2=0 $Y2=0
cc_770 N_A_1201_55#_c_907_n N_A_1017_81#_c_1009_n 2.50685e-19 $X=6.13 $Y=2.21
+ $X2=0 $Y2=0
cc_771 N_A_1201_55#_c_901_n N_A_1017_81#_c_994_n 7.71193e-19 $X=6.26 $Y=1.78
+ $X2=0 $Y2=0
cc_772 N_A_1201_55#_c_904_n N_A_1017_81#_c_994_n 0.020088f $X=6.17 $Y=0.855
+ $X2=0 $Y2=0
cc_773 N_A_1201_55#_c_906_n N_A_1017_81#_c_994_n 0.00291423f $X=6.17 $Y=0.935
+ $X2=0 $Y2=0
cc_774 N_A_1201_55#_c_907_n N_A_1017_81#_c_995_n 7.82209e-19 $X=6.13 $Y=2.21
+ $X2=0 $Y2=0
cc_775 N_A_1201_55#_c_901_n N_A_1017_81#_c_995_n 0.011116f $X=6.26 $Y=1.78 $X2=0
+ $Y2=0
cc_776 N_A_1201_55#_c_902_n N_A_1017_81#_c_995_n 0.0104262f $X=6.77 $Y=0.855
+ $X2=0 $Y2=0
cc_777 N_A_1201_55#_c_909_n N_A_1017_81#_c_995_n 0.0117696f $X=7.035 $Y=2.035
+ $X2=0 $Y2=0
cc_778 N_A_1201_55#_c_904_n N_A_1017_81#_c_995_n 0.0250033f $X=6.17 $Y=0.855
+ $X2=0 $Y2=0
cc_779 N_A_1201_55#_c_905_n N_A_1017_81#_c_995_n 7.8432e-19 $X=6.17 $Y=1.1 $X2=0
+ $Y2=0
cc_780 N_A_1201_55#_c_911_n N_A_1017_81#_c_995_n 0.0237253f $X=6.205 $Y=1.945
+ $X2=0 $Y2=0
cc_781 N_A_1201_55#_c_902_n N_A_1017_81#_c_996_n 0.0114571f $X=6.77 $Y=0.855
+ $X2=0 $Y2=0
cc_782 N_A_1201_55#_c_909_n N_A_1017_81#_c_996_n 0.00746539f $X=7.035 $Y=2.035
+ $X2=0 $Y2=0
cc_783 N_A_1201_55#_c_901_n N_A_1017_81#_c_998_n 0.00119856f $X=6.26 $Y=1.78
+ $X2=0 $Y2=0
cc_784 N_A_1201_55#_c_902_n N_A_1017_81#_c_998_n 0.0270039f $X=6.77 $Y=0.855
+ $X2=0 $Y2=0
cc_785 N_A_1201_55#_c_909_n N_A_1017_81#_c_998_n 0.0255117f $X=7.035 $Y=2.035
+ $X2=0 $Y2=0
cc_786 N_A_1201_55#_c_904_n N_A_1017_81#_c_998_n 0.00758966f $X=6.17 $Y=0.855
+ $X2=0 $Y2=0
cc_787 N_A_1201_55#_c_905_n N_A_1017_81#_c_998_n 0.00166639f $X=6.17 $Y=1.1
+ $X2=0 $Y2=0
cc_788 N_A_1201_55#_c_902_n N_A_1017_81#_c_999_n 0.0151126f $X=6.77 $Y=0.855
+ $X2=0 $Y2=0
cc_789 N_A_1201_55#_c_904_n N_A_1017_81#_c_999_n 0.00166032f $X=6.17 $Y=0.855
+ $X2=0 $Y2=0
cc_790 N_A_1201_55#_c_905_n N_A_1017_81#_c_999_n 0.0197395f $X=6.17 $Y=1.1 $X2=0
+ $Y2=0
cc_791 N_A_1201_55#_c_906_n N_A_1017_81#_c_999_n 7.97846e-19 $X=6.17 $Y=0.935
+ $X2=0 $Y2=0
cc_792 N_A_1201_55#_c_909_n N_SET_B_c_1169_n 0.00145714f $X=7.035 $Y=2.035 $X2=0
+ $Y2=0
cc_793 N_A_1201_55#_c_910_n N_SET_B_c_1170_n 0.00266484f $X=7.12 $Y=2.495 $X2=0
+ $Y2=0
cc_794 N_A_1201_55#_c_902_n N_SET_B_M1003_g 4.99343e-19 $X=6.77 $Y=0.855 $X2=0
+ $Y2=0
cc_795 N_A_1201_55#_c_903_n N_SET_B_M1003_g 0.00118801f $X=6.935 $Y=0.58 $X2=0
+ $Y2=0
cc_796 N_A_1201_55#_c_909_n N_SET_B_c_1165_n 8.43333e-19 $X=7.035 $Y=2.035 $X2=0
+ $Y2=0
cc_797 N_A_1201_55#_c_909_n N_SET_B_c_1166_n 2.32957e-19 $X=7.035 $Y=2.035 $X2=0
+ $Y2=0
cc_798 N_A_1201_55#_c_907_n N_A_616_74#_c_1323_n 0.0148903f $X=6.13 $Y=2.21
+ $X2=0 $Y2=0
cc_799 N_A_1201_55#_c_907_n N_A_616_74#_c_1324_n 0.0086575f $X=6.13 $Y=2.21
+ $X2=0 $Y2=0
cc_800 N_A_1201_55#_c_907_n N_VPWR_c_1952_n 0.00294083f $X=6.13 $Y=2.21 $X2=0
+ $Y2=0
cc_801 N_A_1201_55#_c_907_n N_VPWR_c_1947_n 9.49986e-19 $X=6.13 $Y=2.21 $X2=0
+ $Y2=0
cc_802 N_A_1201_55#_c_902_n N_VGND_M1019_d 0.00207662f $X=6.77 $Y=0.855 $X2=0
+ $Y2=0
cc_803 N_A_1201_55#_c_904_n N_VGND_M1019_d 0.00147032f $X=6.17 $Y=0.855 $X2=0
+ $Y2=0
cc_804 N_A_1201_55#_c_902_n N_VGND_c_2418_n 0.0161913f $X=6.77 $Y=0.855 $X2=0
+ $Y2=0
cc_805 N_A_1201_55#_c_903_n N_VGND_c_2418_n 0.0168548f $X=6.935 $Y=0.58 $X2=0
+ $Y2=0
cc_806 N_A_1201_55#_c_904_n N_VGND_c_2418_n 0.0104232f $X=6.17 $Y=0.855 $X2=0
+ $Y2=0
cc_807 N_A_1201_55#_c_905_n N_VGND_c_2418_n 6.45517e-19 $X=6.17 $Y=1.1 $X2=0
+ $Y2=0
cc_808 N_A_1201_55#_c_906_n N_VGND_c_2418_n 0.00891712f $X=6.17 $Y=0.935 $X2=0
+ $Y2=0
cc_809 N_A_1201_55#_c_902_n N_VGND_c_2419_n 0.00564835f $X=6.77 $Y=0.855 $X2=0
+ $Y2=0
cc_810 N_A_1201_55#_c_903_n N_VGND_c_2419_n 0.0140506f $X=6.935 $Y=0.58 $X2=0
+ $Y2=0
cc_811 N_A_1201_55#_c_906_n N_VGND_c_2430_n 0.00552345f $X=6.17 $Y=0.935 $X2=0
+ $Y2=0
cc_812 N_A_1201_55#_c_903_n N_VGND_c_2431_n 0.014415f $X=6.935 $Y=0.58 $X2=0
+ $Y2=0
cc_813 N_A_1201_55#_c_902_n N_VGND_c_2444_n 0.00920397f $X=6.77 $Y=0.855 $X2=0
+ $Y2=0
cc_814 N_A_1201_55#_c_903_n N_VGND_c_2444_n 0.0119404f $X=6.935 $Y=0.58 $X2=0
+ $Y2=0
cc_815 N_A_1201_55#_c_904_n N_VGND_c_2444_n 0.0082444f $X=6.17 $Y=0.855 $X2=0
+ $Y2=0
cc_816 N_A_1201_55#_c_906_n N_VGND_c_2444_n 0.00534666f $X=6.17 $Y=0.935 $X2=0
+ $Y2=0
cc_817 N_A_1017_81#_c_1002_n N_SET_B_c_1169_n 0.00873199f $X=6.865 $Y=2.12 $X2=0
+ $Y2=0
cc_818 N_A_1017_81#_c_1005_n N_SET_B_c_1169_n 0.00718294f $X=8.025 $Y=1.79 $X2=0
+ $Y2=0
cc_819 N_A_1017_81#_c_1003_n N_SET_B_c_1170_n 0.0157553f $X=6.865 $Y=2.21 $X2=0
+ $Y2=0
cc_820 N_A_1017_81#_c_1005_n N_SET_B_c_1170_n 0.00705028f $X=8.025 $Y=1.79 $X2=0
+ $Y2=0
cc_821 N_A_1017_81#_c_987_n N_SET_B_M1003_g 0.0395874f $X=7.15 $Y=0.865 $X2=0
+ $Y2=0
cc_822 N_A_1017_81#_c_989_n N_SET_B_M1003_g 0.00633066f $X=8.31 $Y=1.085 $X2=0
+ $Y2=0
cc_823 N_A_1017_81#_c_996_n N_SET_B_M1003_g 0.0161084f $X=7.935 $Y=1.195 $X2=0
+ $Y2=0
cc_824 N_A_1017_81#_c_998_n N_SET_B_M1003_g 0.00100603f $X=6.79 $Y=1.195 $X2=0
+ $Y2=0
cc_825 N_A_1017_81#_c_999_n N_SET_B_M1003_g 0.0103422f $X=6.79 $Y=1.275 $X2=0
+ $Y2=0
cc_826 N_A_1017_81#_c_1000_n N_SET_B_M1003_g 0.00115118f $X=8.1 $Y=1.195 $X2=0
+ $Y2=0
cc_827 N_A_1017_81#_c_1001_n N_SET_B_M1003_g 0.014002f $X=8.475 $Y=1.267 $X2=0
+ $Y2=0
cc_828 N_A_1017_81#_c_988_n N_SET_B_c_1163_n 0.00359996f $X=8.025 $Y=1.7 $X2=0
+ $Y2=0
cc_829 N_A_1017_81#_c_1005_n N_SET_B_c_1163_n 0.00217075f $X=8.025 $Y=1.79 $X2=0
+ $Y2=0
cc_830 N_A_1017_81#_c_990_n N_SET_B_c_1163_n 0.00593846f $X=8.475 $Y=1.7 $X2=0
+ $Y2=0
cc_831 N_A_1017_81#_c_1007_n N_SET_B_c_1163_n 0.00225539f $X=8.475 $Y=1.79 $X2=0
+ $Y2=0
cc_832 N_A_1017_81#_c_996_n N_SET_B_c_1163_n 0.00889936f $X=7.935 $Y=1.195 $X2=0
+ $Y2=0
cc_833 N_A_1017_81#_c_1000_n N_SET_B_c_1163_n 0.00863738f $X=8.1 $Y=1.195 $X2=0
+ $Y2=0
cc_834 N_A_1017_81#_c_1001_n N_SET_B_c_1163_n 8.76419e-19 $X=8.475 $Y=1.267
+ $X2=0 $Y2=0
cc_835 N_A_1017_81#_c_988_n N_SET_B_c_1176_n 2.31912e-19 $X=8.025 $Y=1.7 $X2=0
+ $Y2=0
cc_836 N_A_1017_81#_c_1005_n N_SET_B_c_1176_n 2.31912e-19 $X=8.025 $Y=1.79 $X2=0
+ $Y2=0
cc_837 N_A_1017_81#_c_996_n N_SET_B_c_1176_n 0.00224843f $X=7.935 $Y=1.195 $X2=0
+ $Y2=0
cc_838 N_A_1017_81#_c_998_n N_SET_B_c_1176_n 0.0012711f $X=6.79 $Y=1.195 $X2=0
+ $Y2=0
cc_839 N_A_1017_81#_c_988_n N_SET_B_c_1165_n 0.00254632f $X=8.025 $Y=1.7 $X2=0
+ $Y2=0
cc_840 N_A_1017_81#_c_992_n N_SET_B_c_1165_n 0.00120584f $X=6.79 $Y=1.615 $X2=0
+ $Y2=0
cc_841 N_A_1017_81#_c_996_n N_SET_B_c_1165_n 0.0253086f $X=7.935 $Y=1.195 $X2=0
+ $Y2=0
cc_842 N_A_1017_81#_c_998_n N_SET_B_c_1165_n 0.0174044f $X=6.79 $Y=1.195 $X2=0
+ $Y2=0
cc_843 N_A_1017_81#_c_988_n N_SET_B_c_1166_n 0.014002f $X=8.025 $Y=1.7 $X2=0
+ $Y2=0
cc_844 N_A_1017_81#_c_992_n N_SET_B_c_1166_n 0.0176356f $X=6.79 $Y=1.615 $X2=0
+ $Y2=0
cc_845 N_A_1017_81#_c_996_n N_SET_B_c_1166_n 0.00633174f $X=7.935 $Y=1.195 $X2=0
+ $Y2=0
cc_846 N_A_1017_81#_c_998_n N_SET_B_c_1166_n 4.17584e-19 $X=6.79 $Y=1.195 $X2=0
+ $Y2=0
cc_847 N_A_1017_81#_c_999_n N_SET_B_c_1166_n 6.62393e-19 $X=6.79 $Y=1.275 $X2=0
+ $Y2=0
cc_848 N_A_1017_81#_c_994_n N_A_616_74#_M1002_g 0.00294822f $X=5.475 $Y=0.615
+ $X2=0 $Y2=0
cc_849 N_A_1017_81#_c_1009_n N_A_616_74#_c_1323_n 0.00324522f $X=5.34 $Y=2.415
+ $X2=0 $Y2=0
cc_850 N_A_1017_81#_c_1003_n N_A_616_74#_c_1324_n 0.00739034f $X=6.865 $Y=2.21
+ $X2=0 $Y2=0
cc_851 N_A_1017_81#_c_1005_n N_A_616_74#_c_1324_n 0.00900287f $X=8.025 $Y=1.79
+ $X2=0 $Y2=0
cc_852 N_A_1017_81#_c_1007_n N_A_616_74#_c_1324_n 0.00900015f $X=8.475 $Y=1.79
+ $X2=0 $Y2=0
cc_853 N_A_1017_81#_c_991_n N_A_1823_524#_c_1614_n 6.04331e-19 $X=8.74 $Y=1.085
+ $X2=0 $Y2=0
cc_854 N_A_1017_81#_c_1007_n N_A_1823_524#_c_1636_n 6.66034e-19 $X=8.475 $Y=1.79
+ $X2=0 $Y2=0
cc_855 N_A_1017_81#_c_1003_n N_VPWR_c_1952_n 6.7383e-19 $X=6.865 $Y=2.21 $X2=0
+ $Y2=0
cc_856 N_A_1017_81#_c_1005_n N_VPWR_c_1953_n 0.00344719f $X=8.025 $Y=1.79 $X2=0
+ $Y2=0
cc_857 N_A_1017_81#_c_1005_n N_VPWR_c_1954_n 4.3601e-19 $X=8.025 $Y=1.79 $X2=0
+ $Y2=0
cc_858 N_A_1017_81#_c_1007_n N_VPWR_c_1954_n 0.00762644f $X=8.475 $Y=1.79 $X2=0
+ $Y2=0
cc_859 N_A_1017_81#_c_1005_n N_VPWR_c_1947_n 9.49986e-19 $X=8.025 $Y=1.79 $X2=0
+ $Y2=0
cc_860 N_A_1017_81#_c_1007_n N_VPWR_c_1947_n 8.6132e-19 $X=8.475 $Y=1.79 $X2=0
+ $Y2=0
cc_861 N_A_1017_81#_c_1011_n N_A_288_464#_c_2165_n 0.00512835f $X=5.34 $Y=2.275
+ $X2=0 $Y2=0
cc_862 N_A_1017_81#_c_1011_n N_A_288_464#_c_2172_n 0.048791f $X=5.34 $Y=2.275
+ $X2=0 $Y2=0
cc_863 N_A_1017_81#_c_1005_n N_A_1620_373#_c_2293_n 0.00324443f $X=8.025 $Y=1.79
+ $X2=0 $Y2=0
cc_864 N_A_1017_81#_c_1005_n N_A_1620_373#_c_2289_n 0.00473576f $X=8.025 $Y=1.79
+ $X2=0 $Y2=0
cc_865 N_A_1017_81#_c_1007_n N_A_1620_373#_c_2290_n 0.0142929f $X=8.475 $Y=1.79
+ $X2=0 $Y2=0
cc_866 N_A_1017_81#_c_987_n N_VGND_c_2418_n 0.00324482f $X=7.15 $Y=0.865 $X2=0
+ $Y2=0
cc_867 N_A_1017_81#_c_994_n N_VGND_c_2418_n 0.00331332f $X=5.475 $Y=0.615 $X2=0
+ $Y2=0
cc_868 N_A_1017_81#_c_987_n N_VGND_c_2419_n 0.00222368f $X=7.15 $Y=0.865 $X2=0
+ $Y2=0
cc_869 N_A_1017_81#_c_989_n N_VGND_c_2419_n 0.0112679f $X=8.31 $Y=1.085 $X2=0
+ $Y2=0
cc_870 N_A_1017_81#_c_991_n N_VGND_c_2419_n 4.94598e-19 $X=8.74 $Y=1.085 $X2=0
+ $Y2=0
cc_871 N_A_1017_81#_c_996_n N_VGND_c_2419_n 0.0275558f $X=7.935 $Y=1.195 $X2=0
+ $Y2=0
cc_872 N_A_1017_81#_c_1000_n N_VGND_c_2419_n 0.0243688f $X=8.1 $Y=1.195 $X2=0
+ $Y2=0
cc_873 N_A_1017_81#_c_1001_n N_VGND_c_2419_n 0.00208692f $X=8.475 $Y=1.267 $X2=0
+ $Y2=0
cc_874 N_A_1017_81#_c_989_n N_VGND_c_2420_n 5.01478e-19 $X=8.31 $Y=1.085 $X2=0
+ $Y2=0
cc_875 N_A_1017_81#_c_991_n N_VGND_c_2420_n 0.0114363f $X=8.74 $Y=1.085 $X2=0
+ $Y2=0
cc_876 N_A_1017_81#_c_994_n N_VGND_c_2430_n 0.0127604f $X=5.475 $Y=0.615 $X2=0
+ $Y2=0
cc_877 N_A_1017_81#_c_987_n N_VGND_c_2431_n 0.00434272f $X=7.15 $Y=0.865 $X2=0
+ $Y2=0
cc_878 N_A_1017_81#_c_989_n N_VGND_c_2432_n 0.00383152f $X=8.31 $Y=1.085 $X2=0
+ $Y2=0
cc_879 N_A_1017_81#_c_991_n N_VGND_c_2432_n 0.00383152f $X=8.74 $Y=1.085 $X2=0
+ $Y2=0
cc_880 N_A_1017_81#_c_987_n N_VGND_c_2444_n 0.00825979f $X=7.15 $Y=0.865 $X2=0
+ $Y2=0
cc_881 N_A_1017_81#_c_989_n N_VGND_c_2444_n 0.0075754f $X=8.31 $Y=1.085 $X2=0
+ $Y2=0
cc_882 N_A_1017_81#_c_991_n N_VGND_c_2444_n 0.0075754f $X=8.74 $Y=1.085 $X2=0
+ $Y2=0
cc_883 N_A_1017_81#_c_994_n N_VGND_c_2444_n 0.011834f $X=5.475 $Y=0.615 $X2=0
+ $Y2=0
cc_884 N_A_1017_81#_c_989_n N_A_1677_74#_c_2590_n 0.00190583f $X=8.31 $Y=1.085
+ $X2=0 $Y2=0
cc_885 N_A_1017_81#_c_991_n N_A_1677_74#_c_2590_n 0.00190583f $X=8.74 $Y=1.085
+ $X2=0 $Y2=0
cc_886 N_A_1017_81#_c_1001_n N_A_1677_74#_c_2590_n 0.00425796f $X=8.475 $Y=1.267
+ $X2=0 $Y2=0
cc_887 N_A_1017_81#_c_1001_n N_A_1677_74#_c_2591_n 0.0156828f $X=8.475 $Y=1.267
+ $X2=0 $Y2=0
cc_888 N_A_1017_81#_c_1000_n N_A_1677_74#_c_2592_n 0.0132563f $X=8.1 $Y=1.195
+ $X2=0 $Y2=0
cc_889 N_A_1017_81#_c_1001_n N_A_1677_74#_c_2592_n 0.0096918f $X=8.475 $Y=1.267
+ $X2=0 $Y2=0
cc_890 N_SET_B_c_1170_n N_A_616_74#_c_1324_n 0.00738456f $X=7.345 $Y=2.21 $X2=0
+ $Y2=0
cc_891 N_SET_B_c_1163_n N_A_616_74#_c_1327_n 0.00307872f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_892 N_SET_B_c_1163_n N_A_616_74#_c_1310_n 0.0131967f $X=11.615 $Y=1.665 $X2=0
+ $Y2=0
cc_893 N_SET_B_c_1163_n N_A_616_74#_c_1311_n 0.00448132f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_894 N_SET_B_M1038_g N_A_2191_180#_c_1504_n 0.00916689f $X=11.6 $Y=0.58 $X2=0
+ $Y2=0
cc_895 N_SET_B_c_1163_n N_A_2191_180#_c_1504_n 0.00215544f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_896 N_SET_B_c_1167_n N_A_2191_180#_c_1504_n 0.0231364f $X=11.635 $Y=1.635
+ $X2=0 $Y2=0
cc_897 N_SET_B_c_1168_n N_A_2191_180#_c_1504_n 0.00223173f $X=11.635 $Y=1.635
+ $X2=0 $Y2=0
cc_898 N_SET_B_c_1173_n N_A_2191_180#_c_1513_n 0.0113229f $X=11.515 $Y=2.465
+ $X2=0 $Y2=0
cc_899 N_SET_B_c_1174_n N_A_2191_180#_c_1513_n 0.0231364f $X=11.612 $Y=2.14
+ $X2=0 $Y2=0
cc_900 N_SET_B_M1038_g N_A_2191_180#_c_1505_n 0.0160995f $X=11.6 $Y=0.58 $X2=0
+ $Y2=0
cc_901 N_SET_B_c_1163_n N_A_2191_180#_c_1505_n 0.00661014f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_902 SET_B N_A_2191_180#_c_1505_n 0.00274238f $X=11.675 $Y=1.58 $X2=0 $Y2=0
cc_903 N_SET_B_c_1167_n N_A_2191_180#_c_1505_n 0.00253093f $X=11.635 $Y=1.635
+ $X2=0 $Y2=0
cc_904 N_SET_B_c_1168_n N_A_2191_180#_c_1505_n 0.0139265f $X=11.635 $Y=1.635
+ $X2=0 $Y2=0
cc_905 N_SET_B_M1038_g N_A_2191_180#_c_1506_n 0.0011456f $X=11.6 $Y=0.58 $X2=0
+ $Y2=0
cc_906 N_SET_B_M1038_g N_A_2191_180#_c_1508_n 0.00115306f $X=11.6 $Y=0.58 $X2=0
+ $Y2=0
cc_907 N_SET_B_c_1163_n N_A_2191_180#_c_1508_n 0.00707363f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_908 N_SET_B_M1038_g N_A_2191_180#_c_1509_n 0.0182617f $X=11.6 $Y=0.58 $X2=0
+ $Y2=0
cc_909 N_SET_B_c_1173_n N_A_2191_180#_c_1516_n 6.62644e-19 $X=11.515 $Y=2.465
+ $X2=0 $Y2=0
cc_910 N_SET_B_M1038_g N_A_2191_180#_c_1511_n 0.0225658f $X=11.6 $Y=0.58 $X2=0
+ $Y2=0
cc_911 N_SET_B_M1038_g N_A_1823_524#_M1039_g 0.0230846f $X=11.6 $Y=0.58 $X2=0
+ $Y2=0
cc_912 N_SET_B_c_1174_n N_A_1823_524#_c_1621_n 0.00113802f $X=11.612 $Y=2.14
+ $X2=0 $Y2=0
cc_913 N_SET_B_c_1163_n N_A_1823_524#_c_1629_n 0.00590712f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_914 N_SET_B_M1038_g N_A_1823_524#_c_1616_n 3.68415e-19 $X=11.6 $Y=0.58 $X2=0
+ $Y2=0
cc_915 N_SET_B_c_1163_n N_A_1823_524#_c_1616_n 0.0148238f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_916 N_SET_B_c_1167_n N_A_1823_524#_c_1616_n 3.71364e-19 $X=11.635 $Y=1.635
+ $X2=0 $Y2=0
cc_917 N_SET_B_c_1168_n N_A_1823_524#_c_1616_n 0.00424222f $X=11.635 $Y=1.635
+ $X2=0 $Y2=0
cc_918 N_SET_B_c_1163_n N_A_1823_524#_c_1617_n 0.00898771f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_919 N_SET_B_c_1163_n N_A_1823_524#_c_1618_n 0.0217366f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_920 SET_B N_A_1823_524#_c_1618_n 3.26663e-19 $X=11.675 $Y=1.58 $X2=0 $Y2=0
cc_921 N_SET_B_c_1167_n N_A_1823_524#_c_1618_n 0.00307419f $X=11.635 $Y=1.635
+ $X2=0 $Y2=0
cc_922 N_SET_B_c_1168_n N_A_1823_524#_c_1618_n 0.0201242f $X=11.635 $Y=1.635
+ $X2=0 $Y2=0
cc_923 N_SET_B_c_1172_n N_A_1823_524#_c_1632_n 0.00408774f $X=11.515 $Y=2.375
+ $X2=0 $Y2=0
cc_924 N_SET_B_c_1173_n N_A_1823_524#_c_1632_n 0.00594531f $X=11.515 $Y=2.465
+ $X2=0 $Y2=0
cc_925 N_SET_B_c_1163_n N_A_1823_524#_c_1632_n 0.0111329f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_926 N_SET_B_c_1168_n N_A_1823_524#_c_1632_n 0.0306884f $X=11.635 $Y=1.635
+ $X2=0 $Y2=0
cc_927 N_SET_B_c_1173_n N_A_1823_524#_c_1633_n 0.00900709f $X=11.515 $Y=2.465
+ $X2=0 $Y2=0
cc_928 N_SET_B_M1038_g N_A_1823_524#_c_1619_n 7.62235e-19 $X=11.6 $Y=0.58 $X2=0
+ $Y2=0
cc_929 SET_B N_A_1823_524#_c_1619_n 0.00749737f $X=11.675 $Y=1.58 $X2=0 $Y2=0
cc_930 N_SET_B_c_1167_n N_A_1823_524#_c_1619_n 2.0927e-19 $X=11.635 $Y=1.635
+ $X2=0 $Y2=0
cc_931 N_SET_B_c_1168_n N_A_1823_524#_c_1619_n 0.0504194f $X=11.635 $Y=1.635
+ $X2=0 $Y2=0
cc_932 N_SET_B_M1038_g N_A_1823_524#_c_1620_n 0.0049566f $X=11.6 $Y=0.58 $X2=0
+ $Y2=0
cc_933 SET_B N_A_1823_524#_c_1620_n 0.00436578f $X=11.675 $Y=1.58 $X2=0 $Y2=0
cc_934 N_SET_B_c_1167_n N_A_1823_524#_c_1620_n 0.0313977f $X=11.635 $Y=1.635
+ $X2=0 $Y2=0
cc_935 N_SET_B_c_1168_n N_A_1823_524#_c_1620_n 0.00363171f $X=11.635 $Y=1.635
+ $X2=0 $Y2=0
cc_936 N_SET_B_c_1172_n N_A_1823_524#_c_1635_n 0.00447942f $X=11.515 $Y=2.375
+ $X2=0 $Y2=0
cc_937 N_SET_B_c_1174_n N_A_1823_524#_c_1635_n 5.47225e-19 $X=11.612 $Y=2.14
+ $X2=0 $Y2=0
cc_938 N_SET_B_c_1172_n N_A_1823_524#_c_1638_n 0.00205401f $X=11.515 $Y=2.375
+ $X2=0 $Y2=0
cc_939 N_SET_B_c_1173_n N_A_1823_524#_c_1638_n 0.00294831f $X=11.515 $Y=2.465
+ $X2=0 $Y2=0
cc_940 N_SET_B_c_1174_n N_A_1823_524#_c_1638_n 0.00135736f $X=11.612 $Y=2.14
+ $X2=0 $Y2=0
cc_941 SET_B N_A_1823_524#_c_1638_n 0.00214435f $X=11.675 $Y=1.58 $X2=0 $Y2=0
cc_942 N_SET_B_c_1171_n N_A_1823_524#_c_1700_n 2.0927e-19 $X=11.612 $Y=1.953
+ $X2=0 $Y2=0
cc_943 N_SET_B_c_1170_n N_VPWR_c_1953_n 0.00153105f $X=7.345 $Y=2.21 $X2=0 $Y2=0
cc_944 N_SET_B_c_1163_n N_VPWR_c_1953_n 3.62696e-19 $X=11.615 $Y=1.665 $X2=0
+ $Y2=0
cc_945 N_SET_B_c_1173_n N_VPWR_c_1955_n 0.00402106f $X=11.515 $Y=2.465 $X2=0
+ $Y2=0
cc_946 N_SET_B_c_1173_n N_VPWR_c_1969_n 0.00445602f $X=11.515 $Y=2.465 $X2=0
+ $Y2=0
cc_947 N_SET_B_c_1173_n N_VPWR_c_1947_n 0.0046151f $X=11.515 $Y=2.465 $X2=0
+ $Y2=0
cc_948 N_SET_B_c_1163_n N_A_1620_373#_c_2290_n 0.00155961f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_949 N_SET_B_M1003_g N_VGND_c_2419_n 0.0184827f $X=7.54 $Y=0.58 $X2=0 $Y2=0
cc_950 N_SET_B_M1038_g N_VGND_c_2421_n 0.0175686f $X=11.6 $Y=0.58 $X2=0 $Y2=0
cc_951 N_SET_B_M1003_g N_VGND_c_2431_n 0.00383152f $X=7.54 $Y=0.58 $X2=0 $Y2=0
cc_952 N_SET_B_M1038_g N_VGND_c_2433_n 0.00383152f $X=11.6 $Y=0.58 $X2=0 $Y2=0
cc_953 N_SET_B_M1003_g N_VGND_c_2444_n 0.0075725f $X=7.54 $Y=0.58 $X2=0 $Y2=0
cc_954 N_SET_B_M1038_g N_VGND_c_2444_n 0.00758569f $X=11.6 $Y=0.58 $X2=0 $Y2=0
cc_955 N_SET_B_c_1163_n N_A_1677_74#_c_2591_n 0.0287108f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_956 N_SET_B_c_1163_n N_A_1677_74#_c_2592_n 0.00399518f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_957 N_A_616_74#_M1026_g N_A_2191_180#_c_1504_n 0.0210257f $X=10.67 $Y=0.58
+ $X2=0 $Y2=0
cc_958 N_A_616_74#_M1026_g N_A_2191_180#_c_1508_n 0.00116793f $X=10.67 $Y=0.58
+ $X2=0 $Y2=0
cc_959 N_A_616_74#_M1026_g N_A_2191_180#_c_1509_n 0.0197474f $X=10.67 $Y=0.58
+ $X2=0 $Y2=0
cc_960 N_A_616_74#_M1026_g N_A_2191_180#_c_1511_n 0.0358279f $X=10.67 $Y=0.58
+ $X2=0 $Y2=0
cc_961 N_A_616_74#_c_1324_n N_A_1823_524#_c_1628_n 4.52794e-19 $X=9.395 $Y=3.15
+ $X2=0 $Y2=0
cc_962 N_A_616_74#_c_1325_n N_A_1823_524#_c_1628_n 0.00948523f $X=9.485 $Y=3.035
+ $X2=0 $Y2=0
cc_963 N_A_616_74#_c_1326_n N_A_1823_524#_c_1628_n 0.0100692f $X=9.845 $Y=3.15
+ $X2=0 $Y2=0
cc_964 N_A_616_74#_M1030_g N_A_1823_524#_c_1628_n 0.0133297f $X=9.935 $Y=2.54
+ $X2=0 $Y2=0
cc_965 N_A_616_74#_c_1333_n N_A_1823_524#_c_1628_n 0.0037543f $X=9.485 $Y=3.13
+ $X2=0 $Y2=0
cc_966 N_A_616_74#_M1026_g N_A_1823_524#_c_1613_n 0.00401774f $X=10.67 $Y=0.58
+ $X2=0 $Y2=0
cc_967 N_A_616_74#_M1026_g N_A_1823_524#_c_1615_n 0.0160978f $X=10.67 $Y=0.58
+ $X2=0 $Y2=0
cc_968 N_A_616_74#_c_1310_n N_A_1823_524#_c_1616_n 0.0054437f $X=10.595 $Y=1.52
+ $X2=0 $Y2=0
cc_969 N_A_616_74#_M1026_g N_A_1823_524#_c_1616_n 0.00857875f $X=10.67 $Y=0.58
+ $X2=0 $Y2=0
cc_970 N_A_616_74#_c_1310_n N_A_1823_524#_c_1617_n 0.0191332f $X=10.595 $Y=1.52
+ $X2=0 $Y2=0
cc_971 N_A_616_74#_c_1310_n N_A_1823_524#_c_1618_n 5.03394e-19 $X=10.595 $Y=1.52
+ $X2=0 $Y2=0
cc_972 N_A_616_74#_c_1324_n N_A_1823_524#_c_1636_n 0.00676385f $X=9.395 $Y=3.15
+ $X2=0 $Y2=0
cc_973 N_A_616_74#_c_1325_n N_A_1823_524#_c_1636_n 8.1772e-19 $X=9.485 $Y=3.035
+ $X2=0 $Y2=0
cc_974 N_A_616_74#_c_1333_n N_A_1823_524#_c_1636_n 5.49707e-19 $X=9.485 $Y=3.13
+ $X2=0 $Y2=0
cc_975 N_A_616_74#_c_1335_n N_VPWR_M1028_d 0.00200574f $X=3.885 $Y=1.945 $X2=0
+ $Y2=0
cc_976 N_A_616_74#_c_1317_n N_VPWR_c_1951_n 0.00730018f $X=3.96 $Y=1.765 $X2=0
+ $Y2=0
cc_977 N_A_616_74#_c_1322_n N_VPWR_c_1951_n 0.00213268f $X=4.605 $Y=3.15 $X2=0
+ $Y2=0
cc_978 N_A_616_74#_c_1323_n N_VPWR_c_1952_n 7.32825e-19 $X=5.625 $Y=2.97 $X2=0
+ $Y2=0
cc_979 N_A_616_74#_c_1324_n N_VPWR_c_1952_n 0.0211091f $X=9.395 $Y=3.15 $X2=0
+ $Y2=0
cc_980 N_A_616_74#_c_1332_n N_VPWR_c_1952_n 7.10913e-19 $X=5.625 $Y=3.15 $X2=0
+ $Y2=0
cc_981 N_A_616_74#_c_1324_n N_VPWR_c_1953_n 0.0163491f $X=9.395 $Y=3.15 $X2=0
+ $Y2=0
cc_982 N_A_616_74#_c_1324_n N_VPWR_c_1954_n 0.0249704f $X=9.395 $Y=3.15 $X2=0
+ $Y2=0
cc_983 N_A_616_74#_c_1325_n N_VPWR_c_1954_n 0.00389954f $X=9.485 $Y=3.035 $X2=0
+ $Y2=0
cc_984 N_A_616_74#_c_1324_n N_VPWR_c_1961_n 0.0291914f $X=9.395 $Y=3.15 $X2=0
+ $Y2=0
cc_985 N_A_616_74#_c_1324_n N_VPWR_c_1963_n 0.0198799f $X=9.395 $Y=3.15 $X2=0
+ $Y2=0
cc_986 N_A_616_74#_c_1317_n N_VPWR_c_1967_n 0.00413917f $X=3.96 $Y=1.765 $X2=0
+ $Y2=0
cc_987 N_A_616_74#_c_1322_n N_VPWR_c_1967_n 0.044661f $X=4.605 $Y=3.15 $X2=0
+ $Y2=0
cc_988 N_A_616_74#_c_1324_n N_VPWR_c_1968_n 0.0279463f $X=9.395 $Y=3.15 $X2=0
+ $Y2=0
cc_989 N_A_616_74#_c_1317_n N_VPWR_c_1947_n 0.00818763f $X=3.96 $Y=1.765 $X2=0
+ $Y2=0
cc_990 N_A_616_74#_c_1321_n N_VPWR_c_1947_n 0.0216332f $X=5.535 $Y=3.15 $X2=0
+ $Y2=0
cc_991 N_A_616_74#_c_1322_n N_VPWR_c_1947_n 0.00600633f $X=4.605 $Y=3.15 $X2=0
+ $Y2=0
cc_992 N_A_616_74#_c_1324_n N_VPWR_c_1947_n 0.101935f $X=9.395 $Y=3.15 $X2=0
+ $Y2=0
cc_993 N_A_616_74#_c_1326_n N_VPWR_c_1947_n 0.0129445f $X=9.845 $Y=3.15 $X2=0
+ $Y2=0
cc_994 N_A_616_74#_c_1332_n N_VPWR_c_1947_n 0.00441257f $X=5.625 $Y=3.15 $X2=0
+ $Y2=0
cc_995 N_A_616_74#_c_1333_n N_VPWR_c_1947_n 0.00440873f $X=9.485 $Y=3.13 $X2=0
+ $Y2=0
cc_996 N_A_616_74#_c_1316_n N_A_288_464#_c_2162_n 0.00517647f $X=3.197 $Y=1.01
+ $X2=0 $Y2=0
cc_997 N_A_616_74#_c_1314_n N_A_288_464#_c_2164_n 5.13943e-19 $X=3.09 $Y=1.82
+ $X2=0 $Y2=0
cc_998 N_A_616_74#_M1028_s N_A_288_464#_c_2169_n 0.0110751f $X=3.14 $Y=1.84
+ $X2=0 $Y2=0
cc_999 N_A_616_74#_c_1317_n N_A_288_464#_c_2169_n 0.0154002f $X=3.96 $Y=1.765
+ $X2=0 $Y2=0
cc_1000 N_A_616_74#_c_1306_n N_A_288_464#_c_2169_n 0.00471966f $X=4.45 $Y=1.68
+ $X2=0 $Y2=0
cc_1001 N_A_616_74#_c_1331_n N_A_288_464#_c_2169_n 0.0015154f $X=4.53 $Y=2.045
+ $X2=0 $Y2=0
cc_1002 N_A_616_74#_c_1335_n N_A_288_464#_c_2169_n 0.0609561f $X=3.885 $Y=1.945
+ $X2=0 $Y2=0
cc_1003 N_A_616_74#_M1021_g N_A_288_464#_c_2165_n 0.00124454f $X=3.94 $Y=0.74
+ $X2=0 $Y2=0
cc_1004 N_A_616_74#_c_1305_n N_A_288_464#_c_2165_n 0.00634768f $X=4.45 $Y=1.35
+ $X2=0 $Y2=0
cc_1005 N_A_616_74#_c_1306_n N_A_288_464#_c_2165_n 0.0100578f $X=4.45 $Y=1.68
+ $X2=0 $Y2=0
cc_1006 N_A_616_74#_c_1319_n N_A_288_464#_c_2165_n 0.00523979f $X=4.45 $Y=1.97
+ $X2=0 $Y2=0
cc_1007 N_A_616_74#_c_1307_n N_A_288_464#_c_2165_n 0.00539182f $X=4.935 $Y=1.115
+ $X2=0 $Y2=0
cc_1008 N_A_616_74#_c_1308_n N_A_288_464#_c_2165_n 0.00485757f $X=4.525 $Y=1.115
+ $X2=0 $Y2=0
cc_1009 N_A_616_74#_M1002_g N_A_288_464#_c_2165_n 0.00195875f $X=5.01 $Y=0.615
+ $X2=0 $Y2=0
cc_1010 N_A_616_74#_c_1335_n N_A_288_464#_c_2165_n 0.00568568f $X=3.885 $Y=1.945
+ $X2=0 $Y2=0
cc_1011 N_A_616_74#_c_1315_n N_A_288_464#_c_2165_n 0.0305869f $X=4.05 $Y=1.515
+ $X2=0 $Y2=0
cc_1012 N_A_616_74#_M1028_s N_A_288_464#_c_2171_n 0.00532576f $X=3.14 $Y=1.84
+ $X2=0 $Y2=0
cc_1013 N_A_616_74#_c_1336_n N_A_288_464#_c_2171_n 0.0150765f $X=3.175 $Y=1.945
+ $X2=0 $Y2=0
cc_1014 N_A_616_74#_c_1307_n N_A_288_464#_c_2166_n 0.00779105f $X=4.935 $Y=1.115
+ $X2=0 $Y2=0
cc_1015 N_A_616_74#_c_1308_n N_A_288_464#_c_2166_n 0.00100653f $X=4.525 $Y=1.115
+ $X2=0 $Y2=0
cc_1016 N_A_616_74#_M1002_g N_A_288_464#_c_2166_n 0.00669516f $X=5.01 $Y=0.615
+ $X2=0 $Y2=0
cc_1017 N_A_616_74#_c_1317_n N_A_288_464#_c_2172_n 0.00308619f $X=3.96 $Y=1.765
+ $X2=0 $Y2=0
cc_1018 N_A_616_74#_c_1319_n N_A_288_464#_c_2172_n 0.00233833f $X=4.45 $Y=1.97
+ $X2=0 $Y2=0
cc_1019 N_A_616_74#_c_1320_n N_A_288_464#_c_2172_n 0.0221984f $X=4.53 $Y=3.075
+ $X2=0 $Y2=0
cc_1020 N_A_616_74#_c_1331_n N_A_288_464#_c_2172_n 0.00913348f $X=4.53 $Y=2.045
+ $X2=0 $Y2=0
cc_1021 N_A_616_74#_c_1335_n N_A_288_464#_c_2172_n 0.0132248f $X=3.885 $Y=1.945
+ $X2=0 $Y2=0
cc_1022 N_A_616_74#_c_1324_n N_A_1620_373#_c_2289_n 0.00517428f $X=9.395 $Y=3.15
+ $X2=0 $Y2=0
cc_1023 N_A_616_74#_c_1325_n N_A_1620_373#_c_2290_n 0.0109343f $X=9.485 $Y=3.035
+ $X2=0 $Y2=0
cc_1024 N_A_616_74#_c_1325_n N_A_1620_373#_c_2291_n 0.0156533f $X=9.485 $Y=3.035
+ $X2=0 $Y2=0
cc_1025 N_A_616_74#_c_1328_n N_A_1620_373#_c_2291_n 4.24894e-19 $X=9.935
+ $Y=2.045 $X2=0 $Y2=0
cc_1026 N_A_616_74#_M1030_g N_A_1620_373#_c_2291_n 0.00831143f $X=9.935 $Y=2.54
+ $X2=0 $Y2=0
cc_1027 N_A_616_74#_c_1313_n N_VGND_c_2415_n 0.0270111f $X=3.225 $Y=0.515 $X2=0
+ $Y2=0
cc_1028 N_A_616_74#_c_1313_n N_VGND_c_2416_n 0.0169976f $X=3.225 $Y=0.515 $X2=0
+ $Y2=0
cc_1029 N_A_616_74#_M1021_g N_VGND_c_2417_n 0.0120466f $X=3.94 $Y=0.74 $X2=0
+ $Y2=0
cc_1030 N_A_616_74#_c_1313_n N_VGND_c_2417_n 0.026108f $X=3.225 $Y=0.515 $X2=0
+ $Y2=0
cc_1031 N_A_616_74#_M1021_g N_VGND_c_2430_n 0.00383152f $X=3.94 $Y=0.74 $X2=0
+ $Y2=0
cc_1032 N_A_616_74#_M1002_g N_VGND_c_2430_n 9.34059e-19 $X=5.01 $Y=0.615 $X2=0
+ $Y2=0
cc_1033 N_A_616_74#_M1026_g N_VGND_c_2433_n 0.00461464f $X=10.67 $Y=0.58 $X2=0
+ $Y2=0
cc_1034 N_A_616_74#_M1021_g N_VGND_c_2444_n 0.00762539f $X=3.94 $Y=0.74 $X2=0
+ $Y2=0
cc_1035 N_A_616_74#_M1026_g N_VGND_c_2444_n 0.00909821f $X=10.67 $Y=0.58 $X2=0
+ $Y2=0
cc_1036 N_A_616_74#_c_1313_n N_VGND_c_2444_n 0.0140217f $X=3.225 $Y=0.515 $X2=0
+ $Y2=0
cc_1037 N_A_616_74#_c_1311_n N_A_1677_74#_c_2591_n 0.00197309f $X=10.025 $Y=1.52
+ $X2=0 $Y2=0
cc_1038 N_A_2191_180#_c_1505_n N_A_1823_524#_M1039_g 0.0124612f $X=12.32
+ $Y=0.985 $X2=0 $Y2=0
cc_1039 N_A_2191_180#_c_1506_n N_A_1823_524#_M1039_g 0.0119097f $X=12.485
+ $Y=0.58 $X2=0 $Y2=0
cc_1040 N_A_2191_180#_c_1507_n N_A_1823_524#_M1039_g 0.00896473f $X=12.625
+ $Y=2.18 $X2=0 $Y2=0
cc_1041 N_A_2191_180#_c_1510_n N_A_1823_524#_M1039_g 0.00442658f $X=12.515
+ $Y=0.985 $X2=0 $Y2=0
cc_1042 N_A_2191_180#_c_1514_n N_A_1823_524#_c_1621_n 0.00134849f $X=12.465
+ $Y=2.65 $X2=0 $Y2=0
cc_1043 N_A_2191_180#_c_1507_n N_A_1823_524#_c_1621_n 0.00390512f $X=12.625
+ $Y=2.18 $X2=0 $Y2=0
cc_1044 N_A_2191_180#_c_1517_n N_A_1823_524#_c_1621_n 0.0146625f $X=12.625
+ $Y=2.265 $X2=0 $Y2=0
cc_1045 N_A_2191_180#_c_1514_n N_A_1823_524#_c_1622_n 0.0102336f $X=12.465
+ $Y=2.65 $X2=0 $Y2=0
cc_1046 N_A_2191_180#_c_1516_n N_A_1823_524#_c_1622_n 0.00665776f $X=12.465
+ $Y=2.815 $X2=0 $Y2=0
cc_1047 N_A_2191_180#_c_1507_n N_A_1823_524#_c_1623_n 0.00638826f $X=12.625
+ $Y=2.18 $X2=0 $Y2=0
cc_1048 N_A_2191_180#_c_1517_n N_A_1823_524#_c_1623_n 4.98011e-19 $X=12.625
+ $Y=2.265 $X2=0 $Y2=0
cc_1049 N_A_2191_180#_c_1514_n N_A_1823_524#_c_1624_n 6.52737e-19 $X=12.465
+ $Y=2.65 $X2=0 $Y2=0
cc_1050 N_A_2191_180#_c_1507_n N_A_1823_524#_c_1624_n 0.00108095f $X=12.625
+ $Y=2.18 $X2=0 $Y2=0
cc_1051 N_A_2191_180#_c_1517_n N_A_1823_524#_c_1624_n 0.00147908f $X=12.625
+ $Y=2.265 $X2=0 $Y2=0
cc_1052 N_A_2191_180#_c_1506_n N_A_1823_524#_M1008_g 0.00102192f $X=12.485
+ $Y=0.58 $X2=0 $Y2=0
cc_1053 N_A_2191_180#_c_1507_n N_A_1823_524#_M1008_g 0.00270972f $X=12.625
+ $Y=2.18 $X2=0 $Y2=0
cc_1054 N_A_2191_180#_c_1513_n N_A_1823_524#_c_1628_n 4.31891e-19 $X=11.065
+ $Y=2.465 $X2=0 $Y2=0
cc_1055 N_A_2191_180#_c_1513_n N_A_1823_524#_c_1647_n 7.72678e-19 $X=11.065
+ $Y=2.465 $X2=0 $Y2=0
cc_1056 N_A_2191_180#_c_1508_n N_A_1823_524#_c_1615_n 0.0133926f $X=11.12
+ $Y=0.985 $X2=0 $Y2=0
cc_1057 N_A_2191_180#_c_1504_n N_A_1823_524#_c_1616_n 0.00784384f $X=11.065
+ $Y=2.375 $X2=0 $Y2=0
cc_1058 N_A_2191_180#_c_1508_n N_A_1823_524#_c_1616_n 0.0114201f $X=11.12
+ $Y=0.985 $X2=0 $Y2=0
cc_1059 N_A_2191_180#_c_1504_n N_A_1823_524#_c_1618_n 0.0216535f $X=11.065
+ $Y=2.375 $X2=0 $Y2=0
cc_1060 N_A_2191_180#_c_1504_n N_A_1823_524#_c_1632_n 0.00216439f $X=11.065
+ $Y=2.375 $X2=0 $Y2=0
cc_1061 N_A_2191_180#_c_1513_n N_A_1823_524#_c_1632_n 0.00250678f $X=11.065
+ $Y=2.465 $X2=0 $Y2=0
cc_1062 N_A_2191_180#_c_1513_n N_A_1823_524#_c_1633_n 8.50792e-19 $X=11.065
+ $Y=2.465 $X2=0 $Y2=0
cc_1063 N_A_2191_180#_c_1514_n N_A_1823_524#_c_1633_n 0.00645614f $X=12.465
+ $Y=2.65 $X2=0 $Y2=0
cc_1064 N_A_2191_180#_c_1516_n N_A_1823_524#_c_1633_n 0.0225794f $X=12.465
+ $Y=2.815 $X2=0 $Y2=0
cc_1065 N_A_2191_180#_c_1505_n N_A_1823_524#_c_1619_n 0.0152233f $X=12.32
+ $Y=0.985 $X2=0 $Y2=0
cc_1066 N_A_2191_180#_c_1507_n N_A_1823_524#_c_1619_n 0.0478089f $X=12.625
+ $Y=2.18 $X2=0 $Y2=0
cc_1067 N_A_2191_180#_c_1510_n N_A_1823_524#_c_1619_n 0.0029784f $X=12.515
+ $Y=0.985 $X2=0 $Y2=0
cc_1068 N_A_2191_180#_c_1505_n N_A_1823_524#_c_1620_n 9.74505e-19 $X=12.32
+ $Y=0.985 $X2=0 $Y2=0
cc_1069 N_A_2191_180#_c_1507_n N_A_1823_524#_c_1620_n 0.0225871f $X=12.625
+ $Y=2.18 $X2=0 $Y2=0
cc_1070 N_A_2191_180#_c_1516_n N_A_1823_524#_c_1620_n 0.0033637f $X=12.465
+ $Y=2.815 $X2=0 $Y2=0
cc_1071 N_A_2191_180#_c_1510_n N_A_1823_524#_c_1620_n 0.00760198f $X=12.515
+ $Y=0.985 $X2=0 $Y2=0
cc_1072 N_A_2191_180#_c_1517_n N_A_1823_524#_c_1620_n 0.00234945f $X=12.625
+ $Y=2.265 $X2=0 $Y2=0
cc_1073 N_A_2191_180#_c_1507_n N_A_1823_524#_c_1635_n 0.00726945f $X=12.625
+ $Y=2.18 $X2=0 $Y2=0
cc_1074 N_A_2191_180#_c_1517_n N_A_1823_524#_c_1635_n 0.0102741f $X=12.625
+ $Y=2.265 $X2=0 $Y2=0
cc_1075 N_A_2191_180#_c_1504_n N_A_1823_524#_c_1637_n 0.00183584f $X=11.065
+ $Y=2.375 $X2=0 $Y2=0
cc_1076 N_A_2191_180#_c_1513_n N_A_1823_524#_c_1637_n 0.00631033f $X=11.065
+ $Y=2.465 $X2=0 $Y2=0
cc_1077 N_A_2191_180#_c_1514_n N_A_1823_524#_c_1638_n 0.0108937f $X=12.465
+ $Y=2.65 $X2=0 $Y2=0
cc_1078 N_A_2191_180#_c_1516_n N_A_1823_524#_c_1638_n 0.00572708f $X=12.465
+ $Y=2.815 $X2=0 $Y2=0
cc_1079 N_A_2191_180#_c_1517_n N_A_1823_524#_c_1638_n 0.00337662f $X=12.625
+ $Y=2.265 $X2=0 $Y2=0
cc_1080 N_A_2191_180#_c_1516_n N_A_1823_524#_c_1700_n 0.0045697f $X=12.465
+ $Y=2.815 $X2=0 $Y2=0
cc_1081 N_A_2191_180#_c_1506_n N_A_2580_74#_c_1834_n 0.0463408f $X=12.485
+ $Y=0.58 $X2=0 $Y2=0
cc_1082 N_A_2191_180#_c_1507_n N_A_2580_74#_c_1834_n 0.0197418f $X=12.625
+ $Y=2.18 $X2=0 $Y2=0
cc_1083 N_A_2191_180#_c_1510_n N_A_2580_74#_c_1834_n 0.0150382f $X=12.515
+ $Y=0.985 $X2=0 $Y2=0
cc_1084 N_A_2191_180#_c_1514_n N_A_2580_74#_c_1835_n 0.0042639f $X=12.465
+ $Y=2.65 $X2=0 $Y2=0
cc_1085 N_A_2191_180#_c_1507_n N_A_2580_74#_c_1835_n 0.0186863f $X=12.625
+ $Y=2.18 $X2=0 $Y2=0
cc_1086 N_A_2191_180#_c_1517_n N_A_2580_74#_c_1835_n 0.00615389f $X=12.625
+ $Y=2.265 $X2=0 $Y2=0
cc_1087 N_A_2191_180#_c_1507_n N_A_2580_74#_c_1837_n 0.0211268f $X=12.625
+ $Y=2.18 $X2=0 $Y2=0
cc_1088 N_A_2191_180#_c_1507_n N_VPWR_M1013_d 8.41796e-19 $X=12.625 $Y=2.18
+ $X2=0 $Y2=0
cc_1089 N_A_2191_180#_c_1517_n N_VPWR_M1013_d 0.00301745f $X=12.625 $Y=2.265
+ $X2=0 $Y2=0
cc_1090 N_A_2191_180#_c_1513_n N_VPWR_c_1955_n 0.00711873f $X=11.065 $Y=2.465
+ $X2=0 $Y2=0
cc_1091 N_A_2191_180#_c_1514_n N_VPWR_c_1956_n 0.00940733f $X=12.465 $Y=2.65
+ $X2=0 $Y2=0
cc_1092 N_A_2191_180#_c_1516_n N_VPWR_c_1956_n 0.0255186f $X=12.465 $Y=2.815
+ $X2=0 $Y2=0
cc_1093 N_A_2191_180#_c_1513_n N_VPWR_c_1968_n 0.00413917f $X=11.065 $Y=2.465
+ $X2=0 $Y2=0
cc_1094 N_A_2191_180#_c_1516_n N_VPWR_c_1969_n 0.0172262f $X=12.465 $Y=2.815
+ $X2=0 $Y2=0
cc_1095 N_A_2191_180#_c_1513_n N_VPWR_c_1947_n 0.00418005f $X=11.065 $Y=2.465
+ $X2=0 $Y2=0
cc_1096 N_A_2191_180#_c_1516_n N_VPWR_c_1947_n 0.0144762f $X=12.465 $Y=2.815
+ $X2=0 $Y2=0
cc_1097 N_A_2191_180#_c_1513_n A_2103_508# 0.00231449f $X=11.065 $Y=2.465
+ $X2=-0.19 $Y2=-0.245
cc_1098 N_A_2191_180#_c_1505_n N_VGND_c_2421_n 0.0314789f $X=12.32 $Y=0.985
+ $X2=0 $Y2=0
cc_1099 N_A_2191_180#_c_1506_n N_VGND_c_2421_n 0.0135447f $X=12.485 $Y=0.58
+ $X2=0 $Y2=0
cc_1100 N_A_2191_180#_c_1511_n N_VGND_c_2421_n 0.00204005f $X=11.12 $Y=0.9 $X2=0
+ $Y2=0
cc_1101 N_A_2191_180#_c_1506_n N_VGND_c_2426_n 0.0172816f $X=12.485 $Y=0.58
+ $X2=0 $Y2=0
cc_1102 N_A_2191_180#_c_1511_n N_VGND_c_2433_n 0.00461464f $X=11.12 $Y=0.9 $X2=0
+ $Y2=0
cc_1103 N_A_2191_180#_c_1506_n N_VGND_c_2444_n 0.0142302f $X=12.485 $Y=0.58
+ $X2=0 $Y2=0
cc_1104 N_A_2191_180#_c_1511_n N_VGND_c_2444_n 0.00910057f $X=11.12 $Y=0.9 $X2=0
+ $Y2=0
cc_1105 N_A_1823_524#_M1008_g N_A_2580_74#_M1000_g 0.0327036f $X=13.26 $Y=0.74
+ $X2=0 $Y2=0
cc_1106 N_A_1823_524#_M1008_g N_A_2580_74#_c_1838_n 0.00190507f $X=13.26 $Y=0.74
+ $X2=0 $Y2=0
cc_1107 N_A_1823_524#_c_1626_n N_A_2580_74#_c_1838_n 0.0190051f $X=13.48
+ $Y=2.045 $X2=0 $Y2=0
cc_1108 N_A_1823_524#_c_1627_n N_A_2580_74#_c_1838_n 0.00577778f $X=13.26
+ $Y=1.967 $X2=0 $Y2=0
cc_1109 N_A_1823_524#_M1008_g N_A_2580_74#_c_1830_n 0.00187313f $X=13.26 $Y=0.74
+ $X2=0 $Y2=0
cc_1110 N_A_1823_524#_M1039_g N_A_2580_74#_c_1834_n 0.00167283f $X=12.27 $Y=0.58
+ $X2=0 $Y2=0
cc_1111 N_A_1823_524#_M1008_g N_A_2580_74#_c_1834_n 0.0176758f $X=13.26 $Y=0.74
+ $X2=0 $Y2=0
cc_1112 N_A_1823_524#_c_1624_n N_A_2580_74#_c_1835_n 0.00595084f $X=13.03
+ $Y=2.045 $X2=0 $Y2=0
cc_1113 N_A_1823_524#_M1008_g N_A_2580_74#_c_1835_n 0.00732029f $X=13.26 $Y=0.74
+ $X2=0 $Y2=0
cc_1114 N_A_1823_524#_c_1626_n N_A_2580_74#_c_1835_n 0.00495772f $X=13.48
+ $Y=2.045 $X2=0 $Y2=0
cc_1115 N_A_1823_524#_c_1627_n N_A_2580_74#_c_1835_n 0.0128793f $X=13.26
+ $Y=1.967 $X2=0 $Y2=0
cc_1116 N_A_1823_524#_c_1620_n N_A_2580_74#_c_1835_n 7.80167e-19 $X=12.205
+ $Y=1.505 $X2=0 $Y2=0
cc_1117 N_A_1823_524#_c_1627_n N_A_2580_74#_c_1836_n 0.00852046f $X=13.26
+ $Y=1.967 $X2=0 $Y2=0
cc_1118 N_A_1823_524#_c_1623_n N_A_2580_74#_c_1837_n 0.00771468f $X=12.94
+ $Y=1.965 $X2=0 $Y2=0
cc_1119 N_A_1823_524#_M1008_g N_A_2580_74#_c_1837_n 0.0198504f $X=13.26 $Y=0.74
+ $X2=0 $Y2=0
cc_1120 N_A_1823_524#_c_1620_n N_A_2580_74#_c_1837_n 0.00125585f $X=12.205
+ $Y=1.505 $X2=0 $Y2=0
cc_1121 N_A_1823_524#_c_1636_n N_VPWR_c_1954_n 0.0316308f $X=9.26 $Y=2.79 $X2=0
+ $Y2=0
cc_1122 N_A_1823_524#_c_1632_n N_VPWR_c_1955_n 0.0173769f $X=11.575 $Y=2.395
+ $X2=0 $Y2=0
cc_1123 N_A_1823_524#_c_1633_n N_VPWR_c_1955_n 0.0221564f $X=11.74 $Y=2.75 $X2=0
+ $Y2=0
cc_1124 N_A_1823_524#_c_1622_n N_VPWR_c_1956_n 0.00601163f $X=12.525 $Y=2.465
+ $X2=0 $Y2=0
cc_1125 N_A_1823_524#_c_1623_n N_VPWR_c_1956_n 0.00575399f $X=12.94 $Y=1.965
+ $X2=0 $Y2=0
cc_1126 N_A_1823_524#_c_1624_n N_VPWR_c_1956_n 0.0095306f $X=13.03 $Y=2.045
+ $X2=0 $Y2=0
cc_1127 N_A_1823_524#_c_1626_n N_VPWR_c_1956_n 4.674e-19 $X=13.48 $Y=2.045 $X2=0
+ $Y2=0
cc_1128 N_A_1823_524#_c_1624_n N_VPWR_c_1957_n 5.9374e-19 $X=13.03 $Y=2.045
+ $X2=0 $Y2=0
cc_1129 N_A_1823_524#_c_1626_n N_VPWR_c_1957_n 0.0151699f $X=13.48 $Y=2.045
+ $X2=0 $Y2=0
cc_1130 N_A_1823_524#_c_1627_n N_VPWR_c_1957_n 4.25443e-19 $X=13.26 $Y=1.967
+ $X2=0 $Y2=0
cc_1131 N_A_1823_524#_c_1628_n N_VPWR_c_1968_n 0.0663726f $X=10.045 $Y=2.967
+ $X2=0 $Y2=0
cc_1132 N_A_1823_524#_c_1636_n N_VPWR_c_1968_n 0.018469f $X=9.26 $Y=2.79 $X2=0
+ $Y2=0
cc_1133 N_A_1823_524#_c_1622_n N_VPWR_c_1969_n 0.00348254f $X=12.525 $Y=2.465
+ $X2=0 $Y2=0
cc_1134 N_A_1823_524#_c_1633_n N_VPWR_c_1969_n 0.014274f $X=11.74 $Y=2.75 $X2=0
+ $Y2=0
cc_1135 N_A_1823_524#_c_1624_n N_VPWR_c_1970_n 0.00413917f $X=13.03 $Y=2.045
+ $X2=0 $Y2=0
cc_1136 N_A_1823_524#_c_1626_n N_VPWR_c_1970_n 0.00413917f $X=13.48 $Y=2.045
+ $X2=0 $Y2=0
cc_1137 N_A_1823_524#_c_1622_n N_VPWR_c_1947_n 0.00585102f $X=12.525 $Y=2.465
+ $X2=0 $Y2=0
cc_1138 N_A_1823_524#_c_1624_n N_VPWR_c_1947_n 0.00817726f $X=13.03 $Y=2.045
+ $X2=0 $Y2=0
cc_1139 N_A_1823_524#_c_1626_n N_VPWR_c_1947_n 0.00817726f $X=13.48 $Y=2.045
+ $X2=0 $Y2=0
cc_1140 N_A_1823_524#_c_1628_n N_VPWR_c_1947_n 0.035213f $X=10.045 $Y=2.967
+ $X2=0 $Y2=0
cc_1141 N_A_1823_524#_c_1629_n N_VPWR_c_1947_n 0.00535163f $X=10.935 $Y=2.395
+ $X2=0 $Y2=0
cc_1142 N_A_1823_524#_c_1632_n N_VPWR_c_1947_n 0.0152923f $X=11.575 $Y=2.395
+ $X2=0 $Y2=0
cc_1143 N_A_1823_524#_c_1633_n N_VPWR_c_1947_n 0.011923f $X=11.74 $Y=2.75 $X2=0
+ $Y2=0
cc_1144 N_A_1823_524#_c_1636_n N_VPWR_c_1947_n 0.00943811f $X=9.26 $Y=2.79 $X2=0
+ $Y2=0
cc_1145 N_A_1823_524#_c_1637_n N_VPWR_c_1947_n 0.00501343f $X=11.02 $Y=2.395
+ $X2=0 $Y2=0
cc_1146 N_A_1823_524#_c_1628_n N_A_1620_373#_M1016_d 0.00199159f $X=10.045
+ $Y=2.967 $X2=0 $Y2=0
cc_1147 N_A_1823_524#_M1016_s N_A_1620_373#_c_2290_n 0.00549258f $X=9.115
+ $Y=2.62 $X2=0 $Y2=0
cc_1148 N_A_1823_524#_c_1628_n N_A_1620_373#_c_2290_n 0.00341576f $X=10.045
+ $Y=2.967 $X2=0 $Y2=0
cc_1149 N_A_1823_524#_c_1636_n N_A_1620_373#_c_2290_n 0.0131939f $X=9.26 $Y=2.79
+ $X2=0 $Y2=0
cc_1150 N_A_1823_524#_c_1628_n N_A_1620_373#_c_2291_n 0.0162931f $X=10.045
+ $Y=2.967 $X2=0 $Y2=0
cc_1151 N_A_1823_524#_c_1628_n A_2103_508# 0.00581768f $X=10.045 $Y=2.967
+ $X2=-0.19 $Y2=-0.245
cc_1152 N_A_1823_524#_c_1629_n A_2103_508# 0.0284228f $X=10.935 $Y=2.395
+ $X2=-0.19 $Y2=-0.245
cc_1153 N_A_1823_524#_c_1626_n N_Q_c_2339_n 2.70969e-19 $X=13.48 $Y=2.045 $X2=0
+ $Y2=0
cc_1154 N_A_1823_524#_c_1627_n N_Q_c_2339_n 8.6525e-19 $X=13.26 $Y=1.967 $X2=0
+ $Y2=0
cc_1155 N_A_1823_524#_c_1626_n N_Q_c_2340_n 2.75868e-19 $X=13.48 $Y=2.045 $X2=0
+ $Y2=0
cc_1156 N_A_1823_524#_c_1612_n N_VGND_c_2420_n 0.0346868f $X=9.515 $Y=0.515
+ $X2=0 $Y2=0
cc_1157 N_A_1823_524#_c_1614_n N_VGND_c_2420_n 0.0121616f $X=9.68 $Y=0.34 $X2=0
+ $Y2=0
cc_1158 N_A_1823_524#_M1039_g N_VGND_c_2421_n 0.00600886f $X=12.27 $Y=0.58 $X2=0
+ $Y2=0
cc_1159 N_A_1823_524#_M1008_g N_VGND_c_2422_n 0.00728495f $X=13.26 $Y=0.74 $X2=0
+ $Y2=0
cc_1160 N_A_1823_524#_M1039_g N_VGND_c_2426_n 0.00434272f $X=12.27 $Y=0.58 $X2=0
+ $Y2=0
cc_1161 N_A_1823_524#_M1008_g N_VGND_c_2426_n 0.00434272f $X=13.26 $Y=0.74 $X2=0
+ $Y2=0
cc_1162 N_A_1823_524#_c_1613_n N_VGND_c_2433_n 0.0569302f $X=10.21 $Y=0.34 $X2=0
+ $Y2=0
cc_1163 N_A_1823_524#_c_1614_n N_VGND_c_2433_n 0.0235818f $X=9.68 $Y=0.34 $X2=0
+ $Y2=0
cc_1164 N_A_1823_524#_M1039_g N_VGND_c_2444_n 0.00826973f $X=12.27 $Y=0.58 $X2=0
+ $Y2=0
cc_1165 N_A_1823_524#_M1008_g N_VGND_c_2444_n 0.00825771f $X=13.26 $Y=0.74 $X2=0
+ $Y2=0
cc_1166 N_A_1823_524#_c_1613_n N_VGND_c_2444_n 0.0314975f $X=10.21 $Y=0.34 $X2=0
+ $Y2=0
cc_1167 N_A_1823_524#_c_1614_n N_VGND_c_2444_n 0.0127177f $X=9.68 $Y=0.34 $X2=0
+ $Y2=0
cc_1168 N_A_1823_524#_c_1613_n N_A_1677_74#_M1010_s 0.00168754f $X=10.21 $Y=0.34
+ $X2=0 $Y2=0
cc_1169 N_A_1823_524#_c_1612_n N_A_1677_74#_c_2591_n 0.0232012f $X=9.515
+ $Y=0.515 $X2=0 $Y2=0
cc_1170 N_A_1823_524#_c_1615_n N_A_1677_74#_c_2591_n 0.0133511f $X=10.375
+ $Y=0.515 $X2=0 $Y2=0
cc_1171 N_A_1823_524#_c_1613_n N_A_1677_74#_c_2593_n 0.0126419f $X=10.21 $Y=0.34
+ $X2=0 $Y2=0
cc_1172 N_A_1823_524#_c_1615_n N_A_1677_74#_c_2593_n 0.0218734f $X=10.375
+ $Y=0.515 $X2=0 $Y2=0
cc_1173 N_A_2580_74#_c_1835_n N_VPWR_c_1956_n 0.029359f $X=13.255 $Y=2.265 $X2=0
+ $Y2=0
cc_1174 N_A_2580_74#_c_1838_n N_VPWR_c_1957_n 0.00643415f $X=13.985 $Y=1.765
+ $X2=0 $Y2=0
cc_1175 N_A_2580_74#_c_1830_n N_VPWR_c_1957_n 0.00404999f $X=14.975 $Y=1.395
+ $X2=0 $Y2=0
cc_1176 N_A_2580_74#_c_1835_n N_VPWR_c_1957_n 0.0573751f $X=13.255 $Y=2.265
+ $X2=0 $Y2=0
cc_1177 N_A_2580_74#_c_1836_n N_VPWR_c_1957_n 0.0131456f $X=14.53 $Y=1.485 $X2=0
+ $Y2=0
cc_1178 N_A_2580_74#_c_1838_n N_VPWR_c_1958_n 5.25817e-19 $X=13.985 $Y=1.765
+ $X2=0 $Y2=0
cc_1179 N_A_2580_74#_c_1839_n N_VPWR_c_1958_n 0.0106094f $X=14.435 $Y=1.765
+ $X2=0 $Y2=0
cc_1180 N_A_2580_74#_c_1840_n N_VPWR_c_1958_n 0.0109773f $X=14.885 $Y=1.765
+ $X2=0 $Y2=0
cc_1181 N_A_2580_74#_c_1843_n N_VPWR_c_1958_n 5.26866e-19 $X=15.335 $Y=1.765
+ $X2=0 $Y2=0
cc_1182 N_A_2580_74#_c_1840_n N_VPWR_c_1960_n 5.78844e-19 $X=14.885 $Y=1.765
+ $X2=0 $Y2=0
cc_1183 N_A_2580_74#_c_1843_n N_VPWR_c_1960_n 0.0154543f $X=15.335 $Y=1.765
+ $X2=0 $Y2=0
cc_1184 N_A_2580_74#_c_1835_n N_VPWR_c_1970_n 0.00749631f $X=13.255 $Y=2.265
+ $X2=0 $Y2=0
cc_1185 N_A_2580_74#_c_1838_n N_VPWR_c_1971_n 0.00445602f $X=13.985 $Y=1.765
+ $X2=0 $Y2=0
cc_1186 N_A_2580_74#_c_1839_n N_VPWR_c_1971_n 0.00413917f $X=14.435 $Y=1.765
+ $X2=0 $Y2=0
cc_1187 N_A_2580_74#_c_1840_n N_VPWR_c_1972_n 0.00413917f $X=14.885 $Y=1.765
+ $X2=0 $Y2=0
cc_1188 N_A_2580_74#_c_1843_n N_VPWR_c_1972_n 0.00413917f $X=15.335 $Y=1.765
+ $X2=0 $Y2=0
cc_1189 N_A_2580_74#_c_1838_n N_VPWR_c_1947_n 0.00857585f $X=13.985 $Y=1.765
+ $X2=0 $Y2=0
cc_1190 N_A_2580_74#_c_1839_n N_VPWR_c_1947_n 0.00817726f $X=14.435 $Y=1.765
+ $X2=0 $Y2=0
cc_1191 N_A_2580_74#_c_1840_n N_VPWR_c_1947_n 0.00817726f $X=14.885 $Y=1.765
+ $X2=0 $Y2=0
cc_1192 N_A_2580_74#_c_1843_n N_VPWR_c_1947_n 0.00817726f $X=15.335 $Y=1.765
+ $X2=0 $Y2=0
cc_1193 N_A_2580_74#_c_1835_n N_VPWR_c_1947_n 0.0062048f $X=13.255 $Y=2.265
+ $X2=0 $Y2=0
cc_1194 N_A_2580_74#_M1000_g N_Q_c_2330_n 0.00599748f $X=13.76 $Y=0.74 $X2=0
+ $Y2=0
cc_1195 N_A_2580_74#_M1015_g N_Q_c_2330_n 0.00400087f $X=14.345 $Y=0.74 $X2=0
+ $Y2=0
cc_1196 N_A_2580_74#_c_1838_n N_Q_c_2339_n 0.00839931f $X=13.985 $Y=1.765 $X2=0
+ $Y2=0
cc_1197 N_A_2580_74#_c_1830_n N_Q_c_2339_n 0.00682234f $X=14.975 $Y=1.395 $X2=0
+ $Y2=0
cc_1198 N_A_2580_74#_c_1836_n N_Q_c_2339_n 0.0235455f $X=14.53 $Y=1.485 $X2=0
+ $Y2=0
cc_1199 N_A_2580_74#_c_1838_n N_Q_c_2340_n 0.0088579f $X=13.985 $Y=1.765 $X2=0
+ $Y2=0
cc_1200 N_A_2580_74#_c_1839_n N_Q_c_2340_n 3.88029e-19 $X=14.435 $Y=1.765 $X2=0
+ $Y2=0
cc_1201 N_A_2580_74#_M1015_g N_Q_c_2331_n 0.0151786f $X=14.345 $Y=0.74 $X2=0
+ $Y2=0
cc_1202 N_A_2580_74#_M1023_g N_Q_c_2331_n 0.0143475f $X=14.845 $Y=0.74 $X2=0
+ $Y2=0
cc_1203 N_A_2580_74#_c_1830_n N_Q_c_2331_n 0.00383291f $X=14.975 $Y=1.395 $X2=0
+ $Y2=0
cc_1204 N_A_2580_74#_c_1836_n N_Q_c_2331_n 0.0347268f $X=14.53 $Y=1.485 $X2=0
+ $Y2=0
cc_1205 N_A_2580_74#_M1000_g N_Q_c_2332_n 0.00219788f $X=13.76 $Y=0.74 $X2=0
+ $Y2=0
cc_1206 N_A_2580_74#_c_1830_n N_Q_c_2332_n 0.00649429f $X=14.975 $Y=1.395 $X2=0
+ $Y2=0
cc_1207 N_A_2580_74#_c_1836_n N_Q_c_2332_n 0.0278315f $X=14.53 $Y=1.485 $X2=0
+ $Y2=0
cc_1208 N_A_2580_74#_c_1839_n N_Q_c_2341_n 0.0176407f $X=14.435 $Y=1.765 $X2=0
+ $Y2=0
cc_1209 N_A_2580_74#_c_1840_n N_Q_c_2341_n 0.0192773f $X=14.885 $Y=1.765 $X2=0
+ $Y2=0
cc_1210 N_A_2580_74#_c_1830_n N_Q_c_2341_n 0.00966048f $X=14.975 $Y=1.395 $X2=0
+ $Y2=0
cc_1211 N_A_2580_74#_c_1836_n N_Q_c_2341_n 0.0286254f $X=14.53 $Y=1.485 $X2=0
+ $Y2=0
cc_1212 N_A_2580_74#_M1015_g N_Q_c_2333_n 6.22327e-19 $X=14.345 $Y=0.74 $X2=0
+ $Y2=0
cc_1213 N_A_2580_74#_M1023_g N_Q_c_2333_n 0.00926373f $X=14.845 $Y=0.74 $X2=0
+ $Y2=0
cc_1214 N_A_2580_74#_M1027_g N_Q_c_2333_n 0.00788812f $X=15.275 $Y=0.74 $X2=0
+ $Y2=0
cc_1215 N_A_2580_74#_c_1840_n N_Q_c_2342_n 0.00567416f $X=14.885 $Y=1.765 $X2=0
+ $Y2=0
cc_1216 N_A_2580_74#_c_1843_n N_Q_c_2342_n 0.0029216f $X=15.335 $Y=1.765 $X2=0
+ $Y2=0
cc_1217 N_A_2580_74#_c_1832_n N_Q_c_2334_n 0.0049963f $X=15.335 $Y=1.675 $X2=0
+ $Y2=0
cc_1218 N_A_2580_74#_c_1843_n N_Q_c_2334_n 0.0113109f $X=15.335 $Y=1.765 $X2=0
+ $Y2=0
cc_1219 N_A_2580_74#_M1027_g N_Q_c_2335_n 0.00737919f $X=15.275 $Y=0.74 $X2=0
+ $Y2=0
cc_1220 N_A_2580_74#_c_1833_n N_Q_c_2335_n 0.00847991f $X=15.312 $Y=1.395 $X2=0
+ $Y2=0
cc_1221 N_A_2580_74#_M1015_g N_Q_c_2376_n 8.81603e-19 $X=14.345 $Y=0.74 $X2=0
+ $Y2=0
cc_1222 N_A_2580_74#_M1023_g N_Q_c_2376_n 0.00666364f $X=14.845 $Y=0.74 $X2=0
+ $Y2=0
cc_1223 N_A_2580_74#_c_1829_n N_Q_c_2376_n 0.00742135f $X=15.2 $Y=1.395 $X2=0
+ $Y2=0
cc_1224 N_A_2580_74#_c_1830_n N_Q_c_2376_n 0.00426636f $X=14.975 $Y=1.395 $X2=0
+ $Y2=0
cc_1225 N_A_2580_74#_M1027_g N_Q_c_2376_n 0.0114488f $X=15.275 $Y=0.74 $X2=0
+ $Y2=0
cc_1226 N_A_2580_74#_c_1833_n N_Q_c_2376_n 9.29092e-19 $X=15.312 $Y=1.395 $X2=0
+ $Y2=0
cc_1227 N_A_2580_74#_c_1836_n N_Q_c_2376_n 0.0083343f $X=14.53 $Y=1.485 $X2=0
+ $Y2=0
cc_1228 N_A_2580_74#_c_1840_n N_Q_c_2336_n 0.0014206f $X=14.885 $Y=1.765 $X2=0
+ $Y2=0
cc_1229 N_A_2580_74#_c_1829_n N_Q_c_2336_n 0.00220067f $X=15.2 $Y=1.395 $X2=0
+ $Y2=0
cc_1230 N_A_2580_74#_c_1830_n N_Q_c_2336_n 0.0041705f $X=14.975 $Y=1.395 $X2=0
+ $Y2=0
cc_1231 N_A_2580_74#_c_1843_n N_Q_c_2336_n 0.0054475f $X=15.335 $Y=1.765 $X2=0
+ $Y2=0
cc_1232 N_A_2580_74#_c_1836_n N_Q_c_2336_n 0.00211413f $X=14.53 $Y=1.485 $X2=0
+ $Y2=0
cc_1233 N_A_2580_74#_c_1833_n Q 0.00709893f $X=15.312 $Y=1.395 $X2=0 $Y2=0
cc_1234 N_A_2580_74#_M1000_g N_VGND_c_2422_n 0.013974f $X=13.76 $Y=0.74 $X2=0
+ $Y2=0
cc_1235 N_A_2580_74#_M1015_g N_VGND_c_2422_n 7.39638e-19 $X=14.345 $Y=0.74 $X2=0
+ $Y2=0
cc_1236 N_A_2580_74#_c_1834_n N_VGND_c_2422_n 0.0308484f $X=13.045 $Y=0.515
+ $X2=0 $Y2=0
cc_1237 N_A_2580_74#_c_1836_n N_VGND_c_2422_n 0.0266086f $X=14.53 $Y=1.485 $X2=0
+ $Y2=0
cc_1238 N_A_2580_74#_M1000_g N_VGND_c_2423_n 5.94884e-19 $X=13.76 $Y=0.74 $X2=0
+ $Y2=0
cc_1239 N_A_2580_74#_M1015_g N_VGND_c_2423_n 0.0103873f $X=14.345 $Y=0.74 $X2=0
+ $Y2=0
cc_1240 N_A_2580_74#_M1023_g N_VGND_c_2423_n 0.00417204f $X=14.845 $Y=0.74 $X2=0
+ $Y2=0
cc_1241 N_A_2580_74#_M1027_g N_VGND_c_2425_n 0.0178469f $X=15.275 $Y=0.74 $X2=0
+ $Y2=0
cc_1242 N_A_2580_74#_c_1834_n N_VGND_c_2426_n 0.0145639f $X=13.045 $Y=0.515
+ $X2=0 $Y2=0
cc_1243 N_A_2580_74#_M1000_g N_VGND_c_2434_n 0.00383152f $X=13.76 $Y=0.74 $X2=0
+ $Y2=0
cc_1244 N_A_2580_74#_M1015_g N_VGND_c_2434_n 0.00383152f $X=14.345 $Y=0.74 $X2=0
+ $Y2=0
cc_1245 N_A_2580_74#_M1023_g N_VGND_c_2435_n 0.00434272f $X=14.845 $Y=0.74 $X2=0
+ $Y2=0
cc_1246 N_A_2580_74#_M1027_g N_VGND_c_2435_n 0.00434272f $X=15.275 $Y=0.74 $X2=0
+ $Y2=0
cc_1247 N_A_2580_74#_M1000_g N_VGND_c_2444_n 0.00758887f $X=13.76 $Y=0.74 $X2=0
+ $Y2=0
cc_1248 N_A_2580_74#_M1015_g N_VGND_c_2444_n 0.00758887f $X=14.345 $Y=0.74 $X2=0
+ $Y2=0
cc_1249 N_A_2580_74#_M1023_g N_VGND_c_2444_n 0.00820718f $X=14.845 $Y=0.74 $X2=0
+ $Y2=0
cc_1250 N_A_2580_74#_M1027_g N_VGND_c_2444_n 0.00823934f $X=15.275 $Y=0.74 $X2=0
+ $Y2=0
cc_1251 N_A_2580_74#_c_1834_n N_VGND_c_2444_n 0.0119984f $X=13.045 $Y=0.515
+ $X2=0 $Y2=0
cc_1252 N_VPWR_c_1948_n N_A_288_464#_c_2173_n 0.00764771f $X=0.72 $Y=2.78 $X2=0
+ $Y2=0
cc_1253 N_VPWR_c_1966_n N_A_288_464#_c_2173_n 0.0222791f $X=2.56 $Y=3.33 $X2=0
+ $Y2=0
cc_1254 N_VPWR_c_1947_n N_A_288_464#_c_2173_n 0.0261026f $X=15.6 $Y=3.33 $X2=0
+ $Y2=0
cc_1255 N_VPWR_M1001_d N_A_288_464#_c_2168_n 0.00951605f $X=2.49 $Y=2.32 $X2=0
+ $Y2=0
cc_1256 N_VPWR_c_1949_n N_A_288_464#_c_2168_n 0.0253286f $X=2.725 $Y=2.995 $X2=0
+ $Y2=0
cc_1257 N_VPWR_c_1950_n N_A_288_464#_c_2168_n 0.00194063f $X=3.57 $Y=3.33 $X2=0
+ $Y2=0
cc_1258 N_VPWR_c_1966_n N_A_288_464#_c_2168_n 0.00229351f $X=2.56 $Y=3.33 $X2=0
+ $Y2=0
cc_1259 N_VPWR_c_1947_n N_A_288_464#_c_2168_n 0.00899875f $X=15.6 $Y=3.33 $X2=0
+ $Y2=0
cc_1260 N_VPWR_M1028_d N_A_288_464#_c_2169_n 0.00395001f $X=3.585 $Y=1.84 $X2=0
+ $Y2=0
cc_1261 N_VPWR_c_1951_n N_A_288_464#_c_2169_n 0.0171894f $X=3.735 $Y=2.78 $X2=0
+ $Y2=0
cc_1262 N_VPWR_c_1949_n N_A_288_464#_c_2194_n 0.00578857f $X=2.725 $Y=2.995
+ $X2=0 $Y2=0
cc_1263 N_VPWR_c_1966_n N_A_288_464#_c_2194_n 0.00469602f $X=2.56 $Y=3.33 $X2=0
+ $Y2=0
cc_1264 N_VPWR_c_1947_n N_A_288_464#_c_2194_n 0.00571824f $X=15.6 $Y=3.33 $X2=0
+ $Y2=0
cc_1265 N_VPWR_c_1950_n N_A_288_464#_c_2171_n 0.00302288f $X=3.57 $Y=3.33 $X2=0
+ $Y2=0
cc_1266 N_VPWR_c_1951_n N_A_288_464#_c_2171_n 0.00308348f $X=3.735 $Y=2.78 $X2=0
+ $Y2=0
cc_1267 N_VPWR_c_1947_n N_A_288_464#_c_2171_n 0.00485809f $X=15.6 $Y=3.33 $X2=0
+ $Y2=0
cc_1268 N_VPWR_c_1953_n N_A_1620_373#_c_2289_n 0.0273167f $X=7.8 $Y=2.505 $X2=0
+ $Y2=0
cc_1269 N_VPWR_c_1954_n N_A_1620_373#_c_2289_n 0.00993345f $X=8.7 $Y=2.55 $X2=0
+ $Y2=0
cc_1270 N_VPWR_c_1963_n N_A_1620_373#_c_2289_n 0.00577068f $X=8.535 $Y=3.33
+ $X2=0 $Y2=0
cc_1271 N_VPWR_c_1947_n N_A_1620_373#_c_2289_n 0.00739579f $X=15.6 $Y=3.33 $X2=0
+ $Y2=0
cc_1272 N_VPWR_M1047_s N_A_1620_373#_c_2290_n 0.00512955f $X=8.55 $Y=1.865 $X2=0
+ $Y2=0
cc_1273 N_VPWR_c_1954_n N_A_1620_373#_c_2290_n 0.0220323f $X=8.7 $Y=2.55 $X2=0
+ $Y2=0
cc_1274 N_VPWR_c_1955_n A_2103_508# 0.0126284f $X=11.29 $Y=2.815 $X2=-0.19
+ $Y2=-0.245
cc_1275 N_VPWR_c_1968_n A_2103_508# 0.0173016f $X=11.125 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_1276 N_VPWR_c_1947_n A_2103_508# 0.0147808f $X=15.6 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_1277 N_VPWR_c_1957_n N_Q_c_2340_n 0.03041f $X=13.705 $Y=2.265 $X2=0 $Y2=0
cc_1278 N_VPWR_c_1958_n N_Q_c_2340_n 0.0255358f $X=14.66 $Y=2.405 $X2=0 $Y2=0
cc_1279 N_VPWR_c_1971_n N_Q_c_2340_n 0.0123628f $X=14.495 $Y=3.33 $X2=0 $Y2=0
cc_1280 N_VPWR_c_1947_n N_Q_c_2340_n 0.0101999f $X=15.6 $Y=3.33 $X2=0 $Y2=0
cc_1281 N_VPWR_M1037_s N_Q_c_2341_n 0.00201799f $X=14.51 $Y=1.84 $X2=0 $Y2=0
cc_1282 N_VPWR_c_1958_n N_Q_c_2341_n 0.0179913f $X=14.66 $Y=2.405 $X2=0 $Y2=0
cc_1283 N_VPWR_c_1958_n N_Q_c_2342_n 0.0430177f $X=14.66 $Y=2.405 $X2=0 $Y2=0
cc_1284 N_VPWR_c_1960_n N_Q_c_2342_n 0.0540587f $X=15.56 $Y=2.115 $X2=0 $Y2=0
cc_1285 N_VPWR_c_1972_n N_Q_c_2342_n 0.00749631f $X=15.395 $Y=3.33 $X2=0 $Y2=0
cc_1286 N_VPWR_c_1947_n N_Q_c_2342_n 0.0062048f $X=15.6 $Y=3.33 $X2=0 $Y2=0
cc_1287 N_VPWR_c_1960_n N_Q_c_2334_n 0.00462998f $X=15.56 $Y=2.115 $X2=0 $Y2=0
cc_1288 N_VPWR_c_1960_n N_Q_c_2336_n 0.0145667f $X=15.56 $Y=2.115 $X2=0 $Y2=0
cc_1289 N_VPWR_c_1960_n N_Q_c_2338_n 0.0207054f $X=15.56 $Y=2.115 $X2=0 $Y2=0
cc_1290 N_A_288_464#_c_2173_n A_414_464# 0.00525631f $X=2.215 $Y=2.785 $X2=-0.19
+ $Y2=-0.245
cc_1291 N_A_288_464#_c_2164_n A_414_464# 0.00140003f $X=2.3 $Y=2.49 $X2=-0.19
+ $Y2=-0.245
cc_1292 N_A_288_464#_c_2194_n A_414_464# 0.00344777f $X=2.3 $Y=2.575 $X2=-0.19
+ $Y2=-0.245
cc_1293 N_A_288_464#_c_2182_n N_VGND_c_2415_n 0.010729f $X=1.875 $Y=0.575 $X2=0
+ $Y2=0
cc_1294 N_A_288_464#_c_2182_n N_VGND_c_2429_n 0.0142996f $X=1.875 $Y=0.575 $X2=0
+ $Y2=0
cc_1295 N_A_288_464#_c_2182_n N_VGND_c_2444_n 0.0165485f $X=1.875 $Y=0.575 $X2=0
+ $Y2=0
cc_1296 N_Q_c_2331_n N_VGND_M1015_s 0.00250873f $X=14.895 $Y=1.065 $X2=0 $Y2=0
cc_1297 N_Q_c_2330_n N_VGND_c_2422_n 0.0458088f $X=14.06 $Y=0.515 $X2=0 $Y2=0
cc_1298 N_Q_c_2332_n N_VGND_c_2422_n 0.0116373f $X=14.225 $Y=1.065 $X2=0 $Y2=0
cc_1299 N_Q_c_2330_n N_VGND_c_2423_n 0.0180508f $X=14.06 $Y=0.515 $X2=0 $Y2=0
cc_1300 N_Q_c_2331_n N_VGND_c_2423_n 0.0209867f $X=14.895 $Y=1.065 $X2=0 $Y2=0
cc_1301 N_Q_c_2333_n N_VGND_c_2423_n 0.0180508f $X=15.06 $Y=0.515 $X2=0 $Y2=0
cc_1302 N_Q_c_2333_n N_VGND_c_2425_n 0.0288948f $X=15.06 $Y=0.515 $X2=0 $Y2=0
cc_1303 N_Q_c_2335_n N_VGND_c_2425_n 0.0277188f $X=15.485 $Y=1.355 $X2=0 $Y2=0
cc_1304 N_Q_c_2330_n N_VGND_c_2434_n 0.0146357f $X=14.06 $Y=0.515 $X2=0 $Y2=0
cc_1305 N_Q_c_2333_n N_VGND_c_2435_n 0.0144922f $X=15.06 $Y=0.515 $X2=0 $Y2=0
cc_1306 N_Q_c_2330_n N_VGND_c_2444_n 0.0121141f $X=14.06 $Y=0.515 $X2=0 $Y2=0
cc_1307 N_Q_c_2333_n N_VGND_c_2444_n 0.0118826f $X=15.06 $Y=0.515 $X2=0 $Y2=0
cc_1308 N_VGND_c_2419_n N_A_1677_74#_c_2590_n 0.0238508f $X=8.095 $Y=0.495 $X2=0
+ $Y2=0
cc_1309 N_VGND_c_2420_n N_A_1677_74#_c_2590_n 0.0218329f $X=8.955 $Y=0.515 $X2=0
+ $Y2=0
cc_1310 N_VGND_c_2432_n N_A_1677_74#_c_2590_n 0.00749631f $X=8.79 $Y=0 $X2=0
+ $Y2=0
cc_1311 N_VGND_c_2444_n N_A_1677_74#_c_2590_n 0.0062048f $X=15.6 $Y=0 $X2=0
+ $Y2=0
cc_1312 N_VGND_c_2420_n N_A_1677_74#_c_2591_n 0.0243991f $X=8.955 $Y=0.515 $X2=0
+ $Y2=0
