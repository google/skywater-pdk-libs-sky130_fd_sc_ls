* File: sky130_fd_sc_ls__sdfrtp_4.pxi.spice
* Created: Fri Aug 28 14:03:32 2020
* 
x_PM_SKY130_FD_SC_LS__SDFRTP_4%A_27_74# N_A_27_74#_M1036_s N_A_27_74#_M1023_s
+ N_A_27_74#_c_302_n N_A_27_74#_c_303_n N_A_27_74#_M1005_g N_A_27_74#_c_309_n
+ N_A_27_74#_M1014_g N_A_27_74#_c_304_n N_A_27_74#_c_305_n N_A_27_74#_c_311_n
+ N_A_27_74#_c_306_n N_A_27_74#_c_312_n N_A_27_74#_c_307_n N_A_27_74#_c_313_n
+ N_A_27_74#_c_314_n N_A_27_74#_c_308_n PM_SKY130_FD_SC_LS__SDFRTP_4%A_27_74#
x_PM_SKY130_FD_SC_LS__SDFRTP_4%SCE N_SCE_c_393_n N_SCE_M1036_g N_SCE_c_394_n
+ N_SCE_M1023_g N_SCE_c_395_n N_SCE_c_396_n N_SCE_M1026_g N_SCE_c_385_n
+ N_SCE_M1037_g N_SCE_c_387_n N_SCE_c_388_n N_SCE_c_389_n N_SCE_c_390_n SCE SCE
+ SCE N_SCE_c_391_n SCE N_SCE_c_392_n PM_SKY130_FD_SC_LS__SDFRTP_4%SCE
x_PM_SKY130_FD_SC_LS__SDFRTP_4%D N_D_M1006_g N_D_c_471_n N_D_c_476_n N_D_M1002_g
+ D N_D_c_472_n N_D_c_473_n N_D_c_474_n PM_SKY130_FD_SC_LS__SDFRTP_4%D
x_PM_SKY130_FD_SC_LS__SDFRTP_4%SCD N_SCD_c_521_n N_SCD_M1029_g N_SCD_M1040_g
+ N_SCD_c_518_n SCD SCD N_SCD_c_520_n PM_SKY130_FD_SC_LS__SDFRTP_4%SCD
x_PM_SKY130_FD_SC_LS__SDFRTP_4%CLK N_CLK_c_560_n N_CLK_M1010_g N_CLK_M1030_g CLK
+ PM_SKY130_FD_SC_LS__SDFRTP_4%CLK
x_PM_SKY130_FD_SC_LS__SDFRTP_4%A_1034_392# N_A_1034_392#_M1013_d
+ N_A_1034_392#_M1034_d N_A_1034_392#_c_635_n N_A_1034_392#_c_636_n
+ N_A_1034_392#_M1000_g N_A_1034_392#_c_614_n N_A_1034_392#_M1041_g
+ N_A_1034_392#_c_616_n N_A_1034_392#_M1003_g N_A_1034_392#_c_617_n
+ N_A_1034_392#_c_618_n N_A_1034_392#_c_638_n N_A_1034_392#_M1018_g
+ N_A_1034_392#_c_619_n N_A_1034_392#_c_620_n N_A_1034_392#_c_621_n
+ N_A_1034_392#_c_622_n N_A_1034_392#_c_623_n N_A_1034_392#_c_624_n
+ N_A_1034_392#_c_625_n N_A_1034_392#_c_678_p N_A_1034_392#_c_626_n
+ N_A_1034_392#_c_627_n N_A_1034_392#_c_628_n N_A_1034_392#_c_629_n
+ N_A_1034_392#_c_665_p N_A_1034_392#_c_642_n N_A_1034_392#_c_630_n
+ N_A_1034_392#_c_631_n N_A_1034_392#_c_632_n N_A_1034_392#_c_633_n
+ N_A_1034_392#_c_634_n PM_SKY130_FD_SC_LS__SDFRTP_4%A_1034_392#
x_PM_SKY130_FD_SC_LS__SDFRTP_4%A_1367_112# N_A_1367_112#_M1019_d
+ N_A_1367_112#_M1031_d N_A_1367_112#_M1044_g N_A_1367_112#_c_848_n
+ N_A_1367_112#_c_849_n N_A_1367_112#_M1009_g N_A_1367_112#_c_844_n
+ N_A_1367_112#_c_845_n N_A_1367_112#_c_863_n N_A_1367_112#_c_846_n
+ N_A_1367_112#_c_847_n N_A_1367_112#_c_853_n N_A_1367_112#_c_874_n
+ N_A_1367_112#_c_876_n PM_SKY130_FD_SC_LS__SDFRTP_4%A_1367_112#
x_PM_SKY130_FD_SC_LS__SDFRTP_4%RESET_B N_RESET_B_c_953_n N_RESET_B_M1012_g
+ N_RESET_B_c_964_n N_RESET_B_M1045_g N_RESET_B_c_955_n N_RESET_B_c_956_n
+ N_RESET_B_M1024_g N_RESET_B_c_958_n N_RESET_B_c_959_n N_RESET_B_c_965_n
+ N_RESET_B_M1001_g N_RESET_B_c_960_n N_RESET_B_M1038_g N_RESET_B_c_968_n
+ N_RESET_B_c_969_n N_RESET_B_M1015_g N_RESET_B_c_962_n N_RESET_B_c_970_n
+ N_RESET_B_c_971_n N_RESET_B_c_972_n N_RESET_B_c_973_n N_RESET_B_c_974_n
+ RESET_B N_RESET_B_c_976_n N_RESET_B_c_977_n N_RESET_B_c_978_n
+ N_RESET_B_c_979_n N_RESET_B_c_980_n PM_SKY130_FD_SC_LS__SDFRTP_4%RESET_B
x_PM_SKY130_FD_SC_LS__SDFRTP_4%A_1236_138# N_A_1236_138#_M1032_d
+ N_A_1236_138#_M1000_d N_A_1236_138#_M1001_d N_A_1236_138#_M1019_g
+ N_A_1236_138#_c_1180_n N_A_1236_138#_c_1188_n N_A_1236_138#_M1031_g
+ N_A_1236_138#_c_1189_n N_A_1236_138#_c_1202_n N_A_1236_138#_c_1181_n
+ N_A_1236_138#_c_1225_n N_A_1236_138#_c_1182_n N_A_1236_138#_c_1183_n
+ N_A_1236_138#_c_1184_n N_A_1236_138#_c_1185_n N_A_1236_138#_c_1186_n
+ N_A_1236_138#_c_1193_n PM_SKY130_FD_SC_LS__SDFRTP_4%A_1236_138#
x_PM_SKY130_FD_SC_LS__SDFRTP_4%A_837_98# N_A_837_98#_M1010_s N_A_837_98#_M1030_s
+ N_A_837_98#_M1034_g N_A_837_98#_M1013_g N_A_837_98#_c_1314_n
+ N_A_837_98#_c_1315_n N_A_837_98#_c_1316_n N_A_837_98#_c_1329_n
+ N_A_837_98#_c_1330_n N_A_837_98#_c_1317_n N_A_837_98#_c_1318_n
+ N_A_837_98#_M1032_g N_A_837_98#_c_1331_n N_A_837_98#_c_1332_n
+ N_A_837_98#_c_1333_n N_A_837_98#_M1008_g N_A_837_98#_c_1334_n
+ N_A_837_98#_c_1335_n N_A_837_98#_c_1336_n N_A_837_98#_M1042_g
+ N_A_837_98#_c_1319_n N_A_837_98#_c_1320_n N_A_837_98#_M1027_g
+ N_A_837_98#_c_1340_n N_A_837_98#_c_1347_n N_A_837_98#_c_1341_n
+ N_A_837_98#_c_1351_n N_A_837_98#_c_1353_n N_A_837_98#_c_1322_n
+ N_A_837_98#_c_1323_n N_A_837_98#_c_1342_n N_A_837_98#_c_1324_n
+ N_A_837_98#_c_1325_n N_A_837_98#_c_1326_n
+ PM_SKY130_FD_SC_LS__SDFRTP_4%A_837_98#
x_PM_SKY130_FD_SC_LS__SDFRTP_4%A_2003_48# N_A_2003_48#_M1020_d
+ N_A_2003_48#_M1015_d N_A_2003_48#_M1021_g N_A_2003_48#_c_1520_n
+ N_A_2003_48#_c_1529_n N_A_2003_48#_M1043_g N_A_2003_48#_c_1521_n
+ N_A_2003_48#_c_1522_n N_A_2003_48#_c_1523_n N_A_2003_48#_c_1524_n
+ N_A_2003_48#_c_1525_n N_A_2003_48#_c_1530_n N_A_2003_48#_c_1526_n
+ N_A_2003_48#_c_1527_n PM_SKY130_FD_SC_LS__SDFRTP_4%A_2003_48#
x_PM_SKY130_FD_SC_LS__SDFRTP_4%A_1745_74# N_A_1745_74#_M1003_d
+ N_A_1745_74#_M1042_d N_A_1745_74#_c_1608_n N_A_1745_74#_M1020_g
+ N_A_1745_74#_c_1609_n N_A_1745_74#_c_1624_n N_A_1745_74#_c_1625_n
+ N_A_1745_74#_M1035_g N_A_1745_74#_c_1610_n N_A_1745_74#_c_1626_n
+ N_A_1745_74#_M1033_g N_A_1745_74#_c_1611_n N_A_1745_74#_M1011_g
+ N_A_1745_74#_c_1612_n N_A_1745_74#_c_1613_n N_A_1745_74#_c_1628_n
+ N_A_1745_74#_M1046_g N_A_1745_74#_c_1614_n N_A_1745_74#_c_1615_n
+ N_A_1745_74#_c_1616_n N_A_1745_74#_c_1641_n N_A_1745_74#_c_1630_n
+ N_A_1745_74#_c_1617_n N_A_1745_74#_c_1618_n N_A_1745_74#_c_1619_n
+ N_A_1745_74#_c_1632_n N_A_1745_74#_c_1633_n N_A_1745_74#_c_1634_n
+ N_A_1745_74#_c_1620_n N_A_1745_74#_c_1621_n N_A_1745_74#_c_1622_n
+ PM_SKY130_FD_SC_LS__SDFRTP_4%A_1745_74#
x_PM_SKY130_FD_SC_LS__SDFRTP_4%A_2339_74# N_A_2339_74#_M1011_s
+ N_A_2339_74#_M1033_d N_A_2339_74#_c_1772_n N_A_2339_74#_M1007_g
+ N_A_2339_74#_c_1773_n N_A_2339_74#_c_1774_n N_A_2339_74#_c_1775_n
+ N_A_2339_74#_M1016_g N_A_2339_74#_c_1783_n N_A_2339_74#_M1004_g
+ N_A_2339_74#_c_1784_n N_A_2339_74#_M1017_g N_A_2339_74#_c_1785_n
+ N_A_2339_74#_M1025_g N_A_2339_74#_c_1776_n N_A_2339_74#_M1022_g
+ N_A_2339_74#_c_1786_n N_A_2339_74#_M1039_g N_A_2339_74#_c_1777_n
+ N_A_2339_74#_M1028_g N_A_2339_74#_c_1778_n N_A_2339_74#_c_1779_n
+ N_A_2339_74#_c_1780_n N_A_2339_74#_c_1781_n N_A_2339_74#_c_1782_n
+ PM_SKY130_FD_SC_LS__SDFRTP_4%A_2339_74#
x_PM_SKY130_FD_SC_LS__SDFRTP_4%VPWR N_VPWR_M1023_d N_VPWR_M1029_d N_VPWR_M1030_d
+ N_VPWR_M1009_d N_VPWR_M1031_s N_VPWR_M1043_d N_VPWR_M1035_d N_VPWR_M1046_s
+ N_VPWR_M1017_d N_VPWR_M1039_d N_VPWR_c_1890_n N_VPWR_c_1891_n N_VPWR_c_1892_n
+ N_VPWR_c_1893_n N_VPWR_c_1894_n N_VPWR_c_1895_n N_VPWR_c_1896_n
+ N_VPWR_c_1897_n N_VPWR_c_1898_n N_VPWR_c_1899_n N_VPWR_c_1900_n
+ N_VPWR_c_1901_n N_VPWR_c_1902_n N_VPWR_c_1903_n N_VPWR_c_1904_n
+ N_VPWR_c_1905_n VPWR N_VPWR_c_1906_n N_VPWR_c_1907_n N_VPWR_c_1908_n
+ N_VPWR_c_1909_n N_VPWR_c_1910_n N_VPWR_c_1911_n N_VPWR_c_1912_n
+ N_VPWR_c_1913_n N_VPWR_c_1914_n N_VPWR_c_1915_n N_VPWR_c_1916_n
+ N_VPWR_c_1917_n N_VPWR_c_1918_n N_VPWR_c_1889_n
+ PM_SKY130_FD_SC_LS__SDFRTP_4%VPWR
x_PM_SKY130_FD_SC_LS__SDFRTP_4%A_415_81# N_A_415_81#_M1006_d N_A_415_81#_M1032_s
+ N_A_415_81#_M1002_d N_A_415_81#_M1045_d N_A_415_81#_M1000_s
+ N_A_415_81#_c_2083_n N_A_415_81#_c_2099_n N_A_415_81#_c_2084_n
+ N_A_415_81#_c_2085_n N_A_415_81#_c_2091_n N_A_415_81#_c_2086_n
+ N_A_415_81#_c_2092_n N_A_415_81#_c_2087_n N_A_415_81#_c_2088_n
+ N_A_415_81#_c_2093_n N_A_415_81#_c_2094_n N_A_415_81#_c_2089_n
+ N_A_415_81#_c_2096_n N_A_415_81#_c_2097_n N_A_415_81#_c_2098_n
+ N_A_415_81#_c_2135_n PM_SKY130_FD_SC_LS__SDFRTP_4%A_415_81#
x_PM_SKY130_FD_SC_LS__SDFRTP_4%Q N_Q_M1007_s N_Q_M1022_s N_Q_M1004_s N_Q_M1025_s
+ N_Q_c_2245_n N_Q_c_2256_n N_Q_c_2260_n N_Q_c_2249_n N_Q_c_2250_n N_Q_c_2251_n
+ N_Q_c_2252_n N_Q_c_2246_n N_Q_c_2247_n Q PM_SKY130_FD_SC_LS__SDFRTP_4%Q
x_PM_SKY130_FD_SC_LS__SDFRTP_4%VGND N_VGND_M1036_d N_VGND_M1012_d N_VGND_M1010_d
+ N_VGND_M1024_d N_VGND_M1021_d N_VGND_M1011_d N_VGND_M1016_d N_VGND_M1028_d
+ N_VGND_c_2312_n N_VGND_c_2313_n N_VGND_c_2314_n N_VGND_c_2315_n
+ N_VGND_c_2316_n N_VGND_c_2317_n N_VGND_c_2318_n N_VGND_c_2319_n
+ N_VGND_c_2320_n N_VGND_c_2321_n VGND N_VGND_c_2322_n N_VGND_c_2323_n
+ N_VGND_c_2324_n N_VGND_c_2325_n N_VGND_c_2326_n N_VGND_c_2327_n
+ N_VGND_c_2328_n N_VGND_c_2329_n N_VGND_c_2330_n N_VGND_c_2331_n
+ N_VGND_c_2332_n N_VGND_c_2333_n N_VGND_c_2334_n
+ PM_SKY130_FD_SC_LS__SDFRTP_4%VGND
x_PM_SKY130_FD_SC_LS__SDFRTP_4%noxref_24 N_noxref_24_M1005_s N_noxref_24_M1040_d
+ N_noxref_24_c_2457_n N_noxref_24_c_2475_n N_noxref_24_c_2458_n
+ PM_SKY130_FD_SC_LS__SDFRTP_4%noxref_24
cc_1 VNB N_A_27_74#_c_302_n 0.0258189f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=1.01
cc_2 VNB N_A_27_74#_c_303_n 0.0213547f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.935
cc_3 VNB N_A_27_74#_c_304_n 0.0257773f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=0.58
cc_4 VNB N_A_27_74#_c_305_n 0.0190417f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=2.005
cc_5 VNB N_A_27_74#_c_306_n 0.00987534f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.1
cc_6 VNB N_A_27_74#_c_307_n 0.018224f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.1
cc_7 VNB N_A_27_74#_c_308_n 0.0395906f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.01
cc_8 VNB N_SCE_M1036_g 0.0668709f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_SCE_c_385_n 0.0558046f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.935
cc_10 VNB N_SCE_M1037_g 0.0220088f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=0.58
cc_11 VNB N_SCE_c_387_n 0.00775502f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=2.005
cc_12 VNB N_SCE_c_388_n 0.0420954f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.175
cc_13 VNB N_SCE_c_389_n 0.0130109f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.465
cc_14 VNB N_SCE_c_390_n 0.00601274f $X=-0.19 $Y=-0.245 $X2=0.365 $Y2=1.1
cc_15 VNB N_SCE_c_391_n 0.0106235f $X=-0.19 $Y=-0.245 $X2=2.535 $Y2=1.995
cc_16 VNB N_SCE_c_392_n 0.00168276f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_D_c_471_n 0.027915f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_D_c_472_n 0.0381078f $X=-0.19 $Y=-0.245 $X2=2.495 $Y2=2.245
cc_19 VNB N_D_c_473_n 0.00727955f $X=-0.19 $Y=-0.245 $X2=2.495 $Y2=2.64
cc_20 VNB N_D_c_474_n 0.0173744f $X=-0.19 $Y=-0.245 $X2=2.495 $Y2=2.64
cc_21 VNB N_SCD_M1040_g 0.0396526f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_SCD_c_518_n 0.00374897f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.615
cc_23 VNB SCD 0.00354477f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.615
cc_24 VNB N_SCD_c_520_n 0.0154615f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.58
cc_25 VNB N_CLK_c_560_n 0.095406f $X=-0.19 $Y=-0.245 $X2=0.135 $Y2=0.37
cc_26 VNB CLK 0.0139448f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.615
cc_27 VNB N_A_1034_392#_c_614_n 0.00991128f $X=-0.19 $Y=-0.245 $X2=2.495
+ $Y2=2.245
cc_28 VNB N_A_1034_392#_M1041_g 0.0361107f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.58
cc_29 VNB N_A_1034_392#_c_616_n 0.0168538f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_1034_392#_c_617_n 0.0237434f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.175
cc_31 VNB N_A_1034_392#_c_618_n 0.00657402f $X=-0.19 $Y=-0.245 $X2=0.28
+ $Y2=2.465
cc_32 VNB N_A_1034_392#_c_619_n 0.00764076f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_1034_392#_c_620_n 8.1098e-19 $X=-0.19 $Y=-0.245 $X2=0.445 $Y2=2.09
cc_34 VNB N_A_1034_392#_c_621_n 0.0325626f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.1
cc_35 VNB N_A_1034_392#_c_622_n 0.00467722f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.09
cc_36 VNB N_A_1034_392#_c_623_n 0.00130626f $X=-0.19 $Y=-0.245 $X2=2.54
+ $Y2=1.995
cc_37 VNB N_A_1034_392#_c_624_n 0.00176975f $X=-0.19 $Y=-0.245 $X2=2.535
+ $Y2=1.995
cc_38 VNB N_A_1034_392#_c_625_n 0.00102705f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_1034_392#_c_626_n 0.00657839f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_1034_392#_c_627_n 0.00209509f $X=-0.19 $Y=-0.245 $X2=2.535
+ $Y2=1.995
cc_41 VNB N_A_1034_392#_c_628_n 0.00144678f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_1034_392#_c_629_n 0.005194f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_1034_392#_c_630_n 0.00223099f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_1034_392#_c_631_n 0.00756725f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_1034_392#_c_632_n 0.0332641f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_1034_392#_c_633_n 0.00593212f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_1034_392#_c_634_n 0.00982041f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_1367_112#_M1044_g 0.0347927f $X=-0.19 $Y=-0.245 $X2=1.485
+ $Y2=0.935
cc_49 VNB N_A_1367_112#_c_844_n 0.00473079f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_1367_112#_c_845_n 0.0144435f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=1.265
cc_51 VNB N_A_1367_112#_c_846_n 0.00556937f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_1367_112#_c_847_n 0.00450848f $X=-0.19 $Y=-0.245 $X2=0.365 $Y2=1.1
cc_53 VNB N_RESET_B_c_953_n 0.0312683f $X=-0.19 $Y=-0.245 $X2=0.135 $Y2=2.32
cc_54 VNB N_RESET_B_M1012_g 0.0189594f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_RESET_B_c_955_n 0.267881f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.615
cc_56 VNB N_RESET_B_c_956_n 0.012806f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.615
cc_57 VNB N_RESET_B_M1024_g 0.0336923f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.935
cc_58 VNB N_RESET_B_c_958_n 0.0238599f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.58
cc_59 VNB N_RESET_B_c_959_n 0.00691999f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=0.58
cc_60 VNB N_RESET_B_c_960_n 0.0181108f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.465
cc_61 VNB N_RESET_B_M1038_g 0.0569134f $X=-0.19 $Y=-0.245 $X2=0.365 $Y2=1.1
cc_62 VNB N_RESET_B_c_962_n 0.00908099f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.09
cc_63 VNB N_A_1236_138#_M1019_g 0.0225417f $X=-0.19 $Y=-0.245 $X2=2.495
+ $Y2=2.245
cc_64 VNB N_A_1236_138#_c_1180_n 0.0164115f $X=-0.19 $Y=-0.245 $X2=2.495
+ $Y2=2.64
cc_65 VNB N_A_1236_138#_c_1181_n 0.00367242f $X=-0.19 $Y=-0.245 $X2=0.975
+ $Y2=1.1
cc_66 VNB N_A_1236_138#_c_1182_n 5.47792e-19 $X=-0.19 $Y=-0.245 $X2=2.375
+ $Y2=2.09
cc_67 VNB N_A_1236_138#_c_1183_n 0.00176601f $X=-0.19 $Y=-0.245 $X2=0.445
+ $Y2=2.09
cc_68 VNB N_A_1236_138#_c_1184_n 0.00526285f $X=-0.19 $Y=-0.245 $X2=0.28
+ $Y2=2.09
cc_69 VNB N_A_1236_138#_c_1185_n 0.0281158f $X=-0.19 $Y=-0.245 $X2=2.54
+ $Y2=1.995
cc_70 VNB N_A_1236_138#_c_1186_n 0.00176618f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_837_98#_c_1314_n 0.0127498f $X=-0.19 $Y=-0.245 $X2=2.495 $Y2=2.64
cc_72 VNB N_A_837_98#_c_1315_n 0.0234148f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.58
cc_73 VNB N_A_837_98#_c_1316_n 0.00893594f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=0.58
cc_74 VNB N_A_837_98#_c_1317_n 0.0269744f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=2.005
cc_75 VNB N_A_837_98#_c_1318_n 0.0150195f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.465
cc_76 VNB N_A_837_98#_c_1319_n 0.019724f $X=-0.19 $Y=-0.245 $X2=2.54 $Y2=2.09
cc_77 VNB N_A_837_98#_c_1320_n 0.00441832f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_837_98#_M1027_g 0.0510568f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.1
cc_79 VNB N_A_837_98#_c_1322_n 0.00106022f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_837_98#_c_1323_n 0.00252759f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_837_98#_c_1324_n 0.00710906f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_837_98#_c_1325_n 0.0250817f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_837_98#_c_1326_n 0.0154349f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_2003_48#_M1021_g 0.0340019f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.935
cc_85 VNB N_A_2003_48#_c_1520_n 0.0060931f $X=-0.19 $Y=-0.245 $X2=2.495
+ $Y2=2.245
cc_86 VNB N_A_2003_48#_c_1521_n 0.0178026f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.58
cc_87 VNB N_A_2003_48#_c_1522_n 0.00567377f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_2003_48#_c_1523_n 0.00480935f $X=-0.19 $Y=-0.245 $X2=0.365 $Y2=1.1
cc_89 VNB N_A_2003_48#_c_1524_n 0.00289977f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.1
cc_90 VNB N_A_2003_48#_c_1525_n 0.031198f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.1
cc_91 VNB N_A_2003_48#_c_1526_n 0.00270148f $X=-0.19 $Y=-0.245 $X2=2.54
+ $Y2=1.995
cc_92 VNB N_A_2003_48#_c_1527_n 0.00662489f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_1745_74#_c_1608_n 0.021255f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=1.01
cc_94 VNB N_A_1745_74#_c_1609_n 0.00668157f $X=-0.19 $Y=-0.245 $X2=2.495
+ $Y2=2.245
cc_95 VNB N_A_1745_74#_c_1610_n 0.0250522f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=0.58
cc_96 VNB N_A_1745_74#_c_1611_n 0.0185474f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.465
cc_97 VNB N_A_1745_74#_c_1612_n 0.0159493f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.1
cc_98 VNB N_A_1745_74#_c_1613_n 0.014028f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.1
cc_99 VNB N_A_1745_74#_c_1614_n 0.0143997f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.1
cc_100 VNB N_A_1745_74#_c_1615_n 0.00251602f $X=-0.19 $Y=-0.245 $X2=0.28
+ $Y2=2.09
cc_101 VNB N_A_1745_74#_c_1616_n 0.00496366f $X=-0.19 $Y=-0.245 $X2=2.54
+ $Y2=1.995
cc_102 VNB N_A_1745_74#_c_1617_n 0.00146437f $X=-0.19 $Y=-0.245 $X2=2.535
+ $Y2=1.995
cc_103 VNB N_A_1745_74#_c_1618_n 0.00359384f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_A_1745_74#_c_1619_n 0.0291774f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_A_1745_74#_c_1620_n 0.00123798f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_A_1745_74#_c_1621_n 0.00179963f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_A_1745_74#_c_1622_n 0.0646681f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_A_2339_74#_c_1772_n 0.0177259f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=1.01
cc_109 VNB N_A_2339_74#_c_1773_n 0.0142247f $X=-0.19 $Y=-0.245 $X2=1.485
+ $Y2=0.615
cc_110 VNB N_A_2339_74#_c_1774_n 0.00638412f $X=-0.19 $Y=-0.245 $X2=1.485
+ $Y2=0.615
cc_111 VNB N_A_2339_74#_c_1775_n 0.021315f $X=-0.19 $Y=-0.245 $X2=2.495
+ $Y2=2.245
cc_112 VNB N_A_2339_74#_c_1776_n 0.0221017f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_A_2339_74#_c_1777_n 0.0216728f $X=-0.19 $Y=-0.245 $X2=2.375
+ $Y2=2.09
cc_114 VNB N_A_2339_74#_c_1778_n 0.00311192f $X=-0.19 $Y=-0.245 $X2=2.535
+ $Y2=1.995
cc_115 VNB N_A_2339_74#_c_1779_n 0.00104691f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_A_2339_74#_c_1780_n 0.00999107f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_A_2339_74#_c_1781_n 0.00570341f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_A_2339_74#_c_1782_n 0.14135f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_VPWR_c_1889_n 0.621437f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_A_415_81#_c_2083_n 0.00667808f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_A_415_81#_c_2084_n 0.0157401f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_A_415_81#_c_2085_n 0.00481408f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.1
cc_123 VNB N_A_415_81#_c_2086_n 0.0028959f $X=-0.19 $Y=-0.245 $X2=2.535
+ $Y2=1.995
cc_124 VNB N_A_415_81#_c_2087_n 0.00513426f $X=-0.19 $Y=-0.245 $X2=0.975
+ $Y2=1.01
cc_125 VNB N_A_415_81#_c_2088_n 0.00196739f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_A_415_81#_c_2089_n 0.00250836f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_Q_c_2245_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.935
cc_128 VNB N_Q_c_2246_n 0.00178889f $X=-0.19 $Y=-0.245 $X2=2.535 $Y2=1.995
cc_129 VNB N_Q_c_2247_n 0.00200996f $X=-0.19 $Y=-0.245 $X2=2.54 $Y2=2.09
cc_130 VNB Q 0.0195094f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.01
cc_131 VNB N_VGND_c_2312_n 0.0110567f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.1
cc_132 VNB N_VGND_c_2313_n 0.0136116f $X=-0.19 $Y=-0.245 $X2=0.445 $Y2=2.09
cc_133 VNB N_VGND_c_2314_n 0.0151298f $X=-0.19 $Y=-0.245 $X2=2.535 $Y2=1.995
cc_134 VNB N_VGND_c_2315_n 0.0574849f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_VGND_c_2316_n 0.00428891f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_VGND_c_2317_n 0.00497485f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_VGND_c_2318_n 0.0120272f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB N_VGND_c_2319_n 0.0413125f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VNB N_VGND_c_2320_n 0.0653362f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_VGND_c_2321_n 0.00432799f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_141 VNB N_VGND_c_2322_n 0.0173909f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_142 VNB N_VGND_c_2323_n 0.0187711f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_143 VNB N_VGND_c_2324_n 0.0602754f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_144 VNB N_VGND_c_2325_n 0.0428668f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_145 VNB N_VGND_c_2326_n 0.0151727f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_146 VNB N_VGND_c_2327_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_147 VNB N_VGND_c_2328_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_148 VNB N_VGND_c_2329_n 0.0142666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_149 VNB N_VGND_c_2330_n 0.00808418f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_150 VNB N_VGND_c_2331_n 0.00481148f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_151 VNB N_VGND_c_2332_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_152 VNB N_VGND_c_2333_n 0.0272142f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_153 VNB N_VGND_c_2334_n 0.765689f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_154 VNB N_noxref_24_c_2457_n 0.0168149f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=1.01
cc_155 VNB N_noxref_24_c_2458_n 0.00655627f $X=-0.19 $Y=-0.245 $X2=2.495
+ $Y2=2.64
cc_156 VPB N_A_27_74#_c_309_n 0.051379f $X=-0.19 $Y=1.66 $X2=2.495 $Y2=2.245
cc_157 VPB N_A_27_74#_c_305_n 0.016494f $X=-0.19 $Y=1.66 $X2=0.2 $Y2=2.005
cc_158 VPB N_A_27_74#_c_311_n 0.0338402f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.465
cc_159 VPB N_A_27_74#_c_312_n 0.0350559f $X=-0.19 $Y=1.66 $X2=2.375 $Y2=2.09
cc_160 VPB N_A_27_74#_c_313_n 0.0129728f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.09
cc_161 VPB N_A_27_74#_c_314_n 0.00601783f $X=-0.19 $Y=1.66 $X2=2.535 $Y2=1.995
cc_162 VPB N_SCE_c_393_n 0.0264922f $X=-0.19 $Y=1.66 $X2=0.135 $Y2=2.32
cc_163 VPB N_SCE_c_394_n 0.0318721f $X=-0.19 $Y=1.66 $X2=1.41 $Y2=1.01
cc_164 VPB N_SCE_c_395_n 0.0231924f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.615
cc_165 VPB N_SCE_c_396_n 0.0275749f $X=-0.19 $Y=1.66 $X2=2.495 $Y2=2.245
cc_166 VPB N_SCE_c_387_n 0.00782879f $X=-0.19 $Y=1.66 $X2=0.2 $Y2=2.005
cc_167 VPB N_SCE_c_388_n 0.0410982f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.175
cc_168 VPB N_SCE_c_390_n 0.00293105f $X=-0.19 $Y=1.66 $X2=0.365 $Y2=1.1
cc_169 VPB N_SCE_c_392_n 0.00270951f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_170 VPB N_D_c_471_n 0.0301353f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_171 VPB N_D_c_476_n 0.0220363f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_172 VPB N_SCD_c_521_n 0.0170214f $X=-0.19 $Y=1.66 $X2=0.135 $Y2=0.37
cc_173 VPB N_SCD_c_518_n 0.0470646f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.615
cc_174 VPB SCD 0.00449661f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.615
cc_175 VPB N_CLK_c_560_n 0.00770267f $X=-0.19 $Y=1.66 $X2=0.135 $Y2=0.37
cc_176 VPB N_CLK_M1030_g 0.0230821f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_177 VPB N_A_1034_392#_c_635_n 0.0145245f $X=-0.19 $Y=1.66 $X2=1.14 $Y2=1.01
cc_178 VPB N_A_1034_392#_c_636_n 0.0198142f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.935
cc_179 VPB N_A_1034_392#_c_614_n 0.0146437f $X=-0.19 $Y=1.66 $X2=2.495 $Y2=2.245
cc_180 VPB N_A_1034_392#_c_638_n 0.057308f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.465
cc_181 VPB N_A_1034_392#_c_623_n 0.00475099f $X=-0.19 $Y=1.66 $X2=2.54 $Y2=1.995
cc_182 VPB N_A_1034_392#_c_624_n 0.00196266f $X=-0.19 $Y=1.66 $X2=2.535
+ $Y2=1.995
cc_183 VPB N_A_1034_392#_c_629_n 0.00112381f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_184 VPB N_A_1034_392#_c_642_n 0.00501177f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_185 VPB N_A_1034_392#_c_634_n 0.0202385f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_186 VPB N_A_1367_112#_c_848_n 0.0136749f $X=-0.19 $Y=1.66 $X2=2.495 $Y2=2.245
cc_187 VPB N_A_1367_112#_c_849_n 0.0212139f $X=-0.19 $Y=1.66 $X2=2.495 $Y2=2.64
cc_188 VPB N_A_1367_112#_c_844_n 0.00199812f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_189 VPB N_A_1367_112#_c_845_n 0.0359673f $X=-0.19 $Y=1.66 $X2=0.2 $Y2=1.265
cc_190 VPB N_A_1367_112#_c_847_n 7.08723e-19 $X=-0.19 $Y=1.66 $X2=0.365 $Y2=1.1
cc_191 VPB N_A_1367_112#_c_853_n 0.00336227f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.1
cc_192 VPB N_RESET_B_c_953_n 0.0101791f $X=-0.19 $Y=1.66 $X2=0.135 $Y2=2.32
cc_193 VPB N_RESET_B_c_964_n 0.0216256f $X=-0.19 $Y=1.66 $X2=1.41 $Y2=1.01
cc_194 VPB N_RESET_B_c_965_n 0.0167099f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_195 VPB N_RESET_B_c_960_n 0.0106437f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.465
cc_196 VPB N_RESET_B_M1038_g 0.00996849f $X=-0.19 $Y=1.66 $X2=0.365 $Y2=1.1
cc_197 VPB N_RESET_B_c_968_n 0.0149978f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.1
cc_198 VPB N_RESET_B_c_969_n 0.0251375f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_199 VPB N_RESET_B_c_970_n 0.0200891f $X=-0.19 $Y=1.66 $X2=2.54 $Y2=1.995
cc_200 VPB N_RESET_B_c_971_n 0.00163741f $X=-0.19 $Y=1.66 $X2=2.535 $Y2=1.995
cc_201 VPB N_RESET_B_c_972_n 0.0213442f $X=-0.19 $Y=1.66 $X2=2.535 $Y2=1.995
cc_202 VPB N_RESET_B_c_973_n 0.00238517f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_203 VPB N_RESET_B_c_974_n 0.00204342f $X=-0.19 $Y=1.66 $X2=2.535 $Y2=1.995
cc_204 VPB RESET_B 0.00336207f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_205 VPB N_RESET_B_c_976_n 0.0658019f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_206 VPB N_RESET_B_c_977_n 0.00235058f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_207 VPB N_RESET_B_c_978_n 0.0621565f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_208 VPB N_RESET_B_c_979_n 0.00478311f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_209 VPB N_RESET_B_c_980_n 0.0461401f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_210 VPB N_A_1236_138#_c_1180_n 0.0157054f $X=-0.19 $Y=1.66 $X2=2.495 $Y2=2.64
cc_211 VPB N_A_1236_138#_c_1188_n 0.0155175f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=0.58
cc_212 VPB N_A_1236_138#_c_1189_n 0.00306925f $X=-0.19 $Y=1.66 $X2=0.2 $Y2=1.265
cc_213 VPB N_A_1236_138#_c_1181_n 0.00749107f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.1
cc_214 VPB N_A_1236_138#_c_1182_n 0.0121924f $X=-0.19 $Y=1.66 $X2=2.375 $Y2=2.09
cc_215 VPB N_A_1236_138#_c_1185_n 0.00783535f $X=-0.19 $Y=1.66 $X2=2.54
+ $Y2=1.995
cc_216 VPB N_A_1236_138#_c_1193_n 0.00186797f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_217 VPB N_A_837_98#_M1034_g 0.020297f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.935
cc_218 VPB N_A_837_98#_c_1316_n 0.07521f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=0.58
cc_219 VPB N_A_837_98#_c_1329_n 0.0586461f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_220 VPB N_A_837_98#_c_1330_n 0.0123764f $X=-0.19 $Y=1.66 $X2=0.2 $Y2=1.265
cc_221 VPB N_A_837_98#_c_1331_n 0.00718351f $X=-0.19 $Y=1.66 $X2=0.365 $Y2=1.1
cc_222 VPB N_A_837_98#_c_1332_n 0.0163876f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.1
cc_223 VPB N_A_837_98#_c_1333_n 0.0160547f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.1
cc_224 VPB N_A_837_98#_c_1334_n 0.186352f $X=-0.19 $Y=1.66 $X2=2.375 $Y2=2.09
cc_225 VPB N_A_837_98#_c_1335_n 0.00735052f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.1
cc_226 VPB N_A_837_98#_c_1336_n 0.0131075f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.09
cc_227 VPB N_A_837_98#_M1042_g 0.0082806f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_228 VPB N_A_837_98#_c_1319_n 0.0195614f $X=-0.19 $Y=1.66 $X2=2.54 $Y2=2.09
cc_229 VPB N_A_837_98#_c_1320_n 0.00360844f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_230 VPB N_A_837_98#_c_1340_n 0.0089864f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_231 VPB N_A_837_98#_c_1341_n 0.00353228f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_232 VPB N_A_837_98#_c_1342_n 0.00280642f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_233 VPB N_A_837_98#_c_1324_n 0.00157987f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_234 VPB N_A_837_98#_c_1325_n 0.00618994f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_235 VPB N_A_2003_48#_c_1520_n 0.0412197f $X=-0.19 $Y=1.66 $X2=2.495 $Y2=2.245
cc_236 VPB N_A_2003_48#_c_1529_n 0.0232955f $X=-0.19 $Y=1.66 $X2=2.495 $Y2=2.64
cc_237 VPB N_A_2003_48#_c_1530_n 0.00836779f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.09
cc_238 VPB N_A_2003_48#_c_1526_n 0.0185734f $X=-0.19 $Y=1.66 $X2=2.54 $Y2=1.995
cc_239 VPB N_A_1745_74#_c_1609_n 3.48694e-19 $X=-0.19 $Y=1.66 $X2=2.495
+ $Y2=2.245
cc_240 VPB N_A_1745_74#_c_1624_n 0.0451105f $X=-0.19 $Y=1.66 $X2=2.495 $Y2=2.64
cc_241 VPB N_A_1745_74#_c_1625_n 0.0242804f $X=-0.19 $Y=1.66 $X2=2.495 $Y2=2.64
cc_242 VPB N_A_1745_74#_c_1626_n 0.0157526f $X=-0.19 $Y=1.66 $X2=0.2 $Y2=1.265
cc_243 VPB N_A_1745_74#_c_1613_n 0.0115338f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.1
cc_244 VPB N_A_1745_74#_c_1628_n 0.0157765f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_245 VPB N_A_1745_74#_c_1615_n 0.00496747f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.09
cc_246 VPB N_A_1745_74#_c_1630_n 0.00176961f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_247 VPB N_A_1745_74#_c_1618_n 0.00118746f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_248 VPB N_A_1745_74#_c_1632_n 0.0080022f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_249 VPB N_A_1745_74#_c_1633_n 0.00237571f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_250 VPB N_A_1745_74#_c_1634_n 0.00700686f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_251 VPB N_A_2339_74#_c_1783_n 0.0160879f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=0.935
cc_252 VPB N_A_2339_74#_c_1784_n 0.0148316f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_253 VPB N_A_2339_74#_c_1785_n 0.0143946f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.175
cc_254 VPB N_A_2339_74#_c_1786_n 0.0165543f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.1
cc_255 VPB N_A_2339_74#_c_1779_n 0.00394633f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_256 VPB N_A_2339_74#_c_1782_n 0.0271172f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_257 VPB N_VPWR_c_1890_n 0.0066125f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.09
cc_258 VPB N_VPWR_c_1891_n 0.00396467f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_259 VPB N_VPWR_c_1892_n 0.013846f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_260 VPB N_VPWR_c_1893_n 0.0230775f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_261 VPB N_VPWR_c_1894_n 0.0142717f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_262 VPB N_VPWR_c_1895_n 0.0137486f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_263 VPB N_VPWR_c_1896_n 0.0277893f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_264 VPB N_VPWR_c_1897_n 0.0214037f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_265 VPB N_VPWR_c_1898_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_266 VPB N_VPWR_c_1899_n 0.00508939f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_267 VPB N_VPWR_c_1900_n 0.0115177f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_268 VPB N_VPWR_c_1901_n 0.0443867f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_269 VPB N_VPWR_c_1902_n 0.0349943f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_270 VPB N_VPWR_c_1903_n 0.00601569f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_271 VPB N_VPWR_c_1904_n 0.0520927f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_272 VPB N_VPWR_c_1905_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_273 VPB N_VPWR_c_1906_n 0.0191816f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_274 VPB N_VPWR_c_1907_n 0.0457766f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_275 VPB N_VPWR_c_1908_n 0.0593f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_276 VPB N_VPWR_c_1909_n 0.0245819f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_277 VPB N_VPWR_c_1910_n 0.0218508f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_278 VPB N_VPWR_c_1911_n 0.0173667f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_279 VPB N_VPWR_c_1912_n 0.0312859f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_280 VPB N_VPWR_c_1913_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_281 VPB N_VPWR_c_1914_n 0.00463502f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_282 VPB N_VPWR_c_1915_n 0.00223798f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_283 VPB N_VPWR_c_1916_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_284 VPB N_VPWR_c_1917_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_285 VPB N_VPWR_c_1918_n 0.00460249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_286 VPB N_VPWR_c_1889_n 0.136411f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_287 VPB N_A_415_81#_c_2085_n 0.00482721f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.1
cc_288 VPB N_A_415_81#_c_2091_n 0.00312097f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.1
cc_289 VPB N_A_415_81#_c_2092_n 0.00523828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_290 VPB N_A_415_81#_c_2093_n 0.00723707f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.1
cc_291 VPB N_A_415_81#_c_2094_n 0.00195598f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_292 VPB N_A_415_81#_c_2089_n 0.00581282f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_293 VPB N_A_415_81#_c_2096_n 0.00257025f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_294 VPB N_A_415_81#_c_2097_n 0.0106179f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_295 VPB N_A_415_81#_c_2098_n 0.00833017f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_296 VPB N_Q_c_2249_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.175
cc_297 VPB N_Q_c_2250_n 0.0023624f $X=-0.19 $Y=1.66 $X2=0.365 $Y2=1.1
cc_298 VPB N_Q_c_2251_n 0.00183442f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.1
cc_299 VPB N_Q_c_2252_n 0.00221952f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_300 VPB Q 0.0136248f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.01
cc_301 N_A_27_74#_c_312_n N_SCE_c_393_n 0.0121883f $X=2.375 $Y=2.09 $X2=0 $Y2=0
cc_302 N_A_27_74#_c_313_n N_SCE_c_393_n 0.00496169f $X=0.28 $Y=2.09 $X2=0 $Y2=0
cc_303 N_A_27_74#_c_304_n N_SCE_M1036_g 0.00686809f $X=0.28 $Y=0.58 $X2=0 $Y2=0
cc_304 N_A_27_74#_c_305_n N_SCE_M1036_g 0.00830473f $X=0.2 $Y=2.005 $X2=0 $Y2=0
cc_305 N_A_27_74#_c_306_n N_SCE_M1036_g 0.0281157f $X=0.975 $Y=1.1 $X2=0 $Y2=0
cc_306 N_A_27_74#_c_308_n N_SCE_M1036_g 0.0181297f $X=0.975 $Y=1.01 $X2=0 $Y2=0
cc_307 N_A_27_74#_c_311_n N_SCE_c_394_n 0.0173713f $X=0.28 $Y=2.465 $X2=0 $Y2=0
cc_308 N_A_27_74#_c_312_n N_SCE_c_394_n 0.00721429f $X=2.375 $Y=2.09 $X2=0 $Y2=0
cc_309 N_A_27_74#_c_313_n N_SCE_c_394_n 4.59028e-19 $X=0.28 $Y=2.09 $X2=0 $Y2=0
cc_310 N_A_27_74#_c_312_n N_SCE_c_395_n 0.0100663f $X=2.375 $Y=2.09 $X2=0 $Y2=0
cc_311 N_A_27_74#_c_312_n N_SCE_c_396_n 0.00784761f $X=2.375 $Y=2.09 $X2=0 $Y2=0
cc_312 N_A_27_74#_c_309_n N_SCE_c_385_n 0.0165585f $X=2.495 $Y=2.245 $X2=0 $Y2=0
cc_313 N_A_27_74#_c_314_n N_SCE_c_385_n 3.29506e-19 $X=2.535 $Y=1.995 $X2=0
+ $Y2=0
cc_314 N_A_27_74#_c_305_n N_SCE_c_387_n 0.0158921f $X=0.2 $Y=2.005 $X2=0 $Y2=0
cc_315 N_A_27_74#_c_306_n N_SCE_c_387_n 0.00162366f $X=0.975 $Y=1.1 $X2=0 $Y2=0
cc_316 N_A_27_74#_c_302_n N_SCE_c_388_n 0.0106974f $X=1.41 $Y=1.01 $X2=0 $Y2=0
cc_317 N_A_27_74#_c_306_n N_SCE_c_388_n 0.00180358f $X=0.975 $Y=1.1 $X2=0 $Y2=0
cc_318 N_A_27_74#_c_312_n N_SCE_c_388_n 0.0170396f $X=2.375 $Y=2.09 $X2=0 $Y2=0
cc_319 N_A_27_74#_c_308_n N_SCE_c_388_n 0.0175645f $X=0.975 $Y=1.01 $X2=0 $Y2=0
cc_320 N_A_27_74#_c_309_n N_SCE_c_389_n 3.4369e-19 $X=2.495 $Y=2.245 $X2=0 $Y2=0
cc_321 N_A_27_74#_c_312_n N_SCE_c_389_n 0.0253366f $X=2.375 $Y=2.09 $X2=0 $Y2=0
cc_322 N_A_27_74#_c_314_n N_SCE_c_389_n 0.00219771f $X=2.535 $Y=1.995 $X2=0
+ $Y2=0
cc_323 N_A_27_74#_c_309_n N_SCE_c_390_n 0.0010238f $X=2.495 $Y=2.245 $X2=0 $Y2=0
cc_324 N_A_27_74#_c_314_n N_SCE_c_390_n 0.0242771f $X=2.535 $Y=1.995 $X2=0 $Y2=0
cc_325 N_A_27_74#_c_302_n N_SCE_c_391_n 0.00818136f $X=1.41 $Y=1.01 $X2=0 $Y2=0
cc_326 N_A_27_74#_c_305_n N_SCE_c_391_n 0.0170838f $X=0.2 $Y=2.005 $X2=0 $Y2=0
cc_327 N_A_27_74#_c_306_n N_SCE_c_391_n 0.0353374f $X=0.975 $Y=1.1 $X2=0 $Y2=0
cc_328 N_A_27_74#_c_312_n N_SCE_c_391_n 0.0893268f $X=2.375 $Y=2.09 $X2=0 $Y2=0
cc_329 N_A_27_74#_c_308_n N_SCE_c_391_n 0.00202099f $X=0.975 $Y=1.01 $X2=0 $Y2=0
cc_330 N_A_27_74#_c_309_n N_D_c_471_n 0.0188152f $X=2.495 $Y=2.245 $X2=0 $Y2=0
cc_331 N_A_27_74#_c_312_n N_D_c_471_n 0.0091263f $X=2.375 $Y=2.09 $X2=0 $Y2=0
cc_332 N_A_27_74#_c_314_n N_D_c_471_n 0.00124819f $X=2.535 $Y=1.995 $X2=0 $Y2=0
cc_333 N_A_27_74#_c_309_n N_D_c_476_n 0.0140909f $X=2.495 $Y=2.245 $X2=0 $Y2=0
cc_334 N_A_27_74#_c_312_n N_D_c_476_n 0.00753484f $X=2.375 $Y=2.09 $X2=0 $Y2=0
cc_335 N_A_27_74#_c_302_n N_D_c_472_n 0.00979811f $X=1.41 $Y=1.01 $X2=0 $Y2=0
cc_336 N_A_27_74#_c_306_n N_D_c_472_n 2.46751e-19 $X=0.975 $Y=1.1 $X2=0 $Y2=0
cc_337 N_A_27_74#_c_308_n N_D_c_472_n 0.00223479f $X=0.975 $Y=1.01 $X2=0 $Y2=0
cc_338 N_A_27_74#_c_303_n N_D_c_473_n 0.00580814f $X=1.485 $Y=0.935 $X2=0 $Y2=0
cc_339 N_A_27_74#_c_306_n N_D_c_473_n 0.0143876f $X=0.975 $Y=1.1 $X2=0 $Y2=0
cc_340 N_A_27_74#_c_308_n N_D_c_473_n 8.79717e-19 $X=0.975 $Y=1.01 $X2=0 $Y2=0
cc_341 N_A_27_74#_c_303_n N_D_c_474_n 0.0224455f $X=1.485 $Y=0.935 $X2=0 $Y2=0
cc_342 N_A_27_74#_c_309_n N_SCD_c_521_n 0.0258628f $X=2.495 $Y=2.245 $X2=-0.19
+ $Y2=-0.245
cc_343 N_A_27_74#_c_309_n N_SCD_c_518_n 0.0208734f $X=2.495 $Y=2.245 $X2=0 $Y2=0
cc_344 N_A_27_74#_c_314_n N_SCD_c_518_n 0.00250603f $X=2.535 $Y=1.995 $X2=0
+ $Y2=0
cc_345 N_A_27_74#_c_309_n SCD 4.02276e-19 $X=2.495 $Y=2.245 $X2=0 $Y2=0
cc_346 N_A_27_74#_c_314_n SCD 0.0195546f $X=2.535 $Y=1.995 $X2=0 $Y2=0
cc_347 N_A_27_74#_c_309_n N_VPWR_c_1890_n 0.00141778f $X=2.495 $Y=2.245 $X2=0
+ $Y2=0
cc_348 N_A_27_74#_c_311_n N_VPWR_c_1906_n 0.0145938f $X=0.28 $Y=2.465 $X2=0
+ $Y2=0
cc_349 N_A_27_74#_c_309_n N_VPWR_c_1907_n 0.00445602f $X=2.495 $Y=2.245 $X2=0
+ $Y2=0
cc_350 N_A_27_74#_c_311_n N_VPWR_c_1912_n 0.0247088f $X=0.28 $Y=2.465 $X2=0
+ $Y2=0
cc_351 N_A_27_74#_c_312_n N_VPWR_c_1912_n 0.0746993f $X=2.375 $Y=2.09 $X2=0
+ $Y2=0
cc_352 N_A_27_74#_c_309_n N_VPWR_c_1889_n 0.00448781f $X=2.495 $Y=2.245 $X2=0
+ $Y2=0
cc_353 N_A_27_74#_c_311_n N_VPWR_c_1889_n 0.0120466f $X=0.28 $Y=2.465 $X2=0
+ $Y2=0
cc_354 N_A_27_74#_c_309_n N_A_415_81#_c_2099_n 0.0101811f $X=2.495 $Y=2.245
+ $X2=0 $Y2=0
cc_355 N_A_27_74#_c_314_n N_A_415_81#_c_2099_n 0.0180834f $X=2.535 $Y=1.995
+ $X2=0 $Y2=0
cc_356 N_A_27_74#_c_309_n N_A_415_81#_c_2096_n 0.00974144f $X=2.495 $Y=2.245
+ $X2=0 $Y2=0
cc_357 N_A_27_74#_c_312_n N_A_415_81#_c_2096_n 0.0189432f $X=2.375 $Y=2.09 $X2=0
+ $Y2=0
cc_358 N_A_27_74#_c_314_n N_A_415_81#_c_2096_n 0.00295889f $X=2.535 $Y=1.995
+ $X2=0 $Y2=0
cc_359 N_A_27_74#_c_303_n N_VGND_c_2312_n 0.00287309f $X=1.485 $Y=0.935 $X2=0
+ $Y2=0
cc_360 N_A_27_74#_c_304_n N_VGND_c_2312_n 0.0156021f $X=0.28 $Y=0.58 $X2=0 $Y2=0
cc_361 N_A_27_74#_c_306_n N_VGND_c_2312_n 0.0254818f $X=0.975 $Y=1.1 $X2=0 $Y2=0
cc_362 N_A_27_74#_c_308_n N_VGND_c_2312_n 0.00149092f $X=0.975 $Y=1.01 $X2=0
+ $Y2=0
cc_363 N_A_27_74#_c_303_n N_VGND_c_2320_n 9.09582e-19 $X=1.485 $Y=0.935 $X2=0
+ $Y2=0
cc_364 N_A_27_74#_c_304_n N_VGND_c_2322_n 0.011066f $X=0.28 $Y=0.58 $X2=0 $Y2=0
cc_365 N_A_27_74#_c_304_n N_VGND_c_2334_n 0.00915947f $X=0.28 $Y=0.58 $X2=0
+ $Y2=0
cc_366 N_A_27_74#_c_303_n N_noxref_24_c_2457_n 0.011495f $X=1.485 $Y=0.935 $X2=0
+ $Y2=0
cc_367 N_A_27_74#_c_303_n N_noxref_24_c_2458_n 0.00899724f $X=1.485 $Y=0.935
+ $X2=0 $Y2=0
cc_368 N_A_27_74#_c_306_n N_noxref_24_c_2458_n 0.00178881f $X=0.975 $Y=1.1 $X2=0
+ $Y2=0
cc_369 N_A_27_74#_c_308_n N_noxref_24_c_2458_n 0.00859402f $X=0.975 $Y=1.01
+ $X2=0 $Y2=0
cc_370 N_SCE_c_388_n N_D_c_471_n 0.0203026f $X=1.535 $Y=1.67 $X2=0 $Y2=0
cc_371 N_SCE_c_389_n N_D_c_471_n 0.0146216f $X=2.405 $Y=1.575 $X2=0 $Y2=0
cc_372 N_SCE_c_390_n N_D_c_471_n 3.20022e-19 $X=2.565 $Y=1.425 $X2=0 $Y2=0
cc_373 N_SCE_c_392_n N_D_c_471_n 0.00479409f $X=1.795 $Y=1.662 $X2=0 $Y2=0
cc_374 N_SCE_c_395_n N_D_c_476_n 0.0203026f $X=1.625 $Y=2.155 $X2=0 $Y2=0
cc_375 N_SCE_c_396_n N_D_c_476_n 0.0373591f $X=1.625 $Y=2.245 $X2=0 $Y2=0
cc_376 N_SCE_c_385_n N_D_c_472_n 0.0227885f $X=2.785 $Y=1.05 $X2=0 $Y2=0
cc_377 N_SCE_M1037_g N_D_c_472_n 0.00179056f $X=2.785 $Y=0.615 $X2=0 $Y2=0
cc_378 N_SCE_c_390_n N_D_c_472_n 0.00147436f $X=2.565 $Y=1.425 $X2=0 $Y2=0
cc_379 N_SCE_c_392_n N_D_c_472_n 0.00411836f $X=1.795 $Y=1.662 $X2=0 $Y2=0
cc_380 N_SCE_c_385_n N_D_c_473_n 9.80386e-19 $X=2.785 $Y=1.05 $X2=0 $Y2=0
cc_381 N_SCE_M1037_g N_D_c_473_n 4.78719e-19 $X=2.785 $Y=0.615 $X2=0 $Y2=0
cc_382 N_SCE_c_388_n N_D_c_473_n 0.00106377f $X=1.535 $Y=1.67 $X2=0 $Y2=0
cc_383 N_SCE_c_391_n N_D_c_473_n 0.0344941f $X=1.623 $Y=1.662 $X2=0 $Y2=0
cc_384 N_SCE_M1037_g N_D_c_474_n 0.00976046f $X=2.785 $Y=0.615 $X2=0 $Y2=0
cc_385 N_SCE_c_385_n N_SCD_M1040_g 0.0083988f $X=2.785 $Y=1.05 $X2=0 $Y2=0
cc_386 N_SCE_M1037_g N_SCD_M1040_g 0.0576059f $X=2.785 $Y=0.615 $X2=0 $Y2=0
cc_387 N_SCE_c_390_n N_SCD_M1040_g 0.00357167f $X=2.565 $Y=1.425 $X2=0 $Y2=0
cc_388 N_SCE_c_390_n SCD 0.014834f $X=2.565 $Y=1.425 $X2=0 $Y2=0
cc_389 N_SCE_c_385_n N_SCD_c_520_n 0.00942916f $X=2.785 $Y=1.05 $X2=0 $Y2=0
cc_390 N_SCE_c_390_n N_SCD_c_520_n 0.0024124f $X=2.565 $Y=1.425 $X2=0 $Y2=0
cc_391 N_SCE_c_394_n N_VPWR_c_1906_n 0.00445602f $X=0.505 $Y=2.245 $X2=0 $Y2=0
cc_392 N_SCE_c_396_n N_VPWR_c_1907_n 0.00415318f $X=1.625 $Y=2.245 $X2=0 $Y2=0
cc_393 N_SCE_c_394_n N_VPWR_c_1912_n 0.017697f $X=0.505 $Y=2.245 $X2=0 $Y2=0
cc_394 N_SCE_c_396_n N_VPWR_c_1912_n 0.0163904f $X=1.625 $Y=2.245 $X2=0 $Y2=0
cc_395 N_SCE_c_394_n N_VPWR_c_1889_n 0.00865213f $X=0.505 $Y=2.245 $X2=0 $Y2=0
cc_396 N_SCE_c_396_n N_VPWR_c_1889_n 0.00817532f $X=1.625 $Y=2.245 $X2=0 $Y2=0
cc_397 N_SCE_c_385_n N_A_415_81#_c_2083_n 0.0072321f $X=2.785 $Y=1.05 $X2=0
+ $Y2=0
cc_398 N_SCE_M1037_g N_A_415_81#_c_2083_n 0.0127864f $X=2.785 $Y=0.615 $X2=0
+ $Y2=0
cc_399 N_SCE_c_389_n N_A_415_81#_c_2083_n 0.0041139f $X=2.405 $Y=1.575 $X2=0
+ $Y2=0
cc_400 N_SCE_c_390_n N_A_415_81#_c_2083_n 0.0198392f $X=2.565 $Y=1.425 $X2=0
+ $Y2=0
cc_401 N_SCE_c_385_n N_A_415_81#_c_2084_n 0.0056718f $X=2.785 $Y=1.05 $X2=0
+ $Y2=0
cc_402 N_SCE_M1037_g N_A_415_81#_c_2084_n 0.00612765f $X=2.785 $Y=0.615 $X2=0
+ $Y2=0
cc_403 N_SCE_c_396_n N_A_415_81#_c_2096_n 0.00182961f $X=1.625 $Y=2.245 $X2=0
+ $Y2=0
cc_404 N_SCE_M1036_g N_VGND_c_2312_n 0.0129468f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_405 N_SCE_M1037_g N_VGND_c_2320_n 9.15902e-19 $X=2.785 $Y=0.615 $X2=0 $Y2=0
cc_406 N_SCE_M1036_g N_VGND_c_2322_n 0.00383152f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_407 N_SCE_M1036_g N_VGND_c_2334_n 0.00761198f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_408 N_SCE_c_385_n N_noxref_24_c_2457_n 3.08157e-19 $X=2.785 $Y=1.05 $X2=0
+ $Y2=0
cc_409 N_SCE_M1037_g N_noxref_24_c_2457_n 0.0119336f $X=2.785 $Y=0.615 $X2=0
+ $Y2=0
cc_410 N_SCE_M1036_g N_noxref_24_c_2458_n 9.19966e-19 $X=0.495 $Y=0.58 $X2=0
+ $Y2=0
cc_411 N_D_c_476_n N_VPWR_c_1907_n 0.00445602f $X=2.045 $Y=2.245 $X2=0 $Y2=0
cc_412 N_D_c_476_n N_VPWR_c_1912_n 0.00236192f $X=2.045 $Y=2.245 $X2=0 $Y2=0
cc_413 N_D_c_476_n N_VPWR_c_1889_n 0.00858241f $X=2.045 $Y=2.245 $X2=0 $Y2=0
cc_414 N_D_c_472_n N_A_415_81#_c_2083_n 0.00121844f $X=1.935 $Y=1.1 $X2=0 $Y2=0
cc_415 N_D_c_473_n N_A_415_81#_c_2083_n 0.0115884f $X=1.935 $Y=1.1 $X2=0 $Y2=0
cc_416 N_D_c_474_n N_A_415_81#_c_2083_n 0.00599383f $X=1.952 $Y=0.935 $X2=0
+ $Y2=0
cc_417 N_D_c_476_n N_A_415_81#_c_2096_n 0.0112736f $X=2.045 $Y=2.245 $X2=0 $Y2=0
cc_418 N_D_c_474_n N_VGND_c_2320_n 9.15902e-19 $X=1.952 $Y=0.935 $X2=0 $Y2=0
cc_419 N_D_c_472_n N_noxref_24_c_2457_n 0.00121903f $X=1.935 $Y=1.1 $X2=0 $Y2=0
cc_420 N_D_c_473_n N_noxref_24_c_2457_n 0.014028f $X=1.935 $Y=1.1 $X2=0 $Y2=0
cc_421 N_D_c_474_n N_noxref_24_c_2457_n 0.0125454f $X=1.952 $Y=0.935 $X2=0 $Y2=0
cc_422 N_D_c_474_n N_noxref_24_c_2458_n 0.00108287f $X=1.952 $Y=0.935 $X2=0
+ $Y2=0
cc_423 N_D_c_473_n noxref_25 0.00395662f $X=1.935 $Y=1.1 $X2=-0.19 $Y2=-0.245
cc_424 SCD N_RESET_B_c_953_n 0.00216554f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_425 N_SCD_c_520_n N_RESET_B_c_953_n 0.021668f $X=3.105 $Y=1.605 $X2=0 $Y2=0
cc_426 N_SCD_M1040_g N_RESET_B_M1012_g 0.0149708f $X=3.145 $Y=0.615 $X2=0 $Y2=0
cc_427 N_SCD_c_521_n N_RESET_B_c_964_n 0.0163024f $X=3.035 $Y=2.245 $X2=0 $Y2=0
cc_428 N_SCD_M1040_g N_RESET_B_c_962_n 0.0219591f $X=3.145 $Y=0.615 $X2=0 $Y2=0
cc_429 N_SCD_c_518_n N_RESET_B_c_976_n 0.0259291f $X=3.105 $Y=1.945 $X2=0 $Y2=0
cc_430 N_SCD_c_521_n N_VPWR_c_1890_n 0.0100582f $X=3.035 $Y=2.245 $X2=0 $Y2=0
cc_431 N_SCD_c_521_n N_VPWR_c_1907_n 0.00413917f $X=3.035 $Y=2.245 $X2=0 $Y2=0
cc_432 N_SCD_c_521_n N_VPWR_c_1889_n 0.00409681f $X=3.035 $Y=2.245 $X2=0 $Y2=0
cc_433 N_SCD_M1040_g N_A_415_81#_c_2083_n 0.00136969f $X=3.145 $Y=0.615 $X2=0
+ $Y2=0
cc_434 N_SCD_c_521_n N_A_415_81#_c_2099_n 0.0130079f $X=3.035 $Y=2.245 $X2=0
+ $Y2=0
cc_435 N_SCD_c_518_n N_A_415_81#_c_2099_n 7.93085e-19 $X=3.105 $Y=1.945 $X2=0
+ $Y2=0
cc_436 SCD N_A_415_81#_c_2099_n 0.0212424f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_437 N_SCD_M1040_g N_A_415_81#_c_2084_n 0.0124831f $X=3.145 $Y=0.615 $X2=0
+ $Y2=0
cc_438 SCD N_A_415_81#_c_2084_n 0.0147205f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_439 N_SCD_c_520_n N_A_415_81#_c_2084_n 0.00124535f $X=3.105 $Y=1.605 $X2=0
+ $Y2=0
cc_440 N_SCD_c_521_n N_A_415_81#_c_2085_n 0.00151656f $X=3.035 $Y=2.245 $X2=0
+ $Y2=0
cc_441 N_SCD_M1040_g N_A_415_81#_c_2085_n 0.00668437f $X=3.145 $Y=0.615 $X2=0
+ $Y2=0
cc_442 N_SCD_c_518_n N_A_415_81#_c_2085_n 0.00180807f $X=3.105 $Y=1.945 $X2=0
+ $Y2=0
cc_443 SCD N_A_415_81#_c_2085_n 0.0562719f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_444 N_SCD_c_520_n N_A_415_81#_c_2085_n 0.00193985f $X=3.105 $Y=1.605 $X2=0
+ $Y2=0
cc_445 N_SCD_c_521_n N_A_415_81#_c_2096_n 0.00167919f $X=3.035 $Y=2.245 $X2=0
+ $Y2=0
cc_446 N_SCD_c_521_n N_A_415_81#_c_2097_n 0.0010086f $X=3.035 $Y=2.245 $X2=0
+ $Y2=0
cc_447 N_SCD_M1040_g N_VGND_c_2320_n 9.15902e-19 $X=3.145 $Y=0.615 $X2=0 $Y2=0
cc_448 N_SCD_M1040_g N_noxref_24_c_2457_n 0.0107463f $X=3.145 $Y=0.615 $X2=0
+ $Y2=0
cc_449 N_CLK_c_560_n N_A_1034_392#_c_619_n 8.17254e-19 $X=4.605 $Y=1.41 $X2=0
+ $Y2=0
cc_450 N_CLK_M1030_g N_A_1034_392#_c_623_n 8.77169e-19 $X=4.645 $Y=2.46 $X2=0
+ $Y2=0
cc_451 N_CLK_c_560_n N_RESET_B_c_953_n 0.0241646f $X=4.605 $Y=1.41 $X2=0 $Y2=0
cc_452 CLK N_RESET_B_c_953_n 0.00303155f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_453 N_CLK_c_560_n N_RESET_B_c_955_n 0.0101115f $X=4.605 $Y=1.41 $X2=0 $Y2=0
cc_454 N_CLK_c_560_n N_RESET_B_c_970_n 0.00229617f $X=4.605 $Y=1.41 $X2=0 $Y2=0
cc_455 N_CLK_M1030_g N_RESET_B_c_970_n 0.00240204f $X=4.645 $Y=2.46 $X2=0 $Y2=0
cc_456 CLK N_RESET_B_c_970_n 0.00556699f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_457 N_CLK_c_560_n N_RESET_B_c_971_n 0.00134728f $X=4.605 $Y=1.41 $X2=0 $Y2=0
cc_458 CLK N_RESET_B_c_971_n 0.00376241f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_459 N_CLK_c_560_n N_RESET_B_c_976_n 0.0168483f $X=4.605 $Y=1.41 $X2=0 $Y2=0
cc_460 N_CLK_M1030_g N_RESET_B_c_976_n 0.00526706f $X=4.645 $Y=2.46 $X2=0 $Y2=0
cc_461 CLK N_RESET_B_c_976_n 9.14892e-19 $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_462 N_CLK_c_560_n N_RESET_B_c_977_n 0.00211095f $X=4.605 $Y=1.41 $X2=0 $Y2=0
cc_463 CLK N_RESET_B_c_977_n 0.0174898f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_464 CLK N_A_837_98#_M1010_s 0.00275914f $X=3.995 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_465 N_CLK_M1030_g N_A_837_98#_M1034_g 0.0407453f $X=4.645 $Y=2.46 $X2=0 $Y2=0
cc_466 N_CLK_c_560_n N_A_837_98#_c_1347_n 0.00591117f $X=4.605 $Y=1.41 $X2=0
+ $Y2=0
cc_467 N_CLK_c_560_n N_A_837_98#_c_1341_n 0.00172667f $X=4.605 $Y=1.41 $X2=0
+ $Y2=0
cc_468 N_CLK_M1030_g N_A_837_98#_c_1341_n 0.0123157f $X=4.645 $Y=2.46 $X2=0
+ $Y2=0
cc_469 CLK N_A_837_98#_c_1341_n 0.00625715f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_470 N_CLK_c_560_n N_A_837_98#_c_1351_n 0.0106749f $X=4.605 $Y=1.41 $X2=0
+ $Y2=0
cc_471 CLK N_A_837_98#_c_1351_n 0.00710736f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_472 N_CLK_c_560_n N_A_837_98#_c_1353_n 0.00382755f $X=4.605 $Y=1.41 $X2=0
+ $Y2=0
cc_473 CLK N_A_837_98#_c_1353_n 0.00911074f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_474 N_CLK_c_560_n N_A_837_98#_c_1322_n 0.00416568f $X=4.605 $Y=1.41 $X2=0
+ $Y2=0
cc_475 CLK N_A_837_98#_c_1322_n 0.0141873f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_476 N_CLK_c_560_n N_A_837_98#_c_1323_n 0.00694556f $X=4.605 $Y=1.41 $X2=0
+ $Y2=0
cc_477 CLK N_A_837_98#_c_1323_n 0.00725176f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_478 N_CLK_c_560_n N_A_837_98#_c_1342_n 0.00527775f $X=4.605 $Y=1.41 $X2=0
+ $Y2=0
cc_479 N_CLK_M1030_g N_A_837_98#_c_1342_n 4.68575e-19 $X=4.645 $Y=2.46 $X2=0
+ $Y2=0
cc_480 CLK N_A_837_98#_c_1342_n 0.0105132f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_481 N_CLK_c_560_n N_A_837_98#_c_1324_n 0.00758375f $X=4.605 $Y=1.41 $X2=0
+ $Y2=0
cc_482 CLK N_A_837_98#_c_1324_n 0.0155168f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_483 N_CLK_c_560_n N_A_837_98#_c_1325_n 0.0223101f $X=4.605 $Y=1.41 $X2=0
+ $Y2=0
cc_484 N_CLK_c_560_n N_A_837_98#_c_1326_n 0.02115f $X=4.605 $Y=1.41 $X2=0 $Y2=0
cc_485 N_CLK_M1030_g N_VPWR_c_1891_n 0.0164315f $X=4.645 $Y=2.46 $X2=0 $Y2=0
cc_486 N_CLK_M1030_g N_VPWR_c_1902_n 0.00303184f $X=4.645 $Y=2.46 $X2=0 $Y2=0
cc_487 N_CLK_M1030_g N_VPWR_c_1889_n 0.00397656f $X=4.645 $Y=2.46 $X2=0 $Y2=0
cc_488 N_CLK_c_560_n N_A_415_81#_c_2085_n 6.01825e-19 $X=4.605 $Y=1.41 $X2=0
+ $Y2=0
cc_489 CLK N_A_415_81#_c_2085_n 0.0250371f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_490 N_CLK_M1030_g N_A_415_81#_c_2091_n 0.00649883f $X=4.645 $Y=2.46 $X2=0
+ $Y2=0
cc_491 N_CLK_M1030_g N_A_415_81#_c_2097_n 0.0119582f $X=4.645 $Y=2.46 $X2=0
+ $Y2=0
cc_492 N_CLK_c_560_n N_A_415_81#_c_2098_n 4.49597e-19 $X=4.605 $Y=1.41 $X2=0
+ $Y2=0
cc_493 N_CLK_M1030_g N_A_415_81#_c_2098_n 0.00460785f $X=4.645 $Y=2.46 $X2=0
+ $Y2=0
cc_494 N_CLK_M1030_g N_A_415_81#_c_2135_n 0.00438299f $X=4.645 $Y=2.46 $X2=0
+ $Y2=0
cc_495 N_CLK_c_560_n N_VGND_c_2313_n 0.00375111f $X=4.605 $Y=1.41 $X2=0 $Y2=0
cc_496 CLK N_VGND_c_2313_n 0.00712523f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_497 N_CLK_c_560_n N_VGND_c_2314_n 0.00386191f $X=4.605 $Y=1.41 $X2=0 $Y2=0
cc_498 N_CLK_c_560_n N_VGND_c_2334_n 9.39239e-19 $X=4.605 $Y=1.41 $X2=0 $Y2=0
cc_499 N_A_1034_392#_c_626_n N_A_1367_112#_M1019_d 0.00224844f $X=8.825 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_500 N_A_1034_392#_M1041_g N_A_1367_112#_M1044_g 0.0328999f $X=6.535 $Y=0.9
+ $X2=0 $Y2=0
cc_501 N_A_1034_392#_c_621_n N_A_1367_112#_M1044_g 0.00321205f $X=7.055 $Y=0.415
+ $X2=0 $Y2=0
cc_502 N_A_1034_392#_c_631_n N_A_1367_112#_M1044_g 0.00342215f $X=7.14 $Y=0.415
+ $X2=0 $Y2=0
cc_503 N_A_1034_392#_c_635_n N_A_1367_112#_c_848_n 0.00142315f $X=6.135 $Y=2.15
+ $X2=0 $Y2=0
cc_504 N_A_1034_392#_c_636_n N_A_1367_112#_c_849_n 0.00142315f $X=6.135 $Y=2.24
+ $X2=0 $Y2=0
cc_505 N_A_1034_392#_c_635_n N_A_1367_112#_c_845_n 3.5795e-19 $X=6.135 $Y=2.15
+ $X2=0 $Y2=0
cc_506 N_A_1034_392#_c_614_n N_A_1367_112#_c_845_n 0.0328999f $X=6.46 $Y=1.66
+ $X2=0 $Y2=0
cc_507 N_A_1034_392#_c_634_n N_A_1367_112#_c_845_n 0.0023084f $X=6.065 $Y=1.66
+ $X2=0 $Y2=0
cc_508 N_A_1034_392#_c_625_n N_A_1367_112#_c_863_n 0.00761753f $X=7.93 $Y=0.665
+ $X2=0 $Y2=0
cc_509 N_A_1034_392#_c_631_n N_A_1367_112#_c_863_n 0.00974988f $X=7.14 $Y=0.415
+ $X2=0 $Y2=0
cc_510 N_A_1034_392#_c_618_n N_A_1367_112#_c_846_n 0.00476106f $X=8.725 $Y=1.16
+ $X2=0 $Y2=0
cc_511 N_A_1034_392#_c_629_n N_A_1367_112#_c_846_n 0.00539231f $X=9.33 $Y=2.065
+ $X2=0 $Y2=0
cc_512 N_A_1034_392#_c_633_n N_A_1367_112#_c_846_n 0.0108396f $X=9.33 $Y=1.07
+ $X2=0 $Y2=0
cc_513 N_A_1034_392#_c_618_n N_A_1367_112#_c_847_n 0.00855892f $X=8.725 $Y=1.16
+ $X2=0 $Y2=0
cc_514 N_A_1034_392#_c_629_n N_A_1367_112#_c_847_n 0.0129187f $X=9.33 $Y=2.065
+ $X2=0 $Y2=0
cc_515 N_A_1034_392#_c_633_n N_A_1367_112#_c_847_n 0.0180376f $X=9.33 $Y=1.07
+ $X2=0 $Y2=0
cc_516 N_A_1034_392#_c_638_n N_A_1367_112#_c_853_n 0.00106238f $X=9.835 $Y=2.465
+ $X2=0 $Y2=0
cc_517 N_A_1034_392#_c_629_n N_A_1367_112#_c_853_n 0.0240786f $X=9.33 $Y=2.065
+ $X2=0 $Y2=0
cc_518 N_A_1034_392#_c_665_p N_A_1367_112#_c_853_n 0.0118335f $X=9.415 $Y=2.222
+ $X2=0 $Y2=0
cc_519 N_A_1034_392#_c_625_n N_A_1367_112#_c_874_n 0.0484504f $X=7.93 $Y=0.665
+ $X2=0 $Y2=0
cc_520 N_A_1034_392#_c_626_n N_A_1367_112#_c_874_n 0.00422751f $X=8.825 $Y=0.34
+ $X2=0 $Y2=0
cc_521 N_A_1034_392#_c_616_n N_A_1367_112#_c_876_n 0.00932475f $X=8.65 $Y=1.085
+ $X2=0 $Y2=0
cc_522 N_A_1034_392#_c_618_n N_A_1367_112#_c_876_n 2.66567e-19 $X=8.725 $Y=1.16
+ $X2=0 $Y2=0
cc_523 N_A_1034_392#_c_626_n N_A_1367_112#_c_876_n 0.02112f $X=8.825 $Y=0.34
+ $X2=0 $Y2=0
cc_524 N_A_1034_392#_c_628_n N_A_1367_112#_c_876_n 0.0232075f $X=8.91 $Y=0.905
+ $X2=0 $Y2=0
cc_525 N_A_1034_392#_c_633_n N_A_1367_112#_c_876_n 0.0158476f $X=9.33 $Y=1.07
+ $X2=0 $Y2=0
cc_526 N_A_1034_392#_M1041_g N_RESET_B_c_955_n 0.00526413f $X=6.535 $Y=0.9 $X2=0
+ $Y2=0
cc_527 N_A_1034_392#_c_621_n N_RESET_B_c_955_n 0.0257323f $X=7.055 $Y=0.415
+ $X2=0 $Y2=0
cc_528 N_A_1034_392#_c_622_n N_RESET_B_c_955_n 0.009452f $X=5.62 $Y=0.415 $X2=0
+ $Y2=0
cc_529 N_A_1034_392#_c_631_n N_RESET_B_c_955_n 0.00184232f $X=7.14 $Y=0.415
+ $X2=0 $Y2=0
cc_530 N_A_1034_392#_c_625_n N_RESET_B_M1024_g 0.0116325f $X=7.93 $Y=0.665 $X2=0
+ $Y2=0
cc_531 N_A_1034_392#_c_678_p N_RESET_B_M1024_g 0.0035287f $X=8.015 $Y=0.58 $X2=0
+ $Y2=0
cc_532 N_A_1034_392#_c_627_n N_RESET_B_M1024_g 6.46496e-19 $X=8.1 $Y=0.34 $X2=0
+ $Y2=0
cc_533 N_A_1034_392#_c_631_n N_RESET_B_M1024_g 0.0104865f $X=7.14 $Y=0.415 $X2=0
+ $Y2=0
cc_534 N_A_1034_392#_c_635_n N_RESET_B_c_970_n 0.00393395f $X=6.135 $Y=2.15
+ $X2=0 $Y2=0
cc_535 N_A_1034_392#_c_614_n N_RESET_B_c_970_n 0.00414957f $X=6.46 $Y=1.66 $X2=0
+ $Y2=0
cc_536 N_A_1034_392#_c_623_n N_RESET_B_c_970_n 0.0385239f $X=5.655 $Y=1.75 $X2=0
+ $Y2=0
cc_537 N_A_1034_392#_c_624_n N_RESET_B_c_970_n 0.0163211f $X=6.065 $Y=1.75 $X2=0
+ $Y2=0
cc_538 N_A_1034_392#_c_634_n N_RESET_B_c_970_n 0.00388711f $X=6.065 $Y=1.66
+ $X2=0 $Y2=0
cc_539 N_A_1034_392#_c_638_n N_RESET_B_c_972_n 0.00245933f $X=9.835 $Y=2.465
+ $X2=0 $Y2=0
cc_540 N_A_1034_392#_c_629_n N_RESET_B_c_972_n 0.0104861f $X=9.33 $Y=2.065 $X2=0
+ $Y2=0
cc_541 N_A_1034_392#_c_665_p N_RESET_B_c_972_n 0.00467739f $X=9.415 $Y=2.222
+ $X2=0 $Y2=0
cc_542 N_A_1034_392#_c_642_n N_RESET_B_c_972_n 0.0172592f $X=9.79 $Y=2.215 $X2=0
+ $Y2=0
cc_543 N_A_1034_392#_c_616_n N_A_1236_138#_M1019_g 0.0216734f $X=8.65 $Y=1.085
+ $X2=0 $Y2=0
cc_544 N_A_1034_392#_c_625_n N_A_1236_138#_M1019_g 0.00459622f $X=7.93 $Y=0.665
+ $X2=0 $Y2=0
cc_545 N_A_1034_392#_c_626_n N_A_1236_138#_M1019_g 0.00898149f $X=8.825 $Y=0.34
+ $X2=0 $Y2=0
cc_546 N_A_1034_392#_c_627_n N_A_1236_138#_M1019_g 0.00298755f $X=8.1 $Y=0.34
+ $X2=0 $Y2=0
cc_547 N_A_1034_392#_c_618_n N_A_1236_138#_c_1180_n 0.0121912f $X=8.725 $Y=1.16
+ $X2=0 $Y2=0
cc_548 N_A_1034_392#_c_629_n N_A_1236_138#_c_1180_n 3.24532e-19 $X=9.33 $Y=2.065
+ $X2=0 $Y2=0
cc_549 N_A_1034_392#_c_636_n N_A_1236_138#_c_1189_n 0.00181918f $X=6.135 $Y=2.24
+ $X2=0 $Y2=0
cc_550 N_A_1034_392#_c_614_n N_A_1236_138#_c_1189_n 7.58927e-19 $X=6.46 $Y=1.66
+ $X2=0 $Y2=0
cc_551 N_A_1034_392#_M1041_g N_A_1236_138#_c_1202_n 0.0106114f $X=6.535 $Y=0.9
+ $X2=0 $Y2=0
cc_552 N_A_1034_392#_c_621_n N_A_1236_138#_c_1202_n 0.0143503f $X=7.055 $Y=0.415
+ $X2=0 $Y2=0
cc_553 N_A_1034_392#_c_635_n N_A_1236_138#_c_1181_n 3.69789e-19 $X=6.135 $Y=2.15
+ $X2=0 $Y2=0
cc_554 N_A_1034_392#_M1041_g N_A_1236_138#_c_1181_n 0.00662576f $X=6.535 $Y=0.9
+ $X2=0 $Y2=0
cc_555 N_A_1034_392#_c_614_n N_A_1236_138#_c_1186_n 4.38542e-19 $X=6.46 $Y=1.66
+ $X2=0 $Y2=0
cc_556 N_A_1034_392#_M1041_g N_A_1236_138#_c_1186_n 0.00504454f $X=6.535 $Y=0.9
+ $X2=0 $Y2=0
cc_557 N_A_1034_392#_c_621_n N_A_1236_138#_c_1186_n 0.0236154f $X=7.055 $Y=0.415
+ $X2=0 $Y2=0
cc_558 N_A_1034_392#_c_631_n N_A_1236_138#_c_1186_n 0.00224505f $X=7.14 $Y=0.415
+ $X2=0 $Y2=0
cc_559 N_A_1034_392#_c_623_n N_A_837_98#_M1034_g 0.00700429f $X=5.655 $Y=1.75
+ $X2=0 $Y2=0
cc_560 N_A_1034_392#_c_620_n N_A_837_98#_c_1314_n 0.00550212f $X=5.535 $Y=1.585
+ $X2=0 $Y2=0
cc_561 N_A_1034_392#_c_623_n N_A_837_98#_c_1314_n 0.00160082f $X=5.655 $Y=1.75
+ $X2=0 $Y2=0
cc_562 N_A_1034_392#_c_630_n N_A_837_98#_c_1314_n 0.00512277f $X=5.407 $Y=1.24
+ $X2=0 $Y2=0
cc_563 N_A_1034_392#_c_620_n N_A_837_98#_c_1315_n 0.0113002f $X=5.535 $Y=1.585
+ $X2=0 $Y2=0
cc_564 N_A_1034_392#_c_621_n N_A_837_98#_c_1315_n 0.00377769f $X=7.055 $Y=0.415
+ $X2=0 $Y2=0
cc_565 N_A_1034_392#_c_624_n N_A_837_98#_c_1315_n 0.00129942f $X=6.065 $Y=1.75
+ $X2=0 $Y2=0
cc_566 N_A_1034_392#_c_630_n N_A_837_98#_c_1315_n 0.0030377f $X=5.407 $Y=1.24
+ $X2=0 $Y2=0
cc_567 N_A_1034_392#_c_635_n N_A_837_98#_c_1316_n 0.0108355f $X=6.135 $Y=2.15
+ $X2=0 $Y2=0
cc_568 N_A_1034_392#_c_636_n N_A_837_98#_c_1316_n 0.0129473f $X=6.135 $Y=2.24
+ $X2=0 $Y2=0
cc_569 N_A_1034_392#_c_620_n N_A_837_98#_c_1316_n 0.00115334f $X=5.535 $Y=1.585
+ $X2=0 $Y2=0
cc_570 N_A_1034_392#_c_623_n N_A_837_98#_c_1316_n 0.0209904f $X=5.655 $Y=1.75
+ $X2=0 $Y2=0
cc_571 N_A_1034_392#_c_624_n N_A_837_98#_c_1316_n 0.00625338f $X=6.065 $Y=1.75
+ $X2=0 $Y2=0
cc_572 N_A_1034_392#_c_634_n N_A_837_98#_c_1316_n 0.021378f $X=6.065 $Y=1.66
+ $X2=0 $Y2=0
cc_573 N_A_1034_392#_c_636_n N_A_837_98#_c_1329_n 0.0103438f $X=6.135 $Y=2.24
+ $X2=0 $Y2=0
cc_574 N_A_1034_392#_c_621_n N_A_837_98#_c_1317_n 0.00133044f $X=7.055 $Y=0.415
+ $X2=0 $Y2=0
cc_575 N_A_1034_392#_c_624_n N_A_837_98#_c_1317_n 0.00334396f $X=6.065 $Y=1.75
+ $X2=0 $Y2=0
cc_576 N_A_1034_392#_c_634_n N_A_837_98#_c_1317_n 0.0143634f $X=6.065 $Y=1.66
+ $X2=0 $Y2=0
cc_577 N_A_1034_392#_M1041_g N_A_837_98#_c_1318_n 0.0184816f $X=6.535 $Y=0.9
+ $X2=0 $Y2=0
cc_578 N_A_1034_392#_c_619_n N_A_837_98#_c_1318_n 0.0041298f $X=5.37 $Y=0.745
+ $X2=0 $Y2=0
cc_579 N_A_1034_392#_c_621_n N_A_837_98#_c_1318_n 0.00357604f $X=7.055 $Y=0.415
+ $X2=0 $Y2=0
cc_580 N_A_1034_392#_c_636_n N_A_837_98#_c_1331_n 0.0024093f $X=6.135 $Y=2.24
+ $X2=0 $Y2=0
cc_581 N_A_1034_392#_c_636_n N_A_837_98#_c_1333_n 0.0137651f $X=6.135 $Y=2.24
+ $X2=0 $Y2=0
cc_582 N_A_1034_392#_c_614_n N_A_837_98#_c_1333_n 0.00158155f $X=6.46 $Y=1.66
+ $X2=0 $Y2=0
cc_583 N_A_1034_392#_c_638_n N_A_837_98#_c_1335_n 0.00689629f $X=9.835 $Y=2.465
+ $X2=0 $Y2=0
cc_584 N_A_1034_392#_c_638_n N_A_837_98#_M1042_g 0.0151225f $X=9.835 $Y=2.465
+ $X2=0 $Y2=0
cc_585 N_A_1034_392#_c_629_n N_A_837_98#_M1042_g 0.00774077f $X=9.33 $Y=2.065
+ $X2=0 $Y2=0
cc_586 N_A_1034_392#_c_665_p N_A_837_98#_M1042_g 0.00196389f $X=9.415 $Y=2.222
+ $X2=0 $Y2=0
cc_587 N_A_1034_392#_c_638_n N_A_837_98#_c_1319_n 0.00483103f $X=9.835 $Y=2.465
+ $X2=0 $Y2=0
cc_588 N_A_1034_392#_c_629_n N_A_837_98#_c_1319_n 0.0123734f $X=9.33 $Y=2.065
+ $X2=0 $Y2=0
cc_589 N_A_1034_392#_c_642_n N_A_837_98#_c_1319_n 0.00422095f $X=9.79 $Y=2.215
+ $X2=0 $Y2=0
cc_590 N_A_1034_392#_c_632_n N_A_837_98#_c_1319_n 0.00922521f $X=9.25 $Y=1.07
+ $X2=0 $Y2=0
cc_591 N_A_1034_392#_c_617_n N_A_837_98#_c_1320_n 0.00922521f $X=9.085 $Y=1.16
+ $X2=0 $Y2=0
cc_592 N_A_1034_392#_c_633_n N_A_837_98#_c_1320_n 0.00132052f $X=9.33 $Y=1.07
+ $X2=0 $Y2=0
cc_593 N_A_1034_392#_c_626_n N_A_837_98#_M1027_g 0.0039082f $X=8.825 $Y=0.34
+ $X2=0 $Y2=0
cc_594 N_A_1034_392#_c_628_n N_A_837_98#_M1027_g 0.00172497f $X=8.91 $Y=0.905
+ $X2=0 $Y2=0
cc_595 N_A_1034_392#_c_629_n N_A_837_98#_M1027_g 0.00175577f $X=9.33 $Y=2.065
+ $X2=0 $Y2=0
cc_596 N_A_1034_392#_c_632_n N_A_837_98#_M1027_g 0.0213739f $X=9.25 $Y=1.07
+ $X2=0 $Y2=0
cc_597 N_A_1034_392#_c_633_n N_A_837_98#_M1027_g 3.81838e-19 $X=9.33 $Y=1.07
+ $X2=0 $Y2=0
cc_598 N_A_1034_392#_c_630_n N_A_837_98#_c_1351_n 0.0116128f $X=5.407 $Y=1.24
+ $X2=0 $Y2=0
cc_599 N_A_1034_392#_c_620_n N_A_837_98#_c_1322_n 0.005941f $X=5.535 $Y=1.585
+ $X2=0 $Y2=0
cc_600 N_A_1034_392#_c_630_n N_A_837_98#_c_1322_n 0.00923218f $X=5.407 $Y=1.24
+ $X2=0 $Y2=0
cc_601 N_A_1034_392#_c_623_n N_A_837_98#_c_1342_n 0.00278431f $X=5.655 $Y=1.75
+ $X2=0 $Y2=0
cc_602 N_A_1034_392#_c_620_n N_A_837_98#_c_1324_n 0.0129947f $X=5.535 $Y=1.585
+ $X2=0 $Y2=0
cc_603 N_A_1034_392#_c_623_n N_A_837_98#_c_1324_n 0.0350942f $X=5.655 $Y=1.75
+ $X2=0 $Y2=0
cc_604 N_A_1034_392#_c_630_n N_A_837_98#_c_1324_n 0.00449451f $X=5.407 $Y=1.24
+ $X2=0 $Y2=0
cc_605 N_A_1034_392#_c_623_n N_A_837_98#_c_1325_n 0.00427453f $X=5.655 $Y=1.75
+ $X2=0 $Y2=0
cc_606 N_A_1034_392#_c_619_n N_A_837_98#_c_1326_n 0.00772518f $X=5.37 $Y=0.745
+ $X2=0 $Y2=0
cc_607 N_A_1034_392#_c_620_n N_A_837_98#_c_1326_n 0.00129629f $X=5.535 $Y=1.585
+ $X2=0 $Y2=0
cc_608 N_A_1034_392#_c_622_n N_A_837_98#_c_1326_n 0.00126334f $X=5.62 $Y=0.415
+ $X2=0 $Y2=0
cc_609 N_A_1034_392#_c_630_n N_A_837_98#_c_1326_n 0.00474804f $X=5.407 $Y=1.24
+ $X2=0 $Y2=0
cc_610 N_A_1034_392#_c_638_n N_A_2003_48#_c_1520_n 0.0213667f $X=9.835 $Y=2.465
+ $X2=0 $Y2=0
cc_611 N_A_1034_392#_c_642_n N_A_2003_48#_c_1520_n 3.86848e-19 $X=9.79 $Y=2.215
+ $X2=0 $Y2=0
cc_612 N_A_1034_392#_c_638_n N_A_2003_48#_c_1529_n 0.0337241f $X=9.835 $Y=2.465
+ $X2=0 $Y2=0
cc_613 N_A_1034_392#_c_626_n N_A_1745_74#_M1003_d 0.00191611f $X=8.825 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_614 N_A_1034_392#_c_628_n N_A_1745_74#_M1003_d 0.0113939f $X=8.91 $Y=0.905
+ $X2=-0.19 $Y2=-0.245
cc_615 N_A_1034_392#_c_633_n N_A_1745_74#_M1003_d 0.00132295f $X=9.33 $Y=1.07
+ $X2=-0.19 $Y2=-0.245
cc_616 N_A_1034_392#_c_629_n N_A_1745_74#_M1042_d 0.00800505f $X=9.33 $Y=2.065
+ $X2=0 $Y2=0
cc_617 N_A_1034_392#_c_665_p N_A_1745_74#_M1042_d 0.00493868f $X=9.415 $Y=2.222
+ $X2=0 $Y2=0
cc_618 N_A_1034_392#_c_642_n N_A_1745_74#_M1042_d 0.0018712f $X=9.79 $Y=2.215
+ $X2=0 $Y2=0
cc_619 N_A_1034_392#_c_616_n N_A_1745_74#_c_1641_n 6.35408e-19 $X=8.65 $Y=1.085
+ $X2=0 $Y2=0
cc_620 N_A_1034_392#_c_626_n N_A_1745_74#_c_1641_n 0.00169523f $X=8.825 $Y=0.34
+ $X2=0 $Y2=0
cc_621 N_A_1034_392#_c_628_n N_A_1745_74#_c_1641_n 0.0248143f $X=8.91 $Y=0.905
+ $X2=0 $Y2=0
cc_622 N_A_1034_392#_c_632_n N_A_1745_74#_c_1641_n 0.00569557f $X=9.25 $Y=1.07
+ $X2=0 $Y2=0
cc_623 N_A_1034_392#_c_633_n N_A_1745_74#_c_1641_n 0.0194065f $X=9.33 $Y=1.07
+ $X2=0 $Y2=0
cc_624 N_A_1034_392#_c_638_n N_A_1745_74#_c_1630_n 0.0210277f $X=9.835 $Y=2.465
+ $X2=0 $Y2=0
cc_625 N_A_1034_392#_c_665_p N_A_1745_74#_c_1630_n 0.0118084f $X=9.415 $Y=2.222
+ $X2=0 $Y2=0
cc_626 N_A_1034_392#_c_642_n N_A_1745_74#_c_1630_n 0.0365613f $X=9.79 $Y=2.215
+ $X2=0 $Y2=0
cc_627 N_A_1034_392#_c_628_n N_A_1745_74#_c_1617_n 0.00376918f $X=8.91 $Y=0.905
+ $X2=0 $Y2=0
cc_628 N_A_1034_392#_c_629_n N_A_1745_74#_c_1618_n 0.0357282f $X=9.33 $Y=2.065
+ $X2=0 $Y2=0
cc_629 N_A_1034_392#_c_632_n N_A_1745_74#_c_1618_n 5.18898e-19 $X=9.25 $Y=1.07
+ $X2=0 $Y2=0
cc_630 N_A_1034_392#_c_633_n N_A_1745_74#_c_1618_n 0.014106f $X=9.33 $Y=1.07
+ $X2=0 $Y2=0
cc_631 N_A_1034_392#_c_638_n N_A_1745_74#_c_1632_n 0.00349139f $X=9.835 $Y=2.465
+ $X2=0 $Y2=0
cc_632 N_A_1034_392#_c_642_n N_A_1745_74#_c_1632_n 0.0123723f $X=9.79 $Y=2.215
+ $X2=0 $Y2=0
cc_633 N_A_1034_392#_c_638_n N_A_1745_74#_c_1633_n 9.40099e-19 $X=9.835 $Y=2.465
+ $X2=0 $Y2=0
cc_634 N_A_1034_392#_c_629_n N_A_1745_74#_c_1633_n 0.0141964f $X=9.33 $Y=2.065
+ $X2=0 $Y2=0
cc_635 N_A_1034_392#_c_642_n N_A_1745_74#_c_1633_n 0.0119213f $X=9.79 $Y=2.215
+ $X2=0 $Y2=0
cc_636 N_A_1034_392#_c_638_n N_A_1745_74#_c_1634_n 0.00429238f $X=9.835 $Y=2.465
+ $X2=0 $Y2=0
cc_637 N_A_1034_392#_c_642_n N_A_1745_74#_c_1634_n 0.0246458f $X=9.79 $Y=2.215
+ $X2=0 $Y2=0
cc_638 N_A_1034_392#_c_628_n N_A_1745_74#_c_1620_n 7.09256e-19 $X=8.91 $Y=0.905
+ $X2=0 $Y2=0
cc_639 N_A_1034_392#_c_632_n N_A_1745_74#_c_1620_n 5.62433e-19 $X=9.25 $Y=1.07
+ $X2=0 $Y2=0
cc_640 N_A_1034_392#_c_633_n N_A_1745_74#_c_1620_n 0.0131492f $X=9.33 $Y=1.07
+ $X2=0 $Y2=0
cc_641 N_A_1034_392#_c_638_n N_VPWR_c_1904_n 0.00304676f $X=9.835 $Y=2.465 $X2=0
+ $Y2=0
cc_642 N_A_1034_392#_c_636_n N_VPWR_c_1889_n 9.39239e-19 $X=6.135 $Y=2.24 $X2=0
+ $Y2=0
cc_643 N_A_1034_392#_c_638_n N_VPWR_c_1889_n 0.00375679f $X=9.835 $Y=2.465 $X2=0
+ $Y2=0
cc_644 N_A_1034_392#_M1034_d N_A_415_81#_c_2091_n 0.00710909f $X=5.17 $Y=1.96
+ $X2=0 $Y2=0
cc_645 N_A_1034_392#_c_623_n N_A_415_81#_c_2091_n 0.0323397f $X=5.655 $Y=1.75
+ $X2=0 $Y2=0
cc_646 N_A_1034_392#_c_624_n N_A_415_81#_c_2091_n 0.00139329f $X=6.065 $Y=1.75
+ $X2=0 $Y2=0
cc_647 N_A_1034_392#_M1041_g N_A_415_81#_c_2086_n 2.59435e-19 $X=6.535 $Y=0.9
+ $X2=0 $Y2=0
cc_648 N_A_1034_392#_c_619_n N_A_415_81#_c_2086_n 0.0457818f $X=5.37 $Y=0.745
+ $X2=0 $Y2=0
cc_649 N_A_1034_392#_c_621_n N_A_415_81#_c_2086_n 0.0158801f $X=7.055 $Y=0.415
+ $X2=0 $Y2=0
cc_650 N_A_1034_392#_c_636_n N_A_415_81#_c_2092_n 0.00777844f $X=6.135 $Y=2.24
+ $X2=0 $Y2=0
cc_651 N_A_1034_392#_c_624_n N_A_415_81#_c_2092_n 0.00139775f $X=6.065 $Y=1.75
+ $X2=0 $Y2=0
cc_652 N_A_1034_392#_M1041_g N_A_415_81#_c_2087_n 0.00656958f $X=6.535 $Y=0.9
+ $X2=0 $Y2=0
cc_653 N_A_1034_392#_c_624_n N_A_415_81#_c_2087_n 0.0156466f $X=6.065 $Y=1.75
+ $X2=0 $Y2=0
cc_654 N_A_1034_392#_c_634_n N_A_415_81#_c_2087_n 0.00606607f $X=6.065 $Y=1.66
+ $X2=0 $Y2=0
cc_655 N_A_1034_392#_c_620_n N_A_415_81#_c_2088_n 0.0133096f $X=5.535 $Y=1.585
+ $X2=0 $Y2=0
cc_656 N_A_1034_392#_c_624_n N_A_415_81#_c_2088_n 0.0167772f $X=6.065 $Y=1.75
+ $X2=0 $Y2=0
cc_657 N_A_1034_392#_c_634_n N_A_415_81#_c_2088_n 5.99815e-19 $X=6.065 $Y=1.66
+ $X2=0 $Y2=0
cc_658 N_A_1034_392#_c_635_n N_A_415_81#_c_2093_n 0.00332822f $X=6.135 $Y=2.15
+ $X2=0 $Y2=0
cc_659 N_A_1034_392#_c_636_n N_A_415_81#_c_2093_n 0.00876113f $X=6.135 $Y=2.24
+ $X2=0 $Y2=0
cc_660 N_A_1034_392#_c_614_n N_A_415_81#_c_2093_n 0.00252722f $X=6.46 $Y=1.66
+ $X2=0 $Y2=0
cc_661 N_A_1034_392#_c_624_n N_A_415_81#_c_2093_n 0.00797914f $X=6.065 $Y=1.75
+ $X2=0 $Y2=0
cc_662 N_A_1034_392#_c_635_n N_A_415_81#_c_2094_n 0.00108341f $X=6.135 $Y=2.15
+ $X2=0 $Y2=0
cc_663 N_A_1034_392#_c_636_n N_A_415_81#_c_2094_n 0.00170504f $X=6.135 $Y=2.24
+ $X2=0 $Y2=0
cc_664 N_A_1034_392#_c_623_n N_A_415_81#_c_2094_n 0.0132392f $X=5.655 $Y=1.75
+ $X2=0 $Y2=0
cc_665 N_A_1034_392#_c_624_n N_A_415_81#_c_2094_n 0.0167298f $X=6.065 $Y=1.75
+ $X2=0 $Y2=0
cc_666 N_A_1034_392#_c_634_n N_A_415_81#_c_2094_n 0.00323194f $X=6.065 $Y=1.66
+ $X2=0 $Y2=0
cc_667 N_A_1034_392#_c_635_n N_A_415_81#_c_2089_n 0.00366894f $X=6.135 $Y=2.15
+ $X2=0 $Y2=0
cc_668 N_A_1034_392#_c_614_n N_A_415_81#_c_2089_n 0.0107867f $X=6.46 $Y=1.66
+ $X2=0 $Y2=0
cc_669 N_A_1034_392#_M1041_g N_A_415_81#_c_2089_n 0.00503924f $X=6.535 $Y=0.9
+ $X2=0 $Y2=0
cc_670 N_A_1034_392#_c_624_n N_A_415_81#_c_2089_n 0.0256546f $X=6.065 $Y=1.75
+ $X2=0 $Y2=0
cc_671 N_A_1034_392#_c_634_n N_A_415_81#_c_2089_n 0.00187233f $X=6.065 $Y=1.66
+ $X2=0 $Y2=0
cc_672 N_A_1034_392#_c_625_n N_VGND_M1024_d 0.0162233f $X=7.93 $Y=0.665 $X2=0
+ $Y2=0
cc_673 N_A_1034_392#_c_678_p N_VGND_M1024_d 0.00247125f $X=8.015 $Y=0.58 $X2=0
+ $Y2=0
cc_674 N_A_1034_392#_c_627_n N_VGND_M1024_d 6.8704e-19 $X=8.1 $Y=0.34 $X2=0
+ $Y2=0
cc_675 N_A_1034_392#_c_619_n N_VGND_c_2314_n 0.0135513f $X=5.37 $Y=0.745 $X2=0
+ $Y2=0
cc_676 N_A_1034_392#_c_622_n N_VGND_c_2314_n 0.0148789f $X=5.62 $Y=0.415 $X2=0
+ $Y2=0
cc_677 N_A_1034_392#_c_621_n N_VGND_c_2315_n 0.0628116f $X=7.055 $Y=0.415 $X2=0
+ $Y2=0
cc_678 N_A_1034_392#_c_622_n N_VGND_c_2315_n 0.0196297f $X=5.62 $Y=0.415 $X2=0
+ $Y2=0
cc_679 N_A_1034_392#_c_625_n N_VGND_c_2315_n 0.00392706f $X=7.93 $Y=0.665 $X2=0
+ $Y2=0
cc_680 N_A_1034_392#_c_631_n N_VGND_c_2315_n 0.00786741f $X=7.14 $Y=0.415 $X2=0
+ $Y2=0
cc_681 N_A_1034_392#_c_616_n N_VGND_c_2324_n 0.00278271f $X=8.65 $Y=1.085 $X2=0
+ $Y2=0
cc_682 N_A_1034_392#_c_625_n N_VGND_c_2324_n 0.00335833f $X=7.93 $Y=0.665 $X2=0
+ $Y2=0
cc_683 N_A_1034_392#_c_626_n N_VGND_c_2324_n 0.0579202f $X=8.825 $Y=0.34 $X2=0
+ $Y2=0
cc_684 N_A_1034_392#_c_627_n N_VGND_c_2324_n 0.0118998f $X=8.1 $Y=0.34 $X2=0
+ $Y2=0
cc_685 N_A_1034_392#_c_625_n N_VGND_c_2329_n 0.0246013f $X=7.93 $Y=0.665 $X2=0
+ $Y2=0
cc_686 N_A_1034_392#_c_627_n N_VGND_c_2329_n 0.0135791f $X=8.1 $Y=0.34 $X2=0
+ $Y2=0
cc_687 N_A_1034_392#_c_631_n N_VGND_c_2329_n 0.00555628f $X=7.14 $Y=0.415 $X2=0
+ $Y2=0
cc_688 N_A_1034_392#_c_616_n N_VGND_c_2334_n 0.00358928f $X=8.65 $Y=1.085 $X2=0
+ $Y2=0
cc_689 N_A_1034_392#_c_621_n N_VGND_c_2334_n 0.0456845f $X=7.055 $Y=0.415 $X2=0
+ $Y2=0
cc_690 N_A_1034_392#_c_622_n N_VGND_c_2334_n 0.0135126f $X=5.62 $Y=0.415 $X2=0
+ $Y2=0
cc_691 N_A_1034_392#_c_625_n N_VGND_c_2334_n 0.012145f $X=7.93 $Y=0.665 $X2=0
+ $Y2=0
cc_692 N_A_1034_392#_c_626_n N_VGND_c_2334_n 0.0324872f $X=8.825 $Y=0.34 $X2=0
+ $Y2=0
cc_693 N_A_1034_392#_c_627_n N_VGND_c_2334_n 0.00655543f $X=8.1 $Y=0.34 $X2=0
+ $Y2=0
cc_694 N_A_1034_392#_c_631_n N_VGND_c_2334_n 0.0055105f $X=7.14 $Y=0.415 $X2=0
+ $Y2=0
cc_695 N_A_1034_392#_c_631_n A_1397_138# 0.00203667f $X=7.14 $Y=0.415 $X2=-0.19
+ $Y2=-0.245
cc_696 N_A_1367_112#_M1044_g N_RESET_B_c_955_n 0.00526413f $X=6.91 $Y=0.9 $X2=0
+ $Y2=0
cc_697 N_A_1367_112#_M1044_g N_RESET_B_M1024_g 0.0394201f $X=6.91 $Y=0.9 $X2=0
+ $Y2=0
cc_698 N_A_1367_112#_c_844_n N_RESET_B_M1024_g 0.00515512f $X=7.19 $Y=1.78 $X2=0
+ $Y2=0
cc_699 N_A_1367_112#_c_863_n N_RESET_B_M1024_g 0.00422682f $X=7.325 $Y=1.005
+ $X2=0 $Y2=0
cc_700 N_A_1367_112#_c_874_n N_RESET_B_M1024_g 0.0067801f $X=8.27 $Y=0.842 $X2=0
+ $Y2=0
cc_701 N_A_1367_112#_c_874_n N_RESET_B_c_958_n 0.00975109f $X=8.27 $Y=0.842
+ $X2=0 $Y2=0
cc_702 N_A_1367_112#_c_844_n N_RESET_B_c_959_n 0.00753567f $X=7.19 $Y=1.78 $X2=0
+ $Y2=0
cc_703 N_A_1367_112#_c_845_n N_RESET_B_c_959_n 0.00620241f $X=7.19 $Y=1.78 $X2=0
+ $Y2=0
cc_704 N_A_1367_112#_c_849_n N_RESET_B_c_965_n 0.0123322f $X=7.025 $Y=2.24 $X2=0
+ $Y2=0
cc_705 N_A_1367_112#_M1044_g N_RESET_B_c_960_n 0.00326496f $X=6.91 $Y=0.9 $X2=0
+ $Y2=0
cc_706 N_A_1367_112#_c_844_n N_RESET_B_c_960_n 0.00113842f $X=7.19 $Y=1.78 $X2=0
+ $Y2=0
cc_707 N_A_1367_112#_c_845_n N_RESET_B_c_960_n 0.0110407f $X=7.19 $Y=1.78 $X2=0
+ $Y2=0
cc_708 N_A_1367_112#_c_848_n N_RESET_B_c_970_n 0.0105234f $X=7.025 $Y=2.15 $X2=0
+ $Y2=0
cc_709 N_A_1367_112#_c_844_n N_RESET_B_c_970_n 0.009228f $X=7.19 $Y=1.78 $X2=0
+ $Y2=0
cc_710 N_A_1367_112#_c_845_n N_RESET_B_c_970_n 0.00237054f $X=7.19 $Y=1.78 $X2=0
+ $Y2=0
cc_711 N_A_1367_112#_c_847_n N_RESET_B_c_972_n 0.00727956f $X=8.9 $Y=1.575 $X2=0
+ $Y2=0
cc_712 N_A_1367_112#_c_853_n N_RESET_B_c_972_n 0.030687f $X=8.9 $Y=1.88 $X2=0
+ $Y2=0
cc_713 N_A_1367_112#_c_848_n N_RESET_B_c_978_n 0.00683215f $X=7.025 $Y=2.15
+ $X2=0 $Y2=0
cc_714 N_A_1367_112#_c_845_n N_RESET_B_c_978_n 0.00760267f $X=7.19 $Y=1.78 $X2=0
+ $Y2=0
cc_715 N_A_1367_112#_c_846_n N_A_1236_138#_M1019_g 0.00313626f $X=8.57 $Y=1.405
+ $X2=0 $Y2=0
cc_716 N_A_1367_112#_c_874_n N_A_1236_138#_M1019_g 0.0131882f $X=8.27 $Y=0.842
+ $X2=0 $Y2=0
cc_717 N_A_1367_112#_c_846_n N_A_1236_138#_c_1180_n 0.00107505f $X=8.57 $Y=1.405
+ $X2=0 $Y2=0
cc_718 N_A_1367_112#_c_847_n N_A_1236_138#_c_1180_n 0.0131822f $X=8.9 $Y=1.575
+ $X2=0 $Y2=0
cc_719 N_A_1367_112#_c_853_n N_A_1236_138#_c_1180_n 0.00530481f $X=8.9 $Y=1.88
+ $X2=0 $Y2=0
cc_720 N_A_1367_112#_c_876_n N_A_1236_138#_c_1180_n 0.00405015f $X=8.57 $Y=0.842
+ $X2=0 $Y2=0
cc_721 N_A_1367_112#_c_853_n N_A_1236_138#_c_1188_n 0.0151257f $X=8.9 $Y=1.88
+ $X2=0 $Y2=0
cc_722 N_A_1367_112#_M1044_g N_A_1236_138#_c_1202_n 0.00463522f $X=6.91 $Y=0.9
+ $X2=0 $Y2=0
cc_723 N_A_1367_112#_c_863_n N_A_1236_138#_c_1202_n 0.0130756f $X=7.325 $Y=1.005
+ $X2=0 $Y2=0
cc_724 N_A_1367_112#_M1044_g N_A_1236_138#_c_1181_n 0.00936736f $X=6.91 $Y=0.9
+ $X2=0 $Y2=0
cc_725 N_A_1367_112#_c_848_n N_A_1236_138#_c_1181_n 0.0045184f $X=7.025 $Y=2.15
+ $X2=0 $Y2=0
cc_726 N_A_1367_112#_c_849_n N_A_1236_138#_c_1181_n 9.21498e-19 $X=7.025 $Y=2.24
+ $X2=0 $Y2=0
cc_727 N_A_1367_112#_c_844_n N_A_1236_138#_c_1181_n 0.062072f $X=7.19 $Y=1.78
+ $X2=0 $Y2=0
cc_728 N_A_1367_112#_c_845_n N_A_1236_138#_c_1181_n 0.0104152f $X=7.19 $Y=1.78
+ $X2=0 $Y2=0
cc_729 N_A_1367_112#_c_863_n N_A_1236_138#_c_1181_n 0.00114989f $X=7.325
+ $Y=1.005 $X2=0 $Y2=0
cc_730 N_A_1367_112#_c_849_n N_A_1236_138#_c_1225_n 0.0109144f $X=7.025 $Y=2.24
+ $X2=0 $Y2=0
cc_731 N_A_1367_112#_c_844_n N_A_1236_138#_c_1225_n 0.00526266f $X=7.19 $Y=1.78
+ $X2=0 $Y2=0
cc_732 N_A_1367_112#_c_845_n N_A_1236_138#_c_1225_n 0.00311782f $X=7.19 $Y=1.78
+ $X2=0 $Y2=0
cc_733 N_A_1367_112#_c_848_n N_A_1236_138#_c_1182_n 0.00204704f $X=7.025 $Y=2.15
+ $X2=0 $Y2=0
cc_734 N_A_1367_112#_c_849_n N_A_1236_138#_c_1182_n 0.00139157f $X=7.025 $Y=2.24
+ $X2=0 $Y2=0
cc_735 N_A_1367_112#_c_844_n N_A_1236_138#_c_1182_n 0.0274325f $X=7.19 $Y=1.78
+ $X2=0 $Y2=0
cc_736 N_A_1367_112#_c_845_n N_A_1236_138#_c_1182_n 0.00208168f $X=7.19 $Y=1.78
+ $X2=0 $Y2=0
cc_737 N_A_1367_112#_c_844_n N_A_1236_138#_c_1183_n 0.0268297f $X=7.19 $Y=1.78
+ $X2=0 $Y2=0
cc_738 N_A_1367_112#_c_874_n N_A_1236_138#_c_1183_n 0.0133196f $X=8.27 $Y=0.842
+ $X2=0 $Y2=0
cc_739 N_A_1367_112#_c_846_n N_A_1236_138#_c_1184_n 0.0115079f $X=8.57 $Y=1.405
+ $X2=0 $Y2=0
cc_740 N_A_1367_112#_c_847_n N_A_1236_138#_c_1184_n 0.0142233f $X=8.9 $Y=1.575
+ $X2=0 $Y2=0
cc_741 N_A_1367_112#_c_874_n N_A_1236_138#_c_1184_n 0.0443118f $X=8.27 $Y=0.842
+ $X2=0 $Y2=0
cc_742 N_A_1367_112#_c_846_n N_A_1236_138#_c_1185_n 0.00161618f $X=8.57 $Y=1.405
+ $X2=0 $Y2=0
cc_743 N_A_1367_112#_c_847_n N_A_1236_138#_c_1185_n 3.02987e-19 $X=8.9 $Y=1.575
+ $X2=0 $Y2=0
cc_744 N_A_1367_112#_c_874_n N_A_1236_138#_c_1185_n 0.00252719f $X=8.27 $Y=0.842
+ $X2=0 $Y2=0
cc_745 N_A_1367_112#_c_876_n N_A_1236_138#_c_1185_n 0.00137742f $X=8.57 $Y=0.842
+ $X2=0 $Y2=0
cc_746 N_A_1367_112#_M1044_g N_A_1236_138#_c_1186_n 0.00105321f $X=6.91 $Y=0.9
+ $X2=0 $Y2=0
cc_747 N_A_1367_112#_c_849_n N_A_1236_138#_c_1193_n 0.0060004f $X=7.025 $Y=2.24
+ $X2=0 $Y2=0
cc_748 N_A_1367_112#_c_849_n N_A_837_98#_c_1331_n 0.00323347f $X=7.025 $Y=2.24
+ $X2=0 $Y2=0
cc_749 N_A_1367_112#_c_849_n N_A_837_98#_c_1333_n 0.0307207f $X=7.025 $Y=2.24
+ $X2=0 $Y2=0
cc_750 N_A_1367_112#_c_849_n N_A_837_98#_c_1334_n 0.0100502f $X=7.025 $Y=2.24
+ $X2=0 $Y2=0
cc_751 N_A_1367_112#_c_853_n N_A_837_98#_c_1334_n 0.00400096f $X=8.9 $Y=1.88
+ $X2=0 $Y2=0
cc_752 N_A_1367_112#_c_853_n N_A_837_98#_c_1335_n 5.08057e-19 $X=8.9 $Y=1.88
+ $X2=0 $Y2=0
cc_753 N_A_1367_112#_c_853_n N_A_837_98#_M1042_g 0.014001f $X=8.9 $Y=1.88 $X2=0
+ $Y2=0
cc_754 N_A_1367_112#_c_847_n N_A_837_98#_c_1320_n 0.0021457f $X=8.9 $Y=1.575
+ $X2=0 $Y2=0
cc_755 N_A_1367_112#_c_853_n N_A_837_98#_c_1320_n 0.00289869f $X=8.9 $Y=1.88
+ $X2=0 $Y2=0
cc_756 N_A_1367_112#_c_853_n N_A_1745_74#_c_1630_n 0.0146147f $X=8.9 $Y=1.88
+ $X2=0 $Y2=0
cc_757 N_A_1367_112#_c_849_n N_VPWR_c_1892_n 0.00433246f $X=7.025 $Y=2.24 $X2=0
+ $Y2=0
cc_758 N_A_1367_112#_c_847_n N_VPWR_c_1894_n 0.00369686f $X=8.9 $Y=1.575 $X2=0
+ $Y2=0
cc_759 N_A_1367_112#_c_853_n N_VPWR_c_1894_n 0.064586f $X=8.9 $Y=1.88 $X2=0
+ $Y2=0
cc_760 N_A_1367_112#_c_876_n N_VPWR_c_1894_n 0.00374786f $X=8.57 $Y=0.842 $X2=0
+ $Y2=0
cc_761 N_A_1367_112#_c_853_n N_VPWR_c_1904_n 0.00748753f $X=8.9 $Y=1.88 $X2=0
+ $Y2=0
cc_762 N_A_1367_112#_c_849_n N_VPWR_c_1889_n 9.39239e-19 $X=7.025 $Y=2.24 $X2=0
+ $Y2=0
cc_763 N_A_1367_112#_c_853_n N_VPWR_c_1889_n 0.00904755f $X=8.9 $Y=1.88 $X2=0
+ $Y2=0
cc_764 N_A_1367_112#_M1044_g N_A_415_81#_c_2089_n 2.91755e-19 $X=6.91 $Y=0.9
+ $X2=0 $Y2=0
cc_765 N_A_1367_112#_c_845_n N_A_415_81#_c_2089_n 6.15582e-19 $X=7.19 $Y=1.78
+ $X2=0 $Y2=0
cc_766 N_A_1367_112#_c_874_n N_VGND_M1024_d 0.0155117f $X=8.27 $Y=0.842 $X2=0
+ $Y2=0
cc_767 N_A_1367_112#_c_863_n A_1397_138# 0.00260878f $X=7.325 $Y=1.005 $X2=-0.19
+ $Y2=-0.245
cc_768 N_RESET_B_c_958_n N_A_1236_138#_M1019_g 0.00269339f $X=7.595 $Y=1.26
+ $X2=0 $Y2=0
cc_769 N_RESET_B_c_972_n N_A_1236_138#_c_1180_n 3.01246e-19 $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_770 N_RESET_B_c_972_n N_A_1236_138#_c_1188_n 0.00699288f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_771 N_RESET_B_c_970_n N_A_1236_138#_c_1189_n 0.00819966f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_772 N_RESET_B_M1024_g N_A_1236_138#_c_1202_n 2.03434e-19 $X=7.3 $Y=0.9 $X2=0
+ $Y2=0
cc_773 N_RESET_B_M1024_g N_A_1236_138#_c_1181_n 2.11405e-19 $X=7.3 $Y=0.9 $X2=0
+ $Y2=0
cc_774 N_RESET_B_c_970_n N_A_1236_138#_c_1181_n 0.0241128f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_775 N_RESET_B_c_970_n N_A_1236_138#_c_1225_n 0.020887f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_776 N_RESET_B_c_965_n N_A_1236_138#_c_1182_n 0.0179696f $X=7.665 $Y=2.24
+ $X2=0 $Y2=0
cc_777 N_RESET_B_c_960_n N_A_1236_138#_c_1182_n 0.0117416f $X=7.67 $Y=1.82 $X2=0
+ $Y2=0
cc_778 N_RESET_B_c_970_n N_A_1236_138#_c_1182_n 0.0257004f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_779 N_RESET_B_c_973_n N_A_1236_138#_c_1182_n 0.0106292f $X=8.065 $Y=2.035
+ $X2=0 $Y2=0
cc_780 N_RESET_B_c_974_n N_A_1236_138#_c_1182_n 0.0363198f $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_781 N_RESET_B_c_978_n N_A_1236_138#_c_1182_n 0.020253f $X=7.67 $Y=2.03 $X2=0
+ $Y2=0
cc_782 N_RESET_B_c_958_n N_A_1236_138#_c_1183_n 0.00569114f $X=7.595 $Y=1.26
+ $X2=0 $Y2=0
cc_783 N_RESET_B_c_960_n N_A_1236_138#_c_1183_n 0.00438308f $X=7.67 $Y=1.82
+ $X2=0 $Y2=0
cc_784 N_RESET_B_c_958_n N_A_1236_138#_c_1184_n 0.00188178f $X=7.595 $Y=1.26
+ $X2=0 $Y2=0
cc_785 N_RESET_B_c_960_n N_A_1236_138#_c_1184_n 0.00586797f $X=7.67 $Y=1.82
+ $X2=0 $Y2=0
cc_786 N_RESET_B_c_970_n N_A_1236_138#_c_1184_n 0.00357593f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_787 N_RESET_B_c_972_n N_A_1236_138#_c_1184_n 0.00641796f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_788 N_RESET_B_c_973_n N_A_1236_138#_c_1184_n 0.00373314f $X=8.065 $Y=2.035
+ $X2=0 $Y2=0
cc_789 N_RESET_B_c_974_n N_A_1236_138#_c_1184_n 0.0158779f $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_790 N_RESET_B_c_978_n N_A_1236_138#_c_1184_n 0.00716371f $X=7.67 $Y=2.03
+ $X2=0 $Y2=0
cc_791 N_RESET_B_c_958_n N_A_1236_138#_c_1185_n 0.0194698f $X=7.595 $Y=1.26
+ $X2=0 $Y2=0
cc_792 N_RESET_B_c_972_n N_A_1236_138#_c_1185_n 0.00591166f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_793 N_RESET_B_c_974_n N_A_1236_138#_c_1185_n 6.12607e-19 $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_794 N_RESET_B_c_978_n N_A_1236_138#_c_1185_n 0.00918526f $X=7.67 $Y=2.03
+ $X2=0 $Y2=0
cc_795 N_RESET_B_c_970_n N_A_837_98#_M1030_s 0.00168963f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_796 N_RESET_B_c_970_n N_A_837_98#_M1034_g 0.00360859f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_797 N_RESET_B_c_970_n N_A_837_98#_c_1316_n 0.00172072f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_798 N_RESET_B_c_955_n N_A_837_98#_c_1318_n 0.00526413f $X=7.225 $Y=0.18 $X2=0
+ $Y2=0
cc_799 N_RESET_B_c_970_n N_A_837_98#_c_1333_n 0.00378573f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_800 N_RESET_B_c_965_n N_A_837_98#_c_1334_n 0.0100134f $X=7.665 $Y=2.24 $X2=0
+ $Y2=0
cc_801 N_RESET_B_c_972_n N_A_837_98#_M1042_g 0.0124871f $X=10.655 $Y=2.035 $X2=0
+ $Y2=0
cc_802 N_RESET_B_c_972_n N_A_837_98#_c_1319_n 0.00423021f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_803 N_RESET_B_c_970_n N_A_837_98#_c_1341_n 0.0131961f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_804 N_RESET_B_c_955_n N_A_837_98#_c_1351_n 0.0011436f $X=7.225 $Y=0.18 $X2=0
+ $Y2=0
cc_805 N_RESET_B_c_955_n N_A_837_98#_c_1323_n 0.00701575f $X=7.225 $Y=0.18 $X2=0
+ $Y2=0
cc_806 N_RESET_B_c_970_n N_A_837_98#_c_1342_n 0.0118682f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_807 N_RESET_B_c_971_n N_A_837_98#_c_1342_n 0.00275582f $X=4.225 $Y=2.035
+ $X2=0 $Y2=0
cc_808 N_RESET_B_c_976_n N_A_837_98#_c_1342_n 0.00285508f $X=3.605 $Y=2.037
+ $X2=0 $Y2=0
cc_809 N_RESET_B_c_977_n N_A_837_98#_c_1342_n 0.0238091f $X=3.95 $Y=1.995 $X2=0
+ $Y2=0
cc_810 N_RESET_B_c_970_n N_A_837_98#_c_1324_n 0.0164918f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_811 N_RESET_B_c_970_n N_A_837_98#_c_1325_n 0.00111147f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_812 N_RESET_B_c_955_n N_A_837_98#_c_1326_n 0.0102196f $X=7.225 $Y=0.18 $X2=0
+ $Y2=0
cc_813 N_RESET_B_M1038_g N_A_2003_48#_M1021_g 0.0216011f $X=10.63 $Y=0.58 $X2=0
+ $Y2=0
cc_814 N_RESET_B_c_968_n N_A_2003_48#_c_1520_n 0.00394367f $X=10.94 $Y=2.375
+ $X2=0 $Y2=0
cc_815 N_RESET_B_c_972_n N_A_2003_48#_c_1520_n 0.00331802f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_816 N_RESET_B_c_979_n N_A_2003_48#_c_1520_n 0.00106389f $X=10.75 $Y=1.985
+ $X2=0 $Y2=0
cc_817 N_RESET_B_c_980_n N_A_2003_48#_c_1520_n 0.029932f $X=10.94 $Y=1.985 $X2=0
+ $Y2=0
cc_818 N_RESET_B_c_969_n N_A_2003_48#_c_1529_n 0.0126655f $X=10.94 $Y=2.465
+ $X2=0 $Y2=0
cc_819 N_RESET_B_M1038_g N_A_2003_48#_c_1521_n 0.0128807f $X=10.63 $Y=0.58 $X2=0
+ $Y2=0
cc_820 N_RESET_B_c_972_n N_A_2003_48#_c_1521_n 0.00879069f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_821 RESET_B N_A_2003_48#_c_1521_n 0.00259932f $X=10.715 $Y=1.95 $X2=0 $Y2=0
cc_822 N_RESET_B_c_979_n N_A_2003_48#_c_1521_n 0.0152297f $X=10.75 $Y=1.985
+ $X2=0 $Y2=0
cc_823 N_RESET_B_c_980_n N_A_2003_48#_c_1521_n 0.00391331f $X=10.94 $Y=1.985
+ $X2=0 $Y2=0
cc_824 N_RESET_B_M1038_g N_A_2003_48#_c_1522_n 9.6789e-19 $X=10.63 $Y=0.58 $X2=0
+ $Y2=0
cc_825 N_RESET_B_M1038_g N_A_2003_48#_c_1524_n 0.00118187f $X=10.63 $Y=0.58
+ $X2=0 $Y2=0
cc_826 N_RESET_B_c_972_n N_A_2003_48#_c_1524_n 0.00250381f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_827 N_RESET_B_M1038_g N_A_2003_48#_c_1525_n 0.029932f $X=10.63 $Y=0.58 $X2=0
+ $Y2=0
cc_828 N_RESET_B_c_969_n N_A_2003_48#_c_1530_n 0.00739105f $X=10.94 $Y=2.465
+ $X2=0 $Y2=0
cc_829 N_RESET_B_M1038_g N_A_2003_48#_c_1526_n 0.00453304f $X=10.63 $Y=0.58
+ $X2=0 $Y2=0
cc_830 N_RESET_B_c_969_n N_A_2003_48#_c_1526_n 0.00121218f $X=10.94 $Y=2.465
+ $X2=0 $Y2=0
cc_831 RESET_B N_A_2003_48#_c_1526_n 0.00621393f $X=10.715 $Y=1.95 $X2=0 $Y2=0
cc_832 N_RESET_B_c_979_n N_A_2003_48#_c_1526_n 0.0154382f $X=10.75 $Y=1.985
+ $X2=0 $Y2=0
cc_833 N_RESET_B_c_980_n N_A_2003_48#_c_1526_n 0.0101596f $X=10.94 $Y=1.985
+ $X2=0 $Y2=0
cc_834 N_RESET_B_c_972_n N_A_1745_74#_M1042_d 0.00323029f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_835 N_RESET_B_M1038_g N_A_1745_74#_c_1608_n 0.0694909f $X=10.63 $Y=0.58 $X2=0
+ $Y2=0
cc_836 N_RESET_B_c_980_n N_A_1745_74#_c_1624_n 0.00857472f $X=10.94 $Y=1.985
+ $X2=0 $Y2=0
cc_837 N_RESET_B_c_968_n N_A_1745_74#_c_1625_n 0.00857472f $X=10.94 $Y=2.375
+ $X2=0 $Y2=0
cc_838 N_RESET_B_c_969_n N_A_1745_74#_c_1625_n 0.010499f $X=10.94 $Y=2.465 $X2=0
+ $Y2=0
cc_839 N_RESET_B_M1038_g N_A_1745_74#_c_1614_n 0.00550286f $X=10.63 $Y=0.58
+ $X2=0 $Y2=0
cc_840 N_RESET_B_c_972_n N_A_1745_74#_c_1630_n 0.00708586f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_841 N_RESET_B_M1038_g N_A_1745_74#_c_1619_n 0.0150978f $X=10.63 $Y=0.58 $X2=0
+ $Y2=0
cc_842 N_RESET_B_M1038_g N_A_1745_74#_c_1632_n 8.1654e-19 $X=10.63 $Y=0.58 $X2=0
+ $Y2=0
cc_843 N_RESET_B_c_972_n N_A_1745_74#_c_1632_n 0.0117357f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_844 N_RESET_B_c_979_n N_A_1745_74#_c_1632_n 0.00391217f $X=10.75 $Y=1.985
+ $X2=0 $Y2=0
cc_845 N_RESET_B_c_972_n N_A_1745_74#_c_1633_n 0.00499654f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_846 N_RESET_B_c_968_n N_A_1745_74#_c_1634_n 0.00158772f $X=10.94 $Y=2.375
+ $X2=0 $Y2=0
cc_847 N_RESET_B_c_969_n N_A_1745_74#_c_1634_n 2.73747e-19 $X=10.94 $Y=2.465
+ $X2=0 $Y2=0
cc_848 N_RESET_B_c_972_n N_A_1745_74#_c_1634_n 0.0200435f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_849 RESET_B N_A_1745_74#_c_1634_n 4.97327e-19 $X=10.715 $Y=1.95 $X2=0 $Y2=0
cc_850 N_RESET_B_c_979_n N_A_1745_74#_c_1634_n 0.00972451f $X=10.75 $Y=1.985
+ $X2=0 $Y2=0
cc_851 N_RESET_B_c_980_n N_A_1745_74#_c_1634_n 8.72425e-19 $X=10.94 $Y=1.985
+ $X2=0 $Y2=0
cc_852 N_RESET_B_M1038_g N_A_1745_74#_c_1621_n 0.00118187f $X=10.63 $Y=0.58
+ $X2=0 $Y2=0
cc_853 N_RESET_B_c_980_n N_A_1745_74#_c_1622_n 0.00231637f $X=10.94 $Y=1.985
+ $X2=0 $Y2=0
cc_854 N_RESET_B_c_970_n N_VPWR_M1030_d 0.00315295f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_855 N_RESET_B_c_972_n N_VPWR_M1031_s 0.00641842f $X=10.655 $Y=2.035 $X2=0
+ $Y2=0
cc_856 N_RESET_B_c_964_n N_VPWR_c_1890_n 0.00548967f $X=3.605 $Y=2.245 $X2=0
+ $Y2=0
cc_857 N_RESET_B_c_965_n N_VPWR_c_1892_n 0.00421039f $X=7.665 $Y=2.24 $X2=0
+ $Y2=0
cc_858 N_RESET_B_c_970_n N_VPWR_c_1892_n 7.46496e-19 $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_859 N_RESET_B_c_965_n N_VPWR_c_1894_n 0.00486917f $X=7.665 $Y=2.24 $X2=0
+ $Y2=0
cc_860 N_RESET_B_c_960_n N_VPWR_c_1894_n 0.00160044f $X=7.67 $Y=1.82 $X2=0 $Y2=0
cc_861 N_RESET_B_c_972_n N_VPWR_c_1894_n 0.0183166f $X=10.655 $Y=2.035 $X2=0
+ $Y2=0
cc_862 N_RESET_B_c_973_n N_VPWR_c_1894_n 5.40997e-19 $X=8.065 $Y=2.035 $X2=0
+ $Y2=0
cc_863 N_RESET_B_c_974_n N_VPWR_c_1894_n 0.0179605f $X=7.92 $Y=2.035 $X2=0 $Y2=0
cc_864 N_RESET_B_c_978_n N_VPWR_c_1894_n 0.00312179f $X=7.67 $Y=2.03 $X2=0 $Y2=0
cc_865 N_RESET_B_c_969_n N_VPWR_c_1895_n 0.00816134f $X=10.94 $Y=2.465 $X2=0
+ $Y2=0
cc_866 N_RESET_B_c_972_n N_VPWR_c_1895_n 0.00540169f $X=10.655 $Y=2.035 $X2=0
+ $Y2=0
cc_867 RESET_B N_VPWR_c_1895_n 0.00113612f $X=10.715 $Y=1.95 $X2=0 $Y2=0
cc_868 N_RESET_B_c_979_n N_VPWR_c_1895_n 0.00684931f $X=10.75 $Y=1.985 $X2=0
+ $Y2=0
cc_869 N_RESET_B_c_980_n N_VPWR_c_1895_n 0.00269311f $X=10.94 $Y=1.985 $X2=0
+ $Y2=0
cc_870 N_RESET_B_c_964_n N_VPWR_c_1902_n 0.00388952f $X=3.605 $Y=2.245 $X2=0
+ $Y2=0
cc_871 N_RESET_B_c_969_n N_VPWR_c_1909_n 0.00445602f $X=10.94 $Y=2.465 $X2=0
+ $Y2=0
cc_872 N_RESET_B_c_964_n N_VPWR_c_1889_n 0.00420469f $X=3.605 $Y=2.245 $X2=0
+ $Y2=0
cc_873 N_RESET_B_c_965_n N_VPWR_c_1889_n 9.39239e-19 $X=7.665 $Y=2.24 $X2=0
+ $Y2=0
cc_874 N_RESET_B_c_969_n N_VPWR_c_1889_n 0.0089746f $X=10.94 $Y=2.465 $X2=0
+ $Y2=0
cc_875 N_RESET_B_c_953_n N_A_415_81#_c_2084_n 0.00193822f $X=3.555 $Y=1.83 $X2=0
+ $Y2=0
cc_876 N_RESET_B_M1012_g N_A_415_81#_c_2084_n 0.00887388f $X=3.575 $Y=0.615
+ $X2=0 $Y2=0
cc_877 N_RESET_B_c_962_n N_A_415_81#_c_2084_n 0.00666445f $X=3.565 $Y=1.06 $X2=0
+ $Y2=0
cc_878 N_RESET_B_c_953_n N_A_415_81#_c_2085_n 0.0252779f $X=3.555 $Y=1.83 $X2=0
+ $Y2=0
cc_879 N_RESET_B_c_964_n N_A_415_81#_c_2085_n 0.00445911f $X=3.605 $Y=2.245
+ $X2=0 $Y2=0
cc_880 N_RESET_B_c_971_n N_A_415_81#_c_2085_n 0.00108729f $X=4.225 $Y=2.035
+ $X2=0 $Y2=0
cc_881 N_RESET_B_c_976_n N_A_415_81#_c_2085_n 0.0152319f $X=3.605 $Y=2.037 $X2=0
+ $Y2=0
cc_882 N_RESET_B_c_977_n N_A_415_81#_c_2085_n 0.0228135f $X=3.95 $Y=1.995 $X2=0
+ $Y2=0
cc_883 N_RESET_B_c_970_n N_A_415_81#_c_2091_n 0.00485112f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_884 N_RESET_B_c_970_n N_A_415_81#_c_2092_n 0.0021067f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_885 N_RESET_B_c_970_n N_A_415_81#_c_2087_n 0.0037715f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_886 N_RESET_B_c_970_n N_A_415_81#_c_2093_n 0.0160834f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_887 N_RESET_B_c_970_n N_A_415_81#_c_2094_n 0.0155324f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_888 N_RESET_B_c_970_n N_A_415_81#_c_2089_n 0.011933f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_889 N_RESET_B_c_964_n N_A_415_81#_c_2097_n 0.0197998f $X=3.605 $Y=2.245 $X2=0
+ $Y2=0
cc_890 N_RESET_B_c_971_n N_A_415_81#_c_2097_n 4.98701e-19 $X=4.225 $Y=2.035
+ $X2=0 $Y2=0
cc_891 N_RESET_B_c_976_n N_A_415_81#_c_2097_n 0.00783424f $X=3.605 $Y=2.037
+ $X2=0 $Y2=0
cc_892 N_RESET_B_c_977_n N_A_415_81#_c_2097_n 0.0168153f $X=3.95 $Y=1.995 $X2=0
+ $Y2=0
cc_893 N_RESET_B_c_970_n N_A_415_81#_c_2098_n 0.00682901f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_894 N_RESET_B_c_971_n N_A_415_81#_c_2098_n 0.00378634f $X=4.225 $Y=2.035
+ $X2=0 $Y2=0
cc_895 N_RESET_B_c_976_n N_A_415_81#_c_2098_n 0.0025272f $X=3.605 $Y=2.037 $X2=0
+ $Y2=0
cc_896 N_RESET_B_c_977_n N_A_415_81#_c_2098_n 0.00812968f $X=3.95 $Y=1.995 $X2=0
+ $Y2=0
cc_897 N_RESET_B_c_970_n N_A_415_81#_c_2135_n 0.0133121f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_898 N_RESET_B_M1012_g N_VGND_c_2313_n 0.00348169f $X=3.575 $Y=0.615 $X2=0
+ $Y2=0
cc_899 N_RESET_B_c_955_n N_VGND_c_2313_n 0.0231933f $X=7.225 $Y=0.18 $X2=0 $Y2=0
cc_900 N_RESET_B_c_955_n N_VGND_c_2314_n 0.02563f $X=7.225 $Y=0.18 $X2=0 $Y2=0
cc_901 N_RESET_B_c_955_n N_VGND_c_2315_n 0.0529861f $X=7.225 $Y=0.18 $X2=0 $Y2=0
cc_902 N_RESET_B_M1038_g N_VGND_c_2316_n 0.0101056f $X=10.63 $Y=0.58 $X2=0 $Y2=0
cc_903 N_RESET_B_c_956_n N_VGND_c_2320_n 0.00659533f $X=3.65 $Y=0.18 $X2=0 $Y2=0
cc_904 N_RESET_B_c_955_n N_VGND_c_2323_n 0.0211036f $X=7.225 $Y=0.18 $X2=0 $Y2=0
cc_905 N_RESET_B_M1038_g N_VGND_c_2325_n 0.00383152f $X=10.63 $Y=0.58 $X2=0
+ $Y2=0
cc_906 N_RESET_B_c_955_n N_VGND_c_2329_n 0.0108145f $X=7.225 $Y=0.18 $X2=0 $Y2=0
cc_907 N_RESET_B_c_955_n N_VGND_c_2334_n 0.0859068f $X=7.225 $Y=0.18 $X2=0 $Y2=0
cc_908 N_RESET_B_c_956_n N_VGND_c_2334_n 0.0113881f $X=3.65 $Y=0.18 $X2=0 $Y2=0
cc_909 N_RESET_B_M1038_g N_VGND_c_2334_n 0.0075694f $X=10.63 $Y=0.58 $X2=0 $Y2=0
cc_910 N_RESET_B_M1012_g N_noxref_24_c_2457_n 0.00165018f $X=3.575 $Y=0.615
+ $X2=0 $Y2=0
cc_911 N_A_1236_138#_c_1189_n N_A_837_98#_c_1329_n 0.00405916f $X=6.715 $Y=2.59
+ $X2=0 $Y2=0
cc_912 N_A_1236_138#_c_1186_n N_A_837_98#_c_1318_n 0.0049036f $X=6.32 $Y=0.87
+ $X2=0 $Y2=0
cc_913 N_A_1236_138#_c_1189_n N_A_837_98#_c_1331_n 6.3693e-19 $X=6.715 $Y=2.59
+ $X2=0 $Y2=0
cc_914 N_A_1236_138#_c_1193_n N_A_837_98#_c_1331_n 3.29021e-19 $X=6.8 $Y=2.537
+ $X2=0 $Y2=0
cc_915 N_A_1236_138#_c_1189_n N_A_837_98#_c_1333_n 0.0126759f $X=6.715 $Y=2.59
+ $X2=0 $Y2=0
cc_916 N_A_1236_138#_c_1181_n N_A_837_98#_c_1333_n 0.00130784f $X=6.8 $Y=2.32
+ $X2=0 $Y2=0
cc_917 N_A_1236_138#_c_1188_n N_A_837_98#_c_1334_n 0.0103487f $X=8.675 $Y=1.66
+ $X2=0 $Y2=0
cc_918 N_A_1236_138#_c_1225_n N_A_837_98#_c_1334_n 0.00319775f $X=7.495 $Y=2.405
+ $X2=0 $Y2=0
cc_919 N_A_1236_138#_c_1182_n N_A_837_98#_c_1334_n 0.00775183f $X=7.58 $Y=2.32
+ $X2=0 $Y2=0
cc_920 N_A_1236_138#_c_1193_n N_A_837_98#_c_1334_n 0.00142193f $X=6.8 $Y=2.537
+ $X2=0 $Y2=0
cc_921 N_A_1236_138#_c_1188_n N_A_837_98#_c_1335_n 0.00230914f $X=8.675 $Y=1.66
+ $X2=0 $Y2=0
cc_922 N_A_1236_138#_c_1188_n N_A_837_98#_M1042_g 0.00599467f $X=8.675 $Y=1.66
+ $X2=0 $Y2=0
cc_923 N_A_1236_138#_c_1180_n N_A_837_98#_c_1320_n 0.00718094f $X=8.585 $Y=1.52
+ $X2=0 $Y2=0
cc_924 N_A_1236_138#_c_1225_n N_VPWR_M1009_d 0.00824542f $X=7.495 $Y=2.405 $X2=0
+ $Y2=0
cc_925 N_A_1236_138#_c_1182_n N_VPWR_M1009_d 3.72881e-19 $X=7.58 $Y=2.32 $X2=0
+ $Y2=0
cc_926 N_A_1236_138#_c_1225_n N_VPWR_c_1892_n 0.0249179f $X=7.495 $Y=2.405 $X2=0
+ $Y2=0
cc_927 N_A_1236_138#_c_1182_n N_VPWR_c_1892_n 0.00848094f $X=7.58 $Y=2.32 $X2=0
+ $Y2=0
cc_928 N_A_1236_138#_c_1193_n N_VPWR_c_1892_n 0.00558555f $X=6.8 $Y=2.537 $X2=0
+ $Y2=0
cc_929 N_A_1236_138#_c_1182_n N_VPWR_c_1893_n 0.00731736f $X=7.58 $Y=2.32 $X2=0
+ $Y2=0
cc_930 N_A_1236_138#_c_1180_n N_VPWR_c_1894_n 0.00426403f $X=8.585 $Y=1.52 $X2=0
+ $Y2=0
cc_931 N_A_1236_138#_c_1188_n N_VPWR_c_1894_n 0.00771875f $X=8.675 $Y=1.66 $X2=0
+ $Y2=0
cc_932 N_A_1236_138#_c_1182_n N_VPWR_c_1894_n 0.0227303f $X=7.58 $Y=2.32 $X2=0
+ $Y2=0
cc_933 N_A_1236_138#_c_1189_n N_VPWR_c_1908_n 0.00990874f $X=6.715 $Y=2.59 $X2=0
+ $Y2=0
cc_934 N_A_1236_138#_c_1193_n N_VPWR_c_1908_n 0.00390498f $X=6.8 $Y=2.537 $X2=0
+ $Y2=0
cc_935 N_A_1236_138#_c_1188_n N_VPWR_c_1889_n 9.39239e-19 $X=8.675 $Y=1.66 $X2=0
+ $Y2=0
cc_936 N_A_1236_138#_c_1189_n N_VPWR_c_1889_n 0.0123809f $X=6.715 $Y=2.59 $X2=0
+ $Y2=0
cc_937 N_A_1236_138#_c_1225_n N_VPWR_c_1889_n 0.00931484f $X=7.495 $Y=2.405
+ $X2=0 $Y2=0
cc_938 N_A_1236_138#_c_1182_n N_VPWR_c_1889_n 0.0155791f $X=7.58 $Y=2.32 $X2=0
+ $Y2=0
cc_939 N_A_1236_138#_c_1193_n N_VPWR_c_1889_n 0.00468883f $X=6.8 $Y=2.537 $X2=0
+ $Y2=0
cc_940 N_A_1236_138#_c_1186_n N_A_415_81#_c_2086_n 0.0157845f $X=6.32 $Y=0.87
+ $X2=0 $Y2=0
cc_941 N_A_1236_138#_c_1189_n N_A_415_81#_c_2092_n 0.0139505f $X=6.715 $Y=2.59
+ $X2=0 $Y2=0
cc_942 N_A_1236_138#_c_1181_n N_A_415_81#_c_2092_n 0.00162745f $X=6.8 $Y=2.32
+ $X2=0 $Y2=0
cc_943 N_A_1236_138#_c_1202_n N_A_415_81#_c_2087_n 0.00571315f $X=6.715 $Y=0.99
+ $X2=0 $Y2=0
cc_944 N_A_1236_138#_c_1181_n N_A_415_81#_c_2087_n 0.0135846f $X=6.8 $Y=2.32
+ $X2=0 $Y2=0
cc_945 N_A_1236_138#_c_1186_n N_A_415_81#_c_2087_n 0.0203409f $X=6.32 $Y=0.87
+ $X2=0 $Y2=0
cc_946 N_A_1236_138#_c_1189_n N_A_415_81#_c_2093_n 0.0210559f $X=6.715 $Y=2.59
+ $X2=0 $Y2=0
cc_947 N_A_1236_138#_c_1181_n N_A_415_81#_c_2093_n 0.0141771f $X=6.8 $Y=2.32
+ $X2=0 $Y2=0
cc_948 N_A_1236_138#_c_1181_n N_A_415_81#_c_2089_n 0.0485656f $X=6.8 $Y=2.32
+ $X2=0 $Y2=0
cc_949 N_A_1236_138#_c_1193_n A_1342_463# 0.00298041f $X=6.8 $Y=2.537 $X2=-0.19
+ $Y2=-0.245
cc_950 N_A_1236_138#_M1019_g N_VGND_c_2324_n 0.00278271f $X=8.175 $Y=0.74 $X2=0
+ $Y2=0
cc_951 N_A_1236_138#_M1019_g N_VGND_c_2329_n 0.00118431f $X=8.175 $Y=0.74 $X2=0
+ $Y2=0
cc_952 N_A_1236_138#_M1019_g N_VGND_c_2334_n 0.00358928f $X=8.175 $Y=0.74 $X2=0
+ $Y2=0
cc_953 N_A_1236_138#_c_1202_n A_1322_138# 0.00343237f $X=6.715 $Y=0.99 $X2=-0.19
+ $Y2=-0.245
cc_954 N_A_1236_138#_c_1181_n A_1322_138# 3.8017e-19 $X=6.8 $Y=2.32 $X2=-0.19
+ $Y2=-0.245
cc_955 N_A_837_98#_M1027_g N_A_2003_48#_M1021_g 0.0336121f $X=9.7 $Y=0.58 $X2=0
+ $Y2=0
cc_956 N_A_837_98#_c_1319_n N_A_2003_48#_c_1520_n 0.00387806f $X=9.625 $Y=1.585
+ $X2=0 $Y2=0
cc_957 N_A_837_98#_M1027_g N_A_2003_48#_c_1524_n 0.00111235f $X=9.7 $Y=0.58
+ $X2=0 $Y2=0
cc_958 N_A_837_98#_c_1319_n N_A_2003_48#_c_1525_n 0.0336121f $X=9.625 $Y=1.585
+ $X2=0 $Y2=0
cc_959 N_A_837_98#_M1027_g N_A_1745_74#_c_1641_n 0.0163048f $X=9.7 $Y=0.58 $X2=0
+ $Y2=0
cc_960 N_A_837_98#_c_1335_n N_A_1745_74#_c_1630_n 0.00242116f $X=9.125 $Y=2.9
+ $X2=0 $Y2=0
cc_961 N_A_837_98#_M1042_g N_A_1745_74#_c_1630_n 0.00427038f $X=9.125 $Y=2.235
+ $X2=0 $Y2=0
cc_962 N_A_837_98#_M1027_g N_A_1745_74#_c_1617_n 0.00585097f $X=9.7 $Y=0.58
+ $X2=0 $Y2=0
cc_963 N_A_837_98#_c_1319_n N_A_1745_74#_c_1618_n 0.00934901f $X=9.625 $Y=1.585
+ $X2=0 $Y2=0
cc_964 N_A_837_98#_M1027_g N_A_1745_74#_c_1618_n 0.0140808f $X=9.7 $Y=0.58 $X2=0
+ $Y2=0
cc_965 N_A_837_98#_M1027_g N_A_1745_74#_c_1619_n 0.00333053f $X=9.7 $Y=0.58
+ $X2=0 $Y2=0
cc_966 N_A_837_98#_c_1319_n N_A_1745_74#_c_1632_n 3.21304e-19 $X=9.625 $Y=1.585
+ $X2=0 $Y2=0
cc_967 N_A_837_98#_M1027_g N_A_1745_74#_c_1620_n 0.00274755f $X=9.7 $Y=0.58
+ $X2=0 $Y2=0
cc_968 N_A_837_98#_c_1341_n N_VPWR_M1030_d 2.73365e-19 $X=4.805 $Y=1.905 $X2=0
+ $Y2=0
cc_969 N_A_837_98#_c_1324_n N_VPWR_M1030_d 0.00163893f $X=5.115 $Y=1.61 $X2=0
+ $Y2=0
cc_970 N_A_837_98#_M1034_g N_VPWR_c_1891_n 0.00850453f $X=5.095 $Y=2.46 $X2=0
+ $Y2=0
cc_971 N_A_837_98#_c_1316_n N_VPWR_c_1891_n 0.00158412f $X=5.615 $Y=3.075 $X2=0
+ $Y2=0
cc_972 N_A_837_98#_c_1330_n N_VPWR_c_1891_n 0.00232909f $X=5.69 $Y=3.15 $X2=0
+ $Y2=0
cc_973 N_A_837_98#_c_1331_n N_VPWR_c_1892_n 0.0060536f $X=6.635 $Y=2.9 $X2=0
+ $Y2=0
cc_974 N_A_837_98#_c_1334_n N_VPWR_c_1892_n 0.0264476f $X=9.035 $Y=3.15 $X2=0
+ $Y2=0
cc_975 N_A_837_98#_c_1334_n N_VPWR_c_1893_n 0.0260616f $X=9.035 $Y=3.15 $X2=0
+ $Y2=0
cc_976 N_A_837_98#_c_1334_n N_VPWR_c_1894_n 0.0170937f $X=9.035 $Y=3.15 $X2=0
+ $Y2=0
cc_977 N_A_837_98#_c_1335_n N_VPWR_c_1894_n 0.00527525f $X=9.125 $Y=2.9 $X2=0
+ $Y2=0
cc_978 N_A_837_98#_c_1334_n N_VPWR_c_1904_n 0.0212209f $X=9.035 $Y=3.15 $X2=0
+ $Y2=0
cc_979 N_A_837_98#_M1034_g N_VPWR_c_1908_n 0.00303678f $X=5.095 $Y=2.46 $X2=0
+ $Y2=0
cc_980 N_A_837_98#_c_1330_n N_VPWR_c_1908_n 0.0467195f $X=5.69 $Y=3.15 $X2=0
+ $Y2=0
cc_981 N_A_837_98#_M1034_g N_VPWR_c_1889_n 0.00394737f $X=5.095 $Y=2.46 $X2=0
+ $Y2=0
cc_982 N_A_837_98#_c_1329_n N_VPWR_c_1889_n 0.0245043f $X=6.545 $Y=3.15 $X2=0
+ $Y2=0
cc_983 N_A_837_98#_c_1330_n N_VPWR_c_1889_n 0.00688721f $X=5.69 $Y=3.15 $X2=0
+ $Y2=0
cc_984 N_A_837_98#_c_1334_n N_VPWR_c_1889_n 0.0714547f $X=9.035 $Y=3.15 $X2=0
+ $Y2=0
cc_985 N_A_837_98#_c_1340_n N_VPWR_c_1889_n 0.00495681f $X=6.635 $Y=3.15 $X2=0
+ $Y2=0
cc_986 N_A_837_98#_M1034_g N_A_415_81#_c_2091_n 0.0142972f $X=5.095 $Y=2.46
+ $X2=0 $Y2=0
cc_987 N_A_837_98#_c_1316_n N_A_415_81#_c_2091_n 0.0135518f $X=5.615 $Y=3.075
+ $X2=0 $Y2=0
cc_988 N_A_837_98#_c_1324_n N_A_415_81#_c_2091_n 0.0051603f $X=5.115 $Y=1.61
+ $X2=0 $Y2=0
cc_989 N_A_837_98#_c_1317_n N_A_415_81#_c_2086_n 0.00728271f $X=6.03 $Y=1.26
+ $X2=0 $Y2=0
cc_990 N_A_837_98#_c_1318_n N_A_415_81#_c_2086_n 0.00400671f $X=6.105 $Y=1.185
+ $X2=0 $Y2=0
cc_991 N_A_837_98#_c_1316_n N_A_415_81#_c_2092_n 0.00867519f $X=5.615 $Y=3.075
+ $X2=0 $Y2=0
cc_992 N_A_837_98#_c_1329_n N_A_415_81#_c_2092_n 0.00566688f $X=6.545 $Y=3.15
+ $X2=0 $Y2=0
cc_993 N_A_837_98#_c_1333_n N_A_415_81#_c_2092_n 5.20664e-19 $X=6.635 $Y=2.81
+ $X2=0 $Y2=0
cc_994 N_A_837_98#_c_1317_n N_A_415_81#_c_2087_n 0.0110024f $X=6.03 $Y=1.26
+ $X2=0 $Y2=0
cc_995 N_A_837_98#_c_1315_n N_A_415_81#_c_2088_n 0.00185966f $X=5.615 $Y=1.56
+ $X2=0 $Y2=0
cc_996 N_A_837_98#_c_1317_n N_A_415_81#_c_2088_n 0.0051163f $X=6.03 $Y=1.26
+ $X2=0 $Y2=0
cc_997 N_A_837_98#_c_1333_n N_A_415_81#_c_2093_n 6.723e-19 $X=6.635 $Y=2.81
+ $X2=0 $Y2=0
cc_998 N_A_837_98#_c_1316_n N_A_415_81#_c_2094_n 0.00159754f $X=5.615 $Y=3.075
+ $X2=0 $Y2=0
cc_999 N_A_837_98#_c_1315_n N_A_415_81#_c_2089_n 0.00407901f $X=5.615 $Y=1.56
+ $X2=0 $Y2=0
cc_1000 N_A_837_98#_M1030_s N_A_415_81#_c_2098_n 0.00816674f $X=4.275 $Y=1.96
+ $X2=0 $Y2=0
cc_1001 N_A_837_98#_c_1341_n N_A_415_81#_c_2098_n 5.63361e-19 $X=4.805 $Y=1.905
+ $X2=0 $Y2=0
cc_1002 N_A_837_98#_c_1342_n N_A_415_81#_c_2098_n 0.0130406f $X=4.425 $Y=1.905
+ $X2=0 $Y2=0
cc_1003 N_A_837_98#_c_1341_n N_A_415_81#_c_2135_n 0.00376251f $X=4.805 $Y=1.905
+ $X2=0 $Y2=0
cc_1004 N_A_837_98#_c_1351_n N_VGND_M1010_d 0.0076493f $X=4.805 $Y=1.005 $X2=0
+ $Y2=0
cc_1005 N_A_837_98#_c_1322_n N_VGND_M1010_d 0.0061573f $X=4.89 $Y=1.41 $X2=0
+ $Y2=0
cc_1006 N_A_837_98#_c_1323_n N_VGND_c_2313_n 0.0166884f $X=4.45 $Y=0.65 $X2=0
+ $Y2=0
cc_1007 N_A_837_98#_c_1351_n N_VGND_c_2314_n 0.0208234f $X=4.805 $Y=1.005 $X2=0
+ $Y2=0
cc_1008 N_A_837_98#_c_1323_n N_VGND_c_2314_n 0.00898519f $X=4.45 $Y=0.65 $X2=0
+ $Y2=0
cc_1009 N_A_837_98#_c_1324_n N_VGND_c_2314_n 0.00161245f $X=5.115 $Y=1.61 $X2=0
+ $Y2=0
cc_1010 N_A_837_98#_c_1325_n N_VGND_c_2314_n 4.02857e-19 $X=5.115 $Y=1.485 $X2=0
+ $Y2=0
cc_1011 N_A_837_98#_c_1326_n N_VGND_c_2314_n 0.00213166f $X=5.115 $Y=1.41 $X2=0
+ $Y2=0
cc_1012 N_A_837_98#_M1027_g N_VGND_c_2316_n 0.00156589f $X=9.7 $Y=0.58 $X2=0
+ $Y2=0
cc_1013 N_A_837_98#_c_1323_n N_VGND_c_2323_n 0.00802673f $X=4.45 $Y=0.65 $X2=0
+ $Y2=0
cc_1014 N_A_837_98#_M1027_g N_VGND_c_2324_n 0.00320499f $X=9.7 $Y=0.58 $X2=0
+ $Y2=0
cc_1015 N_A_837_98#_M1027_g N_VGND_c_2334_n 0.00443186f $X=9.7 $Y=0.58 $X2=0
+ $Y2=0
cc_1016 N_A_837_98#_c_1323_n N_VGND_c_2334_n 0.00988116f $X=4.45 $Y=0.65 $X2=0
+ $Y2=0
cc_1017 N_A_837_98#_c_1326_n N_VGND_c_2334_n 8.45315e-19 $X=5.115 $Y=1.41 $X2=0
+ $Y2=0
cc_1018 N_A_2003_48#_c_1522_n N_A_1745_74#_c_1608_n 0.00593167f $X=11.415
+ $Y=0.55 $X2=0 $Y2=0
cc_1019 N_A_2003_48#_c_1523_n N_A_1745_74#_c_1608_n 0.00443992f $X=11.5 $Y=1.385
+ $X2=0 $Y2=0
cc_1020 N_A_2003_48#_c_1527_n N_A_1745_74#_c_1609_n 0.00146716f $X=11.5 $Y=1.47
+ $X2=0 $Y2=0
cc_1021 N_A_2003_48#_c_1526_n N_A_1745_74#_c_1625_n 0.00555199f $X=11.165
+ $Y=2.52 $X2=0 $Y2=0
cc_1022 N_A_2003_48#_c_1523_n N_A_1745_74#_c_1610_n 0.00271488f $X=11.5 $Y=1.385
+ $X2=0 $Y2=0
cc_1023 N_A_2003_48#_c_1527_n N_A_1745_74#_c_1612_n 4.51356e-19 $X=11.5 $Y=1.47
+ $X2=0 $Y2=0
cc_1024 N_A_2003_48#_c_1523_n N_A_1745_74#_c_1614_n 0.00311356f $X=11.5 $Y=1.385
+ $X2=0 $Y2=0
cc_1025 N_A_2003_48#_c_1526_n N_A_1745_74#_c_1614_n 0.0136035f $X=11.165 $Y=2.52
+ $X2=0 $Y2=0
cc_1026 N_A_2003_48#_c_1527_n N_A_1745_74#_c_1614_n 0.0149058f $X=11.5 $Y=1.47
+ $X2=0 $Y2=0
cc_1027 N_A_2003_48#_M1021_g N_A_1745_74#_c_1641_n 0.00125881f $X=10.09 $Y=0.58
+ $X2=0 $Y2=0
cc_1028 N_A_2003_48#_c_1529_n N_A_1745_74#_c_1630_n 0.0108165f $X=10.255
+ $Y=2.465 $X2=0 $Y2=0
cc_1029 N_A_2003_48#_M1021_g N_A_1745_74#_c_1617_n 9.29499e-19 $X=10.09 $Y=0.58
+ $X2=0 $Y2=0
cc_1030 N_A_2003_48#_M1021_g N_A_1745_74#_c_1618_n 0.00223708f $X=10.09 $Y=0.58
+ $X2=0 $Y2=0
cc_1031 N_A_2003_48#_c_1520_n N_A_1745_74#_c_1618_n 0.00234903f $X=10.255
+ $Y=2.375 $X2=0 $Y2=0
cc_1032 N_A_2003_48#_c_1524_n N_A_1745_74#_c_1618_n 0.0167585f $X=10.18 $Y=1.39
+ $X2=0 $Y2=0
cc_1033 N_A_2003_48#_M1021_g N_A_1745_74#_c_1619_n 0.0143799f $X=10.09 $Y=0.58
+ $X2=0 $Y2=0
cc_1034 N_A_2003_48#_c_1521_n N_A_1745_74#_c_1619_n 0.0259611f $X=11.16 $Y=1.47
+ $X2=0 $Y2=0
cc_1035 N_A_2003_48#_c_1524_n N_A_1745_74#_c_1619_n 0.0242156f $X=10.18 $Y=1.39
+ $X2=0 $Y2=0
cc_1036 N_A_2003_48#_c_1525_n N_A_1745_74#_c_1619_n 0.001245f $X=10.18 $Y=1.39
+ $X2=0 $Y2=0
cc_1037 N_A_2003_48#_c_1520_n N_A_1745_74#_c_1632_n 0.00995549f $X=10.255
+ $Y=2.375 $X2=0 $Y2=0
cc_1038 N_A_2003_48#_c_1524_n N_A_1745_74#_c_1632_n 0.0210104f $X=10.18 $Y=1.39
+ $X2=0 $Y2=0
cc_1039 N_A_2003_48#_c_1525_n N_A_1745_74#_c_1632_n 0.00106876f $X=10.18 $Y=1.39
+ $X2=0 $Y2=0
cc_1040 N_A_2003_48#_c_1520_n N_A_1745_74#_c_1634_n 0.0141267f $X=10.255
+ $Y=2.375 $X2=0 $Y2=0
cc_1041 N_A_2003_48#_c_1529_n N_A_1745_74#_c_1634_n 0.00550853f $X=10.255
+ $Y=2.465 $X2=0 $Y2=0
cc_1042 N_A_2003_48#_c_1521_n N_A_1745_74#_c_1621_n 0.0247317f $X=11.16 $Y=1.47
+ $X2=0 $Y2=0
cc_1043 N_A_2003_48#_c_1522_n N_A_1745_74#_c_1621_n 0.014253f $X=11.415 $Y=0.55
+ $X2=0 $Y2=0
cc_1044 N_A_2003_48#_c_1523_n N_A_1745_74#_c_1621_n 0.0236842f $X=11.5 $Y=1.385
+ $X2=0 $Y2=0
cc_1045 N_A_2003_48#_c_1521_n N_A_1745_74#_c_1622_n 0.0121221f $X=11.16 $Y=1.47
+ $X2=0 $Y2=0
cc_1046 N_A_2003_48#_c_1522_n N_A_1745_74#_c_1622_n 0.00619797f $X=11.415
+ $Y=0.55 $X2=0 $Y2=0
cc_1047 N_A_2003_48#_c_1523_n N_A_1745_74#_c_1622_n 0.0191241f $X=11.5 $Y=1.385
+ $X2=0 $Y2=0
cc_1048 N_A_2003_48#_c_1522_n N_A_2339_74#_c_1778_n 0.026931f $X=11.415 $Y=0.55
+ $X2=0 $Y2=0
cc_1049 N_A_2003_48#_c_1523_n N_A_2339_74#_c_1778_n 0.0405862f $X=11.5 $Y=1.385
+ $X2=0 $Y2=0
cc_1050 N_A_2003_48#_c_1523_n N_A_2339_74#_c_1780_n 0.00909743f $X=11.5 $Y=1.385
+ $X2=0 $Y2=0
cc_1051 N_A_2003_48#_c_1526_n N_A_2339_74#_c_1780_n 0.00195796f $X=11.165
+ $Y=2.52 $X2=0 $Y2=0
cc_1052 N_A_2003_48#_c_1527_n N_A_2339_74#_c_1780_n 0.0157384f $X=11.5 $Y=1.47
+ $X2=0 $Y2=0
cc_1053 N_A_2003_48#_c_1529_n N_VPWR_c_1895_n 0.00888901f $X=10.255 $Y=2.465
+ $X2=0 $Y2=0
cc_1054 N_A_2003_48#_c_1530_n N_VPWR_c_1895_n 0.0309795f $X=11.165 $Y=2.75 $X2=0
+ $Y2=0
cc_1055 N_A_2003_48#_c_1526_n N_VPWR_c_1896_n 0.057723f $X=11.165 $Y=2.52 $X2=0
+ $Y2=0
cc_1056 N_A_2003_48#_c_1529_n N_VPWR_c_1904_n 0.00341164f $X=10.255 $Y=2.465
+ $X2=0 $Y2=0
cc_1057 N_A_2003_48#_c_1530_n N_VPWR_c_1909_n 0.0143991f $X=11.165 $Y=2.75 $X2=0
+ $Y2=0
cc_1058 N_A_2003_48#_c_1529_n N_VPWR_c_1889_n 0.00538309f $X=10.255 $Y=2.465
+ $X2=0 $Y2=0
cc_1059 N_A_2003_48#_c_1530_n N_VPWR_c_1889_n 0.0119711f $X=11.165 $Y=2.75 $X2=0
+ $Y2=0
cc_1060 N_A_2003_48#_M1021_g N_VGND_c_2316_n 0.00986387f $X=10.09 $Y=0.58 $X2=0
+ $Y2=0
cc_1061 N_A_2003_48#_c_1522_n N_VGND_c_2316_n 0.0104724f $X=11.415 $Y=0.55 $X2=0
+ $Y2=0
cc_1062 N_A_2003_48#_M1021_g N_VGND_c_2324_n 0.00383152f $X=10.09 $Y=0.58 $X2=0
+ $Y2=0
cc_1063 N_A_2003_48#_c_1522_n N_VGND_c_2325_n 0.0191719f $X=11.415 $Y=0.55 $X2=0
+ $Y2=0
cc_1064 N_A_2003_48#_M1021_g N_VGND_c_2334_n 0.0075725f $X=10.09 $Y=0.58 $X2=0
+ $Y2=0
cc_1065 N_A_2003_48#_c_1522_n N_VGND_c_2334_n 0.0192149f $X=11.415 $Y=0.55 $X2=0
+ $Y2=0
cc_1066 N_A_1745_74#_c_1611_n N_A_2339_74#_c_1772_n 0.00970941f $X=12.055
+ $Y=1.185 $X2=0 $Y2=0
cc_1067 N_A_1745_74#_c_1613_n N_A_2339_74#_c_1774_n 0.00924572f $X=12.415
+ $Y=1.69 $X2=0 $Y2=0
cc_1068 N_A_1745_74#_c_1616_n N_A_2339_74#_c_1774_n 0.00970941f $X=12.055
+ $Y=1.26 $X2=0 $Y2=0
cc_1069 N_A_1745_74#_c_1628_n N_A_2339_74#_c_1783_n 0.0130951f $X=12.49 $Y=1.765
+ $X2=0 $Y2=0
cc_1070 N_A_1745_74#_c_1608_n N_A_2339_74#_c_1778_n 5.54394e-19 $X=10.99 $Y=0.9
+ $X2=0 $Y2=0
cc_1071 N_A_1745_74#_c_1610_n N_A_2339_74#_c_1778_n 0.00765913f $X=11.98 $Y=1.26
+ $X2=0 $Y2=0
cc_1072 N_A_1745_74#_c_1611_n N_A_2339_74#_c_1778_n 0.0035045f $X=12.055
+ $Y=1.185 $X2=0 $Y2=0
cc_1073 N_A_1745_74#_c_1622_n N_A_2339_74#_c_1778_n 8.98164e-19 $X=11.535
+ $Y=1.117 $X2=0 $Y2=0
cc_1074 N_A_1745_74#_c_1609_n N_A_2339_74#_c_1779_n 0.00115484f $X=11.475
+ $Y=1.665 $X2=0 $Y2=0
cc_1075 N_A_1745_74#_c_1626_n N_A_2339_74#_c_1779_n 0.0135732f $X=12.04 $Y=1.765
+ $X2=0 $Y2=0
cc_1076 N_A_1745_74#_c_1612_n N_A_2339_74#_c_1779_n 6.63362e-19 $X=12.055
+ $Y=1.615 $X2=0 $Y2=0
cc_1077 N_A_1745_74#_c_1613_n N_A_2339_74#_c_1779_n 0.0137178f $X=12.415 $Y=1.69
+ $X2=0 $Y2=0
cc_1078 N_A_1745_74#_c_1628_n N_A_2339_74#_c_1779_n 0.0135773f $X=12.49 $Y=1.765
+ $X2=0 $Y2=0
cc_1079 N_A_1745_74#_c_1615_n N_A_2339_74#_c_1779_n 0.00313656f $X=12.04 $Y=1.69
+ $X2=0 $Y2=0
cc_1080 N_A_1745_74#_c_1609_n N_A_2339_74#_c_1780_n 2.72834e-19 $X=11.475
+ $Y=1.665 $X2=0 $Y2=0
cc_1081 N_A_1745_74#_c_1610_n N_A_2339_74#_c_1780_n 0.00807224f $X=11.98 $Y=1.26
+ $X2=0 $Y2=0
cc_1082 N_A_1745_74#_c_1612_n N_A_2339_74#_c_1780_n 0.0179017f $X=12.055
+ $Y=1.615 $X2=0 $Y2=0
cc_1083 N_A_1745_74#_c_1613_n N_A_2339_74#_c_1780_n 0.00885109f $X=12.415
+ $Y=1.69 $X2=0 $Y2=0
cc_1084 N_A_1745_74#_c_1614_n N_A_2339_74#_c_1780_n 0.00110135f $X=11.475
+ $Y=1.575 $X2=0 $Y2=0
cc_1085 N_A_1745_74#_c_1615_n N_A_2339_74#_c_1780_n 0.00144773f $X=12.04 $Y=1.69
+ $X2=0 $Y2=0
cc_1086 N_A_1745_74#_c_1616_n N_A_2339_74#_c_1780_n 0.00802343f $X=12.055
+ $Y=1.26 $X2=0 $Y2=0
cc_1087 N_A_1745_74#_c_1612_n N_A_2339_74#_c_1782_n 0.00212764f $X=12.055
+ $Y=1.615 $X2=0 $Y2=0
cc_1088 N_A_1745_74#_c_1613_n N_A_2339_74#_c_1782_n 0.00620598f $X=12.415
+ $Y=1.69 $X2=0 $Y2=0
cc_1089 N_A_1745_74#_c_1630_n N_VPWR_c_1895_n 0.0271933f $X=10.125 $Y=2.715
+ $X2=0 $Y2=0
cc_1090 N_A_1745_74#_c_1634_n N_VPWR_c_1895_n 0.00221611f $X=10.21 $Y=2.55 $X2=0
+ $Y2=0
cc_1091 N_A_1745_74#_c_1624_n N_VPWR_c_1896_n 0.0068494f $X=11.475 $Y=2.375
+ $X2=0 $Y2=0
cc_1092 N_A_1745_74#_c_1625_n N_VPWR_c_1896_n 0.0116785f $X=11.475 $Y=2.465
+ $X2=0 $Y2=0
cc_1093 N_A_1745_74#_c_1610_n N_VPWR_c_1896_n 0.00368592f $X=11.98 $Y=1.26 $X2=0
+ $Y2=0
cc_1094 N_A_1745_74#_c_1626_n N_VPWR_c_1896_n 0.00713044f $X=12.04 $Y=1.765
+ $X2=0 $Y2=0
cc_1095 N_A_1745_74#_c_1628_n N_VPWR_c_1897_n 0.0107123f $X=12.49 $Y=1.765 $X2=0
+ $Y2=0
cc_1096 N_A_1745_74#_c_1630_n N_VPWR_c_1904_n 0.0274709f $X=10.125 $Y=2.715
+ $X2=0 $Y2=0
cc_1097 N_A_1745_74#_c_1625_n N_VPWR_c_1909_n 0.00461464f $X=11.475 $Y=2.465
+ $X2=0 $Y2=0
cc_1098 N_A_1745_74#_c_1626_n N_VPWR_c_1910_n 0.00393873f $X=12.04 $Y=1.765
+ $X2=0 $Y2=0
cc_1099 N_A_1745_74#_c_1628_n N_VPWR_c_1910_n 0.00393873f $X=12.49 $Y=1.765
+ $X2=0 $Y2=0
cc_1100 N_A_1745_74#_c_1625_n N_VPWR_c_1889_n 0.00990964f $X=11.475 $Y=2.465
+ $X2=0 $Y2=0
cc_1101 N_A_1745_74#_c_1626_n N_VPWR_c_1889_n 0.00462577f $X=12.04 $Y=1.765
+ $X2=0 $Y2=0
cc_1102 N_A_1745_74#_c_1628_n N_VPWR_c_1889_n 0.00462577f $X=12.49 $Y=1.765
+ $X2=0 $Y2=0
cc_1103 N_A_1745_74#_c_1630_n N_VPWR_c_1889_n 0.0333279f $X=10.125 $Y=2.715
+ $X2=0 $Y2=0
cc_1104 N_A_1745_74#_c_1630_n A_1982_508# 0.00498821f $X=10.125 $Y=2.715
+ $X2=-0.19 $Y2=-0.245
cc_1105 N_A_1745_74#_c_1608_n N_VGND_c_2316_n 0.00154514f $X=10.99 $Y=0.9 $X2=0
+ $Y2=0
cc_1106 N_A_1745_74#_c_1641_n N_VGND_c_2316_n 0.011455f $X=9.585 $Y=0.57 $X2=0
+ $Y2=0
cc_1107 N_A_1745_74#_c_1619_n N_VGND_c_2316_n 0.0267689f $X=10.915 $Y=0.97 $X2=0
+ $Y2=0
cc_1108 N_A_1745_74#_c_1611_n N_VGND_c_2317_n 0.0149682f $X=12.055 $Y=1.185
+ $X2=0 $Y2=0
cc_1109 N_A_1745_74#_c_1641_n N_VGND_c_2324_n 0.0190071f $X=9.585 $Y=0.57 $X2=0
+ $Y2=0
cc_1110 N_A_1745_74#_c_1608_n N_VGND_c_2325_n 0.00433941f $X=10.99 $Y=0.9 $X2=0
+ $Y2=0
cc_1111 N_A_1745_74#_c_1611_n N_VGND_c_2325_n 0.00383152f $X=12.055 $Y=1.185
+ $X2=0 $Y2=0
cc_1112 N_A_1745_74#_c_1608_n N_VGND_c_2334_n 0.00822721f $X=10.99 $Y=0.9 $X2=0
+ $Y2=0
cc_1113 N_A_1745_74#_c_1611_n N_VGND_c_2334_n 0.00762539f $X=12.055 $Y=1.185
+ $X2=0 $Y2=0
cc_1114 N_A_1745_74#_c_1641_n N_VGND_c_2334_n 0.0200126f $X=9.585 $Y=0.57 $X2=0
+ $Y2=0
cc_1115 N_A_2339_74#_c_1779_n N_VPWR_c_1896_n 0.059064f $X=12.265 $Y=1.985 $X2=0
+ $Y2=0
cc_1116 N_A_2339_74#_c_1780_n N_VPWR_c_1896_n 0.0106252f $X=12.43 $Y=1.435 $X2=0
+ $Y2=0
cc_1117 N_A_2339_74#_c_1773_n N_VPWR_c_1897_n 9.84896e-19 $X=12.84 $Y=1.3 $X2=0
+ $Y2=0
cc_1118 N_A_2339_74#_c_1783_n N_VPWR_c_1897_n 0.0091433f $X=13.025 $Y=1.765
+ $X2=0 $Y2=0
cc_1119 N_A_2339_74#_c_1779_n N_VPWR_c_1897_n 0.0579567f $X=12.265 $Y=1.985
+ $X2=0 $Y2=0
cc_1120 N_A_2339_74#_c_1781_n N_VPWR_c_1897_n 0.0181117f $X=13.685 $Y=1.435
+ $X2=0 $Y2=0
cc_1121 N_A_2339_74#_c_1782_n N_VPWR_c_1897_n 0.00116289f $X=14.375 $Y=1.495
+ $X2=0 $Y2=0
cc_1122 N_A_2339_74#_c_1783_n N_VPWR_c_1898_n 0.00445602f $X=13.025 $Y=1.765
+ $X2=0 $Y2=0
cc_1123 N_A_2339_74#_c_1784_n N_VPWR_c_1898_n 0.00445602f $X=13.475 $Y=1.765
+ $X2=0 $Y2=0
cc_1124 N_A_2339_74#_c_1784_n N_VPWR_c_1899_n 0.00653972f $X=13.475 $Y=1.765
+ $X2=0 $Y2=0
cc_1125 N_A_2339_74#_c_1785_n N_VPWR_c_1899_n 0.0140029f $X=13.925 $Y=1.765
+ $X2=0 $Y2=0
cc_1126 N_A_2339_74#_c_1786_n N_VPWR_c_1899_n 5.97443e-19 $X=14.375 $Y=1.765
+ $X2=0 $Y2=0
cc_1127 N_A_2339_74#_c_1786_n N_VPWR_c_1901_n 0.00671837f $X=14.375 $Y=1.765
+ $X2=0 $Y2=0
cc_1128 N_A_2339_74#_c_1779_n N_VPWR_c_1910_n 0.00664674f $X=12.265 $Y=1.985
+ $X2=0 $Y2=0
cc_1129 N_A_2339_74#_c_1785_n N_VPWR_c_1911_n 0.00413917f $X=13.925 $Y=1.765
+ $X2=0 $Y2=0
cc_1130 N_A_2339_74#_c_1786_n N_VPWR_c_1911_n 0.00461464f $X=14.375 $Y=1.765
+ $X2=0 $Y2=0
cc_1131 N_A_2339_74#_c_1783_n N_VPWR_c_1889_n 0.00862391f $X=13.025 $Y=1.765
+ $X2=0 $Y2=0
cc_1132 N_A_2339_74#_c_1784_n N_VPWR_c_1889_n 0.00857589f $X=13.475 $Y=1.765
+ $X2=0 $Y2=0
cc_1133 N_A_2339_74#_c_1785_n N_VPWR_c_1889_n 0.00817726f $X=13.925 $Y=1.765
+ $X2=0 $Y2=0
cc_1134 N_A_2339_74#_c_1786_n N_VPWR_c_1889_n 0.00911437f $X=14.375 $Y=1.765
+ $X2=0 $Y2=0
cc_1135 N_A_2339_74#_c_1779_n N_VPWR_c_1889_n 0.00995652f $X=12.265 $Y=1.985
+ $X2=0 $Y2=0
cc_1136 N_A_2339_74#_c_1772_n N_Q_c_2245_n 0.00667713f $X=12.485 $Y=1.225 $X2=0
+ $Y2=0
cc_1137 N_A_2339_74#_c_1775_n N_Q_c_2245_n 0.0125407f $X=12.915 $Y=1.225 $X2=0
+ $Y2=0
cc_1138 N_A_2339_74#_c_1775_n N_Q_c_2256_n 0.0131906f $X=12.915 $Y=1.225 $X2=0
+ $Y2=0
cc_1139 N_A_2339_74#_c_1776_n N_Q_c_2256_n 0.0164113f $X=13.955 $Y=1.225 $X2=0
+ $Y2=0
cc_1140 N_A_2339_74#_c_1781_n N_Q_c_2256_n 0.0693421f $X=13.685 $Y=1.435 $X2=0
+ $Y2=0
cc_1141 N_A_2339_74#_c_1782_n N_Q_c_2256_n 0.0179128f $X=14.375 $Y=1.495 $X2=0
+ $Y2=0
cc_1142 N_A_2339_74#_c_1772_n N_Q_c_2260_n 0.00205797f $X=12.485 $Y=1.225 $X2=0
+ $Y2=0
cc_1143 N_A_2339_74#_c_1773_n N_Q_c_2260_n 0.00210982f $X=12.84 $Y=1.3 $X2=0
+ $Y2=0
cc_1144 N_A_2339_74#_c_1775_n N_Q_c_2260_n 7.32094e-19 $X=12.915 $Y=1.225 $X2=0
+ $Y2=0
cc_1145 N_A_2339_74#_c_1781_n N_Q_c_2260_n 0.0218379f $X=13.685 $Y=1.435 $X2=0
+ $Y2=0
cc_1146 N_A_2339_74#_c_1783_n N_Q_c_2249_n 0.0117913f $X=13.025 $Y=1.765 $X2=0
+ $Y2=0
cc_1147 N_A_2339_74#_c_1784_n N_Q_c_2249_n 0.0130095f $X=13.475 $Y=1.765 $X2=0
+ $Y2=0
cc_1148 N_A_2339_74#_c_1785_n N_Q_c_2249_n 7.91051e-19 $X=13.925 $Y=1.765 $X2=0
+ $Y2=0
cc_1149 N_A_2339_74#_c_1784_n N_Q_c_2250_n 0.0120074f $X=13.475 $Y=1.765 $X2=0
+ $Y2=0
cc_1150 N_A_2339_74#_c_1785_n N_Q_c_2250_n 0.0157775f $X=13.925 $Y=1.765 $X2=0
+ $Y2=0
cc_1151 N_A_2339_74#_c_1781_n N_Q_c_2250_n 0.0321534f $X=13.685 $Y=1.435 $X2=0
+ $Y2=0
cc_1152 N_A_2339_74#_c_1782_n N_Q_c_2250_n 0.00943636f $X=14.375 $Y=1.495 $X2=0
+ $Y2=0
cc_1153 N_A_2339_74#_c_1783_n N_Q_c_2251_n 0.0033048f $X=13.025 $Y=1.765 $X2=0
+ $Y2=0
cc_1154 N_A_2339_74#_c_1784_n N_Q_c_2251_n 0.00132156f $X=13.475 $Y=1.765 $X2=0
+ $Y2=0
cc_1155 N_A_2339_74#_c_1779_n N_Q_c_2251_n 0.00129097f $X=12.265 $Y=1.985 $X2=0
+ $Y2=0
cc_1156 N_A_2339_74#_c_1781_n N_Q_c_2251_n 0.0276943f $X=13.685 $Y=1.435 $X2=0
+ $Y2=0
cc_1157 N_A_2339_74#_c_1782_n N_Q_c_2251_n 0.00739484f $X=14.375 $Y=1.495 $X2=0
+ $Y2=0
cc_1158 N_A_2339_74#_c_1785_n N_Q_c_2252_n 0.00471332f $X=13.925 $Y=1.765 $X2=0
+ $Y2=0
cc_1159 N_A_2339_74#_c_1786_n N_Q_c_2252_n 4.03081e-19 $X=14.375 $Y=1.765 $X2=0
+ $Y2=0
cc_1160 N_A_2339_74#_c_1776_n N_Q_c_2246_n 3.92031e-19 $X=13.955 $Y=1.225 $X2=0
+ $Y2=0
cc_1161 N_A_2339_74#_c_1777_n N_Q_c_2246_n 3.92313e-19 $X=14.385 $Y=1.225 $X2=0
+ $Y2=0
cc_1162 N_A_2339_74#_c_1776_n N_Q_c_2247_n 0.00272065f $X=13.955 $Y=1.225 $X2=0
+ $Y2=0
cc_1163 N_A_2339_74#_c_1777_n N_Q_c_2247_n 0.00240279f $X=14.385 $Y=1.225 $X2=0
+ $Y2=0
cc_1164 N_A_2339_74#_c_1781_n N_Q_c_2247_n 0.00167694f $X=13.685 $Y=1.435 $X2=0
+ $Y2=0
cc_1165 N_A_2339_74#_c_1782_n N_Q_c_2247_n 0.00901833f $X=14.375 $Y=1.495 $X2=0
+ $Y2=0
cc_1166 N_A_2339_74#_c_1786_n Q 0.0145189f $X=14.375 $Y=1.765 $X2=0 $Y2=0
cc_1167 N_A_2339_74#_c_1781_n Q 0.0194661f $X=13.685 $Y=1.435 $X2=0 $Y2=0
cc_1168 N_A_2339_74#_c_1782_n Q 0.050284f $X=14.375 $Y=1.495 $X2=0 $Y2=0
cc_1169 N_A_2339_74#_c_1772_n N_VGND_c_2317_n 0.00182441f $X=12.485 $Y=1.225
+ $X2=0 $Y2=0
cc_1170 N_A_2339_74#_c_1778_n N_VGND_c_2317_n 0.0266033f $X=11.84 $Y=0.515 $X2=0
+ $Y2=0
cc_1171 N_A_2339_74#_c_1780_n N_VGND_c_2317_n 0.0191073f $X=12.43 $Y=1.435 $X2=0
+ $Y2=0
cc_1172 N_A_2339_74#_c_1776_n N_VGND_c_2319_n 4.98647e-19 $X=13.955 $Y=1.225
+ $X2=0 $Y2=0
cc_1173 N_A_2339_74#_c_1777_n N_VGND_c_2319_n 0.0149937f $X=14.385 $Y=1.225
+ $X2=0 $Y2=0
cc_1174 N_A_2339_74#_c_1778_n N_VGND_c_2325_n 0.00749631f $X=11.84 $Y=0.515
+ $X2=0 $Y2=0
cc_1175 N_A_2339_74#_c_1776_n N_VGND_c_2326_n 0.00383152f $X=13.955 $Y=1.225
+ $X2=0 $Y2=0
cc_1176 N_A_2339_74#_c_1777_n N_VGND_c_2326_n 0.00383152f $X=14.385 $Y=1.225
+ $X2=0 $Y2=0
cc_1177 N_A_2339_74#_c_1772_n N_VGND_c_2332_n 0.00434272f $X=12.485 $Y=1.225
+ $X2=0 $Y2=0
cc_1178 N_A_2339_74#_c_1775_n N_VGND_c_2332_n 0.00434272f $X=12.915 $Y=1.225
+ $X2=0 $Y2=0
cc_1179 N_A_2339_74#_c_1775_n N_VGND_c_2333_n 0.00452683f $X=12.915 $Y=1.225
+ $X2=0 $Y2=0
cc_1180 N_A_2339_74#_c_1776_n N_VGND_c_2333_n 0.0108787f $X=13.955 $Y=1.225
+ $X2=0 $Y2=0
cc_1181 N_A_2339_74#_c_1777_n N_VGND_c_2333_n 4.44374e-19 $X=14.385 $Y=1.225
+ $X2=0 $Y2=0
cc_1182 N_A_2339_74#_c_1772_n N_VGND_c_2334_n 0.00820158f $X=12.485 $Y=1.225
+ $X2=0 $Y2=0
cc_1183 N_A_2339_74#_c_1775_n N_VGND_c_2334_n 0.00825037f $X=12.915 $Y=1.225
+ $X2=0 $Y2=0
cc_1184 N_A_2339_74#_c_1776_n N_VGND_c_2334_n 0.00752925f $X=13.955 $Y=1.225
+ $X2=0 $Y2=0
cc_1185 N_A_2339_74#_c_1777_n N_VGND_c_2334_n 0.0075754f $X=14.385 $Y=1.225
+ $X2=0 $Y2=0
cc_1186 N_A_2339_74#_c_1778_n N_VGND_c_2334_n 0.0062048f $X=11.84 $Y=0.515 $X2=0
+ $Y2=0
cc_1187 N_VPWR_M1029_d N_A_415_81#_c_2099_n 0.0108376f $X=3.11 $Y=2.32 $X2=0
+ $Y2=0
cc_1188 N_VPWR_c_1890_n N_A_415_81#_c_2099_n 0.0214041f $X=3.26 $Y=2.79 $X2=0
+ $Y2=0
cc_1189 N_VPWR_c_1889_n N_A_415_81#_c_2099_n 0.0231955f $X=14.64 $Y=3.33 $X2=0
+ $Y2=0
cc_1190 N_VPWR_M1030_d N_A_415_81#_c_2091_n 0.00468818f $X=4.72 $Y=1.96 $X2=0
+ $Y2=0
cc_1191 N_VPWR_c_1891_n N_A_415_81#_c_2091_n 0.0166205f $X=4.87 $Y=2.835 $X2=0
+ $Y2=0
cc_1192 N_VPWR_c_1902_n N_A_415_81#_c_2091_n 7.47605e-19 $X=4.705 $Y=3.33 $X2=0
+ $Y2=0
cc_1193 N_VPWR_c_1908_n N_A_415_81#_c_2091_n 0.00916817f $X=7.17 $Y=3.33 $X2=0
+ $Y2=0
cc_1194 N_VPWR_c_1889_n N_A_415_81#_c_2091_n 0.0194223f $X=14.64 $Y=3.33 $X2=0
+ $Y2=0
cc_1195 N_VPWR_c_1908_n N_A_415_81#_c_2092_n 0.00746747f $X=7.17 $Y=3.33 $X2=0
+ $Y2=0
cc_1196 N_VPWR_c_1889_n N_A_415_81#_c_2092_n 0.00906023f $X=14.64 $Y=3.33 $X2=0
+ $Y2=0
cc_1197 N_VPWR_c_1890_n N_A_415_81#_c_2096_n 0.00713257f $X=3.26 $Y=2.79 $X2=0
+ $Y2=0
cc_1198 N_VPWR_c_1907_n N_A_415_81#_c_2096_n 0.0144799f $X=3.095 $Y=3.33 $X2=0
+ $Y2=0
cc_1199 N_VPWR_c_1912_n N_A_415_81#_c_2096_n 0.0198341f $X=1.4 $Y=2.465 $X2=0
+ $Y2=0
cc_1200 N_VPWR_c_1889_n N_A_415_81#_c_2096_n 0.0119509f $X=14.64 $Y=3.33 $X2=0
+ $Y2=0
cc_1201 N_VPWR_M1029_d N_A_415_81#_c_2097_n 8.56696e-19 $X=3.11 $Y=2.32 $X2=0
+ $Y2=0
cc_1202 N_VPWR_c_1890_n N_A_415_81#_c_2097_n 0.02127f $X=3.26 $Y=2.79 $X2=0
+ $Y2=0
cc_1203 N_VPWR_c_1902_n N_A_415_81#_c_2097_n 0.0166211f $X=4.705 $Y=3.33 $X2=0
+ $Y2=0
cc_1204 N_VPWR_c_1889_n N_A_415_81#_c_2097_n 0.019787f $X=14.64 $Y=3.33 $X2=0
+ $Y2=0
cc_1205 N_VPWR_c_1902_n N_A_415_81#_c_2098_n 0.00886067f $X=4.705 $Y=3.33 $X2=0
+ $Y2=0
cc_1206 N_VPWR_c_1889_n N_A_415_81#_c_2098_n 0.0167394f $X=14.64 $Y=3.33 $X2=0
+ $Y2=0
cc_1207 N_VPWR_c_1897_n N_Q_c_2249_n 0.0697297f $X=12.8 $Y=1.985 $X2=0 $Y2=0
cc_1208 N_VPWR_c_1898_n N_Q_c_2249_n 0.014552f $X=13.615 $Y=3.33 $X2=0 $Y2=0
cc_1209 N_VPWR_c_1899_n N_Q_c_2249_n 0.058364f $X=13.7 $Y=2.275 $X2=0 $Y2=0
cc_1210 N_VPWR_c_1889_n N_Q_c_2249_n 0.0119791f $X=14.64 $Y=3.33 $X2=0 $Y2=0
cc_1211 N_VPWR_M1017_d N_Q_c_2250_n 0.00222494f $X=13.55 $Y=1.84 $X2=0 $Y2=0
cc_1212 N_VPWR_c_1899_n N_Q_c_2250_n 0.0154248f $X=13.7 $Y=2.275 $X2=0 $Y2=0
cc_1213 N_VPWR_c_1897_n N_Q_c_2251_n 0.00857239f $X=12.8 $Y=1.985 $X2=0 $Y2=0
cc_1214 N_VPWR_c_1899_n N_Q_c_2252_n 0.0565072f $X=13.7 $Y=2.275 $X2=0 $Y2=0
cc_1215 N_VPWR_c_1901_n N_Q_c_2252_n 0.00140347f $X=14.6 $Y=2.275 $X2=0 $Y2=0
cc_1216 N_VPWR_c_1911_n N_Q_c_2252_n 0.00950426f $X=14.47 $Y=3.33 $X2=0 $Y2=0
cc_1217 N_VPWR_c_1889_n N_Q_c_2252_n 0.0078668f $X=14.64 $Y=3.33 $X2=0 $Y2=0
cc_1218 N_VPWR_M1039_d Q 0.0031824f $X=14.45 $Y=1.84 $X2=0 $Y2=0
cc_1219 N_VPWR_c_1901_n Q 0.0222952f $X=14.6 $Y=2.275 $X2=0 $Y2=0
cc_1220 N_A_415_81#_c_2099_n A_514_464# 0.0139074f $X=3.445 $Y=2.43 $X2=-0.19
+ $Y2=-0.245
cc_1221 N_A_415_81#_M1006_d N_noxref_24_c_2457_n 0.0094466f $X=2.075 $Y=0.405
+ $X2=0 $Y2=0
cc_1222 N_A_415_81#_c_2083_n N_noxref_24_c_2457_n 0.028856f $X=2.565 $Y=0.72
+ $X2=0 $Y2=0
cc_1223 N_A_415_81#_c_2084_n N_noxref_24_c_2457_n 0.0132335f $X=3.445 $Y=1.005
+ $X2=0 $Y2=0
cc_1224 N_A_415_81#_c_2084_n N_noxref_24_c_2475_n 0.0153497f $X=3.445 $Y=1.005
+ $X2=0 $Y2=0
cc_1225 N_Q_c_2256_n N_VGND_M1016_d 0.019527f $X=14.085 $Y=1.015 $X2=0 $Y2=0
cc_1226 N_Q_c_2245_n N_VGND_c_2317_n 0.0224879f $X=12.7 $Y=0.515 $X2=0 $Y2=0
cc_1227 N_Q_c_2246_n N_VGND_c_2319_n 0.0214745f $X=14.17 $Y=0.515 $X2=0 $Y2=0
cc_1228 N_Q_c_2247_n N_VGND_c_2319_n 0.00176181f $X=14.17 $Y=1.3 $X2=0 $Y2=0
cc_1229 Q N_VGND_c_2319_n 0.0295377f $X=14.555 $Y=1.58 $X2=0 $Y2=0
cc_1230 N_Q_c_2246_n N_VGND_c_2326_n 0.00749631f $X=14.17 $Y=0.515 $X2=0 $Y2=0
cc_1231 N_Q_c_2245_n N_VGND_c_2332_n 0.0144922f $X=12.7 $Y=0.515 $X2=0 $Y2=0
cc_1232 N_Q_c_2245_n N_VGND_c_2333_n 0.0163053f $X=12.7 $Y=0.515 $X2=0 $Y2=0
cc_1233 N_Q_c_2256_n N_VGND_c_2333_n 0.0647108f $X=14.085 $Y=1.015 $X2=0 $Y2=0
cc_1234 N_Q_c_2246_n N_VGND_c_2333_n 0.0171417f $X=14.17 $Y=0.515 $X2=0 $Y2=0
cc_1235 N_Q_c_2245_n N_VGND_c_2334_n 0.0118826f $X=12.7 $Y=0.515 $X2=0 $Y2=0
cc_1236 N_Q_c_2246_n N_VGND_c_2334_n 0.0062048f $X=14.17 $Y=0.515 $X2=0 $Y2=0
cc_1237 N_VGND_c_2313_n N_noxref_24_c_2457_n 0.0134202f $X=3.79 $Y=0.585 $X2=0
+ $Y2=0
cc_1238 N_VGND_c_2320_n N_noxref_24_c_2457_n 0.134533f $X=3.67 $Y=0 $X2=0 $Y2=0
cc_1239 N_VGND_c_2334_n N_noxref_24_c_2457_n 0.0779011f $X=14.64 $Y=0 $X2=0
+ $Y2=0
cc_1240 N_VGND_c_2312_n N_noxref_24_c_2458_n 0.0259561f $X=0.71 $Y=0.555 $X2=0
+ $Y2=0
cc_1241 N_VGND_c_2320_n N_noxref_24_c_2458_n 0.0225398f $X=3.67 $Y=0 $X2=0 $Y2=0
cc_1242 N_VGND_c_2334_n N_noxref_24_c_2458_n 0.0125704f $X=14.64 $Y=0 $X2=0
+ $Y2=0
cc_1243 N_noxref_24_c_2457_n noxref_25 0.00373495f $X=3.225 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_1244 N_noxref_24_c_2457_n noxref_26 0.0017247f $X=3.225 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
