# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ls__sdlclkp_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ls__sdlclkp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.160000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN GATE
    ANTENNAGATEAREA  0.208500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.795000 1.630000 1.300000 2.150000 ;
    END
  END GATE
  PIN GCLK
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.210000 1.820000 7.565000 2.980000 ;
        RECT 7.295000 0.350000 7.625000 1.130000 ;
        RECT 7.395000 1.130000 7.565000 1.820000 ;
    END
  END GCLK
  PIN SCE
    ANTENNAGATEAREA  0.208500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.290000 0.550000 1.960000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.498000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 5.335000 1.180000 5.665000 1.550000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 8.160000 0.085000 ;
        RECT 0.115000  0.085000 0.365000 1.120000 ;
        RECT 1.055000  0.085000 1.385000 0.370000 ;
        RECT 3.870000  0.085000 4.040000 0.735000 ;
        RECT 5.530000  0.085000 5.860000 1.010000 ;
        RECT 6.865000  0.085000 7.115000 0.790000 ;
        RECT 7.805000  0.085000 8.055000 1.130000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
        RECT 6.395000 -0.085000 6.565000 0.085000 ;
        RECT 6.875000 -0.085000 7.045000 0.085000 ;
        RECT 7.355000 -0.085000 7.525000 0.085000 ;
        RECT 7.835000 -0.085000 8.005000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.160000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 8.160000 3.415000 ;
        RECT 0.105000 2.130000 0.435000 3.245000 ;
        RECT 1.485000 2.660000 1.815000 3.245000 ;
        RECT 3.990000 2.095000 4.240000 3.245000 ;
        RECT 5.510000 2.560000 5.840000 3.245000 ;
        RECT 6.710000 2.140000 7.040000 3.245000 ;
        RECT 7.740000 1.820000 7.990000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
        RECT 6.395000 3.245000 6.565000 3.415000 ;
        RECT 6.875000 3.245000 7.045000 3.415000 ;
        RECT 7.355000 3.245000 7.525000 3.415000 ;
        RECT 7.835000 3.245000 8.005000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 8.160000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.545000 0.540000 2.375000 0.710000 ;
      RECT 0.545000 0.710000 0.890000 1.120000 ;
      RECT 0.720000 1.120000 0.890000 1.220000 ;
      RECT 0.720000 1.220000 1.640000 1.390000 ;
      RECT 0.945000 2.320000 2.800000 2.490000 ;
      RECT 0.945000 2.490000 1.275000 2.980000 ;
      RECT 1.470000 1.390000 1.640000 2.320000 ;
      RECT 1.565000 0.880000 1.980000 1.050000 ;
      RECT 1.810000 1.050000 1.980000 1.545000 ;
      RECT 1.810000 1.545000 3.020000 1.715000 ;
      RECT 1.810000 1.715000 2.340000 2.150000 ;
      RECT 2.125000 0.350000 2.375000 0.540000 ;
      RECT 2.150000 1.030000 2.715000 1.200000 ;
      RECT 2.150000 1.200000 2.480000 1.360000 ;
      RECT 2.545000 0.255000 3.700000 0.425000 ;
      RECT 2.545000 0.425000 2.715000 1.030000 ;
      RECT 2.550000 1.885000 2.800000 2.320000 ;
      RECT 2.550000 2.490000 2.800000 2.755000 ;
      RECT 2.690000 1.385000 3.020000 1.545000 ;
      RECT 2.885000 0.595000 3.360000 0.845000 ;
      RECT 3.000000 2.235000 3.360000 2.695000 ;
      RECT 3.190000 0.845000 3.360000 1.245000 ;
      RECT 3.190000 1.245000 4.485000 1.415000 ;
      RECT 3.190000 1.415000 3.360000 2.235000 ;
      RECT 3.530000 0.425000 3.700000 0.905000 ;
      RECT 3.530000 0.905000 4.380000 1.075000 ;
      RECT 3.530000 1.585000 3.860000 1.755000 ;
      RECT 3.530000 1.755000 4.825000 1.925000 ;
      RECT 4.155000 1.415000 4.485000 1.585000 ;
      RECT 4.210000 0.255000 5.360000 0.425000 ;
      RECT 4.210000 0.425000 4.380000 0.905000 ;
      RECT 4.440000 1.925000 4.825000 2.220000 ;
      RECT 4.440000 2.220000 6.005000 2.390000 ;
      RECT 4.440000 2.390000 4.825000 2.920000 ;
      RECT 4.550000 0.595000 4.825000 1.075000 ;
      RECT 4.655000 1.075000 4.825000 1.755000 ;
      RECT 4.995000 0.425000 5.360000 1.010000 ;
      RECT 4.995000 1.010000 5.165000 1.720000 ;
      RECT 4.995000 1.720000 5.310000 2.050000 ;
      RECT 5.835000 1.300000 6.530000 1.630000 ;
      RECT 5.835000 1.630000 6.005000 2.220000 ;
      RECT 6.175000 1.800000 7.040000 1.970000 ;
      RECT 6.175000 1.970000 6.505000 2.890000 ;
      RECT 6.325000 0.350000 6.655000 0.960000 ;
      RECT 6.325000 0.960000 7.040000 1.130000 ;
      RECT 6.870000 1.130000 7.040000 1.300000 ;
      RECT 6.870000 1.300000 7.225000 1.630000 ;
      RECT 6.870000 1.630000 7.040000 1.800000 ;
  END
END sky130_fd_sc_ls__sdlclkp_2
