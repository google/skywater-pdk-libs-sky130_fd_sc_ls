* File: sky130_fd_sc_ls__a211o_4.spice
* Created: Wed Sep  2 10:47:26 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__a211o_4.pex.spice"
.subckt sky130_fd_sc_ls__a211o_4  VNB VPB B1 C1 A1 A2 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A2	A2
* A1	A1
* C1	C1
* B1	B1
* VPB	VPB
* VNB	VNB
MM1001 N_X_M1001_d N_A_105_280#_M1001_g N_VGND_M1001_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1961 PD=1.02 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75004.4 A=0.111 P=1.78 MULT=1
MM1010 N_X_M1001_d N_A_105_280#_M1010_g N_VGND_M1010_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75004 A=0.111 P=1.78 MULT=1
MM1011 N_X_M1011_d N_A_105_280#_M1011_g N_VGND_M1010_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75003.6 A=0.111 P=1.78 MULT=1
MM1018 N_X_M1011_d N_A_105_280#_M1018_g N_VGND_M1018_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.130894 PD=1.02 PS=1.15826 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75003.1 A=0.111 P=1.78 MULT=1
MM1005 N_A_105_280#_M1005_d N_B1_M1005_g N_VGND_M1018_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.113206 PD=0.92 PS=1.00174 NRD=0 NRS=11.712 M=1 R=4.26667
+ SA=75002 SB=75003.1 A=0.096 P=1.58 MULT=1
MM1020 N_VGND_M1020_d N_C1_M1020_g N_A_105_280#_M1005_d VNB NSHORT L=0.15 W=0.64
+ AD=0.114925 AS=0.0896 PD=1.05 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75002.4
+ SB=75002.7 A=0.096 P=1.58 MULT=1
MM1021 N_VGND_M1020_d N_C1_M1021_g N_A_105_280#_M1021_s VNB NSHORT L=0.15 W=0.64
+ AD=0.114925 AS=0.110562 PD=1.05 PS=1.04 NRD=12.18 NRS=4.68 M=1 R=4.26667
+ SA=75002.6 SB=75002.5 A=0.096 P=1.58 MULT=1
MM1015 N_A_105_280#_M1021_s N_B1_M1015_g N_VGND_M1015_s VNB NSHORT L=0.15 W=0.64
+ AD=0.110562 AS=0.2304 PD=1.04 PS=1.36 NRD=3.744 NRS=0 M=1 R=4.26667 SA=75002.7
+ SB=75002.4 A=0.096 P=1.58 MULT=1
MM1000 N_A_1064_123#_M1000_d N_A2_M1000_g N_VGND_M1015_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.2304 PD=0.92 PS=1.36 NRD=0 NRS=82.5 M=1 R=4.26667
+ SA=75003.6 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1002 N_A_105_280#_M1002_d N_A1_M1002_g N_A_1064_123#_M1000_d VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75004
+ SB=75001.1 A=0.096 P=1.58 MULT=1
MM1017 N_A_105_280#_M1002_d N_A1_M1017_g N_A_1064_123#_M1017_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75004.4 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1022 N_A_1064_123#_M1017_s N_A2_M1022_g N_VGND_M1022_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75004.9 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1008 N_VPWR_M1008_d N_A_105_280#_M1008_g N_X_M1008_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.308 AS=0.168 PD=2.79 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75001.5 A=0.168 P=2.54 MULT=1
MM1013 N_VPWR_M1013_d N_A_105_280#_M1013_g N_X_M1008_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.6 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1016 N_VPWR_M1013_d N_A_105_280#_M1016_g N_X_M1016_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75000.6 A=0.168 P=2.54 MULT=1
MM1019 N_VPWR_M1019_d N_A_105_280#_M1019_g N_X_M1016_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.308 AS=0.168 PD=2.79 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.5 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1003 N_A_517_392#_M1003_d N_B1_M1003_g N_A_602_392#_M1003_s VPB PHIGHVT L=0.15
+ W=1 AD=0.275 AS=0.175 PD=2.55 PS=1.35 NRD=1.9503 NRS=11.8003 M=1 R=6.66667
+ SA=75000.2 SB=75003.8 A=0.15 P=2.3 MULT=1
MM1004 N_A_105_280#_M1004_d N_C1_M1004_g N_A_602_392#_M1003_s VPB PHIGHVT L=0.15
+ W=1 AD=0.15 AS=0.175 PD=1.3 PS=1.35 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75000.7 SB=75003.3 A=0.15 P=2.3 MULT=1
MM1009 N_A_105_280#_M1004_d N_C1_M1009_g N_A_602_392#_M1009_s VPB PHIGHVT L=0.15
+ W=1 AD=0.15 AS=0.1625 PD=1.3 PS=1.325 NRD=1.9503 NRS=3.9203 M=1 R=6.66667
+ SA=75001.1 SB=75002.8 A=0.15 P=2.3 MULT=1
MM1023 N_A_517_392#_M1023_d N_B1_M1023_g N_A_602_392#_M1009_s VPB PHIGHVT L=0.15
+ W=1 AD=0.1525 AS=0.1625 PD=1.305 PS=1.325 NRD=1.9503 NRS=4.9053 M=1 R=6.66667
+ SA=75001.6 SB=75002.4 A=0.15 P=2.3 MULT=1
MM1006 N_VPWR_M1006_d N_A2_M1006_g N_A_517_392#_M1023_d VPB PHIGHVT L=0.15 W=1
+ AD=0.3275 AS=0.1525 PD=1.655 PS=1.305 NRD=2.9353 NRS=2.9353 M=1 R=6.66667
+ SA=75002.1 SB=75001.9 A=0.15 P=2.3 MULT=1
MM1007 N_VPWR_M1006_d N_A1_M1007_g N_A_517_392#_M1007_s VPB PHIGHVT L=0.15 W=1
+ AD=0.3275 AS=0.15 PD=1.655 PS=1.3 NRD=2.9353 NRS=1.9503 M=1 R=6.66667
+ SA=75002.9 SB=75001.1 A=0.15 P=2.3 MULT=1
MM1012 N_VPWR_M1012_d N_A1_M1012_g N_A_517_392#_M1007_s VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75003.3
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1014 N_VPWR_M1012_d N_A2_M1014_g N_A_517_392#_M1014_s VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.275 PD=1.3 PS=2.55 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75003.8
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX24_noxref VNB VPB NWDIODE A=14.0988 P=18.88
*
.include "sky130_fd_sc_ls__a211o_4.pxi.spice"
*
.ends
*
*
