* File: sky130_fd_sc_ls__dlrtp_1.pxi.spice
* Created: Fri Aug 28 13:19:09 2020
* 
x_PM_SKY130_FD_SC_LS__DLRTP_1%D N_D_c_137_n N_D_c_138_n N_D_M1011_g N_D_M1016_g
+ D N_D_c_135_n N_D_c_136_n PM_SKY130_FD_SC_LS__DLRTP_1%D
x_PM_SKY130_FD_SC_LS__DLRTP_1%GATE N_GATE_c_167_n N_GATE_c_168_n N_GATE_M1008_g
+ N_GATE_M1002_g GATE N_GATE_c_166_n PM_SKY130_FD_SC_LS__DLRTP_1%GATE
x_PM_SKY130_FD_SC_LS__DLRTP_1%A_216_424# N_A_216_424#_M1002_d
+ N_A_216_424#_M1008_d N_A_216_424#_c_204_n N_A_216_424#_c_205_n
+ N_A_216_424#_c_221_n N_A_216_424#_M1015_g N_A_216_424#_M1010_g
+ N_A_216_424#_c_222_n N_A_216_424#_M1001_g N_A_216_424#_c_223_n
+ N_A_216_424#_c_224_n N_A_216_424#_M1006_g N_A_216_424#_c_208_n
+ N_A_216_424#_c_225_n N_A_216_424#_c_209_n N_A_216_424#_c_226_n
+ N_A_216_424#_c_210_n N_A_216_424#_c_211_n N_A_216_424#_c_212_n
+ N_A_216_424#_c_213_n N_A_216_424#_c_214_n N_A_216_424#_c_215_n
+ N_A_216_424#_c_216_n N_A_216_424#_c_217_n N_A_216_424#_c_218_n
+ N_A_216_424#_c_219_n PM_SKY130_FD_SC_LS__DLRTP_1%A_216_424#
x_PM_SKY130_FD_SC_LS__DLRTP_1%A_27_424# N_A_27_424#_M1016_s N_A_27_424#_M1011_s
+ N_A_27_424#_M1017_g N_A_27_424#_c_354_n N_A_27_424#_M1004_g
+ N_A_27_424#_c_355_n N_A_27_424#_c_360_n N_A_27_424#_c_361_n
+ N_A_27_424#_c_362_n N_A_27_424#_c_363_n N_A_27_424#_c_356_n
+ N_A_27_424#_c_357_n PM_SKY130_FD_SC_LS__DLRTP_1%A_27_424#
x_PM_SKY130_FD_SC_LS__DLRTP_1%A_363_74# N_A_363_74#_M1010_s N_A_363_74#_M1015_s
+ N_A_363_74#_M1018_g N_A_363_74#_c_451_n N_A_363_74#_M1009_g
+ N_A_363_74#_c_444_n N_A_363_74#_c_445_n N_A_363_74#_c_446_n
+ N_A_363_74#_c_503_n N_A_363_74#_c_447_n N_A_363_74#_c_454_n
+ N_A_363_74#_c_455_n N_A_363_74#_c_456_n N_A_363_74#_c_457_n
+ N_A_363_74#_c_489_n N_A_363_74#_c_448_n N_A_363_74#_c_449_n
+ N_A_363_74#_c_450_n PM_SKY130_FD_SC_LS__DLRTP_1%A_363_74#
x_PM_SKY130_FD_SC_LS__DLRTP_1%A_817_48# N_A_817_48#_M1014_s N_A_817_48#_M1019_d
+ N_A_817_48#_c_557_n N_A_817_48#_M1007_g N_A_817_48#_c_567_n
+ N_A_817_48#_M1005_g N_A_817_48#_c_558_n N_A_817_48#_c_559_n
+ N_A_817_48#_M1013_g N_A_817_48#_c_560_n N_A_817_48#_M1012_g
+ N_A_817_48#_c_561_n N_A_817_48#_c_570_n N_A_817_48#_c_562_n
+ N_A_817_48#_c_571_n N_A_817_48#_c_563_n N_A_817_48#_c_564_n
+ N_A_817_48#_c_565_n N_A_817_48#_c_572_n N_A_817_48#_c_566_n
+ PM_SKY130_FD_SC_LS__DLRTP_1%A_817_48#
x_PM_SKY130_FD_SC_LS__DLRTP_1%A_643_74# N_A_643_74#_M1018_d N_A_643_74#_M1001_d
+ N_A_643_74#_c_669_n N_A_643_74#_M1019_g N_A_643_74#_M1014_g
+ N_A_643_74#_c_664_n N_A_643_74#_c_665_n N_A_643_74#_c_666_n
+ N_A_643_74#_c_673_n N_A_643_74#_c_674_n N_A_643_74#_c_667_n
+ N_A_643_74#_c_689_n N_A_643_74#_c_675_n N_A_643_74#_c_668_n
+ PM_SKY130_FD_SC_LS__DLRTP_1%A_643_74#
x_PM_SKY130_FD_SC_LS__DLRTP_1%RESET_B N_RESET_B_M1003_g N_RESET_B_c_747_n
+ N_RESET_B_M1000_g RESET_B N_RESET_B_c_748_n
+ PM_SKY130_FD_SC_LS__DLRTP_1%RESET_B
x_PM_SKY130_FD_SC_LS__DLRTP_1%VPWR N_VPWR_M1011_d N_VPWR_M1015_d N_VPWR_M1005_d
+ N_VPWR_M1000_d N_VPWR_c_783_n N_VPWR_c_784_n N_VPWR_c_785_n N_VPWR_c_786_n
+ N_VPWR_c_787_n VPWR N_VPWR_c_788_n N_VPWR_c_789_n N_VPWR_c_790_n
+ N_VPWR_c_791_n N_VPWR_c_782_n N_VPWR_c_793_n N_VPWR_c_794_n N_VPWR_c_795_n
+ PM_SKY130_FD_SC_LS__DLRTP_1%VPWR
x_PM_SKY130_FD_SC_LS__DLRTP_1%Q N_Q_M1013_d N_Q_M1012_d N_Q_c_865_n N_Q_c_866_n
+ N_Q_c_863_n Q PM_SKY130_FD_SC_LS__DLRTP_1%Q
x_PM_SKY130_FD_SC_LS__DLRTP_1%VGND N_VGND_M1016_d N_VGND_M1010_d N_VGND_M1007_d
+ N_VGND_M1003_d N_VGND_c_886_n N_VGND_c_887_n N_VGND_c_888_n N_VGND_c_889_n
+ N_VGND_c_890_n N_VGND_c_891_n N_VGND_c_892_n N_VGND_c_893_n N_VGND_c_894_n
+ N_VGND_c_895_n VGND N_VGND_c_896_n N_VGND_c_897_n N_VGND_c_898_n
+ N_VGND_c_899_n PM_SKY130_FD_SC_LS__DLRTP_1%VGND
cc_1 VNB N_D_M1016_g 0.0302124f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=0.835
cc_2 VNB N_D_c_135_n 0.00715327f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_3 VNB N_D_c_136_n 0.0657379f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.54
cc_4 VNB N_GATE_M1002_g 0.0370084f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=0.835
cc_5 VNB GATE 0.00257351f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_6 VNB N_GATE_c_166_n 0.0243966f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.465
cc_7 VNB N_A_216_424#_c_204_n 0.0178334f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=0.835
cc_8 VNB N_A_216_424#_c_205_n 0.00889432f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_9 VNB N_A_216_424#_M1010_g 0.0363752f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.3
cc_10 VNB N_A_216_424#_M1006_g 0.0350581f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_216_424#_c_208_n 0.0103796f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_216_424#_c_209_n 0.0100621f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_216_424#_c_210_n 0.00636311f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_216_424#_c_211_n 0.00612679f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_216_424#_c_212_n 0.00201944f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_216_424#_c_213_n 0.0114186f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_216_424#_c_214_n 0.00449969f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_216_424#_c_215_n 0.00669166f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_216_424#_c_216_n 0.00498474f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_216_424#_c_217_n 0.0454379f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_216_424#_c_218_n 0.00422813f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_216_424#_c_219_n 0.0277565f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_27_424#_M1017_g 0.0349143f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_27_424#_c_354_n 0.0281964f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_27_424#_c_355_n 0.00520606f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.465
cc_26 VNB N_A_27_424#_c_356_n 0.0305779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_27_424#_c_357_n 0.0016951f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_363_74#_c_444_n 0.00268395f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_29 VNB N_A_363_74#_c_445_n 0.0198185f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.54
cc_30 VNB N_A_363_74#_c_446_n 0.00250666f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.3
cc_31 VNB N_A_363_74#_c_447_n 0.00315036f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_363_74#_c_448_n 0.0062466f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_363_74#_c_449_n 0.0315985f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_363_74#_c_450_n 0.0176429f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_817_48#_c_557_n 0.0174955f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=0.835
cc_36 VNB N_A_817_48#_c_558_n 0.0398073f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_37 VNB N_A_817_48#_c_559_n 0.0223702f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.54
cc_38 VNB N_A_817_48#_c_560_n 0.042037f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_817_48#_c_561_n 0.0294045f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_817_48#_c_562_n 0.00937344f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_817_48#_c_563_n 0.0147792f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_817_48#_c_564_n 0.00368394f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_817_48#_c_565_n 0.00566982f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_817_48#_c_566_n 0.00351959f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_643_74#_M1014_g 0.0329854f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.54
cc_46 VNB N_A_643_74#_c_664_n 0.0213847f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_47 VNB N_A_643_74#_c_665_n 0.0063868f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.54
cc_48 VNB N_A_643_74#_c_666_n 0.0126245f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.665
cc_49 VNB N_A_643_74#_c_667_n 0.00108293f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_643_74#_c_668_n 0.00575851f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_RESET_B_M1003_g 0.0237015f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.045
cc_52 VNB N_RESET_B_c_747_n 0.0268847f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.54
cc_53 VNB N_RESET_B_c_748_n 0.00165846f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.54
cc_54 VNB N_VPWR_c_782_n 0.283096f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_Q_c_863_n 0.0390828f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.54
cc_56 VNB Q 0.030012f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.3
cc_57 VNB N_VGND_c_886_n 0.0139492f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.54
cc_58 VNB N_VGND_c_887_n 0.00396956f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.665
cc_59 VNB N_VGND_c_888_n 0.0167618f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_889_n 0.00647919f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_890_n 0.0276506f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_891_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_892_n 0.0371416f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_893_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_894_n 0.0306291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_895_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_896_n 0.0362066f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_897_n 0.0234371f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_898_n 0.394164f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_899_n 0.00702378f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VPB N_D_c_137_n 0.0141841f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.955
cc_72 VPB N_D_c_138_n 0.0291586f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.045
cc_73 VPB N_D_c_135_n 0.00850726f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_74 VPB N_D_c_136_n 0.00693093f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.54
cc_75 VPB N_GATE_c_167_n 0.0113323f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.955
cc_76 VPB N_GATE_c_168_n 0.0259175f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.045
cc_77 VPB N_GATE_c_166_n 0.0104858f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.465
cc_78 VPB N_A_216_424#_c_205_n 9.19396e-19 $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_79 VPB N_A_216_424#_c_221_n 0.0279015f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 VPB N_A_216_424#_c_222_n 0.0148588f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_A_216_424#_c_223_n 0.0305493f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 VPB N_A_216_424#_c_224_n 0.0104348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 VPB N_A_216_424#_c_225_n 0.0120067f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_84 VPB N_A_216_424#_c_226_n 0.00394235f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_A_216_424#_c_214_n 0.00312026f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_A_216_424#_c_217_n 0.00892495f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_A_216_424#_c_219_n 0.00937713f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_A_27_424#_c_354_n 0.0284933f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_A_27_424#_c_355_n 0.00414363f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.465
cc_90 VPB N_A_27_424#_c_360_n 0.00887864f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB N_A_27_424#_c_361_n 0.00128825f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_92 VPB N_A_27_424#_c_362_n 0.0187571f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_A_27_424#_c_363_n 0.0225001f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB N_A_363_74#_c_451_n 0.0659882f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_95 VPB N_A_363_74#_c_444_n 0.00227193f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_96 VPB N_A_363_74#_c_447_n 0.00231101f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_A_363_74#_c_454_n 0.00619746f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_A_363_74#_c_455_n 0.00206083f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB N_A_363_74#_c_456_n 0.00176728f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 VPB N_A_363_74#_c_457_n 0.00227301f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB N_A_817_48#_c_567_n 0.0580525f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_102 VPB N_A_817_48#_c_558_n 0.0272908f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_103 VPB N_A_817_48#_c_560_n 0.0296776f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB N_A_817_48#_c_570_n 0.00407784f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_105 VPB N_A_817_48#_c_571_n 0.00289722f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_A_817_48#_c_572_n 0.00775618f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB N_A_817_48#_c_566_n 0.00253524f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_A_643_74#_c_669_n 0.0171772f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=0.835
cc_109 VPB N_A_643_74#_c_664_n 0.0179659f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_110 VPB N_A_643_74#_c_665_n 0.0107054f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.54
cc_111 VPB N_A_643_74#_c_666_n 5.50244e-19 $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.665
cc_112 VPB N_A_643_74#_c_673_n 0.0289585f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_A_643_74#_c_674_n 0.00442299f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_A_643_74#_c_675_n 0.002928f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_A_643_74#_c_668_n 0.00315278f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_RESET_B_c_747_n 0.0360911f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.54
cc_117 VPB N_RESET_B_c_748_n 0.0038344f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.54
cc_118 VPB N_VPWR_c_783_n 0.00651803f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.54
cc_119 VPB N_VPWR_c_784_n 0.0132002f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.665
cc_120 VPB N_VPWR_c_785_n 0.0137717f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_786_n 0.0185677f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_787_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_788_n 0.0191515f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_789_n 0.0438518f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_790_n 0.0436723f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_791_n 0.0198718f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_782_n 0.0932277f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_793_n 0.00614151f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_794_n 0.00700711f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_795_n 0.0180078f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_Q_c_865_n 0.041687f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_Q_c_866_n 0.0138263f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_133 VPB N_Q_c_863_n 0.00777792f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.54
cc_134 N_D_c_137_n N_GATE_c_167_n 0.00411146f $X=0.505 $Y=1.955 $X2=0 $Y2=0
cc_135 N_D_c_138_n N_GATE_c_168_n 0.0314038f $X=0.505 $Y=2.045 $X2=0 $Y2=0
cc_136 N_D_M1016_g N_GATE_M1002_g 0.0162965f $X=0.6 $Y=0.835 $X2=0 $Y2=0
cc_137 N_D_c_136_n GATE 3.32426e-19 $X=0.505 $Y=1.54 $X2=0 $Y2=0
cc_138 N_D_c_136_n N_GATE_c_166_n 0.0117846f $X=0.505 $Y=1.54 $X2=0 $Y2=0
cc_139 N_D_c_137_n N_A_27_424#_c_355_n 0.00870199f $X=0.505 $Y=1.955 $X2=0 $Y2=0
cc_140 N_D_c_138_n N_A_27_424#_c_355_n 0.00754651f $X=0.505 $Y=2.045 $X2=0 $Y2=0
cc_141 N_D_M1016_g N_A_27_424#_c_355_n 0.00990189f $X=0.6 $Y=0.835 $X2=0 $Y2=0
cc_142 N_D_c_135_n N_A_27_424#_c_355_n 0.0343288f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_143 N_D_c_136_n N_A_27_424#_c_355_n 0.0148841f $X=0.505 $Y=1.54 $X2=0 $Y2=0
cc_144 N_D_c_138_n N_A_27_424#_c_362_n 0.00733505f $X=0.505 $Y=2.045 $X2=0 $Y2=0
cc_145 N_D_c_138_n N_A_27_424#_c_363_n 0.0237728f $X=0.505 $Y=2.045 $X2=0 $Y2=0
cc_146 N_D_c_135_n N_A_27_424#_c_363_n 0.0147162f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_147 N_D_c_136_n N_A_27_424#_c_363_n 0.00275636f $X=0.505 $Y=1.54 $X2=0 $Y2=0
cc_148 N_D_M1016_g N_A_27_424#_c_356_n 0.0202375f $X=0.6 $Y=0.835 $X2=0 $Y2=0
cc_149 N_D_c_135_n N_A_27_424#_c_356_n 0.0131784f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_150 N_D_c_136_n N_A_27_424#_c_356_n 0.00817663f $X=0.505 $Y=1.54 $X2=0 $Y2=0
cc_151 N_D_c_138_n N_VPWR_c_783_n 0.00452824f $X=0.505 $Y=2.045 $X2=0 $Y2=0
cc_152 N_D_c_138_n N_VPWR_c_788_n 0.00445602f $X=0.505 $Y=2.045 $X2=0 $Y2=0
cc_153 N_D_c_138_n N_VPWR_c_782_n 0.00441841f $X=0.505 $Y=2.045 $X2=0 $Y2=0
cc_154 N_D_M1016_g N_VGND_c_886_n 0.0042545f $X=0.6 $Y=0.835 $X2=0 $Y2=0
cc_155 N_D_M1016_g N_VGND_c_890_n 0.00340649f $X=0.6 $Y=0.835 $X2=0 $Y2=0
cc_156 N_D_M1016_g N_VGND_c_898_n 0.00487769f $X=0.6 $Y=0.835 $X2=0 $Y2=0
cc_157 N_GATE_c_168_n N_A_216_424#_c_225_n 0.00670055f $X=1.005 $Y=2.045 $X2=0
+ $Y2=0
cc_158 GATE N_A_216_424#_c_225_n 0.00971996f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_159 N_GATE_c_166_n N_A_216_424#_c_225_n 0.00288243f $X=1.185 $Y=1.615 $X2=0
+ $Y2=0
cc_160 N_GATE_M1002_g N_A_216_424#_c_209_n 0.00634199f $X=1.185 $Y=0.74 $X2=0
+ $Y2=0
cc_161 N_GATE_c_167_n N_A_216_424#_c_226_n 0.00537f $X=1.005 $Y=1.955 $X2=0
+ $Y2=0
cc_162 N_GATE_M1002_g N_A_216_424#_c_213_n 0.00469117f $X=1.185 $Y=0.74 $X2=0
+ $Y2=0
cc_163 GATE N_A_216_424#_c_213_n 0.00257643f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_164 GATE N_A_216_424#_c_214_n 0.027849f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_165 N_GATE_c_166_n N_A_216_424#_c_214_n 0.00638325f $X=1.185 $Y=1.615 $X2=0
+ $Y2=0
cc_166 N_GATE_M1002_g N_A_216_424#_c_215_n 0.00531887f $X=1.185 $Y=0.74 $X2=0
+ $Y2=0
cc_167 GATE N_A_216_424#_c_219_n 0.00100641f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_168 N_GATE_c_166_n N_A_216_424#_c_219_n 0.0181923f $X=1.185 $Y=1.615 $X2=0
+ $Y2=0
cc_169 N_GATE_c_168_n N_A_27_424#_c_355_n 4.55856e-19 $X=1.005 $Y=2.045 $X2=0
+ $Y2=0
cc_170 N_GATE_M1002_g N_A_27_424#_c_355_n 0.00541079f $X=1.185 $Y=0.74 $X2=0
+ $Y2=0
cc_171 GATE N_A_27_424#_c_355_n 0.0208665f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_172 N_GATE_c_166_n N_A_27_424#_c_355_n 0.00690299f $X=1.185 $Y=1.615 $X2=0
+ $Y2=0
cc_173 N_GATE_c_168_n N_A_27_424#_c_360_n 0.0160006f $X=1.005 $Y=2.045 $X2=0
+ $Y2=0
cc_174 GATE N_A_27_424#_c_360_n 0.00481059f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_175 N_GATE_c_166_n N_A_27_424#_c_360_n 9.54685e-19 $X=1.185 $Y=1.615 $X2=0
+ $Y2=0
cc_176 N_GATE_c_168_n N_A_27_424#_c_362_n 6.02639e-19 $X=1.005 $Y=2.045 $X2=0
+ $Y2=0
cc_177 N_GATE_c_168_n N_A_27_424#_c_363_n 0.00559067f $X=1.005 $Y=2.045 $X2=0
+ $Y2=0
cc_178 N_GATE_c_168_n N_VPWR_c_783_n 0.0172571f $X=1.005 $Y=2.045 $X2=0 $Y2=0
cc_179 N_GATE_c_168_n N_VPWR_c_789_n 0.00413917f $X=1.005 $Y=2.045 $X2=0 $Y2=0
cc_180 N_GATE_c_168_n N_VPWR_c_782_n 0.00403443f $X=1.005 $Y=2.045 $X2=0 $Y2=0
cc_181 N_GATE_M1002_g N_VGND_c_886_n 0.00522565f $X=1.185 $Y=0.74 $X2=0 $Y2=0
cc_182 GATE N_VGND_c_886_n 0.00653399f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_183 N_GATE_c_166_n N_VGND_c_886_n 0.00366723f $X=1.185 $Y=1.615 $X2=0 $Y2=0
cc_184 N_GATE_M1002_g N_VGND_c_896_n 0.00434272f $X=1.185 $Y=0.74 $X2=0 $Y2=0
cc_185 N_GATE_M1002_g N_VGND_c_898_n 0.00830282f $X=1.185 $Y=0.74 $X2=0 $Y2=0
cc_186 N_A_216_424#_M1010_g N_A_27_424#_M1017_g 0.0310105f $X=2.24 $Y=0.74 $X2=0
+ $Y2=0
cc_187 N_A_216_424#_c_210_n N_A_27_424#_M1017_g 0.0111444f $X=2.85 $Y=0.855
+ $X2=0 $Y2=0
cc_188 N_A_216_424#_c_212_n N_A_27_424#_M1017_g 0.0011351f $X=3.02 $Y=0.34 $X2=0
+ $Y2=0
cc_189 N_A_216_424#_c_205_n N_A_27_424#_c_354_n 0.00960669f $X=2.185 $Y=1.795
+ $X2=0 $Y2=0
cc_190 N_A_216_424#_c_221_n N_A_27_424#_c_354_n 0.0227353f $X=2.185 $Y=1.885
+ $X2=0 $Y2=0
cc_191 N_A_216_424#_c_222_n N_A_27_424#_c_354_n 0.0467548f $X=3.185 $Y=1.885
+ $X2=0 $Y2=0
cc_192 N_A_216_424#_c_224_n N_A_27_424#_c_354_n 0.0101123f $X=3.275 $Y=1.765
+ $X2=0 $Y2=0
cc_193 N_A_216_424#_c_208_n N_A_27_424#_c_354_n 0.00863303f $X=2.205 $Y=1.525
+ $X2=0 $Y2=0
cc_194 N_A_216_424#_c_225_n N_A_27_424#_c_355_n 0.00548169f $X=1.455 $Y=2.095
+ $X2=0 $Y2=0
cc_195 N_A_216_424#_M1008_d N_A_27_424#_c_360_n 0.0146511f $X=1.08 $Y=2.12 $X2=0
+ $Y2=0
cc_196 N_A_216_424#_c_221_n N_A_27_424#_c_360_n 0.0170279f $X=2.185 $Y=1.885
+ $X2=0 $Y2=0
cc_197 N_A_216_424#_c_225_n N_A_27_424#_c_360_n 0.0368524f $X=1.455 $Y=2.095
+ $X2=0 $Y2=0
cc_198 N_A_216_424#_c_214_n N_A_27_424#_c_360_n 0.00485156f $X=1.665 $Y=1.615
+ $X2=0 $Y2=0
cc_199 N_A_216_424#_c_219_n N_A_27_424#_c_360_n 0.0012498f $X=1.665 $Y=1.525
+ $X2=0 $Y2=0
cc_200 N_A_216_424#_c_221_n N_A_27_424#_c_361_n 0.00655929f $X=2.185 $Y=1.885
+ $X2=0 $Y2=0
cc_201 N_A_216_424#_c_222_n N_A_27_424#_c_361_n 2.95897e-19 $X=3.185 $Y=1.885
+ $X2=0 $Y2=0
cc_202 N_A_216_424#_c_225_n N_A_27_424#_c_363_n 0.00516371f $X=1.455 $Y=2.095
+ $X2=0 $Y2=0
cc_203 N_A_216_424#_c_205_n N_A_27_424#_c_357_n 7.0957e-19 $X=2.185 $Y=1.795
+ $X2=0 $Y2=0
cc_204 N_A_216_424#_c_208_n N_A_27_424#_c_357_n 5.7423e-19 $X=2.205 $Y=1.525
+ $X2=0 $Y2=0
cc_205 N_A_216_424#_c_210_n N_A_363_74#_M1010_s 0.00989832f $X=2.85 $Y=0.855
+ $X2=-0.19 $Y2=-0.245
cc_206 N_A_216_424#_c_222_n N_A_363_74#_c_451_n 0.0221638f $X=3.185 $Y=1.885
+ $X2=0 $Y2=0
cc_207 N_A_216_424#_c_223_n N_A_363_74#_c_451_n 0.0139957f $X=3.695 $Y=1.765
+ $X2=0 $Y2=0
cc_208 N_A_216_424#_c_217_n N_A_363_74#_c_451_n 0.00367833f $X=3.93 $Y=1.39
+ $X2=0 $Y2=0
cc_209 N_A_216_424#_c_204_n N_A_363_74#_c_444_n 0.00704085f $X=2.095 $Y=1.525
+ $X2=0 $Y2=0
cc_210 N_A_216_424#_c_205_n N_A_363_74#_c_444_n 0.00476942f $X=2.185 $Y=1.795
+ $X2=0 $Y2=0
cc_211 N_A_216_424#_c_221_n N_A_363_74#_c_444_n 0.00706564f $X=2.185 $Y=1.885
+ $X2=0 $Y2=0
cc_212 N_A_216_424#_M1010_g N_A_363_74#_c_444_n 0.00581595f $X=2.24 $Y=0.74
+ $X2=0 $Y2=0
cc_213 N_A_216_424#_c_208_n N_A_363_74#_c_444_n 0.00421753f $X=2.205 $Y=1.525
+ $X2=0 $Y2=0
cc_214 N_A_216_424#_c_225_n N_A_363_74#_c_444_n 0.00229425f $X=1.455 $Y=2.095
+ $X2=0 $Y2=0
cc_215 N_A_216_424#_c_226_n N_A_363_74#_c_444_n 0.00822192f $X=1.54 $Y=1.97
+ $X2=0 $Y2=0
cc_216 N_A_216_424#_c_214_n N_A_363_74#_c_444_n 0.0244847f $X=1.665 $Y=1.615
+ $X2=0 $Y2=0
cc_217 N_A_216_424#_c_215_n N_A_363_74#_c_444_n 0.00729783f $X=1.642 $Y=1.45
+ $X2=0 $Y2=0
cc_218 N_A_216_424#_c_219_n N_A_363_74#_c_444_n 0.00107984f $X=1.665 $Y=1.525
+ $X2=0 $Y2=0
cc_219 N_A_216_424#_M1010_g N_A_363_74#_c_445_n 0.0128205f $X=2.24 $Y=0.74 $X2=0
+ $Y2=0
cc_220 N_A_216_424#_c_210_n N_A_363_74#_c_445_n 0.0120886f $X=2.85 $Y=0.855
+ $X2=0 $Y2=0
cc_221 N_A_216_424#_c_204_n N_A_363_74#_c_446_n 7.98985e-19 $X=2.095 $Y=1.525
+ $X2=0 $Y2=0
cc_222 N_A_216_424#_M1010_g N_A_363_74#_c_446_n 0.00369563f $X=2.24 $Y=0.74
+ $X2=0 $Y2=0
cc_223 N_A_216_424#_c_210_n N_A_363_74#_c_446_n 0.0686872f $X=2.85 $Y=0.855
+ $X2=0 $Y2=0
cc_224 N_A_216_424#_c_213_n N_A_363_74#_c_446_n 0.0142477f $X=1.43 $Y=0.855
+ $X2=0 $Y2=0
cc_225 N_A_216_424#_c_214_n N_A_363_74#_c_446_n 0.00254949f $X=1.665 $Y=1.615
+ $X2=0 $Y2=0
cc_226 N_A_216_424#_c_219_n N_A_363_74#_c_446_n 0.00611482f $X=1.665 $Y=1.525
+ $X2=0 $Y2=0
cc_227 N_A_216_424#_c_222_n N_A_363_74#_c_447_n 0.00195025f $X=3.185 $Y=1.885
+ $X2=0 $Y2=0
cc_228 N_A_216_424#_c_224_n N_A_363_74#_c_447_n 0.00644006f $X=3.275 $Y=1.765
+ $X2=0 $Y2=0
cc_229 N_A_216_424#_c_222_n N_A_363_74#_c_454_n 0.0132479f $X=3.185 $Y=1.885
+ $X2=0 $Y2=0
cc_230 N_A_216_424#_c_222_n N_A_363_74#_c_456_n 5.05727e-19 $X=3.185 $Y=1.885
+ $X2=0 $Y2=0
cc_231 N_A_216_424#_c_204_n N_A_363_74#_c_457_n 0.00481994f $X=2.095 $Y=1.525
+ $X2=0 $Y2=0
cc_232 N_A_216_424#_c_221_n N_A_363_74#_c_457_n 0.00435584f $X=2.185 $Y=1.885
+ $X2=0 $Y2=0
cc_233 N_A_216_424#_c_225_n N_A_363_74#_c_457_n 0.0172708f $X=1.455 $Y=2.095
+ $X2=0 $Y2=0
cc_234 N_A_216_424#_c_214_n N_A_363_74#_c_457_n 0.00198601f $X=1.665 $Y=1.615
+ $X2=0 $Y2=0
cc_235 N_A_216_424#_c_219_n N_A_363_74#_c_457_n 2.26279e-19 $X=1.665 $Y=1.525
+ $X2=0 $Y2=0
cc_236 N_A_216_424#_c_222_n N_A_363_74#_c_489_n 0.00783807f $X=3.185 $Y=1.885
+ $X2=0 $Y2=0
cc_237 N_A_216_424#_c_224_n N_A_363_74#_c_448_n 9.08332e-19 $X=3.275 $Y=1.765
+ $X2=0 $Y2=0
cc_238 N_A_216_424#_c_224_n N_A_363_74#_c_449_n 0.0166643f $X=3.275 $Y=1.765
+ $X2=0 $Y2=0
cc_239 N_A_216_424#_M1006_g N_A_363_74#_c_449_n 0.011696f $X=3.77 $Y=0.58 $X2=0
+ $Y2=0
cc_240 N_A_216_424#_M1006_g N_A_363_74#_c_450_n 0.0168057f $X=3.77 $Y=0.58 $X2=0
+ $Y2=0
cc_241 N_A_216_424#_c_211_n N_A_363_74#_c_450_n 0.0132006f $X=3.835 $Y=0.34
+ $X2=0 $Y2=0
cc_242 N_A_216_424#_c_218_n N_A_363_74#_c_450_n 9.76507e-19 $X=3.965 $Y=1.225
+ $X2=0 $Y2=0
cc_243 N_A_216_424#_M1006_g N_A_817_48#_c_557_n 0.0385805f $X=3.77 $Y=0.58 $X2=0
+ $Y2=0
cc_244 N_A_216_424#_c_211_n N_A_817_48#_c_557_n 0.00133249f $X=3.835 $Y=0.34
+ $X2=0 $Y2=0
cc_245 N_A_216_424#_c_218_n N_A_817_48#_c_557_n 0.00729255f $X=3.965 $Y=1.225
+ $X2=0 $Y2=0
cc_246 N_A_216_424#_M1006_g N_A_817_48#_c_558_n 0.00426541f $X=3.77 $Y=0.58
+ $X2=0 $Y2=0
cc_247 N_A_216_424#_c_216_n N_A_817_48#_c_558_n 0.00197074f $X=3.93 $Y=1.39
+ $X2=0 $Y2=0
cc_248 N_A_216_424#_c_217_n N_A_817_48#_c_558_n 0.0287556f $X=3.93 $Y=1.39 $X2=0
+ $Y2=0
cc_249 N_A_216_424#_c_218_n N_A_817_48#_c_558_n 0.00399793f $X=3.965 $Y=1.225
+ $X2=0 $Y2=0
cc_250 N_A_216_424#_c_217_n N_A_817_48#_c_561_n 6.79409e-19 $X=3.93 $Y=1.39
+ $X2=0 $Y2=0
cc_251 N_A_216_424#_c_211_n N_A_643_74#_M1018_d 0.00417255f $X=3.835 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_252 N_A_216_424#_c_223_n N_A_643_74#_c_666_n 0.00639741f $X=3.695 $Y=1.765
+ $X2=0 $Y2=0
cc_253 N_A_216_424#_M1006_g N_A_643_74#_c_666_n 0.0129937f $X=3.77 $Y=0.58 $X2=0
+ $Y2=0
cc_254 N_A_216_424#_c_218_n N_A_643_74#_c_666_n 0.0457738f $X=3.965 $Y=1.225
+ $X2=0 $Y2=0
cc_255 N_A_216_424#_c_223_n N_A_643_74#_c_673_n 0.00141716f $X=3.695 $Y=1.765
+ $X2=0 $Y2=0
cc_256 N_A_216_424#_c_216_n N_A_643_74#_c_673_n 0.020194f $X=3.93 $Y=1.39 $X2=0
+ $Y2=0
cc_257 N_A_216_424#_c_217_n N_A_643_74#_c_673_n 0.0114646f $X=3.93 $Y=1.39 $X2=0
+ $Y2=0
cc_258 N_A_216_424#_c_223_n N_A_643_74#_c_674_n 0.0135404f $X=3.695 $Y=1.765
+ $X2=0 $Y2=0
cc_259 N_A_216_424#_c_224_n N_A_643_74#_c_674_n 0.00102705f $X=3.275 $Y=1.765
+ $X2=0 $Y2=0
cc_260 N_A_216_424#_M1006_g N_A_643_74#_c_667_n 0.00278503f $X=3.77 $Y=0.58
+ $X2=0 $Y2=0
cc_261 N_A_216_424#_c_211_n N_A_643_74#_c_667_n 0.0279134f $X=3.835 $Y=0.34
+ $X2=0 $Y2=0
cc_262 N_A_216_424#_c_218_n N_A_643_74#_c_667_n 0.0170435f $X=3.965 $Y=1.225
+ $X2=0 $Y2=0
cc_263 N_A_216_424#_c_222_n N_A_643_74#_c_689_n 0.00390285f $X=3.185 $Y=1.885
+ $X2=0 $Y2=0
cc_264 N_A_216_424#_c_223_n N_A_643_74#_c_689_n 0.00164154f $X=3.695 $Y=1.765
+ $X2=0 $Y2=0
cc_265 N_A_216_424#_c_222_n N_A_643_74#_c_675_n 0.00607504f $X=3.185 $Y=1.885
+ $X2=0 $Y2=0
cc_266 N_A_216_424#_c_223_n N_A_643_74#_c_675_n 0.00151884f $X=3.695 $Y=1.765
+ $X2=0 $Y2=0
cc_267 N_A_216_424#_c_216_n N_A_643_74#_c_668_n 0.00226545f $X=3.93 $Y=1.39
+ $X2=0 $Y2=0
cc_268 N_A_216_424#_c_221_n N_VPWR_c_784_n 0.00581666f $X=2.185 $Y=1.885 $X2=0
+ $Y2=0
cc_269 N_A_216_424#_c_222_n N_VPWR_c_784_n 2.77559e-19 $X=3.185 $Y=1.885 $X2=0
+ $Y2=0
cc_270 N_A_216_424#_c_221_n N_VPWR_c_789_n 0.00469064f $X=2.185 $Y=1.885 $X2=0
+ $Y2=0
cc_271 N_A_216_424#_c_222_n N_VPWR_c_790_n 0.00278271f $X=3.185 $Y=1.885 $X2=0
+ $Y2=0
cc_272 N_A_216_424#_c_221_n N_VPWR_c_782_n 0.0049649f $X=2.185 $Y=1.885 $X2=0
+ $Y2=0
cc_273 N_A_216_424#_c_222_n N_VPWR_c_782_n 0.00354422f $X=3.185 $Y=1.885 $X2=0
+ $Y2=0
cc_274 N_A_216_424#_c_210_n N_VGND_M1010_d 0.00508382f $X=2.85 $Y=0.855 $X2=0
+ $Y2=0
cc_275 N_A_216_424#_c_209_n N_VGND_c_886_n 0.0300165f $X=1.4 $Y=0.515 $X2=0
+ $Y2=0
cc_276 N_A_216_424#_M1010_g N_VGND_c_887_n 0.0126864f $X=2.24 $Y=0.74 $X2=0
+ $Y2=0
cc_277 N_A_216_424#_c_209_n N_VGND_c_887_n 0.00713841f $X=1.4 $Y=0.515 $X2=0
+ $Y2=0
cc_278 N_A_216_424#_c_210_n N_VGND_c_887_n 0.0210746f $X=2.85 $Y=0.855 $X2=0
+ $Y2=0
cc_279 N_A_216_424#_c_212_n N_VGND_c_887_n 0.0118766f $X=3.02 $Y=0.34 $X2=0
+ $Y2=0
cc_280 N_A_216_424#_M1006_g N_VGND_c_888_n 5.44443e-19 $X=3.77 $Y=0.58 $X2=0
+ $Y2=0
cc_281 N_A_216_424#_c_211_n N_VGND_c_888_n 0.0123564f $X=3.835 $Y=0.34 $X2=0
+ $Y2=0
cc_282 N_A_216_424#_c_218_n N_VGND_c_888_n 0.0246024f $X=3.965 $Y=1.225 $X2=0
+ $Y2=0
cc_283 N_A_216_424#_M1006_g N_VGND_c_892_n 0.00278262f $X=3.77 $Y=0.58 $X2=0
+ $Y2=0
cc_284 N_A_216_424#_c_211_n N_VGND_c_892_n 0.063753f $X=3.835 $Y=0.34 $X2=0
+ $Y2=0
cc_285 N_A_216_424#_c_212_n N_VGND_c_892_n 0.0121935f $X=3.02 $Y=0.34 $X2=0
+ $Y2=0
cc_286 N_A_216_424#_M1010_g N_VGND_c_896_n 0.00398535f $X=2.24 $Y=0.74 $X2=0
+ $Y2=0
cc_287 N_A_216_424#_c_209_n N_VGND_c_896_n 0.0172412f $X=1.4 $Y=0.515 $X2=0
+ $Y2=0
cc_288 N_A_216_424#_M1010_g N_VGND_c_898_n 0.00388856f $X=2.24 $Y=0.74 $X2=0
+ $Y2=0
cc_289 N_A_216_424#_M1006_g N_VGND_c_898_n 0.00354801f $X=3.77 $Y=0.58 $X2=0
+ $Y2=0
cc_290 N_A_216_424#_c_209_n N_VGND_c_898_n 0.0142144f $X=1.4 $Y=0.515 $X2=0
+ $Y2=0
cc_291 N_A_216_424#_c_210_n N_VGND_c_898_n 0.0302804f $X=2.85 $Y=0.855 $X2=0
+ $Y2=0
cc_292 N_A_216_424#_c_211_n N_VGND_c_898_n 0.0358785f $X=3.835 $Y=0.34 $X2=0
+ $Y2=0
cc_293 N_A_216_424#_c_212_n N_VGND_c_898_n 0.00661049f $X=3.02 $Y=0.34 $X2=0
+ $Y2=0
cc_294 N_A_216_424#_c_210_n A_565_74# 0.00142466f $X=2.85 $Y=0.855 $X2=-0.19
+ $Y2=-0.245
cc_295 N_A_216_424#_c_211_n A_769_74# 5.0299e-19 $X=3.835 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_296 N_A_216_424#_c_218_n A_769_74# 0.003195f $X=3.965 $Y=1.225 $X2=-0.19
+ $Y2=-0.245
cc_297 N_A_27_424#_c_360_n N_A_363_74#_M1015_s 0.00808827f $X=2.525 $Y=2.475
+ $X2=0 $Y2=0
cc_298 N_A_27_424#_M1017_g N_A_363_74#_c_444_n 8.66064e-19 $X=2.75 $Y=0.69 $X2=0
+ $Y2=0
cc_299 N_A_27_424#_c_354_n N_A_363_74#_c_444_n 0.00120795f $X=2.765 $Y=1.885
+ $X2=0 $Y2=0
cc_300 N_A_27_424#_c_357_n N_A_363_74#_c_444_n 0.0219835f $X=2.69 $Y=1.635 $X2=0
+ $Y2=0
cc_301 N_A_27_424#_M1017_g N_A_363_74#_c_445_n 0.0101442f $X=2.75 $Y=0.69 $X2=0
+ $Y2=0
cc_302 N_A_27_424#_c_354_n N_A_363_74#_c_445_n 0.00122335f $X=2.765 $Y=1.885
+ $X2=0 $Y2=0
cc_303 N_A_27_424#_c_357_n N_A_363_74#_c_445_n 0.0228816f $X=2.69 $Y=1.635 $X2=0
+ $Y2=0
cc_304 N_A_27_424#_c_354_n N_A_363_74#_c_503_n 0.00829007f $X=2.765 $Y=1.885
+ $X2=0 $Y2=0
cc_305 N_A_27_424#_c_360_n N_A_363_74#_c_503_n 0.0113396f $X=2.525 $Y=2.475
+ $X2=0 $Y2=0
cc_306 N_A_27_424#_c_361_n N_A_363_74#_c_503_n 0.0148899f $X=2.61 $Y=2.39 $X2=0
+ $Y2=0
cc_307 N_A_27_424#_c_354_n N_A_363_74#_c_447_n 0.00674556f $X=2.765 $Y=1.885
+ $X2=0 $Y2=0
cc_308 N_A_27_424#_c_361_n N_A_363_74#_c_447_n 0.00736754f $X=2.61 $Y=2.39 $X2=0
+ $Y2=0
cc_309 N_A_27_424#_c_357_n N_A_363_74#_c_447_n 0.0248017f $X=2.69 $Y=1.635 $X2=0
+ $Y2=0
cc_310 N_A_27_424#_c_354_n N_A_363_74#_c_455_n 0.00142562f $X=2.765 $Y=1.885
+ $X2=0 $Y2=0
cc_311 N_A_27_424#_c_360_n N_A_363_74#_c_457_n 0.0230736f $X=2.525 $Y=2.475
+ $X2=0 $Y2=0
cc_312 N_A_27_424#_c_361_n N_A_363_74#_c_457_n 0.00840135f $X=2.61 $Y=2.39 $X2=0
+ $Y2=0
cc_313 N_A_27_424#_c_354_n N_A_363_74#_c_489_n 0.00129794f $X=2.765 $Y=1.885
+ $X2=0 $Y2=0
cc_314 N_A_27_424#_c_361_n N_A_363_74#_c_489_n 0.0105035f $X=2.61 $Y=2.39 $X2=0
+ $Y2=0
cc_315 N_A_27_424#_M1017_g N_A_363_74#_c_448_n 0.0044995f $X=2.75 $Y=0.69 $X2=0
+ $Y2=0
cc_316 N_A_27_424#_M1017_g N_A_363_74#_c_450_n 0.0597211f $X=2.75 $Y=0.69 $X2=0
+ $Y2=0
cc_317 N_A_27_424#_c_360_n N_VPWR_M1011_d 0.00762644f $X=2.525 $Y=2.475
+ $X2=-0.19 $Y2=-0.245
cc_318 N_A_27_424#_c_363_n N_VPWR_M1011_d 0.00452151f $X=0.715 $Y=2.33 $X2=-0.19
+ $Y2=-0.245
cc_319 N_A_27_424#_c_360_n N_VPWR_M1015_d 0.0119854f $X=2.525 $Y=2.475 $X2=0
+ $Y2=0
cc_320 N_A_27_424#_c_361_n N_VPWR_M1015_d 0.00516029f $X=2.61 $Y=2.39 $X2=0
+ $Y2=0
cc_321 N_A_27_424#_c_362_n N_VPWR_c_783_n 0.0101711f $X=0.28 $Y=2.265 $X2=0
+ $Y2=0
cc_322 N_A_27_424#_c_363_n N_VPWR_c_783_n 0.0200525f $X=0.715 $Y=2.33 $X2=0
+ $Y2=0
cc_323 N_A_27_424#_c_354_n N_VPWR_c_784_n 0.00721133f $X=2.765 $Y=1.885 $X2=0
+ $Y2=0
cc_324 N_A_27_424#_c_360_n N_VPWR_c_784_n 0.0250318f $X=2.525 $Y=2.475 $X2=0
+ $Y2=0
cc_325 N_A_27_424#_c_362_n N_VPWR_c_788_n 0.0140991f $X=0.28 $Y=2.265 $X2=0
+ $Y2=0
cc_326 N_A_27_424#_c_354_n N_VPWR_c_790_n 0.00413917f $X=2.765 $Y=1.885 $X2=0
+ $Y2=0
cc_327 N_A_27_424#_c_354_n N_VPWR_c_782_n 0.00817532f $X=2.765 $Y=1.885 $X2=0
+ $Y2=0
cc_328 N_A_27_424#_c_360_n N_VPWR_c_782_n 0.0508607f $X=2.525 $Y=2.475 $X2=0
+ $Y2=0
cc_329 N_A_27_424#_c_362_n N_VPWR_c_782_n 0.0118561f $X=0.28 $Y=2.265 $X2=0
+ $Y2=0
cc_330 N_A_27_424#_c_363_n N_VPWR_c_782_n 0.00713309f $X=0.715 $Y=2.33 $X2=0
+ $Y2=0
cc_331 N_A_27_424#_c_356_n N_VGND_c_886_n 0.0230738f $X=0.63 $Y=0.835 $X2=0
+ $Y2=0
cc_332 N_A_27_424#_M1017_g N_VGND_c_887_n 0.00507404f $X=2.75 $Y=0.69 $X2=0
+ $Y2=0
cc_333 N_A_27_424#_c_356_n N_VGND_c_890_n 0.0118661f $X=0.63 $Y=0.835 $X2=0
+ $Y2=0
cc_334 N_A_27_424#_M1017_g N_VGND_c_892_n 0.00444681f $X=2.75 $Y=0.69 $X2=0
+ $Y2=0
cc_335 N_A_27_424#_M1017_g N_VGND_c_898_n 0.00427328f $X=2.75 $Y=0.69 $X2=0
+ $Y2=0
cc_336 N_A_27_424#_c_356_n N_VGND_c_898_n 0.0158184f $X=0.63 $Y=0.835 $X2=0
+ $Y2=0
cc_337 N_A_363_74#_c_451_n N_A_817_48#_c_567_n 0.0295462f $X=3.72 $Y=2.465 $X2=0
+ $Y2=0
cc_338 N_A_363_74#_c_454_n N_A_817_48#_c_567_n 0.00173515f $X=3.715 $Y=2.99
+ $X2=0 $Y2=0
cc_339 N_A_363_74#_c_456_n N_A_817_48#_c_567_n 0.00943145f $X=3.88 $Y=2.215
+ $X2=0 $Y2=0
cc_340 N_A_363_74#_c_451_n N_A_817_48#_c_570_n 0.00120301f $X=3.72 $Y=2.465
+ $X2=0 $Y2=0
cc_341 N_A_363_74#_c_456_n N_A_817_48#_c_570_n 0.0177637f $X=3.88 $Y=2.215 $X2=0
+ $Y2=0
cc_342 N_A_363_74#_c_454_n N_A_643_74#_M1001_d 0.00444187f $X=3.715 $Y=2.99
+ $X2=0 $Y2=0
cc_343 N_A_363_74#_c_447_n N_A_643_74#_c_666_n 0.0136696f $X=3.11 $Y=1.97 $X2=0
+ $Y2=0
cc_344 N_A_363_74#_c_448_n N_A_643_74#_c_666_n 0.0254068f $X=3.175 $Y=1.195
+ $X2=0 $Y2=0
cc_345 N_A_363_74#_c_449_n N_A_643_74#_c_666_n 0.00244597f $X=3.23 $Y=1.285
+ $X2=0 $Y2=0
cc_346 N_A_363_74#_c_450_n N_A_643_74#_c_666_n 0.00351644f $X=3.23 $Y=1.12 $X2=0
+ $Y2=0
cc_347 N_A_363_74#_c_456_n N_A_643_74#_c_673_n 0.0262119f $X=3.88 $Y=2.215 $X2=0
+ $Y2=0
cc_348 N_A_363_74#_c_451_n N_A_643_74#_c_674_n 0.0043573f $X=3.72 $Y=2.465 $X2=0
+ $Y2=0
cc_349 N_A_363_74#_c_447_n N_A_643_74#_c_674_n 0.0130064f $X=3.11 $Y=1.97 $X2=0
+ $Y2=0
cc_350 N_A_363_74#_c_448_n N_A_643_74#_c_667_n 0.00806711f $X=3.175 $Y=1.195
+ $X2=0 $Y2=0
cc_351 N_A_363_74#_c_449_n N_A_643_74#_c_667_n 0.00341895f $X=3.23 $Y=1.285
+ $X2=0 $Y2=0
cc_352 N_A_363_74#_c_450_n N_A_643_74#_c_667_n 0.00935059f $X=3.23 $Y=1.12 $X2=0
+ $Y2=0
cc_353 N_A_363_74#_c_451_n N_A_643_74#_c_689_n 0.00213143f $X=3.72 $Y=2.465
+ $X2=0 $Y2=0
cc_354 N_A_363_74#_c_454_n N_A_643_74#_c_689_n 0.017233f $X=3.715 $Y=2.99 $X2=0
+ $Y2=0
cc_355 N_A_363_74#_c_451_n N_A_643_74#_c_675_n 0.00387176f $X=3.72 $Y=2.465
+ $X2=0 $Y2=0
cc_356 N_A_363_74#_c_447_n N_A_643_74#_c_675_n 0.00535072f $X=3.11 $Y=1.97 $X2=0
+ $Y2=0
cc_357 N_A_363_74#_c_456_n N_A_643_74#_c_675_n 0.0482168f $X=3.88 $Y=2.215 $X2=0
+ $Y2=0
cc_358 N_A_363_74#_c_489_n N_A_643_74#_c_675_n 0.0123438f $X=3.11 $Y=2.055 $X2=0
+ $Y2=0
cc_359 N_A_363_74#_c_503_n N_VPWR_c_784_n 0.0114807f $X=2.99 $Y=2.905 $X2=0
+ $Y2=0
cc_360 N_A_363_74#_c_455_n N_VPWR_c_784_n 0.0126996f $X=3.075 $Y=2.99 $X2=0
+ $Y2=0
cc_361 N_A_363_74#_c_451_n N_VPWR_c_790_n 0.00278193f $X=3.72 $Y=2.465 $X2=0
+ $Y2=0
cc_362 N_A_363_74#_c_454_n N_VPWR_c_790_n 0.0638747f $X=3.715 $Y=2.99 $X2=0
+ $Y2=0
cc_363 N_A_363_74#_c_455_n N_VPWR_c_790_n 0.0121867f $X=3.075 $Y=2.99 $X2=0
+ $Y2=0
cc_364 N_A_363_74#_c_451_n N_VPWR_c_782_n 0.00356236f $X=3.72 $Y=2.465 $X2=0
+ $Y2=0
cc_365 N_A_363_74#_c_454_n N_VPWR_c_782_n 0.0355129f $X=3.715 $Y=2.99 $X2=0
+ $Y2=0
cc_366 N_A_363_74#_c_455_n N_VPWR_c_782_n 0.00660921f $X=3.075 $Y=2.99 $X2=0
+ $Y2=0
cc_367 N_A_363_74#_c_451_n N_VPWR_c_795_n 4.04476e-19 $X=3.72 $Y=2.465 $X2=0
+ $Y2=0
cc_368 N_A_363_74#_c_454_n N_VPWR_c_795_n 0.00796977f $X=3.715 $Y=2.99 $X2=0
+ $Y2=0
cc_369 N_A_363_74#_c_456_n N_VPWR_c_795_n 0.0109526f $X=3.88 $Y=2.215 $X2=0
+ $Y2=0
cc_370 N_A_363_74#_c_503_n A_568_392# 0.0112933f $X=2.99 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_371 N_A_363_74#_c_455_n A_568_392# 5.72894e-19 $X=3.075 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_372 N_A_363_74#_c_489_n A_568_392# 0.00678783f $X=3.11 $Y=2.055 $X2=-0.19
+ $Y2=-0.245
cc_373 N_A_363_74#_c_454_n A_759_508# 9.16612e-19 $X=3.715 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_374 N_A_363_74#_c_456_n A_759_508# 0.00589473f $X=3.88 $Y=2.215 $X2=-0.19
+ $Y2=-0.245
cc_375 N_A_363_74#_c_450_n N_VGND_c_887_n 2.63324e-19 $X=3.23 $Y=1.12 $X2=0
+ $Y2=0
cc_376 N_A_363_74#_c_450_n N_VGND_c_892_n 0.00278271f $X=3.23 $Y=1.12 $X2=0
+ $Y2=0
cc_377 N_A_363_74#_c_450_n N_VGND_c_898_n 0.00354802f $X=3.23 $Y=1.12 $X2=0
+ $Y2=0
cc_378 N_A_817_48#_c_567_n N_A_643_74#_c_669_n 0.0209772f $X=4.375 $Y=2.465
+ $X2=0 $Y2=0
cc_379 N_A_817_48#_c_558_n N_A_643_74#_c_669_n 0.00324263f $X=4.38 $Y=2.05 $X2=0
+ $Y2=0
cc_380 N_A_817_48#_c_570_n N_A_643_74#_c_669_n 0.00985012f $X=5.095 $Y=2.222
+ $X2=0 $Y2=0
cc_381 N_A_817_48#_c_571_n N_A_643_74#_c_669_n 0.00325694f $X=5.41 $Y=2.465
+ $X2=0 $Y2=0
cc_382 N_A_817_48#_c_572_n N_A_643_74#_c_669_n 0.0197382f $X=5.41 $Y=2.115 $X2=0
+ $Y2=0
cc_383 N_A_817_48#_c_566_n N_A_643_74#_c_669_n 0.00206502f $X=5.335 $Y=1.95
+ $X2=0 $Y2=0
cc_384 N_A_817_48#_c_561_n N_A_643_74#_M1014_g 0.00808109f $X=4.38 $Y=0.94 $X2=0
+ $Y2=0
cc_385 N_A_817_48#_c_562_n N_A_643_74#_M1014_g 0.012954f $X=4.935 $Y=0.515 $X2=0
+ $Y2=0
cc_386 N_A_817_48#_c_565_n N_A_643_74#_M1014_g 0.0127642f $X=5.017 $Y=1.095
+ $X2=0 $Y2=0
cc_387 N_A_817_48#_c_566_n N_A_643_74#_M1014_g 0.009378f $X=5.335 $Y=1.95 $X2=0
+ $Y2=0
cc_388 N_A_817_48#_c_558_n N_A_643_74#_c_664_n 0.0217577f $X=4.38 $Y=2.05 $X2=0
+ $Y2=0
cc_389 N_A_817_48#_c_570_n N_A_643_74#_c_664_n 0.00511011f $X=5.095 $Y=2.222
+ $X2=0 $Y2=0
cc_390 N_A_817_48#_c_565_n N_A_643_74#_c_664_n 0.00709268f $X=5.017 $Y=1.095
+ $X2=0 $Y2=0
cc_391 N_A_817_48#_c_558_n N_A_643_74#_c_665_n 0.00108219f $X=4.38 $Y=2.05 $X2=0
+ $Y2=0
cc_392 N_A_817_48#_c_566_n N_A_643_74#_c_665_n 0.0118583f $X=5.335 $Y=1.95 $X2=0
+ $Y2=0
cc_393 N_A_817_48#_c_567_n N_A_643_74#_c_673_n 0.00474613f $X=4.375 $Y=2.465
+ $X2=0 $Y2=0
cc_394 N_A_817_48#_c_558_n N_A_643_74#_c_673_n 0.01626f $X=4.38 $Y=2.05 $X2=0
+ $Y2=0
cc_395 N_A_817_48#_c_570_n N_A_643_74#_c_673_n 0.0265217f $X=5.095 $Y=2.222
+ $X2=0 $Y2=0
cc_396 N_A_817_48#_c_558_n N_A_643_74#_c_668_n 0.00167293f $X=4.38 $Y=2.05 $X2=0
+ $Y2=0
cc_397 N_A_817_48#_c_570_n N_A_643_74#_c_668_n 0.0217299f $X=5.095 $Y=2.222
+ $X2=0 $Y2=0
cc_398 N_A_817_48#_c_565_n N_A_643_74#_c_668_n 0.00890275f $X=5.017 $Y=1.095
+ $X2=0 $Y2=0
cc_399 N_A_817_48#_c_566_n N_A_643_74#_c_668_n 0.0301206f $X=5.335 $Y=1.95 $X2=0
+ $Y2=0
cc_400 N_A_817_48#_c_559_n N_RESET_B_M1003_g 0.0290173f $X=6.05 $Y=1.22 $X2=0
+ $Y2=0
cc_401 N_A_817_48#_c_562_n N_RESET_B_M1003_g 0.00222669f $X=4.935 $Y=0.515 $X2=0
+ $Y2=0
cc_402 N_A_817_48#_c_563_n N_RESET_B_M1003_g 0.0144185f $X=5.975 $Y=1.095 $X2=0
+ $Y2=0
cc_403 N_A_817_48#_c_564_n N_RESET_B_M1003_g 9.9568e-19 $X=6.14 $Y=1.385 $X2=0
+ $Y2=0
cc_404 N_A_817_48#_c_566_n N_RESET_B_M1003_g 0.00330038f $X=5.335 $Y=1.95 $X2=0
+ $Y2=0
cc_405 N_A_817_48#_c_560_n N_RESET_B_c_747_n 0.0458717f $X=6.215 $Y=1.765 $X2=0
+ $Y2=0
cc_406 N_A_817_48#_c_571_n N_RESET_B_c_747_n 0.00614465f $X=5.41 $Y=2.465 $X2=0
+ $Y2=0
cc_407 N_A_817_48#_c_563_n N_RESET_B_c_747_n 0.00124498f $X=5.975 $Y=1.095 $X2=0
+ $Y2=0
cc_408 N_A_817_48#_c_564_n N_RESET_B_c_747_n 6.9668e-19 $X=6.14 $Y=1.385 $X2=0
+ $Y2=0
cc_409 N_A_817_48#_c_572_n N_RESET_B_c_747_n 0.00560137f $X=5.41 $Y=2.115 $X2=0
+ $Y2=0
cc_410 N_A_817_48#_c_566_n N_RESET_B_c_747_n 0.00512023f $X=5.335 $Y=1.95 $X2=0
+ $Y2=0
cc_411 N_A_817_48#_c_560_n N_RESET_B_c_748_n 0.00345786f $X=6.215 $Y=1.765 $X2=0
+ $Y2=0
cc_412 N_A_817_48#_c_563_n N_RESET_B_c_748_n 0.0247205f $X=5.975 $Y=1.095 $X2=0
+ $Y2=0
cc_413 N_A_817_48#_c_564_n N_RESET_B_c_748_n 0.0126449f $X=6.14 $Y=1.385 $X2=0
+ $Y2=0
cc_414 N_A_817_48#_c_572_n N_RESET_B_c_748_n 0.0123116f $X=5.41 $Y=2.115 $X2=0
+ $Y2=0
cc_415 N_A_817_48#_c_566_n N_RESET_B_c_748_n 0.0327282f $X=5.335 $Y=1.95 $X2=0
+ $Y2=0
cc_416 N_A_817_48#_c_570_n N_VPWR_M1005_d 0.0061068f $X=5.095 $Y=2.222 $X2=0
+ $Y2=0
cc_417 N_A_817_48#_c_560_n N_VPWR_c_785_n 0.0137142f $X=6.215 $Y=1.765 $X2=0
+ $Y2=0
cc_418 N_A_817_48#_c_564_n N_VPWR_c_785_n 0.00434026f $X=6.14 $Y=1.385 $X2=0
+ $Y2=0
cc_419 N_A_817_48#_c_572_n N_VPWR_c_785_n 0.0407271f $X=5.41 $Y=2.115 $X2=0
+ $Y2=0
cc_420 N_A_817_48#_c_571_n N_VPWR_c_786_n 0.0145938f $X=5.41 $Y=2.465 $X2=0
+ $Y2=0
cc_421 N_A_817_48#_c_567_n N_VPWR_c_790_n 0.00415318f $X=4.375 $Y=2.465 $X2=0
+ $Y2=0
cc_422 N_A_817_48#_c_560_n N_VPWR_c_791_n 0.00445602f $X=6.215 $Y=1.765 $X2=0
+ $Y2=0
cc_423 N_A_817_48#_c_567_n N_VPWR_c_782_n 0.00851322f $X=4.375 $Y=2.465 $X2=0
+ $Y2=0
cc_424 N_A_817_48#_c_560_n N_VPWR_c_782_n 0.00862211f $X=6.215 $Y=1.765 $X2=0
+ $Y2=0
cc_425 N_A_817_48#_c_571_n N_VPWR_c_782_n 0.0120466f $X=5.41 $Y=2.465 $X2=0
+ $Y2=0
cc_426 N_A_817_48#_c_567_n N_VPWR_c_795_n 0.0193947f $X=4.375 $Y=2.465 $X2=0
+ $Y2=0
cc_427 N_A_817_48#_c_570_n N_VPWR_c_795_n 0.0328403f $X=5.095 $Y=2.222 $X2=0
+ $Y2=0
cc_428 N_A_817_48#_c_571_n N_VPWR_c_795_n 0.0144922f $X=5.41 $Y=2.465 $X2=0
+ $Y2=0
cc_429 N_A_817_48#_c_563_n N_Q_M1013_d 0.00234008f $X=5.975 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_430 N_A_817_48#_c_560_n N_Q_c_865_n 0.0117221f $X=6.215 $Y=1.765 $X2=0 $Y2=0
cc_431 N_A_817_48#_c_560_n N_Q_c_866_n 0.0044665f $X=6.215 $Y=1.765 $X2=0 $Y2=0
cc_432 N_A_817_48#_c_564_n N_Q_c_866_n 0.00104962f $X=6.14 $Y=1.385 $X2=0 $Y2=0
cc_433 N_A_817_48#_c_559_n N_Q_c_863_n 0.00443182f $X=6.05 $Y=1.22 $X2=0 $Y2=0
cc_434 N_A_817_48#_c_560_n N_Q_c_863_n 0.0152363f $X=6.215 $Y=1.765 $X2=0 $Y2=0
cc_435 N_A_817_48#_c_563_n N_Q_c_863_n 0.0141806f $X=5.975 $Y=1.095 $X2=0 $Y2=0
cc_436 N_A_817_48#_c_564_n N_Q_c_863_n 0.0278652f $X=6.14 $Y=1.385 $X2=0 $Y2=0
cc_437 N_A_817_48#_c_559_n Q 0.00864397f $X=6.05 $Y=1.22 $X2=0 $Y2=0
cc_438 N_A_817_48#_c_560_n Q 0.00106205f $X=6.215 $Y=1.765 $X2=0 $Y2=0
cc_439 N_A_817_48#_c_563_n Q 0.0116838f $X=5.975 $Y=1.095 $X2=0 $Y2=0
cc_440 N_A_817_48#_c_563_n N_VGND_M1003_d 0.00261503f $X=5.975 $Y=1.095 $X2=0
+ $Y2=0
cc_441 N_A_817_48#_c_557_n N_VGND_c_888_n 0.0115327f $X=4.16 $Y=0.865 $X2=0
+ $Y2=0
cc_442 N_A_817_48#_c_561_n N_VGND_c_888_n 0.01149f $X=4.38 $Y=0.94 $X2=0 $Y2=0
cc_443 N_A_817_48#_c_562_n N_VGND_c_888_n 0.0310125f $X=4.935 $Y=0.515 $X2=0
+ $Y2=0
cc_444 N_A_817_48#_c_559_n N_VGND_c_889_n 0.00569497f $X=6.05 $Y=1.22 $X2=0
+ $Y2=0
cc_445 N_A_817_48#_c_562_n N_VGND_c_889_n 0.0155235f $X=4.935 $Y=0.515 $X2=0
+ $Y2=0
cc_446 N_A_817_48#_c_563_n N_VGND_c_889_n 0.0218003f $X=5.975 $Y=1.095 $X2=0
+ $Y2=0
cc_447 N_A_817_48#_c_557_n N_VGND_c_892_n 0.00383152f $X=4.16 $Y=0.865 $X2=0
+ $Y2=0
cc_448 N_A_817_48#_c_562_n N_VGND_c_894_n 0.0145639f $X=4.935 $Y=0.515 $X2=0
+ $Y2=0
cc_449 N_A_817_48#_c_559_n N_VGND_c_897_n 0.00434272f $X=6.05 $Y=1.22 $X2=0
+ $Y2=0
cc_450 N_A_817_48#_c_557_n N_VGND_c_898_n 0.0075725f $X=4.16 $Y=0.865 $X2=0
+ $Y2=0
cc_451 N_A_817_48#_c_559_n N_VGND_c_898_n 0.00825201f $X=6.05 $Y=1.22 $X2=0
+ $Y2=0
cc_452 N_A_817_48#_c_562_n N_VGND_c_898_n 0.0119984f $X=4.935 $Y=0.515 $X2=0
+ $Y2=0
cc_453 N_A_817_48#_c_563_n A_1045_74# 0.0048076f $X=5.975 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_454 N_A_643_74#_M1014_g N_RESET_B_M1003_g 0.0564763f $X=5.15 $Y=0.74 $X2=0
+ $Y2=0
cc_455 N_A_643_74#_c_669_n N_RESET_B_c_747_n 0.0207328f $X=5.135 $Y=1.885 $X2=0
+ $Y2=0
cc_456 N_A_643_74#_M1014_g N_RESET_B_c_747_n 0.020603f $X=5.15 $Y=0.74 $X2=0
+ $Y2=0
cc_457 N_A_643_74#_c_665_n N_RESET_B_c_747_n 0.00751679f $X=5.135 $Y=1.677 $X2=0
+ $Y2=0
cc_458 N_A_643_74#_M1014_g N_RESET_B_c_748_n 3.79805e-19 $X=5.15 $Y=0.74 $X2=0
+ $Y2=0
cc_459 N_A_643_74#_c_665_n N_RESET_B_c_748_n 3.27182e-19 $X=5.135 $Y=1.677 $X2=0
+ $Y2=0
cc_460 N_A_643_74#_c_669_n N_VPWR_c_786_n 0.00415318f $X=5.135 $Y=1.885 $X2=0
+ $Y2=0
cc_461 N_A_643_74#_c_669_n N_VPWR_c_782_n 0.00818241f $X=5.135 $Y=1.885 $X2=0
+ $Y2=0
cc_462 N_A_643_74#_c_669_n N_VPWR_c_795_n 0.0143972f $X=5.135 $Y=1.885 $X2=0
+ $Y2=0
cc_463 N_A_643_74#_M1014_g N_VGND_c_888_n 0.00370782f $X=5.15 $Y=0.74 $X2=0
+ $Y2=0
cc_464 N_A_643_74#_M1014_g N_VGND_c_889_n 0.00194806f $X=5.15 $Y=0.74 $X2=0
+ $Y2=0
cc_465 N_A_643_74#_M1014_g N_VGND_c_894_n 0.00434272f $X=5.15 $Y=0.74 $X2=0
+ $Y2=0
cc_466 N_A_643_74#_M1014_g N_VGND_c_898_n 0.00825979f $X=5.15 $Y=0.74 $X2=0
+ $Y2=0
cc_467 N_RESET_B_c_747_n N_VPWR_c_785_n 0.00856778f $X=5.635 $Y=1.885 $X2=0
+ $Y2=0
cc_468 N_RESET_B_c_748_n N_VPWR_c_785_n 0.00163024f $X=5.6 $Y=1.515 $X2=0 $Y2=0
cc_469 N_RESET_B_c_747_n N_VPWR_c_786_n 0.00445602f $X=5.635 $Y=1.885 $X2=0
+ $Y2=0
cc_470 N_RESET_B_c_747_n N_VPWR_c_782_n 0.00858558f $X=5.635 $Y=1.885 $X2=0
+ $Y2=0
cc_471 N_RESET_B_c_747_n N_VPWR_c_795_n 4.22856e-19 $X=5.635 $Y=1.885 $X2=0
+ $Y2=0
cc_472 N_RESET_B_c_747_n N_Q_c_866_n 8.13355e-19 $X=5.635 $Y=1.885 $X2=0 $Y2=0
cc_473 N_RESET_B_M1003_g N_VGND_c_889_n 0.0138667f $X=5.54 $Y=0.74 $X2=0 $Y2=0
cc_474 N_RESET_B_M1003_g N_VGND_c_894_n 0.00383152f $X=5.54 $Y=0.74 $X2=0 $Y2=0
cc_475 N_RESET_B_M1003_g N_VGND_c_898_n 0.0075725f $X=5.54 $Y=0.74 $X2=0 $Y2=0
cc_476 N_VPWR_c_791_n N_Q_c_865_n 0.0159324f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_477 N_VPWR_c_782_n N_Q_c_865_n 0.0131546f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_478 N_VPWR_c_785_n N_Q_c_866_n 0.0710027f $X=5.91 $Y=2.115 $X2=0 $Y2=0
cc_479 Q N_VGND_c_889_n 0.0196681f $X=6.395 $Y=0.47 $X2=0 $Y2=0
cc_480 Q N_VGND_c_897_n 0.0233346f $X=6.395 $Y=0.47 $X2=0 $Y2=0
cc_481 Q N_VGND_c_898_n 0.0194239f $X=6.395 $Y=0.47 $X2=0 $Y2=0
