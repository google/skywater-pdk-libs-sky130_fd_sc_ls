* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__a222o_2 A1 A2 B1 B2 C1 C2 VGND VNB VPB VPWR X
M1000 X a_27_82# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=1.16865e+12p ps=9.01e+06u
M1001 a_114_82# C1 a_27_82# VNB nshort w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=4.832e+11p ps=4.07e+06u
M1002 X a_27_82# VGND VNB nshort w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=9.428e+11p ps=7.49e+06u
M1003 a_27_82# A1 a_557_74# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=3.795e+11p ps=3.77e+06u
M1004 VPWR a_27_82# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_116_392# B1 a_639_368# VPB phighvt w=1e+06u l=150000u
+  ad=6e+11p pd=5.2e+06u as=9.635e+11p ps=6.17e+06u
M1006 VGND a_27_82# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND B2 a_775_74# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=1.536e+11p ps=1.76e+06u
M1008 a_639_368# A1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_775_74# B1 a_27_82# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_639_368# B2 a_116_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND C2 a_114_82# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_27_82# C2 a_116_392# VPB phighvt w=1e+06u l=150000u
+  ad=5.9e+11p pd=5.18e+06u as=0p ps=0u
M1013 a_116_392# C1 a_27_82# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR A2 a_639_368# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_557_74# A2 VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
