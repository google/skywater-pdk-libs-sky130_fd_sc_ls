* File: sky130_fd_sc_ls__o311a_4.pxi.spice
* Created: Fri Aug 28 13:51:41 2020
* 
x_PM_SKY130_FD_SC_LS__O311A_4%A_83_244# N_A_83_244#_M1008_d N_A_83_244#_M1011_s
+ N_A_83_244#_M1015_d N_A_83_244#_M1000_d N_A_83_244#_c_158_n
+ N_A_83_244#_M1009_g N_A_83_244#_c_148_n N_A_83_244#_M1004_g
+ N_A_83_244#_c_159_n N_A_83_244#_M1010_g N_A_83_244#_c_149_n
+ N_A_83_244#_M1005_g N_A_83_244#_c_160_n N_A_83_244#_M1013_g
+ N_A_83_244#_c_150_n N_A_83_244#_M1021_g N_A_83_244#_c_161_n
+ N_A_83_244#_M1019_g N_A_83_244#_c_151_n N_A_83_244#_M1026_g
+ N_A_83_244#_c_288_p N_A_83_244#_c_152_n N_A_83_244#_c_153_n
+ N_A_83_244#_c_163_n N_A_83_244#_c_242_p N_A_83_244#_c_164_n
+ N_A_83_244#_c_165_n N_A_83_244#_c_166_n N_A_83_244#_c_167_n
+ N_A_83_244#_c_154_n N_A_83_244#_c_155_n N_A_83_244#_c_156_n
+ N_A_83_244#_c_170_n N_A_83_244#_c_171_n N_A_83_244#_c_157_n
+ N_A_83_244#_c_172_n PM_SKY130_FD_SC_LS__O311A_4%A_83_244#
x_PM_SKY130_FD_SC_LS__O311A_4%B1 N_B1_c_337_n N_B1_c_349_n N_B1_M1011_g
+ N_B1_c_338_n N_B1_M1003_g N_B1_c_350_n N_B1_M1022_g N_B1_c_351_n N_B1_c_352_n
+ N_B1_M1024_g N_B1_c_341_n N_B1_c_342_n N_B1_c_343_n N_B1_c_381_n B1
+ N_B1_c_344_n N_B1_c_345_n N_B1_c_346_n N_B1_c_347_n
+ PM_SKY130_FD_SC_LS__O311A_4%B1
x_PM_SKY130_FD_SC_LS__O311A_4%C1 N_C1_c_454_n N_C1_M1007_g N_C1_c_447_n
+ N_C1_c_456_n N_C1_M1015_g N_C1_M1008_g N_C1_c_449_n N_C1_c_450_n N_C1_M1017_g
+ N_C1_c_452_n C1 PM_SKY130_FD_SC_LS__O311A_4%C1
x_PM_SKY130_FD_SC_LS__O311A_4%A3 N_A3_M1012_g N_A3_c_524_n N_A3_M1000_g
+ N_A3_c_525_n N_A3_M1023_g N_A3_M1018_g A3 N_A3_c_523_n
+ PM_SKY130_FD_SC_LS__O311A_4%A3
x_PM_SKY130_FD_SC_LS__O311A_4%A2 N_A2_c_579_n N_A2_c_590_n N_A2_M1001_g
+ N_A2_M1006_g N_A2_c_581_n N_A2_c_592_n N_A2_M1020_g N_A2_c_582_n N_A2_M1014_g
+ N_A2_c_583_n N_A2_c_584_n N_A2_c_585_n A2 A2 N_A2_c_587_n N_A2_c_588_n
+ PM_SKY130_FD_SC_LS__O311A_4%A2
x_PM_SKY130_FD_SC_LS__O311A_4%A1 N_A1_M1002_g N_A1_c_662_n N_A1_M1016_g
+ N_A1_c_663_n N_A1_M1027_g N_A1_M1025_g A1 A1 N_A1_c_661_n
+ PM_SKY130_FD_SC_LS__O311A_4%A1
x_PM_SKY130_FD_SC_LS__O311A_4%VPWR N_VPWR_M1009_s N_VPWR_M1010_s N_VPWR_M1019_s
+ N_VPWR_M1007_s N_VPWR_M1022_d N_VPWR_M1016_d N_VPWR_c_717_n N_VPWR_c_718_n
+ N_VPWR_c_719_n N_VPWR_c_720_n N_VPWR_c_721_n N_VPWR_c_722_n N_VPWR_c_723_n
+ N_VPWR_c_724_n N_VPWR_c_795_n N_VPWR_c_725_n N_VPWR_c_726_n N_VPWR_c_727_n
+ N_VPWR_c_760_n VPWR N_VPWR_c_728_n N_VPWR_c_729_n N_VPWR_c_730_n
+ N_VPWR_c_716_n N_VPWR_c_732_n N_VPWR_c_733_n N_VPWR_c_734_n
+ PM_SKY130_FD_SC_LS__O311A_4%VPWR
x_PM_SKY130_FD_SC_LS__O311A_4%X N_X_M1004_d N_X_M1021_d N_X_M1009_d N_X_M1013_d
+ N_X_c_843_n N_X_c_844_n N_X_c_845_n N_X_c_850_n N_X_c_846_n N_X_c_851_n
+ N_X_c_868_n N_X_c_852_n N_X_c_847_n N_X_c_877_n N_X_c_882_n X N_X_c_849_n
+ PM_SKY130_FD_SC_LS__O311A_4%X
x_PM_SKY130_FD_SC_LS__O311A_4%A_1034_392# N_A_1034_392#_M1000_s
+ N_A_1034_392#_M1023_s N_A_1034_392#_M1020_s N_A_1034_392#_c_912_n
+ N_A_1034_392#_c_913_n N_A_1034_392#_c_914_n N_A_1034_392#_c_915_n
+ PM_SKY130_FD_SC_LS__O311A_4%A_1034_392#
x_PM_SKY130_FD_SC_LS__O311A_4%A_1338_392# N_A_1338_392#_M1001_d
+ N_A_1338_392#_M1027_s N_A_1338_392#_c_948_n N_A_1338_392#_c_950_n
+ PM_SKY130_FD_SC_LS__O311A_4%A_1338_392#
x_PM_SKY130_FD_SC_LS__O311A_4%VGND N_VGND_M1004_s N_VGND_M1005_s N_VGND_M1026_s
+ N_VGND_M1012_s N_VGND_M1006_s N_VGND_M1025_s N_VGND_c_959_n N_VGND_c_960_n
+ N_VGND_c_961_n N_VGND_c_962_n N_VGND_c_963_n N_VGND_c_964_n N_VGND_c_965_n
+ N_VGND_c_966_n N_VGND_c_967_n VGND N_VGND_c_968_n N_VGND_c_969_n
+ N_VGND_c_970_n N_VGND_c_971_n N_VGND_c_972_n N_VGND_c_973_n N_VGND_c_974_n
+ N_VGND_c_975_n N_VGND_c_976_n N_VGND_c_977_n PM_SKY130_FD_SC_LS__O311A_4%VGND
x_PM_SKY130_FD_SC_LS__O311A_4%A_564_78# N_A_564_78#_M1003_s N_A_564_78#_M1024_s
+ N_A_564_78#_M1018_d N_A_564_78#_M1002_d N_A_564_78#_M1014_d
+ N_A_564_78#_c_1058_n N_A_564_78#_c_1059_n N_A_564_78#_c_1060_n
+ N_A_564_78#_c_1068_n N_A_564_78#_c_1069_n N_A_564_78#_c_1061_n
+ N_A_564_78#_c_1090_n N_A_564_78#_c_1062_n N_A_564_78#_c_1094_n
+ N_A_564_78#_c_1063_n N_A_564_78#_c_1064_n N_A_564_78#_c_1065_n
+ N_A_564_78#_c_1103_n PM_SKY130_FD_SC_LS__O311A_4%A_564_78#
x_PM_SKY130_FD_SC_LS__O311A_4%A_651_78# N_A_651_78#_M1003_d N_A_651_78#_M1017_s
+ N_A_651_78#_c_1141_n N_A_651_78#_c_1146_n N_A_651_78#_c_1147_n
+ N_A_651_78#_c_1144_n PM_SKY130_FD_SC_LS__O311A_4%A_651_78#
cc_1 VNB N_A_83_244#_c_148_n 0.0190025f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.22
cc_2 VNB N_A_83_244#_c_149_n 0.0186851f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.22
cc_3 VNB N_A_83_244#_c_150_n 0.0197981f $X=-0.19 $Y=-0.245 $X2=1.69 $Y2=1.22
cc_4 VNB N_A_83_244#_c_151_n 0.0202546f $X=-0.19 $Y=-0.245 $X2=2.19 $Y2=1.22
cc_5 VNB N_A_83_244#_c_152_n 0.00234403f $X=-0.19 $Y=-0.245 $X2=2.18 $Y2=1.55
cc_6 VNB N_A_83_244#_c_153_n 0.00110322f $X=-0.19 $Y=-0.245 $X2=2.18 $Y2=1.72
cc_7 VNB N_A_83_244#_c_154_n 0.0140254f $X=-0.19 $Y=-0.245 $X2=5.53 $Y2=1.215
cc_8 VNB N_A_83_244#_c_155_n 0.00295206f $X=-0.19 $Y=-0.245 $X2=5.615 $Y2=1.95
cc_9 VNB N_A_83_244#_c_156_n 0.137576f $X=-0.19 $Y=-0.245 $X2=2.1 $Y2=1.385
cc_10 VNB N_A_83_244#_c_157_n 0.00329916f $X=-0.19 $Y=-0.245 $X2=4.42 $Y2=1.1
cc_11 VNB N_B1_c_337_n 0.00845064f $X=-0.19 $Y=-0.245 $X2=2.67 $Y2=1.96
cc_12 VNB N_B1_c_338_n 0.0295471f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_B1_M1003_g 0.0296011f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_B1_M1024_g 0.0336185f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.765
cc_15 VNB N_B1_c_341_n 0.0178364f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_16 VNB N_B1_c_342_n 0.0190135f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.22
cc_17 VNB N_B1_c_343_n 0.00185509f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_18 VNB N_B1_c_344_n 0.0332696f $X=-0.19 $Y=-0.245 $X2=2.09 $Y2=2.4
cc_19 VNB N_B1_c_345_n 0.0186746f $X=-0.19 $Y=-0.245 $X2=1.42 $Y2=1.385
cc_20 VNB N_B1_c_346_n 0.00294754f $X=-0.19 $Y=-0.245 $X2=1.42 $Y2=1.385
cc_21 VNB N_B1_c_347_n 0.0136793f $X=-0.19 $Y=-0.245 $X2=2.655 $Y2=1.805
cc_22 VNB N_C1_c_447_n 0.00717907f $X=-0.19 $Y=-0.245 $X2=5.765 $Y2=1.96
cc_23 VNB N_C1_M1008_g 0.0330506f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_C1_c_449_n 0.0298624f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_25 VNB N_C1_c_450_n 0.0523893f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_26 VNB N_C1_M1017_g 0.0255349f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.74
cc_27 VNB N_C1_c_452_n 0.00526697f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.765
cc_28 VNB C1 0.00394353f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_29 VNB N_A3_M1012_g 0.0333241f $X=-0.19 $Y=-0.245 $X2=4.105 $Y2=1.96
cc_30 VNB N_A3_M1018_g 0.0326426f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_31 VNB A3 0.00245697f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_32 VNB N_A3_c_523_n 0.0324948f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.22
cc_33 VNB N_A2_c_579_n 0.00663167f $X=-0.19 $Y=-0.245 $X2=2.67 $Y2=1.96
cc_34 VNB N_A2_M1006_g 0.0219897f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A2_c_581_n 0.00517465f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A2_c_582_n 0.0217296f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_37 VNB N_A2_c_583_n 0.0157023f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.74
cc_38 VNB N_A2_c_584_n 0.0121784f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.765
cc_39 VNB N_A2_c_585_n 0.0286154f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_40 VNB A2 0.00829845f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_41 VNB N_A2_c_587_n 0.0610218f $X=-0.19 $Y=-0.245 $X2=2.09 $Y2=2.4
cc_42 VNB N_A2_c_588_n 0.0101455f $X=-0.19 $Y=-0.245 $X2=2.095 $Y2=1.385
cc_43 VNB N_A1_M1002_g 0.0348369f $X=-0.19 $Y=-0.245 $X2=4.105 $Y2=1.96
cc_44 VNB N_A1_M1025_g 0.0334816f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_45 VNB A1 0.00223017f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.22
cc_46 VNB N_A1_c_661_n 0.0248414f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_47 VNB N_VPWR_c_716_n 0.362705f $X=-0.19 $Y=-0.245 $X2=5.925 $Y2=2.115
cc_48 VNB N_X_c_843_n 0.00277475f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_49 VNB N_X_c_844_n 0.00221303f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_50 VNB N_X_c_845_n 0.00932569f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.22
cc_51 VNB N_X_c_846_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=1.455 $Y2=1.765
cc_52 VNB N_X_c_847_n 0.00280594f $X=-0.19 $Y=-0.245 $X2=1.42 $Y2=1.385
cc_53 VNB X 0.00825292f $X=-0.19 $Y=-0.245 $X2=2.82 $Y2=2.815
cc_54 VNB N_X_c_849_n 0.00941127f $X=-0.19 $Y=-0.245 $X2=2.985 $Y2=2.035
cc_55 VNB N_VGND_c_959_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.765
cc_56 VNB N_VGND_c_960_n 0.035825f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_57 VNB N_VGND_c_961_n 0.00962229f $X=-0.19 $Y=-0.245 $X2=1.455 $Y2=1.765
cc_58 VNB N_VGND_c_962_n 0.0130012f $X=-0.19 $Y=-0.245 $X2=1.69 $Y2=0.74
cc_59 VNB N_VGND_c_963_n 0.00960417f $X=-0.19 $Y=-0.245 $X2=2.09 $Y2=2.4
cc_60 VNB N_VGND_c_964_n 0.00909146f $X=-0.19 $Y=-0.245 $X2=2.095 $Y2=1.385
cc_61 VNB N_VGND_c_965_n 0.0043117f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_966_n 0.0185368f $X=-0.19 $Y=-0.245 $X2=2.655 $Y2=1.805
cc_63 VNB N_VGND_c_967_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=2.265 $Y2=1.805
cc_64 VNB N_VGND_c_968_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=2.82 $Y2=2.815
cc_65 VNB N_VGND_c_969_n 0.075059f $X=-0.19 $Y=-0.245 $X2=4.42 $Y2=2.055
cc_66 VNB N_VGND_c_970_n 0.0187933f $X=-0.19 $Y=-0.245 $X2=2.1 $Y2=1.385
cc_67 VNB N_VGND_c_971_n 0.0186685f $X=-0.19 $Y=-0.245 $X2=2.82 $Y2=2.105
cc_68 VNB N_VGND_c_972_n 0.0175226f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_973_n 0.475145f $X=-0.19 $Y=-0.245 $X2=5.615 $Y2=2.075
cc_70 VNB N_VGND_c_974_n 0.00875182f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.492
cc_71 VNB N_VGND_c_975_n 0.00632279f $X=-0.19 $Y=-0.245 $X2=1.69 $Y2=1.492
cc_72 VNB N_VGND_c_976_n 0.00632279f $X=-0.19 $Y=-0.245 $X2=2.19 $Y2=1.492
cc_73 VNB N_VGND_c_977_n 0.00626177f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_564_78#_c_1058_n 0.00479371f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.74
cc_75 VNB N_A_564_78#_c_1059_n 0.0219218f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_76 VNB N_A_564_78#_c_1060_n 0.00443708f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_77 VNB N_A_564_78#_c_1061_n 0.00252909f $X=-0.19 $Y=-0.245 $X2=1.69 $Y2=0.74
cc_78 VNB N_A_564_78#_c_1062_n 0.00373444f $X=-0.19 $Y=-0.245 $X2=2.19 $Y2=0.74
cc_79 VNB N_A_564_78#_c_1063_n 0.00716619f $X=-0.19 $Y=-0.245 $X2=1.42 $Y2=1.385
cc_80 VNB N_A_564_78#_c_1064_n 0.018815f $X=-0.19 $Y=-0.245 $X2=2.18 $Y2=1.55
cc_81 VNB N_A_564_78#_c_1065_n 0.0100504f $X=-0.19 $Y=-0.245 $X2=2.82 $Y2=2.12
cc_82 VPB N_A_83_244#_c_158_n 0.0174338f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_83 VPB N_A_83_244#_c_159_n 0.0153284f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.765
cc_84 VPB N_A_83_244#_c_160_n 0.0160808f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=1.765
cc_85 VPB N_A_83_244#_c_161_n 0.0164176f $X=-0.19 $Y=1.66 $X2=2.09 $Y2=1.765
cc_86 VPB N_A_83_244#_c_153_n 5.97158e-19 $X=-0.19 $Y=1.66 $X2=2.18 $Y2=1.72
cc_87 VPB N_A_83_244#_c_163_n 0.00586895f $X=-0.19 $Y=1.66 $X2=2.655 $Y2=1.805
cc_88 VPB N_A_83_244#_c_164_n 0.00292509f $X=-0.19 $Y=1.66 $X2=2.82 $Y2=2.815
cc_89 VPB N_A_83_244#_c_165_n 0.00719187f $X=-0.19 $Y=1.66 $X2=4.09 $Y2=2.035
cc_90 VPB N_A_83_244#_c_166_n 0.00289722f $X=-0.19 $Y=1.66 $X2=4.255 $Y2=2.815
cc_91 VPB N_A_83_244#_c_167_n 0.00596316f $X=-0.19 $Y=1.66 $X2=5.53 $Y2=2.055
cc_92 VPB N_A_83_244#_c_155_n 0.00447657f $X=-0.19 $Y=1.66 $X2=5.615 $Y2=1.95
cc_93 VPB N_A_83_244#_c_156_n 0.0298911f $X=-0.19 $Y=1.66 $X2=2.1 $Y2=1.385
cc_94 VPB N_A_83_244#_c_170_n 0.00488608f $X=-0.19 $Y=1.66 $X2=2.82 $Y2=1.805
cc_95 VPB N_A_83_244#_c_171_n 0.00283403f $X=-0.19 $Y=1.66 $X2=4.255 $Y2=2.105
cc_96 VPB N_A_83_244#_c_172_n 0.00278108f $X=-0.19 $Y=1.66 $X2=5.615 $Y2=2.075
cc_97 VPB N_B1_c_337_n 0.00758951f $X=-0.19 $Y=1.66 $X2=2.67 $Y2=1.96
cc_98 VPB N_B1_c_349_n 0.0224491f $X=-0.19 $Y=1.66 $X2=4.105 $Y2=1.96
cc_99 VPB N_B1_c_350_n 0.0197945f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 VPB N_B1_c_351_n 0.024119f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_101 VPB N_B1_c_352_n 0.0120048f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=1.22
cc_102 VPB N_B1_c_345_n 0.0192611f $X=-0.19 $Y=1.66 $X2=1.42 $Y2=1.385
cc_103 VPB N_B1_c_346_n 0.00280541f $X=-0.19 $Y=1.66 $X2=1.42 $Y2=1.385
cc_104 VPB N_C1_c_454_n 0.0182745f $X=-0.19 $Y=1.66 $X2=4.2 $Y2=0.39
cc_105 VPB N_C1_c_447_n 0.0080547f $X=-0.19 $Y=1.66 $X2=5.765 $Y2=1.96
cc_106 VPB N_C1_c_456_n 0.0184202f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB N_C1_c_450_n 0.0351936f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_108 VPB N_C1_c_452_n 0.0138017f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.765
cc_109 VPB C1 0.00342808f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_110 VPB N_A3_c_524_n 0.0182977f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_A3_c_525_n 0.0155268f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB A3 0.00202188f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_113 VPB N_A3_c_523_n 0.0331596f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=1.22
cc_114 VPB N_A2_c_579_n 0.00818609f $X=-0.19 $Y=1.66 $X2=2.67 $Y2=1.96
cc_115 VPB N_A2_c_590_n 0.0221167f $X=-0.19 $Y=1.66 $X2=4.105 $Y2=1.96
cc_116 VPB N_A2_c_581_n 0.00737402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_A2_c_592_n 0.0283248f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB A2 0.0100864f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=0.74
cc_119 VPB N_A1_c_662_n 0.0157463f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_A1_c_663_n 0.0150726f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB A1 0.00221652f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=1.22
cc_122 VPB N_A1_c_661_n 0.0360023f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=0.74
cc_123 VPB N_VPWR_c_717_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.765
cc_124 VPB N_VPWR_c_718_n 0.0570389f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_125 VPB N_VPWR_c_719_n 0.00651803f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=2.4
cc_126 VPB N_VPWR_c_720_n 0.0210836f $X=-0.19 $Y=1.66 $X2=2.09 $Y2=1.765
cc_127 VPB N_VPWR_c_721_n 0.00655695f $X=-0.19 $Y=1.66 $X2=2.19 $Y2=0.74
cc_128 VPB N_VPWR_c_722_n 0.00966671f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_723_n 0.00129618f $X=-0.19 $Y=1.66 $X2=2.18 $Y2=1.72
cc_130 VPB N_VPWR_c_724_n 0.0121876f $X=-0.19 $Y=1.66 $X2=2.655 $Y2=1.805
cc_131 VPB N_VPWR_c_725_n 0.0185368f $X=-0.19 $Y=1.66 $X2=4.255 $Y2=2.815
cc_132 VPB N_VPWR_c_726_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_727_n 0.00737409f $X=-0.19 $Y=1.66 $X2=5.53 $Y2=2.055
cc_134 VPB N_VPWR_c_728_n 0.0196495f $X=-0.19 $Y=1.66 $X2=5.615 $Y2=1.3
cc_135 VPB N_VPWR_c_729_n 0.0209234f $X=-0.19 $Y=1.66 $X2=2.82 $Y2=1.805
cc_136 VPB N_VPWR_c_730_n 0.09008f $X=-0.19 $Y=1.66 $X2=5.925 $Y2=2.075
cc_137 VPB N_VPWR_c_716_n 0.0960589f $X=-0.19 $Y=1.66 $X2=5.925 $Y2=2.115
cc_138 VPB N_VPWR_c_732_n 0.00614127f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=1.492
cc_139 VPB N_VPWR_c_733_n 0.00614127f $X=-0.19 $Y=1.66 $X2=2.1 $Y2=1.492
cc_140 VPB N_VPWR_c_734_n 0.013162f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_141 VPB N_X_c_850_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.765
cc_142 VPB N_X_c_851_n 0.00726759f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=2.4
cc_143 VPB N_X_c_852_n 0.00329673f $X=-0.19 $Y=1.66 $X2=2.09 $Y2=2.4
cc_144 VPB N_A_1034_392#_c_912_n 0.017826f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_145 VPB N_A_1034_392#_c_913_n 0.0356091f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=0.74
cc_146 VPB N_A_1034_392#_c_914_n 0.00259481f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=0.74
cc_147 VPB N_A_1034_392#_c_915_n 0.00220046f $X=-0.19 $Y=1.66 $X2=1.455
+ $Y2=1.765
cc_148 N_A_83_244#_c_161_n N_B1_c_337_n 0.00415746f $X=2.09 $Y=1.765 $X2=0 $Y2=0
cc_149 N_A_83_244#_c_153_n N_B1_c_337_n 0.00328959f $X=2.18 $Y=1.72 $X2=0 $Y2=0
cc_150 N_A_83_244#_c_163_n N_B1_c_337_n 0.00427622f $X=2.655 $Y=1.805 $X2=0
+ $Y2=0
cc_151 N_A_83_244#_c_156_n N_B1_c_337_n 0.00746893f $X=2.1 $Y=1.385 $X2=0 $Y2=0
cc_152 N_A_83_244#_c_170_n N_B1_c_337_n 0.00178391f $X=2.82 $Y=1.805 $X2=0 $Y2=0
cc_153 N_A_83_244#_c_161_n N_B1_c_349_n 0.0186898f $X=2.09 $Y=1.765 $X2=0 $Y2=0
cc_154 N_A_83_244#_c_163_n N_B1_c_349_n 0.00898996f $X=2.655 $Y=1.805 $X2=0
+ $Y2=0
cc_155 N_A_83_244#_c_164_n N_B1_c_349_n 0.0086908f $X=2.82 $Y=2.815 $X2=0 $Y2=0
cc_156 N_A_83_244#_c_170_n N_B1_c_349_n 0.00678377f $X=2.82 $Y=1.805 $X2=0 $Y2=0
cc_157 N_A_83_244#_c_165_n N_B1_c_338_n 0.00263013f $X=4.09 $Y=2.035 $X2=0 $Y2=0
cc_158 N_A_83_244#_c_170_n N_B1_c_338_n 0.00181329f $X=2.82 $Y=1.805 $X2=0 $Y2=0
cc_159 N_A_83_244#_c_166_n N_B1_c_350_n 0.00453404f $X=4.255 $Y=2.815 $X2=0
+ $Y2=0
cc_160 N_A_83_244#_c_167_n N_B1_c_350_n 0.0170971f $X=5.53 $Y=2.055 $X2=0 $Y2=0
cc_161 N_A_83_244#_c_171_n N_B1_c_350_n 6.46971e-19 $X=4.255 $Y=2.105 $X2=0
+ $Y2=0
cc_162 N_A_83_244#_c_167_n N_B1_c_351_n 0.0175206f $X=5.53 $Y=2.055 $X2=0 $Y2=0
cc_163 N_A_83_244#_c_154_n N_B1_c_351_n 4.31824e-19 $X=5.53 $Y=1.215 $X2=0 $Y2=0
cc_164 N_A_83_244#_c_154_n N_B1_M1024_g 0.0147682f $X=5.53 $Y=1.215 $X2=0 $Y2=0
cc_165 N_A_83_244#_c_155_n N_B1_M1024_g 0.00309212f $X=5.615 $Y=1.95 $X2=0 $Y2=0
cc_166 N_A_83_244#_c_170_n N_B1_c_341_n 0.002856f $X=2.82 $Y=1.805 $X2=0 $Y2=0
cc_167 N_A_83_244#_c_157_n N_B1_c_341_n 0.013759f $X=4.42 $Y=1.1 $X2=0 $Y2=0
cc_168 N_A_83_244#_c_151_n N_B1_c_342_n 0.00371662f $X=2.19 $Y=1.22 $X2=0 $Y2=0
cc_169 N_A_83_244#_c_152_n N_B1_c_342_n 0.0204545f $X=2.18 $Y=1.55 $X2=0 $Y2=0
cc_170 N_A_83_244#_c_163_n N_B1_c_342_n 0.010768f $X=2.655 $Y=1.805 $X2=0 $Y2=0
cc_171 N_A_83_244#_c_156_n N_B1_c_342_n 4.17118e-19 $X=2.1 $Y=1.385 $X2=0 $Y2=0
cc_172 N_A_83_244#_c_170_n N_B1_c_342_n 0.0220402f $X=2.82 $Y=1.805 $X2=0 $Y2=0
cc_173 N_A_83_244#_c_157_n N_B1_c_343_n 0.00254877f $X=4.42 $Y=1.1 $X2=0 $Y2=0
cc_174 N_A_83_244#_c_165_n N_B1_c_381_n 0.00433757f $X=4.09 $Y=2.035 $X2=0 $Y2=0
cc_175 N_A_83_244#_c_171_n N_B1_c_381_n 0.00420141f $X=4.255 $Y=2.105 $X2=0
+ $Y2=0
cc_176 N_A_83_244#_c_152_n N_B1_c_344_n 4.16751e-19 $X=2.18 $Y=1.55 $X2=0 $Y2=0
cc_177 N_A_83_244#_c_156_n N_B1_c_344_n 0.0182576f $X=2.1 $Y=1.385 $X2=0 $Y2=0
cc_178 N_A_83_244#_c_170_n N_B1_c_344_n 0.00118721f $X=2.82 $Y=1.805 $X2=0 $Y2=0
cc_179 N_A_83_244#_c_154_n N_B1_c_345_n 0.00417712f $X=5.53 $Y=1.215 $X2=0 $Y2=0
cc_180 N_A_83_244#_c_155_n N_B1_c_345_n 0.00230015f $X=5.615 $Y=1.95 $X2=0 $Y2=0
cc_181 N_A_83_244#_c_167_n N_B1_c_346_n 0.0324034f $X=5.53 $Y=2.055 $X2=0 $Y2=0
cc_182 N_A_83_244#_c_155_n N_B1_c_346_n 0.0257722f $X=5.615 $Y=1.95 $X2=0 $Y2=0
cc_183 N_A_83_244#_c_167_n N_B1_c_347_n 0.0208365f $X=5.53 $Y=2.055 $X2=0 $Y2=0
cc_184 N_A_83_244#_c_154_n N_B1_c_347_n 0.0575594f $X=5.53 $Y=1.215 $X2=0 $Y2=0
cc_185 N_A_83_244#_c_171_n N_B1_c_347_n 0.0143391f $X=4.255 $Y=2.105 $X2=0 $Y2=0
cc_186 N_A_83_244#_c_157_n N_B1_c_347_n 0.0198993f $X=4.42 $Y=1.1 $X2=0 $Y2=0
cc_187 N_A_83_244#_c_165_n N_C1_c_454_n 0.0164477f $X=4.09 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_188 N_A_83_244#_c_170_n N_C1_c_454_n 0.0131838f $X=2.82 $Y=1.805 $X2=-0.19
+ $Y2=-0.245
cc_189 N_A_83_244#_c_165_n N_C1_c_447_n 0.0100309f $X=4.09 $Y=2.035 $X2=0 $Y2=0
cc_190 N_A_83_244#_c_165_n N_C1_c_456_n 0.0151009f $X=4.09 $Y=2.035 $X2=0 $Y2=0
cc_191 N_A_83_244#_c_166_n N_C1_c_456_n 0.0135822f $X=4.255 $Y=2.815 $X2=0 $Y2=0
cc_192 N_A_83_244#_c_171_n N_C1_c_456_n 0.00210498f $X=4.255 $Y=2.105 $X2=0
+ $Y2=0
cc_193 N_A_83_244#_c_157_n N_C1_M1008_g 0.00560337f $X=4.42 $Y=1.1 $X2=0 $Y2=0
cc_194 N_A_83_244#_c_157_n N_C1_c_449_n 0.00502784f $X=4.42 $Y=1.1 $X2=0 $Y2=0
cc_195 N_A_83_244#_c_165_n N_C1_c_450_n 0.00512687f $X=4.09 $Y=2.035 $X2=0 $Y2=0
cc_196 N_A_83_244#_c_171_n N_C1_c_450_n 0.00283621f $X=4.255 $Y=2.105 $X2=0
+ $Y2=0
cc_197 N_A_83_244#_c_154_n N_C1_M1017_g 0.00993727f $X=5.53 $Y=1.215 $X2=0 $Y2=0
cc_198 N_A_83_244#_c_157_n N_C1_M1017_g 0.00384839f $X=4.42 $Y=1.1 $X2=0 $Y2=0
cc_199 N_A_83_244#_c_165_n N_C1_c_452_n 0.00123317f $X=4.09 $Y=2.035 $X2=0 $Y2=0
cc_200 N_A_83_244#_c_170_n N_C1_c_452_n 0.00376272f $X=2.82 $Y=1.805 $X2=0 $Y2=0
cc_201 N_A_83_244#_c_165_n C1 0.0270133f $X=4.09 $Y=2.035 $X2=0 $Y2=0
cc_202 N_A_83_244#_c_170_n C1 0.00217232f $X=2.82 $Y=1.805 $X2=0 $Y2=0
cc_203 N_A_83_244#_c_154_n N_A3_M1012_g 0.00854518f $X=5.53 $Y=1.215 $X2=0 $Y2=0
cc_204 N_A_83_244#_c_155_n N_A3_M1012_g 0.0037207f $X=5.615 $Y=1.95 $X2=0 $Y2=0
cc_205 N_A_83_244#_c_155_n N_A3_c_524_n 0.00240123f $X=5.615 $Y=1.95 $X2=0 $Y2=0
cc_206 N_A_83_244#_c_172_n N_A3_c_524_n 0.0151432f $X=5.615 $Y=2.075 $X2=0 $Y2=0
cc_207 N_A_83_244#_c_155_n N_A3_c_525_n 3.4268e-19 $X=5.615 $Y=1.95 $X2=0 $Y2=0
cc_208 N_A_83_244#_c_172_n N_A3_c_525_n 0.00365356f $X=5.615 $Y=2.075 $X2=0
+ $Y2=0
cc_209 N_A_83_244#_c_154_n N_A3_M1018_g 8.93268e-19 $X=5.53 $Y=1.215 $X2=0 $Y2=0
cc_210 N_A_83_244#_c_155_n N_A3_M1018_g 6.3266e-19 $X=5.615 $Y=1.95 $X2=0 $Y2=0
cc_211 N_A_83_244#_c_155_n A3 0.0258311f $X=5.615 $Y=1.95 $X2=0 $Y2=0
cc_212 N_A_83_244#_c_172_n A3 0.0187927f $X=5.615 $Y=2.075 $X2=0 $Y2=0
cc_213 N_A_83_244#_c_155_n N_A3_c_523_n 0.0138241f $X=5.615 $Y=1.95 $X2=0 $Y2=0
cc_214 N_A_83_244#_c_172_n N_A3_c_523_n 0.00619154f $X=5.615 $Y=2.075 $X2=0
+ $Y2=0
cc_215 N_A_83_244#_c_172_n N_A2_c_590_n 2.93601e-19 $X=5.615 $Y=2.075 $X2=0
+ $Y2=0
cc_216 N_A_83_244#_c_163_n N_VPWR_M1019_s 0.00174335f $X=2.655 $Y=1.805 $X2=0
+ $Y2=0
cc_217 N_A_83_244#_c_242_p N_VPWR_M1019_s 4.75633e-19 $X=2.265 $Y=1.805 $X2=0
+ $Y2=0
cc_218 N_A_83_244#_c_165_n N_VPWR_M1007_s 0.00951299f $X=4.09 $Y=2.035 $X2=0
+ $Y2=0
cc_219 N_A_83_244#_c_167_n N_VPWR_M1022_d 0.0061135f $X=5.53 $Y=2.055 $X2=0
+ $Y2=0
cc_220 N_A_83_244#_c_158_n N_VPWR_c_718_n 0.0100916f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_221 N_A_83_244#_c_159_n N_VPWR_c_719_n 0.00809349f $X=0.955 $Y=1.765 $X2=0
+ $Y2=0
cc_222 N_A_83_244#_c_160_n N_VPWR_c_719_n 0.0132474f $X=1.455 $Y=1.765 $X2=0
+ $Y2=0
cc_223 N_A_83_244#_c_161_n N_VPWR_c_719_n 6.37802e-19 $X=2.09 $Y=1.765 $X2=0
+ $Y2=0
cc_224 N_A_83_244#_c_160_n N_VPWR_c_720_n 0.00413917f $X=1.455 $Y=1.765 $X2=0
+ $Y2=0
cc_225 N_A_83_244#_c_161_n N_VPWR_c_720_n 0.00413917f $X=2.09 $Y=1.765 $X2=0
+ $Y2=0
cc_226 N_A_83_244#_c_160_n N_VPWR_c_721_n 7.08771e-19 $X=1.455 $Y=1.765 $X2=0
+ $Y2=0
cc_227 N_A_83_244#_c_161_n N_VPWR_c_721_n 0.0151624f $X=2.09 $Y=1.765 $X2=0
+ $Y2=0
cc_228 N_A_83_244#_c_163_n N_VPWR_c_721_n 0.0167214f $X=2.655 $Y=1.805 $X2=0
+ $Y2=0
cc_229 N_A_83_244#_c_242_p N_VPWR_c_721_n 0.00501415f $X=2.265 $Y=1.805 $X2=0
+ $Y2=0
cc_230 N_A_83_244#_c_156_n N_VPWR_c_721_n 2.52799e-19 $X=2.1 $Y=1.385 $X2=0
+ $Y2=0
cc_231 N_A_83_244#_c_170_n N_VPWR_c_721_n 0.0344647f $X=2.82 $Y=1.805 $X2=0
+ $Y2=0
cc_232 N_A_83_244#_c_164_n N_VPWR_c_722_n 0.0435091f $X=2.82 $Y=2.815 $X2=0
+ $Y2=0
cc_233 N_A_83_244#_c_165_n N_VPWR_c_722_n 0.0499208f $X=4.09 $Y=2.035 $X2=0
+ $Y2=0
cc_234 N_A_83_244#_c_166_n N_VPWR_c_722_n 0.026775f $X=4.255 $Y=2.815 $X2=0
+ $Y2=0
cc_235 N_A_83_244#_c_167_n N_VPWR_c_723_n 0.022153f $X=5.53 $Y=2.055 $X2=0 $Y2=0
cc_236 N_A_83_244#_c_166_n N_VPWR_c_724_n 0.0172628f $X=4.255 $Y=2.815 $X2=0
+ $Y2=0
cc_237 N_A_83_244#_c_166_n N_VPWR_c_725_n 0.0145938f $X=4.255 $Y=2.815 $X2=0
+ $Y2=0
cc_238 N_A_83_244#_M1000_d N_VPWR_c_727_n 0.00416858f $X=5.765 $Y=1.96 $X2=0
+ $Y2=0
cc_239 N_A_83_244#_c_167_n N_VPWR_c_727_n 0.0360999f $X=5.53 $Y=2.055 $X2=0
+ $Y2=0
cc_240 N_A_83_244#_c_172_n N_VPWR_c_727_n 0.0271143f $X=5.615 $Y=2.075 $X2=0
+ $Y2=0
cc_241 N_A_83_244#_c_172_n N_VPWR_c_760_n 0.0134407f $X=5.615 $Y=2.075 $X2=0
+ $Y2=0
cc_242 N_A_83_244#_c_158_n N_VPWR_c_728_n 0.00445602f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_243 N_A_83_244#_c_159_n N_VPWR_c_728_n 0.00445602f $X=0.955 $Y=1.765 $X2=0
+ $Y2=0
cc_244 N_A_83_244#_c_164_n N_VPWR_c_729_n 0.0145938f $X=2.82 $Y=2.815 $X2=0
+ $Y2=0
cc_245 N_A_83_244#_c_158_n N_VPWR_c_716_n 0.00861084f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_246 N_A_83_244#_c_159_n N_VPWR_c_716_n 0.00857378f $X=0.955 $Y=1.765 $X2=0
+ $Y2=0
cc_247 N_A_83_244#_c_160_n N_VPWR_c_716_n 0.00819232f $X=1.455 $Y=1.765 $X2=0
+ $Y2=0
cc_248 N_A_83_244#_c_161_n N_VPWR_c_716_n 0.00819232f $X=2.09 $Y=1.765 $X2=0
+ $Y2=0
cc_249 N_A_83_244#_c_164_n N_VPWR_c_716_n 0.0120466f $X=2.82 $Y=2.815 $X2=0
+ $Y2=0
cc_250 N_A_83_244#_c_166_n N_VPWR_c_716_n 0.0120466f $X=4.255 $Y=2.815 $X2=0
+ $Y2=0
cc_251 N_A_83_244#_c_148_n N_X_c_843_n 0.00853575f $X=0.565 $Y=1.22 $X2=0 $Y2=0
cc_252 N_A_83_244#_c_156_n N_X_c_843_n 0.00729077f $X=2.1 $Y=1.385 $X2=0 $Y2=0
cc_253 N_A_83_244#_c_156_n N_X_c_844_n 0.0148828f $X=2.1 $Y=1.385 $X2=0 $Y2=0
cc_254 N_A_83_244#_c_158_n N_X_c_850_n 0.0127167f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_255 N_A_83_244#_c_159_n N_X_c_850_n 0.0130478f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_256 N_A_83_244#_c_160_n N_X_c_850_n 2.20633e-19 $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_257 N_A_83_244#_c_148_n N_X_c_846_n 0.00682285f $X=0.565 $Y=1.22 $X2=0 $Y2=0
cc_258 N_A_83_244#_c_149_n N_X_c_846_n 0.00905927f $X=0.995 $Y=1.22 $X2=0 $Y2=0
cc_259 N_A_83_244#_c_150_n N_X_c_846_n 9.02751e-19 $X=1.69 $Y=1.22 $X2=0 $Y2=0
cc_260 N_A_83_244#_c_159_n N_X_c_851_n 0.0100072f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_261 N_A_83_244#_c_160_n N_X_c_851_n 0.0115773f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_262 N_A_83_244#_c_161_n N_X_c_851_n 0.00121932f $X=2.09 $Y=1.765 $X2=0 $Y2=0
cc_263 N_A_83_244#_c_288_p N_X_c_851_n 0.0504201f $X=2.095 $Y=1.385 $X2=0 $Y2=0
cc_264 N_A_83_244#_c_242_p N_X_c_851_n 0.0130909f $X=2.265 $Y=1.805 $X2=0 $Y2=0
cc_265 N_A_83_244#_c_156_n N_X_c_851_n 0.0217655f $X=2.1 $Y=1.385 $X2=0 $Y2=0
cc_266 N_A_83_244#_c_149_n N_X_c_868_n 0.0150208f $X=0.995 $Y=1.22 $X2=0 $Y2=0
cc_267 N_A_83_244#_c_150_n N_X_c_868_n 0.0128484f $X=1.69 $Y=1.22 $X2=0 $Y2=0
cc_268 N_A_83_244#_c_288_p N_X_c_868_n 0.0574982f $X=2.095 $Y=1.385 $X2=0 $Y2=0
cc_269 N_A_83_244#_c_156_n N_X_c_868_n 0.0140022f $X=2.1 $Y=1.385 $X2=0 $Y2=0
cc_270 N_A_83_244#_c_160_n N_X_c_852_n 0.0076539f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_271 N_A_83_244#_c_161_n N_X_c_852_n 0.0137838f $X=2.09 $Y=1.765 $X2=0 $Y2=0
cc_272 N_A_83_244#_c_149_n N_X_c_847_n 8.98498e-19 $X=0.995 $Y=1.22 $X2=0 $Y2=0
cc_273 N_A_83_244#_c_150_n N_X_c_847_n 0.00833812f $X=1.69 $Y=1.22 $X2=0 $Y2=0
cc_274 N_A_83_244#_c_151_n N_X_c_847_n 0.00282572f $X=2.19 $Y=1.22 $X2=0 $Y2=0
cc_275 N_A_83_244#_c_158_n N_X_c_877_n 0.00397951f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_276 N_A_83_244#_c_159_n N_X_c_877_n 0.00145848f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_277 N_A_83_244#_c_160_n N_X_c_877_n 3.30248e-19 $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_278 N_A_83_244#_c_288_p N_X_c_877_n 0.00300848f $X=2.095 $Y=1.385 $X2=0 $Y2=0
cc_279 N_A_83_244#_c_156_n N_X_c_877_n 0.0258447f $X=2.1 $Y=1.385 $X2=0 $Y2=0
cc_280 N_A_83_244#_c_148_n N_X_c_882_n 0.010085f $X=0.565 $Y=1.22 $X2=0 $Y2=0
cc_281 N_A_83_244#_c_149_n N_X_c_882_n 0.0059694f $X=0.995 $Y=1.22 $X2=0 $Y2=0
cc_282 N_A_83_244#_c_150_n N_X_c_882_n 7.97311e-19 $X=1.69 $Y=1.22 $X2=0 $Y2=0
cc_283 N_A_83_244#_c_288_p N_X_c_882_n 0.00438389f $X=2.095 $Y=1.385 $X2=0 $Y2=0
cc_284 N_A_83_244#_c_156_n N_X_c_882_n 0.0115825f $X=2.1 $Y=1.385 $X2=0 $Y2=0
cc_285 N_A_83_244#_c_156_n X 0.00815293f $X=2.1 $Y=1.385 $X2=0 $Y2=0
cc_286 N_A_83_244#_c_167_n N_A_1034_392#_M1000_s 0.0115931f $X=5.53 $Y=2.055
+ $X2=-0.19 $Y2=-0.245
cc_287 N_A_83_244#_c_172_n N_A_1034_392#_M1000_s 7.96863e-19 $X=5.615 $Y=2.075
+ $X2=-0.19 $Y2=-0.245
cc_288 N_A_83_244#_M1000_d N_A_1034_392#_c_914_n 0.00468183f $X=5.765 $Y=1.96
+ $X2=0 $Y2=0
cc_289 N_A_83_244#_c_148_n N_VGND_c_960_n 0.00874433f $X=0.565 $Y=1.22 $X2=0
+ $Y2=0
cc_290 N_A_83_244#_c_149_n N_VGND_c_961_n 0.00458165f $X=0.995 $Y=1.22 $X2=0
+ $Y2=0
cc_291 N_A_83_244#_c_150_n N_VGND_c_961_n 0.00458165f $X=1.69 $Y=1.22 $X2=0
+ $Y2=0
cc_292 N_A_83_244#_c_150_n N_VGND_c_962_n 5.20559e-19 $X=1.69 $Y=1.22 $X2=0
+ $Y2=0
cc_293 N_A_83_244#_c_151_n N_VGND_c_962_n 0.0127541f $X=2.19 $Y=1.22 $X2=0 $Y2=0
cc_294 N_A_83_244#_c_152_n N_VGND_c_962_n 0.00198701f $X=2.18 $Y=1.55 $X2=0
+ $Y2=0
cc_295 N_A_83_244#_c_163_n N_VGND_c_962_n 0.00637024f $X=2.655 $Y=1.805 $X2=0
+ $Y2=0
cc_296 N_A_83_244#_c_150_n N_VGND_c_966_n 0.00434272f $X=1.69 $Y=1.22 $X2=0
+ $Y2=0
cc_297 N_A_83_244#_c_151_n N_VGND_c_966_n 0.00383152f $X=2.19 $Y=1.22 $X2=0
+ $Y2=0
cc_298 N_A_83_244#_c_148_n N_VGND_c_968_n 0.00434272f $X=0.565 $Y=1.22 $X2=0
+ $Y2=0
cc_299 N_A_83_244#_c_149_n N_VGND_c_968_n 0.00434272f $X=0.995 $Y=1.22 $X2=0
+ $Y2=0
cc_300 N_A_83_244#_c_148_n N_VGND_c_973_n 0.00823934f $X=0.565 $Y=1.22 $X2=0
+ $Y2=0
cc_301 N_A_83_244#_c_149_n N_VGND_c_973_n 0.00822147f $X=0.995 $Y=1.22 $X2=0
+ $Y2=0
cc_302 N_A_83_244#_c_150_n N_VGND_c_973_n 0.00822805f $X=1.69 $Y=1.22 $X2=0
+ $Y2=0
cc_303 N_A_83_244#_c_151_n N_VGND_c_973_n 0.00758198f $X=2.19 $Y=1.22 $X2=0
+ $Y2=0
cc_304 N_A_83_244#_M1008_d N_A_564_78#_c_1059_n 0.00362444f $X=4.2 $Y=0.39 $X2=0
+ $Y2=0
cc_305 N_A_83_244#_c_151_n N_A_564_78#_c_1060_n 6.04331e-19 $X=2.19 $Y=1.22
+ $X2=0 $Y2=0
cc_306 N_A_83_244#_c_154_n N_A_564_78#_c_1068_n 0.0250317f $X=5.53 $Y=1.215
+ $X2=0 $Y2=0
cc_307 N_A_83_244#_c_154_n N_A_564_78#_c_1069_n 0.00781674f $X=5.53 $Y=1.215
+ $X2=0 $Y2=0
cc_308 N_A_83_244#_M1008_d N_A_651_78#_c_1141_n 0.00846345f $X=4.2 $Y=0.39 $X2=0
+ $Y2=0
cc_309 N_A_83_244#_c_154_n N_A_651_78#_c_1141_n 0.00580809f $X=5.53 $Y=1.215
+ $X2=0 $Y2=0
cc_310 N_A_83_244#_c_157_n N_A_651_78#_c_1141_n 0.0191183f $X=4.42 $Y=1.1 $X2=0
+ $Y2=0
cc_311 N_A_83_244#_c_154_n N_A_651_78#_c_1144_n 0.0207769f $X=5.53 $Y=1.215
+ $X2=0 $Y2=0
cc_312 N_B1_c_349_n N_C1_c_454_n 0.0151231f $X=2.595 $Y=1.885 $X2=-0.19
+ $Y2=-0.245
cc_313 N_B1_c_341_n N_C1_c_447_n 0.00655544f $X=3.995 $Y=1.18 $X2=0 $Y2=0
cc_314 N_B1_c_350_n N_C1_c_456_n 0.0202053f $X=4.53 $Y=1.885 $X2=0 $Y2=0
cc_315 N_B1_c_341_n N_C1_M1008_g 0.00910008f $X=3.995 $Y=1.18 $X2=0 $Y2=0
cc_316 N_B1_c_343_n N_C1_M1008_g 0.0018481f $X=4.08 $Y=1.47 $X2=0 $Y2=0
cc_317 N_B1_c_352_n N_C1_c_449_n 0.017407f $X=4.62 $Y=1.785 $X2=0 $Y2=0
cc_318 N_B1_c_347_n N_C1_c_449_n 0.011782f $X=4.925 $Y=1.635 $X2=0 $Y2=0
cc_319 N_B1_c_338_n N_C1_c_450_n 0.00351212f $X=3.105 $Y=1.295 $X2=0 $Y2=0
cc_320 N_B1_c_352_n N_C1_c_450_n 0.00987319f $X=4.62 $Y=1.785 $X2=0 $Y2=0
cc_321 N_B1_c_341_n N_C1_c_450_n 0.0166594f $X=3.995 $Y=1.18 $X2=0 $Y2=0
cc_322 N_B1_c_342_n N_C1_c_450_n 0.00191437f $X=2.91 $Y=1.18 $X2=0 $Y2=0
cc_323 N_B1_c_343_n N_C1_c_450_n 0.0149951f $X=4.08 $Y=1.47 $X2=0 $Y2=0
cc_324 N_B1_c_381_n N_C1_c_450_n 0.00808787f $X=4.165 $Y=1.555 $X2=0 $Y2=0
cc_325 N_B1_c_344_n N_C1_c_450_n 0.00217919f $X=2.67 $Y=1.295 $X2=0 $Y2=0
cc_326 N_B1_c_347_n N_C1_c_450_n 0.0066652f $X=4.925 $Y=1.635 $X2=0 $Y2=0
cc_327 N_B1_M1024_g N_C1_M1017_g 0.0392884f $X=5.145 $Y=0.71 $X2=0 $Y2=0
cc_328 N_B1_c_337_n N_C1_c_452_n 0.00883637f $X=2.595 $Y=1.795 $X2=0 $Y2=0
cc_329 N_B1_c_338_n N_C1_c_452_n 0.0108268f $X=3.105 $Y=1.295 $X2=0 $Y2=0
cc_330 N_B1_c_341_n N_C1_c_452_n 0.00107758f $X=3.995 $Y=1.18 $X2=0 $Y2=0
cc_331 N_B1_c_352_n C1 2.06767e-19 $X=4.62 $Y=1.785 $X2=0 $Y2=0
cc_332 N_B1_c_341_n C1 0.0256488f $X=3.995 $Y=1.18 $X2=0 $Y2=0
cc_333 N_B1_c_342_n C1 0.00418748f $X=2.91 $Y=1.18 $X2=0 $Y2=0
cc_334 N_B1_c_343_n C1 0.00247156f $X=4.08 $Y=1.47 $X2=0 $Y2=0
cc_335 N_B1_c_381_n C1 0.0135996f $X=4.165 $Y=1.555 $X2=0 $Y2=0
cc_336 N_B1_c_344_n C1 4.39048e-19 $X=2.67 $Y=1.295 $X2=0 $Y2=0
cc_337 N_B1_M1024_g N_A3_M1012_g 0.0247641f $X=5.145 $Y=0.71 $X2=0 $Y2=0
cc_338 N_B1_c_345_n N_A3_c_523_n 0.0215643f $X=5.195 $Y=1.635 $X2=0 $Y2=0
cc_339 N_B1_c_346_n N_A3_c_523_n 3.58845e-19 $X=5.195 $Y=1.635 $X2=0 $Y2=0
cc_340 N_B1_c_349_n N_VPWR_c_721_n 0.00808974f $X=2.595 $Y=1.885 $X2=0 $Y2=0
cc_341 N_B1_c_349_n N_VPWR_c_722_n 6.90782e-19 $X=2.595 $Y=1.885 $X2=0 $Y2=0
cc_342 N_B1_c_350_n N_VPWR_c_723_n 0.00240559f $X=4.53 $Y=1.885 $X2=0 $Y2=0
cc_343 N_B1_c_350_n N_VPWR_c_724_n 0.00920476f $X=4.53 $Y=1.885 $X2=0 $Y2=0
cc_344 N_B1_c_350_n N_VPWR_c_725_n 0.00413917f $X=4.53 $Y=1.885 $X2=0 $Y2=0
cc_345 N_B1_c_349_n N_VPWR_c_729_n 0.00445602f $X=2.595 $Y=1.885 $X2=0 $Y2=0
cc_346 N_B1_c_349_n N_VPWR_c_716_n 0.0085864f $X=2.595 $Y=1.885 $X2=0 $Y2=0
cc_347 N_B1_c_350_n N_VPWR_c_716_n 0.00818241f $X=4.53 $Y=1.885 $X2=0 $Y2=0
cc_348 N_B1_M1003_g N_VGND_c_962_n 0.00493098f $X=3.18 $Y=0.71 $X2=0 $Y2=0
cc_349 N_B1_c_342_n N_VGND_c_962_n 0.00534492f $X=2.91 $Y=1.18 $X2=0 $Y2=0
cc_350 N_B1_c_344_n N_VGND_c_962_n 5.0064e-19 $X=2.67 $Y=1.295 $X2=0 $Y2=0
cc_351 N_B1_M1003_g N_VGND_c_969_n 9.78591e-19 $X=3.18 $Y=0.71 $X2=0 $Y2=0
cc_352 N_B1_M1024_g N_VGND_c_969_n 9.59479e-19 $X=5.145 $Y=0.71 $X2=0 $Y2=0
cc_353 N_B1_M1003_g N_A_564_78#_c_1058_n 0.0134061f $X=3.18 $Y=0.71 $X2=0 $Y2=0
cc_354 N_B1_c_341_n N_A_564_78#_c_1058_n 0.0153407f $X=3.995 $Y=1.18 $X2=0 $Y2=0
cc_355 N_B1_c_342_n N_A_564_78#_c_1058_n 0.00980495f $X=2.91 $Y=1.18 $X2=0 $Y2=0
cc_356 N_B1_c_344_n N_A_564_78#_c_1058_n 0.00164878f $X=2.67 $Y=1.295 $X2=0
+ $Y2=0
cc_357 N_B1_M1003_g N_A_564_78#_c_1059_n 0.0111614f $X=3.18 $Y=0.71 $X2=0 $Y2=0
cc_358 N_B1_M1024_g N_A_564_78#_c_1059_n 0.0144367f $X=5.145 $Y=0.71 $X2=0 $Y2=0
cc_359 N_B1_c_341_n N_A_564_78#_c_1059_n 0.0033315f $X=3.995 $Y=1.18 $X2=0 $Y2=0
cc_360 N_B1_M1003_g N_A_564_78#_c_1060_n 0.00406839f $X=3.18 $Y=0.71 $X2=0 $Y2=0
cc_361 N_B1_c_341_n N_A_651_78#_c_1141_n 0.00392744f $X=3.995 $Y=1.18 $X2=0
+ $Y2=0
cc_362 N_B1_c_341_n N_A_651_78#_c_1146_n 0.0534009f $X=3.995 $Y=1.18 $X2=0 $Y2=0
cc_363 N_B1_c_341_n N_A_651_78#_c_1147_n 0.00440496f $X=3.995 $Y=1.18 $X2=0
+ $Y2=0
cc_364 N_B1_M1024_g N_A_651_78#_c_1144_n 0.00436944f $X=5.145 $Y=0.71 $X2=0
+ $Y2=0
cc_365 N_C1_c_454_n N_VPWR_c_722_n 0.0132956f $X=3.165 $Y=1.885 $X2=0 $Y2=0
cc_366 N_C1_c_456_n N_VPWR_c_722_n 0.00266023f $X=4.03 $Y=1.885 $X2=0 $Y2=0
cc_367 N_C1_c_456_n N_VPWR_c_724_n 4.49956e-19 $X=4.03 $Y=1.885 $X2=0 $Y2=0
cc_368 N_C1_c_456_n N_VPWR_c_725_n 0.00445602f $X=4.03 $Y=1.885 $X2=0 $Y2=0
cc_369 N_C1_c_454_n N_VPWR_c_729_n 0.00413917f $X=3.165 $Y=1.885 $X2=0 $Y2=0
cc_370 N_C1_c_454_n N_VPWR_c_716_n 0.00818781f $X=3.165 $Y=1.885 $X2=0 $Y2=0
cc_371 N_C1_c_456_n N_VPWR_c_716_n 0.00860197f $X=4.03 $Y=1.885 $X2=0 $Y2=0
cc_372 N_C1_M1008_g N_VGND_c_969_n 9.59479e-19 $X=4.125 $Y=0.71 $X2=0 $Y2=0
cc_373 N_C1_M1017_g N_VGND_c_969_n 9.59479e-19 $X=4.715 $Y=0.71 $X2=0 $Y2=0
cc_374 N_C1_M1008_g N_A_564_78#_c_1059_n 0.013136f $X=4.125 $Y=0.71 $X2=0 $Y2=0
cc_375 N_C1_M1017_g N_A_564_78#_c_1059_n 0.0110839f $X=4.715 $Y=0.71 $X2=0 $Y2=0
cc_376 N_C1_M1008_g N_A_651_78#_c_1141_n 0.00973441f $X=4.125 $Y=0.71 $X2=0
+ $Y2=0
cc_377 N_C1_c_449_n N_A_651_78#_c_1141_n 0.00128534f $X=4.64 $Y=1.395 $X2=0
+ $Y2=0
cc_378 N_C1_M1017_g N_A_651_78#_c_1141_n 0.0095672f $X=4.715 $Y=0.71 $X2=0 $Y2=0
cc_379 N_C1_c_450_n N_A_651_78#_c_1146_n 8.49316e-19 $X=4.2 $Y=1.395 $X2=0 $Y2=0
cc_380 N_C1_M1008_g N_A_651_78#_c_1147_n 0.00460933f $X=4.125 $Y=0.71 $X2=0
+ $Y2=0
cc_381 N_C1_M1017_g N_A_651_78#_c_1147_n 7.12735e-19 $X=4.715 $Y=0.71 $X2=0
+ $Y2=0
cc_382 N_C1_M1008_g N_A_651_78#_c_1144_n 8.54543e-19 $X=4.125 $Y=0.71 $X2=0
+ $Y2=0
cc_383 N_C1_M1017_g N_A_651_78#_c_1144_n 0.00532525f $X=4.715 $Y=0.71 $X2=0
+ $Y2=0
cc_384 A3 N_A2_c_579_n 0.00131728f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_385 N_A3_c_523_n N_A2_c_579_n 0.0257444f $X=6.16 $Y=1.652 $X2=0 $Y2=0
cc_386 N_A3_c_525_n N_A2_c_590_n 0.0335496f $X=6.16 $Y=1.885 $X2=0 $Y2=0
cc_387 N_A3_M1018_g N_A2_M1006_g 0.0143172f $X=6.21 $Y=0.71 $X2=0 $Y2=0
cc_388 N_A3_M1018_g N_A2_c_584_n 0.00186424f $X=6.21 $Y=0.71 $X2=0 $Y2=0
cc_389 A3 N_A2_c_584_n 0.00592112f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_390 N_A3_M1018_g N_A2_c_585_n 0.00930097f $X=6.21 $Y=0.71 $X2=0 $Y2=0
cc_391 N_A3_c_524_n N_VPWR_c_723_n 0.00129988f $X=5.69 $Y=1.885 $X2=0 $Y2=0
cc_392 N_A3_c_524_n N_VPWR_c_724_n 0.00721881f $X=5.69 $Y=1.885 $X2=0 $Y2=0
cc_393 N_A3_c_524_n N_VPWR_c_727_n 0.0130736f $X=5.69 $Y=1.885 $X2=0 $Y2=0
cc_394 N_A3_c_525_n N_VPWR_c_727_n 0.0132346f $X=6.16 $Y=1.885 $X2=0 $Y2=0
cc_395 A3 N_VPWR_c_727_n 0.002553f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_396 N_A3_c_525_n N_VPWR_c_760_n 0.0068898f $X=6.16 $Y=1.885 $X2=0 $Y2=0
cc_397 N_A3_c_524_n N_VPWR_c_730_n 0.00294338f $X=5.69 $Y=1.885 $X2=0 $Y2=0
cc_398 N_A3_c_525_n N_VPWR_c_730_n 0.00292731f $X=6.16 $Y=1.885 $X2=0 $Y2=0
cc_399 N_A3_c_524_n N_VPWR_c_716_n 0.00366792f $X=5.69 $Y=1.885 $X2=0 $Y2=0
cc_400 N_A3_c_525_n N_VPWR_c_716_n 0.00361322f $X=6.16 $Y=1.885 $X2=0 $Y2=0
cc_401 N_A3_c_524_n N_A_1034_392#_c_914_n 0.0160323f $X=5.69 $Y=1.885 $X2=0
+ $Y2=0
cc_402 N_A3_c_525_n N_A_1034_392#_c_914_n 0.00975758f $X=6.16 $Y=1.885 $X2=0
+ $Y2=0
cc_403 N_A3_c_524_n N_A_1034_392#_c_915_n 5.32047e-19 $X=5.69 $Y=1.885 $X2=0
+ $Y2=0
cc_404 N_A3_c_525_n N_A_1034_392#_c_915_n 0.00427068f $X=6.16 $Y=1.885 $X2=0
+ $Y2=0
cc_405 N_A3_M1012_g N_VGND_c_963_n 0.00123358f $X=5.675 $Y=0.71 $X2=0 $Y2=0
cc_406 N_A3_M1018_g N_VGND_c_963_n 0.00328128f $X=6.21 $Y=0.71 $X2=0 $Y2=0
cc_407 N_A3_M1012_g N_VGND_c_969_n 0.00563421f $X=5.675 $Y=0.71 $X2=0 $Y2=0
cc_408 N_A3_M1018_g N_VGND_c_970_n 0.00542877f $X=6.21 $Y=0.71 $X2=0 $Y2=0
cc_409 N_A3_M1012_g N_VGND_c_973_n 0.00539454f $X=5.675 $Y=0.71 $X2=0 $Y2=0
cc_410 N_A3_M1018_g N_VGND_c_973_n 0.00539454f $X=6.21 $Y=0.71 $X2=0 $Y2=0
cc_411 N_A3_M1012_g N_A_564_78#_c_1059_n 0.00134496f $X=5.675 $Y=0.71 $X2=0
+ $Y2=0
cc_412 N_A3_M1012_g N_A_564_78#_c_1069_n 0.0117498f $X=5.675 $Y=0.71 $X2=0 $Y2=0
cc_413 N_A3_M1018_g N_A_564_78#_c_1069_n 0.0117966f $X=6.21 $Y=0.71 $X2=0 $Y2=0
cc_414 A3 N_A_564_78#_c_1069_n 0.0101563f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_415 N_A3_c_523_n N_A_564_78#_c_1069_n 0.00183128f $X=6.16 $Y=1.652 $X2=0
+ $Y2=0
cc_416 N_A3_M1012_g N_A_564_78#_c_1061_n 3.19102e-19 $X=5.675 $Y=0.71 $X2=0
+ $Y2=0
cc_417 N_A3_M1018_g N_A_564_78#_c_1061_n 0.0062568f $X=6.21 $Y=0.71 $X2=0 $Y2=0
cc_418 N_A3_M1012_g N_A_564_78#_c_1065_n 4.15266e-19 $X=5.675 $Y=0.71 $X2=0
+ $Y2=0
cc_419 N_A3_M1018_g N_A_564_78#_c_1065_n 0.00322051f $X=6.21 $Y=0.71 $X2=0 $Y2=0
cc_420 N_A2_M1006_g N_A1_M1002_g 0.0226082f $X=6.645 $Y=0.71 $X2=0 $Y2=0
cc_421 N_A2_c_583_n N_A1_M1002_g 0.0111072f $X=8.205 $Y=1.215 $X2=0 $Y2=0
cc_422 N_A2_c_584_n N_A1_M1002_g 0.00473006f $X=6.935 $Y=1.215 $X2=0 $Y2=0
cc_423 N_A2_c_585_n N_A1_M1002_g 0.0172628f $X=6.69 $Y=1.385 $X2=0 $Y2=0
cc_424 N_A2_c_590_n N_A1_c_662_n 0.0278948f $X=6.615 $Y=1.885 $X2=0 $Y2=0
cc_425 N_A2_c_592_n N_A1_c_663_n 0.0173635f $X=8.105 $Y=1.885 $X2=0 $Y2=0
cc_426 N_A2_c_582_n N_A1_M1025_g 0.0236478f $X=8.145 $Y=1.14 $X2=0 $Y2=0
cc_427 N_A2_c_583_n N_A1_M1025_g 0.0109343f $X=8.205 $Y=1.215 $X2=0 $Y2=0
cc_428 A2 N_A1_M1025_g 7.75467e-19 $X=8.315 $Y=1.21 $X2=0 $Y2=0
cc_429 N_A2_c_587_n N_A1_M1025_g 0.016557f $X=8.145 $Y=1.35 $X2=0 $Y2=0
cc_430 N_A2_c_579_n A1 0.00142776f $X=6.615 $Y=1.795 $X2=0 $Y2=0
cc_431 N_A2_c_581_n A1 0.00548689f $X=8.105 $Y=1.795 $X2=0 $Y2=0
cc_432 N_A2_c_592_n A1 5.49111e-19 $X=8.105 $Y=1.885 $X2=0 $Y2=0
cc_433 N_A2_c_583_n A1 0.0698037f $X=8.205 $Y=1.215 $X2=0 $Y2=0
cc_434 N_A2_c_584_n A1 0.00677213f $X=6.935 $Y=1.215 $X2=0 $Y2=0
cc_435 A2 A1 0.0258837f $X=8.315 $Y=1.21 $X2=0 $Y2=0
cc_436 N_A2_c_587_n A1 0.00199873f $X=8.145 $Y=1.35 $X2=0 $Y2=0
cc_437 N_A2_c_579_n N_A1_c_661_n 0.0124598f $X=6.615 $Y=1.795 $X2=0 $Y2=0
cc_438 N_A2_c_592_n N_A1_c_661_n 0.00430036f $X=8.105 $Y=1.885 $X2=0 $Y2=0
cc_439 N_A2_c_583_n N_A1_c_661_n 0.00448411f $X=8.205 $Y=1.215 $X2=0 $Y2=0
cc_440 N_A2_c_587_n N_A1_c_661_n 0.0181313f $X=8.145 $Y=1.35 $X2=0 $Y2=0
cc_441 N_A2_c_590_n N_VPWR_c_795_n 0.019104f $X=6.615 $Y=1.885 $X2=0 $Y2=0
cc_442 N_A2_c_583_n N_VPWR_c_795_n 0.00415351f $X=8.205 $Y=1.215 $X2=0 $Y2=0
cc_443 N_A2_c_585_n N_VPWR_c_795_n 8.09603e-19 $X=6.69 $Y=1.385 $X2=0 $Y2=0
cc_444 N_A2_c_590_n N_VPWR_c_760_n 0.00921443f $X=6.615 $Y=1.885 $X2=0 $Y2=0
cc_445 N_A2_c_584_n N_VPWR_c_760_n 0.01474f $X=6.935 $Y=1.215 $X2=0 $Y2=0
cc_446 N_A2_c_590_n N_VPWR_c_730_n 0.00278271f $X=6.615 $Y=1.885 $X2=0 $Y2=0
cc_447 N_A2_c_592_n N_VPWR_c_730_n 0.00278271f $X=8.105 $Y=1.885 $X2=0 $Y2=0
cc_448 N_A2_c_590_n N_VPWR_c_716_n 0.00355006f $X=6.615 $Y=1.885 $X2=0 $Y2=0
cc_449 N_A2_c_592_n N_VPWR_c_716_n 0.00357673f $X=8.105 $Y=1.885 $X2=0 $Y2=0
cc_450 N_A2_c_590_n N_A_1034_392#_c_912_n 0.00902645f $X=6.615 $Y=1.885 $X2=0
+ $Y2=0
cc_451 N_A2_c_592_n N_A_1034_392#_c_912_n 0.01424f $X=8.105 $Y=1.885 $X2=0 $Y2=0
cc_452 A2 N_A_1034_392#_c_913_n 0.0256065f $X=8.315 $Y=1.21 $X2=0 $Y2=0
cc_453 N_A2_c_587_n N_A_1034_392#_c_913_n 0.00125053f $X=8.145 $Y=1.35 $X2=0
+ $Y2=0
cc_454 N_A2_c_590_n N_A_1034_392#_c_915_n 0.00554574f $X=6.615 $Y=1.885 $X2=0
+ $Y2=0
cc_455 N_A2_M1006_g N_VGND_c_964_n 0.00320426f $X=6.645 $Y=0.71 $X2=0 $Y2=0
cc_456 N_A2_c_582_n N_VGND_c_965_n 0.00926362f $X=8.145 $Y=1.14 $X2=0 $Y2=0
cc_457 N_A2_M1006_g N_VGND_c_970_n 0.00537471f $X=6.645 $Y=0.71 $X2=0 $Y2=0
cc_458 N_A2_c_582_n N_VGND_c_972_n 0.00468165f $X=8.145 $Y=1.14 $X2=0 $Y2=0
cc_459 N_A2_M1006_g N_VGND_c_973_n 0.00539454f $X=6.645 $Y=0.71 $X2=0 $Y2=0
cc_460 N_A2_c_582_n N_VGND_c_973_n 0.00453141f $X=8.145 $Y=1.14 $X2=0 $Y2=0
cc_461 N_A2_M1006_g N_A_564_78#_c_1061_n 0.00643859f $X=6.645 $Y=0.71 $X2=0
+ $Y2=0
cc_462 N_A2_M1006_g N_A_564_78#_c_1090_n 0.00925963f $X=6.645 $Y=0.71 $X2=0
+ $Y2=0
cc_463 N_A2_c_583_n N_A_564_78#_c_1090_n 0.0206132f $X=8.205 $Y=1.215 $X2=0
+ $Y2=0
cc_464 N_A2_c_584_n N_A_564_78#_c_1090_n 0.020703f $X=6.935 $Y=1.215 $X2=0 $Y2=0
cc_465 N_A2_c_585_n N_A_564_78#_c_1090_n 4.79388e-19 $X=6.69 $Y=1.385 $X2=0
+ $Y2=0
cc_466 N_A2_c_582_n N_A_564_78#_c_1094_n 0.00949048f $X=8.145 $Y=1.14 $X2=0
+ $Y2=0
cc_467 N_A2_c_583_n N_A_564_78#_c_1094_n 0.0380593f $X=8.205 $Y=1.215 $X2=0
+ $Y2=0
cc_468 N_A2_c_588_n N_A_564_78#_c_1094_n 0.00365309f $X=8.37 $Y=1.3 $X2=0 $Y2=0
cc_469 N_A2_c_587_n N_A_564_78#_c_1063_n 0.00189009f $X=8.145 $Y=1.35 $X2=0
+ $Y2=0
cc_470 N_A2_c_588_n N_A_564_78#_c_1063_n 0.022669f $X=8.37 $Y=1.3 $X2=0 $Y2=0
cc_471 N_A2_c_582_n N_A_564_78#_c_1064_n 8.90981e-19 $X=8.145 $Y=1.14 $X2=0
+ $Y2=0
cc_472 N_A2_M1006_g N_A_564_78#_c_1065_n 0.00273654f $X=6.645 $Y=0.71 $X2=0
+ $Y2=0
cc_473 N_A2_c_584_n N_A_564_78#_c_1065_n 0.00581955f $X=6.935 $Y=1.215 $X2=0
+ $Y2=0
cc_474 N_A2_c_585_n N_A_564_78#_c_1065_n 3.50288e-19 $X=6.69 $Y=1.385 $X2=0
+ $Y2=0
cc_475 N_A2_c_583_n N_A_564_78#_c_1103_n 0.0242243f $X=8.205 $Y=1.215 $X2=0
+ $Y2=0
cc_476 N_A1_c_662_n N_VPWR_c_795_n 0.017314f $X=7.185 $Y=1.885 $X2=0 $Y2=0
cc_477 N_A1_c_663_n N_VPWR_c_795_n 0.00517585f $X=7.635 $Y=1.885 $X2=0 $Y2=0
cc_478 A1 N_VPWR_c_795_n 0.0318171f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_479 N_A1_c_661_n N_VPWR_c_795_n 0.00624074f $X=7.635 $Y=1.677 $X2=0 $Y2=0
cc_480 N_A1_c_662_n N_VPWR_c_760_n 4.34929e-19 $X=7.185 $Y=1.885 $X2=0 $Y2=0
cc_481 N_A1_c_662_n N_VPWR_c_730_n 0.00278271f $X=7.185 $Y=1.885 $X2=0 $Y2=0
cc_482 N_A1_c_663_n N_VPWR_c_730_n 0.00278271f $X=7.635 $Y=1.885 $X2=0 $Y2=0
cc_483 N_A1_c_662_n N_VPWR_c_716_n 0.00354878f $X=7.185 $Y=1.885 $X2=0 $Y2=0
cc_484 N_A1_c_663_n N_VPWR_c_716_n 0.00354083f $X=7.635 $Y=1.885 $X2=0 $Y2=0
cc_485 N_A1_c_662_n N_A_1034_392#_c_912_n 0.00995575f $X=7.185 $Y=1.885 $X2=0
+ $Y2=0
cc_486 N_A1_c_663_n N_A_1034_392#_c_912_n 0.00948594f $X=7.635 $Y=1.885 $X2=0
+ $Y2=0
cc_487 N_A1_c_662_n N_A_1034_392#_c_915_n 4.89504e-19 $X=7.185 $Y=1.885 $X2=0
+ $Y2=0
cc_488 N_A1_c_662_n N_A_1338_392#_c_948_n 0.00853169f $X=7.185 $Y=1.885 $X2=0
+ $Y2=0
cc_489 N_A1_c_663_n N_A_1338_392#_c_948_n 0.0126242f $X=7.635 $Y=1.885 $X2=0
+ $Y2=0
cc_490 N_A1_c_663_n N_A_1338_392#_c_950_n 0.00529359f $X=7.635 $Y=1.885 $X2=0
+ $Y2=0
cc_491 A1 N_A_1338_392#_c_950_n 0.0191734f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_492 N_A1_M1002_g N_VGND_c_964_n 0.00195239f $X=7.17 $Y=0.71 $X2=0 $Y2=0
cc_493 N_A1_M1002_g N_VGND_c_965_n 3.31989e-19 $X=7.17 $Y=0.71 $X2=0 $Y2=0
cc_494 N_A1_M1025_g N_VGND_c_965_n 0.0061006f $X=7.7 $Y=0.71 $X2=0 $Y2=0
cc_495 N_A1_M1002_g N_VGND_c_971_n 0.00562069f $X=7.17 $Y=0.71 $X2=0 $Y2=0
cc_496 N_A1_M1025_g N_VGND_c_971_n 0.00524507f $X=7.7 $Y=0.71 $X2=0 $Y2=0
cc_497 N_A1_M1002_g N_VGND_c_973_n 0.00539454f $X=7.17 $Y=0.71 $X2=0 $Y2=0
cc_498 N_A1_M1025_g N_VGND_c_973_n 0.00507087f $X=7.7 $Y=0.71 $X2=0 $Y2=0
cc_499 N_A1_M1002_g N_A_564_78#_c_1061_n 3.25679e-19 $X=7.17 $Y=0.71 $X2=0 $Y2=0
cc_500 N_A1_M1002_g N_A_564_78#_c_1090_n 0.010115f $X=7.17 $Y=0.71 $X2=0 $Y2=0
cc_501 N_A1_M1002_g N_A_564_78#_c_1062_n 3.71344e-19 $X=7.17 $Y=0.71 $X2=0 $Y2=0
cc_502 N_A1_M1025_g N_A_564_78#_c_1062_n 3.6365e-19 $X=7.7 $Y=0.71 $X2=0 $Y2=0
cc_503 N_A1_M1025_g N_A_564_78#_c_1094_n 0.00962899f $X=7.7 $Y=0.71 $X2=0 $Y2=0
cc_504 N_A1_M1002_g N_A_564_78#_c_1065_n 4.20891e-19 $X=7.17 $Y=0.71 $X2=0 $Y2=0
cc_505 N_VPWR_c_718_n N_X_c_844_n 7.22336e-19 $X=0.28 $Y=1.985 $X2=0 $Y2=0
cc_506 N_VPWR_c_718_n N_X_c_845_n 0.0210943f $X=0.28 $Y=1.985 $X2=0 $Y2=0
cc_507 N_VPWR_c_719_n N_X_c_850_n 0.0353111f $X=1.23 $Y=2.145 $X2=0 $Y2=0
cc_508 N_VPWR_c_728_n N_X_c_850_n 0.014552f $X=1.065 $Y=3.33 $X2=0 $Y2=0
cc_509 N_VPWR_c_716_n N_X_c_850_n 0.0119791f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_510 N_VPWR_M1010_s N_X_c_851_n 0.00250873f $X=1.03 $Y=1.84 $X2=0 $Y2=0
cc_511 N_VPWR_c_719_n N_X_c_851_n 0.0202249f $X=1.23 $Y=2.145 $X2=0 $Y2=0
cc_512 N_VPWR_c_719_n N_X_c_852_n 0.0353111f $X=1.23 $Y=2.145 $X2=0 $Y2=0
cc_513 N_VPWR_c_720_n N_X_c_852_n 0.0146357f $X=2.15 $Y=3.33 $X2=0 $Y2=0
cc_514 N_VPWR_c_721_n N_X_c_852_n 0.0523615f $X=2.315 $Y=2.145 $X2=0 $Y2=0
cc_515 N_VPWR_c_716_n N_X_c_852_n 0.0121141f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_516 N_VPWR_c_718_n N_X_c_877_n 0.0778054f $X=0.28 $Y=1.985 $X2=0 $Y2=0
cc_517 N_VPWR_c_727_n N_A_1034_392#_M1000_s 0.0109768f $X=6.38 $Y=2.255
+ $X2=-0.19 $Y2=-0.245
cc_518 N_VPWR_c_727_n N_A_1034_392#_M1023_s 0.00423011f $X=6.38 $Y=2.255 $X2=0
+ $Y2=0
cc_519 N_VPWR_c_760_n N_A_1034_392#_M1023_s 0.0103806f $X=6.55 $Y=2.255 $X2=0
+ $Y2=0
cc_520 N_VPWR_M1016_d N_A_1034_392#_c_912_n 0.00198204f $X=7.26 $Y=1.96 $X2=0
+ $Y2=0
cc_521 N_VPWR_c_795_n N_A_1034_392#_c_912_n 0.00413192f $X=7.41 $Y=2.18 $X2=0
+ $Y2=0
cc_522 N_VPWR_c_730_n N_A_1034_392#_c_912_n 0.0236566f $X=8.4 $Y=3.33 $X2=0
+ $Y2=0
cc_523 N_VPWR_c_716_n N_A_1034_392#_c_912_n 0.0128296f $X=8.4 $Y=3.33 $X2=0
+ $Y2=0
cc_524 N_VPWR_c_724_n N_A_1034_392#_c_914_n 0.0177419f $X=4.755 $Y=3.245 $X2=0
+ $Y2=0
cc_525 N_VPWR_c_727_n N_A_1034_392#_c_914_n 0.0403132f $X=6.38 $Y=2.255 $X2=0
+ $Y2=0
cc_526 N_VPWR_c_730_n N_A_1034_392#_c_914_n 0.036799f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_527 N_VPWR_c_716_n N_A_1034_392#_c_914_n 0.0363629f $X=8.4 $Y=3.33 $X2=0
+ $Y2=0
cc_528 N_VPWR_c_760_n N_A_1034_392#_c_915_n 0.0403132f $X=6.55 $Y=2.255 $X2=0
+ $Y2=0
cc_529 N_VPWR_c_730_n N_A_1034_392#_c_915_n 0.126554f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_530 N_VPWR_c_716_n N_A_1034_392#_c_915_n 0.0716645f $X=8.4 $Y=3.33 $X2=0
+ $Y2=0
cc_531 N_VPWR_c_795_n N_A_1338_392#_M1001_d 0.0102016f $X=7.41 $Y=2.18 $X2=-0.19
+ $Y2=-0.245
cc_532 N_VPWR_M1016_d N_A_1338_392#_c_948_n 0.0038712f $X=7.26 $Y=1.96 $X2=0
+ $Y2=0
cc_533 N_VPWR_c_795_n N_A_1338_392#_c_948_n 0.0503517f $X=7.41 $Y=2.18 $X2=0
+ $Y2=0
cc_534 N_VPWR_c_795_n N_A_1338_392#_c_950_n 0.0301137f $X=7.41 $Y=2.18 $X2=0
+ $Y2=0
cc_535 N_X_c_868_n N_VGND_M1005_s 0.0111557f $X=1.74 $Y=0.965 $X2=0 $Y2=0
cc_536 N_X_c_843_n N_VGND_c_960_n 0.00682786f $X=0.615 $Y=1.225 $X2=0 $Y2=0
cc_537 N_X_c_846_n N_VGND_c_960_n 0.0240168f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_538 N_X_c_849_n N_VGND_c_960_n 0.0207054f $X=0.24 $Y=1.31 $X2=0 $Y2=0
cc_539 N_X_c_846_n N_VGND_c_961_n 0.0132122f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_540 N_X_c_868_n N_VGND_c_961_n 0.0310653f $X=1.74 $Y=0.965 $X2=0 $Y2=0
cc_541 N_X_c_847_n N_VGND_c_961_n 0.0132122f $X=1.905 $Y=0.515 $X2=0 $Y2=0
cc_542 N_X_c_847_n N_VGND_c_962_n 0.0206774f $X=1.905 $Y=0.515 $X2=0 $Y2=0
cc_543 N_X_c_847_n N_VGND_c_966_n 0.0145947f $X=1.905 $Y=0.515 $X2=0 $Y2=0
cc_544 N_X_c_846_n N_VGND_c_968_n 0.0144922f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_545 N_X_c_846_n N_VGND_c_973_n 0.0118826f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_546 N_X_c_847_n N_VGND_c_973_n 0.0120104f $X=1.905 $Y=0.515 $X2=0 $Y2=0
cc_547 N_A_1034_392#_c_912_n N_A_1338_392#_M1001_d 0.0034401f $X=8.195 $Y=2.99
+ $X2=-0.19 $Y2=1.66
cc_548 N_A_1034_392#_c_912_n N_A_1338_392#_M1027_s 0.00219003f $X=8.195 $Y=2.99
+ $X2=0 $Y2=0
cc_549 N_A_1034_392#_c_912_n N_A_1338_392#_c_948_n 0.0682877f $X=8.195 $Y=2.99
+ $X2=0 $Y2=0
cc_550 N_VGND_c_962_n N_A_564_78#_c_1058_n 0.0336755f $X=2.405 $Y=0.515 $X2=0
+ $Y2=0
cc_551 N_VGND_c_963_n N_A_564_78#_c_1059_n 0.0118455f $X=5.93 $Y=0.535 $X2=0
+ $Y2=0
cc_552 N_VGND_c_969_n N_A_564_78#_c_1059_n 0.161196f $X=5.765 $Y=0 $X2=0 $Y2=0
cc_553 N_VGND_c_973_n N_A_564_78#_c_1059_n 0.0931052f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_554 N_VGND_c_962_n N_A_564_78#_c_1060_n 0.0121617f $X=2.405 $Y=0.515 $X2=0
+ $Y2=0
cc_555 N_VGND_c_969_n N_A_564_78#_c_1060_n 0.0236302f $X=5.765 $Y=0 $X2=0 $Y2=0
cc_556 N_VGND_c_973_n N_A_564_78#_c_1060_n 0.0128247f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_557 N_VGND_M1012_s N_A_564_78#_c_1069_n 0.00786082f $X=5.75 $Y=0.39 $X2=0
+ $Y2=0
cc_558 N_VGND_c_963_n N_A_564_78#_c_1069_n 0.0215299f $X=5.93 $Y=0.535 $X2=0
+ $Y2=0
cc_559 N_VGND_c_973_n N_A_564_78#_c_1069_n 0.0124679f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_560 N_VGND_c_963_n N_A_564_78#_c_1061_n 0.0101711f $X=5.93 $Y=0.535 $X2=0
+ $Y2=0
cc_561 N_VGND_c_964_n N_A_564_78#_c_1061_n 0.0101711f $X=6.93 $Y=0.535 $X2=0
+ $Y2=0
cc_562 N_VGND_c_970_n N_A_564_78#_c_1061_n 0.0134222f $X=6.765 $Y=0 $X2=0 $Y2=0
cc_563 N_VGND_c_973_n N_A_564_78#_c_1061_n 0.0119304f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_564 N_VGND_M1006_s N_A_564_78#_c_1090_n 0.00548639f $X=6.72 $Y=0.39 $X2=0
+ $Y2=0
cc_565 N_VGND_c_964_n N_A_564_78#_c_1090_n 0.0207355f $X=6.93 $Y=0.535 $X2=0
+ $Y2=0
cc_566 N_VGND_c_973_n N_A_564_78#_c_1090_n 0.0124851f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_567 N_VGND_c_964_n N_A_564_78#_c_1062_n 0.012814f $X=6.93 $Y=0.535 $X2=0
+ $Y2=0
cc_568 N_VGND_c_965_n N_A_564_78#_c_1062_n 0.0117536f $X=7.93 $Y=0.535 $X2=0
+ $Y2=0
cc_569 N_VGND_c_971_n N_A_564_78#_c_1062_n 0.0145203f $X=7.765 $Y=0 $X2=0 $Y2=0
cc_570 N_VGND_c_973_n N_A_564_78#_c_1062_n 0.0120696f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_571 N_VGND_M1025_s N_A_564_78#_c_1094_n 0.00381868f $X=7.775 $Y=0.39 $X2=0
+ $Y2=0
cc_572 N_VGND_c_965_n N_A_564_78#_c_1094_n 0.0167502f $X=7.93 $Y=0.535 $X2=0
+ $Y2=0
cc_573 N_VGND_c_973_n N_A_564_78#_c_1094_n 0.0128307f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_574 N_VGND_c_965_n N_A_564_78#_c_1064_n 0.0111714f $X=7.93 $Y=0.535 $X2=0
+ $Y2=0
cc_575 N_VGND_c_972_n N_A_564_78#_c_1064_n 0.0109788f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_576 N_VGND_c_973_n N_A_564_78#_c_1064_n 0.00912577f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_577 N_A_564_78#_c_1059_n N_A_651_78#_M1003_d 0.00807544f $X=5.265 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_578 N_A_564_78#_c_1059_n N_A_651_78#_M1017_s 0.00176461f $X=5.265 $Y=0.34
+ $X2=0 $Y2=0
cc_579 N_A_564_78#_c_1059_n N_A_651_78#_c_1146_n 0.0886249f $X=5.265 $Y=0.34
+ $X2=0 $Y2=0
cc_580 N_A_564_78#_c_1059_n N_A_651_78#_c_1144_n 0.0152459f $X=5.265 $Y=0.34
+ $X2=0 $Y2=0
