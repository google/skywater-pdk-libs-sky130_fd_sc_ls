* File: sky130_fd_sc_ls__mux2_2.spice
* Created: Fri Aug 28 13:29:55 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__mux2_2.pex.spice"
.subckt sky130_fd_sc_ls__mux2_2  VNB VPB A0 A1 S VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* S	S
* A1	A1
* A0	A0
* VPB	VPB
* VNB	VNB
MM1003 N_A_116_368#_M1003_d N_A0_M1003_g N_A_38_74#_M1003_s VNB NSHORT L=0.15
+ W=0.74 AD=0.21275 AS=0.2109 PD=1.315 PS=2.05 NRD=25.128 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75002 A=0.111 P=1.78 MULT=1
MM1006 A_270_74# N_A1_M1006_g N_A_116_368#_M1003_d VNB NSHORT L=0.15 W=0.74
+ AD=0.0888 AS=0.21275 PD=0.98 PS=1.315 NRD=10.536 NRS=22.692 M=1 R=4.93333
+ SA=75000.9 SB=75001.3 A=0.111 P=1.78 MULT=1
MM1010 N_VGND_M1010_d N_S_M1010_g A_270_74# VNB NSHORT L=0.15 W=0.74 AD=0.20535
+ AS=0.0888 PD=1.295 PS=0.98 NRD=0 NRS=10.536 M=1 R=4.93333 SA=75001.3
+ SB=75000.9 A=0.111 P=1.78 MULT=1
MM1005 N_A_38_74#_M1005_d N_A_459_48#_M1005_g N_VGND_M1010_d VNB NSHORT L=0.15
+ W=0.74 AD=0.2183 AS=0.20535 PD=2.07 PS=1.295 NRD=0 NRS=44.592 M=1 R=4.93333
+ SA=75002 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1011 N_VGND_M1011_d N_S_M1011_g N_A_459_48#_M1011_s VNB NSHORT L=0.15 W=0.55
+ AD=0.117568 AS=0.15675 PD=0.984884 PS=1.67 NRD=21.816 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75001.3 A=0.0825 P=1.4 MULT=1
MM1004 N_X_M1004_d N_A_116_368#_M1004_g N_VGND_M1011_d VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.158182 PD=1.02 PS=1.32512 NRD=0 NRS=5.664 M=1 R=4.93333
+ SA=75000.6 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1013 N_X_M1004_d N_A_116_368#_M1013_g N_VGND_M1013_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.2627 PD=1.02 PS=2.19 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.1
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1008 N_A_116_368#_M1008_d N_A0_M1008_g N_A_27_368#_M1008_s VPB PHIGHVT L=0.15
+ W=1 AD=0.15 AS=0.295 PD=1.3 PS=2.59 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75000.7 A=0.15 P=2.3 MULT=1
MM1009 N_A_206_368#_M1009_d N_A1_M1009_g N_A_116_368#_M1008_d VPB PHIGHVT L=0.15
+ W=1 AD=0.295 AS=0.15 PD=2.59 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75000.7 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1000 N_VPWR_M1000_d N_S_M1000_g N_A_27_368#_M1000_s VPB PHIGHVT L=0.15 W=1
+ AD=0.2 AS=0.295 PD=1.4 PS=2.59 NRD=11.8003 NRS=1.9503 M=1 R=6.66667 SA=75000.2
+ SB=75000.8 A=0.15 P=2.3 MULT=1
MM1002 N_A_206_368#_M1002_d N_A_459_48#_M1002_g N_VPWR_M1000_d VPB PHIGHVT
+ L=0.15 W=1 AD=0.295 AS=0.2 PD=2.59 PS=1.4 NRD=1.9503 NRS=11.8003 M=1 R=6.66667
+ SA=75000.8 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1007 N_VPWR_M1007_d N_S_M1007_g N_A_459_48#_M1007_s VPB PHIGHVT L=0.15 W=0.84
+ AD=0.1788 AS=0.2478 PD=1.29857 PS=2.27 NRD=37.0163 NRS=2.3443 M=1 R=5.6
+ SA=75000.2 SB=75001.3 A=0.126 P=1.98 MULT=1
MM1001 N_VPWR_M1007_d N_A_116_368#_M1001_g N_X_M1001_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.2384 AS=0.168 PD=1.73143 PS=1.42 NRD=2.6201 NRS=1.7533 M=1 R=7.46667
+ SA=75000.6 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1012 N_VPWR_M1012_d N_A_116_368#_M1012_g N_X_M1001_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.392 AS=0.168 PD=2.94 PS=1.42 NRD=6.1464 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75000.3 A=0.168 P=2.54 MULT=1
DX14_noxref VNB VPB NWDIODE A=10.5276 P=15.04
c_584 A_270_74# 0 1.6439e-20 $X=1.35 $Y=0.37
*
.include "sky130_fd_sc_ls__mux2_2.pxi.spice"
*
.ends
*
*
