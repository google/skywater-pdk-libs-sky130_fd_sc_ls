# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ls__mux4_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ls__mux4_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  16.80000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A0
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.470000 2.355000 1.800000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.450000 0.890000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.765000 1.260000 9.475000 1.775000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.725000 1.445000 10.435000 1.775000 ;
    END
  END A3
  PIN S0
    ANTENNAGATEAREA  1.263000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.295000 1.435000 8.515000 1.775000 ;
    END
  END S0
  PIN S1
    ANTENNAGATEAREA  0.771000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.150000 1.275000 13.865000 1.300000 ;
        RECT 12.150000 1.300000 12.835000 1.780000 ;
        RECT 12.665000 1.130000 13.865000 1.275000 ;
        RECT 13.540000 1.300000 13.865000 1.550000 ;
    END
  END S1
  PIN X
    ANTENNADIFFAREA  1.086400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 14.875000 1.800000 16.675000 1.970000 ;
        RECT 14.875000 1.970000 15.205000 2.980000 ;
        RECT 15.065000 0.350000 15.315000 0.960000 ;
        RECT 15.065000 0.960000 16.675000 1.130000 ;
        RECT 15.825000 1.970000 16.155000 2.980000 ;
        RECT 15.925000 0.350000 16.175000 0.960000 ;
        RECT 16.445000 1.130000 16.675000 1.800000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 16.800000 0.085000 ;
        RECT  0.115000  0.085000  0.365000 1.030000 ;
        RECT  0.115000  1.030000  1.370000 1.280000 ;
        RECT  1.045000  0.640000  1.370000 1.030000 ;
        RECT  1.980000  0.085000  2.310000 0.450000 ;
        RECT  5.375000  0.085000  5.705000 1.130000 ;
        RECT  8.495000  0.085000  8.825000 0.410000 ;
        RECT  9.435000  0.085000  9.685000 0.750000 ;
        RECT 10.295000  0.085000 10.545000 1.030000 ;
        RECT 14.715000  0.085000 14.885000 1.130000 ;
        RECT 15.495000  0.085000 15.745000 0.790000 ;
        RECT 16.355000  0.085000 16.685000 0.790000 ;
      LAYER mcon ;
        RECT  0.155000 -0.085000  0.325000 0.085000 ;
        RECT  0.635000 -0.085000  0.805000 0.085000 ;
        RECT  1.115000 -0.085000  1.285000 0.085000 ;
        RECT  1.595000 -0.085000  1.765000 0.085000 ;
        RECT  2.075000 -0.085000  2.245000 0.085000 ;
        RECT  2.555000 -0.085000  2.725000 0.085000 ;
        RECT  3.035000 -0.085000  3.205000 0.085000 ;
        RECT  3.515000 -0.085000  3.685000 0.085000 ;
        RECT  3.995000 -0.085000  4.165000 0.085000 ;
        RECT  4.475000 -0.085000  4.645000 0.085000 ;
        RECT  4.955000 -0.085000  5.125000 0.085000 ;
        RECT  5.435000 -0.085000  5.605000 0.085000 ;
        RECT  5.915000 -0.085000  6.085000 0.085000 ;
        RECT  6.395000 -0.085000  6.565000 0.085000 ;
        RECT  6.875000 -0.085000  7.045000 0.085000 ;
        RECT  7.355000 -0.085000  7.525000 0.085000 ;
        RECT  7.835000 -0.085000  8.005000 0.085000 ;
        RECT  8.315000 -0.085000  8.485000 0.085000 ;
        RECT  8.795000 -0.085000  8.965000 0.085000 ;
        RECT  9.275000 -0.085000  9.445000 0.085000 ;
        RECT  9.755000 -0.085000  9.925000 0.085000 ;
        RECT 10.235000 -0.085000 10.405000 0.085000 ;
        RECT 10.715000 -0.085000 10.885000 0.085000 ;
        RECT 11.195000 -0.085000 11.365000 0.085000 ;
        RECT 11.675000 -0.085000 11.845000 0.085000 ;
        RECT 12.155000 -0.085000 12.325000 0.085000 ;
        RECT 12.635000 -0.085000 12.805000 0.085000 ;
        RECT 13.115000 -0.085000 13.285000 0.085000 ;
        RECT 13.595000 -0.085000 13.765000 0.085000 ;
        RECT 14.075000 -0.085000 14.245000 0.085000 ;
        RECT 14.555000 -0.085000 14.725000 0.085000 ;
        RECT 15.035000 -0.085000 15.205000 0.085000 ;
        RECT 15.515000 -0.085000 15.685000 0.085000 ;
        RECT 15.995000 -0.085000 16.165000 0.085000 ;
        RECT 16.475000 -0.085000 16.645000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 16.800000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 3.245000 16.800000 3.415000 ;
        RECT  0.115000 1.950000  0.365000 3.245000 ;
        RECT  1.095000 2.310000  1.345000 3.245000 ;
        RECT  2.045000 2.650000  2.295000 3.245000 ;
        RECT  5.400000 1.820000  5.730000 3.245000 ;
        RECT  8.320000 2.965000  8.650000 3.245000 ;
        RECT  9.390000 2.965000  9.730000 3.245000 ;
        RECT 10.465000 2.285000 10.635000 3.245000 ;
        RECT 14.375000 1.820000 14.705000 3.245000 ;
        RECT 15.405000 2.140000 15.655000 3.245000 ;
        RECT 16.325000 2.140000 16.655000 3.245000 ;
      LAYER mcon ;
        RECT  0.155000 3.245000  0.325000 3.415000 ;
        RECT  0.635000 3.245000  0.805000 3.415000 ;
        RECT  1.115000 3.245000  1.285000 3.415000 ;
        RECT  1.595000 3.245000  1.765000 3.415000 ;
        RECT  2.075000 3.245000  2.245000 3.415000 ;
        RECT  2.555000 3.245000  2.725000 3.415000 ;
        RECT  3.035000 3.245000  3.205000 3.415000 ;
        RECT  3.515000 3.245000  3.685000 3.415000 ;
        RECT  3.995000 3.245000  4.165000 3.415000 ;
        RECT  4.475000 3.245000  4.645000 3.415000 ;
        RECT  4.955000 3.245000  5.125000 3.415000 ;
        RECT  5.435000 3.245000  5.605000 3.415000 ;
        RECT  5.915000 3.245000  6.085000 3.415000 ;
        RECT  6.395000 3.245000  6.565000 3.415000 ;
        RECT  6.875000 3.245000  7.045000 3.415000 ;
        RECT  7.355000 3.245000  7.525000 3.415000 ;
        RECT  7.835000 3.245000  8.005000 3.415000 ;
        RECT  8.315000 3.245000  8.485000 3.415000 ;
        RECT  8.795000 3.245000  8.965000 3.415000 ;
        RECT  9.275000 3.245000  9.445000 3.415000 ;
        RECT  9.755000 3.245000  9.925000 3.415000 ;
        RECT 10.235000 3.245000 10.405000 3.415000 ;
        RECT 10.715000 3.245000 10.885000 3.415000 ;
        RECT 11.195000 3.245000 11.365000 3.415000 ;
        RECT 11.675000 3.245000 11.845000 3.415000 ;
        RECT 12.155000 3.245000 12.325000 3.415000 ;
        RECT 12.635000 3.245000 12.805000 3.415000 ;
        RECT 13.115000 3.245000 13.285000 3.415000 ;
        RECT 13.595000 3.245000 13.765000 3.415000 ;
        RECT 14.075000 3.245000 14.245000 3.415000 ;
        RECT 14.555000 3.245000 14.725000 3.415000 ;
        RECT 15.035000 3.245000 15.205000 3.415000 ;
        RECT 15.515000 3.245000 15.685000 3.415000 ;
        RECT 15.995000 3.245000 16.165000 3.415000 ;
        RECT 16.475000 3.245000 16.645000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 16.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.545000 0.275000  1.810000 0.470000 ;
      RECT  0.545000 0.470000  0.875000 0.860000 ;
      RECT  0.565000 1.950000  0.895000 1.970000 ;
      RECT  0.565000 1.970000  2.695000 2.140000 ;
      RECT  0.565000 2.140000  0.895000 2.980000 ;
      RECT  1.515000 2.310000  3.300000 2.480000 ;
      RECT  1.515000 2.480000  1.845000 2.980000 ;
      RECT  1.550000 0.960000  1.800000 1.130000 ;
      RECT  1.550000 1.130000  2.695000 1.260000 ;
      RECT  1.550000 1.260000  4.205000 1.300000 ;
      RECT  1.575000 0.470000  1.810000 0.620000 ;
      RECT  1.575000 0.620000  2.140000 0.790000 ;
      RECT  1.970000 0.790000  3.380000 0.960000 ;
      RECT  2.525000 1.300000  4.205000 1.430000 ;
      RECT  2.525000 1.600000  4.190000 1.770000 ;
      RECT  2.525000 1.770000  2.695000 1.970000 ;
      RECT  2.525000 2.650000  2.860000 2.905000 ;
      RECT  2.525000 2.905000  4.720000 3.075000 ;
      RECT  2.540000 0.255000  4.715000 0.425000 ;
      RECT  2.540000 0.425000  2.870000 0.620000 ;
      RECT  2.990000 1.940000  3.300000 2.310000 ;
      RECT  3.045000 2.480000  3.300000 2.735000 ;
      RECT  3.050000 0.595000  3.380000 0.790000 ;
      RECT  3.050000 0.960000  3.380000 1.090000 ;
      RECT  3.490000 1.940000  3.820000 2.905000 ;
      RECT  3.605000 0.425000  3.775000 1.090000 ;
      RECT  3.955000 0.595000  4.205000 1.260000 ;
      RECT  4.020000 1.770000  4.190000 2.735000 ;
      RECT  4.375000 0.425000  4.715000 1.180000 ;
      RECT  4.375000 1.180000  4.545000 1.920000 ;
      RECT  4.375000 1.920000  4.720000 2.905000 ;
      RECT  4.715000 1.350000  5.200000 1.365000 ;
      RECT  4.715000 1.365000  6.705000 1.535000 ;
      RECT  4.715000 1.535000  5.200000 1.680000 ;
      RECT  4.945000 0.350000  5.200000 1.350000 ;
      RECT  4.950000 1.680000  5.200000 2.980000 ;
      RECT  5.935000 0.585000  6.185000 1.025000 ;
      RECT  5.935000 1.025000  7.125000 1.195000 ;
      RECT  5.960000 1.865000  7.125000 1.945000 ;
      RECT  5.960000 1.945000 10.975000 2.035000 ;
      RECT  5.960000 2.035000  6.210000 2.905000 ;
      RECT  6.035000 1.535000  6.705000 1.695000 ;
      RECT  6.365000 0.255000  8.325000 0.425000 ;
      RECT  6.365000 0.425000  6.695000 0.855000 ;
      RECT  6.410000 2.205000  6.740000 2.905000 ;
      RECT  6.410000 2.905000  8.150000 3.075000 ;
      RECT  6.875000 0.595000  7.985000 0.765000 ;
      RECT  6.875000 0.765000  7.125000 1.025000 ;
      RECT  6.875000 1.195000  7.125000 1.265000 ;
      RECT  6.940000 1.265000  7.125000 1.865000 ;
      RECT  6.940000 2.035000 10.975000 2.115000 ;
      RECT  6.940000 2.115000  7.125000 2.735000 ;
      RECT  7.305000 0.935000  7.555000 1.095000 ;
      RECT  7.305000 1.095000  8.325000 1.265000 ;
      RECT  7.310000 2.285000  9.185000 2.455000 ;
      RECT  7.310000 2.455000  7.640000 2.735000 ;
      RECT  7.735000 0.765000  7.985000 0.925000 ;
      RECT  7.980000 2.625000 10.265000 2.795000 ;
      RECT  7.980000 2.795000  8.150000 2.905000 ;
      RECT  8.155000 0.425000  8.325000 0.580000 ;
      RECT  8.155000 0.580000  9.255000 0.750000 ;
      RECT  8.155000 0.920000 10.115000 1.090000 ;
      RECT  8.155000 1.090000  8.325000 1.095000 ;
      RECT  9.005000 0.350000  9.255000 0.580000 ;
      RECT  9.865000 0.350000 10.115000 0.920000 ;
      RECT  9.935000 2.285000 10.265000 2.625000 ;
      RECT  9.935000 2.795000 10.265000 2.980000 ;
      RECT 10.715000 0.255000 11.815000 0.425000 ;
      RECT 10.715000 0.425000 10.885000 1.945000 ;
      RECT 10.805000 2.115000 10.975000 2.905000 ;
      RECT 10.805000 2.905000 12.975000 3.075000 ;
      RECT 11.055000 0.595000 12.675000 0.620000 ;
      RECT 11.055000 0.620000 12.155000 0.765000 ;
      RECT 11.055000 0.765000 11.475000 1.030000 ;
      RECT 11.145000 1.030000 11.475000 2.565000 ;
      RECT 11.145000 2.565000 12.475000 2.735000 ;
      RECT 11.645000 0.935000 13.175000 0.960000 ;
      RECT 11.645000 0.960000 12.495000 1.105000 ;
      RECT 11.645000 1.105000 11.975000 2.395000 ;
      RECT 11.985000 0.255000 14.545000 0.425000 ;
      RECT 11.985000 0.425000 12.675000 0.595000 ;
      RECT 12.145000 1.950000 12.475000 2.060000 ;
      RECT 12.145000 2.060000 13.475000 2.230000 ;
      RECT 12.145000 2.230000 12.475000 2.565000 ;
      RECT 12.325000 0.790000 13.175000 0.935000 ;
      RECT 12.645000 2.400000 12.975000 2.905000 ;
      RECT 12.860000 0.595000 13.175000 0.790000 ;
      RECT 13.005000 1.470000 13.330000 1.720000 ;
      RECT 13.005000 1.720000 14.205000 1.890000 ;
      RECT 13.145000 2.230000 13.475000 2.980000 ;
      RECT 13.345000 0.425000 13.675000 0.960000 ;
      RECT 13.875000 1.890000 14.205000 2.980000 ;
      RECT 13.905000 0.595000 14.205000 0.960000 ;
      RECT 14.035000 0.960000 14.205000 1.720000 ;
      RECT 14.375000 0.425000 14.545000 1.300000 ;
      RECT 14.375000 1.300000 16.210000 1.630000 ;
    LAYER mcon ;
      RECT  4.475000 1.950000  4.645000 2.120000 ;
      RECT 11.675000 1.950000 11.845000 2.120000 ;
    LAYER met1 ;
      RECT  4.415000 1.920000  4.705000 1.965000 ;
      RECT  4.415000 1.965000 11.905000 2.105000 ;
      RECT  4.415000 2.105000  4.705000 2.150000 ;
      RECT 11.615000 1.920000 11.905000 1.965000 ;
      RECT 11.615000 2.105000 11.905000 2.150000 ;
  END
END sky130_fd_sc_ls__mux4_4
