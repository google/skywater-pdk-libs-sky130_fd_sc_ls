* File: sky130_fd_sc_ls__and3b_4.spice
* Created: Fri Aug 28 13:04:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__and3b_4.pex.spice"
.subckt sky130_fd_sc_ls__and3b_4  VNB VPB A_N B C VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* C	C
* B	B
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1019 N_VGND_M1019_d N_A_N_M1019_g N_A_27_74#_M1019_s VNB NSHORT L=0.15 W=0.64
+ AD=0.1888 AS=0.1824 PD=1.87 PS=1.85 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1000 N_A_239_98#_M1000_d N_A_27_74#_M1000_g N_A_298_368#_M1000_s VNB NSHORT
+ L=0.15 W=0.64 AD=0.1824 AS=0.0896 PD=1.85 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1018 N_A_239_98#_M1018_d N_A_27_74#_M1018_g N_A_298_368#_M1000_s VNB NSHORT
+ L=0.15 W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1014 N_A_239_98#_M1018_d N_B_M1014_g N_A_498_98#_M1014_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.112 PD=0.92 PS=0.99 NRD=0 NRS=13.116 M=1 R=4.26667
+ SA=75001.1 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1015 N_A_239_98#_M1015_d N_B_M1015_g N_A_498_98#_M1014_s VNB NSHORT L=0.15
+ W=0.64 AD=0.1824 AS=0.112 PD=1.85 PS=0.99 NRD=0 NRS=0 M=1 R=4.26667 SA=75001.6
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1002 N_A_498_98#_M1002_d N_C_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.1824 PD=0.92 PS=1.85 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75002.5 A=0.096 P=1.58 MULT=1
MM1012 N_A_498_98#_M1002_d N_C_M1012_g N_VGND_M1012_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.12007 PD=0.92 PS=1.02029 NRD=0 NRS=15.468 M=1 R=4.26667
+ SA=75000.6 SB=75002.1 A=0.096 P=1.58 MULT=1
MM1003 N_VGND_M1012_s N_A_298_368#_M1003_g N_X_M1003_s VNB NSHORT L=0.15 W=0.74
+ AD=0.13883 AS=0.1295 PD=1.17971 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1007 N_VGND_M1007_d N_A_298_368#_M1007_g N_X_M1003_s VNB NSHORT L=0.15 W=0.74
+ AD=0.111 AS=0.1295 PD=1.04 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1010 N_VGND_M1007_d N_A_298_368#_M1010_g N_X_M1010_s VNB NSHORT L=0.15 W=0.74
+ AD=0.111 AS=0.1036 PD=1.04 PS=1.02 NRD=3.24 NRS=0 M=1 R=4.93333 SA=75002
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1016 N_VGND_M1016_d N_A_298_368#_M1016_g N_X_M1010_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.4
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1013 N_VPWR_M1013_d N_A_N_M1013_g N_A_27_74#_M1013_s VPB PHIGHVT L=0.15 W=1
+ AD=0.2 AS=0.295 PD=1.4 PS=2.59 NRD=11.8003 NRS=1.9503 M=1 R=6.66667 SA=75000.2
+ SB=75005.4 A=0.15 P=2.3 MULT=1
MM1017 N_A_298_368#_M1017_d N_A_27_74#_M1017_g N_VPWR_M1013_d VPB PHIGHVT L=0.15
+ W=1 AD=0.15 AS=0.2 PD=1.3 PS=1.4 NRD=1.9503 NRS=11.8003 M=1 R=6.66667
+ SA=75000.8 SB=75004.8 A=0.15 P=2.3 MULT=1
MM1020 N_A_298_368#_M1017_d N_A_27_74#_M1020_g N_VPWR_M1020_s VPB PHIGHVT L=0.15
+ W=1 AD=0.15 AS=0.2 PD=1.3 PS=1.4 NRD=1.9503 NRS=11.8003 M=1 R=6.66667
+ SA=75001.2 SB=75004.4 A=0.15 P=2.3 MULT=1
MM1001 N_A_298_368#_M1001_d N_B_M1001_g N_VPWR_M1020_s VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.2 PD=1.3 PS=1.4 NRD=1.9503 NRS=11.8003 M=1 R=6.66667 SA=75001.8
+ SB=75003.8 A=0.15 P=2.3 MULT=1
MM1008 N_A_298_368#_M1001_d N_B_M1008_g N_VPWR_M1008_s VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.23 PD=1.3 PS=1.46 NRD=1.9503 NRS=11.8003 M=1 R=6.66667 SA=75002.2
+ SB=75003.4 A=0.15 P=2.3 MULT=1
MM1004 N_A_298_368#_M1004_d N_C_M1004_g N_VPWR_M1008_s VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.23 PD=1.3 PS=1.46 NRD=1.9503 NRS=23.6203 M=1 R=6.66667 SA=75002.8
+ SB=75002.8 A=0.15 P=2.3 MULT=1
MM1009 N_A_298_368#_M1004_d N_C_M1009_g N_VPWR_M1009_s VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.224717 PD=1.3 PS=1.46698 NRD=1.9503 NRS=19.0302 M=1 R=6.66667
+ SA=75003.3 SB=75002.3 A=0.15 P=2.3 MULT=1
MM1005 N_VPWR_M1009_s N_A_298_368#_M1005_g N_X_M1005_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.251683 AS=0.168 PD=1.64302 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75003.5 SB=75001.7 A=0.168 P=2.54 MULT=1
MM1006 N_VPWR_M1006_d N_A_298_368#_M1006_g N_X_M1005_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.224 AS=0.168 PD=1.52 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75003.9 SB=75001.3 A=0.168 P=2.54 MULT=1
MM1011 N_VPWR_M1006_d N_A_298_368#_M1011_g N_X_M1011_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.224 AS=0.168 PD=1.52 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75004.5 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1021 N_VPWR_M1021_d N_A_298_368#_M1021_g N_X_M1011_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3864 AS=0.168 PD=2.93 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75004.9 SB=75000.3 A=0.168 P=2.54 MULT=1
DX22_noxref VNB VPB NWDIODE A=13.206 P=17.92
*
.include "sky130_fd_sc_ls__and3b_4.pxi.spice"
*
.ends
*
*
