* File: sky130_fd_sc_ls__and3_1.pxi.spice
* Created: Wed Sep  2 10:54:45 2020
* 
x_PM_SKY130_FD_SC_LS__AND3_1%A N_A_c_54_n N_A_c_62_n N_A_M1006_g N_A_c_55_n
+ N_A_M1001_g N_A_c_57_n N_A_c_58_n A N_A_c_60_n PM_SKY130_FD_SC_LS__AND3_1%A
x_PM_SKY130_FD_SC_LS__AND3_1%B N_B_c_98_n N_B_M1004_g N_B_c_99_n N_B_M1002_g B B
+ PM_SKY130_FD_SC_LS__AND3_1%B
x_PM_SKY130_FD_SC_LS__AND3_1%C N_C_c_138_n N_C_M1000_g N_C_M1003_g C
+ PM_SKY130_FD_SC_LS__AND3_1%C
x_PM_SKY130_FD_SC_LS__AND3_1%A_27_398# N_A_27_398#_M1001_s N_A_27_398#_M1006_s
+ N_A_27_398#_M1004_d N_A_27_398#_c_170_n N_A_27_398#_M1007_g
+ N_A_27_398#_c_171_n N_A_27_398#_M1005_g N_A_27_398#_c_172_n
+ N_A_27_398#_c_176_n N_A_27_398#_c_177_n N_A_27_398#_c_178_n
+ N_A_27_398#_c_179_n N_A_27_398#_c_180_n N_A_27_398#_c_181_n
+ N_A_27_398#_c_182_n N_A_27_398#_c_173_n PM_SKY130_FD_SC_LS__AND3_1%A_27_398#
x_PM_SKY130_FD_SC_LS__AND3_1%VPWR N_VPWR_M1006_d N_VPWR_M1000_d N_VPWR_c_243_n
+ N_VPWR_c_244_n VPWR N_VPWR_c_245_n N_VPWR_c_246_n N_VPWR_c_247_n
+ N_VPWR_c_242_n N_VPWR_c_249_n N_VPWR_c_250_n PM_SKY130_FD_SC_LS__AND3_1%VPWR
x_PM_SKY130_FD_SC_LS__AND3_1%X N_X_M1007_d N_X_M1005_d N_X_c_280_n N_X_c_281_n X
+ X X X N_X_c_282_n PM_SKY130_FD_SC_LS__AND3_1%X
x_PM_SKY130_FD_SC_LS__AND3_1%VGND N_VGND_M1003_d N_VGND_c_304_n N_VGND_c_305_n
+ N_VGND_c_306_n VGND N_VGND_c_307_n N_VGND_c_308_n
+ PM_SKY130_FD_SC_LS__AND3_1%VGND
cc_1 VNB N_A_c_54_n 0.00748651f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.825
cc_2 VNB N_A_c_55_n 0.0397668f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=0.57
cc_3 VNB N_A_M1001_g 0.0144312f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1
cc_4 VNB N_A_c_57_n 0.0116107f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.545
cc_5 VNB N_A_c_58_n 0.0424882f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.405
cc_6 VNB A 0.00759927f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=0.47
cc_7 VNB N_A_c_60_n 0.0208892f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=0.462
cc_8 VNB N_B_c_98_n 0.0200688f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_B_c_99_n 0.016463f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.825
cc_10 VNB B 0.00357895f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.41
cc_11 VNB N_C_c_138_n 0.025422f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_C_M1003_g 0.0258025f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.41
cc_13 VNB C 0.00338947f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=0.57
cc_14 VNB N_A_27_398#_c_170_n 0.0220597f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1
cc_15 VNB N_A_27_398#_c_171_n 0.0336918f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.545
cc_16 VNB N_A_27_398#_c_172_n 0.0376576f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_27_398#_c_173_n 0.00166255f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_VPWR_c_242_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_X_c_280_n 0.0234698f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.395
cc_20 VNB N_X_c_281_n 0.0184679f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.412
cc_21 VNB N_X_c_282_n 0.023805f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_304_n 0.0191361f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.41
cc_23 VNB N_VGND_c_305_n 0.0444379f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1
cc_24 VNB N_VGND_c_306_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.395
cc_25 VNB N_VGND_c_307_n 0.0273666f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=0.462
cc_26 VNB N_VGND_c_308_n 0.202229f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VPB N_A_c_54_n 0.0110573f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.825
cc_28 VPB N_A_c_62_n 0.02682f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.915
cc_29 VPB N_B_c_98_n 0.0361793f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_30 VPB B 0.00357649f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.41
cc_31 VPB N_C_c_138_n 0.0428825f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_32 VPB C 0.00203124f $X=-0.19 $Y=1.66 $X2=0.53 $Y2=0.57
cc_33 VPB N_A_27_398#_c_171_n 0.0358952f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.545
cc_34 VPB N_A_27_398#_c_172_n 0.0121764f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_35 VPB N_A_27_398#_c_176_n 0.0311015f $X=-0.19 $Y=1.66 $X2=1.2 $Y2=0.462
cc_36 VPB N_A_27_398#_c_177_n 0.00939188f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_37 VPB N_A_27_398#_c_178_n 0.00302721f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_38 VPB N_A_27_398#_c_179_n 0.00992738f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_39 VPB N_A_27_398#_c_180_n 0.00264418f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_40 VPB N_A_27_398#_c_181_n 0.00719737f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_41 VPB N_A_27_398#_c_182_n 0.00507919f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_42 VPB N_A_27_398#_c_173_n 7.30623e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_43 VPB N_VPWR_c_243_n 0.0170624f $X=-0.19 $Y=1.66 $X2=0.53 $Y2=1.395
cc_44 VPB N_VPWR_c_244_n 0.0097445f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.545
cc_45 VPB N_VPWR_c_245_n 0.0197293f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=0.405
cc_46 VPB N_VPWR_c_246_n 0.0181128f $X=-0.19 $Y=1.66 $X2=1.2 $Y2=0.462
cc_47 VPB N_VPWR_c_247_n 0.017913f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_242_n 0.0658592f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_249_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_250_n 0.0140321f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_51 VPB X 0.00529771f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=0.405
cc_52 VPB X 0.0395498f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_X_c_282_n 0.00896137f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 N_A_c_54_n N_B_c_98_n 0.0156729f $X=0.505 $Y=1.825 $X2=-0.19 $Y2=-0.245
cc_55 N_A_c_62_n N_B_c_98_n 0.0240203f $X=0.505 $Y=1.915 $X2=-0.19 $Y2=-0.245
cc_56 N_A_c_57_n N_B_c_98_n 0.00587736f $X=0.51 $Y=1.545 $X2=-0.19 $Y2=-0.245
cc_57 N_A_c_55_n N_B_c_99_n 0.0011105f $X=0.53 $Y=0.57 $X2=0 $Y2=0
cc_58 N_A_M1001_g N_B_c_99_n 0.0251307f $X=0.53 $Y=1 $X2=0 $Y2=0
cc_59 A N_B_c_99_n 0.00718878f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_60 N_A_c_60_n N_B_c_99_n 0.00365215f $X=1.085 $Y=0.462 $X2=0 $Y2=0
cc_61 N_A_c_54_n B 9.39698e-19 $X=0.505 $Y=1.825 $X2=0 $Y2=0
cc_62 N_A_M1001_g B 0.00222717f $X=0.53 $Y=1 $X2=0 $Y2=0
cc_63 N_A_c_57_n B 4.14418e-19 $X=0.51 $Y=1.545 $X2=0 $Y2=0
cc_64 A B 0.00728026f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_65 N_A_c_60_n B 0.00666142f $X=1.085 $Y=0.462 $X2=0 $Y2=0
cc_66 N_A_c_55_n N_C_M1003_g 7.00286e-19 $X=0.53 $Y=0.57 $X2=0 $Y2=0
cc_67 A N_C_M1003_g 0.00212205f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_68 N_A_c_54_n N_A_27_398#_c_172_n 0.01082f $X=0.505 $Y=1.825 $X2=0 $Y2=0
cc_69 N_A_c_62_n N_A_27_398#_c_172_n 0.00569875f $X=0.505 $Y=1.915 $X2=0 $Y2=0
cc_70 N_A_M1001_g N_A_27_398#_c_172_n 0.0179899f $X=0.53 $Y=1 $X2=0 $Y2=0
cc_71 N_A_c_57_n N_A_27_398#_c_172_n 0.00669835f $X=0.51 $Y=1.545 $X2=0 $Y2=0
cc_72 N_A_c_58_n N_A_27_398#_c_172_n 0.00770329f $X=0.61 $Y=0.405 $X2=0 $Y2=0
cc_73 N_A_c_60_n N_A_27_398#_c_172_n 0.0263323f $X=1.085 $Y=0.462 $X2=0 $Y2=0
cc_74 N_A_c_62_n N_A_27_398#_c_176_n 0.0125247f $X=0.505 $Y=1.915 $X2=0 $Y2=0
cc_75 N_A_c_62_n N_A_27_398#_c_177_n 0.0136156f $X=0.505 $Y=1.915 $X2=0 $Y2=0
cc_76 N_A_c_57_n N_A_27_398#_c_177_n 3.2368e-19 $X=0.51 $Y=1.545 $X2=0 $Y2=0
cc_77 N_A_c_62_n N_A_27_398#_c_178_n 6.37908e-19 $X=0.505 $Y=1.915 $X2=0 $Y2=0
cc_78 N_A_c_62_n N_A_27_398#_c_181_n 0.0033471f $X=0.505 $Y=1.915 $X2=0 $Y2=0
cc_79 N_A_c_62_n N_VPWR_c_243_n 0.0066275f $X=0.505 $Y=1.915 $X2=0 $Y2=0
cc_80 N_A_c_62_n N_VPWR_c_245_n 0.00475875f $X=0.505 $Y=1.915 $X2=0 $Y2=0
cc_81 N_A_c_62_n N_VPWR_c_242_n 0.00505379f $X=0.505 $Y=1.915 $X2=0 $Y2=0
cc_82 A A_233_136# 0.00220589f $X=1.115 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_83 A N_VGND_c_304_n 0.0186975f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_84 N_A_c_58_n N_VGND_c_305_n 0.0116176f $X=0.61 $Y=0.405 $X2=0 $Y2=0
cc_85 N_A_c_60_n N_VGND_c_305_n 0.0795377f $X=1.085 $Y=0.462 $X2=0 $Y2=0
cc_86 N_A_c_55_n N_VGND_c_308_n 0.0073025f $X=0.53 $Y=0.57 $X2=0 $Y2=0
cc_87 N_A_c_58_n N_VGND_c_308_n 0.00773969f $X=0.61 $Y=0.405 $X2=0 $Y2=0
cc_88 N_A_c_60_n N_VGND_c_308_n 0.043082f $X=1.085 $Y=0.462 $X2=0 $Y2=0
cc_89 N_B_c_98_n N_C_c_138_n 0.0385814f $X=1.055 $Y=1.915 $X2=-0.19 $Y2=-0.245
cc_90 B N_C_c_138_n 0.00244375f $X=1.115 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_91 N_B_c_98_n N_C_M1003_g 6.80675e-19 $X=1.055 $Y=1.915 $X2=0 $Y2=0
cc_92 N_B_c_99_n N_C_M1003_g 0.0325782f $X=1.09 $Y=1.43 $X2=0 $Y2=0
cc_93 B N_C_M1003_g 0.0068958f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_94 N_B_c_98_n C 2.8986e-19 $X=1.055 $Y=1.915 $X2=0 $Y2=0
cc_95 B C 0.0268673f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_96 N_B_c_98_n N_A_27_398#_c_172_n 0.00185671f $X=1.055 $Y=1.915 $X2=0 $Y2=0
cc_97 N_B_c_99_n N_A_27_398#_c_172_n 0.00223336f $X=1.09 $Y=1.43 $X2=0 $Y2=0
cc_98 B N_A_27_398#_c_172_n 0.0261437f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_99 N_B_c_98_n N_A_27_398#_c_176_n 6.37052e-19 $X=1.055 $Y=1.915 $X2=0 $Y2=0
cc_100 N_B_c_98_n N_A_27_398#_c_177_n 0.0136649f $X=1.055 $Y=1.915 $X2=0 $Y2=0
cc_101 B N_A_27_398#_c_177_n 0.0212746f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_102 N_B_c_98_n N_A_27_398#_c_178_n 0.0107366f $X=1.055 $Y=1.915 $X2=0 $Y2=0
cc_103 N_B_c_98_n N_A_27_398#_c_182_n 0.0016299f $X=1.055 $Y=1.915 $X2=0 $Y2=0
cc_104 B N_A_27_398#_c_182_n 0.0182697f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_105 N_B_c_98_n N_VPWR_c_243_n 0.0051685f $X=1.055 $Y=1.915 $X2=0 $Y2=0
cc_106 N_B_c_98_n N_VPWR_c_244_n 5.47572e-19 $X=1.055 $Y=1.915 $X2=0 $Y2=0
cc_107 N_B_c_98_n N_VPWR_c_246_n 0.00475875f $X=1.055 $Y=1.915 $X2=0 $Y2=0
cc_108 N_B_c_98_n N_VPWR_c_242_n 0.00505379f $X=1.055 $Y=1.915 $X2=0 $Y2=0
cc_109 B A_121_136# 0.00405918f $X=1.115 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_110 B A_233_136# 0.00359387f $X=1.115 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_111 N_B_c_99_n N_VGND_c_305_n 4.93445e-19 $X=1.09 $Y=1.43 $X2=0 $Y2=0
cc_112 N_C_M1003_g N_A_27_398#_c_170_n 0.0219279f $X=1.565 $Y=0.92 $X2=0 $Y2=0
cc_113 N_C_c_138_n N_A_27_398#_c_171_n 0.0194417f $X=1.505 $Y=1.915 $X2=0 $Y2=0
cc_114 C N_A_27_398#_c_171_n 8.96262e-19 $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_115 N_C_c_138_n N_A_27_398#_c_178_n 9.10391e-19 $X=1.505 $Y=1.915 $X2=0 $Y2=0
cc_116 N_C_c_138_n N_A_27_398#_c_179_n 0.018913f $X=1.505 $Y=1.915 $X2=0 $Y2=0
cc_117 C N_A_27_398#_c_179_n 0.0244211f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_118 N_C_c_138_n N_A_27_398#_c_180_n 0.00369081f $X=1.505 $Y=1.915 $X2=0 $Y2=0
cc_119 N_C_c_138_n N_A_27_398#_c_173_n 8.98411e-19 $X=1.505 $Y=1.915 $X2=0 $Y2=0
cc_120 N_C_M1003_g N_A_27_398#_c_173_n 5.59322e-19 $X=1.565 $Y=0.92 $X2=0 $Y2=0
cc_121 C N_A_27_398#_c_173_n 0.0180069f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_122 N_C_c_138_n N_VPWR_c_244_n 0.0155788f $X=1.505 $Y=1.915 $X2=0 $Y2=0
cc_123 N_C_c_138_n N_VPWR_c_246_n 0.00454039f $X=1.505 $Y=1.915 $X2=0 $Y2=0
cc_124 N_C_c_138_n N_VPWR_c_242_n 0.00475056f $X=1.505 $Y=1.915 $X2=0 $Y2=0
cc_125 N_C_c_138_n N_VGND_c_304_n 8.79027e-19 $X=1.505 $Y=1.915 $X2=0 $Y2=0
cc_126 N_C_M1003_g N_VGND_c_304_n 0.00515513f $X=1.565 $Y=0.92 $X2=0 $Y2=0
cc_127 C N_VGND_c_304_n 0.00681967f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_128 N_C_M1003_g N_VGND_c_305_n 0.00428744f $X=1.565 $Y=0.92 $X2=0 $Y2=0
cc_129 N_C_M1003_g N_VGND_c_308_n 0.00476395f $X=1.565 $Y=0.92 $X2=0 $Y2=0
cc_130 N_A_27_398#_c_177_n N_VPWR_M1006_d 0.00332584f $X=1.115 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_131 N_A_27_398#_c_179_n N_VPWR_M1000_d 0.0132146f $X=2.07 $Y=2.035 $X2=0
+ $Y2=0
cc_132 N_A_27_398#_c_180_n N_VPWR_M1000_d 0.00350977f $X=2.155 $Y=1.95 $X2=0
+ $Y2=0
cc_133 N_A_27_398#_c_176_n N_VPWR_c_243_n 0.021803f $X=0.28 $Y=2.135 $X2=0 $Y2=0
cc_134 N_A_27_398#_c_177_n N_VPWR_c_243_n 0.0232685f $X=1.115 $Y=2.035 $X2=0
+ $Y2=0
cc_135 N_A_27_398#_c_178_n N_VPWR_c_243_n 0.0213364f $X=1.28 $Y=2.135 $X2=0
+ $Y2=0
cc_136 N_A_27_398#_c_171_n N_VPWR_c_244_n 0.0167782f $X=2.375 $Y=1.765 $X2=0
+ $Y2=0
cc_137 N_A_27_398#_c_178_n N_VPWR_c_244_n 0.0242512f $X=1.28 $Y=2.135 $X2=0
+ $Y2=0
cc_138 N_A_27_398#_c_179_n N_VPWR_c_244_n 0.0510726f $X=2.07 $Y=2.035 $X2=0
+ $Y2=0
cc_139 N_A_27_398#_c_173_n N_VPWR_c_244_n 0.00107051f $X=2.235 $Y=1.515 $X2=0
+ $Y2=0
cc_140 N_A_27_398#_c_176_n N_VPWR_c_245_n 0.00953144f $X=0.28 $Y=2.135 $X2=0
+ $Y2=0
cc_141 N_A_27_398#_c_178_n N_VPWR_c_246_n 0.00821887f $X=1.28 $Y=2.135 $X2=0
+ $Y2=0
cc_142 N_A_27_398#_c_171_n N_VPWR_c_247_n 0.00429299f $X=2.375 $Y=1.765 $X2=0
+ $Y2=0
cc_143 N_A_27_398#_c_171_n N_VPWR_c_242_n 0.00851215f $X=2.375 $Y=1.765 $X2=0
+ $Y2=0
cc_144 N_A_27_398#_c_176_n N_VPWR_c_242_n 0.0111133f $X=0.28 $Y=2.135 $X2=0
+ $Y2=0
cc_145 N_A_27_398#_c_178_n N_VPWR_c_242_n 0.00958658f $X=1.28 $Y=2.135 $X2=0
+ $Y2=0
cc_146 N_A_27_398#_c_170_n N_X_c_280_n 0.00624223f $X=2.145 $Y=1.35 $X2=0 $Y2=0
cc_147 N_A_27_398#_c_170_n N_X_c_281_n 0.00220367f $X=2.145 $Y=1.35 $X2=0 $Y2=0
cc_148 N_A_27_398#_c_171_n N_X_c_281_n 0.00382434f $X=2.375 $Y=1.765 $X2=0 $Y2=0
cc_149 N_A_27_398#_c_173_n N_X_c_281_n 0.0131627f $X=2.235 $Y=1.515 $X2=0 $Y2=0
cc_150 N_A_27_398#_c_171_n X 8.50339e-19 $X=2.375 $Y=1.765 $X2=0 $Y2=0
cc_151 N_A_27_398#_c_170_n N_X_c_282_n 0.00426097f $X=2.145 $Y=1.35 $X2=0 $Y2=0
cc_152 N_A_27_398#_c_171_n N_X_c_282_n 0.0117648f $X=2.375 $Y=1.765 $X2=0 $Y2=0
cc_153 N_A_27_398#_c_180_n N_X_c_282_n 0.00759252f $X=2.155 $Y=1.95 $X2=0 $Y2=0
cc_154 N_A_27_398#_c_173_n N_X_c_282_n 0.0223685f $X=2.235 $Y=1.515 $X2=0 $Y2=0
cc_155 N_A_27_398#_c_170_n N_VGND_c_304_n 0.0089425f $X=2.145 $Y=1.35 $X2=0
+ $Y2=0
cc_156 N_A_27_398#_c_170_n N_VGND_c_307_n 0.00467453f $X=2.145 $Y=1.35 $X2=0
+ $Y2=0
cc_157 N_A_27_398#_c_170_n N_VGND_c_308_n 0.00505379f $X=2.145 $Y=1.35 $X2=0
+ $Y2=0
cc_158 N_VPWR_c_244_n X 0.0297014f $X=2.145 $Y=2.375 $X2=0 $Y2=0
cc_159 N_VPWR_c_247_n X 0.0126277f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_160 N_VPWR_c_242_n X 0.0104521f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_161 N_X_c_280_n N_VGND_c_304_n 0.0206774f $X=2.36 $Y=0.645 $X2=0 $Y2=0
cc_162 N_X_c_280_n N_VGND_c_307_n 0.0093375f $X=2.36 $Y=0.645 $X2=0 $Y2=0
cc_163 N_X_c_280_n N_VGND_c_308_n 0.0109911f $X=2.36 $Y=0.645 $X2=0 $Y2=0
