* NGSPICE file created from sky130_fd_sc_ls__nand4bb_2.ext - technology: sky130A

.subckt sky130_fd_sc_ls__nand4bb_2 A_N B_N C D VGND VNB VPB VPWR Y
M1000 a_373_74# a_231_74# a_678_74# VNB nshort w=740000u l=150000u
+  ad=8.504e+11p pd=6.86e+06u as=4.662e+11p ps=4.22e+06u
M1001 Y a_231_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=1.3888e+12p pd=1.144e+07u as=3.0381e+12p ps=1.88e+07u
M1002 a_231_74# B_N VGND VNB nshort w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=5.278e+11p ps=4.3e+06u
M1003 a_886_74# D VGND VNB nshort w=740000u l=150000u
+  ad=6.29e+11p pd=6.14e+06u as=0p ps=0u
M1004 Y C VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND D a_886_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR C Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR a_231_74# Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_373_74# a_27_368# Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.257e+11p ps=2.09e+06u
M1009 Y D VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_231_74# B_N VPWR VPB phighvt w=1e+06u l=150000u
+  ad=3.95e+11p pd=2.79e+06u as=0p ps=0u
M1011 VPWR A_N a_27_368# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.95e+11p ps=2.59e+06u
M1012 Y a_27_368# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_886_74# C a_678_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_678_74# a_231_74# a_373_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR D Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Y a_27_368# a_373_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR a_27_368# Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND A_N a_27_368# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1019 a_678_74# C a_886_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

