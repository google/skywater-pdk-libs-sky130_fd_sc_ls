* File: sky130_fd_sc_ls__xnor2_2.pex.spice
* Created: Wed Sep  2 11:30:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__XNOR2_2%A 1 3 4 6 7 9 10 12 13 15 18 21 22 23 24 26
+ 27 33 34 38
c143 33 0 7.93433e-20 $X=3.12 $Y=1.295
c144 26 0 1.97825e-19 $X=2.975 $Y=1.295
c145 23 0 4.30741e-20 $X=3.355 $Y=1.805
r146 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.69
+ $Y=1.515 $X2=4.69 $Y2=1.515
r147 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.59
+ $Y=1.385 $X2=0.59 $Y2=1.385
r148 34 50 8.44752 $w=3.48e-07 $l=2.55e-07 $layer=LI1_cond $X=3.18 $Y=1.295
+ $X2=3.18 $Y2=1.55
r149 34 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.19
+ $Y=1.385 $X2=3.19 $Y2=1.385
r150 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=1.295
+ $X2=3.12 $Y2=1.295
r151 29 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=1.295
+ $X2=0.72 $Y2=1.295
r152 27 29 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.865 $Y=1.295
+ $X2=0.72 $Y2=1.295
r153 26 33 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.975 $Y=1.295
+ $X2=3.12 $Y2=1.295
r154 26 27 2.61138 $w=1.4e-07 $l=2.11e-06 $layer=MET1_cond $X=2.975 $Y=1.295
+ $X2=0.865 $Y2=1.295
r155 24 54 5.02353 $w=3.4e-07 $l=1.4e-07 $layer=LI1_cond $X=4.65 $Y=1.665
+ $X2=4.65 $Y2=1.805
r156 24 44 5.38235 $w=3.4e-07 $l=1.5e-07 $layer=LI1_cond $X=4.65 $Y=1.665
+ $X2=4.65 $Y2=1.515
r157 22 54 4.80115 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=4.445 $Y=1.805
+ $X2=4.65 $Y2=1.805
r158 22 23 71.1123 $w=1.68e-07 $l=1.09e-06 $layer=LI1_cond $X=4.445 $Y=1.805
+ $X2=3.355 $Y2=1.805
r159 21 23 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.19 $Y=1.72
+ $X2=3.355 $Y2=1.805
r160 21 50 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=3.19 $Y=1.72
+ $X2=3.19 $Y2=1.55
r161 16 43 38.5416 $w=3.03e-07 $l=2.06325e-07 $layer=POLY_cond $X=4.785 $Y=1.35
+ $X2=4.692 $Y2=1.515
r162 16 18 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.785 $Y=1.35
+ $X2=4.785 $Y2=0.74
r163 13 43 52.063 $w=3.03e-07 $l=2.51496e-07 $layer=POLY_cond $X=4.695 $Y=1.765
+ $X2=4.692 $Y2=1.515
r164 13 15 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.695 $Y=1.765
+ $X2=4.695 $Y2=2.4
r165 10 40 38.9026 $w=2.7e-07 $l=1.90526e-07 $layer=POLY_cond $X=3.135 $Y=1.22
+ $X2=3.19 $Y2=1.385
r166 10 12 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.135 $Y=1.22
+ $X2=3.135 $Y2=0.74
r167 7 40 77.2841 $w=2.7e-07 $l=4.15812e-07 $layer=POLY_cond $X=3.115 $Y=1.765
+ $X2=3.19 $Y2=1.385
r168 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.115 $Y=1.765
+ $X2=3.115 $Y2=2.4
r169 4 37 38.9026 $w=2.7e-07 $l=2.05122e-07 $layer=POLY_cond $X=0.68 $Y=1.22
+ $X2=0.59 $Y2=1.385
r170 4 6 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.68 $Y=1.22 $X2=0.68
+ $Y2=0.74
r171 1 37 77.2841 $w=2.7e-07 $l=3.8e-07 $layer=POLY_cond $X=0.59 $Y=1.765
+ $X2=0.59 $Y2=1.385
r172 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.59 $Y=1.765
+ $X2=0.59 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_LS__XNOR2_2%B 3 5 7 8 10 11 13 14 16 17 19 21 24 25 27
+ 28 30 31 32 33 34 36 38 47
c151 31 0 1.11424e-19 $X=5.025 $Y=2.145
c152 21 0 1.97825e-19 $X=1.085 $Y=1.557
r153 47 48 1.65446 $w=4.37e-07 $l=1.5e-08 $layer=POLY_cond $X=4.18 $Y=1.492
+ $X2=4.195 $Y2=1.492
r154 45 47 9.92677 $w=4.37e-07 $l=9e-08 $layer=POLY_cond $X=4.09 $Y=1.492
+ $X2=4.18 $Y2=1.492
r155 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.09
+ $Y=1.385 $X2=4.09 $Y2=1.385
r156 43 45 38.0526 $w=4.37e-07 $l=3.45e-07 $layer=POLY_cond $X=3.745 $Y=1.492
+ $X2=4.09 $Y2=1.492
r157 42 43 1.65446 $w=4.37e-07 $l=1.5e-08 $layer=POLY_cond $X=3.73 $Y=1.492
+ $X2=3.745 $Y2=1.492
r158 38 46 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=4.09 $Y=1.295
+ $X2=4.09 $Y2=1.385
r159 37 38 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=4.09 $Y=1.18
+ $X2=4.09 $Y2=1.295
r160 35 36 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=5.11 $Y=1.18
+ $X2=5.11 $Y2=2.06
r161 34 37 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.255 $Y=1.095
+ $X2=4.09 $Y2=1.18
r162 33 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.025 $Y=1.095
+ $X2=5.11 $Y2=1.18
r163 33 34 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=5.025 $Y=1.095
+ $X2=4.255 $Y2=1.095
r164 31 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.025 $Y=2.145
+ $X2=5.11 $Y2=2.06
r165 31 32 146.791 $w=1.68e-07 $l=2.25e-06 $layer=LI1_cond $X=5.025 $Y=2.145
+ $X2=2.775 $Y2=2.145
r166 30 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.69 $Y=2.06
+ $X2=2.775 $Y2=2.145
r167 29 30 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.69 $Y=1.89
+ $X2=2.69 $Y2=2.06
r168 27 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.605 $Y=1.805
+ $X2=2.69 $Y2=1.89
r169 27 28 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=2.605 $Y=1.805
+ $X2=1.675 $Y2=1.805
r170 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.51
+ $Y=1.515 $X2=1.51 $Y2=1.515
r171 22 28 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.51 $Y=1.72
+ $X2=1.675 $Y2=1.805
r172 22 24 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=1.51 $Y=1.72
+ $X2=1.51 $Y2=1.515
r173 20 25 58.5785 $w=3.3e-07 $l=3.35e-07 $layer=POLY_cond $X=1.175 $Y=1.515
+ $X2=1.51 $Y2=1.515
r174 20 21 5.03009 $w=3.3e-07 $l=1.08995e-07 $layer=POLY_cond $X=1.175 $Y=1.515
+ $X2=1.085 $Y2=1.557
r175 17 48 28.039 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=4.195 $Y=1.765
+ $X2=4.195 $Y2=1.492
r176 17 19 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.195 $Y=1.765
+ $X2=4.195 $Y2=2.4
r177 14 47 28.039 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=4.18 $Y=1.22
+ $X2=4.18 $Y2=1.492
r178 14 16 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.18 $Y=1.22
+ $X2=4.18 $Y2=0.74
r179 11 43 28.039 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=3.745 $Y=1.765
+ $X2=3.745 $Y2=1.492
r180 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.745 $Y=1.765
+ $X2=3.745 $Y2=2.4
r181 8 42 28.039 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=3.73 $Y=1.22
+ $X2=3.73 $Y2=1.492
r182 8 10 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.73 $Y=1.22 $X2=3.73
+ $Y2=0.74
r183 5 21 37.0704 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.085 $Y=1.765
+ $X2=1.085 $Y2=1.557
r184 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.085 $Y=1.765
+ $X2=1.085 $Y2=2.34
r185 1 21 37.0704 $w=1.5e-07 $l=2.14369e-07 $layer=POLY_cond $X=1.07 $Y=1.35
+ $X2=1.085 $Y2=1.557
r186 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.07 $Y=1.35 $X2=1.07
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__XNOR2_2%A_133_368# 1 2 7 9 10 12 13 15 16 18 19 24
+ 28 33 35 40
c99 40 0 2.33841e-19 $X=2.495 $Y=1.492
c100 33 0 1.43539e-19 $X=2.42 $Y=1.385
r101 37 38 1.9127 $w=3.78e-07 $l=1.5e-08 $layer=POLY_cond $X=2.045 $Y=1.492
+ $X2=2.06 $Y2=1.492
r102 34 40 9.56349 $w=3.78e-07 $l=7.5e-08 $layer=POLY_cond $X=2.42 $Y=1.492
+ $X2=2.495 $Y2=1.492
r103 34 38 45.9048 $w=3.78e-07 $l=3.6e-07 $layer=POLY_cond $X=2.42 $Y=1.492
+ $X2=2.06 $Y2=1.492
r104 33 35 17.2988 $w=5.38e-07 $l=5.05e-07 $layer=LI1_cond $X=2.42 $Y=1.28
+ $X2=1.915 $Y2=1.28
r105 33 34 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.42
+ $Y=1.385 $X2=2.42 $Y2=1.385
r106 30 31 6.78944 $w=4.43e-07 $l=8.5e-08 $layer=LI1_cond $X=1.227 $Y=1.095
+ $X2=1.227 $Y2=1.18
r107 28 30 7.63979 $w=4.43e-07 $l=2.95e-07 $layer=LI1_cond $X=1.227 $Y=0.8
+ $X2=1.227 $Y2=1.095
r108 26 30 6.43131 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=1.45 $Y=1.095
+ $X2=1.227 $Y2=1.095
r109 26 35 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=1.45 $Y=1.095
+ $X2=1.915 $Y2=1.095
r110 24 31 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=1.09 $Y=1.82
+ $X2=1.09 $Y2=1.18
r111 19 24 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.005 $Y=1.985
+ $X2=1.09 $Y2=1.82
r112 19 21 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=1.005 $Y=1.985
+ $X2=0.835 $Y2=1.985
r113 16 40 26.7778 $w=3.78e-07 $l=3.62083e-07 $layer=POLY_cond $X=2.705 $Y=1.22
+ $X2=2.495 $Y2=1.492
r114 16 18 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.705 $Y=1.22
+ $X2=2.705 $Y2=0.74
r115 13 40 24.4846 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=2.495 $Y=1.765
+ $X2=2.495 $Y2=1.492
r116 13 15 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.495 $Y=1.765
+ $X2=2.495 $Y2=2.4
r117 10 38 24.4846 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=2.06 $Y=1.22
+ $X2=2.06 $Y2=1.492
r118 10 12 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.06 $Y=1.22
+ $X2=2.06 $Y2=0.74
r119 7 37 24.4846 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=2.045 $Y=1.765
+ $X2=2.045 $Y2=1.492
r120 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.045 $Y=1.765
+ $X2=2.045 $Y2=2.4
r121 2 21 600 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_PDIFF $count=1 $X=0.665
+ $Y=1.84 $X2=0.835 $Y2=1.985
r122 1 28 182 $w=1.7e-07 $l=4.95076e-07 $layer=licon1_NDIFF $count=1 $X=1.145
+ $Y=0.37 $X2=1.285 $Y2=0.8
.ends

.subckt PM_SKY130_FD_SC_LS__XNOR2_2%VPWR 1 2 3 4 13 15 17 21 23 25 27 29 34 46
+ 53 57
r67 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r68 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r69 41 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r70 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r71 38 41 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.56 $Y2=3.33
r72 37 40 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=3.12 $Y=3.33
+ $X2=4.56 $Y2=3.33
r73 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r74 35 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.97 $Y=3.33
+ $X2=2.805 $Y2=3.33
r75 35 37 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=2.97 $Y=3.33 $X2=3.12
+ $Y2=3.33
r76 34 56 4.67153 $w=1.7e-07 $l=2.37e-07 $layer=LI1_cond $X=4.805 $Y=3.33
+ $X2=5.042 $Y2=3.33
r77 34 40 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=4.805 $Y=3.33
+ $X2=4.56 $Y2=3.33
r78 33 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r79 33 44 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.24 $Y2=3.33
r80 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r81 30 43 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.222 $Y2=3.33
r82 30 32 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=1.2 $Y2=3.33
r83 29 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r84 29 46 9.36465 $w=6.43e-07 $l=5.05e-07 $layer=LI1_cond $X=1.552 $Y=3.33
+ $X2=1.552 $Y2=2.825
r85 29 32 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=1.23 $Y=3.33 $X2=1.2
+ $Y2=3.33
r86 27 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r87 27 50 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=1.68 $Y2=3.33
r88 27 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r89 23 56 3.09464 $w=3.3e-07 $l=1.15521e-07 $layer=LI1_cond $X=4.97 $Y=3.245
+ $X2=5.042 $Y2=3.33
r90 23 25 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=4.97 $Y=3.245
+ $X2=4.97 $Y2=2.485
r91 19 53 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.805 $Y=3.245
+ $X2=2.805 $Y2=3.33
r92 19 21 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=2.805 $Y=3.245
+ $X2=2.805 $Y2=2.905
r93 18 29 8.78548 $w=1.7e-07 $l=3.23e-07 $layer=LI1_cond $X=1.875 $Y=3.33
+ $X2=1.552 $Y2=3.33
r94 17 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.64 $Y=3.33
+ $X2=2.805 $Y2=3.33
r95 17 18 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=2.64 $Y=3.33
+ $X2=1.875 $Y2=3.33
r96 13 43 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.222 $Y2=3.33
r97 13 15 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.28 $Y2=2.825
r98 4 25 300 $w=1.7e-07 $l=7.38258e-07 $layer=licon1_PDIFF $count=2 $X=4.77
+ $Y=1.84 $X2=4.97 $Y2=2.485
r99 3 21 600 $w=1.7e-07 $l=1.17665e-06 $layer=licon1_PDIFF $count=1 $X=2.57
+ $Y=1.84 $X2=2.805 $Y2=2.905
r100 2 46 300 $w=1.7e-07 $l=1.26126e-06 $layer=licon1_PDIFF $count=2 $X=1.16
+ $Y=1.84 $X2=1.79 $Y2=2.825
r101 1 15 600 $w=1.7e-07 $l=1.05501e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.825
.ends

.subckt PM_SKY130_FD_SC_LS__XNOR2_2%Y 1 2 3 11 12 13 14 15 17 19 20 23 24 26 31
+ 32 42
r101 35 46 2.51173 $w=3.88e-07 $l=8.5e-08 $layer=LI1_cond $X=2.24 $Y=2.57
+ $X2=2.24 $Y2=2.485
r102 32 39 1.47749 $w=3.88e-07 $l=5e-08 $layer=LI1_cond $X=2.24 $Y=2.775
+ $X2=2.24 $Y2=2.825
r103 32 35 6.05771 $w=3.88e-07 $l=2.05e-07 $layer=LI1_cond $X=2.24 $Y=2.775
+ $X2=2.24 $Y2=2.57
r104 31 46 2.36399 $w=3.88e-07 $l=8e-08 $layer=LI1_cond $X=2.24 $Y=2.405
+ $X2=2.24 $Y2=2.485
r105 31 42 7.68295 $w=3.88e-07 $l=2.6e-07 $layer=LI1_cond $X=2.24 $Y=2.405
+ $X2=2.24 $Y2=2.145
r106 26 29 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=3.97 $Y=2.485 $X2=3.97
+ $Y2=2.565
r107 23 24 10.0285 $w=2.43e-07 $l=1.9e-07 $layer=LI1_cond $X=2.38 $Y=0.377
+ $X2=2.19 $Y2=0.377
r108 21 46 5.6248 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=2.435 $Y=2.485
+ $X2=2.24 $Y2=2.485
r109 20 26 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.805 $Y=2.485
+ $X2=3.97 $Y2=2.485
r110 20 21 89.3797 $w=1.68e-07 $l=1.37e-06 $layer=LI1_cond $X=3.805 $Y=2.485
+ $X2=2.435 $Y2=2.485
r111 19 24 88.4011 $w=1.68e-07 $l=1.355e-06 $layer=LI1_cond $X=0.835 $Y=0.34
+ $X2=2.19 $Y2=0.34
r112 16 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.75 $Y=0.425
+ $X2=0.835 $Y2=0.34
r113 16 17 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=0.75 $Y=0.425
+ $X2=0.75 $Y2=0.84
r114 14 31 5.6248 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=2.045 $Y=2.405
+ $X2=2.24 $Y2=2.405
r115 14 15 116.781 $w=1.68e-07 $l=1.79e-06 $layer=LI1_cond $X=2.045 $Y=2.405
+ $X2=0.255 $Y2=2.405
r116 12 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.665 $Y=0.925
+ $X2=0.75 $Y2=0.84
r117 12 13 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=0.665 $Y=0.925
+ $X2=0.255 $Y2=0.925
r118 11 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.17 $Y=2.32
+ $X2=0.255 $Y2=2.405
r119 10 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.17 $Y=1.01
+ $X2=0.255 $Y2=0.925
r120 10 11 85.4652 $w=1.68e-07 $l=1.31e-06 $layer=LI1_cond $X=0.17 $Y=1.01
+ $X2=0.17 $Y2=2.32
r121 3 29 600 $w=1.7e-07 $l=7.96477e-07 $layer=licon1_PDIFF $count=1 $X=3.82
+ $Y=1.84 $X2=3.97 $Y2=2.565
r122 2 42 400 $w=1.7e-07 $l=3.72525e-07 $layer=licon1_PDIFF $count=1 $X=2.12
+ $Y=1.84 $X2=2.27 $Y2=2.145
r123 2 39 400 $w=1.7e-07 $l=1.05734e-06 $layer=licon1_PDIFF $count=1 $X=2.12
+ $Y=1.84 $X2=2.27 $Y2=2.825
r124 1 23 182 $w=1.7e-07 $l=2.66552e-07 $layer=licon1_NDIFF $count=1 $X=2.135
+ $Y=0.37 $X2=2.38 $Y2=0.415
.ends

.subckt PM_SKY130_FD_SC_LS__XNOR2_2%A_638_368# 1 2 7 11 14
r27 14 16 2.88111 $w=3.38e-07 $l=8.5e-08 $layer=LI1_cond $X=3.43 $Y=2.905
+ $X2=3.43 $Y2=2.99
r28 9 11 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=4.47 $Y=2.905
+ $X2=4.47 $Y2=2.485
r29 8 16 4.80115 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=3.6 $Y=2.99 $X2=3.43
+ $Y2=2.99
r30 7 9 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.305 $Y=2.99
+ $X2=4.47 $Y2=2.905
r31 7 8 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=4.305 $Y=2.99 $X2=3.6
+ $Y2=2.99
r32 2 11 300 $w=1.7e-07 $l=7.38258e-07 $layer=licon1_PDIFF $count=2 $X=4.27
+ $Y=1.84 $X2=4.47 $Y2=2.485
r33 1 14 600 $w=1.7e-07 $l=1.17891e-06 $layer=licon1_PDIFF $count=1 $X=3.19
+ $Y=1.84 $X2=3.43 $Y2=2.905
.ends

.subckt PM_SKY130_FD_SC_LS__XNOR2_2%VGND 1 2 3 10 12 16 20 23 24 25 34 40 41 47
r62 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r63 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r64 41 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.56
+ $Y2=0
r65 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r66 38 47 8.88104 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=4.655 $Y=0 $X2=4.482
+ $Y2=0
r67 38 40 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=4.655 $Y=0 $X2=5.04
+ $Y2=0
r68 37 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r69 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r70 34 47 8.88104 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=4.31 $Y=0 $X2=4.482
+ $Y2=0
r71 34 36 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=4.31 $Y=0 $X2=4.08
+ $Y2=0
r72 33 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r73 32 33 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r74 30 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r75 29 32 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=0.72 $Y=0 $X2=3.12
+ $Y2=0
r76 29 30 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r77 27 44 5.19892 $w=1.7e-07 $l=2.48e-07 $layer=LI1_cond $X=0.495 $Y=0 $X2=0.247
+ $Y2=0
r78 27 29 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.495 $Y=0 $X2=0.72
+ $Y2=0
r79 25 33 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r80 25 30 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.64 $Y=0 $X2=0.72
+ $Y2=0
r81 23 32 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=3.265 $Y=0 $X2=3.12
+ $Y2=0
r82 23 24 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=3.265 $Y=0 $X2=3.432
+ $Y2=0
r83 22 36 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r84 22 24 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=3.6 $Y=0 $X2=3.432
+ $Y2=0
r85 18 47 1.03204 $w=3.45e-07 $l=8.5e-08 $layer=LI1_cond $X=4.482 $Y=0.085
+ $X2=4.482 $Y2=0
r86 18 20 8.35104 $w=3.43e-07 $l=2.5e-07 $layer=LI1_cond $X=4.482 $Y=0.085
+ $X2=4.482 $Y2=0.335
r87 14 24 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=3.432 $Y=0.085
+ $X2=3.432 $Y2=0
r88 14 16 8.60032 $w=3.33e-07 $l=2.5e-07 $layer=LI1_cond $X=3.432 $Y=0.085
+ $X2=3.432 $Y2=0.335
r89 10 44 2.99777 $w=3.8e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.305 $Y=0.085
+ $X2=0.247 $Y2=0
r90 10 12 12.7375 $w=3.78e-07 $l=4.2e-07 $layer=LI1_cond $X=0.305 $Y=0.085
+ $X2=0.305 $Y2=0.505
r91 3 20 182 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_NDIFF $count=1 $X=4.255
+ $Y=0.37 $X2=4.48 $Y2=0.335
r92 2 16 182 $w=1.7e-07 $l=2.36854e-07 $layer=licon1_NDIFF $count=1 $X=3.21
+ $Y=0.37 $X2=3.43 $Y2=0.335
r93 1 12 182 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.36 $X2=0.33 $Y2=0.505
.ends

.subckt PM_SKY130_FD_SC_LS__XNOR2_2%A_340_107# 1 2 3 4 13 17 22 24 30 31 33
c67 1 0 1.43539e-19 $X=1.7 $Y=0.535
r68 33 35 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=5 $Y=0.675 $X2=5
+ $Y2=0.755
r69 29 31 8.48848 $w=3.48e-07 $l=1.65e-07 $layer=LI1_cond $X=3.945 $Y=0.665
+ $X2=4.11 $Y2=0.665
r70 29 30 8.48848 $w=3.48e-07 $l=1.65e-07 $layer=LI1_cond $X=3.945 $Y=0.665
+ $X2=3.78 $Y2=0.665
r71 24 26 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=2.92 $Y=0.515
+ $X2=2.92 $Y2=0.755
r72 20 22 8.85254 $w=2.43e-07 $l=1.65e-07 $layer=LI1_cond $X=1.845 $Y=0.717
+ $X2=2.01 $Y2=0.717
r73 17 35 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.835 $Y=0.755 $X2=5
+ $Y2=0.755
r74 17 31 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=4.835 $Y=0.755
+ $X2=4.11 $Y2=0.755
r75 16 26 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.085 $Y=0.755
+ $X2=2.92 $Y2=0.755
r76 16 30 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=3.085 $Y=0.755
+ $X2=3.78 $Y2=0.755
r77 13 26 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.755 $Y=0.755
+ $X2=2.92 $Y2=0.755
r78 13 22 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=2.755 $Y=0.755
+ $X2=2.01 $Y2=0.755
r79 4 33 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=4.86
+ $Y=0.37 $X2=5 $Y2=0.675
r80 3 29 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=3.805
+ $Y=0.37 $X2=3.945 $Y2=0.675
r81 2 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.78
+ $Y=0.37 $X2=2.92 $Y2=0.515
r82 1 20 182 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_NDIFF $count=1 $X=1.7
+ $Y=0.535 $X2=1.845 $Y2=0.715
.ends

