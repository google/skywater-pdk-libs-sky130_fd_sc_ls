* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__dlrbn_2 D GATE_N RESET_B VGND VNB VPB VPWR Q Q_N
X0 VPWR a_27_112# a_595_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_363_74# a_230_74# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X2 a_592_74# a_230_74# a_670_74# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X3 VPWR a_838_48# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X4 a_363_74# a_230_74# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X5 VGND GATE_N a_230_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X6 VGND a_1446_368# Q_N VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X7 VPWR GATE_N a_230_74# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X8 a_790_74# a_838_48# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 VGND a_838_48# a_1446_368# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X10 VPWR a_670_74# a_838_48# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X11 VGND a_838_48# Q VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X12 VPWR a_1446_368# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X13 a_670_74# a_363_74# a_790_74# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 a_1066_74# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X15 VGND a_27_112# a_592_74# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X16 Q a_838_48# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X17 Q a_838_48# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X18 a_595_392# a_363_74# a_670_74# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 Q_N a_1446_368# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X20 a_27_112# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X21 a_838_48# a_670_74# a_1066_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X22 a_670_74# a_230_74# a_783_508# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X23 VPWR a_838_48# a_1446_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X24 Q_N a_1446_368# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X25 a_783_508# a_838_48# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X26 a_27_112# D VGND VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X27 a_838_48# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
.ends
