* NGSPICE file created from sky130_fd_sc_ls__clkdlyinv3sd3_1.ext - technology: sky130A

.subckt sky130_fd_sc_ls__clkdlyinv3sd3_1 A VGND VNB VPB VPWR Y
M1000 a_288_74# a_28_74# VGND VNB nshort w=420000u l=500000u
+  ad=1.113e+11p pd=1.37e+06u as=2.73e+11p ps=2.98e+06u
M1001 a_288_74# a_28_74# VPWR VPB phighvt w=1e+06u l=500000u
+  ad=2.6e+11p pd=2.52e+06u as=7.148e+11p ps=5.78e+06u
M1002 VGND A a_28_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1003 VPWR A a_28_74# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1004 Y a_288_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1005 Y a_288_74# VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
.ends

