* File: sky130_fd_sc_ls__o311a_2.pxi.spice
* Created: Fri Aug 28 13:51:31 2020
* 
x_PM_SKY130_FD_SC_LS__O311A_2%C1 N_C1_M1000_g N_C1_c_72_n N_C1_M1006_g
+ N_C1_c_69_n N_C1_c_70_n C1 PM_SKY130_FD_SC_LS__O311A_2%C1
x_PM_SKY130_FD_SC_LS__O311A_2%B1 N_B1_M1012_g N_B1_c_97_n N_B1_M1002_g B1
+ N_B1_c_98_n PM_SKY130_FD_SC_LS__O311A_2%B1
x_PM_SKY130_FD_SC_LS__O311A_2%A3 N_A3_M1001_g N_A3_c_129_n N_A3_M1009_g A3
+ N_A3_c_130_n PM_SKY130_FD_SC_LS__O311A_2%A3
x_PM_SKY130_FD_SC_LS__O311A_2%A2 N_A2_c_158_n N_A2_M1005_g N_A2_M1013_g A2 A2 A2
+ A2 N_A2_c_160_n PM_SKY130_FD_SC_LS__O311A_2%A2
x_PM_SKY130_FD_SC_LS__O311A_2%A1 N_A1_c_190_n N_A1_M1011_g N_A1_M1007_g A1
+ N_A1_c_192_n PM_SKY130_FD_SC_LS__O311A_2%A1
x_PM_SKY130_FD_SC_LS__O311A_2%A_32_74# N_A_32_74#_M1000_s N_A_32_74#_M1006_s
+ N_A_32_74#_M1002_d N_A_32_74#_c_225_n N_A_32_74#_M1004_g N_A_32_74#_c_219_n
+ N_A_32_74#_M1003_g N_A_32_74#_c_226_n N_A_32_74#_M1010_g N_A_32_74#_c_220_n
+ N_A_32_74#_M1008_g N_A_32_74#_c_227_n N_A_32_74#_c_221_n N_A_32_74#_c_222_n
+ N_A_32_74#_c_236_n N_A_32_74#_c_258_n N_A_32_74#_c_228_n N_A_32_74#_c_229_n
+ N_A_32_74#_c_223_n N_A_32_74#_c_224_n PM_SKY130_FD_SC_LS__O311A_2%A_32_74#
x_PM_SKY130_FD_SC_LS__O311A_2%VPWR N_VPWR_M1006_d N_VPWR_M1011_d N_VPWR_M1010_s
+ N_VPWR_c_323_n N_VPWR_c_324_n N_VPWR_c_325_n N_VPWR_c_326_n N_VPWR_c_327_n
+ N_VPWR_c_328_n N_VPWR_c_329_n N_VPWR_c_330_n VPWR N_VPWR_c_331_n
+ N_VPWR_c_322_n PM_SKY130_FD_SC_LS__O311A_2%VPWR
x_PM_SKY130_FD_SC_LS__O311A_2%X N_X_M1003_d N_X_M1004_d N_X_c_379_n N_X_c_376_n
+ N_X_c_380_n N_X_c_381_n N_X_c_396_n N_X_c_397_n X X X N_X_c_378_n N_X_c_383_n
+ X PM_SKY130_FD_SC_LS__O311A_2%X
x_PM_SKY130_FD_SC_LS__O311A_2%A_219_74# N_A_219_74#_M1012_d N_A_219_74#_M1013_d
+ N_A_219_74#_c_426_n N_A_219_74#_c_423_n N_A_219_74#_c_424_n
+ PM_SKY130_FD_SC_LS__O311A_2%A_219_74#
x_PM_SKY130_FD_SC_LS__O311A_2%VGND N_VGND_M1001_d N_VGND_M1007_d N_VGND_M1008_s
+ N_VGND_c_451_n N_VGND_c_452_n N_VGND_c_453_n N_VGND_c_454_n N_VGND_c_455_n
+ N_VGND_c_456_n N_VGND_c_457_n VGND N_VGND_c_458_n N_VGND_c_459_n
+ PM_SKY130_FD_SC_LS__O311A_2%VGND
cc_1 VNB N_C1_c_69_n 0.0755182f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.385
cc_2 VNB N_C1_c_70_n 0.0223455f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.22
cc_3 VNB C1 0.0144311f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_B1_M1012_g 0.0252948f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=0.74
cc_5 VNB N_B1_c_97_n 0.0246662f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=2.34
cc_6 VNB N_B1_c_98_n 0.00392806f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_7 VNB N_A3_M1001_g 0.0286878f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=0.74
cc_8 VNB N_A3_c_129_n 0.0262515f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=2.34
cc_9 VNB N_A3_c_130_n 0.00166777f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_10 VNB N_A2_c_158_n 0.0266305f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.22
cc_11 VNB N_A2_M1013_g 0.027243f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=2.34
cc_12 VNB N_A2_c_160_n 0.0016809f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A1_c_190_n 0.0252926f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.22
cc_14 VNB N_A1_M1007_g 0.0257689f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=2.34
cc_15 VNB N_A1_c_192_n 0.00420079f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_16 VNB N_A_32_74#_c_219_n 0.0181781f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_17 VNB N_A_32_74#_c_220_n 0.0181832f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_18 VNB N_A_32_74#_c_221_n 0.00466883f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_32_74#_c_222_n 0.0440786f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_32_74#_c_223_n 0.00348446f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_32_74#_c_224_n 0.0541667f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VPWR_c_322_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_X_c_376_n 0.00208471f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB X 0.0311383f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_X_c_378_n 0.00995846f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_219_74#_c_423_n 0.00284354f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_27 VNB N_A_219_74#_c_424_n 0.00238751f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_451_n 0.00979921f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_29 VNB N_VGND_c_452_n 0.0125758f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_30 VNB N_VGND_c_453_n 0.0227978f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.295
cc_31 VNB N_VGND_c_454_n 0.0173724f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_455_n 0.0481805f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_33 VNB N_VGND_c_456_n 0.0182861f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_457_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_458_n 0.0201153f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_459_n 0.260862f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VPB N_C1_c_72_n 0.020583f $X=-0.19 $Y=1.66 $X2=0.615 $Y2=1.765
cc_38 VPB N_C1_c_69_n 0.00954682f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=1.385
cc_39 VPB N_B1_c_97_n 0.0275526f $X=-0.19 $Y=1.66 $X2=0.615 $Y2=2.34
cc_40 VPB N_B1_c_98_n 0.0034441f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_41 VPB N_A3_c_129_n 0.0283013f $X=-0.19 $Y=1.66 $X2=0.615 $Y2=2.34
cc_42 VPB N_A3_c_130_n 0.00278611f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_43 VPB N_A2_c_158_n 0.0263875f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.22
cc_44 VPB N_A2_c_160_n 0.00259972f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_45 VPB N_A1_c_190_n 0.027881f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.22
cc_46 VPB N_A1_c_192_n 0.00650827f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_47 VPB N_A_32_74#_c_225_n 0.0165084f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_48 VPB N_A_32_74#_c_226_n 0.0165278f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.295
cc_49 VPB N_A_32_74#_c_227_n 0.0319091f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_A_32_74#_c_228_n 0.00382185f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_51 VPB N_A_32_74#_c_229_n 0.0152996f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_A_32_74#_c_223_n 0.00120072f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_A_32_74#_c_224_n 0.014258f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_323_n 0.0168614f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_55 VPB N_VPWR_c_324_n 0.00663353f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.295
cc_56 VPB N_VPWR_c_325_n 0.0136263f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_326_n 0.047631f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_327_n 0.0244728f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_328_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_329_n 0.0472057f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_330_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_331_n 0.0213997f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_322_n 0.0980525f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_X_c_379_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0.615 $Y2=1.22
cc_65 VPB N_X_c_380_n 0.00234139f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_X_c_381_n 0.00284528f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB X 0.00313078f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_X_c_383_n 0.00953878f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 N_C1_c_69_n N_B1_M1012_g 0.0238802f $X=0.525 $Y=1.385 $X2=0 $Y2=0
cc_70 N_C1_c_70_n N_B1_M1012_g 0.0435734f $X=0.615 $Y=1.22 $X2=0 $Y2=0
cc_71 N_C1_c_72_n N_B1_c_97_n 0.0194911f $X=0.615 $Y=1.765 $X2=0 $Y2=0
cc_72 N_C1_c_69_n N_B1_c_97_n 0.00244604f $X=0.525 $Y=1.385 $X2=0 $Y2=0
cc_73 N_C1_c_69_n N_B1_c_98_n 6.43517e-19 $X=0.525 $Y=1.385 $X2=0 $Y2=0
cc_74 N_C1_c_72_n N_A_32_74#_c_227_n 0.0126017f $X=0.615 $Y=1.765 $X2=0 $Y2=0
cc_75 N_C1_c_69_n N_A_32_74#_c_221_n 0.00413135f $X=0.525 $Y=1.385 $X2=0 $Y2=0
cc_76 N_C1_c_70_n N_A_32_74#_c_221_n 0.0296397f $X=0.615 $Y=1.22 $X2=0 $Y2=0
cc_77 C1 N_A_32_74#_c_221_n 0.0200679f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_78 N_C1_c_72_n N_A_32_74#_c_236_n 3.73256e-19 $X=0.615 $Y=1.765 $X2=0 $Y2=0
cc_79 N_C1_c_72_n N_A_32_74#_c_229_n 0.0148691f $X=0.615 $Y=1.765 $X2=0 $Y2=0
cc_80 N_C1_c_69_n N_A_32_74#_c_229_n 0.00599406f $X=0.525 $Y=1.385 $X2=0 $Y2=0
cc_81 C1 N_A_32_74#_c_229_n 0.0125623f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_82 N_C1_c_72_n N_A_32_74#_c_223_n 0.00284738f $X=0.615 $Y=1.765 $X2=0 $Y2=0
cc_83 N_C1_c_69_n N_A_32_74#_c_223_n 0.0213041f $X=0.525 $Y=1.385 $X2=0 $Y2=0
cc_84 N_C1_c_70_n N_A_32_74#_c_223_n 7.45067e-19 $X=0.615 $Y=1.22 $X2=0 $Y2=0
cc_85 C1 N_A_32_74#_c_223_n 0.0265183f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_86 N_C1_c_72_n N_VPWR_c_323_n 0.00798178f $X=0.615 $Y=1.765 $X2=0 $Y2=0
cc_87 N_C1_c_72_n N_VPWR_c_327_n 0.00438942f $X=0.615 $Y=1.765 $X2=0 $Y2=0
cc_88 N_C1_c_72_n N_VPWR_c_322_n 0.00508379f $X=0.615 $Y=1.765 $X2=0 $Y2=0
cc_89 N_C1_c_70_n N_VGND_c_455_n 0.00291513f $X=0.615 $Y=1.22 $X2=0 $Y2=0
cc_90 N_C1_c_70_n N_VGND_c_459_n 0.00362985f $X=0.615 $Y=1.22 $X2=0 $Y2=0
cc_91 N_B1_M1012_g N_A3_M1001_g 0.028005f $X=1.02 $Y=0.74 $X2=0 $Y2=0
cc_92 N_B1_c_97_n N_A3_c_129_n 0.0413102f $X=1.185 $Y=1.765 $X2=0 $Y2=0
cc_93 N_B1_c_98_n N_A3_c_129_n 0.00214941f $X=1.11 $Y=1.515 $X2=0 $Y2=0
cc_94 N_B1_c_97_n N_A3_c_130_n 7.18891e-19 $X=1.185 $Y=1.765 $X2=0 $Y2=0
cc_95 N_B1_c_98_n N_A3_c_130_n 0.0347535f $X=1.11 $Y=1.515 $X2=0 $Y2=0
cc_96 N_B1_c_97_n N_A_32_74#_c_227_n 6.62055e-19 $X=1.185 $Y=1.765 $X2=0 $Y2=0
cc_97 N_B1_M1012_g N_A_32_74#_c_221_n 0.00911188f $X=1.02 $Y=0.74 $X2=0 $Y2=0
cc_98 N_B1_M1012_g N_A_32_74#_c_222_n 0.0154674f $X=1.02 $Y=0.74 $X2=0 $Y2=0
cc_99 N_B1_c_97_n N_A_32_74#_c_222_n 0.00125395f $X=1.185 $Y=1.765 $X2=0 $Y2=0
cc_100 N_B1_c_98_n N_A_32_74#_c_222_n 0.0279742f $X=1.11 $Y=1.515 $X2=0 $Y2=0
cc_101 N_B1_c_97_n N_A_32_74#_c_236_n 0.0166229f $X=1.185 $Y=1.765 $X2=0 $Y2=0
cc_102 N_B1_c_98_n N_A_32_74#_c_236_n 0.0243966f $X=1.11 $Y=1.515 $X2=0 $Y2=0
cc_103 N_B1_c_97_n N_A_32_74#_c_228_n 0.0111304f $X=1.185 $Y=1.765 $X2=0 $Y2=0
cc_104 N_B1_M1012_g N_A_32_74#_c_223_n 0.00530675f $X=1.02 $Y=0.74 $X2=0 $Y2=0
cc_105 N_B1_c_97_n N_A_32_74#_c_223_n 0.00390313f $X=1.185 $Y=1.765 $X2=0 $Y2=0
cc_106 N_B1_c_98_n N_A_32_74#_c_223_n 0.0330201f $X=1.11 $Y=1.515 $X2=0 $Y2=0
cc_107 N_B1_c_97_n N_VPWR_c_323_n 0.00146692f $X=1.185 $Y=1.765 $X2=0 $Y2=0
cc_108 N_B1_c_97_n N_VPWR_c_329_n 0.0049405f $X=1.185 $Y=1.765 $X2=0 $Y2=0
cc_109 N_B1_c_97_n N_VPWR_c_322_n 0.00508379f $X=1.185 $Y=1.765 $X2=0 $Y2=0
cc_110 N_B1_M1012_g N_A_219_74#_c_423_n 0.00577459f $X=1.02 $Y=0.74 $X2=0 $Y2=0
cc_111 N_B1_M1012_g N_VGND_c_455_n 0.00461464f $X=1.02 $Y=0.74 $X2=0 $Y2=0
cc_112 N_B1_M1012_g N_VGND_c_459_n 0.0091035f $X=1.02 $Y=0.74 $X2=0 $Y2=0
cc_113 N_A3_c_129_n N_A2_c_158_n 0.082886f $X=1.725 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_114 N_A3_c_130_n N_A2_c_158_n 0.00130194f $X=1.65 $Y=1.515 $X2=-0.19
+ $Y2=-0.245
cc_115 N_A3_M1001_g N_A2_M1013_g 0.0201424f $X=1.56 $Y=0.74 $X2=0 $Y2=0
cc_116 N_A3_c_129_n N_A2_c_160_n 0.00603367f $X=1.725 $Y=1.765 $X2=0 $Y2=0
cc_117 N_A3_c_130_n N_A2_c_160_n 0.0277335f $X=1.65 $Y=1.515 $X2=0 $Y2=0
cc_118 N_A3_M1001_g N_A_32_74#_c_222_n 0.0121365f $X=1.56 $Y=0.74 $X2=0 $Y2=0
cc_119 N_A3_c_129_n N_A_32_74#_c_222_n 0.00124693f $X=1.725 $Y=1.765 $X2=0 $Y2=0
cc_120 N_A3_c_130_n N_A_32_74#_c_222_n 0.0247243f $X=1.65 $Y=1.515 $X2=0 $Y2=0
cc_121 N_A3_c_129_n N_A_32_74#_c_258_n 0.00332234f $X=1.725 $Y=1.765 $X2=0 $Y2=0
cc_122 N_A3_c_130_n N_A_32_74#_c_258_n 0.0131798f $X=1.65 $Y=1.515 $X2=0 $Y2=0
cc_123 N_A3_c_129_n N_A_32_74#_c_228_n 0.0124764f $X=1.725 $Y=1.765 $X2=0 $Y2=0
cc_124 N_A3_c_129_n N_VPWR_c_323_n 0.00274927f $X=1.725 $Y=1.765 $X2=0 $Y2=0
cc_125 N_A3_c_129_n N_VPWR_c_329_n 0.00445602f $X=1.725 $Y=1.765 $X2=0 $Y2=0
cc_126 N_A3_c_129_n N_VPWR_c_322_n 0.00862959f $X=1.725 $Y=1.765 $X2=0 $Y2=0
cc_127 N_A3_M1001_g N_A_219_74#_c_426_n 0.0101937f $X=1.56 $Y=0.74 $X2=0 $Y2=0
cc_128 N_A3_M1001_g N_A_219_74#_c_423_n 0.00821463f $X=1.56 $Y=0.74 $X2=0 $Y2=0
cc_129 N_A3_M1001_g N_A_219_74#_c_424_n 8.12228e-19 $X=1.56 $Y=0.74 $X2=0 $Y2=0
cc_130 N_A3_M1001_g N_VGND_c_454_n 0.00472847f $X=1.56 $Y=0.74 $X2=0 $Y2=0
cc_131 N_A3_M1001_g N_VGND_c_455_n 0.00324657f $X=1.56 $Y=0.74 $X2=0 $Y2=0
cc_132 N_A3_M1001_g N_VGND_c_459_n 0.00412987f $X=1.56 $Y=0.74 $X2=0 $Y2=0
cc_133 N_A2_c_158_n N_A1_c_190_n 0.0559305f $X=2.145 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_134 N_A2_c_160_n N_A1_c_190_n 0.0123305f $X=2.19 $Y=1.515 $X2=-0.19
+ $Y2=-0.245
cc_135 N_A2_M1013_g N_A1_M1007_g 0.0340316f $X=2.28 $Y=0.74 $X2=0 $Y2=0
cc_136 N_A2_c_158_n N_A1_c_192_n 0.00231886f $X=2.145 $Y=1.765 $X2=0 $Y2=0
cc_137 N_A2_c_160_n N_A1_c_192_n 0.0349694f $X=2.19 $Y=1.515 $X2=0 $Y2=0
cc_138 N_A2_c_158_n N_A_32_74#_c_222_n 0.00124873f $X=2.145 $Y=1.765 $X2=0 $Y2=0
cc_139 N_A2_M1013_g N_A_32_74#_c_222_n 0.0115698f $X=2.28 $Y=0.74 $X2=0 $Y2=0
cc_140 N_A2_c_160_n N_A_32_74#_c_222_n 0.0256551f $X=2.19 $Y=1.515 $X2=0 $Y2=0
cc_141 N_A2_c_158_n N_A_32_74#_c_228_n 0.00120234f $X=2.145 $Y=1.765 $X2=0 $Y2=0
cc_142 N_A2_c_158_n N_VPWR_c_324_n 0.00176709f $X=2.145 $Y=1.765 $X2=0 $Y2=0
cc_143 N_A2_c_160_n N_VPWR_c_324_n 0.038528f $X=2.19 $Y=1.515 $X2=0 $Y2=0
cc_144 N_A2_c_158_n N_VPWR_c_329_n 0.00303293f $X=2.145 $Y=1.765 $X2=0 $Y2=0
cc_145 N_A2_c_160_n N_VPWR_c_329_n 0.00865352f $X=2.19 $Y=1.515 $X2=0 $Y2=0
cc_146 N_A2_c_158_n N_VPWR_c_322_n 0.00372712f $X=2.145 $Y=1.765 $X2=0 $Y2=0
cc_147 N_A2_c_160_n N_VPWR_c_322_n 0.0106888f $X=2.19 $Y=1.515 $X2=0 $Y2=0
cc_148 N_A2_c_160_n A_444_368# 0.0143019f $X=2.19 $Y=1.515 $X2=-0.19 $Y2=-0.245
cc_149 N_A2_M1013_g N_A_219_74#_c_426_n 0.0101837f $X=2.28 $Y=0.74 $X2=0 $Y2=0
cc_150 N_A2_M1013_g N_A_219_74#_c_423_n 8.12228e-19 $X=2.28 $Y=0.74 $X2=0 $Y2=0
cc_151 N_A2_M1013_g N_A_219_74#_c_424_n 0.00810322f $X=2.28 $Y=0.74 $X2=0 $Y2=0
cc_152 N_A2_M1013_g N_VGND_c_454_n 0.00472847f $X=2.28 $Y=0.74 $X2=0 $Y2=0
cc_153 N_A2_M1013_g N_VGND_c_456_n 0.00324657f $X=2.28 $Y=0.74 $X2=0 $Y2=0
cc_154 N_A2_M1013_g N_VGND_c_459_n 0.00412056f $X=2.28 $Y=0.74 $X2=0 $Y2=0
cc_155 N_A1_c_190_n N_A_32_74#_c_225_n 0.0169521f $X=2.685 $Y=1.765 $X2=0 $Y2=0
cc_156 N_A1_M1007_g N_A_32_74#_c_219_n 0.0202161f $X=2.71 $Y=0.74 $X2=0 $Y2=0
cc_157 N_A1_c_190_n N_A_32_74#_c_222_n 0.00253309f $X=2.685 $Y=1.765 $X2=0 $Y2=0
cc_158 N_A1_M1007_g N_A_32_74#_c_222_n 0.0186271f $X=2.71 $Y=0.74 $X2=0 $Y2=0
cc_159 N_A1_c_192_n N_A_32_74#_c_222_n 0.0468355f $X=2.76 $Y=1.515 $X2=0 $Y2=0
cc_160 N_A1_c_190_n N_A_32_74#_c_224_n 0.0187888f $X=2.685 $Y=1.765 $X2=0 $Y2=0
cc_161 N_A1_M1007_g N_A_32_74#_c_224_n 0.00338438f $X=2.71 $Y=0.74 $X2=0 $Y2=0
cc_162 N_A1_c_192_n N_A_32_74#_c_224_n 0.00239804f $X=2.76 $Y=1.515 $X2=0 $Y2=0
cc_163 N_A1_c_190_n N_VPWR_c_324_n 0.020634f $X=2.685 $Y=1.765 $X2=0 $Y2=0
cc_164 N_A1_c_192_n N_VPWR_c_324_n 0.013098f $X=2.76 $Y=1.515 $X2=0 $Y2=0
cc_165 N_A1_c_190_n N_VPWR_c_329_n 0.00413917f $X=2.685 $Y=1.765 $X2=0 $Y2=0
cc_166 N_A1_c_190_n N_VPWR_c_322_n 0.00818558f $X=2.685 $Y=1.765 $X2=0 $Y2=0
cc_167 N_A1_c_190_n N_X_c_379_n 4.83351e-19 $X=2.685 $Y=1.765 $X2=0 $Y2=0
cc_168 N_A1_c_190_n N_X_c_381_n 5.37035e-19 $X=2.685 $Y=1.765 $X2=0 $Y2=0
cc_169 N_A1_c_192_n N_X_c_381_n 0.00264176f $X=2.76 $Y=1.515 $X2=0 $Y2=0
cc_170 N_A1_M1007_g N_A_219_74#_c_424_n 0.00681223f $X=2.71 $Y=0.74 $X2=0 $Y2=0
cc_171 N_A1_M1007_g N_VGND_c_451_n 0.00640249f $X=2.71 $Y=0.74 $X2=0 $Y2=0
cc_172 N_A1_M1007_g N_VGND_c_456_n 0.00434272f $X=2.71 $Y=0.74 $X2=0 $Y2=0
cc_173 N_A1_M1007_g N_VGND_c_459_n 0.00821587f $X=2.71 $Y=0.74 $X2=0 $Y2=0
cc_174 N_A_32_74#_c_236_n N_VPWR_M1006_d 0.0113525f $X=1.335 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_175 N_A_32_74#_c_229_n N_VPWR_M1006_d 0.00334484f $X=0.39 $Y=1.985 $X2=-0.19
+ $Y2=-0.245
cc_176 N_A_32_74#_c_227_n N_VPWR_c_323_n 0.044743f $X=0.39 $Y=2.695 $X2=0 $Y2=0
cc_177 N_A_32_74#_c_236_n N_VPWR_c_323_n 0.0225363f $X=1.335 $Y=2.035 $X2=0
+ $Y2=0
cc_178 N_A_32_74#_c_228_n N_VPWR_c_323_n 0.0270342f $X=1.5 $Y=2.815 $X2=0 $Y2=0
cc_179 N_A_32_74#_c_225_n N_VPWR_c_324_n 0.0126641f $X=3.27 $Y=1.765 $X2=0 $Y2=0
cc_180 N_A_32_74#_c_226_n N_VPWR_c_326_n 0.0227729f $X=3.72 $Y=1.765 $X2=0 $Y2=0
cc_181 N_A_32_74#_c_227_n N_VPWR_c_327_n 0.0111687f $X=0.39 $Y=2.695 $X2=0 $Y2=0
cc_182 N_A_32_74#_c_228_n N_VPWR_c_329_n 0.0145938f $X=1.5 $Y=2.815 $X2=0 $Y2=0
cc_183 N_A_32_74#_c_225_n N_VPWR_c_331_n 0.00445602f $X=3.27 $Y=1.765 $X2=0
+ $Y2=0
cc_184 N_A_32_74#_c_226_n N_VPWR_c_331_n 0.00445602f $X=3.72 $Y=1.765 $X2=0
+ $Y2=0
cc_185 N_A_32_74#_c_225_n N_VPWR_c_322_n 0.00859513f $X=3.27 $Y=1.765 $X2=0
+ $Y2=0
cc_186 N_A_32_74#_c_226_n N_VPWR_c_322_n 0.00860687f $X=3.72 $Y=1.765 $X2=0
+ $Y2=0
cc_187 N_A_32_74#_c_227_n N_VPWR_c_322_n 0.0128476f $X=0.39 $Y=2.695 $X2=0 $Y2=0
cc_188 N_A_32_74#_c_228_n N_VPWR_c_322_n 0.0120466f $X=1.5 $Y=2.815 $X2=0 $Y2=0
cc_189 N_A_32_74#_c_225_n N_X_c_379_n 0.0142282f $X=3.27 $Y=1.765 $X2=0 $Y2=0
cc_190 N_A_32_74#_c_226_n N_X_c_379_n 0.0173715f $X=3.72 $Y=1.765 $X2=0 $Y2=0
cc_191 N_A_32_74#_c_220_n N_X_c_376_n 0.0118569f $X=3.735 $Y=1.22 $X2=0 $Y2=0
cc_192 N_A_32_74#_c_226_n N_X_c_380_n 0.0101222f $X=3.72 $Y=1.765 $X2=0 $Y2=0
cc_193 N_A_32_74#_c_224_n N_X_c_380_n 0.00604231f $X=3.72 $Y=1.492 $X2=0 $Y2=0
cc_194 N_A_32_74#_c_225_n N_X_c_381_n 0.00351555f $X=3.27 $Y=1.765 $X2=0 $Y2=0
cc_195 N_A_32_74#_c_226_n N_X_c_381_n 0.00109449f $X=3.72 $Y=1.765 $X2=0 $Y2=0
cc_196 N_A_32_74#_c_222_n N_X_c_381_n 0.0151207f $X=3.095 $Y=1.095 $X2=0 $Y2=0
cc_197 N_A_32_74#_c_224_n N_X_c_381_n 0.00534575f $X=3.72 $Y=1.492 $X2=0 $Y2=0
cc_198 N_A_32_74#_c_220_n N_X_c_396_n 0.0142632f $X=3.735 $Y=1.22 $X2=0 $Y2=0
cc_199 N_A_32_74#_c_220_n N_X_c_397_n 0.00119573f $X=3.735 $Y=1.22 $X2=0 $Y2=0
cc_200 N_A_32_74#_c_222_n N_X_c_397_n 0.00614869f $X=3.095 $Y=1.095 $X2=0 $Y2=0
cc_201 N_A_32_74#_c_224_n N_X_c_397_n 0.00224023f $X=3.72 $Y=1.492 $X2=0 $Y2=0
cc_202 N_A_32_74#_c_220_n X 0.0220968f $X=3.735 $Y=1.22 $X2=0 $Y2=0
cc_203 N_A_32_74#_c_222_n X 0.0123458f $X=3.095 $Y=1.095 $X2=0 $Y2=0
cc_204 N_A_32_74#_c_221_n A_135_74# 0.00814767f $X=0.69 $Y=1.18 $X2=-0.19
+ $Y2=-0.245
cc_205 N_A_32_74#_c_222_n A_135_74# 0.00427342f $X=3.095 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_206 N_A_32_74#_c_222_n N_A_219_74#_M1012_d 0.00389656f $X=3.095 $Y=1.095
+ $X2=-0.19 $Y2=-0.245
cc_207 N_A_32_74#_c_222_n N_A_219_74#_M1013_d 0.00176461f $X=3.095 $Y=1.095
+ $X2=0 $Y2=0
cc_208 N_A_32_74#_c_222_n N_A_219_74#_c_426_n 0.0500659f $X=3.095 $Y=1.095 $X2=0
+ $Y2=0
cc_209 N_A_32_74#_c_221_n N_A_219_74#_c_423_n 0.0216996f $X=0.69 $Y=1.18 $X2=0
+ $Y2=0
cc_210 N_A_32_74#_c_222_n N_A_219_74#_c_423_n 0.0213487f $X=3.095 $Y=1.095 $X2=0
+ $Y2=0
cc_211 N_A_32_74#_c_222_n N_A_219_74#_c_424_n 0.0167101f $X=3.095 $Y=1.095 $X2=0
+ $Y2=0
cc_212 N_A_32_74#_c_222_n N_VGND_M1001_d 0.00600992f $X=3.095 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_213 N_A_32_74#_c_222_n N_VGND_M1007_d 0.00426848f $X=3.095 $Y=1.095 $X2=0
+ $Y2=0
cc_214 N_A_32_74#_c_219_n N_VGND_c_451_n 0.00845049f $X=3.305 $Y=1.22 $X2=0
+ $Y2=0
cc_215 N_A_32_74#_c_222_n N_VGND_c_451_n 0.0262206f $X=3.095 $Y=1.095 $X2=0
+ $Y2=0
cc_216 N_A_32_74#_c_220_n N_VGND_c_453_n 0.00957981f $X=3.735 $Y=1.22 $X2=0
+ $Y2=0
cc_217 N_A_32_74#_c_221_n N_VGND_c_455_n 0.0249477f $X=0.69 $Y=1.18 $X2=0 $Y2=0
cc_218 N_A_32_74#_c_219_n N_VGND_c_458_n 0.00461464f $X=3.305 $Y=1.22 $X2=0
+ $Y2=0
cc_219 N_A_32_74#_c_220_n N_VGND_c_458_n 0.00434272f $X=3.735 $Y=1.22 $X2=0
+ $Y2=0
cc_220 N_A_32_74#_c_219_n N_VGND_c_459_n 0.00910098f $X=3.305 $Y=1.22 $X2=0
+ $Y2=0
cc_221 N_A_32_74#_c_220_n N_VGND_c_459_n 0.00442526f $X=3.735 $Y=1.22 $X2=0
+ $Y2=0
cc_222 N_A_32_74#_c_221_n N_VGND_c_459_n 0.0203135f $X=0.69 $Y=1.18 $X2=0 $Y2=0
cc_223 N_VPWR_c_324_n N_X_c_379_n 0.0586183f $X=2.91 $Y=2.115 $X2=0 $Y2=0
cc_224 N_VPWR_c_326_n N_X_c_379_n 0.0353111f $X=3.995 $Y=2.145 $X2=0 $Y2=0
cc_225 N_VPWR_c_331_n N_X_c_379_n 0.014552f $X=3.83 $Y=3.33 $X2=0 $Y2=0
cc_226 N_VPWR_c_322_n N_X_c_379_n 0.0119791f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_227 N_VPWR_M1010_s N_X_c_380_n 0.00119058f $X=3.795 $Y=1.84 $X2=0 $Y2=0
cc_228 N_VPWR_c_326_n N_X_c_380_n 0.00915704f $X=3.995 $Y=2.145 $X2=0 $Y2=0
cc_229 N_VPWR_M1010_s N_X_c_383_n 0.00235172f $X=3.795 $Y=1.84 $X2=0 $Y2=0
cc_230 N_VPWR_c_326_n N_X_c_383_n 0.0175586f $X=3.995 $Y=2.145 $X2=0 $Y2=0
cc_231 N_X_c_396_n N_VGND_M1008_s 0.00306514f $X=3.965 $Y=0.93 $X2=0 $Y2=0
cc_232 X N_VGND_M1008_s 0.0013398f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_233 N_X_c_378_n N_VGND_M1008_s 0.00521203f $X=4.08 $Y=1.05 $X2=0 $Y2=0
cc_234 N_X_c_376_n N_VGND_c_451_n 0.0135169f $X=3.52 $Y=0.515 $X2=0 $Y2=0
cc_235 N_X_c_376_n N_VGND_c_453_n 0.00978743f $X=3.52 $Y=0.515 $X2=0 $Y2=0
cc_236 N_X_c_396_n N_VGND_c_453_n 0.00664376f $X=3.965 $Y=0.93 $X2=0 $Y2=0
cc_237 N_X_c_378_n N_VGND_c_453_n 0.0169147f $X=4.08 $Y=1.05 $X2=0 $Y2=0
cc_238 N_X_c_376_n N_VGND_c_458_n 0.0110175f $X=3.52 $Y=0.515 $X2=0 $Y2=0
cc_239 N_X_c_376_n N_VGND_c_459_n 0.0090528f $X=3.52 $Y=0.515 $X2=0 $Y2=0
cc_240 N_X_c_396_n N_VGND_c_459_n 0.00573789f $X=3.965 $Y=0.93 $X2=0 $Y2=0
cc_241 N_X_c_378_n N_VGND_c_459_n 9.73527e-19 $X=4.08 $Y=1.05 $X2=0 $Y2=0
cc_242 N_A_219_74#_c_426_n N_VGND_M1001_d 0.0112181f $X=2.33 $Y=0.755 $X2=-0.19
+ $Y2=-0.245
cc_243 N_A_219_74#_c_424_n N_VGND_c_451_n 0.0191765f $X=2.495 $Y=0.595 $X2=0
+ $Y2=0
cc_244 N_A_219_74#_c_426_n N_VGND_c_454_n 0.0351355f $X=2.33 $Y=0.755 $X2=0
+ $Y2=0
cc_245 N_A_219_74#_c_423_n N_VGND_c_454_n 0.00617451f $X=1.345 $Y=0.595 $X2=0
+ $Y2=0
cc_246 N_A_219_74#_c_424_n N_VGND_c_454_n 0.00617451f $X=2.495 $Y=0.595 $X2=0
+ $Y2=0
cc_247 N_A_219_74#_c_426_n N_VGND_c_455_n 0.00237563f $X=2.33 $Y=0.755 $X2=0
+ $Y2=0
cc_248 N_A_219_74#_c_423_n N_VGND_c_455_n 0.0142249f $X=1.345 $Y=0.595 $X2=0
+ $Y2=0
cc_249 N_A_219_74#_c_426_n N_VGND_c_456_n 0.00237563f $X=2.33 $Y=0.755 $X2=0
+ $Y2=0
cc_250 N_A_219_74#_c_424_n N_VGND_c_456_n 0.0141563f $X=2.495 $Y=0.595 $X2=0
+ $Y2=0
cc_251 N_A_219_74#_c_426_n N_VGND_c_459_n 0.0107664f $X=2.33 $Y=0.755 $X2=0
+ $Y2=0
cc_252 N_A_219_74#_c_423_n N_VGND_c_459_n 0.011867f $X=1.345 $Y=0.595 $X2=0
+ $Y2=0
cc_253 N_A_219_74#_c_424_n N_VGND_c_459_n 0.0117515f $X=2.495 $Y=0.595 $X2=0
+ $Y2=0
