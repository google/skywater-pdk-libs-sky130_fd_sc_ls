* File: sky130_fd_sc_ls__fa_1.spice
* Created: Wed Sep  2 11:07:31 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__fa_1.pex.spice"
.subckt sky130_fd_sc_ls__fa_1  VNB VPB A CIN B SUM VPWR COUT VGND
* 
* VGND	VGND
* COUT	COUT
* VPWR	VPWR
* SUM	SUM
* B	B
* CIN	CIN
* A	A
* VPB	VPB
* VNB	VNB
MM1024 N_VGND_M1024_d N_A_69_260#_M1024_g N_SUM_M1024_s VNB NSHORT L=0.15 W=0.74
+ AD=0.205457 AS=0.2109 PD=1.49609 PS=2.05 NRD=36.096 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75006 A=0.111 P=1.78 MULT=1
MM1008 A_237_75# N_A_M1008_g N_VGND_M1024_d VNB NSHORT L=0.15 W=0.64 AD=0.0768
+ AS=0.177693 PD=0.88 PS=1.29391 NRD=12.18 NRS=18.744 M=1 R=4.26667 SA=75000.8
+ SB=75006.3 A=0.096 P=1.58 MULT=1
MM1025 A_315_75# N_B_M1025_g A_237_75# VNB NSHORT L=0.15 W=0.64 AD=0.0768
+ AS=0.0768 PD=0.88 PS=0.88 NRD=12.18 NRS=12.18 M=1 R=4.26667 SA=75001.2
+ SB=75005.9 A=0.096 P=1.58 MULT=1
MM1026 N_A_69_260#_M1026_d N_CIN_M1026_g A_315_75# VNB NSHORT L=0.15 W=0.64
+ AD=0.1248 AS=0.0768 PD=1.03 PS=0.88 NRD=0 NRS=12.18 M=1 R=4.26667 SA=75001.6
+ SB=75005.5 A=0.096 P=1.58 MULT=1
MM1004 N_A_501_75#_M1004_d N_A_465_249#_M1004_g N_A_69_260#_M1026_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.1152 AS=0.1248 PD=1 PS=1.03 NRD=7.488 NRS=20.616 M=1
+ R=4.26667 SA=75002.1 SB=75005 A=0.096 P=1.58 MULT=1
MM1012 N_VGND_M1012_d N_B_M1012_g N_A_501_75#_M1004_d VNB NSHORT L=0.15 W=0.64
+ AD=0.169075 AS=0.1152 PD=1.275 PS=1 NRD=39.216 NRS=0 M=1 R=4.26667 SA=75002.7
+ SB=75004.5 A=0.096 P=1.58 MULT=1
MM1015 N_A_501_75#_M1015_d N_A_M1015_g N_VGND_M1012_d VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.169075 PD=0.92 PS=1.275 NRD=0 NRS=39.216 M=1 R=4.26667
+ SA=75003.2 SB=75003.9 A=0.096 P=1.58 MULT=1
MM1002 N_VGND_M1002_d N_CIN_M1002_g N_A_501_75#_M1015_d VNB NSHORT L=0.15 W=0.64
+ AD=0.1584 AS=0.0896 PD=1.135 PS=0.92 NRD=26.244 NRS=0 M=1 R=4.26667 SA=75003.7
+ SB=75003.4 A=0.096 P=1.58 MULT=1
MM1027 A_936_75# N_A_M1027_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.64 AD=0.0768
+ AS=0.1584 PD=0.88 PS=1.135 NRD=12.18 NRS=14.052 M=1 R=4.26667 SA=75004.3
+ SB=75002.8 A=0.096 P=1.58 MULT=1
MM1016 N_A_465_249#_M1016_d N_B_M1016_g A_936_75# VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.0768 PD=0.92 PS=0.88 NRD=0 NRS=12.18 M=1 R=4.26667 SA=75004.7
+ SB=75002.4 A=0.096 P=1.58 MULT=1
MM1020 N_A_1100_75#_M1020_d N_CIN_M1020_g N_A_465_249#_M1016_d VNB NSHORT L=0.15
+ W=0.64 AD=0.3596 AS=0.0896 PD=1.73 PS=0.92 NRD=95.028 NRS=0 M=1 R=4.26667
+ SA=75005.1 SB=75002 A=0.096 P=1.58 MULT=1
MM1018 N_VGND_M1018_d N_A_M1018_g N_A_1100_75#_M1020_d VNB NSHORT L=0.15 W=0.64
+ AD=0.212275 AS=0.3596 PD=1.41 PS=1.73 NRD=51.876 NRS=2.808 M=1 R=4.26667
+ SA=75006.2 SB=75000.9 A=0.096 P=1.58 MULT=1
MM1013 N_A_1100_75#_M1013_d N_B_M1013_g N_VGND_M1018_d VNB NSHORT L=0.15 W=0.64
+ AD=0.1696 AS=0.212275 PD=1.81 PS=1.41 NRD=0 NRS=51.876 M=1 R=4.26667
+ SA=75006.9 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1017 N_COUT_M1017_d N_A_465_249#_M1017_g N_VGND_M1017_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1998 AS=0.1961 PD=2.02 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1021 N_VPWR_M1021_d N_A_69_260#_M1021_g N_SUM_M1021_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.210264 AS=0.3192 PD=1.56906 PS=2.81 NRD=1.7533 NRS=1.7533 M=1
+ R=7.46667 SA=75000.2 SB=75004.9 A=0.168 P=2.54 MULT=1
MM1011 A_217_368# N_A_M1011_g N_VPWR_M1021_d VPB PHIGHVT L=0.15 W=1 AD=0.186687
+ AS=0.187736 PD=1.46 PS=1.40094 NRD=25.9252 NRS=15.0902 M=1 R=6.66667
+ SA=75000.7 SB=75004.9 A=0.15 P=2.3 MULT=1
MM1005 A_318_389# N_B_M1005_g A_217_368# VPB PHIGHVT L=0.15 W=1 AD=0.195875
+ AS=0.186687 PD=1.565 PS=1.46 NRD=27.7376 NRS=25.9252 M=1 R=6.66667 SA=75001.1
+ SB=75004.5 A=0.15 P=2.3 MULT=1
MM1000 N_A_69_260#_M1000_d N_CIN_M1000_g A_318_389# VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.195875 PD=1.3 PS=1.565 NRD=1.9503 NRS=27.7376 M=1 R=6.66667
+ SA=75001.4 SB=75005.1 A=0.15 P=2.3 MULT=1
MM1006 N_A_509_347#_M1006_d N_A_465_249#_M1006_g N_A_69_260#_M1000_d VPB PHIGHVT
+ L=0.15 W=1 AD=0.1675 AS=0.15 PD=1.335 PS=1.3 NRD=1.9503 NRS=1.9503 M=1
+ R=6.66667 SA=75001.9 SB=75004.6 A=0.15 P=2.3 MULT=1
MM1019 N_VPWR_M1019_d N_B_M1019_g N_A_509_347#_M1006_d VPB PHIGHVT L=0.15 W=1
+ AD=0.243637 AS=0.1675 PD=1.64 PS=1.335 NRD=37.1542 NRS=2.2852 M=1 R=6.66667
+ SA=75002.3 SB=75004.1 A=0.15 P=2.3 MULT=1
MM1003 N_A_509_347#_M1003_d N_A_M1003_g N_VPWR_M1019_d VPB PHIGHVT L=0.15 W=1
+ AD=0.1775 AS=0.243637 PD=1.355 PS=1.64 NRD=0 NRS=37.1542 M=1 R=6.66667
+ SA=75002.9 SB=75003.5 A=0.15 P=2.3 MULT=1
MM1007 N_VPWR_M1007_d N_CIN_M1007_g N_A_509_347#_M1003_d VPB PHIGHVT L=0.15 W=1
+ AD=0.155 AS=0.1775 PD=1.31 PS=1.355 NRD=1.9503 NRS=12.7853 M=1 R=6.66667
+ SA=75003.4 SB=75003 A=0.15 P=2.3 MULT=1
MM1009 A_916_347# N_A_M1009_g N_VPWR_M1007_d VPB PHIGHVT L=0.15 W=1 AD=0.1775
+ AS=0.155 PD=1.355 PS=1.31 NRD=24.1128 NRS=3.9203 M=1 R=6.66667 SA=75003.9
+ SB=75002.6 A=0.15 P=2.3 MULT=1
MM1010 N_A_465_249#_M1010_d N_B_M1010_g A_916_347# VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.1775 PD=1.3 PS=1.355 NRD=1.9503 NRS=24.1128 M=1 R=6.66667
+ SA=75004.4 SB=75002.1 A=0.15 P=2.3 MULT=1
MM1014 N_A_1107_347#_M1014_d N_CIN_M1014_g N_A_465_249#_M1010_d VPB PHIGHVT
+ L=0.15 W=1 AD=0.2225 AS=0.15 PD=1.445 PS=1.3 NRD=30.535 NRS=1.9503 M=1
+ R=6.66667 SA=75004.9 SB=75001.6 A=0.15 P=2.3 MULT=1
MM1022 N_VPWR_M1022_d N_A_M1022_g N_A_1107_347#_M1014_d VPB PHIGHVT L=0.15 W=1
+ AD=0.349062 AS=0.2225 PD=1.76 PS=1.445 NRD=2.9353 NRS=1.9503 M=1 R=6.66667
+ SA=75005.4 SB=75001 A=0.15 P=2.3 MULT=1
MM1001 N_A_1107_347#_M1001_d N_B_M1001_g N_VPWR_M1022_d VPB PHIGHVT L=0.15 W=1
+ AD=0.335 AS=0.349062 PD=2.67 PS=1.76 NRD=9.8303 NRS=2.9353 M=1 R=6.66667
+ SA=75005.9 SB=75000.3 A=0.15 P=2.3 MULT=1
MM1023 N_COUT_M1023_d N_A_465_249#_M1023_g N_VPWR_M1023_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.3192 AS=0.3304 PD=2.81 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.2 A=0.168 P=2.54 MULT=1
DX28_noxref VNB VPB NWDIODE A=17.4051 P=21.97
c_77 VNB 0 1.97438e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_ls__fa_1.pxi.spice"
*
.ends
*
*
