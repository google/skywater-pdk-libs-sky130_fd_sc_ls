* NGSPICE file created from sky130_fd_sc_ls__o41ai_1.ext - technology: sky130A

.subckt sky130_fd_sc_ls__o41ai_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
M1000 a_157_74# A1 VGND VNB nshort w=740000u l=150000u
+  ad=7.104e+11p pd=6.36e+06u as=6.327e+11p ps=4.67e+06u
M1001 Y B1 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.92e+11p pd=2.94e+06u as=9.072e+11p ps=6.1e+06u
M1002 a_157_74# A3 VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_260_368# A4 Y VPB phighvt w=1.12e+06u l=150000u
+  ad=3.808e+11p pd=2.92e+06u as=0p ps=0u
M1004 VPWR A1 a_472_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=4.704e+11p ps=3.08e+06u
M1005 a_472_368# A2 a_358_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=4.704e+11p ps=3.08e+06u
M1006 VGND A2 a_157_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND A4 a_157_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_157_74# B1 Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1009 a_358_368# A3 a_260_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

