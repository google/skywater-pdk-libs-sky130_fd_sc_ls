* File: sky130_fd_sc_ls__dlrtn_4.spice
* Created: Fri Aug 28 13:19:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__dlrtn_4.pex.spice"
.subckt sky130_fd_sc_ls__dlrtn_4  VNB VPB D GATE_N RESET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* RESET_B	RESET_B
* GATE_N	GATE_N
* D	D
* VPB	VPB
* VNB	VNB
MM1025 N_VGND_M1025_d N_D_M1025_g N_A_27_136#_M1025_s VNB NSHORT L=0.15 W=0.55
+ AD=0.171076 AS=0.15675 PD=1.27054 PS=1.67 NRD=55.86 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75000.9 A=0.0825 P=1.4 MULT=1
MM1002 N_A_232_98#_M1002_d N_GATE_N_M1002_g N_VGND_M1025_d VNB NSHORT L=0.15
+ W=0.74 AD=0.2886 AS=0.230174 PD=2.26 PS=1.70946 NRD=8.1 NRS=41.52 M=1
+ R=4.93333 SA=75000.7 SB=75000.3 A=0.111 P=1.78 MULT=1
MM1021 N_VGND_M1021_d N_A_232_98#_M1021_g N_A_348_392#_M1021_s VNB NSHORT L=0.15
+ W=0.74 AD=0.421076 AS=0.2109 PD=2.11812 PS=2.05 NRD=83.352 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001.6 A=0.111 P=1.78 MULT=1
MM1018 A_666_74# N_A_27_136#_M1018_g N_VGND_M1021_d VNB NSHORT L=0.15 W=0.64
+ AD=0.0768 AS=0.364174 PD=0.88 PS=1.83188 NRD=12.18 NRS=15.936 M=1 R=4.26667
+ SA=75001.2 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1017 N_A_639_392#_M1017_d N_A_232_98#_M1017_g A_666_74# VNB NSHORT L=0.15
+ W=0.64 AD=0.115623 AS=0.0768 PD=1.16528 PS=0.88 NRD=8.436 NRS=12.18 M=1
+ R=4.26667 SA=75001.6 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1007 A_839_74# N_A_348_392#_M1007_g N_A_639_392#_M1017_d VNB NSHORT L=0.15
+ W=0.42 AD=0.05775 AS=0.0758774 PD=0.695 PS=0.764717 NRD=23.568 NRS=0 M=1 R=2.8
+ SA=75002 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1016 N_VGND_M1016_d N_A_888_406#_M1016_g A_839_74# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.05775 PD=1.41 PS=0.695 NRD=0 NRS=23.568 M=1 R=2.8 SA=75002.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1010 N_A_1035_74#_M1010_d N_A_639_392#_M1010_g N_A_888_406#_M1010_s VNB NSHORT
+ L=0.15 W=0.64 AD=0.1824 AS=0.0896 PD=1.85 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1026 N_A_1035_74#_M1026_d N_A_639_392#_M1026_g N_A_888_406#_M1010_s VNB NSHORT
+ L=0.15 W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1000 N_A_1035_74#_M1026_d N_RESET_B_M1000_g N_VGND_M1000_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.1 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1023 N_A_1035_74#_M1023_d N_RESET_B_M1023_g N_VGND_M1000_s VNB NSHORT L=0.15
+ W=0.64 AD=0.1824 AS=0.0896 PD=1.85 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.5 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1003 N_VGND_M1003_d N_A_888_406#_M1003_g N_Q_M1003_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.5 A=0.111 P=1.78 MULT=1
MM1011 N_VGND_M1011_d N_A_888_406#_M1011_g N_Q_M1003_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1024 N_VGND_M1011_d N_A_888_406#_M1024_g N_Q_M1024_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1029 N_VGND_M1029_d N_A_888_406#_M1029_g N_Q_M1024_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1014 N_VPWR_M1014_d N_D_M1014_g N_A_27_136#_M1014_s VPB PHIGHVT L=0.15 W=0.84
+ AD=0.168 AS=0.2478 PD=1.24 PS=2.27 NRD=14.0658 NRS=2.3443 M=1 R=5.6 SA=75000.2
+ SB=75000.8 A=0.126 P=1.98 MULT=1
MM1027 N_A_232_98#_M1027_d N_GATE_N_M1027_g N_VPWR_M1014_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.2478 AS=0.168 PD=2.27 PS=1.24 NRD=2.3443 NRS=14.0658 M=1 R=5.6
+ SA=75000.8 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1012 N_VPWR_M1012_d N_A_232_98#_M1012_g N_A_348_392#_M1012_s VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.235793 AS=0.2478 PD=1.53391 PS=2.27 NRD=52.9142 NRS=2.3443
+ M=1 R=5.6 SA=75000.2 SB=75003.2 A=0.126 P=1.98 MULT=1
MM1006 A_561_392# N_A_27_136#_M1006_g N_VPWR_M1012_d VPB PHIGHVT L=0.15 W=1
+ AD=0.12 AS=0.280707 PD=1.24 PS=1.82609 NRD=12.7853 NRS=19.6803 M=1 R=6.66667
+ SA=75000.8 SB=75003.1 A=0.15 P=2.3 MULT=1
MM1019 N_A_639_392#_M1019_d N_A_348_392#_M1019_g A_561_392# VPB PHIGHVT L=0.15
+ W=1 AD=0.237394 AS=0.12 PD=1.95775 PS=1.24 NRD=1.9503 NRS=12.7853 M=1
+ R=6.66667 SA=75001.1 SB=75002.7 A=0.15 P=2.3 MULT=1
MM1005 A_747_504# N_A_232_98#_M1005_g N_A_639_392#_M1019_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1512 AS=0.0997056 PD=1.14 PS=0.822254 NRD=143.042 NRS=85.5374 M=1
+ R=2.8 SA=75001.6 SB=75005.5 A=0.063 P=1.14 MULT=1
MM1020 N_VPWR_M1020_d N_A_888_406#_M1020_g A_747_504# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1421 AS=0.1512 PD=1.06 PS=1.14 NRD=4.6886 NRS=143.042 M=1 R=2.8
+ SA=75002.5 SB=75004.7 A=0.063 P=1.14 MULT=1
MM1001 N_A_888_406#_M1001_d N_A_639_392#_M1001_g N_VPWR_M1020_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.126 AS=0.2842 PD=1.14 PS=2.12 NRD=2.3443 NRS=14.0658 M=1
+ R=5.6 SA=75001.8 SB=75003.8 A=0.126 P=1.98 MULT=1
MM1008 N_A_888_406#_M1001_d N_A_639_392#_M1008_g N_VPWR_M1008_s VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.126 AS=0.147 PD=1.14 PS=1.19 NRD=2.3443 NRS=14.0658 M=1
+ R=5.6 SA=75002.2 SB=75003.3 A=0.126 P=1.98 MULT=1
MM1009 N_VPWR_M1008_s N_RESET_B_M1009_g N_A_888_406#_M1009_s VPB PHIGHVT L=0.15
+ W=0.84 AD=0.147 AS=0.1554 PD=1.19 PS=1.21 NRD=2.3443 NRS=14.0658 M=1 R=5.6
+ SA=75002.7 SB=75002.8 A=0.126 P=1.98 MULT=1
MM1015 N_VPWR_M1015_d N_RESET_B_M1015_g N_A_888_406#_M1009_s VPB PHIGHVT L=0.15
+ W=0.84 AD=0.189086 AS=0.1554 PD=1.33286 PS=1.21 NRD=22.261 NRS=7.0329 M=1
+ R=5.6 SA=75003.2 SB=75002.3 A=0.126 P=1.98 MULT=1
MM1004 N_VPWR_M1015_d N_A_888_406#_M1004_g N_Q_M1004_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.252114 AS=0.168 PD=1.77714 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75002.9 SB=75001.7 A=0.168 P=2.54 MULT=1
MM1013 N_VPWR_M1013_d N_A_888_406#_M1013_g N_Q_M1004_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.196 AS=0.168 PD=1.47 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75003.4 SB=75001.3 A=0.168 P=2.54 MULT=1
MM1022 N_VPWR_M1013_d N_A_888_406#_M1022_g N_Q_M1022_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.196 AS=0.224 PD=1.47 PS=1.52 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75003.9 SB=75000.8 A=0.168 P=2.54 MULT=1
MM1028 N_VPWR_M1028_d N_A_888_406#_M1028_g N_Q_M1022_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.224 PD=2.83 PS=1.52 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75004.4 SB=75000.2 A=0.168 P=2.54 MULT=1
DX30_noxref VNB VPB NWDIODE A=18.5628 P=23.68
*
.include "sky130_fd_sc_ls__dlrtn_4.pxi.spice"
*
.ends
*
*
