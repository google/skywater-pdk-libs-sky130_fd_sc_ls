* File: sky130_fd_sc_ls__fa_2.pex.spice
* Created: Fri Aug 28 13:25:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__FA_2%A 3 5 7 8 10 11 13 14 16 17 19 22 24 26 27 28
+ 29 30 31 32 38 40 43 47 50 56
c225 56 0 1.40112e-19 $X=6.43 $Y=1.515
c226 47 0 1.68414e-19 $X=0.27 $Y=1.465
c227 32 0 2.13543e-19 $X=4.225 $Y=1.665
c228 31 0 1.49152e-19 $X=6.335 $Y=1.665
c229 30 0 1.12499e-19 $X=2.785 $Y=1.665
c230 28 0 1.73388e-19 $X=0.385 $Y=1.665
c231 22 0 1.1376e-19 $X=6.34 $Y=0.765
c232 11 0 1.6514e-19 $X=2.765 $Y=1.66
r233 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.43
+ $Y=1.515 $X2=6.43 $Y2=1.515
r234 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.36
+ $Y=1.41 $X2=4.36 $Y2=1.41
r235 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.84
+ $Y=1.41 $X2=2.84 $Y2=1.41
r236 47 60 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=0.27 $Y=1.465 $X2=0.27
+ $Y2=1.665
r237 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.465 $X2=0.27 $Y2=1.465
r238 43 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=1.665
+ $X2=0.24 $Y2=1.665
r239 40 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=1.665
+ $X2=6.48 $Y2=1.665
r240 38 53 8.69211 $w=3.93e-07 $l=2.8e-07 $layer=LI1_cond $X=4.08 $Y=1.512
+ $X2=4.36 $Y2=1.512
r241 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=1.665
+ $X2=4.08 $Y2=1.665
r242 35 50 8.16535 $w=3.81e-07 $l=3.11288e-07 $layer=LI1_cond $X=2.64 $Y=1.665
+ $X2=2.765 $Y2=1.41
r243 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=1.665
+ $X2=2.64 $Y2=1.665
r244 32 37 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.225 $Y=1.665
+ $X2=4.08 $Y2=1.665
r245 31 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.335 $Y=1.665
+ $X2=6.48 $Y2=1.665
r246 31 32 2.61138 $w=1.4e-07 $l=2.11e-06 $layer=MET1_cond $X=6.335 $Y=1.665
+ $X2=4.225 $Y2=1.665
r247 30 34 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.785 $Y=1.665
+ $X2=2.64 $Y2=1.665
r248 29 37 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.935 $Y=1.665
+ $X2=4.08 $Y2=1.665
r249 29 30 1.42326 $w=1.4e-07 $l=1.15e-06 $layer=MET1_cond $X=3.935 $Y=1.665
+ $X2=2.785 $Y2=1.665
r250 28 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.385 $Y=1.665
+ $X2=0.24 $Y2=1.665
r251 27 34 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.495 $Y=1.665
+ $X2=2.64 $Y2=1.665
r252 27 28 2.61138 $w=1.4e-07 $l=2.11e-06 $layer=MET1_cond $X=2.495 $Y=1.665
+ $X2=0.385 $Y2=1.665
r253 24 55 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=6.355 $Y=1.765
+ $X2=6.43 $Y2=1.515
r254 24 26 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.355 $Y=1.765
+ $X2=6.355 $Y2=2.34
r255 20 55 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=6.34 $Y=1.35
+ $X2=6.43 $Y2=1.515
r256 20 22 299.968 $w=1.5e-07 $l=5.85e-07 $layer=POLY_cond $X=6.34 $Y=1.35
+ $X2=6.34 $Y2=0.765
r257 17 52 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=4.45 $Y=1.245
+ $X2=4.36 $Y2=1.41
r258 17 19 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.45 $Y=1.245
+ $X2=4.45 $Y2=0.765
r259 14 52 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=4.435 $Y=1.66
+ $X2=4.36 $Y2=1.41
r260 14 16 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=4.435 $Y=1.66
+ $X2=4.435 $Y2=2.235
r261 11 49 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=2.765 $Y=1.66
+ $X2=2.84 $Y2=1.41
r262 11 13 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.765 $Y=1.66
+ $X2=2.765 $Y2=2.235
r263 8 49 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=2.75 $Y=1.245
+ $X2=2.84 $Y2=1.41
r264 8 10 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.75 $Y=1.245
+ $X2=2.75 $Y2=0.765
r265 5 46 63.2057 $w=3.69e-07 $l=4.20416e-07 $layer=POLY_cond $X=0.505 $Y=1.815
+ $X2=0.35 $Y2=1.465
r266 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.505 $Y=1.815
+ $X2=0.505 $Y2=2.39
r267 1 46 39.0404 $w=3.69e-07 $l=2.26164e-07 $layer=POLY_cond $X=0.495 $Y=1.3
+ $X2=0.35 $Y2=1.465
r268 1 3 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=0.495 $Y=1.3
+ $X2=0.495 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LS__FA_2%CIN 1 3 4 6 7 9 10 12 13 15 16 18 19 25 26 27
+ 29 30 31 34 38 42 43 49 53 56 60
c172 38 0 1.12499e-19 $X=3.38 $Y=1.41
c173 34 0 1.35287e-19 $X=5.47 $Y=1.41
c174 13 0 1.22946e-19 $X=5.395 $Y=1.66
c175 7 0 1.14658e-19 $X=3.34 $Y=1.66
c176 4 0 1.91229e-19 $X=1.86 $Y=1.245
r177 54 56 2.94811 $w=2.13e-07 $l=5.5e-08 $layer=LI1_cond $X=3.545 $Y=2.042
+ $X2=3.6 $Y2=2.042
r178 53 60 0.428816 $w=2.13e-07 $l=8e-09 $layer=LI1_cond $X=4.088 $Y=2.042
+ $X2=4.08 $Y2=2.042
r179 48 49 34.3324 $w=3.58e-07 $l=2.55e-07 $layer=POLY_cond $X=1.605 $Y=1.452
+ $X2=1.86 $Y2=1.452
r180 43 53 2.14263 $w=2.53e-07 $l=1.12406e-07 $layer=LI1_cond $X=4.126 $Y=1.947
+ $X2=4.088 $Y2=2.042
r181 43 60 2.09048 $w=2.13e-07 $l=3.9e-08 $layer=LI1_cond $X=4.041 $Y=2.042
+ $X2=4.08 $Y2=2.042
r182 42 54 4.65272 $w=1.92e-07 $l=8.5e-08 $layer=LI1_cond $X=3.46 $Y=2.042
+ $X2=3.545 $Y2=2.042
r183 42 43 22.8345 $w=2.13e-07 $l=4.26e-07 $layer=LI1_cond $X=3.615 $Y=2.042
+ $X2=4.041 $Y2=2.042
r184 42 56 0.80403 $w=2.13e-07 $l=1.5e-08 $layer=LI1_cond $X=3.615 $Y=2.042
+ $X2=3.6 $Y2=2.042
r185 38 41 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.38 $Y=1.41
+ $X2=3.38 $Y2=1.575
r186 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.38
+ $Y=1.41 $X2=3.38 $Y2=1.41
r187 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.47
+ $Y=1.41 $X2=5.47 $Y2=1.41
r188 32 34 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=5.47 $Y=1.745
+ $X2=5.47 $Y2=1.41
r189 31 43 21.0404 $w=2.53e-07 $l=4.63825e-07 $layer=LI1_cond $X=4.535 $Y=1.83
+ $X2=4.126 $Y2=1.947
r190 30 32 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.305 $Y=1.83
+ $X2=5.47 $Y2=1.745
r191 30 31 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=5.305 $Y=1.83
+ $X2=4.535 $Y2=1.83
r192 29 42 1.79375 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=3.46 $Y=1.935
+ $X2=3.46 $Y2=2.042
r193 29 41 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=3.46 $Y=1.935
+ $X2=3.46 $Y2=1.575
r194 26 42 4.65272 $w=1.92e-07 $l=8.84308e-08 $layer=LI1_cond $X=3.375 $Y=2.035
+ $X2=3.46 $Y2=2.042
r195 26 27 75.0267 $w=1.68e-07 $l=1.15e-06 $layer=LI1_cond $X=3.375 $Y=2.035
+ $X2=2.225 $Y2=2.035
r196 25 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.14 $Y=1.95
+ $X2=2.225 $Y2=2.035
r197 24 25 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=2.14 $Y=1.575
+ $X2=2.14 $Y2=1.95
r198 22 49 2.69274 $w=3.58e-07 $l=2e-08 $layer=POLY_cond $X=1.88 $Y=1.452
+ $X2=1.86 $Y2=1.452
r199 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.88
+ $Y=1.41 $X2=1.88 $Y2=1.41
r200 19 24 7.64049 $w=3.15e-07 $l=1.95944e-07 $layer=LI1_cond $X=2.055 $Y=1.417
+ $X2=2.14 $Y2=1.575
r201 19 21 6.40246 $w=3.13e-07 $l=1.75e-07 $layer=LI1_cond $X=2.055 $Y=1.417
+ $X2=1.88 $Y2=1.417
r202 16 35 38.5562 $w=2.99e-07 $l=1.88348e-07 $layer=POLY_cond $X=5.52 $Y=1.245
+ $X2=5.47 $Y2=1.41
r203 16 18 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.52 $Y=1.245
+ $X2=5.52 $Y2=0.765
r204 13 35 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=5.395 $Y=1.66
+ $X2=5.47 $Y2=1.41
r205 13 15 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.395 $Y=1.66
+ $X2=5.395 $Y2=2.235
r206 10 39 38.5562 $w=2.99e-07 $l=1.88348e-07 $layer=POLY_cond $X=3.43 $Y=1.245
+ $X2=3.38 $Y2=1.41
r207 10 12 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.43 $Y=1.245
+ $X2=3.43 $Y2=0.765
r208 7 39 52.2586 $w=2.99e-07 $l=2.69258e-07 $layer=POLY_cond $X=3.34 $Y=1.66
+ $X2=3.38 $Y2=1.41
r209 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.34 $Y=1.66
+ $X2=3.34 $Y2=2.235
r210 4 49 23.1716 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.86 $Y=1.245
+ $X2=1.86 $Y2=1.452
r211 4 6 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.86 $Y=1.245 $X2=1.86
+ $Y2=0.765
r212 1 48 23.1716 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.605 $Y=1.66
+ $X2=1.605 $Y2=1.452
r213 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.605 $Y=1.66
+ $X2=1.605 $Y2=2.235
.ends

.subckt PM_SKY130_FD_SC_LS__FA_2%A_336_347# 1 2 7 9 10 12 13 15 16 18 19 22 23
+ 25 26 28 29 31 32 33 35 38 40 44 47 50 53 58 60 61 65
c199 44 0 9.88845e-20 $X=4.93 $Y=1.41
r200 66 69 15.6607 $w=2.77e-07 $l=9e-08 $layer=POLY_cond $X=7 $Y=1.42 $X2=7
+ $Y2=1.33
r201 65 66 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7 $Y=1.42
+ $X2=7 $Y2=1.42
r202 62 65 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=6.85 $Y=1.42 $X2=7
+ $Y2=1.42
r203 55 58 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=1.8 $Y=2.455 $X2=2
+ $Y2=2.455
r204 51 53 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.46 $Y=1.83
+ $X2=1.8 $Y2=1.83
r205 50 62 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.85 $Y=1.255
+ $X2=6.85 $Y2=1.42
r206 49 50 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=6.85 $Y=1.09
+ $X2=6.85 $Y2=1.255
r207 48 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.095 $Y=1.005
+ $X2=4.93 $Y2=1.005
r208 47 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.765 $Y=1.005
+ $X2=6.85 $Y2=1.09
r209 47 48 108.952 $w=1.68e-07 $l=1.67e-06 $layer=LI1_cond $X=6.765 $Y=1.005
+ $X2=5.095 $Y2=1.005
r210 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.93
+ $Y=1.41 $X2=4.93 $Y2=1.41
r211 42 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.93 $Y=1.09
+ $X2=4.93 $Y2=1.005
r212 42 44 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=4.93 $Y=1.09
+ $X2=4.93 $Y2=1.41
r213 41 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.31 $Y=1.005
+ $X2=2.145 $Y2=1.005
r214 40 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.765 $Y=1.005
+ $X2=4.93 $Y2=1.005
r215 40 41 160.166 $w=1.68e-07 $l=2.455e-06 $layer=LI1_cond $X=4.765 $Y=1.005
+ $X2=2.31 $Y2=1.005
r216 36 60 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.145 $Y=0.92
+ $X2=2.145 $Y2=1.005
r217 36 38 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=2.145 $Y=0.92
+ $X2=2.145 $Y2=0.54
r218 35 55 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.8 $Y=2.29 $X2=1.8
+ $Y2=2.455
r219 34 53 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.8 $Y=1.915
+ $X2=1.8 $Y2=1.83
r220 34 35 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.8 $Y=1.915
+ $X2=1.8 $Y2=2.29
r221 32 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.98 $Y=1.005
+ $X2=2.145 $Y2=1.005
r222 32 33 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=1.98 $Y=1.005
+ $X2=1.545 $Y2=1.005
r223 31 51 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.46 $Y=1.745
+ $X2=1.46 $Y2=1.83
r224 30 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.46 $Y=1.09
+ $X2=1.545 $Y2=1.005
r225 30 31 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=1.46 $Y=1.09
+ $X2=1.46 $Y2=1.745
r226 26 29 18.8402 $w=1.65e-07 $l=8.21584e-08 $layer=POLY_cond $X=7.485 $Y=1.255
+ $X2=7.47 $Y2=1.33
r227 26 28 157.453 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=7.485 $Y=1.255
+ $X2=7.485 $Y2=0.765
r228 23 25 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.47 $Y=1.765
+ $X2=7.47 $Y2=2.4
r229 22 23 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=7.47 $Y=1.675
+ $X2=7.47 $Y2=1.765
r230 21 29 18.8402 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=7.47 $Y=1.405
+ $X2=7.47 $Y2=1.33
r231 21 22 104.952 $w=1.8e-07 $l=2.7e-07 $layer=POLY_cond $X=7.47 $Y=1.405
+ $X2=7.47 $Y2=1.675
r232 20 69 17.1008 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.165 $Y=1.33
+ $X2=7 $Y2=1.33
r233 19 29 6.66866 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=7.38 $Y=1.33 $X2=7.47
+ $Y2=1.33
r234 19 20 110.245 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=7.38 $Y=1.33
+ $X2=7.165 $Y2=1.33
r235 16 69 23.1145 $w=2.77e-07 $l=9.87421e-08 $layer=POLY_cond $X=7.055 $Y=1.255
+ $X2=7 $Y2=1.33
r236 16 18 157.453 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=7.055 $Y=1.255
+ $X2=7.055 $Y2=0.765
r237 13 66 70.0964 $w=2.77e-07 $l=3.80657e-07 $layer=POLY_cond $X=6.925 $Y=1.765
+ $X2=7 $Y2=1.42
r238 13 15 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.925 $Y=1.765
+ $X2=6.925 $Y2=2.4
r239 10 45 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=5.02 $Y=1.245
+ $X2=4.93 $Y2=1.41
r240 10 12 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.02 $Y=1.245
+ $X2=5.02 $Y2=0.765
r241 7 45 52.2586 $w=2.99e-07 $l=2.7157e-07 $layer=POLY_cond $X=4.885 $Y=1.66
+ $X2=4.93 $Y2=1.41
r242 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=4.885 $Y=1.66
+ $X2=4.885 $Y2=2.235
r243 2 58 600 $w=1.7e-07 $l=8.65332e-07 $layer=licon1_PDIFF $count=1 $X=1.68
+ $Y=1.735 $X2=2 $Y2=2.455
r244 1 38 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=1.935
+ $Y=0.395 $X2=2.145 $Y2=0.54
.ends

.subckt PM_SKY130_FD_SC_LS__FA_2%B 1 3 4 5 6 9 10 11 12 13 14 15 16 19 22 23 25
+ 26 27 30 33 34 36 37 38 41 44 45 46 47 48 50 51 58 61 65
c198 58 0 1.73388e-19 $X=1 $Y=1.41
c199 41 0 1.40112e-19 $X=5.935 $Y=2.34
r200 61 65 6.56993 $w=2.28e-07 $l=1.15e-07 $layer=LI1_cond $X=0.72 $Y=2.035
+ $X2=0.72 $Y2=1.92
r201 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1 $Y=1.41
+ $X2=1 $Y2=1.41
r202 55 58 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=0.75 $Y=1.41 $X2=1
+ $Y2=1.41
r203 53 55 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.75 $Y=1.575
+ $X2=0.75 $Y2=1.41
r204 53 65 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.75 $Y=1.575
+ $X2=0.75 $Y2=1.92
r205 44 50 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=5.95 $Y=0.765
+ $X2=5.95 $Y2=1.21
r206 39 51 93.4966 $w=1.8e-07 $l=2.35e-07 $layer=POLY_cond $X=5.935 $Y=2.915
+ $X2=5.935 $Y2=3.15
r207 39 41 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.935 $Y=2.915
+ $X2=5.935 $Y2=2.34
r208 38 41 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.935 $Y=1.765
+ $X2=5.935 $Y2=2.34
r209 37 38 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.935 $Y=1.675
+ $X2=5.935 $Y2=1.765
r210 36 50 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.935 $Y=1.3
+ $X2=5.935 $Y2=1.21
r211 36 37 145.766 $w=1.8e-07 $l=3.75e-07 $layer=POLY_cond $X=5.935 $Y=1.3
+ $X2=5.935 $Y2=1.675
r212 35 48 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.935 $Y=3.15
+ $X2=3.845 $Y2=3.15
r213 34 51 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=5.845 $Y=3.15
+ $X2=5.935 $Y2=3.15
r214 34 35 979.383 $w=1.5e-07 $l=1.91e-06 $layer=POLY_cond $X=5.845 $Y=3.15
+ $X2=3.935 $Y2=3.15
r215 33 47 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=3.86 $Y=0.765
+ $X2=3.86 $Y2=1.21
r216 28 48 74.0611 $w=1.8e-07 $l=1.85e-07 $layer=POLY_cond $X=3.845 $Y=2.965
+ $X2=3.845 $Y2=3.15
r217 28 30 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.845 $Y=2.965
+ $X2=3.845 $Y2=2.39
r218 27 30 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.845 $Y=1.815
+ $X2=3.845 $Y2=2.39
r219 26 27 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.845 $Y=1.725
+ $X2=3.845 $Y2=1.815
r220 25 47 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.845 $Y=1.3
+ $X2=3.845 $Y2=1.21
r221 25 26 165.202 $w=1.8e-07 $l=4.25e-07 $layer=POLY_cond $X=3.845 $Y=1.3
+ $X2=3.845 $Y2=1.725
r222 24 46 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.435 $Y=3.15
+ $X2=2.345 $Y2=3.15
r223 23 48 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.755 $Y=3.15
+ $X2=3.845 $Y2=3.15
r224 23 24 676.851 $w=1.5e-07 $l=1.32e-06 $layer=POLY_cond $X=3.755 $Y=3.15
+ $X2=2.435 $Y2=3.15
r225 22 45 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.36 $Y=0.765
+ $X2=2.36 $Y2=1.21
r226 17 19 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.345 $Y=2.81
+ $X2=2.345 $Y2=2.235
r227 16 19 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.345 $Y=1.66
+ $X2=2.345 $Y2=2.235
r228 15 46 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=2.345 $Y=3.075
+ $X2=2.345 $Y2=3.15
r229 14 17 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.345 $Y=2.9
+ $X2=2.345 $Y2=2.81
r230 14 15 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=2.345 $Y=2.9
+ $X2=2.345 $Y2=3.075
r231 13 16 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.345 $Y=1.57
+ $X2=2.345 $Y2=1.66
r232 12 45 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.345 $Y=1.3
+ $X2=2.345 $Y2=1.21
r233 12 13 104.952 $w=1.8e-07 $l=2.7e-07 $layer=POLY_cond $X=2.345 $Y=1.3
+ $X2=2.345 $Y2=1.57
r234 10 46 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.255 $Y=3.15
+ $X2=2.345 $Y2=3.15
r235 10 11 517.894 $w=1.5e-07 $l=1.01e-06 $layer=POLY_cond $X=2.255 $Y=3.15
+ $X2=1.245 $Y2=3.15
r236 7 9 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.155 $Y=2.81
+ $X2=1.155 $Y2=2.235
r237 6 59 50.8664 $w=3.35e-07 $l=3.05369e-07 $layer=POLY_cond $X=1.155 $Y=1.66
+ $X2=1.032 $Y2=1.41
r238 6 9 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.155 $Y=1.66
+ $X2=1.155 $Y2=2.235
r239 5 11 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=1.155 $Y=3.075
+ $X2=1.245 $Y2=3.15
r240 4 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.155 $Y=2.9 $X2=1.155
+ $Y2=2.81
r241 4 5 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=1.155 $Y=2.9
+ $X2=1.155 $Y2=3.075
r242 1 59 38.6365 $w=3.35e-07 $l=2.12238e-07 $layer=POLY_cond $X=1.14 $Y=1.245
+ $X2=1.032 $Y2=1.41
r243 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.14 $Y=1.245 $X2=1.14
+ $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LS__FA_2%A_992_347# 1 2 7 9 12 14 17 18 20 23 25 26 28
+ 33 35 40 45 47
c119 35 0 1.49152e-19 $X=5.17 $Y=2.195
c120 33 0 1.3983e-19 $X=7.965 $Y=2.32
r121 46 49 13.6845 $w=3.17e-07 $l=9e-08 $layer=POLY_cond $X=8.087 $Y=1.485
+ $X2=8.087 $Y2=1.395
r122 45 48 8.49906 $w=3.53e-07 $l=1.65e-07 $layer=LI1_cond $X=8.057 $Y=1.485
+ $X2=8.057 $Y2=1.65
r123 45 47 8.49906 $w=3.53e-07 $l=1.65e-07 $layer=LI1_cond $X=8.057 $Y=1.485
+ $X2=8.057 $Y2=1.32
r124 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.07
+ $Y=1.485 $X2=8.07 $Y2=1.485
r125 40 42 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=5.305 $Y=0.56
+ $X2=5.305 $Y2=0.66
r126 35 37 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=5.17 $Y=2.195
+ $X2=5.17 $Y2=2.405
r127 33 48 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.965 $Y=2.32
+ $X2=7.965 $Y2=1.65
r128 30 47 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=7.965 $Y=0.745
+ $X2=7.965 $Y2=1.32
r129 29 42 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.47 $Y=0.66
+ $X2=5.305 $Y2=0.66
r130 28 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.88 $Y=0.66
+ $X2=7.965 $Y2=0.745
r131 28 29 157.23 $w=1.68e-07 $l=2.41e-06 $layer=LI1_cond $X=7.88 $Y=0.66
+ $X2=5.47 $Y2=0.66
r132 27 37 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.335 $Y=2.405
+ $X2=5.17 $Y2=2.405
r133 26 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.88 $Y=2.405
+ $X2=7.965 $Y2=2.32
r134 26 27 166.037 $w=1.68e-07 $l=2.545e-06 $layer=LI1_cond $X=7.88 $Y=2.405
+ $X2=5.335 $Y2=2.405
r135 21 25 18.8402 $w=1.65e-07 $l=8.21584e-08 $layer=POLY_cond $X=8.625 $Y=1.32
+ $X2=8.61 $Y2=1.395
r136 21 23 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=8.625 $Y=1.32
+ $X2=8.625 $Y2=0.765
r137 18 20 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.61 $Y=1.765
+ $X2=8.61 $Y2=2.4
r138 17 18 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=8.61 $Y=1.675
+ $X2=8.61 $Y2=1.765
r139 16 25 18.8402 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=8.61 $Y=1.47
+ $X2=8.61 $Y2=1.395
r140 16 17 79.6855 $w=1.8e-07 $l=2.05e-07 $layer=POLY_cond $X=8.61 $Y=1.47
+ $X2=8.61 $Y2=1.675
r141 15 49 20.269 $w=1.5e-07 $l=1.83e-07 $layer=POLY_cond $X=8.27 $Y=1.395
+ $X2=8.087 $Y2=1.395
r142 14 25 6.66866 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=8.52 $Y=1.395
+ $X2=8.61 $Y2=1.395
r143 14 15 128.191 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=8.52 $Y=1.395
+ $X2=8.27 $Y2=1.395
r144 10 49 24.856 $w=3.17e-07 $l=1.40584e-07 $layer=POLY_cond $X=8.195 $Y=1.32
+ $X2=8.087 $Y2=1.395
r145 10 12 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=8.195 $Y=1.32
+ $X2=8.195 $Y2=0.765
r146 7 46 56.0264 $w=3.17e-07 $l=3.14388e-07 $layer=POLY_cond $X=8.16 $Y=1.765
+ $X2=8.087 $Y2=1.485
r147 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.16 $Y=1.765
+ $X2=8.16 $Y2=2.4
r148 2 35 300 $w=1.7e-07 $l=5.55158e-07 $layer=licon1_PDIFF $count=2 $X=4.96
+ $Y=1.735 $X2=5.17 $Y2=2.195
r149 1 40 182 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_NDIFF $count=1 $X=5.095
+ $Y=0.395 $X2=5.305 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_LS__FA_2%A_27_378# 1 2 9 13 16 18
c34 16 0 1.68414e-19 $X=0.28 $Y=2.405
r35 18 20 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=1.38 $Y=2.25
+ $X2=1.38 $Y2=2.405
r36 14 16 3.9231 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=0.445 $Y=2.405
+ $X2=0.27 $Y2=2.405
r37 13 20 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.215 $Y=2.405
+ $X2=1.38 $Y2=2.405
r38 13 14 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.215 $Y=2.405
+ $X2=0.445 $Y2=2.405
r39 7 16 2.80976 $w=3.4e-07 $l=8.9861e-08 $layer=LI1_cond $X=0.26 $Y=2.32
+ $X2=0.27 $Y2=2.405
r40 7 9 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=0.26 $Y=2.32 $X2=0.26
+ $Y2=2.035
r41 2 18 300 $w=1.7e-07 $l=5.85214e-07 $layer=licon1_PDIFF $count=2 $X=1.23
+ $Y=1.735 $X2=1.38 $Y2=2.25
r42 1 16 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.89 $X2=0.28 $Y2=2.405
r43 1 9 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.89 $X2=0.26 $Y2=2.035
.ends

.subckt PM_SKY130_FD_SC_LS__FA_2%VPWR 1 2 3 4 5 6 21 25 29 33 35 37 42 43 45 46
+ 47 49 61 72 76 82 85 88 96
r115 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r116 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r117 88 91 11.8458 $w=5.18e-07 $l=5.15e-07 $layer=LI1_cond $X=7.79 $Y=2.815
+ $X2=7.79 $Y2=3.33
r118 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r119 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r120 80 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=8.88 $Y2=3.33
r121 80 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=7.92 $Y2=3.33
r122 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33 $X2=8.4
+ $Y2=3.33
r123 77 91 7.40362 $w=1.7e-07 $l=2.6e-07 $layer=LI1_cond $X=8.05 $Y=3.33
+ $X2=7.79 $Y2=3.33
r124 77 79 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=8.05 $Y=3.33
+ $X2=8.4 $Y2=3.33
r125 76 95 4.0045 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=8.75 $Y=3.33
+ $X2=8.935 $Y2=3.33
r126 76 79 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=8.75 $Y=3.33
+ $X2=8.4 $Y2=3.33
r127 75 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r128 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r129 72 91 7.40362 $w=1.7e-07 $l=2.6e-07 $layer=LI1_cond $X=7.53 $Y=3.33
+ $X2=7.79 $Y2=3.33
r130 72 74 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=7.53 $Y=3.33 $X2=7.44
+ $Y2=3.33
r131 71 75 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=7.44 $Y2=3.33
r132 70 71 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r133 67 70 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.56 $Y=3.33
+ $X2=6.48 $Y2=3.33
r134 65 85 9.56655 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=4.29 $Y=3.33
+ $X2=4.097 $Y2=3.33
r135 65 67 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=4.29 $Y=3.33
+ $X2=4.56 $Y2=3.33
r136 64 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r137 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r138 61 85 9.56655 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=3.905 $Y=3.33
+ $X2=4.097 $Y2=3.33
r139 61 63 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.905 $Y=3.33
+ $X2=3.6 $Y2=3.33
r140 60 64 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r141 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r142 57 60 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r143 57 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r144 56 59 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r145 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r146 54 82 9.73034 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=1.01 $Y=3.33
+ $X2=0.812 $Y2=3.33
r147 54 56 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.01 $Y=3.33
+ $X2=1.2 $Y2=3.33
r148 52 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r149 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r150 49 82 9.73034 $w=1.7e-07 $l=1.97e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.812 $Y2=3.33
r151 49 51 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.24 $Y2=3.33
r152 47 71 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=6.48 $Y2=3.33
r153 47 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r154 47 67 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r155 45 70 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=6.535 $Y=3.33
+ $X2=6.48 $Y2=3.33
r156 45 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.535 $Y=3.33
+ $X2=6.7 $Y2=3.33
r157 44 74 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=6.865 $Y=3.33
+ $X2=7.44 $Y2=3.33
r158 44 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.865 $Y=3.33
+ $X2=6.7 $Y2=3.33
r159 42 59 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.825 $Y=3.33
+ $X2=2.64 $Y2=3.33
r160 42 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.825 $Y=3.33
+ $X2=2.99 $Y2=3.33
r161 41 63 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=3.155 $Y=3.33
+ $X2=3.6 $Y2=3.33
r162 41 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.155 $Y=3.33
+ $X2=2.99 $Y2=3.33
r163 37 40 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=8.875 $Y=1.985
+ $X2=8.875 $Y2=2.815
r164 35 95 3.13866 $w=2.5e-07 $l=1.11018e-07 $layer=LI1_cond $X=8.875 $Y=3.245
+ $X2=8.935 $Y2=3.33
r165 35 40 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=8.875 $Y=3.245
+ $X2=8.875 $Y2=2.815
r166 31 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.7 $Y=3.245 $X2=6.7
+ $Y2=3.33
r167 31 33 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=6.7 $Y=3.245
+ $X2=6.7 $Y2=2.78
r168 27 85 1.35792 $w=3.85e-07 $l=8.5e-08 $layer=LI1_cond $X=4.097 $Y=3.245
+ $X2=4.097 $Y2=3.33
r169 27 29 14.9668 $w=3.83e-07 $l=5e-07 $layer=LI1_cond $X=4.097 $Y=3.245
+ $X2=4.097 $Y2=2.745
r170 23 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.99 $Y=3.245
+ $X2=2.99 $Y2=3.33
r171 23 25 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=2.99 $Y=3.245
+ $X2=2.99 $Y2=2.455
r172 19 82 1.43204 $w=3.95e-07 $l=8.5e-08 $layer=LI1_cond $X=0.812 $Y=3.245
+ $X2=0.812 $Y2=3.33
r173 19 21 14.5879 $w=3.93e-07 $l=5e-07 $layer=LI1_cond $X=0.812 $Y=3.245
+ $X2=0.812 $Y2=2.745
r174 6 40 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=8.685
+ $Y=1.84 $X2=8.835 $Y2=2.815
r175 6 37 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=8.685
+ $Y=1.84 $X2=8.835 $Y2=1.985
r176 5 88 600 $w=1.7e-07 $l=1.09064e-06 $layer=licon1_PDIFF $count=1 $X=7.545
+ $Y=1.84 $X2=7.79 $Y2=2.815
r177 4 33 600 $w=1.7e-07 $l=1.06649e-06 $layer=licon1_PDIFF $count=1 $X=6.43
+ $Y=1.84 $X2=6.7 $Y2=2.78
r178 3 29 600 $w=1.7e-07 $l=9.3843e-07 $layer=licon1_PDIFF $count=1 $X=3.92
+ $Y=1.89 $X2=4.095 $Y2=2.745
r179 2 25 600 $w=1.7e-07 $l=7.91454e-07 $layer=licon1_PDIFF $count=1 $X=2.84
+ $Y=1.735 $X2=2.99 $Y2=2.455
r180 1 21 600 $w=1.7e-07 $l=9.63159e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.89 $X2=0.81 $Y2=2.745
.ends

.subckt PM_SKY130_FD_SC_LS__FA_2%A_683_347# 1 2 9 15 16
c34 15 0 1.22946e-19 $X=4.66 $Y=2.44
c35 9 0 1.6514e-19 $X=3.57 $Y=2.405
r36 15 16 9.39634 $w=4.78e-07 $l=1.65e-07 $layer=LI1_cond $X=4.66 $Y=2.515
+ $X2=4.495 $Y2=2.515
r37 9 12 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=3.57 $Y=2.405 $X2=3.57
+ $Y2=2.485
r38 8 9 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.735 $Y=2.405
+ $X2=3.57 $Y2=2.405
r39 8 16 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=3.735 $Y=2.405
+ $X2=4.495 $Y2=2.405
r40 2 15 600 $w=1.7e-07 $l=7.76386e-07 $layer=licon1_PDIFF $count=1 $X=4.51
+ $Y=1.735 $X2=4.66 $Y2=2.44
r41 1 12 600 $w=1.7e-07 $l=8.23863e-07 $layer=licon1_PDIFF $count=1 $X=3.415
+ $Y=1.735 $X2=3.57 $Y2=2.485
.ends

.subckt PM_SKY130_FD_SC_LS__FA_2%COUT 1 2 7 12 13 16
c29 7 0 1.1376e-19 $X=7.385 $Y=1
r30 13 16 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.47 $Y=1.985
+ $X2=7.385 $Y2=1.985
r31 13 16 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=7.37 $Y=1.985
+ $X2=7.385 $Y2=1.985
r32 13 18 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=7.37 $Y=1.985
+ $X2=7.195 $Y2=1.985
r33 12 13 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.47 $Y=1.82
+ $X2=7.47 $Y2=1.985
r34 11 12 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=7.47 $Y=1.085
+ $X2=7.47 $Y2=1.82
r35 7 11 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.385 $Y=1
+ $X2=7.47 $Y2=1.085
r36 7 9 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=7.385 $Y=1 $X2=7.27
+ $Y2=1
r37 2 18 600 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=1 $X=7 $Y=1.84
+ $X2=7.195 $Y2=1.985
r38 1 9 182 $w=1.7e-07 $l=6.71361e-07 $layer=licon1_NDIFF $count=1 $X=7.13
+ $Y=0.395 $X2=7.27 $Y2=1
.ends

.subckt PM_SKY130_FD_SC_LS__FA_2%SUM 1 2 9 13 14 15 16 23 32
r40 21 23 1.2336 $w=3.53e-07 $l=3.8e-08 $layer=LI1_cond $X=8.397 $Y=1.997
+ $X2=8.397 $Y2=2.035
r41 15 16 12.0114 $w=3.53e-07 $l=3.7e-07 $layer=LI1_cond $X=8.397 $Y=2.405
+ $X2=8.397 $Y2=2.775
r42 14 21 0.779116 $w=3.53e-07 $l=2.4e-08 $layer=LI1_cond $X=8.397 $Y=1.973
+ $X2=8.397 $Y2=1.997
r43 14 32 8.1095 $w=3.53e-07 $l=1.53e-07 $layer=LI1_cond $X=8.397 $Y=1.973
+ $X2=8.397 $Y2=1.82
r44 14 15 11.2647 $w=3.53e-07 $l=3.47e-07 $layer=LI1_cond $X=8.397 $Y=2.058
+ $X2=8.397 $Y2=2.405
r45 14 23 0.746653 $w=3.53e-07 $l=2.3e-08 $layer=LI1_cond $X=8.397 $Y=2.058
+ $X2=8.397 $Y2=2.035
r46 13 32 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.49 $Y=1.15
+ $X2=8.49 $Y2=1.82
r47 7 13 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=8.41 $Y=0.985
+ $X2=8.41 $Y2=1.15
r48 7 9 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=8.41 $Y=0.985
+ $X2=8.41 $Y2=0.54
r49 2 14 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=8.235
+ $Y=1.84 $X2=8.385 $Y2=1.985
r50 2 16 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=8.235
+ $Y=1.84 $X2=8.385 $Y2=2.815
r51 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.27
+ $Y=0.395 $X2=8.41 $Y2=0.54
.ends

.subckt PM_SKY130_FD_SC_LS__FA_2%A_27_79# 1 2 9 11 12 14 15 17
c36 11 0 1.91229e-19 $X=1.035 $Y=0.99
r37 15 17 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.205 $Y=0.585
+ $X2=1.5 $Y2=0.585
r38 13 15 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.12 $Y=0.75
+ $X2=1.205 $Y2=0.585
r39 13 14 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=1.12 $Y=0.75
+ $X2=1.12 $Y2=0.905
r40 11 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.035 $Y=0.99
+ $X2=1.12 $Y2=0.905
r41 11 12 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=1.035 $Y=0.99
+ $X2=0.445 $Y2=0.99
r42 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=0.905
+ $X2=0.445 $Y2=0.99
r43 7 9 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=0.28 $Y=0.905
+ $X2=0.28 $Y2=0.54
r44 2 17 182 $w=1.7e-07 $l=3.67933e-07 $layer=licon1_NDIFF $count=1 $X=1.215
+ $Y=0.395 $X2=1.5 $Y2=0.585
r45 1 9 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.395 $X2=0.28 $Y2=0.54
.ends

.subckt PM_SKY130_FD_SC_LS__FA_2%VGND 1 2 3 4 5 6 21 25 27 29 31 33 38 46 51 56
+ 61 67 70 74 88 95
r100 94 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r101 88 91 8.50545 $w=4.48e-07 $l=3.2e-07 $layer=LI1_cond $X=7.84 $Y=0 $X2=7.84
+ $Y2=0.32
r102 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r103 74 77 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=4.155 $Y=0
+ $X2=4.155 $Y2=0.325
r104 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r105 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r106 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r107 65 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=8.88
+ $Y2=0
r108 65 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=7.92
+ $Y2=0
r109 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r110 62 88 6.50032 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=8.065 $Y=0 $X2=7.84
+ $Y2=0
r111 62 64 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=8.065 $Y=0 $X2=8.4
+ $Y2=0
r112 61 94 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=8.755 $Y=0
+ $X2=8.937 $Y2=0
r113 61 64 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=8.755 $Y=0 $X2=8.4
+ $Y2=0
r114 60 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=7.92
+ $Y2=0
r115 60 82 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=6.48
+ $Y2=0
r116 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r117 57 59 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=6.925 $Y=0
+ $X2=7.44 $Y2=0
r118 56 88 6.50032 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=7.615 $Y=0 $X2=7.84
+ $Y2=0
r119 56 59 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=7.615 $Y=0
+ $X2=7.44 $Y2=0
r120 52 74 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.32 $Y=0 $X2=4.155
+ $Y2=0
r121 52 54 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=4.32 $Y=0 $X2=4.56
+ $Y2=0
r122 51 84 8.41198 $w=4.53e-07 $l=3.2e-07 $layer=LI1_cond $X=6.697 $Y=0
+ $X2=6.697 $Y2=0.32
r123 51 57 6.56868 $w=1.7e-07 $l=2.28e-07 $layer=LI1_cond $X=6.697 $Y=0
+ $X2=6.925 $Y2=0
r124 51 82 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r125 51 54 124.61 $w=1.68e-07 $l=1.91e-06 $layer=LI1_cond $X=6.47 $Y=0 $X2=4.56
+ $Y2=0
r126 50 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r127 50 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r128 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r129 47 70 11.4275 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=3.31 $Y=0 $X2=3.055
+ $Y2=0
r130 47 49 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=3.31 $Y=0 $X2=3.6
+ $Y2=0
r131 46 74 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.99 $Y=0 $X2=4.155
+ $Y2=0
r132 46 49 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=3.99 $Y=0 $X2=3.6
+ $Y2=0
r133 45 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r134 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r135 42 45 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r136 42 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r137 41 44 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r138 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r139 39 67 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.865 $Y=0 $X2=0.74
+ $Y2=0
r140 39 41 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.865 $Y=0 $X2=1.2
+ $Y2=0
r141 38 70 11.4275 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=2.8 $Y=0 $X2=3.055
+ $Y2=0
r142 38 44 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=2.8 $Y=0 $X2=2.64
+ $Y2=0
r143 36 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r144 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r145 33 67 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.74
+ $Y2=0
r146 33 35 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=0
+ $X2=0.24 $Y2=0
r147 31 82 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.56 $Y=0
+ $X2=6.48 $Y2=0
r148 31 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r149 31 54 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r150 27 94 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=8.88 $Y=0.085
+ $X2=8.937 $Y2=0
r151 27 29 20.9745 $w=2.48e-07 $l=4.55e-07 $layer=LI1_cond $X=8.88 $Y=0.085
+ $X2=8.88 $Y2=0.54
r152 23 70 2.12513 $w=5.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.055 $Y=0.085
+ $X2=3.055 $Y2=0
r153 23 25 10.6709 $w=5.08e-07 $l=4.55e-07 $layer=LI1_cond $X=3.055 $Y=0.085
+ $X2=3.055 $Y2=0.54
r154 19 67 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.74 $Y=0.085
+ $X2=0.74 $Y2=0
r155 19 21 21.6659 $w=2.48e-07 $l=4.7e-07 $layer=LI1_cond $X=0.74 $Y=0.085
+ $X2=0.74 $Y2=0.555
r156 6 29 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.7
+ $Y=0.395 $X2=8.84 $Y2=0.54
r157 5 91 182 $w=1.7e-07 $l=3.15278e-07 $layer=licon1_NDIFF $count=1 $X=7.56
+ $Y=0.395 $X2=7.84 $Y2=0.32
r158 4 84 182 $w=1.7e-07 $l=3.15278e-07 $layer=licon1_NDIFF $count=1 $X=6.415
+ $Y=0.395 $X2=6.695 $Y2=0.32
r159 3 77 182 $w=1.7e-07 $l=2.52587e-07 $layer=licon1_NDIFF $count=1 $X=3.935
+ $Y=0.395 $X2=4.155 $Y2=0.325
r160 2 25 182 $w=1.7e-07 $l=2.93684e-07 $layer=licon1_NDIFF $count=1 $X=2.825
+ $Y=0.395 $X2=3.055 $Y2=0.54
r161 1 21 182 $w=1.7e-07 $l=2.78747e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.395 $X2=0.78 $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_LS__FA_2%A_701_79# 1 2 10 15 16
r29 15 16 10.9068 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=4.735 $Y=0.585
+ $X2=4.5 $Y2=0.585
r30 10 12 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=3.645 $Y=0.56
+ $X2=3.645 $Y2=0.665
r31 8 12 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.81 $Y=0.665
+ $X2=3.645 $Y2=0.665
r32 8 16 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.81 $Y=0.665 $X2=4.5
+ $Y2=0.665
r33 2 15 182 $w=1.7e-07 $l=2.89828e-07 $layer=licon1_NDIFF $count=1 $X=4.525
+ $Y=0.395 $X2=4.735 $Y2=0.585
r34 1 10 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=3.505
+ $Y=0.395 $X2=3.645 $Y2=0.56
.ends

