* File: sky130_fd_sc_ls__o31a_2.spice
* Created: Wed Sep  2 11:22:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__o31a_2.pex.spice"
.subckt sky130_fd_sc_ls__o31a_2  VNB VPB A1 A2 A3 B1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B1	B1
* A3	A3
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1005 N_X_M1005_d N_A_55_264#_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.2627 PD=1.02 PS=2.19 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75000.3
+ SB=75003 A=0.111 P=1.78 MULT=1
MM1006 N_X_M1005_d N_A_55_264#_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1554 PD=1.02 PS=1.16 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75000.7
+ SB=75002.6 A=0.111 P=1.78 MULT=1
MM1010 N_A_328_74#_M1010_d N_A1_M1010_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.74
+ AD=0.12765 AS=0.1554 PD=1.085 PS=1.16 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.3
+ SB=75002 A=0.111 P=1.78 MULT=1
MM1000 N_VGND_M1000_d N_A2_M1000_g N_A_328_74#_M1010_d VNB NSHORT L=0.15 W=0.74
+ AD=0.1554 AS=0.12765 PD=1.16 PS=1.085 NRD=5.664 NRS=10.536 M=1 R=4.93333
+ SA=75001.8 SB=75001.5 A=0.111 P=1.78 MULT=1
MM1009 N_A_328_74#_M1009_d N_A3_M1009_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.74
+ AD=0.18315 AS=0.1554 PD=1.235 PS=1.16 NRD=17.016 NRS=17.016 M=1 R=4.93333
+ SA=75002.3 SB=75000.9 A=0.111 P=1.78 MULT=1
MM1002 N_A_55_264#_M1002_d N_B1_M1002_g N_A_328_74#_M1009_d VNB NSHORT L=0.15
+ W=0.74 AD=0.2627 AS=0.18315 PD=2.19 PS=1.235 NRD=11.34 NRS=17.832 M=1
+ R=4.93333 SA=75003 SB=75000.3 A=0.111 P=1.78 MULT=1
MM1007 N_VPWR_M1007_d N_A_55_264#_M1007_g N_X_M1007_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.1988 PD=2.83 PS=1.475 NRD=1.7533 NRS=6.1464 M=1 R=7.46667
+ SA=75000.2 SB=75002.8 A=0.168 P=2.54 MULT=1
MM1008 N_VPWR_M1008_d N_A_55_264#_M1008_g N_X_M1007_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.278309 AS=0.1988 PD=1.70642 PS=1.475 NRD=18.4589 NRS=7.0329 M=1 R=7.46667
+ SA=75000.7 SB=75002.3 A=0.168 P=2.54 MULT=1
MM1004 A_346_392# N_A1_M1004_g N_VPWR_M1008_d VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.248491 PD=1.27 PS=1.52358 NRD=15.7403 NRS=21.67 M=1 R=6.66667 SA=75001.4
+ SB=75001.9 A=0.15 P=2.3 MULT=1
MM1001 A_430_392# N_A2_M1001_g A_346_392# VPB PHIGHVT L=0.15 W=1 AD=0.21
+ AS=0.135 PD=1.42 PS=1.27 NRD=30.5153 NRS=15.7403 M=1 R=6.66667 SA=75001.8
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1011 N_A_55_264#_M1011_d N_A3_M1011_g A_430_392# VPB PHIGHVT L=0.15 W=1
+ AD=0.195 AS=0.21 PD=1.39 PS=1.42 NRD=13.7703 NRS=30.5153 M=1 R=6.66667
+ SA=75002.4 SB=75000.9 A=0.15 P=2.3 MULT=1
MM1003 N_VPWR_M1003_d N_B1_M1003_g N_A_55_264#_M1011_d VPB PHIGHVT L=0.15 W=1
+ AD=0.445 AS=0.195 PD=2.89 PS=1.39 NRD=31.5003 NRS=7.8603 M=1 R=6.66667
+ SA=75002.9 SB=75000.4 A=0.15 P=2.3 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8492 P=12.16
*
.include "sky130_fd_sc_ls__o31a_2.pxi.spice"
*
.ends
*
*
