* File: sky130_fd_sc_ls__a311o_1.pxi.spice
* Created: Wed Sep  2 10:51:29 2020
* 
x_PM_SKY130_FD_SC_LS__A311O_1%A_89_270# N_A_89_270#_M1004_d N_A_89_270#_M1000_d
+ N_A_89_270#_M1007_d N_A_89_270#_c_75_n N_A_89_270#_M1010_g N_A_89_270#_c_76_n
+ N_A_89_270#_M1003_g N_A_89_270#_c_77_n N_A_89_270#_c_78_n N_A_89_270#_c_79_n
+ N_A_89_270#_c_86_n N_A_89_270#_c_80_n N_A_89_270#_c_81_n N_A_89_270#_c_87_n
+ N_A_89_270#_c_82_n N_A_89_270#_c_83_n PM_SKY130_FD_SC_LS__A311O_1%A_89_270#
x_PM_SKY130_FD_SC_LS__A311O_1%A3 N_A3_c_171_n N_A3_M1009_g N_A3_M1001_g A3
+ PM_SKY130_FD_SC_LS__A311O_1%A3
x_PM_SKY130_FD_SC_LS__A311O_1%A2 N_A2_c_201_n N_A2_M1002_g N_A2_M1008_g A2
+ PM_SKY130_FD_SC_LS__A311O_1%A2
x_PM_SKY130_FD_SC_LS__A311O_1%A1 N_A1_M1004_g N_A1_c_233_n N_A1_c_234_n
+ N_A1_c_239_n N_A1_M1005_g A1 A1 N_A1_c_235_n N_A1_c_236_n N_A1_c_237_n
+ PM_SKY130_FD_SC_LS__A311O_1%A1
x_PM_SKY130_FD_SC_LS__A311O_1%B1 N_B1_M1011_g N_B1_c_285_n N_B1_c_290_n
+ N_B1_M1006_g N_B1_c_286_n B1 N_B1_c_288_n PM_SKY130_FD_SC_LS__A311O_1%B1
x_PM_SKY130_FD_SC_LS__A311O_1%C1 N_C1_c_328_n N_C1_c_335_n N_C1_M1007_g
+ N_C1_M1000_g N_C1_c_330_n N_C1_c_331_n C1 N_C1_c_332_n N_C1_c_333_n
+ PM_SKY130_FD_SC_LS__A311O_1%C1
x_PM_SKY130_FD_SC_LS__A311O_1%X N_X_M1003_s N_X_M1010_s N_X_c_371_n N_X_c_372_n
+ X X X X N_X_c_373_n PM_SKY130_FD_SC_LS__A311O_1%X
x_PM_SKY130_FD_SC_LS__A311O_1%VPWR N_VPWR_M1010_d N_VPWR_M1002_d N_VPWR_c_393_n
+ N_VPWR_c_394_n N_VPWR_c_395_n N_VPWR_c_396_n VPWR N_VPWR_c_397_n
+ N_VPWR_c_392_n N_VPWR_c_399_n PM_SKY130_FD_SC_LS__A311O_1%VPWR
x_PM_SKY130_FD_SC_LS__A311O_1%A_258_392# N_A_258_392#_M1009_d
+ N_A_258_392#_M1005_d N_A_258_392#_c_433_n N_A_258_392#_c_434_n
+ N_A_258_392#_c_435_n N_A_258_392#_c_436_n N_A_258_392#_c_437_n
+ PM_SKY130_FD_SC_LS__A311O_1%A_258_392#
x_PM_SKY130_FD_SC_LS__A311O_1%VGND N_VGND_M1003_d N_VGND_M1011_d N_VGND_c_472_n
+ N_VGND_c_473_n N_VGND_c_474_n N_VGND_c_475_n VGND N_VGND_c_476_n
+ N_VGND_c_477_n N_VGND_c_478_n N_VGND_c_479_n PM_SKY130_FD_SC_LS__A311O_1%VGND
cc_1 VNB N_A_89_270#_c_75_n 0.0294182f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.765
cc_2 VNB N_A_89_270#_c_76_n 0.0215076f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=1.35
cc_3 VNB N_A_89_270#_c_77_n 0.0109532f $X=-0.19 $Y=-0.245 $X2=2.24 $Y2=1.195
cc_4 VNB N_A_89_270#_c_78_n 0.00627074f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=1.195
cc_5 VNB N_A_89_270#_c_79_n 0.0106288f $X=-0.19 $Y=-0.245 $X2=3.245 $Y2=1.53
cc_6 VNB N_A_89_270#_c_80_n 0.0175711f $X=-0.19 $Y=-0.245 $X2=3.41 $Y2=1.105
cc_7 VNB N_A_89_270#_c_81_n 0.003271f $X=-0.19 $Y=-0.245 $X2=2.405 $Y2=1.005
cc_8 VNB N_A_89_270#_c_82_n 0.00228403f $X=-0.19 $Y=-0.245 $X2=3.34 $Y2=1.94
cc_9 VNB N_A_89_270#_c_83_n 0.00770964f $X=-0.19 $Y=-0.245 $X2=3.41 $Y2=1.53
cc_10 VNB N_A3_c_171_n 0.019133f $X=-0.19 $Y=-0.245 $X2=2.265 $Y2=0.615
cc_11 VNB N_A3_M1001_g 0.0239645f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB A3 9.08959e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A2_c_201_n 0.0160683f $X=-0.19 $Y=-0.245 $X2=2.265 $Y2=0.615
cc_14 VNB N_A2_M1008_g 0.0208933f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB A2 0.00320338f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A1_M1004_g 0.00828724f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A1_c_233_n 0.00553125f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A1_c_234_n 0.011874f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A1_c_235_n 0.0466861f $X=-0.19 $Y=-0.245 $X2=2.24 $Y2=1.195
cc_20 VNB N_A1_c_236_n 9.2097e-19 $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=1.195
cc_21 VNB N_A1_c_237_n 0.00608405f $X=-0.19 $Y=-0.245 $X2=3.34 $Y2=2.175
cc_22 VNB N_B1_M1011_g 0.00907604f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_B1_c_285_n 0.00809716f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_B1_c_286_n 0.00997949f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=2.4
cc_25 VNB B1 0.00737349f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=2.4
cc_26 VNB N_B1_c_288_n 0.0353796f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=0.87
cc_27 VNB N_C1_c_328_n 0.0103317f $X=-0.19 $Y=-0.245 $X2=3.27 $Y2=0.615
cc_28 VNB N_C1_M1000_g 0.0111186f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_C1_c_330_n 0.0199393f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=2.4
cc_30 VNB N_C1_c_331_n 0.0137028f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=0.87
cc_31 VNB N_C1_c_332_n 0.0599949f $X=-0.19 $Y=-0.245 $X2=3.245 $Y2=1.53
cc_32 VNB N_C1_c_333_n 0.0126535f $X=-0.19 $Y=-0.245 $X2=2.57 $Y2=1.53
cc_33 VNB N_X_c_371_n 0.0182499f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_X_c_372_n 0.0228556f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=2.4
cc_35 VNB N_X_c_373_n 0.0234973f $X=-0.19 $Y=-0.245 $X2=2.405 $Y2=1.005
cc_36 VNB N_VPWR_c_392_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=1.515
cc_37 VNB N_VGND_c_472_n 0.0203545f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_473_n 0.00567404f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=2.4
cc_39 VNB N_VGND_c_474_n 0.0256231f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=0.87
cc_40 VNB N_VGND_c_475_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=0.87
cc_41 VNB N_VGND_c_476_n 0.0507439f $X=-0.19 $Y=-0.245 $X2=3.41 $Y2=1.445
cc_42 VNB N_VGND_c_477_n 0.0181991f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=1.195
cc_43 VNB N_VGND_c_478_n 0.249518f $X=-0.19 $Y=-0.245 $X2=0.712 $Y2=1.515
cc_44 VNB N_VGND_c_479_n 0.00270401f $X=-0.19 $Y=-0.245 $X2=2.405 $Y2=1.005
cc_45 VPB N_A_89_270#_c_75_n 0.034419f $X=-0.19 $Y=1.66 $X2=0.535 $Y2=1.765
cc_46 VPB N_A_89_270#_c_78_n 0.00421697f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=1.195
cc_47 VPB N_A_89_270#_c_86_n 0.0405767f $X=-0.19 $Y=1.66 $X2=3.27 $Y2=2.815
cc_48 VPB N_A_89_270#_c_87_n 0.0116412f $X=-0.19 $Y=1.66 $X2=3.27 $Y2=2.105
cc_49 VPB N_A_89_270#_c_82_n 0.0159605f $X=-0.19 $Y=1.66 $X2=3.34 $Y2=1.94
cc_50 VPB N_A3_c_171_n 0.0387189f $X=-0.19 $Y=1.66 $X2=2.265 $Y2=0.615
cc_51 VPB A3 8.81819e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_A2_c_201_n 0.0340515f $X=-0.19 $Y=1.66 $X2=2.265 $Y2=0.615
cc_53 VPB A2 0.00214309f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_A1_c_234_n 0.00734272f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_A1_c_239_n 0.0227973f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_B1_c_285_n 0.00727124f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_B1_c_290_n 0.021758f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_C1_c_328_n 0.00771927f $X=-0.19 $Y=1.66 $X2=3.27 $Y2=0.615
cc_59 VPB N_C1_c_335_n 0.0256513f $X=-0.19 $Y=1.66 $X2=3.12 $Y2=1.96
cc_60 VPB X 0.00695105f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=1.195
cc_61 VPB X 0.0408286f $X=-0.19 $Y=1.66 $X2=3.41 $Y2=1.105
cc_62 VPB N_X_c_373_n 0.00919396f $X=-0.19 $Y=1.66 $X2=2.405 $Y2=1.005
cc_63 VPB N_VPWR_c_393_n 0.0142889f $X=-0.19 $Y=1.66 $X2=0.535 $Y2=2.4
cc_64 VPB N_VPWR_c_394_n 0.0093235f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=1.195
cc_65 VPB N_VPWR_c_395_n 0.0196495f $X=-0.19 $Y=1.66 $X2=3.34 $Y2=2.175
cc_66 VPB N_VPWR_c_396_n 0.00555219f $X=-0.19 $Y=1.66 $X2=3.34 $Y2=2.815
cc_67 VPB N_VPWR_c_397_n 0.0514544f $X=-0.19 $Y=1.66 $X2=0.645 $Y2=1.515
cc_68 VPB N_VPWR_c_392_n 0.0795417f $X=-0.19 $Y=1.66 $X2=0.645 $Y2=1.515
cc_69 VPB N_VPWR_c_399_n 0.028772f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_A_258_392#_c_433_n 0.0041202f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_A_258_392#_c_434_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_A_258_392#_c_435_n 0.00465816f $X=-0.19 $Y=1.66 $X2=0.535 $Y2=2.4
cc_73 VPB N_A_258_392#_c_436_n 0.00339359f $X=-0.19 $Y=1.66 $X2=0.735 $Y2=1.35
cc_74 VPB N_A_258_392#_c_437_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0.735 $Y2=0.87
cc_75 N_A_89_270#_c_75_n N_A3_c_171_n 0.0356408f $X=0.535 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_76 N_A_89_270#_c_77_n N_A3_c_171_n 0.00302456f $X=2.24 $Y=1.195 $X2=-0.19
+ $Y2=-0.245
cc_77 N_A_89_270#_c_78_n N_A3_c_171_n 0.00163481f $X=0.945 $Y=1.195 $X2=-0.19
+ $Y2=-0.245
cc_78 N_A_89_270#_c_76_n N_A3_M1001_g 0.0233429f $X=0.735 $Y=1.35 $X2=0 $Y2=0
cc_79 N_A_89_270#_c_77_n N_A3_M1001_g 0.0154265f $X=2.24 $Y=1.195 $X2=0 $Y2=0
cc_80 N_A_89_270#_c_78_n N_A3_M1001_g 0.00384761f $X=0.945 $Y=1.195 $X2=0 $Y2=0
cc_81 N_A_89_270#_c_75_n A3 7.01218e-19 $X=0.535 $Y=1.765 $X2=0 $Y2=0
cc_82 N_A_89_270#_c_77_n A3 0.0181696f $X=2.24 $Y=1.195 $X2=0 $Y2=0
cc_83 N_A_89_270#_c_78_n A3 0.0184377f $X=0.945 $Y=1.195 $X2=0 $Y2=0
cc_84 N_A_89_270#_c_77_n N_A2_c_201_n 0.00427213f $X=2.24 $Y=1.195 $X2=-0.19
+ $Y2=-0.245
cc_85 N_A_89_270#_c_77_n N_A2_M1008_g 0.0122853f $X=2.24 $Y=1.195 $X2=0 $Y2=0
cc_86 N_A_89_270#_c_81_n N_A2_M1008_g 0.00218849f $X=2.405 $Y=1.005 $X2=0 $Y2=0
cc_87 N_A_89_270#_c_77_n A2 0.0250329f $X=2.24 $Y=1.195 $X2=0 $Y2=0
cc_88 N_A_89_270#_c_81_n A2 0.00718333f $X=2.405 $Y=1.005 $X2=0 $Y2=0
cc_89 N_A_89_270#_c_77_n N_A1_M1004_g 0.0111197f $X=2.24 $Y=1.195 $X2=0 $Y2=0
cc_90 N_A_89_270#_c_81_n N_A1_M1004_g 0.00877504f $X=2.405 $Y=1.005 $X2=0 $Y2=0
cc_91 N_A_89_270#_c_81_n N_A1_c_233_n 0.00358622f $X=2.405 $Y=1.005 $X2=0 $Y2=0
cc_92 N_A_89_270#_c_81_n N_A1_c_234_n 0.00652803f $X=2.405 $Y=1.005 $X2=0 $Y2=0
cc_93 N_A_89_270#_c_77_n N_A1_c_235_n 3.32499e-19 $X=2.24 $Y=1.195 $X2=0 $Y2=0
cc_94 N_A_89_270#_c_81_n N_A1_c_235_n 2.43363e-19 $X=2.405 $Y=1.005 $X2=0 $Y2=0
cc_95 N_A_89_270#_M1004_d N_A1_c_236_n 6.27105e-19 $X=2.265 $Y=0.615 $X2=0 $Y2=0
cc_96 N_A_89_270#_c_77_n N_A1_c_236_n 0.00623312f $X=2.24 $Y=1.195 $X2=0 $Y2=0
cc_97 N_A_89_270#_c_81_n N_A1_c_236_n 0.00288651f $X=2.405 $Y=1.005 $X2=0 $Y2=0
cc_98 N_A_89_270#_c_77_n N_A1_c_237_n 0.0113079f $X=2.24 $Y=1.195 $X2=0 $Y2=0
cc_99 N_A_89_270#_c_80_n N_B1_M1011_g 4.84241e-19 $X=3.41 $Y=1.105 $X2=0 $Y2=0
cc_100 N_A_89_270#_c_81_n N_B1_M1011_g 0.00848117f $X=2.405 $Y=1.005 $X2=0 $Y2=0
cc_101 N_A_89_270#_c_79_n N_B1_c_285_n 0.0107926f $X=3.245 $Y=1.53 $X2=0 $Y2=0
cc_102 N_A_89_270#_c_81_n N_B1_c_285_n 0.00197044f $X=2.405 $Y=1.005 $X2=0 $Y2=0
cc_103 N_A_89_270#_c_87_n N_B1_c_290_n 0.0029031f $X=3.27 $Y=2.105 $X2=0 $Y2=0
cc_104 N_A_89_270#_c_79_n N_B1_c_286_n 0.00839397f $X=3.245 $Y=1.53 $X2=0 $Y2=0
cc_105 N_A_89_270#_c_80_n N_B1_c_286_n 2.58467e-19 $X=3.41 $Y=1.105 $X2=0 $Y2=0
cc_106 N_A_89_270#_c_81_n N_B1_c_286_n 0.00446272f $X=2.405 $Y=1.005 $X2=0 $Y2=0
cc_107 N_A_89_270#_c_81_n B1 0.00186884f $X=2.405 $Y=1.005 $X2=0 $Y2=0
cc_108 N_A_89_270#_c_79_n N_C1_c_328_n 0.0134659f $X=3.245 $Y=1.53 $X2=0 $Y2=0
cc_109 N_A_89_270#_c_82_n N_C1_c_328_n 0.0108566f $X=3.34 $Y=1.94 $X2=0 $Y2=0
cc_110 N_A_89_270#_c_86_n N_C1_c_335_n 0.0136119f $X=3.27 $Y=2.815 $X2=0 $Y2=0
cc_111 N_A_89_270#_c_87_n N_C1_c_335_n 0.00503781f $X=3.27 $Y=2.105 $X2=0 $Y2=0
cc_112 N_A_89_270#_c_82_n N_C1_c_335_n 0.00210336f $X=3.34 $Y=1.94 $X2=0 $Y2=0
cc_113 N_A_89_270#_c_80_n N_C1_M1000_g 0.00737166f $X=3.41 $Y=1.105 $X2=0 $Y2=0
cc_114 N_A_89_270#_c_81_n N_C1_M1000_g 5.26759e-19 $X=2.405 $Y=1.005 $X2=0 $Y2=0
cc_115 N_A_89_270#_c_79_n N_C1_c_330_n 0.00906085f $X=3.245 $Y=1.53 $X2=0 $Y2=0
cc_116 N_A_89_270#_c_80_n N_C1_c_330_n 0.00493627f $X=3.41 $Y=1.105 $X2=0 $Y2=0
cc_117 N_A_89_270#_c_81_n N_C1_c_330_n 4.1554e-19 $X=2.405 $Y=1.005 $X2=0 $Y2=0
cc_118 N_A_89_270#_c_87_n N_C1_c_330_n 6.35295e-19 $X=3.27 $Y=2.105 $X2=0 $Y2=0
cc_119 N_A_89_270#_c_83_n N_C1_c_330_n 0.00141795f $X=3.41 $Y=1.53 $X2=0 $Y2=0
cc_120 N_A_89_270#_c_80_n N_C1_c_332_n 0.00363944f $X=3.41 $Y=1.105 $X2=0 $Y2=0
cc_121 N_A_89_270#_M1000_d N_C1_c_333_n 0.00273424f $X=3.27 $Y=0.615 $X2=0 $Y2=0
cc_122 N_A_89_270#_c_80_n N_C1_c_333_n 0.00981852f $X=3.41 $Y=1.105 $X2=0 $Y2=0
cc_123 N_A_89_270#_c_75_n N_X_c_371_n 0.0019783f $X=0.535 $Y=1.765 $X2=0 $Y2=0
cc_124 N_A_89_270#_c_78_n N_X_c_371_n 0.00920337f $X=0.945 $Y=1.195 $X2=0 $Y2=0
cc_125 N_A_89_270#_c_76_n N_X_c_372_n 4.43891e-19 $X=0.735 $Y=1.35 $X2=0 $Y2=0
cc_126 N_A_89_270#_c_75_n X 0.00320178f $X=0.535 $Y=1.765 $X2=0 $Y2=0
cc_127 N_A_89_270#_c_75_n X 0.0102397f $X=0.535 $Y=1.765 $X2=0 $Y2=0
cc_128 N_A_89_270#_c_75_n N_X_c_373_n 0.0135477f $X=0.535 $Y=1.765 $X2=0 $Y2=0
cc_129 N_A_89_270#_c_76_n N_X_c_373_n 0.00256161f $X=0.735 $Y=1.35 $X2=0 $Y2=0
cc_130 N_A_89_270#_c_78_n N_X_c_373_n 0.0299346f $X=0.945 $Y=1.195 $X2=0 $Y2=0
cc_131 N_A_89_270#_c_75_n N_VPWR_c_393_n 0.0124634f $X=0.535 $Y=1.765 $X2=0
+ $Y2=0
cc_132 N_A_89_270#_c_77_n N_VPWR_c_393_n 0.00508495f $X=2.24 $Y=1.195 $X2=0
+ $Y2=0
cc_133 N_A_89_270#_c_78_n N_VPWR_c_393_n 0.0178289f $X=0.945 $Y=1.195 $X2=0
+ $Y2=0
cc_134 N_A_89_270#_c_86_n N_VPWR_c_397_n 0.0208407f $X=3.27 $Y=2.815 $X2=0 $Y2=0
cc_135 N_A_89_270#_c_75_n N_VPWR_c_392_n 0.00862284f $X=0.535 $Y=1.765 $X2=0
+ $Y2=0
cc_136 N_A_89_270#_c_86_n N_VPWR_c_392_n 0.0172173f $X=3.27 $Y=2.815 $X2=0 $Y2=0
cc_137 N_A_89_270#_c_75_n N_VPWR_c_399_n 0.00445602f $X=0.535 $Y=1.765 $X2=0
+ $Y2=0
cc_138 N_A_89_270#_c_77_n N_A_258_392#_c_433_n 0.00649318f $X=2.24 $Y=1.195
+ $X2=0 $Y2=0
cc_139 N_A_89_270#_c_77_n N_A_258_392#_c_435_n 0.00880952f $X=2.24 $Y=1.195
+ $X2=0 $Y2=0
cc_140 N_A_89_270#_c_81_n N_A_258_392#_c_435_n 0.00103949f $X=2.405 $Y=1.005
+ $X2=0 $Y2=0
cc_141 N_A_89_270#_c_79_n N_A_258_392#_c_436_n 0.00117705f $X=3.245 $Y=1.53
+ $X2=0 $Y2=0
cc_142 N_A_89_270#_c_81_n N_A_258_392#_c_436_n 0.0178798f $X=2.405 $Y=1.005
+ $X2=0 $Y2=0
cc_143 N_A_89_270#_c_87_n N_A_258_392#_c_436_n 0.00597484f $X=3.27 $Y=2.105
+ $X2=0 $Y2=0
cc_144 N_A_89_270#_c_87_n N_A_258_392#_c_437_n 0.0270074f $X=3.27 $Y=2.105 $X2=0
+ $Y2=0
cc_145 N_A_89_270#_c_77_n N_VGND_M1003_d 0.00177524f $X=2.24 $Y=1.195 $X2=-0.19
+ $Y2=-0.245
cc_146 N_A_89_270#_c_78_n N_VGND_M1003_d 8.58534e-19 $X=0.945 $Y=1.195 $X2=-0.19
+ $Y2=-0.245
cc_147 N_A_89_270#_c_76_n N_VGND_c_472_n 0.0140304f $X=0.735 $Y=1.35 $X2=0 $Y2=0
cc_148 N_A_89_270#_c_77_n N_VGND_c_472_n 0.0136318f $X=2.24 $Y=1.195 $X2=0 $Y2=0
cc_149 N_A_89_270#_c_78_n N_VGND_c_472_n 0.00890417f $X=0.945 $Y=1.195 $X2=0
+ $Y2=0
cc_150 N_A_89_270#_c_79_n N_VGND_c_473_n 0.0212375f $X=3.245 $Y=1.53 $X2=0 $Y2=0
cc_151 N_A_89_270#_c_81_n N_VGND_c_473_n 6.88425e-19 $X=2.405 $Y=1.005 $X2=0
+ $Y2=0
cc_152 N_A_89_270#_c_76_n N_VGND_c_474_n 0.00405273f $X=0.735 $Y=1.35 $X2=0
+ $Y2=0
cc_153 N_A_89_270#_c_76_n N_VGND_c_478_n 0.00424518f $X=0.735 $Y=1.35 $X2=0
+ $Y2=0
cc_154 N_A_89_270#_c_81_n N_VGND_c_478_n 0.00775516f $X=2.405 $Y=1.005 $X2=0
+ $Y2=0
cc_155 N_A_89_270#_c_77_n A_264_120# 0.00756132f $X=2.24 $Y=1.195 $X2=-0.19
+ $Y2=-0.245
cc_156 N_A_89_270#_c_77_n A_359_123# 0.00335572f $X=2.24 $Y=1.195 $X2=-0.19
+ $Y2=-0.245
cc_157 N_A3_c_171_n N_A2_c_201_n 0.0349921f $X=1.215 $Y=1.885 $X2=-0.19
+ $Y2=-0.245
cc_158 A3 N_A2_c_201_n 4.06578e-19 $X=1.115 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_159 N_A3_M1001_g N_A2_M1008_g 0.0378038f $X=1.245 $Y=0.92 $X2=0 $Y2=0
cc_160 N_A3_c_171_n A2 0.00187659f $X=1.215 $Y=1.885 $X2=0 $Y2=0
cc_161 A3 A2 0.0226838f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_162 N_A3_M1001_g N_A1_c_237_n 0.00181953f $X=1.245 $Y=0.92 $X2=0 $Y2=0
cc_163 N_A3_c_171_n X 5.80701e-19 $X=1.215 $Y=1.885 $X2=0 $Y2=0
cc_164 N_A3_c_171_n N_VPWR_c_393_n 0.0134421f $X=1.215 $Y=1.885 $X2=0 $Y2=0
cc_165 N_A3_c_171_n N_VPWR_c_395_n 0.00445602f $X=1.215 $Y=1.885 $X2=0 $Y2=0
cc_166 N_A3_c_171_n N_VPWR_c_392_n 0.00858778f $X=1.215 $Y=1.885 $X2=0 $Y2=0
cc_167 N_A3_c_171_n N_A_258_392#_c_433_n 0.00292136f $X=1.215 $Y=1.885 $X2=0
+ $Y2=0
cc_168 A3 N_A_258_392#_c_433_n 0.00747456f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_169 N_A3_c_171_n N_A_258_392#_c_434_n 0.00874253f $X=1.215 $Y=1.885 $X2=0
+ $Y2=0
cc_170 N_A3_M1001_g N_VGND_c_472_n 0.00343181f $X=1.245 $Y=0.92 $X2=0 $Y2=0
cc_171 N_A3_M1001_g N_VGND_c_476_n 0.00428744f $X=1.245 $Y=0.92 $X2=0 $Y2=0
cc_172 N_A3_M1001_g N_VGND_c_478_n 0.00476395f $X=1.245 $Y=0.92 $X2=0 $Y2=0
cc_173 N_A2_M1008_g N_A1_M1004_g 0.0378467f $X=1.72 $Y=0.935 $X2=0 $Y2=0
cc_174 N_A2_c_201_n N_A1_c_234_n 0.0242473f $X=1.665 $Y=1.885 $X2=0 $Y2=0
cc_175 A2 N_A1_c_234_n 0.00167797f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_176 N_A2_c_201_n N_A1_c_239_n 0.021479f $X=1.665 $Y=1.885 $X2=0 $Y2=0
cc_177 N_A2_M1008_g N_A1_c_235_n 0.00129249f $X=1.72 $Y=0.935 $X2=0 $Y2=0
cc_178 N_A2_M1008_g N_A1_c_237_n 0.0113054f $X=1.72 $Y=0.935 $X2=0 $Y2=0
cc_179 N_A2_c_201_n N_VPWR_c_394_n 0.00556651f $X=1.665 $Y=1.885 $X2=0 $Y2=0
cc_180 N_A2_c_201_n N_VPWR_c_395_n 0.00445602f $X=1.665 $Y=1.885 $X2=0 $Y2=0
cc_181 N_A2_c_201_n N_VPWR_c_392_n 0.00858505f $X=1.665 $Y=1.885 $X2=0 $Y2=0
cc_182 N_A2_c_201_n N_A_258_392#_c_433_n 9.73076e-19 $X=1.665 $Y=1.885 $X2=0
+ $Y2=0
cc_183 A2 N_A_258_392#_c_433_n 0.00334681f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_184 N_A2_c_201_n N_A_258_392#_c_434_n 0.0107586f $X=1.665 $Y=1.885 $X2=0
+ $Y2=0
cc_185 N_A2_c_201_n N_A_258_392#_c_435_n 0.0163754f $X=1.665 $Y=1.885 $X2=0
+ $Y2=0
cc_186 A2 N_A_258_392#_c_435_n 0.0220075f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_187 N_A2_c_201_n N_A_258_392#_c_437_n 5.94528e-19 $X=1.665 $Y=1.885 $X2=0
+ $Y2=0
cc_188 N_A2_M1008_g N_VGND_c_476_n 6.8294e-19 $X=1.72 $Y=0.935 $X2=0 $Y2=0
cc_189 N_A1_M1004_g N_B1_M1011_g 0.0198607f $X=2.19 $Y=0.935 $X2=0 $Y2=0
cc_190 N_A1_c_236_n N_B1_M1011_g 5.66657e-19 $X=2.17 $Y=0.34 $X2=0 $Y2=0
cc_191 N_A1_c_234_n N_B1_c_285_n 0.0101876f $X=2.205 $Y=1.795 $X2=0 $Y2=0
cc_192 N_A1_c_239_n N_B1_c_290_n 0.0191663f $X=2.205 $Y=1.885 $X2=0 $Y2=0
cc_193 N_A1_c_233_n N_B1_c_286_n 0.00777372f $X=2.205 $Y=1.42 $X2=0 $Y2=0
cc_194 N_A1_M1004_g B1 3.45758e-19 $X=2.19 $Y=0.935 $X2=0 $Y2=0
cc_195 N_A1_c_235_n B1 0.00143004f $X=2.17 $Y=0.34 $X2=0 $Y2=0
cc_196 N_A1_c_236_n B1 0.0285655f $X=2.17 $Y=0.34 $X2=0 $Y2=0
cc_197 N_A1_c_235_n N_B1_c_288_n 0.0213815f $X=2.17 $Y=0.34 $X2=0 $Y2=0
cc_198 N_A1_c_236_n N_B1_c_288_n 3.01834e-19 $X=2.17 $Y=0.34 $X2=0 $Y2=0
cc_199 N_A1_c_239_n N_VPWR_c_394_n 0.0072001f $X=2.205 $Y=1.885 $X2=0 $Y2=0
cc_200 N_A1_c_239_n N_VPWR_c_397_n 0.00445602f $X=2.205 $Y=1.885 $X2=0 $Y2=0
cc_201 N_A1_c_239_n N_VPWR_c_392_n 0.00857833f $X=2.205 $Y=1.885 $X2=0 $Y2=0
cc_202 N_A1_c_239_n N_A_258_392#_c_434_n 6.89398e-19 $X=2.205 $Y=1.885 $X2=0
+ $Y2=0
cc_203 N_A1_c_239_n N_A_258_392#_c_435_n 0.014741f $X=2.205 $Y=1.885 $X2=0 $Y2=0
cc_204 N_A1_c_239_n N_A_258_392#_c_436_n 0.00145363f $X=2.205 $Y=1.885 $X2=0
+ $Y2=0
cc_205 N_A1_c_239_n N_A_258_392#_c_437_n 0.010265f $X=2.205 $Y=1.885 $X2=0 $Y2=0
cc_206 N_A1_c_237_n N_VGND_c_472_n 0.00827599f $X=2.005 $Y=0.555 $X2=0 $Y2=0
cc_207 N_A1_c_235_n N_VGND_c_476_n 0.0066215f $X=2.17 $Y=0.34 $X2=0 $Y2=0
cc_208 N_A1_c_236_n N_VGND_c_476_n 0.0215843f $X=2.17 $Y=0.34 $X2=0 $Y2=0
cc_209 N_A1_c_237_n N_VGND_c_476_n 0.0132973f $X=2.005 $Y=0.555 $X2=0 $Y2=0
cc_210 N_A1_c_235_n N_VGND_c_478_n 0.00960263f $X=2.17 $Y=0.34 $X2=0 $Y2=0
cc_211 N_A1_c_236_n N_VGND_c_478_n 0.0110944f $X=2.17 $Y=0.34 $X2=0 $Y2=0
cc_212 N_A1_c_237_n N_VGND_c_478_n 0.0147336f $X=2.005 $Y=0.555 $X2=0 $Y2=0
cc_213 N_A1_c_237_n A_264_120# 0.00131491f $X=2.005 $Y=0.555 $X2=-0.19
+ $Y2=-0.245
cc_214 N_A1_c_236_n A_359_123# 0.00103536f $X=2.17 $Y=0.34 $X2=-0.19 $Y2=-0.245
cc_215 N_A1_c_237_n A_359_123# 0.00273639f $X=2.005 $Y=0.555 $X2=-0.19
+ $Y2=-0.245
cc_216 N_B1_c_285_n N_C1_c_328_n 0.0118625f $X=2.655 $Y=1.795 $X2=0 $Y2=0
cc_217 N_B1_c_290_n N_C1_c_335_n 0.0718606f $X=2.655 $Y=1.885 $X2=0 $Y2=0
cc_218 N_B1_M1011_g N_C1_M1000_g 0.0179711f $X=2.62 $Y=0.935 $X2=0 $Y2=0
cc_219 B1 N_C1_M1000_g 4.01526e-19 $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_220 N_B1_c_286_n N_C1_c_330_n 0.0118625f $X=2.645 $Y=1.48 $X2=0 $Y2=0
cc_221 B1 N_C1_c_331_n 2.72693e-19 $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_222 N_B1_c_288_n N_C1_c_331_n 0.0179383f $X=2.71 $Y=0.34 $X2=0 $Y2=0
cc_223 N_B1_c_290_n N_VPWR_c_397_n 0.00445602f $X=2.655 $Y=1.885 $X2=0 $Y2=0
cc_224 N_B1_c_290_n N_VPWR_c_392_n 0.00857948f $X=2.655 $Y=1.885 $X2=0 $Y2=0
cc_225 N_B1_c_290_n N_A_258_392#_c_436_n 0.00401345f $X=2.655 $Y=1.885 $X2=0
+ $Y2=0
cc_226 N_B1_c_290_n N_A_258_392#_c_437_n 0.0143199f $X=2.655 $Y=1.885 $X2=0
+ $Y2=0
cc_227 N_B1_M1011_g N_VGND_c_473_n 0.00474594f $X=2.62 $Y=0.935 $X2=0 $Y2=0
cc_228 B1 N_VGND_c_473_n 0.0304236f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_229 N_B1_c_288_n N_VGND_c_473_n 0.00291452f $X=2.71 $Y=0.34 $X2=0 $Y2=0
cc_230 B1 N_VGND_c_476_n 0.0227602f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_231 N_B1_c_288_n N_VGND_c_476_n 0.00659434f $X=2.71 $Y=0.34 $X2=0 $Y2=0
cc_232 B1 N_VGND_c_478_n 0.011864f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_233 N_B1_c_288_n N_VGND_c_478_n 0.00886835f $X=2.71 $Y=0.34 $X2=0 $Y2=0
cc_234 N_C1_c_335_n N_VPWR_c_397_n 0.00445602f $X=3.045 $Y=1.885 $X2=0 $Y2=0
cc_235 N_C1_c_335_n N_VPWR_c_392_n 0.00862666f $X=3.045 $Y=1.885 $X2=0 $Y2=0
cc_236 N_C1_c_335_n N_A_258_392#_c_436_n 5.02024e-19 $X=3.045 $Y=1.885 $X2=0
+ $Y2=0
cc_237 N_C1_c_335_n N_A_258_392#_c_437_n 0.00240695f $X=3.045 $Y=1.885 $X2=0
+ $Y2=0
cc_238 N_C1_M1000_g N_VGND_c_473_n 0.0170264f $X=3.195 $Y=0.935 $X2=0 $Y2=0
cc_239 N_C1_c_330_n N_VGND_c_473_n 0.00343901f $X=3.195 $Y=1.405 $X2=0 $Y2=0
cc_240 N_C1_c_331_n N_VGND_c_473_n 0.0116775f $X=3.27 $Y=0.34 $X2=0 $Y2=0
cc_241 N_C1_c_333_n N_VGND_c_473_n 0.030194f $X=3.55 $Y=0.34 $X2=0 $Y2=0
cc_242 N_C1_c_331_n N_VGND_c_477_n 0.011998f $X=3.27 $Y=0.34 $X2=0 $Y2=0
cc_243 N_C1_c_333_n N_VGND_c_477_n 0.0215843f $X=3.55 $Y=0.34 $X2=0 $Y2=0
cc_244 N_C1_c_331_n N_VGND_c_478_n 0.00332328f $X=3.27 $Y=0.34 $X2=0 $Y2=0
cc_245 N_C1_c_332_n N_VGND_c_478_n 0.0149884f $X=3.55 $Y=0.34 $X2=0 $Y2=0
cc_246 N_C1_c_333_n N_VGND_c_478_n 0.0110944f $X=3.55 $Y=0.34 $X2=0 $Y2=0
cc_247 X N_VPWR_c_393_n 0.039791f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_248 X N_VPWR_c_392_n 0.0127853f $X=0.24 $Y=2.035 $X2=0 $Y2=0
cc_249 X N_VPWR_c_399_n 0.0154862f $X=0.24 $Y=2.035 $X2=0 $Y2=0
cc_250 N_X_c_372_n N_VGND_c_472_n 0.017215f $X=0.52 $Y=0.645 $X2=0 $Y2=0
cc_251 N_X_c_372_n N_VGND_c_474_n 0.00710472f $X=0.52 $Y=0.645 $X2=0 $Y2=0
cc_252 N_X_c_372_n N_VGND_c_478_n 0.00832885f $X=0.52 $Y=0.645 $X2=0 $Y2=0
cc_253 N_VPWR_c_393_n N_A_258_392#_c_433_n 0.00755647f $X=0.875 $Y=2.115 $X2=0
+ $Y2=0
cc_254 N_VPWR_c_393_n N_A_258_392#_c_434_n 0.0330629f $X=0.875 $Y=2.115 $X2=0
+ $Y2=0
cc_255 N_VPWR_c_394_n N_A_258_392#_c_434_n 0.0468234f $X=1.91 $Y=2.455 $X2=0
+ $Y2=0
cc_256 N_VPWR_c_395_n N_A_258_392#_c_434_n 0.014552f $X=1.805 $Y=3.33 $X2=0
+ $Y2=0
cc_257 N_VPWR_c_392_n N_A_258_392#_c_434_n 0.0119791f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_258 N_VPWR_M1002_d N_A_258_392#_c_435_n 0.00344568f $X=1.74 $Y=1.96 $X2=0
+ $Y2=0
cc_259 N_VPWR_c_394_n N_A_258_392#_c_435_n 0.0217227f $X=1.91 $Y=2.455 $X2=0
+ $Y2=0
cc_260 N_VPWR_c_394_n N_A_258_392#_c_437_n 0.0266656f $X=1.91 $Y=2.455 $X2=0
+ $Y2=0
cc_261 N_VPWR_c_397_n N_A_258_392#_c_437_n 0.014552f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_262 N_VPWR_c_392_n N_A_258_392#_c_437_n 0.0119791f $X=3.6 $Y=3.33 $X2=0 $Y2=0
