* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__dfxbp_2 CLK D VGND VNB VPB VPWR Q Q_N
M1000 a_1248_128# a_27_74# a_1000_424# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=3.9205e+11p ps=3.36e+06u
M1001 a_558_445# a_206_368# a_451_503# VPB phighvt w=420000u l=150000u
+  ad=2.394e+11p pd=1.98e+06u as=2.1245e+11p ps=2.19e+06u
M1002 Q a_1290_102# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=2.84038e+12p ps=2.25e+07u
M1003 VGND a_753_284# a_717_102# VNB nshort w=420000u l=150000u
+  ad=2.10485e+12p pd=1.739e+07u as=1.008e+11p ps=1.32e+06u
M1004 Q a_1290_102# VGND VNB nshort w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1005 VPWR a_1290_102# a_1835_368# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.95e+11p ps=2.59e+06u
M1006 Q_N a_1835_368# VGND VNB nshort w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1007 a_753_284# a_558_445# VGND VNB nshort w=550000u l=150000u
+  ad=3.87e+11p pd=2.98e+06u as=0p ps=0u
M1008 VGND a_1835_368# Q_N VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR a_1000_424# a_1290_102# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=2.52e+11p ps=2.28e+06u
M1010 VGND a_1290_102# a_1248_128# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_206_368# a_27_74# VGND VNB nshort w=740000u l=150000u
+  ad=3.252e+11p pd=2.59e+06u as=0p ps=0u
M1012 VPWR a_1835_368# Q_N VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.36e+11p ps=2.84e+06u
M1013 a_1290_102# a_1000_424# VPWR VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_1000_424# a_206_368# a_753_284# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND a_1290_102# Q VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_717_102# a_206_368# a_558_445# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.66075e+11p ps=1.73e+06u
M1017 VGND a_1290_102# a_1835_368# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1018 VPWR a_753_284# a_702_445# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1019 VPWR a_1290_102# a_1208_479# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.785e+11p ps=1.69e+06u
M1020 Q_N a_1835_368# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_753_284# a_558_445# VPWR VPB phighvt w=840000u l=150000u
+  ad=2.52e+11p pd=2.28e+06u as=0p ps=0u
M1022 VPWR CLK a_27_74# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.304e+11p ps=2.83e+06u
M1023 a_206_368# a_27_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=0p ps=0u
M1024 a_702_445# a_27_74# a_558_445# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VGND a_1000_424# a_1290_102# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1026 a_1000_424# a_27_74# a_753_284# VPB phighvt w=840000u l=150000u
+  ad=4.851e+11p pd=3.46e+06u as=0p ps=0u
M1027 a_451_503# D VGND VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1028 a_451_503# D VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VGND CLK a_27_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1030 a_558_445# a_27_74# a_451_503# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VPWR a_1290_102# Q VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_1208_479# a_206_368# a_1000_424# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
