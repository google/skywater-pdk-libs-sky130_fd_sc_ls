* File: sky130_fd_sc_ls__o2bb2ai_1.pex.spice
* Created: Fri Aug 28 13:50:33 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__O2BB2AI_1%A1_N 3 6 7 9 12 14 20
c32 14 0 1.98144e-19 $X=0.24 $Y=1.295
c33 12 0 4.06224e-20 $X=0.58 $Y=1.765
r34 17 20 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=0.27 $Y=1.345
+ $X2=0.495 $Y2=1.345
r35 14 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.345 $X2=0.27 $Y2=1.345
r36 10 12 43.5851 $w=1.5e-07 $l=8.5e-08 $layer=POLY_cond $X=0.495 $Y=1.765
+ $X2=0.58 $Y2=1.765
r37 7 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.58 $Y=1.84 $X2=0.58
+ $Y2=1.765
r38 7 9 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.58 $Y=1.84 $X2=0.58
+ $Y2=2.335
r39 6 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.495 $Y=1.69
+ $X2=0.495 $Y2=1.765
r40 5 20 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.51
+ $X2=0.495 $Y2=1.345
r41 5 6 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=0.495 $Y=1.51
+ $X2=0.495 $Y2=1.69
r42 1 20 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.18
+ $X2=0.495 $Y2=1.345
r43 1 3 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=0.495 $Y=1.18
+ $X2=0.495 $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_LS__O2BB2AI_1%A2_N 1 3 4 5 6 8 9 13
c40 13 0 1.00927e-19 $X=0.945 $Y=1.285
c41 4 0 1.98144e-19 $X=1.03 $Y=1.45
r42 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.945
+ $Y=1.285 $X2=0.945 $Y2=1.285
r43 9 13 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=0.72 $Y=1.285
+ $X2=0.945 $Y2=1.285
r44 6 8 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.03 $Y=1.84 $X2=1.03
+ $Y2=2.335
r45 5 6 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.03 $Y=1.75 $X2=1.03
+ $Y2=1.84
r46 4 12 33.9921 $w=3.34e-07 $l=2.0106e-07 $layer=POLY_cond $X=1.03 $Y=1.45
+ $X2=0.95 $Y2=1.285
r47 4 5 116.613 $w=1.8e-07 $l=3e-07 $layer=POLY_cond $X=1.03 $Y=1.45 $X2=1.03
+ $Y2=1.75
r48 1 12 38.6287 $w=3.34e-07 $l=1.94808e-07 $layer=POLY_cond $X=0.885 $Y=1.12
+ $X2=0.95 $Y2=1.285
r49 1 3 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=0.885 $Y=1.12
+ $X2=0.885 $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_LS__O2BB2AI_1%A_131_383# 1 2 9 11 13 14 15 18 20 21 25
+ 29 31
c72 29 0 4.06224e-20 $X=1.525 $Y=1.515
c73 15 0 1.44605e-19 $X=1.925 $Y=1.557
c74 14 0 1.00927e-19 $X=1.835 $Y=1.515
c75 11 0 5.15112e-20 $X=1.925 $Y=1.765
c76 9 0 5.70837e-20 $X=1.91 $Y=0.74
r77 29 32 5.21343 $w=4.18e-07 $l=1.9e-07 $layer=LI1_cond $X=1.48 $Y=1.515
+ $X2=1.48 $Y2=1.705
r78 29 31 8.7366 $w=4.18e-07 $l=1.65e-07 $layer=LI1_cond $X=1.48 $Y=1.515
+ $X2=1.48 $Y2=1.35
r79 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.525
+ $Y=1.515 $X2=1.525 $Y2=1.515
r80 27 31 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=1.355 $Y=0.95
+ $X2=1.355 $Y2=1.35
r81 25 27 15.9428 $w=5.03e-07 $l=4.35e-07 $layer=LI1_cond $X=1.187 $Y=0.515
+ $X2=1.187 $Y2=0.95
r82 20 32 6.07598 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=1.27 $Y=1.705
+ $X2=1.48 $Y2=1.705
r83 20 21 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.27 $Y=1.705 $X2=0.97
+ $Y2=1.705
r84 16 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.805 $Y=1.79
+ $X2=0.97 $Y2=1.705
r85 16 18 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=0.805 $Y=1.79
+ $X2=0.805 $Y2=2.06
r86 14 30 54.207 $w=3.3e-07 $l=3.1e-07 $layer=POLY_cond $X=1.835 $Y=1.515
+ $X2=1.525 $Y2=1.515
r87 14 15 5.03009 $w=3.3e-07 $l=1.08995e-07 $layer=POLY_cond $X=1.835 $Y=1.515
+ $X2=1.925 $Y2=1.557
r88 11 15 37.0704 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.925 $Y=1.765
+ $X2=1.925 $Y2=1.557
r89 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.925 $Y=1.765
+ $X2=1.925 $Y2=2.4
r90 7 15 37.0704 $w=1.5e-07 $l=2.14369e-07 $layer=POLY_cond $X=1.91 $Y=1.35
+ $X2=1.925 $Y2=1.557
r91 7 9 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.91 $Y=1.35 $X2=1.91
+ $Y2=0.74
r92 2 18 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=0.655
+ $Y=1.915 $X2=0.805 $Y2=2.06
r93 1 25 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.96
+ $Y=0.37 $X2=1.1 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__O2BB2AI_1%B2 1 3 6 8
c35 8 0 1.08595e-19 $X=2.64 $Y=1.665
r36 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.39
+ $Y=1.465 $X2=2.39 $Y2=1.465
r37 8 12 6.22958 $w=4.78e-07 $l=2.5e-07 $layer=LI1_cond $X=2.64 $Y=1.54 $X2=2.39
+ $Y2=1.54
r38 4 11 38.6549 $w=2.86e-07 $l=1.74714e-07 $layer=POLY_cond $X=2.41 $Y=1.3
+ $X2=2.39 $Y2=1.465
r39 4 6 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.41 $Y=1.3 $X2=2.41
+ $Y2=0.74
r40 1 11 61.4066 $w=2.86e-07 $l=3.07409e-07 $layer=POLY_cond $X=2.375 $Y=1.765
+ $X2=2.39 $Y2=1.465
r41 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.375 $Y=1.765
+ $X2=2.375 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__O2BB2AI_1%B1 3 5 7 8 12
r23 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.09
+ $Y=1.465 $X2=3.09 $Y2=1.465
r24 8 12 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=3.09 $Y=1.665 $X2=3.09
+ $Y2=1.465
r25 5 11 55.8528 $w=4e-07 $l=3.69459e-07 $layer=POLY_cond $X=2.855 $Y=1.765
+ $X2=3.01 $Y2=1.465
r26 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.855 $Y=1.765
+ $X2=2.855 $Y2=2.4
r27 1 11 39.5853 $w=4e-07 $l=2.38642e-07 $layer=POLY_cond $X=2.84 $Y=1.3
+ $X2=3.01 $Y2=1.465
r28 1 3 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.84 $Y=1.3 $X2=2.84
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__O2BB2AI_1%VPWR 1 2 3 10 12 14 18 25 27 31 33 42 48
r38 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r39 42 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r40 40 45 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r41 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r42 37 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r43 36 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r44 34 42 11.9488 $w=1.7e-07 $l=2.75e-07 $layer=LI1_cond $X=1.69 $Y=3.33
+ $X2=1.415 $Y2=3.33
r45 34 36 61.9786 $w=1.68e-07 $l=9.5e-07 $layer=LI1_cond $X=1.69 $Y=3.33
+ $X2=2.64 $Y2=3.33
r46 33 47 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=2.995 $Y=3.33
+ $X2=3.177 $Y2=3.33
r47 33 36 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=2.995 $Y=3.33
+ $X2=2.64 $Y2=3.33
r48 31 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r49 31 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r50 31 42 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r51 27 30 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=3.12 $Y=2.115 $X2=3.12
+ $Y2=2.815
r52 25 47 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=3.12 $Y=3.245
+ $X2=3.177 $Y2=3.33
r53 25 30 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=3.12 $Y=3.245
+ $X2=3.12 $Y2=2.815
r54 21 24 8.37255 $w=5.48e-07 $l=3.85e-07 $layer=LI1_cond $X=1.415 $Y=2.43
+ $X2=1.415 $Y2=2.815
r55 18 21 8.04635 $w=5.48e-07 $l=3.7e-07 $layer=LI1_cond $X=1.415 $Y=2.06
+ $X2=1.415 $Y2=2.43
r56 16 42 2.31338 $w=5.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.415 $Y=3.245
+ $X2=1.415 $Y2=3.33
r57 16 24 9.35116 $w=5.48e-07 $l=4.3e-07 $layer=LI1_cond $X=1.415 $Y=3.245
+ $X2=1.415 $Y2=2.815
r58 15 39 4.67962 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=0.47 $Y=3.33
+ $X2=0.235 $Y2=3.33
r59 14 42 11.9488 $w=1.7e-07 $l=2.75e-07 $layer=LI1_cond $X=1.14 $Y=3.33
+ $X2=1.415 $Y2=3.33
r60 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.14 $Y=3.33
+ $X2=0.47 $Y2=3.33
r61 10 39 3.08656 $w=3.3e-07 $l=1.14782e-07 $layer=LI1_cond $X=0.305 $Y=3.245
+ $X2=0.235 $Y2=3.33
r62 10 12 41.3832 $w=3.28e-07 $l=1.185e-06 $layer=LI1_cond $X=0.305 $Y=3.245
+ $X2=0.305 $Y2=2.06
r63 3 30 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.93
+ $Y=1.84 $X2=3.08 $Y2=2.815
r64 3 27 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=2.93
+ $Y=1.84 $X2=3.08 $Y2=2.115
r65 2 24 600 $w=5.2e-07 $l=1.1225e-06 $layer=licon1_PDIFF $count=1 $X=1.105
+ $Y=1.915 $X2=1.605 $Y2=2.815
r66 2 21 600 $w=5.2e-07 $l=7.22997e-07 $layer=licon1_PDIFF $count=1 $X=1.105
+ $Y=1.915 $X2=1.605 $Y2=2.43
r67 2 21 600 $w=5.2e-07 $l=5.85214e-07 $layer=licon1_PDIFF $count=1 $X=1.105
+ $Y=1.915 $X2=1.255 $Y2=2.43
r68 2 18 600 $w=5.2e-07 $l=3.75566e-07 $layer=licon1_PDIFF $count=1 $X=1.105
+ $Y=1.915 $X2=1.415 $Y2=2.06
r69 1 12 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.16
+ $Y=1.915 $X2=0.305 $Y2=2.06
.ends

.subckt PM_SKY130_FD_SC_LS__O2BB2AI_1%Y 1 2 9 15 19 20 21 22
c35 15 0 1.44605e-19 $X=1.945 $Y=1.095
r36 21 22 9.72635 $w=4.53e-07 $l=3.7e-07 $layer=LI1_cond $X=2.087 $Y=2.405
+ $X2=2.087 $Y2=2.775
r37 19 20 9.25191 $w=4.53e-07 $l=1.65e-07 $layer=LI1_cond $X=2.087 $Y=2.115
+ $X2=2.087 $Y2=1.95
r38 17 21 5.99354 $w=4.53e-07 $l=2.28e-07 $layer=LI1_cond $X=2.087 $Y=2.177
+ $X2=2.087 $Y2=2.405
r39 17 19 1.62982 $w=4.53e-07 $l=6.2e-08 $layer=LI1_cond $X=2.087 $Y=2.177
+ $X2=2.087 $Y2=2.115
r40 11 15 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.945 $Y=1.18
+ $X2=1.945 $Y2=1.095
r41 11 20 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.945 $Y=1.18
+ $X2=1.945 $Y2=1.95
r42 7 15 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=1.735 $Y=1.095
+ $X2=1.945 $Y2=1.095
r43 7 9 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=1.735 $Y=1.01
+ $X2=1.735 $Y2=0.515
r44 2 22 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2 $Y=1.84
+ $X2=2.15 $Y2=2.815
r45 2 19 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=2 $Y=1.84
+ $X2=2.15 $Y2=2.115
r46 1 9 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=1.55
+ $Y=0.37 $X2=1.695 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__O2BB2AI_1%VGND 1 2 7 9 13 16 17 18 28 29
r35 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r36 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r37 26 29 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r38 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r39 23 33 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r40 22 25 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.72 $Y=0 $X2=2.16
+ $Y2=0
r41 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r42 20 32 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.222
+ $Y2=0
r43 20 22 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.72
+ $Y2=0
r44 18 26 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r45 18 23 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r46 16 25 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=2.54 $Y=0 $X2=2.16
+ $Y2=0
r47 16 17 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.54 $Y=0 $X2=2.625
+ $Y2=0
r48 15 28 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=2.71 $Y=0 $X2=3.12
+ $Y2=0
r49 15 17 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.71 $Y=0 $X2=2.625
+ $Y2=0
r50 11 17 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.625 $Y=0.085
+ $X2=2.625 $Y2=0
r51 11 13 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=2.625 $Y=0.085
+ $X2=2.625 $Y2=0.57
r52 7 32 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.222 $Y2=0
r53 7 9 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.28 $Y=0.085 $X2=0.28
+ $Y2=0.515
r54 2 13 182 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=1 $X=2.485
+ $Y=0.37 $X2=2.625 $Y2=0.57
r55 1 9 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__O2BB2AI_1%A_397_74# 1 2 7 11 14
r25 14 15 19.8022 $w=2.68e-07 $l=4.35e-07 $layer=LI1_cond $X=2.2 $Y=0.61 $X2=2.2
+ $Y2=1.045
r26 9 11 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=3.055 $Y=0.96
+ $X2=3.055 $Y2=0.515
r27 8 15 3.40055 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=2.37 $Y=1.045 $X2=2.2
+ $Y2=1.045
r28 7 9 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.89 $Y=1.045
+ $X2=3.055 $Y2=0.96
r29 7 8 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.89 $Y=1.045 $X2=2.37
+ $Y2=1.045
r30 2 11 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.915
+ $Y=0.37 $X2=3.055 $Y2=0.515
r31 1 14 182 $w=1.7e-07 $l=3.28634e-07 $layer=licon1_NDIFF $count=1 $X=1.985
+ $Y=0.37 $X2=2.195 $Y2=0.61
.ends

