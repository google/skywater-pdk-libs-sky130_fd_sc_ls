* File: sky130_fd_sc_ls__nand3_1.spice
* Created: Wed Sep  2 11:12:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__nand3_1.pex.spice"
.subckt sky130_fd_sc_ls__nand3_1  VNB VPB C B A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* B	B
* C	C
* VPB	VPB
* VNB	VNB
MM1001 A_155_74# N_C_M1001_g N_VGND_M1001_s VNB NSHORT L=0.15 W=0.74 AD=0.0888
+ AS=0.2109 PD=0.98 PS=2.05 NRD=10.536 NRS=0 M=1 R=4.93333 SA=75000.2 SB=75001.2
+ A=0.111 P=1.78 MULT=1
MM1000 A_233_74# N_B_M1000_g A_155_74# VNB NSHORT L=0.15 W=0.74 AD=0.1554
+ AS=0.0888 PD=1.16 PS=0.98 NRD=25.128 NRS=10.536 M=1 R=4.93333 SA=75000.6
+ SB=75000.8 A=0.111 P=1.78 MULT=1
MM1005 N_Y_M1005_d N_A_M1005_g A_233_74# VNB NSHORT L=0.15 W=0.74 AD=0.2109
+ AS=0.1554 PD=2.05 PS=1.16 NRD=0 NRS=25.128 M=1 R=4.93333 SA=75001.2 SB=75000.2
+ A=0.111 P=1.78 MULT=1
MM1003 N_Y_M1003_d N_C_M1003_g N_VPWR_M1003_s VPB PHIGHVT L=0.15 W=1.12 AD=0.168
+ AS=0.42 PD=1.42 PS=2.99 NRD=1.7533 NRS=15.8191 M=1 R=7.46667 SA=75000.3
+ SB=75001.2 A=0.168 P=2.54 MULT=1
MM1004 N_VPWR_M1004_d N_B_M1004_g N_Y_M1003_d VPB PHIGHVT L=0.15 W=1.12
+ AD=0.2352 AS=0.168 PD=1.54 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75000.8 A=0.168 P=2.54 MULT=1
MM1002 N_Y_M1002_d N_A_M1002_g N_VPWR_M1004_d VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.2352 PD=2.83 PS=1.54 NRD=1.7533 NRS=14.0658 M=1 R=7.46667
+ SA=75001.3 SB=75000.2 A=0.168 P=2.54 MULT=1
DX6_noxref VNB VPB NWDIODE A=5.1708 P=9.28
*
.include "sky130_fd_sc_ls__nand3_1.pxi.spice"
*
.ends
*
*
