* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
M1000 VPWR RESET_B a_30_78# VPB phighvt w=420000u l=150000u
+  ad=1.91035e+12p pd=1.728e+07u as=2.415e+11p ps=2.83e+06u
M1001 a_1468_493# a_490_390# a_1266_74# VPB phighvt w=420000u l=150000u
+  ad=1.134e+11p pd=1.38e+06u as=4.603e+11p ps=3.46e+06u
M1002 VGND a_1864_409# Q VNB nshort w=740000u l=150000u
+  ad=1.38578e+12p pd=1.21e+07u as=2.109e+11p ps=2.05e+06u
M1003 VPWR a_830_359# a_785_457# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1004 VGND RESET_B a_894_138# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1005 a_830_359# a_695_457# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=3.8125e+11p pd=3.01e+06u as=0p ps=0u
M1006 VPWR CLK a_306_96# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=3.1e+11p ps=2.62e+06u
M1007 VPWR a_1864_409# Q VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.808e+11p ps=2.92e+06u
M1008 VGND RESET_B a_117_78# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1009 a_695_457# a_490_390# a_30_78# VPB phighvt w=420000u l=150000u
+  ad=2.499e+11p pd=2.87e+06u as=0p ps=0u
M1010 a_1518_203# RESET_B VPWR VPB phighvt w=420000u l=150000u
+  ad=1.26e+11p pd=1.44e+06u as=0p ps=0u
M1011 a_490_390# a_306_96# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.85e+11p pd=2.57e+06u as=0p ps=0u
M1012 a_894_138# a_830_359# a_816_138# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1013 a_1864_409# a_1266_74# VPWR VPB phighvt w=840000u l=150000u
+  ad=2.478e+11p pd=2.27e+06u as=0p ps=0u
M1014 VGND a_1518_203# a_1476_81# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1015 a_1266_74# a_306_96# a_830_359# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_1476_81# a_306_96# a_1266_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=4.58e+11p ps=3.28e+06u
M1017 a_1518_203# a_1266_74# a_1656_81# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=8.82e+10p ps=1.26e+06u
M1018 a_30_78# D VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_785_457# a_306_96# a_695_457# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_117_78# D a_30_78# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=2.394e+11p ps=2.82e+06u
M1021 VPWR a_1266_74# a_1518_203# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_1266_74# a_490_390# a_830_359# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=4.921e+11p ps=2.81e+06u
M1023 a_1864_409# a_1266_74# VGND VNB nshort w=550000u l=150000u
+  ad=1.5675e+11p pd=1.67e+06u as=0p ps=0u
M1024 VPWR a_1518_203# a_1468_493# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_490_390# a_306_96# VGND VNB nshort w=740000u l=150000u
+  ad=2.183e+11p pd=2.07e+06u as=0p ps=0u
M1026 a_830_359# a_695_457# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_816_138# a_490_390# a_695_457# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.47e+11p ps=1.54e+06u
M1028 a_1656_81# RESET_B VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_695_457# RESET_B VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VGND CLK a_306_96# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.646e+11p ps=2.4e+06u
M1031 a_695_457# a_306_96# a_30_78# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
