* File: sky130_fd_sc_ls__a32oi_4.pxi.spice
* Created: Wed Sep  2 10:53:19 2020
* 
x_PM_SKY130_FD_SC_LS__A32OI_4%B2 N_B2_M1009_g N_B2_c_150_n N_B2_M1000_g
+ N_B2_M1013_g N_B2_c_151_n N_B2_M1021_g N_B2_M1029_g N_B2_c_152_n N_B2_M1024_g
+ N_B2_c_153_n N_B2_M1032_g N_B2_M1033_g B2 B2 B2 B2 N_B2_c_149_n
+ PM_SKY130_FD_SC_LS__A32OI_4%B2
x_PM_SKY130_FD_SC_LS__A32OI_4%B1 N_B1_M1014_g N_B1_c_229_n N_B1_M1010_g
+ N_B1_M1023_g N_B1_c_230_n N_B1_M1015_g N_B1_M1030_g N_B1_c_231_n N_B1_M1025_g
+ N_B1_M1037_g N_B1_c_232_n N_B1_M1034_g B1 B1 B1 B1 B1 N_B1_c_228_n
+ PM_SKY130_FD_SC_LS__A32OI_4%B1
x_PM_SKY130_FD_SC_LS__A32OI_4%A1 N_A1_c_319_n N_A1_M1007_g N_A1_M1005_g
+ N_A1_c_320_n N_A1_M1012_g N_A1_M1022_g N_A1_c_321_n N_A1_M1016_g N_A1_M1031_g
+ N_A1_c_322_n N_A1_M1026_g N_A1_M1038_g A1 A1 A1 N_A1_c_317_n N_A1_c_318_n
+ PM_SKY130_FD_SC_LS__A32OI_4%A1
x_PM_SKY130_FD_SC_LS__A32OI_4%A2 N_A2_M1003_g N_A2_c_400_n N_A2_M1001_g
+ N_A2_M1006_g N_A2_c_401_n N_A2_M1011_g N_A2_M1018_g N_A2_c_402_n N_A2_M1017_g
+ N_A2_M1019_g N_A2_c_403_n N_A2_M1028_g A2 A2 A2 A2 N_A2_c_399_n
+ PM_SKY130_FD_SC_LS__A32OI_4%A2
x_PM_SKY130_FD_SC_LS__A32OI_4%A3 N_A3_c_490_n N_A3_M1002_g N_A3_M1004_g
+ N_A3_c_491_n N_A3_M1008_g N_A3_M1020_g N_A3_c_492_n N_A3_M1027_g N_A3_M1035_g
+ N_A3_c_493_n N_A3_M1036_g N_A3_M1039_g A3 A3 A3 A3 N_A3_c_489_n
+ PM_SKY130_FD_SC_LS__A32OI_4%A3
x_PM_SKY130_FD_SC_LS__A32OI_4%A_27_368# N_A_27_368#_M1000_d N_A_27_368#_M1021_d
+ N_A_27_368#_M1032_d N_A_27_368#_M1015_s N_A_27_368#_M1034_s
+ N_A_27_368#_M1012_s N_A_27_368#_M1026_s N_A_27_368#_M1011_d
+ N_A_27_368#_M1028_d N_A_27_368#_M1008_s N_A_27_368#_M1036_s
+ N_A_27_368#_c_568_n N_A_27_368#_c_569_n N_A_27_368#_c_570_n
+ N_A_27_368#_c_667_p N_A_27_368#_c_571_n N_A_27_368#_c_592_n
+ N_A_27_368#_c_572_n N_A_27_368#_c_596_n N_A_27_368#_c_573_n
+ N_A_27_368#_c_675_p N_A_27_368#_c_603_n N_A_27_368#_c_604_n
+ N_A_27_368#_c_606_n N_A_27_368#_c_614_n N_A_27_368#_c_618_n
+ N_A_27_368#_c_623_n N_A_27_368#_c_574_n N_A_27_368#_c_630_n
+ N_A_27_368#_c_575_n N_A_27_368#_c_635_n N_A_27_368#_c_576_n
+ N_A_27_368#_c_650_n N_A_27_368#_c_577_n N_A_27_368#_c_578_n
+ N_A_27_368#_c_579_n N_A_27_368#_c_580_n N_A_27_368#_c_581_n
+ N_A_27_368#_c_582_n N_A_27_368#_c_583_n N_A_27_368#_c_638_n
+ N_A_27_368#_c_640_n N_A_27_368#_c_659_n PM_SKY130_FD_SC_LS__A32OI_4%A_27_368#
x_PM_SKY130_FD_SC_LS__A32OI_4%Y N_Y_M1014_s N_Y_M1030_s N_Y_M1005_s N_Y_M1031_s
+ N_Y_M1000_s N_Y_M1024_s N_Y_M1010_d N_Y_M1025_d N_Y_c_748_n N_Y_c_752_n
+ N_Y_c_740_n N_Y_c_768_n N_Y_c_772_n N_Y_c_741_n N_Y_c_753_n N_Y_c_757_n
+ N_Y_c_742_n N_Y_c_780_n N_Y_c_743_n N_Y_c_785_n N_Y_c_744_n Y Y Y N_Y_c_745_n
+ N_Y_c_746_n PM_SKY130_FD_SC_LS__A32OI_4%Y
x_PM_SKY130_FD_SC_LS__A32OI_4%VPWR N_VPWR_M1007_d N_VPWR_M1016_d N_VPWR_M1001_s
+ N_VPWR_M1017_s N_VPWR_M1002_d N_VPWR_M1027_d N_VPWR_c_866_n N_VPWR_c_867_n
+ N_VPWR_c_868_n N_VPWR_c_869_n N_VPWR_c_870_n N_VPWR_c_871_n N_VPWR_c_872_n
+ N_VPWR_c_873_n N_VPWR_c_874_n N_VPWR_c_875_n N_VPWR_c_876_n N_VPWR_c_877_n
+ N_VPWR_c_878_n N_VPWR_c_879_n N_VPWR_c_880_n N_VPWR_c_881_n VPWR
+ N_VPWR_c_882_n N_VPWR_c_883_n N_VPWR_c_865_n N_VPWR_c_885_n
+ PM_SKY130_FD_SC_LS__A32OI_4%VPWR
x_PM_SKY130_FD_SC_LS__A32OI_4%A_27_74# N_A_27_74#_M1009_d N_A_27_74#_M1013_d
+ N_A_27_74#_M1033_d N_A_27_74#_M1023_d N_A_27_74#_M1037_d N_A_27_74#_c_996_n
+ N_A_27_74#_c_997_n N_A_27_74#_c_998_n N_A_27_74#_c_999_n N_A_27_74#_c_1000_n
+ N_A_27_74#_c_1001_n N_A_27_74#_c_1002_n N_A_27_74#_c_1003_n
+ N_A_27_74#_c_1004_n N_A_27_74#_c_1005_n N_A_27_74#_c_1006_n
+ PM_SKY130_FD_SC_LS__A32OI_4%A_27_74#
x_PM_SKY130_FD_SC_LS__A32OI_4%VGND N_VGND_M1009_s N_VGND_M1029_s N_VGND_M1004_d
+ N_VGND_M1020_d N_VGND_M1039_d N_VGND_c_1070_n N_VGND_c_1071_n N_VGND_c_1072_n
+ N_VGND_c_1073_n N_VGND_c_1074_n N_VGND_c_1075_n VGND N_VGND_c_1076_n
+ N_VGND_c_1077_n N_VGND_c_1078_n N_VGND_c_1079_n N_VGND_c_1080_n
+ N_VGND_c_1081_n N_VGND_c_1082_n N_VGND_c_1083_n N_VGND_c_1084_n
+ N_VGND_c_1085_n PM_SKY130_FD_SC_LS__A32OI_4%VGND
x_PM_SKY130_FD_SC_LS__A32OI_4%A_868_74# N_A_868_74#_M1005_d N_A_868_74#_M1022_d
+ N_A_868_74#_M1038_d N_A_868_74#_M1006_d N_A_868_74#_M1019_d
+ N_A_868_74#_c_1182_n N_A_868_74#_c_1183_n N_A_868_74#_c_1184_n
+ PM_SKY130_FD_SC_LS__A32OI_4%A_868_74#
x_PM_SKY130_FD_SC_LS__A32OI_4%A_1313_74# N_A_1313_74#_M1003_s
+ N_A_1313_74#_M1018_s N_A_1313_74#_M1004_s N_A_1313_74#_M1035_s
+ N_A_1313_74#_c_1222_n N_A_1313_74#_c_1223_n N_A_1313_74#_c_1224_n
+ N_A_1313_74#_c_1225_n N_A_1313_74#_c_1226_n N_A_1313_74#_c_1227_n
+ N_A_1313_74#_c_1228_n N_A_1313_74#_c_1229_n
+ PM_SKY130_FD_SC_LS__A32OI_4%A_1313_74#
cc_1 VNB N_B2_M1009_g 0.0336211f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_B2_M1013_g 0.0234867f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_3 VNB N_B2_M1029_g 0.0234201f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=0.74
cc_4 VNB N_B2_M1033_g 0.0245585f $X=-0.19 $Y=-0.245 $X2=1.92 $Y2=0.74
cc_5 VNB B2 0.0166475f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_6 VNB N_B2_c_149_n 0.0772304f $X=-0.19 $Y=-0.245 $X2=1.905 $Y2=1.557
cc_7 VNB N_B1_M1014_g 0.022921f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_8 VNB N_B1_M1023_g 0.0232068f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_9 VNB N_B1_M1030_g 0.0231908f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=0.74
cc_10 VNB N_B1_M1037_g 0.030436f $X=-0.19 $Y=-0.245 $X2=1.905 $Y2=2.4
cc_11 VNB B1 0.0107199f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_B1_c_228_n 0.0811167f $X=-0.19 $Y=-0.245 $X2=1.92 $Y2=1.557
cc_13 VNB N_A1_M1005_g 0.0318671f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.4
cc_14 VNB N_A1_M1022_g 0.0242232f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.4
cc_15 VNB N_A1_M1031_g 0.0233769f $X=-0.19 $Y=-0.245 $X2=1.455 $Y2=2.4
cc_16 VNB N_A1_M1038_g 0.0238886f $X=-0.19 $Y=-0.245 $X2=1.92 $Y2=0.74
cc_17 VNB N_A1_c_317_n 0.00260092f $X=-0.19 $Y=-0.245 $X2=1.605 $Y2=1.557
cc_18 VNB N_A1_c_318_n 0.0810377f $X=-0.19 $Y=-0.245 $X2=1.605 $Y2=1.515
cc_19 VNB N_A2_M1003_g 0.0238306f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_20 VNB N_A2_M1006_g 0.0230765f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_21 VNB N_A2_M1018_g 0.0230833f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=0.74
cc_22 VNB N_A2_M1019_g 0.0306791f $X=-0.19 $Y=-0.245 $X2=1.905 $Y2=2.4
cc_23 VNB A2 0.00526789f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_24 VNB N_A2_c_399_n 0.0802905f $X=-0.19 $Y=-0.245 $X2=1.605 $Y2=1.515
cc_25 VNB N_A3_M1004_g 0.0305493f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.4
cc_26 VNB N_A3_M1020_g 0.0224899f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.4
cc_27 VNB N_A3_M1035_g 0.0224899f $X=-0.19 $Y=-0.245 $X2=1.455 $Y2=2.4
cc_28 VNB N_A3_M1039_g 0.031746f $X=-0.19 $Y=-0.245 $X2=1.92 $Y2=0.74
cc_29 VNB A3 0.016914f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_30 VNB N_A3_c_489_n 0.0831316f $X=-0.19 $Y=-0.245 $X2=1.905 $Y2=1.557
cc_31 VNB N_Y_c_740_n 0.00392452f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_Y_c_741_n 0.0109512f $X=-0.19 $Y=-0.245 $X2=1.605 $Y2=1.515
cc_33 VNB N_Y_c_742_n 0.00229834f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.565
cc_34 VNB N_Y_c_743_n 0.00104729f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=1.565
cc_35 VNB N_Y_c_744_n 0.0096783f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_Y_c_745_n 0.0236767f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_Y_c_746_n 0.00229613f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VPWR_c_865_n 0.442315f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_27_74#_c_996_n 0.0277086f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_27_74#_c_997_n 0.00317099f $X=-0.19 $Y=-0.245 $X2=1.455 $Y2=2.4
cc_41 VNB N_A_27_74#_c_998_n 0.0104987f $X=-0.19 $Y=-0.245 $X2=1.455 $Y2=2.4
cc_42 VNB N_A_27_74#_c_999_n 0.00178908f $X=-0.19 $Y=-0.245 $X2=1.905 $Y2=2.4
cc_43 VNB N_A_27_74#_c_1000_n 0.00822418f $X=-0.19 $Y=-0.245 $X2=1.92 $Y2=0.74
cc_44 VNB N_A_27_74#_c_1001_n 0.0029327f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_45 VNB N_A_27_74#_c_1002_n 0.00218829f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_27_74#_c_1003_n 0.00199363f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_27_74#_c_1004_n 0.00127131f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_27_74#_c_1005_n 0.00240889f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.557
cc_49 VNB N_A_27_74#_c_1006_n 0.00747294f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.557
cc_50 VNB N_VGND_c_1070_n 0.00568581f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_1071_n 0.00544084f $X=-0.19 $Y=-0.245 $X2=1.905 $Y2=1.765
cc_52 VNB N_VGND_c_1072_n 0.0115972f $X=-0.19 $Y=-0.245 $X2=1.92 $Y2=0.74
cc_53 VNB N_VGND_c_1073_n 0.00250542f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_54 VNB N_VGND_c_1074_n 0.0120272f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_55 VNB N_VGND_c_1075_n 0.0416027f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_1076_n 0.0191515f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.557
cc_57 VNB N_VGND_c_1077_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.557
cc_58 VNB N_VGND_c_1078_n 0.159911f $X=-0.19 $Y=-0.245 $X2=1.605 $Y2=1.515
cc_59 VNB N_VGND_c_1079_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_1080_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_1081_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_1082_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_1083_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_1084_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_1085_n 0.562946f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_868_74#_c_1182_n 0.00799024f $X=-0.19 $Y=-0.245 $X2=1.905 $Y2=2.4
cc_67 VNB N_A_868_74#_c_1183_n 0.00583627f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_68 VNB N_A_868_74#_c_1184_n 0.0171655f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_69 VNB N_A_1313_74#_c_1222_n 0.0180757f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=1.35
cc_70 VNB N_A_1313_74#_c_1223_n 0.00178908f $X=-0.19 $Y=-0.245 $X2=1.455
+ $Y2=1.765
cc_71 VNB N_A_1313_74#_c_1224_n 0.00527187f $X=-0.19 $Y=-0.245 $X2=1.455 $Y2=2.4
cc_72 VNB N_A_1313_74#_c_1225_n 0.00178908f $X=-0.19 $Y=-0.245 $X2=1.92 $Y2=1.35
cc_73 VNB N_A_1313_74#_c_1226_n 0.00526132f $X=-0.19 $Y=-0.245 $X2=0.635
+ $Y2=1.58
cc_74 VNB N_A_1313_74#_c_1227_n 0.0034448f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_75 VNB N_A_1313_74#_c_1228_n 0.00114016f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_1313_74#_c_1229_n 0.00127131f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VPB N_B2_c_150_n 0.0189957f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.765
cc_78 VPB N_B2_c_151_n 0.0150113f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.765
cc_79 VPB N_B2_c_152_n 0.014664f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=1.765
cc_80 VPB N_B2_c_153_n 0.0152777f $X=-0.19 $Y=1.66 $X2=1.905 $Y2=1.765
cc_81 VPB B2 0.0182603f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.58
cc_82 VPB N_B2_c_149_n 0.049934f $X=-0.19 $Y=1.66 $X2=1.905 $Y2=1.557
cc_83 VPB N_B1_c_229_n 0.0155385f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.765
cc_84 VPB N_B1_c_230_n 0.0154316f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.765
cc_85 VPB N_B1_c_231_n 0.0154273f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=1.765
cc_86 VPB N_B1_c_232_n 0.0163905f $X=-0.19 $Y=1.66 $X2=1.92 $Y2=0.74
cc_87 VPB B1 0.0164154f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_B1_c_228_n 0.0532671f $X=-0.19 $Y=1.66 $X2=1.92 $Y2=1.557
cc_89 VPB N_A1_c_319_n 0.0168644f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.35
cc_90 VPB N_A1_c_320_n 0.0158891f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=1.35
cc_91 VPB N_A1_c_321_n 0.0162341f $X=-0.19 $Y=1.66 $X2=1.425 $Y2=1.35
cc_92 VPB N_A1_c_322_n 0.0166827f $X=-0.19 $Y=1.66 $X2=1.905 $Y2=1.765
cc_93 VPB N_A1_c_317_n 0.010258f $X=-0.19 $Y=1.66 $X2=1.605 $Y2=1.557
cc_94 VPB N_A1_c_318_n 0.0524412f $X=-0.19 $Y=1.66 $X2=1.605 $Y2=1.515
cc_95 VPB N_A2_c_400_n 0.0166169f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.765
cc_96 VPB N_A2_c_401_n 0.0161673f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.765
cc_97 VPB N_A2_c_402_n 0.0158891f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=1.765
cc_98 VPB N_A2_c_403_n 0.0160527f $X=-0.19 $Y=1.66 $X2=1.92 $Y2=0.74
cc_99 VPB A2 0.0136348f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.58
cc_100 VPB N_A2_c_399_n 0.0529013f $X=-0.19 $Y=1.66 $X2=1.605 $Y2=1.515
cc_101 VPB N_A3_c_490_n 0.0165793f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.35
cc_102 VPB N_A3_c_491_n 0.015774f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=1.35
cc_103 VPB N_A3_c_492_n 0.0166601f $X=-0.19 $Y=1.66 $X2=1.425 $Y2=1.35
cc_104 VPB N_A3_c_493_n 0.0216202f $X=-0.19 $Y=1.66 $X2=1.905 $Y2=1.765
cc_105 VPB A3 0.0174223f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.58
cc_106 VPB N_A3_c_489_n 0.0547351f $X=-0.19 $Y=1.66 $X2=1.905 $Y2=1.557
cc_107 VPB N_A_27_368#_c_568_n 0.0366851f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_A_27_368#_c_569_n 0.00291212f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.515
cc_109 VPB N_A_27_368#_c_570_n 0.00988933f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.515
cc_110 VPB N_A_27_368#_c_571_n 0.0028338f $X=-0.19 $Y=1.66 $X2=1.605 $Y2=1.557
cc_111 VPB N_A_27_368#_c_572_n 0.00273412f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_A_27_368#_c_573_n 0.00672073f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_A_27_368#_c_574_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_A_27_368#_c_575_n 0.00289722f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_A_27_368#_c_576_n 0.00289722f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_A_27_368#_c_577_n 0.00739392f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_A_27_368#_c_578_n 0.0353617f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_A_27_368#_c_579_n 0.00123754f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_A_27_368#_c_580_n 0.0022931f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_A_27_368#_c_581_n 0.0022931f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_A_27_368#_c_582_n 0.00257417f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_A_27_368#_c_583_n 0.00265997f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_Y_c_741_n 0.00374514f $X=-0.19 $Y=1.66 $X2=1.605 $Y2=1.515
cc_124 VPB N_VPWR_c_866_n 0.00581944f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=2.4
cc_125 VPB N_VPWR_c_867_n 0.00830446f $X=-0.19 $Y=1.66 $X2=1.92 $Y2=1.35
cc_126 VPB N_VPWR_c_868_n 0.00830302f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_127 VPB N_VPWR_c_869_n 0.00526854f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_870_n 0.00526854f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.557
cc_129 VPB N_VPWR_c_871_n 0.00904197f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.515
cc_130 VPB N_VPWR_c_872_n 0.107585f $X=-0.19 $Y=1.66 $X2=1.425 $Y2=1.557
cc_131 VPB N_VPWR_c_873_n 0.00614127f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=1.557
cc_132 VPB N_VPWR_c_874_n 0.0186948f $X=-0.19 $Y=1.66 $X2=1.605 $Y2=1.515
cc_133 VPB N_VPWR_c_875_n 0.00632158f $X=-0.19 $Y=1.66 $X2=1.605 $Y2=1.515
cc_134 VPB N_VPWR_c_876_n 0.0186748f $X=-0.19 $Y=1.66 $X2=1.92 $Y2=1.557
cc_135 VPB N_VPWR_c_877_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.565
cc_136 VPB N_VPWR_c_878_n 0.0186948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_VPWR_c_879_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.565
cc_138 VPB N_VPWR_c_880_n 0.0185368f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_881_n 0.00614127f $X=-0.19 $Y=1.66 $X2=1.2 $Y2=1.565
cc_140 VPB N_VPWR_c_882_n 0.0185368f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_883_n 0.0194498f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_142 VPB N_VPWR_c_865_n 0.102671f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_143 VPB N_VPWR_c_885_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_144 N_B2_M1033_g N_B1_M1014_g 0.0168335f $X=1.92 $Y=0.74 $X2=0 $Y2=0
cc_145 N_B2_c_153_n N_B1_c_229_n 0.0312239f $X=1.905 $Y=1.765 $X2=0 $Y2=0
cc_146 B2 B1 0.0289875f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_147 N_B2_c_149_n B1 0.00471138f $X=1.905 $Y=1.557 $X2=0 $Y2=0
cc_148 B2 N_B1_c_228_n 2.25699e-19 $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_149 N_B2_c_149_n N_B1_c_228_n 0.0197022f $X=1.905 $Y=1.557 $X2=0 $Y2=0
cc_150 N_B2_c_150_n N_A_27_368#_c_568_n 0.0103707f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_151 N_B2_c_151_n N_A_27_368#_c_568_n 9.23286e-19 $X=1.005 $Y=1.765 $X2=0
+ $Y2=0
cc_152 B2 N_A_27_368#_c_568_n 0.025553f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_153 N_B2_c_150_n N_A_27_368#_c_569_n 0.0114142f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_154 N_B2_c_151_n N_A_27_368#_c_569_n 0.0130825f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_155 N_B2_c_150_n N_A_27_368#_c_570_n 0.00253309f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_156 N_B2_c_152_n N_A_27_368#_c_571_n 0.0128349f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_157 N_B2_c_153_n N_A_27_368#_c_571_n 0.013793f $X=1.905 $Y=1.765 $X2=0 $Y2=0
cc_158 N_B2_c_151_n N_Y_c_748_n 0.0120074f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_159 N_B2_c_152_n N_Y_c_748_n 0.0120074f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_160 B2 N_Y_c_748_n 0.0393875f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_161 N_B2_c_149_n N_Y_c_748_n 0.00130859f $X=1.905 $Y=1.557 $X2=0 $Y2=0
cc_162 N_B2_c_153_n N_Y_c_752_n 0.0163125f $X=1.905 $Y=1.765 $X2=0 $Y2=0
cc_163 N_B2_c_151_n N_Y_c_753_n 0.00887901f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_164 N_B2_c_152_n N_Y_c_753_n 5.7112e-19 $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_165 B2 N_Y_c_753_n 0.0252536f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_166 N_B2_c_149_n N_Y_c_753_n 0.00166699f $X=1.905 $Y=1.557 $X2=0 $Y2=0
cc_167 N_B2_c_151_n N_Y_c_757_n 5.7112e-19 $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_168 N_B2_c_152_n N_Y_c_757_n 0.00891808f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_169 N_B2_c_153_n N_Y_c_757_n 0.00946786f $X=1.905 $Y=1.765 $X2=0 $Y2=0
cc_170 B2 N_Y_c_757_n 0.0210582f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_171 N_B2_c_149_n N_Y_c_757_n 0.00137451f $X=1.905 $Y=1.557 $X2=0 $Y2=0
cc_172 N_B2_c_150_n N_VPWR_c_872_n 0.00278262f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_173 N_B2_c_151_n N_VPWR_c_872_n 0.00278271f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_174 N_B2_c_152_n N_VPWR_c_872_n 0.00278271f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_175 N_B2_c_153_n N_VPWR_c_872_n 0.00278271f $X=1.905 $Y=1.765 $X2=0 $Y2=0
cc_176 N_B2_c_150_n N_VPWR_c_865_n 0.0035775f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_177 N_B2_c_151_n N_VPWR_c_865_n 0.0035424f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_178 N_B2_c_152_n N_VPWR_c_865_n 0.00353823f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_179 N_B2_c_153_n N_VPWR_c_865_n 0.00354337f $X=1.905 $Y=1.765 $X2=0 $Y2=0
cc_180 N_B2_M1009_g N_A_27_74#_c_996_n 0.0101077f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_181 N_B2_M1013_g N_A_27_74#_c_996_n 9.62944e-19 $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_182 N_B2_M1009_g N_A_27_74#_c_997_n 0.0115433f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_183 N_B2_M1013_g N_A_27_74#_c_997_n 0.0134851f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_184 B2 N_A_27_74#_c_997_n 0.0510636f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_185 N_B2_c_149_n N_A_27_74#_c_997_n 0.00381149f $X=1.905 $Y=1.557 $X2=0 $Y2=0
cc_186 N_B2_M1009_g N_A_27_74#_c_998_n 0.00214722f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_187 B2 N_A_27_74#_c_998_n 0.0286342f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_188 N_B2_M1013_g N_A_27_74#_c_999_n 3.92313e-19 $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_189 N_B2_M1029_g N_A_27_74#_c_999_n 3.92313e-19 $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_190 N_B2_M1029_g N_A_27_74#_c_1000_n 0.0134594f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_191 N_B2_M1033_g N_A_27_74#_c_1000_n 0.0185515f $X=1.92 $Y=0.74 $X2=0 $Y2=0
cc_192 B2 N_A_27_74#_c_1000_n 0.0377574f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_193 N_B2_c_149_n N_A_27_74#_c_1000_n 0.00369939f $X=1.905 $Y=1.557 $X2=0
+ $Y2=0
cc_194 N_B2_M1033_g N_A_27_74#_c_1002_n 0.00109794f $X=1.92 $Y=0.74 $X2=0 $Y2=0
cc_195 B2 N_A_27_74#_c_1004_n 0.0146029f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_196 N_B2_c_149_n N_A_27_74#_c_1004_n 0.00232957f $X=1.905 $Y=1.557 $X2=0
+ $Y2=0
cc_197 N_B2_M1009_g N_VGND_c_1070_n 0.00571035f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_198 N_B2_M1013_g N_VGND_c_1070_n 0.0103415f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_199 N_B2_M1029_g N_VGND_c_1070_n 4.71636e-19 $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_200 N_B2_M1013_g N_VGND_c_1071_n 4.71636e-19 $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_201 N_B2_M1029_g N_VGND_c_1071_n 0.01032f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_202 N_B2_M1033_g N_VGND_c_1071_n 0.00397166f $X=1.92 $Y=0.74 $X2=0 $Y2=0
cc_203 N_B2_M1009_g N_VGND_c_1076_n 0.00434272f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_204 N_B2_M1013_g N_VGND_c_1077_n 0.00383152f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_205 N_B2_M1029_g N_VGND_c_1077_n 0.00383152f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_206 N_B2_M1033_g N_VGND_c_1078_n 0.00461464f $X=1.92 $Y=0.74 $X2=0 $Y2=0
cc_207 N_B2_M1009_g N_VGND_c_1085_n 0.00824376f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_208 N_B2_M1013_g N_VGND_c_1085_n 0.0075754f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_209 N_B2_M1029_g N_VGND_c_1085_n 0.0075754f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_210 N_B2_M1033_g N_VGND_c_1085_n 0.00908708f $X=1.92 $Y=0.74 $X2=0 $Y2=0
cc_211 N_B1_c_232_n N_A1_c_319_n 0.02625f $X=3.905 $Y=1.765 $X2=-0.19 $Y2=-0.245
cc_212 B1 N_A1_c_317_n 0.0305566f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_213 N_B1_c_228_n N_A1_c_317_n 0.00132015f $X=3.8 $Y=1.515 $X2=0 $Y2=0
cc_214 B1 N_A1_c_318_n 0.00193892f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_215 N_B1_c_228_n N_A1_c_318_n 0.00934408f $X=3.8 $Y=1.515 $X2=0 $Y2=0
cc_216 N_B1_c_229_n N_A_27_368#_c_592_n 0.00769091f $X=2.405 $Y=1.765 $X2=0
+ $Y2=0
cc_217 N_B1_c_230_n N_A_27_368#_c_592_n 5.85804e-19 $X=2.905 $Y=1.765 $X2=0
+ $Y2=0
cc_218 N_B1_c_229_n N_A_27_368#_c_572_n 0.0111147f $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_219 N_B1_c_230_n N_A_27_368#_c_572_n 0.014127f $X=2.905 $Y=1.765 $X2=0 $Y2=0
cc_220 N_B1_c_231_n N_A_27_368#_c_596_n 0.00769091f $X=3.405 $Y=1.765 $X2=0
+ $Y2=0
cc_221 N_B1_c_232_n N_A_27_368#_c_596_n 5.85804e-19 $X=3.905 $Y=1.765 $X2=0
+ $Y2=0
cc_222 N_B1_c_231_n N_A_27_368#_c_573_n 0.0111147f $X=3.405 $Y=1.765 $X2=0 $Y2=0
cc_223 N_B1_c_232_n N_A_27_368#_c_573_n 0.0143028f $X=3.905 $Y=1.765 $X2=0 $Y2=0
cc_224 N_B1_c_229_n N_A_27_368#_c_580_n 0.00189622f $X=2.405 $Y=1.765 $X2=0
+ $Y2=0
cc_225 N_B1_c_231_n N_A_27_368#_c_581_n 0.00193739f $X=3.405 $Y=1.765 $X2=0
+ $Y2=0
cc_226 N_B1_c_229_n N_Y_c_752_n 0.0153714f $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_227 B1 N_Y_c_752_n 0.0330918f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_228 N_B1_M1023_g N_Y_c_740_n 0.014265f $X=2.78 $Y=0.74 $X2=0 $Y2=0
cc_229 N_B1_M1030_g N_Y_c_740_n 0.0146892f $X=3.28 $Y=0.74 $X2=0 $Y2=0
cc_230 B1 N_Y_c_740_n 0.115026f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_231 N_B1_c_228_n N_Y_c_740_n 0.00644215f $X=3.8 $Y=1.515 $X2=0 $Y2=0
cc_232 N_B1_c_230_n N_Y_c_768_n 0.0122806f $X=2.905 $Y=1.765 $X2=0 $Y2=0
cc_233 N_B1_c_231_n N_Y_c_768_n 0.0154321f $X=3.405 $Y=1.765 $X2=0 $Y2=0
cc_234 B1 N_Y_c_768_n 0.046015f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_235 N_B1_c_228_n N_Y_c_768_n 0.00157913f $X=3.8 $Y=1.515 $X2=0 $Y2=0
cc_236 N_B1_c_232_n N_Y_c_772_n 0.0127987f $X=3.905 $Y=1.765 $X2=0 $Y2=0
cc_237 B1 N_Y_c_772_n 0.0248711f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_238 N_B1_c_229_n N_Y_c_757_n 4.54023e-19 $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_239 N_B1_M1014_g N_Y_c_742_n 0.00904704f $X=2.35 $Y=0.74 $X2=0 $Y2=0
cc_240 N_B1_M1023_g N_Y_c_742_n 0.00906556f $X=2.78 $Y=0.74 $X2=0 $Y2=0
cc_241 N_B1_M1030_g N_Y_c_742_n 9.11723e-19 $X=3.28 $Y=0.74 $X2=0 $Y2=0
cc_242 B1 N_Y_c_742_n 0.0276216f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_243 N_B1_c_228_n N_Y_c_742_n 0.00231547f $X=3.8 $Y=1.515 $X2=0 $Y2=0
cc_244 N_B1_c_230_n N_Y_c_780_n 0.00891158f $X=2.905 $Y=1.765 $X2=0 $Y2=0
cc_245 N_B1_c_231_n N_Y_c_780_n 4.54023e-19 $X=3.405 $Y=1.765 $X2=0 $Y2=0
cc_246 B1 N_Y_c_780_n 0.025478f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_247 N_B1_c_228_n N_Y_c_780_n 0.00167458f $X=3.8 $Y=1.515 $X2=0 $Y2=0
cc_248 N_B1_M1037_g N_Y_c_743_n 0.00820324f $X=3.71 $Y=0.74 $X2=0 $Y2=0
cc_249 N_B1_c_232_n N_Y_c_785_n 0.00920253f $X=3.905 $Y=1.765 $X2=0 $Y2=0
cc_250 B1 N_Y_c_785_n 0.025478f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_251 N_B1_c_228_n N_Y_c_785_n 0.00167176f $X=3.8 $Y=1.515 $X2=0 $Y2=0
cc_252 N_B1_M1037_g N_Y_c_745_n 0.00954049f $X=3.71 $Y=0.74 $X2=0 $Y2=0
cc_253 N_B1_c_228_n N_Y_c_745_n 0.00533187f $X=3.8 $Y=1.515 $X2=0 $Y2=0
cc_254 N_B1_c_232_n N_VPWR_c_866_n 2.60283e-19 $X=3.905 $Y=1.765 $X2=0 $Y2=0
cc_255 N_B1_c_229_n N_VPWR_c_872_n 0.00278257f $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_256 N_B1_c_230_n N_VPWR_c_872_n 0.00278271f $X=2.905 $Y=1.765 $X2=0 $Y2=0
cc_257 N_B1_c_231_n N_VPWR_c_872_n 0.00278257f $X=3.405 $Y=1.765 $X2=0 $Y2=0
cc_258 N_B1_c_232_n N_VPWR_c_872_n 0.00278271f $X=3.905 $Y=1.765 $X2=0 $Y2=0
cc_259 N_B1_c_229_n N_VPWR_c_865_n 0.00354797f $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_260 N_B1_c_230_n N_VPWR_c_865_n 0.00354745f $X=2.905 $Y=1.765 $X2=0 $Y2=0
cc_261 N_B1_c_231_n N_VPWR_c_865_n 0.00354744f $X=3.405 $Y=1.765 $X2=0 $Y2=0
cc_262 N_B1_c_232_n N_VPWR_c_865_n 0.00355815f $X=3.905 $Y=1.765 $X2=0 $Y2=0
cc_263 N_B1_M1014_g N_A_27_74#_c_1000_n 5.7591e-19 $X=2.35 $Y=0.74 $X2=0 $Y2=0
cc_264 B1 N_A_27_74#_c_1000_n 0.0156959f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_265 N_B1_M1014_g N_A_27_74#_c_1001_n 0.0119575f $X=2.35 $Y=0.74 $X2=0 $Y2=0
cc_266 N_B1_M1023_g N_A_27_74#_c_1001_n 0.00934417f $X=2.78 $Y=0.74 $X2=0 $Y2=0
cc_267 N_B1_M1030_g N_A_27_74#_c_1003_n 0.00805131f $X=3.28 $Y=0.74 $X2=0 $Y2=0
cc_268 N_B1_M1037_g N_A_27_74#_c_1003_n 0.0092831f $X=3.71 $Y=0.74 $X2=0 $Y2=0
cc_269 N_B1_M1023_g N_A_27_74#_c_1005_n 4.46617e-19 $X=2.78 $Y=0.74 $X2=0 $Y2=0
cc_270 N_B1_M1030_g N_A_27_74#_c_1005_n 0.00767662f $X=3.28 $Y=0.74 $X2=0 $Y2=0
cc_271 N_B1_M1037_g N_A_27_74#_c_1005_n 9.18514e-19 $X=3.71 $Y=0.74 $X2=0 $Y2=0
cc_272 N_B1_M1030_g N_A_27_74#_c_1006_n 9.18514e-19 $X=3.28 $Y=0.74 $X2=0 $Y2=0
cc_273 N_B1_M1037_g N_A_27_74#_c_1006_n 0.0087405f $X=3.71 $Y=0.74 $X2=0 $Y2=0
cc_274 N_B1_M1014_g N_VGND_c_1078_n 0.00278271f $X=2.35 $Y=0.74 $X2=0 $Y2=0
cc_275 N_B1_M1023_g N_VGND_c_1078_n 0.00278271f $X=2.78 $Y=0.74 $X2=0 $Y2=0
cc_276 N_B1_M1030_g N_VGND_c_1078_n 0.00279469f $X=3.28 $Y=0.74 $X2=0 $Y2=0
cc_277 N_B1_M1037_g N_VGND_c_1078_n 0.00279469f $X=3.71 $Y=0.74 $X2=0 $Y2=0
cc_278 N_B1_M1014_g N_VGND_c_1085_n 0.00353526f $X=2.35 $Y=0.74 $X2=0 $Y2=0
cc_279 N_B1_M1023_g N_VGND_c_1085_n 0.00354087f $X=2.78 $Y=0.74 $X2=0 $Y2=0
cc_280 N_B1_M1030_g N_VGND_c_1085_n 0.00353176f $X=3.28 $Y=0.74 $X2=0 $Y2=0
cc_281 N_B1_M1037_g N_VGND_c_1085_n 0.00357517f $X=3.71 $Y=0.74 $X2=0 $Y2=0
cc_282 N_B1_M1037_g N_A_868_74#_c_1182_n 0.00378887f $X=3.71 $Y=0.74 $X2=0 $Y2=0
cc_283 N_A1_M1038_g N_A2_M1003_g 0.0246394f $X=6.06 $Y=0.74 $X2=0 $Y2=0
cc_284 N_A1_c_322_n N_A2_c_400_n 0.022874f $X=6.045 $Y=1.765 $X2=0 $Y2=0
cc_285 N_A1_c_318_n N_A2_c_399_n 0.0246394f $X=6.045 $Y=1.557 $X2=0 $Y2=0
cc_286 N_A1_c_319_n N_A_27_368#_c_573_n 0.00183777f $X=4.545 $Y=1.765 $X2=0
+ $Y2=0
cc_287 N_A1_c_319_n N_A_27_368#_c_603_n 0.00733034f $X=4.545 $Y=1.765 $X2=0
+ $Y2=0
cc_288 N_A1_c_319_n N_A_27_368#_c_604_n 0.0155721f $X=4.545 $Y=1.765 $X2=0 $Y2=0
cc_289 N_A1_c_320_n N_A_27_368#_c_604_n 0.0120693f $X=5.045 $Y=1.765 $X2=0 $Y2=0
cc_290 N_A1_c_321_n N_A_27_368#_c_606_n 0.0123082f $X=5.495 $Y=1.765 $X2=0 $Y2=0
cc_291 N_A1_c_322_n N_A_27_368#_c_606_n 0.0123082f $X=6.045 $Y=1.765 $X2=0 $Y2=0
cc_292 N_A1_c_319_n N_A_27_368#_c_582_n 8.30643e-19 $X=4.545 $Y=1.765 $X2=0
+ $Y2=0
cc_293 N_A1_c_320_n N_A_27_368#_c_582_n 0.00726618f $X=5.045 $Y=1.765 $X2=0
+ $Y2=0
cc_294 N_A1_c_321_n N_A_27_368#_c_582_n 0.00746197f $X=5.495 $Y=1.765 $X2=0
+ $Y2=0
cc_295 N_A1_c_322_n N_A_27_368#_c_582_n 5.94284e-19 $X=6.045 $Y=1.765 $X2=0
+ $Y2=0
cc_296 N_A1_c_321_n N_A_27_368#_c_583_n 5.94284e-19 $X=5.495 $Y=1.765 $X2=0
+ $Y2=0
cc_297 N_A1_c_322_n N_A_27_368#_c_583_n 0.00746247f $X=6.045 $Y=1.765 $X2=0
+ $Y2=0
cc_298 N_A1_c_319_n N_Y_c_772_n 0.0117971f $X=4.545 $Y=1.765 $X2=0 $Y2=0
cc_299 N_A1_c_320_n N_Y_c_772_n 0.0110052f $X=5.045 $Y=1.765 $X2=0 $Y2=0
cc_300 N_A1_c_321_n N_Y_c_772_n 0.0112441f $X=5.495 $Y=1.765 $X2=0 $Y2=0
cc_301 N_A1_c_322_n N_Y_c_772_n 0.0153546f $X=6.045 $Y=1.765 $X2=0 $Y2=0
cc_302 N_A1_c_317_n N_Y_c_772_n 0.0940576f $X=5.64 $Y=1.515 $X2=0 $Y2=0
cc_303 N_A1_c_318_n N_Y_c_772_n 0.00861095f $X=6.045 $Y=1.557 $X2=0 $Y2=0
cc_304 N_A1_c_322_n N_Y_c_741_n 0.00423837f $X=6.045 $Y=1.765 $X2=0 $Y2=0
cc_305 N_A1_M1038_g N_Y_c_741_n 0.0100753f $X=6.06 $Y=0.74 $X2=0 $Y2=0
cc_306 N_A1_c_317_n N_Y_c_741_n 0.0192759f $X=5.64 $Y=1.515 $X2=0 $Y2=0
cc_307 N_A1_c_319_n N_Y_c_785_n 8.85902e-19 $X=4.545 $Y=1.765 $X2=0 $Y2=0
cc_308 N_A1_M1022_g N_Y_c_744_n 0.0122111f $X=5.2 $Y=0.74 $X2=0 $Y2=0
cc_309 N_A1_M1031_g N_Y_c_744_n 0.014039f $X=5.63 $Y=0.74 $X2=0 $Y2=0
cc_310 N_A1_M1038_g N_Y_c_744_n 0.0177212f $X=6.06 $Y=0.74 $X2=0 $Y2=0
cc_311 N_A1_c_317_n N_Y_c_744_n 0.0426866f $X=5.64 $Y=1.515 $X2=0 $Y2=0
cc_312 N_A1_c_318_n N_Y_c_744_n 0.00610369f $X=6.045 $Y=1.557 $X2=0 $Y2=0
cc_313 N_A1_M1005_g N_Y_c_745_n 0.0138679f $X=4.7 $Y=0.74 $X2=0 $Y2=0
cc_314 N_A1_c_317_n N_Y_c_745_n 0.0556202f $X=5.64 $Y=1.515 $X2=0 $Y2=0
cc_315 N_A1_c_318_n N_Y_c_745_n 0.00442419f $X=6.045 $Y=1.557 $X2=0 $Y2=0
cc_316 N_A1_M1022_g N_Y_c_746_n 0.0034533f $X=5.2 $Y=0.74 $X2=0 $Y2=0
cc_317 N_A1_M1031_g N_Y_c_746_n 2.36785e-19 $X=5.63 $Y=0.74 $X2=0 $Y2=0
cc_318 N_A1_c_318_n N_Y_c_746_n 0.00416755f $X=6.045 $Y=1.557 $X2=0 $Y2=0
cc_319 N_A1_c_319_n N_VPWR_c_866_n 0.00763441f $X=4.545 $Y=1.765 $X2=0 $Y2=0
cc_320 N_A1_c_320_n N_VPWR_c_866_n 0.00367221f $X=5.045 $Y=1.765 $X2=0 $Y2=0
cc_321 N_A1_c_321_n N_VPWR_c_867_n 0.00396235f $X=5.495 $Y=1.765 $X2=0 $Y2=0
cc_322 N_A1_c_322_n N_VPWR_c_867_n 0.00396235f $X=6.045 $Y=1.765 $X2=0 $Y2=0
cc_323 N_A1_c_319_n N_VPWR_c_872_n 0.00413917f $X=4.545 $Y=1.765 $X2=0 $Y2=0
cc_324 N_A1_c_320_n N_VPWR_c_874_n 0.00445602f $X=5.045 $Y=1.765 $X2=0 $Y2=0
cc_325 N_A1_c_321_n N_VPWR_c_874_n 0.00445602f $X=5.495 $Y=1.765 $X2=0 $Y2=0
cc_326 N_A1_c_322_n N_VPWR_c_876_n 0.00445602f $X=6.045 $Y=1.765 $X2=0 $Y2=0
cc_327 N_A1_c_319_n N_VPWR_c_865_n 0.00819257f $X=4.545 $Y=1.765 $X2=0 $Y2=0
cc_328 N_A1_c_320_n N_VPWR_c_865_n 0.00857378f $X=5.045 $Y=1.765 $X2=0 $Y2=0
cc_329 N_A1_c_321_n N_VPWR_c_865_n 0.00857797f $X=5.495 $Y=1.765 $X2=0 $Y2=0
cc_330 N_A1_c_322_n N_VPWR_c_865_n 0.0085797f $X=6.045 $Y=1.765 $X2=0 $Y2=0
cc_331 N_A1_M1005_g N_A_27_74#_c_1006_n 0.00314096f $X=4.7 $Y=0.74 $X2=0 $Y2=0
cc_332 N_A1_M1005_g N_VGND_c_1078_n 0.00292759f $X=4.7 $Y=0.74 $X2=0 $Y2=0
cc_333 N_A1_M1022_g N_VGND_c_1078_n 0.00291649f $X=5.2 $Y=0.74 $X2=0 $Y2=0
cc_334 N_A1_M1031_g N_VGND_c_1078_n 0.00291649f $X=5.63 $Y=0.74 $X2=0 $Y2=0
cc_335 N_A1_M1038_g N_VGND_c_1078_n 0.00291649f $X=6.06 $Y=0.74 $X2=0 $Y2=0
cc_336 N_A1_M1005_g N_VGND_c_1085_n 0.00363814f $X=4.7 $Y=0.74 $X2=0 $Y2=0
cc_337 N_A1_M1022_g N_VGND_c_1085_n 0.00359779f $X=5.2 $Y=0.74 $X2=0 $Y2=0
cc_338 N_A1_M1031_g N_VGND_c_1085_n 0.00359121f $X=5.63 $Y=0.74 $X2=0 $Y2=0
cc_339 N_A1_M1038_g N_VGND_c_1085_n 0.00359219f $X=6.06 $Y=0.74 $X2=0 $Y2=0
cc_340 N_A1_M1005_g N_A_868_74#_c_1182_n 0.00792667f $X=4.7 $Y=0.74 $X2=0 $Y2=0
cc_341 N_A1_M1022_g N_A_868_74#_c_1182_n 8.9082e-19 $X=5.2 $Y=0.74 $X2=0 $Y2=0
cc_342 N_A1_M1005_g N_A_868_74#_c_1184_n 0.0114225f $X=4.7 $Y=0.74 $X2=0 $Y2=0
cc_343 N_A1_M1022_g N_A_868_74#_c_1184_n 0.0107985f $X=5.2 $Y=0.74 $X2=0 $Y2=0
cc_344 N_A1_M1031_g N_A_868_74#_c_1184_n 0.010218f $X=5.63 $Y=0.74 $X2=0 $Y2=0
cc_345 N_A1_M1038_g N_A_868_74#_c_1184_n 0.010213f $X=6.06 $Y=0.74 $X2=0 $Y2=0
cc_346 N_A1_M1038_g N_A_1313_74#_c_1226_n 2.90368e-19 $X=6.06 $Y=0.74 $X2=0
+ $Y2=0
cc_347 N_A2_c_403_n N_A3_c_490_n 0.0244158f $X=7.995 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_348 A2 N_A3_c_490_n 0.00175333f $X=8.315 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_349 A2 A3 0.0278076f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_350 A2 N_A3_c_489_n 0.0135526f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_351 N_A2_c_399_n N_A3_c_489_n 0.0114182f $X=7.92 $Y=1.515 $X2=0 $Y2=0
cc_352 N_A2_c_400_n N_A_27_368#_c_614_n 0.0173825f $X=6.505 $Y=1.765 $X2=0 $Y2=0
cc_353 N_A2_c_401_n N_A_27_368#_c_614_n 0.013783f $X=7.045 $Y=1.765 $X2=0 $Y2=0
cc_354 A2 N_A_27_368#_c_614_n 0.011627f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_355 N_A2_c_399_n N_A_27_368#_c_614_n 0.0039109f $X=7.92 $Y=1.515 $X2=0 $Y2=0
cc_356 N_A2_c_400_n N_A_27_368#_c_618_n 7.68695e-19 $X=6.505 $Y=1.765 $X2=0
+ $Y2=0
cc_357 N_A2_c_401_n N_A_27_368#_c_618_n 0.00374425f $X=7.045 $Y=1.765 $X2=0
+ $Y2=0
cc_358 N_A2_c_402_n N_A_27_368#_c_618_n 4.27055e-19 $X=7.495 $Y=1.765 $X2=0
+ $Y2=0
cc_359 A2 N_A_27_368#_c_618_n 0.0237598f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_360 N_A2_c_399_n N_A_27_368#_c_618_n 0.00143843f $X=7.92 $Y=1.515 $X2=0 $Y2=0
cc_361 N_A2_c_400_n N_A_27_368#_c_623_n 7.70272e-19 $X=6.505 $Y=1.765 $X2=0
+ $Y2=0
cc_362 N_A2_c_401_n N_A_27_368#_c_623_n 0.0032203f $X=7.045 $Y=1.765 $X2=0 $Y2=0
cc_363 N_A2_c_402_n N_A_27_368#_c_623_n 0.00324175f $X=7.495 $Y=1.765 $X2=0
+ $Y2=0
cc_364 N_A2_c_403_n N_A_27_368#_c_623_n 4.53245e-19 $X=7.995 $Y=1.765 $X2=0
+ $Y2=0
cc_365 N_A2_c_400_n N_A_27_368#_c_574_n 5.48808e-19 $X=6.505 $Y=1.765 $X2=0
+ $Y2=0
cc_366 N_A2_c_401_n N_A_27_368#_c_574_n 0.0070355f $X=7.045 $Y=1.765 $X2=0 $Y2=0
cc_367 N_A2_c_402_n N_A_27_368#_c_574_n 0.00532707f $X=7.495 $Y=1.765 $X2=0
+ $Y2=0
cc_368 N_A2_c_402_n N_A_27_368#_c_630_n 0.0122806f $X=7.495 $Y=1.765 $X2=0 $Y2=0
cc_369 N_A2_c_403_n N_A_27_368#_c_630_n 0.0153714f $X=7.995 $Y=1.765 $X2=0 $Y2=0
cc_370 A2 N_A_27_368#_c_630_n 0.046015f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_371 N_A2_c_399_n N_A_27_368#_c_630_n 0.00157631f $X=7.92 $Y=1.515 $X2=0 $Y2=0
cc_372 N_A2_c_403_n N_A_27_368#_c_575_n 0.00464047f $X=7.995 $Y=1.765 $X2=0
+ $Y2=0
cc_373 A2 N_A_27_368#_c_635_n 0.00580317f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_374 N_A2_c_400_n N_A_27_368#_c_583_n 0.00654007f $X=6.505 $Y=1.765 $X2=0
+ $Y2=0
cc_375 N_A2_c_401_n N_A_27_368#_c_583_n 5.85239e-19 $X=7.045 $Y=1.765 $X2=0
+ $Y2=0
cc_376 N_A2_c_401_n N_A_27_368#_c_638_n 2.24111e-19 $X=7.045 $Y=1.765 $X2=0
+ $Y2=0
cc_377 N_A2_c_402_n N_A_27_368#_c_638_n 0.00162804f $X=7.495 $Y=1.765 $X2=0
+ $Y2=0
cc_378 A2 N_A_27_368#_c_640_n 0.0254782f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_379 N_A2_c_400_n N_Y_c_772_n 0.0052808f $X=6.505 $Y=1.765 $X2=0 $Y2=0
cc_380 N_A2_M1003_g N_Y_c_741_n 0.00901187f $X=6.49 $Y=0.74 $X2=0 $Y2=0
cc_381 N_A2_c_400_n N_Y_c_741_n 0.00413128f $X=6.505 $Y=1.765 $X2=0 $Y2=0
cc_382 A2 N_Y_c_741_n 0.0189003f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_383 N_A2_M1003_g N_Y_c_744_n 0.0030096f $X=6.49 $Y=0.74 $X2=0 $Y2=0
cc_384 N_A2_c_400_n N_VPWR_c_868_n 0.00202193f $X=6.505 $Y=1.765 $X2=0 $Y2=0
cc_385 N_A2_c_401_n N_VPWR_c_868_n 0.00390537f $X=7.045 $Y=1.765 $X2=0 $Y2=0
cc_386 N_A2_c_402_n N_VPWR_c_869_n 0.00548145f $X=7.495 $Y=1.765 $X2=0 $Y2=0
cc_387 N_A2_c_403_n N_VPWR_c_869_n 0.0107303f $X=7.995 $Y=1.765 $X2=0 $Y2=0
cc_388 N_A2_c_400_n N_VPWR_c_876_n 0.00456932f $X=6.505 $Y=1.765 $X2=0 $Y2=0
cc_389 N_A2_c_401_n N_VPWR_c_878_n 0.00445602f $X=7.045 $Y=1.765 $X2=0 $Y2=0
cc_390 N_A2_c_402_n N_VPWR_c_878_n 0.00445602f $X=7.495 $Y=1.765 $X2=0 $Y2=0
cc_391 N_A2_c_403_n N_VPWR_c_880_n 0.00413917f $X=7.995 $Y=1.765 $X2=0 $Y2=0
cc_392 N_A2_c_400_n N_VPWR_c_865_n 0.00890567f $X=6.505 $Y=1.765 $X2=0 $Y2=0
cc_393 N_A2_c_401_n N_VPWR_c_865_n 0.00857717f $X=7.045 $Y=1.765 $X2=0 $Y2=0
cc_394 N_A2_c_402_n N_VPWR_c_865_n 0.00857378f $X=7.495 $Y=1.765 $X2=0 $Y2=0
cc_395 N_A2_c_403_n N_VPWR_c_865_n 0.00818241f $X=7.995 $Y=1.765 $X2=0 $Y2=0
cc_396 N_A2_M1019_g N_VGND_c_1072_n 0.00708914f $X=7.785 $Y=0.74 $X2=0 $Y2=0
cc_397 N_A2_M1003_g N_VGND_c_1078_n 0.00291649f $X=6.49 $Y=0.74 $X2=0 $Y2=0
cc_398 N_A2_M1006_g N_VGND_c_1078_n 0.00291649f $X=6.92 $Y=0.74 $X2=0 $Y2=0
cc_399 N_A2_M1018_g N_VGND_c_1078_n 0.00291649f $X=7.355 $Y=0.74 $X2=0 $Y2=0
cc_400 N_A2_M1019_g N_VGND_c_1078_n 0.00291649f $X=7.785 $Y=0.74 $X2=0 $Y2=0
cc_401 N_A2_M1003_g N_VGND_c_1085_n 0.00359219f $X=6.49 $Y=0.74 $X2=0 $Y2=0
cc_402 N_A2_M1006_g N_VGND_c_1085_n 0.00359171f $X=6.92 $Y=0.74 $X2=0 $Y2=0
cc_403 N_A2_M1018_g N_VGND_c_1085_n 0.00359171f $X=7.355 $Y=0.74 $X2=0 $Y2=0
cc_404 N_A2_M1019_g N_VGND_c_1085_n 0.0036412f $X=7.785 $Y=0.74 $X2=0 $Y2=0
cc_405 N_A2_M1018_g N_A_868_74#_c_1183_n 3.85913e-19 $X=7.355 $Y=0.74 $X2=0
+ $Y2=0
cc_406 N_A2_M1019_g N_A_868_74#_c_1183_n 0.00311138f $X=7.785 $Y=0.74 $X2=0
+ $Y2=0
cc_407 N_A2_M1003_g N_A_868_74#_c_1184_n 0.0142216f $X=6.49 $Y=0.74 $X2=0 $Y2=0
cc_408 N_A2_M1006_g N_A_868_74#_c_1184_n 0.0106163f $X=6.92 $Y=0.74 $X2=0 $Y2=0
cc_409 N_A2_M1018_g N_A_868_74#_c_1184_n 0.010696f $X=7.355 $Y=0.74 $X2=0 $Y2=0
cc_410 N_A2_M1019_g N_A_868_74#_c_1184_n 0.00974906f $X=7.785 $Y=0.74 $X2=0
+ $Y2=0
cc_411 N_A2_M1019_g N_A_1313_74#_c_1222_n 0.0103942f $X=7.785 $Y=0.74 $X2=0
+ $Y2=0
cc_412 N_A2_c_399_n N_A_1313_74#_c_1222_n 0.00566818f $X=7.92 $Y=1.515 $X2=0
+ $Y2=0
cc_413 N_A2_M1003_g N_A_1313_74#_c_1226_n 0.00669488f $X=6.49 $Y=0.74 $X2=0
+ $Y2=0
cc_414 N_A2_M1006_g N_A_1313_74#_c_1226_n 0.0037133f $X=6.92 $Y=0.74 $X2=0 $Y2=0
cc_415 N_A2_M1018_g N_A_1313_74#_c_1226_n 3.85091e-19 $X=7.355 $Y=0.74 $X2=0
+ $Y2=0
cc_416 A2 N_A_1313_74#_c_1226_n 0.140642f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_417 N_A2_c_399_n N_A_1313_74#_c_1226_n 0.00377477f $X=7.92 $Y=1.515 $X2=0
+ $Y2=0
cc_418 N_A2_M1006_g N_A_1313_74#_c_1227_n 0.0116925f $X=6.92 $Y=0.74 $X2=0 $Y2=0
cc_419 N_A2_M1018_g N_A_1313_74#_c_1227_n 0.0140807f $X=7.355 $Y=0.74 $X2=0
+ $Y2=0
cc_420 N_A2_c_399_n N_A_1313_74#_c_1227_n 0.00503527f $X=7.92 $Y=1.515 $X2=0
+ $Y2=0
cc_421 N_A2_M1019_g N_A_1313_74#_c_1228_n 0.00945167f $X=7.785 $Y=0.74 $X2=0
+ $Y2=0
cc_422 N_A3_c_490_n N_A_27_368#_c_575_n 0.0102085f $X=8.495 $Y=1.765 $X2=0 $Y2=0
cc_423 N_A3_c_491_n N_A_27_368#_c_575_n 6.21762e-19 $X=8.995 $Y=1.765 $X2=0
+ $Y2=0
cc_424 N_A3_c_490_n N_A_27_368#_c_635_n 0.0137905f $X=8.495 $Y=1.765 $X2=0 $Y2=0
cc_425 N_A3_c_491_n N_A_27_368#_c_635_n 0.0154321f $X=8.995 $Y=1.765 $X2=0 $Y2=0
cc_426 A3 N_A_27_368#_c_635_n 0.022737f $X=10.235 $Y=1.58 $X2=0 $Y2=0
cc_427 N_A3_c_489_n N_A_27_368#_c_635_n 0.00598447f $X=10.05 $Y=1.557 $X2=0
+ $Y2=0
cc_428 N_A3_c_491_n N_A_27_368#_c_576_n 0.00464047f $X=8.995 $Y=1.765 $X2=0
+ $Y2=0
cc_429 N_A3_c_492_n N_A_27_368#_c_576_n 0.0103256f $X=9.495 $Y=1.765 $X2=0 $Y2=0
cc_430 N_A3_c_493_n N_A_27_368#_c_576_n 6.62391e-19 $X=10.05 $Y=1.765 $X2=0
+ $Y2=0
cc_431 N_A3_c_492_n N_A_27_368#_c_650_n 0.0125417f $X=9.495 $Y=1.765 $X2=0 $Y2=0
cc_432 N_A3_c_493_n N_A_27_368#_c_650_n 0.0125417f $X=10.05 $Y=1.765 $X2=0 $Y2=0
cc_433 A3 N_A_27_368#_c_650_n 0.0477508f $X=10.235 $Y=1.58 $X2=0 $Y2=0
cc_434 N_A3_c_489_n N_A_27_368#_c_650_n 0.00187375f $X=10.05 $Y=1.557 $X2=0
+ $Y2=0
cc_435 N_A3_c_493_n N_A_27_368#_c_577_n 4.27055e-19 $X=10.05 $Y=1.765 $X2=0
+ $Y2=0
cc_436 A3 N_A_27_368#_c_577_n 0.0260502f $X=10.235 $Y=1.58 $X2=0 $Y2=0
cc_437 N_A3_c_492_n N_A_27_368#_c_578_n 6.66225e-19 $X=9.495 $Y=1.765 $X2=0
+ $Y2=0
cc_438 N_A3_c_493_n N_A_27_368#_c_578_n 0.0105634f $X=10.05 $Y=1.765 $X2=0 $Y2=0
cc_439 N_A3_c_490_n N_A_27_368#_c_640_n 4.27055e-19 $X=8.495 $Y=1.765 $X2=0
+ $Y2=0
cc_440 N_A3_c_492_n N_A_27_368#_c_659_n 4.27055e-19 $X=9.495 $Y=1.765 $X2=0
+ $Y2=0
cc_441 A3 N_A_27_368#_c_659_n 0.025478f $X=10.235 $Y=1.58 $X2=0 $Y2=0
cc_442 N_A3_c_489_n N_A_27_368#_c_659_n 0.00166999f $X=10.05 $Y=1.557 $X2=0
+ $Y2=0
cc_443 N_A3_c_490_n N_VPWR_c_869_n 5.07678e-19 $X=8.495 $Y=1.765 $X2=0 $Y2=0
cc_444 N_A3_c_490_n N_VPWR_c_870_n 0.00548145f $X=8.495 $Y=1.765 $X2=0 $Y2=0
cc_445 N_A3_c_491_n N_VPWR_c_870_n 0.0107303f $X=8.995 $Y=1.765 $X2=0 $Y2=0
cc_446 N_A3_c_492_n N_VPWR_c_870_n 5.07678e-19 $X=9.495 $Y=1.765 $X2=0 $Y2=0
cc_447 N_A3_c_492_n N_VPWR_c_871_n 0.00603556f $X=9.495 $Y=1.765 $X2=0 $Y2=0
cc_448 N_A3_c_493_n N_VPWR_c_871_n 0.00736167f $X=10.05 $Y=1.765 $X2=0 $Y2=0
cc_449 N_A3_c_490_n N_VPWR_c_880_n 0.00445602f $X=8.495 $Y=1.765 $X2=0 $Y2=0
cc_450 N_A3_c_491_n N_VPWR_c_882_n 0.00413917f $X=8.995 $Y=1.765 $X2=0 $Y2=0
cc_451 N_A3_c_492_n N_VPWR_c_882_n 0.00445602f $X=9.495 $Y=1.765 $X2=0 $Y2=0
cc_452 N_A3_c_493_n N_VPWR_c_883_n 0.00445602f $X=10.05 $Y=1.765 $X2=0 $Y2=0
cc_453 N_A3_c_490_n N_VPWR_c_865_n 0.00857893f $X=8.495 $Y=1.765 $X2=0 $Y2=0
cc_454 N_A3_c_491_n N_VPWR_c_865_n 0.00818187f $X=8.995 $Y=1.765 $X2=0 $Y2=0
cc_455 N_A3_c_492_n N_VPWR_c_865_n 0.00858298f $X=9.495 $Y=1.765 $X2=0 $Y2=0
cc_456 N_A3_c_493_n N_VPWR_c_865_n 0.0086146f $X=10.05 $Y=1.765 $X2=0 $Y2=0
cc_457 N_A3_M1004_g N_VGND_c_1072_n 0.0120602f $X=8.775 $Y=0.74 $X2=0 $Y2=0
cc_458 N_A3_M1020_g N_VGND_c_1072_n 4.71636e-19 $X=9.205 $Y=0.74 $X2=0 $Y2=0
cc_459 N_A3_M1004_g N_VGND_c_1073_n 4.71636e-19 $X=8.775 $Y=0.74 $X2=0 $Y2=0
cc_460 N_A3_M1020_g N_VGND_c_1073_n 0.0103289f $X=9.205 $Y=0.74 $X2=0 $Y2=0
cc_461 N_A3_M1035_g N_VGND_c_1073_n 0.0103289f $X=9.635 $Y=0.74 $X2=0 $Y2=0
cc_462 N_A3_M1039_g N_VGND_c_1073_n 4.71636e-19 $X=10.065 $Y=0.74 $X2=0 $Y2=0
cc_463 N_A3_M1035_g N_VGND_c_1075_n 5.67074e-19 $X=9.635 $Y=0.74 $X2=0 $Y2=0
cc_464 N_A3_M1039_g N_VGND_c_1075_n 0.015057f $X=10.065 $Y=0.74 $X2=0 $Y2=0
cc_465 A3 N_VGND_c_1075_n 0.023775f $X=10.235 $Y=1.58 $X2=0 $Y2=0
cc_466 N_A3_M1004_g N_VGND_c_1079_n 0.00383152f $X=8.775 $Y=0.74 $X2=0 $Y2=0
cc_467 N_A3_M1020_g N_VGND_c_1079_n 0.00383152f $X=9.205 $Y=0.74 $X2=0 $Y2=0
cc_468 N_A3_M1035_g N_VGND_c_1080_n 0.00383152f $X=9.635 $Y=0.74 $X2=0 $Y2=0
cc_469 N_A3_M1039_g N_VGND_c_1080_n 0.00383152f $X=10.065 $Y=0.74 $X2=0 $Y2=0
cc_470 N_A3_M1004_g N_VGND_c_1085_n 0.0075754f $X=8.775 $Y=0.74 $X2=0 $Y2=0
cc_471 N_A3_M1020_g N_VGND_c_1085_n 0.0075754f $X=9.205 $Y=0.74 $X2=0 $Y2=0
cc_472 N_A3_M1035_g N_VGND_c_1085_n 0.0075754f $X=9.635 $Y=0.74 $X2=0 $Y2=0
cc_473 N_A3_M1039_g N_VGND_c_1085_n 0.0075754f $X=10.065 $Y=0.74 $X2=0 $Y2=0
cc_474 N_A3_M1004_g N_A_868_74#_c_1183_n 7.60322e-19 $X=8.775 $Y=0.74 $X2=0
+ $Y2=0
cc_475 N_A3_M1004_g N_A_1313_74#_c_1222_n 0.0169578f $X=8.775 $Y=0.74 $X2=0
+ $Y2=0
cc_476 A3 N_A_1313_74#_c_1222_n 0.010384f $X=10.235 $Y=1.58 $X2=0 $Y2=0
cc_477 N_A3_c_489_n N_A_1313_74#_c_1222_n 0.00608292f $X=10.05 $Y=1.557 $X2=0
+ $Y2=0
cc_478 N_A3_M1004_g N_A_1313_74#_c_1223_n 3.92313e-19 $X=8.775 $Y=0.74 $X2=0
+ $Y2=0
cc_479 N_A3_M1020_g N_A_1313_74#_c_1223_n 3.92313e-19 $X=9.205 $Y=0.74 $X2=0
+ $Y2=0
cc_480 N_A3_M1020_g N_A_1313_74#_c_1224_n 0.0130453f $X=9.205 $Y=0.74 $X2=0
+ $Y2=0
cc_481 N_A3_M1035_g N_A_1313_74#_c_1224_n 0.0128967f $X=9.635 $Y=0.74 $X2=0
+ $Y2=0
cc_482 N_A3_M1039_g N_A_1313_74#_c_1224_n 0.00174382f $X=10.065 $Y=0.74 $X2=0
+ $Y2=0
cc_483 A3 N_A_1313_74#_c_1224_n 0.0663371f $X=10.235 $Y=1.58 $X2=0 $Y2=0
cc_484 N_A3_c_489_n N_A_1313_74#_c_1224_n 0.0047849f $X=10.05 $Y=1.557 $X2=0
+ $Y2=0
cc_485 N_A3_M1035_g N_A_1313_74#_c_1225_n 3.92313e-19 $X=9.635 $Y=0.74 $X2=0
+ $Y2=0
cc_486 N_A3_M1039_g N_A_1313_74#_c_1225_n 3.92313e-19 $X=10.065 $Y=0.74 $X2=0
+ $Y2=0
cc_487 A3 N_A_1313_74#_c_1229_n 0.0146029f $X=10.235 $Y=1.58 $X2=0 $Y2=0
cc_488 N_A3_c_489_n N_A_1313_74#_c_1229_n 0.00272398f $X=10.05 $Y=1.557 $X2=0
+ $Y2=0
cc_489 N_A_27_368#_c_569_n N_Y_M1000_s 0.00245557f $X=1.145 $Y=2.99 $X2=0 $Y2=0
cc_490 N_A_27_368#_c_571_n N_Y_M1024_s 0.00197722f $X=2.015 $Y=2.99 $X2=0 $Y2=0
cc_491 N_A_27_368#_c_572_n N_Y_M1010_d 0.00250873f $X=3.015 $Y=2.99 $X2=0 $Y2=0
cc_492 N_A_27_368#_c_573_n N_Y_M1025_d 0.00250873f $X=4.015 $Y=2.99 $X2=0 $Y2=0
cc_493 N_A_27_368#_M1021_d N_Y_c_748_n 0.00408911f $X=1.08 $Y=1.84 $X2=0 $Y2=0
cc_494 N_A_27_368#_c_667_p N_Y_c_748_n 0.0136682f $X=1.23 $Y=2.455 $X2=0 $Y2=0
cc_495 N_A_27_368#_M1032_d N_Y_c_752_n 0.00524356f $X=1.98 $Y=1.84 $X2=0 $Y2=0
cc_496 N_A_27_368#_c_592_n N_Y_c_752_n 0.0202249f $X=2.18 $Y=2.455 $X2=0 $Y2=0
cc_497 N_A_27_368#_M1015_s N_Y_c_768_n 0.00455969f $X=2.98 $Y=1.84 $X2=0 $Y2=0
cc_498 N_A_27_368#_c_596_n N_Y_c_768_n 0.0202249f $X=3.18 $Y=2.455 $X2=0 $Y2=0
cc_499 N_A_27_368#_M1034_s N_Y_c_772_n 0.0152091f $X=3.98 $Y=1.84 $X2=0 $Y2=0
cc_500 N_A_27_368#_M1012_s N_Y_c_772_n 0.00359365f $X=5.12 $Y=1.84 $X2=0 $Y2=0
cc_501 N_A_27_368#_M1026_s N_Y_c_772_n 0.00452588f $X=6.12 $Y=1.84 $X2=0 $Y2=0
cc_502 N_A_27_368#_c_675_p N_Y_c_772_n 0.0250584f $X=4.18 $Y=2.46 $X2=0 $Y2=0
cc_503 N_A_27_368#_c_604_n N_Y_c_772_n 0.0413277f $X=5.105 $Y=2.375 $X2=0 $Y2=0
cc_504 N_A_27_368#_c_606_n N_Y_c_772_n 0.039006f $X=6.105 $Y=2.375 $X2=0 $Y2=0
cc_505 N_A_27_368#_c_582_n N_Y_c_772_n 0.0173542f $X=5.27 $Y=2.455 $X2=0 $Y2=0
cc_506 N_A_27_368#_c_583_n N_Y_c_772_n 0.0164906f $X=6.27 $Y=2.455 $X2=0 $Y2=0
cc_507 N_A_27_368#_M1026_s N_Y_c_741_n 0.00270113f $X=6.12 $Y=1.84 $X2=0 $Y2=0
cc_508 N_A_27_368#_c_569_n N_Y_c_753_n 0.0185424f $X=1.145 $Y=2.99 $X2=0 $Y2=0
cc_509 N_A_27_368#_c_667_p N_Y_c_753_n 0.0289859f $X=1.23 $Y=2.455 $X2=0 $Y2=0
cc_510 N_A_27_368#_c_667_p N_Y_c_757_n 0.0289859f $X=1.23 $Y=2.455 $X2=0 $Y2=0
cc_511 N_A_27_368#_c_571_n N_Y_c_757_n 0.0160777f $X=2.015 $Y=2.99 $X2=0 $Y2=0
cc_512 N_A_27_368#_c_572_n N_Y_c_780_n 0.018923f $X=3.015 $Y=2.99 $X2=0 $Y2=0
cc_513 N_A_27_368#_c_573_n N_Y_c_785_n 0.018923f $X=4.015 $Y=2.99 $X2=0 $Y2=0
cc_514 N_A_27_368#_c_604_n N_VPWR_M1007_d 0.00481401f $X=5.105 $Y=2.375
+ $X2=-0.19 $Y2=1.66
cc_515 N_A_27_368#_c_606_n N_VPWR_M1016_d 0.00620588f $X=6.105 $Y=2.375 $X2=0
+ $Y2=0
cc_516 N_A_27_368#_c_614_n N_VPWR_M1001_s 0.00771636f $X=7.105 $Y=2.375 $X2=0
+ $Y2=0
cc_517 N_A_27_368#_c_630_n N_VPWR_M1017_s 0.00455969f $X=8.105 $Y=2.035 $X2=0
+ $Y2=0
cc_518 N_A_27_368#_c_635_n N_VPWR_M1002_d 0.00508935f $X=9.105 $Y=2.035 $X2=0
+ $Y2=0
cc_519 N_A_27_368#_c_650_n N_VPWR_M1027_d 0.00604077f $X=10.11 $Y=2.035 $X2=0
+ $Y2=0
cc_520 N_A_27_368#_c_573_n N_VPWR_c_866_n 0.0103383f $X=4.015 $Y=2.99 $X2=0
+ $Y2=0
cc_521 N_A_27_368#_c_603_n N_VPWR_c_866_n 0.0153822f $X=4.18 $Y=2.905 $X2=0
+ $Y2=0
cc_522 N_A_27_368#_c_604_n N_VPWR_c_866_n 0.0202249f $X=5.105 $Y=2.375 $X2=0
+ $Y2=0
cc_523 N_A_27_368#_c_582_n N_VPWR_c_866_n 0.0139233f $X=5.27 $Y=2.455 $X2=0
+ $Y2=0
cc_524 N_A_27_368#_c_606_n N_VPWR_c_867_n 0.0232685f $X=6.105 $Y=2.375 $X2=0
+ $Y2=0
cc_525 N_A_27_368#_c_582_n N_VPWR_c_867_n 0.0139233f $X=5.27 $Y=2.455 $X2=0
+ $Y2=0
cc_526 N_A_27_368#_c_583_n N_VPWR_c_867_n 0.0139233f $X=6.27 $Y=2.455 $X2=0
+ $Y2=0
cc_527 N_A_27_368#_c_614_n N_VPWR_c_868_n 0.022455f $X=7.105 $Y=2.375 $X2=0
+ $Y2=0
cc_528 N_A_27_368#_c_574_n N_VPWR_c_868_n 0.0139233f $X=7.27 $Y=2.815 $X2=0
+ $Y2=0
cc_529 N_A_27_368#_c_583_n N_VPWR_c_868_n 0.0139233f $X=6.27 $Y=2.455 $X2=0
+ $Y2=0
cc_530 N_A_27_368#_c_574_n N_VPWR_c_869_n 0.0202646f $X=7.27 $Y=2.815 $X2=0
+ $Y2=0
cc_531 N_A_27_368#_c_630_n N_VPWR_c_869_n 0.0202249f $X=8.105 $Y=2.035 $X2=0
+ $Y2=0
cc_532 N_A_27_368#_c_575_n N_VPWR_c_869_n 0.0266809f $X=8.27 $Y=2.815 $X2=0
+ $Y2=0
cc_533 N_A_27_368#_c_575_n N_VPWR_c_870_n 0.0266809f $X=8.27 $Y=2.815 $X2=0
+ $Y2=0
cc_534 N_A_27_368#_c_635_n N_VPWR_c_870_n 0.0202249f $X=9.105 $Y=2.035 $X2=0
+ $Y2=0
cc_535 N_A_27_368#_c_576_n N_VPWR_c_870_n 0.0266809f $X=9.27 $Y=2.815 $X2=0
+ $Y2=0
cc_536 N_A_27_368#_c_576_n N_VPWR_c_871_n 0.0266809f $X=9.27 $Y=2.815 $X2=0
+ $Y2=0
cc_537 N_A_27_368#_c_650_n N_VPWR_c_871_n 0.0236753f $X=10.11 $Y=2.035 $X2=0
+ $Y2=0
cc_538 N_A_27_368#_c_578_n N_VPWR_c_871_n 0.0260697f $X=10.275 $Y=2.815 $X2=0
+ $Y2=0
cc_539 N_A_27_368#_c_569_n N_VPWR_c_872_n 0.0441932f $X=1.145 $Y=2.99 $X2=0
+ $Y2=0
cc_540 N_A_27_368#_c_570_n N_VPWR_c_872_n 0.0236215f $X=0.445 $Y=2.99 $X2=0
+ $Y2=0
cc_541 N_A_27_368#_c_571_n N_VPWR_c_872_n 0.0441612f $X=2.015 $Y=2.99 $X2=0
+ $Y2=0
cc_542 N_A_27_368#_c_572_n N_VPWR_c_872_n 0.0422753f $X=3.015 $Y=2.99 $X2=0
+ $Y2=0
cc_543 N_A_27_368#_c_573_n N_VPWR_c_872_n 0.0659319f $X=4.015 $Y=2.99 $X2=0
+ $Y2=0
cc_544 N_A_27_368#_c_579_n N_VPWR_c_872_n 0.0121867f $X=1.23 $Y=2.99 $X2=0 $Y2=0
cc_545 N_A_27_368#_c_580_n N_VPWR_c_872_n 0.0236039f $X=2.18 $Y=2.99 $X2=0 $Y2=0
cc_546 N_A_27_368#_c_581_n N_VPWR_c_872_n 0.0236039f $X=3.18 $Y=2.99 $X2=0 $Y2=0
cc_547 N_A_27_368#_c_582_n N_VPWR_c_874_n 0.0145674f $X=5.27 $Y=2.455 $X2=0
+ $Y2=0
cc_548 N_A_27_368#_c_583_n N_VPWR_c_876_n 0.0145974f $X=6.27 $Y=2.455 $X2=0
+ $Y2=0
cc_549 N_A_27_368#_c_574_n N_VPWR_c_878_n 0.014552f $X=7.27 $Y=2.815 $X2=0 $Y2=0
cc_550 N_A_27_368#_c_575_n N_VPWR_c_880_n 0.0145938f $X=8.27 $Y=2.815 $X2=0
+ $Y2=0
cc_551 N_A_27_368#_c_576_n N_VPWR_c_882_n 0.0145938f $X=9.27 $Y=2.815 $X2=0
+ $Y2=0
cc_552 N_A_27_368#_c_578_n N_VPWR_c_883_n 0.0145938f $X=10.275 $Y=2.815 $X2=0
+ $Y2=0
cc_553 N_A_27_368#_c_569_n N_VPWR_c_865_n 0.0249913f $X=1.145 $Y=2.99 $X2=0
+ $Y2=0
cc_554 N_A_27_368#_c_570_n N_VPWR_c_865_n 0.0127839f $X=0.445 $Y=2.99 $X2=0
+ $Y2=0
cc_555 N_A_27_368#_c_571_n N_VPWR_c_865_n 0.0249452f $X=2.015 $Y=2.99 $X2=0
+ $Y2=0
cc_556 N_A_27_368#_c_572_n N_VPWR_c_865_n 0.0238861f $X=3.015 $Y=2.99 $X2=0
+ $Y2=0
cc_557 N_A_27_368#_c_573_n N_VPWR_c_865_n 0.0367158f $X=4.015 $Y=2.99 $X2=0
+ $Y2=0
cc_558 N_A_27_368#_c_574_n N_VPWR_c_865_n 0.0119791f $X=7.27 $Y=2.815 $X2=0
+ $Y2=0
cc_559 N_A_27_368#_c_575_n N_VPWR_c_865_n 0.0120466f $X=8.27 $Y=2.815 $X2=0
+ $Y2=0
cc_560 N_A_27_368#_c_576_n N_VPWR_c_865_n 0.0120466f $X=9.27 $Y=2.815 $X2=0
+ $Y2=0
cc_561 N_A_27_368#_c_578_n N_VPWR_c_865_n 0.0120466f $X=10.275 $Y=2.815 $X2=0
+ $Y2=0
cc_562 N_A_27_368#_c_579_n N_VPWR_c_865_n 0.00660921f $X=1.23 $Y=2.99 $X2=0
+ $Y2=0
cc_563 N_A_27_368#_c_580_n N_VPWR_c_865_n 0.012761f $X=2.18 $Y=2.99 $X2=0 $Y2=0
cc_564 N_A_27_368#_c_581_n N_VPWR_c_865_n 0.012761f $X=3.18 $Y=2.99 $X2=0 $Y2=0
cc_565 N_A_27_368#_c_582_n N_VPWR_c_865_n 0.0119851f $X=5.27 $Y=2.455 $X2=0
+ $Y2=0
cc_566 N_A_27_368#_c_583_n N_VPWR_c_865_n 0.0120334f $X=6.27 $Y=2.455 $X2=0
+ $Y2=0
cc_567 N_Y_c_772_n N_VPWR_M1007_d 0.0045658f $X=6.18 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_568 N_Y_c_772_n N_VPWR_M1016_d 0.0063196f $X=6.18 $Y=2.035 $X2=0 $Y2=0
cc_569 N_Y_c_740_n N_A_27_74#_M1023_d 0.00255298f $X=3.51 $Y=1.03 $X2=0 $Y2=0
cc_570 N_Y_c_745_n N_A_27_74#_M1037_d 0.00372475f $X=4.82 $Y=0.975 $X2=0 $Y2=0
cc_571 N_Y_c_742_n N_A_27_74#_c_1000_n 0.009209f $X=2.565 $Y=0.86 $X2=0 $Y2=0
cc_572 N_Y_M1014_s N_A_27_74#_c_1001_n 0.00176461f $X=2.425 $Y=0.37 $X2=0 $Y2=0
cc_573 N_Y_c_740_n N_A_27_74#_c_1001_n 0.0039879f $X=3.51 $Y=1.03 $X2=0 $Y2=0
cc_574 N_Y_c_742_n N_A_27_74#_c_1001_n 0.0158692f $X=2.565 $Y=0.86 $X2=0 $Y2=0
cc_575 N_Y_M1030_s N_A_27_74#_c_1003_n 0.00285125f $X=3.355 $Y=0.37 $X2=0 $Y2=0
cc_576 N_Y_c_740_n N_A_27_74#_c_1003_n 0.0108211f $X=3.51 $Y=1.03 $X2=0 $Y2=0
cc_577 N_Y_c_745_n N_A_27_74#_c_1003_n 0.0012223f $X=4.82 $Y=0.975 $X2=0 $Y2=0
cc_578 N_Y_c_740_n N_A_27_74#_c_1005_n 0.0211547f $X=3.51 $Y=1.03 $X2=0 $Y2=0
cc_579 N_Y_c_745_n N_A_27_74#_c_1006_n 0.0139452f $X=4.82 $Y=0.975 $X2=0 $Y2=0
cc_580 N_Y_c_745_n N_A_868_74#_M1005_d 0.00299905f $X=4.82 $Y=0.975 $X2=-0.19
+ $Y2=-0.245
cc_581 N_Y_c_744_n N_A_868_74#_M1022_d 0.00177442f $X=6.18 $Y=0.95 $X2=0 $Y2=0
cc_582 N_Y_c_744_n N_A_868_74#_M1038_d 0.00535397f $X=6.18 $Y=0.95 $X2=0 $Y2=0
cc_583 N_Y_c_745_n N_A_868_74#_c_1182_n 0.0214055f $X=4.82 $Y=0.975 $X2=0 $Y2=0
cc_584 N_Y_M1005_s N_A_868_74#_c_1184_n 0.00254491f $X=4.775 $Y=0.37 $X2=0 $Y2=0
cc_585 N_Y_M1031_s N_A_868_74#_c_1184_n 0.00179007f $X=5.705 $Y=0.37 $X2=0 $Y2=0
cc_586 N_Y_c_744_n N_A_868_74#_c_1184_n 0.0127448f $X=6.18 $Y=0.95 $X2=0 $Y2=0
cc_587 N_Y_c_745_n N_A_868_74#_c_1184_n 0.00412076f $X=4.82 $Y=0.975 $X2=0 $Y2=0
cc_588 N_Y_c_746_n N_A_868_74#_c_1184_n 0.0755709f $X=5.15 $Y=0.975 $X2=0 $Y2=0
cc_589 N_Y_c_741_n N_A_1313_74#_c_1226_n 0.00356311f $X=6.265 $Y=1.95 $X2=0
+ $Y2=0
cc_590 N_Y_c_744_n N_A_1313_74#_c_1226_n 0.0284876f $X=6.18 $Y=0.95 $X2=0 $Y2=0
cc_591 N_A_27_74#_c_997_n N_VGND_M1009_s 0.00250873f $X=1.125 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_592 N_A_27_74#_c_1000_n N_VGND_M1029_s 0.00245557f $X=2.05 $Y=1.095 $X2=0
+ $Y2=0
cc_593 N_A_27_74#_c_996_n N_VGND_c_1070_n 0.0191765f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_594 N_A_27_74#_c_997_n N_VGND_c_1070_n 0.0210288f $X=1.125 $Y=1.095 $X2=0
+ $Y2=0
cc_595 N_A_27_74#_c_999_n N_VGND_c_1070_n 0.0182488f $X=1.21 $Y=0.515 $X2=0
+ $Y2=0
cc_596 N_A_27_74#_c_999_n N_VGND_c_1071_n 0.0182488f $X=1.21 $Y=0.515 $X2=0
+ $Y2=0
cc_597 N_A_27_74#_c_1000_n N_VGND_c_1071_n 0.020622f $X=2.05 $Y=1.095 $X2=0
+ $Y2=0
cc_598 N_A_27_74#_c_1002_n N_VGND_c_1071_n 0.00779323f $X=2.22 $Y=0.34 $X2=0
+ $Y2=0
cc_599 N_A_27_74#_c_996_n N_VGND_c_1076_n 0.0145639f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_600 N_A_27_74#_c_999_n N_VGND_c_1077_n 0.00749631f $X=1.21 $Y=0.515 $X2=0
+ $Y2=0
cc_601 N_A_27_74#_c_1001_n N_VGND_c_1078_n 0.042902f $X=2.9 $Y=0.34 $X2=0 $Y2=0
cc_602 N_A_27_74#_c_1002_n N_VGND_c_1078_n 0.0121867f $X=2.22 $Y=0.34 $X2=0
+ $Y2=0
cc_603 N_A_27_74#_c_1003_n N_VGND_c_1078_n 0.033414f $X=3.76 $Y=0.34 $X2=0 $Y2=0
cc_604 N_A_27_74#_c_1005_n N_VGND_c_1078_n 0.0227371f $X=3.065 $Y=0.34 $X2=0
+ $Y2=0
cc_605 N_A_27_74#_c_1006_n N_VGND_c_1078_n 0.0227371f $X=3.925 $Y=0.34 $X2=0
+ $Y2=0
cc_606 N_A_27_74#_c_996_n N_VGND_c_1085_n 0.0119984f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_607 N_A_27_74#_c_999_n N_VGND_c_1085_n 0.0062048f $X=1.21 $Y=0.515 $X2=0
+ $Y2=0
cc_608 N_A_27_74#_c_1001_n N_VGND_c_1085_n 0.0241973f $X=2.9 $Y=0.34 $X2=0 $Y2=0
cc_609 N_A_27_74#_c_1002_n N_VGND_c_1085_n 0.00660921f $X=2.22 $Y=0.34 $X2=0
+ $Y2=0
cc_610 N_A_27_74#_c_1003_n N_VGND_c_1085_n 0.0187892f $X=3.76 $Y=0.34 $X2=0
+ $Y2=0
cc_611 N_A_27_74#_c_1005_n N_VGND_c_1085_n 0.0125119f $X=3.065 $Y=0.34 $X2=0
+ $Y2=0
cc_612 N_A_27_74#_c_1006_n N_VGND_c_1085_n 0.0125119f $X=3.925 $Y=0.34 $X2=0
+ $Y2=0
cc_613 N_A_27_74#_c_1006_n N_A_868_74#_c_1182_n 0.0242706f $X=3.925 $Y=0.34
+ $X2=0 $Y2=0
cc_614 N_VGND_c_1078_n N_A_868_74#_c_1182_n 0.0142249f $X=8.395 $Y=0 $X2=0 $Y2=0
cc_615 N_VGND_c_1085_n N_A_868_74#_c_1182_n 0.011867f $X=10.32 $Y=0 $X2=0 $Y2=0
cc_616 N_VGND_c_1072_n N_A_868_74#_c_1183_n 0.0231578f $X=8.56 $Y=0.595 $X2=0
+ $Y2=0
cc_617 N_VGND_c_1078_n N_A_868_74#_c_1184_n 0.142724f $X=8.395 $Y=0 $X2=0 $Y2=0
cc_618 N_VGND_c_1085_n N_A_868_74#_c_1184_n 0.120136f $X=10.32 $Y=0 $X2=0 $Y2=0
cc_619 N_VGND_M1004_d N_A_1313_74#_c_1222_n 0.00299905f $X=8.415 $Y=0.37 $X2=0
+ $Y2=0
cc_620 N_VGND_c_1072_n N_A_1313_74#_c_1222_n 0.0219827f $X=8.56 $Y=0.595 $X2=0
+ $Y2=0
cc_621 N_VGND_c_1072_n N_A_1313_74#_c_1223_n 0.0182488f $X=8.56 $Y=0.595 $X2=0
+ $Y2=0
cc_622 N_VGND_c_1073_n N_A_1313_74#_c_1223_n 0.0182488f $X=9.42 $Y=0.595 $X2=0
+ $Y2=0
cc_623 N_VGND_c_1079_n N_A_1313_74#_c_1223_n 0.00749631f $X=9.255 $Y=0 $X2=0
+ $Y2=0
cc_624 N_VGND_c_1085_n N_A_1313_74#_c_1223_n 0.0062048f $X=10.32 $Y=0 $X2=0
+ $Y2=0
cc_625 N_VGND_M1020_d N_A_1313_74#_c_1224_n 0.00176461f $X=9.28 $Y=0.37 $X2=0
+ $Y2=0
cc_626 N_VGND_c_1073_n N_A_1313_74#_c_1224_n 0.0171619f $X=9.42 $Y=0.595 $X2=0
+ $Y2=0
cc_627 N_VGND_c_1075_n N_A_1313_74#_c_1224_n 0.00517071f $X=10.28 $Y=0.515 $X2=0
+ $Y2=0
cc_628 N_VGND_c_1073_n N_A_1313_74#_c_1225_n 0.0182488f $X=9.42 $Y=0.595 $X2=0
+ $Y2=0
cc_629 N_VGND_c_1075_n N_A_1313_74#_c_1225_n 0.0243418f $X=10.28 $Y=0.515 $X2=0
+ $Y2=0
cc_630 N_VGND_c_1080_n N_A_1313_74#_c_1225_n 0.00749631f $X=10.115 $Y=0 $X2=0
+ $Y2=0
cc_631 N_VGND_c_1085_n N_A_1313_74#_c_1225_n 0.0062048f $X=10.32 $Y=0 $X2=0
+ $Y2=0
cc_632 N_A_868_74#_c_1184_n N_A_1313_74#_M1003_s 0.00179007f $X=7.835 $Y=0.515
+ $X2=-0.19 $Y2=-0.245
cc_633 N_A_868_74#_c_1184_n N_A_1313_74#_M1018_s 0.00212678f $X=7.835 $Y=0.515
+ $X2=0 $Y2=0
cc_634 N_A_868_74#_M1019_d N_A_1313_74#_c_1222_n 0.00388574f $X=7.86 $Y=0.37
+ $X2=0 $Y2=0
cc_635 N_A_868_74#_c_1183_n N_A_1313_74#_c_1222_n 0.0127309f $X=8 $Y=0.515 $X2=0
+ $Y2=0
cc_636 N_A_868_74#_c_1184_n N_A_1313_74#_c_1222_n 0.00339963f $X=7.835 $Y=0.515
+ $X2=0 $Y2=0
cc_637 N_A_868_74#_c_1184_n N_A_1313_74#_c_1226_n 0.0163588f $X=7.835 $Y=0.515
+ $X2=0 $Y2=0
cc_638 N_A_868_74#_M1006_d N_A_1313_74#_c_1227_n 0.00217299f $X=6.995 $Y=0.37
+ $X2=0 $Y2=0
cc_639 N_A_868_74#_c_1184_n N_A_1313_74#_c_1227_n 0.0336602f $X=7.835 $Y=0.515
+ $X2=0 $Y2=0
