* File: sky130_fd_sc_ls__or2b_4.pxi.spice
* Created: Wed Sep  2 11:24:38 2020
* 
x_PM_SKY130_FD_SC_LS__OR2B_4%A_81_296# N_A_81_296#_M1004_d N_A_81_296#_M1009_d
+ N_A_81_296#_M1001_d N_A_81_296#_M1008_g N_A_81_296#_c_129_n
+ N_A_81_296#_M1000_g N_A_81_296#_c_114_n N_A_81_296#_M1011_g
+ N_A_81_296#_c_130_n N_A_81_296#_M1003_g N_A_81_296#_c_131_n
+ N_A_81_296#_M1012_g N_A_81_296#_M1014_g N_A_81_296#_c_132_n
+ N_A_81_296#_M1013_g N_A_81_296#_M1015_g N_A_81_296#_c_118_n
+ N_A_81_296#_c_119_n N_A_81_296#_c_120_n N_A_81_296#_c_121_n
+ N_A_81_296#_c_122_n N_A_81_296#_c_123_n N_A_81_296#_c_124_n
+ N_A_81_296#_c_125_n N_A_81_296#_c_126_n N_A_81_296#_c_127_n
+ N_A_81_296#_c_128_n PM_SKY130_FD_SC_LS__OR2B_4%A_81_296#
x_PM_SKY130_FD_SC_LS__OR2B_4%A N_A_M1004_g N_A_c_260_n N_A_c_267_n N_A_M1002_g
+ N_A_c_261_n N_A_c_262_n N_A_M1007_g N_A_M1010_g N_A_c_264_n A A
+ PM_SKY130_FD_SC_LS__OR2B_4%A
x_PM_SKY130_FD_SC_LS__OR2B_4%A_676_48# N_A_676_48#_M1016_d N_A_676_48#_M1006_d
+ N_A_676_48#_M1009_g N_A_676_48#_c_319_n N_A_676_48#_c_320_n
+ N_A_676_48#_c_321_n N_A_676_48#_c_332_n N_A_676_48#_M1001_g
+ N_A_676_48#_M1017_g N_A_676_48#_c_323_n N_A_676_48#_c_324_n
+ N_A_676_48#_M1005_g N_A_676_48#_c_325_n N_A_676_48#_c_326_n
+ N_A_676_48#_c_327_n N_A_676_48#_c_328_n N_A_676_48#_c_329_n
+ N_A_676_48#_c_330_n PM_SKY130_FD_SC_LS__OR2B_4%A_676_48#
x_PM_SKY130_FD_SC_LS__OR2B_4%B_N N_B_N_c_405_n N_B_N_M1016_g N_B_N_c_406_n
+ N_B_N_c_407_n N_B_N_c_410_n N_B_N_M1006_g N_B_N_c_408_n B_N B_N N_B_N_c_409_n
+ PM_SKY130_FD_SC_LS__OR2B_4%B_N
x_PM_SKY130_FD_SC_LS__OR2B_4%VPWR N_VPWR_M1000_s N_VPWR_M1003_s N_VPWR_M1013_s
+ N_VPWR_M1007_s N_VPWR_M1006_s N_VPWR_c_442_n N_VPWR_c_443_n N_VPWR_c_444_n
+ N_VPWR_c_445_n N_VPWR_c_446_n N_VPWR_c_447_n N_VPWR_c_448_n N_VPWR_c_449_n
+ N_VPWR_c_450_n N_VPWR_c_451_n VPWR N_VPWR_c_452_n N_VPWR_c_453_n
+ N_VPWR_c_454_n N_VPWR_c_441_n N_VPWR_c_456_n N_VPWR_c_457_n
+ PM_SKY130_FD_SC_LS__OR2B_4%VPWR
x_PM_SKY130_FD_SC_LS__OR2B_4%X N_X_M1008_s N_X_M1014_s N_X_M1000_d N_X_M1012_d
+ N_X_c_521_n N_X_c_522_n N_X_c_523_n N_X_c_528_n N_X_c_524_n N_X_c_529_n
+ N_X_c_530_n N_X_c_525_n N_X_c_526_n N_X_c_531_n X PM_SKY130_FD_SC_LS__OR2B_4%X
x_PM_SKY130_FD_SC_LS__OR2B_4%A_489_392# N_A_489_392#_M1002_d
+ N_A_489_392#_M1001_s N_A_489_392#_M1005_s N_A_489_392#_c_594_n
+ N_A_489_392#_c_595_n N_A_489_392#_c_596_n N_A_489_392#_c_597_n
+ N_A_489_392#_c_598_n N_A_489_392#_c_599_n N_A_489_392#_c_600_n
+ N_A_489_392#_c_601_n PM_SKY130_FD_SC_LS__OR2B_4%A_489_392#
x_PM_SKY130_FD_SC_LS__OR2B_4%VGND N_VGND_M1008_d N_VGND_M1011_d N_VGND_M1015_d
+ N_VGND_M1010_s N_VGND_M1017_s N_VGND_c_647_n N_VGND_c_648_n N_VGND_c_649_n
+ N_VGND_c_650_n N_VGND_c_651_n N_VGND_c_652_n VGND N_VGND_c_653_n
+ N_VGND_c_654_n N_VGND_c_655_n N_VGND_c_656_n N_VGND_c_657_n N_VGND_c_658_n
+ N_VGND_c_659_n N_VGND_c_660_n N_VGND_c_661_n N_VGND_c_662_n
+ PM_SKY130_FD_SC_LS__OR2B_4%VGND
cc_1 VNB N_A_81_296#_M1008_g 0.0363403f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_A_81_296#_c_114_n 0.014897f $X=-0.19 $Y=-0.245 $X2=0.85 $Y2=1.555
cc_3 VNB N_A_81_296#_M1011_g 0.021162f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.74
cc_4 VNB N_A_81_296#_M1014_g 0.0220733f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=0.74
cc_5 VNB N_A_81_296#_M1015_g 0.0223805f $X=-0.19 $Y=-0.245 $X2=1.88 $Y2=0.74
cc_6 VNB N_A_81_296#_c_118_n 0.014013f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.555
cc_7 VNB N_A_81_296#_c_119_n 0.0021705f $X=-0.19 $Y=-0.245 $X2=1.975 $Y2=1.465
cc_8 VNB N_A_81_296#_c_120_n 0.00687872f $X=-0.19 $Y=-0.245 $X2=2.475 $Y2=1.195
cc_9 VNB N_A_81_296#_c_121_n 0.00553968f $X=-0.19 $Y=-0.245 $X2=2.64 $Y2=0.515
cc_10 VNB N_A_81_296#_c_122_n 0.0119082f $X=-0.19 $Y=-0.245 $X2=3.505 $Y2=1.195
cc_11 VNB N_A_81_296#_c_123_n 0.00307801f $X=-0.19 $Y=-0.245 $X2=3.67 $Y2=0.515
cc_12 VNB N_A_81_296#_c_124_n 3.78434e-19 $X=-0.19 $Y=-0.245 $X2=4.04 $Y2=2.08
cc_13 VNB N_A_81_296#_c_125_n 0.00796175f $X=-0.19 $Y=-0.245 $X2=2.06 $Y2=1.195
cc_14 VNB N_A_81_296#_c_126_n 0.00312763f $X=-0.19 $Y=-0.245 $X2=2.64 $Y2=1.195
cc_15 VNB N_A_81_296#_c_127_n 0.007464f $X=-0.19 $Y=-0.245 $X2=3.63 $Y2=1.28
cc_16 VNB N_A_81_296#_c_128_n 0.0735405f $X=-0.19 $Y=-0.245 $X2=1.845 $Y2=1.532
cc_17 VNB N_A_M1004_g 0.0360123f $X=-0.19 $Y=-0.245 $X2=3.89 $Y2=1.935
cc_18 VNB N_A_c_260_n 0.00382132f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_c_261_n 0.00993221f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.48
cc_20 VNB N_A_c_262_n 0.0148358f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_21 VNB N_A_M1010_g 0.0365137f $X=-0.19 $Y=-0.245 $X2=0.85 $Y2=1.555
cc_22 VNB N_A_c_264_n 0.006075f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.3
cc_23 VNB A 0.0049455f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.74
cc_24 VNB N_A_676_48#_M1009_g 0.0331319f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_676_48#_c_319_n 0.0119927f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_26 VNB N_A_676_48#_c_320_n 0.0101155f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_27 VNB N_A_676_48#_c_321_n 0.00403268f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.765
cc_28 VNB N_A_676_48#_M1017_g 0.035707f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.74
cc_29 VNB N_A_676_48#_c_323_n 0.0121834f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_676_48#_c_324_n 0.0237216f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=2.4
cc_31 VNB N_A_676_48#_c_325_n 0.00374105f $X=-0.19 $Y=-0.245 $X2=1.395 $Y2=2.4
cc_32 VNB N_A_676_48#_c_326_n 0.00141541f $X=-0.19 $Y=-0.245 $X2=1.395 $Y2=2.4
cc_33 VNB N_A_676_48#_c_327_n 0.0385846f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=0.74
cc_34 VNB N_A_676_48#_c_328_n 0.0379768f $X=-0.19 $Y=-0.245 $X2=1.88 $Y2=1.3
cc_35 VNB N_A_676_48#_c_329_n 0.00186199f $X=-0.19 $Y=-0.245 $X2=1.975 $Y2=1.465
cc_36 VNB N_A_676_48#_c_330_n 0.00618737f $X=-0.19 $Y=-0.245 $X2=1.11 $Y2=1.465
cc_37 VNB N_B_N_c_405_n 0.0204172f $X=-0.19 $Y=-0.245 $X2=2.43 $Y2=0.37
cc_38 VNB N_B_N_c_406_n 0.0538601f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_B_N_c_407_n 0.00815644f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_B_N_c_408_n 0.00703507f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.48
cc_41 VNB N_B_N_c_409_n 0.0316413f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_42 VNB N_VPWR_c_441_n 0.243291f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.532
cc_43 VNB N_X_c_521_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_44 VNB N_X_c_522_n 0.0041248f $X=-0.19 $Y=-0.245 $X2=0.85 $Y2=1.555
cc_45 VNB N_X_c_523_n 0.00156967f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.555
cc_46 VNB N_X_c_524_n 0.0060023f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=2.4
cc_47 VNB N_X_c_525_n 0.00280814f $X=-0.19 $Y=-0.245 $X2=1.88 $Y2=0.74
cc_48 VNB N_X_c_526_n 0.0182272f $X=-0.19 $Y=-0.245 $X2=1.975 $Y2=1.465
cc_49 VNB N_VGND_c_647_n 0.010678f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_50 VNB N_VGND_c_648_n 0.0354929f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.555
cc_51 VNB N_VGND_c_649_n 0.00509474f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_650_n 0.00577125f $X=-0.19 $Y=-0.245 $X2=1.395 $Y2=1.765
cc_53 VNB N_VGND_c_651_n 0.00558127f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=0.74
cc_54 VNB N_VGND_c_652_n 0.00923674f $X=-0.19 $Y=-0.245 $X2=1.845 $Y2=2.4
cc_55 VNB N_VGND_c_653_n 0.0172524f $X=-0.19 $Y=-0.245 $X2=1.88 $Y2=0.74
cc_56 VNB N_VGND_c_654_n 0.018682f $X=-0.19 $Y=-0.245 $X2=1.11 $Y2=1.465
cc_57 VNB N_VGND_c_655_n 0.0193334f $X=-0.19 $Y=-0.245 $X2=1.79 $Y2=1.465
cc_58 VNB N_VGND_c_656_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=2.64 $Y2=0.515
cc_59 VNB N_VGND_c_657_n 0.0401986f $X=-0.19 $Y=-0.245 $X2=4.04 $Y2=2.08
cc_60 VNB N_VGND_c_658_n 0.324755f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_659_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=3.63 $Y2=1.28
cc_62 VNB N_VGND_c_660_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=1.532
cc_63 VNB N_VGND_c_661_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=1.532
cc_64 VNB N_VGND_c_662_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=1.88 $Y2=1.532
cc_65 VPB N_A_81_296#_c_129_n 0.018685f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.765
cc_66 VPB N_A_81_296#_c_130_n 0.0147054f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=1.765
cc_67 VPB N_A_81_296#_c_131_n 0.0152275f $X=-0.19 $Y=1.66 $X2=1.395 $Y2=1.765
cc_68 VPB N_A_81_296#_c_132_n 0.01624f $X=-0.19 $Y=1.66 $X2=1.845 $Y2=1.765
cc_69 VPB N_A_81_296#_c_118_n 0.00997134f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.555
cc_70 VPB N_A_81_296#_c_124_n 0.00237762f $X=-0.19 $Y=1.66 $X2=4.04 $Y2=2.08
cc_71 VPB N_A_81_296#_c_128_n 0.0199032f $X=-0.19 $Y=1.66 $X2=1.845 $Y2=1.532
cc_72 VPB N_A_c_260_n 0.00756645f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_A_c_267_n 0.0228348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_A_c_262_n 0.039148f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_75 VPB A 0.00637848f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=0.74
cc_76 VPB N_A_676_48#_c_321_n 0.00686816f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.765
cc_77 VPB N_A_676_48#_c_332_n 0.0251503f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_78 VPB N_A_676_48#_c_324_n 0.0431377f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=2.4
cc_79 VPB N_A_676_48#_c_328_n 0.0561025f $X=-0.19 $Y=1.66 $X2=1.88 $Y2=1.3
cc_80 VPB N_A_676_48#_c_329_n 0.00251184f $X=-0.19 $Y=1.66 $X2=1.975 $Y2=1.465
cc_81 VPB N_B_N_c_410_n 0.0222313f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 VPB N_B_N_c_408_n 0.028679f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.48
cc_83 VPB B_N 0.00252041f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_84 VPB N_VPWR_c_442_n 0.0116916f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_85 VPB N_VPWR_c_443_n 0.0578904f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.555
cc_86 VPB N_VPWR_c_444_n 0.00504372f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=2.4
cc_87 VPB N_VPWR_c_445_n 0.00961427f $X=-0.19 $Y=1.66 $X2=1.395 $Y2=2.4
cc_88 VPB N_VPWR_c_446_n 0.0153769f $X=-0.19 $Y=1.66 $X2=1.845 $Y2=2.4
cc_89 VPB N_VPWR_c_447_n 0.0182617f $X=-0.19 $Y=1.66 $X2=1.88 $Y2=0.74
cc_90 VPB N_VPWR_c_448_n 0.0162121f $X=-0.19 $Y=1.66 $X2=1.11 $Y2=1.465
cc_91 VPB N_VPWR_c_449_n 0.00460249f $X=-0.19 $Y=1.66 $X2=1.11 $Y2=1.465
cc_92 VPB N_VPWR_c_450_n 0.0206041f $X=-0.19 $Y=1.66 $X2=1.79 $Y2=1.465
cc_93 VPB N_VPWR_c_451_n 0.0047828f $X=-0.19 $Y=1.66 $X2=1.79 $Y2=1.465
cc_94 VPB N_VPWR_c_452_n 0.020445f $X=-0.19 $Y=1.66 $X2=3.63 $Y2=1.11
cc_95 VPB N_VPWR_c_453_n 0.0413605f $X=-0.19 $Y=1.66 $X2=4 $Y2=1.45
cc_96 VPB N_VPWR_c_454_n 0.0177091f $X=-0.19 $Y=1.66 $X2=4 $Y2=1.28
cc_97 VPB N_VPWR_c_441_n 0.0981373f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.532
cc_98 VPB N_VPWR_c_456_n 0.0047828f $X=-0.19 $Y=1.66 $X2=1.845 $Y2=1.532
cc_99 VPB N_VPWR_c_457_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 VPB N_X_c_523_n 0.00252918f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.555
cc_101 VPB N_X_c_528_n 0.00207077f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=0.74
cc_102 VPB N_X_c_529_n 0.00419778f $X=-0.19 $Y=1.66 $X2=1.395 $Y2=2.4
cc_103 VPB N_X_c_530_n 0.00257348f $X=-0.19 $Y=1.66 $X2=1.425 $Y2=0.74
cc_104 VPB N_X_c_531_n 6.78741e-19 $X=-0.19 $Y=1.66 $X2=1.11 $Y2=1.465
cc_105 VPB N_A_489_392#_c_594_n 0.00303533f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.48
cc_106 VPB N_A_489_392#_c_595_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_107 VPB N_A_489_392#_c_596_n 0.0147762f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.765
cc_108 VPB N_A_489_392#_c_597_n 0.0034702f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_109 VPB N_A_489_392#_c_598_n 0.00741598f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.3
cc_110 VPB N_A_489_392#_c_599_n 0.00912105f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=0.74
cc_111 VPB N_A_489_392#_c_600_n 0.00391062f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=0.74
cc_112 VPB N_A_489_392#_c_601_n 0.00960504f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=2.4
cc_113 N_A_81_296#_M1015_g N_A_M1004_g 0.0123298f $X=1.88 $Y=0.74 $X2=0 $Y2=0
cc_114 N_A_81_296#_c_120_n N_A_M1004_g 0.0190817f $X=2.475 $Y=1.195 $X2=0 $Y2=0
cc_115 N_A_81_296#_c_121_n N_A_M1004_g 0.00597167f $X=2.64 $Y=0.515 $X2=0 $Y2=0
cc_116 N_A_81_296#_c_125_n N_A_M1004_g 0.00587547f $X=2.06 $Y=1.195 $X2=0 $Y2=0
cc_117 N_A_81_296#_c_132_n N_A_c_260_n 0.00437886f $X=1.845 $Y=1.765 $X2=0 $Y2=0
cc_118 N_A_81_296#_c_128_n N_A_c_260_n 0.00524362f $X=1.845 $Y=1.532 $X2=0 $Y2=0
cc_119 N_A_81_296#_c_132_n N_A_c_267_n 0.015849f $X=1.845 $Y=1.765 $X2=0 $Y2=0
cc_120 N_A_81_296#_c_126_n N_A_c_261_n 0.00685796f $X=2.64 $Y=1.195 $X2=0 $Y2=0
cc_121 N_A_81_296#_c_121_n N_A_M1010_g 0.0105092f $X=2.64 $Y=0.515 $X2=0 $Y2=0
cc_122 N_A_81_296#_c_122_n N_A_M1010_g 0.0155134f $X=3.505 $Y=1.195 $X2=0 $Y2=0
cc_123 N_A_81_296#_c_123_n N_A_M1010_g 7.89164e-19 $X=3.67 $Y=0.515 $X2=0 $Y2=0
cc_124 N_A_81_296#_c_127_n N_A_M1010_g 8.03754e-19 $X=3.63 $Y=1.28 $X2=0 $Y2=0
cc_125 N_A_81_296#_c_128_n N_A_c_264_n 0.0123298f $X=1.845 $Y=1.532 $X2=0 $Y2=0
cc_126 N_A_81_296#_c_122_n A 0.0325657f $X=3.505 $Y=1.195 $X2=0 $Y2=0
cc_127 N_A_81_296#_c_124_n A 0.00993913f $X=4.04 $Y=2.08 $X2=0 $Y2=0
cc_128 N_A_81_296#_c_125_n A 0.00800544f $X=2.06 $Y=1.195 $X2=0 $Y2=0
cc_129 N_A_81_296#_c_126_n A 0.0235756f $X=2.64 $Y=1.195 $X2=0 $Y2=0
cc_130 N_A_81_296#_c_122_n N_A_676_48#_M1009_g 0.0126768f $X=3.505 $Y=1.195
+ $X2=0 $Y2=0
cc_131 N_A_81_296#_c_123_n N_A_676_48#_M1009_g 0.0105052f $X=3.67 $Y=0.515 $X2=0
+ $Y2=0
cc_132 N_A_81_296#_c_127_n N_A_676_48#_M1009_g 0.00726533f $X=3.63 $Y=1.28 $X2=0
+ $Y2=0
cc_133 N_A_81_296#_c_127_n N_A_676_48#_c_319_n 0.00705335f $X=3.63 $Y=1.28 $X2=0
+ $Y2=0
cc_134 N_A_81_296#_c_127_n N_A_676_48#_c_320_n 4.99147e-19 $X=3.63 $Y=1.28 $X2=0
+ $Y2=0
cc_135 N_A_81_296#_c_124_n N_A_676_48#_c_321_n 0.00546594f $X=4.04 $Y=2.08 $X2=0
+ $Y2=0
cc_136 N_A_81_296#_c_124_n N_A_676_48#_c_332_n 0.0177535f $X=4.04 $Y=2.08 $X2=0
+ $Y2=0
cc_137 N_A_81_296#_c_123_n N_A_676_48#_M1017_g 0.00232377f $X=3.67 $Y=0.515
+ $X2=0 $Y2=0
cc_138 N_A_81_296#_c_127_n N_A_676_48#_M1017_g 0.0190269f $X=3.63 $Y=1.28 $X2=0
+ $Y2=0
cc_139 N_A_81_296#_c_124_n N_A_676_48#_c_323_n 0.00638285f $X=4.04 $Y=2.08 $X2=0
+ $Y2=0
cc_140 N_A_81_296#_c_127_n N_A_676_48#_c_323_n 0.00304884f $X=3.63 $Y=1.28 $X2=0
+ $Y2=0
cc_141 N_A_81_296#_c_124_n N_A_676_48#_c_324_n 0.00899763f $X=4.04 $Y=2.08 $X2=0
+ $Y2=0
cc_142 N_A_81_296#_c_124_n N_A_676_48#_c_325_n 0.00478313f $X=4.04 $Y=2.08 $X2=0
+ $Y2=0
cc_143 N_A_81_296#_c_127_n N_A_676_48#_c_325_n 0.00692478f $X=3.63 $Y=1.28 $X2=0
+ $Y2=0
cc_144 N_A_81_296#_c_124_n N_A_676_48#_c_329_n 0.0245536f $X=4.04 $Y=2.08 $X2=0
+ $Y2=0
cc_145 N_A_81_296#_c_127_n N_A_676_48#_c_329_n 3.96184e-19 $X=3.63 $Y=1.28 $X2=0
+ $Y2=0
cc_146 N_A_81_296#_c_127_n N_A_676_48#_c_330_n 0.00914716f $X=3.63 $Y=1.28 $X2=0
+ $Y2=0
cc_147 N_A_81_296#_c_129_n N_VPWR_c_443_n 0.0175194f $X=0.495 $Y=1.765 $X2=0
+ $Y2=0
cc_148 N_A_81_296#_c_130_n N_VPWR_c_443_n 6.37978e-19 $X=0.945 $Y=1.765 $X2=0
+ $Y2=0
cc_149 N_A_81_296#_c_118_n N_VPWR_c_443_n 4.5868e-19 $X=0.495 $Y=1.555 $X2=0
+ $Y2=0
cc_150 N_A_81_296#_c_129_n N_VPWR_c_444_n 5.83721e-19 $X=0.495 $Y=1.765 $X2=0
+ $Y2=0
cc_151 N_A_81_296#_c_130_n N_VPWR_c_444_n 0.0133451f $X=0.945 $Y=1.765 $X2=0
+ $Y2=0
cc_152 N_A_81_296#_c_131_n N_VPWR_c_444_n 0.00630489f $X=1.395 $Y=1.765 $X2=0
+ $Y2=0
cc_153 N_A_81_296#_c_132_n N_VPWR_c_445_n 0.00658808f $X=1.845 $Y=1.765 $X2=0
+ $Y2=0
cc_154 N_A_81_296#_c_120_n N_VPWR_c_445_n 0.00279228f $X=2.475 $Y=1.195 $X2=0
+ $Y2=0
cc_155 N_A_81_296#_c_125_n N_VPWR_c_445_n 0.00923179f $X=2.06 $Y=1.195 $X2=0
+ $Y2=0
cc_156 N_A_81_296#_c_129_n N_VPWR_c_448_n 0.00413917f $X=0.495 $Y=1.765 $X2=0
+ $Y2=0
cc_157 N_A_81_296#_c_130_n N_VPWR_c_448_n 0.00413917f $X=0.945 $Y=1.765 $X2=0
+ $Y2=0
cc_158 N_A_81_296#_c_131_n N_VPWR_c_450_n 0.00445602f $X=1.395 $Y=1.765 $X2=0
+ $Y2=0
cc_159 N_A_81_296#_c_132_n N_VPWR_c_450_n 0.00445602f $X=1.845 $Y=1.765 $X2=0
+ $Y2=0
cc_160 N_A_81_296#_c_129_n N_VPWR_c_441_n 0.00817726f $X=0.495 $Y=1.765 $X2=0
+ $Y2=0
cc_161 N_A_81_296#_c_130_n N_VPWR_c_441_n 0.00817726f $X=0.945 $Y=1.765 $X2=0
+ $Y2=0
cc_162 N_A_81_296#_c_131_n N_VPWR_c_441_n 0.00857589f $X=1.395 $Y=1.765 $X2=0
+ $Y2=0
cc_163 N_A_81_296#_c_132_n N_VPWR_c_441_n 0.00858305f $X=1.845 $Y=1.765 $X2=0
+ $Y2=0
cc_164 N_A_81_296#_M1008_g N_X_c_521_n 0.00760419f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_165 N_A_81_296#_M1011_g N_X_c_521_n 3.97481e-19 $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_166 N_A_81_296#_M1008_g N_X_c_522_n 0.0127847f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_167 N_A_81_296#_M1011_g N_X_c_522_n 0.00591885f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_168 N_A_81_296#_c_119_n N_X_c_522_n 0.00968248f $X=1.975 $Y=1.465 $X2=0 $Y2=0
cc_169 N_A_81_296#_M1008_g N_X_c_523_n 0.00168928f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_170 N_A_81_296#_c_129_n N_X_c_523_n 8.41678e-19 $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_171 N_A_81_296#_c_114_n N_X_c_523_n 0.0167821f $X=0.85 $Y=1.555 $X2=0 $Y2=0
cc_172 N_A_81_296#_c_130_n N_X_c_523_n 7.79736e-19 $X=0.945 $Y=1.765 $X2=0 $Y2=0
cc_173 N_A_81_296#_c_118_n N_X_c_523_n 0.00337535f $X=0.495 $Y=1.555 $X2=0 $Y2=0
cc_174 N_A_81_296#_c_119_n N_X_c_523_n 0.0169058f $X=1.975 $Y=1.465 $X2=0 $Y2=0
cc_175 N_A_81_296#_c_128_n N_X_c_523_n 0.0037137f $X=1.845 $Y=1.532 $X2=0 $Y2=0
cc_176 N_A_81_296#_c_129_n N_X_c_528_n 3.83425e-19 $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_177 N_A_81_296#_c_130_n N_X_c_528_n 0.00454228f $X=0.945 $Y=1.765 $X2=0 $Y2=0
cc_178 N_A_81_296#_M1011_g N_X_c_524_n 0.0142725f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_179 N_A_81_296#_M1014_g N_X_c_524_n 0.0124749f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_180 N_A_81_296#_c_119_n N_X_c_524_n 0.066849f $X=1.975 $Y=1.465 $X2=0 $Y2=0
cc_181 N_A_81_296#_c_121_n N_X_c_524_n 0.00420057f $X=2.64 $Y=0.515 $X2=0 $Y2=0
cc_182 N_A_81_296#_c_125_n N_X_c_524_n 0.00159809f $X=2.06 $Y=1.195 $X2=0 $Y2=0
cc_183 N_A_81_296#_c_128_n N_X_c_524_n 0.00672345f $X=1.845 $Y=1.532 $X2=0 $Y2=0
cc_184 N_A_81_296#_c_114_n N_X_c_529_n 0.00153296f $X=0.85 $Y=1.555 $X2=0 $Y2=0
cc_185 N_A_81_296#_c_130_n N_X_c_529_n 0.0141989f $X=0.945 $Y=1.765 $X2=0 $Y2=0
cc_186 N_A_81_296#_c_131_n N_X_c_529_n 0.0128953f $X=1.395 $Y=1.765 $X2=0 $Y2=0
cc_187 N_A_81_296#_c_132_n N_X_c_529_n 0.00388538f $X=1.845 $Y=1.765 $X2=0 $Y2=0
cc_188 N_A_81_296#_c_119_n N_X_c_529_n 0.0652037f $X=1.975 $Y=1.465 $X2=0 $Y2=0
cc_189 N_A_81_296#_c_128_n N_X_c_529_n 0.015756f $X=1.845 $Y=1.532 $X2=0 $Y2=0
cc_190 N_A_81_296#_c_130_n N_X_c_530_n 7.68526e-19 $X=0.945 $Y=1.765 $X2=0 $Y2=0
cc_191 N_A_81_296#_c_131_n N_X_c_530_n 0.012705f $X=1.395 $Y=1.765 $X2=0 $Y2=0
cc_192 N_A_81_296#_c_132_n N_X_c_530_n 0.0113906f $X=1.845 $Y=1.765 $X2=0 $Y2=0
cc_193 N_A_81_296#_M1011_g N_X_c_525_n 9.72214e-19 $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_194 N_A_81_296#_M1014_g N_X_c_525_n 0.00910117f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_195 N_A_81_296#_M1015_g N_X_c_525_n 4.71232e-19 $X=1.88 $Y=0.74 $X2=0 $Y2=0
cc_196 N_A_81_296#_M1008_g N_X_c_526_n 0.0182661f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_197 N_A_81_296#_c_118_n N_X_c_526_n 4.20821e-19 $X=0.495 $Y=1.555 $X2=0 $Y2=0
cc_198 N_A_81_296#_c_129_n N_X_c_531_n 8.24092e-19 $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_199 N_A_81_296#_c_114_n N_X_c_531_n 0.00102339f $X=0.85 $Y=1.555 $X2=0 $Y2=0
cc_200 N_A_81_296#_c_120_n N_A_489_392#_c_594_n 0.00136603f $X=2.475 $Y=1.195
+ $X2=0 $Y2=0
cc_201 N_A_81_296#_c_126_n N_A_489_392#_c_594_n 0.00178483f $X=2.64 $Y=1.195
+ $X2=0 $Y2=0
cc_202 N_A_81_296#_c_122_n N_A_489_392#_c_596_n 0.00530457f $X=3.505 $Y=1.195
+ $X2=0 $Y2=0
cc_203 N_A_81_296#_c_122_n N_A_489_392#_c_597_n 0.00237093f $X=3.505 $Y=1.195
+ $X2=0 $Y2=0
cc_204 N_A_81_296#_c_124_n N_A_489_392#_c_597_n 0.0144861f $X=4.04 $Y=2.08 $X2=0
+ $Y2=0
cc_205 N_A_81_296#_c_127_n N_A_489_392#_c_597_n 0.00708319f $X=3.63 $Y=1.28
+ $X2=0 $Y2=0
cc_206 N_A_81_296#_c_124_n N_A_489_392#_c_598_n 0.0403584f $X=4.04 $Y=2.08 $X2=0
+ $Y2=0
cc_207 N_A_81_296#_M1001_d N_A_489_392#_c_599_n 0.00222494f $X=3.89 $Y=1.935
+ $X2=0 $Y2=0
cc_208 N_A_81_296#_c_124_n N_A_489_392#_c_599_n 0.0144323f $X=4.04 $Y=2.08 $X2=0
+ $Y2=0
cc_209 N_A_81_296#_c_124_n N_A_489_392#_c_601_n 0.0529704f $X=4.04 $Y=2.08 $X2=0
+ $Y2=0
cc_210 N_A_81_296#_c_125_n N_VGND_M1015_d 0.00184398f $X=2.06 $Y=1.195 $X2=0
+ $Y2=0
cc_211 N_A_81_296#_M1008_g N_VGND_c_648_n 0.00351842f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_212 N_A_81_296#_M1008_g N_VGND_c_649_n 4.94543e-19 $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_213 N_A_81_296#_M1011_g N_VGND_c_649_n 0.00916944f $X=0.925 $Y=0.74 $X2=0
+ $Y2=0
cc_214 N_A_81_296#_M1014_g N_VGND_c_649_n 0.00393745f $X=1.425 $Y=0.74 $X2=0
+ $Y2=0
cc_215 N_A_81_296#_M1015_g N_VGND_c_650_n 0.00193131f $X=1.88 $Y=0.74 $X2=0
+ $Y2=0
cc_216 N_A_81_296#_c_120_n N_VGND_c_650_n 0.0103909f $X=2.475 $Y=1.195 $X2=0
+ $Y2=0
cc_217 N_A_81_296#_c_121_n N_VGND_c_650_n 0.0229287f $X=2.64 $Y=0.515 $X2=0
+ $Y2=0
cc_218 N_A_81_296#_c_125_n N_VGND_c_650_n 0.0132288f $X=2.06 $Y=1.195 $X2=0
+ $Y2=0
cc_219 N_A_81_296#_c_121_n N_VGND_c_651_n 0.0404434f $X=2.64 $Y=0.515 $X2=0
+ $Y2=0
cc_220 N_A_81_296#_c_122_n N_VGND_c_651_n 0.0238718f $X=3.505 $Y=1.195 $X2=0
+ $Y2=0
cc_221 N_A_81_296#_c_123_n N_VGND_c_651_n 0.0220066f $X=3.67 $Y=0.515 $X2=0
+ $Y2=0
cc_222 N_A_81_296#_c_123_n N_VGND_c_652_n 0.025828f $X=3.67 $Y=0.515 $X2=0 $Y2=0
cc_223 N_A_81_296#_c_127_n N_VGND_c_652_n 0.0132716f $X=3.63 $Y=1.28 $X2=0 $Y2=0
cc_224 N_A_81_296#_M1008_g N_VGND_c_653_n 0.00434272f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_225 N_A_81_296#_M1011_g N_VGND_c_653_n 0.00383152f $X=0.925 $Y=0.74 $X2=0
+ $Y2=0
cc_226 N_A_81_296#_M1014_g N_VGND_c_654_n 0.00434272f $X=1.425 $Y=0.74 $X2=0
+ $Y2=0
cc_227 N_A_81_296#_M1015_g N_VGND_c_654_n 0.00461464f $X=1.88 $Y=0.74 $X2=0
+ $Y2=0
cc_228 N_A_81_296#_c_121_n N_VGND_c_655_n 0.0146357f $X=2.64 $Y=0.515 $X2=0
+ $Y2=0
cc_229 N_A_81_296#_c_123_n N_VGND_c_656_n 0.0109942f $X=3.67 $Y=0.515 $X2=0
+ $Y2=0
cc_230 N_A_81_296#_M1008_g N_VGND_c_658_n 0.00823942f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_231 N_A_81_296#_M1011_g N_VGND_c_658_n 0.0075754f $X=0.925 $Y=0.74 $X2=0
+ $Y2=0
cc_232 N_A_81_296#_M1014_g N_VGND_c_658_n 0.00820964f $X=1.425 $Y=0.74 $X2=0
+ $Y2=0
cc_233 N_A_81_296#_M1015_g N_VGND_c_658_n 0.00908295f $X=1.88 $Y=0.74 $X2=0
+ $Y2=0
cc_234 N_A_81_296#_c_121_n N_VGND_c_658_n 0.0121141f $X=2.64 $Y=0.515 $X2=0
+ $Y2=0
cc_235 N_A_81_296#_c_123_n N_VGND_c_658_n 0.00904371f $X=3.67 $Y=0.515 $X2=0
+ $Y2=0
cc_236 N_A_M1010_g N_A_676_48#_M1009_g 0.0160624f $X=2.955 $Y=0.69 $X2=0 $Y2=0
cc_237 N_A_c_262_n N_A_676_48#_c_320_n 0.0160624f $X=2.82 $Y=1.885 $X2=0 $Y2=0
cc_238 A N_A_676_48#_c_320_n 0.00232169f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_239 N_A_c_262_n N_A_676_48#_c_321_n 0.0019669f $X=2.82 $Y=1.885 $X2=0 $Y2=0
cc_240 A N_A_676_48#_c_321_n 0.00179353f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_241 N_A_c_267_n N_VPWR_c_445_n 0.0122091f $X=2.37 $Y=1.885 $X2=0 $Y2=0
cc_242 N_A_c_262_n N_VPWR_c_446_n 0.00714506f $X=2.82 $Y=1.885 $X2=0 $Y2=0
cc_243 N_A_c_267_n N_VPWR_c_452_n 0.00445602f $X=2.37 $Y=1.885 $X2=0 $Y2=0
cc_244 N_A_c_262_n N_VPWR_c_452_n 0.00445602f $X=2.82 $Y=1.885 $X2=0 $Y2=0
cc_245 N_A_c_267_n N_VPWR_c_441_n 0.00858193f $X=2.37 $Y=1.885 $X2=0 $Y2=0
cc_246 N_A_c_262_n N_VPWR_c_441_n 0.00862391f $X=2.82 $Y=1.885 $X2=0 $Y2=0
cc_247 N_A_M1004_g N_X_c_524_n 2.21979e-19 $X=2.355 $Y=0.69 $X2=0 $Y2=0
cc_248 N_A_c_267_n N_X_c_529_n 6.537e-19 $X=2.37 $Y=1.885 $X2=0 $Y2=0
cc_249 N_A_c_267_n N_A_489_392#_c_594_n 0.00289977f $X=2.37 $Y=1.885 $X2=0 $Y2=0
cc_250 N_A_c_261_n N_A_489_392#_c_594_n 3.09627e-19 $X=2.7 $Y=1.515 $X2=0 $Y2=0
cc_251 N_A_c_262_n N_A_489_392#_c_594_n 0.00168072f $X=2.82 $Y=1.885 $X2=0 $Y2=0
cc_252 A N_A_489_392#_c_594_n 0.0204727f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_253 N_A_c_267_n N_A_489_392#_c_595_n 0.00910879f $X=2.37 $Y=1.885 $X2=0 $Y2=0
cc_254 N_A_c_262_n N_A_489_392#_c_595_n 0.0114329f $X=2.82 $Y=1.885 $X2=0 $Y2=0
cc_255 N_A_c_262_n N_A_489_392#_c_596_n 0.0175384f $X=2.82 $Y=1.885 $X2=0 $Y2=0
cc_256 A N_A_489_392#_c_596_n 0.0360063f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_257 N_A_c_262_n N_A_489_392#_c_597_n 8.62857e-19 $X=2.82 $Y=1.885 $X2=0 $Y2=0
cc_258 N_A_c_262_n N_A_489_392#_c_598_n 0.00327785f $X=2.82 $Y=1.885 $X2=0 $Y2=0
cc_259 N_A_M1004_g N_VGND_c_650_n 0.0107172f $X=2.355 $Y=0.69 $X2=0 $Y2=0
cc_260 N_A_M1010_g N_VGND_c_650_n 6.11496e-19 $X=2.955 $Y=0.69 $X2=0 $Y2=0
cc_261 N_A_M1004_g N_VGND_c_651_n 6.29519e-19 $X=2.355 $Y=0.69 $X2=0 $Y2=0
cc_262 N_A_M1010_g N_VGND_c_651_n 0.0112125f $X=2.955 $Y=0.69 $X2=0 $Y2=0
cc_263 N_A_M1004_g N_VGND_c_655_n 0.00383152f $X=2.355 $Y=0.69 $X2=0 $Y2=0
cc_264 N_A_M1010_g N_VGND_c_655_n 0.00383152f $X=2.955 $Y=0.69 $X2=0 $Y2=0
cc_265 N_A_M1004_g N_VGND_c_658_n 0.00758997f $X=2.355 $Y=0.69 $X2=0 $Y2=0
cc_266 N_A_M1010_g N_VGND_c_658_n 0.00758997f $X=2.955 $Y=0.69 $X2=0 $Y2=0
cc_267 N_A_676_48#_M1017_g N_B_N_c_405_n 0.0196085f $X=3.885 $Y=0.69 $X2=-0.19
+ $Y2=-0.245
cc_268 N_A_676_48#_c_326_n N_B_N_c_405_n 0.00686389f $X=4.53 $Y=0.95 $X2=-0.19
+ $Y2=-0.245
cc_269 N_A_676_48#_c_330_n N_B_N_c_405_n 0.00308772f $X=4.46 $Y=1.445 $X2=-0.19
+ $Y2=-0.245
cc_270 N_A_676_48#_c_327_n N_B_N_c_406_n 0.0253584f $X=5.405 $Y=0.65 $X2=0 $Y2=0
cc_271 N_A_676_48#_c_328_n N_B_N_c_406_n 0.0196942f $X=5.49 $Y=2.105 $X2=0 $Y2=0
cc_272 N_A_676_48#_c_330_n N_B_N_c_406_n 0.0113271f $X=4.46 $Y=1.445 $X2=0 $Y2=0
cc_273 N_A_676_48#_c_324_n N_B_N_c_407_n 0.0206227f $X=4.265 $Y=1.86 $X2=0 $Y2=0
cc_274 N_A_676_48#_c_329_n N_B_N_c_407_n 9.63591e-19 $X=4.46 $Y=1.61 $X2=0 $Y2=0
cc_275 N_A_676_48#_c_330_n N_B_N_c_407_n 0.00296893f $X=4.46 $Y=1.445 $X2=0
+ $Y2=0
cc_276 N_A_676_48#_c_324_n N_B_N_c_408_n 3.70002e-19 $X=4.265 $Y=1.86 $X2=0
+ $Y2=0
cc_277 N_A_676_48#_c_328_n N_B_N_c_408_n 0.0107489f $X=5.49 $Y=2.105 $X2=0 $Y2=0
cc_278 N_A_676_48#_c_324_n B_N 0.00149938f $X=4.265 $Y=1.86 $X2=0 $Y2=0
cc_279 N_A_676_48#_c_327_n B_N 0.0282282f $X=5.405 $Y=0.65 $X2=0 $Y2=0
cc_280 N_A_676_48#_c_328_n B_N 0.0517945f $X=5.49 $Y=2.105 $X2=0 $Y2=0
cc_281 N_A_676_48#_c_330_n B_N 0.0330704f $X=4.46 $Y=1.445 $X2=0 $Y2=0
cc_282 N_A_676_48#_c_324_n N_B_N_c_409_n 0.0149629f $X=4.265 $Y=1.86 $X2=0 $Y2=0
cc_283 N_A_676_48#_c_329_n N_B_N_c_409_n 0.00134012f $X=4.46 $Y=1.61 $X2=0 $Y2=0
cc_284 N_A_676_48#_c_330_n N_B_N_c_409_n 0.0045702f $X=4.46 $Y=1.445 $X2=0 $Y2=0
cc_285 N_A_676_48#_c_332_n N_VPWR_c_446_n 5.31157e-19 $X=3.815 $Y=1.86 $X2=0
+ $Y2=0
cc_286 N_A_676_48#_c_324_n N_VPWR_c_447_n 0.00212399f $X=4.265 $Y=1.86 $X2=0
+ $Y2=0
cc_287 N_A_676_48#_c_328_n N_VPWR_c_447_n 0.0684217f $X=5.49 $Y=2.105 $X2=0
+ $Y2=0
cc_288 N_A_676_48#_c_332_n N_VPWR_c_453_n 9.44495e-19 $X=3.815 $Y=1.86 $X2=0
+ $Y2=0
cc_289 N_A_676_48#_c_324_n N_VPWR_c_453_n 9.63649e-19 $X=4.265 $Y=1.86 $X2=0
+ $Y2=0
cc_290 N_A_676_48#_c_328_n N_VPWR_c_454_n 0.011066f $X=5.49 $Y=2.105 $X2=0 $Y2=0
cc_291 N_A_676_48#_c_328_n N_VPWR_c_441_n 0.00915947f $X=5.49 $Y=2.105 $X2=0
+ $Y2=0
cc_292 N_A_676_48#_c_320_n N_A_489_392#_c_596_n 0.00111948f $X=3.53 $Y=1.52
+ $X2=0 $Y2=0
cc_293 N_A_676_48#_c_320_n N_A_489_392#_c_597_n 0.00633348f $X=3.53 $Y=1.52
+ $X2=0 $Y2=0
cc_294 N_A_676_48#_c_332_n N_A_489_392#_c_597_n 0.00124547f $X=3.815 $Y=1.86
+ $X2=0 $Y2=0
cc_295 N_A_676_48#_c_332_n N_A_489_392#_c_599_n 0.0151379f $X=3.815 $Y=1.86
+ $X2=0 $Y2=0
cc_296 N_A_676_48#_c_324_n N_A_489_392#_c_599_n 0.0148754f $X=4.265 $Y=1.86
+ $X2=0 $Y2=0
cc_297 N_A_676_48#_c_332_n N_A_489_392#_c_601_n 7.35453e-19 $X=3.815 $Y=1.86
+ $X2=0 $Y2=0
cc_298 N_A_676_48#_c_324_n N_A_489_392#_c_601_n 0.0133693f $X=4.265 $Y=1.86
+ $X2=0 $Y2=0
cc_299 N_A_676_48#_c_329_n N_A_489_392#_c_601_n 0.0229155f $X=4.46 $Y=1.61 $X2=0
+ $Y2=0
cc_300 N_A_676_48#_M1009_g N_VGND_c_651_n 0.00476029f $X=3.455 $Y=0.69 $X2=0
+ $Y2=0
cc_301 N_A_676_48#_M1009_g N_VGND_c_652_n 5.56357e-19 $X=3.455 $Y=0.69 $X2=0
+ $Y2=0
cc_302 N_A_676_48#_M1017_g N_VGND_c_652_n 0.0117552f $X=3.885 $Y=0.69 $X2=0
+ $Y2=0
cc_303 N_A_676_48#_c_323_n N_VGND_c_652_n 0.00602973f $X=4.175 $Y=1.52 $X2=0
+ $Y2=0
cc_304 N_A_676_48#_c_326_n N_VGND_c_652_n 0.0260683f $X=4.53 $Y=0.95 $X2=0 $Y2=0
cc_305 N_A_676_48#_c_330_n N_VGND_c_652_n 0.00351404f $X=4.46 $Y=1.445 $X2=0
+ $Y2=0
cc_306 N_A_676_48#_M1009_g N_VGND_c_656_n 0.00434272f $X=3.455 $Y=0.69 $X2=0
+ $Y2=0
cc_307 N_A_676_48#_M1017_g N_VGND_c_656_n 0.00383152f $X=3.885 $Y=0.69 $X2=0
+ $Y2=0
cc_308 N_A_676_48#_c_326_n N_VGND_c_657_n 0.00840325f $X=4.53 $Y=0.95 $X2=0
+ $Y2=0
cc_309 N_A_676_48#_c_327_n N_VGND_c_657_n 0.0454555f $X=5.405 $Y=0.65 $X2=0
+ $Y2=0
cc_310 N_A_676_48#_M1009_g N_VGND_c_658_n 0.00820772f $X=3.455 $Y=0.69 $X2=0
+ $Y2=0
cc_311 N_A_676_48#_M1017_g N_VGND_c_658_n 0.0075754f $X=3.885 $Y=0.69 $X2=0
+ $Y2=0
cc_312 N_A_676_48#_c_326_n N_VGND_c_658_n 0.00689675f $X=4.53 $Y=0.95 $X2=0
+ $Y2=0
cc_313 N_A_676_48#_c_327_n N_VGND_c_658_n 0.037886f $X=5.405 $Y=0.65 $X2=0 $Y2=0
cc_314 N_B_N_c_410_n N_VPWR_c_447_n 0.0186373f $X=5.265 $Y=1.885 $X2=0 $Y2=0
cc_315 N_B_N_c_408_n N_VPWR_c_447_n 0.00197705f $X=5.115 $Y=1.58 $X2=0 $Y2=0
cc_316 B_N N_VPWR_c_447_n 0.0233678f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_317 N_B_N_c_410_n N_VPWR_c_454_n 0.00413917f $X=5.265 $Y=1.885 $X2=0 $Y2=0
cc_318 N_B_N_c_410_n N_VPWR_c_441_n 0.00821187f $X=5.265 $Y=1.885 $X2=0 $Y2=0
cc_319 N_B_N_c_410_n N_A_489_392#_c_599_n 5.9004e-19 $X=5.265 $Y=1.885 $X2=0
+ $Y2=0
cc_320 N_B_N_c_410_n N_A_489_392#_c_601_n 3.68457e-19 $X=5.265 $Y=1.885 $X2=0
+ $Y2=0
cc_321 N_B_N_c_405_n N_VGND_c_652_n 0.00676331f $X=4.385 $Y=1.085 $X2=0 $Y2=0
cc_322 N_B_N_c_405_n N_VGND_c_657_n 0.00433139f $X=4.385 $Y=1.085 $X2=0 $Y2=0
cc_323 N_B_N_c_405_n N_VGND_c_658_n 0.00822102f $X=4.385 $Y=1.085 $X2=0 $Y2=0
cc_324 N_VPWR_c_443_n N_X_c_528_n 0.0386303f $X=0.27 $Y=1.985 $X2=0 $Y2=0
cc_325 N_VPWR_c_444_n N_X_c_528_n 0.0542575f $X=1.17 $Y=2.305 $X2=0 $Y2=0
cc_326 N_VPWR_c_448_n N_X_c_528_n 0.00883494f $X=1.005 $Y=3.33 $X2=0 $Y2=0
cc_327 N_VPWR_c_441_n N_X_c_528_n 0.0073128f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_328 N_VPWR_M1003_s N_X_c_529_n 0.00222494f $X=1.02 $Y=1.84 $X2=0 $Y2=0
cc_329 N_VPWR_c_444_n N_X_c_529_n 0.0154248f $X=1.17 $Y=2.305 $X2=0 $Y2=0
cc_330 N_VPWR_c_445_n N_X_c_529_n 0.00213573f $X=2.07 $Y=2.105 $X2=0 $Y2=0
cc_331 N_VPWR_c_444_n N_X_c_530_n 0.0563525f $X=1.17 $Y=2.305 $X2=0 $Y2=0
cc_332 N_VPWR_c_445_n N_X_c_530_n 0.0677182f $X=2.07 $Y=2.105 $X2=0 $Y2=0
cc_333 N_VPWR_c_450_n N_X_c_530_n 0.014552f $X=1.985 $Y=3.33 $X2=0 $Y2=0
cc_334 N_VPWR_c_441_n N_X_c_530_n 0.0119791f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_335 N_VPWR_c_443_n N_X_c_526_n 0.0143443f $X=0.27 $Y=1.985 $X2=0 $Y2=0
cc_336 N_VPWR_c_443_n N_X_c_531_n 0.00654085f $X=0.27 $Y=1.985 $X2=0 $Y2=0
cc_337 N_VPWR_c_445_n N_A_489_392#_c_594_n 0.0123566f $X=2.07 $Y=2.105 $X2=0
+ $Y2=0
cc_338 N_VPWR_c_445_n N_A_489_392#_c_595_n 0.0587921f $X=2.07 $Y=2.105 $X2=0
+ $Y2=0
cc_339 N_VPWR_c_446_n N_A_489_392#_c_595_n 0.0462948f $X=3.045 $Y=2.455 $X2=0
+ $Y2=0
cc_340 N_VPWR_c_452_n N_A_489_392#_c_595_n 0.014552f $X=2.96 $Y=3.33 $X2=0 $Y2=0
cc_341 N_VPWR_c_441_n N_A_489_392#_c_595_n 0.0119791f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_342 N_VPWR_M1007_s N_A_489_392#_c_596_n 0.00359549f $X=2.895 $Y=1.96 $X2=0
+ $Y2=0
cc_343 N_VPWR_c_446_n N_A_489_392#_c_596_n 0.0202669f $X=3.045 $Y=2.455 $X2=0
+ $Y2=0
cc_344 N_VPWR_c_446_n N_A_489_392#_c_598_n 0.0416236f $X=3.045 $Y=2.455 $X2=0
+ $Y2=0
cc_345 N_VPWR_c_447_n N_A_489_392#_c_599_n 0.0125437f $X=5.04 $Y=2.125 $X2=0
+ $Y2=0
cc_346 N_VPWR_c_453_n N_A_489_392#_c_599_n 0.0654702f $X=4.875 $Y=3.33 $X2=0
+ $Y2=0
cc_347 N_VPWR_c_441_n N_A_489_392#_c_599_n 0.0372602f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_348 N_VPWR_c_446_n N_A_489_392#_c_600_n 0.0124983f $X=3.045 $Y=2.455 $X2=0
+ $Y2=0
cc_349 N_VPWR_c_453_n N_A_489_392#_c_600_n 0.0179217f $X=4.875 $Y=3.33 $X2=0
+ $Y2=0
cc_350 N_VPWR_c_441_n N_A_489_392#_c_600_n 0.00971942f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_351 N_VPWR_c_447_n N_A_489_392#_c_601_n 0.0656672f $X=5.04 $Y=2.125 $X2=0
+ $Y2=0
cc_352 N_X_c_524_n N_VGND_M1011_d 0.00266f $X=1.475 $Y=1.045 $X2=0 $Y2=0
cc_353 N_X_c_521_n N_VGND_c_648_n 0.0216462f $X=0.71 $Y=0.515 $X2=0 $Y2=0
cc_354 N_X_c_526_n N_VGND_c_648_n 0.0201602f $X=0.545 $Y=1.295 $X2=0 $Y2=0
cc_355 N_X_c_521_n N_VGND_c_649_n 0.0156021f $X=0.71 $Y=0.515 $X2=0 $Y2=0
cc_356 N_X_c_524_n N_VGND_c_649_n 0.018932f $X=1.475 $Y=1.045 $X2=0 $Y2=0
cc_357 N_X_c_525_n N_VGND_c_649_n 0.0163623f $X=1.64 $Y=0.515 $X2=0 $Y2=0
cc_358 N_X_c_525_n N_VGND_c_650_n 0.022799f $X=1.64 $Y=0.515 $X2=0 $Y2=0
cc_359 N_X_c_521_n N_VGND_c_653_n 0.0109942f $X=0.71 $Y=0.515 $X2=0 $Y2=0
cc_360 N_X_c_525_n N_VGND_c_654_n 0.0145639f $X=1.64 $Y=0.515 $X2=0 $Y2=0
cc_361 N_X_c_521_n N_VGND_c_658_n 0.00904371f $X=0.71 $Y=0.515 $X2=0 $Y2=0
cc_362 N_X_c_525_n N_VGND_c_658_n 0.0119984f $X=1.64 $Y=0.515 $X2=0 $Y2=0
