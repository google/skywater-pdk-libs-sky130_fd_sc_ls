* File: sky130_fd_sc_ls__mux2i_1.pex.spice
* Created: Wed Sep  2 11:10:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__MUX2I_1%S 3 5 7 8 11 12 14 15 17 19 20 21 22 23 27
c64 15 0 1.0697e-19 $X=1.485 $Y=1.185
c65 5 0 8.19203e-20 $X=0.495 $Y=2.045
r66 27 28 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.385
+ $Y=1.35 $X2=0.385 $Y2=1.35
r67 23 28 8.54164 $w=4.23e-07 $l=3.15e-07 $layer=LI1_cond $X=0.337 $Y=1.665
+ $X2=0.337 $Y2=1.35
r68 22 28 1.4914 $w=4.23e-07 $l=5.5e-08 $layer=LI1_cond $X=0.337 $Y=1.295
+ $X2=0.337 $Y2=1.35
r69 20 27 54.4068 $w=3.5e-07 $l=3.3e-07 $layer=POLY_cond $X=0.395 $Y=1.68
+ $X2=0.395 $Y2=1.35
r70 18 27 2.47304 $w=3.5e-07 $l=1.5e-08 $layer=POLY_cond $X=0.395 $Y=1.335
+ $X2=0.395 $Y2=1.35
r71 18 19 13.0992 $w=2.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.395 $Y=1.335
+ $X2=0.395 $Y2=1.26
r72 15 21 18.8402 $w=1.65e-07 $l=8.21584e-08 $layer=POLY_cond $X=1.485 $Y=1.185
+ $X2=1.47 $Y2=1.26
r73 15 17 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.485 $Y=1.185
+ $X2=1.485 $Y2=0.74
r74 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.47 $Y=1.765
+ $X2=1.47 $Y2=2.4
r75 11 12 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.47 $Y=1.675 $X2=1.47
+ $Y2=1.765
r76 10 21 18.8402 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=1.47 $Y=1.335
+ $X2=1.47 $Y2=1.26
r77 10 11 132.161 $w=1.8e-07 $l=3.4e-07 $layer=POLY_cond $X=1.47 $Y=1.335
+ $X2=1.47 $Y2=1.675
r78 9 19 12.7694 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=0.57 $Y=1.26
+ $X2=0.395 $Y2=1.26
r79 8 21 6.66866 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=1.38 $Y=1.26 $X2=1.47
+ $Y2=1.26
r80 8 9 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=1.38 $Y=1.26 $X2=0.57
+ $Y2=1.26
r81 5 20 67.4061 $w=2.61e-07 $l=4.11977e-07 $layer=POLY_cond $X=0.495 $Y=2.045
+ $X2=0.395 $Y2=1.68
r82 5 7 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.495 $Y=2.045
+ $X2=0.495 $Y2=2.54
r83 1 19 13.0992 $w=2.5e-07 $l=1.32288e-07 $layer=POLY_cond $X=0.495 $Y=1.185
+ $X2=0.395 $Y2=1.26
r84 1 3 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=0.495 $Y=1.185
+ $X2=0.495 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_LS__MUX2I_1%A_114_74# 1 2 7 9 12 17 20 23 27 28 29 30
c71 17 0 1.0697e-19 $X=0.805 $Y=1.35
r72 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.965
+ $Y=1.515 $X2=1.965 $Y2=1.515
r73 30 33 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=1.965 $Y=1.435
+ $X2=1.965 $Y2=1.515
r74 27 28 8.46614 $w=3.33e-07 $l=1.65e-07 $layer=LI1_cond $X=0.722 $Y=2.265
+ $X2=0.722 $Y2=2.1
r75 23 25 11.6528 $w=3.43e-07 $l=2.6e-07 $layer=LI1_cond $X=0.717 $Y=0.645
+ $X2=0.717 $Y2=0.905
r76 21 29 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.89 $Y=1.435
+ $X2=0.805 $Y2=1.435
r77 20 30 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.8 $Y=1.435
+ $X2=1.965 $Y2=1.435
r78 20 21 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=1.8 $Y=1.435 $X2=0.89
+ $Y2=1.435
r79 18 29 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.805 $Y=1.52
+ $X2=0.805 $Y2=1.435
r80 18 28 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=0.805 $Y=1.52
+ $X2=0.805 $Y2=2.1
r81 17 29 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.805 $Y=1.35
+ $X2=0.805 $Y2=1.435
r82 17 25 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=0.805 $Y=1.35
+ $X2=0.805 $Y2=0.905
r83 10 34 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=2.055 $Y=1.35
+ $X2=1.965 $Y2=1.515
r84 10 12 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.055 $Y=1.35
+ $X2=2.055 $Y2=0.74
r85 7 34 52.2586 $w=2.99e-07 $l=2.7157e-07 $layer=POLY_cond $X=1.92 $Y=1.765
+ $X2=1.965 $Y2=1.515
r86 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.92 $Y=1.765
+ $X2=1.92 $Y2=2.4
r87 2 27 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=0.57
+ $Y=2.12 $X2=0.72 $Y2=2.265
r88 1 23 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_LS__MUX2I_1%A0 3 5 7 8 12 13
r34 12 14 31.861 $w=2.95e-07 $l=1.95e-07 $layer=POLY_cond $X=2.7 $Y=1.557
+ $X2=2.895 $Y2=1.557
r35 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.7
+ $Y=1.515 $X2=2.7 $Y2=1.515
r36 8 13 5.08431 $w=3.38e-07 $l=1.5e-07 $layer=LI1_cond $X=2.695 $Y=1.665
+ $X2=2.695 $Y2=1.515
r37 5 14 18.5736 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.895 $Y=1.765
+ $X2=2.895 $Y2=1.557
r38 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.895 $Y=1.765
+ $X2=2.895 $Y2=2.4
r39 1 12 41.6644 $w=2.95e-07 $l=3.43235e-07 $layer=POLY_cond $X=2.445 $Y=1.35
+ $X2=2.7 $Y2=1.557
r40 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.445 $Y=1.35
+ $X2=2.445 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__MUX2I_1%A1 1 3 4 6 7
r20 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.56
+ $Y=1.385 $X2=3.56 $Y2=1.385
r21 7 11 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=3.56 $Y=1.295 $X2=3.56
+ $Y2=1.385
r22 4 10 66.8857 $w=3.73e-07 $l=4.40227e-07 $layer=POLY_cond $X=3.345 $Y=1.765
+ $X2=3.475 $Y2=1.385
r23 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.345 $Y=1.765
+ $X2=3.345 $Y2=2.4
r24 1 10 39.1028 $w=3.73e-07 $l=2.43926e-07 $layer=POLY_cond $X=3.3 $Y=1.22
+ $X2=3.475 $Y2=1.385
r25 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.3 $Y=1.22 $X2=3.3
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__MUX2I_1%VPWR 1 2 7 9 13 15 17 27 28 34
r37 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r38 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r39 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r40 25 28 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.6 $Y2=3.33
r41 24 27 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=3.6 $Y2=3.33
r42 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r43 22 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.86 $Y=3.33
+ $X2=1.695 $Y2=3.33
r44 22 24 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.86 $Y=3.33 $X2=2.16
+ $Y2=3.33
r45 21 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r46 21 32 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.24 $Y2=3.33
r47 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r48 18 31 4.02368 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=0.355 $Y=3.33
+ $X2=0.177 $Y2=3.33
r49 18 20 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=0.355 $Y=3.33
+ $X2=1.2 $Y2=3.33
r50 17 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.53 $Y=3.33
+ $X2=1.695 $Y2=3.33
r51 17 20 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.53 $Y=3.33 $X2=1.2
+ $Y2=3.33
r52 15 25 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.16 $Y2=3.33
r53 15 35 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r54 11 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.695 $Y=3.245
+ $X2=1.695 $Y2=3.33
r55 11 13 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=1.695 $Y=3.245
+ $X2=1.695 $Y2=2.455
r56 7 31 3.11948 $w=2.5e-07 $l=1.08305e-07 $layer=LI1_cond $X=0.23 $Y=3.245
+ $X2=0.177 $Y2=3.33
r57 7 9 45.1758 $w=2.48e-07 $l=9.8e-07 $layer=LI1_cond $X=0.23 $Y=3.245 $X2=0.23
+ $Y2=2.265
r58 2 13 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=1.545
+ $Y=1.84 $X2=1.695 $Y2=2.455
r59 1 9 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.12 $X2=0.27 $Y2=2.265
.ends

.subckt PM_SKY130_FD_SC_LS__MUX2I_1%A_223_368# 1 2 7 9 11 18
c30 7 0 8.19203e-20 $X=1.205 $Y=2.12
r31 12 16 3.99177 $w=1.7e-07 $l=1.5411e-07 $layer=LI1_cond $X=1.33 $Y=2.035
+ $X2=1.205 $Y2=1.97
r32 11 18 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.505 $Y=2.035
+ $X2=2.67 $Y2=2.035
r33 11 12 76.6578 $w=1.68e-07 $l=1.175e-06 $layer=LI1_cond $X=2.505 $Y=2.035
+ $X2=1.33 $Y2=2.035
r34 7 16 3.1514 $w=2.5e-07 $l=1.5e-07 $layer=LI1_cond $X=1.205 $Y=2.12 $X2=1.205
+ $Y2=1.97
r35 7 9 12.9074 $w=2.48e-07 $l=2.8e-07 $layer=LI1_cond $X=1.205 $Y=2.12
+ $X2=1.205 $Y2=2.4
r36 2 18 300 $w=1.7e-07 $l=3.33729e-07 $layer=licon1_PDIFF $count=2 $X=2.54
+ $Y=1.84 $X2=2.67 $Y2=2.115
r37 1 16 600 $w=1.7e-07 $l=1.99687e-07 $layer=licon1_PDIFF $count=1 $X=1.115
+ $Y=1.84 $X2=1.245 $Y2=1.985
r38 1 9 300 $w=1.7e-07 $l=6.21611e-07 $layer=licon1_PDIFF $count=2 $X=1.115
+ $Y=1.84 $X2=1.245 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__MUX2I_1%A_399_368# 1 2 9 11 12 15
r25 15 18 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=3.57 $Y=1.985
+ $X2=3.57 $Y2=2.815
r26 13 18 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=3.57 $Y=2.905 $X2=3.57
+ $Y2=2.815
r27 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.405 $Y=2.99
+ $X2=3.57 $Y2=2.905
r28 11 12 71.4385 $w=1.68e-07 $l=1.095e-06 $layer=LI1_cond $X=3.405 $Y=2.99
+ $X2=2.31 $Y2=2.99
r29 7 12 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.185 $Y=2.905
+ $X2=2.31 $Y2=2.99
r30 7 9 20.744 $w=2.48e-07 $l=4.5e-07 $layer=LI1_cond $X=2.185 $Y=2.905
+ $X2=2.185 $Y2=2.455
r31 2 18 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=3.42
+ $Y=1.84 $X2=3.57 $Y2=2.815
r32 2 15 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=3.42
+ $Y=1.84 $X2=3.57 $Y2=1.985
r33 1 9 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=1.995
+ $Y=1.84 $X2=2.145 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_LS__MUX2I_1%Y 1 2 7 9 11 14
r21 11 14 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=3.035 $Y=0.87
+ $X2=2.64 $Y2=0.87
r22 11 13 2.73294 $w=3.3e-07 $l=9.5e-08 $layer=LI1_cond $X=3.035 $Y=0.87
+ $X2=3.13 $Y2=0.87
r23 7 13 4.74669 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=3.13 $Y=1.035
+ $X2=3.13 $Y2=0.87
r24 7 9 55.4545 $w=1.88e-07 $l=9.5e-07 $layer=LI1_cond $X=3.13 $Y=1.035 $X2=3.13
+ $Y2=1.985
r25 2 9 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=2.97
+ $Y=1.84 $X2=3.12 $Y2=1.985
r26 1 13 91 $w=1.7e-07 $l=7.75709e-07 $layer=licon1_NDIFF $count=2 $X=2.52
+ $Y=0.37 $X2=3.085 $Y2=0.87
.ends

.subckt PM_SKY130_FD_SC_LS__MUX2I_1%VGND 1 2 7 9 13 15 17 27 28 34
r36 34 35 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r37 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r38 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r39 25 28 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.6
+ $Y2=0
r40 24 27 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.16 $Y=0 $X2=3.6
+ $Y2=0
r41 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r42 22 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.935 $Y=0 $X2=1.77
+ $Y2=0
r43 22 24 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=1.935 $Y=0 $X2=2.16
+ $Y2=0
r44 21 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r45 21 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r46 20 21 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r47 18 31 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=0 $X2=0.182
+ $Y2=0
r48 18 20 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=0 $X2=0.72
+ $Y2=0
r49 17 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.605 $Y=0 $X2=1.77
+ $Y2=0
r50 17 20 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=1.605 $Y=0 $X2=0.72
+ $Y2=0
r51 15 25 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.16
+ $Y2=0
r52 15 35 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r53 11 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.77 $Y=0.085
+ $X2=1.77 $Y2=0
r54 11 13 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=1.77 $Y=0.085
+ $X2=1.77 $Y2=0.675
r55 7 31 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.182 $Y2=0
r56 7 9 25.8147 $w=2.48e-07 $l=5.6e-07 $layer=LI1_cond $X=0.24 $Y=0.085 $X2=0.24
+ $Y2=0.645
r57 2 13 182 $w=1.7e-07 $l=3.96327e-07 $layer=licon1_NDIFF $count=1 $X=1.56
+ $Y=0.37 $X2=1.77 $Y2=0.675
r58 1 9 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_LS__MUX2I_1%A_225_74# 1 2 9 11 12 14 15 16 20
r48 15 20 4.62824 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=3.395 $Y=0.435
+ $X2=3.537 $Y2=0.435
r49 15 16 73.0695 $w=1.68e-07 $l=1.12e-06 $layer=LI1_cond $X=3.395 $Y=0.435
+ $X2=2.275 $Y2=0.435
r50 13 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.19 $Y=0.52
+ $X2=2.275 $Y2=0.435
r51 13 14 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=2.19 $Y=0.52
+ $X2=2.19 $Y2=1.01
r52 11 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.105 $Y=1.095
+ $X2=2.19 $Y2=1.01
r53 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.105 $Y=1.095
+ $X2=1.435 $Y2=1.095
r54 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.27 $Y=1.01
+ $X2=1.435 $Y2=1.095
r55 7 9 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=1.27 $Y=1.01 $X2=1.27
+ $Y2=0.515
r56 2 20 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=3.375
+ $Y=0.37 $X2=3.515 $Y2=0.495
r57 1 9 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=1.125
+ $Y=0.37 $X2=1.27 $Y2=0.515
.ends

