* File: sky130_fd_sc_ls__sdfrtp_2.pex.spice
* Created: Wed Sep  2 11:27:23 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__SDFRTP_2%A_27_74# 1 2 7 9 11 12 14 17 20 23 27 30 32
+ 33 35 40
c80 35 0 9.95498e-21 $X=2.5 $Y=1.995
c81 30 0 2.73032e-20 $X=2.375 $Y=2.09
c82 12 0 1.82457e-19 $X=2.485 $Y=2.245
c83 9 0 3.56444e-20 $X=1.485 $Y=0.935
r84 35 38 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=2.54 $Y=1.995
+ $X2=2.54 $Y2=2.09
r85 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.5
+ $Y=1.995 $X2=2.5 $Y2=1.995
r86 31 33 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.445 $Y=2.09
+ $X2=0.28 $Y2=2.09
r87 30 38 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.375 $Y=2.09
+ $X2=2.54 $Y2=2.09
r88 30 31 125.914 $w=1.68e-07 $l=1.93e-06 $layer=LI1_cond $X=2.375 $Y=2.09
+ $X2=0.445 $Y2=2.09
r89 28 40 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.975 $Y=1.1 $X2=0.975
+ $Y2=1.01
r90 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.975
+ $Y=1.1 $X2=0.975 $Y2=1.1
r91 25 32 0.221902 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=0.365 $Y=1.1
+ $X2=0.24 $Y2=1.1
r92 25 27 21.3027 $w=3.28e-07 $l=6.1e-07 $layer=LI1_cond $X=0.365 $Y=1.1
+ $X2=0.975 $Y2=1.1
r93 21 33 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.28 $Y=2.175
+ $X2=0.28 $Y2=2.09
r94 21 23 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=0.28 $Y=2.175
+ $X2=0.28 $Y2=2.465
r95 20 33 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=0.2 $Y=2.005
+ $X2=0.28 $Y2=2.09
r96 19 32 7.38875 $w=2.1e-07 $l=1.83916e-07 $layer=LI1_cond $X=0.2 $Y=1.265
+ $X2=0.24 $Y2=1.1
r97 19 20 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=0.2 $Y=1.265 $X2=0.2
+ $Y2=2.005
r98 15 32 7.38875 $w=2.1e-07 $l=1.65e-07 $layer=LI1_cond $X=0.24 $Y=0.935
+ $X2=0.24 $Y2=1.1
r99 15 17 16.3647 $w=2.48e-07 $l=3.55e-07 $layer=LI1_cond $X=0.24 $Y=0.935
+ $X2=0.24 $Y2=0.58
r100 12 36 52.2586 $w=2.99e-07 $l=2.57391e-07 $layer=POLY_cond $X=2.485 $Y=2.245
+ $X2=2.5 $Y2=1.995
r101 12 14 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.485 $Y=2.245
+ $X2=2.485 $Y2=2.64
r102 9 11 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.485 $Y=0.935
+ $X2=1.485 $Y2=0.615
r103 8 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.14 $Y=1.01
+ $X2=0.975 $Y2=1.01
r104 7 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.41 $Y=1.01
+ $X2=1.485 $Y2=0.935
r105 7 8 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=1.41 $Y=1.01 $X2=1.14
+ $Y2=1.01
r106 2 23 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.32 $X2=0.28 $Y2=2.465
r107 1 17 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTP_2%SCE 2 5 7 9 11 12 14 19 21 22 23 24 25 28
+ 29 30 31 42
c79 28 0 2.07913e-19 $X=2.51 $Y=1.425
r80 39 40 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.45
+ $Y=1.67 $X2=1.45 $Y2=1.67
r81 36 39 118.906 $w=3.3e-07 $l=6.8e-07 $layer=POLY_cond $X=0.77 $Y=1.67
+ $X2=1.45 $Y2=1.67
r82 31 40 7.68295 $w=3.43e-07 $l=2.3e-07 $layer=LI1_cond $X=1.68 $Y=1.662
+ $X2=1.45 $Y2=1.662
r83 30 40 8.35104 $w=3.43e-07 $l=2.5e-07 $layer=LI1_cond $X=1.2 $Y=1.662
+ $X2=1.45 $Y2=1.662
r84 29 30 16.034 $w=3.43e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.662 $X2=1.2
+ $Y2=1.662
r85 29 36 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.77
+ $Y=1.67 $X2=0.77 $Y2=1.67
r86 28 42 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.51 $Y=1.425
+ $X2=2.51 $Y2=1.26
r87 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.51
+ $Y=1.425 $X2=2.51 $Y2=1.425
r88 25 31 11.7917 $w=3.43e-07 $l=3.53e-07 $layer=LI1_cond $X=2.033 $Y=1.662
+ $X2=1.68 $Y2=1.662
r89 25 27 16.9138 $w=3.45e-07 $l=5.31398e-07 $layer=LI1_cond $X=2.033 $Y=1.662
+ $X2=2.51 $Y2=1.547
r90 24 42 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=2.6 $Y=1.05 $X2=2.6
+ $Y2=1.26
r91 23 24 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=2.625 $Y=0.9 $X2=2.625
+ $Y2=1.05
r92 22 39 14.8632 $w=3.3e-07 $l=8.5e-08 $layer=POLY_cond $X=1.535 $Y=1.67
+ $X2=1.45 $Y2=1.67
r93 20 36 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=0.595 $Y=1.67
+ $X2=0.77 $Y2=1.67
r94 20 21 3.90195 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.595 $Y=1.67
+ $X2=0.505 $Y2=1.67
r95 19 23 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.65 $Y=0.615
+ $X2=2.65 $Y2=0.9
r96 12 14 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.625 $Y=2.245
+ $X2=1.625 $Y2=2.64
r97 11 12 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.625 $Y=2.155
+ $X2=1.625 $Y2=2.245
r98 10 22 30.0773 $w=3.3e-07 $l=2.05122e-07 $layer=POLY_cond $X=1.625 $Y=1.835
+ $X2=1.535 $Y2=1.67
r99 10 11 124.387 $w=1.8e-07 $l=3.2e-07 $layer=POLY_cond $X=1.625 $Y=1.835
+ $X2=1.625 $Y2=2.155
r100 7 9 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.505 $Y=2.245
+ $X2=0.505 $Y2=2.64
r101 3 21 34.7346 $w=1.65e-07 $l=1.69926e-07 $layer=POLY_cond $X=0.495 $Y=1.505
+ $X2=0.505 $Y2=1.67
r102 3 5 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=0.495 $Y=1.505
+ $X2=0.495 $Y2=0.58
r103 2 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.505 $Y=2.155
+ $X2=0.505 $Y2=2.245
r104 1 21 34.7346 $w=1.65e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.835
+ $X2=0.505 $Y2=1.67
r105 1 2 124.387 $w=1.8e-07 $l=3.2e-07 $layer=POLY_cond $X=0.505 $Y=1.835
+ $X2=0.505 $Y2=2.155
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTP_2%D 3 5 8 9 10 13 15
c44 10 0 1.7437e-20 $X=1.68 $Y=0.925
c45 9 0 9.95498e-21 $X=2.04 $Y=2.245
r46 13 16 42.5558 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=1.947 $Y=1.1
+ $X2=1.947 $Y2=1.265
r47 13 15 46.504 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=1.947 $Y=1.1
+ $X2=1.947 $Y2=0.935
r48 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.935
+ $Y=1.1 $X2=1.935 $Y2=1.1
r49 10 14 4.76417 $w=6.53e-07 $l=2.55e-07 $layer=LI1_cond $X=1.68 $Y=0.93
+ $X2=1.935 $Y2=0.93
r50 8 9 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.045 $Y=2.64
+ $X2=2.045 $Y2=2.245
r51 5 9 36.7214 $w=1.7e-07 $l=8.5e-08 $layer=POLY_cond $X=2.04 $Y=2.16 $X2=2.04
+ $Y2=2.245
r52 5 16 378.412 $w=1.7e-07 $l=8.95e-07 $layer=POLY_cond $X=2.04 $Y=2.16
+ $X2=2.04 $Y2=1.265
r53 3 15 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.875 $Y=0.615
+ $X2=1.875 $Y2=0.935
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTP_2%SCD 3 6 10 11 12 13 18 26
c43 12 0 3.4563e-19 $X=3.12 $Y=1.665
c44 6 0 1.49819e-19 $X=3.04 $Y=0.615
r45 26 27 1.39543 $w=3.98e-07 $l=3.5e-08 $layer=LI1_cond $X=3.075 $Y=2.035
+ $X2=3.075 $Y2=2
r46 13 26 0.720277 $w=3.98e-07 $l=2.5e-08 $layer=LI1_cond $X=3.075 $Y=2.06
+ $X2=3.075 $Y2=2.035
r47 13 27 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=3.11 $Y=1.975
+ $X2=3.11 $Y2=2
r48 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.11 $Y=1.605
+ $X2=3.11 $Y2=1.975
r49 12 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.05
+ $Y=1.605 $X2=3.05 $Y2=1.605
r50 10 18 83.0591 $w=3.3e-07 $l=4.75e-07 $layer=POLY_cond $X=3.05 $Y=2.08
+ $X2=3.05 $Y2=1.605
r51 10 11 38.3209 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.05 $Y=2.08
+ $X2=3.05 $Y2=2.245
r52 9 18 38.0424 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.05 $Y=1.44
+ $X2=3.05 $Y2=1.605
r53 6 9 423.032 $w=1.5e-07 $l=8.25e-07 $layer=POLY_cond $X=3.04 $Y=0.615
+ $X2=3.04 $Y2=1.44
r54 3 11 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.035 $Y=2.64
+ $X2=3.035 $Y2=2.245
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTP_2%CLK 1 2 3 5 7 10 12 13 16 19
c54 16 0 1.89542e-19 $X=4.08 $Y=1.295
c55 13 0 1.4151e-19 $X=4.62 $Y=1.885
r56 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.95
+ $Y=1.115 $X2=3.95 $Y2=1.115
r57 16 20 6.1 $w=3.6e-07 $l=1.8e-07 $layer=LI1_cond $X=3.99 $Y=1.295 $X2=3.99
+ $Y2=1.115
r58 11 19 51.5841 $w=3.3e-07 $l=2.95e-07 $layer=POLY_cond $X=3.95 $Y=1.41
+ $X2=3.95 $Y2=1.115
r59 10 13 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=4.645 $Y=2.46
+ $X2=4.645 $Y2=1.885
r60 7 13 37.4512 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=4.62 $Y=1.785 $X2=4.62
+ $Y2=1.885
r61 6 12 23.6879 $w=1.75e-07 $l=1.05e-07 $layer=POLY_cond $X=4.62 $Y=1.62
+ $X2=4.62 $Y2=1.515
r62 6 7 54.7102 $w=2e-07 $l=1.65e-07 $layer=POLY_cond $X=4.62 $Y=1.62 $X2=4.62
+ $Y2=1.785
r63 3 12 23.6879 $w=1.75e-07 $l=1.16833e-07 $layer=POLY_cond $X=4.595 $Y=1.41
+ $X2=4.62 $Y2=1.515
r64 3 5 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=4.595 $Y=1.41
+ $X2=4.595 $Y2=0.965
r65 2 11 28.6974 $w=2.1e-07 $l=2.11069e-07 $layer=POLY_cond $X=4.115 $Y=1.515
+ $X2=3.95 $Y2=1.41
r66 1 12 2.7459 $w=2.1e-07 $l=1e-07 $layer=POLY_cond $X=4.52 $Y=1.515 $X2=4.62
+ $Y2=1.515
r67 1 2 127.894 $w=2.1e-07 $l=4.05e-07 $layer=POLY_cond $X=4.52 $Y=1.515
+ $X2=4.115 $Y2=1.515
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTP_2%A_1034_392# 1 2 8 9 11 12 16 18 20 21 22 23
+ 25 26 33 35 36 37 38 40 44 45 46 48 49 50 52 53 54 57 60 64 68
c207 57 0 8.16714e-20 $X=9.645 $Y=1.17
c208 54 0 9.62383e-20 $X=9.26 $Y=1.17
c209 53 0 1.18082e-19 $X=9.785 $Y=1.17
c210 46 0 1.61901e-19 $X=7.22 $Y=0.665
c211 23 0 4.68929e-20 $X=10.11 $Y=2.465
c212 21 0 2.95884e-20 $X=9.48 $Y=1.26
c213 9 0 1.58245e-19 $X=6.135 $Y=2.21
r214 63 64 9.72653 $w=4.03e-07 $l=2.15e-07 $layer=LI1_cond $X=5.422 $Y=1.07
+ $X2=5.422 $Y2=1.285
r215 60 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.95
+ $Y=2.165 $X2=9.95 $Y2=2.165
r216 58 60 36.0954 $w=2.63e-07 $l=8.3e-07 $layer=LI1_cond $X=9.917 $Y=1.335
+ $X2=9.917 $Y2=2.165
r217 57 74 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=9.645 $Y=1.17
+ $X2=9.645 $Y2=1.26
r218 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.645
+ $Y=1.17 $X2=9.645 $Y2=1.17
r219 54 56 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=9.26 $Y=1.17
+ $X2=9.645 $Y2=1.17
r220 53 58 6.92284 $w=3.3e-07 $l=2.21371e-07 $layer=LI1_cond $X=9.785 $Y=1.17
+ $X2=9.917 $Y2=1.335
r221 53 56 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=9.785 $Y=1.17
+ $X2=9.645 $Y2=1.17
r222 52 54 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.175 $Y=1.005
+ $X2=9.26 $Y2=1.17
r223 51 52 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=9.175 $Y=0.425
+ $X2=9.175 $Y2=1.005
r224 49 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.09 $Y=0.34
+ $X2=9.175 $Y2=0.425
r225 49 50 64.5882 $w=1.68e-07 $l=9.9e-07 $layer=LI1_cond $X=9.09 $Y=0.34
+ $X2=8.1 $Y2=0.34
r226 47 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.015 $Y=0.425
+ $X2=8.1 $Y2=0.34
r227 47 48 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=8.015 $Y=0.425
+ $X2=8.015 $Y2=0.58
r228 45 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.93 $Y=0.665
+ $X2=8.015 $Y2=0.58
r229 45 46 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=7.93 $Y=0.665
+ $X2=7.22 $Y2=0.665
r230 44 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.135 $Y=0.58
+ $X2=7.22 $Y2=0.665
r231 43 44 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=7.135 $Y=0.425
+ $X2=7.135 $Y2=0.58
r232 41 71 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.085 $Y=1.71
+ $X2=6.085 $Y2=1.875
r233 41 68 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=6.085 $Y=1.71
+ $X2=6.085 $Y2=1.635
r234 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.085
+ $Y=1.71 $X2=6.085 $Y2=1.71
r235 38 40 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=5.63 $Y=1.71
+ $X2=6.085 $Y2=1.71
r236 36 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.05 $Y=0.34
+ $X2=7.135 $Y2=0.425
r237 36 37 93.2941 $w=1.68e-07 $l=1.43e-06 $layer=LI1_cond $X=7.05 $Y=0.34
+ $X2=5.62 $Y2=0.34
r238 35 38 10.1667 $w=1.78e-07 $l=1.65e-07 $layer=LI1_cond $X=5.54 $Y=1.545
+ $X2=5.54 $Y2=1.71
r239 35 64 16.0202 $w=1.78e-07 $l=2.6e-07 $layer=LI1_cond $X=5.54 $Y=1.545
+ $X2=5.54 $Y2=1.285
r240 33 63 8.25206 $w=4.03e-07 $l=2.9e-07 $layer=LI1_cond $X=5.417 $Y=0.78
+ $X2=5.417 $Y2=1.07
r241 30 37 8.41448 $w=1.7e-07 $l=2.41793e-07 $layer=LI1_cond $X=5.417 $Y=0.425
+ $X2=5.62 $Y2=0.34
r242 30 33 10.1017 $w=4.03e-07 $l=3.55e-07 $layer=LI1_cond $X=5.417 $Y=0.425
+ $X2=5.417 $Y2=0.78
r243 26 38 23.1061 $w=1.78e-07 $l=3.75e-07 $layer=LI1_cond $X=5.54 $Y=2.085
+ $X2=5.54 $Y2=1.71
r244 26 28 5.76222 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=5.45 $Y=2.085
+ $X2=5.32 $Y2=2.085
r245 23 61 57.5457 $w=3.46e-07 $l=3.54119e-07 $layer=POLY_cond $X=10.11 $Y=2.465
+ $X2=9.992 $Y2=2.165
r246 23 25 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=10.11 $Y=2.465
+ $X2=10.11 $Y2=2.75
r247 21 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.48 $Y=1.26
+ $X2=9.645 $Y2=1.26
r248 21 22 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=9.48 $Y=1.26
+ $X2=9.12 $Y2=1.26
r249 18 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.045 $Y=1.185
+ $X2=9.12 $Y2=1.26
r250 18 20 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=9.045 $Y=1.185
+ $X2=9.045 $Y2=0.74
r251 14 16 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=6.525 $Y=1.545
+ $X2=6.525 $Y2=0.805
r252 13 68 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.25 $Y=1.635
+ $X2=6.085 $Y2=1.635
r253 12 14 27.2212 $w=1.8e-07 $l=1.21861e-07 $layer=POLY_cond $X=6.45 $Y=1.635
+ $X2=6.525 $Y2=1.545
r254 12 13 77.7419 $w=1.8e-07 $l=2e-07 $layer=POLY_cond $X=6.45 $Y=1.635
+ $X2=6.25 $Y2=1.635
r255 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.135 $Y=2.21
+ $X2=6.135 $Y2=2.495
r256 8 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.135 $Y=2.12 $X2=6.135
+ $Y2=2.21
r257 8 71 95.2339 $w=1.8e-07 $l=2.45e-07 $layer=POLY_cond $X=6.135 $Y=2.12
+ $X2=6.135 $Y2=1.875
r258 2 28 600 $w=1.7e-07 $l=2.33238e-07 $layer=licon1_PDIFF $count=1 $X=5.17
+ $Y=1.96 $X2=5.32 $Y2=2.13
r259 1 33 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=5.22
+ $Y=0.595 $X2=5.36 $Y2=0.78
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTP_2%A_1367_93# 1 2 9 13 17 18 21 26 30 31 34 35
c100 9 0 1.43931e-19 $X=6.91 $Y=0.805
r101 36 38 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=6.91 $Y=1.64
+ $X2=6.945 $Y2=1.64
r102 34 35 8.52431 $w=3.63e-07 $l=1.65e-07 $layer=LI1_cond $X=8.932 $Y=1.88
+ $X2=8.932 $Y2=1.715
r103 29 31 1.93306 $w=4.93e-07 $l=8e-08 $layer=LI1_cond $X=8.755 $Y=0.842
+ $X2=8.835 $Y2=0.842
r104 29 30 17.2188 $w=4.93e-07 $l=4.85e-07 $layer=LI1_cond $X=8.755 $Y=0.842
+ $X2=8.27 $Y2=0.842
r105 24 34 0.536754 $w=3.63e-07 $l=1.7e-08 $layer=LI1_cond $X=8.932 $Y=1.897
+ $X2=8.932 $Y2=1.88
r106 24 26 10.6719 $w=3.63e-07 $l=3.38e-07 $layer=LI1_cond $X=8.932 $Y=1.897
+ $X2=8.932 $Y2=2.235
r107 22 31 7.09362 $w=1.7e-07 $l=2.48e-07 $layer=LI1_cond $X=8.835 $Y=1.09
+ $X2=8.835 $Y2=0.842
r108 22 35 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=8.835 $Y=1.09
+ $X2=8.835 $Y2=1.715
r109 21 30 65.5668 $w=1.68e-07 $l=1.005e-06 $layer=LI1_cond $X=7.265 $Y=1.005
+ $X2=8.27 $Y2=1.005
r110 18 38 34.9723 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=7.145 $Y=1.64
+ $X2=6.945 $Y2=1.64
r111 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.145
+ $Y=1.64 $X2=7.145 $Y2=1.64
r112 15 21 7.07814 $w=1.7e-07 $l=1.56844e-07 $layer=LI1_cond $X=7.145 $Y=1.09
+ $X2=7.265 $Y2=1.005
r113 15 17 26.4102 $w=2.38e-07 $l=5.5e-07 $layer=LI1_cond $X=7.145 $Y=1.09
+ $X2=7.145 $Y2=1.64
r114 11 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.945 $Y=1.805
+ $X2=6.945 $Y2=1.64
r115 11 13 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.945 $Y=1.805
+ $X2=6.945 $Y2=2.495
r116 7 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.91 $Y=1.475
+ $X2=6.91 $Y2=1.64
r117 7 9 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=6.91 $Y=1.475
+ $X2=6.91 $Y2=0.805
r118 2 34 600 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=1 $X=8.715
+ $Y=1.735 $X2=8.95 $Y2=1.88
r119 2 26 300 $w=1.7e-07 $l=6.06218e-07 $layer=licon1_PDIFF $count=2 $X=8.715
+ $Y=1.735 $X2=8.95 $Y2=2.235
r120 1 29 182 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_NDIFF $count=1 $X=8.615
+ $Y=0.37 $X2=8.755 $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTP_2%RESET_B 4 7 8 9 10 11 15 16 18 20 23 26 27
+ 29 32 35 37 38 39 40 47 48 52 54 60 68
c220 52 0 1.4151e-19 $X=3.95 $Y=1.995
c221 40 0 1.09002e-19 $X=8.545 $Y=2.035
c222 37 0 6.54652e-20 $X=8.255 $Y=2.035
c223 32 0 9.37604e-20 $X=3.56 $Y=2.245
c224 27 0 1.84389e-19 $X=11.35 $Y=2.465
c225 15 0 1.75393e-19 $X=7.3 $Y=0.805
r226 60 62 11.8137 $w=3.06e-07 $l=7.5e-08 $layer=POLY_cond $X=11.275 $Y=2.07
+ $X2=11.35 $Y2=2.07
r227 60 68 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.275
+ $Y=2.07 $X2=11.275 $Y2=2.07
r228 58 60 22.0523 $w=3.06e-07 $l=1.4e-07 $layer=POLY_cond $X=11.135 $Y=2.07
+ $X2=11.275 $Y2=2.07
r229 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.86
+ $Y=1.96 $X2=7.86 $Y2=1.96
r230 54 56 39.5449 $w=3.23e-07 $l=2.65e-07 $layer=POLY_cond $X=7.595 $Y=2.002
+ $X2=7.86 $Y2=2.002
r231 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.95
+ $Y=1.995 $X2=3.95 $Y2=1.995
r232 48 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=2.035
+ $X2=11.28 $Y2=2.035
r233 47 57 17.5301 $w=3.53e-07 $l=5.4e-07 $layer=LI1_cond $X=8.4 $Y=1.972
+ $X2=7.86 $Y2=1.972
r234 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=2.035
+ $X2=8.4 $Y2=2.035
r235 42 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=2.035
+ $X2=4.08 $Y2=2.035
r236 40 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.545 $Y=2.035
+ $X2=8.4 $Y2=2.035
r237 39 48 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=11.135 $Y=2.035
+ $X2=11.28 $Y2=2.035
r238 39 40 3.20544 $w=1.4e-07 $l=2.59e-06 $layer=MET1_cond $X=11.135 $Y=2.035
+ $X2=8.545 $Y2=2.035
r239 38 42 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.225 $Y=2.035
+ $X2=4.08 $Y2=2.035
r240 37 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.255 $Y=2.035
+ $X2=8.4 $Y2=2.035
r241 37 38 4.98761 $w=1.4e-07 $l=4.03e-06 $layer=MET1_cond $X=8.255 $Y=2.035
+ $X2=4.225 $Y2=2.035
r242 33 35 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=7.3 $Y=1.19
+ $X2=7.595 $Y2=1.19
r243 27 29 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=11.35 $Y=2.465
+ $X2=11.35 $Y2=2.75
r244 26 27 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=11.35 $Y=2.375
+ $X2=11.35 $Y2=2.465
r245 25 62 15.178 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=11.35 $Y=2.235
+ $X2=11.35 $Y2=2.07
r246 25 26 54.4194 $w=1.8e-07 $l=1.4e-07 $layer=POLY_cond $X=11.35 $Y=2.235
+ $X2=11.35 $Y2=2.375
r247 21 58 19.4347 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.135 $Y=1.905
+ $X2=11.135 $Y2=2.07
r248 21 23 679.415 $w=1.5e-07 $l=1.325e-06 $layer=POLY_cond $X=11.135 $Y=1.905
+ $X2=11.135 $Y2=0.58
r249 20 54 20.7134 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.595 $Y=1.795
+ $X2=7.595 $Y2=2.002
r250 19 35 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.595 $Y=1.265
+ $X2=7.595 $Y2=1.19
r251 19 20 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=7.595 $Y=1.265
+ $X2=7.595 $Y2=1.795
r252 16 54 29.8452 $w=3.23e-07 $l=2.91314e-07 $layer=POLY_cond $X=7.395 $Y=2.21
+ $X2=7.595 $Y2=2.002
r253 16 18 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.395 $Y=2.21
+ $X2=7.395 $Y2=2.495
r254 13 33 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.3 $Y=1.115
+ $X2=7.3 $Y2=1.19
r255 13 15 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=7.3 $Y=1.115
+ $X2=7.3 $Y2=0.805
r256 12 15 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=7.3 $Y=0.255
+ $X2=7.3 $Y2=0.805
r257 11 32 67.3007 $w=2.7e-07 $l=2.5e-07 $layer=POLY_cond $X=3.56 $Y=1.995
+ $X2=3.56 $Y2=2.245
r258 11 31 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.56 $Y=1.995
+ $X2=3.56 $Y2=1.83
r259 10 51 2.92121 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=3.93 $Y=1.995
+ $X2=3.95 $Y2=1.995
r260 10 11 41.0924 $w=3.3e-07 $l=2.35e-07 $layer=POLY_cond $X=3.93 $Y=1.995
+ $X2=3.695 $Y2=1.995
r261 8 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.225 $Y=0.18
+ $X2=7.3 $Y2=0.255
r262 8 9 1871.6 $w=1.5e-07 $l=3.65e-06 $layer=POLY_cond $X=7.225 $Y=0.18
+ $X2=3.575 $Y2=0.18
r263 7 32 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.605 $Y=2.64
+ $X2=3.605 $Y2=2.245
r264 4 31 623.011 $w=1.5e-07 $l=1.215e-06 $layer=POLY_cond $X=3.5 $Y=0.615
+ $X2=3.5 $Y2=1.83
r265 1 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.5 $Y=0.255
+ $X2=3.575 $Y2=0.18
r266 1 4 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=3.5 $Y=0.255 $X2=3.5
+ $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTP_2%A_1234_119# 1 2 3 12 14 16 18 19 23 26 28
+ 29 32 35 37 41 45 46 48 49
c126 45 0 7.56682e-20 $X=6.77 $Y=2.075
c127 26 0 1.75393e-19 $X=6.77 $Y=1.985
c128 23 0 1.51844e-20 $X=6.685 $Y=0.945
c129 19 0 1.58245e-19 $X=6.685 $Y=2.555
c130 12 0 9.62383e-20 $X=8.54 $Y=0.74
r131 48 49 10.0337 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=7.6 $Y=2.53 $X2=7.6
+ $Y2=2.32
r132 41 43 4.78707 $w=3.23e-07 $l=1.35e-07 $layer=LI1_cond $X=6.307 $Y=0.81
+ $X2=6.307 $Y2=0.945
r133 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.255
+ $Y=1.41 $X2=8.255 $Y2=1.41
r134 35 37 26.2838 $w=2.83e-07 $l=6.5e-07 $layer=LI1_cond $X=7.605 $Y=1.402
+ $X2=8.255 $Y2=1.402
r135 33 46 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=7.52 $Y=2.165 $X2=7.52
+ $Y2=2.075
r136 33 49 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=7.52 $Y=2.165
+ $X2=7.52 $Y2=2.32
r137 32 46 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=7.52 $Y=1.985 $X2=7.52
+ $Y2=2.075
r138 31 35 7.39867 $w=2.85e-07 $l=1.80566e-07 $layer=LI1_cond $X=7.52 $Y=1.545
+ $X2=7.605 $Y2=1.402
r139 31 32 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=7.52 $Y=1.545
+ $X2=7.52 $Y2=1.985
r140 30 45 1.13756 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=6.855 $Y=2.075
+ $X2=6.77 $Y2=2.075
r141 29 46 1.13756 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=7.435 $Y=2.075
+ $X2=7.52 $Y2=2.075
r142 29 30 35.7374 $w=1.78e-07 $l=5.8e-07 $layer=LI1_cond $X=7.435 $Y=2.075
+ $X2=6.855 $Y2=2.075
r143 27 45 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=6.77 $Y=2.165 $X2=6.77
+ $Y2=2.075
r144 27 28 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=6.77 $Y=2.165
+ $X2=6.77 $Y2=2.385
r145 26 45 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=6.77 $Y=1.985 $X2=6.77
+ $Y2=2.075
r146 25 26 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=6.77 $Y=1.03
+ $X2=6.77 $Y2=1.985
r147 24 43 4.53325 $w=1.7e-07 $l=1.63e-07 $layer=LI1_cond $X=6.47 $Y=0.945
+ $X2=6.307 $Y2=0.945
r148 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.685 $Y=0.945
+ $X2=6.77 $Y2=1.03
r149 23 24 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=6.685 $Y=0.945
+ $X2=6.47 $Y2=0.945
r150 19 28 7.85115 $w=3.4e-07 $l=2.08207e-07 $layer=LI1_cond $X=6.685 $Y=2.555
+ $X2=6.77 $Y2=2.385
r151 19 21 11.016 $w=3.38e-07 $l=3.25e-07 $layer=LI1_cond $X=6.685 $Y=2.555
+ $X2=6.36 $Y2=2.555
r152 18 38 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=8.465 $Y=1.41
+ $X2=8.255 $Y2=1.41
r153 14 18 64.0286 $w=1.97e-07 $l=2.70647e-07 $layer=POLY_cond $X=8.64 $Y=1.66
+ $X2=8.597 $Y2=1.41
r154 14 16 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=8.64 $Y=1.66
+ $X2=8.64 $Y2=2.235
r155 10 18 43.2316 $w=1.97e-07 $l=1.9139e-07 $layer=POLY_cond $X=8.54 $Y=1.245
+ $X2=8.597 $Y2=1.41
r156 10 12 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=8.54 $Y=1.245
+ $X2=8.54 $Y2=0.74
r157 3 48 600 $w=1.7e-07 $l=3.11087e-07 $layer=licon1_PDIFF $count=1 $X=7.47
+ $Y=2.285 $X2=7.62 $Y2=2.53
r158 2 21 600 $w=1.7e-07 $l=3.36749e-07 $layer=licon1_PDIFF $count=1 $X=6.21
+ $Y=2.285 $X2=6.36 $Y2=2.555
r159 1 41 182 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=1 $X=6.17
+ $Y=0.595 $X2=6.31 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTP_2%A_835_98# 1 2 7 9 10 12 14 15 16 17 19 21
+ 24 26 31 32 33 35 38 40 41 45 48 50 54 57
c180 57 0 1.89542e-19 $X=5.115 $Y=1.635
c181 54 0 9.37604e-20 $X=4.93 $Y=1.852
c182 24 0 7.56682e-20 $X=6.585 $Y=2.495
c183 19 0 1.51844e-20 $X=6.095 $Y=1.115
c184 7 0 1.94423e-19 $X=5.095 $Y=1.875
r185 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.115
+ $Y=1.635 $X2=5.115 $Y2=1.635
r186 54 56 5.21247 $w=4.33e-07 $l=2.95354e-07 $layer=LI1_cond $X=4.93 $Y=1.852
+ $X2=5.115 $Y2=1.635
r187 53 54 14.3695 $w=4.33e-07 $l=5.1e-07 $layer=LI1_cond $X=4.42 $Y=1.852
+ $X2=4.93 $Y2=1.852
r188 48 54 4.44229 $w=2.3e-07 $l=3.97e-07 $layer=LI1_cond $X=4.93 $Y=1.455
+ $X2=4.93 $Y2=1.852
r189 47 50 24.8067 $w=3e-07 $l=7.35989e-07 $layer=LI1_cond $X=4.93 $Y=1.08
+ $X2=4.32 $Y2=0.802
r190 47 48 18.7898 $w=2.28e-07 $l=3.75e-07 $layer=LI1_cond $X=4.93 $Y=1.08
+ $X2=4.93 $Y2=1.455
r191 43 45 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=10.125 $Y=1.055
+ $X2=10.315 $Y2=1.055
r192 36 45 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.315 $Y=0.98
+ $X2=10.315 $Y2=1.055
r193 36 38 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=10.315 $Y=0.98
+ $X2=10.315 $Y2=0.58
r194 34 43 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.125 $Y=1.13
+ $X2=10.125 $Y2=1.055
r195 34 35 228.181 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=10.125 $Y=1.13
+ $X2=10.125 $Y2=1.575
r196 32 35 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.05 $Y=1.65
+ $X2=10.125 $Y2=1.575
r197 32 33 358.936 $w=1.5e-07 $l=7e-07 $layer=POLY_cond $X=10.05 $Y=1.65
+ $X2=9.35 $Y2=1.65
r198 29 41 97.3837 $w=1.8e-07 $l=2.45e-07 $layer=POLY_cond $X=9.26 $Y=2.905
+ $X2=9.26 $Y2=3.15
r199 29 31 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=9.26 $Y=2.905
+ $X2=9.26 $Y2=2.33
r200 28 33 26.9307 $w=1.5e-07 $l=1.43091e-07 $layer=POLY_cond $X=9.26 $Y=1.755
+ $X2=9.35 $Y2=1.65
r201 28 31 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=9.26 $Y=1.755
+ $X2=9.26 $Y2=2.33
r202 27 40 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.66 $Y=3.15
+ $X2=6.585 $Y2=3.15
r203 26 41 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=9.17 $Y=3.15 $X2=9.26
+ $Y2=3.15
r204 26 27 1287.04 $w=1.5e-07 $l=2.51e-06 $layer=POLY_cond $X=9.17 $Y=3.15
+ $X2=6.66 $Y2=3.15
r205 22 40 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.585 $Y=3.075
+ $X2=6.585 $Y2=3.15
r206 22 24 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.585 $Y=3.075
+ $X2=6.585 $Y2=2.495
r207 19 21 99.6133 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=6.095 $Y=1.115
+ $X2=6.095 $Y2=0.805
r208 18 57 37.7859 $w=5.23e-07 $l=5.69122e-07 $layer=POLY_cond $X=5.71 $Y=1.225
+ $X2=5.33 $Y2=1.635
r209 17 19 28.2037 $w=2.2e-07 $l=1.42653e-07 $layer=POLY_cond $X=6.02 $Y=1.225
+ $X2=6.095 $Y2=1.115
r210 17 18 90.4236 $w=2.2e-07 $l=3.1e-07 $layer=POLY_cond $X=6.02 $Y=1.225
+ $X2=5.71 $Y2=1.225
r211 15 40 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.51 $Y=3.15
+ $X2=6.585 $Y2=3.15
r212 15 16 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=6.51 $Y=3.15
+ $X2=5.69 $Y2=3.15
r213 14 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.615 $Y=3.075
+ $X2=5.69 $Y2=3.15
r214 13 57 46.2206 $w=2.61e-07 $l=3.86814e-07 $layer=POLY_cond $X=5.615 $Y=1.875
+ $X2=5.33 $Y2=1.635
r215 13 14 615.319 $w=1.5e-07 $l=1.2e-06 $layer=POLY_cond $X=5.615 $Y=1.875
+ $X2=5.615 $Y2=3.075
r216 10 18 44.3687 $w=5.23e-07 $l=6.50961e-07 $layer=POLY_cond $X=5.145 $Y=1.41
+ $X2=5.71 $Y2=1.225
r217 10 12 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=5.145 $Y=1.41
+ $X2=5.145 $Y2=0.965
r218 7 57 46.2206 $w=2.61e-07 $l=3.37639e-07 $layer=POLY_cond $X=5.095 $Y=1.875
+ $X2=5.33 $Y2=1.635
r219 7 9 187.98 $w=1.5e-07 $l=5.85e-07 $layer=POLY_cond $X=5.095 $Y=1.875
+ $X2=5.095 $Y2=2.46
r220 2 53 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=4.275
+ $Y=1.96 $X2=4.42 $Y2=2.085
r221 1 50 182 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_NDIFF $count=1 $X=4.175
+ $Y=0.49 $X2=4.32 $Y2=0.665
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTP_2%A_2082_446# 1 2 7 9 12 14 18 19 20 22 23 26
+ 30 32 33 35 37 38
c122 23 0 4.68929e-20 $X=10.85 $Y=2.475
c123 18 0 2.97873e-19 $X=10.685 $Y=2.215
c124 12 0 1.18082e-19 $X=10.705 $Y=0.58
r125 38 41 5.42589 $w=4.1e-07 $l=4e-08 $layer=POLY_cond $X=10.645 $Y=1.535
+ $X2=10.645 $Y2=1.575
r126 38 44 45.9078 $w=4.1e-07 $l=1.65e-07 $layer=POLY_cond $X=10.645 $Y=1.535
+ $X2=10.645 $Y2=1.37
r127 37 40 5.16612 $w=2.88e-07 $l=1.3e-07 $layer=LI1_cond $X=10.705 $Y=1.535
+ $X2=10.705 $Y2=1.665
r128 37 38 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=10.685
+ $Y=1.535 $X2=10.685 $Y2=1.535
r129 34 35 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=12.145 $Y=0.94
+ $X2=12.145 $Y2=1.58
r130 32 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=12.06 $Y=0.855
+ $X2=12.145 $Y2=0.94
r131 32 33 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=12.06 $Y=0.855
+ $X2=11.875 $Y2=0.855
r132 28 33 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=11.71 $Y=0.77
+ $X2=11.875 $Y2=0.855
r133 28 30 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=11.71 $Y=0.77
+ $X2=11.71 $Y2=0.58
r134 24 26 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=11.575 $Y=2.56
+ $X2=11.575 $Y2=2.75
r135 22 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=11.41 $Y=2.475
+ $X2=11.575 $Y2=2.56
r136 22 23 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=11.41 $Y=2.475
+ $X2=10.85 $Y2=2.475
r137 21 40 3.86198 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=10.85 $Y=1.665
+ $X2=10.705 $Y2=1.665
r138 20 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=12.06 $Y=1.665
+ $X2=12.145 $Y2=1.58
r139 20 21 78.9412 $w=1.68e-07 $l=1.21e-06 $layer=LI1_cond $X=12.06 $Y=1.665
+ $X2=10.85 $Y2=1.665
r140 19 41 86.8143 $w=4.1e-07 $l=6.4e-07 $layer=POLY_cond $X=10.645 $Y=2.215
+ $X2=10.645 $Y2=1.575
r141 18 19 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=10.685
+ $Y=2.215 $X2=10.685 $Y2=2.215
r142 16 23 7.43784 $w=1.7e-07 $l=1.8262e-07 $layer=LI1_cond $X=10.705 $Y=2.39
+ $X2=10.85 $Y2=2.475
r143 16 18 6.9544 $w=2.88e-07 $l=1.75e-07 $layer=LI1_cond $X=10.705 $Y=2.39
+ $X2=10.705 $Y2=2.215
r144 15 40 3.37785 $w=2.88e-07 $l=8.5e-08 $layer=LI1_cond $X=10.705 $Y=1.75
+ $X2=10.705 $Y2=1.665
r145 15 18 18.4788 $w=2.88e-07 $l=4.65e-07 $layer=LI1_cond $X=10.705 $Y=1.75
+ $X2=10.705 $Y2=2.215
r146 14 19 2.03471 $w=4.1e-07 $l=1.5e-08 $layer=POLY_cond $X=10.645 $Y=2.23
+ $X2=10.645 $Y2=2.215
r147 12 44 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=10.705 $Y=0.58
+ $X2=10.705 $Y2=1.37
r148 7 14 32.8319 $w=3.45e-07 $l=2.98831e-07 $layer=POLY_cond $X=10.5 $Y=2.465
+ $X2=10.645 $Y2=2.23
r149 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=10.5 $Y=2.465 $X2=10.5
+ $Y2=2.75
r150 2 26 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=11.425
+ $Y=2.54 $X2=11.575 $Y2=2.75
r151 1 30 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=11.57
+ $Y=0.37 $X2=11.71 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTP_2%A_1824_74# 1 2 9 11 12 13 15 18 19 21 22 24
+ 25 27 28 29 32 34 38 39 43 45 50 53 54 55
c144 53 0 6.53658e-20 $X=10.305 $Y=1.115
c145 43 0 1.63056e-20 $X=10.305 $Y=1.03
c146 32 0 2.95884e-20 $X=9.485 $Y=2.005
c147 28 0 6.36774e-20 $X=11.8 $Y=1.665
r148 54 55 8.67671 $w=2.98e-07 $l=1.7e-07 $layer=LI1_cond $X=11.02 $Y=1.22
+ $X2=11.19 $Y2=1.22
r149 51 58 15.7174 $w=2.76e-07 $l=9e-08 $layer=POLY_cond $X=11.725 $Y=1.26
+ $X2=11.815 $Y2=1.26
r150 50 55 20.5519 $w=2.98e-07 $l=5.35e-07 $layer=LI1_cond $X=11.725 $Y=1.26
+ $X2=11.19 $Y2=1.26
r151 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.725
+ $Y=1.26 $X2=11.725 $Y2=1.26
r152 47 53 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.39 $Y=1.115
+ $X2=10.305 $Y2=1.115
r153 47 54 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=10.39 $Y=1.115
+ $X2=11.02 $Y2=1.115
r154 44 53 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.305 $Y=1.2
+ $X2=10.305 $Y2=1.115
r155 44 45 86.1176 $w=1.68e-07 $l=1.32e-06 $layer=LI1_cond $X=10.305 $Y=1.2
+ $X2=10.305 $Y2=2.52
r156 43 53 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.305 $Y=1.03
+ $X2=10.305 $Y2=1.115
r157 42 43 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=10.305 $Y=0.81
+ $X2=10.305 $Y2=1.03
r158 39 41 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=9.6 $Y=2.685
+ $X2=9.885 $Y2=2.685
r159 38 45 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=10.22 $Y=2.685
+ $X2=10.305 $Y2=2.52
r160 38 41 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=10.22 $Y=2.685
+ $X2=9.885 $Y2=2.685
r161 34 42 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=10.22 $Y=0.645
+ $X2=10.305 $Y2=0.81
r162 34 36 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=10.22 $Y=0.645
+ $X2=10.1 $Y2=0.645
r163 30 39 6.87623 $w=3.3e-07 $l=2.24332e-07 $layer=LI1_cond $X=9.46 $Y=2.52
+ $X2=9.6 $Y2=2.685
r164 30 32 21.1967 $w=2.78e-07 $l=5.15e-07 $layer=LI1_cond $X=9.46 $Y=2.52
+ $X2=9.46 $Y2=2.005
r165 25 29 34.7346 $w=1.65e-07 $l=1.9e-07 $layer=POLY_cond $X=12.485 $Y=1.095
+ $X2=12.295 $Y2=1.095
r166 25 27 130.14 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=12.485 $Y=1.095
+ $X2=12.485 $Y2=0.69
r167 22 24 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=12.385 $Y=1.885
+ $X2=12.385 $Y2=2.46
r168 21 22 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=12.385 $Y=1.795
+ $X2=12.385 $Y2=1.885
r169 20 29 34.7346 $w=1.65e-07 $l=3.7229e-07 $layer=POLY_cond $X=12.385 $Y=1.425
+ $X2=12.295 $Y2=1.095
r170 20 21 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=12.385 $Y=1.425
+ $X2=12.385 $Y2=1.795
r171 19 58 12.3868 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=11.89 $Y=1.26
+ $X2=11.815 $Y2=1.26
r172 18 29 3.90195 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=12.295 $Y=1.26
+ $X2=12.295 $Y2=1.095
r173 18 19 70.8188 $w=3.3e-07 $l=4.05e-07 $layer=POLY_cond $X=12.295 $Y=1.26
+ $X2=11.89 $Y2=1.26
r174 16 58 17.0164 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.815 $Y=1.425
+ $X2=11.815 $Y2=1.26
r175 16 28 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=11.815 $Y=1.425
+ $X2=11.815 $Y2=1.665
r176 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=11.8 $Y=2.465
+ $X2=11.8 $Y2=2.75
r177 12 13 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=11.8 $Y=2.375
+ $X2=11.8 $Y2=2.465
r178 11 28 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=11.8 $Y=1.755
+ $X2=11.8 $Y2=1.665
r179 11 12 241 $w=1.8e-07 $l=6.2e-07 $layer=POLY_cond $X=11.8 $Y=1.755 $X2=11.8
+ $Y2=2.375
r180 7 51 40.1667 $w=2.76e-07 $l=3.01413e-07 $layer=POLY_cond $X=11.495 $Y=1.095
+ $X2=11.725 $Y2=1.26
r181 7 9 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=11.495 $Y=1.095
+ $X2=11.495 $Y2=0.58
r182 2 41 300 $w=1.7e-07 $l=1.09603e-06 $layer=licon1_PDIFF $count=2 $X=9.335
+ $Y=1.83 $X2=9.885 $Y2=2.685
r183 2 32 300 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=2 $X=9.335
+ $Y=1.83 $X2=9.485 $Y2=2.005
r184 1 36 91 $w=1.7e-07 $l=1.10901e-06 $layer=licon1_NDIFF $count=2 $X=9.12
+ $Y=0.37 $X2=10.1 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTP_2%A_2492_392# 1 2 7 9 12 14 16 19 23 25 29 35
+ 38 39 43
r62 43 44 7.77419 $w=3.72e-07 $l=6e-08 $layer=POLY_cond $X=13.845 $Y=1.532
+ $X2=13.905 $Y2=1.532
r63 42 43 47.9409 $w=3.72e-07 $l=3.7e-07 $layer=POLY_cond $X=13.475 $Y=1.532
+ $X2=13.845 $Y2=1.532
r64 41 42 10.3656 $w=3.72e-07 $l=8e-08 $layer=POLY_cond $X=13.395 $Y=1.532
+ $X2=13.475 $Y2=1.532
r65 36 41 26.5618 $w=3.72e-07 $l=2.05e-07 $layer=POLY_cond $X=13.19 $Y=1.532
+ $X2=13.395 $Y2=1.532
r66 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.19
+ $Y=1.465 $X2=13.19 $Y2=1.465
r67 33 39 0.144206 $w=3.3e-07 $l=1.3e-07 $layer=LI1_cond $X=12.865 $Y=1.465
+ $X2=12.735 $Y2=1.465
r68 33 35 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=12.865 $Y=1.465
+ $X2=13.19 $Y2=1.465
r69 31 39 7.25953 $w=2.15e-07 $l=1.86145e-07 $layer=LI1_cond $X=12.69 $Y=1.63
+ $X2=12.735 $Y2=1.465
r70 31 38 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=12.69 $Y=1.63
+ $X2=12.69 $Y2=1.94
r71 27 39 7.25953 $w=2.15e-07 $l=1.65e-07 $layer=LI1_cond $X=12.735 $Y=1.3
+ $X2=12.735 $Y2=1.465
r72 27 29 34.7949 $w=2.58e-07 $l=7.85e-07 $layer=LI1_cond $X=12.735 $Y=1.3
+ $X2=12.735 $Y2=0.515
r73 23 38 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=12.61 $Y=2.105
+ $X2=12.61 $Y2=1.94
r74 23 25 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=12.61 $Y=2.105
+ $X2=12.61 $Y2=2.815
r75 17 44 24.0971 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=13.905 $Y=1.3
+ $X2=13.905 $Y2=1.532
r76 17 19 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=13.905 $Y=1.3
+ $X2=13.905 $Y2=0.74
r77 14 43 24.0971 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=13.845 $Y=1.765
+ $X2=13.845 $Y2=1.532
r78 14 16 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=13.845 $Y=1.765
+ $X2=13.845 $Y2=2.4
r79 10 42 24.0971 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=13.475 $Y=1.3
+ $X2=13.475 $Y2=1.532
r80 10 12 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=13.475 $Y=1.3
+ $X2=13.475 $Y2=0.74
r81 7 41 24.0971 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=13.395 $Y=1.765
+ $X2=13.395 $Y2=1.532
r82 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=13.395 $Y=1.765
+ $X2=13.395 $Y2=2.4
r83 2 25 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=12.46
+ $Y=1.96 $X2=12.61 $Y2=2.815
r84 2 23 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=12.46
+ $Y=1.96 $X2=12.61 $Y2=2.105
r85 1 29 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=12.56
+ $Y=0.37 $X2=12.7 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTP_2%VPWR 1 2 3 4 5 6 7 8 9 30 34 38 42 46 52 56
+ 58 63 64 66 67 69 70 71 73 78 96 100 112 116 122 129 132 135 142 146
c172 42 0 6.54652e-20 $X=8.415 $Y=2.425
c173 2 0 1.19423e-19 $X=3.11 $Y=2.32
r174 145 146 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.16 $Y=3.33
+ $X2=14.16 $Y2=3.33
r175 142 143 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=3.33
+ $X2=13.2 $Y2=3.33
r176 138 139 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r177 135 138 9.05853 $w=6.78e-07 $l=5.15e-07 $layer=LI1_cond $X=10.9 $Y=2.815
+ $X2=10.9 $Y2=3.33
r178 132 133 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r179 129 130 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r180 125 126 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r181 122 125 11.1084 $w=9.48e-07 $l=8.65e-07 $layer=LI1_cond $X=1.09 $Y=2.465
+ $X2=1.09 $Y2=3.33
r182 120 146 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=3.33
+ $X2=14.16 $Y2=3.33
r183 120 143 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=3.33
+ $X2=13.2 $Y2=3.33
r184 119 120 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=3.33
+ $X2=13.68 $Y2=3.33
r185 117 142 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.335 $Y=3.33
+ $X2=13.17 $Y2=3.33
r186 117 119 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=13.335 $Y=3.33
+ $X2=13.68 $Y2=3.33
r187 116 145 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=13.955 $Y=3.33
+ $X2=14.177 $Y2=3.33
r188 116 119 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=13.955 $Y=3.33
+ $X2=13.68 $Y2=3.33
r189 115 143 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=13.2 $Y2=3.33
r190 114 115 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r191 112 142 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.005 $Y=3.33
+ $X2=13.17 $Y2=3.33
r192 112 114 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=13.005 $Y=3.33
+ $X2=12.72 $Y2=3.33
r193 111 115 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=12.72 $Y2=3.33
r194 111 139 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=10.8 $Y2=3.33
r195 110 111 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r196 108 138 9.13095 $w=1.7e-07 $l=3.4e-07 $layer=LI1_cond $X=11.24 $Y=3.33
+ $X2=10.9 $Y2=3.33
r197 108 110 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=11.24 $Y=3.33
+ $X2=11.76 $Y2=3.33
r198 107 139 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=10.8 $Y2=3.33
r199 106 107 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r200 104 107 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=10.32 $Y2=3.33
r201 104 133 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=8.4 $Y2=3.33
r202 103 106 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=8.88 $Y=3.33
+ $X2=10.32 $Y2=3.33
r203 103 104 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r204 101 132 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=8.58 $Y=3.33
+ $X2=8.412 $Y2=3.33
r205 101 103 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=8.58 $Y=3.33
+ $X2=8.88 $Y2=3.33
r206 100 138 9.13095 $w=1.7e-07 $l=3.4e-07 $layer=LI1_cond $X=10.56 $Y=3.33
+ $X2=10.9 $Y2=3.33
r207 100 106 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=10.56 $Y=3.33
+ $X2=10.32 $Y2=3.33
r208 99 133 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r209 98 99 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r210 96 132 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=8.245 $Y=3.33
+ $X2=8.412 $Y2=3.33
r211 96 98 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=8.245 $Y=3.33
+ $X2=7.92 $Y2=3.33
r212 94 95 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r213 92 95 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=6.96 $Y2=3.33
r214 91 94 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=5.04 $Y=3.33
+ $X2=6.96 $Y2=3.33
r215 91 92 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r216 89 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r217 88 89 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r218 86 89 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r219 86 130 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r220 85 88 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.6 $Y=3.33 $X2=4.56
+ $Y2=3.33
r221 85 86 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r222 83 129 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.425 $Y=3.33
+ $X2=3.26 $Y2=3.33
r223 83 85 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.425 $Y=3.33
+ $X2=3.6 $Y2=3.33
r224 82 130 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=3.12 $Y2=3.33
r225 82 126 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r226 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r227 79 125 11.3727 $w=1.7e-07 $l=4.75e-07 $layer=LI1_cond $X=1.565 $Y=3.33
+ $X2=1.09 $Y2=3.33
r228 79 81 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=1.565 $Y=3.33
+ $X2=1.68 $Y2=3.33
r229 78 129 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.095 $Y=3.33
+ $X2=3.26 $Y2=3.33
r230 78 81 92.3155 $w=1.68e-07 $l=1.415e-06 $layer=LI1_cond $X=3.095 $Y=3.33
+ $X2=1.68 $Y2=3.33
r231 76 126 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r232 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r233 73 125 11.3727 $w=1.7e-07 $l=4.75e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=1.09 $Y2=3.33
r234 73 75 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.24 $Y2=3.33
r235 71 99 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=7.2 $Y=3.33
+ $X2=7.92 $Y2=3.33
r236 71 95 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=7.2 $Y=3.33
+ $X2=6.96 $Y2=3.33
r237 69 110 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=11.945 $Y=3.33
+ $X2=11.76 $Y2=3.33
r238 69 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.945 $Y=3.33
+ $X2=12.11 $Y2=3.33
r239 68 114 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=12.275 $Y=3.33
+ $X2=12.72 $Y2=3.33
r240 68 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.275 $Y=3.33
+ $X2=12.11 $Y2=3.33
r241 66 94 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=7.025 $Y=3.33
+ $X2=6.96 $Y2=3.33
r242 66 67 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=7.025 $Y=3.33
+ $X2=7.145 $Y2=3.33
r243 65 98 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=7.265 $Y=3.33
+ $X2=7.92 $Y2=3.33
r244 65 67 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=7.265 $Y=3.33
+ $X2=7.145 $Y2=3.33
r245 63 88 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=4.705 $Y=3.33
+ $X2=4.56 $Y2=3.33
r246 63 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.705 $Y=3.33
+ $X2=4.87 $Y2=3.33
r247 62 91 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=5.035 $Y=3.33
+ $X2=5.04 $Y2=3.33
r248 62 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.035 $Y=3.33
+ $X2=4.87 $Y2=3.33
r249 58 61 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=14.12 $Y=1.985
+ $X2=14.12 $Y2=2.815
r250 56 145 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=14.12 $Y=3.245
+ $X2=14.177 $Y2=3.33
r251 56 61 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=14.12 $Y=3.245
+ $X2=14.12 $Y2=2.815
r252 52 55 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=13.17 $Y=1.985
+ $X2=13.17 $Y2=2.815
r253 50 142 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.17 $Y=3.245
+ $X2=13.17 $Y2=3.33
r254 50 55 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=13.17 $Y=3.245
+ $X2=13.17 $Y2=2.815
r255 46 49 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=12.11 $Y=2.105
+ $X2=12.11 $Y2=2.815
r256 44 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.11 $Y=3.245
+ $X2=12.11 $Y2=3.33
r257 44 49 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=12.11 $Y=3.245
+ $X2=12.11 $Y2=2.815
r258 40 132 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=8.412 $Y=3.245
+ $X2=8.412 $Y2=3.33
r259 40 42 28.2091 $w=3.33e-07 $l=8.2e-07 $layer=LI1_cond $X=8.412 $Y=3.245
+ $X2=8.412 $Y2=2.425
r260 36 67 0.135687 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=7.145 $Y=3.245
+ $X2=7.145 $Y2=3.33
r261 36 38 31.9323 $w=2.38e-07 $l=6.65e-07 $layer=LI1_cond $X=7.145 $Y=3.245
+ $X2=7.145 $Y2=2.58
r262 32 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.87 $Y=3.245
+ $X2=4.87 $Y2=3.33
r263 32 34 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=4.87 $Y=3.245
+ $X2=4.87 $Y2=2.835
r264 28 129 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.26 $Y=3.245
+ $X2=3.26 $Y2=3.33
r265 28 30 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.26 $Y=3.245
+ $X2=3.26 $Y2=2.815
r266 9 61 400 $w=1.7e-07 $l=1.07034e-06 $layer=licon1_PDIFF $count=1 $X=13.92
+ $Y=1.84 $X2=14.12 $Y2=2.815
r267 9 58 400 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=1 $X=13.92
+ $Y=1.84 $X2=14.12 $Y2=1.985
r268 8 55 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=13.025
+ $Y=1.84 $X2=13.17 $Y2=2.815
r269 8 52 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=13.025
+ $Y=1.84 $X2=13.17 $Y2=1.985
r270 7 49 600 $w=1.7e-07 $l=3.745e-07 $layer=licon1_PDIFF $count=1 $X=11.875
+ $Y=2.54 $X2=12.11 $Y2=2.815
r271 7 46 300 $w=1.7e-07 $l=5.39861e-07 $layer=licon1_PDIFF $count=2 $X=11.875
+ $Y=2.54 $X2=12.11 $Y2=2.105
r272 6 135 300 $w=1.7e-07 $l=6.22495e-07 $layer=licon1_PDIFF $count=2 $X=10.575
+ $Y=2.54 $X2=11.075 $Y2=2.815
r273 5 42 600 $w=1.7e-07 $l=7.59045e-07 $layer=licon1_PDIFF $count=1 $X=8.27
+ $Y=1.735 $X2=8.415 $Y2=2.425
r274 4 38 600 $w=1.7e-07 $l=3.62319e-07 $layer=licon1_PDIFF $count=1 $X=7.02
+ $Y=2.285 $X2=7.17 $Y2=2.58
r275 3 34 600 $w=1.7e-07 $l=9.47035e-07 $layer=licon1_PDIFF $count=1 $X=4.72
+ $Y=1.96 $X2=4.87 $Y2=2.835
r276 2 30 600 $w=1.7e-07 $l=5.65044e-07 $layer=licon1_PDIFF $count=1 $X=3.11
+ $Y=2.32 $X2=3.26 $Y2=2.815
r277 1 122 150 $w=1.7e-07 $l=8.8955e-07 $layer=licon1_PDIFF $count=4 $X=0.58
+ $Y=2.32 $X2=1.4 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTP_2%A_390_81# 1 2 3 4 5 18 22 25 26 27 28 32 35
+ 37 38 39 40 41 43 45
c156 38 0 1.43931e-19 $X=6.345 $Y=1.285
c157 26 0 1.94423e-19 $X=4.555 $Y=2.52
c158 25 0 1.19423e-19 $X=3.53 $Y=2.33
r159 42 43 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=6.43 $Y=1.37
+ $X2=6.43 $Y2=2.045
r160 40 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.345 $Y=2.13
+ $X2=6.43 $Y2=2.045
r161 40 41 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=6.345 $Y=2.13
+ $X2=6.075 $Y2=2.13
r162 38 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.345 $Y=1.285
+ $X2=6.43 $Y2=1.37
r163 38 39 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=6.345 $Y=1.285
+ $X2=5.975 $Y2=1.285
r164 37 52 3.21189 $w=2.5e-07 $l=1.7e-07 $layer=LI1_cond $X=5.95 $Y=2.385
+ $X2=5.95 $Y2=2.555
r165 36 41 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.95 $Y=2.215
+ $X2=6.075 $Y2=2.13
r166 36 37 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=5.95 $Y=2.215
+ $X2=5.95 $Y2=2.385
r167 35 39 6.81835 $w=1.7e-07 $l=1.23386e-07 $layer=LI1_cond $X=5.887 $Y=1.2
+ $X2=5.975 $Y2=1.285
r168 35 50 12.9922 $w=1.73e-07 $l=2.05e-07 $layer=LI1_cond $X=5.887 $Y=1.2
+ $X2=5.887 $Y2=0.995
r169 30 50 5.54545 $w=1.78e-07 $l=9e-08 $layer=LI1_cond $X=5.885 $Y=0.905
+ $X2=5.885 $Y2=0.995
r170 30 32 5.85354 $w=1.78e-07 $l=9.5e-08 $layer=LI1_cond $X=5.885 $Y=0.905
+ $X2=5.885 $Y2=0.81
r171 28 52 3.74091 $w=1.95e-07 $l=1.57321e-07 $layer=LI1_cond $X=5.825 $Y=2.482
+ $X2=5.95 $Y2=2.555
r172 28 29 67.1142 $w=1.93e-07 $l=1.18e-06 $layer=LI1_cond $X=5.825 $Y=2.482
+ $X2=4.645 $Y2=2.482
r173 27 49 15.7795 $w=4.05e-07 $l=4.82804e-07 $layer=LI1_cond $X=4.25 $Y=2.52
+ $X2=3.83 $Y2=2.655
r174 26 29 5.46269 $w=2.01e-07 $l=1.07331e-07 $layer=LI1_cond $X=4.555 $Y=2.52
+ $X2=4.645 $Y2=2.482
r175 26 27 16.9136 $w=1.98e-07 $l=3.05e-07 $layer=LI1_cond $X=4.555 $Y=2.52
+ $X2=4.25 $Y2=2.52
r176 25 49 9.03704 $w=4.05e-07 $l=4.50694e-07 $layer=LI1_cond $X=3.53 $Y=2.33
+ $X2=3.83 $Y2=2.655
r177 24 46 6.07598 $w=1.7e-07 $l=3.38e-07 $layer=LI1_cond $X=3.53 $Y=1.27
+ $X2=3.53 $Y2=0.932
r178 24 25 69.1551 $w=1.68e-07 $l=1.06e-06 $layer=LI1_cond $X=3.53 $Y=1.27
+ $X2=3.53 $Y2=2.33
r179 23 45 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.425 $Y=2.43
+ $X2=2.26 $Y2=2.43
r180 22 25 6.7671 $w=4.05e-07 $l=1.36015e-07 $layer=LI1_cond $X=3.445 $Y=2.43
+ $X2=3.53 $Y2=2.33
r181 22 23 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=3.445 $Y=2.43
+ $X2=2.425 $Y2=2.43
r182 18 46 23.6232 $w=4.2e-07 $l=8.44373e-07 $layer=LI1_cond $X=2.785 $Y=0.72
+ $X2=3.53 $Y2=0.932
r183 18 20 16.1342 $w=2.48e-07 $l=3.5e-07 $layer=LI1_cond $X=2.785 $Y=0.72
+ $X2=2.435 $Y2=0.72
r184 5 52 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=5.765
+ $Y=2.285 $X2=5.91 $Y2=2.495
r185 4 49 300 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=2 $X=3.68
+ $Y=2.32 $X2=3.83 $Y2=2.475
r186 3 45 300 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=2 $X=2.12
+ $Y=2.32 $X2=2.26 $Y2=2.475
r187 2 32 182 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_NDIFF $count=1 $X=5.755
+ $Y=0.595 $X2=5.88 $Y2=0.81
r188 1 20 182 $w=1.7e-07 $l=6.07124e-07 $layer=licon1_NDIFF $count=1 $X=1.95
+ $Y=0.405 $X2=2.435 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTP_2%Q 1 2 9 13 14 15 29
r21 20 29 1.74613 $w=3.28e-07 $l=5e-08 $layer=LI1_cond $X=13.69 $Y=1.245
+ $X2=13.69 $Y2=1.295
r22 15 31 3.97298 $w=3.28e-07 $l=9.8e-08 $layer=LI1_cond $X=13.69 $Y=1.312
+ $X2=13.69 $Y2=1.41
r23 15 29 0.593683 $w=3.28e-07 $l=1.7e-08 $layer=LI1_cond $X=13.69 $Y=1.312
+ $X2=13.69 $Y2=1.295
r24 15 20 0.628605 $w=3.28e-07 $l=1.8e-08 $layer=LI1_cond $X=13.69 $Y=1.227
+ $X2=13.69 $Y2=1.245
r25 14 15 10.5466 $w=3.28e-07 $l=3.02e-07 $layer=LI1_cond $X=13.69 $Y=0.925
+ $X2=13.69 $Y2=1.227
r26 13 14 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=13.69 $Y=0.515
+ $X2=13.69 $Y2=0.925
r27 9 11 36.7895 $w=2.58e-07 $l=8.3e-07 $layer=LI1_cond $X=13.655 $Y=1.985
+ $X2=13.655 $Y2=2.815
r28 9 31 25.4867 $w=2.58e-07 $l=5.75e-07 $layer=LI1_cond $X=13.655 $Y=1.985
+ $X2=13.655 $Y2=1.41
r29 2 11 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=13.47
+ $Y=1.84 $X2=13.62 $Y2=2.815
r30 2 9 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=13.47
+ $Y=1.84 $X2=13.62 $Y2=1.985
r31 1 13 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=13.55
+ $Y=0.37 $X2=13.69 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTP_2%VGND 1 2 3 4 5 6 7 8 27 31 35 39 43 47 49
+ 51 54 55 57 58 59 61 76 80 85 90 95 101 105 111 114 117 121
c139 121 0 3.56444e-20 $X=14.16 $Y=0
c140 31 0 1.49819e-19 $X=3.76 $Y=0.565
r141 120 121 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.16 $Y=0
+ $X2=14.16 $Y2=0
r142 117 118 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=0
+ $X2=13.2 $Y2=0
r143 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r144 111 112 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=10.8 $Y=0
+ $X2=10.8 $Y2=0
r145 105 108 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=7.595 $Y=0
+ $X2=7.595 $Y2=0.325
r146 105 106 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r147 101 102 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0
+ $X2=0.72 $Y2=0
r148 99 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=0
+ $X2=14.16 $Y2=0
r149 99 118 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=0
+ $X2=13.2 $Y2=0
r150 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=0
+ $X2=13.68 $Y2=0
r151 96 117 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.345 $Y=0
+ $X2=13.22 $Y2=0
r152 96 98 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=13.345 $Y=0
+ $X2=13.68 $Y2=0
r153 95 120 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=14.035 $Y=0
+ $X2=14.217 $Y2=0
r154 95 98 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=14.035 $Y=0
+ $X2=13.68 $Y2=0
r155 94 118 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=0
+ $X2=13.2 $Y2=0
r156 94 115 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=0
+ $X2=12.24 $Y2=0
r157 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r158 91 114 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.435 $Y=0
+ $X2=12.27 $Y2=0
r159 91 93 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=12.435 $Y=0
+ $X2=12.72 $Y2=0
r160 90 117 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.095 $Y=0
+ $X2=13.22 $Y2=0
r161 90 93 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=13.095 $Y=0
+ $X2=12.72 $Y2=0
r162 89 115 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=12.24 $Y2=0
r163 89 112 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=10.8 $Y2=0
r164 88 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r165 86 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.085 $Y=0
+ $X2=10.92 $Y2=0
r166 86 88 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=11.085 $Y=0
+ $X2=11.76 $Y2=0
r167 85 114 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.105 $Y=0
+ $X2=12.27 $Y2=0
r168 85 88 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=12.105 $Y=0
+ $X2=11.76 $Y2=0
r169 84 112 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=7.92 $Y=0
+ $X2=10.8 $Y2=0
r170 84 106 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0
+ $X2=7.44 $Y2=0
r171 83 84 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r172 81 105 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.76 $Y=0
+ $X2=7.595 $Y2=0
r173 81 83 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=7.76 $Y=0 $X2=7.92
+ $Y2=0
r174 80 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.755 $Y=0
+ $X2=10.92 $Y2=0
r175 80 83 184.957 $w=1.68e-07 $l=2.835e-06 $layer=LI1_cond $X=10.755 $Y=0
+ $X2=7.92 $Y2=0
r176 78 79 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r177 76 105 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.43 $Y=0
+ $X2=7.595 $Y2=0
r178 76 78 155.925 $w=1.68e-07 $l=2.39e-06 $layer=LI1_cond $X=7.43 $Y=0 $X2=5.04
+ $Y2=0
r179 75 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r180 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r181 72 75 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r182 71 72 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r183 69 72 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=3.6
+ $Y2=0
r184 69 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r185 68 71 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=3.6
+ $Y2=0
r186 68 69 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r187 66 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.875 $Y=0
+ $X2=0.71 $Y2=0
r188 66 68 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=1.2
+ $Y2=0
r189 64 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0
+ $X2=0.72 $Y2=0
r190 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r191 61 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.545 $Y=0
+ $X2=0.71 $Y2=0
r192 61 63 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0
+ $X2=0.24 $Y2=0
r193 59 106 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=7.2 $Y=0
+ $X2=7.44 $Y2=0
r194 59 79 0.602067 $w=4.9e-07 $l=2.16e-06 $layer=MET1_cond $X=7.2 $Y=0 $X2=5.04
+ $Y2=0
r195 57 74 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=4.705 $Y=0
+ $X2=4.56 $Y2=0
r196 57 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.705 $Y=0 $X2=4.87
+ $Y2=0
r197 56 78 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=5.035 $Y=0 $X2=5.04
+ $Y2=0
r198 56 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.035 $Y=0 $X2=4.87
+ $Y2=0
r199 54 71 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=3.61 $Y=0 $X2=3.6
+ $Y2=0
r200 54 55 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.61 $Y=0 $X2=3.745
+ $Y2=0
r201 53 74 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.88 $Y=0 $X2=4.56
+ $Y2=0
r202 53 55 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.88 $Y=0 $X2=3.745
+ $Y2=0
r203 49 120 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=14.16 $Y=0.085
+ $X2=14.217 $Y2=0
r204 49 51 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=14.16 $Y=0.085
+ $X2=14.16 $Y2=0.515
r205 45 117 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=13.22 $Y=0.085
+ $X2=13.22 $Y2=0
r206 45 47 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=13.22 $Y=0.085
+ $X2=13.22 $Y2=0.515
r207 41 114 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.27 $Y=0.085
+ $X2=12.27 $Y2=0
r208 41 43 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=12.27 $Y=0.085
+ $X2=12.27 $Y2=0.515
r209 37 111 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.92 $Y=0.085
+ $X2=10.92 $Y2=0
r210 37 39 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=10.92 $Y=0.085
+ $X2=10.92 $Y2=0.58
r211 33 58 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.87 $Y=0.085
+ $X2=4.87 $Y2=0
r212 33 35 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=4.87 $Y=0.085
+ $X2=4.87 $Y2=0.625
r213 29 55 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.745 $Y=0.085
+ $X2=3.745 $Y2=0
r214 29 31 20.4879 $w=2.68e-07 $l=4.8e-07 $layer=LI1_cond $X=3.745 $Y=0.085
+ $X2=3.745 $Y2=0.565
r215 25 101 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0
r216 25 27 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0.555
r217 8 51 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=13.98
+ $Y=0.37 $X2=14.12 $Y2=0.515
r218 7 47 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=13.115
+ $Y=0.37 $X2=13.26 $Y2=0.515
r219 6 43 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=12.125
+ $Y=0.37 $X2=12.27 $Y2=0.515
r220 5 39 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=10.78
+ $Y=0.37 $X2=10.92 $Y2=0.58
r221 4 108 182 $w=1.7e-07 $l=3.63731e-07 $layer=licon1_NDIFF $count=1 $X=7.375
+ $Y=0.595 $X2=7.595 $Y2=0.325
r222 3 35 182 $w=1.7e-07 $l=2.14476e-07 $layer=licon1_NDIFF $count=1 $X=4.67
+ $Y=0.595 $X2=4.87 $Y2=0.625
r223 2 31 182 $w=1.7e-07 $l=2.52636e-07 $layer=licon1_NDIFF $count=1 $X=3.575
+ $Y=0.405 $X2=3.76 $Y2=0.565
r224 1 27 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTP_2%noxref_24 1 2 7 11 13
r26 13 16 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=1.27 $Y=0.34
+ $X2=1.27 $Y2=0.55
r27 9 11 6.72258 $w=2.38e-07 $l=1.4e-07 $layer=LI1_cond $X=3.31 $Y=0.425
+ $X2=3.31 $Y2=0.565
r28 8 13 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.435 $Y=0.34
+ $X2=1.27 $Y2=0.34
r29 7 9 7.07814 $w=1.7e-07 $l=1.56844e-07 $layer=LI1_cond $X=3.19 $Y=0.34
+ $X2=3.31 $Y2=0.425
r30 7 8 114.497 $w=1.68e-07 $l=1.755e-06 $layer=LI1_cond $X=3.19 $Y=0.34
+ $X2=1.435 $Y2=0.34
r31 2 11 182 $w=1.7e-07 $l=2.26274e-07 $layer=licon1_NDIFF $count=1 $X=3.115
+ $Y=0.405 $X2=3.275 $Y2=0.565
r32 1 16 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=1.125
+ $Y=0.405 $X2=1.27 $Y2=0.55
.ends

