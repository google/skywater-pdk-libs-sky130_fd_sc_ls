* File: sky130_fd_sc_ls__clkinv_8.pex.spice
* Created: Wed Sep  2 10:59:04 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__CLKINV_8%A 3 5 7 8 10 11 13 14 16 17 19 22 24 26 29
+ 31 33 36 38 40 43 45 47 50 52 54 57 59 61 62 64 67 69 70 71 72 73 74 75 106
+ 107
r200 107 108 1.98626 $w=3.64e-07 $l=1.5e-08 $layer=POLY_cond $X=5.73 $Y=1.557
+ $X2=5.745 $Y2=1.557
r201 105 107 23.8352 $w=3.64e-07 $l=1.8e-07 $layer=POLY_cond $X=5.55 $Y=1.557
+ $X2=5.73 $Y2=1.557
r202 105 106 19.3707 $w=1.7e-07 $l=1.275e-06 $layer=licon1_POLY $count=7 $X=5.55
+ $Y=1.515 $X2=5.55 $Y2=1.515
r203 103 105 35.7527 $w=3.64e-07 $l=2.7e-07 $layer=POLY_cond $X=5.28 $Y=1.557
+ $X2=5.55 $Y2=1.557
r204 102 103 4.63462 $w=3.64e-07 $l=3.5e-08 $layer=POLY_cond $X=5.245 $Y=1.557
+ $X2=5.28 $Y2=1.557
r205 101 102 61.5742 $w=3.64e-07 $l=4.65e-07 $layer=POLY_cond $X=4.78 $Y=1.557
+ $X2=5.245 $Y2=1.557
r206 100 101 13.9038 $w=3.64e-07 $l=1.05e-07 $layer=POLY_cond $X=4.675 $Y=1.557
+ $X2=4.78 $Y2=1.557
r207 99 100 45.6841 $w=3.64e-07 $l=3.45e-07 $layer=POLY_cond $X=4.33 $Y=1.557
+ $X2=4.675 $Y2=1.557
r208 98 99 11.2555 $w=3.64e-07 $l=8.5e-08 $layer=POLY_cond $X=4.245 $Y=1.557
+ $X2=4.33 $Y2=1.557
r209 97 98 54.9533 $w=3.64e-07 $l=4.15e-07 $layer=POLY_cond $X=3.83 $Y=1.557
+ $X2=4.245 $Y2=1.557
r210 96 97 20.5247 $w=3.64e-07 $l=1.55e-07 $layer=POLY_cond $X=3.675 $Y=1.557
+ $X2=3.83 $Y2=1.557
r211 95 96 39.0632 $w=3.64e-07 $l=2.95e-07 $layer=POLY_cond $X=3.38 $Y=1.557
+ $X2=3.675 $Y2=1.557
r212 94 95 17.8764 $w=3.64e-07 $l=1.35e-07 $layer=POLY_cond $X=3.245 $Y=1.557
+ $X2=3.38 $Y2=1.557
r213 93 94 48.3324 $w=3.64e-07 $l=3.65e-07 $layer=POLY_cond $X=2.88 $Y=1.557
+ $X2=3.245 $Y2=1.557
r214 92 93 27.1456 $w=3.64e-07 $l=2.05e-07 $layer=POLY_cond $X=2.675 $Y=1.557
+ $X2=2.88 $Y2=1.557
r215 91 92 32.4423 $w=3.64e-07 $l=2.45e-07 $layer=POLY_cond $X=2.43 $Y=1.557
+ $X2=2.675 $Y2=1.557
r216 90 91 66.2088 $w=3.64e-07 $l=5e-07 $layer=POLY_cond $X=1.93 $Y=1.557
+ $X2=2.43 $Y2=1.557
r217 89 90 59.5879 $w=3.64e-07 $l=4.5e-07 $layer=POLY_cond $X=1.48 $Y=1.557
+ $X2=1.93 $Y2=1.557
r218 88 89 66.2088 $w=3.64e-07 $l=5e-07 $layer=POLY_cond $X=0.98 $Y=1.557
+ $X2=1.48 $Y2=1.557
r219 86 88 25.1593 $w=3.64e-07 $l=1.9e-07 $layer=POLY_cond $X=0.79 $Y=1.557
+ $X2=0.98 $Y2=1.557
r220 86 87 19.3707 $w=1.7e-07 $l=1.275e-06 $layer=licon1_POLY $count=7 $X=0.79
+ $Y=1.515 $X2=0.79 $Y2=1.515
r221 84 86 34.4286 $w=3.64e-07 $l=2.6e-07 $layer=POLY_cond $X=0.53 $Y=1.557
+ $X2=0.79 $Y2=1.557
r222 83 84 1.98626 $w=3.64e-07 $l=1.5e-08 $layer=POLY_cond $X=0.515 $Y=1.557
+ $X2=0.53 $Y2=1.557
r223 75 106 39.3975 $w=4.28e-07 $l=1.47e-06 $layer=LI1_cond $X=4.08 $Y=1.565
+ $X2=5.55 $Y2=1.565
r224 74 75 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=3.6 $Y=1.565
+ $X2=4.08 $Y2=1.565
r225 73 74 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=3.12 $Y=1.565
+ $X2=3.6 $Y2=1.565
r226 72 73 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=2.64 $Y=1.565
+ $X2=3.12 $Y2=1.565
r227 71 72 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=2.16 $Y=1.565
+ $X2=2.64 $Y2=1.565
r228 70 71 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=1.565
+ $X2=2.16 $Y2=1.565
r229 69 70 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.565
+ $X2=1.68 $Y2=1.565
r230 69 87 10.9884 $w=4.28e-07 $l=4.1e-07 $layer=LI1_cond $X=1.2 $Y=1.565
+ $X2=0.79 $Y2=1.565
r231 65 108 23.572 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.745 $Y=1.35
+ $X2=5.745 $Y2=1.557
r232 65 67 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=5.745 $Y=1.35
+ $X2=5.745 $Y2=0.61
r233 62 107 23.572 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=5.73 $Y=1.765
+ $X2=5.73 $Y2=1.557
r234 62 64 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.73 $Y=1.765
+ $X2=5.73 $Y2=2.4
r235 59 103 23.572 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=5.28 $Y=1.765
+ $X2=5.28 $Y2=1.557
r236 59 61 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.28 $Y=1.765
+ $X2=5.28 $Y2=2.4
r237 55 102 23.572 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.245 $Y=1.35
+ $X2=5.245 $Y2=1.557
r238 55 57 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=5.245 $Y=1.35
+ $X2=5.245 $Y2=0.61
r239 52 101 23.572 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=4.78 $Y=1.765
+ $X2=4.78 $Y2=1.557
r240 52 54 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.78 $Y=1.765
+ $X2=4.78 $Y2=2.4
r241 48 100 23.572 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.675 $Y=1.35
+ $X2=4.675 $Y2=1.557
r242 48 50 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=4.675 $Y=1.35
+ $X2=4.675 $Y2=0.61
r243 45 99 23.572 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=4.33 $Y=1.765
+ $X2=4.33 $Y2=1.557
r244 45 47 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.33 $Y=1.765
+ $X2=4.33 $Y2=2.4
r245 41 98 23.572 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.245 $Y=1.35
+ $X2=4.245 $Y2=1.557
r246 41 43 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=4.245 $Y=1.35
+ $X2=4.245 $Y2=0.61
r247 38 97 23.572 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.83 $Y=1.765
+ $X2=3.83 $Y2=1.557
r248 38 40 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.83 $Y=1.765
+ $X2=3.83 $Y2=2.4
r249 34 96 23.572 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.675 $Y=1.35
+ $X2=3.675 $Y2=1.557
r250 34 36 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=3.675 $Y=1.35
+ $X2=3.675 $Y2=0.61
r251 31 95 23.572 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.38 $Y=1.765
+ $X2=3.38 $Y2=1.557
r252 31 33 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.38 $Y=1.765
+ $X2=3.38 $Y2=2.4
r253 27 94 23.572 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.245 $Y=1.35
+ $X2=3.245 $Y2=1.557
r254 27 29 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=3.245 $Y=1.35
+ $X2=3.245 $Y2=0.61
r255 24 93 23.572 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.88 $Y=1.765
+ $X2=2.88 $Y2=1.557
r256 24 26 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.88 $Y=1.765
+ $X2=2.88 $Y2=2.4
r257 20 92 23.572 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.675 $Y=1.35
+ $X2=2.675 $Y2=1.557
r258 20 22 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=2.675 $Y=1.35
+ $X2=2.675 $Y2=0.61
r259 17 91 23.572 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.43 $Y=1.765
+ $X2=2.43 $Y2=1.557
r260 17 19 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.43 $Y=1.765
+ $X2=2.43 $Y2=2.4
r261 14 90 23.572 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.93 $Y=1.765
+ $X2=1.93 $Y2=1.557
r262 14 16 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.93 $Y=1.765
+ $X2=1.93 $Y2=2.4
r263 11 89 23.572 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.48 $Y=1.765
+ $X2=1.48 $Y2=1.557
r264 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.48 $Y=1.765
+ $X2=1.48 $Y2=2.4
r265 8 88 23.572 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.98 $Y=1.765
+ $X2=0.98 $Y2=1.557
r266 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.98 $Y=1.765
+ $X2=0.98 $Y2=2.4
r267 5 84 23.572 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.53 $Y=1.765
+ $X2=0.53 $Y2=1.557
r268 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.53 $Y=1.765
+ $X2=0.53 $Y2=2.4
r269 1 83 23.572 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.515 $Y=1.35
+ $X2=0.515 $Y2=1.557
r270 1 3 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=0.515 $Y=1.35
+ $X2=0.515 $Y2=0.61
.ends

.subckt PM_SKY130_FD_SC_LS__CLKINV_8%VPWR 1 2 3 4 5 6 7 22 24 26 30 34 38 42 46
+ 48 50 52 54 59 64 69 74 83 86 89 92 95 99
r98 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r99 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r100 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r101 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r102 83 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r103 81 84 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r104 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r105 78 99 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33 $X2=6
+ $Y2=3.33
r106 78 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=5.04 $Y2=3.33
r107 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r108 75 95 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.17 $Y=3.33
+ $X2=5.045 $Y2=3.33
r109 75 77 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=5.17 $Y=3.33
+ $X2=5.52 $Y2=3.33
r110 74 98 4.0045 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=5.87 $Y=3.33
+ $X2=6.055 $Y2=3.33
r111 74 77 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=5.87 $Y=3.33
+ $X2=5.52 $Y2=3.33
r112 73 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r113 73 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r114 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r115 70 92 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.22 $Y=3.33
+ $X2=4.095 $Y2=3.33
r116 70 72 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=4.22 $Y=3.33
+ $X2=4.56 $Y2=3.33
r117 69 95 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.92 $Y=3.33
+ $X2=5.045 $Y2=3.33
r118 69 72 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=4.92 $Y=3.33
+ $X2=4.56 $Y2=3.33
r119 68 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r120 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r121 65 89 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.27 $Y=3.33
+ $X2=3.145 $Y2=3.33
r122 65 67 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=3.27 $Y=3.33
+ $X2=3.6 $Y2=3.33
r123 64 92 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.97 $Y=3.33
+ $X2=4.095 $Y2=3.33
r124 64 67 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.97 $Y=3.33 $X2=3.6
+ $Y2=3.33
r125 63 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r126 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r127 60 86 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.32 $Y=3.33
+ $X2=2.195 $Y2=3.33
r128 60 62 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2.32 $Y=3.33
+ $X2=2.64 $Y2=3.33
r129 59 89 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.02 $Y=3.33
+ $X2=3.145 $Y2=3.33
r130 59 62 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=3.02 $Y=3.33
+ $X2=2.64 $Y2=3.33
r131 58 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r132 58 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r133 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r134 55 83 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.37 $Y=3.33
+ $X2=1.245 $Y2=3.33
r135 55 57 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1.37 $Y=3.33
+ $X2=1.68 $Y2=3.33
r136 54 86 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.07 $Y=3.33
+ $X2=2.195 $Y2=3.33
r137 54 57 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=2.07 $Y=3.33
+ $X2=1.68 $Y2=3.33
r138 52 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r139 52 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r140 52 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r141 48 98 3.13866 $w=2.5e-07 $l=1.11018e-07 $layer=LI1_cond $X=5.995 $Y=3.245
+ $X2=6.055 $Y2=3.33
r142 48 50 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=5.995 $Y=3.245
+ $X2=5.995 $Y2=2.455
r143 44 95 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.045 $Y=3.245
+ $X2=5.045 $Y2=3.33
r144 44 46 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=5.045 $Y=3.245
+ $X2=5.045 $Y2=2.455
r145 40 92 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.095 $Y=3.245
+ $X2=4.095 $Y2=3.33
r146 40 42 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=4.095 $Y=3.245
+ $X2=4.095 $Y2=2.455
r147 36 89 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.145 $Y=3.245
+ $X2=3.145 $Y2=3.33
r148 36 38 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=3.145 $Y=3.245
+ $X2=3.145 $Y2=2.455
r149 32 86 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.195 $Y=3.245
+ $X2=2.195 $Y2=3.33
r150 32 34 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=2.195 $Y=3.245
+ $X2=2.195 $Y2=2.455
r151 28 83 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.245 $Y=3.245
+ $X2=1.245 $Y2=3.33
r152 28 30 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=1.245 $Y=3.245
+ $X2=1.245 $Y2=2.455
r153 27 80 4.23679 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=0.39 $Y=3.33
+ $X2=0.195 $Y2=3.33
r154 26 83 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.12 $Y=3.33
+ $X2=1.245 $Y2=3.33
r155 26 27 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.12 $Y=3.33
+ $X2=0.39 $Y2=3.33
r156 22 80 3.08525 $w=2.75e-07 $l=1.09864e-07 $layer=LI1_cond $X=0.252 $Y=3.245
+ $X2=0.195 $Y2=3.33
r157 22 24 33.1065 $w=2.73e-07 $l=7.9e-07 $layer=LI1_cond $X=0.252 $Y=3.245
+ $X2=0.252 $Y2=2.455
r158 7 50 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=5.805
+ $Y=1.84 $X2=5.955 $Y2=2.455
r159 6 46 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=4.855
+ $Y=1.84 $X2=5.005 $Y2=2.455
r160 5 42 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=3.905
+ $Y=1.84 $X2=4.055 $Y2=2.455
r161 4 38 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=2.955
+ $Y=1.84 $X2=3.105 $Y2=2.455
r162 3 34 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=2.005
+ $Y=1.84 $X2=2.155 $Y2=2.455
r163 2 30 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=1.055
+ $Y=1.84 $X2=1.205 $Y2=2.455
r164 1 24 300 $w=1.7e-07 $l=6.8815e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.84 $X2=0.29 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_LS__CLKINV_8%Y 1 2 3 4 5 6 7 8 9 10 32 35 37 38 39 40 43
+ 45 49 51 53 57 61 63 65 69 73 75 77 81 85 87 89 99 102 104 105 107 108 110 111
+ 113 116
r193 115 116 32.8196 $w=2.28e-07 $l=6.55e-07 $layer=LI1_cond $X=6 $Y=1.95 $X2=6
+ $Y2=1.295
r194 114 116 5.76222 $w=2.28e-07 $l=1.15e-07 $layer=LI1_cond $X=6 $Y=1.18 $X2=6
+ $Y2=1.295
r195 101 102 10.933 $w=7.18e-07 $l=1.65e-07 $layer=LI1_cond $X=2.46 $Y=0.82
+ $X2=2.625 $Y2=0.82
r196 94 97 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.37 $Y=2.035
+ $X2=0.755 $Y2=2.035
r197 90 113 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.67 $Y=2.035
+ $X2=5.505 $Y2=2.035
r198 89 115 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=5.885 $Y=2.035
+ $X2=6 $Y2=1.95
r199 89 90 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=5.885 $Y=2.035
+ $X2=5.67 $Y2=2.035
r200 88 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.625 $Y=1.095
+ $X2=5.46 $Y2=1.095
r201 87 114 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=5.885 $Y=1.095
+ $X2=6 $Y2=1.18
r202 87 88 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=5.885 $Y=1.095
+ $X2=5.625 $Y2=1.095
r203 83 113 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.505 $Y=2.12
+ $X2=5.505 $Y2=2.035
r204 83 85 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=5.505 $Y=2.12
+ $X2=5.505 $Y2=2.815
r205 79 111 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.46 $Y=1.01
+ $X2=5.46 $Y2=1.095
r206 79 81 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=5.46 $Y=1.01 $X2=5.46
+ $Y2=0.61
r207 78 110 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.72 $Y=2.035
+ $X2=4.555 $Y2=2.035
r208 77 113 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.34 $Y=2.035
+ $X2=5.505 $Y2=2.035
r209 77 78 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=5.34 $Y=2.035
+ $X2=4.72 $Y2=2.035
r210 76 108 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.625 $Y=1.095
+ $X2=4.46 $Y2=1.095
r211 75 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.295 $Y=1.095
+ $X2=5.46 $Y2=1.095
r212 75 76 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.295 $Y=1.095
+ $X2=4.625 $Y2=1.095
r213 71 110 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.555 $Y=2.12
+ $X2=4.555 $Y2=2.035
r214 71 73 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=4.555 $Y=2.12
+ $X2=4.555 $Y2=2.815
r215 67 108 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.46 $Y=1.01
+ $X2=4.46 $Y2=1.095
r216 67 69 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=4.46 $Y=1.01 $X2=4.46
+ $Y2=0.61
r217 66 107 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.77 $Y=2.035
+ $X2=3.605 $Y2=2.035
r218 65 110 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.39 $Y=2.035
+ $X2=4.555 $Y2=2.035
r219 65 66 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=4.39 $Y=2.035
+ $X2=3.77 $Y2=2.035
r220 64 105 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.625 $Y=1.095
+ $X2=3.46 $Y2=1.095
r221 63 108 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.295 $Y=1.095
+ $X2=4.46 $Y2=1.095
r222 63 64 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.295 $Y=1.095
+ $X2=3.625 $Y2=1.095
r223 59 107 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.605 $Y=2.12
+ $X2=3.605 $Y2=2.035
r224 59 61 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=3.605 $Y=2.12
+ $X2=3.605 $Y2=2.815
r225 55 105 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.46 $Y=1.01
+ $X2=3.46 $Y2=1.095
r226 55 57 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=3.46 $Y=1.01 $X2=3.46
+ $Y2=0.61
r227 54 104 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.82 $Y=2.035
+ $X2=2.655 $Y2=2.035
r228 53 107 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.44 $Y=2.035
+ $X2=3.605 $Y2=2.035
r229 53 54 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=3.44 $Y=2.035
+ $X2=2.82 $Y2=2.035
r230 51 105 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.295 $Y=1.095
+ $X2=3.46 $Y2=1.095
r231 51 102 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.295 $Y=1.095
+ $X2=2.625 $Y2=1.095
r232 47 104 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.655 $Y=2.12
+ $X2=2.655 $Y2=2.035
r233 47 49 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=2.655 $Y=2.12
+ $X2=2.655 $Y2=2.815
r234 46 99 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.87 $Y=2.035
+ $X2=1.705 $Y2=2.035
r235 45 104 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.49 $Y=2.035
+ $X2=2.655 $Y2=2.035
r236 45 46 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=2.49 $Y=2.035
+ $X2=1.87 $Y2=2.035
r237 41 99 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.705 $Y=2.12
+ $X2=1.705 $Y2=2.035
r238 41 43 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=1.705 $Y=2.12
+ $X2=1.705 $Y2=2.815
r239 40 93 4.93733 $w=7.2e-07 $l=1.95e-07 $layer=LI1_cond $X=0.975 $Y=0.82
+ $X2=0.78 $Y2=0.82
r240 39 101 3.23938 $w=7.18e-07 $l=1.95e-07 $layer=LI1_cond $X=2.265 $Y=0.82
+ $X2=2.46 $Y2=0.82
r241 39 40 21.4297 $w=7.18e-07 $l=1.29e-06 $layer=LI1_cond $X=2.265 $Y=0.82
+ $X2=0.975 $Y2=0.82
r242 38 97 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=0.92 $Y=2.035
+ $X2=0.755 $Y2=2.035
r243 37 99 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.54 $Y=2.035
+ $X2=1.705 $Y2=2.035
r244 37 38 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=1.54 $Y=2.035
+ $X2=0.92 $Y2=2.035
r245 35 97 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=0.755 $Y=2.815
+ $X2=0.755 $Y2=2.12
r246 32 94 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.37 $Y=1.95
+ $X2=0.37 $Y2=2.035
r247 31 93 10.9693 $w=4.56e-07 $l=5.61872e-07 $layer=LI1_cond $X=0.37 $Y=1.18
+ $X2=0.78 $Y2=0.82
r248 31 32 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=0.37 $Y=1.18
+ $X2=0.37 $Y2=1.95
r249 10 113 400 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=5.355
+ $Y=1.84 $X2=5.505 $Y2=2.035
r250 10 85 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=5.355
+ $Y=1.84 $X2=5.505 $Y2=2.815
r251 9 110 400 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=4.405
+ $Y=1.84 $X2=4.555 $Y2=2.035
r252 9 73 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=4.405
+ $Y=1.84 $X2=4.555 $Y2=2.815
r253 8 107 400 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=3.455
+ $Y=1.84 $X2=3.605 $Y2=2.035
r254 8 61 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=3.455
+ $Y=1.84 $X2=3.605 $Y2=2.815
r255 7 104 400 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=2.505
+ $Y=1.84 $X2=2.655 $Y2=2.035
r256 7 49 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.505
+ $Y=1.84 $X2=2.655 $Y2=2.815
r257 6 99 400 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=1.555
+ $Y=1.84 $X2=1.705 $Y2=2.035
r258 6 43 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.555
+ $Y=1.84 $X2=1.705 $Y2=2.815
r259 5 97 400 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=0.605
+ $Y=1.84 $X2=0.755 $Y2=2.035
r260 5 35 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=0.605
+ $Y=1.84 $X2=0.755 $Y2=2.815
r261 4 81 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=5.32
+ $Y=0.4 $X2=5.46 $Y2=0.61
r262 3 69 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.32
+ $Y=0.4 $X2=4.46 $Y2=0.61
r263 2 57 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.32
+ $Y=0.4 $X2=3.46 $Y2=0.61
r264 1 101 72.8 $w=1.7e-07 $l=1.97931e-06 $layer=licon1_NDIFF $count=2 $X=0.59
+ $Y=0.4 $X2=2.46 $Y2=0.625
r265 1 93 72.8 $w=1.7e-07 $l=3.05573e-07 $layer=licon1_NDIFF $count=2 $X=0.59
+ $Y=0.4 $X2=0.78 $Y2=0.625
.ends

.subckt PM_SKY130_FD_SC_LS__CLKINV_8%VGND 1 2 3 4 5 16 18 22 26 30 32 34 37 38
+ 40 41 42 54 58 67 71
r55 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r56 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r57 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r58 62 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r59 62 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r60 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r61 59 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.125 $Y=0 $X2=4.96
+ $Y2=0
r62 59 61 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=5.125 $Y=0 $X2=5.52
+ $Y2=0
r63 58 70 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=5.795 $Y=0 $X2=6.017
+ $Y2=0
r64 58 61 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=5.795 $Y=0 $X2=5.52
+ $Y2=0
r65 57 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r66 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r67 54 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.795 $Y=0 $X2=4.96
+ $Y2=0
r68 54 56 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=4.795 $Y=0 $X2=4.56
+ $Y2=0
r69 53 57 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r70 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r71 49 50 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r72 47 50 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=0.72 $Y=0 $X2=2.64
+ $Y2=0
r73 47 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r74 46 49 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.72 $Y=0 $X2=2.64
+ $Y2=0
r75 46 47 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r76 44 64 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.222
+ $Y2=0
r77 44 46 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.72
+ $Y2=0
r78 42 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r79 42 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r80 40 52 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=3.795 $Y=0 $X2=3.6
+ $Y2=0
r81 40 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.795 $Y=0 $X2=3.96
+ $Y2=0
r82 39 56 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=4.125 $Y=0 $X2=4.56
+ $Y2=0
r83 39 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.125 $Y=0 $X2=3.96
+ $Y2=0
r84 37 49 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=2.795 $Y=0 $X2=2.64
+ $Y2=0
r85 37 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.795 $Y=0 $X2=2.96
+ $Y2=0
r86 36 52 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=3.125 $Y=0 $X2=3.6
+ $Y2=0
r87 36 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.125 $Y=0 $X2=2.96
+ $Y2=0
r88 32 70 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=5.96 $Y=0.085
+ $X2=6.017 $Y2=0
r89 32 34 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=5.96 $Y=0.085
+ $X2=5.96 $Y2=0.61
r90 28 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.96 $Y=0.085
+ $X2=4.96 $Y2=0
r91 28 30 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=4.96 $Y=0.085
+ $X2=4.96 $Y2=0.61
r92 24 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.96 $Y=0.085
+ $X2=3.96 $Y2=0
r93 24 26 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=3.96 $Y=0.085
+ $X2=3.96 $Y2=0.61
r94 20 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.96 $Y=0.085
+ $X2=2.96 $Y2=0
r95 20 22 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=2.96 $Y=0.085
+ $X2=2.96 $Y2=0.61
r96 16 64 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.222 $Y2=0
r97 16 18 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.28 $Y2=0.61
r98 5 34 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=5.82
+ $Y=0.4 $X2=5.96 $Y2=0.61
r99 4 30 182 $w=1.7e-07 $l=2.96985e-07 $layer=licon1_NDIFF $count=1 $X=4.75
+ $Y=0.4 $X2=4.96 $Y2=0.61
r100 3 26 182 $w=1.7e-07 $l=2.96985e-07 $layer=licon1_NDIFF $count=1 $X=3.75
+ $Y=0.4 $X2=3.96 $Y2=0.61
r101 2 22 182 $w=1.7e-07 $l=2.96985e-07 $layer=licon1_NDIFF $count=1 $X=2.75
+ $Y=0.4 $X2=2.96 $Y2=0.61
r102 1 18 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.4 $X2=0.28 $Y2=0.61
.ends

