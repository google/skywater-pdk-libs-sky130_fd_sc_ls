# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ls__a2bb2o_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ls__a2bb2o_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1_N
    ANTENNAGATEAREA  0.232500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.070000 1.180000 1.335000 1.620000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.232500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.545000 1.180000 1.850000 1.620000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485000 0.255000 4.195000 0.670000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.875000 1.450000 3.235000 1.780000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.504100 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.420000 0.590000 1.150000 ;
        RECT 0.125000 1.150000 0.295000 1.820000 ;
        RECT 0.125000 1.820000 0.560000 2.980000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.465000  1.320000 0.900000 1.650000 ;
      RECT 0.730000  1.650000 0.900000 1.790000 ;
      RECT 0.730000  1.790000 2.190000 1.960000 ;
      RECT 0.760000  2.130000 1.090000 3.245000 ;
      RECT 0.770000  0.085000 1.100000 1.010000 ;
      RECT 1.285000  0.255000 2.595000 0.520000 ;
      RECT 1.285000  0.520000 1.590000 1.010000 ;
      RECT 1.325000  1.960000 1.495000 2.905000 ;
      RECT 1.325000  2.905000 2.515000 3.075000 ;
      RECT 1.665000  2.130000 2.530000 2.300000 ;
      RECT 1.665000  2.300000 1.995000 2.735000 ;
      RECT 1.760000  0.690000 2.935000 0.860000 ;
      RECT 2.020000  1.030000 2.900000 1.210000 ;
      RECT 2.020000  1.210000 2.190000 1.790000 ;
      RECT 2.185000  2.470000 2.515000 2.905000 ;
      RECT 2.360000  1.450000 2.665000 1.780000 ;
      RECT 2.360000  1.780000 2.530000 2.130000 ;
      RECT 2.715000  1.950000 3.895000 2.120000 ;
      RECT 2.715000  2.120000 2.885000 2.980000 ;
      RECT 2.765000  0.085000 2.935000 0.690000 ;
      RECT 3.085000  2.290000 3.445000 3.245000 ;
      RECT 3.145000  0.085000 3.315000 0.840000 ;
      RECT 3.145000  0.840000 3.870000 1.010000 ;
      RECT 3.540000  1.010000 3.870000 1.290000 ;
      RECT 3.645000  1.940000 3.895000 1.950000 ;
      RECT 3.645000  2.120000 3.895000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_ls__a2bb2o_1
END LIBRARY
