* File: sky130_fd_sc_ls__or2_4.pex.spice
* Created: Wed Sep  2 11:24:18 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__OR2_4%A_83_260# 1 2 9 11 13 16 18 20 23 25 27 28 30
+ 33 35 43 47 49 51 54 55 57 58 62 71
c135 71 0 1.44954e-19 $X=1.855 $Y=1.532
r136 71 72 1.83969 $w=3.93e-07 $l=1.5e-08 $layer=POLY_cond $X=1.855 $Y=1.532
+ $X2=1.87 $Y2=1.532
r137 68 69 6.13232 $w=3.93e-07 $l=5e-08 $layer=POLY_cond $X=1.355 $Y=1.532
+ $X2=1.405 $Y2=1.532
r138 67 68 49.0585 $w=3.93e-07 $l=4e-07 $layer=POLY_cond $X=0.955 $Y=1.532
+ $X2=1.355 $Y2=1.532
r139 66 67 3.67939 $w=3.93e-07 $l=3e-08 $layer=POLY_cond $X=0.925 $Y=1.532
+ $X2=0.955 $Y2=1.532
r140 63 64 1.22646 $w=3.93e-07 $l=1e-08 $layer=POLY_cond $X=0.495 $Y=1.532
+ $X2=0.505 $Y2=1.532
r141 56 57 72.4171 $w=1.68e-07 $l=1.11e-06 $layer=LI1_cond $X=4.15 $Y=1.18
+ $X2=4.15 $Y2=2.29
r142 54 57 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.065 $Y=2.375
+ $X2=4.15 $Y2=2.29
r143 54 55 54.4759 $w=1.68e-07 $l=8.35e-07 $layer=LI1_cond $X=4.065 $Y=2.375
+ $X2=3.23 $Y2=2.375
r144 51 55 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.105 $Y=2.46
+ $X2=3.23 $Y2=2.375
r145 51 53 2.44 $w=2.5e-07 $l=5e-08 $layer=LI1_cond $X=3.105 $Y=2.46 $X2=3.105
+ $Y2=2.51
r146 50 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.75 $Y=1.095
+ $X2=2.585 $Y2=1.095
r147 49 56 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.065 $Y=1.095
+ $X2=4.15 $Y2=1.18
r148 49 50 85.7914 $w=1.68e-07 $l=1.315e-06 $layer=LI1_cond $X=4.065 $Y=1.095
+ $X2=2.75 $Y2=1.095
r149 45 62 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.585 $Y=1.01
+ $X2=2.585 $Y2=1.095
r150 45 47 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=2.585 $Y=1.01
+ $X2=2.585 $Y2=0.515
r151 44 58 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.04 $Y=1.095
+ $X2=1.955 $Y2=1.095
r152 43 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.42 $Y=1.095
+ $X2=2.585 $Y2=1.095
r153 43 44 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=2.42 $Y=1.095
+ $X2=2.04 $Y2=1.095
r154 42 71 9.19847 $w=3.93e-07 $l=7.5e-08 $layer=POLY_cond $X=1.78 $Y=1.532
+ $X2=1.855 $Y2=1.532
r155 42 69 45.9924 $w=3.93e-07 $l=3.75e-07 $layer=POLY_cond $X=1.78 $Y=1.532
+ $X2=1.405 $Y2=1.532
r156 41 42 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.78
+ $Y=1.465 $X2=1.78 $Y2=1.465
r157 38 66 20.2366 $w=3.93e-07 $l=1.65e-07 $layer=POLY_cond $X=0.76 $Y=1.532
+ $X2=0.925 $Y2=1.532
r158 38 64 31.2748 $w=3.93e-07 $l=2.55e-07 $layer=POLY_cond $X=0.76 $Y=1.532
+ $X2=0.505 $Y2=1.532
r159 37 41 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=0.76 $Y=1.465
+ $X2=1.78 $Y2=1.465
r160 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.76
+ $Y=1.465 $X2=0.76 $Y2=1.465
r161 35 58 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.955 $Y=1.465
+ $X2=1.955 $Y2=1.095
r162 35 41 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=1.87 $Y=1.465
+ $X2=1.78 $Y2=1.465
r163 31 72 25.4309 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=1.87 $Y=1.3
+ $X2=1.87 $Y2=1.532
r164 31 33 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.87 $Y=1.3
+ $X2=1.87 $Y2=0.74
r165 28 71 25.4309 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=1.855 $Y=1.765
+ $X2=1.855 $Y2=1.532
r166 28 30 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.855 $Y=1.765
+ $X2=1.855 $Y2=2.4
r167 25 69 25.4309 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=1.405 $Y=1.765
+ $X2=1.405 $Y2=1.532
r168 25 27 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.405 $Y=1.765
+ $X2=1.405 $Y2=2.4
r169 21 68 25.4309 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=1.355 $Y=1.3
+ $X2=1.355 $Y2=1.532
r170 21 23 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.355 $Y=1.3
+ $X2=1.355 $Y2=0.74
r171 18 67 25.4309 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=0.955 $Y=1.765
+ $X2=0.955 $Y2=1.532
r172 18 20 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.955 $Y=1.765
+ $X2=0.955 $Y2=2.4
r173 14 66 25.4309 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=0.925 $Y=1.3
+ $X2=0.925 $Y2=1.532
r174 14 16 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.925 $Y=1.3
+ $X2=0.925 $Y2=0.74
r175 11 64 25.4309 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=1.532
r176 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.4
r177 7 63 25.4309 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=0.495 $Y=1.3
+ $X2=0.495 $Y2=1.532
r178 7 9 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.495 $Y=1.3
+ $X2=0.495 $Y2=0.74
r179 2 53 600 $w=1.7e-07 $l=6.40625e-07 $layer=licon1_PDIFF $count=1 $X=2.915
+ $Y=1.94 $X2=3.065 $Y2=2.51
r180 1 47 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.445
+ $Y=0.37 $X2=2.585 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__OR2_4%A 3 5 7 8 10 11 15 18
c75 15 0 1.16609e-19 $X=3.755 $Y=1.615
c76 8 0 9.52465e-20 $X=3.79 $Y=1.865
r77 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.375
+ $Y=1.515 $X2=2.375 $Y2=1.515
r78 18 22 3.84454 $w=4.76e-07 $l=1.5e-07 $layer=LI1_cond $X=2.482 $Y=1.665
+ $X2=2.482 $Y2=1.515
r79 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.755
+ $Y=1.615 $X2=3.755 $Y2=1.615
r80 13 15 12.658 $w=3.03e-07 $l=3.35e-07 $layer=LI1_cond $X=3.742 $Y=1.95
+ $X2=3.742 $Y2=1.615
r81 12 18 9.48319 $w=4.76e-07 $l=4.8776e-07 $layer=LI1_cond $X=2.755 $Y=2.035
+ $X2=2.482 $Y2=1.665
r82 11 13 7.55824 $w=1.7e-07 $l=1.898e-07 $layer=LI1_cond $X=3.59 $Y=2.035
+ $X2=3.742 $Y2=1.95
r83 11 12 54.4759 $w=1.68e-07 $l=8.35e-07 $layer=LI1_cond $X=3.59 $Y=2.035
+ $X2=2.755 $Y2=2.035
r84 8 16 52.2586 $w=2.99e-07 $l=2.66927e-07 $layer=POLY_cond $X=3.79 $Y=1.865
+ $X2=3.755 $Y2=1.615
r85 8 10 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.79 $Y=1.865
+ $X2=3.79 $Y2=2.44
r86 5 21 71.0994 $w=2.76e-07 $l=3.57421e-07 $layer=POLY_cond $X=2.39 $Y=1.865
+ $X2=2.375 $Y2=1.515
r87 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.39 $Y=1.865
+ $X2=2.39 $Y2=2.44
r88 1 21 38.7914 $w=2.76e-07 $l=1.67481e-07 $layer=POLY_cond $X=2.37 $Y=1.35
+ $X2=2.375 $Y2=1.515
r89 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.37 $Y=1.35 $X2=2.37
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__OR2_4%B 1 3 6 8 10 11 16
r46 16 18 28.8623 $w=3.34e-07 $l=2e-07 $layer=POLY_cond $X=3.09 $Y=1.657
+ $X2=3.29 $Y2=1.657
r47 14 16 33.9132 $w=3.34e-07 $l=2.35e-07 $layer=POLY_cond $X=2.855 $Y=1.657
+ $X2=3.09 $Y2=1.657
r48 13 14 2.16467 $w=3.34e-07 $l=1.5e-08 $layer=POLY_cond $X=2.84 $Y=1.657
+ $X2=2.855 $Y2=1.657
r49 11 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.09
+ $Y=1.615 $X2=3.09 $Y2=1.615
r50 8 18 21.5099 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.29 $Y=1.865
+ $X2=3.29 $Y2=1.657
r51 8 10 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.29 $Y=1.865
+ $X2=3.29 $Y2=2.44
r52 4 14 21.5099 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.855 $Y=1.45
+ $X2=2.855 $Y2=1.657
r53 4 6 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=2.855 $Y=1.45
+ $X2=2.855 $Y2=0.74
r54 1 13 21.5099 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.84 $Y=1.865
+ $X2=2.84 $Y2=1.657
r55 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.84 $Y=1.865
+ $X2=2.84 $Y2=2.44
.ends

.subckt PM_SKY130_FD_SC_LS__OR2_4%VPWR 1 2 3 4 13 15 19 23 25 27 30 31 32 38 42
+ 54 58
r62 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r63 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r64 49 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r65 48 49 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r66 46 49 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r67 45 48 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.64 $Y=3.33 $X2=3.6
+ $Y2=3.33
r68 45 46 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r69 43 54 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.245 $Y=3.33
+ $X2=2.12 $Y2=3.33
r70 43 45 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=2.245 $Y=3.33
+ $X2=2.64 $Y2=3.33
r71 42 57 4.22425 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=3.93 $Y=3.33
+ $X2=4.125 $Y2=3.33
r72 42 48 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=3.93 $Y=3.33 $X2=3.6
+ $Y2=3.33
r73 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r74 38 54 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.995 $Y=3.33
+ $X2=2.12 $Y2=3.33
r75 38 40 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.995 $Y=3.33
+ $X2=1.68 $Y2=3.33
r76 37 41 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r77 37 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r78 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r79 34 51 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.182 $Y2=3.33
r80 34 36 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.72 $Y2=3.33
r81 32 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r82 32 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r83 32 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r84 30 36 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.095 $Y=3.33
+ $X2=0.72 $Y2=3.33
r85 30 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.095 $Y=3.33
+ $X2=1.18 $Y2=3.33
r86 29 40 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=1.265 $Y=3.33
+ $X2=1.68 $Y2=3.33
r87 29 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.265 $Y=3.33
+ $X2=1.18 $Y2=3.33
r88 25 57 3.09779 $w=2.75e-07 $l=1.1025e-07 $layer=LI1_cond $X=4.067 $Y=3.245
+ $X2=4.125 $Y2=3.33
r89 25 27 18.8582 $w=2.73e-07 $l=4.5e-07 $layer=LI1_cond $X=4.067 $Y=3.245
+ $X2=4.067 $Y2=2.795
r90 21 54 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.12 $Y=3.245
+ $X2=2.12 $Y2=3.33
r91 21 23 44.2538 $w=2.48e-07 $l=9.6e-07 $layer=LI1_cond $X=2.12 $Y=3.245
+ $X2=2.12 $Y2=2.285
r92 17 31 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.18 $Y=3.245
+ $X2=1.18 $Y2=3.33
r93 17 19 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=1.18 $Y=3.245
+ $X2=1.18 $Y2=2.305
r94 13 51 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.182 $Y2=3.33
r95 13 15 43.3319 $w=2.48e-07 $l=9.4e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.24 $Y2=2.305
r96 4 27 600 $w=1.7e-07 $l=9.31571e-07 $layer=licon1_PDIFF $count=1 $X=3.865
+ $Y=1.94 $X2=4.025 $Y2=2.795
r97 3 23 300 $w=1.7e-07 $l=5.14563e-07 $layer=licon1_PDIFF $count=2 $X=1.93
+ $Y=1.84 $X2=2.08 $Y2=2.285
r98 2 19 300 $w=1.7e-07 $l=5.34766e-07 $layer=licon1_PDIFF $count=2 $X=1.03
+ $Y=1.84 $X2=1.18 $Y2=2.305
r99 1 15 300 $w=1.7e-07 $l=5.32588e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.305
.ends

.subckt PM_SKY130_FD_SC_LS__OR2_4%X 1 2 3 4 13 14 15 16 19 23 27 29 33 37 43 44
+ 45 46
c80 13 0 2.19366e-19 $X=0.545 $Y=1.045
r81 45 46 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=1.295
+ $X2=0.24 $Y2=1.665
r82 42 46 6.76434 $w=2.28e-07 $l=1.35e-07 $layer=LI1_cond $X=0.24 $Y=1.8
+ $X2=0.24 $Y2=1.665
r83 41 45 8.26753 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.24 $Y=1.13
+ $X2=0.24 $Y2=1.295
r84 37 39 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=1.63 $Y=1.985
+ $X2=1.63 $Y2=2.815
r85 35 37 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=1.63 $Y=1.97
+ $X2=1.63 $Y2=1.985
r86 31 33 17.3843 $w=2.93e-07 $l=4.45e-07 $layer=LI1_cond $X=1.552 $Y=0.96
+ $X2=1.552 $Y2=0.515
r87 30 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=1.885
+ $X2=0.73 $Y2=1.885
r88 29 35 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.465 $Y=1.885
+ $X2=1.63 $Y2=1.97
r89 29 30 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.465 $Y=1.885
+ $X2=0.895 $Y2=1.885
r90 28 43 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.795 $Y=1.045
+ $X2=0.67 $Y2=1.045
r91 27 31 7.47753 $w=1.7e-07 $l=1.84673e-07 $layer=LI1_cond $X=1.405 $Y=1.045
+ $X2=1.552 $Y2=0.96
r92 27 28 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=1.405 $Y=1.045
+ $X2=0.795 $Y2=1.045
r93 23 25 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=0.73 $Y=1.985
+ $X2=0.73 $Y2=2.815
r94 21 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=1.97 $X2=0.73
+ $Y2=1.885
r95 21 23 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=0.73 $Y=1.97
+ $X2=0.73 $Y2=1.985
r96 17 43 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.67 $Y=0.96
+ $X2=0.67 $Y2=1.045
r97 17 19 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=0.67 $Y=0.96
+ $X2=0.67 $Y2=0.515
r98 16 42 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.355 $Y=1.885
+ $X2=0.24 $Y2=1.8
r99 15 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.565 $Y=1.885
+ $X2=0.73 $Y2=1.885
r100 15 16 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=0.565 $Y=1.885
+ $X2=0.355 $Y2=1.885
r101 14 41 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.355 $Y=1.045
+ $X2=0.24 $Y2=1.13
r102 13 43 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.545 $Y=1.045
+ $X2=0.67 $Y2=1.045
r103 13 14 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=0.545 $Y=1.045
+ $X2=0.355 $Y2=1.045
r104 4 39 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.48
+ $Y=1.84 $X2=1.63 $Y2=2.815
r105 4 37 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.48
+ $Y=1.84 $X2=1.63 $Y2=1.985
r106 3 25 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.84 $X2=0.73 $Y2=2.815
r107 3 23 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.84 $X2=0.73 $Y2=1.985
r108 2 33 91 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=2 $X=1.43
+ $Y=0.37 $X2=1.59 $Y2=0.515
r109 1 19 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__OR2_4%A_493_388# 1 2 9 11 12 14
c32 11 0 9.52465e-20 $X=3.4 $Y=2.99
c33 2 0 1.16609e-19 $X=3.365 $Y=1.94
r34 14 16 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=3.565 $Y=2.795
+ $X2=3.565 $Y2=2.99
r35 11 16 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.4 $Y=2.99
+ $X2=3.565 $Y2=2.99
r36 11 12 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=3.4 $Y=2.99 $X2=2.78
+ $Y2=2.99
r37 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.615 $Y=2.905
+ $X2=2.78 $Y2=2.99
r38 7 9 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=2.615 $Y=2.905
+ $X2=2.615 $Y2=2.455
r39 2 14 600 $w=1.7e-07 $l=9.4975e-07 $layer=licon1_PDIFF $count=1 $X=3.365
+ $Y=1.94 $X2=3.565 $Y2=2.795
r40 1 9 300 $w=1.7e-07 $l=5.85214e-07 $layer=licon1_PDIFF $count=2 $X=2.465
+ $Y=1.94 $X2=2.615 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_LS__OR2_4%VGND 1 2 3 4 13 15 19 23 26 27 28 34 38 47 55
+ 58
c55 1 0 7.44113e-20 $X=0.135 $Y=0.37
r56 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r57 55 57 0.778422 $w=8.62e-07 $l=5.5e-08 $layer=LI1_cond $X=4.025 $Y=0.377
+ $X2=4.08 $Y2=0.377
r58 53 58 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r59 52 55 12.8086 $w=8.62e-07 $l=9.05e-07 $layer=LI1_cond $X=3.12 $Y=0.377
+ $X2=4.025 $Y2=0.377
r60 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r61 50 52 0.707657 $w=8.62e-07 $l=5e-08 $layer=LI1_cond $X=3.07 $Y=0.377
+ $X2=3.12 $Y2=0.377
r62 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r63 42 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r64 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r65 39 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.25 $Y=0 $X2=2.085
+ $Y2=0
r66 39 41 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=2.25 $Y=0 $X2=2.64
+ $Y2=0
r67 38 50 11.8328 $w=8.62e-07 $l=4.45734e-07 $layer=LI1_cond $X=2.92 $Y=0
+ $X2=3.07 $Y2=0.377
r68 38 41 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=2.92 $Y=0 $X2=2.64
+ $Y2=0
r69 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r70 34 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.92 $Y=0 $X2=2.085
+ $Y2=0
r71 34 36 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r72 33 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r73 33 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r74 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r75 30 44 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=0 $X2=0.182
+ $Y2=0
r76 30 32 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=0 $X2=0.72
+ $Y2=0
r77 28 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r78 28 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r79 28 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r80 26 32 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.975 $Y=0 $X2=0.72
+ $Y2=0
r81 26 27 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.975 $Y=0 $X2=1.1
+ $Y2=0
r82 25 36 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=1.225 $Y=0 $X2=1.68
+ $Y2=0
r83 25 27 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.225 $Y=0 $X2=1.1
+ $Y2=0
r84 21 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.085 $Y=0.085
+ $X2=2.085 $Y2=0
r85 21 23 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=2.085 $Y=0.085
+ $X2=2.085 $Y2=0.675
r86 17 27 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=0.085
+ $X2=1.1 $Y2=0
r87 17 19 22.3574 $w=2.48e-07 $l=4.85e-07 $layer=LI1_cond $X=1.1 $Y=0.085
+ $X2=1.1 $Y2=0.57
r88 13 44 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.182 $Y2=0
r89 13 15 22.3574 $w=2.48e-07 $l=4.85e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.24 $Y2=0.57
r90 4 55 121.333 $w=1.7e-07 $l=1.23814e-06 $layer=licon1_NDIFF $count=1 $X=2.93
+ $Y=0.37 $X2=4.025 $Y2=0.675
r91 4 50 121.333 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=2.93
+ $Y=0.37 $X2=3.07 $Y2=0.675
r92 3 23 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=1.945
+ $Y=0.37 $X2=2.085 $Y2=0.675
r93 2 19 182 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=1 $X=1 $Y=0.37
+ $X2=1.14 $Y2=0.57
r94 1 15 182 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.57
.ends

