* File: sky130_fd_sc_ls__sdfbbp_1.pxi.spice
* Created: Wed Sep  2 11:26:46 2020
* 
x_PM_SKY130_FD_SC_LS__SDFBBP_1%SCD N_SCD_c_329_n N_SCD_c_334_n N_SCD_M1026_g
+ N_SCD_M1006_g SCD SCD N_SCD_c_330_n N_SCD_c_331_n N_SCD_c_332_n
+ PM_SKY130_FD_SC_LS__SDFBBP_1%SCD
x_PM_SKY130_FD_SC_LS__SDFBBP_1%D N_D_M1009_g N_D_c_359_n N_D_c_360_n N_D_M1010_g
+ D N_D_c_358_n PM_SKY130_FD_SC_LS__SDFBBP_1%D
x_PM_SKY130_FD_SC_LS__SDFBBP_1%A_341_93# N_A_341_93#_M1041_d N_A_341_93#_M1027_d
+ N_A_341_93#_M1012_g N_A_341_93#_c_409_n N_A_341_93#_M1019_g
+ N_A_341_93#_c_403_n N_A_341_93#_c_404_n N_A_341_93#_c_405_n
+ N_A_341_93#_c_406_n N_A_341_93#_c_411_n N_A_341_93#_c_412_n
+ N_A_341_93#_c_413_n N_A_341_93#_c_414_n N_A_341_93#_c_407_n
+ N_A_341_93#_c_408_n PM_SKY130_FD_SC_LS__SDFBBP_1%A_341_93#
x_PM_SKY130_FD_SC_LS__SDFBBP_1%SCE N_SCE_M1029_g N_SCE_c_493_n N_SCE_M1018_g
+ N_SCE_c_485_n N_SCE_c_486_n N_SCE_M1041_g N_SCE_c_488_n N_SCE_c_489_n
+ N_SCE_c_490_n N_SCE_c_495_n N_SCE_M1027_g SCE PM_SKY130_FD_SC_LS__SDFBBP_1%SCE
x_PM_SKY130_FD_SC_LS__SDFBBP_1%CLK N_CLK_c_568_n N_CLK_M1042_g N_CLK_c_571_n
+ N_CLK_M1040_g CLK N_CLK_c_570_n PM_SKY130_FD_SC_LS__SDFBBP_1%CLK
x_PM_SKY130_FD_SC_LS__SDFBBP_1%A_1250_231# N_A_1250_231#_M1015_d
+ N_A_1250_231#_M1024_d N_A_1250_231#_M1046_g N_A_1250_231#_c_612_n
+ N_A_1250_231#_c_622_n N_A_1250_231#_M1045_g N_A_1250_231#_c_613_n
+ N_A_1250_231#_M1034_g N_A_1250_231#_c_614_n N_A_1250_231#_c_615_n
+ N_A_1250_231#_M1013_g N_A_1250_231#_c_616_n N_A_1250_231#_c_617_n
+ N_A_1250_231#_c_652_p N_A_1250_231#_c_624_n N_A_1250_231#_c_625_n
+ N_A_1250_231#_c_626_n N_A_1250_231#_c_618_n N_A_1250_231#_c_627_n
+ N_A_1250_231#_c_687_p N_A_1250_231#_c_630_p N_A_1250_231#_c_673_p
+ N_A_1250_231#_c_619_n N_A_1250_231#_c_620_n
+ PM_SKY130_FD_SC_LS__SDFBBP_1%A_1250_231#
x_PM_SKY130_FD_SC_LS__SDFBBP_1%SET_B N_SET_B_M1022_g N_SET_B_c_772_n
+ N_SET_B_M1024_g N_SET_B_M1002_g N_SET_B_c_774_n N_SET_B_M1037_g
+ N_SET_B_c_778_n N_SET_B_c_779_n N_SET_B_c_780_n N_SET_B_c_781_n
+ N_SET_B_c_804_n N_SET_B_c_806_n N_SET_B_c_782_n N_SET_B_c_783_n
+ N_SET_B_c_784_n N_SET_B_c_785_n N_SET_B_c_786_n N_SET_B_c_787_n
+ N_SET_B_c_810_p N_SET_B_c_788_n N_SET_B_c_789_n SET_B
+ PM_SKY130_FD_SC_LS__SDFBBP_1%SET_B
x_PM_SKY130_FD_SC_LS__SDFBBP_1%A_1092_96# N_A_1092_96#_M1035_d
+ N_A_1092_96#_M1014_d N_A_1092_96#_M1015_g N_A_1092_96#_c_940_n
+ N_A_1092_96#_c_951_n N_A_1092_96#_M1039_g N_A_1092_96#_c_952_n
+ N_A_1092_96#_c_941_n N_A_1092_96#_c_953_n N_A_1092_96#_c_942_n
+ N_A_1092_96#_c_943_n N_A_1092_96#_c_944_n N_A_1092_96#_c_945_n
+ N_A_1092_96#_c_946_n N_A_1092_96#_c_947_n N_A_1092_96#_c_948_n
+ N_A_1092_96#_c_955_n N_A_1092_96#_c_949_n
+ PM_SKY130_FD_SC_LS__SDFBBP_1%A_1092_96#
x_PM_SKY130_FD_SC_LS__SDFBBP_1%A_1625_93# N_A_1625_93#_M1007_s
+ N_A_1625_93#_M1028_s N_A_1625_93#_M1016_g N_A_1625_93#_c_1059_n
+ N_A_1625_93#_c_1074_n N_A_1625_93#_M1033_g N_A_1625_93#_c_1060_n
+ N_A_1625_93#_c_1076_n N_A_1625_93#_M1017_g N_A_1625_93#_c_1061_n
+ N_A_1625_93#_M1043_g N_A_1625_93#_c_1062_n N_A_1625_93#_c_1063_n
+ N_A_1625_93#_c_1064_n N_A_1625_93#_c_1065_n N_A_1625_93#_c_1066_n
+ N_A_1625_93#_c_1067_n N_A_1625_93#_c_1068_n N_A_1625_93#_c_1069_n
+ N_A_1625_93#_c_1070_n N_A_1625_93#_c_1071_n N_A_1625_93#_c_1072_n
+ PM_SKY130_FD_SC_LS__SDFBBP_1%A_1625_93#
x_PM_SKY130_FD_SC_LS__SDFBBP_1%A_622_98# N_A_622_98#_M1042_s N_A_622_98#_M1040_s
+ N_A_622_98#_c_1196_n N_A_622_98#_M1000_g N_A_622_98#_c_1197_n
+ N_A_622_98#_M1004_g N_A_622_98#_c_1198_n N_A_622_98#_c_1199_n
+ N_A_622_98#_c_1200_n N_A_622_98#_c_1201_n N_A_622_98#_c_1202_n
+ N_A_622_98#_c_1220_n N_A_622_98#_c_1221_n N_A_622_98#_c_1203_n
+ N_A_622_98#_M1035_g N_A_622_98#_c_1222_n N_A_622_98#_c_1223_n
+ N_A_622_98#_c_1224_n N_A_622_98#_M1005_g N_A_622_98#_c_1225_n
+ N_A_622_98#_c_1204_n N_A_622_98#_M1008_g N_A_622_98#_M1023_g
+ N_A_622_98#_c_1205_n N_A_622_98#_c_1228_n N_A_622_98#_c_1206_n
+ N_A_622_98#_c_1207_n N_A_622_98#_c_1230_n N_A_622_98#_c_1231_n
+ N_A_622_98#_c_1232_n N_A_622_98#_c_1261_n N_A_622_98#_c_1233_n
+ N_A_622_98#_c_1208_n N_A_622_98#_c_1209_n N_A_622_98#_c_1210_n
+ N_A_622_98#_c_1211_n N_A_622_98#_c_1212_n N_A_622_98#_c_1213_n
+ N_A_622_98#_c_1235_n N_A_622_98#_c_1214_n N_A_622_98#_c_1215_n
+ N_A_622_98#_c_1216_n N_A_622_98#_c_1217_n
+ PM_SKY130_FD_SC_LS__SDFBBP_1%A_622_98#
x_PM_SKY130_FD_SC_LS__SDFBBP_1%A_877_98# N_A_877_98#_M1000_d N_A_877_98#_M1004_d
+ N_A_877_98#_c_1440_n N_A_877_98#_M1014_g N_A_877_98#_c_1441_n
+ N_A_877_98#_M1030_g N_A_877_98#_c_1443_n N_A_877_98#_c_1444_n
+ N_A_877_98#_M1001_g N_A_877_98#_c_1453_n N_A_877_98#_M1020_g
+ N_A_877_98#_c_1446_n N_A_877_98#_c_1447_n N_A_877_98#_c_1448_n
+ N_A_877_98#_c_1455_n N_A_877_98#_c_1449_n N_A_877_98#_c_1450_n
+ N_A_877_98#_c_1457_n N_A_877_98#_c_1458_n N_A_877_98#_c_1451_n
+ PM_SKY130_FD_SC_LS__SDFBBP_1%A_877_98#
x_PM_SKY130_FD_SC_LS__SDFBBP_1%A_2037_442# N_A_2037_442#_M1031_d
+ N_A_2037_442#_M1037_d N_A_2037_442#_c_1601_n N_A_2037_442#_M1036_g
+ N_A_2037_442#_M1047_g N_A_2037_442#_c_1591_n N_A_2037_442#_M1032_g
+ N_A_2037_442#_c_1592_n N_A_2037_442#_M1021_g N_A_2037_442#_c_1593_n
+ N_A_2037_442#_c_1594_n N_A_2037_442#_c_1595_n N_A_2037_442#_c_1605_n
+ N_A_2037_442#_c_1606_n N_A_2037_442#_c_1596_n N_A_2037_442#_M1025_g
+ N_A_2037_442#_c_1607_n N_A_2037_442#_M1011_g N_A_2037_442#_c_1597_n
+ N_A_2037_442#_c_1608_n N_A_2037_442#_c_1598_n N_A_2037_442#_c_1610_n
+ N_A_2037_442#_c_1626_n N_A_2037_442#_c_1599_n N_A_2037_442#_c_1612_n
+ N_A_2037_442#_c_1613_n N_A_2037_442#_c_1614_n N_A_2037_442#_c_1655_n
+ N_A_2037_442#_c_1600_n PM_SKY130_FD_SC_LS__SDFBBP_1%A_2037_442#
x_PM_SKY130_FD_SC_LS__SDFBBP_1%A_1878_420# N_A_1878_420#_M1001_d
+ N_A_1878_420#_M1008_d N_A_1878_420#_c_1772_n N_A_1878_420#_M1031_g
+ N_A_1878_420#_c_1773_n N_A_1878_420#_c_1774_n N_A_1878_420#_c_1783_n
+ N_A_1878_420#_M1044_g N_A_1878_420#_c_1775_n N_A_1878_420#_c_1776_n
+ N_A_1878_420#_c_1777_n N_A_1878_420#_c_1784_n N_A_1878_420#_c_1785_n
+ N_A_1878_420#_c_1778_n N_A_1878_420#_c_1787_n N_A_1878_420#_c_1779_n
+ N_A_1878_420#_c_1780_n N_A_1878_420#_c_1781_n
+ PM_SKY130_FD_SC_LS__SDFBBP_1%A_1878_420#
x_PM_SKY130_FD_SC_LS__SDFBBP_1%RESET_B N_RESET_B_c_1889_n N_RESET_B_M1028_g
+ N_RESET_B_c_1890_n N_RESET_B_M1007_g RESET_B
+ PM_SKY130_FD_SC_LS__SDFBBP_1%RESET_B
x_PM_SKY130_FD_SC_LS__SDFBBP_1%A_2881_74# N_A_2881_74#_M1025_s
+ N_A_2881_74#_M1011_s N_A_2881_74#_c_1921_n N_A_2881_74#_M1003_g
+ N_A_2881_74#_c_1923_n N_A_2881_74#_M1038_g N_A_2881_74#_c_1924_n
+ N_A_2881_74#_c_1928_n N_A_2881_74#_c_1925_n N_A_2881_74#_c_1926_n
+ PM_SKY130_FD_SC_LS__SDFBBP_1%A_2881_74#
x_PM_SKY130_FD_SC_LS__SDFBBP_1%A_27_464# N_A_27_464#_M1026_s N_A_27_464#_M1019_d
+ N_A_27_464#_c_1971_n N_A_27_464#_c_1981_n N_A_27_464#_c_1972_n
+ N_A_27_464#_c_1973_n N_A_27_464#_c_1974_n N_A_27_464#_c_1975_n
+ PM_SKY130_FD_SC_LS__SDFBBP_1%A_27_464#
x_PM_SKY130_FD_SC_LS__SDFBBP_1%VPWR N_VPWR_M1026_d N_VPWR_M1027_s N_VPWR_M1040_d
+ N_VPWR_M1045_d N_VPWR_M1033_d N_VPWR_M1036_d N_VPWR_M1017_d N_VPWR_M1028_d
+ N_VPWR_M1011_d N_VPWR_c_2013_n N_VPWR_c_2014_n N_VPWR_c_2015_n N_VPWR_c_2016_n
+ N_VPWR_c_2017_n N_VPWR_c_2018_n N_VPWR_c_2019_n N_VPWR_c_2020_n
+ N_VPWR_c_2021_n N_VPWR_c_2022_n N_VPWR_c_2023_n N_VPWR_c_2024_n
+ N_VPWR_c_2025_n N_VPWR_c_2026_n VPWR N_VPWR_c_2027_n N_VPWR_c_2028_n
+ N_VPWR_c_2029_n N_VPWR_c_2030_n N_VPWR_c_2031_n N_VPWR_c_2032_n
+ N_VPWR_c_2012_n N_VPWR_c_2034_n N_VPWR_c_2035_n N_VPWR_c_2036_n
+ N_VPWR_c_2037_n N_VPWR_c_2038_n N_VPWR_c_2039_n N_VPWR_c_2040_n
+ PM_SKY130_FD_SC_LS__SDFBBP_1%VPWR
x_PM_SKY130_FD_SC_LS__SDFBBP_1%A_197_119# N_A_197_119#_M1029_d
+ N_A_197_119#_M1035_s N_A_197_119#_M1010_d N_A_197_119#_M1014_s
+ N_A_197_119#_c_2192_n N_A_197_119#_c_2193_n N_A_197_119#_c_2194_n
+ N_A_197_119#_c_2207_n N_A_197_119#_c_2208_n N_A_197_119#_c_2209_n
+ N_A_197_119#_c_2195_n N_A_197_119#_c_2196_n N_A_197_119#_c_2197_n
+ N_A_197_119#_c_2198_n N_A_197_119#_c_2199_n N_A_197_119#_c_2272_n
+ N_A_197_119#_c_2211_n N_A_197_119#_c_2200_n N_A_197_119#_c_2201_n
+ N_A_197_119#_c_2202_n N_A_197_119#_c_2212_n N_A_197_119#_c_2213_n
+ N_A_197_119#_c_2203_n N_A_197_119#_c_2204_n N_A_197_119#_c_2205_n
+ N_A_197_119#_c_2206_n PM_SKY130_FD_SC_LS__SDFBBP_1%A_197_119#
x_PM_SKY130_FD_SC_LS__SDFBBP_1%Q_N N_Q_N_M1032_d N_Q_N_M1021_d N_Q_N_c_2376_n
+ N_Q_N_c_2378_n N_Q_N_c_2377_n Q_N Q_N Q_N PM_SKY130_FD_SC_LS__SDFBBP_1%Q_N
x_PM_SKY130_FD_SC_LS__SDFBBP_1%Q N_Q_M1003_d N_Q_M1038_d Q Q Q Q Q Q Q
+ PM_SKY130_FD_SC_LS__SDFBBP_1%Q
x_PM_SKY130_FD_SC_LS__SDFBBP_1%VGND N_VGND_M1006_s N_VGND_M1012_d N_VGND_M1042_d
+ N_VGND_M1046_d N_VGND_M1013_s N_VGND_M1047_d N_VGND_M1007_d N_VGND_M1025_d
+ N_VGND_c_2429_n N_VGND_c_2430_n N_VGND_c_2431_n N_VGND_c_2432_n
+ N_VGND_c_2433_n N_VGND_c_2434_n N_VGND_c_2435_n N_VGND_c_2436_n
+ N_VGND_c_2437_n N_VGND_c_2438_n N_VGND_c_2439_n N_VGND_c_2440_n
+ N_VGND_c_2441_n N_VGND_c_2442_n N_VGND_c_2443_n N_VGND_c_2444_n
+ N_VGND_c_2445_n N_VGND_c_2446_n N_VGND_c_2447_n VGND N_VGND_c_2448_n
+ N_VGND_c_2449_n N_VGND_c_2450_n N_VGND_c_2451_n N_VGND_c_2452_n
+ N_VGND_c_2453_n PM_SKY130_FD_SC_LS__SDFBBP_1%VGND
x_PM_SKY130_FD_SC_LS__SDFBBP_1%A_1418_125# N_A_1418_125#_M1022_d
+ N_A_1418_125#_M1016_d N_A_1418_125#_c_2600_n N_A_1418_125#_c_2601_n
+ N_A_1418_125#_c_2602_n N_A_1418_125#_c_2603_n
+ PM_SKY130_FD_SC_LS__SDFBBP_1%A_1418_125#
x_PM_SKY130_FD_SC_LS__SDFBBP_1%A_2271_74# N_A_2271_74#_M1002_d
+ N_A_2271_74#_M1043_d N_A_2271_74#_c_2628_n N_A_2271_74#_c_2626_n
+ N_A_2271_74#_c_2627_n N_A_2271_74#_c_2633_n
+ PM_SKY130_FD_SC_LS__SDFBBP_1%A_2271_74#
cc_1 VNB N_SCD_c_329_n 0.0299743f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.948
cc_2 VNB N_SCD_c_330_n 0.0225775f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.29
cc_3 VNB N_SCD_c_331_n 0.0240257f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.29
cc_4 VNB N_SCD_c_332_n 0.021308f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.125
cc_5 VNB N_D_M1009_g 0.036595f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.245
cc_6 VNB N_D_c_358_n 0.0178857f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.125
cc_7 VNB N_A_341_93#_M1012_g 0.0181701f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_8 VNB N_A_341_93#_c_403_n 0.0211159f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.29
cc_9 VNB N_A_341_93#_c_404_n 0.0070293f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.29
cc_10 VNB N_A_341_93#_c_405_n 0.0178377f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.97
cc_11 VNB N_A_341_93#_c_406_n 0.00480727f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.295
cc_12 VNB N_A_341_93#_c_407_n 0.00834216f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_341_93#_c_408_n 0.00230615f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_SCE_M1029_g 0.0600402f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.64
cc_15 VNB N_SCE_c_485_n 0.119631f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.805
cc_16 VNB N_SCE_c_486_n 0.0125534f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_17 VNB N_SCE_M1041_g 0.0424886f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.29
cc_18 VNB N_SCE_c_488_n 0.0341067f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.29
cc_19 VNB N_SCE_c_489_n 0.0082902f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.29
cc_20 VNB N_SCE_c_490_n 0.0144311f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.97
cc_21 VNB SCE 0.00729349f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_CLK_c_568_n 0.0209923f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.312
cc_23 VNB CLK 0.00149658f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.805
cc_24 VNB N_CLK_c_570_n 0.0473525f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_1250_231#_c_612_n 0.011191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_1250_231#_c_613_n 0.0442235f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.29
cc_27 VNB N_A_1250_231#_c_614_n 0.025206f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.97
cc_28 VNB N_A_1250_231#_c_615_n 0.0145459f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.29
cc_29 VNB N_A_1250_231#_c_616_n 0.00148285f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_1250_231#_c_617_n 0.0350307f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.97
cc_31 VNB N_A_1250_231#_c_618_n 0.00379322f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_1250_231#_c_619_n 0.00429347f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_1250_231#_c_620_n 0.017055f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_SET_B_M1022_g 0.0236098f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.245
cc_35 VNB N_SET_B_c_772_n 0.0324133f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.64
cc_36 VNB N_SET_B_M1002_g 0.0296477f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_37 VNB N_SET_B_c_774_n 0.0161335f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB SET_B 0.00293766f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_1092_96#_c_940_n 0.00435109f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_1092_96#_c_941_n 0.00502195f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.29
cc_41 VNB N_A_1092_96#_c_942_n 0.00978809f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_1092_96#_c_943_n 0.00738082f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.97
cc_43 VNB N_A_1092_96#_c_944_n 0.00937933f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_1092_96#_c_945_n 5.02483e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_1092_96#_c_946_n 0.00185291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_1092_96#_c_947_n 0.0330562f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_1092_96#_c_948_n 0.00329536f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_1092_96#_c_949_n 0.0150638f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_1625_93#_c_1059_n 0.00427417f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_1625_93#_c_1060_n 0.00560626f $X=-0.19 $Y=-0.245 $X2=0.407
+ $Y2=1.125
cc_51 VNB N_A_1625_93#_c_1061_n 0.0196411f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.29
cc_52 VNB N_A_1625_93#_c_1062_n 0.0103489f $X=-0.19 $Y=-0.245 $X2=0.337
+ $Y2=1.665
cc_53 VNB N_A_1625_93#_c_1063_n 0.00307309f $X=-0.19 $Y=-0.245 $X2=0.337
+ $Y2=1.97
cc_54 VNB N_A_1625_93#_c_1064_n 0.0102643f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_1625_93#_c_1065_n 0.0281833f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_1625_93#_c_1066_n 0.00316019f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_1625_93#_c_1067_n 0.00529492f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_1625_93#_c_1068_n 0.00558243f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_1625_93#_c_1069_n 0.00711735f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_1625_93#_c_1070_n 0.0472107f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_1625_93#_c_1071_n 0.0297949f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_1625_93#_c_1072_n 0.0162149f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_622_98#_c_1196_n 0.0205215f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.805
cc_64 VNB N_A_622_98#_c_1197_n 0.0192311f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_65 VNB N_A_622_98#_c_1198_n 0.0131244f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.29
cc_66 VNB N_A_622_98#_c_1199_n 0.0519925f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.125
cc_67 VNB N_A_622_98#_c_1200_n 0.00632024f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.97
cc_68 VNB N_A_622_98#_c_1201_n 0.0279179f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.97
cc_69 VNB N_A_622_98#_c_1202_n 0.0110612f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.29
cc_70 VNB N_A_622_98#_c_1203_n 0.0150535f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_622_98#_c_1204_n 0.0110666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_622_98#_c_1205_n 0.00456748f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_622_98#_c_1206_n 0.00270253f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_622_98#_c_1207_n 0.0103991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_622_98#_c_1208_n 0.00140895f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_622_98#_c_1209_n 0.0072384f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_622_98#_c_1210_n 0.00159638f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_622_98#_c_1211_n 9.35272e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_622_98#_c_1212_n 0.0409235f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_622_98#_c_1213_n 0.00110081f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_622_98#_c_1214_n 0.00578366f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_622_98#_c_1215_n 0.00276655f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_622_98#_c_1216_n 0.00283386f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_622_98#_c_1217_n 0.0177786f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_877_98#_c_1440_n 0.0264225f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.805
cc_86 VNB N_A_877_98#_c_1441_n 0.0295705f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_87 VNB N_A_877_98#_M1030_g 0.0387224f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.29
cc_88 VNB N_A_877_98#_c_1443_n 0.277845f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.125
cc_89 VNB N_A_877_98#_c_1444_n 0.012806f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.97
cc_90 VNB N_A_877_98#_M1001_g 0.0231085f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_877_98#_c_1446_n 0.0254326f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_877_98#_c_1447_n 0.0201749f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_877_98#_c_1448_n 8.29766e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_877_98#_c_1449_n 0.00188683f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_877_98#_c_1450_n 0.00319436f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_877_98#_c_1451_n 0.00104269f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_2037_442#_M1047_g 0.0660669f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_A_2037_442#_c_1591_n 0.0218739f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.29
cc_99 VNB N_A_2037_442#_c_1592_n 0.0267693f $X=-0.19 $Y=-0.245 $X2=0.407
+ $Y2=1.97
cc_100 VNB N_A_2037_442#_c_1593_n 0.013428f $X=-0.19 $Y=-0.245 $X2=0.337
+ $Y2=1.29
cc_101 VNB N_A_2037_442#_c_1594_n 0.0103711f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_A_2037_442#_c_1595_n 0.0385556f $X=-0.19 $Y=-0.245 $X2=0.337
+ $Y2=1.665
cc_103 VNB N_A_2037_442#_c_1596_n 0.0209162f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_A_2037_442#_c_1597_n 0.0180758f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_A_2037_442#_c_1598_n 0.00361747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_A_2037_442#_c_1599_n 2.54044e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_A_2037_442#_c_1600_n 0.0038611f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_A_1878_420#_c_1772_n 0.0170847f $X=-0.19 $Y=-0.245 $X2=0.52
+ $Y2=0.805
cc_109 VNB N_A_1878_420#_c_1773_n 0.0365731f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.58
cc_110 VNB N_A_1878_420#_c_1774_n 0.00109646f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_A_1878_420#_c_1775_n 0.00339841f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.97
cc_112 VNB N_A_1878_420#_c_1776_n 0.0168291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_A_1878_420#_c_1777_n 0.0112033f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_A_1878_420#_c_1778_n 0.00596049f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_A_1878_420#_c_1779_n 0.00263867f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_A_1878_420#_c_1780_n 0.00373872f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_A_1878_420#_c_1781_n 0.0062116f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_RESET_B_c_1889_n 0.0331418f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.312
cc_119 VNB N_RESET_B_c_1890_n 0.0191296f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.64
cc_120 VNB RESET_B 0.00507151f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.805
cc_121 VNB N_A_2881_74#_c_1921_n 0.0319612f $X=-0.19 $Y=-0.245 $X2=0.52
+ $Y2=0.805
cc_122 VNB N_A_2881_74#_M1003_g 0.0336849f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB N_A_2881_74#_c_1923_n 0.018961f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.29
cc_124 VNB N_A_2881_74#_c_1924_n 0.00727279f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.97
cc_125 VNB N_A_2881_74#_c_1925_n 0.00322927f $X=-0.19 $Y=-0.245 $X2=0.337
+ $Y2=1.97
cc_126 VNB N_A_2881_74#_c_1926_n 0.0205386f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_VPWR_c_2012_n 0.661241f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_A_197_119#_c_2192_n 0.00522969f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.29
cc_129 VNB N_A_197_119#_c_2193_n 0.0113434f $X=-0.19 $Y=-0.245 $X2=0.407
+ $Y2=1.97
cc_130 VNB N_A_197_119#_c_2194_n 0.00690269f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.97
cc_131 VNB N_A_197_119#_c_2195_n 0.00301188f $X=-0.19 $Y=-0.245 $X2=0.337
+ $Y2=1.97
cc_132 VNB N_A_197_119#_c_2196_n 0.00354417f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_A_197_119#_c_2197_n 0.0288489f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_A_197_119#_c_2198_n 0.00159638f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_A_197_119#_c_2199_n 4.70669e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_A_197_119#_c_2200_n 0.00116096f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_A_197_119#_c_2201_n 0.00806298f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB N_A_197_119#_c_2202_n 0.00224477f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VNB N_A_197_119#_c_2203_n 0.00535167f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_A_197_119#_c_2204_n 0.00634509f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_141 VNB N_A_197_119#_c_2205_n 0.0032067f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_142 VNB N_A_197_119#_c_2206_n 0.0049218f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_143 VNB N_Q_N_c_2376_n 0.0124108f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_144 VNB N_Q_N_c_2377_n 0.0024989f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.125
cc_145 VNB Q 0.0551271f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.805
cc_146 VNB N_VGND_c_2429_n 0.0130142f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_147 VNB N_VGND_c_2430_n 0.0375162f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_148 VNB N_VGND_c_2431_n 0.0115598f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_149 VNB N_VGND_c_2432_n 0.0111314f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_150 VNB N_VGND_c_2433_n 0.00960112f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_151 VNB N_VGND_c_2434_n 0.00833696f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_152 VNB N_VGND_c_2435_n 0.0105017f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_153 VNB N_VGND_c_2436_n 0.0199168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_154 VNB N_VGND_c_2437_n 0.0101645f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_155 VNB N_VGND_c_2438_n 0.0405226f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_156 VNB N_VGND_c_2439_n 0.00332923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_157 VNB N_VGND_c_2440_n 0.0628821f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_158 VNB N_VGND_c_2441_n 0.00523215f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_159 VNB N_VGND_c_2442_n 0.0512358f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_160 VNB N_VGND_c_2443_n 0.00332923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_161 VNB N_VGND_c_2444_n 0.0405127f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_162 VNB N_VGND_c_2445_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_163 VNB N_VGND_c_2446_n 0.0546501f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_164 VNB N_VGND_c_2447_n 0.00567425f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_165 VNB N_VGND_c_2448_n 0.0409263f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_166 VNB N_VGND_c_2449_n 0.0354411f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_167 VNB N_VGND_c_2450_n 0.0190734f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_168 VNB N_VGND_c_2451_n 0.813184f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_169 VNB N_VGND_c_2452_n 0.00631593f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_170 VNB N_VGND_c_2453_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_171 VNB N_A_1418_125#_c_2600_n 0.00487644f $X=-0.19 $Y=-0.245 $X2=0.52
+ $Y2=0.805
cc_172 VNB N_A_1418_125#_c_2601_n 0.00158793f $X=-0.19 $Y=-0.245 $X2=0.407
+ $Y2=1.29
cc_173 VNB N_A_1418_125#_c_2602_n 0.00603259f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.29
cc_174 VNB N_A_1418_125#_c_2603_n 0.00709193f $X=-0.19 $Y=-0.245 $X2=0.407
+ $Y2=1.125
cc_175 VNB N_A_2271_74#_c_2626_n 0.0094573f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_176 VNB N_A_2271_74#_c_2627_n 0.00203831f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_177 VPB N_SCD_c_329_n 0.0245355f $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.948
cc_178 VPB N_SCD_c_334_n 0.0535941f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.245
cc_179 VPB N_SCD_c_331_n 0.0209678f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.29
cc_180 VPB N_D_c_359_n 0.0178017f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.125
cc_181 VPB N_D_c_360_n 0.0198219f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=0.805
cc_182 VPB N_D_c_358_n 0.0222605f $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.125
cc_183 VPB N_A_341_93#_c_409_n 0.0450815f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_184 VPB N_A_341_93#_c_405_n 0.00965853f $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.97
cc_185 VPB N_A_341_93#_c_411_n 0.00930676f $X=-0.19 $Y=1.66 $X2=0.337 $Y2=1.97
cc_186 VPB N_A_341_93#_c_412_n 0.00836781f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_187 VPB N_A_341_93#_c_413_n 0.0181357f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_188 VPB N_A_341_93#_c_414_n 0.0453272f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_189 VPB N_A_341_93#_c_407_n 0.00297857f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_190 VPB N_SCE_M1029_g 0.00456256f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.64
cc_191 VPB N_SCE_c_493_n 0.0546516f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.64
cc_192 VPB N_SCE_c_490_n 0.0314782f $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.97
cc_193 VPB N_SCE_c_495_n 0.0272508f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.97
cc_194 VPB SCE 0.00698056f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_195 VPB N_CLK_c_571_n 0.0200933f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.64
cc_196 VPB CLK 0.00305837f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=0.805
cc_197 VPB N_CLK_c_570_n 0.0198164f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_198 VPB N_A_1250_231#_c_612_n 0.018996f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_199 VPB N_A_1250_231#_c_622_n 0.0248493f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_200 VPB N_A_1250_231#_c_613_n 0.0280871f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.29
cc_201 VPB N_A_1250_231#_c_624_n 0.00152427f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_202 VPB N_A_1250_231#_c_625_n 0.0118339f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_203 VPB N_A_1250_231#_c_626_n 0.00428337f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_204 VPB N_A_1250_231#_c_627_n 0.00110086f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_205 VPB N_SET_B_c_772_n 0.0393336f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.64
cc_206 VPB N_SET_B_c_774_n 0.0358814f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_207 VPB N_SET_B_c_778_n 0.00407861f $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.125
cc_208 VPB N_SET_B_c_779_n 0.0177039f $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.97
cc_209 VPB N_SET_B_c_780_n 0.00177503f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.97
cc_210 VPB N_SET_B_c_781_n 0.00388944f $X=-0.19 $Y=1.66 $X2=0.337 $Y2=1.29
cc_211 VPB N_SET_B_c_782_n 0.00179506f $X=-0.19 $Y=1.66 $X2=0.337 $Y2=1.665
cc_212 VPB N_SET_B_c_783_n 0.00724703f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_213 VPB N_SET_B_c_784_n 0.00254398f $X=-0.19 $Y=1.66 $X2=0.337 $Y2=1.97
cc_214 VPB N_SET_B_c_785_n 0.00214602f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_215 VPB N_SET_B_c_786_n 0.0123352f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_216 VPB N_SET_B_c_787_n 0.00322848f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_217 VPB N_SET_B_c_788_n 0.00366606f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_218 VPB N_SET_B_c_789_n 0.00295066f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_219 VPB SET_B 0.00298333f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_220 VPB N_A_1092_96#_c_940_n 0.00406303f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_221 VPB N_A_1092_96#_c_951_n 0.0193276f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_222 VPB N_A_1092_96#_c_952_n 0.00227653f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.29
cc_223 VPB N_A_1092_96#_c_953_n 0.00362539f $X=-0.19 $Y=1.66 $X2=0.337 $Y2=1.295
cc_224 VPB N_A_1092_96#_c_942_n 0.0152188f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_225 VPB N_A_1092_96#_c_955_n 0.00172346f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_226 VPB N_A_1625_93#_c_1059_n 0.00398537f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_227 VPB N_A_1625_93#_c_1074_n 0.0182282f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_228 VPB N_A_1625_93#_c_1060_n 0.00723134f $X=-0.19 $Y=1.66 $X2=0.407
+ $Y2=1.125
cc_229 VPB N_A_1625_93#_c_1076_n 0.022882f $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.97
cc_230 VPB N_A_1625_93#_c_1069_n 0.0170231f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_231 VPB N_A_622_98#_c_1197_n 0.0280526f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_232 VPB N_A_622_98#_c_1200_n 0.0803312f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.97
cc_233 VPB N_A_622_98#_c_1220_n 0.070684f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_234 VPB N_A_622_98#_c_1221_n 0.0123767f $X=-0.19 $Y=1.66 $X2=0.337 $Y2=1.295
cc_235 VPB N_A_622_98#_c_1222_n 0.00656267f $X=-0.19 $Y=1.66 $X2=0.337 $Y2=1.97
cc_236 VPB N_A_622_98#_c_1223_n 0.0329654f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_237 VPB N_A_622_98#_c_1224_n 0.0148684f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_238 VPB N_A_622_98#_c_1225_n 0.2555f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_239 VPB N_A_622_98#_c_1204_n 0.0335846f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_240 VPB N_A_622_98#_M1008_g 0.00917622f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_241 VPB N_A_622_98#_c_1228_n 0.00898827f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_242 VPB N_A_622_98#_c_1207_n 0.00469044f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_243 VPB N_A_622_98#_c_1230_n 0.0150216f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_244 VPB N_A_622_98#_c_1231_n 0.00386124f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_245 VPB N_A_622_98#_c_1232_n 0.0124161f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_246 VPB N_A_622_98#_c_1233_n 0.00342379f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_247 VPB N_A_622_98#_c_1208_n 0.00167683f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_248 VPB N_A_622_98#_c_1235_n 0.00177302f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_249 VPB N_A_622_98#_c_1214_n 5.76242e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_250 VPB N_A_877_98#_c_1440_n 0.0444048f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=0.805
cc_251 VPB N_A_877_98#_c_1453_n 0.0301827f $X=-0.19 $Y=1.66 $X2=0.337 $Y2=1.295
cc_252 VPB N_A_877_98#_c_1447_n 0.0285716f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_253 VPB N_A_877_98#_c_1455_n 0.00317395f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_254 VPB N_A_877_98#_c_1450_n 0.00544687f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_255 VPB N_A_877_98#_c_1457_n 0.00217276f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_256 VPB N_A_877_98#_c_1458_n 0.00134775f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_257 VPB N_A_877_98#_c_1451_n 2.87022e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_258 VPB N_A_2037_442#_c_1601_n 0.0150669f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=0.805
cc_259 VPB N_A_2037_442#_M1047_g 0.0228768f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_260 VPB N_A_2037_442#_c_1592_n 0.0244998f $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.97
cc_261 VPB N_A_2037_442#_c_1594_n 0.0131366f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_262 VPB N_A_2037_442#_c_1605_n 0.0437592f $X=-0.19 $Y=1.66 $X2=0.337 $Y2=1.97
cc_263 VPB N_A_2037_442#_c_1606_n 0.00987561f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_264 VPB N_A_2037_442#_c_1607_n 0.0204901f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_265 VPB N_A_2037_442#_c_1608_n 0.00321393f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_266 VPB N_A_2037_442#_c_1598_n 0.00245711f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_267 VPB N_A_2037_442#_c_1610_n 0.0126556f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_268 VPB N_A_2037_442#_c_1599_n 0.00176643f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_269 VPB N_A_2037_442#_c_1612_n 0.00613952f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_270 VPB N_A_2037_442#_c_1613_n 0.066091f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_271 VPB N_A_2037_442#_c_1614_n 0.00220763f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_272 VPB N_A_1878_420#_c_1774_n 0.00773295f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_273 VPB N_A_1878_420#_c_1783_n 0.0224225f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_274 VPB N_A_1878_420#_c_1784_n 0.00262024f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_275 VPB N_A_1878_420#_c_1785_n 0.00246477f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_276 VPB N_A_1878_420#_c_1778_n 5.70636e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_277 VPB N_A_1878_420#_c_1787_n 0.00347891f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_278 VPB N_RESET_B_c_1889_n 0.028975f $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.312
cc_279 VPB N_A_2881_74#_c_1923_n 0.0299957f $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.29
cc_280 VPB N_A_2881_74#_c_1928_n 0.0151144f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_281 VPB N_A_2881_74#_c_1925_n 8.90107e-19 $X=-0.19 $Y=1.66 $X2=0.337 $Y2=1.97
cc_282 VPB N_A_2881_74#_c_1926_n 0.00503556f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_283 VPB N_A_27_464#_c_1971_n 0.0101407f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_284 VPB N_A_27_464#_c_1972_n 0.00696227f $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.29
cc_285 VPB N_A_27_464#_c_1973_n 0.00213961f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.29
cc_286 VPB N_A_27_464#_c_1974_n 0.00364112f $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.97
cc_287 VPB N_A_27_464#_c_1975_n 0.0315505f $X=-0.19 $Y=1.66 $X2=0.337 $Y2=1.29
cc_288 VPB N_VPWR_c_2013_n 0.00662307f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_289 VPB N_VPWR_c_2014_n 0.0129036f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_290 VPB N_VPWR_c_2015_n 0.00799266f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_291 VPB N_VPWR_c_2016_n 0.018036f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_292 VPB N_VPWR_c_2017_n 0.00413849f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_293 VPB N_VPWR_c_2018_n 0.0282121f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_294 VPB N_VPWR_c_2019_n 0.0326941f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_295 VPB N_VPWR_c_2020_n 0.00996174f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_296 VPB N_VPWR_c_2021_n 0.0691689f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_297 VPB N_VPWR_c_2022_n 0.00436868f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_298 VPB N_VPWR_c_2023_n 0.0342772f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_299 VPB N_VPWR_c_2024_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_300 VPB N_VPWR_c_2025_n 0.0226891f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_301 VPB N_VPWR_c_2026_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_302 VPB N_VPWR_c_2027_n 0.0191515f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_303 VPB N_VPWR_c_2028_n 0.0382186f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_304 VPB N_VPWR_c_2029_n 0.0358621f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_305 VPB N_VPWR_c_2030_n 0.0325825f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_306 VPB N_VPWR_c_2031_n 0.0353089f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_307 VPB N_VPWR_c_2032_n 0.0197098f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_308 VPB N_VPWR_c_2012_n 0.168359f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_309 VPB N_VPWR_c_2034_n 0.00615051f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_310 VPB N_VPWR_c_2035_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_311 VPB N_VPWR_c_2036_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_312 VPB N_VPWR_c_2037_n 0.00490136f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_313 VPB N_VPWR_c_2038_n 0.0410497f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_314 VPB N_VPWR_c_2039_n 0.027589f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_315 VPB N_VPWR_c_2040_n 0.00497514f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_316 VPB N_A_197_119#_c_2207_n 0.00108792f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_317 VPB N_A_197_119#_c_2208_n 0.0043045f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_318 VPB N_A_197_119#_c_2209_n 0.00134561f $X=-0.19 $Y=1.66 $X2=0.337
+ $Y2=1.665
cc_319 VPB N_A_197_119#_c_2195_n 0.00307007f $X=-0.19 $Y=1.66 $X2=0.337 $Y2=1.97
cc_320 VPB N_A_197_119#_c_2211_n 0.00744044f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_321 VPB N_A_197_119#_c_2212_n 0.00517366f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_322 VPB N_A_197_119#_c_2213_n 0.00380491f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_323 VPB N_A_197_119#_c_2203_n 0.00353661f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_324 VPB N_Q_N_c_2378_n 0.00231862f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.29
cc_325 VPB N_Q_N_c_2377_n 9.54076e-19 $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.125
cc_326 VPB Q_N 0.0153067f $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.97
cc_327 VPB Q 0.054161f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=0.805
cc_328 N_SCD_c_331_n N_SCE_M1029_g 0.00215162f $X=0.385 $Y=1.29 $X2=0 $Y2=0
cc_329 N_SCD_c_332_n N_SCE_M1029_g 0.0682973f $X=0.407 $Y=1.125 $X2=0 $Y2=0
cc_330 N_SCD_c_329_n N_SCE_c_493_n 0.0204388f $X=0.407 $Y=1.948 $X2=0 $Y2=0
cc_331 N_SCD_c_334_n N_SCE_c_493_n 0.0261117f $X=0.505 $Y=2.245 $X2=0 $Y2=0
cc_332 N_SCD_c_331_n N_SCE_c_493_n 0.00129746f $X=0.385 $Y=1.29 $X2=0 $Y2=0
cc_333 N_SCD_c_329_n SCE 0.0027259f $X=0.407 $Y=1.948 $X2=0 $Y2=0
cc_334 N_SCD_c_331_n SCE 0.0319671f $X=0.385 $Y=1.29 $X2=0 $Y2=0
cc_335 N_SCD_c_334_n N_A_27_464#_c_1971_n 0.0111273f $X=0.505 $Y=2.245 $X2=0
+ $Y2=0
cc_336 N_SCD_c_331_n N_A_27_464#_c_1971_n 0.00788818f $X=0.385 $Y=1.29 $X2=0
+ $Y2=0
cc_337 N_SCD_c_334_n N_A_27_464#_c_1975_n 0.00968942f $X=0.505 $Y=2.245 $X2=0
+ $Y2=0
cc_338 N_SCD_c_331_n N_A_27_464#_c_1975_n 0.0287832f $X=0.385 $Y=1.29 $X2=0
+ $Y2=0
cc_339 N_SCD_c_334_n N_VPWR_c_2013_n 0.0050377f $X=0.505 $Y=2.245 $X2=0 $Y2=0
cc_340 N_SCD_c_334_n N_VPWR_c_2027_n 0.00445602f $X=0.505 $Y=2.245 $X2=0 $Y2=0
cc_341 N_SCD_c_334_n N_VPWR_c_2012_n 0.00459495f $X=0.505 $Y=2.245 $X2=0 $Y2=0
cc_342 N_SCD_c_331_n N_A_197_119#_c_2192_n 0.00215723f $X=0.385 $Y=1.29 $X2=0
+ $Y2=0
cc_343 N_SCD_c_331_n N_A_197_119#_c_2194_n 0.00655282f $X=0.385 $Y=1.29 $X2=0
+ $Y2=0
cc_344 N_SCD_c_330_n N_VGND_c_2430_n 0.00158682f $X=0.385 $Y=1.29 $X2=0 $Y2=0
cc_345 N_SCD_c_331_n N_VGND_c_2430_n 0.0263818f $X=0.385 $Y=1.29 $X2=0 $Y2=0
cc_346 N_SCD_c_332_n N_VGND_c_2430_n 0.012236f $X=0.407 $Y=1.125 $X2=0 $Y2=0
cc_347 N_SCD_c_332_n N_VGND_c_2438_n 0.0035863f $X=0.407 $Y=1.125 $X2=0 $Y2=0
cc_348 N_SCD_c_332_n N_VGND_c_2451_n 0.00401353f $X=0.407 $Y=1.125 $X2=0 $Y2=0
cc_349 N_D_M1009_g N_A_341_93#_M1012_g 0.050569f $X=1.42 $Y=0.805 $X2=0 $Y2=0
cc_350 N_D_c_359_n N_A_341_93#_c_409_n 0.0100047f $X=1.435 $Y=2.155 $X2=0 $Y2=0
cc_351 N_D_c_360_n N_A_341_93#_c_409_n 0.0178411f $X=1.435 $Y=2.245 $X2=0 $Y2=0
cc_352 N_D_c_358_n N_A_341_93#_c_404_n 0.00439424f $X=1.61 $Y=1.69 $X2=0 $Y2=0
cc_353 N_D_M1009_g N_A_341_93#_c_405_n 0.00208748f $X=1.42 $Y=0.805 $X2=0 $Y2=0
cc_354 D N_A_341_93#_c_405_n 3.54127e-19 $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_355 N_D_c_358_n N_A_341_93#_c_405_n 0.0176055f $X=1.61 $Y=1.69 $X2=0 $Y2=0
cc_356 N_D_M1009_g N_SCE_M1029_g 0.0344736f $X=1.42 $Y=0.805 $X2=0 $Y2=0
cc_357 D N_SCE_M1029_g 2.70819e-19 $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_358 N_D_c_359_n N_SCE_c_493_n 0.00824688f $X=1.435 $Y=2.155 $X2=0 $Y2=0
cc_359 N_D_c_360_n N_SCE_c_493_n 0.033628f $X=1.435 $Y=2.245 $X2=0 $Y2=0
cc_360 N_D_c_358_n N_SCE_c_493_n 0.0198435f $X=1.61 $Y=1.69 $X2=0 $Y2=0
cc_361 N_D_M1009_g N_SCE_c_485_n 0.0103003f $X=1.42 $Y=0.805 $X2=0 $Y2=0
cc_362 D SCE 0.0248041f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_363 N_D_c_358_n SCE 0.00579035f $X=1.61 $Y=1.69 $X2=0 $Y2=0
cc_364 N_D_c_360_n N_A_27_464#_c_1971_n 0.00142944f $X=1.435 $Y=2.245 $X2=0
+ $Y2=0
cc_365 N_D_c_360_n N_A_27_464#_c_1981_n 0.00393698f $X=1.435 $Y=2.245 $X2=0
+ $Y2=0
cc_366 N_D_c_360_n N_A_27_464#_c_1972_n 0.0129513f $X=1.435 $Y=2.245 $X2=0 $Y2=0
cc_367 N_D_c_360_n N_A_27_464#_c_1974_n 5.94448e-19 $X=1.435 $Y=2.245 $X2=0
+ $Y2=0
cc_368 N_D_c_360_n N_VPWR_c_2013_n 2.78881e-19 $X=1.435 $Y=2.245 $X2=0 $Y2=0
cc_369 N_D_c_360_n N_VPWR_c_2028_n 0.00278271f $X=1.435 $Y=2.245 $X2=0 $Y2=0
cc_370 N_D_c_360_n N_VPWR_c_2012_n 0.00353713f $X=1.435 $Y=2.245 $X2=0 $Y2=0
cc_371 N_D_M1009_g N_A_197_119#_c_2192_n 0.0129351f $X=1.42 $Y=0.805 $X2=0 $Y2=0
cc_372 N_D_M1009_g N_A_197_119#_c_2193_n 0.0138039f $X=1.42 $Y=0.805 $X2=0 $Y2=0
cc_373 D N_A_197_119#_c_2193_n 0.0231488f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_374 N_D_c_358_n N_A_197_119#_c_2193_n 0.00524488f $X=1.61 $Y=1.69 $X2=0 $Y2=0
cc_375 N_D_M1009_g N_A_197_119#_c_2194_n 0.00377559f $X=1.42 $Y=0.805 $X2=0
+ $Y2=0
cc_376 N_D_c_360_n N_A_197_119#_c_2207_n 0.00822785f $X=1.435 $Y=2.245 $X2=0
+ $Y2=0
cc_377 D N_A_197_119#_c_2208_n 0.0014655f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_378 N_D_c_358_n N_A_197_119#_c_2208_n 7.19666e-19 $X=1.61 $Y=1.69 $X2=0 $Y2=0
cc_379 N_D_c_359_n N_A_197_119#_c_2209_n 0.0048136f $X=1.435 $Y=2.155 $X2=0
+ $Y2=0
cc_380 N_D_c_360_n N_A_197_119#_c_2209_n 0.00125422f $X=1.435 $Y=2.245 $X2=0
+ $Y2=0
cc_381 D N_A_197_119#_c_2209_n 0.0210226f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_382 N_D_c_358_n N_A_197_119#_c_2209_n 0.00512292f $X=1.61 $Y=1.69 $X2=0 $Y2=0
cc_383 N_D_M1009_g N_A_197_119#_c_2195_n 0.00327089f $X=1.42 $Y=0.805 $X2=0
+ $Y2=0
cc_384 N_D_c_359_n N_A_197_119#_c_2195_n 0.00159203f $X=1.435 $Y=2.155 $X2=0
+ $Y2=0
cc_385 D N_A_197_119#_c_2195_n 0.0246554f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_386 N_D_c_358_n N_A_197_119#_c_2195_n 0.00199864f $X=1.61 $Y=1.69 $X2=0 $Y2=0
cc_387 N_D_M1009_g N_VGND_c_2431_n 0.00175435f $X=1.42 $Y=0.805 $X2=0 $Y2=0
cc_388 N_D_M1009_g N_VGND_c_2451_n 9.39239e-19 $X=1.42 $Y=0.805 $X2=0 $Y2=0
cc_389 N_A_341_93#_M1012_g N_SCE_c_485_n 0.0103107f $X=1.78 $Y=0.805 $X2=0 $Y2=0
cc_390 N_A_341_93#_M1012_g N_SCE_M1041_g 0.00805388f $X=1.78 $Y=0.805 $X2=0
+ $Y2=0
cc_391 N_A_341_93#_c_403_n N_SCE_M1041_g 0.00805231f $X=2.015 $Y=1.24 $X2=0
+ $Y2=0
cc_392 N_A_341_93#_c_408_n N_SCE_M1041_g 0.00701634f $X=2.735 $Y=1.035 $X2=0
+ $Y2=0
cc_393 N_A_341_93#_c_413_n N_SCE_c_488_n 4.75164e-19 $X=2.43 $Y=1.995 $X2=0
+ $Y2=0
cc_394 N_A_341_93#_c_407_n N_SCE_c_488_n 0.0147593f $X=2.527 $Y=1.83 $X2=0 $Y2=0
cc_395 N_A_341_93#_c_408_n N_SCE_c_488_n 0.00307297f $X=2.735 $Y=1.035 $X2=0
+ $Y2=0
cc_396 N_A_341_93#_c_405_n N_SCE_c_489_n 0.00805231f $X=2.09 $Y=1.83 $X2=0 $Y2=0
cc_397 N_A_341_93#_c_413_n N_SCE_c_489_n 0.0012634f $X=2.43 $Y=1.995 $X2=0 $Y2=0
cc_398 N_A_341_93#_c_414_n N_SCE_c_489_n 0.00596612f $X=2.43 $Y=1.995 $X2=0
+ $Y2=0
cc_399 N_A_341_93#_c_405_n N_SCE_c_490_n 0.00409988f $X=2.09 $Y=1.83 $X2=0 $Y2=0
cc_400 N_A_341_93#_c_414_n N_SCE_c_490_n 0.0249515f $X=2.43 $Y=1.995 $X2=0 $Y2=0
cc_401 N_A_341_93#_c_407_n N_SCE_c_490_n 0.00610297f $X=2.527 $Y=1.83 $X2=0
+ $Y2=0
cc_402 N_A_341_93#_c_411_n N_SCE_c_495_n 0.0216638f $X=2.955 $Y=2.265 $X2=0
+ $Y2=0
cc_403 N_A_341_93#_c_412_n N_SCE_c_495_n 0.0126551f $X=3.12 $Y=2.465 $X2=0 $Y2=0
cc_404 N_A_341_93#_c_413_n N_SCE_c_495_n 0.00731794f $X=2.43 $Y=1.995 $X2=0
+ $Y2=0
cc_405 N_A_341_93#_c_411_n N_CLK_c_571_n 3.52096e-19 $X=2.955 $Y=2.265 $X2=0
+ $Y2=0
cc_406 N_A_341_93#_c_412_n N_CLK_c_571_n 0.00114899f $X=3.12 $Y=2.465 $X2=0
+ $Y2=0
cc_407 N_A_341_93#_c_406_n N_A_622_98#_c_1206_n 0.0141509f $X=2.695 $Y=0.815
+ $X2=0 $Y2=0
cc_408 N_A_341_93#_c_407_n N_A_622_98#_c_1207_n 0.0393014f $X=2.527 $Y=1.83
+ $X2=0 $Y2=0
cc_409 N_A_341_93#_c_411_n N_A_622_98#_c_1230_n 0.0020737f $X=2.955 $Y=2.265
+ $X2=0 $Y2=0
cc_410 N_A_341_93#_c_411_n N_A_622_98#_c_1231_n 0.0158349f $X=2.955 $Y=2.265
+ $X2=0 $Y2=0
cc_411 N_A_341_93#_c_413_n N_A_622_98#_c_1231_n 0.0101803f $X=2.43 $Y=1.995
+ $X2=0 $Y2=0
cc_412 N_A_341_93#_c_411_n N_A_622_98#_c_1232_n 0.0118844f $X=2.955 $Y=2.265
+ $X2=0 $Y2=0
cc_413 N_A_341_93#_c_412_n N_A_622_98#_c_1232_n 0.0424401f $X=3.12 $Y=2.465
+ $X2=0 $Y2=0
cc_414 N_A_341_93#_c_408_n N_A_622_98#_c_1213_n 0.0141509f $X=2.735 $Y=1.035
+ $X2=0 $Y2=0
cc_415 N_A_341_93#_c_409_n N_A_27_464#_c_1972_n 0.0137419f $X=1.885 $Y=2.245
+ $X2=0 $Y2=0
cc_416 N_A_341_93#_c_409_n N_A_27_464#_c_1974_n 0.0163176f $X=1.885 $Y=2.245
+ $X2=0 $Y2=0
cc_417 N_A_341_93#_c_413_n N_VPWR_M1027_s 0.0029325f $X=2.43 $Y=1.995 $X2=0
+ $Y2=0
cc_418 N_A_341_93#_c_409_n N_VPWR_c_2014_n 0.00155687f $X=1.885 $Y=2.245 $X2=0
+ $Y2=0
cc_419 N_A_341_93#_c_412_n N_VPWR_c_2014_n 0.030873f $X=3.12 $Y=2.465 $X2=0
+ $Y2=0
cc_420 N_A_341_93#_c_413_n N_VPWR_c_2014_n 0.0222424f $X=2.43 $Y=1.995 $X2=0
+ $Y2=0
cc_421 N_A_341_93#_c_414_n N_VPWR_c_2014_n 5.39441e-19 $X=2.43 $Y=1.995 $X2=0
+ $Y2=0
cc_422 N_A_341_93#_c_409_n N_VPWR_c_2028_n 0.00278257f $X=1.885 $Y=2.245 $X2=0
+ $Y2=0
cc_423 N_A_341_93#_c_412_n N_VPWR_c_2029_n 0.0145938f $X=3.12 $Y=2.465 $X2=0
+ $Y2=0
cc_424 N_A_341_93#_c_409_n N_VPWR_c_2012_n 0.00358707f $X=1.885 $Y=2.245 $X2=0
+ $Y2=0
cc_425 N_A_341_93#_c_412_n N_VPWR_c_2012_n 0.0120466f $X=3.12 $Y=2.465 $X2=0
+ $Y2=0
cc_426 N_A_341_93#_M1012_g N_A_197_119#_c_2192_n 0.00205619f $X=1.78 $Y=0.805
+ $X2=0 $Y2=0
cc_427 N_A_341_93#_c_403_n N_A_197_119#_c_2193_n 0.00251998f $X=2.015 $Y=1.24
+ $X2=0 $Y2=0
cc_428 N_A_341_93#_c_404_n N_A_197_119#_c_2193_n 0.0102501f $X=1.855 $Y=1.24
+ $X2=0 $Y2=0
cc_429 N_A_341_93#_c_409_n N_A_197_119#_c_2207_n 0.00631246f $X=1.885 $Y=2.245
+ $X2=0 $Y2=0
cc_430 N_A_341_93#_c_413_n N_A_197_119#_c_2207_n 0.00561945f $X=2.43 $Y=1.995
+ $X2=0 $Y2=0
cc_431 N_A_341_93#_c_409_n N_A_197_119#_c_2208_n 0.0195349f $X=1.885 $Y=2.245
+ $X2=0 $Y2=0
cc_432 N_A_341_93#_c_413_n N_A_197_119#_c_2208_n 0.0138837f $X=2.43 $Y=1.995
+ $X2=0 $Y2=0
cc_433 N_A_341_93#_c_409_n N_A_197_119#_c_2195_n 0.00581324f $X=1.885 $Y=2.245
+ $X2=0 $Y2=0
cc_434 N_A_341_93#_c_403_n N_A_197_119#_c_2195_n 8.20788e-19 $X=2.015 $Y=1.24
+ $X2=0 $Y2=0
cc_435 N_A_341_93#_c_405_n N_A_197_119#_c_2195_n 0.0140014f $X=2.09 $Y=1.83
+ $X2=0 $Y2=0
cc_436 N_A_341_93#_c_413_n N_A_197_119#_c_2195_n 0.0143835f $X=2.43 $Y=1.995
+ $X2=0 $Y2=0
cc_437 N_A_341_93#_c_407_n N_A_197_119#_c_2195_n 0.0146195f $X=2.527 $Y=1.83
+ $X2=0 $Y2=0
cc_438 N_A_341_93#_M1012_g N_A_197_119#_c_2196_n 0.00356535f $X=1.78 $Y=0.805
+ $X2=0 $Y2=0
cc_439 N_A_341_93#_c_403_n N_A_197_119#_c_2196_n 4.69448e-19 $X=2.015 $Y=1.24
+ $X2=0 $Y2=0
cc_440 N_A_341_93#_c_408_n N_A_197_119#_c_2196_n 0.0241746f $X=2.735 $Y=1.035
+ $X2=0 $Y2=0
cc_441 N_A_341_93#_c_406_n N_A_197_119#_c_2197_n 0.0189979f $X=2.695 $Y=0.815
+ $X2=0 $Y2=0
cc_442 N_A_341_93#_c_403_n N_A_197_119#_c_2204_n 0.00919997f $X=2.015 $Y=1.24
+ $X2=0 $Y2=0
cc_443 N_A_341_93#_c_405_n N_A_197_119#_c_2204_n 0.00391173f $X=2.09 $Y=1.83
+ $X2=0 $Y2=0
cc_444 N_A_341_93#_c_413_n N_A_197_119#_c_2204_n 0.00512817f $X=2.43 $Y=1.995
+ $X2=0 $Y2=0
cc_445 N_A_341_93#_c_414_n N_A_197_119#_c_2204_n 0.0038267f $X=2.43 $Y=1.995
+ $X2=0 $Y2=0
cc_446 N_A_341_93#_c_407_n N_A_197_119#_c_2204_n 0.0121121f $X=2.527 $Y=1.83
+ $X2=0 $Y2=0
cc_447 N_A_341_93#_M1012_g N_VGND_c_2431_n 0.0116571f $X=1.78 $Y=0.805 $X2=0
+ $Y2=0
cc_448 N_A_341_93#_c_403_n N_VGND_c_2431_n 0.00484302f $X=2.015 $Y=1.24 $X2=0
+ $Y2=0
cc_449 N_A_341_93#_M1012_g N_VGND_c_2451_n 7.88961e-19 $X=1.78 $Y=0.805 $X2=0
+ $Y2=0
cc_450 N_SCE_c_488_n N_CLK_c_568_n 0.00424269f $X=2.805 $Y=1.38 $X2=-0.19
+ $Y2=-0.245
cc_451 N_SCE_c_490_n N_CLK_c_570_n 0.00424269f $X=2.895 $Y=2.155 $X2=0 $Y2=0
cc_452 N_SCE_c_488_n N_A_622_98#_c_1207_n 0.00776119f $X=2.805 $Y=1.38 $X2=0
+ $Y2=0
cc_453 N_SCE_c_490_n N_A_622_98#_c_1231_n 0.00423256f $X=2.895 $Y=2.155 $X2=0
+ $Y2=0
cc_454 N_SCE_c_490_n N_A_622_98#_c_1232_n 0.00438614f $X=2.895 $Y=2.155 $X2=0
+ $Y2=0
cc_455 N_SCE_c_495_n N_A_622_98#_c_1232_n 0.00171231f $X=2.895 $Y=2.245 $X2=0
+ $Y2=0
cc_456 N_SCE_c_493_n N_A_27_464#_c_1971_n 0.0137462f $X=1.015 $Y=2.245 $X2=0
+ $Y2=0
cc_457 SCE N_A_27_464#_c_1971_n 0.0333898f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_458 N_SCE_c_493_n N_A_27_464#_c_1973_n 0.00120849f $X=1.015 $Y=2.245 $X2=0
+ $Y2=0
cc_459 N_SCE_c_493_n N_A_27_464#_c_1975_n 4.44963e-19 $X=1.015 $Y=2.245 $X2=0
+ $Y2=0
cc_460 N_SCE_c_493_n N_VPWR_c_2013_n 0.00561513f $X=1.015 $Y=2.245 $X2=0 $Y2=0
cc_461 N_SCE_c_495_n N_VPWR_c_2014_n 0.00729942f $X=2.895 $Y=2.245 $X2=0 $Y2=0
cc_462 N_SCE_c_493_n N_VPWR_c_2028_n 0.00444681f $X=1.015 $Y=2.245 $X2=0 $Y2=0
cc_463 N_SCE_c_495_n N_VPWR_c_2029_n 0.00445602f $X=2.895 $Y=2.245 $X2=0 $Y2=0
cc_464 N_SCE_c_493_n N_VPWR_c_2012_n 0.00448284f $X=1.015 $Y=2.245 $X2=0 $Y2=0
cc_465 N_SCE_c_495_n N_VPWR_c_2012_n 0.00867193f $X=2.895 $Y=2.245 $X2=0 $Y2=0
cc_466 N_SCE_M1029_g N_A_197_119#_c_2192_n 0.00633736f $X=0.91 $Y=0.805 $X2=0
+ $Y2=0
cc_467 N_SCE_c_485_n N_A_197_119#_c_2192_n 0.00555293f $X=2.405 $Y=0.18 $X2=0
+ $Y2=0
cc_468 N_SCE_M1029_g N_A_197_119#_c_2194_n 0.00253737f $X=0.91 $Y=0.805 $X2=0
+ $Y2=0
cc_469 N_SCE_c_493_n N_A_197_119#_c_2194_n 4.6141e-19 $X=1.015 $Y=2.245 $X2=0
+ $Y2=0
cc_470 SCE N_A_197_119#_c_2194_n 0.0203976f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_471 N_SCE_c_493_n N_A_197_119#_c_2207_n 7.49884e-19 $X=1.015 $Y=2.245 $X2=0
+ $Y2=0
cc_472 N_SCE_c_493_n N_A_197_119#_c_2209_n 5.28301e-19 $X=1.015 $Y=2.245 $X2=0
+ $Y2=0
cc_473 SCE N_A_197_119#_c_2209_n 0.00511267f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_474 N_SCE_c_489_n N_A_197_119#_c_2195_n 4.11552e-19 $X=2.555 $Y=1.38 $X2=0
+ $Y2=0
cc_475 SCE N_A_197_119#_c_2195_n 0.00539731f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_476 N_SCE_M1041_g N_A_197_119#_c_2196_n 0.0224621f $X=2.48 $Y=0.805 $X2=0
+ $Y2=0
cc_477 N_SCE_M1041_g N_A_197_119#_c_2197_n 0.0132477f $X=2.48 $Y=0.805 $X2=0
+ $Y2=0
cc_478 N_SCE_c_485_n N_A_197_119#_c_2198_n 0.0030135f $X=2.405 $Y=0.18 $X2=0
+ $Y2=0
cc_479 N_SCE_M1041_g N_A_197_119#_c_2198_n 0.00319103f $X=2.48 $Y=0.805 $X2=0
+ $Y2=0
cc_480 N_SCE_M1041_g N_A_197_119#_c_2204_n 0.00249837f $X=2.48 $Y=0.805 $X2=0
+ $Y2=0
cc_481 N_SCE_c_489_n N_A_197_119#_c_2204_n 0.00154215f $X=2.555 $Y=1.38 $X2=0
+ $Y2=0
cc_482 N_SCE_M1029_g N_VGND_c_2430_n 0.00166246f $X=0.91 $Y=0.805 $X2=0 $Y2=0
cc_483 N_SCE_c_486_n N_VGND_c_2430_n 0.00977077f $X=0.985 $Y=0.18 $X2=0 $Y2=0
cc_484 N_SCE_c_485_n N_VGND_c_2431_n 0.0210723f $X=2.405 $Y=0.18 $X2=0 $Y2=0
cc_485 N_SCE_M1041_g N_VGND_c_2431_n 0.00260915f $X=2.48 $Y=0.805 $X2=0 $Y2=0
cc_486 N_SCE_c_486_n N_VGND_c_2438_n 0.03227f $X=0.985 $Y=0.18 $X2=0 $Y2=0
cc_487 N_SCE_c_485_n N_VGND_c_2448_n 0.012994f $X=2.405 $Y=0.18 $X2=0 $Y2=0
cc_488 N_SCE_c_485_n N_VGND_c_2451_n 0.0501808f $X=2.405 $Y=0.18 $X2=0 $Y2=0
cc_489 N_SCE_c_486_n N_VGND_c_2451_n 0.0116041f $X=0.985 $Y=0.18 $X2=0 $Y2=0
cc_490 N_CLK_c_568_n N_A_622_98#_c_1196_n 0.0141211f $X=3.47 $Y=1.34 $X2=0 $Y2=0
cc_491 CLK N_A_622_98#_c_1196_n 0.00301156f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_492 N_CLK_c_571_n N_A_622_98#_c_1197_n 0.0205083f $X=3.905 $Y=1.765 $X2=0
+ $Y2=0
cc_493 CLK N_A_622_98#_c_1197_n 2.47524e-19 $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_494 N_CLK_c_570_n N_A_622_98#_c_1197_n 0.0201929f $X=3.595 $Y=1.505 $X2=0
+ $Y2=0
cc_495 N_CLK_c_568_n N_A_622_98#_c_1207_n 0.0117849f $X=3.47 $Y=1.34 $X2=0 $Y2=0
cc_496 N_CLK_c_571_n N_A_622_98#_c_1207_n 0.00165935f $X=3.905 $Y=1.765 $X2=0
+ $Y2=0
cc_497 CLK N_A_622_98#_c_1207_n 0.0367217f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_498 N_CLK_c_570_n N_A_622_98#_c_1207_n 0.0022226f $X=3.595 $Y=1.505 $X2=0
+ $Y2=0
cc_499 CLK N_A_622_98#_c_1230_n 0.00650302f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_500 N_CLK_c_570_n N_A_622_98#_c_1230_n 0.00207629f $X=3.595 $Y=1.505 $X2=0
+ $Y2=0
cc_501 N_CLK_c_571_n N_A_622_98#_c_1232_n 0.0122184f $X=3.905 $Y=1.765 $X2=0
+ $Y2=0
cc_502 N_CLK_c_571_n N_A_622_98#_c_1261_n 0.0153482f $X=3.905 $Y=1.765 $X2=0
+ $Y2=0
cc_503 N_CLK_c_571_n N_A_622_98#_c_1233_n 0.00169707f $X=3.905 $Y=1.765 $X2=0
+ $Y2=0
cc_504 N_CLK_c_570_n N_A_622_98#_c_1233_n 0.00220016f $X=3.595 $Y=1.505 $X2=0
+ $Y2=0
cc_505 N_CLK_c_571_n N_A_622_98#_c_1235_n 9.07447e-19 $X=3.905 $Y=1.765 $X2=0
+ $Y2=0
cc_506 CLK N_A_622_98#_c_1235_n 0.0208593f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_507 N_CLK_c_570_n N_A_622_98#_c_1235_n 0.00340098f $X=3.595 $Y=1.505 $X2=0
+ $Y2=0
cc_508 CLK N_A_622_98#_c_1214_n 0.0169888f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_509 N_CLK_c_570_n N_A_622_98#_c_1214_n 0.00345208f $X=3.595 $Y=1.505 $X2=0
+ $Y2=0
cc_510 N_CLK_c_571_n N_A_877_98#_c_1457_n 7.96058e-19 $X=3.905 $Y=1.765 $X2=0
+ $Y2=0
cc_511 N_CLK_c_571_n N_VPWR_c_2015_n 0.00556363f $X=3.905 $Y=1.765 $X2=0 $Y2=0
cc_512 N_CLK_c_571_n N_VPWR_c_2029_n 0.00445602f $X=3.905 $Y=1.765 $X2=0 $Y2=0
cc_513 N_CLK_c_571_n N_VPWR_c_2012_n 0.00862475f $X=3.905 $Y=1.765 $X2=0 $Y2=0
cc_514 N_CLK_c_568_n N_A_197_119#_c_2197_n 0.010802f $X=3.47 $Y=1.34 $X2=0 $Y2=0
cc_515 N_CLK_c_568_n N_A_197_119#_c_2199_n 0.0108329f $X=3.47 $Y=1.34 $X2=0
+ $Y2=0
cc_516 N_CLK_c_568_n N_A_197_119#_c_2272_n 0.00619015f $X=3.47 $Y=1.34 $X2=0
+ $Y2=0
cc_517 CLK N_A_197_119#_c_2272_n 0.00553438f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_518 N_CLK_c_570_n N_A_197_119#_c_2272_n 5.34366e-19 $X=3.595 $Y=1.505 $X2=0
+ $Y2=0
cc_519 CLK N_A_197_119#_c_2205_n 0.00365142f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_520 N_CLK_c_570_n N_A_197_119#_c_2205_n 0.00684242f $X=3.595 $Y=1.505 $X2=0
+ $Y2=0
cc_521 CLK N_VGND_M1042_d 0.00322771f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_522 N_CLK_c_568_n N_VGND_c_2432_n 4.29002e-19 $X=3.47 $Y=1.34 $X2=0 $Y2=0
cc_523 N_CLK_c_568_n N_VGND_c_2448_n 7.44058e-19 $X=3.47 $Y=1.34 $X2=0 $Y2=0
cc_524 N_A_1250_231#_c_616_n N_SET_B_M1022_g 0.00343382f $X=6.415 $Y=1.32 $X2=0
+ $Y2=0
cc_525 N_A_1250_231#_c_617_n N_SET_B_M1022_g 0.00913261f $X=6.415 $Y=1.32 $X2=0
+ $Y2=0
cc_526 N_A_1250_231#_c_630_p N_SET_B_M1022_g 0.0134669f $X=7.82 $Y=0.777 $X2=0
+ $Y2=0
cc_527 N_A_1250_231#_c_620_n N_SET_B_M1022_g 0.0138644f $X=6.415 $Y=1.155 $X2=0
+ $Y2=0
cc_528 N_A_1250_231#_c_612_n N_SET_B_c_772_n 0.00874645f $X=6.45 $Y=1.93 $X2=0
+ $Y2=0
cc_529 N_A_1250_231#_c_622_n N_SET_B_c_772_n 0.00589544f $X=6.45 $Y=2.02 $X2=0
+ $Y2=0
cc_530 N_A_1250_231#_c_624_n N_SET_B_c_772_n 0.00627137f $X=7.6 $Y=2.04 $X2=0
+ $Y2=0
cc_531 N_A_1250_231#_c_626_n N_SET_B_c_772_n 0.00154481f $X=7.765 $Y=1.91 $X2=0
+ $Y2=0
cc_532 N_A_1250_231#_c_612_n N_SET_B_c_778_n 0.00327819f $X=6.45 $Y=1.93 $X2=0
+ $Y2=0
cc_533 N_A_1250_231#_c_622_n N_SET_B_c_778_n 0.00142598f $X=6.45 $Y=2.02 $X2=0
+ $Y2=0
cc_534 N_A_1250_231#_c_624_n N_SET_B_c_778_n 0.0547143f $X=7.6 $Y=2.04 $X2=0
+ $Y2=0
cc_535 N_A_1250_231#_c_626_n N_SET_B_c_778_n 0.0135401f $X=7.765 $Y=1.91 $X2=0
+ $Y2=0
cc_536 N_A_1250_231#_c_624_n N_SET_B_c_779_n 0.0230707f $X=7.6 $Y=2.04 $X2=0
+ $Y2=0
cc_537 N_A_1250_231#_c_613_n N_SET_B_c_804_n 0.0152788f $X=8.755 $Y=1.82 $X2=0
+ $Y2=0
cc_538 N_A_1250_231#_c_625_n N_SET_B_c_804_n 0.0514033f $X=8.685 $Y=1.91 $X2=0
+ $Y2=0
cc_539 N_A_1250_231#_c_625_n N_SET_B_c_806_n 0.0120411f $X=8.685 $Y=1.91 $X2=0
+ $Y2=0
cc_540 N_A_1250_231#_c_613_n N_SET_B_c_782_n 0.00366867f $X=8.755 $Y=1.82 $X2=0
+ $Y2=0
cc_541 N_A_1250_231#_c_624_n N_A_1092_96#_c_951_n 0.0101997f $X=7.6 $Y=2.04
+ $X2=0 $Y2=0
cc_542 N_A_1250_231#_c_625_n N_A_1092_96#_c_951_n 0.0126355f $X=8.685 $Y=1.91
+ $X2=0 $Y2=0
cc_543 N_A_1250_231#_c_626_n N_A_1092_96#_c_951_n 0.00190786f $X=7.765 $Y=1.91
+ $X2=0 $Y2=0
cc_544 N_A_1250_231#_c_622_n N_A_1092_96#_c_952_n 0.00103236f $X=6.45 $Y=2.02
+ $X2=0 $Y2=0
cc_545 N_A_1250_231#_c_612_n N_A_1092_96#_c_941_n 0.00337742f $X=6.45 $Y=1.93
+ $X2=0 $Y2=0
cc_546 N_A_1250_231#_c_616_n N_A_1092_96#_c_941_n 0.0426566f $X=6.415 $Y=1.32
+ $X2=0 $Y2=0
cc_547 N_A_1250_231#_c_617_n N_A_1092_96#_c_941_n 0.0022803f $X=6.415 $Y=1.32
+ $X2=0 $Y2=0
cc_548 N_A_1250_231#_c_652_p N_A_1092_96#_c_941_n 0.00350049f $X=6.535 $Y=0.815
+ $X2=0 $Y2=0
cc_549 N_A_1250_231#_c_620_n N_A_1092_96#_c_941_n 0.00183057f $X=6.415 $Y=1.155
+ $X2=0 $Y2=0
cc_550 N_A_1250_231#_c_612_n N_A_1092_96#_c_953_n 0.00557547f $X=6.45 $Y=1.93
+ $X2=0 $Y2=0
cc_551 N_A_1250_231#_c_622_n N_A_1092_96#_c_953_n 0.00147337f $X=6.45 $Y=2.02
+ $X2=0 $Y2=0
cc_552 N_A_1250_231#_c_612_n N_A_1092_96#_c_942_n 0.0193831f $X=6.45 $Y=1.93
+ $X2=0 $Y2=0
cc_553 N_A_1250_231#_c_616_n N_A_1092_96#_c_942_n 0.0183691f $X=6.415 $Y=1.32
+ $X2=0 $Y2=0
cc_554 N_A_1250_231#_c_617_n N_A_1092_96#_c_942_n 0.00371918f $X=6.415 $Y=1.32
+ $X2=0 $Y2=0
cc_555 N_A_1250_231#_c_612_n N_A_1092_96#_c_943_n 0.00189752f $X=6.45 $Y=1.93
+ $X2=0 $Y2=0
cc_556 N_A_1250_231#_c_616_n N_A_1092_96#_c_943_n 0.0179367f $X=6.415 $Y=1.32
+ $X2=0 $Y2=0
cc_557 N_A_1250_231#_c_617_n N_A_1092_96#_c_943_n 0.00191992f $X=6.415 $Y=1.32
+ $X2=0 $Y2=0
cc_558 N_A_1250_231#_M1015_d N_A_1092_96#_c_944_n 0.00118937f $X=7.845 $Y=0.595
+ $X2=0 $Y2=0
cc_559 N_A_1250_231#_c_626_n N_A_1092_96#_c_944_n 0.00533796f $X=7.765 $Y=1.91
+ $X2=0 $Y2=0
cc_560 N_A_1250_231#_c_630_p N_A_1092_96#_c_944_n 0.0589129f $X=7.82 $Y=0.777
+ $X2=0 $Y2=0
cc_561 N_A_1250_231#_c_616_n N_A_1092_96#_c_945_n 0.0141814f $X=6.415 $Y=1.32
+ $X2=0 $Y2=0
cc_562 N_A_1250_231#_c_617_n N_A_1092_96#_c_945_n 7.47272e-19 $X=6.415 $Y=1.32
+ $X2=0 $Y2=0
cc_563 N_A_1250_231#_c_630_p N_A_1092_96#_c_945_n 0.013831f $X=7.82 $Y=0.777
+ $X2=0 $Y2=0
cc_564 N_A_1250_231#_c_620_n N_A_1092_96#_c_945_n 3.08362e-19 $X=6.415 $Y=1.155
+ $X2=0 $Y2=0
cc_565 N_A_1250_231#_c_625_n N_A_1092_96#_c_946_n 0.00843521f $X=8.685 $Y=1.91
+ $X2=0 $Y2=0
cc_566 N_A_1250_231#_c_626_n N_A_1092_96#_c_946_n 0.0119991f $X=7.765 $Y=1.91
+ $X2=0 $Y2=0
cc_567 N_A_1250_231#_c_626_n N_A_1092_96#_c_947_n 0.00112764f $X=7.765 $Y=1.91
+ $X2=0 $Y2=0
cc_568 N_A_1250_231#_c_630_p N_A_1092_96#_c_947_n 4.0724e-19 $X=7.82 $Y=0.777
+ $X2=0 $Y2=0
cc_569 N_A_1250_231#_c_673_p N_A_1092_96#_c_947_n 2.23578e-19 $X=8.15 $Y=0.777
+ $X2=0 $Y2=0
cc_570 N_A_1250_231#_c_652_p N_A_1092_96#_c_948_n 0.0108489f $X=6.535 $Y=0.815
+ $X2=0 $Y2=0
cc_571 N_A_1250_231#_c_620_n N_A_1092_96#_c_948_n 0.00290069f $X=6.415 $Y=1.155
+ $X2=0 $Y2=0
cc_572 N_A_1250_231#_c_630_p N_A_1092_96#_c_949_n 0.00885154f $X=7.82 $Y=0.777
+ $X2=0 $Y2=0
cc_573 N_A_1250_231#_c_673_p N_A_1092_96#_c_949_n 0.00424303f $X=8.15 $Y=0.777
+ $X2=0 $Y2=0
cc_574 N_A_1250_231#_c_613_n N_A_1625_93#_c_1059_n 0.00924456f $X=8.755 $Y=1.82
+ $X2=0 $Y2=0
cc_575 N_A_1250_231#_c_627_n N_A_1625_93#_c_1059_n 0.00138492f $X=8.85 $Y=1.825
+ $X2=0 $Y2=0
cc_576 N_A_1250_231#_c_613_n N_A_1625_93#_c_1074_n 0.0240739f $X=8.755 $Y=1.82
+ $X2=0 $Y2=0
cc_577 N_A_1250_231#_c_624_n N_A_1625_93#_c_1074_n 0.0010532f $X=7.6 $Y=2.04
+ $X2=0 $Y2=0
cc_578 N_A_1250_231#_c_625_n N_A_1625_93#_c_1074_n 0.0120766f $X=8.685 $Y=1.91
+ $X2=0 $Y2=0
cc_579 N_A_1250_231#_c_613_n N_A_1625_93#_c_1065_n 0.006929f $X=8.755 $Y=1.82
+ $X2=0 $Y2=0
cc_580 N_A_1250_231#_c_614_n N_A_1625_93#_c_1065_n 0.0162501f $X=9.25 $Y=1.295
+ $X2=0 $Y2=0
cc_581 N_A_1250_231#_c_625_n N_A_1625_93#_c_1065_n 0.00469137f $X=8.685 $Y=1.91
+ $X2=0 $Y2=0
cc_582 N_A_1250_231#_c_618_n N_A_1625_93#_c_1065_n 0.00534822f $X=8.685 $Y=0.815
+ $X2=0 $Y2=0
cc_583 N_A_1250_231#_c_687_p N_A_1625_93#_c_1065_n 0.0216998f $X=8.85 $Y=1.5
+ $X2=0 $Y2=0
cc_584 N_A_1250_231#_c_619_n N_A_1625_93#_c_1065_n 0.0137054f $X=8.85 $Y=1.335
+ $X2=0 $Y2=0
cc_585 N_A_1250_231#_c_613_n N_A_1625_93#_c_1066_n 8.06207e-19 $X=8.755 $Y=1.82
+ $X2=0 $Y2=0
cc_586 N_A_1250_231#_c_625_n N_A_1625_93#_c_1066_n 0.00245941f $X=8.685 $Y=1.91
+ $X2=0 $Y2=0
cc_587 N_A_1250_231#_c_618_n N_A_1625_93#_c_1066_n 0.00316048f $X=8.685 $Y=0.815
+ $X2=0 $Y2=0
cc_588 N_A_1250_231#_c_687_p N_A_1625_93#_c_1066_n 0.00132788f $X=8.85 $Y=1.5
+ $X2=0 $Y2=0
cc_589 N_A_1250_231#_c_619_n N_A_1625_93#_c_1066_n 0.00132903f $X=8.85 $Y=1.335
+ $X2=0 $Y2=0
cc_590 N_A_1250_231#_c_613_n N_A_1625_93#_c_1067_n 0.00204231f $X=8.755 $Y=1.82
+ $X2=0 $Y2=0
cc_591 N_A_1250_231#_c_625_n N_A_1625_93#_c_1067_n 0.0212526f $X=8.685 $Y=1.91
+ $X2=0 $Y2=0
cc_592 N_A_1250_231#_c_673_p N_A_1625_93#_c_1067_n 0.0155144f $X=8.15 $Y=0.777
+ $X2=0 $Y2=0
cc_593 N_A_1250_231#_c_619_n N_A_1625_93#_c_1067_n 0.0295318f $X=8.85 $Y=1.335
+ $X2=0 $Y2=0
cc_594 N_A_1250_231#_c_613_n N_A_1625_93#_c_1071_n 0.0213532f $X=8.755 $Y=1.82
+ $X2=0 $Y2=0
cc_595 N_A_1250_231#_c_625_n N_A_1625_93#_c_1071_n 9.74547e-19 $X=8.685 $Y=1.91
+ $X2=0 $Y2=0
cc_596 N_A_1250_231#_c_618_n N_A_1625_93#_c_1071_n 8.36667e-19 $X=8.685 $Y=0.815
+ $X2=0 $Y2=0
cc_597 N_A_1250_231#_c_619_n N_A_1625_93#_c_1071_n 4.08406e-19 $X=8.85 $Y=1.335
+ $X2=0 $Y2=0
cc_598 N_A_1250_231#_c_613_n N_A_1625_93#_c_1072_n 0.00110147f $X=8.755 $Y=1.82
+ $X2=0 $Y2=0
cc_599 N_A_1250_231#_c_618_n N_A_1625_93#_c_1072_n 0.00999322f $X=8.685 $Y=0.815
+ $X2=0 $Y2=0
cc_600 N_A_1250_231#_c_673_p N_A_1625_93#_c_1072_n 0.00434626f $X=8.15 $Y=0.777
+ $X2=0 $Y2=0
cc_601 N_A_1250_231#_c_619_n N_A_1625_93#_c_1072_n 0.00762936f $X=8.85 $Y=1.335
+ $X2=0 $Y2=0
cc_602 N_A_1250_231#_c_622_n N_A_622_98#_c_1222_n 0.00284772f $X=6.45 $Y=2.02
+ $X2=0 $Y2=0
cc_603 N_A_1250_231#_c_622_n N_A_622_98#_c_1224_n 0.0274712f $X=6.45 $Y=2.02
+ $X2=0 $Y2=0
cc_604 N_A_1250_231#_c_622_n N_A_622_98#_c_1225_n 0.00495681f $X=6.45 $Y=2.02
+ $X2=0 $Y2=0
cc_605 N_A_1250_231#_c_613_n N_A_622_98#_c_1225_n 0.0104018f $X=8.755 $Y=1.82
+ $X2=0 $Y2=0
cc_606 N_A_1250_231#_c_613_n N_A_622_98#_c_1204_n 0.0135472f $X=8.755 $Y=1.82
+ $X2=0 $Y2=0
cc_607 N_A_1250_231#_c_614_n N_A_622_98#_c_1204_n 0.00988849f $X=9.25 $Y=1.295
+ $X2=0 $Y2=0
cc_608 N_A_1250_231#_c_625_n N_A_622_98#_c_1204_n 0.00254788f $X=8.685 $Y=1.91
+ $X2=0 $Y2=0
cc_609 N_A_1250_231#_c_627_n N_A_622_98#_c_1204_n 0.00150525f $X=8.85 $Y=1.825
+ $X2=0 $Y2=0
cc_610 N_A_1250_231#_c_613_n N_A_622_98#_M1008_g 0.0195888f $X=8.755 $Y=1.82
+ $X2=0 $Y2=0
cc_611 N_A_1250_231#_c_613_n N_A_622_98#_c_1208_n 4.51932e-19 $X=8.755 $Y=1.82
+ $X2=0 $Y2=0
cc_612 N_A_1250_231#_c_625_n N_A_622_98#_c_1208_n 0.00741276f $X=8.685 $Y=1.91
+ $X2=0 $Y2=0
cc_613 N_A_1250_231#_c_627_n N_A_622_98#_c_1208_n 0.0145976f $X=8.85 $Y=1.825
+ $X2=0 $Y2=0
cc_614 N_A_1250_231#_c_615_n N_A_622_98#_c_1215_n 0.00468731f $X=9.325 $Y=1.22
+ $X2=0 $Y2=0
cc_615 N_A_1250_231#_c_619_n N_A_622_98#_c_1215_n 0.0055458f $X=8.85 $Y=1.335
+ $X2=0 $Y2=0
cc_616 N_A_1250_231#_c_613_n N_A_622_98#_c_1216_n 0.00530265f $X=8.755 $Y=1.82
+ $X2=0 $Y2=0
cc_617 N_A_1250_231#_c_614_n N_A_622_98#_c_1216_n 0.00592053f $X=9.25 $Y=1.295
+ $X2=0 $Y2=0
cc_618 N_A_1250_231#_c_687_p N_A_622_98#_c_1216_n 0.0145976f $X=8.85 $Y=1.5
+ $X2=0 $Y2=0
cc_619 N_A_1250_231#_c_612_n N_A_877_98#_c_1441_n 7.51872e-19 $X=6.45 $Y=1.93
+ $X2=0 $Y2=0
cc_620 N_A_1250_231#_c_616_n N_A_877_98#_M1030_g 5.48859e-19 $X=6.415 $Y=1.32
+ $X2=0 $Y2=0
cc_621 N_A_1250_231#_c_617_n N_A_877_98#_M1030_g 0.013411f $X=6.415 $Y=1.32
+ $X2=0 $Y2=0
cc_622 N_A_1250_231#_c_620_n N_A_877_98#_M1030_g 0.0226694f $X=6.415 $Y=1.155
+ $X2=0 $Y2=0
cc_623 N_A_1250_231#_c_615_n N_A_877_98#_c_1443_n 0.0103107f $X=9.325 $Y=1.22
+ $X2=0 $Y2=0
cc_624 N_A_1250_231#_c_652_p N_A_877_98#_c_1443_n 5.19956e-19 $X=6.535 $Y=0.815
+ $X2=0 $Y2=0
cc_625 N_A_1250_231#_c_618_n N_A_877_98#_c_1443_n 0.00256696f $X=8.685 $Y=0.815
+ $X2=0 $Y2=0
cc_626 N_A_1250_231#_c_630_p N_A_877_98#_c_1443_n 0.0029304f $X=7.82 $Y=0.777
+ $X2=0 $Y2=0
cc_627 N_A_1250_231#_c_620_n N_A_877_98#_c_1443_n 0.00852452f $X=6.415 $Y=1.155
+ $X2=0 $Y2=0
cc_628 N_A_1250_231#_c_615_n N_A_877_98#_M1001_g 0.027011f $X=9.325 $Y=1.22
+ $X2=0 $Y2=0
cc_629 N_A_1250_231#_c_614_n N_A_877_98#_c_1446_n 0.027011f $X=9.25 $Y=1.295
+ $X2=0 $Y2=0
cc_630 N_A_1250_231#_c_613_n N_A_1878_420#_c_1784_n 5.45049e-19 $X=8.755 $Y=1.82
+ $X2=0 $Y2=0
cc_631 N_A_1250_231#_c_625_n N_VPWR_M1033_d 0.0026214f $X=8.685 $Y=1.91 $X2=0
+ $Y2=0
cc_632 N_A_1250_231#_c_622_n N_VPWR_c_2016_n 0.0107964f $X=6.45 $Y=2.02 $X2=0
+ $Y2=0
cc_633 N_A_1250_231#_c_613_n N_VPWR_c_2017_n 0.00505774f $X=8.755 $Y=1.82 $X2=0
+ $Y2=0
cc_634 N_A_1250_231#_c_622_n N_VPWR_c_2012_n 9.72468e-19 $X=6.45 $Y=2.02 $X2=0
+ $Y2=0
cc_635 N_A_1250_231#_c_613_n N_VPWR_c_2012_n 9.14192e-19 $X=8.755 $Y=1.82 $X2=0
+ $Y2=0
cc_636 N_A_1250_231#_c_612_n N_A_197_119#_c_2203_n 7.3128e-19 $X=6.45 $Y=1.93
+ $X2=0 $Y2=0
cc_637 N_A_1250_231#_c_625_n A_1580_379# 0.00165852f $X=8.685 $Y=1.91 $X2=-0.19
+ $Y2=-0.245
cc_638 N_A_1250_231#_c_625_n A_1766_379# 0.00263617f $X=8.685 $Y=1.91 $X2=-0.19
+ $Y2=-0.245
cc_639 N_A_1250_231#_c_616_n N_VGND_M1046_d 0.00212348f $X=6.415 $Y=1.32 $X2=0
+ $Y2=0
cc_640 N_A_1250_231#_c_652_p N_VGND_M1046_d 4.09279e-19 $X=6.535 $Y=0.815 $X2=0
+ $Y2=0
cc_641 N_A_1250_231#_c_630_p N_VGND_M1046_d 0.0117278f $X=7.82 $Y=0.777 $X2=0
+ $Y2=0
cc_642 N_A_1250_231#_c_617_n N_VGND_c_2433_n 2.19791e-19 $X=6.415 $Y=1.32 $X2=0
+ $Y2=0
cc_643 N_A_1250_231#_c_652_p N_VGND_c_2433_n 0.0037988f $X=6.535 $Y=0.815 $X2=0
+ $Y2=0
cc_644 N_A_1250_231#_c_630_p N_VGND_c_2433_n 0.0273008f $X=7.82 $Y=0.777 $X2=0
+ $Y2=0
cc_645 N_A_1250_231#_c_620_n N_VGND_c_2433_n 0.00113285f $X=6.415 $Y=1.155 $X2=0
+ $Y2=0
cc_646 N_A_1250_231#_c_614_n N_VGND_c_2434_n 0.00781231f $X=9.25 $Y=1.295 $X2=0
+ $Y2=0
cc_647 N_A_1250_231#_c_615_n N_VGND_c_2434_n 0.0101025f $X=9.325 $Y=1.22 $X2=0
+ $Y2=0
cc_648 N_A_1250_231#_c_618_n N_VGND_c_2434_n 0.0145003f $X=8.685 $Y=0.815 $X2=0
+ $Y2=0
cc_649 N_A_1250_231#_c_619_n N_VGND_c_2434_n 0.011381f $X=8.85 $Y=1.335 $X2=0
+ $Y2=0
cc_650 N_A_1250_231#_c_652_p N_VGND_c_2440_n 0.00245352f $X=6.535 $Y=0.815 $X2=0
+ $Y2=0
cc_651 N_A_1250_231#_c_618_n N_VGND_c_2442_n 0.0023514f $X=8.685 $Y=0.815 $X2=0
+ $Y2=0
cc_652 N_A_1250_231#_c_630_p N_VGND_c_2442_n 0.00281701f $X=7.82 $Y=0.777 $X2=0
+ $Y2=0
cc_653 N_A_1250_231#_c_615_n N_VGND_c_2451_n 7.88961e-19 $X=9.325 $Y=1.22 $X2=0
+ $Y2=0
cc_654 N_A_1250_231#_c_652_p N_VGND_c_2451_n 0.00481003f $X=6.535 $Y=0.815 $X2=0
+ $Y2=0
cc_655 N_A_1250_231#_c_618_n N_VGND_c_2451_n 0.00348353f $X=8.685 $Y=0.815 $X2=0
+ $Y2=0
cc_656 N_A_1250_231#_c_630_p N_VGND_c_2451_n 0.00828529f $X=7.82 $Y=0.777 $X2=0
+ $Y2=0
cc_657 N_A_1250_231#_c_620_n N_VGND_c_2451_n 9.49986e-19 $X=6.415 $Y=1.155 $X2=0
+ $Y2=0
cc_658 N_A_1250_231#_c_630_p N_A_1418_125#_M1022_d 0.0116116f $X=7.82 $Y=0.777
+ $X2=-0.19 $Y2=-0.245
cc_659 N_A_1250_231#_c_618_n N_A_1418_125#_M1016_d 0.00991095f $X=8.685 $Y=0.815
+ $X2=0 $Y2=0
cc_660 N_A_1250_231#_c_619_n N_A_1418_125#_M1016_d 0.00353615f $X=8.85 $Y=1.335
+ $X2=0 $Y2=0
cc_661 N_A_1250_231#_c_630_p N_A_1418_125#_c_2600_n 0.0355643f $X=7.82 $Y=0.777
+ $X2=0 $Y2=0
cc_662 N_A_1250_231#_c_615_n N_A_1418_125#_c_2602_n 4.33749e-19 $X=9.325 $Y=1.22
+ $X2=0 $Y2=0
cc_663 N_A_1250_231#_c_618_n N_A_1418_125#_c_2602_n 0.0279844f $X=8.685 $Y=0.815
+ $X2=0 $Y2=0
cc_664 N_A_1250_231#_c_618_n N_A_1418_125#_c_2603_n 0.00722944f $X=8.685
+ $Y=0.815 $X2=0 $Y2=0
cc_665 N_A_1250_231#_c_630_p N_A_1418_125#_c_2603_n 0.00722944f $X=7.82 $Y=0.777
+ $X2=0 $Y2=0
cc_666 N_A_1250_231#_c_673_p N_A_1418_125#_c_2603_n 0.0190774f $X=8.15 $Y=0.777
+ $X2=0 $Y2=0
cc_667 N_SET_B_c_772_n N_A_1092_96#_c_940_n 0.00873347f $X=7.285 $Y=1.82 $X2=0
+ $Y2=0
cc_668 N_SET_B_c_778_n N_A_1092_96#_c_940_n 8.15264e-19 $X=7.18 $Y=2.905 $X2=0
+ $Y2=0
cc_669 N_SET_B_c_810_p N_A_1092_96#_c_940_n 4.19145e-19 $X=7.21 $Y=1.535 $X2=0
+ $Y2=0
cc_670 N_SET_B_c_772_n N_A_1092_96#_c_951_n 0.0164604f $X=7.285 $Y=1.82 $X2=0
+ $Y2=0
cc_671 N_SET_B_c_778_n N_A_1092_96#_c_951_n 7.67235e-19 $X=7.18 $Y=2.905 $X2=0
+ $Y2=0
cc_672 N_SET_B_c_779_n N_A_1092_96#_c_951_n 0.00347797f $X=7.935 $Y=2.99 $X2=0
+ $Y2=0
cc_673 N_SET_B_c_781_n N_A_1092_96#_c_951_n 0.00343421f $X=8.02 $Y=2.905 $X2=0
+ $Y2=0
cc_674 N_SET_B_c_772_n N_A_1092_96#_c_942_n 0.00104761f $X=7.285 $Y=1.82 $X2=0
+ $Y2=0
cc_675 N_SET_B_c_778_n N_A_1092_96#_c_942_n 0.0117718f $X=7.18 $Y=2.905 $X2=0
+ $Y2=0
cc_676 N_SET_B_M1022_g N_A_1092_96#_c_943_n 0.00657656f $X=7.015 $Y=0.9 $X2=0
+ $Y2=0
cc_677 N_SET_B_c_810_p N_A_1092_96#_c_943_n 0.0183734f $X=7.21 $Y=1.535 $X2=0
+ $Y2=0
cc_678 N_SET_B_M1022_g N_A_1092_96#_c_944_n 0.0147347f $X=7.015 $Y=0.9 $X2=0
+ $Y2=0
cc_679 N_SET_B_c_772_n N_A_1092_96#_c_944_n 0.00737349f $X=7.285 $Y=1.82 $X2=0
+ $Y2=0
cc_680 N_SET_B_c_810_p N_A_1092_96#_c_944_n 0.0250891f $X=7.21 $Y=1.535 $X2=0
+ $Y2=0
cc_681 N_SET_B_M1022_g N_A_1092_96#_c_946_n 8.70544e-19 $X=7.015 $Y=0.9 $X2=0
+ $Y2=0
cc_682 N_SET_B_c_772_n N_A_1092_96#_c_946_n 9.34747e-19 $X=7.285 $Y=1.82 $X2=0
+ $Y2=0
cc_683 N_SET_B_c_810_p N_A_1092_96#_c_946_n 0.0110904f $X=7.21 $Y=1.535 $X2=0
+ $Y2=0
cc_684 N_SET_B_M1022_g N_A_1092_96#_c_947_n 0.00304624f $X=7.015 $Y=0.9 $X2=0
+ $Y2=0
cc_685 N_SET_B_c_772_n N_A_1092_96#_c_947_n 0.013649f $X=7.285 $Y=1.82 $X2=0
+ $Y2=0
cc_686 N_SET_B_c_810_p N_A_1092_96#_c_947_n 6.09509e-19 $X=7.21 $Y=1.535 $X2=0
+ $Y2=0
cc_687 N_SET_B_M1022_g N_A_1092_96#_c_949_n 0.0139641f $X=7.015 $Y=0.9 $X2=0
+ $Y2=0
cc_688 N_SET_B_c_781_n N_A_1625_93#_c_1074_n 0.00658823f $X=8.02 $Y=2.905 $X2=0
+ $Y2=0
cc_689 N_SET_B_c_804_n N_A_1625_93#_c_1074_n 0.0144616f $X=8.855 $Y=2.25 $X2=0
+ $Y2=0
cc_690 N_SET_B_M1002_g N_A_1625_93#_c_1065_n 0.00150429f $X=11.28 $Y=0.74 $X2=0
+ $Y2=0
cc_691 N_SET_B_c_774_n N_A_1625_93#_c_1065_n 0.00458846f $X=11.295 $Y=1.885
+ $X2=0 $Y2=0
cc_692 N_SET_B_c_786_n N_A_1625_93#_c_1065_n 0.00707697f $X=11.055 $Y=1.775
+ $X2=0 $Y2=0
cc_693 N_SET_B_c_787_n N_A_1625_93#_c_1065_n 0.00102133f $X=10.295 $Y=1.775
+ $X2=0 $Y2=0
cc_694 SET_B N_A_1625_93#_c_1065_n 0.00802342f $X=11.195 $Y=1.95 $X2=0 $Y2=0
cc_695 N_SET_B_c_772_n N_A_622_98#_c_1225_n 0.00915973f $X=7.285 $Y=1.82 $X2=0
+ $Y2=0
cc_696 N_SET_B_c_779_n N_A_622_98#_c_1225_n 0.0158397f $X=7.935 $Y=2.99 $X2=0
+ $Y2=0
cc_697 N_SET_B_c_780_n N_A_622_98#_c_1225_n 0.00328385f $X=7.265 $Y=2.99 $X2=0
+ $Y2=0
cc_698 N_SET_B_c_783_n N_A_622_98#_c_1225_n 0.00977019f $X=10.095 $Y=2.99 $X2=0
+ $Y2=0
cc_699 N_SET_B_c_784_n N_A_622_98#_c_1225_n 0.00420304f $X=9.025 $Y=2.99 $X2=0
+ $Y2=0
cc_700 N_SET_B_c_804_n N_A_622_98#_M1008_g 0.00163974f $X=8.855 $Y=2.25 $X2=0
+ $Y2=0
cc_701 N_SET_B_c_782_n N_A_622_98#_M1008_g 0.00723827f $X=8.94 $Y=2.905 $X2=0
+ $Y2=0
cc_702 N_SET_B_c_783_n N_A_622_98#_M1008_g 0.0116574f $X=10.095 $Y=2.99 $X2=0
+ $Y2=0
cc_703 N_SET_B_M1022_g N_A_877_98#_c_1443_n 0.00848668f $X=7.015 $Y=0.9 $X2=0
+ $Y2=0
cc_704 N_SET_B_c_783_n N_A_877_98#_c_1453_n 0.0109203f $X=10.095 $Y=2.99 $X2=0
+ $Y2=0
cc_705 N_SET_B_c_785_n N_A_877_98#_c_1453_n 0.00661524f $X=10.18 $Y=2.905 $X2=0
+ $Y2=0
cc_706 N_SET_B_c_787_n N_A_877_98#_c_1447_n 0.00151263f $X=10.295 $Y=1.775 $X2=0
+ $Y2=0
cc_707 N_SET_B_c_788_n N_A_877_98#_c_1447_n 0.00297299f $X=10.195 $Y=2.015 $X2=0
+ $Y2=0
cc_708 N_SET_B_c_789_n N_A_877_98#_c_1447_n 0.00152793f $X=10.195 $Y=2.185 $X2=0
+ $Y2=0
cc_709 N_SET_B_c_783_n N_A_2037_442#_c_1601_n 0.00498681f $X=10.095 $Y=2.99
+ $X2=0 $Y2=0
cc_710 N_SET_B_c_785_n N_A_2037_442#_c_1601_n 0.0140746f $X=10.18 $Y=2.905 $X2=0
+ $Y2=0
cc_711 N_SET_B_M1002_g N_A_2037_442#_M1047_g 0.0263216f $X=11.28 $Y=0.74 $X2=0
+ $Y2=0
cc_712 N_SET_B_c_774_n N_A_2037_442#_M1047_g 0.0372135f $X=11.295 $Y=1.885 $X2=0
+ $Y2=0
cc_713 N_SET_B_c_786_n N_A_2037_442#_M1047_g 0.0125961f $X=11.055 $Y=1.775 $X2=0
+ $Y2=0
cc_714 N_SET_B_c_788_n N_A_2037_442#_M1047_g 0.00452974f $X=10.195 $Y=2.015
+ $X2=0 $Y2=0
cc_715 SET_B N_A_2037_442#_M1047_g 0.00606634f $X=11.195 $Y=1.95 $X2=0 $Y2=0
cc_716 N_SET_B_c_774_n N_A_2037_442#_c_1608_n 0.0143477f $X=11.295 $Y=1.885
+ $X2=0 $Y2=0
cc_717 N_SET_B_c_786_n N_A_2037_442#_c_1608_n 0.00928944f $X=11.055 $Y=1.775
+ $X2=0 $Y2=0
cc_718 SET_B N_A_2037_442#_c_1608_n 0.0200692f $X=11.195 $Y=1.95 $X2=0 $Y2=0
cc_719 SET_B N_A_2037_442#_c_1598_n 0.0067676f $X=11.195 $Y=1.95 $X2=0 $Y2=0
cc_720 N_SET_B_c_774_n N_A_2037_442#_c_1626_n 0.00624182f $X=11.295 $Y=1.885
+ $X2=0 $Y2=0
cc_721 SET_B N_A_2037_442#_c_1626_n 0.0148744f $X=11.195 $Y=1.95 $X2=0 $Y2=0
cc_722 N_SET_B_c_774_n N_A_2037_442#_c_1612_n 0.00139265f $X=11.295 $Y=1.885
+ $X2=0 $Y2=0
cc_723 N_SET_B_c_785_n N_A_2037_442#_c_1612_n 0.019698f $X=10.18 $Y=2.905 $X2=0
+ $Y2=0
cc_724 N_SET_B_c_786_n N_A_2037_442#_c_1612_n 0.0250442f $X=11.055 $Y=1.775
+ $X2=0 $Y2=0
cc_725 N_SET_B_c_789_n N_A_2037_442#_c_1612_n 0.0117952f $X=10.195 $Y=2.185
+ $X2=0 $Y2=0
cc_726 SET_B N_A_2037_442#_c_1612_n 0.00671591f $X=11.195 $Y=1.95 $X2=0 $Y2=0
cc_727 N_SET_B_c_785_n N_A_2037_442#_c_1613_n 0.00821331f $X=10.18 $Y=2.905
+ $X2=0 $Y2=0
cc_728 N_SET_B_c_786_n N_A_2037_442#_c_1613_n 0.00675887f $X=11.055 $Y=1.775
+ $X2=0 $Y2=0
cc_729 N_SET_B_c_789_n N_A_2037_442#_c_1613_n 0.0030167f $X=10.195 $Y=2.185
+ $X2=0 $Y2=0
cc_730 N_SET_B_c_774_n N_A_2037_442#_c_1614_n 0.0070934f $X=11.295 $Y=1.885
+ $X2=0 $Y2=0
cc_731 N_SET_B_c_783_n N_A_1878_420#_M1008_d 0.00296216f $X=10.095 $Y=2.99 $X2=0
+ $Y2=0
cc_732 N_SET_B_M1002_g N_A_1878_420#_c_1772_n 0.0123775f $X=11.28 $Y=0.74 $X2=0
+ $Y2=0
cc_733 N_SET_B_M1002_g N_A_1878_420#_c_1773_n 0.0138767f $X=11.28 $Y=0.74 $X2=0
+ $Y2=0
cc_734 N_SET_B_c_774_n N_A_1878_420#_c_1773_n 0.0151932f $X=11.295 $Y=1.885
+ $X2=0 $Y2=0
cc_735 SET_B N_A_1878_420#_c_1773_n 0.00112454f $X=11.195 $Y=1.95 $X2=0 $Y2=0
cc_736 N_SET_B_c_774_n N_A_1878_420#_c_1783_n 0.0174703f $X=11.295 $Y=1.885
+ $X2=0 $Y2=0
cc_737 SET_B N_A_1878_420#_c_1783_n 9.37463e-19 $X=11.195 $Y=1.95 $X2=0 $Y2=0
cc_738 N_SET_B_c_786_n N_A_1878_420#_c_1776_n 0.0294373f $X=11.055 $Y=1.775
+ $X2=0 $Y2=0
cc_739 N_SET_B_c_787_n N_A_1878_420#_c_1776_n 0.0133014f $X=10.295 $Y=1.775
+ $X2=0 $Y2=0
cc_740 N_SET_B_c_789_n N_A_1878_420#_c_1776_n 0.00116624f $X=10.195 $Y=2.185
+ $X2=0 $Y2=0
cc_741 N_SET_B_M1002_g N_A_1878_420#_c_1777_n 0.01317f $X=11.28 $Y=0.74 $X2=0
+ $Y2=0
cc_742 N_SET_B_c_774_n N_A_1878_420#_c_1777_n 0.00427702f $X=11.295 $Y=1.885
+ $X2=0 $Y2=0
cc_743 N_SET_B_c_786_n N_A_1878_420#_c_1777_n 0.00554997f $X=11.055 $Y=1.775
+ $X2=0 $Y2=0
cc_744 SET_B N_A_1878_420#_c_1777_n 0.0222931f $X=11.195 $Y=1.95 $X2=0 $Y2=0
cc_745 N_SET_B_c_804_n N_A_1878_420#_c_1784_n 0.00834819f $X=8.855 $Y=2.25 $X2=0
+ $Y2=0
cc_746 N_SET_B_c_782_n N_A_1878_420#_c_1784_n 0.0176104f $X=8.94 $Y=2.905 $X2=0
+ $Y2=0
cc_747 N_SET_B_c_783_n N_A_1878_420#_c_1784_n 0.0320856f $X=10.095 $Y=2.99 $X2=0
+ $Y2=0
cc_748 N_SET_B_c_785_n N_A_1878_420#_c_1784_n 0.0276978f $X=10.18 $Y=2.905 $X2=0
+ $Y2=0
cc_749 N_SET_B_c_787_n N_A_1878_420#_c_1785_n 0.00104181f $X=10.295 $Y=1.775
+ $X2=0 $Y2=0
cc_750 N_SET_B_c_788_n N_A_1878_420#_c_1785_n 0.00974859f $X=10.195 $Y=2.015
+ $X2=0 $Y2=0
cc_751 N_SET_B_c_789_n N_A_1878_420#_c_1785_n 0.0276978f $X=10.195 $Y=2.185
+ $X2=0 $Y2=0
cc_752 N_SET_B_c_787_n N_A_1878_420#_c_1787_n 0.013235f $X=10.295 $Y=1.775 $X2=0
+ $Y2=0
cc_753 N_SET_B_M1002_g N_A_1878_420#_c_1780_n 0.00220582f $X=11.28 $Y=0.74 $X2=0
+ $Y2=0
cc_754 N_SET_B_c_774_n N_A_1878_420#_c_1780_n 0.00102095f $X=11.295 $Y=1.885
+ $X2=0 $Y2=0
cc_755 N_SET_B_c_786_n N_A_1878_420#_c_1780_n 0.0116578f $X=11.055 $Y=1.775
+ $X2=0 $Y2=0
cc_756 N_SET_B_M1002_g N_A_1878_420#_c_1781_n 9.59139e-19 $X=11.28 $Y=0.74 $X2=0
+ $Y2=0
cc_757 N_SET_B_c_774_n N_A_1878_420#_c_1781_n 3.95637e-19 $X=11.295 $Y=1.885
+ $X2=0 $Y2=0
cc_758 SET_B N_A_1878_420#_c_1781_n 0.00188563f $X=11.195 $Y=1.95 $X2=0 $Y2=0
cc_759 N_SET_B_c_778_n N_VPWR_M1045_d 0.00938801f $X=7.18 $Y=2.905 $X2=0 $Y2=0
cc_760 N_SET_B_c_804_n N_VPWR_M1033_d 0.00516133f $X=8.855 $Y=2.25 $X2=0 $Y2=0
cc_761 SET_B N_VPWR_M1036_d 0.00332263f $X=11.195 $Y=1.95 $X2=0 $Y2=0
cc_762 N_SET_B_c_772_n N_VPWR_c_2016_n 0.003189f $X=7.285 $Y=1.82 $X2=0 $Y2=0
cc_763 N_SET_B_c_778_n N_VPWR_c_2016_n 0.0639085f $X=7.18 $Y=2.905 $X2=0 $Y2=0
cc_764 N_SET_B_c_780_n N_VPWR_c_2016_n 0.0150385f $X=7.265 $Y=2.99 $X2=0 $Y2=0
cc_765 N_SET_B_c_779_n N_VPWR_c_2017_n 0.0130647f $X=7.935 $Y=2.99 $X2=0 $Y2=0
cc_766 N_SET_B_c_781_n N_VPWR_c_2017_n 0.0256951f $X=8.02 $Y=2.905 $X2=0 $Y2=0
cc_767 N_SET_B_c_804_n N_VPWR_c_2017_n 0.0205394f $X=8.855 $Y=2.25 $X2=0 $Y2=0
cc_768 N_SET_B_c_782_n N_VPWR_c_2017_n 0.0217628f $X=8.94 $Y=2.905 $X2=0 $Y2=0
cc_769 N_SET_B_c_784_n N_VPWR_c_2017_n 0.0151624f $X=9.025 $Y=2.99 $X2=0 $Y2=0
cc_770 N_SET_B_c_774_n N_VPWR_c_2023_n 0.00461464f $X=11.295 $Y=1.885 $X2=0
+ $Y2=0
cc_771 N_SET_B_c_779_n N_VPWR_c_2030_n 0.0546768f $X=7.935 $Y=2.99 $X2=0 $Y2=0
cc_772 N_SET_B_c_780_n N_VPWR_c_2030_n 0.0115893f $X=7.265 $Y=2.99 $X2=0 $Y2=0
cc_773 N_SET_B_c_774_n N_VPWR_c_2012_n 0.0047002f $X=11.295 $Y=1.885 $X2=0 $Y2=0
cc_774 N_SET_B_c_779_n N_VPWR_c_2012_n 0.028344f $X=7.935 $Y=2.99 $X2=0 $Y2=0
cc_775 N_SET_B_c_780_n N_VPWR_c_2012_n 0.00583135f $X=7.265 $Y=2.99 $X2=0 $Y2=0
cc_776 N_SET_B_c_783_n N_VPWR_c_2012_n 0.0451852f $X=10.095 $Y=2.99 $X2=0 $Y2=0
cc_777 N_SET_B_c_784_n N_VPWR_c_2012_n 0.00583135f $X=9.025 $Y=2.99 $X2=0 $Y2=0
cc_778 N_SET_B_c_783_n N_VPWR_c_2038_n 0.0805277f $X=10.095 $Y=2.99 $X2=0 $Y2=0
cc_779 N_SET_B_c_784_n N_VPWR_c_2038_n 0.0115893f $X=9.025 $Y=2.99 $X2=0 $Y2=0
cc_780 N_SET_B_c_774_n N_VPWR_c_2039_n 0.0134607f $X=11.295 $Y=1.885 $X2=0 $Y2=0
cc_781 N_SET_B_c_783_n N_VPWR_c_2039_n 0.0151761f $X=10.095 $Y=2.99 $X2=0 $Y2=0
cc_782 N_SET_B_c_785_n N_VPWR_c_2039_n 0.0193067f $X=10.18 $Y=2.905 $X2=0 $Y2=0
cc_783 N_SET_B_c_781_n A_1580_379# 0.00601775f $X=8.02 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_784 N_SET_B_c_804_n A_1580_379# 3.41682e-19 $X=8.855 $Y=2.25 $X2=-0.19
+ $Y2=-0.245
cc_785 N_SET_B_c_806_n A_1580_379# 0.00193591f $X=8.105 $Y=2.25 $X2=-0.19
+ $Y2=-0.245
cc_786 N_SET_B_c_804_n A_1766_379# 0.00387807f $X=8.855 $Y=2.25 $X2=-0.19
+ $Y2=-0.245
cc_787 N_SET_B_c_782_n A_1766_379# 0.0088731f $X=8.94 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_788 N_SET_B_c_783_n A_1766_379# 0.00602618f $X=10.095 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_789 N_SET_B_c_783_n A_1986_504# 0.00408264f $X=10.095 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_790 N_SET_B_c_785_n A_1986_504# 0.00375007f $X=10.18 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_791 N_SET_B_M1022_g N_VGND_c_2433_n 7.8833e-19 $X=7.015 $Y=0.9 $X2=0 $Y2=0
cc_792 N_SET_B_M1002_g N_VGND_c_2435_n 0.0013418f $X=11.28 $Y=0.74 $X2=0 $Y2=0
cc_793 N_SET_B_M1002_g N_VGND_c_2446_n 0.00430908f $X=11.28 $Y=0.74 $X2=0 $Y2=0
cc_794 N_SET_B_M1022_g N_VGND_c_2451_n 9.49986e-19 $X=7.015 $Y=0.9 $X2=0 $Y2=0
cc_795 N_SET_B_M1002_g N_VGND_c_2451_n 0.00816573f $X=11.28 $Y=0.74 $X2=0 $Y2=0
cc_796 N_SET_B_M1022_g N_A_1418_125#_c_2600_n 8.42727e-19 $X=7.015 $Y=0.9 $X2=0
+ $Y2=0
cc_797 N_SET_B_M1002_g N_A_2271_74#_c_2628_n 0.0067893f $X=11.28 $Y=0.74 $X2=0
+ $Y2=0
cc_798 N_SET_B_M1002_g N_A_2271_74#_c_2627_n 0.00325143f $X=11.28 $Y=0.74 $X2=0
+ $Y2=0
cc_799 N_A_1092_96#_c_940_n N_A_1625_93#_c_1059_n 0.00699503f $X=7.825 $Y=1.73
+ $X2=0 $Y2=0
cc_800 N_A_1092_96#_c_951_n N_A_1625_93#_c_1074_n 0.0499177f $X=7.825 $Y=1.82
+ $X2=0 $Y2=0
cc_801 N_A_1092_96#_c_944_n N_A_1625_93#_c_1066_n 3.76443e-19 $X=7.585 $Y=1.155
+ $X2=0 $Y2=0
cc_802 N_A_1092_96#_c_946_n N_A_1625_93#_c_1066_n 8.94149e-19 $X=7.75 $Y=1.42
+ $X2=0 $Y2=0
cc_803 N_A_1092_96#_c_944_n N_A_1625_93#_c_1067_n 0.00393432f $X=7.585 $Y=1.155
+ $X2=0 $Y2=0
cc_804 N_A_1092_96#_c_946_n N_A_1625_93#_c_1067_n 0.0211611f $X=7.75 $Y=1.42
+ $X2=0 $Y2=0
cc_805 N_A_1092_96#_c_947_n N_A_1625_93#_c_1067_n 0.00114848f $X=7.75 $Y=1.42
+ $X2=0 $Y2=0
cc_806 N_A_1092_96#_c_946_n N_A_1625_93#_c_1071_n 0.00114936f $X=7.75 $Y=1.42
+ $X2=0 $Y2=0
cc_807 N_A_1092_96#_c_947_n N_A_1625_93#_c_1071_n 0.0201104f $X=7.75 $Y=1.42
+ $X2=0 $Y2=0
cc_808 N_A_1092_96#_c_944_n N_A_1625_93#_c_1072_n 0.00328085f $X=7.585 $Y=1.155
+ $X2=0 $Y2=0
cc_809 N_A_1092_96#_c_949_n N_A_1625_93#_c_1072_n 0.0184197f $X=7.75 $Y=1.255
+ $X2=0 $Y2=0
cc_810 N_A_1092_96#_c_952_n N_A_622_98#_c_1220_n 0.00662969f $X=5.955 $Y=2.37
+ $X2=0 $Y2=0
cc_811 N_A_1092_96#_c_941_n N_A_622_98#_c_1203_n 5.10155e-19 $X=6.04 $Y=1.655
+ $X2=0 $Y2=0
cc_812 N_A_1092_96#_c_948_n N_A_622_98#_c_1203_n 0.00214566f $X=5.67 $Y=0.655
+ $X2=0 $Y2=0
cc_813 N_A_1092_96#_c_952_n N_A_622_98#_c_1222_n 0.00153106f $X=5.955 $Y=2.37
+ $X2=0 $Y2=0
cc_814 N_A_1092_96#_c_952_n N_A_622_98#_c_1224_n 0.0100254f $X=5.955 $Y=2.37
+ $X2=0 $Y2=0
cc_815 N_A_1092_96#_c_953_n N_A_622_98#_c_1224_n 0.00982558f $X=6.04 $Y=2.205
+ $X2=0 $Y2=0
cc_816 N_A_1092_96#_c_951_n N_A_622_98#_c_1225_n 0.00882199f $X=7.825 $Y=1.82
+ $X2=0 $Y2=0
cc_817 N_A_1092_96#_c_953_n N_A_877_98#_c_1440_n 0.00117754f $X=6.04 $Y=2.205
+ $X2=0 $Y2=0
cc_818 N_A_1092_96#_c_952_n N_A_877_98#_c_1441_n 0.00412455f $X=5.955 $Y=2.37
+ $X2=0 $Y2=0
cc_819 N_A_1092_96#_c_941_n N_A_877_98#_c_1441_n 0.00336206f $X=6.04 $Y=1.655
+ $X2=0 $Y2=0
cc_820 N_A_1092_96#_c_948_n N_A_877_98#_c_1441_n 7.30194e-19 $X=5.67 $Y=0.655
+ $X2=0 $Y2=0
cc_821 N_A_1092_96#_c_941_n N_A_877_98#_M1030_g 0.0104792f $X=6.04 $Y=1.655
+ $X2=0 $Y2=0
cc_822 N_A_1092_96#_c_948_n N_A_877_98#_M1030_g 0.0183636f $X=5.67 $Y=0.655
+ $X2=0 $Y2=0
cc_823 N_A_1092_96#_c_948_n N_A_877_98#_c_1443_n 0.00139736f $X=5.67 $Y=0.655
+ $X2=0 $Y2=0
cc_824 N_A_1092_96#_c_949_n N_A_877_98#_c_1443_n 0.00880557f $X=7.75 $Y=1.255
+ $X2=0 $Y2=0
cc_825 N_A_1092_96#_c_952_n N_VPWR_c_2016_n 0.00668433f $X=5.955 $Y=2.37 $X2=0
+ $Y2=0
cc_826 N_A_1092_96#_c_953_n N_VPWR_c_2016_n 0.00283451f $X=6.04 $Y=2.205 $X2=0
+ $Y2=0
cc_827 N_A_1092_96#_c_942_n N_VPWR_c_2016_n 0.0191398f $X=6.705 $Y=1.74 $X2=0
+ $Y2=0
cc_828 N_A_1092_96#_c_952_n N_VPWR_c_2012_n 0.0187254f $X=5.955 $Y=2.37 $X2=0
+ $Y2=0
cc_829 N_A_1092_96#_c_953_n N_A_197_119#_c_2211_n 0.00470927f $X=6.04 $Y=2.205
+ $X2=0 $Y2=0
cc_830 N_A_1092_96#_c_941_n N_A_197_119#_c_2200_n 0.00391399f $X=6.04 $Y=1.655
+ $X2=0 $Y2=0
cc_831 N_A_1092_96#_c_941_n N_A_197_119#_c_2201_n 0.0136046f $X=6.04 $Y=1.655
+ $X2=0 $Y2=0
cc_832 N_A_1092_96#_c_948_n N_A_197_119#_c_2201_n 0.0218829f $X=5.67 $Y=0.655
+ $X2=0 $Y2=0
cc_833 N_A_1092_96#_c_952_n N_A_197_119#_c_2212_n 0.0168758f $X=5.955 $Y=2.37
+ $X2=0 $Y2=0
cc_834 N_A_1092_96#_c_953_n N_A_197_119#_c_2212_n 0.0141453f $X=6.04 $Y=2.205
+ $X2=0 $Y2=0
cc_835 N_A_1092_96#_c_941_n N_A_197_119#_c_2203_n 0.032757f $X=6.04 $Y=1.655
+ $X2=0 $Y2=0
cc_836 N_A_1092_96#_c_953_n N_A_197_119#_c_2203_n 0.00293665f $X=6.04 $Y=2.205
+ $X2=0 $Y2=0
cc_837 N_A_1092_96#_c_955_n N_A_197_119#_c_2203_n 0.0143579f $X=6.04 $Y=1.74
+ $X2=0 $Y2=0
cc_838 N_A_1092_96#_c_948_n N_A_197_119#_c_2206_n 0.0154541f $X=5.67 $Y=0.655
+ $X2=0 $Y2=0
cc_839 N_A_1092_96#_c_945_n N_VGND_M1046_d 0.00309396f $X=6.875 $Y=1.155 $X2=0
+ $Y2=0
cc_840 N_A_1092_96#_c_948_n N_VGND_c_2433_n 0.00286827f $X=5.67 $Y=0.655 $X2=0
+ $Y2=0
cc_841 N_A_1092_96#_c_948_n N_VGND_c_2440_n 0.0139308f $X=5.67 $Y=0.655 $X2=0
+ $Y2=0
cc_842 N_A_1092_96#_c_948_n N_VGND_c_2451_n 0.0179751f $X=5.67 $Y=0.655 $X2=0
+ $Y2=0
cc_843 N_A_1092_96#_c_941_n A_1192_96# 0.00157575f $X=6.04 $Y=1.655 $X2=-0.19
+ $Y2=-0.245
cc_844 N_A_1092_96#_c_948_n A_1192_96# 0.00348804f $X=5.67 $Y=0.655 $X2=-0.19
+ $Y2=-0.245
cc_845 N_A_1092_96#_c_944_n N_A_1418_125#_M1022_d 0.00592612f $X=7.585 $Y=1.155
+ $X2=-0.19 $Y2=-0.245
cc_846 N_A_1092_96#_c_949_n N_A_1418_125#_c_2601_n 0.00278649f $X=7.75 $Y=1.255
+ $X2=0 $Y2=0
cc_847 N_A_1092_96#_c_949_n N_A_1418_125#_c_2603_n 0.00399463f $X=7.75 $Y=1.255
+ $X2=0 $Y2=0
cc_848 N_A_1625_93#_c_1074_n N_A_622_98#_c_1225_n 0.0104018f $X=8.245 $Y=1.82
+ $X2=0 $Y2=0
cc_849 N_A_1625_93#_c_1065_n N_A_622_98#_c_1211_n 0.00851227f $X=12.575 $Y=1.295
+ $X2=0 $Y2=0
cc_850 N_A_1625_93#_c_1065_n N_A_622_98#_c_1212_n 0.00605232f $X=12.575 $Y=1.295
+ $X2=0 $Y2=0
cc_851 N_A_1625_93#_c_1065_n N_A_622_98#_c_1215_n 0.0146673f $X=12.575 $Y=1.295
+ $X2=0 $Y2=0
cc_852 N_A_1625_93#_c_1065_n N_A_622_98#_c_1216_n 0.0150214f $X=12.575 $Y=1.295
+ $X2=0 $Y2=0
cc_853 N_A_1625_93#_c_1072_n N_A_877_98#_c_1443_n 0.00880557f $X=8.29 $Y=1.255
+ $X2=0 $Y2=0
cc_854 N_A_1625_93#_c_1065_n N_A_877_98#_c_1446_n 0.0121899f $X=12.575 $Y=1.295
+ $X2=0 $Y2=0
cc_855 N_A_1625_93#_c_1065_n N_A_2037_442#_M1047_g 0.00283763f $X=12.575
+ $Y=1.295 $X2=0 $Y2=0
cc_856 N_A_1625_93#_c_1069_n N_A_2037_442#_c_1592_n 2.27331e-19 $X=12.72
+ $Y=1.295 $X2=0 $Y2=0
cc_857 N_A_1625_93#_c_1060_n N_A_2037_442#_c_1598_n 0.00547592f $X=12.235
+ $Y=1.795 $X2=0 $Y2=0
cc_858 N_A_1625_93#_c_1076_n N_A_2037_442#_c_1598_n 0.00522828f $X=12.235
+ $Y=1.885 $X2=0 $Y2=0
cc_859 N_A_1625_93#_c_1061_n N_A_2037_442#_c_1598_n 0.00611109f $X=12.25 $Y=1.22
+ $X2=0 $Y2=0
cc_860 N_A_1625_93#_c_1062_n N_A_2037_442#_c_1598_n 0.00863047f $X=12.145 $Y=1.4
+ $X2=0 $Y2=0
cc_861 N_A_1625_93#_c_1063_n N_A_2037_442#_c_1598_n 0.00546445f $X=12.81 $Y=1.18
+ $X2=0 $Y2=0
cc_862 N_A_1625_93#_c_1065_n N_A_2037_442#_c_1598_n 0.0228634f $X=12.575
+ $Y=1.295 $X2=0 $Y2=0
cc_863 N_A_1625_93#_c_1068_n N_A_2037_442#_c_1598_n 4.47366e-19 $X=12.72
+ $Y=1.295 $X2=0 $Y2=0
cc_864 N_A_1625_93#_c_1069_n N_A_2037_442#_c_1598_n 0.0386818f $X=12.72 $Y=1.295
+ $X2=0 $Y2=0
cc_865 N_A_1625_93#_M1028_s N_A_2037_442#_c_1610_n 0.0117736f $X=12.86 $Y=1.74
+ $X2=0 $Y2=0
cc_866 N_A_1625_93#_c_1076_n N_A_2037_442#_c_1610_n 0.0134212f $X=12.235
+ $Y=1.885 $X2=0 $Y2=0
cc_867 N_A_1625_93#_c_1069_n N_A_2037_442#_c_1610_n 0.0415715f $X=12.72 $Y=1.295
+ $X2=0 $Y2=0
cc_868 N_A_1625_93#_c_1070_n N_A_2037_442#_c_1610_n 0.003784f $X=12.61 $Y=1.385
+ $X2=0 $Y2=0
cc_869 N_A_1625_93#_c_1076_n N_A_2037_442#_c_1626_n 0.0164192f $X=12.235
+ $Y=1.885 $X2=0 $Y2=0
cc_870 N_A_1625_93#_c_1065_n N_A_2037_442#_c_1626_n 0.00804224f $X=12.575
+ $Y=1.295 $X2=0 $Y2=0
cc_871 N_A_1625_93#_c_1069_n N_A_2037_442#_c_1599_n 0.0157594f $X=12.72 $Y=1.295
+ $X2=0 $Y2=0
cc_872 N_A_1625_93#_c_1076_n N_A_2037_442#_c_1614_n 0.00137387f $X=12.235
+ $Y=1.885 $X2=0 $Y2=0
cc_873 N_A_1625_93#_c_1061_n N_A_2037_442#_c_1655_n 0.00571558f $X=12.25 $Y=1.22
+ $X2=0 $Y2=0
cc_874 N_A_1625_93#_c_1065_n N_A_2037_442#_c_1655_n 0.00797186f $X=12.575
+ $Y=1.295 $X2=0 $Y2=0
cc_875 N_A_1625_93#_c_1061_n N_A_1878_420#_c_1772_n 0.020929f $X=12.25 $Y=1.22
+ $X2=0 $Y2=0
cc_876 N_A_1625_93#_c_1060_n N_A_1878_420#_c_1773_n 0.00986205f $X=12.235
+ $Y=1.795 $X2=0 $Y2=0
cc_877 N_A_1625_93#_c_1062_n N_A_1878_420#_c_1773_n 0.0185668f $X=12.145 $Y=1.4
+ $X2=0 $Y2=0
cc_878 N_A_1625_93#_c_1065_n N_A_1878_420#_c_1773_n 0.0023f $X=12.575 $Y=1.295
+ $X2=0 $Y2=0
cc_879 N_A_1625_93#_c_1076_n N_A_1878_420#_c_1774_n 0.00986205f $X=12.235
+ $Y=1.885 $X2=0 $Y2=0
cc_880 N_A_1625_93#_c_1076_n N_A_1878_420#_c_1783_n 0.0624017f $X=12.235
+ $Y=1.885 $X2=0 $Y2=0
cc_881 N_A_1625_93#_c_1065_n N_A_1878_420#_c_1775_n 0.0187205f $X=12.575
+ $Y=1.295 $X2=0 $Y2=0
cc_882 N_A_1625_93#_c_1065_n N_A_1878_420#_c_1776_n 0.0270033f $X=12.575
+ $Y=1.295 $X2=0 $Y2=0
cc_883 N_A_1625_93#_c_1065_n N_A_1878_420#_c_1777_n 0.0291312f $X=12.575
+ $Y=1.295 $X2=0 $Y2=0
cc_884 N_A_1625_93#_c_1065_n N_A_1878_420#_c_1787_n 0.00122709f $X=12.575
+ $Y=1.295 $X2=0 $Y2=0
cc_885 N_A_1625_93#_c_1065_n N_A_1878_420#_c_1779_n 0.0107145f $X=12.575
+ $Y=1.295 $X2=0 $Y2=0
cc_886 N_A_1625_93#_c_1065_n N_A_1878_420#_c_1780_n 0.0159733f $X=12.575
+ $Y=1.295 $X2=0 $Y2=0
cc_887 N_A_1625_93#_c_1062_n N_A_1878_420#_c_1781_n 3.72296e-19 $X=12.145 $Y=1.4
+ $X2=0 $Y2=0
cc_888 N_A_1625_93#_c_1065_n N_A_1878_420#_c_1781_n 0.0211316f $X=12.575
+ $Y=1.295 $X2=0 $Y2=0
cc_889 N_A_1625_93#_c_1064_n N_RESET_B_c_1889_n 0.00113718f $X=13.03 $Y=0.84
+ $X2=-0.19 $Y2=-0.245
cc_890 N_A_1625_93#_c_1069_n N_RESET_B_c_1889_n 0.0123564f $X=12.72 $Y=1.295
+ $X2=-0.19 $Y2=-0.245
cc_891 N_A_1625_93#_c_1070_n N_RESET_B_c_1889_n 0.0149046f $X=12.61 $Y=1.385
+ $X2=-0.19 $Y2=-0.245
cc_892 N_A_1625_93#_c_1063_n N_RESET_B_c_1890_n 0.00480829f $X=12.81 $Y=1.18
+ $X2=0 $Y2=0
cc_893 N_A_1625_93#_c_1064_n N_RESET_B_c_1890_n 4.28014e-19 $X=13.03 $Y=0.84
+ $X2=0 $Y2=0
cc_894 N_A_1625_93#_c_1069_n N_RESET_B_c_1890_n 2.32911e-19 $X=12.72 $Y=1.295
+ $X2=0 $Y2=0
cc_895 N_A_1625_93#_c_1064_n RESET_B 0.00398773f $X=13.03 $Y=0.84 $X2=0 $Y2=0
cc_896 N_A_1625_93#_c_1068_n RESET_B 0.00154479f $X=12.72 $Y=1.295 $X2=0 $Y2=0
cc_897 N_A_1625_93#_c_1069_n RESET_B 0.0355209f $X=12.72 $Y=1.295 $X2=0 $Y2=0
cc_898 N_A_1625_93#_c_1070_n RESET_B 3.25754e-19 $X=12.61 $Y=1.385 $X2=0 $Y2=0
cc_899 N_A_1625_93#_c_1074_n N_VPWR_c_2017_n 0.00531163f $X=8.245 $Y=1.82 $X2=0
+ $Y2=0
cc_900 N_A_1625_93#_c_1076_n N_VPWR_c_2018_n 0.0155839f $X=12.235 $Y=1.885 $X2=0
+ $Y2=0
cc_901 N_A_1625_93#_c_1076_n N_VPWR_c_2023_n 0.00413917f $X=12.235 $Y=1.885
+ $X2=0 $Y2=0
cc_902 N_A_1625_93#_c_1074_n N_VPWR_c_2012_n 9.14192e-19 $X=8.245 $Y=1.82 $X2=0
+ $Y2=0
cc_903 N_A_1625_93#_c_1076_n N_VPWR_c_2012_n 0.00817239f $X=12.235 $Y=1.885
+ $X2=0 $Y2=0
cc_904 N_A_1625_93#_c_1065_n N_VGND_c_2434_n 0.0115947f $X=12.575 $Y=1.295 $X2=0
+ $Y2=0
cc_905 N_A_1625_93#_c_1065_n N_VGND_c_2435_n 0.00191454f $X=12.575 $Y=1.295
+ $X2=0 $Y2=0
cc_906 N_A_1625_93#_c_1064_n N_VGND_c_2436_n 0.012384f $X=13.03 $Y=0.84 $X2=0
+ $Y2=0
cc_907 N_A_1625_93#_c_1061_n N_VGND_c_2446_n 0.00278271f $X=12.25 $Y=1.22 $X2=0
+ $Y2=0
cc_908 N_A_1625_93#_c_1064_n N_VGND_c_2446_n 0.0069583f $X=13.03 $Y=0.84 $X2=0
+ $Y2=0
cc_909 N_A_1625_93#_c_1061_n N_VGND_c_2451_n 0.00359456f $X=12.25 $Y=1.22 $X2=0
+ $Y2=0
cc_910 N_A_1625_93#_c_1064_n N_VGND_c_2451_n 0.0111617f $X=13.03 $Y=0.84 $X2=0
+ $Y2=0
cc_911 N_A_1625_93#_c_1072_n N_A_1418_125#_c_2602_n 0.00339325f $X=8.29 $Y=1.255
+ $X2=0 $Y2=0
cc_912 N_A_1625_93#_c_1072_n N_A_1418_125#_c_2603_n 0.00398082f $X=8.29 $Y=1.255
+ $X2=0 $Y2=0
cc_913 N_A_1625_93#_c_1061_n N_A_2271_74#_c_2628_n 9.0523e-19 $X=12.25 $Y=1.22
+ $X2=0 $Y2=0
cc_914 N_A_1625_93#_c_1065_n N_A_2271_74#_c_2628_n 0.00249118f $X=12.575
+ $Y=1.295 $X2=0 $Y2=0
cc_915 N_A_1625_93#_c_1061_n N_A_2271_74#_c_2626_n 0.0131811f $X=12.25 $Y=1.22
+ $X2=0 $Y2=0
cc_916 N_A_1625_93#_c_1064_n N_A_2271_74#_c_2633_n 0.0268324f $X=13.03 $Y=0.84
+ $X2=0 $Y2=0
cc_917 N_A_1625_93#_c_1065_n N_A_2271_74#_c_2633_n 0.00359698f $X=12.575
+ $Y=1.295 $X2=0 $Y2=0
cc_918 N_A_1625_93#_c_1069_n N_A_2271_74#_c_2633_n 0.00901771f $X=12.72 $Y=1.295
+ $X2=0 $Y2=0
cc_919 N_A_1625_93#_c_1070_n N_A_2271_74#_c_2633_n 0.00328544f $X=12.61 $Y=1.385
+ $X2=0 $Y2=0
cc_920 N_A_622_98#_c_1200_n N_A_877_98#_c_1440_n 0.0185464f $X=4.875 $Y=3.075
+ $X2=0 $Y2=0
cc_921 N_A_622_98#_c_1220_n N_A_877_98#_c_1440_n 0.0103487f $X=5.94 $Y=3.15
+ $X2=0 $Y2=0
cc_922 N_A_622_98#_c_1203_n N_A_877_98#_c_1440_n 0.00523803f $X=5.385 $Y=0.405
+ $X2=0 $Y2=0
cc_923 N_A_622_98#_c_1222_n N_A_877_98#_c_1440_n 0.00938554f $X=6.03 $Y=2.68
+ $X2=0 $Y2=0
cc_924 N_A_622_98#_c_1224_n N_A_877_98#_c_1440_n 0.0106005f $X=6.03 $Y=2.59
+ $X2=0 $Y2=0
cc_925 N_A_622_98#_c_1205_n N_A_877_98#_c_1440_n 0.0214265f $X=4.875 $Y=1.415
+ $X2=0 $Y2=0
cc_926 N_A_622_98#_c_1201_n N_A_877_98#_M1030_g 0.020088f $X=5.31 $Y=0.33 $X2=0
+ $Y2=0
cc_927 N_A_622_98#_c_1210_n N_A_877_98#_c_1443_n 0.0032544f $X=9.615 $Y=0.34
+ $X2=0 $Y2=0
cc_928 N_A_622_98#_c_1217_n N_A_877_98#_c_1443_n 0.00974585f $X=10.32 $Y=0.9
+ $X2=0 $Y2=0
cc_929 N_A_622_98#_c_1209_n N_A_877_98#_M1001_g 0.0124359f $X=10.155 $Y=0.34
+ $X2=0 $Y2=0
cc_930 N_A_622_98#_c_1210_n N_A_877_98#_M1001_g 0.0030674f $X=9.615 $Y=0.34
+ $X2=0 $Y2=0
cc_931 N_A_622_98#_c_1211_n N_A_877_98#_M1001_g 8.16681e-19 $X=10.32 $Y=1.065
+ $X2=0 $Y2=0
cc_932 N_A_622_98#_c_1212_n N_A_877_98#_M1001_g 0.00974585f $X=10.32 $Y=1.065
+ $X2=0 $Y2=0
cc_933 N_A_622_98#_c_1215_n N_A_877_98#_M1001_g 0.0136728f $X=9.435 $Y=1.335
+ $X2=0 $Y2=0
cc_934 N_A_622_98#_c_1225_n N_A_877_98#_c_1453_n 0.00167456f $X=9.225 $Y=3.15
+ $X2=0 $Y2=0
cc_935 N_A_622_98#_M1008_g N_A_877_98#_c_1453_n 0.0161947f $X=9.315 $Y=2.52
+ $X2=0 $Y2=0
cc_936 N_A_622_98#_c_1212_n N_A_877_98#_c_1446_n 6.52121e-19 $X=10.32 $Y=1.065
+ $X2=0 $Y2=0
cc_937 N_A_622_98#_c_1215_n N_A_877_98#_c_1446_n 0.00161516f $X=9.435 $Y=1.335
+ $X2=0 $Y2=0
cc_938 N_A_622_98#_c_1216_n N_A_877_98#_c_1446_n 6.13228e-19 $X=9.435 $Y=1.505
+ $X2=0 $Y2=0
cc_939 N_A_622_98#_c_1204_n N_A_877_98#_c_1447_n 0.022985f $X=9.315 $Y=2.025
+ $X2=0 $Y2=0
cc_940 N_A_622_98#_M1008_g N_A_877_98#_c_1447_n 0.00296877f $X=9.315 $Y=2.52
+ $X2=0 $Y2=0
cc_941 N_A_622_98#_c_1208_n N_A_877_98#_c_1447_n 0.00114988f $X=9.42 $Y=1.775
+ $X2=0 $Y2=0
cc_942 N_A_622_98#_c_1216_n N_A_877_98#_c_1447_n 9.86445e-19 $X=9.435 $Y=1.505
+ $X2=0 $Y2=0
cc_943 N_A_622_98#_c_1196_n N_A_877_98#_c_1448_n 0.00837336f $X=4.31 $Y=1.34
+ $X2=0 $Y2=0
cc_944 N_A_622_98#_c_1197_n N_A_877_98#_c_1448_n 0.00548201f $X=4.355 $Y=1.765
+ $X2=0 $Y2=0
cc_945 N_A_622_98#_c_1199_n N_A_877_98#_c_1448_n 0.00731087f $X=4.875 $Y=1.34
+ $X2=0 $Y2=0
cc_946 N_A_622_98#_c_1214_n N_A_877_98#_c_1448_n 0.0129723f $X=4.4 $Y=1.505
+ $X2=0 $Y2=0
cc_947 N_A_622_98#_c_1197_n N_A_877_98#_c_1455_n 0.0106367f $X=4.355 $Y=1.765
+ $X2=0 $Y2=0
cc_948 N_A_622_98#_c_1200_n N_A_877_98#_c_1455_n 0.0341092f $X=4.875 $Y=3.075
+ $X2=0 $Y2=0
cc_949 N_A_622_98#_c_1196_n N_A_877_98#_c_1449_n 0.00278843f $X=4.31 $Y=1.34
+ $X2=0 $Y2=0
cc_950 N_A_622_98#_c_1198_n N_A_877_98#_c_1449_n 4.56256e-19 $X=4.8 $Y=1.415
+ $X2=0 $Y2=0
cc_951 N_A_622_98#_c_1199_n N_A_877_98#_c_1449_n 0.00849541f $X=4.875 $Y=1.34
+ $X2=0 $Y2=0
cc_952 N_A_622_98#_c_1205_n N_A_877_98#_c_1449_n 0.00112453f $X=4.875 $Y=1.415
+ $X2=0 $Y2=0
cc_953 N_A_622_98#_c_1214_n N_A_877_98#_c_1449_n 0.00174498f $X=4.4 $Y=1.505
+ $X2=0 $Y2=0
cc_954 N_A_622_98#_c_1200_n N_A_877_98#_c_1450_n 0.0047606f $X=4.875 $Y=3.075
+ $X2=0 $Y2=0
cc_955 N_A_622_98#_c_1205_n N_A_877_98#_c_1450_n 0.00281698f $X=4.875 $Y=1.415
+ $X2=0 $Y2=0
cc_956 N_A_622_98#_c_1197_n N_A_877_98#_c_1457_n 0.00587461f $X=4.355 $Y=1.765
+ $X2=0 $Y2=0
cc_957 N_A_622_98#_c_1198_n N_A_877_98#_c_1457_n 0.00373956f $X=4.8 $Y=1.415
+ $X2=0 $Y2=0
cc_958 N_A_622_98#_c_1200_n N_A_877_98#_c_1457_n 0.00777625f $X=4.875 $Y=3.075
+ $X2=0 $Y2=0
cc_959 N_A_622_98#_c_1232_n N_A_877_98#_c_1457_n 0.0048272f $X=3.68 $Y=2.815
+ $X2=0 $Y2=0
cc_960 N_A_622_98#_c_1214_n N_A_877_98#_c_1457_n 0.00966564f $X=4.4 $Y=1.505
+ $X2=0 $Y2=0
cc_961 N_A_622_98#_c_1197_n N_A_877_98#_c_1458_n 0.00111158f $X=4.355 $Y=1.765
+ $X2=0 $Y2=0
cc_962 N_A_622_98#_c_1200_n N_A_877_98#_c_1458_n 0.00456881f $X=4.875 $Y=3.075
+ $X2=0 $Y2=0
cc_963 N_A_622_98#_c_1233_n N_A_877_98#_c_1458_n 0.0051601f $X=4.16 $Y=1.84
+ $X2=0 $Y2=0
cc_964 N_A_622_98#_c_1197_n N_A_877_98#_c_1451_n 9.29283e-19 $X=4.355 $Y=1.765
+ $X2=0 $Y2=0
cc_965 N_A_622_98#_c_1198_n N_A_877_98#_c_1451_n 0.00415752f $X=4.8 $Y=1.415
+ $X2=0 $Y2=0
cc_966 N_A_622_98#_c_1200_n N_A_877_98#_c_1451_n 0.00288841f $X=4.875 $Y=3.075
+ $X2=0 $Y2=0
cc_967 N_A_622_98#_c_1205_n N_A_877_98#_c_1451_n 0.00123591f $X=4.875 $Y=1.415
+ $X2=0 $Y2=0
cc_968 N_A_622_98#_c_1233_n N_A_877_98#_c_1451_n 0.0010093f $X=4.16 $Y=1.84
+ $X2=0 $Y2=0
cc_969 N_A_622_98#_c_1214_n N_A_877_98#_c_1451_n 0.0260033f $X=4.4 $Y=1.505
+ $X2=0 $Y2=0
cc_970 N_A_622_98#_c_1209_n N_A_2037_442#_M1047_g 0.00176953f $X=10.155 $Y=0.34
+ $X2=0 $Y2=0
cc_971 N_A_622_98#_c_1211_n N_A_2037_442#_M1047_g 0.00596986f $X=10.32 $Y=1.065
+ $X2=0 $Y2=0
cc_972 N_A_622_98#_c_1212_n N_A_2037_442#_M1047_g 0.0207114f $X=10.32 $Y=1.065
+ $X2=0 $Y2=0
cc_973 N_A_622_98#_c_1217_n N_A_2037_442#_M1047_g 0.0170701f $X=10.32 $Y=0.9
+ $X2=0 $Y2=0
cc_974 N_A_622_98#_c_1209_n N_A_1878_420#_M1001_d 0.00529413f $X=10.155 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_975 N_A_622_98#_c_1209_n N_A_1878_420#_c_1775_n 0.0140001f $X=10.155 $Y=0.34
+ $X2=0 $Y2=0
cc_976 N_A_622_98#_c_1211_n N_A_1878_420#_c_1775_n 0.0437292f $X=10.32 $Y=1.065
+ $X2=0 $Y2=0
cc_977 N_A_622_98#_c_1215_n N_A_1878_420#_c_1775_n 0.0323996f $X=9.435 $Y=1.335
+ $X2=0 $Y2=0
cc_978 N_A_622_98#_c_1217_n N_A_1878_420#_c_1775_n 0.0053389f $X=10.32 $Y=0.9
+ $X2=0 $Y2=0
cc_979 N_A_622_98#_c_1211_n N_A_1878_420#_c_1776_n 0.0223986f $X=10.32 $Y=1.065
+ $X2=0 $Y2=0
cc_980 N_A_622_98#_c_1212_n N_A_1878_420#_c_1776_n 0.00626155f $X=10.32 $Y=1.065
+ $X2=0 $Y2=0
cc_981 N_A_622_98#_c_1204_n N_A_1878_420#_c_1784_n 0.00127627f $X=9.315 $Y=2.025
+ $X2=0 $Y2=0
cc_982 N_A_622_98#_M1008_g N_A_1878_420#_c_1784_n 0.00986345f $X=9.315 $Y=2.52
+ $X2=0 $Y2=0
cc_983 N_A_622_98#_c_1208_n N_A_1878_420#_c_1784_n 0.0153945f $X=9.42 $Y=1.775
+ $X2=0 $Y2=0
cc_984 N_A_622_98#_c_1216_n N_A_1878_420#_c_1784_n 0.00105518f $X=9.435 $Y=1.505
+ $X2=0 $Y2=0
cc_985 N_A_622_98#_c_1204_n N_A_1878_420#_c_1785_n 0.00150093f $X=9.315 $Y=2.025
+ $X2=0 $Y2=0
cc_986 N_A_622_98#_M1008_g N_A_1878_420#_c_1785_n 0.00142265f $X=9.315 $Y=2.52
+ $X2=0 $Y2=0
cc_987 N_A_622_98#_c_1204_n N_A_1878_420#_c_1778_n 3.46152e-19 $X=9.315 $Y=2.025
+ $X2=0 $Y2=0
cc_988 N_A_622_98#_c_1208_n N_A_1878_420#_c_1778_n 0.0106213f $X=9.42 $Y=1.775
+ $X2=0 $Y2=0
cc_989 N_A_622_98#_c_1204_n N_A_1878_420#_c_1787_n 0.00142581f $X=9.315 $Y=2.025
+ $X2=0 $Y2=0
cc_990 N_A_622_98#_c_1208_n N_A_1878_420#_c_1787_n 0.0200389f $X=9.42 $Y=1.775
+ $X2=0 $Y2=0
cc_991 N_A_622_98#_c_1208_n N_A_1878_420#_c_1779_n 0.00114554f $X=9.42 $Y=1.775
+ $X2=0 $Y2=0
cc_992 N_A_622_98#_c_1216_n N_A_1878_420#_c_1779_n 0.013405f $X=9.435 $Y=1.505
+ $X2=0 $Y2=0
cc_993 N_A_622_98#_c_1212_n N_A_1878_420#_c_1780_n 3.59235e-19 $X=10.32 $Y=1.065
+ $X2=0 $Y2=0
cc_994 N_A_622_98#_c_1261_n N_VPWR_M1040_d 0.00448307f $X=4.075 $Y=1.925 $X2=0
+ $Y2=0
cc_995 N_A_622_98#_c_1197_n N_VPWR_c_2015_n 0.00556363f $X=4.355 $Y=1.765 $X2=0
+ $Y2=0
cc_996 N_A_622_98#_c_1200_n N_VPWR_c_2015_n 0.00225512f $X=4.875 $Y=3.075 $X2=0
+ $Y2=0
cc_997 N_A_622_98#_c_1232_n N_VPWR_c_2015_n 0.0521368f $X=3.68 $Y=2.815 $X2=0
+ $Y2=0
cc_998 N_A_622_98#_c_1261_n N_VPWR_c_2015_n 0.0142476f $X=4.075 $Y=1.925 $X2=0
+ $Y2=0
cc_999 N_A_622_98#_c_1222_n N_VPWR_c_2016_n 0.0118751f $X=6.03 $Y=2.68 $X2=0
+ $Y2=0
cc_1000 N_A_622_98#_c_1225_n N_VPWR_c_2016_n 0.0261591f $X=9.225 $Y=3.15 $X2=0
+ $Y2=0
cc_1001 N_A_622_98#_c_1225_n N_VPWR_c_2017_n 0.0279235f $X=9.225 $Y=3.15 $X2=0
+ $Y2=0
cc_1002 N_A_622_98#_M1008_g N_VPWR_c_2017_n 4.33975e-19 $X=9.315 $Y=2.52 $X2=0
+ $Y2=0
cc_1003 N_A_622_98#_c_1197_n N_VPWR_c_2021_n 0.00445602f $X=4.355 $Y=1.765 $X2=0
+ $Y2=0
cc_1004 N_A_622_98#_c_1221_n N_VPWR_c_2021_n 0.0600202f $X=4.95 $Y=3.15 $X2=0
+ $Y2=0
cc_1005 N_A_622_98#_c_1232_n N_VPWR_c_2029_n 0.0145938f $X=3.68 $Y=2.815 $X2=0
+ $Y2=0
cc_1006 N_A_622_98#_c_1225_n N_VPWR_c_2030_n 0.0337061f $X=9.225 $Y=3.15 $X2=0
+ $Y2=0
cc_1007 N_A_622_98#_c_1197_n N_VPWR_c_2012_n 0.00858307f $X=4.355 $Y=1.765 $X2=0
+ $Y2=0
cc_1008 N_A_622_98#_c_1220_n N_VPWR_c_2012_n 0.0330622f $X=5.94 $Y=3.15 $X2=0
+ $Y2=0
cc_1009 N_A_622_98#_c_1221_n N_VPWR_c_2012_n 0.00774408f $X=4.95 $Y=3.15 $X2=0
+ $Y2=0
cc_1010 N_A_622_98#_c_1225_n N_VPWR_c_2012_n 0.0841862f $X=9.225 $Y=3.15 $X2=0
+ $Y2=0
cc_1011 N_A_622_98#_c_1228_n N_VPWR_c_2012_n 0.00559601f $X=6.03 $Y=3.15 $X2=0
+ $Y2=0
cc_1012 N_A_622_98#_c_1232_n N_VPWR_c_2012_n 0.0120466f $X=3.68 $Y=2.815 $X2=0
+ $Y2=0
cc_1013 N_A_622_98#_c_1225_n N_VPWR_c_2038_n 0.0176167f $X=9.225 $Y=3.15 $X2=0
+ $Y2=0
cc_1014 N_A_622_98#_c_1206_n N_A_197_119#_c_2197_n 0.0189779f $X=3.255 $Y=0.8
+ $X2=0 $Y2=0
cc_1015 N_A_622_98#_c_1196_n N_A_197_119#_c_2199_n 0.00265744f $X=4.31 $Y=1.34
+ $X2=0 $Y2=0
cc_1016 N_A_622_98#_c_1200_n N_A_197_119#_c_2211_n 0.00589152f $X=4.875 $Y=3.075
+ $X2=0 $Y2=0
cc_1017 N_A_622_98#_c_1220_n N_A_197_119#_c_2211_n 0.00641825f $X=5.94 $Y=3.15
+ $X2=0 $Y2=0
cc_1018 N_A_622_98#_c_1222_n N_A_197_119#_c_2211_n 7.62388e-19 $X=6.03 $Y=2.68
+ $X2=0 $Y2=0
cc_1019 N_A_622_98#_c_1224_n N_A_197_119#_c_2211_n 7.5081e-19 $X=6.03 $Y=2.59
+ $X2=0 $Y2=0
cc_1020 N_A_622_98#_c_1199_n N_A_197_119#_c_2200_n 0.00362479f $X=4.875 $Y=1.34
+ $X2=0 $Y2=0
cc_1021 N_A_622_98#_c_1203_n N_A_197_119#_c_2200_n 0.00531745f $X=5.385 $Y=0.405
+ $X2=0 $Y2=0
cc_1022 N_A_622_98#_c_1203_n N_A_197_119#_c_2201_n 0.00664391f $X=5.385 $Y=0.405
+ $X2=0 $Y2=0
cc_1023 N_A_622_98#_c_1199_n N_A_197_119#_c_2202_n 0.00335272f $X=4.875 $Y=1.34
+ $X2=0 $Y2=0
cc_1024 N_A_622_98#_c_1203_n N_A_197_119#_c_2202_n 2.70037e-19 $X=5.385 $Y=0.405
+ $X2=0 $Y2=0
cc_1025 N_A_622_98#_c_1224_n N_A_197_119#_c_2212_n 5.34654e-19 $X=6.03 $Y=2.59
+ $X2=0 $Y2=0
cc_1026 N_A_622_98#_c_1200_n N_A_197_119#_c_2213_n 0.00145939f $X=4.875 $Y=3.075
+ $X2=0 $Y2=0
cc_1027 N_A_622_98#_c_1199_n N_A_197_119#_c_2203_n 0.00358179f $X=4.875 $Y=1.34
+ $X2=0 $Y2=0
cc_1028 N_A_622_98#_c_1196_n N_A_197_119#_c_2205_n 0.0151175f $X=4.31 $Y=1.34
+ $X2=0 $Y2=0
cc_1029 N_A_622_98#_c_1199_n N_A_197_119#_c_2205_n 0.0134424f $X=4.875 $Y=1.34
+ $X2=0 $Y2=0
cc_1030 N_A_622_98#_c_1214_n N_A_197_119#_c_2205_n 0.00841151f $X=4.4 $Y=1.505
+ $X2=0 $Y2=0
cc_1031 N_A_622_98#_c_1196_n N_A_197_119#_c_2206_n 8.60511e-19 $X=4.31 $Y=1.34
+ $X2=0 $Y2=0
cc_1032 N_A_622_98#_c_1199_n N_A_197_119#_c_2206_n 0.00465249f $X=4.875 $Y=1.34
+ $X2=0 $Y2=0
cc_1033 N_A_622_98#_c_1201_n N_A_197_119#_c_2206_n 0.00464948f $X=5.31 $Y=0.33
+ $X2=0 $Y2=0
cc_1034 N_A_622_98#_c_1203_n N_A_197_119#_c_2206_n 0.00457f $X=5.385 $Y=0.405
+ $X2=0 $Y2=0
cc_1035 N_A_622_98#_c_1196_n N_VGND_c_2432_n 0.0041157f $X=4.31 $Y=1.34 $X2=0
+ $Y2=0
cc_1036 N_A_622_98#_c_1202_n N_VGND_c_2432_n 0.00328037f $X=4.95 $Y=0.33 $X2=0
+ $Y2=0
cc_1037 N_A_622_98#_c_1210_n N_VGND_c_2434_n 0.0147452f $X=9.615 $Y=0.34 $X2=0
+ $Y2=0
cc_1038 N_A_622_98#_c_1215_n N_VGND_c_2434_n 0.0289547f $X=9.435 $Y=1.335 $X2=0
+ $Y2=0
cc_1039 N_A_622_98#_c_1216_n N_VGND_c_2434_n 6.49245e-19 $X=9.435 $Y=1.505 $X2=0
+ $Y2=0
cc_1040 N_A_622_98#_c_1209_n N_VGND_c_2435_n 0.00659783f $X=10.155 $Y=0.34 $X2=0
+ $Y2=0
cc_1041 N_A_622_98#_c_1211_n N_VGND_c_2435_n 0.0167158f $X=10.32 $Y=1.065 $X2=0
+ $Y2=0
cc_1042 N_A_622_98#_c_1196_n N_VGND_c_2440_n 0.0038134f $X=4.31 $Y=1.34 $X2=0
+ $Y2=0
cc_1043 N_A_622_98#_c_1202_n N_VGND_c_2440_n 0.0184744f $X=4.95 $Y=0.33 $X2=0
+ $Y2=0
cc_1044 N_A_622_98#_c_1209_n N_VGND_c_2444_n 0.0574379f $X=10.155 $Y=0.34 $X2=0
+ $Y2=0
cc_1045 N_A_622_98#_c_1210_n N_VGND_c_2444_n 0.0115566f $X=9.615 $Y=0.34 $X2=0
+ $Y2=0
cc_1046 N_A_622_98#_c_1217_n N_VGND_c_2444_n 0.00278125f $X=10.32 $Y=0.9 $X2=0
+ $Y2=0
cc_1047 N_A_622_98#_c_1196_n N_VGND_c_2451_n 0.00508379f $X=4.31 $Y=1.34 $X2=0
+ $Y2=0
cc_1048 N_A_622_98#_c_1202_n N_VGND_c_2451_n 0.022448f $X=4.95 $Y=0.33 $X2=0
+ $Y2=0
cc_1049 N_A_622_98#_c_1209_n N_VGND_c_2451_n 0.0317788f $X=10.155 $Y=0.34 $X2=0
+ $Y2=0
cc_1050 N_A_622_98#_c_1210_n N_VGND_c_2451_n 0.00579705f $X=9.615 $Y=0.34 $X2=0
+ $Y2=0
cc_1051 N_A_622_98#_c_1217_n N_VGND_c_2451_n 0.00355513f $X=10.32 $Y=0.9 $X2=0
+ $Y2=0
cc_1052 N_A_622_98#_c_1209_n A_2061_74# 7.09228e-19 $X=10.155 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_1053 N_A_622_98#_c_1211_n A_2061_74# 0.00458877f $X=10.32 $Y=1.065 $X2=-0.19
+ $Y2=-0.245
cc_1054 N_A_877_98#_c_1453_n N_A_2037_442#_c_1601_n 0.0273058f $X=9.855 $Y=2.445
+ $X2=0 $Y2=0
cc_1055 N_A_877_98#_c_1453_n N_A_2037_442#_c_1613_n 0.0118417f $X=9.855 $Y=2.445
+ $X2=0 $Y2=0
cc_1056 N_A_877_98#_c_1447_n N_A_2037_442#_c_1613_n 0.00271626f $X=9.855 $Y=2.18
+ $X2=0 $Y2=0
cc_1057 N_A_877_98#_M1001_g N_A_1878_420#_c_1775_n 0.00163459f $X=9.685 $Y=0.87
+ $X2=0 $Y2=0
cc_1058 N_A_877_98#_c_1446_n N_A_1878_420#_c_1775_n 0.00843523f $X=9.87 $Y=1.295
+ $X2=0 $Y2=0
cc_1059 N_A_877_98#_c_1453_n N_A_1878_420#_c_1784_n 0.0217837f $X=9.855 $Y=2.445
+ $X2=0 $Y2=0
cc_1060 N_A_877_98#_c_1447_n N_A_1878_420#_c_1784_n 0.00226274f $X=9.855 $Y=2.18
+ $X2=0 $Y2=0
cc_1061 N_A_877_98#_c_1447_n N_A_1878_420#_c_1785_n 0.00609352f $X=9.855 $Y=2.18
+ $X2=0 $Y2=0
cc_1062 N_A_877_98#_c_1447_n N_A_1878_420#_c_1778_n 0.00562928f $X=9.855 $Y=2.18
+ $X2=0 $Y2=0
cc_1063 N_A_877_98#_c_1446_n N_A_1878_420#_c_1787_n 0.00105725f $X=9.87 $Y=1.295
+ $X2=0 $Y2=0
cc_1064 N_A_877_98#_c_1447_n N_A_1878_420#_c_1787_n 0.00619513f $X=9.855 $Y=2.18
+ $X2=0 $Y2=0
cc_1065 N_A_877_98#_c_1446_n N_A_1878_420#_c_1779_n 0.00121413f $X=9.87 $Y=1.295
+ $X2=0 $Y2=0
cc_1066 N_A_877_98#_c_1447_n N_A_1878_420#_c_1779_n 0.00777841f $X=9.855 $Y=2.18
+ $X2=0 $Y2=0
cc_1067 N_A_877_98#_c_1455_n N_VPWR_c_2015_n 0.0537794f $X=4.58 $Y=2.815 $X2=0
+ $Y2=0
cc_1068 N_A_877_98#_c_1455_n N_VPWR_c_2021_n 0.0214223f $X=4.58 $Y=2.815 $X2=0
+ $Y2=0
cc_1069 N_A_877_98#_c_1440_n N_VPWR_c_2012_n 9.39239e-19 $X=5.465 $Y=2.02 $X2=0
+ $Y2=0
cc_1070 N_A_877_98#_c_1455_n N_VPWR_c_2012_n 0.0174543f $X=4.58 $Y=2.815 $X2=0
+ $Y2=0
cc_1071 N_A_877_98#_c_1453_n N_VPWR_c_2038_n 9.59479e-19 $X=9.855 $Y=2.445 $X2=0
+ $Y2=0
cc_1072 N_A_877_98#_c_1440_n N_A_197_119#_c_2211_n 0.0116653f $X=5.465 $Y=2.02
+ $X2=0 $Y2=0
cc_1073 N_A_877_98#_c_1457_n N_A_197_119#_c_2211_n 0.0585791f $X=4.58 $Y=2.005
+ $X2=0 $Y2=0
cc_1074 N_A_877_98#_M1030_g N_A_197_119#_c_2200_n 5.35185e-19 $X=5.885 $Y=0.69
+ $X2=0 $Y2=0
cc_1075 N_A_877_98#_c_1448_n N_A_197_119#_c_2200_n 0.00139841f $X=4.735 $Y=1.085
+ $X2=0 $Y2=0
cc_1076 N_A_877_98#_c_1440_n N_A_197_119#_c_2201_n 0.00517817f $X=5.465 $Y=2.02
+ $X2=0 $Y2=0
cc_1077 N_A_877_98#_M1030_g N_A_197_119#_c_2201_n 0.00397398f $X=5.885 $Y=0.69
+ $X2=0 $Y2=0
cc_1078 N_A_877_98#_c_1450_n N_A_197_119#_c_2201_n 0.0082296f $X=5.325 $Y=1.53
+ $X2=0 $Y2=0
cc_1079 N_A_877_98#_c_1440_n N_A_197_119#_c_2202_n 0.00349791f $X=5.465 $Y=2.02
+ $X2=0 $Y2=0
cc_1080 N_A_877_98#_c_1448_n N_A_197_119#_c_2202_n 0.00917765f $X=4.735 $Y=1.085
+ $X2=0 $Y2=0
cc_1081 N_A_877_98#_c_1449_n N_A_197_119#_c_2202_n 0.00143475f $X=4.82 $Y=1.365
+ $X2=0 $Y2=0
cc_1082 N_A_877_98#_c_1450_n N_A_197_119#_c_2202_n 0.013637f $X=5.325 $Y=1.53
+ $X2=0 $Y2=0
cc_1083 N_A_877_98#_c_1440_n N_A_197_119#_c_2212_n 0.0142468f $X=5.465 $Y=2.02
+ $X2=0 $Y2=0
cc_1084 N_A_877_98#_c_1441_n N_A_197_119#_c_2212_n 0.00123656f $X=5.81 $Y=1.44
+ $X2=0 $Y2=0
cc_1085 N_A_877_98#_c_1450_n N_A_197_119#_c_2212_n 0.00282261f $X=5.325 $Y=1.53
+ $X2=0 $Y2=0
cc_1086 N_A_877_98#_c_1440_n N_A_197_119#_c_2213_n 0.00851906f $X=5.465 $Y=2.02
+ $X2=0 $Y2=0
cc_1087 N_A_877_98#_c_1450_n N_A_197_119#_c_2213_n 0.0280456f $X=5.325 $Y=1.53
+ $X2=0 $Y2=0
cc_1088 N_A_877_98#_c_1457_n N_A_197_119#_c_2213_n 0.0147868f $X=4.58 $Y=2.005
+ $X2=0 $Y2=0
cc_1089 N_A_877_98#_c_1440_n N_A_197_119#_c_2203_n 0.011099f $X=5.465 $Y=2.02
+ $X2=0 $Y2=0
cc_1090 N_A_877_98#_c_1441_n N_A_197_119#_c_2203_n 0.0135988f $X=5.81 $Y=1.44
+ $X2=0 $Y2=0
cc_1091 N_A_877_98#_M1030_g N_A_197_119#_c_2203_n 0.00384681f $X=5.885 $Y=0.69
+ $X2=0 $Y2=0
cc_1092 N_A_877_98#_c_1450_n N_A_197_119#_c_2203_n 0.0257448f $X=5.325 $Y=1.53
+ $X2=0 $Y2=0
cc_1093 N_A_877_98#_M1000_d N_A_197_119#_c_2205_n 0.00832489f $X=4.385 $Y=0.49
+ $X2=0 $Y2=0
cc_1094 N_A_877_98#_c_1448_n N_A_197_119#_c_2205_n 0.0364195f $X=4.735 $Y=1.085
+ $X2=0 $Y2=0
cc_1095 N_A_877_98#_c_1450_n N_A_197_119#_c_2205_n 0.00903718f $X=5.325 $Y=1.53
+ $X2=0 $Y2=0
cc_1096 N_A_877_98#_M1030_g N_VGND_c_2433_n 0.00602378f $X=5.885 $Y=0.69 $X2=0
+ $Y2=0
cc_1097 N_A_877_98#_c_1443_n N_VGND_c_2433_n 0.0283099f $X=9.61 $Y=0.18 $X2=0
+ $Y2=0
cc_1098 N_A_877_98#_c_1443_n N_VGND_c_2434_n 0.0210801f $X=9.61 $Y=0.18 $X2=0
+ $Y2=0
cc_1099 N_A_877_98#_M1001_g N_VGND_c_2434_n 0.00149617f $X=9.685 $Y=0.87 $X2=0
+ $Y2=0
cc_1100 N_A_877_98#_c_1444_n N_VGND_c_2440_n 0.0196812f $X=5.96 $Y=0.18 $X2=0
+ $Y2=0
cc_1101 N_A_877_98#_c_1443_n N_VGND_c_2442_n 0.0489606f $X=9.61 $Y=0.18 $X2=0
+ $Y2=0
cc_1102 N_A_877_98#_c_1443_n N_VGND_c_2444_n 0.0131953f $X=9.61 $Y=0.18 $X2=0
+ $Y2=0
cc_1103 N_A_877_98#_c_1443_n N_VGND_c_2451_n 0.0919547f $X=9.61 $Y=0.18 $X2=0
+ $Y2=0
cc_1104 N_A_877_98#_c_1444_n N_VGND_c_2451_n 0.00668353f $X=5.96 $Y=0.18 $X2=0
+ $Y2=0
cc_1105 N_A_877_98#_c_1443_n N_A_1418_125#_c_2600_n 0.0312071f $X=9.61 $Y=0.18
+ $X2=0 $Y2=0
cc_1106 N_A_2037_442#_c_1598_n N_A_1878_420#_c_1772_n 0.00245184f $X=12.13
+ $Y=1.97 $X2=0 $Y2=0
cc_1107 N_A_2037_442#_c_1655_n N_A_1878_420#_c_1772_n 0.00373128f $X=12.035
+ $Y=0.8 $X2=0 $Y2=0
cc_1108 N_A_2037_442#_c_1598_n N_A_1878_420#_c_1773_n 0.00639712f $X=12.13
+ $Y=1.97 $X2=0 $Y2=0
cc_1109 N_A_2037_442#_c_1626_n N_A_1878_420#_c_1773_n 9.21113e-19 $X=12.215
+ $Y=2.225 $X2=0 $Y2=0
cc_1110 N_A_2037_442#_c_1655_n N_A_1878_420#_c_1773_n 0.00250495f $X=12.035
+ $Y=0.8 $X2=0 $Y2=0
cc_1111 N_A_2037_442#_c_1598_n N_A_1878_420#_c_1783_n 7.4532e-19 $X=12.13
+ $Y=1.97 $X2=0 $Y2=0
cc_1112 N_A_2037_442#_c_1626_n N_A_1878_420#_c_1783_n 0.0215607f $X=12.215
+ $Y=2.225 $X2=0 $Y2=0
cc_1113 N_A_2037_442#_c_1614_n N_A_1878_420#_c_1783_n 0.00830144f $X=11.62
+ $Y=2.135 $X2=0 $Y2=0
cc_1114 N_A_2037_442#_M1047_g N_A_1878_420#_c_1776_n 0.00558533f $X=10.77
+ $Y=0.58 $X2=0 $Y2=0
cc_1115 N_A_2037_442#_c_1613_n N_A_1878_420#_c_1776_n 4.02351e-19 $X=10.63
+ $Y=2.195 $X2=0 $Y2=0
cc_1116 N_A_2037_442#_M1047_g N_A_1878_420#_c_1777_n 4.92357e-19 $X=10.77
+ $Y=0.58 $X2=0 $Y2=0
cc_1117 N_A_2037_442#_c_1626_n N_A_1878_420#_c_1777_n 0.00107002f $X=12.215
+ $Y=2.225 $X2=0 $Y2=0
cc_1118 N_A_2037_442#_c_1601_n N_A_1878_420#_c_1784_n 3.04665e-19 $X=10.275
+ $Y=2.445 $X2=0 $Y2=0
cc_1119 N_A_2037_442#_c_1613_n N_A_1878_420#_c_1784_n 2.40682e-19 $X=10.63
+ $Y=2.195 $X2=0 $Y2=0
cc_1120 N_A_2037_442#_M1047_g N_A_1878_420#_c_1780_n 0.017157f $X=10.77 $Y=0.58
+ $X2=0 $Y2=0
cc_1121 N_A_2037_442#_c_1598_n N_A_1878_420#_c_1781_n 0.026731f $X=12.13 $Y=1.97
+ $X2=0 $Y2=0
cc_1122 N_A_2037_442#_c_1626_n N_A_1878_420#_c_1781_n 0.00841365f $X=12.215
+ $Y=2.225 $X2=0 $Y2=0
cc_1123 N_A_2037_442#_c_1592_n N_RESET_B_c_1889_n 0.0490953f $X=13.73 $Y=1.665
+ $X2=-0.19 $Y2=-0.245
cc_1124 N_A_2037_442#_c_1610_n N_RESET_B_c_1889_n 0.0190656f $X=13.53 $Y=2.225
+ $X2=-0.19 $Y2=-0.245
cc_1125 N_A_2037_442#_c_1599_n N_RESET_B_c_1889_n 0.00690416f $X=13.615 $Y=2.14
+ $X2=-0.19 $Y2=-0.245
cc_1126 N_A_2037_442#_c_1600_n N_RESET_B_c_1889_n 0.00193552f $X=13.75 $Y=1.385
+ $X2=-0.19 $Y2=-0.245
cc_1127 N_A_2037_442#_c_1591_n N_RESET_B_c_1890_n 0.0114189f $X=13.72 $Y=1.22
+ $X2=0 $Y2=0
cc_1128 N_A_2037_442#_c_1591_n RESET_B 8.15883e-19 $X=13.72 $Y=1.22 $X2=0 $Y2=0
cc_1129 N_A_2037_442#_c_1592_n RESET_B 3.55566e-19 $X=13.73 $Y=1.665 $X2=0 $Y2=0
cc_1130 N_A_2037_442#_c_1610_n RESET_B 0.00460648f $X=13.53 $Y=2.225 $X2=0 $Y2=0
cc_1131 N_A_2037_442#_c_1600_n RESET_B 0.0261964f $X=13.75 $Y=1.385 $X2=0 $Y2=0
cc_1132 N_A_2037_442#_c_1605_n N_A_2881_74#_c_1921_n 0.00331969f $X=14.76
+ $Y=1.97 $X2=0 $Y2=0
cc_1133 N_A_2037_442#_c_1596_n N_A_2881_74#_M1003_g 0.0183151f $X=14.765
+ $Y=0.995 $X2=0 $Y2=0
cc_1134 N_A_2037_442#_c_1605_n N_A_2881_74#_c_1923_n 0.00540482f $X=14.76
+ $Y=1.97 $X2=0 $Y2=0
cc_1135 N_A_2037_442#_c_1607_n N_A_2881_74#_c_1923_n 0.0167542f $X=14.835
+ $Y=2.045 $X2=0 $Y2=0
cc_1136 N_A_2037_442#_c_1591_n N_A_2881_74#_c_1924_n 7.54105e-19 $X=13.72
+ $Y=1.22 $X2=0 $Y2=0
cc_1137 N_A_2037_442#_c_1595_n N_A_2881_74#_c_1924_n 0.0176565f $X=14.69 $Y=1.07
+ $X2=0 $Y2=0
cc_1138 N_A_2037_442#_c_1596_n N_A_2881_74#_c_1924_n 0.0124552f $X=14.765
+ $Y=0.995 $X2=0 $Y2=0
cc_1139 N_A_2037_442#_c_1597_n N_A_2881_74#_c_1924_n 0.00378707f $X=14.23
+ $Y=1.07 $X2=0 $Y2=0
cc_1140 N_A_2037_442#_c_1592_n N_A_2881_74#_c_1928_n 0.00317173f $X=13.73
+ $Y=1.665 $X2=0 $Y2=0
cc_1141 N_A_2037_442#_c_1605_n N_A_2881_74#_c_1928_n 0.0208441f $X=14.76 $Y=1.97
+ $X2=0 $Y2=0
cc_1142 N_A_2037_442#_c_1607_n N_A_2881_74#_c_1928_n 0.0148293f $X=14.835
+ $Y=2.045 $X2=0 $Y2=0
cc_1143 N_A_2037_442#_c_1594_n N_A_2881_74#_c_1925_n 0.00378707f $X=14.23
+ $Y=1.895 $X2=0 $Y2=0
cc_1144 N_A_2037_442#_c_1595_n N_A_2881_74#_c_1925_n 9.58601e-19 $X=14.69
+ $Y=1.07 $X2=0 $Y2=0
cc_1145 N_A_2037_442#_c_1605_n N_A_2881_74#_c_1925_n 5.31902e-19 $X=14.76
+ $Y=1.97 $X2=0 $Y2=0
cc_1146 N_A_2037_442#_c_1595_n N_A_2881_74#_c_1926_n 0.0212545f $X=14.69 $Y=1.07
+ $X2=0 $Y2=0
cc_1147 N_A_2037_442#_c_1605_n N_A_2881_74#_c_1926_n 0.0214695f $X=14.76 $Y=1.97
+ $X2=0 $Y2=0
cc_1148 N_A_2037_442#_c_1597_n N_A_2881_74#_c_1926_n 0.0195557f $X=14.23 $Y=1.07
+ $X2=0 $Y2=0
cc_1149 N_A_2037_442#_c_1608_n N_VPWR_M1036_d 0.00520498f $X=11.535 $Y=2.405
+ $X2=0 $Y2=0
cc_1150 N_A_2037_442#_c_1610_n N_VPWR_M1017_d 0.00669951f $X=13.53 $Y=2.225
+ $X2=0 $Y2=0
cc_1151 N_A_2037_442#_c_1610_n N_VPWR_M1028_d 0.00906824f $X=13.53 $Y=2.225
+ $X2=0 $Y2=0
cc_1152 N_A_2037_442#_c_1599_n N_VPWR_M1028_d 0.0048099f $X=13.615 $Y=2.14 $X2=0
+ $Y2=0
cc_1153 N_A_2037_442#_c_1610_n N_VPWR_c_2018_n 0.0220389f $X=13.53 $Y=2.225
+ $X2=0 $Y2=0
cc_1154 N_A_2037_442#_c_1626_n N_VPWR_c_2018_n 3.24411e-19 $X=12.215 $Y=2.225
+ $X2=0 $Y2=0
cc_1155 N_A_2037_442#_c_1614_n N_VPWR_c_2018_n 0.0146625f $X=11.62 $Y=2.135
+ $X2=0 $Y2=0
cc_1156 N_A_2037_442#_c_1592_n N_VPWR_c_2019_n 0.0122151f $X=13.73 $Y=1.665
+ $X2=0 $Y2=0
cc_1157 N_A_2037_442#_c_1610_n N_VPWR_c_2019_n 0.0224192f $X=13.53 $Y=2.225
+ $X2=0 $Y2=0
cc_1158 N_A_2037_442#_c_1607_n N_VPWR_c_2020_n 0.0078018f $X=14.835 $Y=2.045
+ $X2=0 $Y2=0
cc_1159 N_A_2037_442#_c_1614_n N_VPWR_c_2023_n 0.0110241f $X=11.62 $Y=2.135
+ $X2=0 $Y2=0
cc_1160 N_A_2037_442#_c_1592_n N_VPWR_c_2031_n 0.00455225f $X=13.73 $Y=1.665
+ $X2=0 $Y2=0
cc_1161 N_A_2037_442#_c_1607_n N_VPWR_c_2031_n 0.00445602f $X=14.835 $Y=2.045
+ $X2=0 $Y2=0
cc_1162 N_A_2037_442#_c_1601_n N_VPWR_c_2012_n 0.00305691f $X=10.275 $Y=2.445
+ $X2=0 $Y2=0
cc_1163 N_A_2037_442#_c_1592_n N_VPWR_c_2012_n 0.00466424f $X=13.73 $Y=1.665
+ $X2=0 $Y2=0
cc_1164 N_A_2037_442#_c_1607_n N_VPWR_c_2012_n 0.00862315f $X=14.835 $Y=2.045
+ $X2=0 $Y2=0
cc_1165 N_A_2037_442#_c_1608_n N_VPWR_c_2012_n 0.0133547f $X=11.535 $Y=2.405
+ $X2=0 $Y2=0
cc_1166 N_A_2037_442#_c_1612_n N_VPWR_c_2012_n 0.00115284f $X=10.63 $Y=2.195
+ $X2=0 $Y2=0
cc_1167 N_A_2037_442#_c_1613_n N_VPWR_c_2012_n 3.16035e-19 $X=10.63 $Y=2.195
+ $X2=0 $Y2=0
cc_1168 N_A_2037_442#_c_1614_n N_VPWR_c_2012_n 0.00909194f $X=11.62 $Y=2.135
+ $X2=0 $Y2=0
cc_1169 N_A_2037_442#_c_1601_n N_VPWR_c_2038_n 0.00360789f $X=10.275 $Y=2.445
+ $X2=0 $Y2=0
cc_1170 N_A_2037_442#_c_1601_n N_VPWR_c_2039_n 0.00906542f $X=10.275 $Y=2.445
+ $X2=0 $Y2=0
cc_1171 N_A_2037_442#_c_1608_n N_VPWR_c_2039_n 0.0283172f $X=11.535 $Y=2.405
+ $X2=0 $Y2=0
cc_1172 N_A_2037_442#_c_1612_n N_VPWR_c_2039_n 0.028442f $X=10.63 $Y=2.195 $X2=0
+ $Y2=0
cc_1173 N_A_2037_442#_c_1613_n N_VPWR_c_2039_n 0.00327848f $X=10.63 $Y=2.195
+ $X2=0 $Y2=0
cc_1174 N_A_2037_442#_c_1614_n N_VPWR_c_2039_n 0.0146722f $X=11.62 $Y=2.135
+ $X2=0 $Y2=0
cc_1175 N_A_2037_442#_c_1626_n A_2384_392# 0.0069385f $X=12.215 $Y=2.225
+ $X2=-0.19 $Y2=-0.245
cc_1176 N_A_2037_442#_c_1591_n N_Q_N_c_2376_n 0.00885704f $X=13.72 $Y=1.22 $X2=0
+ $Y2=0
cc_1177 N_A_2037_442#_c_1592_n N_Q_N_c_2376_n 0.00469661f $X=13.73 $Y=1.665
+ $X2=0 $Y2=0
cc_1178 N_A_2037_442#_c_1596_n N_Q_N_c_2376_n 0.00183613f $X=14.765 $Y=0.995
+ $X2=0 $Y2=0
cc_1179 N_A_2037_442#_c_1597_n N_Q_N_c_2376_n 0.00500792f $X=14.23 $Y=1.07 $X2=0
+ $Y2=0
cc_1180 N_A_2037_442#_c_1600_n N_Q_N_c_2376_n 0.00924171f $X=13.75 $Y=1.385
+ $X2=0 $Y2=0
cc_1181 N_A_2037_442#_c_1592_n N_Q_N_c_2378_n 0.0102635f $X=13.73 $Y=1.665 $X2=0
+ $Y2=0
cc_1182 N_A_2037_442#_c_1593_n N_Q_N_c_2378_n 0.00425199f $X=14.155 $Y=1.295
+ $X2=0 $Y2=0
cc_1183 N_A_2037_442#_c_1594_n N_Q_N_c_2378_n 0.00573682f $X=14.23 $Y=1.895
+ $X2=0 $Y2=0
cc_1184 N_A_2037_442#_c_1606_n N_Q_N_c_2378_n 0.00100169f $X=14.305 $Y=1.97
+ $X2=0 $Y2=0
cc_1185 N_A_2037_442#_c_1599_n N_Q_N_c_2378_n 0.0315553f $X=13.615 $Y=2.14 $X2=0
+ $Y2=0
cc_1186 N_A_2037_442#_c_1600_n N_Q_N_c_2378_n 0.00371067f $X=13.75 $Y=1.385
+ $X2=0 $Y2=0
cc_1187 N_A_2037_442#_c_1591_n N_Q_N_c_2377_n 0.00217368f $X=13.72 $Y=1.22 $X2=0
+ $Y2=0
cc_1188 N_A_2037_442#_c_1592_n N_Q_N_c_2377_n 0.00140406f $X=13.73 $Y=1.665
+ $X2=0 $Y2=0
cc_1189 N_A_2037_442#_c_1593_n N_Q_N_c_2377_n 0.00403922f $X=14.155 $Y=1.295
+ $X2=0 $Y2=0
cc_1190 N_A_2037_442#_c_1594_n N_Q_N_c_2377_n 0.00774786f $X=14.23 $Y=1.895
+ $X2=0 $Y2=0
cc_1191 N_A_2037_442#_c_1597_n N_Q_N_c_2377_n 0.00837031f $X=14.23 $Y=1.07 $X2=0
+ $Y2=0
cc_1192 N_A_2037_442#_c_1599_n N_Q_N_c_2377_n 0.00447794f $X=13.615 $Y=2.14
+ $X2=0 $Y2=0
cc_1193 N_A_2037_442#_c_1600_n N_Q_N_c_2377_n 0.0224758f $X=13.75 $Y=1.385 $X2=0
+ $Y2=0
cc_1194 N_A_2037_442#_c_1606_n Q_N 0.00751751f $X=14.305 $Y=1.97 $X2=0 $Y2=0
cc_1195 N_A_2037_442#_c_1607_n Q_N 0.00182123f $X=14.835 $Y=2.045 $X2=0 $Y2=0
cc_1196 N_A_2037_442#_c_1610_n Q_N 0.0142209f $X=13.53 $Y=2.225 $X2=0 $Y2=0
cc_1197 N_A_2037_442#_c_1605_n Q 6.13961e-19 $X=14.76 $Y=1.97 $X2=0 $Y2=0
cc_1198 N_A_2037_442#_c_1596_n Q 0.00119534f $X=14.765 $Y=0.995 $X2=0 $Y2=0
cc_1199 N_A_2037_442#_c_1607_n Q 4.34701e-19 $X=14.835 $Y=2.045 $X2=0 $Y2=0
cc_1200 N_A_2037_442#_M1047_g N_VGND_c_2435_n 0.0065354f $X=10.77 $Y=0.58 $X2=0
+ $Y2=0
cc_1201 N_A_2037_442#_c_1591_n N_VGND_c_2436_n 0.00899543f $X=13.72 $Y=1.22
+ $X2=0 $Y2=0
cc_1202 N_A_2037_442#_c_1600_n N_VGND_c_2436_n 0.00418987f $X=13.75 $Y=1.385
+ $X2=0 $Y2=0
cc_1203 N_A_2037_442#_c_1596_n N_VGND_c_2437_n 0.00686847f $X=14.765 $Y=0.995
+ $X2=0 $Y2=0
cc_1204 N_A_2037_442#_M1047_g N_VGND_c_2444_n 0.00461464f $X=10.77 $Y=0.58 $X2=0
+ $Y2=0
cc_1205 N_A_2037_442#_c_1591_n N_VGND_c_2449_n 0.00434272f $X=13.72 $Y=1.22
+ $X2=0 $Y2=0
cc_1206 N_A_2037_442#_c_1596_n N_VGND_c_2449_n 0.00434272f $X=14.765 $Y=0.995
+ $X2=0 $Y2=0
cc_1207 N_A_2037_442#_M1047_g N_VGND_c_2451_n 0.00910155f $X=10.77 $Y=0.58 $X2=0
+ $Y2=0
cc_1208 N_A_2037_442#_c_1591_n N_VGND_c_2451_n 0.00830282f $X=13.72 $Y=1.22
+ $X2=0 $Y2=0
cc_1209 N_A_2037_442#_c_1596_n N_VGND_c_2451_n 0.00826607f $X=14.765 $Y=0.995
+ $X2=0 $Y2=0
cc_1210 N_A_2037_442#_c_1655_n N_A_2271_74#_c_2628_n 0.0274769f $X=12.035 $Y=0.8
+ $X2=0 $Y2=0
cc_1211 N_A_2037_442#_M1031_d N_A_2271_74#_c_2626_n 0.00382184f $X=11.785
+ $Y=0.37 $X2=0 $Y2=0
cc_1212 N_A_2037_442#_c_1655_n N_A_2271_74#_c_2626_n 0.0210917f $X=12.035 $Y=0.8
+ $X2=0 $Y2=0
cc_1213 N_A_2037_442#_c_1655_n N_A_2271_74#_c_2633_n 0.0307483f $X=12.035 $Y=0.8
+ $X2=0 $Y2=0
cc_1214 N_A_1878_420#_c_1783_n N_VPWR_c_2018_n 0.00195012f $X=11.845 $Y=1.885
+ $X2=0 $Y2=0
cc_1215 N_A_1878_420#_c_1783_n N_VPWR_c_2023_n 0.00445602f $X=11.845 $Y=1.885
+ $X2=0 $Y2=0
cc_1216 N_A_1878_420#_c_1783_n N_VPWR_c_2012_n 0.00858771f $X=11.845 $Y=1.885
+ $X2=0 $Y2=0
cc_1217 N_A_1878_420#_c_1777_n N_VGND_c_2435_n 0.0186013f $X=11.595 $Y=1.265
+ $X2=0 $Y2=0
cc_1218 N_A_1878_420#_c_1772_n N_VGND_c_2446_n 0.00278247f $X=11.71 $Y=1.22
+ $X2=0 $Y2=0
cc_1219 N_A_1878_420#_c_1772_n N_VGND_c_2451_n 0.00354553f $X=11.71 $Y=1.22
+ $X2=0 $Y2=0
cc_1220 N_A_1878_420#_c_1772_n N_A_2271_74#_c_2628_n 0.00869767f $X=11.71
+ $Y=1.22 $X2=0 $Y2=0
cc_1221 N_A_1878_420#_c_1777_n N_A_2271_74#_c_2628_n 0.0168759f $X=11.595
+ $Y=1.265 $X2=0 $Y2=0
cc_1222 N_A_1878_420#_c_1781_n N_A_2271_74#_c_2628_n 0.00340264f $X=11.735
+ $Y=1.265 $X2=0 $Y2=0
cc_1223 N_A_1878_420#_c_1772_n N_A_2271_74#_c_2626_n 0.0105911f $X=11.71 $Y=1.22
+ $X2=0 $Y2=0
cc_1224 N_A_1878_420#_c_1772_n N_A_2271_74#_c_2627_n 0.00184834f $X=11.71
+ $Y=1.22 $X2=0 $Y2=0
cc_1225 N_RESET_B_c_1889_n N_VPWR_c_2018_n 7.75483e-19 $X=13.215 $Y=1.665 $X2=0
+ $Y2=0
cc_1226 N_RESET_B_c_1889_n N_VPWR_c_2019_n 8.5114e-19 $X=13.215 $Y=1.665 $X2=0
+ $Y2=0
cc_1227 N_RESET_B_c_1889_n N_VPWR_c_2012_n 0.00388259f $X=13.215 $Y=1.665 $X2=0
+ $Y2=0
cc_1228 N_RESET_B_c_1890_n N_Q_N_c_2376_n 3.29774e-19 $X=13.245 $Y=1.22 $X2=0
+ $Y2=0
cc_1229 N_RESET_B_c_1890_n N_VGND_c_2436_n 0.0106582f $X=13.245 $Y=1.22 $X2=0
+ $Y2=0
cc_1230 RESET_B N_VGND_c_2436_n 0.00341404f $X=13.115 $Y=1.21 $X2=0 $Y2=0
cc_1231 N_RESET_B_c_1890_n N_VGND_c_2446_n 0.00318082f $X=13.245 $Y=1.22 $X2=0
+ $Y2=0
cc_1232 N_RESET_B_c_1890_n N_VGND_c_2451_n 0.0037954f $X=13.245 $Y=1.22 $X2=0
+ $Y2=0
cc_1233 N_RESET_B_c_1890_n N_A_2271_74#_c_2633_n 0.00273771f $X=13.245 $Y=1.22
+ $X2=0 $Y2=0
cc_1234 N_A_2881_74#_c_1921_n N_VPWR_c_2020_n 0.00671978f $X=15.255 $Y=1.43
+ $X2=0 $Y2=0
cc_1235 N_A_2881_74#_c_1923_n N_VPWR_c_2020_n 0.0066161f $X=15.345 $Y=1.765
+ $X2=0 $Y2=0
cc_1236 N_A_2881_74#_c_1928_n N_VPWR_c_2020_n 0.0333798f $X=14.61 $Y=2.265 $X2=0
+ $Y2=0
cc_1237 N_A_2881_74#_c_1928_n N_VPWR_c_2031_n 0.0145938f $X=14.61 $Y=2.265 $X2=0
+ $Y2=0
cc_1238 N_A_2881_74#_c_1923_n N_VPWR_c_2032_n 0.00434272f $X=15.345 $Y=1.765
+ $X2=0 $Y2=0
cc_1239 N_A_2881_74#_c_1923_n N_VPWR_c_2012_n 0.00824959f $X=15.345 $Y=1.765
+ $X2=0 $Y2=0
cc_1240 N_A_2881_74#_c_1928_n N_VPWR_c_2012_n 0.0120466f $X=14.61 $Y=2.265 $X2=0
+ $Y2=0
cc_1241 N_A_2881_74#_c_1924_n N_Q_N_c_2376_n 0.0686037f $X=14.55 $Y=0.645 $X2=0
+ $Y2=0
cc_1242 N_A_2881_74#_c_1928_n N_Q_N_c_2378_n 0.0686037f $X=14.61 $Y=2.265 $X2=0
+ $Y2=0
cc_1243 N_A_2881_74#_c_1925_n N_Q_N_c_2377_n 0.0686037f $X=14.68 $Y=1.52 $X2=0
+ $Y2=0
cc_1244 N_A_2881_74#_c_1926_n N_Q_N_c_2377_n 3.41194e-19 $X=14.68 $Y=1.43 $X2=0
+ $Y2=0
cc_1245 N_A_2881_74#_M1003_g Q 0.0262142f $X=15.345 $Y=0.74 $X2=0 $Y2=0
cc_1246 N_A_2881_74#_c_1923_n Q 0.0382855f $X=15.345 $Y=1.765 $X2=0 $Y2=0
cc_1247 N_A_2881_74#_c_1928_n Q 0.0118616f $X=14.61 $Y=2.265 $X2=0 $Y2=0
cc_1248 N_A_2881_74#_c_1925_n Q 0.0096057f $X=14.68 $Y=1.52 $X2=0 $Y2=0
cc_1249 N_A_2881_74#_c_1926_n Q 6.15324e-19 $X=14.68 $Y=1.43 $X2=0 $Y2=0
cc_1250 N_A_2881_74#_c_1921_n N_VGND_c_2437_n 0.0102009f $X=15.255 $Y=1.43 $X2=0
+ $Y2=0
cc_1251 N_A_2881_74#_M1003_g N_VGND_c_2437_n 0.00691628f $X=15.345 $Y=0.74 $X2=0
+ $Y2=0
cc_1252 N_A_2881_74#_c_1924_n N_VGND_c_2437_n 0.0220246f $X=14.55 $Y=0.645 $X2=0
+ $Y2=0
cc_1253 N_A_2881_74#_c_1924_n N_VGND_c_2449_n 0.0118867f $X=14.55 $Y=0.645 $X2=0
+ $Y2=0
cc_1254 N_A_2881_74#_M1003_g N_VGND_c_2450_n 0.00434272f $X=15.345 $Y=0.74 $X2=0
+ $Y2=0
cc_1255 N_A_2881_74#_M1003_g N_VGND_c_2451_n 0.00825042f $X=15.345 $Y=0.74 $X2=0
+ $Y2=0
cc_1256 N_A_2881_74#_c_1924_n N_VGND_c_2451_n 0.00978237f $X=14.55 $Y=0.645
+ $X2=0 $Y2=0
cc_1257 N_A_27_464#_c_1971_n N_VPWR_M1026_d 0.00258237f $X=1.115 $Y=2.39
+ $X2=-0.19 $Y2=1.66
cc_1258 N_A_27_464#_c_1971_n N_VPWR_c_2013_n 0.0198565f $X=1.115 $Y=2.39 $X2=0
+ $Y2=0
cc_1259 N_A_27_464#_c_1973_n N_VPWR_c_2013_n 0.0117236f $X=1.285 $Y=2.99 $X2=0
+ $Y2=0
cc_1260 N_A_27_464#_c_1975_n N_VPWR_c_2013_n 0.0133605f $X=0.28 $Y=2.47 $X2=0
+ $Y2=0
cc_1261 N_A_27_464#_c_1972_n N_VPWR_c_2014_n 0.0119251f $X=1.945 $Y=2.99 $X2=0
+ $Y2=0
cc_1262 N_A_27_464#_c_1974_n N_VPWR_c_2014_n 0.0253882f $X=2.11 $Y=2.75 $X2=0
+ $Y2=0
cc_1263 N_A_27_464#_c_1975_n N_VPWR_c_2027_n 0.014586f $X=0.28 $Y=2.47 $X2=0
+ $Y2=0
cc_1264 N_A_27_464#_c_1972_n N_VPWR_c_2028_n 0.0648791f $X=1.945 $Y=2.99 $X2=0
+ $Y2=0
cc_1265 N_A_27_464#_c_1973_n N_VPWR_c_2028_n 0.0121505f $X=1.285 $Y=2.99 $X2=0
+ $Y2=0
cc_1266 N_A_27_464#_c_1971_n N_VPWR_c_2012_n 0.010659f $X=1.115 $Y=2.39 $X2=0
+ $Y2=0
cc_1267 N_A_27_464#_c_1972_n N_VPWR_c_2012_n 0.0362041f $X=1.945 $Y=2.99 $X2=0
+ $Y2=0
cc_1268 N_A_27_464#_c_1973_n N_VPWR_c_2012_n 0.00660393f $X=1.285 $Y=2.99 $X2=0
+ $Y2=0
cc_1269 N_A_27_464#_c_1975_n N_VPWR_c_2012_n 0.0120436f $X=0.28 $Y=2.47 $X2=0
+ $Y2=0
cc_1270 N_A_27_464#_c_1971_n A_218_464# 0.00155866f $X=1.115 $Y=2.39 $X2=-0.19
+ $Y2=1.66
cc_1271 N_A_27_464#_c_1981_n A_218_464# 0.00558502f $X=1.2 $Y=2.905 $X2=-0.19
+ $Y2=1.66
cc_1272 N_A_27_464#_c_1972_n A_218_464# 6.48644e-19 $X=1.945 $Y=2.99 $X2=-0.19
+ $Y2=1.66
cc_1273 N_A_27_464#_c_1972_n N_A_197_119#_M1010_d 0.00222494f $X=1.945 $Y=2.99
+ $X2=0 $Y2=0
cc_1274 N_A_27_464#_c_1971_n N_A_197_119#_c_2207_n 0.0117279f $X=1.115 $Y=2.39
+ $X2=0 $Y2=0
cc_1275 N_A_27_464#_c_1981_n N_A_197_119#_c_2207_n 0.0159385f $X=1.2 $Y=2.905
+ $X2=0 $Y2=0
cc_1276 N_A_27_464#_c_1972_n N_A_197_119#_c_2207_n 0.014518f $X=1.945 $Y=2.99
+ $X2=0 $Y2=0
cc_1277 N_A_27_464#_c_1974_n N_A_197_119#_c_2207_n 0.014416f $X=2.11 $Y=2.75
+ $X2=0 $Y2=0
cc_1278 N_A_27_464#_c_1974_n N_A_197_119#_c_2208_n 0.00668276f $X=2.11 $Y=2.75
+ $X2=0 $Y2=0
cc_1279 N_VPWR_c_2021_n N_A_197_119#_c_2211_n 0.00751822f $X=6.595 $Y=3.33 $X2=0
+ $Y2=0
cc_1280 N_VPWR_c_2012_n N_A_197_119#_c_2211_n 0.00908407f $X=15.6 $Y=3.33 $X2=0
+ $Y2=0
cc_1281 N_VPWR_c_2019_n Q_N 0.0285837f $X=13.505 $Y=2.645 $X2=0 $Y2=0
cc_1282 N_VPWR_c_2031_n Q_N 0.0131779f $X=14.945 $Y=3.33 $X2=0 $Y2=0
cc_1283 N_VPWR_c_2012_n Q_N 0.0140512f $X=15.6 $Y=3.33 $X2=0 $Y2=0
cc_1284 N_VPWR_c_2020_n Q 0.0606769f $X=15.115 $Y=2.28 $X2=0 $Y2=0
cc_1285 N_VPWR_c_2032_n Q 0.0150101f $X=15.6 $Y=3.33 $X2=0 $Y2=0
cc_1286 N_VPWR_c_2012_n Q 0.0123677f $X=15.6 $Y=3.33 $X2=0 $Y2=0
cc_1287 N_A_197_119#_c_2196_n N_VGND_M1012_d 0.00383506f $X=2.335 $Y=1.185 $X2=0
+ $Y2=0
cc_1288 N_A_197_119#_c_2199_n N_VGND_M1042_d 0.00272968f $X=3.595 $Y=0.66 $X2=0
+ $Y2=0
cc_1289 N_A_197_119#_c_2272_n N_VGND_M1042_d 0.00103672f $X=3.68 $Y=0.745 $X2=0
+ $Y2=0
cc_1290 N_A_197_119#_c_2205_n N_VGND_M1042_d 0.0191365f $X=5.005 $Y=0.645 $X2=0
+ $Y2=0
cc_1291 N_A_197_119#_c_2192_n N_VGND_c_2430_n 0.0055977f $X=1.205 $Y=0.805 $X2=0
+ $Y2=0
cc_1292 N_A_197_119#_c_2192_n N_VGND_c_2431_n 0.0144146f $X=1.205 $Y=0.805 $X2=0
+ $Y2=0
cc_1293 N_A_197_119#_c_2193_n N_VGND_c_2431_n 0.0168484f $X=1.935 $Y=1.27 $X2=0
+ $Y2=0
cc_1294 N_A_197_119#_c_2196_n N_VGND_c_2431_n 0.0445613f $X=2.335 $Y=1.185 $X2=0
+ $Y2=0
cc_1295 N_A_197_119#_c_2198_n N_VGND_c_2431_n 0.0147451f $X=2.42 $Y=0.34 $X2=0
+ $Y2=0
cc_1296 N_A_197_119#_c_2197_n N_VGND_c_2432_n 0.0150381f $X=3.51 $Y=0.34 $X2=0
+ $Y2=0
cc_1297 N_A_197_119#_c_2199_n N_VGND_c_2432_n 0.00511549f $X=3.595 $Y=0.66 $X2=0
+ $Y2=0
cc_1298 N_A_197_119#_c_2205_n N_VGND_c_2432_n 0.0251653f $X=5.005 $Y=0.645 $X2=0
+ $Y2=0
cc_1299 N_A_197_119#_c_2192_n N_VGND_c_2438_n 0.00749591f $X=1.205 $Y=0.805
+ $X2=0 $Y2=0
cc_1300 N_A_197_119#_c_2205_n N_VGND_c_2440_n 0.0125652f $X=5.005 $Y=0.645 $X2=0
+ $Y2=0
cc_1301 N_A_197_119#_c_2206_n N_VGND_c_2440_n 0.00964446f $X=5.25 $Y=0.645 $X2=0
+ $Y2=0
cc_1302 N_A_197_119#_c_2197_n N_VGND_c_2448_n 0.0818011f $X=3.51 $Y=0.34 $X2=0
+ $Y2=0
cc_1303 N_A_197_119#_c_2198_n N_VGND_c_2448_n 0.0115566f $X=2.42 $Y=0.34 $X2=0
+ $Y2=0
cc_1304 N_A_197_119#_c_2205_n N_VGND_c_2448_n 0.00279509f $X=5.005 $Y=0.645
+ $X2=0 $Y2=0
cc_1305 N_A_197_119#_c_2192_n N_VGND_c_2451_n 0.00907254f $X=1.205 $Y=0.805
+ $X2=0 $Y2=0
cc_1306 N_A_197_119#_c_2197_n N_VGND_c_2451_n 0.0469402f $X=3.51 $Y=0.34 $X2=0
+ $Y2=0
cc_1307 N_A_197_119#_c_2198_n N_VGND_c_2451_n 0.00579705f $X=2.42 $Y=0.34 $X2=0
+ $Y2=0
cc_1308 N_A_197_119#_c_2205_n N_VGND_c_2451_n 0.0290319f $X=5.005 $Y=0.645 $X2=0
+ $Y2=0
cc_1309 N_A_197_119#_c_2206_n N_VGND_c_2451_n 0.0110526f $X=5.25 $Y=0.645 $X2=0
+ $Y2=0
cc_1310 N_Q_N_c_2376_n N_VGND_c_2436_n 0.0256095f $X=13.935 $Y=0.515 $X2=0 $Y2=0
cc_1311 N_Q_N_c_2376_n N_VGND_c_2449_n 0.022404f $X=13.935 $Y=0.515 $X2=0 $Y2=0
cc_1312 N_Q_N_c_2376_n N_VGND_c_2451_n 0.018474f $X=13.935 $Y=0.515 $X2=0 $Y2=0
cc_1313 Q N_VGND_c_2437_n 0.0230301f $X=15.515 $Y=0.47 $X2=0 $Y2=0
cc_1314 Q N_VGND_c_2450_n 0.0150101f $X=15.515 $Y=0.47 $X2=0 $Y2=0
cc_1315 Q N_VGND_c_2451_n 0.0123677f $X=15.515 $Y=0.47 $X2=0 $Y2=0
cc_1316 N_VGND_c_2433_n N_A_1418_125#_c_2600_n 0.0163753f $X=6.685 $Y=0.475
+ $X2=0 $Y2=0
cc_1317 N_VGND_c_2442_n N_A_1418_125#_c_2600_n 0.076244f $X=9.025 $Y=0 $X2=0
+ $Y2=0
cc_1318 N_VGND_c_2451_n N_A_1418_125#_c_2600_n 0.0510536f $X=15.6 $Y=0 $X2=0
+ $Y2=0
cc_1319 N_VGND_c_2434_n N_A_1418_125#_c_2602_n 0.0139605f $X=9.11 $Y=0.845 $X2=0
+ $Y2=0
cc_1320 N_VGND_c_2446_n N_A_2271_74#_c_2626_n 0.0580341f $X=13.295 $Y=0 $X2=0
+ $Y2=0
cc_1321 N_VGND_c_2451_n N_A_2271_74#_c_2626_n 0.0326087f $X=15.6 $Y=0 $X2=0
+ $Y2=0
cc_1322 N_VGND_c_2435_n N_A_2271_74#_c_2627_n 0.0112234f $X=11.065 $Y=0.505
+ $X2=0 $Y2=0
cc_1323 N_VGND_c_2446_n N_A_2271_74#_c_2627_n 0.0234809f $X=13.295 $Y=0 $X2=0
+ $Y2=0
cc_1324 N_VGND_c_2451_n N_A_2271_74#_c_2627_n 0.0126009f $X=15.6 $Y=0 $X2=0
+ $Y2=0
