* File: sky130_fd_sc_ls__xor3_2.pxi.spice
* Created: Fri Aug 28 14:11:00 2020
* 
x_PM_SKY130_FD_SC_LS__XOR3_2%A_83_289# N_A_83_289#_M1022_d N_A_83_289#_M1020_d
+ N_A_83_289#_M1006_d N_A_83_289#_M1003_d N_A_83_289#_M1017_g
+ N_A_83_289#_c_197_n N_A_83_289#_M1000_g N_A_83_289#_c_198_n
+ N_A_83_289#_c_204_n N_A_83_289#_c_258_p N_A_83_289#_c_216_p
+ N_A_83_289#_c_199_n N_A_83_289#_c_206_n N_A_83_289#_c_207_n
+ N_A_83_289#_c_208_n N_A_83_289#_c_209_n N_A_83_289#_c_210_n
+ N_A_83_289#_c_200_n N_A_83_289#_c_201_n PM_SKY130_FD_SC_LS__XOR3_2%A_83_289#
x_PM_SKY130_FD_SC_LS__XOR3_2%A N_A_c_305_n N_A_M1006_g N_A_c_306_n N_A_M1022_g A
+ PM_SKY130_FD_SC_LS__XOR3_2%A
x_PM_SKY130_FD_SC_LS__XOR3_2%A_440_315# N_A_440_315#_M1009_s
+ N_A_440_315#_M1011_s N_A_440_315#_c_351_n N_A_440_315#_c_352_n
+ N_A_440_315#_M1015_g N_A_440_315#_M1008_g N_A_440_315#_c_340_n
+ N_A_440_315#_c_341_n N_A_440_315#_c_355_n N_A_440_315#_M1003_g
+ N_A_440_315#_c_342_n N_A_440_315#_M1020_g N_A_440_315#_c_344_n
+ N_A_440_315#_c_345_n N_A_440_315#_c_346_n N_A_440_315#_c_347_n
+ N_A_440_315#_c_348_n N_A_440_315#_c_349_n N_A_440_315#_c_350_n
+ PM_SKY130_FD_SC_LS__XOR3_2%A_440_315#
x_PM_SKY130_FD_SC_LS__XOR3_2%B N_B_c_465_n N_B_M1012_g N_B_c_466_n N_B_c_467_n
+ N_B_M1019_g N_B_c_453_n N_B_c_454_n N_B_c_468_n N_B_c_469_n N_B_c_470_n
+ N_B_M1021_g N_B_c_471_n N_B_M1016_g N_B_c_456_n N_B_c_457_n N_B_c_458_n
+ N_B_c_459_n N_B_c_460_n N_B_c_461_n N_B_M1011_g N_B_c_462_n N_B_M1009_g
+ N_B_c_474_n N_B_c_463_n B PM_SKY130_FD_SC_LS__XOR3_2%B
x_PM_SKY130_FD_SC_LS__XOR3_2%A_1162_379# N_A_1162_379#_M1018_s
+ N_A_1162_379#_M1010_s N_A_1162_379#_c_589_n N_A_1162_379#_M1013_g
+ N_A_1162_379#_M1004_g N_A_1162_379#_c_590_n N_A_1162_379#_c_591_n
+ N_A_1162_379#_c_592_n N_A_1162_379#_c_593_n N_A_1162_379#_c_594_n
+ N_A_1162_379#_c_595_n N_A_1162_379#_c_584_n N_A_1162_379#_c_585_n
+ N_A_1162_379#_c_586_n N_A_1162_379#_c_587_n N_A_1162_379#_c_588_n
+ PM_SKY130_FD_SC_LS__XOR3_2%A_1162_379#
x_PM_SKY130_FD_SC_LS__XOR3_2%C N_C_c_700_n N_C_c_701_n N_C_M1023_g N_C_c_691_n
+ N_C_M1007_g N_C_c_692_n N_C_c_693_n N_C_c_694_n N_C_c_695_n N_C_M1010_g
+ N_C_c_696_n N_C_c_697_n N_C_c_698_n N_C_M1018_g C PM_SKY130_FD_SC_LS__XOR3_2%C
x_PM_SKY130_FD_SC_LS__XOR3_2%A_1195_424# N_A_1195_424#_M1004_d
+ N_A_1195_424#_M1013_d N_A_1195_424#_c_799_n N_A_1195_424#_M1001_g
+ N_A_1195_424#_M1002_g N_A_1195_424#_c_789_n N_A_1195_424#_c_790_n
+ N_A_1195_424#_M1014_g N_A_1195_424#_c_801_n N_A_1195_424#_M1005_g
+ N_A_1195_424#_c_792_n N_A_1195_424#_c_793_n N_A_1195_424#_c_794_n
+ N_A_1195_424#_c_795_n N_A_1195_424#_c_796_n N_A_1195_424#_c_797_n
+ N_A_1195_424#_c_803_n N_A_1195_424#_c_804_n N_A_1195_424#_c_798_n
+ N_A_1195_424#_c_849_p N_A_1195_424#_c_806_n
+ PM_SKY130_FD_SC_LS__XOR3_2%A_1195_424#
x_PM_SKY130_FD_SC_LS__XOR3_2%A_27_134# N_A_27_134#_M1017_s N_A_27_134#_M1008_d
+ N_A_27_134#_M1000_s N_A_27_134#_M1015_d N_A_27_134#_c_900_n
+ N_A_27_134#_c_901_n N_A_27_134#_c_902_n N_A_27_134#_c_903_n
+ N_A_27_134#_c_904_n N_A_27_134#_c_905_n N_A_27_134#_c_906_n
+ N_A_27_134#_c_907_n N_A_27_134#_c_908_n N_A_27_134#_c_913_n
+ N_A_27_134#_c_909_n N_A_27_134#_c_910_n N_A_27_134#_c_911_n
+ PM_SKY130_FD_SC_LS__XOR3_2%A_27_134#
x_PM_SKY130_FD_SC_LS__XOR3_2%VPWR N_VPWR_M1000_d N_VPWR_M1011_d N_VPWR_M1010_d
+ N_VPWR_M1005_s N_VPWR_c_988_n N_VPWR_c_989_n N_VPWR_c_990_n N_VPWR_c_991_n
+ N_VPWR_c_992_n N_VPWR_c_993_n N_VPWR_c_994_n N_VPWR_c_995_n N_VPWR_c_1038_n
+ VPWR N_VPWR_c_996_n N_VPWR_c_997_n N_VPWR_c_998_n N_VPWR_c_999_n
+ N_VPWR_c_1000_n N_VPWR_c_987_n PM_SKY130_FD_SC_LS__XOR3_2%VPWR
x_PM_SKY130_FD_SC_LS__XOR3_2%A_372_419# N_A_372_419#_M1016_d
+ N_A_372_419#_M1004_s N_A_372_419#_M1012_d N_A_372_419#_M1023_d
+ N_A_372_419#_c_1095_n N_A_372_419#_c_1096_n N_A_372_419#_c_1108_n
+ N_A_372_419#_c_1085_n N_A_372_419#_c_1086_n N_A_372_419#_c_1087_n
+ N_A_372_419#_c_1136_n N_A_372_419#_c_1088_n N_A_372_419#_c_1140_n
+ N_A_372_419#_c_1089_n N_A_372_419#_c_1090_n N_A_372_419#_c_1091_n
+ N_A_372_419#_c_1098_n N_A_372_419#_c_1099_n N_A_372_419#_c_1100_n
+ N_A_372_419#_c_1092_n N_A_372_419#_c_1093_n N_A_372_419#_c_1094_n
+ PM_SKY130_FD_SC_LS__XOR3_2%A_372_419#
x_PM_SKY130_FD_SC_LS__XOR3_2%A_416_113# N_A_416_113#_M1019_d
+ N_A_416_113#_M1007_d N_A_416_113#_M1021_d N_A_416_113#_M1013_s
+ N_A_416_113#_c_1232_n N_A_416_113#_c_1233_n N_A_416_113#_c_1234_n
+ N_A_416_113#_c_1241_n N_A_416_113#_c_1242_n N_A_416_113#_c_1235_n
+ N_A_416_113#_c_1236_n N_A_416_113#_c_1291_n N_A_416_113#_c_1292_n
+ N_A_416_113#_c_1237_n N_A_416_113#_c_1238_n N_A_416_113#_c_1243_n
+ N_A_416_113#_c_1261_n N_A_416_113#_c_1244_n N_A_416_113#_c_1245_n
+ N_A_416_113#_c_1246_n N_A_416_113#_c_1239_n N_A_416_113#_c_1240_n
+ PM_SKY130_FD_SC_LS__XOR3_2%A_416_113#
x_PM_SKY130_FD_SC_LS__XOR3_2%X N_X_M1002_s N_X_M1001_d X X X X X X X
+ PM_SKY130_FD_SC_LS__XOR3_2%X
x_PM_SKY130_FD_SC_LS__XOR3_2%VGND N_VGND_M1017_d N_VGND_M1009_d N_VGND_M1018_d
+ N_VGND_M1014_d N_VGND_c_1378_n N_VGND_c_1379_n N_VGND_c_1380_n N_VGND_c_1381_n
+ VGND N_VGND_c_1382_n N_VGND_c_1383_n N_VGND_c_1384_n N_VGND_c_1385_n
+ N_VGND_c_1386_n N_VGND_c_1387_n N_VGND_c_1388_n N_VGND_c_1389_n
+ PM_SKY130_FD_SC_LS__XOR3_2%VGND
cc_1 VNB N_A_83_289#_M1017_g 0.025899f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.99
cc_2 VNB N_A_83_289#_c_197_n 0.0213533f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.86
cc_3 VNB N_A_83_289#_c_198_n 0.00288335f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.61
cc_4 VNB N_A_83_289#_c_199_n 0.00787075f $X=-0.19 $Y=-0.245 $X2=1.54 $Y2=1.165
cc_5 VNB N_A_83_289#_c_200_n 0.00297214f $X=-0.19 $Y=-0.245 $X2=4.06 $Y2=1.905
cc_6 VNB N_A_83_289#_c_201_n 8.48484e-19 $X=-0.19 $Y=-0.245 $X2=4.31 $Y2=1.1
cc_7 VNB N_A_c_305_n 0.0296327f $X=-0.19 $Y=-0.245 $X2=1.4 $Y2=0.67
cc_8 VNB N_A_c_306_n 0.0210019f $X=-0.19 $Y=-0.245 $X2=3.35 $Y2=1.895
cc_9 VNB A 0.00137659f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_440_315#_M1008_g 0.0365935f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.99
cc_11 VNB N_A_440_315#_c_340_n 0.0212262f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_440_315#_c_341_n 0.0123579f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.86
cc_13 VNB N_A_440_315#_c_342_n 0.0108329f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.61
cc_14 VNB N_A_440_315#_M1020_g 0.0193825f $X=-0.19 $Y=-0.245 $X2=1.31 $Y2=2.005
cc_15 VNB N_A_440_315#_c_344_n 0.00889208f $X=-0.19 $Y=-0.245 $X2=1.475 $Y2=2.24
cc_16 VNB N_A_440_315#_c_345_n 0.00122356f $X=-0.19 $Y=-0.245 $X2=1.54 $Y2=1.165
cc_17 VNB N_A_440_315#_c_346_n 0.00935992f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_440_315#_c_347_n 3.26207e-19 $X=-0.19 $Y=-0.245 $X2=3.725 $Y2=2.99
cc_19 VNB N_A_440_315#_c_348_n 0.0065592f $X=-0.19 $Y=-0.245 $X2=3.81 $Y2=2.905
cc_20 VNB N_A_440_315#_c_349_n 0.00140635f $X=-0.19 $Y=-0.245 $X2=4.06 $Y2=2.755
cc_21 VNB N_A_440_315#_c_350_n 0.024011f $X=-0.19 $Y=-0.245 $X2=4.15 $Y2=1.1
cc_22 VNB N_B_M1019_g 0.0412954f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_B_c_453_n 0.0694559f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_B_c_454_n 0.012806f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_B_M1016_g 0.0335493f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.61
cc_26 VNB N_B_c_456_n 0.089017f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.61
cc_27 VNB N_B_c_457_n 0.0180259f $X=-0.19 $Y=-0.245 $X2=1.31 $Y2=2.005
cc_28 VNB N_B_c_458_n 0.00660556f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=2.005
cc_29 VNB N_B_c_459_n 0.0579081f $X=-0.19 $Y=-0.245 $X2=1.475 $Y2=2.905
cc_30 VNB N_B_c_460_n 0.0190806f $X=-0.19 $Y=-0.245 $X2=1.475 $Y2=2.24
cc_31 VNB N_B_c_461_n 0.0504682f $X=-0.19 $Y=-0.245 $X2=1.54 $Y2=1.92
cc_32 VNB N_B_c_462_n 0.0199242f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_B_c_463_n 0.00749069f $X=-0.19 $Y=-0.245 $X2=3.81 $Y2=2.905
cc_34 VNB B 0.0062914f $X=-0.19 $Y=-0.245 $X2=4.31 $Y2=1.905
cc_35 VNB N_A_1162_379#_M1004_g 0.0259339f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_1162_379#_c_584_n 4.38491e-19 $X=-0.19 $Y=-0.245 $X2=1.475
+ $Y2=2.09
cc_37 VNB N_A_1162_379#_c_585_n 0.00454486f $X=-0.19 $Y=-0.245 $X2=1.475
+ $Y2=2.905
cc_38 VNB N_A_1162_379#_c_586_n 0.00752181f $X=-0.19 $Y=-0.245 $X2=1.475
+ $Y2=2.24
cc_39 VNB N_A_1162_379#_c_587_n 0.00213207f $X=-0.19 $Y=-0.245 $X2=1.54
+ $Y2=1.165
cc_40 VNB N_A_1162_379#_c_588_n 0.034674f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_C_c_691_n 0.0206136f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_C_c_692_n 0.0352899f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_C_c_693_n 0.0359362f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_C_c_694_n 0.0206211f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_C_c_695_n 0.0145784f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.445
cc_46 VNB N_C_c_696_n 0.027196f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_C_c_697_n 0.011937f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.86
cc_48 VNB N_C_c_698_n 0.0174959f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=2.435
cc_49 VNB C 7.99339e-19 $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.61
cc_50 VNB N_A_1195_424#_M1002_g 0.0221192f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_1195_424#_c_789_n 0.00970685f $X=-0.19 $Y=-0.245 $X2=0.495
+ $Y2=0.99
cc_52 VNB N_A_1195_424#_c_790_n 0.0151082f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.86
cc_53 VNB N_A_1195_424#_M1014_g 0.0248256f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.92
cc_54 VNB N_A_1195_424#_c_792_n 0.0413116f $X=-0.19 $Y=-0.245 $X2=1.31 $Y2=2.005
cc_55 VNB N_A_1195_424#_c_793_n 0.0105781f $X=-0.19 $Y=-0.245 $X2=0.745
+ $Y2=2.005
cc_56 VNB N_A_1195_424#_c_794_n 0.0124983f $X=-0.19 $Y=-0.245 $X2=1.475 $Y2=2.09
cc_57 VNB N_A_1195_424#_c_795_n 0.00243198f $X=-0.19 $Y=-0.245 $X2=1.475
+ $Y2=2.24
cc_58 VNB N_A_1195_424#_c_796_n 0.00555163f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_1195_424#_c_797_n 0.00493017f $X=-0.19 $Y=-0.245 $X2=3.81
+ $Y2=2.755
cc_60 VNB N_A_1195_424#_c_798_n 0.0010115f $X=-0.19 $Y=-0.245 $X2=4.06 $Y2=2.755
cc_61 VNB N_A_27_134#_c_900_n 0.0122262f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.445
cc_62 VNB N_A_27_134#_c_901_n 0.0103833f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.99
cc_63 VNB N_A_27_134#_c_902_n 0.00553396f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.86
cc_64 VNB N_A_27_134#_c_903_n 0.00184736f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.92
cc_65 VNB N_A_27_134#_c_904_n 0.011717f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.61
cc_66 VNB N_A_27_134#_c_905_n 0.00394375f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.61
cc_67 VNB N_A_27_134#_c_906_n 4.4909e-19 $X=-0.19 $Y=-0.245 $X2=1.31 $Y2=2.005
cc_68 VNB N_A_27_134#_c_907_n 0.00200956f $X=-0.19 $Y=-0.245 $X2=1.475 $Y2=2.905
cc_69 VNB N_A_27_134#_c_908_n 0.00710642f $X=-0.19 $Y=-0.245 $X2=1.54 $Y2=1.92
cc_70 VNB N_A_27_134#_c_909_n 0.0180441f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_27_134#_c_910_n 0.0054336f $X=-0.19 $Y=-0.245 $X2=1.64 $Y2=2.99
cc_72 VNB N_A_27_134#_c_911_n 0.00346141f $X=-0.19 $Y=-0.245 $X2=4.31 $Y2=1.905
cc_73 VNB N_VPWR_c_987_n 0.40251f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_372_419#_c_1085_n 0.00979392f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.61
cc_75 VNB N_A_372_419#_c_1086_n 0.021596f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.61
cc_76 VNB N_A_372_419#_c_1087_n 0.00289389f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_372_419#_c_1088_n 0.00673931f $X=-0.19 $Y=-0.245 $X2=1.475
+ $Y2=2.09
cc_78 VNB N_A_372_419#_c_1089_n 0.00540474f $X=-0.19 $Y=-0.245 $X2=1.475
+ $Y2=2.24
cc_79 VNB N_A_372_419#_c_1090_n 0.0332271f $X=-0.19 $Y=-0.245 $X2=1.54 $Y2=1.92
cc_80 VNB N_A_372_419#_c_1091_n 0.00432252f $X=-0.19 $Y=-0.245 $X2=1.54
+ $Y2=1.165
cc_81 VNB N_A_372_419#_c_1092_n 0.00361673f $X=-0.19 $Y=-0.245 $X2=4.31
+ $Y2=1.905
cc_82 VNB N_A_372_419#_c_1093_n 0.0166275f $X=-0.19 $Y=-0.245 $X2=4.06 $Y2=2.07
cc_83 VNB N_A_372_419#_c_1094_n 0.00844405f $X=-0.19 $Y=-0.245 $X2=4.15 $Y2=1.1
cc_84 VNB N_A_416_113#_c_1232_n 0.00163083f $X=-0.19 $Y=-0.245 $X2=0.495
+ $Y2=0.99
cc_85 VNB N_A_416_113#_c_1233_n 0.0128498f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.86
cc_86 VNB N_A_416_113#_c_1234_n 0.00351336f $X=-0.19 $Y=-0.245 $X2=0.655
+ $Y2=2.435
cc_87 VNB N_A_416_113#_c_1235_n 0.0141251f $X=-0.19 $Y=-0.245 $X2=1.54 $Y2=1.92
cc_88 VNB N_A_416_113#_c_1236_n 0.00344537f $X=-0.19 $Y=-0.245 $X2=1.54
+ $Y2=1.165
cc_89 VNB N_A_416_113#_c_1237_n 0.00643748f $X=-0.19 $Y=-0.245 $X2=3.81
+ $Y2=2.905
cc_90 VNB N_A_416_113#_c_1238_n 0.00230384f $X=-0.19 $Y=-0.245 $X2=4.31
+ $Y2=1.265
cc_91 VNB N_A_416_113#_c_1239_n 0.00505131f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_416_113#_c_1240_n 0.0107302f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB X 0.00248472f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_VGND_c_1378_n 0.00766793f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.99
cc_95 VNB N_VGND_c_1379_n 0.0157044f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=2.435
cc_96 VNB N_VGND_c_1380_n 0.011316f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.61
cc_97 VNB N_VGND_c_1381_n 0.0467556f $X=-0.19 $Y=-0.245 $X2=1.31 $Y2=2.005
cc_98 VNB N_VGND_c_1382_n 0.102977f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_VGND_c_1383_n 0.0640359f $X=-0.19 $Y=-0.245 $X2=4.06 $Y2=2.07
cc_100 VNB N_VGND_c_1384_n 0.0191116f $X=-0.19 $Y=-0.245 $X2=4.15 $Y2=1.1
cc_101 VNB N_VGND_c_1385_n 0.0197198f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_VGND_c_1386_n 0.037346f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_VGND_c_1387_n 0.00477918f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_VGND_c_1388_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_VGND_c_1389_n 0.506431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VPB N_A_83_289#_c_197_n 0.0395778f $X=-0.19 $Y=1.66 $X2=0.655 $Y2=1.86
cc_107 VPB N_A_83_289#_c_198_n 0.00210455f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=1.61
cc_108 VPB N_A_83_289#_c_204_n 0.0085376f $X=-0.19 $Y=1.66 $X2=1.31 $Y2=2.005
cc_109 VPB N_A_83_289#_c_199_n 0.00690601f $X=-0.19 $Y=1.66 $X2=1.54 $Y2=1.165
cc_110 VPB N_A_83_289#_c_206_n 0.0344474f $X=-0.19 $Y=1.66 $X2=3.725 $Y2=2.99
cc_111 VPB N_A_83_289#_c_207_n 0.00255622f $X=-0.19 $Y=1.66 $X2=1.64 $Y2=2.99
cc_112 VPB N_A_83_289#_c_208_n 0.00523651f $X=-0.19 $Y=1.66 $X2=3.81 $Y2=2.905
cc_113 VPB N_A_83_289#_c_209_n 0.00581926f $X=-0.19 $Y=1.66 $X2=1.31 $Y2=1.92
cc_114 VPB N_A_83_289#_c_210_n 0.0104124f $X=-0.19 $Y=1.66 $X2=3.81 $Y2=2.07
cc_115 VPB N_A_83_289#_c_200_n 0.00329913f $X=-0.19 $Y=1.66 $X2=4.06 $Y2=1.905
cc_116 VPB N_A_c_305_n 0.0390865f $X=-0.19 $Y=1.66 $X2=1.4 $Y2=0.67
cc_117 VPB A 0.00190989f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_A_440_315#_c_351_n 0.0158328f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_A_440_315#_c_352_n 0.0203838f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_A_440_315#_c_340_n 0.019913f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_A_440_315#_c_341_n 0.0106007f $X=-0.19 $Y=1.66 $X2=0.655 $Y2=1.86
cc_122 VPB N_A_440_315#_c_355_n 0.0156457f $X=-0.19 $Y=1.66 $X2=0.655 $Y2=2.435
cc_123 VPB N_A_440_315#_c_342_n 0.0127697f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.61
cc_124 VPB N_A_440_315#_c_344_n 0.00873141f $X=-0.19 $Y=1.66 $X2=1.475 $Y2=2.24
cc_125 VPB N_A_440_315#_c_348_n 0.00564133f $X=-0.19 $Y=1.66 $X2=3.81 $Y2=2.905
cc_126 VPB N_A_440_315#_c_349_n 4.64599e-19 $X=-0.19 $Y=1.66 $X2=4.06 $Y2=2.755
cc_127 VPB N_A_440_315#_c_350_n 0.0135441f $X=-0.19 $Y=1.66 $X2=4.15 $Y2=1.1
cc_128 VPB N_B_c_465_n 0.0188478f $X=-0.19 $Y=1.66 $X2=1.4 $Y2=0.67
cc_129 VPB N_B_c_466_n 0.0540201f $X=-0.19 $Y=1.66 $X2=3.35 $Y2=1.895
cc_130 VPB N_B_c_467_n 0.019206f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_B_c_468_n 0.00809905f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_B_c_469_n 0.0134034f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.445
cc_133 VPB N_B_c_470_n 0.0137131f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.99
cc_134 VPB N_B_c_471_n 0.113935f $X=-0.19 $Y=1.66 $X2=0.655 $Y2=1.86
cc_135 VPB N_B_c_458_n 0.0893728f $X=-0.19 $Y=1.66 $X2=0.745 $Y2=2.005
cc_136 VPB N_B_c_461_n 0.0263968f $X=-0.19 $Y=1.66 $X2=1.54 $Y2=1.92
cc_137 VPB N_B_c_474_n 0.0089864f $X=-0.19 $Y=1.66 $X2=3.81 $Y2=2.755
cc_138 VPB N_A_1162_379#_c_589_n 0.0200244f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_A_1162_379#_c_590_n 0.00869713f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.99
cc_140 VPB N_A_1162_379#_c_591_n 0.0289022f $X=-0.19 $Y=1.66 $X2=0.655 $Y2=2.435
cc_141 VPB N_A_1162_379#_c_592_n 0.00327735f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.61
cc_142 VPB N_A_1162_379#_c_593_n 0.0227054f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=1.61
cc_143 VPB N_A_1162_379#_c_594_n 0.00305237f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=1.61
cc_144 VPB N_A_1162_379#_c_595_n 0.0127293f $X=-0.19 $Y=1.66 $X2=1.31 $Y2=2.005
cc_145 VPB N_A_1162_379#_c_584_n 0.00915273f $X=-0.19 $Y=1.66 $X2=1.475 $Y2=2.09
cc_146 VPB N_A_1162_379#_c_587_n 0.00170428f $X=-0.19 $Y=1.66 $X2=1.54 $Y2=1.165
cc_147 VPB N_A_1162_379#_c_588_n 0.0044609f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_148 VPB N_C_c_700_n 0.0164618f $X=-0.19 $Y=1.66 $X2=3.84 $Y2=0.625
cc_149 VPB N_C_c_701_n 0.0261652f $X=-0.19 $Y=1.66 $X2=1.325 $Y2=1.935
cc_150 VPB N_C_c_693_n 0.0137087f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_151 VPB N_C_c_695_n 0.0276861f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.445
cc_152 VPB C 0.00197916f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=1.61
cc_153 VPB N_A_1195_424#_c_799_n 0.0160231f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_154 VPB N_A_1195_424#_c_790_n 0.00111912f $X=-0.19 $Y=1.66 $X2=0.655 $Y2=1.86
cc_155 VPB N_A_1195_424#_c_801_n 0.0258458f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=1.61
cc_156 VPB N_A_1195_424#_c_793_n 0.00769406f $X=-0.19 $Y=1.66 $X2=0.745
+ $Y2=2.005
cc_157 VPB N_A_1195_424#_c_803_n 0.0106241f $X=-0.19 $Y=1.66 $X2=1.31 $Y2=1.92
cc_158 VPB N_A_1195_424#_c_804_n 0.00211174f $X=-0.19 $Y=1.66 $X2=4.06 $Y2=2.07
cc_159 VPB N_A_1195_424#_c_798_n 0.00275279f $X=-0.19 $Y=1.66 $X2=4.06 $Y2=2.755
cc_160 VPB N_A_1195_424#_c_806_n 0.0029919f $X=-0.19 $Y=1.66 $X2=4.31 $Y2=1.1
cc_161 VPB N_A_27_134#_c_906_n 0.00208841f $X=-0.19 $Y=1.66 $X2=1.31 $Y2=2.005
cc_162 VPB N_A_27_134#_c_913_n 0.0381571f $X=-0.19 $Y=1.66 $X2=1.54 $Y2=1.165
cc_163 VPB N_A_27_134#_c_909_n 0.0285695f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_164 VPB N_VPWR_c_988_n 0.0107656f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.99
cc_165 VPB N_VPWR_c_989_n 0.00834949f $X=-0.19 $Y=1.66 $X2=0.655 $Y2=2.435
cc_166 VPB N_VPWR_c_990_n 0.00566488f $X=-0.19 $Y=1.66 $X2=1.31 $Y2=2.005
cc_167 VPB N_VPWR_c_991_n 0.0132563f $X=-0.19 $Y=1.66 $X2=1.475 $Y2=2.905
cc_168 VPB N_VPWR_c_992_n 0.0106521f $X=-0.19 $Y=1.66 $X2=1.475 $Y2=2.24
cc_169 VPB N_VPWR_c_993_n 0.0592421f $X=-0.19 $Y=1.66 $X2=1.54 $Y2=1.92
cc_170 VPB N_VPWR_c_994_n 0.0227085f $X=-0.19 $Y=1.66 $X2=1.64 $Y2=2.99
cc_171 VPB N_VPWR_c_995_n 0.00632158f $X=-0.19 $Y=1.66 $X2=3.81 $Y2=2.755
cc_172 VPB N_VPWR_c_996_n 0.0940373f $X=-0.19 $Y=1.66 $X2=4.15 $Y2=1.1
cc_173 VPB N_VPWR_c_997_n 0.0711821f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_174 VPB N_VPWR_c_998_n 0.0198086f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_175 VPB N_VPWR_c_999_n 0.00460249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_176 VPB N_VPWR_c_1000_n 0.0106494f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_177 VPB N_VPWR_c_987_n 0.112692f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_178 VPB N_A_372_419#_c_1095_n 0.00501008f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.99
cc_179 VPB N_A_372_419#_c_1096_n 8.77792e-19 $X=-0.19 $Y=1.66 $X2=0.655 $Y2=1.86
cc_180 VPB N_A_372_419#_c_1085_n 0.00371521f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=1.61
cc_181 VPB N_A_372_419#_c_1098_n 0.00795012f $X=-0.19 $Y=1.66 $X2=3.725 $Y2=2.99
cc_182 VPB N_A_372_419#_c_1099_n 0.00674591f $X=-0.19 $Y=1.66 $X2=3.81 $Y2=2.755
cc_183 VPB N_A_372_419#_c_1100_n 0.00450367f $X=-0.19 $Y=1.66 $X2=3.81 $Y2=2.905
cc_184 VPB N_A_372_419#_c_1092_n 0.00442062f $X=-0.19 $Y=1.66 $X2=4.31 $Y2=1.905
cc_185 VPB N_A_416_113#_c_1241_n 3.7394e-19 $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.61
cc_186 VPB N_A_416_113#_c_1242_n 0.013813f $X=-0.19 $Y=1.66 $X2=1.475 $Y2=2.09
cc_187 VPB N_A_416_113#_c_1243_n 0.011909f $X=-0.19 $Y=1.66 $X2=1.31 $Y2=1.92
cc_188 VPB N_A_416_113#_c_1244_n 0.00298342f $X=-0.19 $Y=1.66 $X2=4.06 $Y2=2.755
cc_189 VPB N_A_416_113#_c_1245_n 0.00684386f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_190 VPB N_A_416_113#_c_1246_n 0.00925538f $X=-0.19 $Y=1.66 $X2=4.31 $Y2=1.1
cc_191 VPB N_A_416_113#_c_1239_n 0.00151514f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_192 VPB N_A_416_113#_c_1240_n 0.00700164f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_193 VPB X 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_194 N_A_83_289#_M1017_g N_A_c_305_n 8.70324e-19 $X=0.495 $Y=0.99 $X2=-0.19
+ $Y2=-0.245
cc_195 N_A_83_289#_c_197_n N_A_c_305_n 0.0465276f $X=0.655 $Y=1.86 $X2=-0.19
+ $Y2=-0.245
cc_196 N_A_83_289#_c_198_n N_A_c_305_n 0.00284697f $X=0.58 $Y=1.61 $X2=-0.19
+ $Y2=-0.245
cc_197 N_A_83_289#_c_204_n N_A_c_305_n 0.0152386f $X=1.31 $Y=2.005 $X2=-0.19
+ $Y2=-0.245
cc_198 N_A_83_289#_c_216_p N_A_c_305_n 0.0123706f $X=1.475 $Y=2.24 $X2=-0.19
+ $Y2=-0.245
cc_199 N_A_83_289#_c_199_n N_A_c_305_n 0.00619098f $X=1.54 $Y=1.165 $X2=-0.19
+ $Y2=-0.245
cc_200 N_A_83_289#_c_207_n N_A_c_305_n 0.00384879f $X=1.64 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_201 N_A_83_289#_c_209_n N_A_c_305_n 0.00665162f $X=1.31 $Y=1.92 $X2=-0.19
+ $Y2=-0.245
cc_202 N_A_83_289#_M1017_g N_A_c_306_n 0.0147663f $X=0.495 $Y=0.99 $X2=0 $Y2=0
cc_203 N_A_83_289#_c_199_n N_A_c_306_n 0.0111091f $X=1.54 $Y=1.165 $X2=0 $Y2=0
cc_204 N_A_83_289#_M1017_g A 0.00405976f $X=0.495 $Y=0.99 $X2=0 $Y2=0
cc_205 N_A_83_289#_c_197_n A 0.00106229f $X=0.655 $Y=1.86 $X2=0 $Y2=0
cc_206 N_A_83_289#_c_198_n A 0.0192835f $X=0.58 $Y=1.61 $X2=0 $Y2=0
cc_207 N_A_83_289#_c_204_n A 0.0254385f $X=1.31 $Y=2.005 $X2=0 $Y2=0
cc_208 N_A_83_289#_c_199_n A 0.0378672f $X=1.54 $Y=1.165 $X2=0 $Y2=0
cc_209 N_A_83_289#_c_209_n N_A_440_315#_c_351_n 0.00133418f $X=1.31 $Y=1.92
+ $X2=0 $Y2=0
cc_210 N_A_83_289#_c_206_n N_A_440_315#_c_352_n 0.00115048f $X=3.725 $Y=2.99
+ $X2=0 $Y2=0
cc_211 N_A_83_289#_c_199_n N_A_440_315#_c_341_n 0.00853359f $X=1.54 $Y=1.165
+ $X2=0 $Y2=0
cc_212 N_A_83_289#_c_206_n N_A_440_315#_c_355_n 0.00115048f $X=3.725 $Y=2.99
+ $X2=0 $Y2=0
cc_213 N_A_83_289#_c_210_n N_A_440_315#_c_355_n 0.0057628f $X=3.81 $Y=2.07 $X2=0
+ $Y2=0
cc_214 N_A_83_289#_c_200_n N_A_440_315#_M1020_g 4.86955e-19 $X=4.06 $Y=1.905
+ $X2=0 $Y2=0
cc_215 N_A_83_289#_c_201_n N_A_440_315#_M1020_g 0.00119421f $X=4.31 $Y=1.1 $X2=0
+ $Y2=0
cc_216 N_A_83_289#_c_200_n N_A_440_315#_c_345_n 0.00794453f $X=4.06 $Y=1.905
+ $X2=0 $Y2=0
cc_217 N_A_83_289#_M1020_d N_A_440_315#_c_346_n 0.0066978f $X=3.84 $Y=0.625
+ $X2=0 $Y2=0
cc_218 N_A_83_289#_c_201_n N_A_440_315#_c_346_n 0.0483684f $X=4.31 $Y=1.1 $X2=0
+ $Y2=0
cc_219 N_A_83_289#_c_200_n N_A_440_315#_c_348_n 0.102962f $X=4.06 $Y=1.905 $X2=0
+ $Y2=0
cc_220 N_A_83_289#_c_210_n N_A_440_315#_c_349_n 0.0250643f $X=3.81 $Y=2.07 $X2=0
+ $Y2=0
cc_221 N_A_83_289#_c_200_n N_A_440_315#_c_349_n 0.0225071f $X=4.06 $Y=1.905
+ $X2=0 $Y2=0
cc_222 N_A_83_289#_c_210_n N_A_440_315#_c_350_n 0.00811391f $X=3.81 $Y=2.07
+ $X2=0 $Y2=0
cc_223 N_A_83_289#_c_200_n N_A_440_315#_c_350_n 0.00113401f $X=4.06 $Y=1.905
+ $X2=0 $Y2=0
cc_224 N_A_83_289#_c_216_p N_B_c_465_n 0.0106287f $X=1.475 $Y=2.24 $X2=-0.19
+ $Y2=-0.245
cc_225 N_A_83_289#_c_206_n N_B_c_465_n 0.0118001f $X=3.725 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_226 N_A_83_289#_c_209_n N_B_c_465_n 0.00364241f $X=1.31 $Y=1.92 $X2=-0.19
+ $Y2=-0.245
cc_227 N_A_83_289#_c_206_n N_B_c_466_n 0.0156543f $X=3.725 $Y=2.99 $X2=0 $Y2=0
cc_228 N_A_83_289#_c_206_n N_B_c_467_n 0.00566576f $X=3.725 $Y=2.99 $X2=0 $Y2=0
cc_229 N_A_83_289#_c_199_n N_B_M1019_g 9.19484e-19 $X=1.54 $Y=1.165 $X2=0 $Y2=0
cc_230 N_A_83_289#_c_206_n N_B_c_469_n 0.014816f $X=3.725 $Y=2.99 $X2=0 $Y2=0
cc_231 N_A_83_289#_c_206_n N_B_c_471_n 0.0205994f $X=3.725 $Y=2.99 $X2=0 $Y2=0
cc_232 N_A_83_289#_c_210_n N_B_c_471_n 0.00629714f $X=3.81 $Y=2.07 $X2=0 $Y2=0
cc_233 N_A_83_289#_c_200_n N_B_c_457_n 0.0075973f $X=4.06 $Y=1.905 $X2=0 $Y2=0
cc_234 N_A_83_289#_c_201_n N_B_c_457_n 0.00195237f $X=4.31 $Y=1.1 $X2=0 $Y2=0
cc_235 N_A_83_289#_c_206_n N_B_c_458_n 0.00546456f $X=3.725 $Y=2.99 $X2=0 $Y2=0
cc_236 N_A_83_289#_c_208_n N_B_c_458_n 0.00399845f $X=3.81 $Y=2.905 $X2=0 $Y2=0
cc_237 N_A_83_289#_c_210_n N_B_c_458_n 0.0344517f $X=3.81 $Y=2.07 $X2=0 $Y2=0
cc_238 N_A_83_289#_c_200_n N_B_c_458_n 0.00951175f $X=4.06 $Y=1.905 $X2=0 $Y2=0
cc_239 N_A_83_289#_c_201_n N_B_c_459_n 0.00788621f $X=4.31 $Y=1.1 $X2=0 $Y2=0
cc_240 N_A_83_289#_c_258_p N_A_27_134#_M1000_s 0.00279118f $X=0.745 $Y=2.005
+ $X2=0 $Y2=0
cc_241 N_A_83_289#_M1017_g N_A_27_134#_c_900_n 0.00162247f $X=0.495 $Y=0.99
+ $X2=0 $Y2=0
cc_242 N_A_83_289#_M1017_g N_A_27_134#_c_901_n 0.0115093f $X=0.495 $Y=0.99 $X2=0
+ $Y2=0
cc_243 N_A_83_289#_M1022_d N_A_27_134#_c_902_n 0.0132999f $X=1.4 $Y=0.67 $X2=0
+ $Y2=0
cc_244 N_A_83_289#_M1017_g N_A_27_134#_c_902_n 0.0109735f $X=0.495 $Y=0.99 $X2=0
+ $Y2=0
cc_245 N_A_83_289#_c_197_n N_A_27_134#_c_902_n 6.88341e-19 $X=0.655 $Y=1.86
+ $X2=0 $Y2=0
cc_246 N_A_83_289#_c_198_n N_A_27_134#_c_902_n 0.00736351f $X=0.58 $Y=1.61 $X2=0
+ $Y2=0
cc_247 N_A_83_289#_c_199_n N_A_27_134#_c_902_n 0.0135869f $X=1.54 $Y=1.165 $X2=0
+ $Y2=0
cc_248 N_A_83_289#_M1022_d N_A_27_134#_c_903_n 0.00424046f $X=1.4 $Y=0.67 $X2=0
+ $Y2=0
cc_249 N_A_83_289#_c_199_n N_A_27_134#_c_903_n 0.0290186f $X=1.54 $Y=1.165 $X2=0
+ $Y2=0
cc_250 N_A_83_289#_c_199_n N_A_27_134#_c_905_n 0.0143578f $X=1.54 $Y=1.165 $X2=0
+ $Y2=0
cc_251 N_A_83_289#_M1017_g N_A_27_134#_c_908_n 0.00602985f $X=0.495 $Y=0.99
+ $X2=0 $Y2=0
cc_252 N_A_83_289#_c_198_n N_A_27_134#_c_908_n 0.0015079f $X=0.58 $Y=1.61 $X2=0
+ $Y2=0
cc_253 N_A_83_289#_c_197_n N_A_27_134#_c_913_n 0.00830772f $X=0.655 $Y=1.86
+ $X2=0 $Y2=0
cc_254 N_A_83_289#_c_258_p N_A_27_134#_c_913_n 0.0099559f $X=0.745 $Y=2.005
+ $X2=0 $Y2=0
cc_255 N_A_83_289#_M1017_g N_A_27_134#_c_909_n 0.00411368f $X=0.495 $Y=0.99
+ $X2=0 $Y2=0
cc_256 N_A_83_289#_c_197_n N_A_27_134#_c_909_n 0.0125302f $X=0.655 $Y=1.86 $X2=0
+ $Y2=0
cc_257 N_A_83_289#_c_198_n N_A_27_134#_c_909_n 0.0361694f $X=0.58 $Y=1.61 $X2=0
+ $Y2=0
cc_258 N_A_83_289#_c_258_p N_A_27_134#_c_909_n 0.0140831f $X=0.745 $Y=2.005
+ $X2=0 $Y2=0
cc_259 N_A_83_289#_c_204_n N_VPWR_M1000_d 0.00482237f $X=1.31 $Y=2.005 $X2=-0.19
+ $Y2=-0.245
cc_260 N_A_83_289#_c_197_n N_VPWR_c_988_n 0.00786945f $X=0.655 $Y=1.86 $X2=0
+ $Y2=0
cc_261 N_A_83_289#_c_204_n N_VPWR_c_988_n 0.0249771f $X=1.31 $Y=2.005 $X2=0
+ $Y2=0
cc_262 N_A_83_289#_c_216_p N_VPWR_c_988_n 0.0417669f $X=1.475 $Y=2.24 $X2=0
+ $Y2=0
cc_263 N_A_83_289#_c_207_n N_VPWR_c_988_n 0.0119463f $X=1.64 $Y=2.99 $X2=0 $Y2=0
cc_264 N_A_83_289#_c_197_n N_VPWR_c_994_n 0.00544739f $X=0.655 $Y=1.86 $X2=0
+ $Y2=0
cc_265 N_A_83_289#_c_206_n N_VPWR_c_996_n 0.144761f $X=3.725 $Y=2.99 $X2=0 $Y2=0
cc_266 N_A_83_289#_c_207_n N_VPWR_c_996_n 0.0236566f $X=1.64 $Y=2.99 $X2=0 $Y2=0
cc_267 N_A_83_289#_c_210_n N_VPWR_c_996_n 0.0112583f $X=3.81 $Y=2.07 $X2=0 $Y2=0
cc_268 N_A_83_289#_c_197_n N_VPWR_c_987_n 0.00537853f $X=0.655 $Y=1.86 $X2=0
+ $Y2=0
cc_269 N_A_83_289#_c_206_n N_VPWR_c_987_n 0.0758332f $X=3.725 $Y=2.99 $X2=0
+ $Y2=0
cc_270 N_A_83_289#_c_207_n N_VPWR_c_987_n 0.0128296f $X=1.64 $Y=2.99 $X2=0 $Y2=0
cc_271 N_A_83_289#_c_210_n N_VPWR_c_987_n 0.01371f $X=3.81 $Y=2.07 $X2=0 $Y2=0
cc_272 N_A_83_289#_c_206_n N_A_372_419#_M1012_d 0.00229245f $X=3.725 $Y=2.99
+ $X2=0 $Y2=0
cc_273 N_A_83_289#_c_216_p N_A_372_419#_c_1095_n 0.0312812f $X=1.475 $Y=2.24
+ $X2=0 $Y2=0
cc_274 N_A_83_289#_c_209_n N_A_372_419#_c_1095_n 0.00107943f $X=1.31 $Y=1.92
+ $X2=0 $Y2=0
cc_275 N_A_83_289#_M1003_d N_A_372_419#_c_1096_n 0.00343339f $X=3.35 $Y=1.895
+ $X2=0 $Y2=0
cc_276 N_A_83_289#_c_206_n N_A_372_419#_c_1096_n 0.0850674f $X=3.725 $Y=2.99
+ $X2=0 $Y2=0
cc_277 N_A_83_289#_c_210_n N_A_372_419#_c_1096_n 0.0152397f $X=3.81 $Y=2.07
+ $X2=0 $Y2=0
cc_278 N_A_83_289#_c_216_p N_A_372_419#_c_1108_n 0.0118923f $X=1.475 $Y=2.24
+ $X2=0 $Y2=0
cc_279 N_A_83_289#_c_206_n N_A_372_419#_c_1108_n 0.0198506f $X=3.725 $Y=2.99
+ $X2=0 $Y2=0
cc_280 N_A_83_289#_M1003_d N_A_372_419#_c_1085_n 0.0105509f $X=3.35 $Y=1.895
+ $X2=0 $Y2=0
cc_281 N_A_83_289#_c_210_n N_A_372_419#_c_1085_n 0.0514618f $X=3.81 $Y=2.07
+ $X2=0 $Y2=0
cc_282 N_A_83_289#_c_200_n N_A_372_419#_c_1085_n 0.00493854f $X=4.06 $Y=1.905
+ $X2=0 $Y2=0
cc_283 N_A_83_289#_M1003_d N_A_416_113#_c_1243_n 0.0102411f $X=3.35 $Y=1.895
+ $X2=0 $Y2=0
cc_284 N_A_83_289#_c_210_n N_A_416_113#_c_1243_n 0.0691818f $X=3.81 $Y=2.07
+ $X2=0 $Y2=0
cc_285 N_A_83_289#_M1017_g N_VGND_c_1385_n 0.00305419f $X=0.495 $Y=0.99 $X2=0
+ $Y2=0
cc_286 N_A_83_289#_M1017_g N_VGND_c_1389_n 0.00457172f $X=0.495 $Y=0.99 $X2=0
+ $Y2=0
cc_287 N_A_c_305_n N_B_c_465_n 0.0163966f $X=1.25 $Y=1.86 $X2=-0.19 $Y2=-0.245
cc_288 N_A_c_305_n N_B_c_467_n 0.0017072f $X=1.25 $Y=1.86 $X2=0 $Y2=0
cc_289 N_A_c_306_n N_B_M1019_g 0.0120059f $X=1.325 $Y=1.42 $X2=0 $Y2=0
cc_290 N_A_c_305_n N_A_27_134#_c_902_n 0.00104511f $X=1.25 $Y=1.86 $X2=0 $Y2=0
cc_291 N_A_c_306_n N_A_27_134#_c_902_n 0.0172797f $X=1.325 $Y=1.42 $X2=0 $Y2=0
cc_292 A N_A_27_134#_c_902_n 0.01258f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_293 N_A_c_306_n N_A_27_134#_c_903_n 0.00341356f $X=1.325 $Y=1.42 $X2=0 $Y2=0
cc_294 A N_A_27_134#_c_908_n 0.0031593f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_295 N_A_c_305_n N_VPWR_c_988_n 0.00783891f $X=1.25 $Y=1.86 $X2=0 $Y2=0
cc_296 N_A_c_305_n N_VPWR_c_996_n 0.00513163f $X=1.25 $Y=1.86 $X2=0 $Y2=0
cc_297 N_A_c_305_n N_VPWR_c_987_n 0.00484068f $X=1.25 $Y=1.86 $X2=0 $Y2=0
cc_298 A N_VGND_M1017_d 0.00601105f $X=1.115 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_299 N_A_c_306_n N_VGND_c_1382_n 0.00305517f $X=1.325 $Y=1.42 $X2=0 $Y2=0
cc_300 N_A_c_306_n N_VGND_c_1389_n 0.00457172f $X=1.325 $Y=1.42 $X2=0 $Y2=0
cc_301 N_A_440_315#_c_352_n N_B_c_465_n 0.0166387f $X=2.29 $Y=2.02 $X2=-0.19
+ $Y2=-0.245
cc_302 N_A_440_315#_c_352_n N_B_c_466_n 0.00882199f $X=2.29 $Y=2.02 $X2=0 $Y2=0
cc_303 N_A_440_315#_M1008_g N_B_M1019_g 0.0109333f $X=2.505 $Y=0.995 $X2=0 $Y2=0
cc_304 N_A_440_315#_M1008_g N_B_c_453_n 0.00355453f $X=2.505 $Y=0.995 $X2=0
+ $Y2=0
cc_305 N_A_440_315#_c_352_n N_B_c_468_n 0.00278823f $X=2.29 $Y=2.02 $X2=0 $Y2=0
cc_306 N_A_440_315#_c_355_n N_B_c_468_n 0.0022019f $X=3.275 $Y=1.82 $X2=0 $Y2=0
cc_307 N_A_440_315#_c_352_n N_B_c_470_n 0.0201585f $X=2.29 $Y=2.02 $X2=0 $Y2=0
cc_308 N_A_440_315#_c_340_n N_B_c_470_n 0.0097793f $X=3.185 $Y=1.65 $X2=0 $Y2=0
cc_309 N_A_440_315#_c_355_n N_B_c_470_n 0.019149f $X=3.275 $Y=1.82 $X2=0 $Y2=0
cc_310 N_A_440_315#_c_355_n N_B_c_471_n 0.00882199f $X=3.275 $Y=1.82 $X2=0 $Y2=0
cc_311 N_A_440_315#_M1008_g N_B_M1016_g 0.0121494f $X=2.505 $Y=0.995 $X2=0 $Y2=0
cc_312 N_A_440_315#_c_340_n N_B_M1016_g 0.00886717f $X=3.185 $Y=1.65 $X2=0 $Y2=0
cc_313 N_A_440_315#_M1020_g N_B_M1016_g 0.0152172f $X=3.765 $Y=0.945 $X2=0 $Y2=0
cc_314 N_A_440_315#_M1020_g N_B_c_456_n 0.00737859f $X=3.765 $Y=0.945 $X2=0
+ $Y2=0
cc_315 N_A_440_315#_M1020_g N_B_c_457_n 7.80508e-19 $X=3.765 $Y=0.945 $X2=0
+ $Y2=0
cc_316 N_A_440_315#_c_345_n N_B_c_457_n 4.54349e-19 $X=3.81 $Y=1.435 $X2=0 $Y2=0
cc_317 N_A_440_315#_c_348_n N_B_c_457_n 0.00112154f $X=4.665 $Y=1.985 $X2=0
+ $Y2=0
cc_318 N_A_440_315#_c_349_n N_B_c_457_n 3.32909e-19 $X=3.89 $Y=1.57 $X2=0 $Y2=0
cc_319 N_A_440_315#_c_350_n N_B_c_457_n 0.0180459f $X=3.89 $Y=1.57 $X2=0 $Y2=0
cc_320 N_A_440_315#_c_348_n N_B_c_458_n 0.0136292f $X=4.665 $Y=1.985 $X2=0 $Y2=0
cc_321 N_A_440_315#_M1020_g N_B_c_459_n 0.0167537f $X=3.765 $Y=0.945 $X2=0 $Y2=0
cc_322 N_A_440_315#_c_346_n N_B_c_459_n 0.0210838f $X=4.58 $Y=0.68 $X2=0 $Y2=0
cc_323 N_A_440_315#_c_346_n N_B_c_460_n 7.32755e-19 $X=4.58 $Y=0.68 $X2=0 $Y2=0
cc_324 N_A_440_315#_c_348_n N_B_c_460_n 0.0141116f $X=4.665 $Y=1.985 $X2=0 $Y2=0
cc_325 N_A_440_315#_c_348_n N_B_c_461_n 0.0123873f $X=4.665 $Y=1.985 $X2=0 $Y2=0
cc_326 N_A_440_315#_c_348_n N_B_c_462_n 0.00418241f $X=4.665 $Y=1.985 $X2=0
+ $Y2=0
cc_327 N_A_440_315#_c_348_n B 0.0272067f $X=4.665 $Y=1.985 $X2=0 $Y2=0
cc_328 N_A_440_315#_M1008_g N_A_27_134#_c_903_n 0.00139233f $X=2.505 $Y=0.995
+ $X2=0 $Y2=0
cc_329 N_A_440_315#_c_341_n N_A_27_134#_c_904_n 0.00735194f $X=2.58 $Y=1.65
+ $X2=0 $Y2=0
cc_330 N_A_440_315#_c_351_n N_A_27_134#_c_906_n 0.0130602f $X=2.29 $Y=1.93 $X2=0
+ $Y2=0
cc_331 N_A_440_315#_c_352_n N_A_27_134#_c_906_n 0.00948677f $X=2.29 $Y=2.02
+ $X2=0 $Y2=0
cc_332 N_A_440_315#_M1008_g N_A_27_134#_c_906_n 3.68706e-19 $X=2.505 $Y=0.995
+ $X2=0 $Y2=0
cc_333 N_A_440_315#_c_340_n N_A_27_134#_c_906_n 0.00691558f $X=3.185 $Y=1.65
+ $X2=0 $Y2=0
cc_334 N_A_440_315#_c_341_n N_A_27_134#_c_906_n 0.0156112f $X=2.58 $Y=1.65 $X2=0
+ $Y2=0
cc_335 N_A_440_315#_c_355_n N_A_27_134#_c_906_n 7.07311e-19 $X=3.275 $Y=1.82
+ $X2=0 $Y2=0
cc_336 N_A_440_315#_c_344_n N_A_27_134#_c_906_n 4.81873e-19 $X=3.275 $Y=1.65
+ $X2=0 $Y2=0
cc_337 N_A_440_315#_M1008_g N_A_27_134#_c_907_n 0.00622153f $X=2.505 $Y=0.995
+ $X2=0 $Y2=0
cc_338 N_A_440_315#_M1008_g N_A_27_134#_c_910_n 0.0133067f $X=2.505 $Y=0.995
+ $X2=0 $Y2=0
cc_339 N_A_440_315#_M1008_g N_A_27_134#_c_911_n 0.0140064f $X=2.505 $Y=0.995
+ $X2=0 $Y2=0
cc_340 N_A_440_315#_c_340_n N_A_27_134#_c_911_n 0.00629061f $X=3.185 $Y=1.65
+ $X2=0 $Y2=0
cc_341 N_A_440_315#_c_348_n N_VPWR_c_989_n 0.0729754f $X=4.665 $Y=1.985 $X2=0
+ $Y2=0
cc_342 N_A_440_315#_c_348_n N_VPWR_c_996_n 0.00749631f $X=4.665 $Y=1.985 $X2=0
+ $Y2=0
cc_343 N_A_440_315#_c_348_n N_VPWR_c_987_n 0.0062048f $X=4.665 $Y=1.985 $X2=0
+ $Y2=0
cc_344 N_A_440_315#_c_352_n N_A_372_419#_c_1095_n 0.00270318f $X=2.29 $Y=2.02
+ $X2=0 $Y2=0
cc_345 N_A_440_315#_c_352_n N_A_372_419#_c_1096_n 0.0141907f $X=2.29 $Y=2.02
+ $X2=0 $Y2=0
cc_346 N_A_440_315#_c_355_n N_A_372_419#_c_1096_n 0.0121869f $X=3.275 $Y=1.82
+ $X2=0 $Y2=0
cc_347 N_A_440_315#_c_355_n N_A_372_419#_c_1085_n 0.0146066f $X=3.275 $Y=1.82
+ $X2=0 $Y2=0
cc_348 N_A_440_315#_c_342_n N_A_372_419#_c_1085_n 0.0145675f $X=3.69 $Y=1.65
+ $X2=0 $Y2=0
cc_349 N_A_440_315#_M1020_g N_A_372_419#_c_1085_n 0.013414f $X=3.765 $Y=0.945
+ $X2=0 $Y2=0
cc_350 N_A_440_315#_c_344_n N_A_372_419#_c_1085_n 0.00210238f $X=3.275 $Y=1.65
+ $X2=0 $Y2=0
cc_351 N_A_440_315#_c_345_n N_A_372_419#_c_1085_n 0.0471932f $X=3.81 $Y=1.435
+ $X2=0 $Y2=0
cc_352 N_A_440_315#_c_347_n N_A_372_419#_c_1085_n 0.0133618f $X=3.895 $Y=0.68
+ $X2=0 $Y2=0
cc_353 N_A_440_315#_c_349_n N_A_372_419#_c_1085_n 0.0219455f $X=3.89 $Y=1.57
+ $X2=0 $Y2=0
cc_354 N_A_440_315#_M1009_s N_A_372_419#_c_1086_n 0.00231738f $X=4.585 $Y=0.37
+ $X2=0 $Y2=0
cc_355 N_A_440_315#_M1020_g N_A_372_419#_c_1086_n 0.00174767f $X=3.765 $Y=0.945
+ $X2=0 $Y2=0
cc_356 N_A_440_315#_c_346_n N_A_372_419#_c_1086_n 0.0642029f $X=4.58 $Y=0.68
+ $X2=0 $Y2=0
cc_357 N_A_440_315#_c_347_n N_A_372_419#_c_1086_n 0.0129683f $X=3.895 $Y=0.68
+ $X2=0 $Y2=0
cc_358 N_A_440_315#_M1008_g N_A_416_113#_c_1232_n 0.00586918f $X=2.505 $Y=0.995
+ $X2=0 $Y2=0
cc_359 N_A_440_315#_M1008_g N_A_416_113#_c_1233_n 0.0029704f $X=2.505 $Y=0.995
+ $X2=0 $Y2=0
cc_360 N_A_440_315#_c_355_n N_A_416_113#_c_1241_n 0.0041627f $X=3.275 $Y=1.82
+ $X2=0 $Y2=0
cc_361 N_A_440_315#_M1011_s N_A_416_113#_c_1243_n 0.00703981f $X=4.52 $Y=1.84
+ $X2=0 $Y2=0
cc_362 N_A_440_315#_c_355_n N_A_416_113#_c_1243_n 0.00642085f $X=3.275 $Y=1.82
+ $X2=0 $Y2=0
cc_363 N_A_440_315#_c_342_n N_A_416_113#_c_1243_n 0.00372063f $X=3.69 $Y=1.65
+ $X2=0 $Y2=0
cc_364 N_A_440_315#_c_344_n N_A_416_113#_c_1243_n 3.49166e-19 $X=3.275 $Y=1.65
+ $X2=0 $Y2=0
cc_365 N_A_440_315#_c_348_n N_A_416_113#_c_1243_n 0.0195384f $X=4.665 $Y=1.985
+ $X2=0 $Y2=0
cc_366 N_A_440_315#_c_349_n N_A_416_113#_c_1243_n 0.00212633f $X=3.89 $Y=1.57
+ $X2=0 $Y2=0
cc_367 N_A_440_315#_c_350_n N_A_416_113#_c_1243_n 9.6797e-19 $X=3.89 $Y=1.57
+ $X2=0 $Y2=0
cc_368 N_A_440_315#_c_355_n N_A_416_113#_c_1261_n 0.0025958f $X=3.275 $Y=1.82
+ $X2=0 $Y2=0
cc_369 N_A_440_315#_c_351_n N_A_416_113#_c_1244_n 3.71439e-19 $X=2.29 $Y=1.93
+ $X2=0 $Y2=0
cc_370 N_A_440_315#_c_340_n N_A_416_113#_c_1244_n 0.006398f $X=3.185 $Y=1.65
+ $X2=0 $Y2=0
cc_371 N_A_440_315#_c_355_n N_A_416_113#_c_1244_n 0.00252805f $X=3.275 $Y=1.82
+ $X2=0 $Y2=0
cc_372 N_A_440_315#_c_351_n N_A_416_113#_c_1239_n 5.37562e-19 $X=2.29 $Y=1.93
+ $X2=0 $Y2=0
cc_373 N_A_440_315#_M1008_g N_A_416_113#_c_1239_n 0.00190803f $X=2.505 $Y=0.995
+ $X2=0 $Y2=0
cc_374 N_A_440_315#_c_340_n N_A_416_113#_c_1239_n 0.0104884f $X=3.185 $Y=1.65
+ $X2=0 $Y2=0
cc_375 N_A_440_315#_c_355_n N_A_416_113#_c_1239_n 0.0014578f $X=3.275 $Y=1.82
+ $X2=0 $Y2=0
cc_376 N_A_440_315#_c_344_n N_A_416_113#_c_1239_n 0.00584743f $X=3.275 $Y=1.65
+ $X2=0 $Y2=0
cc_377 N_B_c_461_n N_A_1162_379#_c_588_n 0.00261039f $X=4.89 $Y=1.765 $X2=0
+ $Y2=0
cc_378 N_B_M1019_g N_A_27_134#_c_902_n 0.00578498f $X=2.005 $Y=0.885 $X2=0 $Y2=0
cc_379 N_B_M1019_g N_A_27_134#_c_903_n 0.0128816f $X=2.005 $Y=0.885 $X2=0 $Y2=0
cc_380 N_B_M1019_g N_A_27_134#_c_904_n 0.00536183f $X=2.005 $Y=0.885 $X2=0 $Y2=0
cc_381 N_B_c_465_n N_A_27_134#_c_905_n 0.00234227f $X=1.785 $Y=3.01 $X2=0 $Y2=0
cc_382 N_B_c_465_n N_A_27_134#_c_906_n 5.84264e-19 $X=1.785 $Y=3.01 $X2=0 $Y2=0
cc_383 N_B_c_470_n N_A_27_134#_c_906_n 0.00634934f $X=2.74 $Y=2.81 $X2=0 $Y2=0
cc_384 N_B_M1019_g N_A_27_134#_c_907_n 3.62456e-19 $X=2.005 $Y=0.885 $X2=0 $Y2=0
cc_385 N_B_M1016_g N_A_27_134#_c_907_n 3.86096e-19 $X=3.175 $Y=0.885 $X2=0 $Y2=0
cc_386 N_B_M1016_g N_A_27_134#_c_911_n 0.00169191f $X=3.175 $Y=0.885 $X2=0 $Y2=0
cc_387 N_B_c_467_n N_VPWR_c_988_n 0.00239041f $X=1.875 $Y=3.15 $X2=0 $Y2=0
cc_388 N_B_c_471_n N_VPWR_c_989_n 0.00229165f $X=4.295 $Y=3.15 $X2=0 $Y2=0
cc_389 N_B_c_458_n N_VPWR_c_989_n 8.69313e-19 $X=4.37 $Y=3.075 $X2=0 $Y2=0
cc_390 N_B_c_461_n N_VPWR_c_989_n 0.0199133f $X=4.89 $Y=1.765 $X2=0 $Y2=0
cc_391 B N_VPWR_c_989_n 0.0134342f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_392 N_B_c_467_n N_VPWR_c_996_n 0.060425f $X=1.875 $Y=3.15 $X2=0 $Y2=0
cc_393 N_B_c_461_n N_VPWR_c_996_n 0.00413917f $X=4.89 $Y=1.765 $X2=0 $Y2=0
cc_394 N_B_c_466_n N_VPWR_c_987_n 0.0180126f $X=2.65 $Y=3.15 $X2=0 $Y2=0
cc_395 N_B_c_467_n N_VPWR_c_987_n 0.00674619f $X=1.875 $Y=3.15 $X2=0 $Y2=0
cc_396 N_B_c_471_n N_VPWR_c_987_n 0.0436101f $X=4.295 $Y=3.15 $X2=0 $Y2=0
cc_397 N_B_c_461_n N_VPWR_c_987_n 0.0081836f $X=4.89 $Y=1.765 $X2=0 $Y2=0
cc_398 N_B_c_474_n N_VPWR_c_987_n 0.00441524f $X=2.74 $Y=3.15 $X2=0 $Y2=0
cc_399 N_B_c_465_n N_A_372_419#_c_1095_n 0.00536656f $X=1.785 $Y=3.01 $X2=0
+ $Y2=0
cc_400 N_B_c_470_n N_A_372_419#_c_1096_n 0.0149409f $X=2.74 $Y=2.81 $X2=0 $Y2=0
cc_401 N_B_c_465_n N_A_372_419#_c_1108_n 0.00185396f $X=1.785 $Y=3.01 $X2=0
+ $Y2=0
cc_402 N_B_M1016_g N_A_372_419#_c_1085_n 0.00780549f $X=3.175 $Y=0.885 $X2=0
+ $Y2=0
cc_403 N_B_c_456_n N_A_372_419#_c_1086_n 0.0143527f $X=4.36 $Y=0.18 $X2=0 $Y2=0
cc_404 N_B_c_459_n N_A_372_419#_c_1086_n 0.0121042f $X=4.435 $Y=1.22 $X2=0 $Y2=0
cc_405 N_B_c_462_n N_A_372_419#_c_1086_n 0.0134432f $X=4.935 $Y=1.22 $X2=0 $Y2=0
cc_406 N_B_M1016_g N_A_372_419#_c_1087_n 0.00724099f $X=3.175 $Y=0.885 $X2=0
+ $Y2=0
cc_407 N_B_c_456_n N_A_372_419#_c_1087_n 0.00420304f $X=4.36 $Y=0.18 $X2=0 $Y2=0
cc_408 N_B_c_459_n N_A_372_419#_c_1136_n 8.24696e-19 $X=4.435 $Y=1.22 $X2=0
+ $Y2=0
cc_409 N_B_c_462_n N_A_372_419#_c_1136_n 0.00826933f $X=4.935 $Y=1.22 $X2=0
+ $Y2=0
cc_410 N_B_c_461_n N_A_372_419#_c_1088_n 5.83726e-19 $X=4.89 $Y=1.765 $X2=0
+ $Y2=0
cc_411 B N_A_372_419#_c_1088_n 0.0050401f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_412 N_B_c_461_n N_A_372_419#_c_1140_n 6.76062e-19 $X=4.89 $Y=1.765 $X2=0
+ $Y2=0
cc_413 N_B_c_462_n N_A_372_419#_c_1140_n 0.00670237f $X=4.935 $Y=1.22 $X2=0
+ $Y2=0
cc_414 B N_A_372_419#_c_1140_n 0.00729471f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_415 N_B_c_453_n N_A_416_113#_c_1233_n 0.0129409f $X=3.1 $Y=0.18 $X2=0 $Y2=0
cc_416 N_B_M1016_g N_A_416_113#_c_1233_n 0.00870892f $X=3.175 $Y=0.885 $X2=0
+ $Y2=0
cc_417 N_B_M1019_g N_A_416_113#_c_1234_n 0.0064969f $X=2.005 $Y=0.885 $X2=0
+ $Y2=0
cc_418 N_B_c_453_n N_A_416_113#_c_1234_n 0.00305251f $X=3.1 $Y=0.18 $X2=0 $Y2=0
cc_419 N_B_c_462_n N_A_416_113#_c_1236_n 0.00482248f $X=4.935 $Y=1.22 $X2=0
+ $Y2=0
cc_420 B N_A_416_113#_c_1236_n 3.28587e-19 $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_421 N_B_c_457_n N_A_416_113#_c_1243_n 0.00154074f $X=4.37 $Y=1.52 $X2=0 $Y2=0
cc_422 N_B_c_458_n N_A_416_113#_c_1243_n 0.00528025f $X=4.37 $Y=3.075 $X2=0
+ $Y2=0
cc_423 N_B_c_460_n N_A_416_113#_c_1243_n 0.0025141f $X=4.8 $Y=1.295 $X2=0 $Y2=0
cc_424 N_B_c_461_n N_A_416_113#_c_1243_n 0.0106552f $X=4.89 $Y=1.765 $X2=0 $Y2=0
cc_425 B N_A_416_113#_c_1243_n 0.00403396f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_426 N_B_c_470_n N_A_416_113#_c_1244_n 0.00390493f $X=2.74 $Y=2.81 $X2=0 $Y2=0
cc_427 N_B_c_461_n N_A_416_113#_c_1246_n 0.00206878f $X=4.89 $Y=1.765 $X2=0
+ $Y2=0
cc_428 N_B_M1016_g N_A_416_113#_c_1239_n 0.0203921f $X=3.175 $Y=0.885 $X2=0
+ $Y2=0
cc_429 N_B_c_461_n N_A_416_113#_c_1240_n 0.0118769f $X=4.89 $Y=1.765 $X2=0 $Y2=0
cc_430 B N_A_416_113#_c_1240_n 0.020093f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_431 N_B_c_462_n N_VGND_c_1378_n 0.00174649f $X=4.935 $Y=1.22 $X2=0 $Y2=0
cc_432 N_B_c_454_n N_VGND_c_1382_n 0.0625641f $X=2.08 $Y=0.18 $X2=0 $Y2=0
cc_433 N_B_c_462_n N_VGND_c_1382_n 0.00278237f $X=4.935 $Y=1.22 $X2=0 $Y2=0
cc_434 N_B_c_453_n N_VGND_c_1389_n 0.0268561f $X=3.1 $Y=0.18 $X2=0 $Y2=0
cc_435 N_B_c_454_n N_VGND_c_1389_n 0.0104612f $X=2.08 $Y=0.18 $X2=0 $Y2=0
cc_436 N_B_c_456_n N_VGND_c_1389_n 0.0367758f $X=4.36 $Y=0.18 $X2=0 $Y2=0
cc_437 N_B_c_462_n N_VGND_c_1389_n 0.00359083f $X=4.935 $Y=1.22 $X2=0 $Y2=0
cc_438 N_B_c_463_n N_VGND_c_1389_n 0.00512617f $X=3.175 $Y=0.18 $X2=0 $Y2=0
cc_439 N_A_1162_379#_c_590_n N_C_c_700_n 0.00566283f $X=6.155 $Y=1.895 $X2=0
+ $Y2=0
cc_440 N_A_1162_379#_c_592_n N_C_c_700_n 2.17042e-19 $X=6.095 $Y=2.905 $X2=0
+ $Y2=0
cc_441 N_A_1162_379#_c_589_n N_C_c_701_n 0.00977938f $X=5.9 $Y=2.045 $X2=0 $Y2=0
cc_442 N_A_1162_379#_c_591_n N_C_c_701_n 0.00566283f $X=6.155 $Y=1.97 $X2=0
+ $Y2=0
cc_443 N_A_1162_379#_c_592_n N_C_c_701_n 0.00478999f $X=6.095 $Y=2.905 $X2=0
+ $Y2=0
cc_444 N_A_1162_379#_c_593_n N_C_c_701_n 0.0165459f $X=7.28 $Y=2.99 $X2=0 $Y2=0
cc_445 N_A_1162_379#_c_595_n N_C_c_701_n 0.00524322f $X=7.365 $Y=2.905 $X2=0
+ $Y2=0
cc_446 N_A_1162_379#_M1004_g N_C_c_691_n 0.00796138f $X=6.155 $Y=0.855 $X2=0
+ $Y2=0
cc_447 N_A_1162_379#_c_584_n N_C_c_692_n 0.00422824f $X=7.72 $Y=2.195 $X2=0
+ $Y2=0
cc_448 N_A_1162_379#_c_585_n N_C_c_692_n 0.002567f $X=7.9 $Y=1.435 $X2=0 $Y2=0
cc_449 N_A_1162_379#_c_587_n N_C_c_693_n 2.17042e-19 $X=6.015 $Y=1.52 $X2=0
+ $Y2=0
cc_450 N_A_1162_379#_c_588_n N_C_c_693_n 0.0136242f $X=6.015 $Y=1.52 $X2=0 $Y2=0
cc_451 N_A_1162_379#_c_586_n N_C_c_694_n 0.00961036f $X=7.86 $Y=0.6 $X2=0 $Y2=0
cc_452 N_A_1162_379#_c_595_n N_C_c_695_n 0.00233656f $X=7.365 $Y=2.905 $X2=0
+ $Y2=0
cc_453 N_A_1162_379#_c_584_n N_C_c_695_n 0.0364551f $X=7.72 $Y=2.195 $X2=0 $Y2=0
cc_454 N_A_1162_379#_c_585_n N_C_c_695_n 0.0115509f $X=7.9 $Y=1.435 $X2=0 $Y2=0
cc_455 N_A_1162_379#_c_586_n N_C_c_695_n 0.00287098f $X=7.86 $Y=0.6 $X2=0 $Y2=0
cc_456 N_A_1162_379#_c_585_n N_C_c_696_n 5.32204e-19 $X=7.9 $Y=1.435 $X2=0 $Y2=0
cc_457 N_A_1162_379#_c_586_n N_C_c_696_n 0.0128944f $X=7.86 $Y=0.6 $X2=0 $Y2=0
cc_458 N_A_1162_379#_c_586_n N_C_c_697_n 0.00248458f $X=7.86 $Y=0.6 $X2=0 $Y2=0
cc_459 N_A_1162_379#_c_586_n N_C_c_698_n 0.00802643f $X=7.86 $Y=0.6 $X2=0 $Y2=0
cc_460 N_A_1162_379#_c_592_n N_A_1195_424#_M1013_d 0.0136995f $X=6.095 $Y=2.905
+ $X2=0 $Y2=0
cc_461 N_A_1162_379#_c_593_n N_A_1195_424#_M1013_d 0.00919565f $X=7.28 $Y=2.99
+ $X2=0 $Y2=0
cc_462 N_A_1162_379#_c_594_n N_A_1195_424#_M1013_d 4.50551e-19 $X=6.18 $Y=2.99
+ $X2=0 $Y2=0
cc_463 N_A_1162_379#_c_586_n N_A_1195_424#_M1002_g 0.00421174f $X=7.86 $Y=0.6
+ $X2=0 $Y2=0
cc_464 N_A_1162_379#_c_585_n N_A_1195_424#_c_792_n 0.00141437f $X=7.9 $Y=1.435
+ $X2=0 $Y2=0
cc_465 N_A_1162_379#_c_586_n N_A_1195_424#_c_792_n 0.00100179f $X=7.86 $Y=0.6
+ $X2=0 $Y2=0
cc_466 N_A_1162_379#_M1004_g N_A_1195_424#_c_795_n 0.00398659f $X=6.155 $Y=0.855
+ $X2=0 $Y2=0
cc_467 N_A_1162_379#_c_587_n N_A_1195_424#_c_796_n 0.0495155f $X=6.015 $Y=1.52
+ $X2=0 $Y2=0
cc_468 N_A_1162_379#_c_588_n N_A_1195_424#_c_796_n 0.00304279f $X=6.015 $Y=1.52
+ $X2=0 $Y2=0
cc_469 N_A_1162_379#_c_584_n N_A_1195_424#_c_797_n 0.00164698f $X=7.72 $Y=2.195
+ $X2=0 $Y2=0
cc_470 N_A_1162_379#_c_585_n N_A_1195_424#_c_797_n 0.0135398f $X=7.9 $Y=1.435
+ $X2=0 $Y2=0
cc_471 N_A_1162_379#_c_586_n N_A_1195_424#_c_797_n 0.00890402f $X=7.86 $Y=0.6
+ $X2=0 $Y2=0
cc_472 N_A_1162_379#_M1010_s N_A_1195_424#_c_803_n 0.00536549f $X=7.3 $Y=1.84
+ $X2=0 $Y2=0
cc_473 N_A_1162_379#_c_584_n N_A_1195_424#_c_803_n 0.0259303f $X=7.72 $Y=2.195
+ $X2=0 $Y2=0
cc_474 N_A_1162_379#_c_585_n N_A_1195_424#_c_803_n 0.00703403f $X=7.9 $Y=1.435
+ $X2=0 $Y2=0
cc_475 N_A_1162_379#_c_591_n N_A_1195_424#_c_804_n 0.00253348f $X=6.155 $Y=1.97
+ $X2=0 $Y2=0
cc_476 N_A_1162_379#_c_592_n N_A_1195_424#_c_804_n 0.00729123f $X=6.095 $Y=2.905
+ $X2=0 $Y2=0
cc_477 N_A_1162_379#_c_590_n N_A_1195_424#_c_798_n 0.00304279f $X=6.155 $Y=1.895
+ $X2=0 $Y2=0
cc_478 N_A_1162_379#_c_592_n N_A_1195_424#_c_798_n 0.0495155f $X=6.095 $Y=2.905
+ $X2=0 $Y2=0
cc_479 N_A_1162_379#_c_593_n N_A_1195_424#_c_798_n 0.012307f $X=7.28 $Y=2.99
+ $X2=0 $Y2=0
cc_480 N_A_1162_379#_c_584_n N_A_1195_424#_c_806_n 0.00540375f $X=7.72 $Y=2.195
+ $X2=0 $Y2=0
cc_481 N_A_1162_379#_c_589_n N_VPWR_c_989_n 0.00403661f $X=5.9 $Y=2.045 $X2=0
+ $Y2=0
cc_482 N_A_1162_379#_c_591_n N_VPWR_c_989_n 3.50637e-19 $X=6.155 $Y=1.97 $X2=0
+ $Y2=0
cc_483 N_A_1162_379#_c_584_n N_VPWR_c_990_n 0.0501802f $X=7.72 $Y=2.195 $X2=0
+ $Y2=0
cc_484 N_A_1162_379#_c_585_n N_VPWR_c_990_n 0.00322867f $X=7.9 $Y=1.435 $X2=0
+ $Y2=0
cc_485 N_A_1162_379#_c_593_n N_VPWR_c_991_n 0.00703128f $X=7.28 $Y=2.99 $X2=0
+ $Y2=0
cc_486 N_A_1162_379#_c_595_n N_VPWR_c_1038_n 0.0145268f $X=7.365 $Y=2.905 $X2=0
+ $Y2=0
cc_487 N_A_1162_379#_c_589_n N_VPWR_c_997_n 0.00445602f $X=5.9 $Y=2.045 $X2=0
+ $Y2=0
cc_488 N_A_1162_379#_c_593_n N_VPWR_c_997_n 0.0824005f $X=7.28 $Y=2.99 $X2=0
+ $Y2=0
cc_489 N_A_1162_379#_c_594_n N_VPWR_c_997_n 0.0121867f $X=6.18 $Y=2.99 $X2=0
+ $Y2=0
cc_490 N_A_1162_379#_c_589_n N_VPWR_c_987_n 0.00865371f $X=5.9 $Y=2.045 $X2=0
+ $Y2=0
cc_491 N_A_1162_379#_c_593_n N_VPWR_c_987_n 0.0472477f $X=7.28 $Y=2.99 $X2=0
+ $Y2=0
cc_492 N_A_1162_379#_c_594_n N_VPWR_c_987_n 0.00660921f $X=6.18 $Y=2.99 $X2=0
+ $Y2=0
cc_493 N_A_1162_379#_c_584_n N_VPWR_c_987_n 0.0126028f $X=7.72 $Y=2.195 $X2=0
+ $Y2=0
cc_494 N_A_1162_379#_c_593_n N_A_372_419#_M1023_d 0.0031459f $X=7.28 $Y=2.99
+ $X2=0 $Y2=0
cc_495 N_A_1162_379#_M1004_g N_A_372_419#_c_1089_n 0.00442722f $X=6.155 $Y=0.855
+ $X2=0 $Y2=0
cc_496 N_A_1162_379#_M1004_g N_A_372_419#_c_1090_n 0.00730004f $X=6.155 $Y=0.855
+ $X2=0 $Y2=0
cc_497 N_A_1162_379#_c_586_n N_A_372_419#_c_1090_n 0.00472011f $X=7.86 $Y=0.6
+ $X2=0 $Y2=0
cc_498 N_A_1162_379#_c_593_n N_A_372_419#_c_1098_n 0.0160379f $X=7.28 $Y=2.99
+ $X2=0 $Y2=0
cc_499 N_A_1162_379#_c_595_n N_A_372_419#_c_1098_n 0.0119875f $X=7.365 $Y=2.905
+ $X2=0 $Y2=0
cc_500 N_A_1162_379#_c_584_n N_A_372_419#_c_1098_n 0.0235139f $X=7.72 $Y=2.195
+ $X2=0 $Y2=0
cc_501 N_A_1162_379#_M1010_s N_A_372_419#_c_1099_n 0.00358171f $X=7.3 $Y=1.84
+ $X2=0 $Y2=0
cc_502 N_A_1162_379#_c_584_n N_A_372_419#_c_1099_n 0.0204983f $X=7.72 $Y=2.195
+ $X2=0 $Y2=0
cc_503 N_A_1162_379#_M1010_s N_A_372_419#_c_1092_n 2.42835e-19 $X=7.3 $Y=1.84
+ $X2=0 $Y2=0
cc_504 N_A_1162_379#_c_584_n N_A_372_419#_c_1092_n 0.0181633f $X=7.72 $Y=2.195
+ $X2=0 $Y2=0
cc_505 N_A_1162_379#_c_585_n N_A_372_419#_c_1092_n 0.0130101f $X=7.9 $Y=1.435
+ $X2=0 $Y2=0
cc_506 N_A_1162_379#_c_586_n N_A_372_419#_c_1092_n 0.0076654f $X=7.86 $Y=0.6
+ $X2=0 $Y2=0
cc_507 N_A_1162_379#_c_586_n N_A_372_419#_c_1093_n 0.0505046f $X=7.86 $Y=0.6
+ $X2=0 $Y2=0
cc_508 N_A_1162_379#_c_586_n N_A_372_419#_c_1094_n 0.0130296f $X=7.86 $Y=0.6
+ $X2=0 $Y2=0
cc_509 N_A_1162_379#_c_589_n N_A_416_113#_c_1242_n 0.0124279f $X=5.9 $Y=2.045
+ $X2=0 $Y2=0
cc_510 N_A_1162_379#_c_594_n N_A_416_113#_c_1242_n 0.00383537f $X=6.18 $Y=2.99
+ $X2=0 $Y2=0
cc_511 N_A_1162_379#_M1004_g N_A_416_113#_c_1235_n 0.0150552f $X=6.155 $Y=0.855
+ $X2=0 $Y2=0
cc_512 N_A_1162_379#_c_587_n N_A_416_113#_c_1235_n 0.0251443f $X=6.015 $Y=1.52
+ $X2=0 $Y2=0
cc_513 N_A_1162_379#_c_588_n N_A_416_113#_c_1235_n 0.00161433f $X=6.015 $Y=1.52
+ $X2=0 $Y2=0
cc_514 N_A_1162_379#_M1004_g N_A_416_113#_c_1291_n 0.0107362f $X=6.155 $Y=0.855
+ $X2=0 $Y2=0
cc_515 N_A_1162_379#_M1004_g N_A_416_113#_c_1292_n 0.00552867f $X=6.155 $Y=0.855
+ $X2=0 $Y2=0
cc_516 N_A_1162_379#_c_592_n N_A_416_113#_c_1245_n 0.00107267f $X=6.095 $Y=2.905
+ $X2=0 $Y2=0
cc_517 N_A_1162_379#_c_589_n N_A_416_113#_c_1246_n 0.00249396f $X=5.9 $Y=2.045
+ $X2=0 $Y2=0
cc_518 N_A_1162_379#_c_591_n N_A_416_113#_c_1246_n 0.00642395f $X=6.155 $Y=1.97
+ $X2=0 $Y2=0
cc_519 N_A_1162_379#_c_592_n N_A_416_113#_c_1246_n 0.0440127f $X=6.095 $Y=2.905
+ $X2=0 $Y2=0
cc_520 N_A_1162_379#_M1004_g N_A_416_113#_c_1240_n 0.00453554f $X=6.155 $Y=0.855
+ $X2=0 $Y2=0
cc_521 N_A_1162_379#_c_591_n N_A_416_113#_c_1240_n 6.6135e-19 $X=6.155 $Y=1.97
+ $X2=0 $Y2=0
cc_522 N_A_1162_379#_c_592_n N_A_416_113#_c_1240_n 0.0110355f $X=6.095 $Y=2.905
+ $X2=0 $Y2=0
cc_523 N_A_1162_379#_c_587_n N_A_416_113#_c_1240_n 0.0248017f $X=6.015 $Y=1.52
+ $X2=0 $Y2=0
cc_524 N_A_1162_379#_c_588_n N_A_416_113#_c_1240_n 0.00507613f $X=6.015 $Y=1.52
+ $X2=0 $Y2=0
cc_525 N_A_1162_379#_M1004_g N_VGND_c_1378_n 2.09474e-19 $X=6.155 $Y=0.855 $X2=0
+ $Y2=0
cc_526 N_A_1162_379#_c_586_n N_VGND_c_1379_n 0.0415257f $X=7.86 $Y=0.6 $X2=0
+ $Y2=0
cc_527 N_A_1162_379#_M1004_g N_VGND_c_1383_n 6.51701e-19 $X=6.155 $Y=0.855 $X2=0
+ $Y2=0
cc_528 N_A_1162_379#_c_586_n N_VGND_c_1383_n 0.0101731f $X=7.86 $Y=0.6 $X2=0
+ $Y2=0
cc_529 N_A_1162_379#_c_586_n N_VGND_c_1389_n 0.00902782f $X=7.86 $Y=0.6 $X2=0
+ $Y2=0
cc_530 N_C_c_698_n N_A_1195_424#_M1002_g 0.0144313f $X=8.075 $Y=0.885 $X2=0
+ $Y2=0
cc_531 N_C_c_694_n N_A_1195_424#_c_792_n 0.00538345f $X=7.735 $Y=1.355 $X2=0
+ $Y2=0
cc_532 N_C_c_695_n N_A_1195_424#_c_792_n 0.00465864f $X=7.75 $Y=1.765 $X2=0
+ $Y2=0
cc_533 N_C_c_695_n N_A_1195_424#_c_793_n 0.00107388f $X=7.75 $Y=1.765 $X2=0
+ $Y2=0
cc_534 N_C_c_691_n N_A_1195_424#_c_795_n 0.00167979f $X=6.835 $Y=1.355 $X2=0
+ $Y2=0
cc_535 C N_A_1195_424#_c_795_n 0.023585f $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_536 N_C_c_693_n N_A_1195_424#_c_796_n 0.00754199f $X=7.14 $Y=1.43 $X2=0 $Y2=0
cc_537 N_C_c_695_n N_A_1195_424#_c_797_n 3.32685e-19 $X=7.75 $Y=1.765 $X2=0
+ $Y2=0
cc_538 N_C_c_701_n N_A_1195_424#_c_803_n 0.00943359f $X=6.66 $Y=2.045 $X2=0
+ $Y2=0
cc_539 N_C_c_692_n N_A_1195_424#_c_803_n 0.00341283f $X=7.66 $Y=1.43 $X2=0 $Y2=0
cc_540 N_C_c_693_n N_A_1195_424#_c_803_n 8.5126e-19 $X=7.14 $Y=1.43 $X2=0 $Y2=0
cc_541 N_C_c_695_n N_A_1195_424#_c_803_n 0.00360171f $X=7.75 $Y=1.765 $X2=0
+ $Y2=0
cc_542 C N_A_1195_424#_c_803_n 0.00148248f $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_543 N_C_c_700_n N_A_1195_424#_c_804_n 5.51094e-19 $X=6.66 $Y=1.955 $X2=0
+ $Y2=0
cc_544 N_C_c_701_n N_A_1195_424#_c_804_n 0.00156705f $X=6.66 $Y=2.045 $X2=0
+ $Y2=0
cc_545 N_C_c_700_n N_A_1195_424#_c_798_n 0.0110861f $X=6.66 $Y=1.955 $X2=0 $Y2=0
cc_546 N_C_c_701_n N_A_1195_424#_c_798_n 0.012877f $X=6.66 $Y=2.045 $X2=0 $Y2=0
cc_547 N_C_c_693_n N_A_1195_424#_c_798_n 0.0054384f $X=7.14 $Y=1.43 $X2=0 $Y2=0
cc_548 C N_A_1195_424#_c_798_n 0.00784722f $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_549 N_C_c_695_n N_A_1195_424#_c_806_n 0.00206666f $X=7.75 $Y=1.765 $X2=0
+ $Y2=0
cc_550 N_C_c_695_n N_VPWR_c_990_n 0.0156941f $X=7.75 $Y=1.765 $X2=0 $Y2=0
cc_551 N_C_c_701_n N_VPWR_c_997_n 0.00278271f $X=6.66 $Y=2.045 $X2=0 $Y2=0
cc_552 N_C_c_695_n N_VPWR_c_997_n 0.00314304f $X=7.75 $Y=1.765 $X2=0 $Y2=0
cc_553 N_C_c_701_n N_VPWR_c_987_n 0.00360843f $X=6.66 $Y=2.045 $X2=0 $Y2=0
cc_554 N_C_c_695_n N_VPWR_c_987_n 0.00411481f $X=7.75 $Y=1.765 $X2=0 $Y2=0
cc_555 N_C_c_691_n N_A_372_419#_c_1090_n 0.00455332f $X=6.835 $Y=1.355 $X2=0
+ $Y2=0
cc_556 N_C_c_698_n N_A_372_419#_c_1090_n 0.00234865f $X=8.075 $Y=0.885 $X2=0
+ $Y2=0
cc_557 N_C_c_701_n N_A_372_419#_c_1098_n 0.005351f $X=6.66 $Y=2.045 $X2=0 $Y2=0
cc_558 N_C_c_695_n N_A_372_419#_c_1098_n 0.00193717f $X=7.75 $Y=1.765 $X2=0
+ $Y2=0
cc_559 N_C_c_692_n N_A_372_419#_c_1099_n 0.00435379f $X=7.66 $Y=1.43 $X2=0 $Y2=0
cc_560 N_C_c_693_n N_A_372_419#_c_1099_n 0.00112054f $X=7.14 $Y=1.43 $X2=0 $Y2=0
cc_561 N_C_c_695_n N_A_372_419#_c_1099_n 0.00116163f $X=7.75 $Y=1.765 $X2=0
+ $Y2=0
cc_562 C N_A_372_419#_c_1099_n 0.00530888f $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_563 N_C_c_700_n N_A_372_419#_c_1100_n 0.00394113f $X=6.66 $Y=1.955 $X2=0
+ $Y2=0
cc_564 N_C_c_693_n N_A_372_419#_c_1100_n 0.00576853f $X=7.14 $Y=1.43 $X2=0 $Y2=0
cc_565 C N_A_372_419#_c_1100_n 0.0141845f $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_566 N_C_c_700_n N_A_372_419#_c_1092_n 0.00399377f $X=6.66 $Y=1.955 $X2=0
+ $Y2=0
cc_567 N_C_c_691_n N_A_372_419#_c_1092_n 3.87848e-19 $X=6.835 $Y=1.355 $X2=0
+ $Y2=0
cc_568 N_C_c_692_n N_A_372_419#_c_1092_n 0.0133863f $X=7.66 $Y=1.43 $X2=0 $Y2=0
cc_569 N_C_c_693_n N_A_372_419#_c_1092_n 0.00180986f $X=7.14 $Y=1.43 $X2=0 $Y2=0
cc_570 N_C_c_694_n N_A_372_419#_c_1092_n 0.00178741f $X=7.735 $Y=1.355 $X2=0
+ $Y2=0
cc_571 N_C_c_695_n N_A_372_419#_c_1092_n 0.00174209f $X=7.75 $Y=1.765 $X2=0
+ $Y2=0
cc_572 C N_A_372_419#_c_1092_n 0.0307052f $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_573 N_C_c_691_n N_A_372_419#_c_1093_n 0.00692779f $X=6.835 $Y=1.355 $X2=0
+ $Y2=0
cc_574 N_C_c_697_n N_A_372_419#_c_1093_n 0.00547767f $X=7.81 $Y=0.96 $X2=0 $Y2=0
cc_575 N_C_c_698_n N_A_372_419#_c_1093_n 9.09628e-19 $X=8.075 $Y=0.885 $X2=0
+ $Y2=0
cc_576 N_C_c_691_n N_A_372_419#_c_1094_n 0.00194033f $X=6.835 $Y=1.355 $X2=0
+ $Y2=0
cc_577 N_C_c_692_n N_A_372_419#_c_1094_n 0.00513991f $X=7.66 $Y=1.43 $X2=0 $Y2=0
cc_578 N_C_c_694_n N_A_372_419#_c_1094_n 0.00375665f $X=7.735 $Y=1.355 $X2=0
+ $Y2=0
cc_579 C N_A_372_419#_c_1094_n 0.00675568f $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_580 C N_A_416_113#_M1007_d 0.00270076f $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_581 N_C_c_691_n N_A_416_113#_c_1291_n 0.00141899f $X=6.835 $Y=1.355 $X2=0
+ $Y2=0
cc_582 N_C_c_691_n N_A_416_113#_c_1237_n 0.00409002f $X=6.835 $Y=1.355 $X2=0
+ $Y2=0
cc_583 N_C_c_693_n N_A_416_113#_c_1237_n 0.00460589f $X=7.14 $Y=1.43 $X2=0 $Y2=0
cc_584 C N_A_416_113#_c_1237_n 0.0110577f $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_585 N_C_c_691_n N_A_416_113#_c_1238_n 0.0113393f $X=6.835 $Y=1.355 $X2=0
+ $Y2=0
cc_586 C N_A_416_113#_c_1238_n 3.08063e-19 $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_587 N_C_c_694_n N_VGND_c_1379_n 5.24626e-19 $X=7.735 $Y=1.355 $X2=0 $Y2=0
cc_588 N_C_c_698_n N_VGND_c_1379_n 0.00684806f $X=8.075 $Y=0.885 $X2=0 $Y2=0
cc_589 N_C_c_698_n N_VGND_c_1383_n 0.00537471f $X=8.075 $Y=0.885 $X2=0 $Y2=0
cc_590 N_C_c_697_n N_VGND_c_1389_n 0.00289176f $X=7.81 $Y=0.96 $X2=0 $Y2=0
cc_591 N_C_c_698_n N_VGND_c_1389_n 0.00539454f $X=8.075 $Y=0.885 $X2=0 $Y2=0
cc_592 N_A_1195_424#_c_803_n N_VPWR_M1010_d 0.0106335f $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_593 N_A_1195_424#_c_849_p N_VPWR_M1010_d 0.00637365f $X=8.4 $Y=2.035 $X2=0
+ $Y2=0
cc_594 N_A_1195_424#_c_806_n N_VPWR_M1010_d 0.00615745f $X=8.4 $Y=2.035 $X2=0
+ $Y2=0
cc_595 N_A_1195_424#_c_799_n N_VPWR_c_990_n 0.00285753f $X=8.645 $Y=1.765 $X2=0
+ $Y2=0
cc_596 N_A_1195_424#_c_803_n N_VPWR_c_990_n 0.0202422f $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_597 N_A_1195_424#_c_849_p N_VPWR_c_990_n 0.00275409f $X=8.4 $Y=2.035 $X2=0
+ $Y2=0
cc_598 N_A_1195_424#_c_806_n N_VPWR_c_990_n 0.0227956f $X=8.4 $Y=2.035 $X2=0
+ $Y2=0
cc_599 N_A_1195_424#_c_799_n N_VPWR_c_991_n 0.0054453f $X=8.645 $Y=1.765 $X2=0
+ $Y2=0
cc_600 N_A_1195_424#_c_801_n N_VPWR_c_993_n 0.0100916f $X=9.095 $Y=1.765 $X2=0
+ $Y2=0
cc_601 N_A_1195_424#_c_792_n N_VPWR_c_1038_n 0.00133964f $X=8.555 $Y=1.485 $X2=0
+ $Y2=0
cc_602 N_A_1195_424#_c_797_n N_VPWR_c_1038_n 0.00123758f $X=8.36 $Y=1.485 $X2=0
+ $Y2=0
cc_603 N_A_1195_424#_c_803_n N_VPWR_c_1038_n 0.00448577f $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_604 N_A_1195_424#_c_849_p N_VPWR_c_1038_n 0.00428557f $X=8.4 $Y=2.035 $X2=0
+ $Y2=0
cc_605 N_A_1195_424#_c_806_n N_VPWR_c_1038_n 0.0144797f $X=8.4 $Y=2.035 $X2=0
+ $Y2=0
cc_606 N_A_1195_424#_c_799_n N_VPWR_c_998_n 0.00445602f $X=8.645 $Y=1.765 $X2=0
+ $Y2=0
cc_607 N_A_1195_424#_c_801_n N_VPWR_c_998_n 0.00445602f $X=9.095 $Y=1.765 $X2=0
+ $Y2=0
cc_608 N_A_1195_424#_c_799_n N_VPWR_c_987_n 0.00861831f $X=8.645 $Y=1.765 $X2=0
+ $Y2=0
cc_609 N_A_1195_424#_c_801_n N_VPWR_c_987_n 0.00861084f $X=9.095 $Y=1.765 $X2=0
+ $Y2=0
cc_610 N_A_1195_424#_c_803_n N_A_372_419#_c_1098_n 0.0191656f $X=8.255 $Y=2.035
+ $X2=0 $Y2=0
cc_611 N_A_1195_424#_c_804_n N_A_372_419#_c_1098_n 0.0011513f $X=6.625 $Y=2.035
+ $X2=0 $Y2=0
cc_612 N_A_1195_424#_c_798_n N_A_372_419#_c_1098_n 0.0248646f $X=6.48 $Y=2.035
+ $X2=0 $Y2=0
cc_613 N_A_1195_424#_c_803_n N_A_372_419#_c_1099_n 0.0189311f $X=8.255 $Y=2.035
+ $X2=0 $Y2=0
cc_614 N_A_1195_424#_c_803_n N_A_372_419#_c_1100_n 0.00661589f $X=8.255 $Y=2.035
+ $X2=0 $Y2=0
cc_615 N_A_1195_424#_c_804_n N_A_372_419#_c_1100_n 0.00116189f $X=6.625 $Y=2.035
+ $X2=0 $Y2=0
cc_616 N_A_1195_424#_c_798_n N_A_372_419#_c_1100_n 0.0117673f $X=6.48 $Y=2.035
+ $X2=0 $Y2=0
cc_617 N_A_1195_424#_M1004_d N_A_416_113#_c_1235_n 0.00152064f $X=6.23 $Y=0.535
+ $X2=0 $Y2=0
cc_618 N_A_1195_424#_c_795_n N_A_416_113#_c_1235_n 0.0138486f $X=6.62 $Y=1.1
+ $X2=0 $Y2=0
cc_619 N_A_1195_424#_c_796_n N_A_416_113#_c_1235_n 0.00129791f $X=6.527 $Y=1.525
+ $X2=0 $Y2=0
cc_620 N_A_1195_424#_M1004_d N_A_416_113#_c_1291_n 0.00304149f $X=6.23 $Y=0.535
+ $X2=0 $Y2=0
cc_621 N_A_1195_424#_c_795_n N_A_416_113#_c_1291_n 0.00577431f $X=6.62 $Y=1.1
+ $X2=0 $Y2=0
cc_622 N_A_1195_424#_M1004_d N_A_416_113#_c_1292_n 8.211e-19 $X=6.23 $Y=0.535
+ $X2=0 $Y2=0
cc_623 N_A_1195_424#_M1004_d N_A_416_113#_c_1238_n 0.00779558f $X=6.23 $Y=0.535
+ $X2=0 $Y2=0
cc_624 N_A_1195_424#_c_795_n N_A_416_113#_c_1238_n 0.0134906f $X=6.62 $Y=1.1
+ $X2=0 $Y2=0
cc_625 N_A_1195_424#_c_796_n N_A_416_113#_c_1238_n 0.00575786f $X=6.527 $Y=1.525
+ $X2=0 $Y2=0
cc_626 N_A_1195_424#_c_799_n X 0.0157512f $X=8.645 $Y=1.765 $X2=0 $Y2=0
cc_627 N_A_1195_424#_M1002_g X 0.0188787f $X=8.655 $Y=0.76 $X2=0 $Y2=0
cc_628 N_A_1195_424#_c_789_n X 0.008373f $X=9.005 $Y=1.395 $X2=0 $Y2=0
cc_629 N_A_1195_424#_c_790_n X 0.0113269f $X=9.095 $Y=1.675 $X2=0 $Y2=0
cc_630 N_A_1195_424#_M1014_g X 0.0192976f $X=9.085 $Y=0.76 $X2=0 $Y2=0
cc_631 N_A_1195_424#_c_801_n X 0.0221058f $X=9.095 $Y=1.765 $X2=0 $Y2=0
cc_632 N_A_1195_424#_c_793_n X 0.0108716f $X=8.645 $Y=1.542 $X2=0 $Y2=0
cc_633 N_A_1195_424#_c_794_n X 0.00663376f $X=9.095 $Y=1.395 $X2=0 $Y2=0
cc_634 N_A_1195_424#_c_797_n X 0.0506711f $X=8.36 $Y=1.485 $X2=0 $Y2=0
cc_635 N_A_1195_424#_c_849_p X 0.00732723f $X=8.4 $Y=2.035 $X2=0 $Y2=0
cc_636 N_A_1195_424#_M1002_g N_VGND_c_1379_n 0.00969831f $X=8.655 $Y=0.76 $X2=0
+ $Y2=0
cc_637 N_A_1195_424#_c_792_n N_VGND_c_1379_n 0.0029613f $X=8.555 $Y=1.485 $X2=0
+ $Y2=0
cc_638 N_A_1195_424#_c_797_n N_VGND_c_1379_n 0.0278705f $X=8.36 $Y=1.485 $X2=0
+ $Y2=0
cc_639 N_A_1195_424#_M1014_g N_VGND_c_1381_n 0.00650727f $X=9.085 $Y=0.76 $X2=0
+ $Y2=0
cc_640 N_A_1195_424#_M1002_g N_VGND_c_1384_n 0.00537471f $X=8.655 $Y=0.76 $X2=0
+ $Y2=0
cc_641 N_A_1195_424#_M1014_g N_VGND_c_1384_n 0.00537471f $X=9.085 $Y=0.76 $X2=0
+ $Y2=0
cc_642 N_A_1195_424#_M1002_g N_VGND_c_1389_n 0.00539454f $X=8.655 $Y=0.76 $X2=0
+ $Y2=0
cc_643 N_A_1195_424#_M1014_g N_VGND_c_1389_n 0.00539454f $X=9.085 $Y=0.76 $X2=0
+ $Y2=0
cc_644 N_A_27_134#_c_913_n N_VPWR_c_988_n 0.0286637f $X=0.43 $Y=2.425 $X2=0
+ $Y2=0
cc_645 N_A_27_134#_c_913_n N_VPWR_c_994_n 0.0205784f $X=0.43 $Y=2.425 $X2=0
+ $Y2=0
cc_646 N_A_27_134#_c_913_n N_VPWR_c_987_n 0.0184744f $X=0.43 $Y=2.425 $X2=0
+ $Y2=0
cc_647 N_A_27_134#_c_904_n N_A_372_419#_c_1095_n 0.00838799f $X=2.35 $Y=1.48
+ $X2=0 $Y2=0
cc_648 N_A_27_134#_c_905_n N_A_372_419#_c_1095_n 0.00491286f $X=1.965 $Y=1.48
+ $X2=0 $Y2=0
cc_649 N_A_27_134#_c_906_n N_A_372_419#_c_1095_n 0.0127976f $X=2.515 $Y=2.275
+ $X2=0 $Y2=0
cc_650 N_A_27_134#_M1015_d N_A_372_419#_c_1096_n 0.00356186f $X=2.365 $Y=2.095
+ $X2=0 $Y2=0
cc_651 N_A_27_134#_c_906_n N_A_372_419#_c_1096_n 0.0171814f $X=2.515 $Y=2.275
+ $X2=0 $Y2=0
cc_652 N_A_27_134#_c_903_n N_A_416_113#_c_1232_n 0.0140676f $X=1.88 $Y=1.395
+ $X2=0 $Y2=0
cc_653 N_A_27_134#_c_904_n N_A_416_113#_c_1232_n 0.0141889f $X=2.35 $Y=1.48
+ $X2=0 $Y2=0
cc_654 N_A_27_134#_c_911_n N_A_416_113#_c_1232_n 0.0296524f $X=2.79 $Y=0.995
+ $X2=0 $Y2=0
cc_655 N_A_27_134#_M1008_d N_A_416_113#_c_1233_n 0.00913335f $X=2.58 $Y=0.785
+ $X2=0 $Y2=0
cc_656 N_A_27_134#_c_911_n N_A_416_113#_c_1233_n 0.0277569f $X=2.79 $Y=0.995
+ $X2=0 $Y2=0
cc_657 N_A_27_134#_c_906_n N_A_416_113#_c_1261_n 0.00133559f $X=2.515 $Y=2.275
+ $X2=0 $Y2=0
cc_658 N_A_27_134#_c_906_n N_A_416_113#_c_1244_n 0.0341592f $X=2.515 $Y=2.275
+ $X2=0 $Y2=0
cc_659 N_A_27_134#_c_906_n N_A_416_113#_c_1239_n 0.0132323f $X=2.515 $Y=2.275
+ $X2=0 $Y2=0
cc_660 N_A_27_134#_c_907_n N_A_416_113#_c_1239_n 0.00752401f $X=2.595 $Y=1.395
+ $X2=0 $Y2=0
cc_661 N_A_27_134#_c_910_n N_A_416_113#_c_1239_n 0.00844652f $X=2.515 $Y=1.48
+ $X2=0 $Y2=0
cc_662 N_A_27_134#_c_911_n N_A_416_113#_c_1239_n 0.0194534f $X=2.79 $Y=0.995
+ $X2=0 $Y2=0
cc_663 N_A_27_134#_c_902_n N_VGND_M1017_d 0.02171f $X=1.795 $Y=0.745 $X2=-0.19
+ $Y2=-0.245
cc_664 N_A_27_134#_c_902_n N_VGND_c_1382_n 0.0125374f $X=1.795 $Y=0.745 $X2=0
+ $Y2=0
cc_665 N_A_27_134#_c_900_n N_VGND_c_1385_n 0.00698834f $X=0.265 $Y=0.83 $X2=0
+ $Y2=0
cc_666 N_A_27_134#_c_902_n N_VGND_c_1385_n 0.00286374f $X=1.795 $Y=0.745 $X2=0
+ $Y2=0
cc_667 N_A_27_134#_c_902_n N_VGND_c_1386_n 0.0436747f $X=1.795 $Y=0.745 $X2=0
+ $Y2=0
cc_668 N_A_27_134#_c_900_n N_VGND_c_1389_n 0.0107515f $X=0.265 $Y=0.83 $X2=0
+ $Y2=0
cc_669 N_A_27_134#_c_902_n N_VGND_c_1389_n 0.0288798f $X=1.795 $Y=0.745 $X2=0
+ $Y2=0
cc_670 N_VPWR_c_997_n N_A_416_113#_c_1242_n 0.019279f $X=7.975 $Y=3.33 $X2=0
+ $Y2=0
cc_671 N_VPWR_c_987_n N_A_416_113#_c_1242_n 0.0159246f $X=9.36 $Y=3.33 $X2=0
+ $Y2=0
cc_672 N_VPWR_M1011_d N_A_416_113#_c_1243_n 0.00323229f $X=4.965 $Y=1.84 $X2=0
+ $Y2=0
cc_673 N_VPWR_c_989_n N_A_416_113#_c_1243_n 0.0239351f $X=5.115 $Y=1.985 $X2=0
+ $Y2=0
cc_674 N_VPWR_c_989_n N_A_416_113#_c_1245_n 0.00263503f $X=5.115 $Y=1.985 $X2=0
+ $Y2=0
cc_675 N_VPWR_c_989_n N_A_416_113#_c_1246_n 0.0726101f $X=5.115 $Y=1.985 $X2=0
+ $Y2=0
cc_676 N_VPWR_c_989_n N_A_416_113#_c_1240_n 0.00496387f $X=5.115 $Y=1.985 $X2=0
+ $Y2=0
cc_677 N_VPWR_c_990_n X 0.00491762f $X=8.06 $Y=1.985 $X2=0 $Y2=0
cc_678 N_VPWR_c_991_n X 0.0250331f $X=8.252 $Y=3.245 $X2=0 $Y2=0
cc_679 N_VPWR_c_993_n X 0.0778383f $X=9.32 $Y=1.985 $X2=0 $Y2=0
cc_680 N_VPWR_c_998_n X 0.014552f $X=9.235 $Y=3.33 $X2=0 $Y2=0
cc_681 N_VPWR_c_987_n X 0.0119791f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_682 N_VPWR_c_993_n N_VGND_c_1381_n 0.00814581f $X=9.32 $Y=1.985 $X2=0 $Y2=0
cc_683 N_A_372_419#_c_1096_n N_A_416_113#_M1021_d 0.00581781f $X=3.385 $Y=2.65
+ $X2=0 $Y2=0
cc_684 N_A_372_419#_c_1085_n N_A_416_113#_c_1233_n 0.0135079f $X=3.47 $Y=0.71
+ $X2=0 $Y2=0
cc_685 N_A_372_419#_c_1096_n N_A_416_113#_c_1241_n 0.0210759f $X=3.385 $Y=2.65
+ $X2=0 $Y2=0
cc_686 N_A_372_419#_M1004_s N_A_416_113#_c_1235_n 0.00315345f $X=5.805 $Y=0.535
+ $X2=0 $Y2=0
cc_687 N_A_372_419#_c_1088_n N_A_416_113#_c_1235_n 0.00707829f $X=5.775 $Y=0.76
+ $X2=0 $Y2=0
cc_688 N_A_372_419#_c_1089_n N_A_416_113#_c_1235_n 0.0200365f $X=5.9 $Y=0.675
+ $X2=0 $Y2=0
cc_689 N_A_372_419#_c_1090_n N_A_416_113#_c_1235_n 0.00363379f $X=7.435 $Y=0.34
+ $X2=0 $Y2=0
cc_690 N_A_372_419#_c_1088_n N_A_416_113#_c_1236_n 0.0142807f $X=5.775 $Y=0.76
+ $X2=0 $Y2=0
cc_691 N_A_372_419#_c_1090_n N_A_416_113#_c_1292_n 0.0105973f $X=7.435 $Y=0.34
+ $X2=0 $Y2=0
cc_692 N_A_372_419#_c_1093_n N_A_416_113#_c_1237_n 0.0270814f $X=7.52 $Y=1.095
+ $X2=0 $Y2=0
cc_693 N_A_372_419#_c_1090_n N_A_416_113#_c_1238_n 0.0644024f $X=7.435 $Y=0.34
+ $X2=0 $Y2=0
cc_694 N_A_372_419#_c_1096_n N_A_416_113#_c_1243_n 0.00348341f $X=3.385 $Y=2.65
+ $X2=0 $Y2=0
cc_695 N_A_372_419#_c_1085_n N_A_416_113#_c_1243_n 0.0188093f $X=3.47 $Y=0.71
+ $X2=0 $Y2=0
cc_696 N_A_372_419#_c_1096_n N_A_416_113#_c_1261_n 0.00259918f $X=3.385 $Y=2.65
+ $X2=0 $Y2=0
cc_697 N_A_372_419#_c_1085_n N_A_416_113#_c_1261_n 0.00237204f $X=3.47 $Y=0.71
+ $X2=0 $Y2=0
cc_698 N_A_372_419#_c_1085_n N_A_416_113#_c_1239_n 0.112445f $X=3.47 $Y=0.71
+ $X2=0 $Y2=0
cc_699 N_A_372_419#_c_1086_n N_VGND_M1009_d 0.00247003f $X=4.975 $Y=0.34 $X2=0
+ $Y2=0
cc_700 N_A_372_419#_c_1136_n N_VGND_M1009_d 0.00410163f $X=5.06 $Y=0.675 $X2=0
+ $Y2=0
cc_701 N_A_372_419#_c_1088_n N_VGND_M1009_d 0.0200041f $X=5.775 $Y=0.76 $X2=0
+ $Y2=0
cc_702 N_A_372_419#_c_1140_n N_VGND_M1009_d 9.76702e-19 $X=5.145 $Y=0.76 $X2=0
+ $Y2=0
cc_703 N_A_372_419#_c_1086_n N_VGND_c_1378_n 0.0141996f $X=4.975 $Y=0.34 $X2=0
+ $Y2=0
cc_704 N_A_372_419#_c_1136_n N_VGND_c_1378_n 0.00594708f $X=5.06 $Y=0.675 $X2=0
+ $Y2=0
cc_705 N_A_372_419#_c_1088_n N_VGND_c_1378_n 0.0192217f $X=5.775 $Y=0.76 $X2=0
+ $Y2=0
cc_706 N_A_372_419#_c_1089_n N_VGND_c_1378_n 0.00547381f $X=5.9 $Y=0.675 $X2=0
+ $Y2=0
cc_707 N_A_372_419#_c_1091_n N_VGND_c_1378_n 0.0127057f $X=6.025 $Y=0.34 $X2=0
+ $Y2=0
cc_708 N_A_372_419#_c_1090_n N_VGND_c_1379_n 0.00418126f $X=7.435 $Y=0.34 $X2=0
+ $Y2=0
cc_709 N_A_372_419#_c_1086_n N_VGND_c_1382_n 0.102488f $X=4.975 $Y=0.34 $X2=0
+ $Y2=0
cc_710 N_A_372_419#_c_1087_n N_VGND_c_1382_n 0.0115893f $X=3.555 $Y=0.34 $X2=0
+ $Y2=0
cc_711 N_A_372_419#_c_1088_n N_VGND_c_1382_n 0.00270711f $X=5.775 $Y=0.76 $X2=0
+ $Y2=0
cc_712 N_A_372_419#_c_1088_n N_VGND_c_1383_n 0.00350729f $X=5.775 $Y=0.76 $X2=0
+ $Y2=0
cc_713 N_A_372_419#_c_1090_n N_VGND_c_1383_n 0.102958f $X=7.435 $Y=0.34 $X2=0
+ $Y2=0
cc_714 N_A_372_419#_c_1091_n N_VGND_c_1383_n 0.0177305f $X=6.025 $Y=0.34 $X2=0
+ $Y2=0
cc_715 N_A_372_419#_c_1086_n N_VGND_c_1389_n 0.0553628f $X=4.975 $Y=0.34 $X2=0
+ $Y2=0
cc_716 N_A_372_419#_c_1087_n N_VGND_c_1389_n 0.00583135f $X=3.555 $Y=0.34 $X2=0
+ $Y2=0
cc_717 N_A_372_419#_c_1088_n N_VGND_c_1389_n 0.0116289f $X=5.775 $Y=0.76 $X2=0
+ $Y2=0
cc_718 N_A_372_419#_c_1090_n N_VGND_c_1389_n 0.0596141f $X=7.435 $Y=0.34 $X2=0
+ $Y2=0
cc_719 N_A_372_419#_c_1091_n N_VGND_c_1389_n 0.00968346f $X=6.025 $Y=0.34 $X2=0
+ $Y2=0
cc_720 N_A_416_113#_c_1236_n N_VGND_M1009_d 0.00213745f $X=5.68 $Y=1.1 $X2=0
+ $Y2=0
cc_721 N_A_416_113#_c_1233_n N_VGND_c_1382_n 0.0284116f $X=3.045 $Y=0.51 $X2=0
+ $Y2=0
cc_722 N_A_416_113#_c_1234_n N_VGND_c_1382_n 0.00581481f $X=2.305 $Y=0.51 $X2=0
+ $Y2=0
cc_723 N_A_416_113#_c_1233_n N_VGND_c_1389_n 0.0270015f $X=3.045 $Y=0.51 $X2=0
+ $Y2=0
cc_724 N_A_416_113#_c_1234_n N_VGND_c_1389_n 0.00530552f $X=2.305 $Y=0.51 $X2=0
+ $Y2=0
cc_725 X N_VGND_c_1379_n 0.0308484f $X=8.795 $Y=0.47 $X2=0 $Y2=0
cc_726 X N_VGND_c_1381_n 0.0294122f $X=8.795 $Y=0.47 $X2=0 $Y2=0
cc_727 X N_VGND_c_1384_n 0.0134077f $X=8.795 $Y=0.47 $X2=0 $Y2=0
cc_728 X N_VGND_c_1389_n 0.0119261f $X=8.795 $Y=0.47 $X2=0 $Y2=0
