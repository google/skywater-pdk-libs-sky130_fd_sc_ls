* File: sky130_fd_sc_ls__sedfxtp_2.spice
* Created: Fri Aug 28 14:07:33 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__sedfxtp_2.pex.spice"
.subckt sky130_fd_sc_ls__sedfxtp_2  VNB VPB D DE SCD SCE CLK VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* CLK	CLK
* SCE	SCE
* SCD	SCD
* DE	DE
* D	D
* VPB	VPB
* VNB	VNB
MM1005 A_138_74# N_D_M1005_g N_A_40_464#_M1005_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1029 N_VGND_M1029_d N_DE_M1029_g A_138_74# VNB NSHORT L=0.15 W=0.42 AD=0.1197
+ AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.6 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1013 N_VGND_M1013_d N_DE_M1013_g N_A_180_290#_M1013_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75001.7
+ A=0.063 P=1.14 MULT=1
MM1015 A_500_113# N_A_180_290#_M1015_g N_VGND_M1013_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0588 PD=0.66 PS=0.7 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1025 N_A_40_464#_M1025_d N_A_548_87#_M1025_g A_500_113# VNB NSHORT L=0.15
+ W=0.42 AD=0.08925 AS=0.0504 PD=0.845 PS=0.66 NRD=19.992 NRS=18.564 M=1 R=2.8
+ SA=75001 SB=75000.9 A=0.063 P=1.14 MULT=1
MM1026 N_A_693_113#_M1026_d N_A_663_87#_M1026_g N_A_40_464#_M1025_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.1491 AS=0.08925 PD=1.55 PS=0.845 NRD=19.992 NRS=21.42 M=1
+ R=2.8 SA=75001.6 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1031 N_VGND_M1031_d N_SCE_M1031_g N_A_663_87#_M1031_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0735 AS=0.1197 PD=0.77 PS=1.41 NRD=19.992 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1041 A_1068_125# N_SCD_M1041_g N_VGND_M1031_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0735 PD=0.63 PS=0.77 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.7
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1004 N_A_693_113#_M1004_d N_SCE_M1004_g A_1068_125# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1042 N_A_1340_74#_M1042_d N_CLK_M1042_g N_VGND_M1042_s VNB NSHORT L=0.15
+ W=0.74 AD=0.2109 AS=0.2183 PD=2.05 PS=2.07 NRD=0 NRS=0.804 M=1 R=4.93333
+ SA=75000.2 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1024 N_A_1538_74#_M1024_d N_A_1340_74#_M1024_g N_VGND_M1024_s VNB NSHORT
+ L=0.15 W=0.74 AD=0.2109 AS=0.2109 PD=2.05 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1012 N_A_1736_97#_M1012_d N_A_1340_74#_M1012_g N_A_693_113#_M1012_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.1113 AS=0.1197 PD=0.95 PS=1.41 NRD=71.424 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002.3 A=0.063 P=1.14 MULT=1
MM1016 A_1872_97# N_A_1538_74#_M1016_g N_A_1736_97#_M1012_d VNB NSHORT L=0.15
+ W=0.42 AD=0.11235 AS=0.1113 PD=0.955 PS=0.95 NRD=60.708 NRS=0 M=1 R=2.8
+ SA=75000.9 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1019 N_VGND_M1019_d N_A_1979_71#_M1019_g A_1872_97# VNB NSHORT L=0.15 W=0.42
+ AD=0.139472 AS=0.11235 PD=1.00245 PS=0.955 NRD=25.704 NRS=60.708 M=1 R=2.8
+ SA=75001.6 SB=75001 A=0.063 P=1.14 MULT=1
MM1017 N_A_1979_71#_M1017_d N_A_1736_97#_M1017_g N_VGND_M1019_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.1824 AS=0.212528 PD=1.85 PS=1.52755 NRD=0 NRS=48.744 M=1
+ R=4.26667 SA=75001.7 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1039 A_2402_74# N_A_1979_71#_M1039_g N_VGND_M1039_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0672 AS=0.1824 PD=0.85 PS=1.85 NRD=9.372 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75001.9 A=0.096 P=1.58 MULT=1
MM1040 N_A_2474_74#_M1040_d N_A_1538_74#_M1040_g A_2402_74# VNB NSHORT L=0.15
+ W=0.64 AD=0.115623 AS=0.0672 PD=1.16528 PS=0.85 NRD=8.436 NRS=9.372 M=1
+ R=4.26667 SA=75000.6 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1020 A_2569_74# N_A_1340_74#_M1020_g N_A_2474_74#_M1040_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.0758774 PD=0.66 PS=0.764717 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75001 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1021 N_VGND_M1021_d N_A_548_87#_M1021_g A_2569_74# VNB NSHORT L=0.15 W=0.42
+ AD=0.20055 AS=0.0504 PD=1.375 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.4
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1023 N_A_548_87#_M1023_d N_A_2474_74#_M1023_g N_VGND_M1021_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1197 AS=0.20055 PD=1.41 PS=1.375 NRD=0 NRS=19.992 M=1 R=2.8
+ SA=75002.5 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1008 N_Q_M1008_d N_A_2474_74#_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.2627 PD=1.02 PS=2.19 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75000.3
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1036 N_Q_M1008_d N_A_2474_74#_M1036_g N_VGND_M1036_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.2627 PD=1.02 PS=2.19 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75000.7
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1009 A_129_464# N_D_M1009_g N_A_40_464#_M1009_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0864 AS=0.1888 PD=0.91 PS=1.87 NRD=24.625 NRS=3.0732 M=1 R=4.26667
+ SA=75000.2 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1034 N_VPWR_M1034_d N_A_180_290#_M1034_g A_129_464# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1888 AS=0.0864 PD=1.87 PS=0.91 NRD=3.0732 NRS=24.625 M=1 R=4.26667
+ SA=75000.6 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1038 N_VPWR_M1038_d N_DE_M1038_g N_A_180_290#_M1038_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1696 AS=0.1888 PD=1.17 PS=1.87 NRD=73.8553 NRS=3.0732 M=1
+ R=4.26667 SA=75000.2 SB=75001.7 A=0.096 P=1.58 MULT=1
MM1014 A_575_463# N_DE_M1014_g N_VPWR_M1038_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0768 AS=0.1696 PD=0.88 PS=1.17 NRD=19.9955 NRS=3.0732 M=1 R=4.26667
+ SA=75000.9 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1032 N_A_40_464#_M1032_d N_A_548_87#_M1032_g A_575_463# VPB PHIGHVT L=0.15
+ W=0.64 AD=0.096 AS=0.0768 PD=0.94 PS=0.88 NRD=3.0732 NRS=19.9955 M=1 R=4.26667
+ SA=75001.3 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1002 N_A_693_113#_M1002_d N_SCE_M1002_g N_A_40_464#_M1032_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1856 AS=0.096 PD=1.86 PS=0.94 NRD=3.0732 NRS=3.0732 M=1 R=4.26667
+ SA=75001.7 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1003 N_VPWR_M1003_d N_SCE_M1003_g N_A_663_87#_M1003_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1696 AS=0.1856 PD=1.17 PS=1.86 NRD=73.8553 NRS=3.0732 M=1
+ R=4.26667 SA=75000.2 SB=75001.3 A=0.096 P=1.58 MULT=1
MM1018 A_1079_455# N_SCD_M1018_g N_VPWR_M1003_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0864 AS=0.1696 PD=0.91 PS=1.17 NRD=24.625 NRS=3.0732 M=1 R=4.26667
+ SA=75000.9 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1010 N_A_693_113#_M1010_d N_A_663_87#_M1010_g A_1079_455# VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1888 AS=0.0864 PD=1.87 PS=0.91 NRD=3.0732 NRS=24.625 M=1 R=4.26667
+ SA=75001.3 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1011 N_A_1340_74#_M1011_d N_CLK_M1011_g N_VPWR_M1011_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.3304 AS=0.336 PD=2.83 PS=2.84 NRD=1.7533 NRS=2.6201 M=1 R=7.46667
+ SA=75000.2 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1033 N_A_1538_74#_M1033_d N_A_1340_74#_M1033_g N_VPWR_M1033_s VPB PHIGHVT
+ L=0.15 W=1.12 AD=0.3304 AS=0.3304 PD=2.83 PS=2.83 NRD=1.7533 NRS=1.7533 M=1
+ R=7.46667 SA=75000.2 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1000 N_A_1736_97#_M1000_d N_A_1538_74#_M1000_g N_A_693_113#_M1000_s VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.063 AS=0.1239 PD=0.72 PS=1.43 NRD=4.6886 NRS=4.6886
+ M=1 R=2.8 SA=75000.2 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1007 A_1936_508# N_A_1340_74#_M1007_g N_A_1736_97#_M1000_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.084 AS=0.063 PD=0.82 PS=0.72 NRD=68.0044 NRS=4.6886 M=1 R=2.8
+ SA=75000.7 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1001 N_VPWR_M1001_d N_A_1979_71#_M1001_g A_1936_508# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0985833 AS=0.084 PD=0.903333 PS=0.82 NRD=4.6886 NRS=68.0044 M=1 R=2.8
+ SA=75001.2 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1030 N_A_1979_71#_M1030_d N_A_1736_97#_M1030_g N_VPWR_M1001_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.2478 AS=0.197167 PD=2.27 PS=1.80667 NRD=2.3443 NRS=23.443
+ M=1 R=5.6 SA=75000.7 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1028 A_2357_392# N_A_1979_71#_M1028_g N_VPWR_M1028_s VPB PHIGHVT L=0.15 W=1
+ AD=0.405 AS=0.305 PD=1.81 PS=2.61 NRD=68.9303 NRS=2.9353 M=1 R=6.66667
+ SA=75000.2 SB=75001.9 A=0.15 P=2.3 MULT=1
MM1043 N_A_2474_74#_M1043_d N_A_1340_74#_M1043_g A_2357_392# VPB PHIGHVT L=0.15
+ W=1 AD=0.223592 AS=0.405 PD=1.95775 PS=1.81 NRD=19.7 NRS=68.9303 M=1 R=6.66667
+ SA=75001.2 SB=75000.9 A=0.15 P=2.3 MULT=1
MM1006 A_2657_508# N_A_1538_74#_M1006_g N_A_2474_74#_M1043_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0567 AS=0.0939085 PD=0.69 PS=0.822254 NRD=37.5088 NRS=4.6886 M=1
+ R=2.8 SA=75001.7 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1037 N_VPWR_M1037_d N_A_548_87#_M1037_g A_2657_508# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.116292 AS=0.0567 PD=0.950943 PS=0.69 NRD=53.9386 NRS=37.5088 M=1 R=2.8
+ SA=75002.1 SB=75000.9 A=0.063 P=1.14 MULT=1
MM1035 N_A_548_87#_M1035_d N_A_2474_74#_M1035_g N_VPWR_M1037_d VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.1888 AS=0.177208 PD=1.87 PS=1.44906 NRD=3.0732 NRS=50.7866
+ M=1 R=4.26667 SA=75001.9 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1022 N_VPWR_M1022_d N_A_2474_74#_M1022_g N_Q_M1022_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.1764 PD=2.83 PS=1.435 NRD=1.7533 NRS=2.6201 M=1 R=7.46667
+ SA=75000.2 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1027 N_VPWR_M1027_d N_A_2474_74#_M1027_g N_Q_M1022_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.1764 PD=2.83 PS=1.435 NRD=1.7533 NRS=3.5066 M=1 R=7.46667
+ SA=75000.7 SB=75000.2 A=0.168 P=2.54 MULT=1
DX44_noxref VNB VPB NWDIODE A=31.0841 P=37.16
c_173 VNB 0 3.03176e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_ls__sedfxtp_2.pxi.spice"
*
.ends
*
*
