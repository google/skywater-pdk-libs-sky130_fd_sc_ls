* File: sky130_fd_sc_ls__nand4b_2.spice
* Created: Fri Aug 28 13:35:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__nand4b_2.pex.spice"
.subckt sky130_fd_sc_ls__nand4b_2  VNB VPB A_N B C D VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* D	D
* C	C
* B	B
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1015 N_VGND_M1015_d N_A_N_M1015_g N_A_27_74#_M1015_s VNB NSHORT L=0.15 W=0.64
+ AD=0.1726 AS=0.1824 PD=1.85 PS=1.85 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1007 N_A_225_74#_M1007_d N_A_27_74#_M1007_g N_Y_M1007_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1962 AS=0.1147 PD=2.05 PS=1.05 NRD=0 NRS=2.424 M=1 R=4.93333
+ SA=75000.2 SB=75001.7 A=0.111 P=1.78 MULT=1
MM1017 N_A_225_74#_M1017_d N_A_27_74#_M1017_g N_Y_M1007_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1147 PD=1.02 PS=1.05 NRD=0 NRS=2.424 M=1 R=4.93333
+ SA=75000.7 SB=75001.2 A=0.111 P=1.78 MULT=1
MM1002 N_A_225_74#_M1017_d N_B_M1002_g N_A_490_74#_M1002_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1773 PD=1.02 PS=1.28 NRD=0 NRS=13.776 M=1 R=4.93333
+ SA=75001.1 SB=75000.8 A=0.111 P=1.78 MULT=1
MM1013 N_A_225_74#_M1013_d N_B_M1013_g N_A_490_74#_M1002_s VNB NSHORT L=0.15
+ W=0.74 AD=0.197775 AS=0.1773 PD=2.05 PS=1.28 NRD=0 NRS=13.776 M=1 R=4.93333
+ SA=75001.7 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1000 N_A_719_123#_M1000_d N_C_M1000_g N_A_490_74#_M1000_s VNB NSHORT L=0.15
+ W=0.74 AD=0.204075 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001.5 A=0.111 P=1.78 MULT=1
MM1012 N_A_719_123#_M1012_d N_C_M1012_g N_A_490_74#_M1000_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1009 N_A_719_123#_M1012_d N_D_M1009_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.111 PD=1.02 PS=1.04 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1010 N_A_719_123#_M1010_d N_D_M1010_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.111 PD=2.05 PS=1.04 NRD=0 NRS=3.24 M=1 R=4.93333 SA=75001.5
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1014 N_VPWR_M1014_d N_A_N_M1014_g N_A_27_74#_M1014_s VPB PHIGHVT L=0.15 W=1
+ AD=0.200943 AS=0.295 PD=1.42453 PS=2.59 NRD=19.0302 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75004.6 A=0.15 P=2.3 MULT=1
MM1003 N_Y_M1003_d N_A_27_74#_M1003_g N_VPWR_M1014_d VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.225057 PD=1.42 PS=1.59547 NRD=1.7533 NRS=2.6201 M=1 R=7.46667
+ SA=75000.7 SB=75004 A=0.168 P=2.54 MULT=1
MM1006 N_Y_M1003_d N_A_27_74#_M1006_g N_VPWR_M1006_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.3724 PD=1.42 PS=1.785 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.2 SB=75003.6 A=0.168 P=2.54 MULT=1
MM1011 N_Y_M1011_d N_B_M1011_g N_VPWR_M1006_s VPB PHIGHVT L=0.15 W=1.12 AD=0.168
+ AS=0.3724 PD=1.42 PS=1.785 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75002
+ SB=75002.8 A=0.168 P=2.54 MULT=1
MM1016 N_Y_M1011_d N_B_M1016_g N_VPWR_M1016_s VPB PHIGHVT L=0.15 W=1.12 AD=0.168
+ AS=0.224 PD=1.42 PS=1.52 NRD=1.7533 NRS=10.5395 M=1 R=7.46667 SA=75002.4
+ SB=75002.3 A=0.168 P=2.54 MULT=1
MM1001 N_Y_M1001_d N_C_M1001_g N_VPWR_M1016_s VPB PHIGHVT L=0.15 W=1.12 AD=0.168
+ AS=0.224 PD=1.42 PS=1.52 NRD=1.7533 NRS=10.5395 M=1 R=7.46667 SA=75003
+ SB=75001.8 A=0.168 P=2.54 MULT=1
MM1004 N_Y_M1001_d N_C_M1004_g N_VPWR_M1004_s VPB PHIGHVT L=0.15 W=1.12 AD=0.168
+ AS=0.28 PD=1.42 PS=1.62 NRD=1.7533 NRS=21.0987 M=1 R=7.46667 SA=75003.4
+ SB=75001.3 A=0.168 P=2.54 MULT=1
MM1005 N_Y_M1005_d N_D_M1005_g N_VPWR_M1004_s VPB PHIGHVT L=0.15 W=1.12 AD=0.168
+ AS=0.28 PD=1.42 PS=1.62 NRD=1.7533 NRS=17.5724 M=1 R=7.46667 SA=75004.1
+ SB=75000.7 A=0.168 P=2.54 MULT=1
MM1008 N_Y_M1005_d N_D_M1008_g N_VPWR_M1008_s VPB PHIGHVT L=0.15 W=1.12 AD=0.168
+ AS=0.336 PD=1.42 PS=2.84 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75004.5
+ SB=75000.2 A=0.168 P=2.54 MULT=1
DX18_noxref VNB VPB NWDIODE A=11.4204 P=16
*
.include "sky130_fd_sc_ls__nand4b_2.pxi.spice"
*
.ends
*
*
