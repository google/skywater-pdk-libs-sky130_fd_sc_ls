* File: sky130_fd_sc_ls__nand2_1.pxi.spice
* Created: Wed Sep  2 11:11:14 2020
* 
x_PM_SKY130_FD_SC_LS__NAND2_1%B N_B_c_25_n N_B_M1001_g N_B_c_26_n N_B_M1003_g B
+ PM_SKY130_FD_SC_LS__NAND2_1%B
x_PM_SKY130_FD_SC_LS__NAND2_1%A N_A_c_48_n N_A_M1000_g N_A_c_49_n N_A_M1002_g A
+ PM_SKY130_FD_SC_LS__NAND2_1%A
x_PM_SKY130_FD_SC_LS__NAND2_1%VPWR N_VPWR_M1001_s N_VPWR_M1002_d N_VPWR_c_72_n
+ N_VPWR_c_73_n N_VPWR_c_74_n N_VPWR_c_75_n VPWR N_VPWR_c_76_n N_VPWR_c_71_n
+ PM_SKY130_FD_SC_LS__NAND2_1%VPWR
x_PM_SKY130_FD_SC_LS__NAND2_1%Y N_Y_M1000_d N_Y_M1001_d N_Y_c_92_n N_Y_c_93_n Y
+ Y Y Y Y Y N_Y_c_95_n PM_SKY130_FD_SC_LS__NAND2_1%Y
x_PM_SKY130_FD_SC_LS__NAND2_1%VGND N_VGND_M1003_s N_VGND_c_122_n N_VGND_c_123_n
+ VGND N_VGND_c_124_n N_VGND_c_125_n PM_SKY130_FD_SC_LS__NAND2_1%VGND
cc_1 VNB N_B_c_25_n 0.0675637f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.765
cc_2 VNB N_B_c_26_n 0.0207038f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.22
cc_3 VNB B 0.00878284f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_A_c_48_n 0.0221784f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.765
cc_5 VNB N_A_c_49_n 0.0688437f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.22
cc_6 VNB A 0.0096067f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_7 VNB N_VPWR_c_71_n 0.0641695f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_Y_c_92_n 0.0070579f $X=-0.19 $Y=-0.245 $X2=0.345 $Y2=1.385
cc_9 VNB N_Y_c_93_n 0.0213168f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_10 VNB Y 0.00714178f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_Y_c_95_n 6.31494e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_VGND_c_122_n 0.0125057f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.22
cc_13 VNB N_VGND_c_123_n 0.0344105f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.74
cc_14 VNB N_VGND_c_124_n 0.0306085f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.295
cc_15 VNB N_VGND_c_125_n 0.119298f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VPB N_B_c_25_n 0.0291926f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.765
cc_17 VPB N_A_c_49_n 0.0291926f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.22
cc_18 VPB N_VPWR_c_72_n 0.0116916f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_19 VPB N_VPWR_c_73_n 0.0555647f $X=-0.19 $Y=1.66 $X2=0.345 $Y2=1.385
cc_20 VPB N_VPWR_c_74_n 0.0116916f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_21 VPB N_VPWR_c_75_n 0.0555647f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_22 VPB N_VPWR_c_76_n 0.0159778f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_23 VPB N_VPWR_c_71_n 0.0485419f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_24 VPB Y 0.00649418f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_25 N_B_c_26_n N_A_c_48_n 0.0329441f $X=0.51 $Y=1.22 $X2=-0.19 $Y2=-0.245
cc_26 N_B_c_25_n N_A_c_49_n 0.0497587f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_27 B N_A_c_49_n 2.30773e-19 $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_28 N_B_c_25_n N_VPWR_c_73_n 0.0201717f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_29 B N_VPWR_c_73_n 0.0197435f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_30 N_B_c_25_n N_VPWR_c_75_n 6.29256e-19 $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_31 N_B_c_25_n N_VPWR_c_76_n 0.00413917f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_32 N_B_c_25_n N_VPWR_c_71_n 0.0081781f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_33 N_B_c_26_n N_Y_c_92_n 0.00129102f $X=0.51 $Y=1.22 $X2=0 $Y2=0
cc_34 N_B_c_26_n N_Y_c_93_n 0.00138696f $X=0.51 $Y=1.22 $X2=0 $Y2=0
cc_35 N_B_c_25_n Y 0.00633977f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_36 N_B_c_26_n Y 0.00436559f $X=0.51 $Y=1.22 $X2=0 $Y2=0
cc_37 B Y 0.0285816f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_38 N_B_c_26_n N_Y_c_95_n 0.00382427f $X=0.51 $Y=1.22 $X2=0 $Y2=0
cc_39 N_B_c_25_n N_VGND_c_123_n 0.0019927f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_40 N_B_c_26_n N_VGND_c_123_n 0.0166171f $X=0.51 $Y=1.22 $X2=0 $Y2=0
cc_41 B N_VGND_c_123_n 0.0241219f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_42 N_B_c_26_n N_VGND_c_124_n 0.00383152f $X=0.51 $Y=1.22 $X2=0 $Y2=0
cc_43 N_B_c_26_n N_VGND_c_125_n 0.0075725f $X=0.51 $Y=1.22 $X2=0 $Y2=0
cc_44 N_A_c_49_n N_VPWR_c_73_n 6.29256e-19 $X=0.945 $Y=1.765 $X2=0 $Y2=0
cc_45 N_A_c_49_n N_VPWR_c_75_n 0.0201717f $X=0.945 $Y=1.765 $X2=0 $Y2=0
cc_46 A N_VPWR_c_75_n 0.0197435f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_47 N_A_c_49_n N_VPWR_c_76_n 0.00413917f $X=0.945 $Y=1.765 $X2=0 $Y2=0
cc_48 N_A_c_49_n N_VPWR_c_71_n 0.0081781f $X=0.945 $Y=1.765 $X2=0 $Y2=0
cc_49 N_A_c_48_n N_Y_c_92_n 0.0126998f $X=0.9 $Y=1.22 $X2=0 $Y2=0
cc_50 N_A_c_49_n N_Y_c_92_n 0.00167291f $X=0.945 $Y=1.765 $X2=0 $Y2=0
cc_51 A N_Y_c_92_n 0.0207374f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_52 N_A_c_48_n N_Y_c_93_n 0.00922372f $X=0.9 $Y=1.22 $X2=0 $Y2=0
cc_53 N_A_c_48_n Y 6.89533e-19 $X=0.9 $Y=1.22 $X2=0 $Y2=0
cc_54 N_A_c_49_n Y 0.0153569f $X=0.945 $Y=1.765 $X2=0 $Y2=0
cc_55 A Y 0.0271114f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_56 N_A_c_48_n N_Y_c_95_n 0.00776809f $X=0.9 $Y=1.22 $X2=0 $Y2=0
cc_57 N_A_c_48_n N_VGND_c_123_n 0.00208984f $X=0.9 $Y=1.22 $X2=0 $Y2=0
cc_58 N_A_c_48_n N_VGND_c_124_n 0.00434272f $X=0.9 $Y=1.22 $X2=0 $Y2=0
cc_59 N_A_c_48_n N_VGND_c_125_n 0.00451209f $X=0.9 $Y=1.22 $X2=0 $Y2=0
cc_60 N_VPWR_c_73_n Y 0.0450228f $X=0.27 $Y=1.985 $X2=0 $Y2=0
cc_61 N_VPWR_c_75_n Y 0.0450228f $X=1.17 $Y=1.985 $X2=0 $Y2=0
cc_62 N_VPWR_c_76_n Y 0.0101736f $X=1.005 $Y=3.33 $X2=0 $Y2=0
cc_63 N_VPWR_c_71_n Y 0.0084208f $X=1.2 $Y=3.33 $X2=0 $Y2=0
cc_64 N_Y_c_92_n N_VGND_c_123_n 0.0119089f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_65 N_Y_c_93_n N_VGND_c_123_n 0.0155235f $X=1.115 $Y=0.515 $X2=0 $Y2=0
cc_66 N_Y_c_93_n N_VGND_c_124_n 0.0142249f $X=1.115 $Y=0.515 $X2=0 $Y2=0
cc_67 N_Y_c_92_n N_VGND_c_125_n 0.00901755f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_68 N_Y_c_93_n N_VGND_c_125_n 0.011867f $X=1.115 $Y=0.515 $X2=0 $Y2=0
cc_69 N_Y_c_92_n A_117_74# 0.00390405f $X=1.115 $Y=0.84 $X2=-0.19 $Y2=-0.245
cc_70 N_Y_c_95_n A_117_74# 0.00140851f $X=0.72 $Y=1.18 $X2=-0.19 $Y2=-0.245
