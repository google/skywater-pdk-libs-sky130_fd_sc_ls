* File: sky130_fd_sc_ls__a311oi_4.pxi.spice
* Created: Fri Aug 28 12:58:27 2020
* 
x_PM_SKY130_FD_SC_LS__A311OI_4%A3 N_A3_c_155_n N_A3_M1000_g N_A3_M1003_g
+ N_A3_c_156_n N_A3_M1008_g N_A3_M1018_g N_A3_M1023_g N_A3_c_157_n N_A3_M1028_g
+ N_A3_M1026_g N_A3_c_158_n N_A3_M1029_g A3 A3 A3 N_A3_c_159_n N_A3_c_154_n
+ PM_SKY130_FD_SC_LS__A311OI_4%A3
x_PM_SKY130_FD_SC_LS__A311OI_4%A2 N_A2_M1002_g N_A2_c_232_n N_A2_M1005_g
+ N_A2_M1011_g N_A2_c_233_n N_A2_M1016_g N_A2_M1033_g N_A2_c_234_n N_A2_M1024_g
+ N_A2_M1034_g N_A2_c_235_n N_A2_M1031_g A2 A2 A2 A2 N_A2_c_231_n
+ PM_SKY130_FD_SC_LS__A311OI_4%A2
x_PM_SKY130_FD_SC_LS__A311OI_4%A1 N_A1_c_318_n N_A1_M1006_g N_A1_c_310_n
+ N_A1_c_320_n N_A1_M1013_g N_A1_M1007_g N_A1_c_321_n N_A1_M1014_g N_A1_M1012_g
+ N_A1_c_322_n N_A1_M1017_g N_A1_M1021_g N_A1_M1035_g N_A1_c_315_n A1 A1
+ N_A1_c_317_n PM_SKY130_FD_SC_LS__A311OI_4%A1
x_PM_SKY130_FD_SC_LS__A311OI_4%B1 N_B1_c_400_n N_B1_M1001_g N_B1_M1010_g
+ N_B1_c_401_n N_B1_M1009_g N_B1_c_402_n N_B1_M1020_g N_B1_M1019_g N_B1_c_403_n
+ N_B1_M1027_g B1 B1 N_B1_c_398_n N_B1_c_399_n PM_SKY130_FD_SC_LS__A311OI_4%B1
x_PM_SKY130_FD_SC_LS__A311OI_4%C1 N_C1_c_472_n N_C1_M1004_g N_C1_c_479_n
+ N_C1_M1015_g N_C1_c_473_n N_C1_M1030_g N_C1_c_480_n N_C1_M1022_g N_C1_c_481_n
+ N_C1_M1025_g N_C1_c_474_n N_C1_c_475_n N_C1_c_476_n N_C1_c_484_n N_C1_M1032_g
+ C1 C1 N_C1_c_477_n N_C1_c_478_n C1 PM_SKY130_FD_SC_LS__A311OI_4%C1
x_PM_SKY130_FD_SC_LS__A311OI_4%VPWR N_VPWR_M1000_s N_VPWR_M1008_s N_VPWR_M1029_s
+ N_VPWR_M1016_d N_VPWR_M1031_d N_VPWR_M1013_d N_VPWR_M1017_d N_VPWR_c_551_n
+ N_VPWR_c_552_n N_VPWR_c_553_n N_VPWR_c_554_n N_VPWR_c_555_n N_VPWR_c_556_n
+ N_VPWR_c_557_n N_VPWR_c_558_n N_VPWR_c_559_n N_VPWR_c_560_n N_VPWR_c_561_n
+ N_VPWR_c_562_n N_VPWR_c_563_n N_VPWR_c_564_n N_VPWR_c_565_n N_VPWR_c_566_n
+ N_VPWR_c_567_n VPWR N_VPWR_c_568_n N_VPWR_c_569_n N_VPWR_c_550_n
+ N_VPWR_c_571_n N_VPWR_c_572_n PM_SKY130_FD_SC_LS__A311OI_4%VPWR
x_PM_SKY130_FD_SC_LS__A311OI_4%A_114_368# N_A_114_368#_M1000_d
+ N_A_114_368#_M1028_d N_A_114_368#_M1005_s N_A_114_368#_M1024_s
+ N_A_114_368#_M1006_s N_A_114_368#_M1014_s N_A_114_368#_M1001_d
+ N_A_114_368#_M1020_d N_A_114_368#_c_703_n N_A_114_368#_c_692_n
+ N_A_114_368#_c_708_n N_A_114_368#_c_693_n N_A_114_368#_c_714_n
+ N_A_114_368#_c_694_n N_A_114_368#_c_722_n N_A_114_368#_c_695_n
+ N_A_114_368#_c_728_n N_A_114_368#_c_696_n N_A_114_368#_c_738_n
+ N_A_114_368#_c_697_n N_A_114_368#_c_698_n N_A_114_368#_c_806_p
+ N_A_114_368#_c_699_n N_A_114_368#_c_700_n N_A_114_368#_c_809_p
+ N_A_114_368#_c_716_n N_A_114_368#_c_730_n N_A_114_368#_c_732_n
+ N_A_114_368#_c_701_n N_A_114_368#_c_752_n N_A_114_368#_c_702_n
+ PM_SKY130_FD_SC_LS__A311OI_4%A_114_368#
x_PM_SKY130_FD_SC_LS__A311OI_4%A_1213_368# N_A_1213_368#_M1001_s
+ N_A_1213_368#_M1009_s N_A_1213_368#_M1027_s N_A_1213_368#_M1022_s
+ N_A_1213_368#_M1032_s N_A_1213_368#_c_811_n N_A_1213_368#_c_812_n
+ N_A_1213_368#_c_813_n N_A_1213_368#_c_828_n N_A_1213_368#_c_814_n
+ N_A_1213_368#_c_815_n N_A_1213_368#_c_816_n N_A_1213_368#_c_846_n
+ N_A_1213_368#_c_817_n N_A_1213_368#_c_818_n N_A_1213_368#_c_819_n
+ N_A_1213_368#_c_820_n N_A_1213_368#_c_821_n
+ PM_SKY130_FD_SC_LS__A311OI_4%A_1213_368#
x_PM_SKY130_FD_SC_LS__A311OI_4%Y N_Y_M1007_s N_Y_M1012_s N_Y_M1035_s N_Y_M1019_s
+ N_Y_M1030_d N_Y_M1015_d N_Y_M1025_d N_Y_c_896_n N_Y_c_897_n N_Y_c_919_n
+ N_Y_c_898_n N_Y_c_930_n N_Y_c_904_n N_Y_c_905_n N_Y_c_899_n N_Y_c_945_n
+ N_Y_c_900_n N_Y_c_901_n N_Y_c_927_n N_Y_c_907_n Y Y Y N_Y_c_949_n Y
+ N_Y_c_903_n PM_SKY130_FD_SC_LS__A311OI_4%Y
x_PM_SKY130_FD_SC_LS__A311OI_4%A_34_74# N_A_34_74#_M1003_s N_A_34_74#_M1018_s
+ N_A_34_74#_M1026_s N_A_34_74#_M1011_s N_A_34_74#_M1034_s N_A_34_74#_c_995_n
+ N_A_34_74#_c_996_n N_A_34_74#_c_997_n N_A_34_74#_c_998_n N_A_34_74#_c_999_n
+ N_A_34_74#_c_1000_n N_A_34_74#_c_1001_n N_A_34_74#_c_1002_n
+ N_A_34_74#_c_1003_n N_A_34_74#_c_1004_n N_A_34_74#_c_1005_n
+ N_A_34_74#_c_1006_n PM_SKY130_FD_SC_LS__A311OI_4%A_34_74#
x_PM_SKY130_FD_SC_LS__A311OI_4%VGND N_VGND_M1003_d N_VGND_M1023_d N_VGND_M1010_d
+ N_VGND_M1004_s N_VGND_c_1069_n N_VGND_c_1070_n N_VGND_c_1071_n VGND
+ N_VGND_c_1072_n N_VGND_c_1073_n N_VGND_c_1074_n N_VGND_c_1075_n
+ N_VGND_c_1076_n N_VGND_c_1077_n N_VGND_c_1078_n N_VGND_c_1079_n
+ N_VGND_c_1080_n N_VGND_c_1081_n PM_SKY130_FD_SC_LS__A311OI_4%VGND
x_PM_SKY130_FD_SC_LS__A311OI_4%A_465_74# N_A_465_74#_M1002_d N_A_465_74#_M1033_d
+ N_A_465_74#_M1007_d N_A_465_74#_M1021_d N_A_465_74#_c_1158_n
+ N_A_465_74#_c_1159_n N_A_465_74#_c_1160_n N_A_465_74#_c_1161_n
+ N_A_465_74#_c_1162_n PM_SKY130_FD_SC_LS__A311OI_4%A_465_74#
cc_1 VNB N_A3_M1003_g 0.0318708f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=0.74
cc_2 VNB N_A3_M1018_g 0.0230578f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=0.74
cc_3 VNB N_A3_M1023_g 0.0224931f $X=-0.19 $Y=-0.245 $X2=1.39 $Y2=0.74
cc_4 VNB N_A3_M1026_g 0.0229868f $X=-0.19 $Y=-0.245 $X2=1.82 $Y2=0.74
cc_5 VNB N_A3_c_154_n 0.0828315f $X=-0.19 $Y=-0.245 $X2=1.82 $Y2=1.557
cc_6 VNB N_A2_M1002_g 0.0236065f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_7 VNB N_A2_M1011_g 0.0230075f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=2.4
cc_8 VNB N_A2_M1033_g 0.0230075f $X=-0.19 $Y=-0.245 $X2=1.39 $Y2=0.74
cc_9 VNB N_A2_M1034_g 0.0325857f $X=-0.19 $Y=-0.245 $X2=1.82 $Y2=0.74
cc_10 VNB A2 0.00306242f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A2_c_231_n 0.078333f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.565
cc_12 VNB N_A1_c_310_n 0.0137327f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.35
cc_13 VNB N_A1_M1007_g 0.0337355f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=1.35
cc_14 VNB N_A1_M1012_g 0.0234256f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A1_M1021_g 0.0234256f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A1_M1035_g 0.0240737f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_17 VNB N_A1_c_315_n 0.0147873f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_18 VNB A1 0.0109081f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A1_c_317_n 0.0717989f $X=-0.19 $Y=-0.245 $X2=1.82 $Y2=1.557
cc_20 VNB N_B1_M1010_g 0.0261425f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=0.74
cc_21 VNB N_B1_M1019_g 0.0259064f $X=-0.19 $Y=-0.245 $X2=1.39 $Y2=0.74
cc_22 VNB B1 0.00796405f $X=-0.19 $Y=-0.245 $X2=1.82 $Y2=1.35
cc_23 VNB N_B1_c_398_n 0.116403f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.557
cc_24 VNB N_B1_c_399_n 0.00679545f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.557
cc_25 VNB N_C1_c_472_n 0.0168861f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.765
cc_26 VNB N_C1_c_473_n 0.0210077f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_C1_c_474_n 0.0422463f $X=-0.19 $Y=-0.245 $X2=1.39 $Y2=0.74
cc_28 VNB N_C1_c_475_n 0.0882376f $X=-0.19 $Y=-0.245 $X2=1.39 $Y2=0.74
cc_29 VNB N_C1_c_476_n 0.0158274f $X=-0.19 $Y=-0.245 $X2=1.395 $Y2=1.765
cc_30 VNB N_C1_c_477_n 0.0046005f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.557
cc_31 VNB N_C1_c_478_n 0.00623501f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.515
cc_32 VNB N_VPWR_c_550_n 0.422413f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_Y_c_896_n 0.00842476f $X=-0.19 $Y=-0.245 $X2=1.82 $Y2=1.35
cc_34 VNB N_Y_c_897_n 0.00206055f $X=-0.19 $Y=-0.245 $X2=1.845 $Y2=2.4
cc_35 VNB N_Y_c_898_n 0.00206768f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_Y_c_899_n 0.0137919f $X=-0.19 $Y=-0.245 $X2=1.71 $Y2=1.515
cc_37 VNB N_Y_c_900_n 0.00967636f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.565
cc_38 VNB N_Y_c_901_n 0.00828779f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=1.565
cc_39 VNB Y 0.0381136f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_Y_c_903_n 0.0357019f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_34_74#_c_995_n 0.0266107f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_34_74#_c_996_n 0.00273425f $X=-0.19 $Y=-0.245 $X2=1.395 $Y2=2.4
cc_43 VNB N_A_34_74#_c_997_n 0.0126474f $X=-0.19 $Y=-0.245 $X2=1.395 $Y2=2.4
cc_44 VNB N_A_34_74#_c_998_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=1.82 $Y2=0.74
cc_45 VNB N_A_34_74#_c_999_n 0.0036153f $X=-0.19 $Y=-0.245 $X2=1.845 $Y2=1.765
cc_46 VNB N_A_34_74#_c_1000_n 0.00178301f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_47 VNB N_A_34_74#_c_1001_n 0.00226168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_34_74#_c_1002_n 0.00178779f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.557
cc_49 VNB N_A_34_74#_c_1003_n 0.0045734f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.557
cc_50 VNB N_A_34_74#_c_1004_n 0.00275936f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=1.557
cc_51 VNB N_A_34_74#_c_1005_n 0.00228886f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=1.557
cc_52 VNB N_A_34_74#_c_1006_n 0.0156582f $X=-0.19 $Y=-0.245 $X2=1.395 $Y2=1.557
cc_53 VNB N_VGND_c_1069_n 0.00481913f $X=-0.19 $Y=-0.245 $X2=1.39 $Y2=1.35
cc_54 VNB N_VGND_c_1070_n 0.00334323f $X=-0.19 $Y=-0.245 $X2=1.395 $Y2=1.765
cc_55 VNB N_VGND_c_1071_n 0.00332936f $X=-0.19 $Y=-0.245 $X2=1.82 $Y2=0.74
cc_56 VNB N_VGND_c_1072_n 0.0185047f $X=-0.19 $Y=-0.245 $X2=1.845 $Y2=2.4
cc_57 VNB N_VGND_c_1073_n 0.0172524f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_1074_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=1.71 $Y2=1.515
cc_59 VNB N_VGND_c_1075_n 0.0418428f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=1.565
cc_60 VNB N_VGND_c_1076_n 0.525006f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_1077_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_1078_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_1079_n 0.12018f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_1080_n 0.0364641f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_1081_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_465_74#_c_1158_n 0.00199246f $X=-0.19 $Y=-0.245 $X2=1.82 $Y2=1.35
cc_67 VNB N_A_465_74#_c_1159_n 0.00310413f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_465_74#_c_1160_n 0.00161093f $X=-0.19 $Y=-0.245 $X2=1.845
+ $Y2=1.765
cc_69 VNB N_A_465_74#_c_1161_n 0.002374f $X=-0.19 $Y=-0.245 $X2=1.845 $Y2=2.4
cc_70 VNB N_A_465_74#_c_1162_n 0.0338474f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_71 VPB N_A3_c_155_n 0.0177026f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.765
cc_72 VPB N_A3_c_156_n 0.0149991f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=1.765
cc_73 VPB N_A3_c_157_n 0.0149968f $X=-0.19 $Y=1.66 $X2=1.395 $Y2=1.765
cc_74 VPB N_A3_c_158_n 0.0151753f $X=-0.19 $Y=1.66 $X2=1.845 $Y2=1.765
cc_75 VPB N_A3_c_159_n 0.00839387f $X=-0.19 $Y=1.66 $X2=1.71 $Y2=1.515
cc_76 VPB N_A3_c_154_n 0.0503102f $X=-0.19 $Y=1.66 $X2=1.82 $Y2=1.557
cc_77 VPB N_A2_c_232_n 0.0151049f $X=-0.19 $Y=1.66 $X2=0.53 $Y2=0.74
cc_78 VPB N_A2_c_233_n 0.0149968f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=0.74
cc_79 VPB N_A2_c_234_n 0.0149968f $X=-0.19 $Y=1.66 $X2=1.395 $Y2=1.765
cc_80 VPB N_A2_c_235_n 0.0151789f $X=-0.19 $Y=1.66 $X2=1.845 $Y2=1.765
cc_81 VPB A2 0.0107416f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 VPB N_A2_c_231_n 0.04616f $X=-0.19 $Y=1.66 $X2=0.69 $Y2=1.565
cc_83 VPB N_A1_c_318_n 0.015224f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.765
cc_84 VPB N_A1_c_310_n 0.00663083f $X=-0.19 $Y=1.66 $X2=0.53 $Y2=1.35
cc_85 VPB N_A1_c_320_n 0.0150935f $X=-0.19 $Y=1.66 $X2=0.53 $Y2=0.74
cc_86 VPB N_A1_c_321_n 0.0155087f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=0.74
cc_87 VPB N_A1_c_322_n 0.0188209f $X=-0.19 $Y=1.66 $X2=1.395 $Y2=2.4
cc_88 VPB N_A1_c_315_n 0.00613987f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.58
cc_89 VPB A1 0.0125553f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB N_A1_c_317_n 0.0500286f $X=-0.19 $Y=1.66 $X2=1.82 $Y2=1.557
cc_91 VPB N_B1_c_400_n 0.0183434f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.765
cc_92 VPB N_B1_c_401_n 0.0145654f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=1.765
cc_93 VPB N_B1_c_402_n 0.0145655f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=1.35
cc_94 VPB N_B1_c_403_n 0.0147736f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_95 VPB N_B1_c_398_n 0.0264266f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.557
cc_96 VPB N_C1_c_479_n 0.0147569f $X=-0.19 $Y=1.66 $X2=0.53 $Y2=1.35
cc_97 VPB N_C1_c_480_n 0.0141056f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=2.4
cc_98 VPB N_C1_c_481_n 0.0141056f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=0.74
cc_99 VPB N_C1_c_475_n 0.0190645f $X=-0.19 $Y=1.66 $X2=1.39 $Y2=0.74
cc_100 VPB N_C1_c_476_n 0.00117364f $X=-0.19 $Y=1.66 $X2=1.395 $Y2=1.765
cc_101 VPB N_C1_c_484_n 0.0272314f $X=-0.19 $Y=1.66 $X2=1.395 $Y2=2.4
cc_102 VPB N_VPWR_c_551_n 0.0103331f $X=-0.19 $Y=1.66 $X2=1.82 $Y2=1.35
cc_103 VPB N_VPWR_c_552_n 0.0599112f $X=-0.19 $Y=1.66 $X2=1.82 $Y2=0.74
cc_104 VPB N_VPWR_c_553_n 0.00271781f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_105 VPB N_VPWR_c_554_n 0.00261791f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_VPWR_c_555_n 0.00261791f $X=-0.19 $Y=1.66 $X2=0.69 $Y2=1.515
cc_107 VPB N_VPWR_c_556_n 0.00261791f $X=-0.19 $Y=1.66 $X2=1.39 $Y2=1.557
cc_108 VPB N_VPWR_c_557_n 0.00434496f $X=-0.19 $Y=1.66 $X2=1.71 $Y2=1.515
cc_109 VPB N_VPWR_c_558_n 0.0185253f $X=-0.19 $Y=1.66 $X2=1.845 $Y2=1.557
cc_110 VPB N_VPWR_c_559_n 0.012368f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_VPWR_c_560_n 0.0164465f $X=-0.19 $Y=1.66 $X2=1.68 $Y2=1.565
cc_112 VPB N_VPWR_c_561_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_VPWR_c_562_n 0.0164465f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_VPWR_c_563_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_VPWR_c_564_n 0.0164465f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_VPWR_c_565_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_566_n 0.0164465f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_567_n 0.00460249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_568_n 0.0185253f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_569_n 0.0991101f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_550_n 0.113565f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_571_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_572_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_A_114_368#_c_692_n 0.00216998f $X=-0.19 $Y=1.66 $X2=1.845 $Y2=2.4
cc_125 VPB N_A_114_368#_c_693_n 0.00180921f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 VPB N_A_114_368#_c_694_n 0.00180921f $X=-0.19 $Y=1.66 $X2=0.69 $Y2=1.515
cc_127 VPB N_A_114_368#_c_695_n 0.00180921f $X=-0.19 $Y=1.66 $X2=1.71 $Y2=1.515
cc_128 VPB N_A_114_368#_c_696_n 0.00180921f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.565
cc_129 VPB N_A_114_368#_c_697_n 0.00216998f $X=-0.19 $Y=1.66 $X2=1.71 $Y2=1.565
cc_130 VPB N_A_114_368#_c_698_n 0.0107168f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_A_114_368#_c_699_n 0.00230503f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_A_114_368#_c_700_n 0.0015494f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_A_114_368#_c_701_n 0.00226167f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_A_114_368#_c_702_n 0.00297142f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_A_1213_368#_c_811_n 0.00555723f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_A_1213_368#_c_812_n 0.00213603f $X=-0.19 $Y=1.66 $X2=1.395 $Y2=2.4
cc_137 VPB N_A_1213_368#_c_813_n 0.00424137f $X=-0.19 $Y=1.66 $X2=1.395 $Y2=2.4
cc_138 VPB N_A_1213_368#_c_814_n 0.00213603f $X=-0.19 $Y=1.66 $X2=1.845
+ $Y2=1.765
cc_139 VPB N_A_1213_368#_c_815_n 0.00926962f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_140 VPB N_A_1213_368#_c_816_n 0.00213603f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_141 VPB N_A_1213_368#_c_817_n 0.0119677f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=1.557
cc_142 VPB N_A_1213_368#_c_818_n 0.053585f $X=-0.19 $Y=1.66 $X2=1.71 $Y2=1.557
cc_143 VPB N_A_1213_368#_c_819_n 0.0021839f $X=-0.19 $Y=1.66 $X2=1.845 $Y2=1.557
cc_144 VPB N_A_1213_368#_c_820_n 0.0021839f $X=-0.19 $Y=1.66 $X2=0.69 $Y2=1.565
cc_145 VPB N_A_1213_368#_c_821_n 0.0021839f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_146 VPB N_Y_c_904_n 0.00432775f $X=-0.19 $Y=1.66 $X2=1.39 $Y2=1.557
cc_147 VPB N_Y_c_905_n 0.00266714f $X=-0.19 $Y=1.66 $X2=1.395 $Y2=1.557
cc_148 VPB N_Y_c_899_n 0.00115545f $X=-0.19 $Y=1.66 $X2=1.71 $Y2=1.515
cc_149 VPB N_Y_c_907_n 0.00137967f $X=-0.19 $Y=1.66 $X2=1.71 $Y2=1.565
cc_150 N_A3_M1026_g N_A2_M1002_g 0.0195801f $X=1.82 $Y=0.74 $X2=0 $Y2=0
cc_151 N_A3_c_158_n N_A2_c_232_n 0.0264592f $X=1.845 $Y=1.765 $X2=0 $Y2=0
cc_152 N_A3_c_159_n A2 0.0381127f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_153 N_A3_c_154_n A2 0.00337932f $X=1.82 $Y=1.557 $X2=0 $Y2=0
cc_154 N_A3_c_159_n N_A2_c_231_n 3.62763e-19 $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_155 N_A3_c_154_n N_A2_c_231_n 0.0205436f $X=1.82 $Y=1.557 $X2=0 $Y2=0
cc_156 N_A3_c_155_n N_VPWR_c_552_n 0.0110944f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_157 N_A3_c_155_n N_VPWR_c_553_n 5.55114e-19 $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_158 N_A3_c_156_n N_VPWR_c_553_n 0.0111578f $X=0.945 $Y=1.765 $X2=0 $Y2=0
cc_159 N_A3_c_157_n N_VPWR_c_553_n 0.0110266f $X=1.395 $Y=1.765 $X2=0 $Y2=0
cc_160 N_A3_c_158_n N_VPWR_c_553_n 5.35985e-19 $X=1.845 $Y=1.765 $X2=0 $Y2=0
cc_161 N_A3_c_157_n N_VPWR_c_554_n 5.35985e-19 $X=1.395 $Y=1.765 $X2=0 $Y2=0
cc_162 N_A3_c_158_n N_VPWR_c_554_n 0.0109874f $X=1.845 $Y=1.765 $X2=0 $Y2=0
cc_163 N_A3_c_157_n N_VPWR_c_560_n 0.00413917f $X=1.395 $Y=1.765 $X2=0 $Y2=0
cc_164 N_A3_c_158_n N_VPWR_c_560_n 0.00413917f $X=1.845 $Y=1.765 $X2=0 $Y2=0
cc_165 N_A3_c_155_n N_VPWR_c_568_n 0.00445602f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_166 N_A3_c_156_n N_VPWR_c_568_n 0.00413917f $X=0.945 $Y=1.765 $X2=0 $Y2=0
cc_167 N_A3_c_155_n N_VPWR_c_550_n 0.0086105f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_168 N_A3_c_156_n N_VPWR_c_550_n 0.00817726f $X=0.945 $Y=1.765 $X2=0 $Y2=0
cc_169 N_A3_c_157_n N_VPWR_c_550_n 0.00817726f $X=1.395 $Y=1.765 $X2=0 $Y2=0
cc_170 N_A3_c_158_n N_VPWR_c_550_n 0.00817726f $X=1.845 $Y=1.765 $X2=0 $Y2=0
cc_171 N_A3_c_155_n N_A_114_368#_c_703_n 0.00203651f $X=0.495 $Y=1.765 $X2=0
+ $Y2=0
cc_172 N_A3_c_159_n N_A_114_368#_c_703_n 0.0193936f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_173 N_A3_c_154_n N_A_114_368#_c_703_n 0.00124229f $X=1.82 $Y=1.557 $X2=0
+ $Y2=0
cc_174 N_A3_c_155_n N_A_114_368#_c_692_n 0.00955225f $X=0.495 $Y=1.765 $X2=0
+ $Y2=0
cc_175 N_A3_c_156_n N_A_114_368#_c_692_n 0.00605728f $X=0.945 $Y=1.765 $X2=0
+ $Y2=0
cc_176 N_A3_c_156_n N_A_114_368#_c_708_n 0.0126853f $X=0.945 $Y=1.765 $X2=0
+ $Y2=0
cc_177 N_A3_c_157_n N_A_114_368#_c_708_n 0.0126853f $X=1.395 $Y=1.765 $X2=0
+ $Y2=0
cc_178 N_A3_c_159_n N_A_114_368#_c_708_n 0.0477183f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_179 N_A3_c_154_n N_A_114_368#_c_708_n 0.00169151f $X=1.82 $Y=1.557 $X2=0
+ $Y2=0
cc_180 N_A3_c_157_n N_A_114_368#_c_693_n 0.00554978f $X=1.395 $Y=1.765 $X2=0
+ $Y2=0
cc_181 N_A3_c_158_n N_A_114_368#_c_693_n 0.00554978f $X=1.845 $Y=1.765 $X2=0
+ $Y2=0
cc_182 N_A3_c_158_n N_A_114_368#_c_714_n 0.0139644f $X=1.845 $Y=1.765 $X2=0
+ $Y2=0
cc_183 N_A3_c_159_n N_A_114_368#_c_714_n 0.0106982f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_184 N_A3_c_159_n N_A_114_368#_c_716_n 0.0150275f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_185 N_A3_c_154_n N_A_114_368#_c_716_n 0.00104296f $X=1.82 $Y=1.557 $X2=0
+ $Y2=0
cc_186 N_A3_M1003_g N_A_34_74#_c_995_n 0.00159319f $X=0.53 $Y=0.74 $X2=0 $Y2=0
cc_187 N_A3_M1003_g N_A_34_74#_c_996_n 0.0157914f $X=0.53 $Y=0.74 $X2=0 $Y2=0
cc_188 N_A3_M1018_g N_A_34_74#_c_996_n 0.01115f $X=0.96 $Y=0.74 $X2=0 $Y2=0
cc_189 N_A3_c_159_n N_A_34_74#_c_996_n 0.0364045f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_190 N_A3_c_154_n N_A_34_74#_c_996_n 0.00427455f $X=1.82 $Y=1.557 $X2=0 $Y2=0
cc_191 N_A3_M1003_g N_A_34_74#_c_998_n 6.58468e-19 $X=0.53 $Y=0.74 $X2=0 $Y2=0
cc_192 N_A3_M1018_g N_A_34_74#_c_998_n 0.00918302f $X=0.96 $Y=0.74 $X2=0 $Y2=0
cc_193 N_A3_M1023_g N_A_34_74#_c_998_n 3.97481e-19 $X=1.39 $Y=0.74 $X2=0 $Y2=0
cc_194 N_A3_M1023_g N_A_34_74#_c_999_n 0.0130918f $X=1.39 $Y=0.74 $X2=0 $Y2=0
cc_195 N_A3_M1026_g N_A_34_74#_c_999_n 0.0136838f $X=1.82 $Y=0.74 $X2=0 $Y2=0
cc_196 N_A3_c_159_n N_A_34_74#_c_999_n 0.0460928f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_197 N_A3_c_154_n N_A_34_74#_c_999_n 0.00385949f $X=1.82 $Y=1.557 $X2=0 $Y2=0
cc_198 N_A3_M1026_g N_A_34_74#_c_1000_n 3.92313e-19 $X=1.82 $Y=0.74 $X2=0 $Y2=0
cc_199 N_A3_M1018_g N_A_34_74#_c_1002_n 0.00157732f $X=0.96 $Y=0.74 $X2=0 $Y2=0
cc_200 N_A3_c_159_n N_A_34_74#_c_1002_n 0.0213626f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_201 N_A3_c_154_n N_A_34_74#_c_1002_n 0.00232957f $X=1.82 $Y=1.557 $X2=0 $Y2=0
cc_202 N_A3_M1003_g N_VGND_c_1069_n 0.0128874f $X=0.53 $Y=0.74 $X2=0 $Y2=0
cc_203 N_A3_M1018_g N_VGND_c_1069_n 0.00204878f $X=0.96 $Y=0.74 $X2=0 $Y2=0
cc_204 N_A3_M1018_g N_VGND_c_1070_n 5.19194e-19 $X=0.96 $Y=0.74 $X2=0 $Y2=0
cc_205 N_A3_M1023_g N_VGND_c_1070_n 0.0108127f $X=1.39 $Y=0.74 $X2=0 $Y2=0
cc_206 N_A3_M1026_g N_VGND_c_1070_n 0.0107959f $X=1.82 $Y=0.74 $X2=0 $Y2=0
cc_207 N_A3_M1003_g N_VGND_c_1072_n 0.00383152f $X=0.53 $Y=0.74 $X2=0 $Y2=0
cc_208 N_A3_M1018_g N_VGND_c_1073_n 0.00434272f $X=0.96 $Y=0.74 $X2=0 $Y2=0
cc_209 N_A3_M1023_g N_VGND_c_1073_n 0.00383152f $X=1.39 $Y=0.74 $X2=0 $Y2=0
cc_210 N_A3_M1003_g N_VGND_c_1076_n 0.00761312f $X=0.53 $Y=0.74 $X2=0 $Y2=0
cc_211 N_A3_M1018_g N_VGND_c_1076_n 0.00820284f $X=0.96 $Y=0.74 $X2=0 $Y2=0
cc_212 N_A3_M1023_g N_VGND_c_1076_n 0.0075754f $X=1.39 $Y=0.74 $X2=0 $Y2=0
cc_213 N_A3_M1026_g N_VGND_c_1076_n 0.00757637f $X=1.82 $Y=0.74 $X2=0 $Y2=0
cc_214 N_A3_M1026_g N_VGND_c_1079_n 0.00383152f $X=1.82 $Y=0.74 $X2=0 $Y2=0
cc_215 N_A2_c_235_n N_A1_c_318_n 0.0259428f $X=3.645 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_216 A2 N_A1_c_315_n 0.00158372f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_217 N_A2_c_231_n N_A1_c_315_n 0.0128527f $X=3.54 $Y=1.557 $X2=0 $Y2=0
cc_218 N_A2_c_232_n N_VPWR_c_554_n 0.0109874f $X=2.295 $Y=1.765 $X2=0 $Y2=0
cc_219 N_A2_c_233_n N_VPWR_c_554_n 5.35985e-19 $X=2.745 $Y=1.765 $X2=0 $Y2=0
cc_220 N_A2_c_232_n N_VPWR_c_555_n 5.35985e-19 $X=2.295 $Y=1.765 $X2=0 $Y2=0
cc_221 N_A2_c_233_n N_VPWR_c_555_n 0.0110266f $X=2.745 $Y=1.765 $X2=0 $Y2=0
cc_222 N_A2_c_234_n N_VPWR_c_555_n 0.0110266f $X=3.195 $Y=1.765 $X2=0 $Y2=0
cc_223 N_A2_c_235_n N_VPWR_c_555_n 5.35985e-19 $X=3.645 $Y=1.765 $X2=0 $Y2=0
cc_224 N_A2_c_234_n N_VPWR_c_556_n 5.35985e-19 $X=3.195 $Y=1.765 $X2=0 $Y2=0
cc_225 N_A2_c_235_n N_VPWR_c_556_n 0.0109294f $X=3.645 $Y=1.765 $X2=0 $Y2=0
cc_226 N_A2_c_232_n N_VPWR_c_562_n 0.00413917f $X=2.295 $Y=1.765 $X2=0 $Y2=0
cc_227 N_A2_c_233_n N_VPWR_c_562_n 0.00413917f $X=2.745 $Y=1.765 $X2=0 $Y2=0
cc_228 N_A2_c_234_n N_VPWR_c_564_n 0.00413917f $X=3.195 $Y=1.765 $X2=0 $Y2=0
cc_229 N_A2_c_235_n N_VPWR_c_564_n 0.00413917f $X=3.645 $Y=1.765 $X2=0 $Y2=0
cc_230 N_A2_c_232_n N_VPWR_c_550_n 0.00817726f $X=2.295 $Y=1.765 $X2=0 $Y2=0
cc_231 N_A2_c_233_n N_VPWR_c_550_n 0.00817726f $X=2.745 $Y=1.765 $X2=0 $Y2=0
cc_232 N_A2_c_234_n N_VPWR_c_550_n 0.00817726f $X=3.195 $Y=1.765 $X2=0 $Y2=0
cc_233 N_A2_c_235_n N_VPWR_c_550_n 0.00817726f $X=3.645 $Y=1.765 $X2=0 $Y2=0
cc_234 N_A2_c_232_n N_A_114_368#_c_714_n 0.0126342f $X=2.295 $Y=1.765 $X2=0
+ $Y2=0
cc_235 A2 N_A_114_368#_c_714_n 0.0258505f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_236 N_A2_c_232_n N_A_114_368#_c_694_n 0.00554978f $X=2.295 $Y=1.765 $X2=0
+ $Y2=0
cc_237 N_A2_c_233_n N_A_114_368#_c_694_n 0.00554978f $X=2.745 $Y=1.765 $X2=0
+ $Y2=0
cc_238 N_A2_c_233_n N_A_114_368#_c_722_n 0.0126853f $X=2.745 $Y=1.765 $X2=0
+ $Y2=0
cc_239 N_A2_c_234_n N_A_114_368#_c_722_n 0.0126853f $X=3.195 $Y=1.765 $X2=0
+ $Y2=0
cc_240 A2 N_A_114_368#_c_722_n 0.0477183f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_241 N_A2_c_231_n N_A_114_368#_c_722_n 0.00169504f $X=3.54 $Y=1.557 $X2=0
+ $Y2=0
cc_242 N_A2_c_234_n N_A_114_368#_c_695_n 0.00554978f $X=3.195 $Y=1.765 $X2=0
+ $Y2=0
cc_243 N_A2_c_235_n N_A_114_368#_c_695_n 0.00554978f $X=3.645 $Y=1.765 $X2=0
+ $Y2=0
cc_244 N_A2_c_235_n N_A_114_368#_c_728_n 0.0127781f $X=3.645 $Y=1.765 $X2=0
+ $Y2=0
cc_245 A2 N_A_114_368#_c_728_n 0.0136167f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_246 A2 N_A_114_368#_c_730_n 0.0150275f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_247 N_A2_c_231_n N_A_114_368#_c_730_n 0.00104155f $X=3.54 $Y=1.557 $X2=0
+ $Y2=0
cc_248 A2 N_A_114_368#_c_732_n 0.0150275f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_249 N_A2_c_231_n N_A_114_368#_c_732_n 0.00103872f $X=3.54 $Y=1.557 $X2=0
+ $Y2=0
cc_250 N_A2_M1002_g N_A_34_74#_c_1000_n 4.08775e-19 $X=2.25 $Y=0.74 $X2=0 $Y2=0
cc_251 N_A2_M1033_g N_A_34_74#_c_1001_n 0.00914581f $X=3.11 $Y=0.74 $X2=0 $Y2=0
cc_252 N_A2_M1034_g N_A_34_74#_c_1001_n 0.00983999f $X=3.54 $Y=0.74 $X2=0 $Y2=0
cc_253 N_A2_c_231_n N_A_34_74#_c_1001_n 0.00226259f $X=3.54 $Y=1.557 $X2=0 $Y2=0
cc_254 A2 N_A_34_74#_c_1003_n 0.00676262f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_255 N_A2_M1002_g N_A_34_74#_c_1004_n 0.0142123f $X=2.25 $Y=0.74 $X2=0 $Y2=0
cc_256 N_A2_M1011_g N_A_34_74#_c_1004_n 0.00913639f $X=2.68 $Y=0.74 $X2=0 $Y2=0
cc_257 A2 N_A_34_74#_c_1004_n 0.11368f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_258 N_A2_c_231_n N_A_34_74#_c_1004_n 0.00225173f $X=3.54 $Y=1.557 $X2=0 $Y2=0
cc_259 N_A2_M1002_g N_A_34_74#_c_1005_n 6.21182e-19 $X=2.25 $Y=0.74 $X2=0 $Y2=0
cc_260 N_A2_M1011_g N_A_34_74#_c_1005_n 0.0058f $X=2.68 $Y=0.74 $X2=0 $Y2=0
cc_261 N_A2_M1033_g N_A_34_74#_c_1005_n 0.00554487f $X=3.11 $Y=0.74 $X2=0 $Y2=0
cc_262 N_A2_M1034_g N_A_34_74#_c_1005_n 6.0146e-19 $X=3.54 $Y=0.74 $X2=0 $Y2=0
cc_263 N_A2_c_231_n N_A_34_74#_c_1005_n 0.00229127f $X=3.54 $Y=1.557 $X2=0 $Y2=0
cc_264 N_A2_M1033_g N_A_34_74#_c_1006_n 7.02574e-19 $X=3.11 $Y=0.74 $X2=0 $Y2=0
cc_265 N_A2_M1034_g N_A_34_74#_c_1006_n 0.00667962f $X=3.54 $Y=0.74 $X2=0 $Y2=0
cc_266 A2 N_A_34_74#_c_1006_n 0.0101258f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_267 N_A2_c_231_n N_A_34_74#_c_1006_n 0.00355377f $X=3.54 $Y=1.557 $X2=0 $Y2=0
cc_268 N_A2_M1002_g N_VGND_c_1070_n 6.96792e-19 $X=2.25 $Y=0.74 $X2=0 $Y2=0
cc_269 N_A2_M1002_g N_VGND_c_1076_n 0.00817716f $X=2.25 $Y=0.74 $X2=0 $Y2=0
cc_270 N_A2_M1011_g N_VGND_c_1076_n 0.00359121f $X=2.68 $Y=0.74 $X2=0 $Y2=0
cc_271 N_A2_M1033_g N_VGND_c_1076_n 0.00359121f $X=3.11 $Y=0.74 $X2=0 $Y2=0
cc_272 N_A2_M1034_g N_VGND_c_1076_n 0.0036412f $X=3.54 $Y=0.74 $X2=0 $Y2=0
cc_273 N_A2_M1002_g N_VGND_c_1079_n 0.00433162f $X=2.25 $Y=0.74 $X2=0 $Y2=0
cc_274 N_A2_M1011_g N_VGND_c_1079_n 0.00291649f $X=2.68 $Y=0.74 $X2=0 $Y2=0
cc_275 N_A2_M1033_g N_VGND_c_1079_n 0.00291649f $X=3.11 $Y=0.74 $X2=0 $Y2=0
cc_276 N_A2_M1034_g N_VGND_c_1079_n 0.00291649f $X=3.54 $Y=0.74 $X2=0 $Y2=0
cc_277 N_A2_M1002_g N_A_465_74#_c_1158_n 0.00432482f $X=2.25 $Y=0.74 $X2=0 $Y2=0
cc_278 N_A2_M1011_g N_A_465_74#_c_1159_n 0.0111551f $X=2.68 $Y=0.74 $X2=0 $Y2=0
cc_279 N_A2_M1033_g N_A_465_74#_c_1159_n 0.0111551f $X=3.11 $Y=0.74 $X2=0 $Y2=0
cc_280 N_A2_M1034_g N_A_465_74#_c_1162_n 0.0141524f $X=3.54 $Y=0.74 $X2=0 $Y2=0
cc_281 A1 N_B1_c_400_n 5.26509e-19 $X=5.915 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_282 N_A1_M1035_g N_B1_M1010_g 0.0184495f $X=6 $Y=0.74 $X2=0 $Y2=0
cc_283 N_A1_M1035_g N_B1_c_398_n 0.0193595f $X=6 $Y=0.74 $X2=0 $Y2=0
cc_284 A1 N_B1_c_398_n 0.00812377f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_285 A1 N_B1_c_399_n 0.0093478f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_286 N_A1_c_318_n N_VPWR_c_556_n 0.0109874f $X=4.095 $Y=1.765 $X2=0 $Y2=0
cc_287 N_A1_c_320_n N_VPWR_c_556_n 5.35985e-19 $X=4.545 $Y=1.765 $X2=0 $Y2=0
cc_288 N_A1_c_318_n N_VPWR_c_557_n 5.37805e-19 $X=4.095 $Y=1.765 $X2=0 $Y2=0
cc_289 N_A1_c_320_n N_VPWR_c_557_n 0.0106464f $X=4.545 $Y=1.765 $X2=0 $Y2=0
cc_290 N_A1_c_321_n N_VPWR_c_557_n 0.00395359f $X=4.995 $Y=1.765 $X2=0 $Y2=0
cc_291 N_A1_c_321_n N_VPWR_c_558_n 0.00445602f $X=4.995 $Y=1.765 $X2=0 $Y2=0
cc_292 N_A1_c_322_n N_VPWR_c_558_n 0.00413917f $X=5.445 $Y=1.765 $X2=0 $Y2=0
cc_293 N_A1_c_321_n N_VPWR_c_559_n 5.55114e-19 $X=4.995 $Y=1.765 $X2=0 $Y2=0
cc_294 N_A1_c_322_n N_VPWR_c_559_n 0.0121487f $X=5.445 $Y=1.765 $X2=0 $Y2=0
cc_295 N_A1_c_318_n N_VPWR_c_566_n 0.00413917f $X=4.095 $Y=1.765 $X2=0 $Y2=0
cc_296 N_A1_c_320_n N_VPWR_c_566_n 0.00413917f $X=4.545 $Y=1.765 $X2=0 $Y2=0
cc_297 N_A1_c_318_n N_VPWR_c_550_n 0.00817726f $X=4.095 $Y=1.765 $X2=0 $Y2=0
cc_298 N_A1_c_320_n N_VPWR_c_550_n 0.00817726f $X=4.545 $Y=1.765 $X2=0 $Y2=0
cc_299 N_A1_c_321_n N_VPWR_c_550_n 0.00857589f $X=4.995 $Y=1.765 $X2=0 $Y2=0
cc_300 N_A1_c_322_n N_VPWR_c_550_n 0.00817726f $X=5.445 $Y=1.765 $X2=0 $Y2=0
cc_301 N_A1_c_318_n N_A_114_368#_c_728_n 0.0167245f $X=4.095 $Y=1.765 $X2=0
+ $Y2=0
cc_302 N_A1_c_310_n N_A_114_368#_c_728_n 8.52892e-19 $X=4.455 $Y=1.605 $X2=0
+ $Y2=0
cc_303 N_A1_c_318_n N_A_114_368#_c_696_n 0.00576879f $X=4.095 $Y=1.765 $X2=0
+ $Y2=0
cc_304 N_A1_c_320_n N_A_114_368#_c_696_n 0.0039133f $X=4.545 $Y=1.765 $X2=0
+ $Y2=0
cc_305 N_A1_c_310_n N_A_114_368#_c_738_n 8.52892e-19 $X=4.455 $Y=1.605 $X2=0
+ $Y2=0
cc_306 N_A1_c_320_n N_A_114_368#_c_738_n 0.0167755f $X=4.545 $Y=1.765 $X2=0
+ $Y2=0
cc_307 N_A1_c_321_n N_A_114_368#_c_738_n 0.0120074f $X=4.995 $Y=1.765 $X2=0
+ $Y2=0
cc_308 A1 N_A_114_368#_c_738_n 0.0289213f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_309 N_A1_c_317_n N_A_114_368#_c_738_n 0.00130366f $X=5.91 $Y=1.515 $X2=0
+ $Y2=0
cc_310 N_A1_c_320_n N_A_114_368#_c_697_n 6.71799e-19 $X=4.545 $Y=1.765 $X2=0
+ $Y2=0
cc_311 N_A1_c_321_n N_A_114_368#_c_697_n 0.0104892f $X=4.995 $Y=1.765 $X2=0
+ $Y2=0
cc_312 N_A1_c_322_n N_A_114_368#_c_697_n 0.00605728f $X=5.445 $Y=1.765 $X2=0
+ $Y2=0
cc_313 N_A1_c_322_n N_A_114_368#_c_698_n 0.0146058f $X=5.445 $Y=1.765 $X2=0
+ $Y2=0
cc_314 A1 N_A_114_368#_c_698_n 0.059662f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_315 N_A1_c_317_n N_A_114_368#_c_698_n 0.00303269f $X=5.91 $Y=1.515 $X2=0
+ $Y2=0
cc_316 N_A1_c_318_n N_A_114_368#_c_701_n 0.00262483f $X=4.095 $Y=1.765 $X2=0
+ $Y2=0
cc_317 N_A1_c_310_n N_A_114_368#_c_701_n 0.00721924f $X=4.455 $Y=1.605 $X2=0
+ $Y2=0
cc_318 N_A1_c_320_n N_A_114_368#_c_701_n 0.00262483f $X=4.545 $Y=1.765 $X2=0
+ $Y2=0
cc_319 N_A1_c_321_n N_A_114_368#_c_752_n 4.27055e-19 $X=4.995 $Y=1.765 $X2=0
+ $Y2=0
cc_320 A1 N_A_114_368#_c_752_n 0.0193936f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_321 N_A1_c_317_n N_A_114_368#_c_752_n 0.00123522f $X=5.91 $Y=1.515 $X2=0
+ $Y2=0
cc_322 N_A1_c_322_n N_A_1213_368#_c_813_n 5.75404e-19 $X=5.445 $Y=1.765 $X2=0
+ $Y2=0
cc_323 N_A1_M1007_g N_Y_c_896_n 0.0106768f $X=4.71 $Y=0.74 $X2=0 $Y2=0
cc_324 N_A1_M1012_g N_Y_c_896_n 0.0123927f $X=5.14 $Y=0.74 $X2=0 $Y2=0
cc_325 N_A1_M1021_g N_Y_c_896_n 0.0123136f $X=5.57 $Y=0.74 $X2=0 $Y2=0
cc_326 N_A1_M1035_g N_Y_c_896_n 0.0132419f $X=6 $Y=0.74 $X2=0 $Y2=0
cc_327 N_A1_c_317_n N_Y_c_896_n 0.00696502f $X=5.91 $Y=1.515 $X2=0 $Y2=0
cc_328 N_A1_M1035_g N_Y_c_897_n 4.15473e-19 $X=6 $Y=0.74 $X2=0 $Y2=0
cc_329 N_A1_c_310_n N_Y_c_900_n 0.00985076f $X=4.455 $Y=1.605 $X2=0 $Y2=0
cc_330 N_A1_M1007_g N_Y_c_900_n 0.00318903f $X=4.71 $Y=0.74 $X2=0 $Y2=0
cc_331 N_A1_M1012_g N_Y_c_900_n 3.85913e-19 $X=5.14 $Y=0.74 $X2=0 $Y2=0
cc_332 A1 N_Y_c_900_n 0.0949302f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_333 N_A1_M1007_g N_VGND_c_1076_n 0.0036412f $X=4.71 $Y=0.74 $X2=0 $Y2=0
cc_334 N_A1_M1012_g N_VGND_c_1076_n 0.00359121f $X=5.14 $Y=0.74 $X2=0 $Y2=0
cc_335 N_A1_M1021_g N_VGND_c_1076_n 0.00359121f $X=5.57 $Y=0.74 $X2=0 $Y2=0
cc_336 N_A1_M1035_g N_VGND_c_1076_n 0.00449183f $X=6 $Y=0.74 $X2=0 $Y2=0
cc_337 N_A1_M1007_g N_VGND_c_1079_n 0.00291649f $X=4.71 $Y=0.74 $X2=0 $Y2=0
cc_338 N_A1_M1012_g N_VGND_c_1079_n 0.00291649f $X=5.14 $Y=0.74 $X2=0 $Y2=0
cc_339 N_A1_M1021_g N_VGND_c_1079_n 0.00291649f $X=5.57 $Y=0.74 $X2=0 $Y2=0
cc_340 N_A1_M1035_g N_VGND_c_1079_n 0.00433162f $X=6 $Y=0.74 $X2=0 $Y2=0
cc_341 N_A1_M1012_g N_A_465_74#_c_1161_n 3.85913e-19 $X=5.14 $Y=0.74 $X2=0 $Y2=0
cc_342 N_A1_M1021_g N_A_465_74#_c_1161_n 0.00281528f $X=5.57 $Y=0.74 $X2=0 $Y2=0
cc_343 N_A1_M1035_g N_A_465_74#_c_1161_n 0.00420713f $X=6 $Y=0.74 $X2=0 $Y2=0
cc_344 N_A1_M1007_g N_A_465_74#_c_1162_n 0.0136253f $X=4.71 $Y=0.74 $X2=0 $Y2=0
cc_345 N_A1_M1012_g N_A_465_74#_c_1162_n 0.0106927f $X=5.14 $Y=0.74 $X2=0 $Y2=0
cc_346 N_A1_M1021_g N_A_465_74#_c_1162_n 0.00920696f $X=5.57 $Y=0.74 $X2=0 $Y2=0
cc_347 N_B1_M1019_g N_C1_c_472_n 0.0122583f $X=7.71 $Y=0.74 $X2=-0.19 $Y2=-0.245
cc_348 N_B1_c_403_n N_C1_c_479_n 0.0106731f $X=7.765 $Y=1.765 $X2=0 $Y2=0
cc_349 B1 N_C1_c_475_n 8.33085e-19 $X=7.355 $Y=1.21 $X2=0 $Y2=0
cc_350 N_B1_c_398_n N_C1_c_475_n 0.0270603f $X=7.71 $Y=1.542 $X2=0 $Y2=0
cc_351 N_B1_M1019_g N_C1_c_478_n 3.74992e-19 $X=7.71 $Y=0.74 $X2=0 $Y2=0
cc_352 B1 N_C1_c_478_n 0.0168871f $X=7.355 $Y=1.21 $X2=0 $Y2=0
cc_353 N_B1_c_398_n N_C1_c_478_n 4.37969e-19 $X=7.71 $Y=1.542 $X2=0 $Y2=0
cc_354 N_B1_c_400_n N_VPWR_c_559_n 0.00180354f $X=6.415 $Y=1.765 $X2=0 $Y2=0
cc_355 N_B1_c_400_n N_VPWR_c_569_n 0.00278257f $X=6.415 $Y=1.765 $X2=0 $Y2=0
cc_356 N_B1_c_401_n N_VPWR_c_569_n 0.00278257f $X=6.865 $Y=1.765 $X2=0 $Y2=0
cc_357 N_B1_c_402_n N_VPWR_c_569_n 0.00278257f $X=7.315 $Y=1.765 $X2=0 $Y2=0
cc_358 N_B1_c_403_n N_VPWR_c_569_n 0.00278257f $X=7.765 $Y=1.765 $X2=0 $Y2=0
cc_359 N_B1_c_400_n N_VPWR_c_550_n 0.00358623f $X=6.415 $Y=1.765 $X2=0 $Y2=0
cc_360 N_B1_c_401_n N_VPWR_c_550_n 0.00353822f $X=6.865 $Y=1.765 $X2=0 $Y2=0
cc_361 N_B1_c_402_n N_VPWR_c_550_n 0.00353822f $X=7.315 $Y=1.765 $X2=0 $Y2=0
cc_362 N_B1_c_403_n N_VPWR_c_550_n 0.00353905f $X=7.765 $Y=1.765 $X2=0 $Y2=0
cc_363 N_B1_c_400_n N_A_114_368#_c_698_n 0.0175856f $X=6.415 $Y=1.765 $X2=0
+ $Y2=0
cc_364 N_B1_c_401_n N_A_114_368#_c_699_n 0.0176407f $X=6.865 $Y=1.765 $X2=0
+ $Y2=0
cc_365 N_B1_c_402_n N_A_114_368#_c_699_n 0.0176946f $X=7.315 $Y=1.765 $X2=0
+ $Y2=0
cc_366 B1 N_A_114_368#_c_699_n 0.00824106f $X=7.355 $Y=1.21 $X2=0 $Y2=0
cc_367 N_B1_c_398_n N_A_114_368#_c_699_n 0.00875199f $X=7.71 $Y=1.542 $X2=0
+ $Y2=0
cc_368 N_B1_c_399_n N_A_114_368#_c_699_n 0.0432857f $X=7.32 $Y=1.415 $X2=0 $Y2=0
cc_369 B1 N_A_114_368#_c_700_n 0.0197638f $X=7.355 $Y=1.21 $X2=0 $Y2=0
cc_370 N_B1_c_398_n N_A_114_368#_c_700_n 0.00181f $X=7.71 $Y=1.542 $X2=0 $Y2=0
cc_371 N_B1_c_400_n N_A_114_368#_c_702_n 0.00925563f $X=6.415 $Y=1.765 $X2=0
+ $Y2=0
cc_372 N_B1_c_398_n N_A_114_368#_c_702_n 0.0121421f $X=7.71 $Y=1.542 $X2=0 $Y2=0
cc_373 N_B1_c_400_n N_A_1213_368#_c_811_n 0.00749701f $X=6.415 $Y=1.765 $X2=0
+ $Y2=0
cc_374 N_B1_c_401_n N_A_1213_368#_c_811_n 5.44258e-19 $X=6.865 $Y=1.765 $X2=0
+ $Y2=0
cc_375 N_B1_c_400_n N_A_1213_368#_c_812_n 0.0108414f $X=6.415 $Y=1.765 $X2=0
+ $Y2=0
cc_376 N_B1_c_401_n N_A_1213_368#_c_812_n 0.0108414f $X=6.865 $Y=1.765 $X2=0
+ $Y2=0
cc_377 N_B1_c_400_n N_A_1213_368#_c_813_n 0.00262934f $X=6.415 $Y=1.765 $X2=0
+ $Y2=0
cc_378 N_B1_c_400_n N_A_1213_368#_c_828_n 5.44258e-19 $X=6.415 $Y=1.765 $X2=0
+ $Y2=0
cc_379 N_B1_c_401_n N_A_1213_368#_c_828_n 0.00732658f $X=6.865 $Y=1.765 $X2=0
+ $Y2=0
cc_380 N_B1_c_402_n N_A_1213_368#_c_828_n 0.00732658f $X=7.315 $Y=1.765 $X2=0
+ $Y2=0
cc_381 N_B1_c_403_n N_A_1213_368#_c_828_n 5.44258e-19 $X=7.765 $Y=1.765 $X2=0
+ $Y2=0
cc_382 N_B1_c_402_n N_A_1213_368#_c_814_n 0.0108414f $X=7.315 $Y=1.765 $X2=0
+ $Y2=0
cc_383 N_B1_c_403_n N_A_1213_368#_c_814_n 0.0108414f $X=7.765 $Y=1.765 $X2=0
+ $Y2=0
cc_384 N_B1_c_402_n N_A_1213_368#_c_815_n 6.82622e-19 $X=7.315 $Y=1.765 $X2=0
+ $Y2=0
cc_385 N_B1_c_403_n N_A_1213_368#_c_815_n 0.0131042f $X=7.765 $Y=1.765 $X2=0
+ $Y2=0
cc_386 N_B1_c_398_n N_A_1213_368#_c_815_n 7.38909e-19 $X=7.71 $Y=1.542 $X2=0
+ $Y2=0
cc_387 N_B1_c_401_n N_A_1213_368#_c_819_n 0.00175197f $X=6.865 $Y=1.765 $X2=0
+ $Y2=0
cc_388 N_B1_c_402_n N_A_1213_368#_c_819_n 0.00175197f $X=7.315 $Y=1.765 $X2=0
+ $Y2=0
cc_389 N_B1_c_403_n N_A_1213_368#_c_820_n 0.00171731f $X=7.765 $Y=1.765 $X2=0
+ $Y2=0
cc_390 N_B1_M1010_g N_Y_c_897_n 0.0114845f $X=6.43 $Y=0.74 $X2=0 $Y2=0
cc_391 N_B1_M1010_g N_Y_c_919_n 0.0143576f $X=6.43 $Y=0.74 $X2=0 $Y2=0
cc_392 N_B1_M1019_g N_Y_c_919_n 0.0112203f $X=7.71 $Y=0.74 $X2=0 $Y2=0
cc_393 B1 N_Y_c_919_n 0.0268604f $X=7.355 $Y=1.21 $X2=0 $Y2=0
cc_394 N_B1_c_398_n N_Y_c_919_n 0.00966104f $X=7.71 $Y=1.542 $X2=0 $Y2=0
cc_395 N_B1_c_399_n N_Y_c_919_n 0.0436852f $X=7.32 $Y=1.415 $X2=0 $Y2=0
cc_396 N_B1_M1019_g N_Y_c_898_n 0.0109447f $X=7.71 $Y=0.74 $X2=0 $Y2=0
cc_397 N_B1_M1010_g N_Y_c_901_n 0.00755467f $X=6.43 $Y=0.74 $X2=0 $Y2=0
cc_398 N_B1_c_398_n N_Y_c_901_n 0.00138366f $X=7.71 $Y=1.542 $X2=0 $Y2=0
cc_399 N_B1_M1019_g N_Y_c_927_n 0.0024979f $X=7.71 $Y=0.74 $X2=0 $Y2=0
cc_400 B1 N_Y_c_927_n 0.00135505f $X=7.355 $Y=1.21 $X2=0 $Y2=0
cc_401 N_B1_c_398_n N_Y_c_927_n 0.00143832f $X=7.71 $Y=1.542 $X2=0 $Y2=0
cc_402 N_B1_M1019_g N_VGND_c_1071_n 4.39708e-19 $X=7.71 $Y=0.74 $X2=0 $Y2=0
cc_403 N_B1_M1019_g N_VGND_c_1074_n 0.00434272f $X=7.71 $Y=0.74 $X2=0 $Y2=0
cc_404 N_B1_M1010_g N_VGND_c_1076_n 0.00449911f $X=6.43 $Y=0.74 $X2=0 $Y2=0
cc_405 N_B1_M1019_g N_VGND_c_1076_n 0.00449911f $X=7.71 $Y=0.74 $X2=0 $Y2=0
cc_406 N_B1_M1010_g N_VGND_c_1079_n 0.00434272f $X=6.43 $Y=0.74 $X2=0 $Y2=0
cc_407 N_B1_M1010_g N_VGND_c_1080_n 0.0113932f $X=6.43 $Y=0.74 $X2=0 $Y2=0
cc_408 N_B1_M1019_g N_VGND_c_1080_n 0.00963538f $X=7.71 $Y=0.74 $X2=0 $Y2=0
cc_409 N_C1_c_479_n N_VPWR_c_569_n 0.00278257f $X=8.215 $Y=1.765 $X2=0 $Y2=0
cc_410 N_C1_c_480_n N_VPWR_c_569_n 0.00278257f $X=8.665 $Y=1.765 $X2=0 $Y2=0
cc_411 N_C1_c_481_n N_VPWR_c_569_n 0.00278257f $X=9.115 $Y=1.765 $X2=0 $Y2=0
cc_412 N_C1_c_484_n N_VPWR_c_569_n 0.00278257f $X=9.565 $Y=1.765 $X2=0 $Y2=0
cc_413 N_C1_c_479_n N_VPWR_c_550_n 0.00353905f $X=8.215 $Y=1.765 $X2=0 $Y2=0
cc_414 N_C1_c_480_n N_VPWR_c_550_n 0.00353822f $X=8.665 $Y=1.765 $X2=0 $Y2=0
cc_415 N_C1_c_481_n N_VPWR_c_550_n 0.00353822f $X=9.115 $Y=1.765 $X2=0 $Y2=0
cc_416 N_C1_c_484_n N_VPWR_c_550_n 0.00357349f $X=9.565 $Y=1.765 $X2=0 $Y2=0
cc_417 N_C1_c_479_n N_A_1213_368#_c_815_n 0.0133547f $X=8.215 $Y=1.765 $X2=0
+ $Y2=0
cc_418 N_C1_c_480_n N_A_1213_368#_c_815_n 7.22826e-19 $X=8.665 $Y=1.765 $X2=0
+ $Y2=0
cc_419 N_C1_c_475_n N_A_1213_368#_c_815_n 9.43675e-19 $X=9.205 $Y=1.345 $X2=0
+ $Y2=0
cc_420 N_C1_c_478_n N_A_1213_368#_c_815_n 0.00526811f $X=8.47 $Y=1.365 $X2=0
+ $Y2=0
cc_421 N_C1_c_479_n N_A_1213_368#_c_816_n 0.0108414f $X=8.215 $Y=1.765 $X2=0
+ $Y2=0
cc_422 N_C1_c_480_n N_A_1213_368#_c_816_n 0.0108414f $X=8.665 $Y=1.765 $X2=0
+ $Y2=0
cc_423 N_C1_c_479_n N_A_1213_368#_c_846_n 6.41034e-19 $X=8.215 $Y=1.765 $X2=0
+ $Y2=0
cc_424 N_C1_c_480_n N_A_1213_368#_c_846_n 0.0125495f $X=8.665 $Y=1.765 $X2=0
+ $Y2=0
cc_425 N_C1_c_481_n N_A_1213_368#_c_846_n 0.0125495f $X=9.115 $Y=1.765 $X2=0
+ $Y2=0
cc_426 N_C1_c_484_n N_A_1213_368#_c_846_n 6.41034e-19 $X=9.565 $Y=1.765 $X2=0
+ $Y2=0
cc_427 N_C1_c_481_n N_A_1213_368#_c_817_n 0.0108414f $X=9.115 $Y=1.765 $X2=0
+ $Y2=0
cc_428 N_C1_c_484_n N_A_1213_368#_c_817_n 0.0134708f $X=9.565 $Y=1.765 $X2=0
+ $Y2=0
cc_429 N_C1_c_481_n N_A_1213_368#_c_818_n 7.22826e-19 $X=9.115 $Y=1.765 $X2=0
+ $Y2=0
cc_430 N_C1_c_484_n N_A_1213_368#_c_818_n 0.0151366f $X=9.565 $Y=1.765 $X2=0
+ $Y2=0
cc_431 N_C1_c_479_n N_A_1213_368#_c_820_n 0.00171731f $X=8.215 $Y=1.765 $X2=0
+ $Y2=0
cc_432 N_C1_c_480_n N_A_1213_368#_c_821_n 0.00175197f $X=8.665 $Y=1.765 $X2=0
+ $Y2=0
cc_433 N_C1_c_481_n N_A_1213_368#_c_821_n 0.00175197f $X=9.115 $Y=1.765 $X2=0
+ $Y2=0
cc_434 N_C1_c_479_n N_Y_c_930_n 0.00351644f $X=8.215 $Y=1.765 $X2=0 $Y2=0
cc_435 N_C1_c_480_n N_Y_c_930_n 0.006269f $X=8.665 $Y=1.765 $X2=0 $Y2=0
cc_436 N_C1_c_480_n N_Y_c_904_n 0.0101246f $X=8.665 $Y=1.765 $X2=0 $Y2=0
cc_437 N_C1_c_481_n N_Y_c_904_n 0.0101246f $X=9.115 $Y=1.765 $X2=0 $Y2=0
cc_438 N_C1_c_475_n N_Y_c_904_n 0.0148625f $X=9.205 $Y=1.345 $X2=0 $Y2=0
cc_439 N_C1_c_477_n N_Y_c_904_n 0.0408056f $X=8.91 $Y=1.385 $X2=0 $Y2=0
cc_440 N_C1_c_479_n N_Y_c_905_n 0.00212373f $X=8.215 $Y=1.765 $X2=0 $Y2=0
cc_441 N_C1_c_475_n N_Y_c_905_n 0.00243064f $X=9.205 $Y=1.345 $X2=0 $Y2=0
cc_442 N_C1_c_477_n N_Y_c_905_n 0.00463739f $X=8.91 $Y=1.385 $X2=0 $Y2=0
cc_443 N_C1_c_478_n N_Y_c_905_n 0.00982302f $X=8.47 $Y=1.365 $X2=0 $Y2=0
cc_444 N_C1_c_473_n N_Y_c_899_n 0.00275313f $X=8.57 $Y=1.22 $X2=0 $Y2=0
cc_445 N_C1_c_474_n N_Y_c_899_n 0.0226183f $X=9.475 $Y=1.345 $X2=0 $Y2=0
cc_446 N_C1_c_475_n N_Y_c_899_n 0.00479365f $X=9.205 $Y=1.345 $X2=0 $Y2=0
cc_447 N_C1_c_476_n N_Y_c_899_n 0.00598622f $X=9.565 $Y=1.675 $X2=0 $Y2=0
cc_448 N_C1_c_477_n N_Y_c_899_n 0.0273925f $X=8.91 $Y=1.385 $X2=0 $Y2=0
cc_449 N_C1_c_481_n N_Y_c_945_n 0.006269f $X=9.115 $Y=1.765 $X2=0 $Y2=0
cc_450 N_C1_c_484_n N_Y_c_945_n 0.00351644f $X=9.565 $Y=1.765 $X2=0 $Y2=0
cc_451 N_C1_c_484_n N_Y_c_907_n 0.00355831f $X=9.565 $Y=1.765 $X2=0 $Y2=0
cc_452 N_C1_c_474_n Y 0.00678239f $X=9.475 $Y=1.345 $X2=0 $Y2=0
cc_453 N_C1_c_472_n N_Y_c_949_n 0.00985057f $X=8.14 $Y=1.22 $X2=0 $Y2=0
cc_454 N_C1_c_473_n N_Y_c_949_n 0.00961729f $X=8.57 $Y=1.22 $X2=0 $Y2=0
cc_455 N_C1_c_475_n N_Y_c_949_n 6.22937e-19 $X=9.205 $Y=1.345 $X2=0 $Y2=0
cc_456 N_C1_c_477_n N_Y_c_949_n 0.046849f $X=8.91 $Y=1.385 $X2=0 $Y2=0
cc_457 N_C1_c_478_n N_Y_c_949_n 0.0251469f $X=8.47 $Y=1.365 $X2=0 $Y2=0
cc_458 N_C1_c_473_n N_Y_c_903_n 8.21094e-19 $X=8.57 $Y=1.22 $X2=0 $Y2=0
cc_459 N_C1_c_474_n N_Y_c_903_n 7.19437e-19 $X=9.475 $Y=1.345 $X2=0 $Y2=0
cc_460 N_C1_c_475_n N_Y_c_903_n 0.0110987f $X=9.205 $Y=1.345 $X2=0 $Y2=0
cc_461 N_C1_c_472_n N_VGND_c_1071_n 0.00769352f $X=8.14 $Y=1.22 $X2=0 $Y2=0
cc_462 N_C1_c_473_n N_VGND_c_1071_n 0.0105522f $X=8.57 $Y=1.22 $X2=0 $Y2=0
cc_463 N_C1_c_472_n N_VGND_c_1074_n 0.00383152f $X=8.14 $Y=1.22 $X2=0 $Y2=0
cc_464 N_C1_c_473_n N_VGND_c_1075_n 0.00383152f $X=8.57 $Y=1.22 $X2=0 $Y2=0
cc_465 N_C1_c_472_n N_VGND_c_1076_n 0.00384065f $X=8.14 $Y=1.22 $X2=0 $Y2=0
cc_466 N_C1_c_473_n N_VGND_c_1076_n 0.00388966f $X=8.57 $Y=1.22 $X2=0 $Y2=0
cc_467 N_VPWR_c_552_n N_A_114_368#_c_703_n 0.0121024f $X=0.27 $Y=1.985 $X2=0
+ $Y2=0
cc_468 N_VPWR_c_552_n N_A_114_368#_c_692_n 0.0564818f $X=0.27 $Y=1.985 $X2=0
+ $Y2=0
cc_469 N_VPWR_c_553_n N_A_114_368#_c_692_n 0.0462948f $X=1.17 $Y=2.455 $X2=0
+ $Y2=0
cc_470 N_VPWR_c_568_n N_A_114_368#_c_692_n 0.0110241f $X=1.005 $Y=3.33 $X2=0
+ $Y2=0
cc_471 N_VPWR_c_550_n N_A_114_368#_c_692_n 0.00909194f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_472 N_VPWR_M1008_s N_A_114_368#_c_708_n 0.00359365f $X=1.02 $Y=1.84 $X2=0
+ $Y2=0
cc_473 N_VPWR_c_553_n N_A_114_368#_c_708_n 0.0171813f $X=1.17 $Y=2.455 $X2=0
+ $Y2=0
cc_474 N_VPWR_c_553_n N_A_114_368#_c_693_n 0.0449718f $X=1.17 $Y=2.455 $X2=0
+ $Y2=0
cc_475 N_VPWR_c_554_n N_A_114_368#_c_693_n 0.0449718f $X=2.07 $Y=2.455 $X2=0
+ $Y2=0
cc_476 N_VPWR_c_560_n N_A_114_368#_c_693_n 0.00749631f $X=1.905 $Y=3.33 $X2=0
+ $Y2=0
cc_477 N_VPWR_c_550_n N_A_114_368#_c_693_n 0.0062048f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_478 N_VPWR_M1029_s N_A_114_368#_c_714_n 0.00582921f $X=1.92 $Y=1.84 $X2=0
+ $Y2=0
cc_479 N_VPWR_c_554_n N_A_114_368#_c_714_n 0.0171814f $X=2.07 $Y=2.455 $X2=0
+ $Y2=0
cc_480 N_VPWR_c_554_n N_A_114_368#_c_694_n 0.0449718f $X=2.07 $Y=2.455 $X2=0
+ $Y2=0
cc_481 N_VPWR_c_555_n N_A_114_368#_c_694_n 0.0449718f $X=2.97 $Y=2.455 $X2=0
+ $Y2=0
cc_482 N_VPWR_c_562_n N_A_114_368#_c_694_n 0.00749631f $X=2.805 $Y=3.33 $X2=0
+ $Y2=0
cc_483 N_VPWR_c_550_n N_A_114_368#_c_694_n 0.0062048f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_484 N_VPWR_M1016_d N_A_114_368#_c_722_n 0.00359365f $X=2.82 $Y=1.84 $X2=0
+ $Y2=0
cc_485 N_VPWR_c_555_n N_A_114_368#_c_722_n 0.0171813f $X=2.97 $Y=2.455 $X2=0
+ $Y2=0
cc_486 N_VPWR_c_555_n N_A_114_368#_c_695_n 0.0449718f $X=2.97 $Y=2.455 $X2=0
+ $Y2=0
cc_487 N_VPWR_c_556_n N_A_114_368#_c_695_n 0.0449718f $X=3.87 $Y=2.455 $X2=0
+ $Y2=0
cc_488 N_VPWR_c_564_n N_A_114_368#_c_695_n 0.00749631f $X=3.705 $Y=3.33 $X2=0
+ $Y2=0
cc_489 N_VPWR_c_550_n N_A_114_368#_c_695_n 0.0062048f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_490 N_VPWR_M1031_d N_A_114_368#_c_728_n 0.00907415f $X=3.72 $Y=1.84 $X2=0
+ $Y2=0
cc_491 N_VPWR_c_556_n N_A_114_368#_c_728_n 0.0171814f $X=3.87 $Y=2.455 $X2=0
+ $Y2=0
cc_492 N_VPWR_c_556_n N_A_114_368#_c_696_n 0.0449718f $X=3.87 $Y=2.455 $X2=0
+ $Y2=0
cc_493 N_VPWR_c_557_n N_A_114_368#_c_696_n 0.0440249f $X=4.77 $Y=2.455 $X2=0
+ $Y2=0
cc_494 N_VPWR_c_566_n N_A_114_368#_c_696_n 0.00749631f $X=4.605 $Y=3.33 $X2=0
+ $Y2=0
cc_495 N_VPWR_c_550_n N_A_114_368#_c_696_n 0.0062048f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_496 N_VPWR_M1013_d N_A_114_368#_c_738_n 0.00384138f $X=4.62 $Y=1.84 $X2=0
+ $Y2=0
cc_497 N_VPWR_c_557_n N_A_114_368#_c_738_n 0.0154248f $X=4.77 $Y=2.455 $X2=0
+ $Y2=0
cc_498 N_VPWR_c_557_n N_A_114_368#_c_697_n 0.0453479f $X=4.77 $Y=2.455 $X2=0
+ $Y2=0
cc_499 N_VPWR_c_558_n N_A_114_368#_c_697_n 0.0110241f $X=5.505 $Y=3.33 $X2=0
+ $Y2=0
cc_500 N_VPWR_c_559_n N_A_114_368#_c_697_n 0.0462948f $X=5.67 $Y=2.455 $X2=0
+ $Y2=0
cc_501 N_VPWR_c_550_n N_A_114_368#_c_697_n 0.00909194f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_502 N_VPWR_M1017_d N_A_114_368#_c_698_n 0.0050953f $X=5.52 $Y=1.84 $X2=0
+ $Y2=0
cc_503 N_VPWR_c_559_n N_A_114_368#_c_698_n 0.0220544f $X=5.67 $Y=2.455 $X2=0
+ $Y2=0
cc_504 N_VPWR_c_559_n N_A_1213_368#_c_811_n 0.045008f $X=5.67 $Y=2.455 $X2=0
+ $Y2=0
cc_505 N_VPWR_c_569_n N_A_1213_368#_c_812_n 0.03588f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_506 N_VPWR_c_550_n N_A_1213_368#_c_812_n 0.0201952f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_507 N_VPWR_c_559_n N_A_1213_368#_c_813_n 0.0139f $X=5.67 $Y=2.455 $X2=0 $Y2=0
cc_508 N_VPWR_c_569_n N_A_1213_368#_c_813_n 0.0236039f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_509 N_VPWR_c_550_n N_A_1213_368#_c_813_n 0.012761f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_510 N_VPWR_c_569_n N_A_1213_368#_c_814_n 0.03588f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_511 N_VPWR_c_550_n N_A_1213_368#_c_814_n 0.0201952f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_512 N_VPWR_c_569_n N_A_1213_368#_c_816_n 0.03588f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_513 N_VPWR_c_550_n N_A_1213_368#_c_816_n 0.0201952f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_514 N_VPWR_c_569_n N_A_1213_368#_c_817_n 0.0594839f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_515 N_VPWR_c_550_n N_A_1213_368#_c_817_n 0.0329562f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_516 N_VPWR_c_569_n N_A_1213_368#_c_819_n 0.0235512f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_517 N_VPWR_c_550_n N_A_1213_368#_c_819_n 0.0126924f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_518 N_VPWR_c_569_n N_A_1213_368#_c_820_n 0.0235512f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_519 N_VPWR_c_550_n N_A_1213_368#_c_820_n 0.0126924f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_520 N_VPWR_c_569_n N_A_1213_368#_c_821_n 0.0235512f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_521 N_VPWR_c_550_n N_A_1213_368#_c_821_n 0.0126924f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_522 N_VPWR_c_552_n N_A_34_74#_c_997_n 0.00754091f $X=0.27 $Y=1.985 $X2=0
+ $Y2=0
cc_523 N_A_114_368#_c_698_n N_A_1213_368#_M1001_s 0.0102914f $X=6.475 $Y=2.035
+ $X2=-0.19 $Y2=1.66
cc_524 N_A_114_368#_c_699_n N_A_1213_368#_M1009_s 0.00201799f $X=7.425 $Y=1.985
+ $X2=0 $Y2=0
cc_525 N_A_114_368#_c_698_n N_A_1213_368#_c_811_n 0.0195484f $X=6.475 $Y=2.035
+ $X2=0 $Y2=0
cc_526 N_A_114_368#_M1001_d N_A_1213_368#_c_812_n 0.00197722f $X=6.49 $Y=1.84
+ $X2=0 $Y2=0
cc_527 N_A_114_368#_c_806_p N_A_1213_368#_c_812_n 0.014157f $X=6.64 $Y=2.57
+ $X2=0 $Y2=0
cc_528 N_A_114_368#_c_699_n N_A_1213_368#_c_828_n 0.0179913f $X=7.425 $Y=1.985
+ $X2=0 $Y2=0
cc_529 N_A_114_368#_M1020_d N_A_1213_368#_c_814_n 0.00197722f $X=7.39 $Y=1.84
+ $X2=0 $Y2=0
cc_530 N_A_114_368#_c_809_p N_A_1213_368#_c_814_n 0.014157f $X=7.54 $Y=2.57
+ $X2=0 $Y2=0
cc_531 N_A_114_368#_c_700_n N_A_1213_368#_c_815_n 0.0133269f $X=7.54 $Y=2.15
+ $X2=0 $Y2=0
cc_532 N_A_1213_368#_c_816_n N_Y_M1015_d 0.00243452f $X=8.725 $Y=2.99 $X2=0
+ $Y2=0
cc_533 N_A_1213_368#_c_817_n N_Y_M1025_d 0.00243452f $X=9.625 $Y=2.99 $X2=0
+ $Y2=0
cc_534 N_A_1213_368#_c_815_n N_Y_c_930_n 0.0550085f $X=7.99 $Y=1.985 $X2=0 $Y2=0
cc_535 N_A_1213_368#_c_816_n N_Y_c_930_n 0.012787f $X=8.725 $Y=2.99 $X2=0 $Y2=0
cc_536 N_A_1213_368#_c_846_n N_Y_c_930_n 0.0439674f $X=8.89 $Y=2.225 $X2=0 $Y2=0
cc_537 N_A_1213_368#_M1022_s N_Y_c_904_n 0.00197722f $X=8.74 $Y=1.84 $X2=0 $Y2=0
cc_538 N_A_1213_368#_c_846_n N_Y_c_904_n 0.0171813f $X=8.89 $Y=2.225 $X2=0 $Y2=0
cc_539 N_A_1213_368#_c_815_n N_Y_c_905_n 0.00513432f $X=7.99 $Y=1.985 $X2=0
+ $Y2=0
cc_540 N_A_1213_368#_c_846_n N_Y_c_945_n 0.0439674f $X=8.89 $Y=2.225 $X2=0 $Y2=0
cc_541 N_A_1213_368#_c_817_n N_Y_c_945_n 0.012787f $X=9.625 $Y=2.99 $X2=0 $Y2=0
cc_542 N_A_1213_368#_c_818_n N_Y_c_945_n 0.0550085f $X=9.79 $Y=1.985 $X2=0 $Y2=0
cc_543 N_A_1213_368#_c_818_n N_Y_c_907_n 0.00513432f $X=9.79 $Y=1.985 $X2=0
+ $Y2=0
cc_544 N_Y_c_900_n N_A_34_74#_c_1006_n 0.0169912f $X=4.66 $Y=0.95 $X2=0 $Y2=0
cc_545 N_Y_c_919_n N_VGND_M1010_d 0.0286593f $X=7.76 $Y=0.925 $X2=0 $Y2=0
cc_546 N_Y_c_949_n N_VGND_M1004_s 0.00330259f $X=8.7 $Y=0.68 $X2=0 $Y2=0
cc_547 N_Y_c_898_n N_VGND_c_1071_n 0.0121972f $X=7.925 $Y=0.515 $X2=0 $Y2=0
cc_548 N_Y_c_949_n N_VGND_c_1071_n 0.0167019f $X=8.7 $Y=0.68 $X2=0 $Y2=0
cc_549 N_Y_c_903_n N_VGND_c_1071_n 0.0122903f $X=9.425 $Y=0.68 $X2=0 $Y2=0
cc_550 N_Y_c_898_n N_VGND_c_1074_n 0.0110175f $X=7.925 $Y=0.515 $X2=0 $Y2=0
cc_551 N_Y_c_903_n N_VGND_c_1075_n 0.0544421f $X=9.425 $Y=0.68 $X2=0 $Y2=0
cc_552 N_Y_c_896_n N_VGND_c_1076_n 0.00789134f $X=6.13 $Y=0.99 $X2=0 $Y2=0
cc_553 N_Y_c_897_n N_VGND_c_1076_n 0.00904371f $X=6.215 $Y=0.515 $X2=0 $Y2=0
cc_554 N_Y_c_919_n N_VGND_c_1076_n 0.0132757f $X=7.76 $Y=0.925 $X2=0 $Y2=0
cc_555 N_Y_c_898_n N_VGND_c_1076_n 0.0090528f $X=7.925 $Y=0.515 $X2=0 $Y2=0
cc_556 N_Y_c_949_n N_VGND_c_1076_n 0.0116543f $X=8.7 $Y=0.68 $X2=0 $Y2=0
cc_557 N_Y_c_903_n N_VGND_c_1076_n 0.0458137f $X=9.425 $Y=0.68 $X2=0 $Y2=0
cc_558 N_Y_c_897_n N_VGND_c_1079_n 0.0109942f $X=6.215 $Y=0.515 $X2=0 $Y2=0
cc_559 N_Y_c_897_n N_VGND_c_1080_n 0.0124113f $X=6.215 $Y=0.515 $X2=0 $Y2=0
cc_560 N_Y_c_919_n N_VGND_c_1080_n 0.0804627f $X=7.76 $Y=0.925 $X2=0 $Y2=0
cc_561 N_Y_c_898_n N_VGND_c_1080_n 0.0124113f $X=7.925 $Y=0.515 $X2=0 $Y2=0
cc_562 N_Y_c_896_n N_A_465_74#_M1007_d 0.00209854f $X=6.13 $Y=0.99 $X2=0 $Y2=0
cc_563 N_Y_c_896_n N_A_465_74#_M1021_d 0.00177318f $X=6.13 $Y=0.99 $X2=0 $Y2=0
cc_564 N_Y_c_896_n N_A_465_74#_c_1161_n 0.0163856f $X=6.13 $Y=0.99 $X2=0 $Y2=0
cc_565 N_Y_c_897_n N_A_465_74#_c_1161_n 0.0135554f $X=6.215 $Y=0.515 $X2=0 $Y2=0
cc_566 N_Y_M1007_s N_A_465_74#_c_1162_n 0.00332037f $X=4.37 $Y=0.37 $X2=0 $Y2=0
cc_567 N_Y_M1012_s N_A_465_74#_c_1162_n 0.00212678f $X=5.215 $Y=0.37 $X2=0 $Y2=0
cc_568 N_Y_c_896_n N_A_465_74#_c_1162_n 0.0379865f $X=6.13 $Y=0.99 $X2=0 $Y2=0
cc_569 N_Y_c_900_n N_A_465_74#_c_1162_n 0.0208358f $X=4.66 $Y=0.95 $X2=0 $Y2=0
cc_570 N_A_34_74#_c_996_n N_VGND_M1003_d 0.00176461f $X=1.01 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_571 N_A_34_74#_c_999_n N_VGND_M1023_d 0.00176461f $X=1.95 $Y=1.095 $X2=0
+ $Y2=0
cc_572 N_A_34_74#_c_995_n N_VGND_c_1069_n 0.0175587f $X=0.315 $Y=0.515 $X2=0
+ $Y2=0
cc_573 N_A_34_74#_c_996_n N_VGND_c_1069_n 0.0152916f $X=1.01 $Y=1.095 $X2=0
+ $Y2=0
cc_574 N_A_34_74#_c_998_n N_VGND_c_1069_n 0.0175587f $X=1.175 $Y=0.515 $X2=0
+ $Y2=0
cc_575 N_A_34_74#_c_998_n N_VGND_c_1070_n 0.0182902f $X=1.175 $Y=0.515 $X2=0
+ $Y2=0
cc_576 N_A_34_74#_c_999_n N_VGND_c_1070_n 0.0170777f $X=1.95 $Y=1.095 $X2=0
+ $Y2=0
cc_577 N_A_34_74#_c_1000_n N_VGND_c_1070_n 0.0182488f $X=2.035 $Y=0.515 $X2=0
+ $Y2=0
cc_578 N_A_34_74#_c_995_n N_VGND_c_1072_n 0.011066f $X=0.315 $Y=0.515 $X2=0
+ $Y2=0
cc_579 N_A_34_74#_c_998_n N_VGND_c_1073_n 0.0109942f $X=1.175 $Y=0.515 $X2=0
+ $Y2=0
cc_580 N_A_34_74#_c_995_n N_VGND_c_1076_n 0.00915947f $X=0.315 $Y=0.515 $X2=0
+ $Y2=0
cc_581 N_A_34_74#_c_998_n N_VGND_c_1076_n 0.00904371f $X=1.175 $Y=0.515 $X2=0
+ $Y2=0
cc_582 N_A_34_74#_c_1000_n N_VGND_c_1076_n 0.0062048f $X=2.035 $Y=0.515 $X2=0
+ $Y2=0
cc_583 N_A_34_74#_c_1000_n N_VGND_c_1079_n 0.00749631f $X=2.035 $Y=0.515 $X2=0
+ $Y2=0
cc_584 N_A_34_74#_c_1004_n N_A_465_74#_M1002_d 0.00229137f $X=2.73 $Y=0.975
+ $X2=-0.19 $Y2=-0.245
cc_585 N_A_34_74#_c_1001_n N_A_465_74#_M1033_d 0.00229137f $X=3.59 $Y=1.077
+ $X2=0 $Y2=0
cc_586 N_A_34_74#_c_1000_n N_A_465_74#_c_1158_n 0.0134146f $X=2.035 $Y=0.515
+ $X2=0 $Y2=0
cc_587 N_A_34_74#_c_1004_n N_A_465_74#_c_1158_n 0.00971408f $X=2.73 $Y=0.975
+ $X2=0 $Y2=0
cc_588 N_A_34_74#_M1011_s N_A_465_74#_c_1159_n 0.00179007f $X=2.755 $Y=0.37
+ $X2=0 $Y2=0
cc_589 N_A_34_74#_c_1001_n N_A_465_74#_c_1159_n 0.00465091f $X=3.59 $Y=1.077
+ $X2=0 $Y2=0
cc_590 N_A_34_74#_c_1004_n N_A_465_74#_c_1159_n 0.00465091f $X=2.73 $Y=0.975
+ $X2=0 $Y2=0
cc_591 N_A_34_74#_c_1005_n N_A_465_74#_c_1159_n 0.0163588f $X=3.06 $Y=0.975
+ $X2=0 $Y2=0
cc_592 N_A_34_74#_c_1001_n N_A_465_74#_c_1160_n 0.00857327f $X=3.59 $Y=1.077
+ $X2=0 $Y2=0
cc_593 N_A_34_74#_M1034_s N_A_465_74#_c_1162_n 0.0033149f $X=3.615 $Y=0.37 $X2=0
+ $Y2=0
cc_594 N_A_34_74#_c_1001_n N_A_465_74#_c_1162_n 0.00466938f $X=3.59 $Y=1.077
+ $X2=0 $Y2=0
cc_595 N_A_34_74#_c_1006_n N_A_465_74#_c_1162_n 0.0209951f $X=3.755 $Y=0.95
+ $X2=0 $Y2=0
cc_596 N_VGND_c_1076_n N_A_465_74#_c_1158_n 0.126157f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_597 N_VGND_c_1079_n N_A_465_74#_c_1158_n 0.149195f $X=6.55 $Y=0.292 $X2=0
+ $Y2=0
