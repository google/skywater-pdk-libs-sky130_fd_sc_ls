# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ls__dfstp_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ls__dfstp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.04000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.475000 0.980000 0.805000 1.990000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.530100 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.500000 0.350000 10.935000 1.050000 ;
        RECT 10.685000 1.050000 10.935000 2.980000 ;
    END
  END Q
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.080000 1.820000 5.635000 2.150000 ;
        RECT 8.185000 1.130000 8.515000 2.140000 ;
      LAYER mcon ;
        RECT 5.435000 1.950000 5.605000 2.120000 ;
        RECT 8.315000 1.950000 8.485000 2.120000 ;
      LAYER met1 ;
        RECT 5.375000 1.920000 5.665000 1.965000 ;
        RECT 5.375000 1.965000 8.545000 2.105000 ;
        RECT 5.375000 2.105000 5.665000 2.150000 ;
        RECT 8.255000 1.920000 8.545000 1.965000 ;
        RECT 8.255000 2.105000 8.545000 2.150000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.315000 1.180000 1.795000 1.550000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 11.040000 0.085000 ;
        RECT  0.545000  0.085000  0.795000 0.810000 ;
        RECT  1.615000  0.085000  1.785000 1.010000 ;
        RECT  4.065000  0.085000  4.455000 0.680000 ;
        RECT  5.620000  0.085000  5.950000 1.030000 ;
        RECT  7.870000  0.085000  8.760000 0.600000 ;
        RECT 10.000000  0.085000 10.330000 1.030000 ;
      LAYER mcon ;
        RECT  0.155000 -0.085000  0.325000 0.085000 ;
        RECT  0.635000 -0.085000  0.805000 0.085000 ;
        RECT  1.115000 -0.085000  1.285000 0.085000 ;
        RECT  1.595000 -0.085000  1.765000 0.085000 ;
        RECT  2.075000 -0.085000  2.245000 0.085000 ;
        RECT  2.555000 -0.085000  2.725000 0.085000 ;
        RECT  3.035000 -0.085000  3.205000 0.085000 ;
        RECT  3.515000 -0.085000  3.685000 0.085000 ;
        RECT  3.995000 -0.085000  4.165000 0.085000 ;
        RECT  4.475000 -0.085000  4.645000 0.085000 ;
        RECT  4.955000 -0.085000  5.125000 0.085000 ;
        RECT  5.435000 -0.085000  5.605000 0.085000 ;
        RECT  5.915000 -0.085000  6.085000 0.085000 ;
        RECT  6.395000 -0.085000  6.565000 0.085000 ;
        RECT  6.875000 -0.085000  7.045000 0.085000 ;
        RECT  7.355000 -0.085000  7.525000 0.085000 ;
        RECT  7.835000 -0.085000  8.005000 0.085000 ;
        RECT  8.315000 -0.085000  8.485000 0.085000 ;
        RECT  8.795000 -0.085000  8.965000 0.085000 ;
        RECT  9.275000 -0.085000  9.445000 0.085000 ;
        RECT  9.755000 -0.085000  9.925000 0.085000 ;
        RECT 10.235000 -0.085000 10.405000 0.085000 ;
        RECT 10.715000 -0.085000 10.885000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 11.040000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 3.245000 11.040000 3.415000 ;
        RECT  0.555000 2.570000  0.885000 3.245000 ;
        RECT  1.540000 2.570000  1.870000 3.245000 ;
        RECT  3.950000 2.425000  4.230000 3.245000 ;
        RECT  5.535000 2.660000  5.785000 3.245000 ;
        RECT  7.770000 2.650000  7.940000 3.245000 ;
        RECT  8.665000 2.650000  8.915000 3.245000 ;
        RECT 10.155000 1.820000 10.485000 3.245000 ;
      LAYER mcon ;
        RECT  0.155000 3.245000  0.325000 3.415000 ;
        RECT  0.635000 3.245000  0.805000 3.415000 ;
        RECT  1.115000 3.245000  1.285000 3.415000 ;
        RECT  1.595000 3.245000  1.765000 3.415000 ;
        RECT  2.075000 3.245000  2.245000 3.415000 ;
        RECT  2.555000 3.245000  2.725000 3.415000 ;
        RECT  3.035000 3.245000  3.205000 3.415000 ;
        RECT  3.515000 3.245000  3.685000 3.415000 ;
        RECT  3.995000 3.245000  4.165000 3.415000 ;
        RECT  4.475000 3.245000  4.645000 3.415000 ;
        RECT  4.955000 3.245000  5.125000 3.415000 ;
        RECT  5.435000 3.245000  5.605000 3.415000 ;
        RECT  5.915000 3.245000  6.085000 3.415000 ;
        RECT  6.395000 3.245000  6.565000 3.415000 ;
        RECT  6.875000 3.245000  7.045000 3.415000 ;
        RECT  7.355000 3.245000  7.525000 3.415000 ;
        RECT  7.835000 3.245000  8.005000 3.415000 ;
        RECT  8.315000 3.245000  8.485000 3.415000 ;
        RECT  8.795000 3.245000  8.965000 3.415000 ;
        RECT  9.275000 3.245000  9.445000 3.415000 ;
        RECT  9.755000 3.245000  9.925000 3.415000 ;
        RECT 10.235000 3.245000 10.405000 3.415000 ;
        RECT 10.715000 3.245000 10.885000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 11.040000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.105000 0.350000  0.365000 0.810000 ;
      RECT 0.105000 0.810000  0.275000 2.230000 ;
      RECT 0.105000 2.230000  1.760000 2.400000 ;
      RECT 0.105000 2.400000  0.355000 2.980000 ;
      RECT 0.975000 0.350000  1.435000 1.010000 ;
      RECT 0.975000 1.010000  1.145000 1.720000 ;
      RECT 0.975000 1.720000  2.315000 1.890000 ;
      RECT 0.975000 1.890000  1.420000 2.060000 ;
      RECT 1.590000 2.060000  2.660000 2.230000 ;
      RECT 1.965000 0.255000  3.075000 0.425000 ;
      RECT 1.965000 0.425000  2.295000 1.090000 ;
      RECT 1.985000 1.260000  2.315000 1.720000 ;
      RECT 2.070000 2.400000  2.320000 2.905000 ;
      RECT 2.070000 2.905000  3.755000 3.075000 ;
      RECT 2.485000 0.595000  2.735000 0.925000 ;
      RECT 2.485000 0.925000  2.660000 2.060000 ;
      RECT 2.490000 2.230000  2.660000 2.295000 ;
      RECT 2.490000 2.295000  2.910000 2.735000 ;
      RECT 2.830000 1.435000  3.075000 2.105000 ;
      RECT 2.905000 0.425000  3.075000 1.435000 ;
      RECT 3.080000 2.295000  3.415000 2.735000 ;
      RECT 3.245000 0.415000  3.575000 0.850000 ;
      RECT 3.245000 0.850000  4.095000 1.020000 ;
      RECT 3.245000 1.020000  3.415000 2.295000 ;
      RECT 3.585000 1.435000  3.755000 2.085000 ;
      RECT 3.585000 2.085000  4.570000 2.255000 ;
      RECT 3.585000 2.255000  3.755000 2.905000 ;
      RECT 3.925000 1.020000  4.095000 1.345000 ;
      RECT 3.925000 1.345000  6.065000 1.515000 ;
      RECT 4.055000 1.685000  4.385000 1.745000 ;
      RECT 4.055000 1.745000  4.910000 1.915000 ;
      RECT 4.265000 0.860000  5.010000 1.030000 ;
      RECT 4.265000 1.030000  4.625000 1.175000 ;
      RECT 4.400000 2.255000  4.570000 2.905000 ;
      RECT 4.400000 2.905000  5.365000 3.075000 ;
      RECT 4.625000 0.570000  5.010000 0.860000 ;
      RECT 4.740000 1.915000  4.910000 2.320000 ;
      RECT 4.740000 2.320000  5.025000 2.735000 ;
      RECT 4.805000 1.215000  6.065000 1.345000 ;
      RECT 4.805000 1.515000  6.065000 1.545000 ;
      RECT 5.195000 2.320000  5.975000 2.490000 ;
      RECT 5.195000 2.490000  5.365000 2.905000 ;
      RECT 5.805000 1.715000  6.405000 1.885000 ;
      RECT 5.805000 1.885000  5.975000 2.320000 ;
      RECT 6.235000 0.255000  7.325000 0.425000 ;
      RECT 6.235000 0.425000  6.405000 1.120000 ;
      RECT 6.235000 1.120000  6.645000 1.450000 ;
      RECT 6.235000 1.450000  6.405000 1.715000 ;
      RECT 6.475000 2.050000  6.810000 2.625000 ;
      RECT 6.475000 2.625000  7.600000 2.980000 ;
      RECT 6.575000 0.595000  6.985000 0.925000 ;
      RECT 6.575000 1.630000  6.985000 1.800000 ;
      RECT 6.575000 1.800000  6.810000 2.050000 ;
      RECT 6.815000 0.925000  6.985000 1.630000 ;
      RECT 6.980000 1.970000  7.325000 2.140000 ;
      RECT 6.980000 2.140000  7.260000 2.355000 ;
      RECT 7.155000 0.425000  7.325000 1.970000 ;
      RECT 7.430000 2.310000  9.105000 2.480000 ;
      RECT 7.430000 2.480000  7.600000 2.625000 ;
      RECT 7.495000 0.790000  9.260000 0.960000 ;
      RECT 7.495000 0.960000  7.730000 1.555000 ;
      RECT 8.140000 2.480000  8.470000 2.930000 ;
      RECT 8.775000 1.370000  9.105000 2.310000 ;
      RECT 8.930000 0.350000  9.260000 0.790000 ;
      RECT 9.090000 0.960000  9.260000 1.030000 ;
      RECT 9.090000 1.030000  9.445000 1.200000 ;
      RECT 9.115000 2.650000  9.445000 2.980000 ;
      RECT 9.275000 1.200000  9.445000 2.650000 ;
      RECT 9.490000 0.350000  9.820000 0.860000 ;
      RECT 9.635000 0.860000  9.820000 1.220000 ;
      RECT 9.635000 1.220000 10.515000 1.550000 ;
      RECT 9.635000 1.550000  9.965000 2.875000 ;
  END
END sky130_fd_sc_ls__dfstp_1
