* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__nand4b_2 A_N B C D VGND VNB VPB VPWR Y
M1000 a_719_123# C a_490_74# VNB nshort w=740000u l=150000u
+  ad=6.22175e+11p pd=6.14e+06u as=5.618e+11p ps=4.6e+06u
M1001 Y C VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=1.344e+12p pd=1.136e+07u as=2.5148e+12p ps=1.571e+07u
M1002 a_225_74# B a_490_74# VNB nshort w=740000u l=150000u
+  ad=6.01175e+11p pd=6.14e+06u as=0p ps=0u
M1003 Y a_27_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR C Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y D VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR a_27_74# Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_225_74# a_27_74# Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.294e+11p ps=2.1e+06u
M1008 VPWR D Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_719_123# D VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=3.946e+11p ps=3.93e+06u
M1010 VGND D a_719_123# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Y B VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_490_74# C a_719_123# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_490_74# B a_225_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR A_N a_27_74# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.95e+11p ps=2.59e+06u
M1015 VGND A_N a_27_74# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1016 VPWR B Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 Y a_27_74# a_225_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
