* File: sky130_fd_sc_ls__sdfsbp_1.pxi.spice
* Created: Wed Sep  2 11:27:37 2020
* 
x_PM_SKY130_FD_SC_LS__SDFSBP_1%A_27_74# N_A_27_74#_M1033_s N_A_27_74#_M1026_s
+ N_A_27_74#_M1036_g N_A_27_74#_c_302_n N_A_27_74#_M1039_g N_A_27_74#_c_297_n
+ N_A_27_74#_c_298_n N_A_27_74#_c_304_n N_A_27_74#_c_305_n N_A_27_74#_c_299_n
+ N_A_27_74#_c_300_n N_A_27_74#_c_306_n N_A_27_74#_c_301_n N_A_27_74#_c_307_n
+ PM_SKY130_FD_SC_LS__SDFSBP_1%A_27_74#
x_PM_SKY130_FD_SC_LS__SDFSBP_1%SCE N_SCE_c_381_n N_SCE_M1033_g N_SCE_c_382_n
+ N_SCE_M1026_g N_SCE_c_383_n N_SCE_M1027_g N_SCE_M1011_g N_SCE_c_384_n
+ N_SCE_c_376_n N_SCE_c_377_n N_SCE_c_378_n SCE N_SCE_c_379_n N_SCE_c_380_n
+ PM_SKY130_FD_SC_LS__SDFSBP_1%SCE
x_PM_SKY130_FD_SC_LS__SDFSBP_1%D N_D_c_453_n N_D_M1014_g N_D_M1037_g D
+ N_D_c_455_n PM_SKY130_FD_SC_LS__SDFSBP_1%D
x_PM_SKY130_FD_SC_LS__SDFSBP_1%SCD N_SCD_c_486_n N_SCD_M1012_g N_SCD_c_490_n
+ N_SCD_M1031_g N_SCD_c_487_n N_SCD_c_488_n SCD SCD SCD
+ PM_SKY130_FD_SC_LS__SDFSBP_1%SCD
x_PM_SKY130_FD_SC_LS__SDFSBP_1%CLK N_CLK_c_529_n N_CLK_M1022_g N_CLK_c_530_n
+ N_CLK_M1019_g CLK PM_SKY130_FD_SC_LS__SDFSBP_1%CLK
x_PM_SKY130_FD_SC_LS__SDFSBP_1%A_781_74# N_A_781_74#_M1020_d N_A_781_74#_M1029_d
+ N_A_781_74#_c_561_n N_A_781_74#_M1017_g N_A_781_74#_M1004_g
+ N_A_781_74#_M1024_g N_A_781_74#_M1035_g N_A_781_74#_c_564_n
+ N_A_781_74#_c_573_n N_A_781_74#_c_565_n N_A_781_74#_c_566_n
+ N_A_781_74#_c_574_n N_A_781_74#_c_575_n N_A_781_74#_c_567_n
+ N_A_781_74#_c_576_n N_A_781_74#_c_577_n N_A_781_74#_c_578_n
+ N_A_781_74#_c_579_n N_A_781_74#_c_580_n N_A_781_74#_c_581_n
+ N_A_781_74#_c_582_n N_A_781_74#_c_583_n N_A_781_74#_c_584_n
+ N_A_781_74#_c_585_n N_A_781_74#_c_586_n N_A_781_74#_c_568_n
+ N_A_781_74#_c_587_n N_A_781_74#_c_569_n N_A_781_74#_c_570_n
+ N_A_781_74#_c_589_n N_A_781_74#_c_590_n PM_SKY130_FD_SC_LS__SDFSBP_1%A_781_74#
x_PM_SKY130_FD_SC_LS__SDFSBP_1%A_1163_48# N_A_1163_48#_M1041_s
+ N_A_1163_48#_M1040_d N_A_1163_48#_c_771_n N_A_1163_48#_M1002_g
+ N_A_1163_48#_c_772_n N_A_1163_48#_c_777_n N_A_1163_48#_c_778_n
+ N_A_1163_48#_M1025_g N_A_1163_48#_c_773_n N_A_1163_48#_c_774_n
+ N_A_1163_48#_c_779_n N_A_1163_48#_c_780_n N_A_1163_48#_c_775_n
+ PM_SKY130_FD_SC_LS__SDFSBP_1%A_1163_48#
x_PM_SKY130_FD_SC_LS__SDFSBP_1%A_995_74# N_A_995_74#_M1034_d N_A_995_74#_M1017_d
+ N_A_995_74#_c_846_n N_A_995_74#_c_847_n N_A_995_74#_c_859_n
+ N_A_995_74#_M1040_g N_A_995_74#_M1041_g N_A_995_74#_c_860_n
+ N_A_995_74#_M1008_g N_A_995_74#_c_849_n N_A_995_74#_M1023_g
+ N_A_995_74#_c_850_n N_A_995_74#_c_851_n N_A_995_74#_c_852_n
+ N_A_995_74#_c_853_n N_A_995_74#_c_854_n N_A_995_74#_c_855_n
+ N_A_995_74#_c_863_n N_A_995_74#_c_856_n N_A_995_74#_c_857_n
+ PM_SKY130_FD_SC_LS__SDFSBP_1%A_995_74#
x_PM_SKY130_FD_SC_LS__SDFSBP_1%SET_B N_SET_B_M1010_g N_SET_B_c_984_n
+ N_SET_B_c_999_n N_SET_B_M1013_g N_SET_B_c_985_n N_SET_B_M1007_g
+ N_SET_B_c_986_n N_SET_B_c_987_n N_SET_B_c_1000_n N_SET_B_c_1001_n
+ N_SET_B_M1015_g N_SET_B_c_988_n N_SET_B_c_1003_n N_SET_B_c_989_n
+ N_SET_B_c_990_n N_SET_B_c_991_n N_SET_B_c_992_n N_SET_B_c_993_n SET_B
+ N_SET_B_c_995_n N_SET_B_c_996_n N_SET_B_c_997_n
+ PM_SKY130_FD_SC_LS__SDFSBP_1%SET_B
x_PM_SKY130_FD_SC_LS__SDFSBP_1%A_594_74# N_A_594_74#_M1022_s N_A_594_74#_M1019_s
+ N_A_594_74#_c_1139_n N_A_594_74#_M1020_g N_A_594_74#_c_1140_n
+ N_A_594_74#_M1029_g N_A_594_74#_c_1141_n N_A_594_74#_c_1142_n
+ N_A_594_74#_c_1143_n N_A_594_74#_c_1154_n N_A_594_74#_c_1155_n
+ N_A_594_74#_M1034_g N_A_594_74#_c_1156_n N_A_594_74#_M1018_g
+ N_A_594_74#_c_1157_n N_A_594_74#_M1000_g N_A_594_74#_M1009_g
+ N_A_594_74#_c_1146_n N_A_594_74#_c_1159_n N_A_594_74#_c_1147_n
+ N_A_594_74#_c_1161_n N_A_594_74#_c_1148_n N_A_594_74#_c_1149_n
+ N_A_594_74#_c_1163_n N_A_594_74#_c_1164_n N_A_594_74#_c_1150_n
+ N_A_594_74#_c_1151_n N_A_594_74#_c_1166_n N_A_594_74#_c_1167_n
+ PM_SKY130_FD_SC_LS__SDFSBP_1%A_594_74#
x_PM_SKY130_FD_SC_LS__SDFSBP_1%A_1924_48# N_A_1924_48#_M1003_d
+ N_A_1924_48#_M1032_s N_A_1924_48#_M1001_g N_A_1924_48#_c_1319_n
+ N_A_1924_48#_c_1332_n N_A_1924_48#_c_1333_n N_A_1924_48#_c_1334_n
+ N_A_1924_48#_M1006_g N_A_1924_48#_c_1320_n N_A_1924_48#_c_1321_n
+ N_A_1924_48#_c_1322_n N_A_1924_48#_c_1335_n N_A_1924_48#_c_1323_n
+ N_A_1924_48#_c_1324_n N_A_1924_48#_c_1325_n N_A_1924_48#_c_1326_n
+ N_A_1924_48#_c_1327_n N_A_1924_48#_c_1336_n N_A_1924_48#_c_1337_n
+ N_A_1924_48#_c_1338_n N_A_1924_48#_c_1328_n N_A_1924_48#_c_1367_n
+ N_A_1924_48#_c_1329_n N_A_1924_48#_c_1330_n
+ PM_SKY130_FD_SC_LS__SDFSBP_1%A_1924_48#
x_PM_SKY130_FD_SC_LS__SDFSBP_1%A_1762_74# N_A_1762_74#_M1024_d
+ N_A_1762_74#_M1035_d N_A_1762_74#_M1015_d N_A_1762_74#_c_1455_n
+ N_A_1762_74#_M1003_g N_A_1762_74#_c_1456_n N_A_1762_74#_c_1470_n
+ N_A_1762_74#_c_1471_n N_A_1762_74#_M1032_g N_A_1762_74#_M1005_g
+ N_A_1762_74#_c_1458_n N_A_1762_74#_c_1459_n N_A_1762_74#_c_1474_n
+ N_A_1762_74#_M1038_g N_A_1762_74#_c_1460_n N_A_1762_74#_M1016_g
+ N_A_1762_74#_c_1476_n N_A_1762_74#_M1030_g N_A_1762_74#_c_1462_n
+ N_A_1762_74#_c_1463_n N_A_1762_74#_c_1464_n N_A_1762_74#_c_1465_n
+ N_A_1762_74#_c_1466_n N_A_1762_74#_c_1481_n N_A_1762_74#_c_1482_n
+ N_A_1762_74#_c_1467_n N_A_1762_74#_c_1568_n N_A_1762_74#_c_1468_n
+ N_A_1762_74#_c_1484_n N_A_1762_74#_c_1469_n N_A_1762_74#_c_1486_n
+ N_A_1762_74#_c_1487_n N_A_1762_74#_c_1488_n
+ PM_SKY130_FD_SC_LS__SDFSBP_1%A_1762_74#
x_PM_SKY130_FD_SC_LS__SDFSBP_1%A_2556_112# N_A_2556_112#_M1016_s
+ N_A_2556_112#_M1030_s N_A_2556_112#_c_1654_n N_A_2556_112#_M1021_g
+ N_A_2556_112#_M1028_g N_A_2556_112#_c_1649_n N_A_2556_112#_c_1650_n
+ N_A_2556_112#_c_1651_n N_A_2556_112#_c_1652_n N_A_2556_112#_c_1653_n
+ PM_SKY130_FD_SC_LS__SDFSBP_1%A_2556_112#
x_PM_SKY130_FD_SC_LS__SDFSBP_1%VPWR N_VPWR_M1026_d N_VPWR_M1031_d N_VPWR_M1019_d
+ N_VPWR_M1025_d N_VPWR_M1013_d N_VPWR_M1006_d N_VPWR_M1032_d N_VPWR_M1030_d
+ N_VPWR_c_1696_n N_VPWR_c_1697_n N_VPWR_c_1698_n N_VPWR_c_1699_n
+ N_VPWR_c_1700_n N_VPWR_c_1701_n N_VPWR_c_1702_n N_VPWR_c_1703_n
+ N_VPWR_c_1704_n N_VPWR_c_1705_n N_VPWR_c_1706_n N_VPWR_c_1707_n
+ N_VPWR_c_1708_n N_VPWR_c_1709_n N_VPWR_c_1710_n VPWR N_VPWR_c_1711_n
+ N_VPWR_c_1712_n N_VPWR_c_1713_n N_VPWR_c_1714_n N_VPWR_c_1715_n
+ N_VPWR_c_1695_n N_VPWR_c_1717_n N_VPWR_c_1718_n N_VPWR_c_1719_n
+ N_VPWR_c_1720_n N_VPWR_c_1721_n PM_SKY130_FD_SC_LS__SDFSBP_1%VPWR
x_PM_SKY130_FD_SC_LS__SDFSBP_1%A_290_464# N_A_290_464#_M1037_d
+ N_A_290_464#_M1034_s N_A_290_464#_M1014_d N_A_290_464#_M1017_s
+ N_A_290_464#_c_1869_n N_A_290_464#_c_1856_n N_A_290_464#_c_1857_n
+ N_A_290_464#_c_1858_n N_A_290_464#_c_1872_n N_A_290_464#_c_1859_n
+ N_A_290_464#_c_1876_n N_A_290_464#_c_1863_n N_A_290_464#_c_1864_n
+ N_A_290_464#_c_1860_n N_A_290_464#_c_1866_n N_A_290_464#_c_1877_n
+ N_A_290_464#_c_1879_n N_A_290_464#_c_1950_n N_A_290_464#_c_1861_n
+ N_A_290_464#_c_1867_n PM_SKY130_FD_SC_LS__SDFSBP_1%A_290_464#
x_PM_SKY130_FD_SC_LS__SDFSBP_1%A_1600_347# N_A_1600_347#_M1008_d
+ N_A_1600_347#_M1009_d N_A_1600_347#_c_1982_n N_A_1600_347#_c_1983_n
+ N_A_1600_347#_c_1984_n PM_SKY130_FD_SC_LS__SDFSBP_1%A_1600_347#
x_PM_SKY130_FD_SC_LS__SDFSBP_1%A_1712_374# N_A_1712_374#_M1035_s
+ N_A_1712_374#_M1006_s N_A_1712_374#_c_2018_n N_A_1712_374#_c_2019_n
+ N_A_1712_374#_c_2020_n PM_SKY130_FD_SC_LS__SDFSBP_1%A_1712_374#
x_PM_SKY130_FD_SC_LS__SDFSBP_1%Q_N N_Q_N_M1005_d N_Q_N_M1038_d N_Q_N_c_2055_n
+ N_Q_N_c_2056_n N_Q_N_c_2052_n Q_N Q_N Q_N PM_SKY130_FD_SC_LS__SDFSBP_1%Q_N
x_PM_SKY130_FD_SC_LS__SDFSBP_1%Q N_Q_M1028_d N_Q_M1021_d Q Q Q Q Q Q Q
+ PM_SKY130_FD_SC_LS__SDFSBP_1%Q
x_PM_SKY130_FD_SC_LS__SDFSBP_1%VGND N_VGND_M1033_d N_VGND_M1012_d N_VGND_M1022_d
+ N_VGND_M1002_d N_VGND_M1010_d N_VGND_M1007_d N_VGND_M1005_s N_VGND_M1016_d
+ N_VGND_c_2101_n N_VGND_c_2102_n N_VGND_c_2103_n N_VGND_c_2104_n
+ N_VGND_c_2105_n N_VGND_c_2106_n N_VGND_c_2107_n N_VGND_c_2108_n
+ N_VGND_c_2109_n N_VGND_c_2110_n VGND N_VGND_c_2111_n N_VGND_c_2112_n
+ N_VGND_c_2113_n N_VGND_c_2114_n N_VGND_c_2115_n N_VGND_c_2116_n
+ N_VGND_c_2117_n N_VGND_c_2118_n N_VGND_c_2119_n N_VGND_c_2120_n
+ N_VGND_c_2121_n N_VGND_c_2122_n N_VGND_c_2123_n N_VGND_c_2124_n
+ PM_SKY130_FD_SC_LS__SDFSBP_1%VGND
cc_1 VNB N_A_27_74#_M1036_g 0.0215636f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=0.58
cc_2 VNB N_A_27_74#_c_297_n 0.0260478f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=0.58
cc_3 VNB N_A_27_74#_c_298_n 0.0186355f $X=-0.19 $Y=-0.245 $X2=0.225 $Y2=2.29
cc_4 VNB N_A_27_74#_c_299_n 0.0084149f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.115
cc_5 VNB N_A_27_74#_c_300_n 0.0327363f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.115
cc_6 VNB N_A_27_74#_c_301_n 0.0182839f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.115
cc_7 VNB N_SCE_M1033_g 0.0641507f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_SCE_M1011_g 0.035064f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_SCE_c_376_n 0.0234769f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=2.46
cc_10 VNB N_SCE_c_377_n 0.00280342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_SCE_c_378_n 0.0318809f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=2.375
cc_12 VNB N_SCE_c_379_n 0.0201092f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.995
cc_13 VNB N_SCE_c_380_n 0.00254062f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=0.95
cc_14 VNB N_D_M1037_g 0.062081f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_SCD_c_486_n 0.0176451f $X=-0.19 $Y=-0.245 $X2=0.135 $Y2=0.37
cc_16 VNB N_SCD_c_487_n 0.0589035f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=0.95
cc_17 VNB N_SCD_c_488_n 0.0257799f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=0.58
cc_18 VNB SCD 0.00577239f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=0.58
cc_19 VNB N_CLK_c_529_n 0.0191493f $X=-0.19 $Y=-0.245 $X2=0.135 $Y2=0.37
cc_20 VNB N_CLK_c_530_n 0.0430831f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB CLK 0.00704257f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=0.95
cc_22 VNB N_A_781_74#_c_561_n 0.0279286f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=0.95
cc_23 VNB N_A_781_74#_M1004_g 0.0623484f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=0.95
cc_24 VNB N_A_781_74#_M1024_g 0.0315835f $X=-0.19 $Y=-0.245 $X2=0.225 $Y2=1.28
cc_25 VNB N_A_781_74#_c_564_n 0.00580499f $X=-0.19 $Y=-0.245 $X2=0.365 $Y2=2.375
cc_26 VNB N_A_781_74#_c_565_n 0.0155903f $X=-0.19 $Y=-0.245 $X2=1.92 $Y2=2.29
cc_27 VNB N_A_781_74#_c_566_n 0.00279267f $X=-0.19 $Y=-0.245 $X2=1.92 $Y2=1.995
cc_28 VNB N_A_781_74#_c_567_n 0.0011848f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_781_74#_c_568_n 0.00602655f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_781_74#_c_569_n 0.00206749f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_781_74#_c_570_n 0.0289989f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_1163_48#_c_771_n 0.0183276f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=0.95
cc_33 VNB N_A_1163_48#_c_772_n 0.00595723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_1163_48#_c_773_n 0.0254327f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=0.58
cc_35 VNB N_A_1163_48#_c_774_n 0.0220946f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_1163_48#_c_775_n 0.0607898f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.995
cc_37 VNB N_A_995_74#_c_846_n 0.0386116f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=0.95
cc_38 VNB N_A_995_74#_c_847_n 0.00326225f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=0.58
cc_39 VNB N_A_995_74#_M1041_g 0.0341535f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=0.95
cc_40 VNB N_A_995_74#_c_849_n 0.0189909f $X=-0.19 $Y=-0.245 $X2=0.225 $Y2=2.29
cc_41 VNB N_A_995_74#_c_850_n 0.00687291f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=2.375
cc_42 VNB N_A_995_74#_c_851_n 0.00207814f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.115
cc_43 VNB N_A_995_74#_c_852_n 0.0252332f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.115
cc_44 VNB N_A_995_74#_c_853_n 0.0198101f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_995_74#_c_854_n 0.00264222f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.995
cc_46 VNB N_A_995_74#_c_855_n 0.0646933f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_995_74#_c_856_n 0.00350923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_995_74#_c_857_n 0.0124973f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_SET_B_M1010_g 0.0406873f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_SET_B_c_984_n 0.00252704f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_SET_B_c_985_n 0.018015f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_SET_B_c_986_n 0.0242576f $X=-0.19 $Y=-0.245 $X2=2.005 $Y2=2.64
cc_53 VNB N_SET_B_c_987_n 0.00843777f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=0.95
cc_54 VNB N_SET_B_c_988_n 0.0174838f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=2.375
cc_55 VNB N_SET_B_c_989_n 0.00206835f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.115
cc_56 VNB N_SET_B_c_990_n 0.0249121f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.115
cc_57 VNB N_SET_B_c_991_n 0.00828735f $X=-0.19 $Y=-0.245 $X2=1.92 $Y2=2.29
cc_58 VNB N_SET_B_c_992_n 0.0184503f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.995
cc_59 VNB N_SET_B_c_993_n 0.00180662f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.995
cc_60 VNB SET_B 0.00199056f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=0.95
cc_61 VNB N_SET_B_c_995_n 0.0274525f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_SET_B_c_996_n 0.00167402f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_SET_B_c_997_n 0.0163976f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_594_74#_c_1139_n 0.0206133f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=0.95
cc_65 VNB N_A_594_74#_c_1140_n 0.0262063f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_594_74#_c_1141_n 0.0266552f $X=-0.19 $Y=-0.245 $X2=2.005 $Y2=2.64
cc_67 VNB N_A_594_74#_c_1142_n 0.00499256f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=0.58
cc_68 VNB N_A_594_74#_c_1143_n 0.028937f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_594_74#_M1034_g 0.0243464f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_594_74#_M1000_g 0.0562556f $X=-0.19 $Y=-0.245 $X2=1.92 $Y2=1.995
cc_71 VNB N_A_594_74#_c_1146_n 0.0256095f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.115
cc_72 VNB N_A_594_74#_c_1147_n 0.00599737f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_594_74#_c_1148_n 0.00880724f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_594_74#_c_1149_n 0.0115805f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_594_74#_c_1150_n 0.00306961f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_594_74#_c_1151_n 0.0016464f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_1924_48#_c_1319_n 0.0161449f $X=-0.19 $Y=-0.245 $X2=2.005
+ $Y2=2.245
cc_78 VNB N_A_1924_48#_c_1320_n 0.0183699f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_1924_48#_c_1321_n 0.0165713f $X=-0.19 $Y=-0.245 $X2=0.225 $Y2=1.28
cc_80 VNB N_A_1924_48#_c_1322_n 0.0230002f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=2.465
cc_81 VNB N_A_1924_48#_c_1323_n 0.0243895f $X=-0.19 $Y=-0.245 $X2=1.795
+ $Y2=2.375
cc_82 VNB N_A_1924_48#_c_1324_n 0.007537f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.115
cc_83 VNB N_A_1924_48#_c_1325_n 0.00286542f $X=-0.19 $Y=-0.245 $X2=1.92 $Y2=2.29
cc_84 VNB N_A_1924_48#_c_1326_n 0.02238f $X=-0.19 $Y=-0.245 $X2=1.92 $Y2=1.995
cc_85 VNB N_A_1924_48#_c_1327_n 0.00154245f $X=-0.19 $Y=-0.245 $X2=1.96
+ $Y2=1.995
cc_86 VNB N_A_1924_48#_c_1328_n 0.00143741f $X=-0.19 $Y=-0.245 $X2=1.96
+ $Y2=1.995
cc_87 VNB N_A_1924_48#_c_1329_n 0.0181664f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_1924_48#_c_1330_n 0.00510964f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_1762_74#_c_1455_n 0.0200354f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_1762_74#_c_1456_n 0.0358613f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=0.95
cc_91 VNB N_A_1762_74#_M1005_g 0.0507407f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.465
cc_92 VNB N_A_1762_74#_c_1458_n 0.00339118f $X=-0.19 $Y=-0.245 $X2=1.795
+ $Y2=2.375
cc_93 VNB N_A_1762_74#_c_1459_n 0.00451186f $X=-0.19 $Y=-0.245 $X2=0.365
+ $Y2=2.375
cc_94 VNB N_A_1762_74#_c_1460_n 0.0212456f $X=-0.19 $Y=-0.245 $X2=0.975
+ $Y2=1.115
cc_95 VNB N_A_1762_74#_M1016_g 0.0436388f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.995
cc_96 VNB N_A_1762_74#_c_1462_n 0.0283734f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_1762_74#_c_1463_n 0.00147097f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_A_1762_74#_c_1464_n 0.0100433f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_A_1762_74#_c_1465_n 0.00551873f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_A_1762_74#_c_1466_n 0.00171038f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_A_1762_74#_c_1467_n 0.00153994f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_A_1762_74#_c_1468_n 0.00938966f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_A_1762_74#_c_1469_n 0.00483919f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_A_2556_112#_c_1649_n 0.0615125f $X=-0.19 $Y=-0.245 $X2=0.28
+ $Y2=0.95
cc_105 VNB N_A_2556_112#_c_1650_n 0.023668f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=0.58
cc_106 VNB N_A_2556_112#_c_1651_n 0.0138984f $X=-0.19 $Y=-0.245 $X2=0.28
+ $Y2=0.58
cc_107 VNB N_A_2556_112#_c_1652_n 0.0023636f $X=-0.19 $Y=-0.245 $X2=0.225
+ $Y2=1.28
cc_108 VNB N_A_2556_112#_c_1653_n 0.0096015f $X=-0.19 $Y=-0.245 $X2=0.28
+ $Y2=2.465
cc_109 VNB N_VPWR_c_1695_n 0.601534f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_A_290_464#_c_1856_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0.225
+ $Y2=2.29
cc_111 VNB N_A_290_464#_c_1857_n 0.0125835f $X=-0.19 $Y=-0.245 $X2=0.24
+ $Y2=2.465
cc_112 VNB N_A_290_464#_c_1858_n 0.0033344f $X=-0.19 $Y=-0.245 $X2=0.28
+ $Y2=2.465
cc_113 VNB N_A_290_464#_c_1859_n 0.0044818f $X=-0.19 $Y=-0.245 $X2=0.445
+ $Y2=1.115
cc_114 VNB N_A_290_464#_c_1860_n 0.00566544f $X=-0.19 $Y=-0.245 $X2=1.96
+ $Y2=1.995
cc_115 VNB N_A_290_464#_c_1861_n 0.00460204f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_Q_N_c_2052_n 0.0103864f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=0.58
cc_117 VNB Q_N 0.0150197f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=0.58
cc_118 VNB Q_N 0.00781016f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.115
cc_119 VNB Q 0.0547356f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=0.95
cc_120 VNB N_VGND_c_2101_n 0.00982527f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.115
cc_121 VNB N_VGND_c_2102_n 0.0109164f $X=-0.19 $Y=-0.245 $X2=1.92 $Y2=2.29
cc_122 VNB N_VGND_c_2103_n 0.00600048f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB N_VGND_c_2104_n 0.0120969f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=0.95
cc_124 VNB N_VGND_c_2105_n 0.0194709f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_2106_n 0.0169908f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_2107_n 0.0411304f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_VGND_c_2108_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_2109_n 0.0596655f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_2110_n 0.00670466f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_2111_n 0.0191515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_2112_n 0.0207541f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_VGND_c_2113_n 0.0583309f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_VGND_c_2114_n 0.0206359f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_VGND_c_2115_n 0.0415877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_VGND_c_2116_n 0.0191124f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_VGND_c_2117_n 0.816858f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_VGND_c_2118_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB N_VGND_c_2119_n 0.00615422f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VNB N_VGND_c_2120_n 0.0324822f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_VGND_c_2121_n 0.0266754f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_141 VNB N_VGND_c_2122_n 0.0210309f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_142 VNB N_VGND_c_2123_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_143 VNB N_VGND_c_2124_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_144 VPB N_A_27_74#_c_302_n 0.0541961f $X=-0.19 $Y=1.66 $X2=2.005 $Y2=2.245
cc_145 VPB N_A_27_74#_c_298_n 0.031974f $X=-0.19 $Y=1.66 $X2=0.225 $Y2=2.29
cc_146 VPB N_A_27_74#_c_304_n 0.0214709f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.465
cc_147 VPB N_A_27_74#_c_305_n 0.012344f $X=-0.19 $Y=1.66 $X2=1.795 $Y2=2.375
cc_148 VPB N_A_27_74#_c_306_n 0.0031701f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=1.995
cc_149 VPB N_A_27_74#_c_307_n 0.00836023f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=2.375
cc_150 VPB N_SCE_c_381_n 0.0178302f $X=-0.19 $Y=1.66 $X2=0.135 $Y2=2.32
cc_151 VPB N_SCE_c_382_n 0.0245127f $X=-0.19 $Y=1.66 $X2=1.065 $Y2=0.95
cc_152 VPB N_SCE_c_383_n 0.0247295f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_153 VPB N_SCE_c_384_n 0.0119787f $X=-0.19 $Y=1.66 $X2=0.225 $Y2=2.29
cc_154 VPB N_SCE_c_379_n 0.0291654f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=1.995
cc_155 VPB N_SCE_c_380_n 0.00166152f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=0.95
cc_156 VPB N_D_c_453_n 0.0524344f $X=-0.19 $Y=1.66 $X2=0.135 $Y2=0.37
cc_157 VPB N_D_M1037_g 0.00913433f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_158 VPB N_D_c_455_n 0.00879535f $X=-0.19 $Y=1.66 $X2=2.005 $Y2=2.64
cc_159 VPB N_SCD_c_490_n 0.05567f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_160 VPB N_SCD_c_488_n 0.0258678f $X=-0.19 $Y=1.66 $X2=1.065 $Y2=0.58
cc_161 VPB SCD 0.00195322f $X=-0.19 $Y=1.66 $X2=1.065 $Y2=0.58
cc_162 VPB N_CLK_c_530_n 0.0259476f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_163 VPB N_A_781_74#_c_561_n 0.057004f $X=-0.19 $Y=1.66 $X2=1.065 $Y2=0.95
cc_164 VPB N_A_781_74#_M1004_g 0.00176557f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=0.95
cc_165 VPB N_A_781_74#_c_573_n 0.0032477f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.115
cc_166 VPB N_A_781_74#_c_574_n 0.0227564f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=1.995
cc_167 VPB N_A_781_74#_c_575_n 0.00300349f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=1.995
cc_168 VPB N_A_781_74#_c_576_n 0.0012556f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=2.375
cc_169 VPB N_A_781_74#_c_577_n 0.00866264f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_170 VPB N_A_781_74#_c_578_n 0.00151842f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_171 VPB N_A_781_74#_c_579_n 0.0238633f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_172 VPB N_A_781_74#_c_580_n 0.00244172f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_173 VPB N_A_781_74#_c_581_n 0.0158392f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_174 VPB N_A_781_74#_c_582_n 0.00177503f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_175 VPB N_A_781_74#_c_583_n 0.00331582f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_176 VPB N_A_781_74#_c_584_n 0.0108876f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_177 VPB N_A_781_74#_c_585_n 0.00198955f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_178 VPB N_A_781_74#_c_586_n 0.00110243f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_179 VPB N_A_781_74#_c_587_n 0.0375924f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_180 VPB N_A_781_74#_c_570_n 0.0156063f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_181 VPB N_A_781_74#_c_589_n 0.0209911f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_182 VPB N_A_781_74#_c_590_n 0.0166888f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_183 VPB N_A_1163_48#_c_772_n 0.026024f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_184 VPB N_A_1163_48#_c_777_n 0.0121868f $X=-0.19 $Y=1.66 $X2=2.005 $Y2=2.245
cc_185 VPB N_A_1163_48#_c_778_n 0.0218752f $X=-0.19 $Y=1.66 $X2=2.005 $Y2=2.64
cc_186 VPB N_A_1163_48#_c_779_n 0.0122379f $X=-0.19 $Y=1.66 $X2=0.225 $Y2=2.29
cc_187 VPB N_A_1163_48#_c_780_n 0.00796129f $X=-0.19 $Y=1.66 $X2=0.445 $Y2=1.115
cc_188 VPB N_A_995_74#_c_847_n 0.0290728f $X=-0.19 $Y=1.66 $X2=1.065 $Y2=0.58
cc_189 VPB N_A_995_74#_c_859_n 0.021231f $X=-0.19 $Y=1.66 $X2=1.065 $Y2=0.58
cc_190 VPB N_A_995_74#_c_860_n 0.0155299f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=0.58
cc_191 VPB N_A_995_74#_c_851_n 0.00921853f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.115
cc_192 VPB N_A_995_74#_c_855_n 0.0076642f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_193 VPB N_A_995_74#_c_863_n 6.03504e-19 $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.115
cc_194 VPB N_SET_B_c_984_n 0.0304546f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_195 VPB N_SET_B_c_999_n 0.0198914f $X=-0.19 $Y=1.66 $X2=1.065 $Y2=0.95
cc_196 VPB N_SET_B_c_1000_n 0.030436f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=2.46
cc_197 VPB N_SET_B_c_1001_n 0.0261518f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=2.465
cc_198 VPB N_SET_B_c_988_n 0.00938523f $X=-0.19 $Y=1.66 $X2=1.795 $Y2=2.375
cc_199 VPB N_SET_B_c_1003_n 0.0223163f $X=-0.19 $Y=1.66 $X2=0.365 $Y2=2.375
cc_200 VPB N_SET_B_c_989_n 0.00200906f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.115
cc_201 VPB N_SET_B_c_991_n 0.00616409f $X=-0.19 $Y=1.66 $X2=1.92 $Y2=2.29
cc_202 VPB N_SET_B_c_992_n 0.0153051f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=1.995
cc_203 VPB N_SET_B_c_993_n 0.00200016f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=1.995
cc_204 VPB SET_B 0.00172634f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=0.95
cc_205 VPB N_SET_B_c_995_n 0.00506136f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_206 VPB N_SET_B_c_996_n 0.00239196f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_207 VPB N_A_594_74#_c_1140_n 0.0211645f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_208 VPB N_A_594_74#_c_1142_n 0.073806f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=0.58
cc_209 VPB N_A_594_74#_c_1154_n 0.0626965f $X=-0.19 $Y=1.66 $X2=0.225 $Y2=2.29
cc_210 VPB N_A_594_74#_c_1155_n 0.012371f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=2.46
cc_211 VPB N_A_594_74#_c_1156_n 0.0148406f $X=-0.19 $Y=1.66 $X2=0.365 $Y2=2.375
cc_212 VPB N_A_594_74#_c_1157_n 0.280761f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.115
cc_213 VPB N_A_594_74#_M1009_g 0.00938516f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=2.375
cc_214 VPB N_A_594_74#_c_1159_n 0.0250393f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=1.995
cc_215 VPB N_A_594_74#_c_1147_n 0.0125719f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_216 VPB N_A_594_74#_c_1161_n 0.0250273f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_217 VPB N_A_594_74#_c_1149_n 0.00355531f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_218 VPB N_A_594_74#_c_1163_n 0.00550874f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_219 VPB N_A_594_74#_c_1164_n 0.0043601f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_220 VPB N_A_594_74#_c_1150_n 0.00165316f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_221 VPB N_A_594_74#_c_1166_n 0.00586251f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_222 VPB N_A_594_74#_c_1167_n 0.00108998f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_223 VPB N_A_1924_48#_c_1319_n 0.0311874f $X=-0.19 $Y=1.66 $X2=2.005 $Y2=2.245
cc_224 VPB N_A_1924_48#_c_1332_n 0.0214933f $X=-0.19 $Y=1.66 $X2=2.005 $Y2=2.64
cc_225 VPB N_A_1924_48#_c_1333_n 0.0111365f $X=-0.19 $Y=1.66 $X2=2.005 $Y2=2.64
cc_226 VPB N_A_1924_48#_c_1334_n 0.0183376f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=0.95
cc_227 VPB N_A_1924_48#_c_1335_n 0.0212763f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.465
cc_228 VPB N_A_1924_48#_c_1336_n 0.0104353f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=1.115
cc_229 VPB N_A_1924_48#_c_1337_n 0.00493064f $X=-0.19 $Y=1.66 $X2=0.975
+ $Y2=1.115
cc_230 VPB N_A_1924_48#_c_1338_n 0.00379531f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=0.95
cc_231 VPB N_A_1924_48#_c_1328_n 9.10193e-19 $X=-0.19 $Y=1.66 $X2=1.96 $Y2=1.995
cc_232 VPB N_A_1762_74#_c_1470_n 0.0178657f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=0.58
cc_233 VPB N_A_1762_74#_c_1471_n 0.0252856f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_234 VPB N_A_1762_74#_c_1458_n 0.00412669f $X=-0.19 $Y=1.66 $X2=1.795
+ $Y2=2.375
cc_235 VPB N_A_1762_74#_c_1459_n 0.0238984f $X=-0.19 $Y=1.66 $X2=0.365 $Y2=2.375
cc_236 VPB N_A_1762_74#_c_1474_n 0.0196801f $X=-0.19 $Y=1.66 $X2=0.445 $Y2=1.115
cc_237 VPB N_A_1762_74#_c_1460_n 0.0287625f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.115
cc_238 VPB N_A_1762_74#_c_1476_n 0.016399f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_239 VPB N_A_1762_74#_c_1463_n 0.0155417f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_240 VPB N_A_1762_74#_c_1464_n 0.0280916f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_241 VPB N_A_1762_74#_c_1465_n 0.00167153f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_242 VPB N_A_1762_74#_c_1466_n 0.0344909f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_243 VPB N_A_1762_74#_c_1481_n 0.00241768f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_244 VPB N_A_1762_74#_c_1482_n 0.0173499f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_245 VPB N_A_1762_74#_c_1467_n 0.00744762f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_246 VPB N_A_1762_74#_c_1484_n 0.00199416f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_247 VPB N_A_1762_74#_c_1469_n 9.77871e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_248 VPB N_A_1762_74#_c_1486_n 0.00354986f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_249 VPB N_A_1762_74#_c_1487_n 0.00808335f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_250 VPB N_A_1762_74#_c_1488_n 0.00551334f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_251 VPB N_A_2556_112#_c_1654_n 0.0206843f $X=-0.19 $Y=1.66 $X2=1.065 $Y2=0.95
cc_252 VPB N_A_2556_112#_c_1649_n 0.00928611f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=0.95
cc_253 VPB N_A_2556_112#_c_1652_n 0.0159542f $X=-0.19 $Y=1.66 $X2=0.225 $Y2=1.28
cc_254 VPB N_VPWR_c_1696_n 0.00396467f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.115
cc_255 VPB N_VPWR_c_1697_n 0.00991012f $X=-0.19 $Y=1.66 $X2=1.92 $Y2=2.29
cc_256 VPB N_VPWR_c_1698_n 0.023804f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=1.995
cc_257 VPB N_VPWR_c_1699_n 0.00396467f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=2.375
cc_258 VPB N_VPWR_c_1700_n 0.00560285f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=1.995
cc_259 VPB N_VPWR_c_1701_n 0.0124734f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_260 VPB N_VPWR_c_1702_n 0.0095499f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_261 VPB N_VPWR_c_1703_n 0.00731223f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_262 VPB N_VPWR_c_1704_n 0.0117659f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_263 VPB N_VPWR_c_1705_n 0.0546187f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_264 VPB N_VPWR_c_1706_n 0.00330333f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_265 VPB N_VPWR_c_1707_n 0.027717f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_266 VPB N_VPWR_c_1708_n 0.00223798f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_267 VPB N_VPWR_c_1709_n 0.0685263f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_268 VPB N_VPWR_c_1710_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_269 VPB N_VPWR_c_1711_n 0.0180274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_270 VPB N_VPWR_c_1712_n 0.0463631f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_271 VPB N_VPWR_c_1713_n 0.0334651f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_272 VPB N_VPWR_c_1714_n 0.0337745f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_273 VPB N_VPWR_c_1715_n 0.0191124f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_274 VPB N_VPWR_c_1695_n 0.137153f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_275 VPB N_VPWR_c_1717_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_276 VPB N_VPWR_c_1718_n 0.00507132f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_277 VPB N_VPWR_c_1719_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_278 VPB N_VPWR_c_1720_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_279 VPB N_VPWR_c_1721_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_280 VPB N_A_290_464#_c_1859_n 0.00530348f $X=-0.19 $Y=1.66 $X2=0.445
+ $Y2=1.115
cc_281 VPB N_A_290_464#_c_1863_n 0.0131901f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.115
cc_282 VPB N_A_290_464#_c_1864_n 0.00351062f $X=-0.19 $Y=1.66 $X2=1.92 $Y2=2.29
cc_283 VPB N_A_290_464#_c_1860_n 0.00402833f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=1.995
cc_284 VPB N_A_290_464#_c_1866_n 0.00473178f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=2.375
cc_285 VPB N_A_290_464#_c_1867_n 0.00812315f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_286 VPB N_A_1600_347#_c_1982_n 0.0116038f $X=-0.19 $Y=1.66 $X2=1.065 $Y2=0.95
cc_287 VPB N_A_1600_347#_c_1983_n 0.0115665f $X=-0.19 $Y=1.66 $X2=1.065 $Y2=0.58
cc_288 VPB N_A_1600_347#_c_1984_n 0.00552071f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=0.58
cc_289 VPB N_A_1712_374#_c_2018_n 0.0265118f $X=-0.19 $Y=1.66 $X2=1.065 $Y2=0.95
cc_290 VPB N_A_1712_374#_c_2019_n 0.0067911f $X=-0.19 $Y=1.66 $X2=2.005
+ $Y2=2.245
cc_291 VPB N_A_1712_374#_c_2020_n 0.0165386f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=0.95
cc_292 VPB N_Q_N_c_2055_n 0.00106684f $X=-0.19 $Y=1.66 $X2=1.065 $Y2=0.58
cc_293 VPB N_Q_N_c_2056_n 0.0023452f $X=-0.19 $Y=1.66 $X2=2.005 $Y2=2.245
cc_294 VPB N_Q_N_c_2052_n 5.04282e-19 $X=-0.19 $Y=1.66 $X2=0.28 $Y2=0.58
cc_295 VPB Q 0.0538644f $X=-0.19 $Y=1.66 $X2=1.065 $Y2=0.95
cc_296 N_A_27_74#_M1036_g N_SCE_M1033_g 0.0154087f $X=1.065 $Y=0.58 $X2=0 $Y2=0
cc_297 N_A_27_74#_c_297_n N_SCE_M1033_g 0.0123507f $X=0.28 $Y=0.58 $X2=0 $Y2=0
cc_298 N_A_27_74#_c_298_n N_SCE_M1033_g 0.00803467f $X=0.225 $Y=2.29 $X2=0 $Y2=0
cc_299 N_A_27_74#_c_299_n N_SCE_M1033_g 0.0168544f $X=0.975 $Y=1.115 $X2=0 $Y2=0
cc_300 N_A_27_74#_c_300_n N_SCE_M1033_g 0.0180926f $X=0.975 $Y=1.115 $X2=0 $Y2=0
cc_301 N_A_27_74#_c_301_n N_SCE_M1033_g 0.00874187f $X=0.28 $Y=1.115 $X2=0 $Y2=0
cc_302 N_A_27_74#_c_298_n N_SCE_c_382_n 0.00168508f $X=0.225 $Y=2.29 $X2=0 $Y2=0
cc_303 N_A_27_74#_c_304_n N_SCE_c_382_n 0.00517645f $X=0.28 $Y=2.465 $X2=0 $Y2=0
cc_304 N_A_27_74#_c_305_n N_SCE_c_382_n 0.0172993f $X=1.795 $Y=2.375 $X2=0 $Y2=0
cc_305 N_A_27_74#_c_305_n N_SCE_c_383_n 0.0172641f $X=1.795 $Y=2.375 $X2=0 $Y2=0
cc_306 N_A_27_74#_c_305_n N_SCE_c_376_n 0.0126508f $X=1.795 $Y=2.375 $X2=0 $Y2=0
cc_307 N_A_27_74#_c_299_n N_SCE_c_376_n 0.0229228f $X=0.975 $Y=1.115 $X2=0 $Y2=0
cc_308 N_A_27_74#_c_300_n N_SCE_c_376_n 0.00422079f $X=0.975 $Y=1.115 $X2=0
+ $Y2=0
cc_309 N_A_27_74#_c_302_n N_SCE_c_377_n 8.97321e-19 $X=2.005 $Y=2.245 $X2=0
+ $Y2=0
cc_310 N_A_27_74#_c_299_n N_SCE_c_377_n 4.79392e-19 $X=0.975 $Y=1.115 $X2=0
+ $Y2=0
cc_311 N_A_27_74#_c_306_n N_SCE_c_377_n 0.0178307f $X=1.96 $Y=1.995 $X2=0 $Y2=0
cc_312 N_A_27_74#_c_302_n N_SCE_c_378_n 0.0192623f $X=2.005 $Y=2.245 $X2=0 $Y2=0
cc_313 N_A_27_74#_c_306_n N_SCE_c_378_n 2.95197e-19 $X=1.96 $Y=1.995 $X2=0 $Y2=0
cc_314 N_A_27_74#_c_298_n N_SCE_c_379_n 0.0246957f $X=0.225 $Y=2.29 $X2=0 $Y2=0
cc_315 N_A_27_74#_c_305_n N_SCE_c_379_n 6.8039e-19 $X=1.795 $Y=2.375 $X2=0 $Y2=0
cc_316 N_A_27_74#_c_299_n N_SCE_c_379_n 0.0014947f $X=0.975 $Y=1.115 $X2=0 $Y2=0
cc_317 N_A_27_74#_c_300_n N_SCE_c_379_n 0.00628947f $X=0.975 $Y=1.115 $X2=0
+ $Y2=0
cc_318 N_A_27_74#_c_301_n N_SCE_c_379_n 2.24402e-19 $X=0.28 $Y=1.115 $X2=0 $Y2=0
cc_319 N_A_27_74#_c_298_n N_SCE_c_380_n 0.030623f $X=0.225 $Y=2.29 $X2=0 $Y2=0
cc_320 N_A_27_74#_c_305_n N_SCE_c_380_n 0.0120121f $X=1.795 $Y=2.375 $X2=0 $Y2=0
cc_321 N_A_27_74#_c_299_n N_SCE_c_380_n 0.0272074f $X=0.975 $Y=1.115 $X2=0 $Y2=0
cc_322 N_A_27_74#_c_302_n N_D_c_453_n 0.0422336f $X=2.005 $Y=2.245 $X2=-0.19
+ $Y2=-0.245
cc_323 N_A_27_74#_c_305_n N_D_c_453_n 0.0196667f $X=1.795 $Y=2.375 $X2=-0.19
+ $Y2=-0.245
cc_324 N_A_27_74#_c_306_n N_D_c_453_n 0.00316692f $X=1.96 $Y=1.995 $X2=-0.19
+ $Y2=-0.245
cc_325 N_A_27_74#_M1036_g N_D_M1037_g 0.0528466f $X=1.065 $Y=0.58 $X2=0 $Y2=0
cc_326 N_A_27_74#_c_299_n N_D_M1037_g 0.0016481f $X=0.975 $Y=1.115 $X2=0 $Y2=0
cc_327 N_A_27_74#_c_302_n N_D_c_455_n 0.00100613f $X=2.005 $Y=2.245 $X2=0 $Y2=0
cc_328 N_A_27_74#_c_305_n N_D_c_455_n 0.0377183f $X=1.795 $Y=2.375 $X2=0 $Y2=0
cc_329 N_A_27_74#_c_306_n N_D_c_455_n 0.018611f $X=1.96 $Y=1.995 $X2=0 $Y2=0
cc_330 N_A_27_74#_c_302_n N_SCD_c_490_n 0.0419256f $X=2.005 $Y=2.245 $X2=0 $Y2=0
cc_331 N_A_27_74#_c_302_n N_SCD_c_488_n 0.0166773f $X=2.005 $Y=2.245 $X2=0 $Y2=0
cc_332 N_A_27_74#_c_306_n N_SCD_c_488_n 2.71882e-19 $X=1.96 $Y=1.995 $X2=0 $Y2=0
cc_333 N_A_27_74#_c_305_n N_VPWR_M1026_d 0.00197722f $X=1.795 $Y=2.375 $X2=-0.19
+ $Y2=-0.245
cc_334 N_A_27_74#_c_304_n N_VPWR_c_1696_n 0.0234974f $X=0.28 $Y=2.465 $X2=0
+ $Y2=0
cc_335 N_A_27_74#_c_305_n N_VPWR_c_1696_n 0.0171814f $X=1.795 $Y=2.375 $X2=0
+ $Y2=0
cc_336 N_A_27_74#_c_304_n N_VPWR_c_1711_n 0.0110674f $X=0.28 $Y=2.465 $X2=0
+ $Y2=0
cc_337 N_A_27_74#_c_302_n N_VPWR_c_1712_n 0.00312371f $X=2.005 $Y=2.245 $X2=0
+ $Y2=0
cc_338 N_A_27_74#_c_302_n N_VPWR_c_1695_n 0.0038838f $X=2.005 $Y=2.245 $X2=0
+ $Y2=0
cc_339 N_A_27_74#_c_304_n N_VPWR_c_1695_n 0.00916f $X=0.28 $Y=2.465 $X2=0 $Y2=0
cc_340 N_A_27_74#_c_305_n A_206_464# 0.00595227f $X=1.795 $Y=2.375 $X2=-0.19
+ $Y2=-0.245
cc_341 N_A_27_74#_c_305_n N_A_290_464#_M1014_d 0.00463034f $X=1.795 $Y=2.375
+ $X2=0 $Y2=0
cc_342 N_A_27_74#_c_305_n N_A_290_464#_c_1869_n 0.0230043f $X=1.795 $Y=2.375
+ $X2=0 $Y2=0
cc_343 N_A_27_74#_M1036_g N_A_290_464#_c_1856_n 0.00194947f $X=1.065 $Y=0.58
+ $X2=0 $Y2=0
cc_344 N_A_27_74#_c_299_n N_A_290_464#_c_1858_n 0.00633768f $X=0.975 $Y=1.115
+ $X2=0 $Y2=0
cc_345 N_A_27_74#_c_302_n N_A_290_464#_c_1872_n 0.00928427f $X=2.005 $Y=2.245
+ $X2=0 $Y2=0
cc_346 N_A_27_74#_c_302_n N_A_290_464#_c_1859_n 0.00313487f $X=2.005 $Y=2.245
+ $X2=0 $Y2=0
cc_347 N_A_27_74#_c_305_n N_A_290_464#_c_1859_n 0.00235958f $X=1.795 $Y=2.375
+ $X2=0 $Y2=0
cc_348 N_A_27_74#_c_306_n N_A_290_464#_c_1859_n 0.0337781f $X=1.96 $Y=1.995
+ $X2=0 $Y2=0
cc_349 N_A_27_74#_c_302_n N_A_290_464#_c_1876_n 0.00297032f $X=2.005 $Y=2.245
+ $X2=0 $Y2=0
cc_350 N_A_27_74#_c_302_n N_A_290_464#_c_1877_n 0.00951864f $X=2.005 $Y=2.245
+ $X2=0 $Y2=0
cc_351 N_A_27_74#_c_305_n N_A_290_464#_c_1877_n 0.0152871f $X=1.795 $Y=2.375
+ $X2=0 $Y2=0
cc_352 N_A_27_74#_c_302_n N_A_290_464#_c_1879_n 0.00179913f $X=2.005 $Y=2.245
+ $X2=0 $Y2=0
cc_353 N_A_27_74#_c_305_n N_A_290_464#_c_1879_n 0.0122365f $X=1.795 $Y=2.375
+ $X2=0 $Y2=0
cc_354 N_A_27_74#_M1036_g N_VGND_c_2101_n 0.00597281f $X=1.065 $Y=0.58 $X2=0
+ $Y2=0
cc_355 N_A_27_74#_c_297_n N_VGND_c_2101_n 0.0169251f $X=0.28 $Y=0.58 $X2=0 $Y2=0
cc_356 N_A_27_74#_c_299_n N_VGND_c_2101_n 0.0268964f $X=0.975 $Y=1.115 $X2=0
+ $Y2=0
cc_357 N_A_27_74#_c_300_n N_VGND_c_2101_n 0.0030881f $X=0.975 $Y=1.115 $X2=0
+ $Y2=0
cc_358 N_A_27_74#_M1036_g N_VGND_c_2107_n 0.00461464f $X=1.065 $Y=0.58 $X2=0
+ $Y2=0
cc_359 N_A_27_74#_c_297_n N_VGND_c_2111_n 0.0145639f $X=0.28 $Y=0.58 $X2=0 $Y2=0
cc_360 N_A_27_74#_M1036_g N_VGND_c_2117_n 0.00909071f $X=1.065 $Y=0.58 $X2=0
+ $Y2=0
cc_361 N_A_27_74#_c_297_n N_VGND_c_2117_n 0.0119984f $X=0.28 $Y=0.58 $X2=0 $Y2=0
cc_362 N_SCE_c_383_n N_D_c_453_n 0.0469524f $X=0.955 $Y=2.245 $X2=-0.19
+ $Y2=-0.245
cc_363 N_SCE_c_376_n N_D_c_453_n 0.00437396f $X=1.795 $Y=1.535 $X2=-0.19
+ $Y2=-0.245
cc_364 N_SCE_c_379_n N_D_c_453_n 0.0196439f $X=0.67 $Y=1.685 $X2=-0.19
+ $Y2=-0.245
cc_365 N_SCE_M1011_g N_D_M1037_g 0.0289627f $X=1.885 $Y=0.58 $X2=0 $Y2=0
cc_366 N_SCE_c_376_n N_D_M1037_g 0.0159859f $X=1.795 $Y=1.535 $X2=0 $Y2=0
cc_367 N_SCE_c_377_n N_D_M1037_g 0.00137327f $X=1.96 $Y=1.425 $X2=0 $Y2=0
cc_368 N_SCE_c_378_n N_D_M1037_g 0.0163018f $X=1.96 $Y=1.425 $X2=0 $Y2=0
cc_369 N_SCE_c_379_n N_D_M1037_g 0.00756384f $X=0.67 $Y=1.685 $X2=0 $Y2=0
cc_370 N_SCE_c_380_n N_D_M1037_g 9.94783e-19 $X=0.67 $Y=1.535 $X2=0 $Y2=0
cc_371 N_SCE_c_376_n N_D_c_455_n 0.0377186f $X=1.795 $Y=1.535 $X2=0 $Y2=0
cc_372 N_SCE_c_379_n N_D_c_455_n 0.0083863f $X=0.67 $Y=1.685 $X2=0 $Y2=0
cc_373 N_SCE_c_380_n N_D_c_455_n 0.00363459f $X=0.67 $Y=1.535 $X2=0 $Y2=0
cc_374 N_SCE_M1011_g N_SCD_c_486_n 0.0397201f $X=1.885 $Y=0.58 $X2=-0.19
+ $Y2=-0.245
cc_375 N_SCE_M1011_g N_SCD_c_487_n 0.00623104f $X=1.885 $Y=0.58 $X2=0 $Y2=0
cc_376 N_SCE_c_377_n N_SCD_c_487_n 2.80393e-19 $X=1.96 $Y=1.425 $X2=0 $Y2=0
cc_377 N_SCE_c_378_n N_SCD_c_487_n 0.0171993f $X=1.96 $Y=1.425 $X2=0 $Y2=0
cc_378 N_SCE_c_382_n N_VPWR_c_1696_n 0.0104494f $X=0.505 $Y=2.245 $X2=0 $Y2=0
cc_379 N_SCE_c_383_n N_VPWR_c_1696_n 0.00994646f $X=0.955 $Y=2.245 $X2=0 $Y2=0
cc_380 N_SCE_c_382_n N_VPWR_c_1711_n 0.00413917f $X=0.505 $Y=2.245 $X2=0 $Y2=0
cc_381 N_SCE_c_383_n N_VPWR_c_1712_n 0.00413917f $X=0.955 $Y=2.245 $X2=0 $Y2=0
cc_382 N_SCE_c_382_n N_VPWR_c_1695_n 0.00821221f $X=0.505 $Y=2.245 $X2=0 $Y2=0
cc_383 N_SCE_c_383_n N_VPWR_c_1695_n 0.00817532f $X=0.955 $Y=2.245 $X2=0 $Y2=0
cc_384 N_SCE_c_383_n N_A_290_464#_c_1869_n 9.43907e-19 $X=0.955 $Y=2.245 $X2=0
+ $Y2=0
cc_385 N_SCE_M1011_g N_A_290_464#_c_1856_n 0.0119647f $X=1.885 $Y=0.58 $X2=0
+ $Y2=0
cc_386 N_SCE_M1011_g N_A_290_464#_c_1857_n 0.0112369f $X=1.885 $Y=0.58 $X2=0
+ $Y2=0
cc_387 N_SCE_c_377_n N_A_290_464#_c_1857_n 0.0153887f $X=1.96 $Y=1.425 $X2=0
+ $Y2=0
cc_388 N_SCE_c_378_n N_A_290_464#_c_1857_n 0.00363502f $X=1.96 $Y=1.425 $X2=0
+ $Y2=0
cc_389 N_SCE_M1011_g N_A_290_464#_c_1858_n 0.00274486f $X=1.885 $Y=0.58 $X2=0
+ $Y2=0
cc_390 N_SCE_c_376_n N_A_290_464#_c_1858_n 0.0143345f $X=1.795 $Y=1.535 $X2=0
+ $Y2=0
cc_391 N_SCE_c_377_n N_A_290_464#_c_1858_n 0.00321217f $X=1.96 $Y=1.425 $X2=0
+ $Y2=0
cc_392 N_SCE_M1011_g N_A_290_464#_c_1859_n 0.00333921f $X=1.885 $Y=0.58 $X2=0
+ $Y2=0
cc_393 N_SCE_c_377_n N_A_290_464#_c_1859_n 0.0266104f $X=1.96 $Y=1.425 $X2=0
+ $Y2=0
cc_394 N_SCE_c_378_n N_A_290_464#_c_1859_n 0.00220024f $X=1.96 $Y=1.425 $X2=0
+ $Y2=0
cc_395 N_SCE_M1033_g N_VGND_c_2101_n 0.00586161f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_396 N_SCE_M1011_g N_VGND_c_2102_n 0.00169331f $X=1.885 $Y=0.58 $X2=0 $Y2=0
cc_397 N_SCE_M1011_g N_VGND_c_2107_n 0.00434272f $X=1.885 $Y=0.58 $X2=0 $Y2=0
cc_398 N_SCE_M1033_g N_VGND_c_2111_n 0.00434272f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_399 N_SCE_M1033_g N_VGND_c_2117_n 0.0082497f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_400 N_SCE_M1011_g N_VGND_c_2117_n 0.00821077f $X=1.885 $Y=0.58 $X2=0 $Y2=0
cc_401 N_D_c_453_n N_VPWR_c_1696_n 0.00159466f $X=1.375 $Y=2.245 $X2=0 $Y2=0
cc_402 N_D_c_453_n N_VPWR_c_1712_n 0.00444752f $X=1.375 $Y=2.245 $X2=0 $Y2=0
cc_403 N_D_c_453_n N_VPWR_c_1695_n 0.00856194f $X=1.375 $Y=2.245 $X2=0 $Y2=0
cc_404 N_D_c_453_n N_A_290_464#_c_1869_n 0.0115882f $X=1.375 $Y=2.245 $X2=0
+ $Y2=0
cc_405 N_D_M1037_g N_A_290_464#_c_1856_n 0.0124194f $X=1.455 $Y=0.58 $X2=0 $Y2=0
cc_406 N_D_M1037_g N_A_290_464#_c_1858_n 0.00512834f $X=1.455 $Y=0.58 $X2=0
+ $Y2=0
cc_407 N_D_M1037_g N_A_290_464#_c_1859_n 0.00342727f $X=1.455 $Y=0.58 $X2=0
+ $Y2=0
cc_408 N_D_c_455_n N_A_290_464#_c_1859_n 0.00111607f $X=1.42 $Y=1.955 $X2=0
+ $Y2=0
cc_409 N_D_M1037_g N_VGND_c_2107_n 0.00434272f $X=1.455 $Y=0.58 $X2=0 $Y2=0
cc_410 N_D_M1037_g N_VGND_c_2117_n 0.00821077f $X=1.455 $Y=0.58 $X2=0 $Y2=0
cc_411 N_SCD_c_487_n N_CLK_c_529_n 0.00165831f $X=2.597 $Y=1.372 $X2=-0.19
+ $Y2=-0.245
cc_412 N_SCD_c_487_n N_CLK_c_530_n 0.00841032f $X=2.597 $Y=1.372 $X2=0 $Y2=0
cc_413 N_SCD_c_488_n N_CLK_c_530_n 0.00583564f $X=2.597 $Y=1.918 $X2=0 $Y2=0
cc_414 N_SCD_c_486_n N_A_594_74#_c_1148_n 0.00350312f $X=2.275 $Y=0.865 $X2=0
+ $Y2=0
cc_415 N_SCD_c_487_n N_A_594_74#_c_1148_n 0.00561892f $X=2.597 $Y=1.372 $X2=0
+ $Y2=0
cc_416 N_SCD_c_487_n N_A_594_74#_c_1149_n 0.00682259f $X=2.597 $Y=1.372 $X2=0
+ $Y2=0
cc_417 SCD N_A_594_74#_c_1149_n 0.0493209f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_418 N_SCD_c_488_n N_A_594_74#_c_1163_n 0.0042094f $X=2.597 $Y=1.918 $X2=0
+ $Y2=0
cc_419 SCD N_A_594_74#_c_1163_n 0.0266661f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_420 N_SCD_c_490_n N_VPWR_c_1697_n 0.00526487f $X=2.425 $Y=2.245 $X2=0 $Y2=0
cc_421 N_SCD_c_490_n N_VPWR_c_1712_n 0.00427116f $X=2.425 $Y=2.245 $X2=0 $Y2=0
cc_422 N_SCD_c_490_n N_VPWR_c_1695_n 0.0045104f $X=2.425 $Y=2.245 $X2=0 $Y2=0
cc_423 N_SCD_c_486_n N_A_290_464#_c_1856_n 0.00199036f $X=2.275 $Y=0.865 $X2=0
+ $Y2=0
cc_424 N_SCD_c_487_n N_A_290_464#_c_1857_n 0.017869f $X=2.597 $Y=1.372 $X2=0
+ $Y2=0
cc_425 N_SCD_c_490_n N_A_290_464#_c_1872_n 0.00557018f $X=2.425 $Y=2.245 $X2=0
+ $Y2=0
cc_426 N_SCD_c_490_n N_A_290_464#_c_1859_n 0.013491f $X=2.425 $Y=2.245 $X2=0
+ $Y2=0
cc_427 N_SCD_c_487_n N_A_290_464#_c_1859_n 0.00695808f $X=2.597 $Y=1.372 $X2=0
+ $Y2=0
cc_428 N_SCD_c_488_n N_A_290_464#_c_1859_n 0.0145162f $X=2.597 $Y=1.918 $X2=0
+ $Y2=0
cc_429 SCD N_A_290_464#_c_1859_n 0.0694511f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_430 N_SCD_c_490_n N_A_290_464#_c_1876_n 0.00661899f $X=2.425 $Y=2.245 $X2=0
+ $Y2=0
cc_431 N_SCD_c_490_n N_A_290_464#_c_1863_n 0.01771f $X=2.425 $Y=2.245 $X2=0
+ $Y2=0
cc_432 SCD N_A_290_464#_c_1863_n 0.0163122f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_433 N_SCD_c_490_n N_A_290_464#_c_1877_n 4.71381e-19 $X=2.425 $Y=2.245 $X2=0
+ $Y2=0
cc_434 N_SCD_c_490_n N_A_290_464#_c_1879_n 0.00171789f $X=2.425 $Y=2.245 $X2=0
+ $Y2=0
cc_435 N_SCD_c_486_n N_VGND_c_2102_n 0.0121542f $X=2.275 $Y=0.865 $X2=0 $Y2=0
cc_436 N_SCD_c_487_n N_VGND_c_2102_n 0.00915488f $X=2.597 $Y=1.372 $X2=0 $Y2=0
cc_437 SCD N_VGND_c_2102_n 0.00453686f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_438 N_SCD_c_486_n N_VGND_c_2107_n 0.00383152f $X=2.275 $Y=0.865 $X2=0 $Y2=0
cc_439 N_SCD_c_486_n N_VGND_c_2117_n 0.0075725f $X=2.275 $Y=0.865 $X2=0 $Y2=0
cc_440 N_CLK_c_529_n N_A_594_74#_c_1139_n 0.0188174f $X=3.33 $Y=1.22 $X2=0 $Y2=0
cc_441 CLK N_A_594_74#_c_1139_n 0.0024284f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_442 N_CLK_c_530_n N_A_594_74#_c_1140_n 0.0650275f $X=3.515 $Y=1.765 $X2=0
+ $Y2=0
cc_443 CLK N_A_594_74#_c_1140_n 0.00149275f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_444 N_CLK_c_529_n N_A_594_74#_c_1148_n 6.68688e-19 $X=3.33 $Y=1.22 $X2=0
+ $Y2=0
cc_445 N_CLK_c_529_n N_A_594_74#_c_1149_n 0.00522155f $X=3.33 $Y=1.22 $X2=0
+ $Y2=0
cc_446 N_CLK_c_530_n N_A_594_74#_c_1149_n 0.00821742f $X=3.515 $Y=1.765 $X2=0
+ $Y2=0
cc_447 CLK N_A_594_74#_c_1149_n 0.028374f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_448 N_CLK_c_530_n N_A_594_74#_c_1164_n 0.00932924f $X=3.515 $Y=1.765 $X2=0
+ $Y2=0
cc_449 N_CLK_c_530_n N_A_594_74#_c_1150_n 0.00274031f $X=3.515 $Y=1.765 $X2=0
+ $Y2=0
cc_450 CLK N_A_594_74#_c_1150_n 0.0267715f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_451 N_CLK_c_530_n N_A_594_74#_c_1166_n 0.00523766f $X=3.515 $Y=1.765 $X2=0
+ $Y2=0
cc_452 CLK N_A_594_74#_c_1166_n 0.0242245f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_453 N_CLK_c_530_n N_A_594_74#_c_1167_n 0.00540192f $X=3.515 $Y=1.765 $X2=0
+ $Y2=0
cc_454 N_CLK_c_530_n N_VPWR_c_1697_n 0.00969005f $X=3.515 $Y=1.765 $X2=0 $Y2=0
cc_455 N_CLK_c_530_n N_VPWR_c_1698_n 0.00413917f $X=3.515 $Y=1.765 $X2=0 $Y2=0
cc_456 N_CLK_c_530_n N_VPWR_c_1699_n 0.0202592f $X=3.515 $Y=1.765 $X2=0 $Y2=0
cc_457 N_CLK_c_530_n N_VPWR_c_1695_n 0.00419307f $X=3.515 $Y=1.765 $X2=0 $Y2=0
cc_458 N_CLK_c_530_n N_A_290_464#_c_1863_n 0.0133694f $X=3.515 $Y=1.765 $X2=0
+ $Y2=0
cc_459 N_CLK_c_529_n N_VGND_c_2102_n 0.00308778f $X=3.33 $Y=1.22 $X2=0 $Y2=0
cc_460 N_CLK_c_529_n N_VGND_c_2103_n 0.0139212f $X=3.33 $Y=1.22 $X2=0 $Y2=0
cc_461 N_CLK_c_530_n N_VGND_c_2103_n 8.2516e-19 $X=3.515 $Y=1.765 $X2=0 $Y2=0
cc_462 CLK N_VGND_c_2103_n 0.0254134f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_463 N_CLK_c_529_n N_VGND_c_2112_n 0.00383152f $X=3.33 $Y=1.22 $X2=0 $Y2=0
cc_464 N_CLK_c_529_n N_VGND_c_2117_n 0.00762539f $X=3.33 $Y=1.22 $X2=0 $Y2=0
cc_465 N_A_781_74#_M1004_g N_A_1163_48#_c_771_n 0.0511043f $X=5.5 $Y=0.58 $X2=0
+ $Y2=0
cc_466 N_A_781_74#_c_577_n N_A_1163_48#_c_772_n 0.00125914f $X=5.725 $Y=2.255
+ $X2=0 $Y2=0
cc_467 N_A_781_74#_c_579_n N_A_1163_48#_c_772_n 0.00428061f $X=6.595 $Y=2.17
+ $X2=0 $Y2=0
cc_468 N_A_781_74#_c_587_n N_A_1163_48#_c_772_n 0.0197055f $X=5.645 $Y=1.855
+ $X2=0 $Y2=0
cc_469 N_A_781_74#_c_577_n N_A_1163_48#_c_777_n 0.0021815f $X=5.725 $Y=2.255
+ $X2=0 $Y2=0
cc_470 N_A_781_74#_c_579_n N_A_1163_48#_c_777_n 0.00620623f $X=6.595 $Y=2.17
+ $X2=0 $Y2=0
cc_471 N_A_781_74#_c_578_n N_A_1163_48#_c_778_n 0.00688986f $X=5.725 $Y=2.905
+ $X2=0 $Y2=0
cc_472 N_A_781_74#_c_579_n N_A_1163_48#_c_778_n 0.0122739f $X=6.595 $Y=2.17
+ $X2=0 $Y2=0
cc_473 N_A_781_74#_c_580_n N_A_1163_48#_c_778_n 0.00352077f $X=6.68 $Y=2.905
+ $X2=0 $Y2=0
cc_474 N_A_781_74#_M1004_g N_A_1163_48#_c_773_n 0.0114125f $X=5.5 $Y=0.58 $X2=0
+ $Y2=0
cc_475 N_A_781_74#_M1004_g N_A_1163_48#_c_774_n 0.00153185f $X=5.5 $Y=0.58 $X2=0
+ $Y2=0
cc_476 N_A_781_74#_c_577_n N_A_1163_48#_c_779_n 0.0133533f $X=5.725 $Y=2.255
+ $X2=0 $Y2=0
cc_477 N_A_781_74#_c_579_n N_A_1163_48#_c_779_n 0.0541693f $X=6.595 $Y=2.17
+ $X2=0 $Y2=0
cc_478 N_A_781_74#_c_587_n N_A_1163_48#_c_779_n 2.73581e-19 $X=5.645 $Y=1.855
+ $X2=0 $Y2=0
cc_479 N_A_781_74#_c_579_n N_A_1163_48#_c_780_n 0.0134997f $X=6.595 $Y=2.17
+ $X2=0 $Y2=0
cc_480 N_A_781_74#_c_580_n N_A_1163_48#_c_780_n 0.0337427f $X=6.68 $Y=2.905
+ $X2=0 $Y2=0
cc_481 N_A_781_74#_c_581_n N_A_1163_48#_c_780_n 0.0130106f $X=7.275 $Y=2.99
+ $X2=0 $Y2=0
cc_482 N_A_781_74#_c_583_n N_A_1163_48#_c_780_n 0.0298578f $X=7.36 $Y=2.905
+ $X2=0 $Y2=0
cc_483 N_A_781_74#_c_585_n N_A_1163_48#_c_780_n 0.0143554f $X=7.445 $Y=2.035
+ $X2=0 $Y2=0
cc_484 N_A_781_74#_c_579_n N_A_995_74#_c_847_n 0.00287465f $X=6.595 $Y=2.17
+ $X2=0 $Y2=0
cc_485 N_A_781_74#_c_579_n N_A_995_74#_c_859_n 0.00361736f $X=6.595 $Y=2.17
+ $X2=0 $Y2=0
cc_486 N_A_781_74#_c_580_n N_A_995_74#_c_859_n 0.0155004f $X=6.68 $Y=2.905 $X2=0
+ $Y2=0
cc_487 N_A_781_74#_c_581_n N_A_995_74#_c_859_n 0.00295621f $X=7.275 $Y=2.99
+ $X2=0 $Y2=0
cc_488 N_A_781_74#_c_583_n N_A_995_74#_c_859_n 0.00101154f $X=7.36 $Y=2.905
+ $X2=0 $Y2=0
cc_489 N_A_781_74#_c_583_n N_A_995_74#_c_860_n 0.0011264f $X=7.36 $Y=2.905 $X2=0
+ $Y2=0
cc_490 N_A_781_74#_c_584_n N_A_995_74#_c_860_n 0.0184984f $X=8.66 $Y=2.035 $X2=0
+ $Y2=0
cc_491 N_A_781_74#_c_586_n N_A_995_74#_c_860_n 0.00319069f $X=8.745 $Y=1.95
+ $X2=0 $Y2=0
cc_492 N_A_781_74#_c_569_n N_A_995_74#_c_860_n 6.95987e-19 $X=8.825 $Y=1.515
+ $X2=0 $Y2=0
cc_493 N_A_781_74#_c_570_n N_A_995_74#_c_860_n 0.00243027f $X=8.825 $Y=1.515
+ $X2=0 $Y2=0
cc_494 N_A_781_74#_M1024_g N_A_995_74#_c_849_n 0.0322153f $X=8.735 $Y=0.69 $X2=0
+ $Y2=0
cc_495 N_A_781_74#_M1004_g N_A_995_74#_c_850_n 0.0256791f $X=5.5 $Y=0.58 $X2=0
+ $Y2=0
cc_496 N_A_781_74#_c_565_n N_A_995_74#_c_850_n 0.00381334f $X=4.86 $Y=0.34 $X2=0
+ $Y2=0
cc_497 N_A_781_74#_c_568_n N_A_995_74#_c_850_n 0.0574008f $X=4.895 $Y=1.37 $X2=0
+ $Y2=0
cc_498 N_A_781_74#_c_561_n N_A_995_74#_c_851_n 0.00961157f $X=4.985 $Y=2.24
+ $X2=0 $Y2=0
cc_499 N_A_781_74#_M1004_g N_A_995_74#_c_851_n 0.00415339f $X=5.5 $Y=0.58 $X2=0
+ $Y2=0
cc_500 N_A_781_74#_c_576_n N_A_995_74#_c_851_n 0.0378893f $X=4.925 $Y=1.535
+ $X2=0 $Y2=0
cc_501 N_A_781_74#_c_577_n N_A_995_74#_c_851_n 0.03794f $X=5.725 $Y=2.255 $X2=0
+ $Y2=0
cc_502 N_A_781_74#_c_578_n N_A_995_74#_c_851_n 0.00571525f $X=5.725 $Y=2.905
+ $X2=0 $Y2=0
cc_503 N_A_781_74#_c_587_n N_A_995_74#_c_851_n 0.00159541f $X=5.645 $Y=1.855
+ $X2=0 $Y2=0
cc_504 N_A_781_74#_c_589_n N_A_995_74#_c_851_n 0.0136656f $X=5.425 $Y=1.855
+ $X2=0 $Y2=0
cc_505 N_A_781_74#_M1004_g N_A_995_74#_c_852_n 0.014507f $X=5.5 $Y=0.58 $X2=0
+ $Y2=0
cc_506 N_A_781_74#_c_577_n N_A_995_74#_c_852_n 0.0210075f $X=5.725 $Y=2.255
+ $X2=0 $Y2=0
cc_507 N_A_781_74#_c_579_n N_A_995_74#_c_852_n 0.00772262f $X=6.595 $Y=2.17
+ $X2=0 $Y2=0
cc_508 N_A_781_74#_c_587_n N_A_995_74#_c_852_n 0.00165663f $X=5.645 $Y=1.855
+ $X2=0 $Y2=0
cc_509 N_A_781_74#_M1024_g N_A_995_74#_c_854_n 0.00114708f $X=8.735 $Y=0.69
+ $X2=0 $Y2=0
cc_510 N_A_781_74#_c_584_n N_A_995_74#_c_854_n 0.00410725f $X=8.66 $Y=2.035
+ $X2=0 $Y2=0
cc_511 N_A_781_74#_c_569_n N_A_995_74#_c_854_n 0.00313951f $X=8.825 $Y=1.515
+ $X2=0 $Y2=0
cc_512 N_A_781_74#_c_584_n N_A_995_74#_c_855_n 0.00789988f $X=8.66 $Y=2.035
+ $X2=0 $Y2=0
cc_513 N_A_781_74#_c_569_n N_A_995_74#_c_855_n 0.00156549f $X=8.825 $Y=1.515
+ $X2=0 $Y2=0
cc_514 N_A_781_74#_c_570_n N_A_995_74#_c_855_n 0.03631f $X=8.825 $Y=1.515 $X2=0
+ $Y2=0
cc_515 N_A_781_74#_c_561_n N_A_995_74#_c_863_n 0.0036212f $X=4.985 $Y=2.24 $X2=0
+ $Y2=0
cc_516 N_A_781_74#_c_574_n N_A_995_74#_c_863_n 0.0248496f $X=5.64 $Y=2.99 $X2=0
+ $Y2=0
cc_517 N_A_781_74#_c_578_n N_A_995_74#_c_863_n 0.0248233f $X=5.725 $Y=2.905
+ $X2=0 $Y2=0
cc_518 N_A_781_74#_c_587_n N_A_995_74#_c_863_n 8.90055e-19 $X=5.645 $Y=1.855
+ $X2=0 $Y2=0
cc_519 N_A_781_74#_c_589_n N_A_995_74#_c_863_n 0.00401388f $X=5.425 $Y=1.855
+ $X2=0 $Y2=0
cc_520 N_A_781_74#_c_561_n N_A_995_74#_c_856_n 0.00130826f $X=4.985 $Y=2.24
+ $X2=0 $Y2=0
cc_521 N_A_781_74#_M1004_g N_A_995_74#_c_856_n 0.00354176f $X=5.5 $Y=0.58 $X2=0
+ $Y2=0
cc_522 N_A_781_74#_c_568_n N_A_995_74#_c_856_n 0.0140925f $X=4.895 $Y=1.37 $X2=0
+ $Y2=0
cc_523 N_A_781_74#_c_583_n N_SET_B_c_984_n 9.69591e-19 $X=7.36 $Y=2.905 $X2=0
+ $Y2=0
cc_524 N_A_781_74#_c_584_n N_SET_B_c_984_n 0.00449499f $X=8.66 $Y=2.035 $X2=0
+ $Y2=0
cc_525 N_A_781_74#_c_585_n N_SET_B_c_984_n 0.00552929f $X=7.445 $Y=2.035 $X2=0
+ $Y2=0
cc_526 N_A_781_74#_c_580_n N_SET_B_c_999_n 2.30666e-19 $X=6.68 $Y=2.905 $X2=0
+ $Y2=0
cc_527 N_A_781_74#_c_583_n N_SET_B_c_999_n 0.0206842f $X=7.36 $Y=2.905 $X2=0
+ $Y2=0
cc_528 N_A_781_74#_c_584_n N_SET_B_c_992_n 0.0395273f $X=8.66 $Y=2.035 $X2=0
+ $Y2=0
cc_529 N_A_781_74#_c_586_n N_SET_B_c_992_n 0.00672398f $X=8.745 $Y=1.95 $X2=0
+ $Y2=0
cc_530 N_A_781_74#_c_569_n N_SET_B_c_992_n 0.0177158f $X=8.825 $Y=1.515 $X2=0
+ $Y2=0
cc_531 N_A_781_74#_c_570_n N_SET_B_c_992_n 0.00477276f $X=8.825 $Y=1.515 $X2=0
+ $Y2=0
cc_532 N_A_781_74#_c_584_n N_SET_B_c_993_n 0.00105565f $X=8.66 $Y=2.035 $X2=0
+ $Y2=0
cc_533 N_A_781_74#_c_585_n N_SET_B_c_993_n 0.00120115f $X=7.445 $Y=2.035 $X2=0
+ $Y2=0
cc_534 N_A_781_74#_c_584_n N_SET_B_c_995_n 6.49836e-19 $X=8.66 $Y=2.035 $X2=0
+ $Y2=0
cc_535 N_A_781_74#_c_584_n N_SET_B_c_996_n 0.0120873f $X=8.66 $Y=2.035 $X2=0
+ $Y2=0
cc_536 N_A_781_74#_c_585_n N_SET_B_c_996_n 0.0100795f $X=7.445 $Y=2.035 $X2=0
+ $Y2=0
cc_537 N_A_781_74#_c_564_n N_A_594_74#_c_1139_n 0.00651805f $X=4.045 $Y=0.505
+ $X2=0 $Y2=0
cc_538 N_A_781_74#_c_566_n N_A_594_74#_c_1139_n 0.00462516f $X=4.21 $Y=0.34
+ $X2=0 $Y2=0
cc_539 N_A_781_74#_c_564_n N_A_594_74#_c_1140_n 0.00163342f $X=4.045 $Y=0.505
+ $X2=0 $Y2=0
cc_540 N_A_781_74#_c_573_n N_A_594_74#_c_1140_n 0.00328099f $X=4.19 $Y=2.765
+ $X2=0 $Y2=0
cc_541 N_A_781_74#_c_575_n N_A_594_74#_c_1140_n 0.00133627f $X=4.355 $Y=2.99
+ $X2=0 $Y2=0
cc_542 N_A_781_74#_c_561_n N_A_594_74#_c_1142_n 0.0193082f $X=4.985 $Y=2.24
+ $X2=0 $Y2=0
cc_543 N_A_781_74#_c_573_n N_A_594_74#_c_1142_n 0.00633501f $X=4.19 $Y=2.765
+ $X2=0 $Y2=0
cc_544 N_A_781_74#_c_574_n N_A_594_74#_c_1142_n 0.0113792f $X=5.64 $Y=2.99 $X2=0
+ $Y2=0
cc_545 N_A_781_74#_c_576_n N_A_594_74#_c_1142_n 3.88824e-19 $X=4.925 $Y=1.535
+ $X2=0 $Y2=0
cc_546 N_A_781_74#_c_561_n N_A_594_74#_c_1143_n 0.0116591f $X=4.985 $Y=2.24
+ $X2=0 $Y2=0
cc_547 N_A_781_74#_c_565_n N_A_594_74#_c_1143_n 0.00253049f $X=4.86 $Y=0.34
+ $X2=0 $Y2=0
cc_548 N_A_781_74#_c_567_n N_A_594_74#_c_1143_n 6.71829e-19 $X=4.895 $Y=1.505
+ $X2=0 $Y2=0
cc_549 N_A_781_74#_c_568_n N_A_594_74#_c_1143_n 0.00664279f $X=4.895 $Y=1.37
+ $X2=0 $Y2=0
cc_550 N_A_781_74#_c_561_n N_A_594_74#_c_1154_n 0.00882199f $X=4.985 $Y=2.24
+ $X2=0 $Y2=0
cc_551 N_A_781_74#_c_574_n N_A_594_74#_c_1154_n 0.0155776f $X=5.64 $Y=2.99 $X2=0
+ $Y2=0
cc_552 N_A_781_74#_M1004_g N_A_594_74#_M1034_g 0.0160063f $X=5.5 $Y=0.58 $X2=0
+ $Y2=0
cc_553 N_A_781_74#_c_564_n N_A_594_74#_M1034_g 0.00301996f $X=4.045 $Y=0.505
+ $X2=0 $Y2=0
cc_554 N_A_781_74#_c_565_n N_A_594_74#_M1034_g 0.010044f $X=4.86 $Y=0.34 $X2=0
+ $Y2=0
cc_555 N_A_781_74#_c_568_n N_A_594_74#_M1034_g 0.0157578f $X=4.895 $Y=1.37 $X2=0
+ $Y2=0
cc_556 N_A_781_74#_c_561_n N_A_594_74#_c_1156_n 0.0116164f $X=4.985 $Y=2.24
+ $X2=0 $Y2=0
cc_557 N_A_781_74#_c_577_n N_A_594_74#_c_1156_n 7.58855e-19 $X=5.725 $Y=2.255
+ $X2=0 $Y2=0
cc_558 N_A_781_74#_c_578_n N_A_594_74#_c_1156_n 0.0148561f $X=5.725 $Y=2.905
+ $X2=0 $Y2=0
cc_559 N_A_781_74#_c_587_n N_A_594_74#_c_1156_n 0.00891023f $X=5.645 $Y=1.855
+ $X2=0 $Y2=0
cc_560 N_A_781_74#_c_574_n N_A_594_74#_c_1157_n 0.00318937f $X=5.64 $Y=2.99
+ $X2=0 $Y2=0
cc_561 N_A_781_74#_c_581_n N_A_594_74#_c_1157_n 0.0121639f $X=7.275 $Y=2.99
+ $X2=0 $Y2=0
cc_562 N_A_781_74#_c_582_n N_A_594_74#_c_1157_n 0.00345098f $X=6.765 $Y=2.99
+ $X2=0 $Y2=0
cc_563 N_A_781_74#_c_590_n N_A_594_74#_c_1157_n 0.00157177f $X=8.825 $Y=1.795
+ $X2=0 $Y2=0
cc_564 N_A_781_74#_M1024_g N_A_594_74#_M1000_g 0.0205499f $X=8.735 $Y=0.69 $X2=0
+ $Y2=0
cc_565 N_A_781_74#_c_569_n N_A_594_74#_M1000_g 4.68509e-19 $X=8.825 $Y=1.515
+ $X2=0 $Y2=0
cc_566 N_A_781_74#_c_570_n N_A_594_74#_M1000_g 0.0242476f $X=8.825 $Y=1.515
+ $X2=0 $Y2=0
cc_567 N_A_781_74#_c_590_n N_A_594_74#_M1009_g 0.0131594f $X=8.825 $Y=1.795
+ $X2=0 $Y2=0
cc_568 N_A_781_74#_c_561_n N_A_594_74#_c_1146_n 0.0423314f $X=4.985 $Y=2.24
+ $X2=0 $Y2=0
cc_569 N_A_781_74#_c_564_n N_A_594_74#_c_1146_n 3.03407e-19 $X=4.045 $Y=0.505
+ $X2=0 $Y2=0
cc_570 N_A_781_74#_c_565_n N_A_594_74#_c_1146_n 5.72887e-19 $X=4.86 $Y=0.34
+ $X2=0 $Y2=0
cc_571 N_A_781_74#_c_567_n N_A_594_74#_c_1146_n 3.88824e-19 $X=4.895 $Y=1.505
+ $X2=0 $Y2=0
cc_572 N_A_781_74#_c_568_n N_A_594_74#_c_1146_n 8.69379e-19 $X=4.895 $Y=1.37
+ $X2=0 $Y2=0
cc_573 N_A_781_74#_c_574_n N_A_594_74#_c_1159_n 0.0171659f $X=5.64 $Y=2.99 $X2=0
+ $Y2=0
cc_574 N_A_781_74#_c_578_n N_A_594_74#_c_1159_n 0.00148788f $X=5.725 $Y=2.905
+ $X2=0 $Y2=0
cc_575 N_A_781_74#_M1029_d N_A_594_74#_c_1164_n 0.00287936f $X=4.04 $Y=1.84
+ $X2=0 $Y2=0
cc_576 N_A_781_74#_c_564_n N_A_594_74#_c_1150_n 0.0216703f $X=4.045 $Y=0.505
+ $X2=0 $Y2=0
cc_577 N_A_781_74#_M1024_g N_A_1762_74#_c_1468_n 0.0185265f $X=8.735 $Y=0.69
+ $X2=0 $Y2=0
cc_578 N_A_781_74#_c_569_n N_A_1762_74#_c_1468_n 0.0100316f $X=8.825 $Y=1.515
+ $X2=0 $Y2=0
cc_579 N_A_781_74#_c_570_n N_A_1762_74#_c_1468_n 0.00130602f $X=8.825 $Y=1.515
+ $X2=0 $Y2=0
cc_580 N_A_781_74#_c_584_n N_A_1762_74#_c_1484_n 0.0116914f $X=8.66 $Y=2.035
+ $X2=0 $Y2=0
cc_581 N_A_781_74#_c_586_n N_A_1762_74#_c_1484_n 0.00619036f $X=8.745 $Y=1.95
+ $X2=0 $Y2=0
cc_582 N_A_781_74#_c_590_n N_A_1762_74#_c_1484_n 0.00419688f $X=8.825 $Y=1.795
+ $X2=0 $Y2=0
cc_583 N_A_781_74#_M1024_g N_A_1762_74#_c_1469_n 0.0041777f $X=8.735 $Y=0.69
+ $X2=0 $Y2=0
cc_584 N_A_781_74#_c_586_n N_A_1762_74#_c_1469_n 0.00405581f $X=8.745 $Y=1.95
+ $X2=0 $Y2=0
cc_585 N_A_781_74#_c_569_n N_A_1762_74#_c_1469_n 0.0195875f $X=8.825 $Y=1.515
+ $X2=0 $Y2=0
cc_586 N_A_781_74#_c_570_n N_A_1762_74#_c_1469_n 0.00247272f $X=8.825 $Y=1.515
+ $X2=0 $Y2=0
cc_587 N_A_781_74#_c_580_n N_VPWR_M1025_d 0.00440946f $X=6.68 $Y=2.905 $X2=0
+ $Y2=0
cc_588 N_A_781_74#_c_584_n N_VPWR_M1013_d 0.00609056f $X=8.66 $Y=2.035 $X2=0
+ $Y2=0
cc_589 N_A_781_74#_c_573_n N_VPWR_c_1699_n 0.0163934f $X=4.19 $Y=2.765 $X2=0
+ $Y2=0
cc_590 N_A_781_74#_c_575_n N_VPWR_c_1699_n 0.0125885f $X=4.355 $Y=2.99 $X2=0
+ $Y2=0
cc_591 N_A_781_74#_c_574_n N_VPWR_c_1700_n 0.00867486f $X=5.64 $Y=2.99 $X2=0
+ $Y2=0
cc_592 N_A_781_74#_c_578_n N_VPWR_c_1700_n 0.0195584f $X=5.725 $Y=2.905 $X2=0
+ $Y2=0
cc_593 N_A_781_74#_c_579_n N_VPWR_c_1700_n 0.017848f $X=6.595 $Y=2.17 $X2=0
+ $Y2=0
cc_594 N_A_781_74#_c_580_n N_VPWR_c_1700_n 0.0363341f $X=6.68 $Y=2.905 $X2=0
+ $Y2=0
cc_595 N_A_781_74#_c_582_n N_VPWR_c_1700_n 0.0147459f $X=6.765 $Y=2.99 $X2=0
+ $Y2=0
cc_596 N_A_781_74#_c_581_n N_VPWR_c_1701_n 0.0143583f $X=7.275 $Y=2.99 $X2=0
+ $Y2=0
cc_597 N_A_781_74#_c_583_n N_VPWR_c_1701_n 0.0431626f $X=7.36 $Y=2.905 $X2=0
+ $Y2=0
cc_598 N_A_781_74#_c_584_n N_VPWR_c_1701_n 0.0129262f $X=8.66 $Y=2.035 $X2=0
+ $Y2=0
cc_599 N_A_781_74#_c_574_n N_VPWR_c_1705_n 0.0933852f $X=5.64 $Y=2.99 $X2=0
+ $Y2=0
cc_600 N_A_781_74#_c_575_n N_VPWR_c_1705_n 0.0175791f $X=4.355 $Y=2.99 $X2=0
+ $Y2=0
cc_601 N_A_781_74#_c_581_n N_VPWR_c_1707_n 0.0443733f $X=7.275 $Y=2.99 $X2=0
+ $Y2=0
cc_602 N_A_781_74#_c_582_n N_VPWR_c_1707_n 0.0115893f $X=6.765 $Y=2.99 $X2=0
+ $Y2=0
cc_603 N_A_781_74#_c_574_n N_VPWR_c_1695_n 0.0489337f $X=5.64 $Y=2.99 $X2=0
+ $Y2=0
cc_604 N_A_781_74#_c_575_n N_VPWR_c_1695_n 0.00965514f $X=4.355 $Y=2.99 $X2=0
+ $Y2=0
cc_605 N_A_781_74#_c_581_n N_VPWR_c_1695_n 0.0229659f $X=7.275 $Y=2.99 $X2=0
+ $Y2=0
cc_606 N_A_781_74#_c_582_n N_VPWR_c_1695_n 0.00583135f $X=6.765 $Y=2.99 $X2=0
+ $Y2=0
cc_607 N_A_781_74#_c_565_n N_A_290_464#_M1034_s 0.00402708f $X=4.86 $Y=0.34
+ $X2=0 $Y2=0
cc_608 N_A_781_74#_M1029_d N_A_290_464#_c_1864_n 0.00620388f $X=4.04 $Y=1.84
+ $X2=0 $Y2=0
cc_609 N_A_781_74#_c_573_n N_A_290_464#_c_1864_n 0.0198453f $X=4.19 $Y=2.765
+ $X2=0 $Y2=0
cc_610 N_A_781_74#_c_574_n N_A_290_464#_c_1864_n 0.00206012f $X=5.64 $Y=2.99
+ $X2=0 $Y2=0
cc_611 N_A_781_74#_c_561_n N_A_290_464#_c_1860_n 0.00505434f $X=4.985 $Y=2.24
+ $X2=0 $Y2=0
cc_612 N_A_781_74#_c_564_n N_A_290_464#_c_1860_n 0.00569556f $X=4.045 $Y=0.505
+ $X2=0 $Y2=0
cc_613 N_A_781_74#_c_567_n N_A_290_464#_c_1860_n 0.0495574f $X=4.895 $Y=1.505
+ $X2=0 $Y2=0
cc_614 N_A_781_74#_c_568_n N_A_290_464#_c_1860_n 0.0228629f $X=4.895 $Y=1.37
+ $X2=0 $Y2=0
cc_615 N_A_781_74#_c_561_n N_A_290_464#_c_1866_n 0.00405887f $X=4.985 $Y=2.24
+ $X2=0 $Y2=0
cc_616 N_A_781_74#_c_573_n N_A_290_464#_c_1866_n 0.0120315f $X=4.19 $Y=2.765
+ $X2=0 $Y2=0
cc_617 N_A_781_74#_c_574_n N_A_290_464#_c_1866_n 0.0231346f $X=5.64 $Y=2.99
+ $X2=0 $Y2=0
cc_618 N_A_781_74#_c_564_n N_A_290_464#_c_1861_n 0.0232909f $X=4.045 $Y=0.505
+ $X2=0 $Y2=0
cc_619 N_A_781_74#_c_565_n N_A_290_464#_c_1861_n 0.0194638f $X=4.86 $Y=0.34
+ $X2=0 $Y2=0
cc_620 N_A_781_74#_c_568_n N_A_290_464#_c_1861_n 0.0240322f $X=4.895 $Y=1.37
+ $X2=0 $Y2=0
cc_621 N_A_781_74#_c_561_n N_A_290_464#_c_1867_n 0.00544732f $X=4.985 $Y=2.24
+ $X2=0 $Y2=0
cc_622 N_A_781_74#_c_574_n N_A_290_464#_c_1867_n 0.00542945f $X=5.64 $Y=2.99
+ $X2=0 $Y2=0
cc_623 N_A_781_74#_c_576_n N_A_290_464#_c_1867_n 0.01419f $X=4.925 $Y=1.535
+ $X2=0 $Y2=0
cc_624 N_A_781_74#_c_578_n A_1133_478# 0.00584471f $X=5.725 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_625 N_A_781_74#_c_584_n N_A_1600_347#_M1008_d 0.00559603f $X=8.66 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_626 N_A_781_74#_c_584_n N_A_1600_347#_c_1982_n 0.028219f $X=8.66 $Y=2.035
+ $X2=0 $Y2=0
cc_627 N_A_781_74#_c_569_n N_A_1600_347#_c_1982_n 0.00163009f $X=8.825 $Y=1.515
+ $X2=0 $Y2=0
cc_628 N_A_781_74#_c_570_n N_A_1600_347#_c_1982_n 8.50223e-19 $X=8.825 $Y=1.515
+ $X2=0 $Y2=0
cc_629 N_A_781_74#_c_590_n N_A_1600_347#_c_1982_n 0.00949462f $X=8.825 $Y=1.795
+ $X2=0 $Y2=0
cc_630 N_A_781_74#_c_584_n N_A_1600_347#_c_1983_n 0.0207253f $X=8.66 $Y=2.035
+ $X2=0 $Y2=0
cc_631 N_A_781_74#_c_590_n N_A_1600_347#_c_1983_n 0.001743f $X=8.825 $Y=1.795
+ $X2=0 $Y2=0
cc_632 N_A_781_74#_c_584_n N_A_1712_374#_M1035_s 0.00458277f $X=8.66 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_633 N_A_781_74#_c_586_n N_A_1712_374#_M1035_s 0.00138884f $X=8.745 $Y=1.95
+ $X2=-0.19 $Y2=-0.245
cc_634 N_A_781_74#_c_590_n N_A_1712_374#_c_2018_n 3.83337e-19 $X=8.825 $Y=1.795
+ $X2=0 $Y2=0
cc_635 N_A_781_74#_c_566_n N_VGND_c_2103_n 0.011924f $X=4.21 $Y=0.34 $X2=0 $Y2=0
cc_636 N_A_781_74#_M1004_g N_VGND_c_2109_n 0.00434272f $X=5.5 $Y=0.58 $X2=0
+ $Y2=0
cc_637 N_A_781_74#_c_565_n N_VGND_c_2109_n 0.0534972f $X=4.86 $Y=0.34 $X2=0
+ $Y2=0
cc_638 N_A_781_74#_c_566_n N_VGND_c_2109_n 0.0235688f $X=4.21 $Y=0.34 $X2=0
+ $Y2=0
cc_639 N_A_781_74#_M1024_g N_VGND_c_2113_n 0.00434272f $X=8.735 $Y=0.69 $X2=0
+ $Y2=0
cc_640 N_A_781_74#_M1004_g N_VGND_c_2117_n 0.00822443f $X=5.5 $Y=0.58 $X2=0
+ $Y2=0
cc_641 N_A_781_74#_M1024_g N_VGND_c_2117_n 0.00822232f $X=8.735 $Y=0.69 $X2=0
+ $Y2=0
cc_642 N_A_781_74#_c_565_n N_VGND_c_2117_n 0.0303548f $X=4.86 $Y=0.34 $X2=0
+ $Y2=0
cc_643 N_A_781_74#_c_566_n N_VGND_c_2117_n 0.0127152f $X=4.21 $Y=0.34 $X2=0
+ $Y2=0
cc_644 N_A_781_74#_M1024_g N_VGND_c_2121_n 0.00164121f $X=8.735 $Y=0.69 $X2=0
+ $Y2=0
cc_645 N_A_1163_48#_c_773_n N_A_995_74#_c_846_n 0.00856703f $X=6.125 $Y=1.635
+ $X2=0 $Y2=0
cc_646 N_A_1163_48#_c_774_n N_A_995_74#_c_846_n 9.45781e-19 $X=6.263 $Y=0.957
+ $X2=0 $Y2=0
cc_647 N_A_1163_48#_c_779_n N_A_995_74#_c_846_n 0.00129303f $X=6.935 $Y=1.802
+ $X2=0 $Y2=0
cc_648 N_A_1163_48#_c_775_n N_A_995_74#_c_846_n 0.00225195f $X=6.32 $Y=1.065
+ $X2=0 $Y2=0
cc_649 N_A_1163_48#_c_772_n N_A_995_74#_c_847_n 0.0132022f $X=6.11 $Y=1.965
+ $X2=0 $Y2=0
cc_650 N_A_1163_48#_c_777_n N_A_995_74#_c_847_n 0.00328197f $X=6.11 $Y=2.15
+ $X2=0 $Y2=0
cc_651 N_A_1163_48#_c_779_n N_A_995_74#_c_847_n 0.0179719f $X=6.935 $Y=1.802
+ $X2=0 $Y2=0
cc_652 N_A_1163_48#_c_780_n N_A_995_74#_c_847_n 0.00576399f $X=7.02 $Y=2.515
+ $X2=0 $Y2=0
cc_653 N_A_1163_48#_c_778_n N_A_995_74#_c_859_n 0.0109309f $X=6.11 $Y=2.24 $X2=0
+ $Y2=0
cc_654 N_A_1163_48#_c_780_n N_A_995_74#_c_859_n 0.00197687f $X=7.02 $Y=2.515
+ $X2=0 $Y2=0
cc_655 N_A_1163_48#_c_774_n N_A_995_74#_M1041_g 0.0162848f $X=6.263 $Y=0.957
+ $X2=0 $Y2=0
cc_656 N_A_1163_48#_c_775_n N_A_995_74#_M1041_g 0.00719364f $X=6.32 $Y=1.065
+ $X2=0 $Y2=0
cc_657 N_A_1163_48#_c_771_n N_A_995_74#_c_850_n 0.00195661f $X=5.89 $Y=0.9 $X2=0
+ $Y2=0
cc_658 N_A_1163_48#_c_773_n N_A_995_74#_c_850_n 5.28691e-19 $X=6.125 $Y=1.635
+ $X2=0 $Y2=0
cc_659 N_A_1163_48#_c_774_n N_A_995_74#_c_850_n 0.0186822f $X=6.263 $Y=0.957
+ $X2=0 $Y2=0
cc_660 N_A_1163_48#_c_775_n N_A_995_74#_c_850_n 2.95653e-19 $X=6.32 $Y=1.065
+ $X2=0 $Y2=0
cc_661 N_A_1163_48#_c_777_n N_A_995_74#_c_851_n 6.0134e-19 $X=6.11 $Y=2.15 $X2=0
+ $Y2=0
cc_662 N_A_1163_48#_c_772_n N_A_995_74#_c_852_n 0.00189647f $X=6.11 $Y=1.965
+ $X2=0 $Y2=0
cc_663 N_A_1163_48#_c_773_n N_A_995_74#_c_852_n 0.0123773f $X=6.125 $Y=1.635
+ $X2=0 $Y2=0
cc_664 N_A_1163_48#_c_774_n N_A_995_74#_c_852_n 0.0607821f $X=6.263 $Y=0.957
+ $X2=0 $Y2=0
cc_665 N_A_1163_48#_c_779_n N_A_995_74#_c_852_n 0.0499605f $X=6.935 $Y=1.802
+ $X2=0 $Y2=0
cc_666 N_A_1163_48#_c_775_n N_A_995_74#_c_852_n 0.00984239f $X=6.32 $Y=1.065
+ $X2=0 $Y2=0
cc_667 N_A_1163_48#_c_773_n N_A_995_74#_c_857_n 6.28152e-19 $X=6.125 $Y=1.635
+ $X2=0 $Y2=0
cc_668 N_A_1163_48#_c_774_n N_A_995_74#_c_857_n 0.0172613f $X=6.263 $Y=0.957
+ $X2=0 $Y2=0
cc_669 N_A_1163_48#_c_779_n N_A_995_74#_c_857_n 0.0307973f $X=6.935 $Y=1.802
+ $X2=0 $Y2=0
cc_670 N_A_1163_48#_c_775_n N_A_995_74#_c_857_n 6.81032e-19 $X=6.32 $Y=1.065
+ $X2=0 $Y2=0
cc_671 N_A_1163_48#_c_774_n N_SET_B_M1010_g 0.00113521f $X=6.263 $Y=0.957 $X2=0
+ $Y2=0
cc_672 N_A_1163_48#_c_779_n N_SET_B_c_984_n 0.00444569f $X=6.935 $Y=1.802 $X2=0
+ $Y2=0
cc_673 N_A_1163_48#_c_780_n N_SET_B_c_984_n 0.00171609f $X=7.02 $Y=2.515 $X2=0
+ $Y2=0
cc_674 N_A_1163_48#_c_780_n N_SET_B_c_999_n 0.00163696f $X=7.02 $Y=2.515 $X2=0
+ $Y2=0
cc_675 N_A_1163_48#_c_779_n N_SET_B_c_993_n 0.00248279f $X=6.935 $Y=1.802 $X2=0
+ $Y2=0
cc_676 N_A_1163_48#_c_779_n N_SET_B_c_996_n 0.00565296f $X=6.935 $Y=1.802 $X2=0
+ $Y2=0
cc_677 N_A_1163_48#_c_778_n N_A_594_74#_c_1156_n 0.0168752f $X=6.11 $Y=2.24
+ $X2=0 $Y2=0
cc_678 N_A_1163_48#_c_778_n N_A_594_74#_c_1157_n 0.010379f $X=6.11 $Y=2.24 $X2=0
+ $Y2=0
cc_679 N_A_1163_48#_c_778_n N_VPWR_c_1700_n 0.00802868f $X=6.11 $Y=2.24 $X2=0
+ $Y2=0
cc_680 N_A_1163_48#_c_778_n N_VPWR_c_1695_n 8.82884e-19 $X=6.11 $Y=2.24 $X2=0
+ $Y2=0
cc_681 N_A_1163_48#_c_774_n N_VGND_M1002_d 0.0034935f $X=6.263 $Y=0.957 $X2=0
+ $Y2=0
cc_682 N_A_1163_48#_c_771_n N_VGND_c_2104_n 0.00891566f $X=5.89 $Y=0.9 $X2=0
+ $Y2=0
cc_683 N_A_1163_48#_c_774_n N_VGND_c_2104_n 0.043708f $X=6.263 $Y=0.957 $X2=0
+ $Y2=0
cc_684 N_A_1163_48#_c_775_n N_VGND_c_2104_n 0.00185009f $X=6.32 $Y=1.065 $X2=0
+ $Y2=0
cc_685 N_A_1163_48#_c_771_n N_VGND_c_2109_n 0.00336577f $X=5.89 $Y=0.9 $X2=0
+ $Y2=0
cc_686 N_A_1163_48#_c_774_n N_VGND_c_2109_n 0.00250183f $X=6.263 $Y=0.957 $X2=0
+ $Y2=0
cc_687 N_A_1163_48#_c_771_n N_VGND_c_2117_n 0.00442062f $X=5.89 $Y=0.9 $X2=0
+ $Y2=0
cc_688 N_A_1163_48#_c_774_n N_VGND_c_2117_n 0.0245359f $X=6.263 $Y=0.957 $X2=0
+ $Y2=0
cc_689 N_A_1163_48#_c_774_n N_VGND_c_2120_n 0.0178253f $X=6.263 $Y=0.957 $X2=0
+ $Y2=0
cc_690 N_A_1163_48#_c_774_n N_VGND_c_2121_n 0.00571502f $X=6.263 $Y=0.957 $X2=0
+ $Y2=0
cc_691 N_A_995_74#_M1041_g N_SET_B_M1010_g 0.0332539f $X=6.98 $Y=0.58 $X2=0
+ $Y2=0
cc_692 N_A_995_74#_c_853_n N_SET_B_M1010_g 0.0165792f $X=7.835 $Y=0.99 $X2=0
+ $Y2=0
cc_693 N_A_995_74#_c_854_n N_SET_B_M1010_g 0.00202609f $X=8 $Y=1.285 $X2=0 $Y2=0
cc_694 N_A_995_74#_c_855_n N_SET_B_M1010_g 0.0044628f $X=8 $Y=1.285 $X2=0 $Y2=0
cc_695 N_A_995_74#_c_857_n N_SET_B_M1010_g 0.00534819f $X=6.89 $Y=1.355 $X2=0
+ $Y2=0
cc_696 N_A_995_74#_c_847_n N_SET_B_c_984_n 0.0061303f $X=6.795 $Y=2.15 $X2=0
+ $Y2=0
cc_697 N_A_995_74#_c_860_n N_SET_B_c_984_n 0.019642f $X=7.925 $Y=1.66 $X2=0
+ $Y2=0
cc_698 N_A_995_74#_c_855_n N_SET_B_c_984_n 0.00285979f $X=8 $Y=1.285 $X2=0 $Y2=0
cc_699 N_A_995_74#_c_859_n N_SET_B_c_999_n 0.0158843f $X=6.795 $Y=2.24 $X2=0
+ $Y2=0
cc_700 N_A_995_74#_c_860_n N_SET_B_c_999_n 0.00990574f $X=7.925 $Y=1.66 $X2=0
+ $Y2=0
cc_701 N_A_995_74#_c_860_n N_SET_B_c_992_n 0.00334164f $X=7.925 $Y=1.66 $X2=0
+ $Y2=0
cc_702 N_A_995_74#_c_853_n N_SET_B_c_992_n 0.00699145f $X=7.835 $Y=0.99 $X2=0
+ $Y2=0
cc_703 N_A_995_74#_c_854_n N_SET_B_c_992_n 0.00966112f $X=8 $Y=1.285 $X2=0 $Y2=0
cc_704 N_A_995_74#_c_855_n N_SET_B_c_992_n 0.0102907f $X=8 $Y=1.285 $X2=0 $Y2=0
cc_705 N_A_995_74#_c_846_n N_SET_B_c_993_n 7.48901e-19 $X=6.795 $Y=1.61 $X2=0
+ $Y2=0
cc_706 N_A_995_74#_c_853_n N_SET_B_c_993_n 0.0010997f $X=7.835 $Y=0.99 $X2=0
+ $Y2=0
cc_707 N_A_995_74#_c_846_n N_SET_B_c_995_n 0.0393842f $X=6.795 $Y=1.61 $X2=0
+ $Y2=0
cc_708 N_A_995_74#_c_853_n N_SET_B_c_995_n 0.00125903f $X=7.835 $Y=0.99 $X2=0
+ $Y2=0
cc_709 N_A_995_74#_c_854_n N_SET_B_c_995_n 7.13996e-19 $X=8 $Y=1.285 $X2=0 $Y2=0
cc_710 N_A_995_74#_c_855_n N_SET_B_c_995_n 0.021177f $X=8 $Y=1.285 $X2=0 $Y2=0
cc_711 N_A_995_74#_c_846_n N_SET_B_c_996_n 0.00180078f $X=6.795 $Y=1.61 $X2=0
+ $Y2=0
cc_712 N_A_995_74#_c_860_n N_SET_B_c_996_n 0.00226078f $X=7.925 $Y=1.66 $X2=0
+ $Y2=0
cc_713 N_A_995_74#_c_853_n N_SET_B_c_996_n 0.0242739f $X=7.835 $Y=0.99 $X2=0
+ $Y2=0
cc_714 N_A_995_74#_c_854_n N_SET_B_c_996_n 0.0129916f $X=8 $Y=1.285 $X2=0 $Y2=0
cc_715 N_A_995_74#_c_855_n N_SET_B_c_996_n 0.00320504f $X=8 $Y=1.285 $X2=0 $Y2=0
cc_716 N_A_995_74#_c_857_n N_SET_B_c_996_n 0.0213842f $X=6.89 $Y=1.355 $X2=0
+ $Y2=0
cc_717 N_A_995_74#_c_850_n N_A_594_74#_M1034_g 0.0026059f $X=5.285 $Y=0.58 $X2=0
+ $Y2=0
cc_718 N_A_995_74#_c_851_n N_A_594_74#_c_1156_n 9.68742e-19 $X=5.285 $Y=2.37
+ $X2=0 $Y2=0
cc_719 N_A_995_74#_c_863_n N_A_594_74#_c_1156_n 0.00355428f $X=5.285 $Y=2.55
+ $X2=0 $Y2=0
cc_720 N_A_995_74#_c_859_n N_A_594_74#_c_1157_n 0.00909901f $X=6.795 $Y=2.24
+ $X2=0 $Y2=0
cc_721 N_A_995_74#_c_860_n N_A_594_74#_c_1157_n 0.0103487f $X=7.925 $Y=1.66
+ $X2=0 $Y2=0
cc_722 N_A_995_74#_c_849_n N_A_1762_74#_c_1468_n 0.0023555f $X=8.345 $Y=1.12
+ $X2=0 $Y2=0
cc_723 N_A_995_74#_c_853_n N_A_1762_74#_c_1468_n 0.00454574f $X=7.835 $Y=0.99
+ $X2=0 $Y2=0
cc_724 N_A_995_74#_c_859_n N_VPWR_c_1700_n 0.00131022f $X=6.795 $Y=2.24 $X2=0
+ $Y2=0
cc_725 N_A_995_74#_c_860_n N_VPWR_c_1701_n 0.00457689f $X=7.925 $Y=1.66 $X2=0
+ $Y2=0
cc_726 N_A_995_74#_c_860_n N_VPWR_c_1695_n 9.39239e-19 $X=7.925 $Y=1.66 $X2=0
+ $Y2=0
cc_727 N_A_995_74#_c_851_n N_A_290_464#_c_1860_n 0.0051899f $X=5.285 $Y=2.37
+ $X2=0 $Y2=0
cc_728 N_A_995_74#_c_863_n N_A_290_464#_c_1866_n 0.0247867f $X=5.285 $Y=2.55
+ $X2=0 $Y2=0
cc_729 N_A_995_74#_c_851_n N_A_290_464#_c_1867_n 0.00876454f $X=5.285 $Y=2.37
+ $X2=0 $Y2=0
cc_730 N_A_995_74#_c_863_n N_A_290_464#_c_1867_n 7.40762e-19 $X=5.285 $Y=2.55
+ $X2=0 $Y2=0
cc_731 N_A_995_74#_c_860_n N_A_1600_347#_c_1983_n 0.00674223f $X=7.925 $Y=1.66
+ $X2=0 $Y2=0
cc_732 N_A_995_74#_c_860_n N_A_1712_374#_c_2020_n 0.00299587f $X=7.925 $Y=1.66
+ $X2=0 $Y2=0
cc_733 N_A_995_74#_c_853_n N_VGND_M1010_d 0.00962076f $X=7.835 $Y=0.99 $X2=0
+ $Y2=0
cc_734 N_A_995_74#_M1041_g N_VGND_c_2104_n 0.00317476f $X=6.98 $Y=0.58 $X2=0
+ $Y2=0
cc_735 N_A_995_74#_c_850_n N_VGND_c_2104_n 0.00319235f $X=5.285 $Y=0.58 $X2=0
+ $Y2=0
cc_736 N_A_995_74#_c_850_n N_VGND_c_2109_n 0.0109942f $X=5.285 $Y=0.58 $X2=0
+ $Y2=0
cc_737 N_A_995_74#_c_849_n N_VGND_c_2113_n 0.00383152f $X=8.345 $Y=1.12 $X2=0
+ $Y2=0
cc_738 N_A_995_74#_M1041_g N_VGND_c_2117_n 0.0082231f $X=6.98 $Y=0.58 $X2=0
+ $Y2=0
cc_739 N_A_995_74#_c_849_n N_VGND_c_2117_n 0.00752635f $X=8.345 $Y=1.12 $X2=0
+ $Y2=0
cc_740 N_A_995_74#_c_850_n N_VGND_c_2117_n 0.00904371f $X=5.285 $Y=0.58 $X2=0
+ $Y2=0
cc_741 N_A_995_74#_M1041_g N_VGND_c_2120_n 0.00433139f $X=6.98 $Y=0.58 $X2=0
+ $Y2=0
cc_742 N_A_995_74#_c_849_n N_VGND_c_2121_n 0.0135277f $X=8.345 $Y=1.12 $X2=0
+ $Y2=0
cc_743 N_A_995_74#_c_853_n N_VGND_c_2121_n 0.0561832f $X=7.835 $Y=0.99 $X2=0
+ $Y2=0
cc_744 N_A_995_74#_c_855_n N_VGND_c_2121_n 0.00421382f $X=8 $Y=1.285 $X2=0 $Y2=0
cc_745 N_SET_B_c_999_n N_A_594_74#_c_1157_n 0.00980497f $X=7.385 $Y=2.24 $X2=0
+ $Y2=0
cc_746 N_SET_B_c_991_n N_A_594_74#_M1000_g 5.49097e-19 $X=10.585 $Y=1.665 $X2=0
+ $Y2=0
cc_747 N_SET_B_c_992_n N_A_594_74#_M1000_g 4.75412e-19 $X=9.695 $Y=1.665 $X2=0
+ $Y2=0
cc_748 SET_B N_A_594_74#_M1000_g 6.71157e-19 $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_749 N_SET_B_c_991_n N_A_594_74#_c_1147_n 9.87584e-19 $X=10.585 $Y=1.665 $X2=0
+ $Y2=0
cc_750 N_SET_B_c_992_n N_A_594_74#_c_1147_n 0.0035987f $X=9.695 $Y=1.665 $X2=0
+ $Y2=0
cc_751 SET_B N_A_594_74#_c_1147_n 7.37013e-19 $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_752 N_SET_B_c_988_n N_A_1924_48#_c_1319_n 0.00789413f $X=10.765 $Y=1.775
+ $X2=0 $Y2=0
cc_753 N_SET_B_c_989_n N_A_1924_48#_c_1319_n 8.51789e-19 $X=10.75 $Y=1.42 $X2=0
+ $Y2=0
cc_754 N_SET_B_c_991_n N_A_1924_48#_c_1319_n 0.0133161f $X=10.585 $Y=1.665 $X2=0
+ $Y2=0
cc_755 SET_B N_A_1924_48#_c_1319_n 0.0020819f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_756 N_SET_B_c_991_n N_A_1924_48#_c_1332_n 0.00262239f $X=10.585 $Y=1.665
+ $X2=0 $Y2=0
cc_757 N_SET_B_c_1001_n N_A_1924_48#_c_1334_n 0.00815304f $X=10.89 $Y=2.465
+ $X2=0 $Y2=0
cc_758 N_SET_B_c_987_n N_A_1924_48#_c_1320_n 0.0101943f $X=10.31 $Y=0.94 $X2=0
+ $Y2=0
cc_759 N_SET_B_c_997_n N_A_1924_48#_c_1320_n 0.00487711f $X=10.75 $Y=1.255 $X2=0
+ $Y2=0
cc_760 N_SET_B_c_985_n N_A_1924_48#_c_1321_n 0.0212296f $X=10.235 $Y=0.865 $X2=0
+ $Y2=0
cc_761 N_SET_B_c_989_n N_A_1924_48#_c_1322_n 0.00158234f $X=10.75 $Y=1.42 $X2=0
+ $Y2=0
cc_762 N_SET_B_c_990_n N_A_1924_48#_c_1322_n 0.00789413f $X=10.75 $Y=1.42 $X2=0
+ $Y2=0
cc_763 N_SET_B_c_991_n N_A_1924_48#_c_1322_n 0.00419833f $X=10.585 $Y=1.665
+ $X2=0 $Y2=0
cc_764 N_SET_B_c_992_n N_A_1924_48#_c_1322_n 0.00205438f $X=9.695 $Y=1.665 $X2=0
+ $Y2=0
cc_765 SET_B N_A_1924_48#_c_1322_n 0.00539133f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_766 N_SET_B_c_1000_n N_A_1924_48#_c_1335_n 0.0150577f $X=10.89 $Y=2.375 $X2=0
+ $Y2=0
cc_767 N_SET_B_c_986_n N_A_1924_48#_c_1323_n 0.0117431f $X=10.55 $Y=0.94 $X2=0
+ $Y2=0
cc_768 N_SET_B_c_987_n N_A_1924_48#_c_1323_n 0.0106933f $X=10.31 $Y=0.94 $X2=0
+ $Y2=0
cc_769 N_SET_B_c_989_n N_A_1924_48#_c_1323_n 0.02412f $X=10.75 $Y=1.42 $X2=0
+ $Y2=0
cc_770 N_SET_B_c_990_n N_A_1924_48#_c_1323_n 0.00273565f $X=10.75 $Y=1.42 $X2=0
+ $Y2=0
cc_771 N_SET_B_c_991_n N_A_1924_48#_c_1323_n 0.0227767f $X=10.585 $Y=1.665 $X2=0
+ $Y2=0
cc_772 SET_B N_A_1924_48#_c_1323_n 6.64033e-19 $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_773 N_SET_B_c_997_n N_A_1924_48#_c_1323_n 0.00520213f $X=10.75 $Y=1.255 $X2=0
+ $Y2=0
cc_774 N_SET_B_c_989_n N_A_1924_48#_c_1325_n 0.00196616f $X=10.75 $Y=1.42 $X2=0
+ $Y2=0
cc_775 N_SET_B_c_997_n N_A_1924_48#_c_1325_n 9.74678e-19 $X=10.75 $Y=1.255 $X2=0
+ $Y2=0
cc_776 N_SET_B_c_989_n N_A_1924_48#_c_1327_n 0.00835006f $X=10.75 $Y=1.42 $X2=0
+ $Y2=0
cc_777 N_SET_B_c_990_n N_A_1924_48#_c_1327_n 6.8943e-19 $X=10.75 $Y=1.42 $X2=0
+ $Y2=0
cc_778 N_SET_B_c_1001_n N_A_1924_48#_c_1336_n 8.72078e-19 $X=10.89 $Y=2.465
+ $X2=0 $Y2=0
cc_779 N_SET_B_c_991_n N_A_1924_48#_c_1367_n 0.00742107f $X=10.585 $Y=1.665
+ $X2=0 $Y2=0
cc_780 N_SET_B_c_992_n N_A_1924_48#_c_1367_n 0.00267727f $X=9.695 $Y=1.665 $X2=0
+ $Y2=0
cc_781 SET_B N_A_1924_48#_c_1367_n 0.00653525f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_782 N_SET_B_c_997_n N_A_1924_48#_c_1367_n 8.32131e-19 $X=10.75 $Y=1.255 $X2=0
+ $Y2=0
cc_783 N_SET_B_c_985_n N_A_1762_74#_c_1455_n 0.00514966f $X=10.235 $Y=0.865
+ $X2=0 $Y2=0
cc_784 N_SET_B_c_989_n N_A_1762_74#_c_1456_n 0.00136743f $X=10.75 $Y=1.42 $X2=0
+ $Y2=0
cc_785 N_SET_B_c_990_n N_A_1762_74#_c_1456_n 0.01211f $X=10.75 $Y=1.42 $X2=0
+ $Y2=0
cc_786 N_SET_B_c_997_n N_A_1762_74#_c_1456_n 0.00524052f $X=10.75 $Y=1.255 $X2=0
+ $Y2=0
cc_787 N_SET_B_c_986_n N_A_1762_74#_c_1462_n 0.00859503f $X=10.55 $Y=0.94 $X2=0
+ $Y2=0
cc_788 N_SET_B_c_990_n N_A_1762_74#_c_1462_n 5.62189e-19 $X=10.75 $Y=1.42 $X2=0
+ $Y2=0
cc_789 N_SET_B_c_988_n N_A_1762_74#_c_1463_n 0.01211f $X=10.765 $Y=1.775 $X2=0
+ $Y2=0
cc_790 N_SET_B_c_1003_n N_A_1762_74#_c_1463_n 0.0100137f $X=10.765 $Y=1.925
+ $X2=0 $Y2=0
cc_791 N_SET_B_c_989_n N_A_1762_74#_c_1463_n 2.72084e-19 $X=10.75 $Y=1.42 $X2=0
+ $Y2=0
cc_792 N_SET_B_c_991_n N_A_1762_74#_c_1481_n 0.0175055f $X=10.585 $Y=1.665 $X2=0
+ $Y2=0
cc_793 N_SET_B_c_992_n N_A_1762_74#_c_1481_n 0.0126053f $X=9.695 $Y=1.665 $X2=0
+ $Y2=0
cc_794 SET_B N_A_1762_74#_c_1481_n 0.008126f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_795 N_SET_B_c_1000_n N_A_1762_74#_c_1482_n 0.0197896f $X=10.89 $Y=2.375 $X2=0
+ $Y2=0
cc_796 N_SET_B_c_1003_n N_A_1762_74#_c_1482_n 0.00251056f $X=10.765 $Y=1.925
+ $X2=0 $Y2=0
cc_797 N_SET_B_c_989_n N_A_1762_74#_c_1482_n 0.0257549f $X=10.75 $Y=1.42 $X2=0
+ $Y2=0
cc_798 N_SET_B_c_991_n N_A_1762_74#_c_1482_n 0.0207168f $X=10.585 $Y=1.665 $X2=0
+ $Y2=0
cc_799 N_SET_B_c_1000_n N_A_1762_74#_c_1467_n 0.00461877f $X=10.89 $Y=2.375
+ $X2=0 $Y2=0
cc_800 N_SET_B_c_988_n N_A_1762_74#_c_1467_n 9.04429e-19 $X=10.765 $Y=1.775
+ $X2=0 $Y2=0
cc_801 N_SET_B_c_1003_n N_A_1762_74#_c_1467_n 0.00657737f $X=10.765 $Y=1.925
+ $X2=0 $Y2=0
cc_802 N_SET_B_c_989_n N_A_1762_74#_c_1467_n 0.0192851f $X=10.75 $Y=1.42 $X2=0
+ $Y2=0
cc_803 N_SET_B_c_992_n N_A_1762_74#_c_1468_n 0.00926935f $X=9.695 $Y=1.665 $X2=0
+ $Y2=0
cc_804 N_SET_B_c_992_n N_A_1762_74#_c_1484_n 0.00844651f $X=9.695 $Y=1.665 $X2=0
+ $Y2=0
cc_805 N_SET_B_c_991_n N_A_1762_74#_c_1469_n 0.00721247f $X=10.585 $Y=1.665
+ $X2=0 $Y2=0
cc_806 N_SET_B_c_992_n N_A_1762_74#_c_1469_n 0.0193428f $X=9.695 $Y=1.665 $X2=0
+ $Y2=0
cc_807 SET_B N_A_1762_74#_c_1469_n 0.00234368f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_808 N_SET_B_c_1000_n N_A_1762_74#_c_1486_n 0.00332493f $X=10.89 $Y=2.375
+ $X2=0 $Y2=0
cc_809 N_SET_B_c_991_n N_A_1762_74#_c_1486_n 0.0133991f $X=10.585 $Y=1.665 $X2=0
+ $Y2=0
cc_810 N_SET_B_c_1001_n N_A_1762_74#_c_1487_n 0.0069352f $X=10.89 $Y=2.465 $X2=0
+ $Y2=0
cc_811 N_SET_B_c_1001_n N_A_1762_74#_c_1488_n 0.00554984f $X=10.89 $Y=2.465
+ $X2=0 $Y2=0
cc_812 N_SET_B_c_992_n N_VPWR_M1013_d 0.00187641f $X=9.695 $Y=1.665 $X2=0 $Y2=0
cc_813 N_SET_B_c_996_n N_VPWR_M1013_d 0.0010181f $X=7.46 $Y=1.41 $X2=0 $Y2=0
cc_814 N_SET_B_c_999_n N_VPWR_c_1701_n 0.00390712f $X=7.385 $Y=2.24 $X2=0 $Y2=0
cc_815 N_SET_B_c_1001_n N_VPWR_c_1702_n 0.00435973f $X=10.89 $Y=2.465 $X2=0
+ $Y2=0
cc_816 N_SET_B_c_1001_n N_VPWR_c_1713_n 0.00445602f $X=10.89 $Y=2.465 $X2=0
+ $Y2=0
cc_817 N_SET_B_c_1001_n N_VPWR_c_1695_n 0.00900303f $X=10.89 $Y=2.465 $X2=0
+ $Y2=0
cc_818 N_SET_B_c_992_n N_A_1600_347#_M1008_d 0.00240778f $X=9.695 $Y=1.665
+ $X2=-0.19 $Y2=-0.245
cc_819 N_SET_B_c_992_n N_A_1600_347#_c_1982_n 0.00584852f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_820 N_SET_B_c_985_n N_VGND_c_2113_n 0.00384553f $X=10.235 $Y=0.865 $X2=0
+ $Y2=0
cc_821 N_SET_B_M1010_g N_VGND_c_2117_n 0.00913019f $X=7.37 $Y=0.58 $X2=0 $Y2=0
cc_822 N_SET_B_c_985_n N_VGND_c_2117_n 0.00758569f $X=10.235 $Y=0.865 $X2=0
+ $Y2=0
cc_823 N_SET_B_M1010_g N_VGND_c_2120_n 0.00461464f $X=7.37 $Y=0.58 $X2=0 $Y2=0
cc_824 N_SET_B_M1010_g N_VGND_c_2121_n 0.00576207f $X=7.37 $Y=0.58 $X2=0 $Y2=0
cc_825 N_SET_B_c_985_n N_VGND_c_2122_n 0.0127134f $X=10.235 $Y=0.865 $X2=0 $Y2=0
cc_826 N_SET_B_c_986_n N_VGND_c_2122_n 0.00878086f $X=10.55 $Y=0.94 $X2=0 $Y2=0
cc_827 N_A_594_74#_M1000_g N_A_1924_48#_c_1319_n 0.00544029f $X=9.305 $Y=0.58
+ $X2=0 $Y2=0
cc_828 N_A_594_74#_M1009_g N_A_1924_48#_c_1319_n 0.0177347f $X=9.44 $Y=2.37
+ $X2=0 $Y2=0
cc_829 N_A_594_74#_c_1147_n N_A_1924_48#_c_1319_n 0.00531267f $X=9.44 $Y=1.72
+ $X2=0 $Y2=0
cc_830 N_A_594_74#_M1000_g N_A_1924_48#_c_1321_n 0.06105f $X=9.305 $Y=0.58 $X2=0
+ $Y2=0
cc_831 N_A_594_74#_M1000_g N_A_1924_48#_c_1367_n 0.00104919f $X=9.305 $Y=0.58
+ $X2=0 $Y2=0
cc_832 N_A_594_74#_M1009_g N_A_1762_74#_c_1481_n 0.00922235f $X=9.44 $Y=2.37
+ $X2=0 $Y2=0
cc_833 N_A_594_74#_M1000_g N_A_1762_74#_c_1468_n 0.0256745f $X=9.305 $Y=0.58
+ $X2=0 $Y2=0
cc_834 N_A_594_74#_M1009_g N_A_1762_74#_c_1484_n 0.00417777f $X=9.44 $Y=2.37
+ $X2=0 $Y2=0
cc_835 N_A_594_74#_M1000_g N_A_1762_74#_c_1469_n 0.0174369f $X=9.305 $Y=0.58
+ $X2=0 $Y2=0
cc_836 N_A_594_74#_M1009_g N_A_1762_74#_c_1469_n 0.00174384f $X=9.44 $Y=2.37
+ $X2=0 $Y2=0
cc_837 N_A_594_74#_c_1147_n N_A_1762_74#_c_1469_n 0.00690274f $X=9.44 $Y=1.72
+ $X2=0 $Y2=0
cc_838 N_A_594_74#_M1009_g N_A_1762_74#_c_1486_n 6.75362e-19 $X=9.44 $Y=2.37
+ $X2=0 $Y2=0
cc_839 N_A_594_74#_c_1164_n N_VPWR_M1019_d 0.00220209f $X=3.885 $Y=1.905 $X2=0
+ $Y2=0
cc_840 N_A_594_74#_c_1140_n N_VPWR_c_1699_n 0.00666461f $X=3.965 $Y=1.765 $X2=0
+ $Y2=0
cc_841 N_A_594_74#_c_1155_n N_VPWR_c_1699_n 0.00246251f $X=4.55 $Y=3.15 $X2=0
+ $Y2=0
cc_842 N_A_594_74#_c_1156_n N_VPWR_c_1700_n 4.8564e-19 $X=5.59 $Y=2.885 $X2=0
+ $Y2=0
cc_843 N_A_594_74#_c_1157_n N_VPWR_c_1700_n 0.0213655f $X=9.35 $Y=3.15 $X2=0
+ $Y2=0
cc_844 N_A_594_74#_c_1159_n N_VPWR_c_1700_n 9.5628e-19 $X=5.59 $Y=3.15 $X2=0
+ $Y2=0
cc_845 N_A_594_74#_c_1157_n N_VPWR_c_1701_n 0.0170937f $X=9.35 $Y=3.15 $X2=0
+ $Y2=0
cc_846 N_A_594_74#_c_1140_n N_VPWR_c_1705_n 0.00413917f $X=3.965 $Y=1.765 $X2=0
+ $Y2=0
cc_847 N_A_594_74#_c_1155_n N_VPWR_c_1705_n 0.043034f $X=4.55 $Y=3.15 $X2=0
+ $Y2=0
cc_848 N_A_594_74#_c_1157_n N_VPWR_c_1707_n 0.0290731f $X=9.35 $Y=3.15 $X2=0
+ $Y2=0
cc_849 N_A_594_74#_c_1157_n N_VPWR_c_1709_n 0.0433129f $X=9.35 $Y=3.15 $X2=0
+ $Y2=0
cc_850 N_A_594_74#_c_1140_n N_VPWR_c_1695_n 0.00818274f $X=3.965 $Y=1.765 $X2=0
+ $Y2=0
cc_851 N_A_594_74#_c_1154_n N_VPWR_c_1695_n 0.0223434f $X=5.5 $Y=3.15 $X2=0
+ $Y2=0
cc_852 N_A_594_74#_c_1155_n N_VPWR_c_1695_n 0.00599976f $X=4.55 $Y=3.15 $X2=0
+ $Y2=0
cc_853 N_A_594_74#_c_1157_n N_VPWR_c_1695_n 0.0988023f $X=9.35 $Y=3.15 $X2=0
+ $Y2=0
cc_854 N_A_594_74#_c_1159_n N_VPWR_c_1695_n 0.0044131f $X=5.59 $Y=3.15 $X2=0
+ $Y2=0
cc_855 N_A_594_74#_c_1161_n N_VPWR_c_1695_n 0.00674811f $X=9.44 $Y=3.15 $X2=0
+ $Y2=0
cc_856 N_A_594_74#_c_1151_n N_A_290_464#_c_1857_n 0.00564313f $X=3.067 $Y=1.01
+ $X2=0 $Y2=0
cc_857 N_A_594_74#_c_1149_n N_A_290_464#_c_1859_n 0.00146536f $X=3.02 $Y=1.82
+ $X2=0 $Y2=0
cc_858 N_A_594_74#_M1019_s N_A_290_464#_c_1863_n 0.00819019f $X=3.15 $Y=1.84
+ $X2=0 $Y2=0
cc_859 N_A_594_74#_c_1163_n N_A_290_464#_c_1863_n 0.014265f $X=3.105 $Y=1.985
+ $X2=0 $Y2=0
cc_860 N_A_594_74#_c_1164_n N_A_290_464#_c_1863_n 0.00535916f $X=3.885 $Y=1.905
+ $X2=0 $Y2=0
cc_861 N_A_594_74#_c_1166_n N_A_290_464#_c_1863_n 0.0223261f $X=3.29 $Y=1.985
+ $X2=0 $Y2=0
cc_862 N_A_594_74#_c_1140_n N_A_290_464#_c_1864_n 0.0145127f $X=3.965 $Y=1.765
+ $X2=0 $Y2=0
cc_863 N_A_594_74#_c_1141_n N_A_290_464#_c_1864_n 0.00236726f $X=4.4 $Y=1.385
+ $X2=0 $Y2=0
cc_864 N_A_594_74#_c_1142_n N_A_290_464#_c_1864_n 0.00401194f $X=4.475 $Y=3.075
+ $X2=0 $Y2=0
cc_865 N_A_594_74#_c_1164_n N_A_290_464#_c_1864_n 0.019495f $X=3.885 $Y=1.905
+ $X2=0 $Y2=0
cc_866 N_A_594_74#_c_1139_n N_A_290_464#_c_1860_n 0.00100658f $X=3.83 $Y=1.22
+ $X2=0 $Y2=0
cc_867 N_A_594_74#_c_1140_n N_A_290_464#_c_1860_n 0.00169219f $X=3.965 $Y=1.765
+ $X2=0 $Y2=0
cc_868 N_A_594_74#_c_1142_n N_A_290_464#_c_1860_n 0.01579f $X=4.475 $Y=3.075
+ $X2=0 $Y2=0
cc_869 N_A_594_74#_c_1143_n N_A_290_464#_c_1860_n 0.00466065f $X=4.825 $Y=1.055
+ $X2=0 $Y2=0
cc_870 N_A_594_74#_M1034_g N_A_290_464#_c_1860_n 0.00101293f $X=4.9 $Y=0.58
+ $X2=0 $Y2=0
cc_871 N_A_594_74#_c_1146_n N_A_290_464#_c_1860_n 0.0200212f $X=4.475 $Y=1.055
+ $X2=0 $Y2=0
cc_872 N_A_594_74#_c_1164_n N_A_290_464#_c_1860_n 0.011652f $X=3.885 $Y=1.905
+ $X2=0 $Y2=0
cc_873 N_A_594_74#_c_1150_n N_A_290_464#_c_1860_n 0.0379515f $X=4.05 $Y=1.385
+ $X2=0 $Y2=0
cc_874 N_A_594_74#_c_1142_n N_A_290_464#_c_1866_n 0.00669365f $X=4.475 $Y=3.075
+ $X2=0 $Y2=0
cc_875 N_A_594_74#_c_1140_n N_A_290_464#_c_1950_n 0.00280588f $X=3.965 $Y=1.765
+ $X2=0 $Y2=0
cc_876 N_A_594_74#_c_1164_n N_A_290_464#_c_1950_n 0.00920256f $X=3.885 $Y=1.905
+ $X2=0 $Y2=0
cc_877 N_A_594_74#_c_1143_n N_A_290_464#_c_1861_n 0.00424734f $X=4.825 $Y=1.055
+ $X2=0 $Y2=0
cc_878 N_A_594_74#_M1034_g N_A_290_464#_c_1861_n 0.00662014f $X=4.9 $Y=0.58
+ $X2=0 $Y2=0
cc_879 N_A_594_74#_c_1146_n N_A_290_464#_c_1861_n 0.00145165f $X=4.475 $Y=1.055
+ $X2=0 $Y2=0
cc_880 N_A_594_74#_c_1142_n N_A_290_464#_c_1867_n 0.00797618f $X=4.475 $Y=3.075
+ $X2=0 $Y2=0
cc_881 N_A_594_74#_c_1157_n N_A_1600_347#_c_1982_n 0.00699557f $X=9.35 $Y=3.15
+ $X2=0 $Y2=0
cc_882 N_A_594_74#_M1009_g N_A_1600_347#_c_1982_n 0.011253f $X=9.44 $Y=2.37
+ $X2=0 $Y2=0
cc_883 N_A_594_74#_c_1147_n N_A_1600_347#_c_1982_n 3.58975e-19 $X=9.44 $Y=1.72
+ $X2=0 $Y2=0
cc_884 N_A_594_74#_c_1157_n N_A_1600_347#_c_1983_n 0.00624256f $X=9.35 $Y=3.15
+ $X2=0 $Y2=0
cc_885 N_A_594_74#_M1009_g N_A_1600_347#_c_1984_n 0.00658375f $X=9.44 $Y=2.37
+ $X2=0 $Y2=0
cc_886 N_A_594_74#_c_1157_n N_A_1712_374#_c_2018_n 0.0102245f $X=9.35 $Y=3.15
+ $X2=0 $Y2=0
cc_887 N_A_594_74#_M1009_g N_A_1712_374#_c_2018_n 0.00550167f $X=9.44 $Y=2.37
+ $X2=0 $Y2=0
cc_888 N_A_594_74#_c_1161_n N_A_1712_374#_c_2018_n 0.0101957f $X=9.44 $Y=3.15
+ $X2=0 $Y2=0
cc_889 N_A_594_74#_M1009_g N_A_1712_374#_c_2019_n 0.00465095f $X=9.44 $Y=2.37
+ $X2=0 $Y2=0
cc_890 N_A_594_74#_c_1157_n N_A_1712_374#_c_2020_n 0.00754643f $X=9.35 $Y=3.15
+ $X2=0 $Y2=0
cc_891 N_A_594_74#_M1009_g N_A_1712_374#_c_2020_n 0.00572817f $X=9.44 $Y=2.37
+ $X2=0 $Y2=0
cc_892 N_A_594_74#_c_1161_n N_A_1712_374#_c_2020_n 3.04883e-19 $X=9.44 $Y=3.15
+ $X2=0 $Y2=0
cc_893 N_A_594_74#_c_1148_n N_VGND_c_2102_n 0.0237473f $X=3.115 $Y=0.505 $X2=0
+ $Y2=0
cc_894 N_A_594_74#_c_1139_n N_VGND_c_2103_n 0.00470925f $X=3.83 $Y=1.22 $X2=0
+ $Y2=0
cc_895 N_A_594_74#_c_1148_n N_VGND_c_2103_n 0.0251347f $X=3.115 $Y=0.505 $X2=0
+ $Y2=0
cc_896 N_A_594_74#_c_1139_n N_VGND_c_2109_n 0.00430908f $X=3.83 $Y=1.22 $X2=0
+ $Y2=0
cc_897 N_A_594_74#_M1034_g N_VGND_c_2109_n 0.00278159f $X=4.9 $Y=0.58 $X2=0
+ $Y2=0
cc_898 N_A_594_74#_c_1148_n N_VGND_c_2112_n 0.0122205f $X=3.115 $Y=0.505 $X2=0
+ $Y2=0
cc_899 N_A_594_74#_M1000_g N_VGND_c_2113_n 0.00292646f $X=9.305 $Y=0.58 $X2=0
+ $Y2=0
cc_900 N_A_594_74#_c_1139_n N_VGND_c_2117_n 0.00821169f $X=3.83 $Y=1.22 $X2=0
+ $Y2=0
cc_901 N_A_594_74#_M1034_g N_VGND_c_2117_n 0.00359882f $X=4.9 $Y=0.58 $X2=0
+ $Y2=0
cc_902 N_A_594_74#_M1000_g N_VGND_c_2117_n 0.00359032f $X=9.305 $Y=0.58 $X2=0
+ $Y2=0
cc_903 N_A_594_74#_c_1148_n N_VGND_c_2117_n 0.00976972f $X=3.115 $Y=0.505 $X2=0
+ $Y2=0
cc_904 N_A_1924_48#_c_1324_n N_A_1762_74#_c_1455_n 0.0142415f $X=11.23 $Y=0.58
+ $X2=0 $Y2=0
cc_905 N_A_1924_48#_c_1325_n N_A_1762_74#_c_1456_n 0.00858132f $X=11.31 $Y=1.3
+ $X2=0 $Y2=0
cc_906 N_A_1924_48#_c_1327_n N_A_1762_74#_c_1456_n 0.0084379f $X=11.395 $Y=1.385
+ $X2=0 $Y2=0
cc_907 N_A_1924_48#_c_1328_n N_A_1762_74#_c_1456_n 6.40251e-19 $X=12.15 $Y=2.18
+ $X2=0 $Y2=0
cc_908 N_A_1924_48#_c_1330_n N_A_1762_74#_c_1456_n 0.00224676f $X=11.23 $Y=0.985
+ $X2=0 $Y2=0
cc_909 N_A_1924_48#_c_1336_n N_A_1762_74#_c_1470_n 0.00475156f $X=11.665 $Y=2.75
+ $X2=0 $Y2=0
cc_910 N_A_1924_48#_c_1337_n N_A_1762_74#_c_1470_n 0.019987f $X=12.065 $Y=2.265
+ $X2=0 $Y2=0
cc_911 N_A_1924_48#_c_1336_n N_A_1762_74#_c_1471_n 0.00510373f $X=11.665 $Y=2.75
+ $X2=0 $Y2=0
cc_912 N_A_1924_48#_c_1325_n N_A_1762_74#_M1005_g 0.00247796f $X=11.31 $Y=1.3
+ $X2=0 $Y2=0
cc_913 N_A_1924_48#_c_1326_n N_A_1762_74#_M1005_g 0.0175404f $X=12.065 $Y=1.385
+ $X2=0 $Y2=0
cc_914 N_A_1924_48#_c_1328_n N_A_1762_74#_M1005_g 0.00604112f $X=12.15 $Y=2.18
+ $X2=0 $Y2=0
cc_915 N_A_1924_48#_c_1328_n N_A_1762_74#_c_1458_n 0.00532618f $X=12.15 $Y=2.18
+ $X2=0 $Y2=0
cc_916 N_A_1924_48#_c_1326_n N_A_1762_74#_c_1459_n 8.26299e-19 $X=12.065
+ $Y=1.385 $X2=0 $Y2=0
cc_917 N_A_1924_48#_c_1337_n N_A_1762_74#_c_1459_n 7.87495e-19 $X=12.065
+ $Y=2.265 $X2=0 $Y2=0
cc_918 N_A_1924_48#_c_1328_n N_A_1762_74#_c_1459_n 0.0128536f $X=12.15 $Y=2.18
+ $X2=0 $Y2=0
cc_919 N_A_1924_48#_c_1337_n N_A_1762_74#_c_1474_n 0.00156231f $X=12.065
+ $Y=2.265 $X2=0 $Y2=0
cc_920 N_A_1924_48#_c_1328_n N_A_1762_74#_c_1474_n 0.0033623f $X=12.15 $Y=2.18
+ $X2=0 $Y2=0
cc_921 N_A_1924_48#_c_1323_n N_A_1762_74#_c_1462_n 0.00958405f $X=11.065
+ $Y=0.985 $X2=0 $Y2=0
cc_922 N_A_1924_48#_c_1324_n N_A_1762_74#_c_1462_n 0.00829222f $X=11.23 $Y=0.58
+ $X2=0 $Y2=0
cc_923 N_A_1924_48#_c_1330_n N_A_1762_74#_c_1462_n 0.00686615f $X=11.23 $Y=0.985
+ $X2=0 $Y2=0
cc_924 N_A_1924_48#_c_1326_n N_A_1762_74#_c_1464_n 0.0110481f $X=12.065 $Y=1.385
+ $X2=0 $Y2=0
cc_925 N_A_1924_48#_c_1337_n N_A_1762_74#_c_1464_n 0.00108592f $X=12.065
+ $Y=2.265 $X2=0 $Y2=0
cc_926 N_A_1924_48#_c_1338_n N_A_1762_74#_c_1464_n 0.00578596f $X=11.75 $Y=2.265
+ $X2=0 $Y2=0
cc_927 N_A_1924_48#_c_1319_n N_A_1762_74#_c_1481_n 0.0110991f $X=9.955 $Y=2.165
+ $X2=0 $Y2=0
cc_928 N_A_1924_48#_c_1322_n N_A_1762_74#_c_1481_n 0.00311771f $X=9.825 $Y=1.405
+ $X2=0 $Y2=0
cc_929 N_A_1924_48#_c_1319_n N_A_1762_74#_c_1482_n 3.79939e-19 $X=9.955 $Y=2.165
+ $X2=0 $Y2=0
cc_930 N_A_1924_48#_c_1332_n N_A_1762_74#_c_1482_n 0.00658213f $X=10.35 $Y=2.24
+ $X2=0 $Y2=0
cc_931 N_A_1924_48#_c_1335_n N_A_1762_74#_c_1482_n 0.0126377f $X=10.44 $Y=2.24
+ $X2=0 $Y2=0
cc_932 N_A_1924_48#_c_1327_n N_A_1762_74#_c_1467_n 0.00457115f $X=11.395
+ $Y=1.385 $X2=0 $Y2=0
cc_933 N_A_1924_48#_c_1338_n N_A_1762_74#_c_1467_n 0.0119447f $X=11.75 $Y=2.265
+ $X2=0 $Y2=0
cc_934 N_A_1924_48#_c_1330_n N_A_1762_74#_c_1467_n 0.00460453f $X=11.23 $Y=0.985
+ $X2=0 $Y2=0
cc_935 N_A_1924_48#_c_1326_n N_A_1762_74#_c_1568_n 0.0375032f $X=12.065 $Y=1.385
+ $X2=0 $Y2=0
cc_936 N_A_1924_48#_c_1327_n N_A_1762_74#_c_1568_n 0.00923271f $X=11.395
+ $Y=1.385 $X2=0 $Y2=0
cc_937 N_A_1924_48#_c_1337_n N_A_1762_74#_c_1568_n 0.0088719f $X=12.065 $Y=2.265
+ $X2=0 $Y2=0
cc_938 N_A_1924_48#_c_1338_n N_A_1762_74#_c_1568_n 0.0179959f $X=11.75 $Y=2.265
+ $X2=0 $Y2=0
cc_939 N_A_1924_48#_c_1328_n N_A_1762_74#_c_1568_n 0.0253686f $X=12.15 $Y=2.18
+ $X2=0 $Y2=0
cc_940 N_A_1924_48#_c_1321_n N_A_1762_74#_c_1468_n 0.00300533f $X=9.785 $Y=0.865
+ $X2=0 $Y2=0
cc_941 N_A_1924_48#_c_1367_n N_A_1762_74#_c_1468_n 0.0189516f $X=9.785 $Y=0.985
+ $X2=0 $Y2=0
cc_942 N_A_1924_48#_c_1319_n N_A_1762_74#_c_1484_n 2.73249e-19 $X=9.955 $Y=2.165
+ $X2=0 $Y2=0
cc_943 N_A_1924_48#_c_1319_n N_A_1762_74#_c_1469_n 0.00185112f $X=9.955 $Y=2.165
+ $X2=0 $Y2=0
cc_944 N_A_1924_48#_c_1329_n N_A_1762_74#_c_1469_n 0.00300533f $X=9.785 $Y=1.065
+ $X2=0 $Y2=0
cc_945 N_A_1924_48#_c_1319_n N_A_1762_74#_c_1486_n 0.0059349f $X=9.955 $Y=2.165
+ $X2=0 $Y2=0
cc_946 N_A_1924_48#_c_1332_n N_A_1762_74#_c_1486_n 0.00552372f $X=10.35 $Y=2.24
+ $X2=0 $Y2=0
cc_947 N_A_1924_48#_c_1333_n N_A_1762_74#_c_1486_n 0.00239652f $X=10.03 $Y=2.24
+ $X2=0 $Y2=0
cc_948 N_A_1924_48#_c_1336_n N_A_1762_74#_c_1488_n 0.0422694f $X=11.665 $Y=2.75
+ $X2=0 $Y2=0
cc_949 N_A_1924_48#_c_1337_n N_VPWR_M1032_d 0.0043753f $X=12.065 $Y=2.265 $X2=0
+ $Y2=0
cc_950 N_A_1924_48#_c_1328_n N_VPWR_M1032_d 0.00765109f $X=12.15 $Y=2.18 $X2=0
+ $Y2=0
cc_951 N_A_1924_48#_c_1334_n N_VPWR_c_1702_n 0.00281001f $X=10.44 $Y=2.465 $X2=0
+ $Y2=0
cc_952 N_A_1924_48#_c_1336_n N_VPWR_c_1703_n 0.0309026f $X=11.665 $Y=2.75 $X2=0
+ $Y2=0
cc_953 N_A_1924_48#_c_1337_n N_VPWR_c_1703_n 0.0246255f $X=12.065 $Y=2.265 $X2=0
+ $Y2=0
cc_954 N_A_1924_48#_c_1334_n N_VPWR_c_1709_n 0.0044313f $X=10.44 $Y=2.465 $X2=0
+ $Y2=0
cc_955 N_A_1924_48#_c_1336_n N_VPWR_c_1713_n 0.011066f $X=11.665 $Y=2.75 $X2=0
+ $Y2=0
cc_956 N_A_1924_48#_c_1334_n N_VPWR_c_1695_n 0.00858246f $X=10.44 $Y=2.465 $X2=0
+ $Y2=0
cc_957 N_A_1924_48#_c_1335_n N_VPWR_c_1695_n 3.30814e-19 $X=10.44 $Y=2.24 $X2=0
+ $Y2=0
cc_958 N_A_1924_48#_c_1336_n N_VPWR_c_1695_n 0.00915947f $X=11.665 $Y=2.75 $X2=0
+ $Y2=0
cc_959 N_A_1924_48#_c_1333_n N_A_1600_347#_c_1984_n 7.2682e-19 $X=10.03 $Y=2.24
+ $X2=0 $Y2=0
cc_960 N_A_1924_48#_c_1334_n N_A_1600_347#_c_1984_n 0.0017475f $X=10.44 $Y=2.465
+ $X2=0 $Y2=0
cc_961 N_A_1924_48#_c_1335_n N_A_1600_347#_c_1984_n 0.00380271f $X=10.44 $Y=2.24
+ $X2=0 $Y2=0
cc_962 N_A_1924_48#_c_1333_n N_A_1712_374#_c_2018_n 0.00406826f $X=10.03 $Y=2.24
+ $X2=0 $Y2=0
cc_963 N_A_1924_48#_c_1334_n N_A_1712_374#_c_2018_n 0.00494591f $X=10.44
+ $Y=2.465 $X2=0 $Y2=0
cc_964 N_A_1924_48#_c_1332_n N_A_1712_374#_c_2019_n 0.00603289f $X=10.35 $Y=2.24
+ $X2=0 $Y2=0
cc_965 N_A_1924_48#_c_1334_n N_A_1712_374#_c_2019_n 0.00486225f $X=10.44
+ $Y=2.465 $X2=0 $Y2=0
cc_966 N_A_1924_48#_c_1335_n N_A_1712_374#_c_2019_n 4.15671e-19 $X=10.44 $Y=2.24
+ $X2=0 $Y2=0
cc_967 N_A_1924_48#_c_1337_n N_Q_N_c_2056_n 0.0115069f $X=12.065 $Y=2.265 $X2=0
+ $Y2=0
cc_968 N_A_1924_48#_c_1326_n N_Q_N_c_2052_n 0.0121685f $X=12.065 $Y=1.385 $X2=0
+ $Y2=0
cc_969 N_A_1924_48#_c_1328_n N_Q_N_c_2052_n 0.0426163f $X=12.15 $Y=2.18 $X2=0
+ $Y2=0
cc_970 N_A_1924_48#_c_1326_n Q_N 0.00999592f $X=12.065 $Y=1.385 $X2=0 $Y2=0
cc_971 N_A_1924_48#_c_1324_n N_VGND_c_2105_n 0.0370462f $X=11.23 $Y=0.58 $X2=0
+ $Y2=0
cc_972 N_A_1924_48#_c_1325_n N_VGND_c_2105_n 0.00382008f $X=11.31 $Y=1.3 $X2=0
+ $Y2=0
cc_973 N_A_1924_48#_c_1326_n N_VGND_c_2105_n 0.0277028f $X=12.065 $Y=1.385 $X2=0
+ $Y2=0
cc_974 N_A_1924_48#_c_1330_n N_VGND_c_2105_n 0.0121589f $X=11.23 $Y=0.985 $X2=0
+ $Y2=0
cc_975 N_A_1924_48#_c_1321_n N_VGND_c_2113_n 0.00461464f $X=9.785 $Y=0.865 $X2=0
+ $Y2=0
cc_976 N_A_1924_48#_c_1324_n N_VGND_c_2114_n 0.0145931f $X=11.23 $Y=0.58 $X2=0
+ $Y2=0
cc_977 N_A_1924_48#_c_1320_n N_VGND_c_2117_n 0.00441445f $X=9.785 $Y=1.03 $X2=0
+ $Y2=0
cc_978 N_A_1924_48#_c_1321_n N_VGND_c_2117_n 0.00910057f $X=9.785 $Y=0.865 $X2=0
+ $Y2=0
cc_979 N_A_1924_48#_c_1324_n N_VGND_c_2117_n 0.0120099f $X=11.23 $Y=0.58 $X2=0
+ $Y2=0
cc_980 N_A_1924_48#_c_1321_n N_VGND_c_2122_n 0.00203578f $X=9.785 $Y=0.865 $X2=0
+ $Y2=0
cc_981 N_A_1924_48#_c_1323_n N_VGND_c_2122_n 0.0374282f $X=11.065 $Y=0.985 $X2=0
+ $Y2=0
cc_982 N_A_1924_48#_c_1324_n N_VGND_c_2122_n 0.0132497f $X=11.23 $Y=0.58 $X2=0
+ $Y2=0
cc_983 N_A_1762_74#_c_1476_n N_A_2556_112#_c_1654_n 0.0189684f $X=13.395 $Y=1.94
+ $X2=0 $Y2=0
cc_984 N_A_1762_74#_c_1466_n N_A_2556_112#_c_1654_n 0.00570196f $X=13.14 $Y=1.79
+ $X2=0 $Y2=0
cc_985 N_A_1762_74#_M1016_g N_A_2556_112#_c_1649_n 0.0212903f $X=13.14 $Y=0.835
+ $X2=0 $Y2=0
cc_986 N_A_1762_74#_c_1466_n N_A_2556_112#_c_1649_n 0.00163137f $X=13.14 $Y=1.79
+ $X2=0 $Y2=0
cc_987 N_A_1762_74#_M1016_g N_A_2556_112#_c_1650_n 0.0093401f $X=13.14 $Y=0.835
+ $X2=0 $Y2=0
cc_988 N_A_1762_74#_M1005_g N_A_2556_112#_c_1651_n 9.40127e-19 $X=12.075 $Y=0.74
+ $X2=0 $Y2=0
cc_989 N_A_1762_74#_c_1460_n N_A_2556_112#_c_1651_n 0.00388219f $X=13.065
+ $Y=1.69 $X2=0 $Y2=0
cc_990 N_A_1762_74#_M1016_g N_A_2556_112#_c_1651_n 0.0367305f $X=13.14 $Y=0.835
+ $X2=0 $Y2=0
cc_991 N_A_1762_74#_c_1474_n N_A_2556_112#_c_1652_n 0.0024952f $X=12.395
+ $Y=1.765 $X2=0 $Y2=0
cc_992 N_A_1762_74#_c_1460_n N_A_2556_112#_c_1652_n 0.00554698f $X=13.065
+ $Y=1.69 $X2=0 $Y2=0
cc_993 N_A_1762_74#_M1016_g N_A_2556_112#_c_1652_n 0.00246233f $X=13.14 $Y=0.835
+ $X2=0 $Y2=0
cc_994 N_A_1762_74#_c_1476_n N_A_2556_112#_c_1652_n 0.00901458f $X=13.395
+ $Y=1.94 $X2=0 $Y2=0
cc_995 N_A_1762_74#_c_1466_n N_A_2556_112#_c_1652_n 0.0170873f $X=13.14 $Y=1.79
+ $X2=0 $Y2=0
cc_996 N_A_1762_74#_c_1466_n N_A_2556_112#_c_1653_n 0.00790181f $X=13.14 $Y=1.79
+ $X2=0 $Y2=0
cc_997 N_A_1762_74#_c_1482_n N_VPWR_c_1702_n 0.0106837f $X=11.11 $Y=2.18 $X2=0
+ $Y2=0
cc_998 N_A_1762_74#_c_1487_n N_VPWR_c_1702_n 0.0300176f $X=11.115 $Y=2.75 $X2=0
+ $Y2=0
cc_999 N_A_1762_74#_c_1471_n N_VPWR_c_1703_n 0.0126536f $X=11.89 $Y=2.465 $X2=0
+ $Y2=0
cc_1000 N_A_1762_74#_c_1474_n N_VPWR_c_1703_n 0.00563594f $X=12.395 $Y=1.765
+ $X2=0 $Y2=0
cc_1001 N_A_1762_74#_c_1476_n N_VPWR_c_1704_n 0.0184604f $X=13.395 $Y=1.94 $X2=0
+ $Y2=0
cc_1002 N_A_1762_74#_c_1466_n N_VPWR_c_1704_n 4.22058e-19 $X=13.14 $Y=1.79 $X2=0
+ $Y2=0
cc_1003 N_A_1762_74#_c_1471_n N_VPWR_c_1713_n 0.00413917f $X=11.89 $Y=2.465
+ $X2=0 $Y2=0
cc_1004 N_A_1762_74#_c_1487_n N_VPWR_c_1713_n 0.0143991f $X=11.115 $Y=2.75 $X2=0
+ $Y2=0
cc_1005 N_A_1762_74#_c_1474_n N_VPWR_c_1714_n 0.00439937f $X=12.395 $Y=1.765
+ $X2=0 $Y2=0
cc_1006 N_A_1762_74#_c_1476_n N_VPWR_c_1714_n 0.00452264f $X=13.395 $Y=1.94
+ $X2=0 $Y2=0
cc_1007 N_A_1762_74#_c_1471_n N_VPWR_c_1695_n 0.00860356f $X=11.89 $Y=2.465
+ $X2=0 $Y2=0
cc_1008 N_A_1762_74#_c_1474_n N_VPWR_c_1695_n 0.00843992f $X=12.395 $Y=1.765
+ $X2=0 $Y2=0
cc_1009 N_A_1762_74#_c_1476_n N_VPWR_c_1695_n 0.00465044f $X=13.395 $Y=1.94
+ $X2=0 $Y2=0
cc_1010 N_A_1762_74#_c_1487_n N_VPWR_c_1695_n 0.0119711f $X=11.115 $Y=2.75 $X2=0
+ $Y2=0
cc_1011 N_A_1762_74#_c_1481_n N_A_1600_347#_M1009_d 0.00446377f $X=10 $Y=2.035
+ $X2=0 $Y2=0
cc_1012 N_A_1762_74#_M1035_d N_A_1600_347#_c_1982_n 0.00516465f $X=8.975 $Y=1.87
+ $X2=0 $Y2=0
cc_1013 N_A_1762_74#_c_1481_n N_A_1600_347#_c_1982_n 0.00723674f $X=10 $Y=2.035
+ $X2=0 $Y2=0
cc_1014 N_A_1762_74#_c_1484_n N_A_1600_347#_c_1982_n 0.0212063f $X=9.21 $Y=2.015
+ $X2=0 $Y2=0
cc_1015 N_A_1762_74#_c_1481_n N_A_1600_347#_c_1984_n 0.0189117f $X=10 $Y=2.035
+ $X2=0 $Y2=0
cc_1016 N_A_1762_74#_c_1486_n N_A_1712_374#_c_2018_n 0.00131213f $X=10.085
+ $Y=2.035 $X2=0 $Y2=0
cc_1017 N_A_1762_74#_c_1482_n N_A_1712_374#_c_2019_n 0.0121645f $X=11.11 $Y=2.18
+ $X2=0 $Y2=0
cc_1018 N_A_1762_74#_c_1486_n N_A_1712_374#_c_2019_n 0.00723033f $X=10.085
+ $Y=2.035 $X2=0 $Y2=0
cc_1019 N_A_1762_74#_c_1474_n N_Q_N_c_2055_n 0.0016734f $X=12.395 $Y=1.765 $X2=0
+ $Y2=0
cc_1020 N_A_1762_74#_c_1460_n N_Q_N_c_2055_n 0.00391459f $X=13.065 $Y=1.69 $X2=0
+ $Y2=0
cc_1021 N_A_1762_74#_c_1476_n N_Q_N_c_2055_n 0.00408934f $X=13.395 $Y=1.94 $X2=0
+ $Y2=0
cc_1022 N_A_1762_74#_c_1466_n N_Q_N_c_2055_n 4.54538e-19 $X=13.14 $Y=1.79 $X2=0
+ $Y2=0
cc_1023 N_A_1762_74#_c_1470_n N_Q_N_c_2056_n 7.36264e-19 $X=11.89 $Y=2.375 $X2=0
+ $Y2=0
cc_1024 N_A_1762_74#_c_1471_n N_Q_N_c_2056_n 3.94152e-19 $X=11.89 $Y=2.465 $X2=0
+ $Y2=0
cc_1025 N_A_1762_74#_c_1474_n N_Q_N_c_2056_n 0.0135312f $X=12.395 $Y=1.765 $X2=0
+ $Y2=0
cc_1026 N_A_1762_74#_M1005_g N_Q_N_c_2052_n 0.00681469f $X=12.075 $Y=0.74 $X2=0
+ $Y2=0
cc_1027 N_A_1762_74#_c_1474_n N_Q_N_c_2052_n 0.00126633f $X=12.395 $Y=1.765
+ $X2=0 $Y2=0
cc_1028 N_A_1762_74#_c_1460_n N_Q_N_c_2052_n 0.0124346f $X=13.065 $Y=1.69 $X2=0
+ $Y2=0
cc_1029 N_A_1762_74#_c_1465_n N_Q_N_c_2052_n 0.00306915f $X=12.395 $Y=1.69 $X2=0
+ $Y2=0
cc_1030 N_A_1762_74#_M1005_g Q_N 0.00766778f $X=12.075 $Y=0.74 $X2=0 $Y2=0
cc_1031 N_A_1762_74#_M1016_g Q_N 0.00756882f $X=13.14 $Y=0.835 $X2=0 $Y2=0
cc_1032 N_A_1762_74#_M1005_g Q_N 0.0034024f $X=12.075 $Y=0.74 $X2=0 $Y2=0
cc_1033 N_A_1762_74#_c_1458_n Q_N 0.00728143f $X=12.32 $Y=1.69 $X2=0 $Y2=0
cc_1034 N_A_1762_74#_c_1476_n Q 6.21038e-19 $X=13.395 $Y=1.94 $X2=0 $Y2=0
cc_1035 N_A_1762_74#_c_1466_n Q 7.9726e-19 $X=13.14 $Y=1.79 $X2=0 $Y2=0
cc_1036 N_A_1762_74#_c_1455_n N_VGND_c_2105_n 0.00389959f $X=11.015 $Y=0.865
+ $X2=0 $Y2=0
cc_1037 N_A_1762_74#_M1005_g N_VGND_c_2105_n 0.0169409f $X=12.075 $Y=0.74 $X2=0
+ $Y2=0
cc_1038 N_A_1762_74#_c_1462_n N_VGND_c_2105_n 0.00114561f $X=11.3 $Y=0.94 $X2=0
+ $Y2=0
cc_1039 N_A_1762_74#_M1016_g N_VGND_c_2106_n 0.0047492f $X=13.14 $Y=0.835 $X2=0
+ $Y2=0
cc_1040 N_A_1762_74#_c_1468_n N_VGND_c_2113_n 0.025983f $X=9.09 $Y=0.515 $X2=0
+ $Y2=0
cc_1041 N_A_1762_74#_c_1455_n N_VGND_c_2114_n 0.00434272f $X=11.015 $Y=0.865
+ $X2=0 $Y2=0
cc_1042 N_A_1762_74#_M1005_g N_VGND_c_2115_n 0.00434272f $X=12.075 $Y=0.74 $X2=0
+ $Y2=0
cc_1043 N_A_1762_74#_M1016_g N_VGND_c_2115_n 0.00340575f $X=13.14 $Y=0.835 $X2=0
+ $Y2=0
cc_1044 N_A_1762_74#_c_1455_n N_VGND_c_2117_n 0.00827575f $X=11.015 $Y=0.865
+ $X2=0 $Y2=0
cc_1045 N_A_1762_74#_M1005_g N_VGND_c_2117_n 0.00830058f $X=12.075 $Y=0.74 $X2=0
+ $Y2=0
cc_1046 N_A_1762_74#_M1016_g N_VGND_c_2117_n 0.00487769f $X=13.14 $Y=0.835 $X2=0
+ $Y2=0
cc_1047 N_A_1762_74#_c_1468_n N_VGND_c_2117_n 0.0210826f $X=9.09 $Y=0.515 $X2=0
+ $Y2=0
cc_1048 N_A_1762_74#_c_1468_n N_VGND_c_2121_n 0.0134766f $X=9.09 $Y=0.515 $X2=0
+ $Y2=0
cc_1049 N_A_1762_74#_c_1455_n N_VGND_c_2122_n 0.00405065f $X=11.015 $Y=0.865
+ $X2=0 $Y2=0
cc_1050 N_A_2556_112#_c_1654_n N_VPWR_c_1704_n 0.00991033f $X=13.9 $Y=1.765
+ $X2=0 $Y2=0
cc_1051 N_A_2556_112#_c_1649_n N_VPWR_c_1704_n 0.00583793f $X=13.81 $Y=1.385
+ $X2=0 $Y2=0
cc_1052 N_A_2556_112#_c_1652_n N_VPWR_c_1704_n 0.059064f $X=13.17 $Y=2.16 $X2=0
+ $Y2=0
cc_1053 N_A_2556_112#_c_1653_n N_VPWR_c_1704_n 0.012653f $X=13.62 $Y=1.385 $X2=0
+ $Y2=0
cc_1054 N_A_2556_112#_c_1652_n N_VPWR_c_1714_n 0.00775887f $X=13.17 $Y=2.16
+ $X2=0 $Y2=0
cc_1055 N_A_2556_112#_c_1654_n N_VPWR_c_1715_n 0.00439937f $X=13.9 $Y=1.765
+ $X2=0 $Y2=0
cc_1056 N_A_2556_112#_c_1654_n N_VPWR_c_1695_n 0.00846965f $X=13.9 $Y=1.765
+ $X2=0 $Y2=0
cc_1057 N_A_2556_112#_c_1652_n N_VPWR_c_1695_n 0.00855956f $X=13.17 $Y=2.16
+ $X2=0 $Y2=0
cc_1058 N_A_2556_112#_c_1652_n N_Q_N_c_2055_n 0.0552255f $X=13.17 $Y=2.16 $X2=0
+ $Y2=0
cc_1059 N_A_2556_112#_c_1651_n N_Q_N_c_2052_n 0.0197595f $X=13.13 $Y=1.55 $X2=0
+ $Y2=0
cc_1060 N_A_2556_112#_c_1652_n N_Q_N_c_2052_n 0.0106741f $X=13.17 $Y=2.16 $X2=0
+ $Y2=0
cc_1061 N_A_2556_112#_c_1651_n Q_N 0.0422235f $X=13.13 $Y=1.55 $X2=0 $Y2=0
cc_1062 N_A_2556_112#_c_1654_n Q 0.0177247f $X=13.9 $Y=1.765 $X2=0 $Y2=0
cc_1063 N_A_2556_112#_c_1649_n Q 0.0268637f $X=13.81 $Y=1.385 $X2=0 $Y2=0
cc_1064 N_A_2556_112#_c_1650_n Q 0.0188373f $X=13.9 $Y=1.22 $X2=0 $Y2=0
cc_1065 N_A_2556_112#_c_1653_n Q 0.026211f $X=13.62 $Y=1.385 $X2=0 $Y2=0
cc_1066 N_A_2556_112#_c_1649_n N_VGND_c_2106_n 0.00760746f $X=13.81 $Y=1.385
+ $X2=0 $Y2=0
cc_1067 N_A_2556_112#_c_1650_n N_VGND_c_2106_n 0.0113395f $X=13.9 $Y=1.22 $X2=0
+ $Y2=0
cc_1068 N_A_2556_112#_c_1651_n N_VGND_c_2106_n 0.0189646f $X=13.13 $Y=1.55 $X2=0
+ $Y2=0
cc_1069 N_A_2556_112#_c_1653_n N_VGND_c_2106_n 0.0265928f $X=13.62 $Y=1.385
+ $X2=0 $Y2=0
cc_1070 N_A_2556_112#_c_1651_n N_VGND_c_2115_n 0.0099752f $X=13.13 $Y=1.55 $X2=0
+ $Y2=0
cc_1071 N_A_2556_112#_c_1650_n N_VGND_c_2116_n 0.00434272f $X=13.9 $Y=1.22 $X2=0
+ $Y2=0
cc_1072 N_A_2556_112#_c_1650_n N_VGND_c_2117_n 0.00828717f $X=13.9 $Y=1.22 $X2=0
+ $Y2=0
cc_1073 N_A_2556_112#_c_1651_n N_VGND_c_2117_n 0.0132953f $X=13.13 $Y=1.55 $X2=0
+ $Y2=0
cc_1074 N_VPWR_c_1696_n N_A_290_464#_c_1869_n 0.0100039f $X=0.73 $Y=2.805 $X2=0
+ $Y2=0
cc_1075 N_VPWR_c_1712_n N_A_290_464#_c_1869_n 0.0174287f $X=2.555 $Y=3.33 $X2=0
+ $Y2=0
cc_1076 N_VPWR_c_1695_n N_A_290_464#_c_1869_n 0.0179948f $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_1077 N_VPWR_c_1712_n N_A_290_464#_c_1872_n 0.00879349f $X=2.555 $Y=3.33 $X2=0
+ $Y2=0
cc_1078 N_VPWR_c_1695_n N_A_290_464#_c_1872_n 0.0130676f $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_1079 N_VPWR_M1031_d N_A_290_464#_c_1863_n 0.00658019f $X=2.5 $Y=2.32 $X2=0
+ $Y2=0
cc_1080 N_VPWR_c_1697_n N_A_290_464#_c_1863_n 0.0208489f $X=2.655 $Y=2.825 $X2=0
+ $Y2=0
cc_1081 N_VPWR_c_1699_n N_A_290_464#_c_1863_n 0.00100103f $X=3.74 $Y=2.78 $X2=0
+ $Y2=0
cc_1082 N_VPWR_c_1695_n N_A_290_464#_c_1863_n 0.0312535f $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_1083 N_VPWR_M1019_d N_A_290_464#_c_1864_n 0.00137078f $X=3.59 $Y=1.84 $X2=0
+ $Y2=0
cc_1084 N_VPWR_c_1699_n N_A_290_464#_c_1864_n 0.00282404f $X=3.74 $Y=2.78 $X2=0
+ $Y2=0
cc_1085 N_VPWR_M1019_d N_A_290_464#_c_1950_n 0.00497294f $X=3.59 $Y=1.84 $X2=0
+ $Y2=0
cc_1086 N_VPWR_c_1699_n N_A_290_464#_c_1950_n 0.0121566f $X=3.74 $Y=2.78 $X2=0
+ $Y2=0
cc_1087 N_VPWR_c_1695_n N_A_290_464#_c_1950_n 5.62582e-19 $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_1088 N_VPWR_c_1695_n N_A_1600_347#_c_1982_n 0.00950249f $X=14.16 $Y=3.33
+ $X2=0 $Y2=0
cc_1089 N_VPWR_c_1701_n N_A_1600_347#_c_1983_n 0.0299903f $X=7.7 $Y=2.525 $X2=0
+ $Y2=0
cc_1090 N_VPWR_c_1709_n N_A_1600_347#_c_1983_n 0.0073103f $X=10.58 $Y=3.33 $X2=0
+ $Y2=0
cc_1091 N_VPWR_c_1695_n N_A_1600_347#_c_1983_n 0.00891228f $X=14.16 $Y=3.33
+ $X2=0 $Y2=0
cc_1092 N_VPWR_c_1702_n N_A_1712_374#_c_2018_n 0.0119328f $X=10.665 $Y=2.75
+ $X2=0 $Y2=0
cc_1093 N_VPWR_c_1709_n N_A_1712_374#_c_2018_n 0.0993421f $X=10.58 $Y=3.33 $X2=0
+ $Y2=0
cc_1094 N_VPWR_c_1695_n N_A_1712_374#_c_2018_n 0.0546301f $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_1095 N_VPWR_c_1702_n N_A_1712_374#_c_2019_n 0.0250721f $X=10.665 $Y=2.75
+ $X2=0 $Y2=0
cc_1096 N_VPWR_c_1709_n N_A_1712_374#_c_2020_n 0.0214714f $X=10.58 $Y=3.33 $X2=0
+ $Y2=0
cc_1097 N_VPWR_c_1695_n N_A_1712_374#_c_2020_n 0.0110721f $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_1098 N_VPWR_c_1703_n N_Q_N_c_2056_n 0.0173822f $X=12.115 $Y=2.75 $X2=0 $Y2=0
cc_1099 N_VPWR_c_1714_n N_Q_N_c_2056_n 0.0112323f $X=13.455 $Y=3.33 $X2=0 $Y2=0
cc_1100 N_VPWR_c_1695_n N_Q_N_c_2056_n 0.00925249f $X=14.16 $Y=3.33 $X2=0 $Y2=0
cc_1101 N_VPWR_c_1704_n Q 0.0378352f $X=13.62 $Y=2.16 $X2=0 $Y2=0
cc_1102 N_VPWR_c_1715_n Q 0.014802f $X=14.16 $Y=3.33 $X2=0 $Y2=0
cc_1103 N_VPWR_c_1695_n Q 0.0122072f $X=14.16 $Y=3.33 $X2=0 $Y2=0
cc_1104 N_A_290_464#_c_1872_n A_416_464# 0.00535326f $X=2.215 $Y=2.715 $X2=-0.19
+ $Y2=-0.245
cc_1105 N_A_290_464#_c_1876_n A_416_464# 0.00156665f $X=2.3 $Y=2.63 $X2=-0.19
+ $Y2=-0.245
cc_1106 N_A_290_464#_c_1879_n A_416_464# 0.00160617f $X=2.3 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_1107 N_A_290_464#_c_1856_n N_VGND_c_2101_n 0.00639088f $X=1.67 $Y=0.58 $X2=0
+ $Y2=0
cc_1108 N_A_290_464#_c_1856_n N_VGND_c_2102_n 0.0126723f $X=1.67 $Y=0.58 $X2=0
+ $Y2=0
cc_1109 N_A_290_464#_c_1857_n N_VGND_c_2102_n 0.00351301f $X=2.215 $Y=1.005
+ $X2=0 $Y2=0
cc_1110 N_A_290_464#_c_1856_n N_VGND_c_2107_n 0.0144922f $X=1.67 $Y=0.58 $X2=0
+ $Y2=0
cc_1111 N_A_290_464#_c_1856_n N_VGND_c_2117_n 0.0118826f $X=1.67 $Y=0.58 $X2=0
+ $Y2=0
cc_1112 N_A_1600_347#_c_1982_n N_A_1712_374#_M1035_s 0.00393221f $X=9.58
+ $Y=2.435 $X2=-0.19 $Y2=1.66
cc_1113 N_A_1600_347#_c_1982_n N_A_1712_374#_c_2018_n 0.023515f $X=9.58 $Y=2.435
+ $X2=0 $Y2=0
cc_1114 N_A_1600_347#_c_1984_n N_A_1712_374#_c_2018_n 0.0186414f $X=9.665
+ $Y=2.51 $X2=0 $Y2=0
cc_1115 N_A_1600_347#_c_1984_n N_A_1712_374#_c_2019_n 0.0146404f $X=9.665
+ $Y=2.51 $X2=0 $Y2=0
cc_1116 N_A_1600_347#_c_1982_n N_A_1712_374#_c_2020_n 0.0253438f $X=9.58
+ $Y=2.435 $X2=0 $Y2=0
cc_1117 N_A_1600_347#_c_1983_n N_A_1712_374#_c_2020_n 0.0045919f $X=8.15
+ $Y=2.435 $X2=0 $Y2=0
cc_1118 Q_N N_VGND_c_2105_n 0.0326809f $X=12.155 $Y=0.47 $X2=0 $Y2=0
cc_1119 Q_N N_VGND_c_2115_n 0.0219264f $X=12.155 $Y=0.47 $X2=0 $Y2=0
cc_1120 Q_N N_VGND_c_2117_n 0.0180924f $X=12.155 $Y=0.47 $X2=0 $Y2=0
cc_1121 Q N_VGND_c_2106_n 0.0271167f $X=14.075 $Y=0.47 $X2=0 $Y2=0
cc_1122 Q N_VGND_c_2116_n 0.014787f $X=14.075 $Y=0.47 $X2=0 $Y2=0
cc_1123 Q N_VGND_c_2117_n 0.012183f $X=14.075 $Y=0.47 $X2=0 $Y2=0
