* File: sky130_fd_sc_ls__dlxbp_1.pex.spice
* Created: Wed Sep  2 11:04:33 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__DLXBP_1%D 2 5 6 8 9 12 14
c40 2 0 1.56139e-19 $X=0.587 $Y=1.713
r41 12 14 46.504 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=0.587 $Y=1.385
+ $X2=0.587 $Y2=1.22
r42 12 13 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.6
+ $Y=1.385 $X2=0.6 $Y2=1.385
r43 9 13 2.14223 $w=6.68e-07 $l=1.2e-07 $layer=LI1_cond $X=0.72 $Y=1.555 $X2=0.6
+ $Y2=1.555
r44 6 8 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.5 $Y=1.99 $X2=0.5
+ $Y2=2.485
r45 5 14 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=0.5 $Y=0.835 $X2=0.5
+ $Y2=1.22
r46 2 6 45.8811 $w=2.91e-07 $l=3.17534e-07 $layer=POLY_cond $X=0.587 $Y=1.713
+ $X2=0.5 $Y2=1.99
r47 1 12 1.95057 $w=3.55e-07 $l=1.2e-08 $layer=POLY_cond $X=0.587 $Y=1.397
+ $X2=0.587 $Y2=1.385
r48 1 2 51.3649 $w=3.55e-07 $l=3.16e-07 $layer=POLY_cond $X=0.587 $Y=1.397
+ $X2=0.587 $Y2=1.713
.ends

.subckt PM_SKY130_FD_SC_LS__DLXBP_1%GATE 3 5 6 8 9 12 14
c40 14 0 3.53875e-20 $X=1.17 $Y=1.22
c41 9 0 7.84293e-20 $X=1.2 $Y=1.295
r42 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.17 $Y=1.385
+ $X2=1.17 $Y2=1.55
r43 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.17 $Y=1.385
+ $X2=1.17 $Y2=1.22
r44 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.17
+ $Y=1.385 $X2=1.17 $Y2=1.385
r45 9 13 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=1.17 $Y=1.295 $X2=1.17
+ $Y2=1.385
r46 6 8 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.11 $Y=1.99 $X2=1.11
+ $Y2=2.485
r47 5 6 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.11 $Y=1.9 $X2=1.11
+ $Y2=1.99
r48 5 15 136.048 $w=1.8e-07 $l=3.5e-07 $layer=POLY_cond $X=1.11 $Y=1.9 $X2=1.11
+ $Y2=1.55
r49 3 14 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.08 $Y=0.74 $X2=1.08
+ $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_LS__DLXBP_1%A_231_74# 1 2 11 13 15 16 18 19 20 24 27 30
+ 31 33 35 36 38 40 41 44
c134 40 0 6.89381e-20 $X=3.91 $Y=0.345
c135 36 0 7.84293e-20 $X=2.165 $Y=1.635
c136 33 0 1.56139e-19 $X=1.675 $Y=1.68
c137 31 0 3.53875e-20 $X=2.91 $Y=0.665
c138 20 0 1.74828e-19 $X=3.335 $Y=1.765
c139 19 0 1.49705e-19 $X=3.925 $Y=1.765
c140 16 0 3.19065e-19 $X=3.245 $Y=1.885
r141 48 49 14.1693 $w=2.54e-07 $l=2.95e-07 $layer=LI1_cond $X=1.295 $Y=1.72
+ $X2=1.59 $Y2=1.72
r142 46 47 13.7503 $w=5.43e-07 $l=3.45e-07 $layer=LI1_cond $X=1.402 $Y=0.665
+ $X2=1.402 $Y2=1.01
r143 44 46 3.18223 $w=5.43e-07 $l=1.45e-07 $layer=LI1_cond $X=1.402 $Y=0.52
+ $X2=1.402 $Y2=0.665
r144 41 57 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.91 $Y=0.345
+ $X2=3.91 $Y2=0.51
r145 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.91
+ $Y=0.345 $X2=3.91 $Y2=0.345
r146 38 52 18.4631 $w=1.68e-07 $l=2.83e-07 $layer=LI1_cond $X=2.995 $Y=0.382
+ $X2=2.995 $Y2=0.665
r147 38 40 37.5109 $w=2.53e-07 $l=8.3e-07 $layer=LI1_cond $X=3.08 $Y=0.382
+ $X2=3.91 $Y2=0.382
r148 35 36 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.165
+ $Y=1.635 $X2=2.165 $Y2=1.635
r149 33 49 4.36065 $w=4.2e-07 $l=1.03078e-07 $layer=LI1_cond $X=1.675 $Y=1.68
+ $X2=1.59 $Y2=1.72
r150 33 35 13.4452 $w=4.18e-07 $l=4.9e-07 $layer=LI1_cond $X=1.675 $Y=1.68
+ $X2=2.165 $Y2=1.68
r151 32 46 7.70116 $w=1.7e-07 $l=2.73e-07 $layer=LI1_cond $X=1.675 $Y=0.665
+ $X2=1.402 $Y2=0.665
r152 31 52 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.91 $Y=0.665
+ $X2=2.995 $Y2=0.665
r153 31 32 80.5722 $w=1.68e-07 $l=1.235e-06 $layer=LI1_cond $X=2.91 $Y=0.665
+ $X2=1.675 $Y2=0.665
r154 30 49 3.08766 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=1.59 $Y=1.47
+ $X2=1.59 $Y2=1.72
r155 30 47 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=1.59 $Y=1.47
+ $X2=1.59 $Y2=1.01
r156 25 48 0.813113 $w=2.5e-07 $l=1.7e-07 $layer=LI1_cond $X=1.295 $Y=1.89
+ $X2=1.295 $Y2=1.72
r157 25 27 14.7513 $w=2.48e-07 $l=3.2e-07 $layer=LI1_cond $X=1.295 $Y=1.89
+ $X2=1.295 $Y2=2.21
r158 24 57 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4 $Y=0.83 $X2=4
+ $Y2=0.51
r159 22 24 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=4 $Y=1.69 $X2=4
+ $Y2=0.83
r160 19 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.925 $Y=1.765
+ $X2=4 $Y2=1.69
r161 19 20 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=3.925 $Y=1.765
+ $X2=3.335 $Y2=1.765
r162 16 20 26.9307 $w=1.5e-07 $l=1.58745e-07 $layer=POLY_cond $X=3.245 $Y=1.885
+ $X2=3.335 $Y2=1.765
r163 16 18 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.245 $Y=1.885
+ $X2=3.245 $Y2=2.46
r164 13 36 37.0704 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.24 $Y=1.885
+ $X2=2.24 $Y2=1.677
r165 13 15 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.24 $Y=1.885
+ $X2=2.24 $Y2=2.38
r166 9 36 37.0704 $w=1.5e-07 $l=2.14369e-07 $layer=POLY_cond $X=2.225 $Y=1.47
+ $X2=2.24 $Y2=1.677
r167 9 11 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.225 $Y=1.47
+ $X2=2.225 $Y2=0.78
r168 2 27 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.185
+ $Y=2.065 $X2=1.335 $Y2=2.21
r169 1 44 91 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=2 $X=1.155
+ $Y=0.37 $X2=1.295 $Y2=0.52
.ends

.subckt PM_SKY130_FD_SC_LS__DLXBP_1%A_27_413# 1 2 7 9 12 17 18 19 21 22 23 26 30
+ 34 35
c95 26 0 3.45399e-19 $X=2.71 $Y=1.635
c96 22 0 1.57288e-19 $X=2.545 $Y=2.145
r97 34 35 8.4794 $w=3.43e-07 $l=1.65e-07 $layer=LI1_cond $X=0.267 $Y=2.225
+ $X2=0.267 $Y2=2.06
r98 32 35 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=0.18 $Y=1.05
+ $X2=0.18 $Y2=2.06
r99 30 32 11.4207 $w=3.53e-07 $l=2.55e-07 $layer=LI1_cond $X=0.272 $Y=0.795
+ $X2=0.272 $Y2=1.05
r100 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.71
+ $Y=1.635 $X2=2.71 $Y2=1.635
r101 24 26 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=2.71 $Y=2.06
+ $X2=2.71 $Y2=1.635
r102 22 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.545 $Y=2.145
+ $X2=2.71 $Y2=2.06
r103 22 23 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=2.545 $Y=2.145
+ $X2=1.76 $Y2=2.145
r104 20 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.675 $Y=2.23
+ $X2=1.76 $Y2=2.145
r105 20 21 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.675 $Y=2.23
+ $X2=1.675 $Y2=2.545
r106 18 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.59 $Y=2.63
+ $X2=1.675 $Y2=2.545
r107 18 19 75.0267 $w=1.68e-07 $l=1.15e-06 $layer=LI1_cond $X=1.59 $Y=2.63
+ $X2=0.44 $Y2=2.63
r108 17 19 7.89393 $w=1.7e-07 $l=2.11268e-07 $layer=LI1_cond $X=0.267 $Y=2.545
+ $X2=0.44 $Y2=2.63
r109 16 34 0.233829 $w=3.43e-07 $l=7e-09 $layer=LI1_cond $X=0.267 $Y=2.232
+ $X2=0.267 $Y2=2.225
r110 16 17 10.4555 $w=3.43e-07 $l=3.13e-07 $layer=LI1_cond $X=0.267 $Y=2.232
+ $X2=0.267 $Y2=2.545
r111 10 27 38.832 $w=3.54e-07 $l=2.18746e-07 $layer=POLY_cond $X=2.87 $Y=1.47
+ $X2=2.745 $Y2=1.635
r112 10 12 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=2.87 $Y=1.47
+ $X2=2.87 $Y2=0.72
r113 7 27 50.4054 $w=3.54e-07 $l=3e-07 $layer=POLY_cond $X=2.855 $Y=1.885
+ $X2=2.745 $Y2=1.635
r114 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.855 $Y=1.885
+ $X2=2.855 $Y2=2.46
r115 2 34 300 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.065 $X2=0.275 $Y2=2.225
r116 1 30 182 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_NDIFF $count=1 $X=0.14
+ $Y=0.56 $X2=0.285 $Y2=0.795
.ends

.subckt PM_SKY130_FD_SC_LS__DLXBP_1%A_373_82# 1 2 9 10 12 13 15 18 19 23 27 31
+ 36 40 42 44
c114 40 0 8.79278e-21 $X=3.35 $Y=1.315
c115 36 0 1.49705e-19 $X=3.28 $Y=1.105
r116 40 44 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.35 $Y=1.315
+ $X2=3.35 $Y2=1.15
r117 39 41 9.33757 $w=4.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.28 $Y=1.315
+ $X2=3.28 $Y2=1.48
r118 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.35
+ $Y=1.315 $X2=3.35 $Y2=1.315
r119 36 39 5.34418 $w=4.68e-07 $l=2.1e-07 $layer=LI1_cond $X=3.28 $Y=1.105
+ $X2=3.28 $Y2=1.315
r120 31 34 3.91831 $w=2.48e-07 $l=8.5e-08 $layer=LI1_cond $X=2.055 $Y=2.525
+ $X2=2.055 $Y2=2.61
r121 27 29 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=2.01 $Y=1.005
+ $X2=2.01 $Y2=1.105
r122 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.935
+ $Y=2.215 $X2=3.935 $Y2=2.215
r123 21 23 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=3.935 $Y=2.44
+ $X2=3.935 $Y2=2.215
r124 20 42 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.215 $Y=2.525
+ $X2=3.13 $Y2=2.525
r125 19 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.77 $Y=2.525
+ $X2=3.935 $Y2=2.44
r126 19 20 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=3.77 $Y=2.525
+ $X2=3.215 $Y2=2.525
r127 18 42 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.13 $Y=2.44
+ $X2=3.13 $Y2=2.525
r128 18 41 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.13 $Y=2.44
+ $X2=3.13 $Y2=1.48
r129 16 31 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.18 $Y=2.525
+ $X2=2.055 $Y2=2.525
r130 15 42 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.045 $Y=2.525
+ $X2=3.13 $Y2=2.525
r131 15 16 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=3.045 $Y=2.525
+ $X2=2.18 $Y2=2.525
r132 14 29 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.175 $Y=1.105
+ $X2=2.01 $Y2=1.105
r133 13 36 6.76998 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=3.045 $Y=1.105
+ $X2=3.28 $Y2=1.105
r134 13 14 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=3.045 $Y=1.105
+ $X2=2.175 $Y2=1.105
r135 10 24 50.1894 $w=3.66e-07 $l=3.02903e-07 $layer=POLY_cond $X=3.775 $Y=2.465
+ $X2=3.892 $Y2=2.215
r136 10 12 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.775 $Y=2.465
+ $X2=3.775 $Y2=2.75
r137 9 44 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.26 $Y=0.72
+ $X2=3.26 $Y2=1.15
r138 2 34 600 $w=1.7e-07 $l=7.18853e-07 $layer=licon1_PDIFF $count=1 $X=1.87
+ $Y=1.96 $X2=2.015 $Y2=2.61
r139 1 27 182 $w=1.7e-07 $l=6.63551e-07 $layer=licon1_NDIFF $count=1 $X=1.865
+ $Y=0.41 $X2=2.01 $Y2=1.005
.ends

.subckt PM_SKY130_FD_SC_LS__DLXBP_1%A_863_98# 1 2 9 11 12 13 15 16 18 21 23 24
+ 25 27 30 33 38 45 48 52 55 57 62 65
c118 48 0 1.88618e-19 $X=5.29 $Y=1.32
c119 33 0 1.77373e-19 $X=6.065 $Y=1.485
c120 23 0 9.14246e-20 $X=6.66 $Y=1.65
c121 9 0 6.89381e-20 $X=4.39 $Y=0.83
r122 62 63 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.61
+ $Y=1.485 $X2=5.61 $Y2=1.485
r123 60 62 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=5.37 $Y=1.485
+ $X2=5.61 $Y2=1.485
r124 58 60 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=5.29 $Y=1.485 $X2=5.37
+ $Y2=1.485
r125 53 65 5.16603 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=5.37 $Y=2.32
+ $X2=5.37 $Y2=2.155
r126 53 55 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=5.37 $Y=2.32
+ $X2=5.37 $Y2=2.815
r127 50 65 5.16603 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=5.37 $Y=1.99
+ $X2=5.37 $Y2=2.155
r128 50 52 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=5.37 $Y=1.99
+ $X2=5.37 $Y2=1.985
r129 49 60 0.716491 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=5.37 $Y=1.65
+ $X2=5.37 $Y2=1.485
r130 49 52 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=5.37 $Y=1.65
+ $X2=5.37 $Y2=1.985
r131 48 58 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.29 $Y=1.32
+ $X2=5.29 $Y2=1.485
r132 48 57 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=5.29 $Y=1.32
+ $X2=5.29 $Y2=1.07
r133 43 57 8.88861 $w=3.53e-07 $l=1.77e-07 $layer=LI1_cond $X=5.197 $Y=0.893
+ $X2=5.197 $Y2=1.07
r134 43 45 12.2711 $w=3.53e-07 $l=3.78e-07 $layer=LI1_cond $X=5.197 $Y=0.893
+ $X2=5.197 $Y2=0.515
r135 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.48
+ $Y=2.155 $X2=4.48 $Y2=2.155
r136 38 65 1.34256 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=5.205 $Y=2.155
+ $X2=5.37 $Y2=2.155
r137 38 40 25.3188 $w=3.28e-07 $l=7.25e-07 $layer=LI1_cond $X=5.205 $Y=2.155
+ $X2=4.48 $Y2=2.155
r138 34 35 2.67778 $w=3.6e-07 $l=2e-08 $layer=POLY_cond $X=6.155 $Y=1.542
+ $X2=6.175 $Y2=1.542
r139 33 63 79.5619 $w=3.3e-07 $l=4.55e-07 $layer=POLY_cond $X=6.065 $Y=1.485
+ $X2=5.61 $Y2=1.485
r140 33 34 12.4725 $w=3.6e-07 $l=1.15022e-07 $layer=POLY_cond $X=6.065 $Y=1.485
+ $X2=6.155 $Y2=1.542
r141 28 37 23.3057 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=6.675 $Y=1.32
+ $X2=6.675 $Y2=1.542
r142 28 30 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.675 $Y=1.32
+ $X2=6.675 $Y2=0.855
r143 25 27 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=6.66 $Y=2.045
+ $X2=6.66 $Y2=2.54
r144 24 25 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.66 $Y=1.955
+ $X2=6.66 $Y2=2.045
r145 23 37 2.00833 $w=3.6e-07 $l=1.5e-08 $layer=POLY_cond $X=6.66 $Y=1.542
+ $X2=6.675 $Y2=1.542
r146 23 35 64.9361 $w=3.6e-07 $l=4.85e-07 $layer=POLY_cond $X=6.66 $Y=1.542
+ $X2=6.175 $Y2=1.542
r147 23 24 118.556 $w=1.8e-07 $l=3.05e-07 $layer=POLY_cond $X=6.66 $Y=1.65
+ $X2=6.66 $Y2=1.955
r148 19 35 23.3057 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=6.175 $Y=1.32
+ $X2=6.175 $Y2=1.542
r149 19 21 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=6.175 $Y=1.32
+ $X2=6.175 $Y2=0.76
r150 16 34 23.3057 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=6.155 $Y=1.765
+ $X2=6.155 $Y2=1.542
r151 16 18 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.155 $Y=1.765
+ $X2=6.155 $Y2=2.4
r152 13 41 66.1563 $w=2.59e-07 $l=3.34066e-07 $layer=POLY_cond $X=4.43 $Y=2.465
+ $X2=4.48 $Y2=2.155
r153 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.43 $Y=2.465
+ $X2=4.43 $Y2=2.75
r154 12 41 2.36368 $w=3.3e-07 $l=8.75758e-08 $layer=POLY_cond $X=4.48 $Y=2.155
+ $X2=4.48 $Y2=2.155
r155 11 32 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.48 $Y=1.975
+ $X2=4.48 $Y2=1.81
r156 11 12 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=4.48 $Y=1.975
+ $X2=4.48 $Y2=2.155
r157 9 32 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=4.39 $Y=0.83
+ $X2=4.39 $Y2=1.81
r158 2 55 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=5.22
+ $Y=1.84 $X2=5.37 $Y2=2.815
r159 2 52 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=5.22
+ $Y=1.84 $X2=5.37 $Y2=1.985
r160 1 45 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.045
+ $Y=0.37 $X2=5.185 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__DLXBP_1%A_664_392# 1 2 9 11 13 14 20 22 23 25 26 30
+ 33
c85 30 0 1.77373e-19 $X=4.87 $Y=1.405
c86 11 0 1.88618e-19 $X=5.145 $Y=1.765
r87 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.87
+ $Y=1.405 $X2=4.87 $Y2=1.405
r88 28 30 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=4.87 $Y=1.65
+ $X2=4.87 $Y2=1.405
r89 27 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.95 $Y=1.735
+ $X2=3.865 $Y2=1.735
r90 26 28 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.705 $Y=1.735
+ $X2=4.87 $Y2=1.65
r91 26 27 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=4.705 $Y=1.735
+ $X2=3.95 $Y2=1.735
r92 25 33 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.865 $Y=1.65
+ $X2=3.865 $Y2=1.735
r93 24 25 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=3.865 $Y=0.85
+ $X2=3.865 $Y2=1.65
r94 22 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.78 $Y=1.735
+ $X2=3.865 $Y2=1.735
r95 22 23 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=3.78 $Y=1.735
+ $X2=3.555 $Y2=1.735
r96 18 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.47 $Y=1.82
+ $X2=3.555 $Y2=1.735
r97 18 20 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=3.47 $Y=1.82
+ $X2=3.47 $Y2=2.105
r98 14 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.78 $Y=0.765
+ $X2=3.865 $Y2=0.85
r99 14 16 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=3.78 $Y=0.765
+ $X2=3.63 $Y2=0.765
r100 11 31 66.7694 $w=3.34e-07 $l=4.38862e-07 $layer=POLY_cond $X=5.145 $Y=1.765
+ $X2=4.97 $Y2=1.405
r101 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.145 $Y=1.765
+ $X2=5.145 $Y2=2.4
r102 7 31 38.6287 $w=3.34e-07 $l=1.65e-07 $layer=POLY_cond $X=4.97 $Y=1.24
+ $X2=4.97 $Y2=1.405
r103 7 9 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=4.97 $Y=1.24 $X2=4.97
+ $Y2=0.74
r104 2 20 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=3.32
+ $Y=1.96 $X2=3.47 $Y2=2.105
r105 1 16 182 $w=1.7e-07 $l=4.90816e-07 $layer=licon1_NDIFF $count=1 $X=3.335
+ $Y=0.4 $X2=3.63 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LS__DLXBP_1%A_1347_424# 1 2 7 9 12 14 15 18 22 28
c44 18 0 9.14246e-20 $X=6.89 $Y=0.855
r45 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.155
+ $Y=1.485 $X2=7.155 $Y2=1.485
r46 26 28 9.35923 $w=3.28e-07 $l=2.68e-07 $layer=LI1_cond $X=6.887 $Y=1.485
+ $X2=7.155 $Y2=1.485
r47 24 26 0.069845 $w=3.28e-07 $l=2e-09 $layer=LI1_cond $X=6.885 $Y=1.485
+ $X2=6.887 $Y2=1.485
r48 20 24 0.716491 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=6.885 $Y=1.65
+ $X2=6.885 $Y2=1.485
r49 20 22 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=6.885 $Y=1.65
+ $X2=6.885 $Y2=2.265
r50 16 26 0.643053 $w=3.35e-07 $l=1.65e-07 $layer=LI1_cond $X=6.887 $Y=1.32
+ $X2=6.887 $Y2=1.485
r51 16 18 15.9966 $w=3.33e-07 $l=4.65e-07 $layer=LI1_cond $X=6.887 $Y=1.32
+ $X2=6.887 $Y2=0.855
r52 14 29 72.5674 $w=3.3e-07 $l=4.15e-07 $layer=POLY_cond $X=7.57 $Y=1.485
+ $X2=7.155 $Y2=1.485
r53 14 15 5.03009 $w=3.3e-07 $l=1.15022e-07 $layer=POLY_cond $X=7.57 $Y=1.485
+ $X2=7.66 $Y2=1.542
r54 10 15 37.0704 $w=1.5e-07 $l=2.24486e-07 $layer=POLY_cond $X=7.665 $Y=1.32
+ $X2=7.66 $Y2=1.542
r55 10 12 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=7.665 $Y=1.32
+ $X2=7.665 $Y2=0.74
r56 7 15 37.0704 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=7.66 $Y=1.765
+ $X2=7.66 $Y2=1.542
r57 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.66 $Y=1.765
+ $X2=7.66 $Y2=2.4
r58 2 22 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=6.735
+ $Y=2.12 $X2=6.885 $Y2=2.265
r59 1 18 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=6.75
+ $Y=0.58 $X2=6.89 $Y2=0.855
.ends

.subckt PM_SKY130_FD_SC_LS__DLXBP_1%VPWR 1 2 3 4 5 20 24 26 30 34 38 43 44 46 47
+ 48 50 69 70 73 76 79
r92 79 80 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r93 76 77 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r94 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r95 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r96 67 70 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.92 $Y2=3.33
r97 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r98 64 67 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.96
+ $Y2=3.33
r99 63 64 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r100 61 64 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33 $X2=6
+ $Y2=3.33
r101 61 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r102 60 63 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=5.04 $Y=3.33 $X2=6
+ $Y2=3.33
r103 60 61 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r104 58 79 11.8853 $w=1.7e-07 $l=2.73e-07 $layer=LI1_cond $X=5.035 $Y=3.33
+ $X2=4.762 $Y2=3.33
r105 58 60 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=5.035 $Y=3.33
+ $X2=5.04 $Y2=3.33
r106 57 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r107 56 57 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r108 54 57 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r109 54 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r110 53 56 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r111 53 54 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r112 51 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.97 $Y=3.33
+ $X2=0.805 $Y2=3.33
r113 51 53 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=0.97 $Y=3.33
+ $X2=1.2 $Y2=3.33
r114 50 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.38 $Y=3.33
+ $X2=2.545 $Y2=3.33
r115 50 56 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=2.38 $Y=3.33
+ $X2=2.16 $Y2=3.33
r116 48 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r117 48 77 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=2.64 $Y2=3.33
r118 46 66 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=7.27 $Y=3.33
+ $X2=6.96 $Y2=3.33
r119 46 47 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.27 $Y=3.33
+ $X2=7.395 $Y2=3.33
r120 45 69 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=7.52 $Y=3.33 $X2=7.92
+ $Y2=3.33
r121 45 47 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.52 $Y=3.33
+ $X2=7.395 $Y2=3.33
r122 43 63 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=6.295 $Y=3.33 $X2=6
+ $Y2=3.33
r123 43 44 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.295 $Y=3.33
+ $X2=6.42 $Y2=3.33
r124 42 66 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=6.545 $Y=3.33
+ $X2=6.96 $Y2=3.33
r125 42 44 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.545 $Y=3.33
+ $X2=6.42 $Y2=3.33
r126 38 41 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=7.395 $Y=1.985
+ $X2=7.395 $Y2=2.815
r127 36 47 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.395 $Y=3.245
+ $X2=7.395 $Y2=3.33
r128 36 41 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=7.395 $Y=3.245
+ $X2=7.395 $Y2=2.815
r129 32 44 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.42 $Y=3.245
+ $X2=6.42 $Y2=3.33
r130 32 34 45.1758 $w=2.48e-07 $l=9.8e-07 $layer=LI1_cond $X=6.42 $Y=3.245
+ $X2=6.42 $Y2=2.265
r131 28 79 2.29102 $w=5.45e-07 $l=8.5e-08 $layer=LI1_cond $X=4.762 $Y=3.245
+ $X2=4.762 $Y2=3.33
r132 28 30 11.7413 $w=5.43e-07 $l=5.35e-07 $layer=LI1_cond $X=4.762 $Y=3.245
+ $X2=4.762 $Y2=2.71
r133 27 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.71 $Y=3.33
+ $X2=2.545 $Y2=3.33
r134 26 79 11.8853 $w=1.7e-07 $l=2.72e-07 $layer=LI1_cond $X=4.49 $Y=3.33
+ $X2=4.762 $Y2=3.33
r135 26 27 116.128 $w=1.68e-07 $l=1.78e-06 $layer=LI1_cond $X=4.49 $Y=3.33
+ $X2=2.71 $Y2=3.33
r136 22 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.545 $Y=3.245
+ $X2=2.545 $Y2=3.33
r137 22 24 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=2.545 $Y=3.245
+ $X2=2.545 $Y2=2.945
r138 18 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.805 $Y=3.245
+ $X2=0.805 $Y2=3.33
r139 18 20 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=0.805 $Y=3.245
+ $X2=0.805 $Y2=3.05
r140 5 41 400 $w=1.7e-07 $l=1.04265e-06 $layer=licon1_PDIFF $count=1 $X=7.295
+ $Y=1.84 $X2=7.435 $Y2=2.815
r141 5 38 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=7.295
+ $Y=1.84 $X2=7.435 $Y2=1.985
r142 4 34 300 $w=1.7e-07 $l=4.94343e-07 $layer=licon1_PDIFF $count=2 $X=6.23
+ $Y=1.84 $X2=6.38 $Y2=2.265
r143 3 30 600 $w=1.7e-07 $l=3.29204e-07 $layer=licon1_PDIFF $count=1 $X=4.505
+ $Y=2.54 $X2=4.76 $Y2=2.71
r144 2 24 600 $w=1.7e-07 $l=1.09397e-06 $layer=licon1_PDIFF $count=1 $X=2.315
+ $Y=1.96 $X2=2.545 $Y2=2.945
r145 1 20 600 $w=1.7e-07 $l=1.09397e-06 $layer=licon1_PDIFF $count=1 $X=0.575
+ $Y=2.065 $X2=0.805 $Y2=3.05
.ends

.subckt PM_SKY130_FD_SC_LS__DLXBP_1%Q 1 2 9 14 15 16 17 28
r39 21 28 2.09535 $w=3.28e-07 $l=6e-08 $layer=LI1_cond $X=5.96 $Y=0.985 $X2=5.96
+ $Y2=0.925
r40 17 30 8.04311 $w=3.28e-07 $l=1.53e-07 $layer=LI1_cond $X=5.96 $Y=0.997
+ $X2=5.96 $Y2=1.15
r41 17 21 0.41907 $w=3.28e-07 $l=1.2e-08 $layer=LI1_cond $X=5.96 $Y=0.997
+ $X2=5.96 $Y2=0.985
r42 17 28 0.453993 $w=3.28e-07 $l=1.3e-08 $layer=LI1_cond $X=5.96 $Y=0.912
+ $X2=5.96 $Y2=0.925
r43 16 17 13.1658 $w=3.28e-07 $l=3.77e-07 $layer=LI1_cond $X=5.96 $Y=0.535
+ $X2=5.96 $Y2=0.912
r44 15 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.04 $Y=1.82
+ $X2=6.04 $Y2=1.15
r45 14 15 8.51103 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=5.945 $Y=1.985
+ $X2=5.945 $Y2=1.82
r46 7 14 0.480185 $w=3.58e-07 $l=1.5e-08 $layer=LI1_cond $X=5.945 $Y=2 $X2=5.945
+ $Y2=1.985
r47 7 9 26.09 $w=3.58e-07 $l=8.15e-07 $layer=LI1_cond $X=5.945 $Y=2 $X2=5.945
+ $Y2=2.815
r48 2 14 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=5.785
+ $Y=1.84 $X2=5.93 $Y2=1.985
r49 2 9 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=5.785
+ $Y=1.84 $X2=5.93 $Y2=2.815
r50 1 16 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.82
+ $Y=0.39 $X2=5.96 $Y2=0.535
.ends

.subckt PM_SKY130_FD_SC_LS__DLXBP_1%Q_N 1 2 7 8 9 10 11 12 13
r14 12 13 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=7.882 $Y=2.405
+ $X2=7.882 $Y2=2.775
r15 11 12 14.4485 $w=3.33e-07 $l=4.2e-07 $layer=LI1_cond $X=7.882 $Y=1.985
+ $X2=7.882 $Y2=2.405
r16 10 11 11.0084 $w=3.33e-07 $l=3.2e-07 $layer=LI1_cond $X=7.882 $Y=1.665
+ $X2=7.882 $Y2=1.985
r17 9 10 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=7.882 $Y=1.295
+ $X2=7.882 $Y2=1.665
r18 8 9 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=7.882 $Y=0.925
+ $X2=7.882 $Y2=1.295
r19 7 8 14.1045 $w=3.33e-07 $l=4.1e-07 $layer=LI1_cond $X=7.882 $Y=0.515
+ $X2=7.882 $Y2=0.925
r20 2 13 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=7.735
+ $Y=1.84 $X2=7.885 $Y2=2.815
r21 2 11 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=7.735
+ $Y=1.84 $X2=7.885 $Y2=1.985
r22 1 7 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.74
+ $Y=0.37 $X2=7.88 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__DLXBP_1%VGND 1 2 3 4 5 18 22 26 30 33 34 35 37 42 50
+ 62 68 69 72 82 85
r85 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r86 82 83 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r87 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r88 69 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=7.44
+ $Y2=0
r89 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r90 66 85 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.535 $Y=0 $X2=7.41
+ $Y2=0
r91 66 68 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=7.535 $Y=0 $X2=7.92
+ $Y2=0
r92 65 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r93 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r94 62 85 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.285 $Y=0 $X2=7.41
+ $Y2=0
r95 62 64 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=7.285 $Y=0 $X2=6.96
+ $Y2=0
r96 61 65 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.96
+ $Y2=0
r97 60 61 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r98 58 61 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=6
+ $Y2=0
r99 58 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.56
+ $Y2=0
r100 57 60 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=5.04 $Y=0 $X2=6
+ $Y2=0
r101 57 58 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r102 55 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.85 $Y=0 $X2=4.685
+ $Y2=0
r103 55 57 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=4.85 $Y=0 $X2=5.04
+ $Y2=0
r104 54 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r105 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r106 51 53 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=2.74 $Y=0 $X2=3.12
+ $Y2=0
r107 50 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.52 $Y=0 $X2=4.685
+ $Y2=0
r108 50 53 91.3369 $w=1.68e-07 $l=1.4e-06 $layer=LI1_cond $X=4.52 $Y=0 $X2=3.12
+ $Y2=0
r109 49 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r110 48 49 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r111 46 49 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r112 46 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r113 45 48 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r114 45 46 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r115 43 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.96 $Y=0 $X2=0.795
+ $Y2=0
r116 43 45 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=0.96 $Y=0 $X2=1.2
+ $Y2=0
r117 42 79 9.72841 $w=3.83e-07 $l=3.25e-07 $layer=LI1_cond $X=2.547 $Y=0
+ $X2=2.547 $Y2=0.325
r118 42 51 5.54671 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=2.547 $Y=0 $X2=2.74
+ $Y2=0
r119 42 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r120 42 48 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=2.355 $Y=0
+ $X2=2.16 $Y2=0
r121 40 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r122 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r123 37 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.63 $Y=0 $X2=0.795
+ $Y2=0
r124 37 39 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=0.63 $Y=0 $X2=0.24
+ $Y2=0
r125 35 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r126 35 54 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.12
+ $Y2=0
r127 33 60 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=6.295 $Y=0 $X2=6
+ $Y2=0
r128 33 34 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.295 $Y=0 $X2=6.42
+ $Y2=0
r129 32 64 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=6.545 $Y=0
+ $X2=6.96 $Y2=0
r130 32 34 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.545 $Y=0 $X2=6.42
+ $Y2=0
r131 28 85 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.41 $Y=0.085
+ $X2=7.41 $Y2=0
r132 28 30 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=7.41 $Y=0.085
+ $X2=7.41 $Y2=0.515
r133 24 34 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.42 $Y=0.085
+ $X2=6.42 $Y2=0
r134 24 26 35.4952 $w=2.48e-07 $l=7.7e-07 $layer=LI1_cond $X=6.42 $Y=0.085
+ $X2=6.42 $Y2=0.855
r135 20 82 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.685 $Y=0.085
+ $X2=4.685 $Y2=0
r136 20 22 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=4.685 $Y=0.085
+ $X2=4.685 $Y2=0.515
r137 16 72 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.795 $Y=0.085
+ $X2=0.795 $Y2=0
r138 16 18 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=0.795 $Y=0.085
+ $X2=0.795 $Y2=0.52
r139 5 30 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=7.305
+ $Y=0.37 $X2=7.45 $Y2=0.515
r140 4 26 182 $w=1.7e-07 $l=5.45527e-07 $layer=licon1_NDIFF $count=1 $X=6.25
+ $Y=0.39 $X2=6.425 $Y2=0.855
r141 3 22 91 $w=1.7e-07 $l=2.67395e-07 $layer=licon1_NDIFF $count=2 $X=4.465
+ $Y=0.62 $X2=4.685 $Y2=0.515
r142 2 79 182 $w=1.7e-07 $l=2.84341e-07 $layer=licon1_NDIFF $count=1 $X=2.3
+ $Y=0.41 $X2=2.545 $Y2=0.325
r143 1 18 91 $w=1.7e-07 $l=2.39165e-07 $layer=licon1_NDIFF $count=2 $X=0.575
+ $Y=0.56 $X2=0.795 $Y2=0.52
.ends

