* File: sky130_fd_sc_ls__maj3_1.pxi.spice
* Created: Wed Sep  2 11:09:48 2020
* 
x_PM_SKY130_FD_SC_LS__MAJ3_1%A_84_74# N_A_84_74#_M1004_d N_A_84_74#_M1008_d
+ N_A_84_74#_M1001_d N_A_84_74#_M1011_d N_A_84_74#_c_69_n N_A_84_74#_M1003_g
+ N_A_84_74#_c_70_n N_A_84_74#_M1009_g N_A_84_74#_c_71_n N_A_84_74#_c_72_n
+ N_A_84_74#_c_73_n N_A_84_74#_c_79_n N_A_84_74#_c_74_n N_A_84_74#_c_104_p
+ N_A_84_74#_c_75_n N_A_84_74#_c_108_p N_A_84_74#_c_81_n N_A_84_74#_c_82_n
+ N_A_84_74#_c_94_p N_A_84_74#_c_76_n PM_SKY130_FD_SC_LS__MAJ3_1%A_84_74#
x_PM_SKY130_FD_SC_LS__MAJ3_1%B N_B_M1004_g N_B_c_183_n N_B_M1001_g N_B_c_180_n
+ N_B_M1013_g N_B_c_184_n N_B_M1010_g B N_B_c_181_n N_B_c_182_n
+ PM_SKY130_FD_SC_LS__MAJ3_1%B
x_PM_SKY130_FD_SC_LS__MAJ3_1%C N_C_c_231_n N_C_M1007_g N_C_c_232_n N_C_M1006_g
+ N_C_c_233_n N_C_M1008_g N_C_c_234_n N_C_M1011_g N_C_c_235_n C N_C_c_236_n
+ PM_SKY130_FD_SC_LS__MAJ3_1%C
x_PM_SKY130_FD_SC_LS__MAJ3_1%A N_A_M1012_g N_A_c_289_n N_A_c_290_n N_A_c_300_n
+ N_A_M1002_g N_A_c_291_n N_A_c_292_n N_A_M1005_g N_A_c_294_n N_A_c_295_n
+ N_A_c_302_n N_A_M1000_g A N_A_c_297_n N_A_c_298_n PM_SKY130_FD_SC_LS__MAJ3_1%A
x_PM_SKY130_FD_SC_LS__MAJ3_1%X N_X_M1003_s N_X_M1009_s N_X_c_368_n N_X_c_369_n X
+ X X N_X_c_370_n PM_SKY130_FD_SC_LS__MAJ3_1%X
x_PM_SKY130_FD_SC_LS__MAJ3_1%VPWR N_VPWR_M1009_d N_VPWR_M1006_d N_VPWR_c_390_n
+ N_VPWR_c_391_n VPWR N_VPWR_c_392_n N_VPWR_c_393_n N_VPWR_c_389_n
+ N_VPWR_c_395_n N_VPWR_c_396_n PM_SKY130_FD_SC_LS__MAJ3_1%VPWR
x_PM_SKY130_FD_SC_LS__MAJ3_1%VGND N_VGND_M1003_d N_VGND_M1007_d N_VGND_c_432_n
+ N_VGND_c_433_n N_VGND_c_449_n N_VGND_c_450_n N_VGND_c_434_n N_VGND_c_435_n
+ VGND N_VGND_c_436_n N_VGND_c_437_n N_VGND_c_438_n N_VGND_c_439_n
+ PM_SKY130_FD_SC_LS__MAJ3_1%VGND
cc_1 VNB N_A_84_74#_c_69_n 0.0215805f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.35
cc_2 VNB N_A_84_74#_c_70_n 0.0269151f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.765
cc_3 VNB N_A_84_74#_c_71_n 0.00825211f $X=-0.19 $Y=-0.245 $X2=1.48 $Y2=1.175
cc_4 VNB N_A_84_74#_c_72_n 0.00591492f $X=-0.19 $Y=-0.245 $X2=0.785 $Y2=1.175
cc_5 VNB N_A_84_74#_c_73_n 0.00347054f $X=-0.19 $Y=-0.245 $X2=1.645 $Y2=0.745
cc_6 VNB N_A_84_74#_c_74_n 0.00257431f $X=-0.19 $Y=-0.245 $X2=1.98 $Y2=1.95
cc_7 VNB N_A_84_74#_c_75_n 9.46947e-19 $X=-0.19 $Y=-0.245 $X2=2.065 $Y2=1.175
cc_8 VNB N_A_84_74#_c_76_n 0.0172793f $X=-0.19 $Y=-0.245 $X2=3.535 $Y2=1.05
cc_9 VNB N_B_M1004_g 0.021382f $X=-0.19 $Y=-0.245 $X2=1.55 $Y2=1.92
cc_10 VNB N_B_c_180_n 0.0152338f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_B_c_181_n 0.00195337f $X=-0.19 $Y=-0.245 $X2=0.785 $Y2=1.175
cc_12 VNB N_B_c_182_n 0.0266992f $X=-0.19 $Y=-0.245 $X2=1.645 $Y2=1.09
cc_13 VNB N_C_c_231_n 0.0134552f $X=-0.19 $Y=-0.245 $X2=1.505 $Y2=0.6
cc_14 VNB N_C_c_232_n 0.0222531f $X=-0.19 $Y=-0.245 $X2=3.41 $Y2=1.92
cc_15 VNB N_C_c_233_n 0.0207444f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_C_c_234_n 0.0216443f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_C_c_235_n 0.0121979f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.87
cc_18 VNB N_C_c_236_n 0.00130225f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_M1012_g 0.0285172f $X=-0.19 $Y=-0.245 $X2=3.41 $Y2=1.92
cc_20 VNB N_A_c_289_n 0.00563382f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_c_290_n 0.0117219f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_c_291_n 0.115517f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_c_292_n 0.011606f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_M1005_g 0.0107186f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.87
cc_25 VNB N_A_c_294_n 0.00491764f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.765
cc_26 VNB N_A_c_295_n 0.00711931f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=2.4
cc_27 VNB A 0.0240534f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_c_297_n 0.0540726f $X=-0.19 $Y=-0.245 $X2=1.98 $Y2=1.95
cc_29 VNB N_A_c_298_n 0.0129204f $X=-0.19 $Y=-0.245 $X2=3.56 $Y2=2.12
cc_30 VNB N_X_c_368_n 0.0241167f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_X_c_369_n 0.00713231f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.35
cc_32 VNB N_X_c_370_n 0.0221111f $X=-0.19 $Y=-0.245 $X2=1.98 $Y2=1.95
cc_33 VNB N_VPWR_c_389_n 0.163682f $X=-0.19 $Y=-0.245 $X2=2.065 $Y2=1.175
cc_34 VNB N_VGND_c_432_n 0.0108282f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_433_n 0.0136584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_434_n 0.0381259f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=2.4
cc_37 VNB N_VGND_c_435_n 0.00229531f $X=-0.19 $Y=-0.245 $X2=1.48 $Y2=1.175
cc_38 VNB N_VGND_c_436_n 0.0195478f $X=-0.19 $Y=-0.245 $X2=1.645 $Y2=0.745
cc_39 VNB N_VGND_c_437_n 0.0337601f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_438_n 0.221862f $X=-0.19 $Y=-0.245 $X2=0.785 $Y2=1.175
cc_41 VNB N_VGND_c_439_n 0.00603779f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.515
cc_42 VPB N_A_84_74#_c_70_n 0.0334283f $X=-0.19 $Y=1.66 $X2=0.55 $Y2=1.765
cc_43 VPB N_A_84_74#_c_72_n 0.00269398f $X=-0.19 $Y=1.66 $X2=0.785 $Y2=1.175
cc_44 VPB N_A_84_74#_c_79_n 0.00315149f $X=-0.19 $Y=1.66 $X2=1.73 $Y2=2.775
cc_45 VPB N_A_84_74#_c_74_n 0.00218641f $X=-0.19 $Y=1.66 $X2=1.98 $Y2=1.95
cc_46 VPB N_A_84_74#_c_81_n 0.00861803f $X=-0.19 $Y=1.66 $X2=3.56 $Y2=2.12
cc_47 VPB N_A_84_74#_c_82_n 0.0340653f $X=-0.19 $Y=1.66 $X2=3.56 $Y2=2.775
cc_48 VPB N_B_c_183_n 0.015006f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 VPB N_B_c_184_n 0.0144655f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_B_c_181_n 0.0102481f $X=-0.19 $Y=1.66 $X2=0.785 $Y2=1.175
cc_51 VPB N_B_c_182_n 0.0293257f $X=-0.19 $Y=1.66 $X2=1.645 $Y2=1.09
cc_52 VPB N_C_c_232_n 0.0320882f $X=-0.19 $Y=1.66 $X2=3.41 $Y2=1.92
cc_53 VPB N_C_c_234_n 0.0393073f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_C_c_235_n 0.00701532f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.87
cc_55 VPB N_C_c_236_n 0.00302418f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_A_c_290_n 0.00463031f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_A_c_300_n 0.0209357f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_A_c_295_n 0.00384606f $X=-0.19 $Y=1.66 $X2=0.55 $Y2=2.4
cc_59 VPB N_A_c_302_n 0.021495f $X=-0.19 $Y=1.66 $X2=0.55 $Y2=2.4
cc_60 VPB X 0.0504915f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.87
cc_61 VPB N_X_c_370_n 0.00919986f $X=-0.19 $Y=1.66 $X2=1.98 $Y2=1.95
cc_62 VPB N_VPWR_c_390_n 0.00803717f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_391_n 0.0106519f $X=-0.19 $Y=1.66 $X2=0.55 $Y2=2.4
cc_64 VPB N_VPWR_c_392_n 0.0435502f $X=-0.19 $Y=1.66 $X2=1.645 $Y2=1.09
cc_65 VPB N_VPWR_c_393_n 0.0315964f $X=-0.19 $Y=1.66 $X2=3.37 $Y2=1.175
cc_66 VPB N_VPWR_c_389_n 0.103296f $X=-0.19 $Y=1.66 $X2=2.065 $Y2=1.175
cc_67 VPB N_VPWR_c_395_n 0.0263192f $X=-0.19 $Y=1.66 $X2=3.56 $Y2=2.12
cc_68 VPB N_VPWR_c_396_n 0.00776418f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 N_A_84_74#_c_71_n N_B_M1004_g 0.0106503f $X=1.48 $Y=1.175 $X2=0 $Y2=0
cc_70 N_A_84_74#_c_73_n N_B_M1004_g 0.00928072f $X=1.645 $Y=0.745 $X2=0 $Y2=0
cc_71 N_A_84_74#_c_74_n N_B_M1004_g 9.50889e-19 $X=1.98 $Y=1.95 $X2=0 $Y2=0
cc_72 N_A_84_74#_c_75_n N_B_M1004_g 0.00112012f $X=2.065 $Y=1.175 $X2=0 $Y2=0
cc_73 N_A_84_74#_c_79_n N_B_c_183_n 2.93854e-19 $X=1.73 $Y=2.775 $X2=0 $Y2=0
cc_74 N_A_84_74#_c_74_n N_B_c_183_n 5.27837e-19 $X=1.98 $Y=1.95 $X2=0 $Y2=0
cc_75 N_A_84_74#_c_73_n N_B_c_180_n 0.00347549f $X=1.645 $Y=0.745 $X2=0 $Y2=0
cc_76 N_A_84_74#_c_74_n N_B_c_180_n 0.00527567f $X=1.98 $Y=1.95 $X2=0 $Y2=0
cc_77 N_A_84_74#_c_75_n N_B_c_180_n 0.0145609f $X=2.065 $Y=1.175 $X2=0 $Y2=0
cc_78 N_A_84_74#_c_79_n N_B_c_184_n 0.0142858f $X=1.73 $Y=2.775 $X2=0 $Y2=0
cc_79 N_A_84_74#_c_74_n N_B_c_184_n 0.00308979f $X=1.98 $Y=1.95 $X2=0 $Y2=0
cc_80 N_A_84_74#_c_94_p N_B_c_184_n 0.0119912f $X=1.73 $Y=2.095 $X2=0 $Y2=0
cc_81 N_A_84_74#_c_70_n N_B_c_181_n 7.27044e-19 $X=0.55 $Y=1.765 $X2=0 $Y2=0
cc_82 N_A_84_74#_c_71_n N_B_c_181_n 0.0453726f $X=1.48 $Y=1.175 $X2=0 $Y2=0
cc_83 N_A_84_74#_c_72_n N_B_c_181_n 0.0136497f $X=0.785 $Y=1.175 $X2=0 $Y2=0
cc_84 N_A_84_74#_c_74_n N_B_c_181_n 0.0222188f $X=1.98 $Y=1.95 $X2=0 $Y2=0
cc_85 N_A_84_74#_c_94_p N_B_c_181_n 0.00856258f $X=1.73 $Y=2.095 $X2=0 $Y2=0
cc_86 N_A_84_74#_c_74_n N_B_c_182_n 0.0138852f $X=1.98 $Y=1.95 $X2=0 $Y2=0
cc_87 N_A_84_74#_c_75_n N_B_c_182_n 0.00539881f $X=2.065 $Y=1.175 $X2=0 $Y2=0
cc_88 N_A_84_74#_c_94_p N_B_c_182_n 0.00795607f $X=1.73 $Y=2.095 $X2=0 $Y2=0
cc_89 N_A_84_74#_c_74_n N_C_c_231_n 0.0042291f $X=1.98 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_90 N_A_84_74#_c_104_p N_C_c_231_n 0.0131284f $X=3.37 $Y=1.175 $X2=-0.19
+ $Y2=-0.245
cc_91 N_A_84_74#_c_79_n N_C_c_232_n 0.00268978f $X=1.73 $Y=2.775 $X2=0 $Y2=0
cc_92 N_A_84_74#_c_74_n N_C_c_232_n 0.00282f $X=1.98 $Y=1.95 $X2=0 $Y2=0
cc_93 N_A_84_74#_c_104_p N_C_c_232_n 0.00501252f $X=3.37 $Y=1.175 $X2=0 $Y2=0
cc_94 N_A_84_74#_c_108_p N_C_c_232_n 0.0159689f $X=3.395 $Y=2.035 $X2=0 $Y2=0
cc_95 N_A_84_74#_c_104_p N_C_c_233_n 0.00928007f $X=3.37 $Y=1.175 $X2=0 $Y2=0
cc_96 N_A_84_74#_c_76_n N_C_c_233_n 0.00674358f $X=3.535 $Y=1.05 $X2=0 $Y2=0
cc_97 N_A_84_74#_c_108_p N_C_c_234_n 0.0118897f $X=3.395 $Y=2.035 $X2=0 $Y2=0
cc_98 N_A_84_74#_c_81_n N_C_c_234_n 0.00414271f $X=3.56 $Y=2.12 $X2=0 $Y2=0
cc_99 N_A_84_74#_c_82_n N_C_c_234_n 0.0146053f $X=3.56 $Y=2.775 $X2=0 $Y2=0
cc_100 N_A_84_74#_c_76_n N_C_c_234_n 0.00405163f $X=3.535 $Y=1.05 $X2=0 $Y2=0
cc_101 N_A_84_74#_c_108_p N_C_c_235_n 0.0381811f $X=3.395 $Y=2.035 $X2=0 $Y2=0
cc_102 N_A_84_74#_c_81_n N_C_c_235_n 0.0122229f $X=3.56 $Y=2.12 $X2=0 $Y2=0
cc_103 N_A_84_74#_c_76_n N_C_c_235_n 0.0137699f $X=3.535 $Y=1.05 $X2=0 $Y2=0
cc_104 N_A_84_74#_c_74_n N_C_c_236_n 0.0228466f $X=1.98 $Y=1.95 $X2=0 $Y2=0
cc_105 N_A_84_74#_c_104_p N_C_c_236_n 0.0728496f $X=3.37 $Y=1.175 $X2=0 $Y2=0
cc_106 N_A_84_74#_c_108_p N_C_c_236_n 0.0330871f $X=3.395 $Y=2.035 $X2=0 $Y2=0
cc_107 N_A_84_74#_c_69_n N_A_M1012_g 0.0199957f $X=0.495 $Y=1.35 $X2=0 $Y2=0
cc_108 N_A_84_74#_c_71_n N_A_M1012_g 0.0179611f $X=1.48 $Y=1.175 $X2=0 $Y2=0
cc_109 N_A_84_74#_c_72_n N_A_M1012_g 0.0055338f $X=0.785 $Y=1.175 $X2=0 $Y2=0
cc_110 N_A_84_74#_c_73_n N_A_M1012_g 0.00182632f $X=1.645 $Y=0.745 $X2=0 $Y2=0
cc_111 N_A_84_74#_c_70_n N_A_c_289_n 0.0197603f $X=0.55 $Y=1.765 $X2=0 $Y2=0
cc_112 N_A_84_74#_c_71_n N_A_c_289_n 8.77498e-19 $X=1.48 $Y=1.175 $X2=0 $Y2=0
cc_113 N_A_84_74#_c_70_n N_A_c_290_n 0.00339363f $X=0.55 $Y=1.765 $X2=0 $Y2=0
cc_114 N_A_84_74#_c_70_n N_A_c_300_n 0.0223224f $X=0.55 $Y=1.765 $X2=0 $Y2=0
cc_115 N_A_84_74#_c_73_n N_A_c_291_n 0.00612247f $X=1.645 $Y=0.745 $X2=0 $Y2=0
cc_116 N_A_84_74#_c_104_p N_A_M1005_g 0.0124955f $X=3.37 $Y=1.175 $X2=0 $Y2=0
cc_117 N_A_84_74#_c_76_n N_A_M1005_g 0.00116861f $X=3.535 $Y=1.05 $X2=0 $Y2=0
cc_118 N_A_84_74#_c_108_p N_A_c_302_n 0.0156091f $X=3.395 $Y=2.035 $X2=0 $Y2=0
cc_119 N_A_84_74#_c_82_n N_A_c_302_n 0.0027017f $X=3.56 $Y=2.775 $X2=0 $Y2=0
cc_120 N_A_84_74#_c_76_n A 0.0178486f $X=3.535 $Y=1.05 $X2=0 $Y2=0
cc_121 N_A_84_74#_c_104_p N_A_c_298_n 0.0147496f $X=3.37 $Y=1.175 $X2=0 $Y2=0
cc_122 N_A_84_74#_c_76_n N_A_c_298_n 0.00467871f $X=3.535 $Y=1.05 $X2=0 $Y2=0
cc_123 N_A_84_74#_c_69_n N_X_c_368_n 0.00692086f $X=0.495 $Y=1.35 $X2=0 $Y2=0
cc_124 N_A_84_74#_c_69_n N_X_c_369_n 0.00300451f $X=0.495 $Y=1.35 $X2=0 $Y2=0
cc_125 N_A_84_74#_c_72_n N_X_c_369_n 0.00152814f $X=0.785 $Y=1.175 $X2=0 $Y2=0
cc_126 N_A_84_74#_c_70_n X 0.012884f $X=0.55 $Y=1.765 $X2=0 $Y2=0
cc_127 N_A_84_74#_c_72_n X 0.00297684f $X=0.785 $Y=1.175 $X2=0 $Y2=0
cc_128 N_A_84_74#_c_69_n N_X_c_370_n 0.0100022f $X=0.495 $Y=1.35 $X2=0 $Y2=0
cc_129 N_A_84_74#_c_70_n N_X_c_370_n 0.00398068f $X=0.55 $Y=1.765 $X2=0 $Y2=0
cc_130 N_A_84_74#_c_72_n N_X_c_370_n 0.0303017f $X=0.785 $Y=1.175 $X2=0 $Y2=0
cc_131 N_A_84_74#_c_108_p N_VPWR_M1006_d 0.00592102f $X=3.395 $Y=2.035 $X2=0
+ $Y2=0
cc_132 N_A_84_74#_c_70_n N_VPWR_c_390_n 0.00993395f $X=0.55 $Y=1.765 $X2=0 $Y2=0
cc_133 N_A_84_74#_c_72_n N_VPWR_c_390_n 0.00696688f $X=0.785 $Y=1.175 $X2=0
+ $Y2=0
cc_134 N_A_84_74#_c_79_n N_VPWR_c_390_n 0.0116001f $X=1.73 $Y=2.775 $X2=0 $Y2=0
cc_135 N_A_84_74#_c_79_n N_VPWR_c_391_n 0.0192031f $X=1.73 $Y=2.775 $X2=0 $Y2=0
cc_136 N_A_84_74#_c_108_p N_VPWR_c_391_n 0.0234793f $X=3.395 $Y=2.035 $X2=0
+ $Y2=0
cc_137 N_A_84_74#_c_82_n N_VPWR_c_391_n 0.00957552f $X=3.56 $Y=2.775 $X2=0 $Y2=0
cc_138 N_A_84_74#_c_79_n N_VPWR_c_392_n 0.0125658f $X=1.73 $Y=2.775 $X2=0 $Y2=0
cc_139 N_A_84_74#_c_82_n N_VPWR_c_393_n 0.0125658f $X=3.56 $Y=2.775 $X2=0 $Y2=0
cc_140 N_A_84_74#_c_70_n N_VPWR_c_389_n 0.00865353f $X=0.55 $Y=1.765 $X2=0 $Y2=0
cc_141 N_A_84_74#_c_79_n N_VPWR_c_389_n 0.011805f $X=1.73 $Y=2.775 $X2=0 $Y2=0
cc_142 N_A_84_74#_c_82_n N_VPWR_c_389_n 0.011805f $X=3.56 $Y=2.775 $X2=0 $Y2=0
cc_143 N_A_84_74#_c_70_n N_VPWR_c_395_n 0.00445602f $X=0.55 $Y=1.765 $X2=0 $Y2=0
cc_144 N_A_84_74#_c_108_p A_406_384# 0.0119045f $X=3.395 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_145 N_A_84_74#_c_108_p A_598_384# 0.00769472f $X=3.395 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_146 N_A_84_74#_c_71_n N_VGND_M1003_d 0.00132837f $X=1.48 $Y=1.175 $X2=-0.19
+ $Y2=-0.245
cc_147 N_A_84_74#_c_72_n N_VGND_M1003_d 0.00248319f $X=0.785 $Y=1.175 $X2=-0.19
+ $Y2=-0.245
cc_148 N_A_84_74#_c_104_p N_VGND_M1007_d 0.00661484f $X=3.37 $Y=1.175 $X2=0
+ $Y2=0
cc_149 N_A_84_74#_c_69_n N_VGND_c_432_n 0.00580418f $X=0.495 $Y=1.35 $X2=0 $Y2=0
cc_150 N_A_84_74#_c_70_n N_VGND_c_432_n 6.00018e-19 $X=0.55 $Y=1.765 $X2=0 $Y2=0
cc_151 N_A_84_74#_c_71_n N_VGND_c_432_n 0.0112589f $X=1.48 $Y=1.175 $X2=0 $Y2=0
cc_152 N_A_84_74#_c_72_n N_VGND_c_432_n 0.0135036f $X=0.785 $Y=1.175 $X2=0 $Y2=0
cc_153 N_A_84_74#_c_73_n N_VGND_c_432_n 0.0105579f $X=1.645 $Y=0.745 $X2=0 $Y2=0
cc_154 N_A_84_74#_c_73_n N_VGND_c_433_n 0.00420212f $X=1.645 $Y=0.745 $X2=0
+ $Y2=0
cc_155 N_A_84_74#_c_104_p N_VGND_c_449_n 0.00820442f $X=3.37 $Y=1.175 $X2=0
+ $Y2=0
cc_156 N_A_84_74#_c_104_p N_VGND_c_450_n 0.02198f $X=3.37 $Y=1.175 $X2=0 $Y2=0
cc_157 N_A_84_74#_c_76_n N_VGND_c_450_n 0.00216203f $X=3.535 $Y=1.05 $X2=0 $Y2=0
cc_158 N_A_84_74#_c_73_n N_VGND_c_434_n 0.00725358f $X=1.645 $Y=0.745 $X2=0
+ $Y2=0
cc_159 N_A_84_74#_c_69_n N_VGND_c_436_n 0.00467453f $X=0.495 $Y=1.35 $X2=0 $Y2=0
cc_160 N_A_84_74#_c_69_n N_VGND_c_438_n 0.00505379f $X=0.495 $Y=1.35 $X2=0 $Y2=0
cc_161 N_A_84_74#_c_73_n N_VGND_c_438_n 0.00890448f $X=1.645 $Y=0.745 $X2=0
+ $Y2=0
cc_162 N_A_84_74#_c_71_n A_223_120# 0.0048076f $X=1.48 $Y=1.175 $X2=-0.19
+ $Y2=-0.245
cc_163 N_A_84_74#_c_104_p A_403_136# 0.0096152f $X=3.37 $Y=1.175 $X2=-0.19
+ $Y2=-0.245
cc_164 N_A_84_74#_c_104_p A_595_136# 0.00453974f $X=3.37 $Y=1.175 $X2=-0.19
+ $Y2=-0.245
cc_165 N_B_c_180_n N_C_c_231_n 0.0451321f $X=1.94 $Y=1.43 $X2=-0.19 $Y2=-0.245
cc_166 N_B_c_184_n N_C_c_232_n 0.0533449f $X=1.955 $Y=1.845 $X2=0 $Y2=0
cc_167 N_B_c_182_n N_C_c_232_n 0.0252957f $X=1.94 $Y=1.637 $X2=0 $Y2=0
cc_168 N_B_c_182_n N_C_c_236_n 3.98061e-19 $X=1.94 $Y=1.637 $X2=0 $Y2=0
cc_169 N_B_M1004_g N_A_M1012_g 0.0437821f $X=1.43 $Y=0.92 $X2=0 $Y2=0
cc_170 N_B_M1004_g N_A_c_289_n 0.0143676f $X=1.43 $Y=0.92 $X2=0 $Y2=0
cc_171 N_B_c_181_n N_A_c_290_n 0.00932579f $X=1.52 $Y=1.595 $X2=0 $Y2=0
cc_172 N_B_c_182_n N_A_c_290_n 0.0143676f $X=1.94 $Y=1.637 $X2=0 $Y2=0
cc_173 N_B_c_183_n N_A_c_300_n 0.0529837f $X=1.475 $Y=1.845 $X2=0 $Y2=0
cc_174 N_B_c_181_n N_A_c_300_n 0.00357958f $X=1.52 $Y=1.595 $X2=0 $Y2=0
cc_175 N_B_c_182_n N_A_c_300_n 0.00500143f $X=1.94 $Y=1.637 $X2=0 $Y2=0
cc_176 N_B_M1004_g N_A_c_291_n 0.0103098f $X=1.43 $Y=0.92 $X2=0 $Y2=0
cc_177 N_B_c_180_n N_A_c_291_n 0.00746712f $X=1.94 $Y=1.43 $X2=0 $Y2=0
cc_178 N_B_c_183_n N_VPWR_c_390_n 0.00339333f $X=1.475 $Y=1.845 $X2=0 $Y2=0
cc_179 N_B_c_184_n N_VPWR_c_391_n 0.00239997f $X=1.955 $Y=1.845 $X2=0 $Y2=0
cc_180 N_B_c_183_n N_VPWR_c_392_n 0.00548708f $X=1.475 $Y=1.845 $X2=0 $Y2=0
cc_181 N_B_c_184_n N_VPWR_c_392_n 0.00534256f $X=1.955 $Y=1.845 $X2=0 $Y2=0
cc_182 N_B_c_183_n N_VPWR_c_389_n 0.00533081f $X=1.475 $Y=1.845 $X2=0 $Y2=0
cc_183 N_B_c_184_n N_VPWR_c_389_n 0.00533081f $X=1.955 $Y=1.845 $X2=0 $Y2=0
cc_184 N_B_M1004_g N_VGND_c_432_n 0.00147743f $X=1.43 $Y=0.92 $X2=0 $Y2=0
cc_185 N_B_c_180_n N_VGND_c_433_n 7.10756e-19 $X=1.94 $Y=1.43 $X2=0 $Y2=0
cc_186 N_B_c_180_n N_VGND_c_449_n 5.65853e-19 $X=1.94 $Y=1.43 $X2=0 $Y2=0
cc_187 N_B_M1004_g N_VGND_c_438_n 9.33152e-19 $X=1.43 $Y=0.92 $X2=0 $Y2=0
cc_188 N_B_c_180_n N_VGND_c_438_n 9.5708e-19 $X=1.94 $Y=1.43 $X2=0 $Y2=0
cc_189 N_C_c_231_n N_A_c_291_n 0.00683881f $X=2.33 $Y=1.4 $X2=0 $Y2=0
cc_190 N_C_c_231_n N_A_M1005_g 0.0240392f $X=2.33 $Y=1.4 $X2=0 $Y2=0
cc_191 N_C_c_232_n N_A_c_294_n 0.0234459f $X=2.375 $Y=1.845 $X2=0 $Y2=0
cc_192 N_C_c_233_n N_A_c_294_n 0.0125649f $X=3.32 $Y=1.43 $X2=0 $Y2=0
cc_193 N_C_c_235_n N_A_c_294_n 0.00424265f $X=3.41 $Y=1.595 $X2=0 $Y2=0
cc_194 N_C_c_234_n N_A_c_295_n 0.0125649f $X=3.335 $Y=1.845 $X2=0 $Y2=0
cc_195 N_C_c_235_n N_A_c_295_n 0.00968576f $X=3.41 $Y=1.595 $X2=0 $Y2=0
cc_196 N_C_c_232_n N_A_c_302_n 0.0265045f $X=2.375 $Y=1.845 $X2=0 $Y2=0
cc_197 N_C_c_234_n N_A_c_302_n 0.0543315f $X=3.335 $Y=1.845 $X2=0 $Y2=0
cc_198 N_C_c_235_n N_A_c_302_n 0.00253689f $X=3.41 $Y=1.595 $X2=0 $Y2=0
cc_199 N_C_c_236_n N_A_c_302_n 5.65769e-19 $X=2.755 $Y=1.605 $X2=0 $Y2=0
cc_200 N_C_c_233_n A 0.00384087f $X=3.32 $Y=1.43 $X2=0 $Y2=0
cc_201 N_C_c_231_n N_A_c_297_n 0.00110103f $X=2.33 $Y=1.4 $X2=0 $Y2=0
cc_202 N_C_c_233_n N_A_c_297_n 0.040752f $X=3.32 $Y=1.43 $X2=0 $Y2=0
cc_203 N_C_c_233_n N_A_c_298_n 0.00756106f $X=3.32 $Y=1.43 $X2=0 $Y2=0
cc_204 N_C_c_232_n N_VPWR_c_391_n 0.0153663f $X=2.375 $Y=1.845 $X2=0 $Y2=0
cc_205 N_C_c_232_n N_VPWR_c_392_n 0.00492531f $X=2.375 $Y=1.845 $X2=0 $Y2=0
cc_206 N_C_c_234_n N_VPWR_c_393_n 0.00534256f $X=3.335 $Y=1.845 $X2=0 $Y2=0
cc_207 N_C_c_232_n N_VPWR_c_389_n 0.00483326f $X=2.375 $Y=1.845 $X2=0 $Y2=0
cc_208 N_C_c_234_n N_VPWR_c_389_n 0.00533081f $X=3.335 $Y=1.845 $X2=0 $Y2=0
cc_209 N_C_c_231_n N_VGND_c_433_n 0.00678491f $X=2.33 $Y=1.4 $X2=0 $Y2=0
cc_210 N_C_c_231_n N_VGND_c_449_n 0.00784325f $X=2.33 $Y=1.4 $X2=0 $Y2=0
cc_211 N_C_c_233_n N_VGND_c_450_n 6.83236e-19 $X=3.32 $Y=1.43 $X2=0 $Y2=0
cc_212 N_C_c_233_n N_VGND_c_437_n 4.78105e-19 $X=3.32 $Y=1.43 $X2=0 $Y2=0
cc_213 N_C_c_231_n N_VGND_c_438_n 3.25407e-19 $X=2.33 $Y=1.4 $X2=0 $Y2=0
cc_214 N_A_M1012_g N_X_c_368_n 8.44714e-19 $X=1.04 $Y=0.92 $X2=0 $Y2=0
cc_215 N_A_c_300_n X 6.52456e-19 $X=1.055 $Y=1.845 $X2=0 $Y2=0
cc_216 N_A_c_300_n N_VPWR_c_390_n 0.0209982f $X=1.055 $Y=1.845 $X2=0 $Y2=0
cc_217 N_A_c_302_n N_VPWR_c_391_n 0.00776455f $X=2.915 $Y=1.845 $X2=0 $Y2=0
cc_218 N_A_c_300_n N_VPWR_c_392_n 0.00510822f $X=1.055 $Y=1.845 $X2=0 $Y2=0
cc_219 N_A_c_302_n N_VPWR_c_393_n 0.00547402f $X=2.915 $Y=1.845 $X2=0 $Y2=0
cc_220 N_A_c_300_n N_VPWR_c_389_n 0.00501096f $X=1.055 $Y=1.845 $X2=0 $Y2=0
cc_221 N_A_c_302_n N_VPWR_c_389_n 0.00533081f $X=2.915 $Y=1.845 $X2=0 $Y2=0
cc_222 N_A_M1012_g N_VGND_c_432_n 0.0223799f $X=1.04 $Y=0.92 $X2=0 $Y2=0
cc_223 N_A_c_292_n N_VGND_c_432_n 0.00786053f $X=1.115 $Y=0.185 $X2=0 $Y2=0
cc_224 N_A_c_291_n N_VGND_c_433_n 0.0157239f $X=2.645 $Y=0.185 $X2=0 $Y2=0
cc_225 N_A_M1005_g N_VGND_c_433_n 0.0029973f $X=2.9 $Y=1 $X2=0 $Y2=0
cc_226 N_A_c_297_n N_VGND_c_433_n 0.00210171f $X=2.81 $Y=0.185 $X2=0 $Y2=0
cc_227 N_A_c_298_n N_VGND_c_433_n 0.0249987f $X=3.485 $Y=0.462 $X2=0 $Y2=0
cc_228 N_A_c_291_n N_VGND_c_450_n 0.00129982f $X=2.645 $Y=0.185 $X2=0 $Y2=0
cc_229 N_A_M1005_g N_VGND_c_450_n 0.00645394f $X=2.9 $Y=1 $X2=0 $Y2=0
cc_230 N_A_c_297_n N_VGND_c_450_n 0.00419722f $X=2.81 $Y=0.185 $X2=0 $Y2=0
cc_231 N_A_c_298_n N_VGND_c_450_n 0.0125685f $X=3.485 $Y=0.462 $X2=0 $Y2=0
cc_232 N_A_c_292_n N_VGND_c_434_n 0.0430809f $X=1.115 $Y=0.185 $X2=0 $Y2=0
cc_233 N_A_c_291_n N_VGND_c_437_n 0.0122079f $X=2.645 $Y=0.185 $X2=0 $Y2=0
cc_234 N_A_c_298_n N_VGND_c_437_n 0.0712235f $X=3.485 $Y=0.462 $X2=0 $Y2=0
cc_235 N_A_c_291_n N_VGND_c_438_n 0.0536057f $X=2.645 $Y=0.185 $X2=0 $Y2=0
cc_236 N_A_c_292_n N_VGND_c_438_n 0.00750358f $X=1.115 $Y=0.185 $X2=0 $Y2=0
cc_237 N_A_c_297_n N_VGND_c_438_n 0.0102245f $X=2.81 $Y=0.185 $X2=0 $Y2=0
cc_238 N_A_c_298_n N_VGND_c_438_n 0.0393319f $X=3.485 $Y=0.462 $X2=0 $Y2=0
cc_239 X N_VPWR_c_390_n 0.0406301f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_240 X N_VPWR_c_389_n 0.0148166f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_241 X N_VPWR_c_395_n 0.0179404f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_242 N_X_c_368_n N_VGND_c_432_n 0.0171569f $X=0.28 $Y=0.645 $X2=0 $Y2=0
cc_243 N_X_c_368_n N_VGND_c_436_n 0.0103924f $X=0.28 $Y=0.645 $X2=0 $Y2=0
cc_244 N_X_c_368_n N_VGND_c_438_n 0.0121284f $X=0.28 $Y=0.645 $X2=0 $Y2=0
