* File: sky130_fd_sc_ls__o2111a_4.spice
* Created: Fri Aug 28 13:42:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__o2111a_4.pex.spice"
.subckt sky130_fd_sc_ls__o2111a_4  VNB VPB D1 C1 B1 A2 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A2	A2
* B1	B1
* C1	C1
* D1	D1
* VPB	VPB
* VNB	VNB
MM1017 N_A_27_74#_M1017_d N_D1_M1017_g N_A_27_392#_M1017_s VNB NSHORT L=0.15
+ W=0.74 AD=0.2146 AS=0.1036 PD=2.06 PS=1.02 NRD=0.804 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001.5 A=0.111 P=1.78 MULT=1
MM1018 N_A_27_74#_M1018_d N_D1_M1018_g N_A_27_392#_M1017_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1002 N_A_287_74#_M1002_d N_C1_M1002_g N_A_27_74#_M1018_d VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.1 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1012 N_A_287_74#_M1002_d N_C1_M1012_g N_A_27_74#_M1012_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.24285 PD=1.02 PS=2.49 NRD=0 NRS=13.776 M=1 R=4.93333
+ SA=75001.5 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1004 N_A_287_74#_M1004_d N_B1_M1004_g N_A_477_198#_M1004_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.21835 PD=1.02 PS=2.21 NRD=0 NRS=6.48 M=1 R=4.93333
+ SA=75000.2 SB=75001.6 A=0.111 P=1.78 MULT=1
MM1025 N_A_287_74#_M1004_d N_B1_M1025_g N_A_477_198#_M1025_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.7 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1011 N_A_477_198#_M1025_s N_A2_M1011_g N_VGND_M1011_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1258 PD=1.02 PS=1.08 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1026 N_A_477_198#_M1026_d N_A2_M1026_g N_VGND_M1011_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2183 AS=0.1258 PD=2.07 PS=1.08 NRD=1.62 NRS=9.72 M=1 R=4.93333 SA=75001.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1006 N_A_477_198#_M1006_d N_A1_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75002.6 A=0.111 P=1.78 MULT=1
MM1019 N_A_477_198#_M1006_d N_A1_M1019_g N_VGND_M1019_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75002.2 A=0.111 P=1.78 MULT=1
MM1010 N_X_M1010_d N_A_27_392#_M1010_g N_VGND_M1019_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.1
+ SB=75001.7 A=0.111 P=1.78 MULT=1
MM1015 N_X_M1010_d N_A_27_392#_M1015_g N_VGND_M1015_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1554 PD=1.02 PS=1.16 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.6
+ SB=75001.3 A=0.111 P=1.78 MULT=1
MM1020 N_X_M1020_d N_A_27_392#_M1020_g N_VGND_M1015_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1554 PD=1.02 PS=1.16 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75002.1
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1022 N_X_M1020_d N_A_27_392#_M1022_g N_VGND_M1022_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.2627 PD=1.02 PS=2.19 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75002.6
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1021 N_A_27_392#_M1021_d N_D1_M1021_g N_VPWR_M1021_s VPB PHIGHVT L=0.15 W=0.84
+ AD=0.2478 AS=0.168 PD=2.27 PS=1.24 NRD=2.3443 NRS=14.0658 M=1 R=5.6 SA=75000.2
+ SB=75003.9 A=0.126 P=1.98 MULT=1
MM1023 N_A_27_392#_M1023_d N_D1_M1023_g N_VPWR_M1021_s VPB PHIGHVT L=0.15 W=0.84
+ AD=0.126 AS=0.168 PD=1.14 PS=1.24 NRD=2.3443 NRS=14.0658 M=1 R=5.6 SA=75000.8
+ SB=75003.3 A=0.126 P=1.98 MULT=1
MM1003 N_A_27_392#_M1023_d N_C1_M1003_g N_VPWR_M1003_s VPB PHIGHVT L=0.15 W=0.84
+ AD=0.126 AS=0.147 PD=1.14 PS=1.19 NRD=2.3443 NRS=14.0658 M=1 R=5.6 SA=75001.2
+ SB=75002.9 A=0.126 P=1.98 MULT=1
MM1027 N_A_27_392#_M1027_d N_C1_M1027_g N_VPWR_M1003_s VPB PHIGHVT L=0.15 W=0.84
+ AD=0.1974 AS=0.147 PD=1.31 PS=1.19 NRD=22.261 NRS=2.3443 M=1 R=5.6 SA=75001.7
+ SB=75002.4 A=0.126 P=1.98 MULT=1
MM1007 N_VPWR_M1007_d N_B1_M1007_g N_A_27_392#_M1027_d VPB PHIGHVT L=0.15 W=0.84
+ AD=0.126 AS=0.1974 PD=1.14 PS=1.31 NRD=2.3443 NRS=22.261 M=1 R=5.6 SA=75002.3
+ SB=75001.8 A=0.126 P=1.98 MULT=1
MM1013 N_VPWR_M1007_d N_B1_M1013_g N_A_27_392#_M1013_s VPB PHIGHVT L=0.15 W=0.84
+ AD=0.126 AS=0.192013 PD=1.14 PS=1.31022 NRD=2.3443 NRS=22.655 M=1 R=5.6
+ SA=75002.8 SB=75001.3 A=0.126 P=1.98 MULT=1
MM1001 N_A_747_392#_M1001_d N_A2_M1001_g N_A_27_392#_M1013_s VPB PHIGHVT L=0.15
+ W=1 AD=0.175 AS=0.228587 PD=1.35 PS=1.55978 NRD=1.9503 NRS=11.8003 M=1
+ R=6.66667 SA=75002.9 SB=75000.7 A=0.15 P=2.3 MULT=1
MM1005 N_A_747_392#_M1001_d N_A2_M1005_g N_A_27_392#_M1005_s VPB PHIGHVT L=0.15
+ W=1 AD=0.175 AS=0.295 PD=1.35 PS=2.59 NRD=11.8003 NRS=1.9503 M=1 R=6.66667
+ SA=75003.4 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1009 N_A_747_392#_M1009_d N_A1_M1009_g N_VPWR_M1009_s VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.345 PD=1.3 PS=2.69 NRD=1.9503 NRS=11.8003 M=1 R=6.66667
+ SA=75000.3 SB=75002.7 A=0.15 P=2.3 MULT=1
MM1016 N_A_747_392#_M1009_d N_A1_M1016_g N_VPWR_M1016_s VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.196604 PD=1.3 PS=1.41981 NRD=1.9503 NRS=18.715 M=1 R=6.66667
+ SA=75000.7 SB=75002.2 A=0.15 P=2.3 MULT=1
MM1000 N_VPWR_M1016_s N_A_27_392#_M1000_g N_X_M1000_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.220196 AS=0.196 PD=1.59019 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75001.1 SB=75001.7 A=0.168 P=2.54 MULT=1
MM1008 N_VPWR_M1008_d N_A_27_392#_M1008_g N_X_M1000_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.6 SB=75001.2 A=0.168 P=2.54 MULT=1
MM1014 N_VPWR_M1008_d N_A_27_392#_M1014_g N_X_M1014_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.1 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1024 N_VPWR_M1024_d N_A_27_392#_M1024_g N_X_M1014_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3864 AS=0.168 PD=2.93 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75002.5 SB=75000.3 A=0.168 P=2.54 MULT=1
DX28_noxref VNB VPB NWDIODE A=15.8844 P=20.8
c_78 VNB 0 5.23076e-20 $X=0 $Y=0
c_148 VPB 0 1.58594e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_ls__o2111a_4.pxi.spice"
*
.ends
*
*
