# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ls__maj3_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ls__maj3_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.160000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.984000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.800000 1.470000 2.275000 1.800000 ;
        RECT 2.105000 1.800000 2.275000 1.875000 ;
        RECT 2.105000 1.875000 4.570000 2.045000 ;
        RECT 4.240000 1.470000 4.570000 1.875000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.984000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.135000 1.130000 3.235000 1.300000 ;
        RECT 1.135000 1.300000 1.465000 1.705000 ;
        RECT 2.525000 1.300000 3.235000 1.705000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.984000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485000 1.130000 4.925000 1.300000 ;
        RECT 3.485000 1.300000 4.010000 1.705000 ;
        RECT 4.755000 1.300000 4.925000 1.470000 ;
        RECT 4.755000 1.470000 5.220000 1.800000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  1.116000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.365000 1.845000 7.515000 2.015000 ;
        RECT 6.365000 2.015000 6.695000 2.980000 ;
        RECT 6.425000 0.475000 6.675000 1.005000 ;
        RECT 6.425000 1.005000 8.035000 1.175000 ;
        RECT 7.345000 1.480000 8.035000 1.650000 ;
        RECT 7.345000 1.650000 7.515000 1.845000 ;
        RECT 7.345000 2.015000 7.515000 2.980000 ;
        RECT 7.805000 1.175000 8.035000 1.480000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 8.160000 0.085000 ;
        RECT 0.115000  0.085000 0.445000 1.285000 ;
        RECT 2.145000  0.085000 2.315000 0.960000 ;
        RECT 4.005000  0.085000 4.335000 0.620000 ;
        RECT 5.955000  0.085000 6.205000 1.175000 ;
        RECT 6.855000  0.085000 7.185000 0.835000 ;
        RECT 7.715000  0.085000 8.045000 0.835000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
        RECT 6.395000 -0.085000 6.565000 0.085000 ;
        RECT 6.875000 -0.085000 7.045000 0.085000 ;
        RECT 7.355000 -0.085000 7.525000 0.085000 ;
        RECT 7.835000 -0.085000 8.005000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.160000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 8.160000 3.415000 ;
        RECT 0.130000 1.940000 0.380000 3.245000 ;
        RECT 2.060000 2.555000 2.320000 3.245000 ;
        RECT 3.990000 2.555000 4.320000 3.245000 ;
        RECT 5.940000 1.940000 6.190000 3.245000 ;
        RECT 6.895000 2.185000 7.145000 3.245000 ;
        RECT 7.715000 1.820000 8.045000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
        RECT 6.395000 3.245000 6.565000 3.415000 ;
        RECT 6.875000 3.245000 7.045000 3.415000 ;
        RECT 7.355000 3.245000 7.525000 3.415000 ;
        RECT 7.835000 3.245000 8.005000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 8.160000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.580000 2.215000 0.910000 2.905000 ;
      RECT 0.580000 2.905000 1.860000 3.075000 ;
      RECT 0.625000 0.265000 1.965000 0.435000 ;
      RECT 0.625000 0.435000 0.955000 0.620000 ;
      RECT 0.795000 0.790000 1.465000 0.960000 ;
      RECT 0.795000 0.960000 0.965000 1.875000 ;
      RECT 0.795000 1.875000 1.410000 2.045000 ;
      RECT 1.095000 2.045000 1.410000 2.215000 ;
      RECT 1.095000 2.215000 5.290000 2.385000 ;
      RECT 1.095000 2.385000 1.350000 2.735000 ;
      RECT 1.135000 0.605000 1.465000 0.790000 ;
      RECT 1.530000 2.555000 1.860000 2.905000 ;
      RECT 1.635000 0.435000 1.965000 0.960000 ;
      RECT 2.490000 2.555000 2.820000 2.905000 ;
      RECT 2.490000 2.905000 3.820000 3.075000 ;
      RECT 2.495000 0.265000 3.825000 0.435000 ;
      RECT 2.495000 0.435000 2.885000 0.935000 ;
      RECT 2.990000 2.385000 3.320000 2.735000 ;
      RECT 3.065000 0.605000 3.315000 0.790000 ;
      RECT 3.065000 0.790000 5.265000 0.960000 ;
      RECT 3.490000 2.555000 3.820000 2.905000 ;
      RECT 3.495000 0.435000 3.825000 0.620000 ;
      RECT 4.505000 0.255000 5.775000 0.425000 ;
      RECT 4.505000 0.425000 4.835000 0.620000 ;
      RECT 4.510000 2.555000 5.740000 2.725000 ;
      RECT 4.510000 2.725000 4.840000 2.980000 ;
      RECT 4.960000 1.970000 5.560000 2.140000 ;
      RECT 4.960000 2.140000 5.290000 2.215000 ;
      RECT 5.095000 0.595000 5.265000 0.790000 ;
      RECT 5.095000 0.960000 5.265000 1.130000 ;
      RECT 5.095000 1.130000 5.560000 1.300000 ;
      RECT 5.390000 1.300000 5.560000 1.345000 ;
      RECT 5.390000 1.345000 7.150000 1.675000 ;
      RECT 5.390000 1.675000 5.560000 1.970000 ;
      RECT 5.410000 2.725000 5.740000 2.980000 ;
      RECT 5.445000 0.425000 5.775000 0.960000 ;
  END
END sky130_fd_sc_ls__maj3_4
