* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__and4b_1 A_N B C D VGND VNB VPB VPWR X
M1000 VGND D a_526_139# VNB nshort w=640000u l=150000u
+  ad=4.5645e+11p pd=3.97e+06u as=3.418e+11p ps=2.55e+06u
M1001 a_448_139# B a_353_124# VNB nshort w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=2.21125e+11p ps=2.08e+06u
M1002 a_353_124# a_27_74# a_226_424# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1003 X a_226_424# VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1004 VPWR B a_226_424# VPB phighvt w=840000u l=150000u
+  ad=1.6114e+12p pd=9.26e+06u as=6.132e+11p ps=4.82e+06u
M1005 a_226_424# a_27_74# VPWR VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_226_424# C VPWR VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR A_N a_27_74# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=2.478e+11p ps=2.27e+06u
M1008 X a_226_424# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=0p ps=0u
M1009 VPWR D a_226_424# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND A_N a_27_74# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1011 a_526_139# C a_448_139# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
