* File: sky130_fd_sc_ls__nor3b_2.spice
* Created: Wed Sep  2 11:15:10 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__nor3b_2.pex.spice"
.subckt sky130_fd_sc_ls__nor3b_2  VNB VPB C_N B A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* B	B
* C_N	C_N
* VPB	VPB
* VNB	VNB
MM1007 N_VGND_M1007_d N_C_N_M1007_g N_A_27_392#_M1007_s VNB NSHORT L=0.15 W=0.64
+ AD=0.136255 AS=0.1824 PD=1.07594 PS=1.85 NRD=13.116 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75004 A=0.096 P=1.58 MULT=1
MM1000 N_VGND_M1007_d N_A_27_392#_M1000_g N_Y_M1000_s VNB NSHORT L=0.15 W=0.74
+ AD=0.157545 AS=0.10915 PD=1.24406 PS=1.035 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75000.7 SB=75003.4 A=0.111 P=1.78 MULT=1
MM1009 N_VGND_M1009_d N_A_27_392#_M1009_g N_Y_M1000_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2664 AS=0.10915 PD=1.46 PS=1.035 NRD=0 NRS=2.424 M=1 R=4.93333 SA=75001.1
+ SB=75003 A=0.111 P=1.78 MULT=1
MM1002 N_Y_M1002_d N_B_M1002_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.74 AD=0.1036
+ AS=0.2664 PD=1.02 PS=1.46 NRD=0 NRS=0 M=1 R=4.93333 SA=75002 SB=75002.1
+ A=0.111 P=1.78 MULT=1
MM1010 N_Y_M1002_d N_B_M1010_g N_VGND_M1010_s VNB NSHORT L=0.15 W=0.74 AD=0.1036
+ AS=0.3108 PD=1.02 PS=1.58 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.4 SB=75001.7
+ A=0.111 P=1.78 MULT=1
MM1004 N_Y_M1004_d N_A_M1004_g N_VGND_M1010_s VNB NSHORT L=0.15 W=0.74 AD=0.1221
+ AS=0.3108 PD=1.07 PS=1.58 NRD=0 NRS=0 M=1 R=4.93333 SA=75003.4 SB=75000.7
+ A=0.111 P=1.78 MULT=1
MM1005 N_Y_M1004_d N_A_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.74 AD=0.1221
+ AS=0.2257 PD=1.07 PS=2.09 NRD=8.1 NRS=3.24 M=1 R=4.93333 SA=75003.9 SB=75000.2
+ A=0.111 P=1.78 MULT=1
MM1011 N_VPWR_M1011_d N_C_N_M1011_g N_A_27_392#_M1011_s VPB PHIGHVT L=0.15 W=1
+ AD=0.29 AS=0.29 PD=2.58 PS=2.58 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75000.2
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1001 N_A_227_368#_M1001_d N_A_27_392#_M1001_g N_Y_M1001_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.3248 AS=0.168 PD=2.82 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1012 N_A_227_368#_M1012_d N_A_27_392#_M1012_g N_Y_M1001_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1006 N_A_495_368#_M1006_d N_B_M1006_g N_A_227_368#_M1012_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1008 N_A_495_368#_M1006_d N_B_M1008_g N_A_227_368#_M1008_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.3248 PD=1.42 PS=2.82 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.6 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1003 N_VPWR_M1003_d N_A_M1003_g N_A_495_368#_M1003_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3248 AS=0.168 PD=2.82 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1013 N_VPWR_M1013_d N_A_M1013_g N_A_495_368#_M1003_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3248 AS=0.168 PD=2.82 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75000.2 A=0.168 P=2.54 MULT=1
DX14_noxref VNB VPB NWDIODE A=9.6348 P=14.08
*
.include "sky130_fd_sc_ls__nor3b_2.pxi.spice"
*
.ends
*
*
