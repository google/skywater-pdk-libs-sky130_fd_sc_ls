# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ls__a21oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_ls__a21oi_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.240000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.925000 1.350000 3.935000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.785000 1.350000 2.275000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.894000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.235000 1.350000 5.245000 1.780000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.478600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525000 0.595000 2.780000 0.880000 ;
        RECT 2.525000 0.880000 4.650000 1.010000 ;
        RECT 2.525000 1.010000 5.590000 1.180000 ;
        RECT 2.525000 1.180000 2.755000 1.950000 ;
        RECT 2.525000 1.950000 5.585000 2.120000 ;
        RECT 4.355000 2.120000 4.685000 2.735000 ;
        RECT 4.400000 0.350000 4.650000 0.880000 ;
        RECT 5.255000 2.120000 5.585000 2.735000 ;
        RECT 5.340000 0.350000 5.590000 1.010000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.240000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 6.240000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.240000 0.085000 ;
      RECT 0.000000  3.245000 6.240000 3.415000 ;
      RECT 0.305000  1.820000 0.555000 1.950000 ;
      RECT 0.305000  1.950000 2.355000 2.120000 ;
      RECT 0.305000  2.120000 0.555000 2.980000 ;
      RECT 0.380000  0.350000 0.630000 1.010000 ;
      RECT 0.380000  1.010000 2.350000 1.180000 ;
      RECT 0.755000  2.290000 1.005000 3.245000 ;
      RECT 0.810000  0.085000 1.140000 0.840000 ;
      RECT 1.205000  2.120000 1.535000 2.980000 ;
      RECT 1.320000  0.350000 1.490000 1.010000 ;
      RECT 1.670000  0.085000 2.000000 0.840000 ;
      RECT 1.735000  2.290000 1.905000 3.245000 ;
      RECT 2.105000  2.120000 2.355000 2.290000 ;
      RECT 2.105000  2.290000 4.155000 2.460000 ;
      RECT 2.105000  2.460000 2.355000 2.980000 ;
      RECT 2.180000  0.255000 4.150000 0.425000 ;
      RECT 2.180000  0.425000 2.350000 1.010000 ;
      RECT 2.555000  2.630000 2.805000 3.245000 ;
      RECT 2.960000  0.425000 3.290000 0.710000 ;
      RECT 3.005000  2.460000 3.335000 2.980000 ;
      RECT 3.535000  2.630000 3.705000 3.245000 ;
      RECT 3.820000  0.425000 4.150000 0.710000 ;
      RECT 3.905000  2.460000 4.155000 2.905000 ;
      RECT 3.905000  2.905000 6.035000 3.075000 ;
      RECT 4.830000  0.085000 5.160000 0.840000 ;
      RECT 4.885000  2.290000 5.055000 2.905000 ;
      RECT 5.785000  1.820000 6.035000 2.905000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
  END
END sky130_fd_sc_ls__a21oi_4
END LIBRARY
