* File: sky130_fd_sc_ls__a22oi_1.pxi.spice
* Created: Wed Sep  2 10:50:31 2020
* 
x_PM_SKY130_FD_SC_LS__A22OI_1%B2 N_B2_c_49_n N_B2_M1004_g N_B2_M1001_g
+ N_B2_c_46_n N_B2_c_47_n B2 B2 PM_SKY130_FD_SC_LS__A22OI_1%B2
x_PM_SKY130_FD_SC_LS__A22OI_1%B1 N_B1_M1000_g N_B1_c_76_n N_B1_M1007_g B1
+ N_B1_c_77_n PM_SKY130_FD_SC_LS__A22OI_1%B1
x_PM_SKY130_FD_SC_LS__A22OI_1%A1 N_A1_M1003_g N_A1_c_109_n N_A1_M1002_g A1
+ N_A1_c_110_n PM_SKY130_FD_SC_LS__A22OI_1%A1
x_PM_SKY130_FD_SC_LS__A22OI_1%A2 N_A2_M1006_g N_A2_c_137_n N_A2_M1005_g A2 A2
+ PM_SKY130_FD_SC_LS__A22OI_1%A2
x_PM_SKY130_FD_SC_LS__A22OI_1%A_71_368# N_A_71_368#_M1004_s N_A_71_368#_M1007_d
+ N_A_71_368#_M1005_d N_A_71_368#_c_161_n N_A_71_368#_c_162_n
+ N_A_71_368#_c_163_n N_A_71_368#_c_173_n N_A_71_368#_c_170_n
+ N_A_71_368#_c_177_n N_A_71_368#_c_164_n N_A_71_368#_c_165_n
+ PM_SKY130_FD_SC_LS__A22OI_1%A_71_368#
x_PM_SKY130_FD_SC_LS__A22OI_1%Y N_Y_M1000_d N_Y_M1004_d N_Y_c_200_n N_Y_c_201_n
+ N_Y_c_202_n N_Y_c_207_n Y Y PM_SKY130_FD_SC_LS__A22OI_1%Y
x_PM_SKY130_FD_SC_LS__A22OI_1%VPWR N_VPWR_M1002_d N_VPWR_c_239_n N_VPWR_c_240_n
+ N_VPWR_c_241_n VPWR N_VPWR_c_242_n N_VPWR_c_238_n
+ PM_SKY130_FD_SC_LS__A22OI_1%VPWR
x_PM_SKY130_FD_SC_LS__A22OI_1%VGND N_VGND_M1001_s N_VGND_M1006_d N_VGND_c_264_n
+ N_VGND_c_265_n N_VGND_c_266_n N_VGND_c_267_n N_VGND_c_268_n N_VGND_c_269_n
+ VGND N_VGND_c_270_n N_VGND_c_271_n PM_SKY130_FD_SC_LS__A22OI_1%VGND
cc_1 VNB N_B2_c_46_n 0.0856761f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.385
cc_2 VNB N_B2_c_47_n 0.018672f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=1.22
cc_3 VNB B2 0.0170831f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_B1_M1000_g 0.0244201f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=2.4
cc_5 VNB N_B1_c_76_n 0.0262555f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=0.74
cc_6 VNB N_B1_c_77_n 0.00166449f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A1_M1003_g 0.0273876f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=2.4
cc_8 VNB N_A1_c_109_n 0.0262417f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=0.74
cc_9 VNB N_A1_c_110_n 0.00689463f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A2_M1006_g 0.0338413f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=2.4
cc_11 VNB N_A2_c_137_n 0.0273588f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=0.74
cc_12 VNB A2 0.0275005f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=1.22
cc_13 VNB N_Y_c_200_n 0.0155629f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=1.385
cc_14 VNB N_Y_c_201_n 0.0028102f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.385
cc_15 VNB N_Y_c_202_n 0.00336771f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB Y 0.00493162f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.665
cc_17 VNB N_VPWR_c_238_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.665
cc_18 VNB N_VGND_c_264_n 0.0285265f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=1.22
cc_19 VNB N_VGND_c_265_n 0.0419806f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_266_n 0.0129628f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_21 VNB N_VGND_c_267_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_268_n 0.0452046f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_269_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_270_n 0.0129628f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_271_n 0.214622f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VPB N_B2_c_49_n 0.0172401f $X=-0.19 $Y=1.66 $X2=0.705 $Y2=1.765
cc_27 VPB N_B2_c_46_n 0.00717166f $X=-0.19 $Y=1.66 $X2=0.615 $Y2=1.385
cc_28 VPB B2 0.0160072f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_29 VPB N_B1_c_76_n 0.0254599f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=0.74
cc_30 VPB N_B1_c_77_n 0.00482805f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_31 VPB N_A1_c_109_n 0.0281172f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=0.74
cc_32 VPB N_A1_c_110_n 0.0023765f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_33 VPB N_A2_c_137_n 0.0338387f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=0.74
cc_34 VPB A2 0.0171206f $X=-0.19 $Y=1.66 $X2=0.705 $Y2=1.22
cc_35 VPB N_A_71_368#_c_161_n 0.0243557f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_36 VPB N_A_71_368#_c_162_n 0.00567337f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_37 VPB N_A_71_368#_c_163_n 0.00987235f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_38 VPB N_A_71_368#_c_164_n 0.0075508f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.665
cc_39 VPB N_A_71_368#_c_165_n 0.0360166f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_40 VPB Y 0.00457769f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.665
cc_41 VPB N_VPWR_c_239_n 0.00960015f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=0.74
cc_42 VPB N_VPWR_c_240_n 0.044794f $X=-0.19 $Y=1.66 $X2=0.705 $Y2=1.22
cc_43 VPB N_VPWR_c_241_n 0.00670627f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_44 VPB N_VPWR_c_242_n 0.0255159f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_45 VPB N_VPWR_c_238_n 0.0734884f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.665
cc_46 N_B2_c_47_n N_B1_M1000_g 0.0432762f $X=0.705 $Y=1.22 $X2=0 $Y2=0
cc_47 N_B2_c_49_n N_B1_c_76_n 0.0208719f $X=0.705 $Y=1.765 $X2=0 $Y2=0
cc_48 N_B2_c_46_n N_B1_c_76_n 0.0472897f $X=0.615 $Y=1.385 $X2=0 $Y2=0
cc_49 N_B2_c_46_n N_B1_c_77_n 6.4876e-19 $X=0.615 $Y=1.385 $X2=0 $Y2=0
cc_50 N_B2_c_49_n N_A_71_368#_c_161_n 0.00766499f $X=0.705 $Y=1.765 $X2=0 $Y2=0
cc_51 B2 N_A_71_368#_c_161_n 0.00493998f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_52 N_B2_c_49_n N_A_71_368#_c_162_n 0.0107904f $X=0.705 $Y=1.765 $X2=0 $Y2=0
cc_53 N_B2_c_49_n N_A_71_368#_c_163_n 0.00262934f $X=0.705 $Y=1.765 $X2=0 $Y2=0
cc_54 N_B2_c_49_n N_A_71_368#_c_170_n 6.22492e-19 $X=0.705 $Y=1.765 $X2=0 $Y2=0
cc_55 N_B2_c_47_n N_Y_c_201_n 0.0133235f $X=0.705 $Y=1.22 $X2=0 $Y2=0
cc_56 N_B2_c_47_n N_Y_c_202_n 0.00217641f $X=0.705 $Y=1.22 $X2=0 $Y2=0
cc_57 N_B2_c_49_n N_Y_c_207_n 0.0163991f $X=0.705 $Y=1.765 $X2=0 $Y2=0
cc_58 N_B2_c_49_n Y 0.00650251f $X=0.705 $Y=1.765 $X2=0 $Y2=0
cc_59 N_B2_c_46_n Y 0.019953f $X=0.615 $Y=1.385 $X2=0 $Y2=0
cc_60 N_B2_c_47_n Y 0.00119049f $X=0.705 $Y=1.22 $X2=0 $Y2=0
cc_61 B2 Y 0.045939f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_62 N_B2_c_49_n N_VPWR_c_240_n 0.00278257f $X=0.705 $Y=1.765 $X2=0 $Y2=0
cc_63 N_B2_c_49_n N_VPWR_c_238_n 0.00357899f $X=0.705 $Y=1.765 $X2=0 $Y2=0
cc_64 N_B2_c_46_n N_VGND_c_264_n 0.00639332f $X=0.615 $Y=1.385 $X2=0 $Y2=0
cc_65 N_B2_c_47_n N_VGND_c_264_n 0.0154153f $X=0.705 $Y=1.22 $X2=0 $Y2=0
cc_66 B2 N_VGND_c_264_n 0.00521723f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_67 N_B2_c_47_n N_VGND_c_268_n 0.00383152f $X=0.705 $Y=1.22 $X2=0 $Y2=0
cc_68 N_B2_c_47_n N_VGND_c_271_n 0.0075694f $X=0.705 $Y=1.22 $X2=0 $Y2=0
cc_69 N_B1_M1000_g N_A1_M1003_g 0.014794f $X=1.08 $Y=0.74 $X2=0 $Y2=0
cc_70 N_B1_c_76_n N_A1_c_109_n 0.0342241f $X=1.155 $Y=1.765 $X2=0 $Y2=0
cc_71 N_B1_c_77_n N_A1_c_109_n 0.00173907f $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_72 N_B1_c_76_n N_A1_c_110_n 0.00128912f $X=1.155 $Y=1.765 $X2=0 $Y2=0
cc_73 N_B1_c_77_n N_A1_c_110_n 0.0277336f $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_74 N_B1_c_76_n N_A_71_368#_c_161_n 5.7112e-19 $X=1.155 $Y=1.765 $X2=0 $Y2=0
cc_75 N_B1_c_76_n N_A_71_368#_c_162_n 0.0124397f $X=1.155 $Y=1.765 $X2=0 $Y2=0
cc_76 N_B1_c_76_n N_A_71_368#_c_173_n 0.0023562f $X=1.155 $Y=1.765 $X2=0 $Y2=0
cc_77 N_B1_c_77_n N_A_71_368#_c_173_n 0.00785128f $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_78 N_B1_c_76_n N_A_71_368#_c_170_n 0.00919154f $X=1.155 $Y=1.765 $X2=0 $Y2=0
cc_79 N_B1_M1000_g N_Y_c_200_n 0.0124193f $X=1.08 $Y=0.74 $X2=0 $Y2=0
cc_80 N_B1_c_76_n N_Y_c_200_n 0.00140923f $X=1.155 $Y=1.765 $X2=0 $Y2=0
cc_81 N_B1_c_77_n N_Y_c_200_n 0.0265531f $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_82 N_B1_M1000_g N_Y_c_202_n 0.012242f $X=1.08 $Y=0.74 $X2=0 $Y2=0
cc_83 N_B1_c_76_n N_Y_c_207_n 0.00222466f $X=1.155 $Y=1.765 $X2=0 $Y2=0
cc_84 N_B1_c_77_n N_Y_c_207_n 7.202e-19 $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_85 N_B1_M1000_g Y 0.00536895f $X=1.08 $Y=0.74 $X2=0 $Y2=0
cc_86 N_B1_c_76_n Y 0.00172537f $X=1.155 $Y=1.765 $X2=0 $Y2=0
cc_87 N_B1_c_77_n Y 0.0334882f $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_88 N_B1_c_76_n N_VPWR_c_240_n 0.00278257f $X=1.155 $Y=1.765 $X2=0 $Y2=0
cc_89 N_B1_c_76_n N_VPWR_c_238_n 0.00354252f $X=1.155 $Y=1.765 $X2=0 $Y2=0
cc_90 N_B1_M1000_g N_VGND_c_264_n 0.00190254f $X=1.08 $Y=0.74 $X2=0 $Y2=0
cc_91 N_B1_M1000_g N_VGND_c_268_n 0.00434272f $X=1.08 $Y=0.74 $X2=0 $Y2=0
cc_92 N_B1_M1000_g N_VGND_c_271_n 0.00821699f $X=1.08 $Y=0.74 $X2=0 $Y2=0
cc_93 N_A1_M1003_g N_A2_M1006_g 0.0328884f $X=1.62 $Y=0.74 $X2=0 $Y2=0
cc_94 N_A1_c_109_n N_A2_c_137_n 0.0493383f $X=1.635 $Y=1.765 $X2=0 $Y2=0
cc_95 N_A1_c_110_n N_A2_c_137_n 7.1218e-19 $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_96 N_A1_c_109_n A2 0.00230997f $X=1.635 $Y=1.765 $X2=0 $Y2=0
cc_97 N_A1_c_110_n A2 0.0366314f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_98 N_A1_c_109_n N_A_71_368#_c_162_n 0.00108743f $X=1.635 $Y=1.765 $X2=0 $Y2=0
cc_99 N_A1_c_109_n N_A_71_368#_c_177_n 0.0142429f $X=1.635 $Y=1.765 $X2=0 $Y2=0
cc_100 N_A1_c_110_n N_A_71_368#_c_177_n 0.0226207f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_101 N_A1_c_109_n N_A_71_368#_c_165_n 8.4516e-19 $X=1.635 $Y=1.765 $X2=0 $Y2=0
cc_102 N_A1_M1003_g N_Y_c_200_n 0.00484582f $X=1.62 $Y=0.74 $X2=0 $Y2=0
cc_103 N_A1_c_110_n N_Y_c_200_n 0.00196319f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_104 N_A1_M1003_g N_Y_c_202_n 0.0144523f $X=1.62 $Y=0.74 $X2=0 $Y2=0
cc_105 N_A1_c_109_n N_VPWR_c_239_n 0.00156185f $X=1.635 $Y=1.765 $X2=0 $Y2=0
cc_106 N_A1_c_109_n N_VPWR_c_240_n 0.00461464f $X=1.635 $Y=1.765 $X2=0 $Y2=0
cc_107 N_A1_c_109_n N_VPWR_c_238_n 0.00908785f $X=1.635 $Y=1.765 $X2=0 $Y2=0
cc_108 N_A1_M1003_g N_VGND_c_265_n 0.00294701f $X=1.62 $Y=0.74 $X2=0 $Y2=0
cc_109 N_A1_M1003_g N_VGND_c_268_n 0.00434272f $X=1.62 $Y=0.74 $X2=0 $Y2=0
cc_110 N_A1_M1003_g N_VGND_c_271_n 0.00823328f $X=1.62 $Y=0.74 $X2=0 $Y2=0
cc_111 N_A2_c_137_n N_A_71_368#_c_177_n 0.0124074f $X=2.175 $Y=1.765 $X2=0 $Y2=0
cc_112 A2 N_A_71_368#_c_177_n 0.0121995f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_113 N_A2_c_137_n N_A_71_368#_c_164_n 0.00124634f $X=2.175 $Y=1.765 $X2=0
+ $Y2=0
cc_114 A2 N_A_71_368#_c_164_n 0.0265363f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_115 N_A2_c_137_n N_A_71_368#_c_165_n 0.0103816f $X=2.175 $Y=1.765 $X2=0 $Y2=0
cc_116 N_A2_M1006_g N_Y_c_200_n 6.02297e-19 $X=2.16 $Y=0.74 $X2=0 $Y2=0
cc_117 N_A2_M1006_g N_Y_c_202_n 0.00204985f $X=2.16 $Y=0.74 $X2=0 $Y2=0
cc_118 N_A2_c_137_n N_VPWR_c_239_n 0.00731029f $X=2.175 $Y=1.765 $X2=0 $Y2=0
cc_119 N_A2_c_137_n N_VPWR_c_242_n 0.00445602f $X=2.175 $Y=1.765 $X2=0 $Y2=0
cc_120 N_A2_c_137_n N_VPWR_c_238_n 0.00861742f $X=2.175 $Y=1.765 $X2=0 $Y2=0
cc_121 N_A2_M1006_g N_VGND_c_265_n 0.022716f $X=2.16 $Y=0.74 $X2=0 $Y2=0
cc_122 N_A2_c_137_n N_VGND_c_265_n 0.00415604f $X=2.175 $Y=1.765 $X2=0 $Y2=0
cc_123 A2 N_VGND_c_265_n 0.0236581f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_124 N_A2_M1006_g N_VGND_c_268_n 0.00383152f $X=2.16 $Y=0.74 $X2=0 $Y2=0
cc_125 N_A2_M1006_g N_VGND_c_271_n 0.00758569f $X=2.16 $Y=0.74 $X2=0 $Y2=0
cc_126 N_A_71_368#_c_162_n N_Y_M1004_d 0.00247267f $X=1.215 $Y=2.99 $X2=0 $Y2=0
cc_127 N_A_71_368#_c_161_n N_Y_c_207_n 0.0300102f $X=0.48 $Y=2.455 $X2=0 $Y2=0
cc_128 N_A_71_368#_c_162_n N_Y_c_207_n 0.0126885f $X=1.215 $Y=2.99 $X2=0 $Y2=0
cc_129 N_A_71_368#_c_173_n N_Y_c_207_n 0.0124534f $X=1.38 $Y=2.12 $X2=0 $Y2=0
cc_130 N_A_71_368#_c_170_n N_Y_c_207_n 0.0400262f $X=1.38 $Y=2.815 $X2=0 $Y2=0
cc_131 N_A_71_368#_c_177_n N_VPWR_M1002_d 0.010589f $X=2.235 $Y=2.035 $X2=-0.19
+ $Y2=1.66
cc_132 N_A_71_368#_c_162_n N_VPWR_c_239_n 0.0101198f $X=1.215 $Y=2.99 $X2=0
+ $Y2=0
cc_133 N_A_71_368#_c_177_n N_VPWR_c_239_n 0.022455f $X=2.235 $Y=2.035 $X2=0
+ $Y2=0
cc_134 N_A_71_368#_c_165_n N_VPWR_c_239_n 0.026688f $X=2.4 $Y=2.815 $X2=0 $Y2=0
cc_135 N_A_71_368#_c_162_n N_VPWR_c_240_n 0.0594839f $X=1.215 $Y=2.99 $X2=0
+ $Y2=0
cc_136 N_A_71_368#_c_163_n N_VPWR_c_240_n 0.0236039f $X=0.645 $Y=2.99 $X2=0
+ $Y2=0
cc_137 N_A_71_368#_c_165_n N_VPWR_c_242_n 0.0145938f $X=2.4 $Y=2.815 $X2=0 $Y2=0
cc_138 N_A_71_368#_c_162_n N_VPWR_c_238_n 0.0329562f $X=1.215 $Y=2.99 $X2=0
+ $Y2=0
cc_139 N_A_71_368#_c_163_n N_VPWR_c_238_n 0.012761f $X=0.645 $Y=2.99 $X2=0 $Y2=0
cc_140 N_A_71_368#_c_165_n N_VPWR_c_238_n 0.0120466f $X=2.4 $Y=2.815 $X2=0 $Y2=0
cc_141 N_Y_c_201_n N_VGND_c_264_n 0.0019893f $X=0.835 $Y=1.095 $X2=0 $Y2=0
cc_142 N_Y_c_202_n N_VGND_c_264_n 0.0167629f $X=1.35 $Y=0.515 $X2=0 $Y2=0
cc_143 N_Y_c_200_n N_VGND_c_265_n 0.00316703f $X=1.13 $Y=1.095 $X2=0 $Y2=0
cc_144 N_Y_c_202_n N_VGND_c_265_n 0.0167858f $X=1.35 $Y=0.515 $X2=0 $Y2=0
cc_145 N_Y_c_202_n N_VGND_c_268_n 0.0194005f $X=1.35 $Y=0.515 $X2=0 $Y2=0
cc_146 N_Y_c_202_n N_VGND_c_271_n 0.0159453f $X=1.35 $Y=0.515 $X2=0 $Y2=0
cc_147 N_Y_c_200_n A_159_74# 0.00366293f $X=1.13 $Y=1.095 $X2=-0.19 $Y2=-0.245
