* File: sky130_fd_sc_ls__nor2_4.pxi.spice
* Created: Wed Sep  2 11:14:05 2020
* 
x_PM_SKY130_FD_SC_LS__NOR2_4%A N_A_c_54_n N_A_M1000_g N_A_c_50_n N_A_M1001_g
+ N_A_c_55_n N_A_M1007_g N_A_c_56_n N_A_M1008_g N_A_c_51_n N_A_M1003_g
+ N_A_c_57_n N_A_M1010_g A A A A N_A_c_53_n PM_SKY130_FD_SC_LS__NOR2_4%A
x_PM_SKY130_FD_SC_LS__NOR2_4%B N_B_c_119_n N_B_M1004_g N_B_c_123_n N_B_M1002_g
+ N_B_c_120_n N_B_M1006_g N_B_c_124_n N_B_M1005_g N_B_c_125_n N_B_M1009_g
+ N_B_c_126_n N_B_M1011_g B B B N_B_c_122_n PM_SKY130_FD_SC_LS__NOR2_4%B
x_PM_SKY130_FD_SC_LS__NOR2_4%A_27_368# N_A_27_368#_M1000_d N_A_27_368#_M1007_d
+ N_A_27_368#_M1010_d N_A_27_368#_M1005_s N_A_27_368#_M1011_s
+ N_A_27_368#_c_181_n N_A_27_368#_c_182_n N_A_27_368#_c_183_n
+ N_A_27_368#_c_184_n N_A_27_368#_c_185_n N_A_27_368#_c_209_n
+ N_A_27_368#_c_186_n N_A_27_368#_c_187_n N_A_27_368#_c_220_n
+ N_A_27_368#_c_188_n N_A_27_368#_c_189_n N_A_27_368#_c_190_n
+ N_A_27_368#_c_191_n PM_SKY130_FD_SC_LS__NOR2_4%A_27_368#
x_PM_SKY130_FD_SC_LS__NOR2_4%VPWR N_VPWR_M1000_s N_VPWR_M1008_s N_VPWR_c_258_n
+ N_VPWR_c_259_n VPWR N_VPWR_c_260_n N_VPWR_c_261_n N_VPWR_c_257_n
+ N_VPWR_c_263_n N_VPWR_c_264_n PM_SKY130_FD_SC_LS__NOR2_4%VPWR
x_PM_SKY130_FD_SC_LS__NOR2_4%Y N_Y_M1001_s N_Y_M1004_d N_Y_M1002_d N_Y_M1009_d
+ N_Y_c_306_n N_Y_c_313_n N_Y_c_307_n N_Y_c_316_n N_Y_c_319_n N_Y_c_321_n
+ N_Y_c_309_n N_Y_c_340_n N_Y_c_308_n N_Y_c_341_n Y PM_SKY130_FD_SC_LS__NOR2_4%Y
x_PM_SKY130_FD_SC_LS__NOR2_4%VGND N_VGND_M1001_d N_VGND_M1003_d N_VGND_M1006_s
+ N_VGND_c_363_n N_VGND_c_364_n N_VGND_c_365_n N_VGND_c_366_n N_VGND_c_367_n
+ VGND N_VGND_c_368_n N_VGND_c_369_n N_VGND_c_370_n
+ PM_SKY130_FD_SC_LS__NOR2_4%VGND
cc_1 VNB N_A_c_50_n 0.0266014f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.22
cc_2 VNB N_A_c_51_n 0.0227304f $X=-0.19 $Y=-0.245 $X2=1.81 $Y2=1.22
cc_3 VNB A 0.0340492f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.21
cc_4 VNB N_A_c_53_n 0.132371f $X=-0.19 $Y=-0.245 $X2=1.81 $Y2=1.492
cc_5 VNB N_B_c_119_n 0.0176155f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_6 VNB N_B_c_120_n 0.0197009f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.765
cc_7 VNB B 0.0270754f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.21
cc_8 VNB N_B_c_122_n 0.174083f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=1.492
cc_9 VNB N_VPWR_c_257_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.492
cc_10 VNB N_Y_c_306_n 0.00695126f $X=-0.19 $Y=-0.245 $X2=1.81 $Y2=1.22
cc_11 VNB N_Y_c_307_n 0.00257348f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.21
cc_12 VNB N_Y_c_308_n 0.00334407f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_VGND_c_363_n 0.0125081f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=1.765
cc_14 VNB N_VGND_c_364_n 0.0352733f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=2.4
cc_15 VNB N_VGND_c_365_n 0.00571115f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=1.765
cc_16 VNB N_VGND_c_366_n 0.0355045f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_17 VNB N_VGND_c_367_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_18 VNB N_VGND_c_368_n 0.0186748f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.385
cc_19 VNB N_VGND_c_369_n 0.082553f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.365
cc_20 VNB N_VGND_c_370_n 0.244311f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VPB N_A_c_54_n 0.0194221f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_22 VPB N_A_c_55_n 0.0149585f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.765
cc_23 VPB N_A_c_56_n 0.0149585f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=1.765
cc_24 VPB N_A_c_57_n 0.0145947f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=1.765
cc_25 VPB N_A_c_53_n 0.0269559f $X=-0.19 $Y=1.66 $X2=1.81 $Y2=1.492
cc_26 VPB N_B_c_123_n 0.0145648f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.22
cc_27 VPB N_B_c_124_n 0.0144861f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=1.765
cc_28 VPB N_B_c_125_n 0.0148581f $X=-0.19 $Y=1.66 $X2=1.81 $Y2=1.22
cc_29 VPB N_B_c_126_n 0.0184944f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=1.765
cc_30 VPB N_B_c_122_n 0.0291543f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=1.492
cc_31 VPB N_A_27_368#_c_181_n 0.0441294f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=2.4
cc_32 VPB N_A_27_368#_c_182_n 0.00219429f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.21
cc_33 VPB N_A_27_368#_c_183_n 0.0106238f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_34 VPB N_A_27_368#_c_184_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_35 VPB N_A_27_368#_c_185_n 0.0133426f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.385
cc_36 VPB N_A_27_368#_c_186_n 0.0026202f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=1.492
cc_37 VPB N_A_27_368#_c_187_n 0.00192911f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.365
cc_38 VPB N_A_27_368#_c_188_n 0.0100303f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_39 VPB N_A_27_368#_c_189_n 0.00313705f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_40 VPB N_A_27_368#_c_190_n 0.00224287f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_41 VPB N_A_27_368#_c_191_n 0.0022931f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_42 VPB N_VPWR_c_258_n 0.00799266f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=2.4
cc_43 VPB N_VPWR_c_259_n 0.00769929f $X=-0.19 $Y=1.66 $X2=1.81 $Y2=0.74
cc_44 VPB N_VPWR_c_260_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_45 VPB N_VPWR_c_261_n 0.0633842f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_257_n 0.0748263f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.492
cc_47 VPB N_VPWR_c_263_n 0.0233502f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.385
cc_48 VPB N_VPWR_c_264_n 0.00324402f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=1.492
cc_49 VPB N_Y_c_309_n 0.0075476f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.385
cc_50 N_A_c_51_n N_B_c_119_n 0.0145322f $X=1.81 $Y=1.22 $X2=-0.19 $Y2=-0.245
cc_51 A N_B_c_119_n 0.0014455f $X=1.595 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_52 N_A_c_57_n N_B_c_123_n 0.00991615f $X=1.855 $Y=1.765 $X2=0 $Y2=0
cc_53 N_A_c_53_n N_B_c_122_n 0.0328797f $X=1.81 $Y=1.492 $X2=0 $Y2=0
cc_54 N_A_c_54_n N_A_27_368#_c_181_n 0.0138448f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_55 N_A_c_55_n N_A_27_368#_c_181_n 7.15508e-19 $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_56 N_A_c_54_n N_A_27_368#_c_182_n 0.00903574f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_57 N_A_c_55_n N_A_27_368#_c_182_n 0.00903574f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_58 A N_A_27_368#_c_182_n 0.042029f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_59 N_A_c_53_n N_A_27_368#_c_182_n 0.00885373f $X=1.81 $Y=1.492 $X2=0 $Y2=0
cc_60 N_A_c_54_n N_A_27_368#_c_183_n 0.00165632f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_61 A N_A_27_368#_c_183_n 0.0282802f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_62 N_A_c_53_n N_A_27_368#_c_183_n 0.00184192f $X=1.81 $Y=1.492 $X2=0 $Y2=0
cc_63 N_A_c_54_n N_A_27_368#_c_184_n 7.15508e-19 $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_64 N_A_c_55_n N_A_27_368#_c_184_n 0.0133148f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_65 N_A_c_56_n N_A_27_368#_c_184_n 0.0133148f $X=1.405 $Y=1.765 $X2=0 $Y2=0
cc_66 N_A_c_57_n N_A_27_368#_c_184_n 7.15508e-19 $X=1.855 $Y=1.765 $X2=0 $Y2=0
cc_67 N_A_c_56_n N_A_27_368#_c_185_n 0.00899835f $X=1.405 $Y=1.765 $X2=0 $Y2=0
cc_68 N_A_c_57_n N_A_27_368#_c_185_n 0.00995664f $X=1.855 $Y=1.765 $X2=0 $Y2=0
cc_69 A N_A_27_368#_c_185_n 0.0334139f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_70 N_A_c_53_n N_A_27_368#_c_185_n 0.0148117f $X=1.81 $Y=1.492 $X2=0 $Y2=0
cc_71 N_A_c_56_n N_A_27_368#_c_209_n 6.9401e-19 $X=1.405 $Y=1.765 $X2=0 $Y2=0
cc_72 N_A_c_57_n N_A_27_368#_c_209_n 0.0120434f $X=1.855 $Y=1.765 $X2=0 $Y2=0
cc_73 N_A_c_57_n N_A_27_368#_c_187_n 0.0032261f $X=1.855 $Y=1.765 $X2=0 $Y2=0
cc_74 N_A_c_55_n N_A_27_368#_c_190_n 0.00109449f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_75 N_A_c_56_n N_A_27_368#_c_190_n 0.00109449f $X=1.405 $Y=1.765 $X2=0 $Y2=0
cc_76 A N_A_27_368#_c_190_n 0.0277828f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_77 N_A_c_53_n N_A_27_368#_c_190_n 0.00501057f $X=1.81 $Y=1.492 $X2=0 $Y2=0
cc_78 N_A_c_54_n N_VPWR_c_258_n 0.00646778f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_79 N_A_c_55_n N_VPWR_c_258_n 0.00646778f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_80 N_A_c_56_n N_VPWR_c_259_n 0.00646778f $X=1.405 $Y=1.765 $X2=0 $Y2=0
cc_81 N_A_c_57_n N_VPWR_c_259_n 0.00491805f $X=1.855 $Y=1.765 $X2=0 $Y2=0
cc_82 N_A_c_55_n N_VPWR_c_260_n 0.00445602f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_83 N_A_c_56_n N_VPWR_c_260_n 0.00445602f $X=1.405 $Y=1.765 $X2=0 $Y2=0
cc_84 N_A_c_57_n N_VPWR_c_261_n 0.0044313f $X=1.855 $Y=1.765 $X2=0 $Y2=0
cc_85 N_A_c_54_n N_VPWR_c_257_n 0.00861084f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_86 N_A_c_55_n N_VPWR_c_257_n 0.00857589f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_87 N_A_c_56_n N_VPWR_c_257_n 0.00857589f $X=1.405 $Y=1.765 $X2=0 $Y2=0
cc_88 N_A_c_57_n N_VPWR_c_257_n 0.00853445f $X=1.855 $Y=1.765 $X2=0 $Y2=0
cc_89 N_A_c_54_n N_VPWR_c_263_n 0.00445602f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_90 N_A_c_50_n N_Y_c_306_n 6.72669e-19 $X=0.52 $Y=1.22 $X2=0 $Y2=0
cc_91 A N_Y_c_306_n 0.0963567f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_92 N_A_c_53_n N_Y_c_306_n 0.00672202f $X=1.81 $Y=1.492 $X2=0 $Y2=0
cc_93 N_A_c_51_n N_Y_c_313_n 0.0125972f $X=1.81 $Y=1.22 $X2=0 $Y2=0
cc_94 N_A_c_53_n N_Y_c_313_n 0.00114846f $X=1.81 $Y=1.492 $X2=0 $Y2=0
cc_95 N_A_c_51_n N_Y_c_307_n 4.29877e-19 $X=1.81 $Y=1.22 $X2=0 $Y2=0
cc_96 N_A_c_51_n N_Y_c_316_n 8.96662e-19 $X=1.81 $Y=1.22 $X2=0 $Y2=0
cc_97 A N_Y_c_316_n 0.00679233f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_98 N_A_c_53_n N_Y_c_316_n 7.28848e-19 $X=1.81 $Y=1.492 $X2=0 $Y2=0
cc_99 A N_Y_c_319_n 0.00406857f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_100 N_A_c_53_n N_Y_c_319_n 0.00132707f $X=1.81 $Y=1.492 $X2=0 $Y2=0
cc_101 N_A_c_57_n N_Y_c_321_n 2.4281e-19 $X=1.855 $Y=1.765 $X2=0 $Y2=0
cc_102 N_A_c_51_n N_Y_c_308_n 6.72669e-19 $X=1.81 $Y=1.22 $X2=0 $Y2=0
cc_103 N_A_c_50_n N_VGND_c_364_n 0.0148927f $X=0.52 $Y=1.22 $X2=0 $Y2=0
cc_104 A N_VGND_c_364_n 0.0273236f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_105 N_A_c_51_n N_VGND_c_365_n 0.0100967f $X=1.81 $Y=1.22 $X2=0 $Y2=0
cc_106 N_A_c_50_n N_VGND_c_366_n 0.00383152f $X=0.52 $Y=1.22 $X2=0 $Y2=0
cc_107 N_A_c_51_n N_VGND_c_366_n 0.00383152f $X=1.81 $Y=1.22 $X2=0 $Y2=0
cc_108 N_A_c_50_n N_VGND_c_370_n 0.00762539f $X=0.52 $Y=1.22 $X2=0 $Y2=0
cc_109 N_A_c_51_n N_VGND_c_370_n 0.00388966f $X=1.81 $Y=1.22 $X2=0 $Y2=0
cc_110 N_B_c_123_n N_A_27_368#_c_185_n 6.42063e-19 $X=2.305 $Y=1.765 $X2=0 $Y2=0
cc_111 N_B_c_122_n N_A_27_368#_c_185_n 3.92385e-19 $X=3.755 $Y=1.492 $X2=0 $Y2=0
cc_112 N_B_c_123_n N_A_27_368#_c_186_n 0.0127563f $X=2.305 $Y=1.765 $X2=0 $Y2=0
cc_113 N_B_c_124_n N_A_27_368#_c_186_n 0.0138537f $X=2.755 $Y=1.765 $X2=0 $Y2=0
cc_114 N_B_c_125_n N_A_27_368#_c_220_n 0.0098831f $X=3.255 $Y=1.765 $X2=0 $Y2=0
cc_115 N_B_c_126_n N_A_27_368#_c_220_n 2.69714e-19 $X=3.755 $Y=1.765 $X2=0 $Y2=0
cc_116 N_B_c_125_n N_A_27_368#_c_188_n 0.0111147f $X=3.255 $Y=1.765 $X2=0 $Y2=0
cc_117 N_B_c_126_n N_A_27_368#_c_188_n 0.0139336f $X=3.755 $Y=1.765 $X2=0 $Y2=0
cc_118 N_B_c_126_n N_A_27_368#_c_189_n 0.00143221f $X=3.755 $Y=1.765 $X2=0 $Y2=0
cc_119 B N_A_27_368#_c_189_n 0.0167379f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_120 N_B_c_122_n N_A_27_368#_c_189_n 0.00612431f $X=3.755 $Y=1.492 $X2=0 $Y2=0
cc_121 N_B_c_125_n N_A_27_368#_c_191_n 0.00193739f $X=3.255 $Y=1.765 $X2=0 $Y2=0
cc_122 N_B_c_123_n N_VPWR_c_261_n 0.00278271f $X=2.305 $Y=1.765 $X2=0 $Y2=0
cc_123 N_B_c_124_n N_VPWR_c_261_n 0.00278271f $X=2.755 $Y=1.765 $X2=0 $Y2=0
cc_124 N_B_c_125_n N_VPWR_c_261_n 0.00278257f $X=3.255 $Y=1.765 $X2=0 $Y2=0
cc_125 N_B_c_126_n N_VPWR_c_261_n 0.00278271f $X=3.755 $Y=1.765 $X2=0 $Y2=0
cc_126 N_B_c_123_n N_VPWR_c_257_n 0.00353907f $X=2.305 $Y=1.765 $X2=0 $Y2=0
cc_127 N_B_c_124_n N_VPWR_c_257_n 0.00354284f $X=2.755 $Y=1.765 $X2=0 $Y2=0
cc_128 N_B_c_125_n N_VPWR_c_257_n 0.00354744f $X=3.255 $Y=1.765 $X2=0 $Y2=0
cc_129 N_B_c_126_n N_VPWR_c_257_n 0.00357961f $X=3.755 $Y=1.765 $X2=0 $Y2=0
cc_130 N_B_c_119_n N_Y_c_313_n 0.0142112f $X=2.29 $Y=1.22 $X2=0 $Y2=0
cc_131 N_B_c_119_n N_Y_c_307_n 0.00694939f $X=2.29 $Y=1.22 $X2=0 $Y2=0
cc_132 N_B_c_120_n N_Y_c_307_n 0.00644058f $X=2.74 $Y=1.22 $X2=0 $Y2=0
cc_133 N_B_c_119_n N_Y_c_316_n 0.00476825f $X=2.29 $Y=1.22 $X2=0 $Y2=0
cc_134 N_B_c_120_n N_Y_c_316_n 0.0142151f $X=2.74 $Y=1.22 $X2=0 $Y2=0
cc_135 B N_Y_c_316_n 0.0137784f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_136 N_B_c_122_n N_Y_c_316_n 0.0174866f $X=3.755 $Y=1.492 $X2=0 $Y2=0
cc_137 B N_Y_c_319_n 0.00682348f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_138 N_B_c_122_n N_Y_c_319_n 0.0228046f $X=3.755 $Y=1.492 $X2=0 $Y2=0
cc_139 N_B_c_123_n N_Y_c_321_n 0.00816264f $X=2.305 $Y=1.765 $X2=0 $Y2=0
cc_140 N_B_c_124_n N_Y_c_321_n 0.00988022f $X=2.755 $Y=1.765 $X2=0 $Y2=0
cc_141 N_B_c_125_n N_Y_c_321_n 2.69714e-19 $X=3.255 $Y=1.765 $X2=0 $Y2=0
cc_142 N_B_c_124_n N_Y_c_309_n 0.0092358f $X=2.755 $Y=1.765 $X2=0 $Y2=0
cc_143 N_B_c_125_n N_Y_c_309_n 0.0114577f $X=3.255 $Y=1.765 $X2=0 $Y2=0
cc_144 N_B_c_126_n N_Y_c_309_n 0.00424884f $X=3.755 $Y=1.765 $X2=0 $Y2=0
cc_145 B N_Y_c_309_n 0.0545029f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_146 N_B_c_122_n N_Y_c_309_n 0.0223156f $X=3.755 $Y=1.492 $X2=0 $Y2=0
cc_147 N_B_c_126_n N_Y_c_340_n 0.00859466f $X=3.755 $Y=1.765 $X2=0 $Y2=0
cc_148 N_B_c_123_n N_Y_c_341_n 0.00210583f $X=2.305 $Y=1.765 $X2=0 $Y2=0
cc_149 N_B_c_124_n N_Y_c_341_n 0.00109449f $X=2.755 $Y=1.765 $X2=0 $Y2=0
cc_150 N_B_c_122_n N_Y_c_341_n 0.00243129f $X=3.755 $Y=1.492 $X2=0 $Y2=0
cc_151 N_B_c_119_n N_VGND_c_365_n 0.00191937f $X=2.29 $Y=1.22 $X2=0 $Y2=0
cc_152 N_B_c_119_n N_VGND_c_368_n 0.00456932f $X=2.29 $Y=1.22 $X2=0 $Y2=0
cc_153 N_B_c_120_n N_VGND_c_368_n 0.00434272f $X=2.74 $Y=1.22 $X2=0 $Y2=0
cc_154 N_B_c_120_n N_VGND_c_369_n 0.00394517f $X=2.74 $Y=1.22 $X2=0 $Y2=0
cc_155 B N_VGND_c_369_n 0.104047f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_156 N_B_c_122_n N_VGND_c_369_n 0.0144527f $X=3.755 $Y=1.492 $X2=0 $Y2=0
cc_157 N_B_c_119_n N_VGND_c_370_n 0.00455422f $X=2.29 $Y=1.22 $X2=0 $Y2=0
cc_158 N_B_c_120_n N_VGND_c_370_n 0.00825234f $X=2.74 $Y=1.22 $X2=0 $Y2=0
cc_159 N_A_27_368#_c_182_n N_VPWR_M1000_s 0.00247267f $X=1.015 $Y=1.805
+ $X2=-0.19 $Y2=1.66
cc_160 N_A_27_368#_c_185_n N_VPWR_M1008_s 0.00247267f $X=1.915 $Y=1.805 $X2=0
+ $Y2=0
cc_161 N_A_27_368#_c_181_n N_VPWR_c_258_n 0.0599532f $X=0.28 $Y=1.985 $X2=0
+ $Y2=0
cc_162 N_A_27_368#_c_182_n N_VPWR_c_258_n 0.0136682f $X=1.015 $Y=1.805 $X2=0
+ $Y2=0
cc_163 N_A_27_368#_c_184_n N_VPWR_c_258_n 0.0599532f $X=1.18 $Y=1.985 $X2=0
+ $Y2=0
cc_164 N_A_27_368#_c_184_n N_VPWR_c_259_n 0.0599532f $X=1.18 $Y=1.985 $X2=0
+ $Y2=0
cc_165 N_A_27_368#_c_185_n N_VPWR_c_259_n 0.0136682f $X=1.915 $Y=1.805 $X2=0
+ $Y2=0
cc_166 N_A_27_368#_c_209_n N_VPWR_c_259_n 0.0543166f $X=2.08 $Y=1.985 $X2=0
+ $Y2=0
cc_167 N_A_27_368#_c_187_n N_VPWR_c_259_n 0.0119328f $X=2.195 $Y=2.99 $X2=0
+ $Y2=0
cc_168 N_A_27_368#_c_184_n N_VPWR_c_260_n 0.014552f $X=1.18 $Y=1.985 $X2=0 $Y2=0
cc_169 N_A_27_368#_c_186_n N_VPWR_c_261_n 0.0422287f $X=2.865 $Y=2.99 $X2=0
+ $Y2=0
cc_170 N_A_27_368#_c_187_n N_VPWR_c_261_n 0.0200196f $X=2.195 $Y=2.99 $X2=0
+ $Y2=0
cc_171 N_A_27_368#_c_188_n N_VPWR_c_261_n 0.0623475f $X=3.865 $Y=2.99 $X2=0
+ $Y2=0
cc_172 N_A_27_368#_c_191_n N_VPWR_c_261_n 0.0236039f $X=3.03 $Y=2.99 $X2=0 $Y2=0
cc_173 N_A_27_368#_c_181_n N_VPWR_c_257_n 0.0120466f $X=0.28 $Y=1.985 $X2=0
+ $Y2=0
cc_174 N_A_27_368#_c_184_n N_VPWR_c_257_n 0.0119791f $X=1.18 $Y=1.985 $X2=0
+ $Y2=0
cc_175 N_A_27_368#_c_186_n N_VPWR_c_257_n 0.0238173f $X=2.865 $Y=2.99 $X2=0
+ $Y2=0
cc_176 N_A_27_368#_c_187_n N_VPWR_c_257_n 0.0108171f $X=2.195 $Y=2.99 $X2=0
+ $Y2=0
cc_177 N_A_27_368#_c_188_n N_VPWR_c_257_n 0.0347719f $X=3.865 $Y=2.99 $X2=0
+ $Y2=0
cc_178 N_A_27_368#_c_191_n N_VPWR_c_257_n 0.012761f $X=3.03 $Y=2.99 $X2=0 $Y2=0
cc_179 N_A_27_368#_c_181_n N_VPWR_c_263_n 0.0145938f $X=0.28 $Y=1.985 $X2=0
+ $Y2=0
cc_180 N_A_27_368#_c_186_n N_Y_M1002_d 0.00197722f $X=2.865 $Y=2.99 $X2=0 $Y2=0
cc_181 N_A_27_368#_c_188_n N_Y_M1009_d 0.00250873f $X=3.865 $Y=2.99 $X2=0 $Y2=0
cc_182 N_A_27_368#_c_186_n N_Y_c_321_n 0.0160777f $X=2.865 $Y=2.99 $X2=0 $Y2=0
cc_183 N_A_27_368#_M1005_s N_Y_c_309_n 0.00250873f $X=2.83 $Y=1.84 $X2=0 $Y2=0
cc_184 N_A_27_368#_c_220_n N_Y_c_309_n 0.0202249f $X=3.03 $Y=2.145 $X2=0 $Y2=0
cc_185 N_A_27_368#_c_189_n N_Y_c_309_n 0.00372299f $X=3.98 $Y=1.985 $X2=0 $Y2=0
cc_186 N_A_27_368#_c_188_n N_Y_c_340_n 0.018923f $X=3.865 $Y=2.99 $X2=0 $Y2=0
cc_187 N_A_27_368#_c_185_n N_Y_c_341_n 0.012724f $X=1.915 $Y=1.805 $X2=0 $Y2=0
cc_188 N_Y_c_313_n N_VGND_M1003_d 0.0103921f $X=2.36 $Y=0.925 $X2=0 $Y2=0
cc_189 N_Y_c_306_n N_VGND_c_364_n 0.0267724f $X=1.355 $Y=0.675 $X2=0 $Y2=0
cc_190 N_Y_c_313_n N_VGND_c_365_n 0.0189346f $X=2.36 $Y=0.925 $X2=0 $Y2=0
cc_191 N_Y_c_307_n N_VGND_c_365_n 0.0127976f $X=2.525 $Y=0.515 $X2=0 $Y2=0
cc_192 N_Y_c_308_n N_VGND_c_365_n 0.0137088f $X=1.69 $Y=0.675 $X2=0 $Y2=0
cc_193 N_Y_c_306_n N_VGND_c_366_n 0.0485195f $X=1.355 $Y=0.675 $X2=0 $Y2=0
cc_194 N_Y_c_307_n N_VGND_c_368_n 0.014552f $X=2.525 $Y=0.515 $X2=0 $Y2=0
cc_195 N_Y_c_307_n N_VGND_c_369_n 0.0193213f $X=2.525 $Y=0.515 $X2=0 $Y2=0
cc_196 N_Y_c_306_n N_VGND_c_370_n 0.0389588f $X=1.355 $Y=0.675 $X2=0 $Y2=0
cc_197 N_Y_c_313_n N_VGND_c_370_n 0.0108653f $X=2.36 $Y=0.925 $X2=0 $Y2=0
cc_198 N_Y_c_307_n N_VGND_c_370_n 0.0119791f $X=2.525 $Y=0.515 $X2=0 $Y2=0
