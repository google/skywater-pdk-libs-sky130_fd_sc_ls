* File: sky130_fd_sc_ls__a32oi_2.pxi.spice
* Created: Fri Aug 28 13:00:45 2020
* 
x_PM_SKY130_FD_SC_LS__A32OI_2%B2 N_B2_M1010_g N_B2_c_104_n N_B2_M1007_g
+ N_B2_M1016_g N_B2_c_105_n N_B2_M1009_g N_B2_c_101_n B2 N_B2_c_102_n
+ N_B2_c_103_n PM_SKY130_FD_SC_LS__A32OI_2%B2
x_PM_SKY130_FD_SC_LS__A32OI_2%B1 N_B1_c_147_n N_B1_M1003_g N_B1_c_151_n
+ N_B1_M1015_g N_B1_c_148_n N_B1_M1008_g N_B1_c_152_n N_B1_M1019_g B1 B1
+ N_B1_c_150_n PM_SKY130_FD_SC_LS__A32OI_2%B1
x_PM_SKY130_FD_SC_LS__A32OI_2%A1 N_A1_c_207_n N_A1_M1004_g N_A1_c_203_n
+ N_A1_M1005_g N_A1_c_204_n N_A1_M1018_g N_A1_c_208_n N_A1_M1017_g A1
+ N_A1_c_206_n PM_SKY130_FD_SC_LS__A32OI_2%A1
x_PM_SKY130_FD_SC_LS__A32OI_2%A2 N_A2_M1013_g N_A2_c_264_n N_A2_M1000_g
+ N_A2_c_265_n N_A2_M1001_g N_A2_M1014_g N_A2_c_260_n N_A2_c_261_n N_A2_c_262_n
+ A2 A2 N_A2_c_263_n PM_SKY130_FD_SC_LS__A32OI_2%A2
x_PM_SKY130_FD_SC_LS__A32OI_2%A3 N_A3_c_320_n N_A3_M1011_g N_A3_c_316_n
+ N_A3_M1002_g N_A3_c_321_n N_A3_M1012_g N_A3_c_317_n N_A3_M1006_g A3
+ N_A3_c_319_n PM_SKY130_FD_SC_LS__A32OI_2%A3
x_PM_SKY130_FD_SC_LS__A32OI_2%A_27_368# N_A_27_368#_M1007_s N_A_27_368#_M1009_s
+ N_A_27_368#_M1019_s N_A_27_368#_M1017_s N_A_27_368#_M1001_d
+ N_A_27_368#_M1012_s N_A_27_368#_c_357_n N_A_27_368#_c_358_n
+ N_A_27_368#_c_359_n N_A_27_368#_c_374_n N_A_27_368#_c_360_n
+ N_A_27_368#_c_413_p N_A_27_368#_c_380_n N_A_27_368#_c_361_n
+ N_A_27_368#_c_385_n N_A_27_368#_c_362_n N_A_27_368#_c_363_n
+ N_A_27_368#_c_364_n N_A_27_368#_c_365_n N_A_27_368#_c_366_n
+ N_A_27_368#_c_383_n PM_SKY130_FD_SC_LS__A32OI_2%A_27_368#
x_PM_SKY130_FD_SC_LS__A32OI_2%Y N_Y_M1003_d N_Y_M1005_d N_Y_M1007_d N_Y_M1015_d
+ N_Y_c_447_n N_Y_c_457_n N_Y_c_448_n N_Y_c_465_n N_Y_c_444_n N_Y_c_449_n
+ N_Y_c_520_p N_Y_c_472_n N_Y_c_450_n N_Y_c_487_n N_Y_c_445_n Y N_Y_c_452_n Y
+ PM_SKY130_FD_SC_LS__A32OI_2%Y
x_PM_SKY130_FD_SC_LS__A32OI_2%VPWR N_VPWR_M1004_d N_VPWR_M1000_s N_VPWR_M1011_d
+ N_VPWR_c_525_n N_VPWR_c_526_n N_VPWR_c_527_n N_VPWR_c_528_n N_VPWR_c_529_n
+ VPWR N_VPWR_c_530_n N_VPWR_c_531_n N_VPWR_c_532_n N_VPWR_c_524_n
+ N_VPWR_c_534_n N_VPWR_c_535_n PM_SKY130_FD_SC_LS__A32OI_2%VPWR
x_PM_SKY130_FD_SC_LS__A32OI_2%A_27_74# N_A_27_74#_M1010_d N_A_27_74#_M1016_d
+ N_A_27_74#_M1008_s N_A_27_74#_c_593_n N_A_27_74#_c_594_n N_A_27_74#_c_595_n
+ N_A_27_74#_c_596_n N_A_27_74#_c_597_n N_A_27_74#_c_598_n
+ PM_SKY130_FD_SC_LS__A32OI_2%A_27_74#
x_PM_SKY130_FD_SC_LS__A32OI_2%VGND N_VGND_M1010_s N_VGND_M1002_s N_VGND_M1006_s
+ N_VGND_c_630_n N_VGND_c_631_n N_VGND_c_632_n N_VGND_c_633_n VGND
+ N_VGND_c_634_n N_VGND_c_635_n N_VGND_c_636_n N_VGND_c_637_n N_VGND_c_638_n
+ N_VGND_c_639_n PM_SKY130_FD_SC_LS__A32OI_2%VGND
x_PM_SKY130_FD_SC_LS__A32OI_2%A_507_74# N_A_507_74#_M1005_s N_A_507_74#_M1018_s
+ N_A_507_74#_M1014_d N_A_507_74#_c_697_n N_A_507_74#_c_698_n
+ N_A_507_74#_c_699_n N_A_507_74#_c_700_n N_A_507_74#_c_701_n
+ N_A_507_74#_c_702_n PM_SKY130_FD_SC_LS__A32OI_2%A_507_74#
x_PM_SKY130_FD_SC_LS__A32OI_2%A_771_74# N_A_771_74#_M1013_s N_A_771_74#_M1002_d
+ N_A_771_74#_c_764_n N_A_771_74#_c_741_n N_A_771_74#_c_742_n
+ N_A_771_74#_c_743_n PM_SKY130_FD_SC_LS__A32OI_2%A_771_74#
cc_1 VNB N_B2_M1010_g 0.0296069f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_B2_M1016_g 0.0221212f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=0.74
cc_3 VNB N_B2_c_101_n 0.00135493f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.465
cc_4 VNB N_B2_c_102_n 0.0565743f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.532
cc_5 VNB N_B2_c_103_n 0.0184277f $X=-0.19 $Y=-0.245 $X2=0.355 $Y2=1.54
cc_6 VNB N_B1_c_147_n 0.0164156f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.3
cc_7 VNB N_B1_c_148_n 0.0207512f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.4
cc_8 VNB B1 0.00940302f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.4
cc_9 VNB N_B1_c_150_n 0.0701358f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_10 VNB N_A1_c_203_n 0.0205288f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A1_c_204_n 0.0164898f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.4
cc_12 VNB A1 0.00441958f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.4
cc_13 VNB N_A1_c_206_n 0.0910124f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_14 VNB N_A2_M1013_g 0.0249505f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_15 VNB N_A2_M1014_g 0.0289552f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.4
cc_16 VNB N_A2_c_260_n 0.00990425f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.465
cc_17 VNB N_A2_c_261_n 0.0161486f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.465
cc_18 VNB N_A2_c_262_n 0.0139879f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.465
cc_19 VNB N_A2_c_263_n 0.00476662f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.532
cc_20 VNB N_A3_c_316_n 0.0192891f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A3_c_317_n 0.0209684f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=0.74
cc_22 VNB A3 0.0140818f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.4
cc_23 VNB N_A3_c_319_n 0.128157f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.465
cc_24 VNB N_Y_c_444_n 0.0117593f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.532
cc_25 VNB N_Y_c_445_n 0.00184708f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB Y 0.00206864f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VPWR_c_524_n 0.263193f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_27_74#_c_593_n 0.0247745f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.765
cc_29 VNB N_A_27_74#_c_594_n 0.00666543f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.4
cc_30 VNB N_A_27_74#_c_595_n 0.00978809f $X=-0.19 $Y=-0.245 $X2=0.355 $Y2=1.465
cc_31 VNB N_A_27_74#_c_596_n 0.00302115f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_32 VNB N_A_27_74#_c_597_n 0.00217191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_27_74#_c_598_n 0.00716337f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.532
cc_34 VNB N_VGND_c_630_n 0.00615265f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.765
cc_35 VNB N_VGND_c_631_n 0.0123645f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.465
cc_36 VNB N_VGND_c_632_n 0.0120272f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.465
cc_37 VNB N_VGND_c_633_n 0.0341338f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_38 VNB N_VGND_c_634_n 0.0173909f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.532
cc_39 VNB N_VGND_c_635_n 0.0965919f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_636_n 0.0172524f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_637_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_638_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_639_n 0.353339f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_507_74#_c_697_n 0.00199363f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=0.74
cc_45 VNB N_A_507_74#_c_698_n 0.00487422f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.4
cc_46 VNB N_A_507_74#_c_699_n 0.00713963f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.465
cc_47 VNB N_A_507_74#_c_700_n 0.00384069f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_48 VNB N_A_507_74#_c_701_n 0.00655402f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.532
cc_49 VNB N_A_507_74#_c_702_n 0.0022203f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.54
cc_50 VNB N_A_771_74#_c_741_n 0.0275552f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_771_74#_c_742_n 0.00341417f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.765
cc_52 VNB N_A_771_74#_c_743_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0.355 $Y2=1.465
cc_53 VPB N_B2_c_104_n 0.0189373f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.765
cc_54 VPB N_B2_c_105_n 0.0151714f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.765
cc_55 VPB N_B2_c_102_n 0.0143874f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.532
cc_56 VPB N_B2_c_103_n 0.0080267f $X=-0.19 $Y=1.66 $X2=0.355 $Y2=1.54
cc_57 VPB N_B1_c_151_n 0.0151927f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_B1_c_152_n 0.0148847f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=0.74
cc_59 VPB N_B1_c_150_n 0.0135068f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_60 VPB N_A1_c_207_n 0.0169296f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.3
cc_61 VPB N_A1_c_208_n 0.01744f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=0.74
cc_62 VPB N_A1_c_206_n 0.0152479f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_63 VPB N_A2_c_264_n 0.0162649f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.765
cc_64 VPB N_A2_c_265_n 0.0169833f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.3
cc_65 VPB N_A2_c_260_n 0.00553092f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.465
cc_66 VPB N_A2_c_261_n 0.010221f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.465
cc_67 VPB N_A2_c_262_n 0.00675179f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.465
cc_68 VPB N_A2_c_263_n 0.00655669f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.532
cc_69 VPB N_A3_c_320_n 0.0169802f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.3
cc_70 VPB N_A3_c_321_n 0.0201263f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=2.4
cc_71 VPB N_A3_c_319_n 0.0162511f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.465
cc_72 VPB N_A_27_368#_c_357_n 0.0366851f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_A_27_368#_c_358_n 0.00269852f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.532
cc_74 VPB N_A_27_368#_c_359_n 0.00988933f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.532
cc_75 VPB N_A_27_368#_c_360_n 0.00603766f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_A_27_368#_c_361_n 0.00247739f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_A_27_368#_c_362_n 0.00616464f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_A_27_368#_c_363_n 0.00406258f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 VPB N_A_27_368#_c_364_n 0.0147997f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 VPB N_A_27_368#_c_365_n 0.0441294f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_A_27_368#_c_366_n 0.0022931f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 VPB N_Y_c_447_n 0.00249201f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.4
cc_83 VPB N_Y_c_448_n 0.00647299f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.465
cc_84 VPB N_Y_c_449_n 0.0107069f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.54
cc_85 VPB N_Y_c_450_n 0.00321873f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB Y 0.00110955f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_Y_c_452_n 0.00194891f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_525_n 0.00684019f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.765
cc_89 VPB N_VPWR_c_526_n 0.00589302f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.465
cc_90 VPB N_VPWR_c_527_n 0.00970163f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_91 VPB N_VPWR_c_528_n 0.021538f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.532
cc_92 VPB N_VPWR_c_529_n 0.00632158f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.532
cc_93 VPB N_VPWR_c_530_n 0.0616751f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_531_n 0.0174563f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_532_n 0.027107f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_524_n 0.0842887f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_534_n 0.0132794f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_535_n 0.00642979f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 N_B2_M1016_g N_B1_c_147_n 0.0167802f $X=0.975 $Y=0.74 $X2=-0.19 $Y2=-0.245
cc_100 N_B2_c_105_n N_B1_c_151_n 0.0289268f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_101 N_B2_M1016_g B1 3.50863e-19 $X=0.975 $Y=0.74 $X2=0 $Y2=0
cc_102 N_B2_c_101_n B1 0.0101592f $X=0.925 $Y=1.465 $X2=0 $Y2=0
cc_103 N_B2_c_102_n B1 9.46057e-19 $X=0.975 $Y=1.532 $X2=0 $Y2=0
cc_104 N_B2_c_101_n N_B1_c_150_n 0.00166525f $X=0.925 $Y=1.465 $X2=0 $Y2=0
cc_105 N_B2_c_102_n N_B1_c_150_n 0.0214874f $X=0.975 $Y=1.532 $X2=0 $Y2=0
cc_106 N_B2_c_104_n N_A_27_368#_c_357_n 0.0105585f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_107 N_B2_c_105_n N_A_27_368#_c_357_n 2.79308e-19 $X=1.005 $Y=1.765 $X2=0
+ $Y2=0
cc_108 N_B2_c_101_n N_A_27_368#_c_357_n 0.00311722f $X=0.925 $Y=1.465 $X2=0
+ $Y2=0
cc_109 N_B2_c_103_n N_A_27_368#_c_357_n 0.0205168f $X=0.355 $Y=1.54 $X2=0 $Y2=0
cc_110 N_B2_c_104_n N_A_27_368#_c_358_n 0.0114142f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_111 N_B2_c_105_n N_A_27_368#_c_358_n 0.0140406f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_112 N_B2_c_104_n N_A_27_368#_c_359_n 0.00253309f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_113 N_B2_c_104_n N_Y_c_447_n 0.0013124f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_114 N_B2_c_105_n N_Y_c_447_n 9.16146e-19 $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_115 N_B2_c_101_n N_Y_c_447_n 0.0277622f $X=0.925 $Y=1.465 $X2=0 $Y2=0
cc_116 N_B2_c_102_n N_Y_c_447_n 0.00806131f $X=0.975 $Y=1.532 $X2=0 $Y2=0
cc_117 N_B2_c_105_n N_Y_c_457_n 0.00911772f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_118 N_B2_c_105_n N_Y_c_448_n 0.01222f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_119 N_B2_c_101_n N_Y_c_448_n 0.0103583f $X=0.925 $Y=1.465 $X2=0 $Y2=0
cc_120 N_B2_c_102_n N_Y_c_448_n 4.55036e-19 $X=0.975 $Y=1.532 $X2=0 $Y2=0
cc_121 N_B2_c_104_n N_VPWR_c_530_n 0.00278262f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_122 N_B2_c_105_n N_VPWR_c_530_n 0.00278271f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_123 N_B2_c_104_n N_VPWR_c_524_n 0.0035775f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_124 N_B2_c_105_n N_VPWR_c_524_n 0.00354754f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_125 N_B2_M1010_g N_A_27_74#_c_593_n 0.00159319f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_126 N_B2_M1010_g N_A_27_74#_c_594_n 0.0128698f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_127 N_B2_M1016_g N_A_27_74#_c_594_n 0.0134606f $X=0.975 $Y=0.74 $X2=0 $Y2=0
cc_128 N_B2_c_101_n N_A_27_74#_c_594_n 0.0535577f $X=0.925 $Y=1.465 $X2=0 $Y2=0
cc_129 N_B2_c_102_n N_A_27_74#_c_594_n 0.00453952f $X=0.975 $Y=1.532 $X2=0 $Y2=0
cc_130 N_B2_c_103_n N_A_27_74#_c_595_n 0.0217492f $X=0.355 $Y=1.54 $X2=0 $Y2=0
cc_131 N_B2_M1016_g N_A_27_74#_c_597_n 0.00106427f $X=0.975 $Y=0.74 $X2=0 $Y2=0
cc_132 N_B2_M1010_g N_VGND_c_630_n 0.0125039f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_133 N_B2_M1016_g N_VGND_c_630_n 0.00182553f $X=0.975 $Y=0.74 $X2=0 $Y2=0
cc_134 N_B2_M1010_g N_VGND_c_634_n 0.00383152f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_135 N_B2_M1016_g N_VGND_c_635_n 0.00461464f $X=0.975 $Y=0.74 $X2=0 $Y2=0
cc_136 N_B2_M1010_g N_VGND_c_639_n 0.00761198f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_137 N_B2_M1016_g N_VGND_c_639_n 0.00908237f $X=0.975 $Y=0.74 $X2=0 $Y2=0
cc_138 N_B1_c_152_n N_A1_c_207_n 0.0240853f $X=2.005 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_139 B1 A1 0.0311944f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_140 N_B1_c_150_n A1 3.24246e-19 $X=2.005 $Y=1.492 $X2=0 $Y2=0
cc_141 B1 N_A1_c_206_n 0.00251916f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_142 N_B1_c_150_n N_A1_c_206_n 0.0280077f $X=2.005 $Y=1.492 $X2=0 $Y2=0
cc_143 N_B1_c_151_n N_A_27_368#_c_374_n 0.0110199f $X=1.505 $Y=1.765 $X2=0 $Y2=0
cc_144 N_B1_c_152_n N_A_27_368#_c_374_n 2.69714e-19 $X=2.005 $Y=1.765 $X2=0
+ $Y2=0
cc_145 N_B1_c_151_n N_A_27_368#_c_360_n 0.0111147f $X=1.505 $Y=1.765 $X2=0 $Y2=0
cc_146 N_B1_c_152_n N_A_27_368#_c_360_n 0.0137852f $X=2.005 $Y=1.765 $X2=0 $Y2=0
cc_147 N_B1_c_151_n N_A_27_368#_c_366_n 0.00189622f $X=1.505 $Y=1.765 $X2=0
+ $Y2=0
cc_148 N_B1_c_151_n N_Y_c_457_n 5.80433e-19 $X=1.505 $Y=1.765 $X2=0 $Y2=0
cc_149 N_B1_c_151_n N_Y_c_448_n 0.0178968f $X=1.505 $Y=1.765 $X2=0 $Y2=0
cc_150 B1 N_Y_c_448_n 0.00593209f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_151 N_B1_c_150_n N_Y_c_448_n 0.00385849f $X=2.005 $Y=1.492 $X2=0 $Y2=0
cc_152 N_B1_c_152_n N_Y_c_465_n 0.00825076f $X=2.005 $Y=1.765 $X2=0 $Y2=0
cc_153 N_B1_c_148_n N_Y_c_444_n 0.0114763f $X=1.835 $Y=1.22 $X2=0 $Y2=0
cc_154 B1 N_Y_c_444_n 0.03567f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_155 N_B1_c_150_n N_Y_c_444_n 0.00154347f $X=2.005 $Y=1.492 $X2=0 $Y2=0
cc_156 N_B1_c_152_n N_Y_c_449_n 0.00919138f $X=2.005 $Y=1.765 $X2=0 $Y2=0
cc_157 B1 N_Y_c_449_n 0.0248442f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_158 N_B1_c_150_n N_Y_c_449_n 0.00527636f $X=2.005 $Y=1.492 $X2=0 $Y2=0
cc_159 N_B1_c_147_n N_Y_c_472_n 0.00608134f $X=1.405 $Y=1.22 $X2=0 $Y2=0
cc_160 N_B1_c_148_n N_Y_c_472_n 0.0100827f $X=1.835 $Y=1.22 $X2=0 $Y2=0
cc_161 B1 N_Y_c_472_n 0.01963f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_162 N_B1_c_150_n N_Y_c_472_n 6.70474e-19 $X=2.005 $Y=1.492 $X2=0 $Y2=0
cc_163 N_B1_c_151_n N_Y_c_450_n 0.00116261f $X=1.505 $Y=1.765 $X2=0 $Y2=0
cc_164 N_B1_c_152_n N_Y_c_450_n 0.00275532f $X=2.005 $Y=1.765 $X2=0 $Y2=0
cc_165 B1 N_Y_c_450_n 0.0279177f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_166 N_B1_c_150_n N_Y_c_450_n 0.00678054f $X=2.005 $Y=1.492 $X2=0 $Y2=0
cc_167 N_B1_c_152_n N_VPWR_c_525_n 3.11624e-19 $X=2.005 $Y=1.765 $X2=0 $Y2=0
cc_168 N_B1_c_151_n N_VPWR_c_530_n 0.00278257f $X=1.505 $Y=1.765 $X2=0 $Y2=0
cc_169 N_B1_c_152_n N_VPWR_c_530_n 0.00278271f $X=2.005 $Y=1.765 $X2=0 $Y2=0
cc_170 N_B1_c_151_n N_VPWR_c_524_n 0.00354797f $X=1.505 $Y=1.765 $X2=0 $Y2=0
cc_171 N_B1_c_152_n N_VPWR_c_524_n 0.00354798f $X=2.005 $Y=1.765 $X2=0 $Y2=0
cc_172 N_B1_c_147_n N_A_27_74#_c_594_n 6.05444e-19 $X=1.405 $Y=1.22 $X2=0 $Y2=0
cc_173 N_B1_c_147_n N_A_27_74#_c_596_n 0.0119575f $X=1.405 $Y=1.22 $X2=0 $Y2=0
cc_174 N_B1_c_148_n N_A_27_74#_c_596_n 0.0107047f $X=1.835 $Y=1.22 $X2=0 $Y2=0
cc_175 N_B1_c_148_n N_A_27_74#_c_598_n 0.00165289f $X=1.835 $Y=1.22 $X2=0 $Y2=0
cc_176 N_B1_c_147_n N_VGND_c_635_n 0.00278271f $X=1.405 $Y=1.22 $X2=0 $Y2=0
cc_177 N_B1_c_148_n N_VGND_c_635_n 0.00278271f $X=1.835 $Y=1.22 $X2=0 $Y2=0
cc_178 N_B1_c_147_n N_VGND_c_639_n 0.00353526f $X=1.405 $Y=1.22 $X2=0 $Y2=0
cc_179 N_B1_c_148_n N_VGND_c_639_n 0.00357518f $X=1.835 $Y=1.22 $X2=0 $Y2=0
cc_180 N_A1_c_204_n N_A2_M1013_g 0.0117174f $X=3.325 $Y=1.22 $X2=0 $Y2=0
cc_181 N_A1_c_206_n N_A2_M1013_g 0.0257905f $X=3.325 $Y=1.492 $X2=0 $Y2=0
cc_182 N_A1_c_208_n N_A2_c_264_n 0.0116278f $X=3.345 $Y=1.765 $X2=0 $Y2=0
cc_183 N_A1_c_206_n N_A2_c_263_n 0.00438872f $X=3.325 $Y=1.492 $X2=0 $Y2=0
cc_184 N_A1_c_207_n N_A_27_368#_c_360_n 0.00108375f $X=2.505 $Y=1.765 $X2=0
+ $Y2=0
cc_185 N_A1_c_207_n N_A_27_368#_c_380_n 0.0142499f $X=2.505 $Y=1.765 $X2=0 $Y2=0
cc_186 N_A1_c_208_n N_A_27_368#_c_380_n 0.0178396f $X=3.345 $Y=1.765 $X2=0 $Y2=0
cc_187 N_A1_c_206_n N_A_27_368#_c_380_n 8.27888e-19 $X=3.325 $Y=1.492 $X2=0
+ $Y2=0
cc_188 N_A1_c_208_n N_A_27_368#_c_383_n 0.0066764f $X=3.345 $Y=1.765 $X2=0 $Y2=0
cc_189 N_A1_c_203_n N_Y_c_444_n 0.0162888f $X=2.895 $Y=1.22 $X2=0 $Y2=0
cc_190 A1 N_Y_c_444_n 0.0256443f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_191 N_A1_c_206_n N_Y_c_444_n 0.00323723f $X=3.325 $Y=1.492 $X2=0 $Y2=0
cc_192 N_A1_c_207_n N_Y_c_449_n 0.00800218f $X=2.505 $Y=1.765 $X2=0 $Y2=0
cc_193 A1 N_Y_c_449_n 0.0244344f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_194 N_A1_c_206_n N_Y_c_449_n 0.0160464f $X=3.325 $Y=1.492 $X2=0 $Y2=0
cc_195 N_A1_c_207_n N_Y_c_450_n 3.22368e-19 $X=2.505 $Y=1.765 $X2=0 $Y2=0
cc_196 N_A1_c_206_n N_Y_c_487_n 0.0077643f $X=3.325 $Y=1.492 $X2=0 $Y2=0
cc_197 N_A1_c_203_n N_Y_c_445_n 0.00251469f $X=2.895 $Y=1.22 $X2=0 $Y2=0
cc_198 N_A1_c_204_n N_Y_c_445_n 0.00224552f $X=3.325 $Y=1.22 $X2=0 $Y2=0
cc_199 A1 N_Y_c_445_n 0.0214567f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_200 N_A1_c_206_n N_Y_c_445_n 0.00306807f $X=3.325 $Y=1.492 $X2=0 $Y2=0
cc_201 N_A1_c_206_n Y 0.0187089f $X=3.325 $Y=1.492 $X2=0 $Y2=0
cc_202 N_A1_c_208_n N_Y_c_452_n 0.0028927f $X=3.345 $Y=1.765 $X2=0 $Y2=0
cc_203 N_A1_c_206_n N_Y_c_452_n 6.9066e-19 $X=3.325 $Y=1.492 $X2=0 $Y2=0
cc_204 N_A1_c_207_n N_VPWR_c_525_n 0.00950907f $X=2.505 $Y=1.765 $X2=0 $Y2=0
cc_205 N_A1_c_208_n N_VPWR_c_525_n 0.0102691f $X=3.345 $Y=1.765 $X2=0 $Y2=0
cc_206 N_A1_c_207_n N_VPWR_c_530_n 0.00429299f $X=2.505 $Y=1.765 $X2=0 $Y2=0
cc_207 N_A1_c_208_n N_VPWR_c_531_n 0.00429299f $X=3.345 $Y=1.765 $X2=0 $Y2=0
cc_208 N_A1_c_207_n N_VPWR_c_524_n 0.00848235f $X=2.505 $Y=1.765 $X2=0 $Y2=0
cc_209 N_A1_c_208_n N_VPWR_c_524_n 0.00847805f $X=3.345 $Y=1.765 $X2=0 $Y2=0
cc_210 N_A1_c_203_n N_A_27_74#_c_598_n 9.7204e-19 $X=2.895 $Y=1.22 $X2=0 $Y2=0
cc_211 N_A1_c_203_n N_VGND_c_635_n 0.00279469f $X=2.895 $Y=1.22 $X2=0 $Y2=0
cc_212 N_A1_c_204_n N_VGND_c_635_n 0.00278247f $X=3.325 $Y=1.22 $X2=0 $Y2=0
cc_213 N_A1_c_203_n N_VGND_c_639_n 0.00357517f $X=2.895 $Y=1.22 $X2=0 $Y2=0
cc_214 N_A1_c_204_n N_VGND_c_639_n 0.00353752f $X=3.325 $Y=1.22 $X2=0 $Y2=0
cc_215 N_A1_c_203_n N_A_507_74#_c_697_n 0.0079299f $X=2.895 $Y=1.22 $X2=0 $Y2=0
cc_216 N_A1_c_204_n N_A_507_74#_c_697_n 0.0100711f $X=3.325 $Y=1.22 $X2=0 $Y2=0
cc_217 N_A1_c_203_n N_A_507_74#_c_698_n 6.12241e-19 $X=2.895 $Y=1.22 $X2=0 $Y2=0
cc_218 N_A1_c_204_n N_A_507_74#_c_698_n 0.010463f $X=3.325 $Y=1.22 $X2=0 $Y2=0
cc_219 N_A1_c_206_n N_A_507_74#_c_698_n 0.0018231f $X=3.325 $Y=1.492 $X2=0 $Y2=0
cc_220 N_A1_c_203_n N_A_507_74#_c_701_n 0.00735466f $X=2.895 $Y=1.22 $X2=0 $Y2=0
cc_221 N_A1_c_204_n N_A_507_74#_c_701_n 5.3819e-19 $X=3.325 $Y=1.22 $X2=0 $Y2=0
cc_222 N_A1_c_204_n N_A_507_74#_c_702_n 0.00194567f $X=3.325 $Y=1.22 $X2=0 $Y2=0
cc_223 N_A2_c_265_n N_A3_c_320_n 0.0216067f $X=4.31 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_224 N_A2_M1014_g N_A3_c_319_n 0.018186f $X=4.325 $Y=0.74 $X2=0 $Y2=0
cc_225 N_A2_c_263_n N_A3_c_319_n 0.00225986f $X=4.21 $Y=1.515 $X2=0 $Y2=0
cc_226 N_A2_c_264_n N_A_27_368#_c_361_n 0.00801929f $X=3.795 $Y=1.765 $X2=0
+ $Y2=0
cc_227 N_A2_c_264_n N_A_27_368#_c_385_n 0.0129284f $X=3.795 $Y=1.765 $X2=0 $Y2=0
cc_228 N_A2_c_265_n N_A_27_368#_c_385_n 0.0162783f $X=4.31 $Y=1.765 $X2=0 $Y2=0
cc_229 N_A2_c_261_n N_A_27_368#_c_385_n 0.00165941f $X=4.22 $Y=1.515 $X2=0 $Y2=0
cc_230 N_A2_c_263_n N_A_27_368#_c_385_n 0.0449973f $X=4.21 $Y=1.515 $X2=0 $Y2=0
cc_231 N_A2_c_265_n N_A_27_368#_c_362_n 0.00497557f $X=4.31 $Y=1.765 $X2=0 $Y2=0
cc_232 N_A2_c_262_n N_A_27_368#_c_362_n 3.89364e-19 $X=4.31 $Y=1.557 $X2=0 $Y2=0
cc_233 N_A2_c_263_n N_A_27_368#_c_362_n 0.00521764f $X=4.21 $Y=1.515 $X2=0 $Y2=0
cc_234 N_A2_c_265_n N_A_27_368#_c_363_n 0.00595854f $X=4.31 $Y=1.765 $X2=0 $Y2=0
cc_235 N_A2_c_264_n N_A_27_368#_c_383_n 0.00299506f $X=3.795 $Y=1.765 $X2=0
+ $Y2=0
cc_236 N_A2_c_265_n N_A_27_368#_c_383_n 6.0668e-19 $X=4.31 $Y=1.765 $X2=0 $Y2=0
cc_237 N_A2_c_263_n N_A_27_368#_c_383_n 0.0193124f $X=4.21 $Y=1.515 $X2=0 $Y2=0
cc_238 N_A2_M1013_g N_Y_c_487_n 4.94418e-19 $X=3.78 $Y=0.74 $X2=0 $Y2=0
cc_239 N_A2_c_263_n Y 0.0234231f $X=4.21 $Y=1.515 $X2=0 $Y2=0
cc_240 N_A2_c_263_n N_Y_c_452_n 0.00420642f $X=4.21 $Y=1.515 $X2=0 $Y2=0
cc_241 N_A2_c_264_n N_VPWR_c_525_n 4.84605e-19 $X=3.795 $Y=1.765 $X2=0 $Y2=0
cc_242 N_A2_c_264_n N_VPWR_c_526_n 0.00558936f $X=3.795 $Y=1.765 $X2=0 $Y2=0
cc_243 N_A2_c_265_n N_VPWR_c_526_n 0.0117108f $X=4.31 $Y=1.765 $X2=0 $Y2=0
cc_244 N_A2_c_265_n N_VPWR_c_528_n 0.00413917f $X=4.31 $Y=1.765 $X2=0 $Y2=0
cc_245 N_A2_c_264_n N_VPWR_c_531_n 0.00445602f $X=3.795 $Y=1.765 $X2=0 $Y2=0
cc_246 N_A2_c_264_n N_VPWR_c_524_n 0.00857592f $X=3.795 $Y=1.765 $X2=0 $Y2=0
cc_247 N_A2_c_265_n N_VPWR_c_524_n 0.0081916f $X=4.31 $Y=1.765 $X2=0 $Y2=0
cc_248 N_A2_M1014_g N_VGND_c_631_n 0.00177115f $X=4.325 $Y=0.74 $X2=0 $Y2=0
cc_249 N_A2_M1013_g N_VGND_c_635_n 0.00278271f $X=3.78 $Y=0.74 $X2=0 $Y2=0
cc_250 N_A2_M1014_g N_VGND_c_635_n 0.00278247f $X=4.325 $Y=0.74 $X2=0 $Y2=0
cc_251 N_A2_M1013_g N_VGND_c_639_n 0.00354791f $X=3.78 $Y=0.74 $X2=0 $Y2=0
cc_252 N_A2_M1014_g N_VGND_c_639_n 0.00359462f $X=4.325 $Y=0.74 $X2=0 $Y2=0
cc_253 N_A2_M1013_g N_A_507_74#_c_698_n 4.70861e-19 $X=3.78 $Y=0.74 $X2=0 $Y2=0
cc_254 N_A2_c_263_n N_A_507_74#_c_698_n 0.0164713f $X=4.21 $Y=1.515 $X2=0 $Y2=0
cc_255 N_A2_M1013_g N_A_507_74#_c_699_n 0.0123067f $X=3.78 $Y=0.74 $X2=0 $Y2=0
cc_256 N_A2_M1014_g N_A_507_74#_c_699_n 0.0124893f $X=4.325 $Y=0.74 $X2=0 $Y2=0
cc_257 N_A2_M1013_g N_A_507_74#_c_700_n 5.11757e-19 $X=3.78 $Y=0.74 $X2=0 $Y2=0
cc_258 N_A2_M1014_g N_A_507_74#_c_700_n 0.00736432f $X=4.325 $Y=0.74 $X2=0 $Y2=0
cc_259 N_A2_M1013_g N_A_507_74#_c_702_n 0.00142735f $X=3.78 $Y=0.74 $X2=0 $Y2=0
cc_260 N_A2_M1014_g N_A_771_74#_c_741_n 0.015237f $X=4.325 $Y=0.74 $X2=0 $Y2=0
cc_261 N_A2_c_263_n N_A_771_74#_c_741_n 0.0124962f $X=4.21 $Y=1.515 $X2=0 $Y2=0
cc_262 N_A2_M1013_g N_A_771_74#_c_742_n 0.00177175f $X=3.78 $Y=0.74 $X2=0 $Y2=0
cc_263 N_A2_c_261_n N_A_771_74#_c_742_n 0.00497826f $X=4.22 $Y=1.515 $X2=0 $Y2=0
cc_264 N_A2_c_263_n N_A_771_74#_c_742_n 0.0279649f $X=4.21 $Y=1.515 $X2=0 $Y2=0
cc_265 N_A3_c_320_n N_A_27_368#_c_362_n 0.0051368f $X=4.935 $Y=1.765 $X2=0 $Y2=0
cc_266 N_A3_c_321_n N_A_27_368#_c_362_n 5.34941e-19 $X=5.485 $Y=1.765 $X2=0
+ $Y2=0
cc_267 N_A3_c_319_n N_A_27_368#_c_362_n 0.00181952f $X=5.745 $Y=1.492 $X2=0
+ $Y2=0
cc_268 N_A3_c_320_n N_A_27_368#_c_363_n 0.0212604f $X=4.935 $Y=1.765 $X2=0 $Y2=0
cc_269 N_A3_c_320_n N_A_27_368#_c_364_n 0.00941072f $X=4.935 $Y=1.765 $X2=0
+ $Y2=0
cc_270 N_A3_c_321_n N_A_27_368#_c_364_n 0.011067f $X=5.485 $Y=1.765 $X2=0 $Y2=0
cc_271 A3 N_A_27_368#_c_364_n 0.00760155f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_272 N_A3_c_319_n N_A_27_368#_c_364_n 0.0278435f $X=5.745 $Y=1.492 $X2=0 $Y2=0
cc_273 N_A3_c_320_n N_A_27_368#_c_365_n 7.10227e-19 $X=4.935 $Y=1.765 $X2=0
+ $Y2=0
cc_274 N_A3_c_321_n N_A_27_368#_c_365_n 0.0136873f $X=5.485 $Y=1.765 $X2=0 $Y2=0
cc_275 N_A3_c_320_n N_VPWR_c_526_n 9.11544e-19 $X=4.935 $Y=1.765 $X2=0 $Y2=0
cc_276 N_A3_c_320_n N_VPWR_c_527_n 0.00874363f $X=4.935 $Y=1.765 $X2=0 $Y2=0
cc_277 N_A3_c_321_n N_VPWR_c_527_n 0.00874363f $X=5.485 $Y=1.765 $X2=0 $Y2=0
cc_278 N_A3_c_320_n N_VPWR_c_528_n 0.00445602f $X=4.935 $Y=1.765 $X2=0 $Y2=0
cc_279 N_A3_c_321_n N_VPWR_c_532_n 0.00445602f $X=5.485 $Y=1.765 $X2=0 $Y2=0
cc_280 N_A3_c_320_n N_VPWR_c_524_n 0.00859231f $X=4.935 $Y=1.765 $X2=0 $Y2=0
cc_281 N_A3_c_321_n N_VPWR_c_524_n 0.00861874f $X=5.485 $Y=1.765 $X2=0 $Y2=0
cc_282 N_A3_c_316_n N_VGND_c_631_n 0.00562548f $X=5.315 $Y=1.22 $X2=0 $Y2=0
cc_283 N_A3_c_316_n N_VGND_c_633_n 5.69925e-19 $X=5.315 $Y=1.22 $X2=0 $Y2=0
cc_284 N_A3_c_317_n N_VGND_c_633_n 0.0122959f $X=5.745 $Y=1.22 $X2=0 $Y2=0
cc_285 A3 N_VGND_c_633_n 0.0251682f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_286 N_A3_c_319_n N_VGND_c_633_n 0.00192797f $X=5.745 $Y=1.492 $X2=0 $Y2=0
cc_287 N_A3_c_316_n N_VGND_c_636_n 0.00434272f $X=5.315 $Y=1.22 $X2=0 $Y2=0
cc_288 N_A3_c_317_n N_VGND_c_636_n 0.00383152f $X=5.745 $Y=1.22 $X2=0 $Y2=0
cc_289 N_A3_c_316_n N_VGND_c_639_n 0.00825283f $X=5.315 $Y=1.22 $X2=0 $Y2=0
cc_290 N_A3_c_317_n N_VGND_c_639_n 0.0075754f $X=5.745 $Y=1.22 $X2=0 $Y2=0
cc_291 N_A3_c_316_n N_A_771_74#_c_741_n 0.0161504f $X=5.315 $Y=1.22 $X2=0 $Y2=0
cc_292 N_A3_c_317_n N_A_771_74#_c_741_n 0.00218762f $X=5.745 $Y=1.22 $X2=0 $Y2=0
cc_293 N_A3_c_319_n N_A_771_74#_c_741_n 0.017248f $X=5.745 $Y=1.492 $X2=0 $Y2=0
cc_294 N_A3_c_316_n N_A_771_74#_c_743_n 0.013408f $X=5.315 $Y=1.22 $X2=0 $Y2=0
cc_295 N_A3_c_317_n N_A_771_74#_c_743_n 3.97481e-19 $X=5.745 $Y=1.22 $X2=0 $Y2=0
cc_296 N_A_27_368#_c_358_n N_Y_M1007_d 0.00245557f $X=1.115 $Y=2.99 $X2=0 $Y2=0
cc_297 N_A_27_368#_c_360_n N_Y_M1015_d 0.00250873f $X=2.115 $Y=2.99 $X2=0 $Y2=0
cc_298 N_A_27_368#_c_358_n N_Y_c_457_n 0.0185424f $X=1.115 $Y=2.99 $X2=0 $Y2=0
cc_299 N_A_27_368#_M1009_s N_Y_c_448_n 0.00250873f $X=1.08 $Y=1.84 $X2=0 $Y2=0
cc_300 N_A_27_368#_c_374_n N_Y_c_448_n 0.0202249f $X=1.28 $Y=2.27 $X2=0 $Y2=0
cc_301 N_A_27_368#_c_360_n N_Y_c_465_n 0.018923f $X=2.115 $Y=2.99 $X2=0 $Y2=0
cc_302 N_A_27_368#_M1019_s N_Y_c_449_n 0.00250873f $X=2.08 $Y=1.84 $X2=0 $Y2=0
cc_303 N_A_27_368#_c_413_p N_Y_c_449_n 0.0192006f $X=2.257 $Y=2.23 $X2=0 $Y2=0
cc_304 N_A_27_368#_c_380_n N_Y_c_449_n 0.0368259f $X=3.405 $Y=2.145 $X2=0 $Y2=0
cc_305 N_A_27_368#_c_380_n N_Y_c_452_n 0.0169206f $X=3.405 $Y=2.145 $X2=0 $Y2=0
cc_306 N_A_27_368#_c_380_n N_VPWR_M1004_d 0.0147605f $X=3.405 $Y=2.145 $X2=-0.19
+ $Y2=1.66
cc_307 N_A_27_368#_c_385_n N_VPWR_M1000_s 0.00489599f $X=4.42 $Y=2.035 $X2=0
+ $Y2=0
cc_308 N_A_27_368#_c_364_n N_VPWR_M1011_d 0.00306736f $X=5.545 $Y=1.805 $X2=0
+ $Y2=0
cc_309 N_A_27_368#_c_360_n N_VPWR_c_525_n 0.0125198f $X=2.115 $Y=2.99 $X2=0
+ $Y2=0
cc_310 N_A_27_368#_c_380_n N_VPWR_c_525_n 0.0481494f $X=3.405 $Y=2.145 $X2=0
+ $Y2=0
cc_311 N_A_27_368#_c_361_n N_VPWR_c_525_n 0.0252395f $X=3.57 $Y=2.465 $X2=0
+ $Y2=0
cc_312 N_A_27_368#_c_361_n N_VPWR_c_526_n 0.0261113f $X=3.57 $Y=2.465 $X2=0
+ $Y2=0
cc_313 N_A_27_368#_c_385_n N_VPWR_c_526_n 0.0214453f $X=4.42 $Y=2.035 $X2=0
+ $Y2=0
cc_314 N_A_27_368#_c_363_n N_VPWR_c_526_n 0.026897f $X=4.585 $Y=2.4 $X2=0 $Y2=0
cc_315 N_A_27_368#_c_363_n N_VPWR_c_527_n 0.0346454f $X=4.585 $Y=2.4 $X2=0 $Y2=0
cc_316 N_A_27_368#_c_364_n N_VPWR_c_527_n 0.0232685f $X=5.545 $Y=1.805 $X2=0
+ $Y2=0
cc_317 N_A_27_368#_c_365_n N_VPWR_c_527_n 0.0353111f $X=5.71 $Y=1.985 $X2=0
+ $Y2=0
cc_318 N_A_27_368#_c_363_n N_VPWR_c_528_n 0.0201714f $X=4.585 $Y=2.4 $X2=0 $Y2=0
cc_319 N_A_27_368#_c_358_n N_VPWR_c_530_n 0.0422607f $X=1.115 $Y=2.99 $X2=0
+ $Y2=0
cc_320 N_A_27_368#_c_359_n N_VPWR_c_530_n 0.0236215f $X=0.445 $Y=2.99 $X2=0
+ $Y2=0
cc_321 N_A_27_368#_c_360_n N_VPWR_c_530_n 0.062706f $X=2.115 $Y=2.99 $X2=0 $Y2=0
cc_322 N_A_27_368#_c_366_n N_VPWR_c_530_n 0.0236039f $X=1.28 $Y=2.99 $X2=0 $Y2=0
cc_323 N_A_27_368#_c_361_n N_VPWR_c_531_n 0.0125859f $X=3.57 $Y=2.465 $X2=0
+ $Y2=0
cc_324 N_A_27_368#_c_365_n N_VPWR_c_532_n 0.0145938f $X=5.71 $Y=1.985 $X2=0
+ $Y2=0
cc_325 N_A_27_368#_c_358_n N_VPWR_c_524_n 0.0238634f $X=1.115 $Y=2.99 $X2=0
+ $Y2=0
cc_326 N_A_27_368#_c_359_n N_VPWR_c_524_n 0.0127839f $X=0.445 $Y=2.99 $X2=0
+ $Y2=0
cc_327 N_A_27_368#_c_360_n N_VPWR_c_524_n 0.0349663f $X=2.115 $Y=2.99 $X2=0
+ $Y2=0
cc_328 N_A_27_368#_c_361_n N_VPWR_c_524_n 0.0103846f $X=3.57 $Y=2.465 $X2=0
+ $Y2=0
cc_329 N_A_27_368#_c_363_n N_VPWR_c_524_n 0.0166633f $X=4.585 $Y=2.4 $X2=0 $Y2=0
cc_330 N_A_27_368#_c_365_n N_VPWR_c_524_n 0.0120466f $X=5.71 $Y=1.985 $X2=0
+ $Y2=0
cc_331 N_A_27_368#_c_366_n N_VPWR_c_524_n 0.012761f $X=1.28 $Y=2.99 $X2=0 $Y2=0
cc_332 N_A_27_368#_c_362_n N_A_771_74#_c_741_n 0.0123321f $X=4.647 $Y=2.12 $X2=0
+ $Y2=0
cc_333 N_A_27_368#_c_364_n N_A_771_74#_c_741_n 0.0242613f $X=5.545 $Y=1.805
+ $X2=0 $Y2=0
cc_334 N_Y_c_449_n N_VPWR_M1004_d 0.00453188f $X=3.005 $Y=1.805 $X2=-0.19
+ $Y2=-0.245
cc_335 N_Y_c_452_n N_VPWR_M1004_d 0.00282171f $X=3.12 $Y=1.72 $X2=-0.19
+ $Y2=-0.245
cc_336 N_Y_c_444_n N_A_27_74#_M1008_s 0.00747698f $X=3.005 $Y=0.925 $X2=0 $Y2=0
cc_337 N_Y_c_448_n N_A_27_74#_c_594_n 0.00590786f $X=1.615 $Y=1.885 $X2=0 $Y2=0
cc_338 N_Y_M1003_d N_A_27_74#_c_596_n 0.00176461f $X=1.48 $Y=0.37 $X2=0 $Y2=0
cc_339 N_Y_c_444_n N_A_27_74#_c_596_n 0.00352531f $X=3.005 $Y=0.925 $X2=0 $Y2=0
cc_340 N_Y_c_472_n N_A_27_74#_c_596_n 0.0154609f $X=1.62 $Y=0.8 $X2=0 $Y2=0
cc_341 N_Y_c_444_n N_A_27_74#_c_598_n 0.0242753f $X=3.005 $Y=0.925 $X2=0 $Y2=0
cc_342 N_Y_c_444_n N_VGND_c_639_n 0.00986599f $X=3.005 $Y=0.925 $X2=0 $Y2=0
cc_343 N_Y_c_444_n N_A_507_74#_M1005_s 0.0052985f $X=3.005 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_344 N_Y_M1005_d N_A_507_74#_c_697_n 0.00176461f $X=2.97 $Y=0.37 $X2=0 $Y2=0
cc_345 N_Y_c_444_n N_A_507_74#_c_697_n 0.0035136f $X=3.005 $Y=0.925 $X2=0 $Y2=0
cc_346 N_Y_c_520_p N_A_507_74#_c_697_n 0.0126348f $X=3.105 $Y=1.01 $X2=0 $Y2=0
cc_347 N_Y_c_445_n N_A_507_74#_c_698_n 0.00523541f $X=3.12 $Y=1.235 $X2=0 $Y2=0
cc_348 N_Y_c_444_n N_A_507_74#_c_701_n 0.0206029f $X=3.005 $Y=0.925 $X2=0 $Y2=0
cc_349 N_Y_c_445_n N_A_771_74#_c_742_n 0.00159757f $X=3.12 $Y=1.235 $X2=0 $Y2=0
cc_350 N_A_27_74#_c_594_n N_VGND_M1010_s 0.00229612f $X=1.105 $Y=1.045 $X2=-0.19
+ $Y2=-0.245
cc_351 N_A_27_74#_c_593_n N_VGND_c_630_n 0.0164982f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_352 N_A_27_74#_c_594_n N_VGND_c_630_n 0.0193595f $X=1.105 $Y=1.045 $X2=0
+ $Y2=0
cc_353 N_A_27_74#_c_597_n N_VGND_c_630_n 0.00814404f $X=1.275 $Y=0.34 $X2=0
+ $Y2=0
cc_354 N_A_27_74#_c_593_n N_VGND_c_634_n 0.011066f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_355 N_A_27_74#_c_596_n N_VGND_c_635_n 0.042902f $X=1.955 $Y=0.34 $X2=0 $Y2=0
cc_356 N_A_27_74#_c_597_n N_VGND_c_635_n 0.0121867f $X=1.275 $Y=0.34 $X2=0 $Y2=0
cc_357 N_A_27_74#_c_598_n N_VGND_c_635_n 0.0226635f $X=2.12 $Y=0.34 $X2=0 $Y2=0
cc_358 N_A_27_74#_c_593_n N_VGND_c_639_n 0.00915947f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_359 N_A_27_74#_c_596_n N_VGND_c_639_n 0.0241973f $X=1.955 $Y=0.34 $X2=0 $Y2=0
cc_360 N_A_27_74#_c_597_n N_VGND_c_639_n 0.00660921f $X=1.275 $Y=0.34 $X2=0
+ $Y2=0
cc_361 N_A_27_74#_c_598_n N_VGND_c_639_n 0.0125932f $X=2.12 $Y=0.34 $X2=0 $Y2=0
cc_362 N_A_27_74#_c_598_n N_A_507_74#_c_701_n 0.0279789f $X=2.12 $Y=0.34 $X2=0
+ $Y2=0
cc_363 N_VGND_c_635_n N_A_507_74#_c_697_n 0.0333877f $X=4.935 $Y=0 $X2=0 $Y2=0
cc_364 N_VGND_c_639_n N_A_507_74#_c_697_n 0.0187857f $X=6 $Y=0 $X2=0 $Y2=0
cc_365 N_VGND_c_631_n N_A_507_74#_c_699_n 0.011925f $X=5.1 $Y=0.675 $X2=0 $Y2=0
cc_366 N_VGND_c_635_n N_A_507_74#_c_699_n 0.065612f $X=4.935 $Y=0 $X2=0 $Y2=0
cc_367 N_VGND_c_639_n N_A_507_74#_c_699_n 0.0365975f $X=6 $Y=0 $X2=0 $Y2=0
cc_368 N_VGND_c_631_n N_A_507_74#_c_700_n 0.0273691f $X=5.1 $Y=0.675 $X2=0 $Y2=0
cc_369 N_VGND_c_635_n N_A_507_74#_c_701_n 0.0225845f $X=4.935 $Y=0 $X2=0 $Y2=0
cc_370 N_VGND_c_639_n N_A_507_74#_c_701_n 0.0124836f $X=6 $Y=0 $X2=0 $Y2=0
cc_371 N_VGND_c_635_n N_A_507_74#_c_702_n 0.0235688f $X=4.935 $Y=0 $X2=0 $Y2=0
cc_372 N_VGND_c_639_n N_A_507_74#_c_702_n 0.0127152f $X=6 $Y=0 $X2=0 $Y2=0
cc_373 N_VGND_M1002_s N_A_771_74#_c_741_n 0.00299905f $X=4.955 $Y=0.37 $X2=0
+ $Y2=0
cc_374 N_VGND_c_631_n N_A_771_74#_c_741_n 0.0201544f $X=5.1 $Y=0.675 $X2=0 $Y2=0
cc_375 N_VGND_c_631_n N_A_771_74#_c_743_n 0.0175587f $X=5.1 $Y=0.675 $X2=0 $Y2=0
cc_376 N_VGND_c_633_n N_A_771_74#_c_743_n 0.0243832f $X=5.96 $Y=0.515 $X2=0
+ $Y2=0
cc_377 N_VGND_c_636_n N_A_771_74#_c_743_n 0.0109942f $X=5.795 $Y=0 $X2=0 $Y2=0
cc_378 N_VGND_c_639_n N_A_771_74#_c_743_n 0.00904371f $X=6 $Y=0 $X2=0 $Y2=0
cc_379 N_A_507_74#_c_699_n N_A_771_74#_M1013_s 0.0030917f $X=4.375 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_380 N_A_507_74#_c_699_n N_A_771_74#_c_764_n 0.0211419f $X=4.375 $Y=0.34 $X2=0
+ $Y2=0
cc_381 N_A_507_74#_M1014_d N_A_771_74#_c_741_n 0.00299905f $X=4.4 $Y=0.37 $X2=0
+ $Y2=0
cc_382 N_A_507_74#_c_699_n N_A_771_74#_c_741_n 0.00304353f $X=4.375 $Y=0.34
+ $X2=0 $Y2=0
cc_383 N_A_507_74#_c_700_n N_A_771_74#_c_741_n 0.021673f $X=4.54 $Y=0.675 $X2=0
+ $Y2=0
cc_384 N_A_507_74#_c_698_n N_A_771_74#_c_742_n 0.00585736f $X=3.54 $Y=0.515
+ $X2=0 $Y2=0
