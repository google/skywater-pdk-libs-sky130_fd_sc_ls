* File: sky130_fd_sc_ls__or4b_4.pex.spice
* Created: Fri Aug 28 14:00:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__OR4B_4%B 2 5 6 8 10 11 13 14 16 20 22 23 27 29 34 41
c77 20 0 1.33875e-19 $X=1.87 $Y=1.385
r78 28 34 4.8455 $w=4.38e-07 $l=1.85e-07 $layer=LI1_cond $X=0.43 $Y=1.33
+ $X2=0.615 $Y2=1.33
r79 27 30 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.43 $Y=1.385
+ $X2=0.43 $Y2=1.55
r80 27 29 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.43 $Y=1.385
+ $X2=0.43 $Y2=1.22
r81 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.43
+ $Y=1.385 $X2=0.43 $Y2=1.385
r82 23 41 7.52572 $w=4.38e-07 $l=1.15e-07 $layer=LI1_cond $X=0.72 $Y=1.33
+ $X2=0.835 $Y2=1.33
r83 23 34 2.75015 $w=4.38e-07 $l=1.05e-07 $layer=LI1_cond $X=0.72 $Y=1.33
+ $X2=0.615 $Y2=1.33
r84 22 28 4.97646 $w=4.38e-07 $l=1.9e-07 $layer=LI1_cond $X=0.24 $Y=1.33
+ $X2=0.43 $Y2=1.33
r85 20 33 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.87 $Y=1.385
+ $X2=1.87 $Y2=1.55
r86 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.87
+ $Y=1.385 $X2=1.87 $Y2=1.385
r87 16 19 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=1.87 $Y=1.195
+ $X2=1.87 $Y2=1.385
r88 14 16 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.705 $Y=1.195
+ $X2=1.87 $Y2=1.195
r89 14 41 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=1.705 $Y=1.195
+ $X2=0.835 $Y2=1.195
r90 11 13 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.905 $Y=1.885
+ $X2=1.905 $Y2=2.46
r91 10 11 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.905 $Y=1.795
+ $X2=1.905 $Y2=1.885
r92 10 33 95.2339 $w=1.8e-07 $l=2.45e-07 $layer=POLY_cond $X=1.905 $Y=1.795
+ $X2=1.905 $Y2=1.55
r93 6 8 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.505 $Y=1.885
+ $X2=0.505 $Y2=2.46
r94 5 29 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.495 $Y=0.74
+ $X2=0.495 $Y2=1.22
r95 2 6 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.505 $Y=1.795 $X2=0.505
+ $Y2=1.885
r96 2 30 95.2339 $w=1.8e-07 $l=2.45e-07 $layer=POLY_cond $X=0.505 $Y=1.795
+ $X2=0.505 $Y2=1.55
.ends

.subckt PM_SKY130_FD_SC_LS__OR4B_4%A 1 3 6 8 10 11 16
c48 1 0 4.75553e-20 $X=0.955 $Y=1.885
r49 16 18 29.0436 $w=3.9e-07 $l=2.35e-07 $layer=POLY_cond $X=1.17 $Y=1.667
+ $X2=1.405 $Y2=1.667
r50 14 16 12.9769 $w=3.9e-07 $l=1.05e-07 $layer=POLY_cond $X=1.065 $Y=1.667
+ $X2=1.17 $Y2=1.667
r51 13 14 13.5949 $w=3.9e-07 $l=1.1e-07 $layer=POLY_cond $X=0.955 $Y=1.667
+ $X2=1.065 $Y2=1.667
r52 11 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.17
+ $Y=1.615 $X2=1.17 $Y2=1.615
r53 8 18 25.2441 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=1.405 $Y=1.885
+ $X2=1.405 $Y2=1.667
r54 8 10 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.405 $Y=1.885
+ $X2=1.405 $Y2=2.46
r55 4 14 25.2441 $w=1.5e-07 $l=2.17e-07 $layer=POLY_cond $X=1.065 $Y=1.45
+ $X2=1.065 $Y2=1.667
r56 4 6 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.065 $Y=1.45
+ $X2=1.065 $Y2=0.74
r57 1 13 25.2441 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=0.955 $Y=1.885
+ $X2=0.955 $Y2=1.667
r58 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.955 $Y=1.885
+ $X2=0.955 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_LS__OR4B_4%C 3 5 6 8 10 11 13 14 15 17 18 20 23 25 30 36
c95 25 0 2.8262e-20 $X=2.41 $Y=1.22
c96 18 0 9.18809e-20 $X=4.08 $Y=1.295
c97 10 0 6.84608e-20 $X=3.805 $Y=1.795
c98 6 0 1.28327e-19 $X=2.405 $Y=1.885
r99 27 30 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=3.805 $Y=1.345
+ $X2=4.03 $Y2=1.345
r100 24 36 4.58497 $w=5.98e-07 $l=2.3e-07 $layer=LI1_cond $X=2.41 $Y=1.48
+ $X2=2.64 $Y2=1.48
r101 23 26 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.41 $Y=1.385
+ $X2=2.41 $Y2=1.55
r102 23 25 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.41 $Y=1.385
+ $X2=2.41 $Y2=1.22
r103 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.41
+ $Y=1.385 $X2=2.41 $Y2=1.385
r104 20 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=1.295
+ $X2=2.64 $Y2=1.295
r105 18 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.03
+ $Y=1.345 $X2=4.03 $Y2=1.345
r106 17 18 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=1.295
+ $X2=4.08 $Y2=1.295
r107 15 20 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.785 $Y=1.295
+ $X2=2.64 $Y2=1.295
r108 14 17 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.935 $Y=1.295
+ $X2=4.08 $Y2=1.295
r109 14 15 1.42326 $w=1.4e-07 $l=1.15e-06 $layer=MET1_cond $X=3.935 $Y=1.295
+ $X2=2.785 $Y2=1.295
r110 11 13 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.805 $Y=1.885
+ $X2=3.805 $Y2=2.46
r111 10 11 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.805 $Y=1.795
+ $X2=3.805 $Y2=1.885
r112 9 27 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.805 $Y=1.51
+ $X2=3.805 $Y2=1.345
r113 9 10 110.782 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=3.805 $Y=1.51
+ $X2=3.805 $Y2=1.795
r114 6 8 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.405 $Y=1.885
+ $X2=2.405 $Y2=2.46
r115 5 6 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.405 $Y=1.795
+ $X2=2.405 $Y2=1.885
r116 5 26 95.2339 $w=1.8e-07 $l=2.45e-07 $layer=POLY_cond $X=2.405 $Y=1.795
+ $X2=2.405 $Y2=1.55
r117 3 25 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.32 $Y=0.74 $X2=2.32
+ $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_LS__OR4B_4%A_563_48# 1 2 9 11 13 14 16 18 21 24 26 27 30
+ 40
c94 40 0 3.30667e-19 $X=3.355 $Y=1.677
r95 40 41 5.79947 $w=3.74e-07 $l=4.5e-08 $layer=POLY_cond $X=3.355 $Y=1.677
+ $X2=3.4 $Y2=1.677
r96 37 38 1.93316 $w=3.74e-07 $l=1.5e-08 $layer=POLY_cond $X=2.89 $Y=1.677
+ $X2=2.905 $Y2=1.677
r97 36 40 1.93316 $w=3.74e-07 $l=1.5e-08 $layer=POLY_cond $X=3.34 $Y=1.677
+ $X2=3.355 $Y2=1.677
r98 36 38 56.0615 $w=3.74e-07 $l=4.35e-07 $layer=POLY_cond $X=3.34 $Y=1.677
+ $X2=2.905 $Y2=1.677
r99 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.34
+ $Y=1.635 $X2=3.34 $Y2=1.635
r100 30 32 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=4.59 $Y=1.985
+ $X2=4.59 $Y2=2.695
r101 28 30 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=4.59 $Y=1.89
+ $X2=4.59 $Y2=1.985
r102 27 35 13.3429 $w=3.68e-07 $l=3.51994e-07 $layer=LI1_cond $X=3.635 $Y=1.805
+ $X2=3.34 $Y2=1.68
r103 26 28 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.425 $Y=1.805
+ $X2=4.59 $Y2=1.89
r104 26 27 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=4.425 $Y=1.805
+ $X2=3.635 $Y2=1.805
r105 21 42 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=3.605 $Y=0.505
+ $X2=3.4 $Y2=0.505
r106 20 24 27.7634 $w=3.28e-07 $l=7.95e-07 $layer=LI1_cond $X=3.605 $Y=0.505
+ $X2=4.4 $Y2=0.505
r107 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.605
+ $Y=0.505 $X2=3.605 $Y2=0.505
r108 18 41 24.2268 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.4 $Y=1.47
+ $X2=3.4 $Y2=1.677
r109 17 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.4 $Y=0.67
+ $X2=3.4 $Y2=0.505
r110 17 18 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=3.4 $Y=0.67 $X2=3.4
+ $Y2=1.47
r111 14 40 24.2268 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.355 $Y=1.885
+ $X2=3.355 $Y2=1.677
r112 14 16 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.355 $Y=1.885
+ $X2=3.355 $Y2=2.46
r113 11 38 24.2268 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.905 $Y=1.885
+ $X2=2.905 $Y2=1.677
r114 11 13 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.905 $Y=1.885
+ $X2=2.905 $Y2=2.46
r115 7 37 24.2268 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.89 $Y=1.47
+ $X2=2.89 $Y2=1.677
r116 7 9 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=2.89 $Y=1.47 $X2=2.89
+ $Y2=0.74
r117 2 32 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=4.445
+ $Y=1.84 $X2=4.59 $Y2=2.695
r118 2 30 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=4.445
+ $Y=1.84 $X2=4.59 $Y2=1.985
r119 1 24 91 $w=1.7e-07 $l=5.88048e-07 $layer=licon1_NDIFF $count=2 $X=3.88
+ $Y=0.36 $X2=4.4 $Y2=0.505
.ends

.subckt PM_SKY130_FD_SC_LS__OR4B_4%D_N 1 3 4 6 7
c36 1 0 5.98002e-20 $X=4.695 $Y=1.22
r37 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.65
+ $Y=1.385 $X2=4.65 $Y2=1.385
r38 7 11 2.80324 $w=3.68e-07 $l=9e-08 $layer=LI1_cond $X=4.63 $Y=1.295 $X2=4.63
+ $Y2=1.385
r39 4 10 70.4572 $w=3.25e-07 $l=4.3589e-07 $layer=POLY_cond $X=4.815 $Y=1.765
+ $X2=4.695 $Y2=1.385
r40 4 6 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=4.815 $Y=1.765
+ $X2=4.815 $Y2=2.34
r41 1 10 38.571 $w=3.25e-07 $l=1.65e-07 $layer=POLY_cond $X=4.695 $Y=1.22
+ $X2=4.695 $Y2=1.385
r42 1 3 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=4.695 $Y=1.22
+ $X2=4.695 $Y2=0.79
.ends

.subckt PM_SKY130_FD_SC_LS__OR4B_4%A_27_74# 1 2 3 4 15 17 19 22 24 26 27 29 32
+ 34 36 39 43 46 47 48 51 55 58 59 62 63 68 71 74 81 91
c194 91 0 1.47325e-19 $X=6.7 $Y=1.542
c195 59 0 1.67773e-19 $X=4.985 $Y=0.925
c196 58 0 9.67228e-20 $X=2.98 $Y=2.02
r197 91 92 0.640957 $w=3.76e-07 $l=5e-09 $layer=POLY_cond $X=6.7 $Y=1.542
+ $X2=6.705 $Y2=1.542
r198 90 91 54.4814 $w=3.76e-07 $l=4.25e-07 $layer=POLY_cond $X=6.275 $Y=1.542
+ $X2=6.7 $Y2=1.542
r199 89 90 3.20479 $w=3.76e-07 $l=2.5e-08 $layer=POLY_cond $X=6.25 $Y=1.542
+ $X2=6.275 $Y2=1.542
r200 86 87 3.20479 $w=3.76e-07 $l=2.5e-08 $layer=POLY_cond $X=5.775 $Y=1.542
+ $X2=5.8 $Y2=1.542
r201 85 86 54.4814 $w=3.76e-07 $l=4.25e-07 $layer=POLY_cond $X=5.35 $Y=1.542
+ $X2=5.775 $Y2=1.542
r202 78 81 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=2.98 $Y=2.105
+ $X2=3.13 $Y2=2.105
r203 76 77 9.78374 $w=3.73e-07 $l=2.05e-07 $layer=LI1_cond $X=3.082 $Y=0.925
+ $X2=3.082 $Y2=1.13
r204 73 74 10.0909 $w=5.88e-07 $l=1.65e-07 $layer=LI1_cond $X=2.035 $Y=0.645
+ $X2=2.2 $Y2=0.645
r205 69 89 33.3298 $w=3.76e-07 $l=2.6e-07 $layer=POLY_cond $X=5.99 $Y=1.542
+ $X2=6.25 $Y2=1.542
r206 69 87 24.3564 $w=3.76e-07 $l=1.9e-07 $layer=POLY_cond $X=5.99 $Y=1.542
+ $X2=5.8 $Y2=1.542
r207 68 69 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=5.99
+ $Y=1.485 $X2=5.99 $Y2=1.485
r208 66 85 5.12766 $w=3.76e-07 $l=4e-08 $layer=POLY_cond $X=5.31 $Y=1.542
+ $X2=5.35 $Y2=1.542
r209 66 83 11.5372 $w=3.76e-07 $l=9e-08 $layer=POLY_cond $X=5.31 $Y=1.542
+ $X2=5.22 $Y2=1.542
r210 65 68 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=5.31 $Y=1.485
+ $X2=5.99 $Y2=1.485
r211 65 66 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=5.31
+ $Y=1.485 $X2=5.31 $Y2=1.485
r212 63 65 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=5.155 $Y=1.485
+ $X2=5.31 $Y2=1.485
r213 62 63 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.07 $Y=1.32
+ $X2=5.155 $Y2=1.485
r214 61 62 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=5.07 $Y=1.01
+ $X2=5.07 $Y2=1.32
r215 60 76 5.38787 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=3.27 $Y=0.925
+ $X2=3.082 $Y2=0.925
r216 59 61 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.985 $Y=0.925
+ $X2=5.07 $Y2=1.01
r217 59 60 111.888 $w=1.68e-07 $l=1.715e-06 $layer=LI1_cond $X=4.985 $Y=0.925
+ $X2=3.27 $Y2=0.925
r218 58 78 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.98 $Y=2.02
+ $X2=2.98 $Y2=2.105
r219 58 77 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=2.98 $Y=2.02
+ $X2=2.98 $Y2=1.13
r220 53 55 7.83661 $w=3.73e-07 $l=2.55e-07 $layer=LI1_cond $X=3.082 $Y=0.77
+ $X2=3.082 $Y2=0.515
r221 51 76 2.15123 $w=3.73e-07 $l=7e-08 $layer=LI1_cond $X=3.082 $Y=0.855
+ $X2=3.082 $Y2=0.925
r222 51 53 2.6122 $w=3.73e-07 $l=8.5e-08 $layer=LI1_cond $X=3.082 $Y=0.855
+ $X2=3.082 $Y2=0.77
r223 51 74 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=2.895 $Y=0.855
+ $X2=2.2 $Y2=0.855
r224 48 71 12.7264 $w=5.88e-07 $l=2.95e-07 $layer=LI1_cond $X=1.41 $Y=0.645
+ $X2=1.115 $Y2=0.645
r225 48 50 4.96677 $w=5.88e-07 $l=2.45e-07 $layer=LI1_cond $X=1.41 $Y=0.645
+ $X2=1.655 $Y2=0.645
r226 47 73 2.63543 $w=5.88e-07 $l=1.3e-07 $layer=LI1_cond $X=1.905 $Y=0.645
+ $X2=2.035 $Y2=0.645
r227 47 50 5.06813 $w=5.88e-07 $l=2.5e-07 $layer=LI1_cond $X=1.905 $Y=0.645
+ $X2=1.655 $Y2=0.645
r228 46 71 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.445 $Y=0.855
+ $X2=1.115 $Y2=0.855
r229 41 46 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=0.77
+ $X2=0.445 $Y2=0.855
r230 41 43 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=0.28 $Y=0.77
+ $X2=0.28 $Y2=0.515
r231 37 92 24.356 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=6.705 $Y=1.32
+ $X2=6.705 $Y2=1.542
r232 37 39 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.705 $Y=1.32
+ $X2=6.705 $Y2=0.74
r233 34 91 24.356 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=6.7 $Y=1.765
+ $X2=6.7 $Y2=1.542
r234 34 36 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.7 $Y=1.765
+ $X2=6.7 $Y2=2.4
r235 30 90 24.356 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=6.275 $Y=1.32
+ $X2=6.275 $Y2=1.542
r236 30 32 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.275 $Y=1.32
+ $X2=6.275 $Y2=0.74
r237 27 89 24.356 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=6.25 $Y=1.765
+ $X2=6.25 $Y2=1.542
r238 27 29 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.25 $Y=1.765
+ $X2=6.25 $Y2=2.4
r239 24 87 24.356 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=5.8 $Y=1.765
+ $X2=5.8 $Y2=1.542
r240 24 26 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.8 $Y=1.765
+ $X2=5.8 $Y2=2.4
r241 20 86 24.356 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=5.775 $Y=1.32
+ $X2=5.775 $Y2=1.542
r242 20 22 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=5.775 $Y=1.32
+ $X2=5.775 $Y2=0.74
r243 17 85 24.356 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=5.35 $Y=1.765
+ $X2=5.35 $Y2=1.542
r244 17 19 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.35 $Y=1.765
+ $X2=5.35 $Y2=2.4
r245 13 83 24.356 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=5.22 $Y=1.32
+ $X2=5.22 $Y2=1.542
r246 13 15 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=5.22 $Y=1.32
+ $X2=5.22 $Y2=0.74
r247 4 81 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.98
+ $Y=1.96 $X2=3.13 $Y2=2.105
r248 3 55 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.965
+ $Y=0.37 $X2=3.105 $Y2=0.515
r249 2 73 91 $w=1.7e-07 $l=9.6478e-07 $layer=licon1_NDIFF $count=2 $X=1.14
+ $Y=0.37 $X2=2.035 $Y2=0.515
r250 2 50 45.5 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_NDIFF $count=4 $X=1.14
+ $Y=0.37 $X2=1.655 $Y2=0.515
r251 1 43 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__OR4B_4%A_27_392# 1 2 3 10 12 14 16 17 20 22 26 30 36
+ 37
c73 22 0 1.30813e-19 $X=3.945 $Y=2.445
c74 16 0 1.33875e-19 $X=2.18 $Y=2.12
c75 10 0 4.75553e-20 $X=0.28 $Y=2.12
r76 28 37 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.07 $Y=2.53 $X2=4.07
+ $Y2=2.445
r77 28 30 13.1378 $w=2.48e-07 $l=2.85e-07 $layer=LI1_cond $X=4.07 $Y=2.53
+ $X2=4.07 $Y2=2.815
r78 24 37 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.07 $Y=2.36 $X2=4.07
+ $Y2=2.445
r79 24 26 6.22319 $w=2.48e-07 $l=1.35e-07 $layer=LI1_cond $X=4.07 $Y=2.36
+ $X2=4.07 $Y2=2.225
r80 23 36 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.345 $Y=2.445
+ $X2=2.18 $Y2=2.445
r81 22 37 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.945 $Y=2.445
+ $X2=4.07 $Y2=2.445
r82 22 23 104.385 $w=1.68e-07 $l=1.6e-06 $layer=LI1_cond $X=3.945 $Y=2.445
+ $X2=2.345 $Y2=2.445
r83 18 36 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.18 $Y=2.53 $X2=2.18
+ $Y2=2.445
r84 18 20 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=2.18 $Y=2.53
+ $X2=2.18 $Y2=2.815
r85 17 36 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.18 $Y=2.36 $X2=2.18
+ $Y2=2.445
r86 16 35 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.18 $Y=2.12 $X2=2.18
+ $Y2=2.035
r87 16 17 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=2.18 $Y=2.12 $X2=2.18
+ $Y2=2.36
r88 15 33 5.07788 $w=1.7e-07 $l=1.67481e-07 $layer=LI1_cond $X=0.445 $Y=2.035
+ $X2=0.28 $Y2=2.03
r89 14 35 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.015 $Y=2.035
+ $X2=2.18 $Y2=2.035
r90 14 15 102.428 $w=1.68e-07 $l=1.57e-06 $layer=LI1_cond $X=2.015 $Y=2.035
+ $X2=0.445 $Y2=2.035
r91 10 33 2.68829 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=0.28 $Y=2.12 $X2=0.28
+ $Y2=2.03
r92 10 12 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=0.28 $Y=2.12
+ $X2=0.28 $Y2=2.815
r93 3 30 600 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=3.88
+ $Y=1.96 $X2=4.03 $Y2=2.815
r94 3 26 600 $w=1.7e-07 $l=3.31625e-07 $layer=licon1_PDIFF $count=1 $X=3.88
+ $Y=1.96 $X2=4.03 $Y2=2.225
r95 2 35 400 $w=1.7e-07 $l=2.66458e-07 $layer=licon1_PDIFF $count=1 $X=1.98
+ $Y=1.96 $X2=2.18 $Y2=2.115
r96 2 20 400 $w=1.7e-07 $l=9.4975e-07 $layer=licon1_PDIFF $count=1 $X=1.98
+ $Y=1.96 $X2=2.18 $Y2=2.815
r97 1 33 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.28 $Y2=2.105
r98 1 12 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.28 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_LS__OR4B_4%A_116_392# 1 2 9 14 16
c23 16 0 1.28327e-19 $X=1.68 $Y=2.455
r24 10 14 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=2.375
+ $X2=0.73 $Y2=2.375
r25 9 16 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.515 $Y=2.375
+ $X2=1.68 $Y2=2.375
r26 9 10 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.515 $Y=2.375
+ $X2=0.815 $Y2=2.375
r27 2 16 300 $w=1.7e-07 $l=5.86536e-07 $layer=licon1_PDIFF $count=2 $X=1.48
+ $Y=1.96 $X2=1.68 $Y2=2.455
r28 1 14 300 $w=1.7e-07 $l=5.65044e-07 $layer=licon1_PDIFF $count=2 $X=0.58
+ $Y=1.96 $X2=0.73 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_LS__OR4B_4%VPWR 1 2 3 4 15 19 25 27 29 31 33 38 43 48 54
+ 57 60 64
r90 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r91 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r92 57 58 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r93 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r94 52 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6.96 $Y2=3.33
r95 52 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33 $X2=6
+ $Y2=3.33
r96 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r97 49 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.19 $Y=3.33
+ $X2=6.025 $Y2=3.33
r98 49 51 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=6.19 $Y=3.33
+ $X2=6.48 $Y2=3.33
r99 48 63 4.746 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=6.76 $Y=3.33 $X2=6.98
+ $Y2=3.33
r100 48 51 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=6.76 $Y=3.33
+ $X2=6.48 $Y2=3.33
r101 47 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33 $X2=6
+ $Y2=3.33
r102 47 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=5.04 $Y2=3.33
r103 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r104 44 57 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.21 $Y=3.33
+ $X2=5.085 $Y2=3.33
r105 44 46 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=5.21 $Y=3.33
+ $X2=5.52 $Y2=3.33
r106 43 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.86 $Y=3.33
+ $X2=6.025 $Y2=3.33
r107 43 46 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=5.86 $Y=3.33
+ $X2=5.52 $Y2=3.33
r108 42 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r109 41 42 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r110 39 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.345 $Y=3.33
+ $X2=1.18 $Y2=3.33
r111 39 41 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.345 $Y=3.33
+ $X2=1.68 $Y2=3.33
r112 38 57 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.96 $Y=3.33
+ $X2=5.085 $Y2=3.33
r113 38 41 213.989 $w=1.68e-07 $l=3.28e-06 $layer=LI1_cond $X=4.96 $Y=3.33
+ $X2=1.68 $Y2=3.33
r114 36 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r115 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r116 33 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.015 $Y=3.33
+ $X2=1.18 $Y2=3.33
r117 33 35 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.015 $Y=3.33
+ $X2=0.72 $Y2=3.33
r118 31 58 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=5.04 $Y2=3.33
r119 31 42 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=1.68 $Y2=3.33
r120 27 63 3.02018 $w=3.3e-07 $l=1.09087e-07 $layer=LI1_cond $X=6.925 $Y=3.245
+ $X2=6.98 $Y2=3.33
r121 27 29 29.3349 $w=3.28e-07 $l=8.4e-07 $layer=LI1_cond $X=6.925 $Y=3.245
+ $X2=6.925 $Y2=2.405
r122 23 60 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.025 $Y=3.245
+ $X2=6.025 $Y2=3.33
r123 23 25 29.3349 $w=3.28e-07 $l=8.4e-07 $layer=LI1_cond $X=6.025 $Y=3.245
+ $X2=6.025 $Y2=2.405
r124 19 22 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=5.085 $Y=1.985
+ $X2=5.085 $Y2=2.815
r125 17 57 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.085 $Y=3.245
+ $X2=5.085 $Y2=3.33
r126 17 22 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=5.085 $Y=3.245
+ $X2=5.085 $Y2=2.815
r127 13 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.18 $Y=3.245
+ $X2=1.18 $Y2=3.33
r128 13 15 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=1.18 $Y=3.245
+ $X2=1.18 $Y2=2.805
r129 4 29 300 $w=1.7e-07 $l=6.3559e-07 $layer=licon1_PDIFF $count=2 $X=6.775
+ $Y=1.84 $X2=6.925 $Y2=2.405
r130 3 25 300 $w=1.7e-07 $l=6.3559e-07 $layer=licon1_PDIFF $count=2 $X=5.875
+ $Y=1.84 $X2=6.025 $Y2=2.405
r131 2 22 600 $w=1.7e-07 $l=1.08616e-06 $layer=licon1_PDIFF $count=1 $X=4.89
+ $Y=1.84 $X2=5.125 $Y2=2.815
r132 2 19 300 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=2 $X=4.89
+ $Y=1.84 $X2=5.125 $Y2=1.985
r133 1 15 600 $w=1.7e-07 $l=9.16938e-07 $layer=licon1_PDIFF $count=1 $X=1.03
+ $Y=1.96 $X2=1.18 $Y2=2.805
.ends

.subckt PM_SKY130_FD_SC_LS__OR4B_4%A_496_392# 1 2 11
r13 8 11 37.0428 $w=2.78e-07 $l=9e-07 $layer=LI1_cond $X=2.68 $Y=2.84 $X2=3.58
+ $Y2=2.84
r14 2 11 600 $w=1.7e-07 $l=9.11921e-07 $layer=licon1_PDIFF $count=1 $X=3.43
+ $Y=1.96 $X2=3.58 $Y2=2.8
r15 1 8 600 $w=1.7e-07 $l=9.34666e-07 $layer=licon1_PDIFF $count=1 $X=2.48
+ $Y=1.96 $X2=2.68 $Y2=2.8
.ends

.subckt PM_SKY130_FD_SC_LS__OR4B_4%X 1 2 3 4 15 17 19 21 22 23 27 33 36 39 40 41
+ 42 43
c77 42 0 1.79001e-19 $X=6.48 $Y=2.035
c78 36 0 1.8329e-19 $X=6.51 $Y=1.82
r79 43 46 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=6.96 $Y=1.985
+ $X2=6.655 $Y2=1.985
r80 42 46 2.3561 $w=3.3e-07 $l=1.48e-07 $layer=LI1_cond $X=6.507 $Y=1.985
+ $X2=6.655 $Y2=1.985
r81 40 41 7.00677 $w=2.88e-07 $l=1.7e-07 $layer=LI1_cond $X=6.49 $Y=1.3 $X2=6.49
+ $Y2=1.47
r82 36 42 3.80668 $w=2.9e-07 $l=1.66493e-07 $layer=LI1_cond $X=6.51 $Y=1.82
+ $X2=6.507 $Y2=1.985
r83 36 41 13.9088 $w=2.88e-07 $l=3.5e-07 $layer=LI1_cond $X=6.51 $Y=1.82
+ $X2=6.51 $Y2=1.47
r84 31 42 3.80668 $w=2.3e-07 $l=1.80291e-07 $layer=LI1_cond $X=6.475 $Y=2.15
+ $X2=6.507 $Y2=1.985
r85 31 33 12.5266 $w=2.28e-07 $l=2.5e-07 $layer=LI1_cond $X=6.475 $Y=2.15
+ $X2=6.475 $Y2=2.4
r86 29 39 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.45 $Y=1.15 $X2=6.45
+ $Y2=1.065
r87 29 40 6.91466 $w=2.48e-07 $l=1.5e-07 $layer=LI1_cond $X=6.45 $Y=1.15
+ $X2=6.45 $Y2=1.3
r88 25 39 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.45 $Y=0.98 $X2=6.45
+ $Y2=1.065
r89 25 27 21.4354 $w=2.48e-07 $l=4.65e-07 $layer=LI1_cond $X=6.45 $Y=0.98
+ $X2=6.45 $Y2=0.515
r90 24 38 3.1563 $w=3.3e-07 $l=1.4e-07 $layer=LI1_cond $X=5.69 $Y=1.985 $X2=5.55
+ $Y2=1.985
r91 23 42 2.3561 $w=3.3e-07 $l=1.47e-07 $layer=LI1_cond $X=6.36 $Y=1.985
+ $X2=6.507 $Y2=1.985
r92 23 24 23.3981 $w=3.28e-07 $l=6.7e-07 $layer=LI1_cond $X=6.36 $Y=1.985
+ $X2=5.69 $Y2=1.985
r93 21 39 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.325 $Y=1.065
+ $X2=6.45 $Y2=1.065
r94 21 22 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.325 $Y=1.065
+ $X2=5.655 $Y2=1.065
r95 17 38 3.71993 $w=2.8e-07 $l=1.65e-07 $layer=LI1_cond $X=5.55 $Y=2.15
+ $X2=5.55 $Y2=1.985
r96 17 19 10.2897 $w=2.78e-07 $l=2.5e-07 $layer=LI1_cond $X=5.55 $Y=2.15
+ $X2=5.55 $Y2=2.4
r97 13 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.49 $Y=0.98
+ $X2=5.655 $Y2=1.065
r98 13 15 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=5.49 $Y=0.98
+ $X2=5.49 $Y2=0.515
r99 4 42 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=6.325
+ $Y=1.84 $X2=6.475 $Y2=1.985
r100 4 33 300 $w=1.7e-07 $l=6.30555e-07 $layer=licon1_PDIFF $count=2 $X=6.325
+ $Y=1.84 $X2=6.475 $Y2=2.4
r101 3 38 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=5.425
+ $Y=1.84 $X2=5.575 $Y2=1.985
r102 3 19 300 $w=1.7e-07 $l=6.30555e-07 $layer=licon1_PDIFF $count=2 $X=5.425
+ $Y=1.84 $X2=5.575 $Y2=2.4
r103 2 27 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.35
+ $Y=0.37 $X2=6.49 $Y2=0.515
r104 1 15 91 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_NDIFF $count=2 $X=5.295
+ $Y=0.37 $X2=5.49 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__OR4B_4%VGND 1 2 3 4 5 18 22 26 30 32 34 36 38 43 51
+ 59 64 70 73 76 79 83
r83 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r84 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r85 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r86 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r87 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r88 68 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6.96
+ $Y2=0
r89 68 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r90 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r91 65 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.155 $Y=0 $X2=5.99
+ $Y2=0
r92 65 67 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=6.155 $Y=0 $X2=6.48
+ $Y2=0
r93 64 82 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=6.755 $Y=0 $X2=6.977
+ $Y2=0
r94 64 67 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.755 $Y=0 $X2=6.48
+ $Y2=0
r95 63 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r96 63 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r97 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r98 60 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.155 $Y=0 $X2=4.99
+ $Y2=0
r99 60 62 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=5.155 $Y=0 $X2=5.52
+ $Y2=0
r100 59 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.825 $Y=0 $X2=5.99
+ $Y2=0
r101 59 62 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.825 $Y=0
+ $X2=5.52 $Y2=0
r102 58 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r103 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r104 55 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r105 54 57 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=3.12 $Y=0 $X2=4.56
+ $Y2=0
r106 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r107 52 73 9.05715 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=2.725 $Y=0
+ $X2=2.547 $Y2=0
r108 52 54 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=2.725 $Y=0
+ $X2=3.12 $Y2=0
r109 51 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.825 $Y=0 $X2=4.99
+ $Y2=0
r110 51 57 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=4.825 $Y=0
+ $X2=4.56 $Y2=0
r111 50 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r112 49 50 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r113 47 50 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r114 47 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r115 46 49 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r116 46 47 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r117 44 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=0.78
+ $Y2=0
r118 44 46 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=1.2
+ $Y2=0
r119 43 73 9.05715 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=2.37 $Y=0 $X2=2.547
+ $Y2=0
r120 43 49 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=2.37 $Y=0 $X2=2.16
+ $Y2=0
r121 41 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r122 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r123 38 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.78
+ $Y2=0
r124 38 40 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=0
+ $X2=0.24 $Y2=0
r125 36 58 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r126 36 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r127 32 82 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=6.92 $Y=0.085
+ $X2=6.977 $Y2=0
r128 32 34 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=6.92 $Y=0.085
+ $X2=6.92 $Y2=0.515
r129 28 79 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.99 $Y=0.085
+ $X2=5.99 $Y2=0
r130 28 30 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=5.99 $Y=0.085
+ $X2=5.99 $Y2=0.58
r131 24 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.99 $Y=0.085
+ $X2=4.99 $Y2=0
r132 24 26 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=4.99 $Y=0.085
+ $X2=4.99 $Y2=0.55
r133 20 73 1.11826 $w=3.55e-07 $l=8.5e-08 $layer=LI1_cond $X=2.547 $Y=0.085
+ $X2=2.547 $Y2=0
r134 20 22 13.9592 $w=3.53e-07 $l=4.3e-07 $layer=LI1_cond $X=2.547 $Y=0.085
+ $X2=2.547 $Y2=0.515
r135 16 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=0.085
+ $X2=0.78 $Y2=0
r136 16 18 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.78 $Y=0.085
+ $X2=0.78 $Y2=0.515
r137 5 34 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.78
+ $Y=0.37 $X2=6.92 $Y2=0.515
r138 4 30 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=5.85
+ $Y=0.37 $X2=5.99 $Y2=0.58
r139 3 26 182 $w=1.7e-07 $l=2.56905e-07 $layer=licon1_NDIFF $count=1 $X=4.77
+ $Y=0.47 $X2=4.99 $Y2=0.55
r140 2 22 182 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_NDIFF $count=1 $X=2.395
+ $Y=0.37 $X2=2.545 $Y2=0.515
r141 1 18 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.78 $Y2=0.515
.ends

