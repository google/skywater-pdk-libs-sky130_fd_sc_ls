* NGSPICE file created from sky130_fd_sc_ls__or3_1.ext - technology: sky130A

.subckt sky130_fd_sc_ls__or3_1 A B C VGND VNB VPB VPWR X
M1000 a_200_368# B a_116_368# VPB phighvt w=1e+06u l=150000u
+  ad=4.2e+11p pd=2.84e+06u as=2.7e+11p ps=2.54e+06u
M1001 VGND A a_27_74# VNB nshort w=550000u l=150000u
+  ad=4.71e+11p pd=4.12e+06u as=5.225e+11p ps=4.1e+06u
M1002 a_27_74# B VGND VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 X a_27_74# VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1004 a_116_368# C a_27_74# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.95e+11p ps=2.59e+06u
M1005 X a_27_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=7.618e+11p ps=3.7e+06u
M1006 VGND C a_27_74# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR A a_200_368# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

