* File: sky130_fd_sc_ls__clkinv_4.pxi.spice
* Created: Wed Sep  2 10:58:57 2020
* 
x_PM_SKY130_FD_SC_LS__CLKINV_4%A N_A_c_63_n N_A_M1000_g N_A_c_55_n N_A_M1001_g
+ N_A_c_65_n N_A_M1002_g N_A_c_66_n N_A_M1003_g N_A_M1004_g N_A_c_67_n
+ N_A_M1005_g N_A_c_68_n N_A_M1006_g N_A_M1007_g N_A_c_69_n N_A_M1008_g
+ N_A_M1009_g N_A_c_60_n A A A A A N_A_c_62_n PM_SKY130_FD_SC_LS__CLKINV_4%A
x_PM_SKY130_FD_SC_LS__CLKINV_4%VPWR N_VPWR_M1000_d N_VPWR_M1002_d N_VPWR_M1005_d
+ N_VPWR_M1008_d N_VPWR_c_164_n N_VPWR_c_165_n N_VPWR_c_166_n N_VPWR_c_167_n
+ N_VPWR_c_168_n N_VPWR_c_169_n N_VPWR_c_170_n N_VPWR_c_171_n VPWR
+ N_VPWR_c_172_n N_VPWR_c_173_n N_VPWR_c_174_n N_VPWR_c_163_n
+ PM_SKY130_FD_SC_LS__CLKINV_4%VPWR
x_PM_SKY130_FD_SC_LS__CLKINV_4%Y N_Y_M1001_d N_Y_M1007_d N_Y_M1000_s N_Y_M1003_s
+ N_Y_M1006_s N_Y_c_216_n N_Y_c_217_n N_Y_c_226_n N_Y_c_240_n N_Y_c_243_n
+ N_Y_c_227_n N_Y_c_218_n N_Y_c_254_n N_Y_c_219_n N_Y_c_228_n N_Y_c_220_n
+ N_Y_c_229_n N_Y_c_221_n N_Y_c_222_n N_Y_c_276_n N_Y_c_223_n N_Y_c_284_n Y
+ PM_SKY130_FD_SC_LS__CLKINV_4%Y
x_PM_SKY130_FD_SC_LS__CLKINV_4%VGND N_VGND_M1001_s N_VGND_M1004_s N_VGND_M1009_s
+ N_VGND_c_324_n N_VGND_c_325_n N_VGND_c_326_n VGND N_VGND_c_327_n
+ N_VGND_c_328_n N_VGND_c_329_n N_VGND_c_330_n N_VGND_c_331_n
+ PM_SKY130_FD_SC_LS__CLKINV_4%VGND
cc_1 VNB N_A_c_55_n 0.0113426f $X=-0.19 $Y=-0.245 $X2=0.865 $Y2=1.605
cc_2 VNB N_A_M1001_g 0.0533591f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=0.61
cc_3 VNB N_A_M1004_g 0.0463332f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=0.61
cc_4 VNB N_A_M1007_g 0.0390581f $X=-0.19 $Y=-0.245 $X2=2.365 $Y2=0.61
cc_5 VNB N_A_M1009_g 0.0454945f $X=-0.19 $Y=-0.245 $X2=2.82 $Y2=0.61
cc_6 VNB N_A_c_60_n 0.0113216f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.605
cc_7 VNB A 0.00410794f $X=-0.19 $Y=-0.245 $X2=2.555 $Y2=1.58
cc_8 VNB N_A_c_62_n 0.101597f $X=-0.19 $Y=-0.245 $X2=2.805 $Y2=1.557
cc_9 VNB N_VPWR_c_163_n 0.143779f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=1.557
cc_10 VNB N_Y_c_216_n 0.0207859f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=0.61
cc_11 VNB N_Y_c_217_n 0.00997995f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_Y_c_218_n 0.00961836f $X=-0.19 $Y=-0.245 $X2=2.805 $Y2=1.765
cc_13 VNB N_Y_c_219_n 0.0047561f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_Y_c_220_n 0.015358f $X=-0.19 $Y=-0.245 $X2=2.075 $Y2=1.58
cc_15 VNB N_Y_c_221_n 0.0110787f $X=-0.19 $Y=-0.245 $X2=1.03 $Y2=1.515
cc_16 VNB N_Y_c_222_n 0.00940303f $X=-0.19 $Y=-0.245 $X2=1.03 $Y2=1.515
cc_17 VNB N_Y_c_223_n 0.00245776f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=1.557
cc_18 VNB Y 0.0243509f $X=-0.19 $Y=-0.245 $X2=2.39 $Y2=1.515
cc_19 VNB N_VGND_c_324_n 0.0138293f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_20 VNB N_VGND_c_325_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=2.4
cc_21 VNB N_VGND_c_326_n 0.0348923f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=1.35
cc_22 VNB N_VGND_c_327_n 0.0299922f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=1.765
cc_23 VNB N_VGND_c_328_n 0.0188284f $X=-0.19 $Y=-0.245 $X2=2.355 $Y2=2.4
cc_24 VNB N_VGND_c_329_n 0.0542217f $X=-0.19 $Y=-0.245 $X2=2.805 $Y2=2.4
cc_25 VNB N_VGND_c_330_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_331_n 0.214061f $X=-0.19 $Y=-0.245 $X2=2.075 $Y2=1.58
cc_27 VPB N_A_c_63_n 0.0168761f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_28 VPB N_A_c_55_n 0.00820074f $X=-0.19 $Y=1.66 $X2=0.865 $Y2=1.605
cc_29 VPB N_A_c_65_n 0.0155086f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.765
cc_30 VPB N_A_c_66_n 0.0155127f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=1.765
cc_31 VPB N_A_c_67_n 0.015892f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=1.765
cc_32 VPB N_A_c_68_n 0.0158874f $X=-0.19 $Y=1.66 $X2=2.355 $Y2=1.765
cc_33 VPB N_A_c_69_n 0.0163319f $X=-0.19 $Y=1.66 $X2=2.805 $Y2=1.765
cc_34 VPB N_A_c_60_n 0.00721598f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.605
cc_35 VPB A 0.0148077f $X=-0.19 $Y=1.66 $X2=2.555 $Y2=1.58
cc_36 VPB N_A_c_62_n 0.0615269f $X=-0.19 $Y=1.66 $X2=2.805 $Y2=1.557
cc_37 VPB N_VPWR_c_164_n 0.0106521f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=1.765
cc_38 VPB N_VPWR_c_165_n 0.0376965f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=2.4
cc_39 VPB N_VPWR_c_166_n 0.00799266f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_40 VPB N_VPWR_c_167_n 0.0082016f $X=-0.19 $Y=1.66 $X2=2.355 $Y2=1.765
cc_41 VPB N_VPWR_c_168_n 0.0121909f $X=-0.19 $Y=1.66 $X2=2.355 $Y2=2.4
cc_42 VPB N_VPWR_c_169_n 0.0384719f $X=-0.19 $Y=1.66 $X2=2.365 $Y2=0.61
cc_43 VPB N_VPWR_c_170_n 0.0206041f $X=-0.19 $Y=1.66 $X2=2.805 $Y2=1.765
cc_44 VPB N_VPWR_c_171_n 0.00324402f $X=-0.19 $Y=1.66 $X2=2.805 $Y2=2.4
cc_45 VPB N_VPWR_c_172_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_173_n 0.0186948f $X=-0.19 $Y=1.66 $X2=2.075 $Y2=1.58
cc_47 VPB N_VPWR_c_174_n 0.0047828f $X=-0.19 $Y=1.66 $X2=1.03 $Y2=1.557
cc_48 VPB N_VPWR_c_163_n 0.0651218f $X=-0.19 $Y=1.66 $X2=1.795 $Y2=1.557
cc_49 VPB N_Y_c_216_n 0.00618364f $X=-0.19 $Y=1.66 $X2=1.795 $Y2=0.61
cc_50 VPB N_Y_c_226_n 0.00257348f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=2.4
cc_51 VPB N_Y_c_227_n 0.00257348f $X=-0.19 $Y=1.66 $X2=2.365 $Y2=0.61
cc_52 VPB N_Y_c_228_n 0.00257348f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_53 VPB N_Y_c_229_n 0.00707089f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB Y 0.0131063f $X=-0.19 $Y=1.66 $X2=2.39 $Y2=1.515
cc_55 N_A_c_63_n N_VPWR_c_165_n 0.00714506f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_56 N_A_c_65_n N_VPWR_c_166_n 0.00486623f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_57 N_A_c_66_n N_VPWR_c_166_n 0.00486623f $X=1.405 $Y=1.765 $X2=0 $Y2=0
cc_58 N_A_c_67_n N_VPWR_c_167_n 0.00534288f $X=1.855 $Y=1.765 $X2=0 $Y2=0
cc_59 N_A_c_68_n N_VPWR_c_167_n 0.00540678f $X=2.355 $Y=1.765 $X2=0 $Y2=0
cc_60 N_A_c_69_n N_VPWR_c_169_n 0.0168809f $X=2.805 $Y=1.765 $X2=0 $Y2=0
cc_61 N_A_c_63_n N_VPWR_c_170_n 0.00445602f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_62 N_A_c_65_n N_VPWR_c_170_n 0.00445602f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_63 N_A_c_66_n N_VPWR_c_172_n 0.00445602f $X=1.405 $Y=1.765 $X2=0 $Y2=0
cc_64 N_A_c_67_n N_VPWR_c_172_n 0.00445602f $X=1.855 $Y=1.765 $X2=0 $Y2=0
cc_65 N_A_c_68_n N_VPWR_c_173_n 0.00445602f $X=2.355 $Y=1.765 $X2=0 $Y2=0
cc_66 N_A_c_69_n N_VPWR_c_173_n 0.00445602f $X=2.805 $Y=1.765 $X2=0 $Y2=0
cc_67 N_A_c_63_n N_VPWR_c_163_n 0.00861084f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_68 N_A_c_65_n N_VPWR_c_163_n 0.00857589f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_69 N_A_c_66_n N_VPWR_c_163_n 0.00857589f $X=1.405 $Y=1.765 $X2=0 $Y2=0
cc_70 N_A_c_67_n N_VPWR_c_163_n 0.0085805f $X=1.855 $Y=1.765 $X2=0 $Y2=0
cc_71 N_A_c_68_n N_VPWR_c_163_n 0.00857378f $X=2.355 $Y=1.765 $X2=0 $Y2=0
cc_72 N_A_c_69_n N_VPWR_c_163_n 0.00860566f $X=2.805 $Y=1.765 $X2=0 $Y2=0
cc_73 N_A_c_63_n N_Y_c_216_n 0.0060862f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_74 N_A_M1001_g N_Y_c_216_n 0.00442873f $X=0.94 $Y=0.61 $X2=0 $Y2=0
cc_75 N_A_c_65_n N_Y_c_216_n 5.77508e-19 $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_76 N_A_c_60_n N_Y_c_216_n 0.00789937f $X=0.505 $Y=1.605 $X2=0 $Y2=0
cc_77 A N_Y_c_216_n 0.0344967f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_78 N_A_c_62_n N_Y_c_216_n 7.51683e-19 $X=2.805 $Y=1.557 $X2=0 $Y2=0
cc_79 N_A_c_63_n N_Y_c_226_n 0.0152303f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_80 N_A_c_65_n N_Y_c_226_n 0.0105292f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_81 N_A_c_66_n N_Y_c_226_n 6.46364e-19 $X=1.405 $Y=1.765 $X2=0 $Y2=0
cc_82 N_A_c_65_n N_Y_c_240_n 0.0120074f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_83 N_A_c_66_n N_Y_c_240_n 0.0120074f $X=1.405 $Y=1.765 $X2=0 $Y2=0
cc_84 N_A_c_62_n N_Y_c_240_n 0.00131635f $X=2.805 $Y=1.557 $X2=0 $Y2=0
cc_85 N_A_c_63_n N_Y_c_243_n 0.0171718f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_86 N_A_c_55_n N_Y_c_243_n 0.0012993f $X=0.865 $Y=1.605 $X2=0 $Y2=0
cc_87 N_A_c_65_n N_Y_c_243_n 4.54092e-19 $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_88 A N_Y_c_243_n 0.0591198f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_89 N_A_c_65_n N_Y_c_227_n 6.45594e-19 $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_90 N_A_c_66_n N_Y_c_227_n 0.0104707f $X=1.405 $Y=1.765 $X2=0 $Y2=0
cc_91 N_A_c_67_n N_Y_c_227_n 0.0107096f $X=1.855 $Y=1.765 $X2=0 $Y2=0
cc_92 N_A_c_68_n N_Y_c_227_n 6.99794e-19 $X=2.355 $Y=1.765 $X2=0 $Y2=0
cc_93 N_A_M1004_g N_Y_c_218_n 0.0118691f $X=1.795 $Y=0.61 $X2=0 $Y2=0
cc_94 N_A_M1007_g N_Y_c_218_n 0.0118691f $X=2.365 $Y=0.61 $X2=0 $Y2=0
cc_95 N_A_c_62_n N_Y_c_218_n 0.00538093f $X=2.805 $Y=1.557 $X2=0 $Y2=0
cc_96 N_A_c_67_n N_Y_c_254_n 0.0122806f $X=1.855 $Y=1.765 $X2=0 $Y2=0
cc_97 N_A_c_68_n N_Y_c_254_n 0.0122806f $X=2.355 $Y=1.765 $X2=0 $Y2=0
cc_98 A N_Y_c_254_n 0.04337f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_99 N_A_c_62_n N_Y_c_254_n 0.00158759f $X=2.805 $Y=1.557 $X2=0 $Y2=0
cc_100 N_A_M1004_g N_Y_c_219_n 6.22763e-19 $X=1.795 $Y=0.61 $X2=0 $Y2=0
cc_101 N_A_M1007_g N_Y_c_219_n 0.0110981f $X=2.365 $Y=0.61 $X2=0 $Y2=0
cc_102 N_A_M1009_g N_Y_c_219_n 0.00547196f $X=2.82 $Y=0.61 $X2=0 $Y2=0
cc_103 N_A_c_67_n N_Y_c_228_n 6.04643e-19 $X=1.855 $Y=1.765 $X2=0 $Y2=0
cc_104 N_A_c_68_n N_Y_c_228_n 0.0102215f $X=2.355 $Y=1.765 $X2=0 $Y2=0
cc_105 N_A_c_69_n N_Y_c_228_n 0.0145698f $X=2.805 $Y=1.765 $X2=0 $Y2=0
cc_106 N_A_M1009_g N_Y_c_220_n 0.018715f $X=2.82 $Y=0.61 $X2=0 $Y2=0
cc_107 A N_Y_c_220_n 6.95742e-19 $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_108 N_A_c_69_n N_Y_c_229_n 0.0172133f $X=2.805 $Y=1.765 $X2=0 $Y2=0
cc_109 A N_Y_c_229_n 6.95742e-19 $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_110 N_A_c_55_n N_Y_c_221_n 0.0012067f $X=0.865 $Y=1.605 $X2=0 $Y2=0
cc_111 N_A_M1001_g N_Y_c_221_n 0.0130527f $X=0.94 $Y=0.61 $X2=0 $Y2=0
cc_112 N_A_c_60_n N_Y_c_221_n 0.00567085f $X=0.505 $Y=1.605 $X2=0 $Y2=0
cc_113 A N_Y_c_221_n 0.144874f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_114 N_A_M1001_g N_Y_c_222_n 0.0256826f $X=0.94 $Y=0.61 $X2=0 $Y2=0
cc_115 N_A_M1004_g N_Y_c_222_n 0.0162981f $X=1.795 $Y=0.61 $X2=0 $Y2=0
cc_116 N_A_M1007_g N_Y_c_222_n 6.05295e-19 $X=2.365 $Y=0.61 $X2=0 $Y2=0
cc_117 N_A_c_62_n N_Y_c_222_n 0.0128478f $X=2.805 $Y=1.557 $X2=0 $Y2=0
cc_118 N_A_c_66_n N_Y_c_276_n 4.27055e-19 $X=1.405 $Y=1.765 $X2=0 $Y2=0
cc_119 N_A_c_67_n N_Y_c_276_n 4.27055e-19 $X=1.855 $Y=1.765 $X2=0 $Y2=0
cc_120 A N_Y_c_276_n 0.0237598f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_121 N_A_c_62_n N_Y_c_276_n 0.00144409f $X=2.805 $Y=1.557 $X2=0 $Y2=0
cc_122 N_A_M1007_g N_Y_c_223_n 0.00294386f $X=2.365 $Y=0.61 $X2=0 $Y2=0
cc_123 N_A_M1009_g N_Y_c_223_n 0.00218126f $X=2.82 $Y=0.61 $X2=0 $Y2=0
cc_124 A N_Y_c_223_n 0.028235f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_125 N_A_c_62_n N_Y_c_223_n 0.00291196f $X=2.805 $Y=1.557 $X2=0 $Y2=0
cc_126 N_A_c_68_n N_Y_c_284_n 4.27055e-19 $X=2.355 $Y=1.765 $X2=0 $Y2=0
cc_127 N_A_c_69_n N_Y_c_284_n 4.27055e-19 $X=2.805 $Y=1.765 $X2=0 $Y2=0
cc_128 A N_Y_c_284_n 0.0237598f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_129 N_A_c_62_n N_Y_c_284_n 0.00144338f $X=2.805 $Y=1.557 $X2=0 $Y2=0
cc_130 N_A_c_69_n Y 0.00663402f $X=2.805 $Y=1.765 $X2=0 $Y2=0
cc_131 N_A_M1009_g Y 0.0180849f $X=2.82 $Y=0.61 $X2=0 $Y2=0
cc_132 A Y 0.0261104f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_133 N_A_M1004_g N_VGND_c_324_n 0.00651086f $X=1.795 $Y=0.61 $X2=0 $Y2=0
cc_134 N_A_M1007_g N_VGND_c_324_n 0.00473938f $X=2.365 $Y=0.61 $X2=0 $Y2=0
cc_135 N_A_M1009_g N_VGND_c_326_n 0.00492488f $X=2.82 $Y=0.61 $X2=0 $Y2=0
cc_136 N_A_M1001_g N_VGND_c_327_n 0.0053111f $X=0.94 $Y=0.61 $X2=0 $Y2=0
cc_137 N_A_M1004_g N_VGND_c_327_n 0.0053111f $X=1.795 $Y=0.61 $X2=0 $Y2=0
cc_138 N_A_M1007_g N_VGND_c_328_n 0.00530655f $X=2.365 $Y=0.61 $X2=0 $Y2=0
cc_139 N_A_M1009_g N_VGND_c_328_n 0.0055601f $X=2.82 $Y=0.61 $X2=0 $Y2=0
cc_140 N_A_M1001_g N_VGND_c_329_n 0.012091f $X=0.94 $Y=0.61 $X2=0 $Y2=0
cc_141 N_A_M1001_g N_VGND_c_331_n 0.00536257f $X=0.94 $Y=0.61 $X2=0 $Y2=0
cc_142 N_A_M1004_g N_VGND_c_331_n 0.00536257f $X=1.795 $Y=0.61 $X2=0 $Y2=0
cc_143 N_A_M1007_g N_VGND_c_331_n 0.00536257f $X=2.365 $Y=0.61 $X2=0 $Y2=0
cc_144 N_A_M1009_g N_VGND_c_331_n 0.00536257f $X=2.82 $Y=0.61 $X2=0 $Y2=0
cc_145 N_VPWR_M1000_d N_Y_c_216_n 0.0045135f $X=0.135 $Y=1.84 $X2=0 $Y2=0
cc_146 N_VPWR_c_165_n N_Y_c_226_n 0.0462948f $X=0.28 $Y=2.455 $X2=0 $Y2=0
cc_147 N_VPWR_c_166_n N_Y_c_226_n 0.0449718f $X=1.18 $Y=2.455 $X2=0 $Y2=0
cc_148 N_VPWR_c_170_n N_Y_c_226_n 0.014552f $X=1.095 $Y=3.33 $X2=0 $Y2=0
cc_149 N_VPWR_c_163_n N_Y_c_226_n 0.0119791f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_150 N_VPWR_M1002_d N_Y_c_240_n 0.00408911f $X=1.03 $Y=1.84 $X2=0 $Y2=0
cc_151 N_VPWR_c_166_n N_Y_c_240_n 0.0136682f $X=1.18 $Y=2.455 $X2=0 $Y2=0
cc_152 N_VPWR_M1000_d N_Y_c_243_n 0.00928011f $X=0.135 $Y=1.84 $X2=0 $Y2=0
cc_153 N_VPWR_c_165_n N_Y_c_243_n 0.00801802f $X=0.28 $Y=2.455 $X2=0 $Y2=0
cc_154 N_VPWR_c_166_n N_Y_c_227_n 0.0449718f $X=1.18 $Y=2.455 $X2=0 $Y2=0
cc_155 N_VPWR_c_167_n N_Y_c_227_n 0.0462948f $X=2.08 $Y=2.455 $X2=0 $Y2=0
cc_156 N_VPWR_c_172_n N_Y_c_227_n 0.014552f $X=1.995 $Y=3.33 $X2=0 $Y2=0
cc_157 N_VPWR_c_163_n N_Y_c_227_n 0.0119791f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_158 N_VPWR_M1005_d N_Y_c_254_n 0.00480741f $X=1.93 $Y=1.84 $X2=0 $Y2=0
cc_159 N_VPWR_c_167_n N_Y_c_254_n 0.0184684f $X=2.08 $Y=2.455 $X2=0 $Y2=0
cc_160 N_VPWR_c_167_n N_Y_c_228_n 0.0266484f $X=2.08 $Y=2.455 $X2=0 $Y2=0
cc_161 N_VPWR_c_169_n N_Y_c_228_n 0.0266809f $X=3.08 $Y=2.455 $X2=0 $Y2=0
cc_162 N_VPWR_c_173_n N_Y_c_228_n 0.014552f $X=2.915 $Y=3.33 $X2=0 $Y2=0
cc_163 N_VPWR_c_163_n N_Y_c_228_n 0.0119791f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_164 N_VPWR_M1008_d N_Y_c_229_n 0.00724473f $X=2.88 $Y=1.84 $X2=0 $Y2=0
cc_165 N_VPWR_c_169_n N_Y_c_229_n 0.0261765f $X=3.08 $Y=2.455 $X2=0 $Y2=0
cc_166 N_VPWR_M1008_d Y 0.00227207f $X=2.88 $Y=1.84 $X2=0 $Y2=0
cc_167 N_Y_c_218_n N_VGND_c_324_n 0.0277029f $X=2.415 $Y=1.095 $X2=0 $Y2=0
cc_168 N_Y_c_219_n N_VGND_c_324_n 0.0188413f $X=2.58 $Y=0.61 $X2=0 $Y2=0
cc_169 N_Y_c_222_n N_VGND_c_324_n 0.0169695f $X=1.745 $Y=0.817 $X2=0 $Y2=0
cc_170 N_Y_c_219_n N_VGND_c_326_n 0.0193875f $X=2.58 $Y=0.61 $X2=0 $Y2=0
cc_171 N_Y_c_220_n N_VGND_c_326_n 0.0290296f $X=3.005 $Y=1.095 $X2=0 $Y2=0
cc_172 N_Y_c_222_n N_VGND_c_327_n 0.0210518f $X=1.745 $Y=0.817 $X2=0 $Y2=0
cc_173 N_Y_c_219_n N_VGND_c_328_n 0.012991f $X=2.58 $Y=0.61 $X2=0 $Y2=0
cc_174 N_Y_c_217_n N_VGND_c_329_n 0.0103794f $X=0.435 $Y=1.095 $X2=0 $Y2=0
cc_175 N_Y_c_221_n N_VGND_c_329_n 0.0207787f $X=0.99 $Y=0.817 $X2=0 $Y2=0
cc_176 N_Y_c_219_n N_VGND_c_331_n 0.0118717f $X=2.58 $Y=0.61 $X2=0 $Y2=0
cc_177 N_Y_c_222_n N_VGND_c_331_n 0.0259639f $X=1.745 $Y=0.817 $X2=0 $Y2=0
