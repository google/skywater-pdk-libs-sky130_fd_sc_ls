* File: sky130_fd_sc_ls__buf_16.spice
* Created: Wed Sep  2 10:56:24 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__buf_16.pex.spice"
.subckt sky130_fd_sc_ls__buf_16  VNB VPB A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1000 N_X_M1000_d N_A_83_260#_M1000_g N_VGND_M1000_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75009.8 A=0.111 P=1.78 MULT=1
MM1004 N_X_M1000_d N_A_83_260#_M1004_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75009.3 A=0.111 P=1.78 MULT=1
MM1008 N_X_M1008_d N_A_83_260#_M1008_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75008.9 A=0.111 P=1.78 MULT=1
MM1010 N_X_M1008_d N_A_83_260#_M1010_g N_VGND_M1010_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75008.5 A=0.111 P=1.78 MULT=1
MM1012 N_X_M1012_d N_A_83_260#_M1012_g N_VGND_M1010_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.9
+ SB=75008 A=0.111 P=1.78 MULT=1
MM1020 N_X_M1012_d N_A_83_260#_M1020_g N_VGND_M1020_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.4
+ SB=75007.6 A=0.111 P=1.78 MULT=1
MM1021 N_X_M1021_d N_A_83_260#_M1021_g N_VGND_M1020_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.8
+ SB=75007.2 A=0.111 P=1.78 MULT=1
MM1024 N_X_M1021_d N_A_83_260#_M1024_g N_VGND_M1024_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75003.2
+ SB=75006.8 A=0.111 P=1.78 MULT=1
MM1025 N_X_M1025_d N_A_83_260#_M1025_g N_VGND_M1024_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75003.6
+ SB=75006.3 A=0.111 P=1.78 MULT=1
MM1026 N_X_M1025_d N_A_83_260#_M1026_g N_VGND_M1026_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1554 PD=1.02 PS=1.16 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75004.1
+ SB=75005.9 A=0.111 P=1.78 MULT=1
MM1032 N_X_M1032_d N_A_83_260#_M1032_g N_VGND_M1026_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1554 PD=1.02 PS=1.16 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75004.6
+ SB=75005.3 A=0.111 P=1.78 MULT=1
MM1033 N_X_M1032_d N_A_83_260#_M1033_g N_VGND_M1033_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1554 PD=1.02 PS=1.16 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75005.1
+ SB=75004.9 A=0.111 P=1.78 MULT=1
MM1036 N_X_M1036_d N_A_83_260#_M1036_g N_VGND_M1033_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1554 PD=1.02 PS=1.16 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75005.6
+ SB=75004.3 A=0.111 P=1.78 MULT=1
MM1037 N_X_M1036_d N_A_83_260#_M1037_g N_VGND_M1037_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1554 PD=1.02 PS=1.16 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75006.1
+ SB=75003.9 A=0.111 P=1.78 MULT=1
MM1038 N_X_M1038_d N_A_83_260#_M1038_g N_VGND_M1037_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1554 PD=1.02 PS=1.16 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75006.6
+ SB=75003.3 A=0.111 P=1.78 MULT=1
MM1039 N_X_M1038_d N_A_83_260#_M1039_g N_VGND_M1039_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75007.1
+ SB=75002.9 A=0.111 P=1.78 MULT=1
MM1005 N_VGND_M1039_s N_A_M1005_g N_A_83_260#_M1005_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75007.5
+ SB=75002.5 A=0.111 P=1.78 MULT=1
MM1011 N_VGND_M1011_d N_A_M1011_g N_A_83_260#_M1005_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75007.9
+ SB=75002 A=0.111 P=1.78 MULT=1
MM1016 N_VGND_M1011_d N_A_M1016_g N_A_83_260#_M1016_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75008.4
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1017 N_VGND_M1017_d N_A_M1017_g N_A_83_260#_M1016_s VNB NSHORT L=0.15 W=0.74
+ AD=0.11655 AS=0.1036 PD=1.055 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75008.8
+ SB=75001.2 A=0.111 P=1.78 MULT=1
MM1040 N_VGND_M1017_d N_A_M1040_g N_A_83_260#_M1040_s VNB NSHORT L=0.15 W=0.74
+ AD=0.11655 AS=0.1295 PD=1.055 PS=1.09 NRD=5.664 NRS=0 M=1 R=4.93333 SA=75009.3
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1043 N_VGND_M1043_d N_A_M1043_g N_A_83_260#_M1040_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.1295 PD=2.05 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75009.8
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1001 N_VPWR_M1001_d N_A_83_260#_M1001_g N_X_M1001_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75009.8 A=0.168 P=2.54 MULT=1
MM1006 N_VPWR_M1006_d N_A_83_260#_M1006_g N_X_M1001_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75009.3 A=0.168 P=2.54 MULT=1
MM1007 N_VPWR_M1006_d N_A_83_260#_M1007_g N_X_M1007_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75008.9 A=0.168 P=2.54 MULT=1
MM1009 N_VPWR_M1009_d N_A_83_260#_M1009_g N_X_M1007_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.196 AS=0.168 PD=1.47 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75001.6 SB=75008.4 A=0.168 P=2.54 MULT=1
MM1013 N_VPWR_M1009_d N_A_83_260#_M1013_g N_X_M1013_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.196 AS=0.168 PD=1.47 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.1 SB=75007.9 A=0.168 P=2.54 MULT=1
MM1014 N_VPWR_M1014_d N_A_83_260#_M1014_g N_X_M1013_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.5 SB=75007.5 A=0.168 P=2.54 MULT=1
MM1018 N_VPWR_M1014_d N_A_83_260#_M1018_g N_X_M1018_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75003
+ SB=75007 A=0.168 P=2.54 MULT=1
MM1022 N_VPWR_M1022_d N_A_83_260#_M1022_g N_X_M1018_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75003.4 SB=75006.6 A=0.168 P=2.54 MULT=1
MM1023 N_VPWR_M1022_d N_A_83_260#_M1023_g N_X_M1023_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75003.9 SB=75006.1 A=0.168 P=2.54 MULT=1
MM1027 N_VPWR_M1027_d N_A_83_260#_M1027_g N_X_M1023_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75004.3 SB=75005.7 A=0.168 P=2.54 MULT=1
MM1028 N_VPWR_M1027_d N_A_83_260#_M1028_g N_X_M1028_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75004.8 SB=75005.2 A=0.168 P=2.54 MULT=1
MM1030 N_VPWR_M1030_d N_A_83_260#_M1030_g N_X_M1028_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75005.2 SB=75004.8 A=0.168 P=2.54 MULT=1
MM1031 N_VPWR_M1030_d N_A_83_260#_M1031_g N_X_M1031_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75005.7 SB=75004.3 A=0.168 P=2.54 MULT=1
MM1034 N_VPWR_M1034_d N_A_83_260#_M1034_g N_X_M1031_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75006.1 SB=75003.9 A=0.168 P=2.54 MULT=1
MM1041 N_VPWR_M1034_d N_A_83_260#_M1041_g N_X_M1041_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75006.6 SB=75003.4 A=0.168 P=2.54 MULT=1
MM1042 N_VPWR_M1042_d N_A_83_260#_M1042_g N_X_M1041_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.196 AS=0.168 PD=1.47 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75007
+ SB=75003 A=0.168 P=2.54 MULT=1
MM1002 N_VPWR_M1042_d N_A_M1002_g N_A_83_260#_M1002_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.196 AS=0.168 PD=1.47 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75007.5 SB=75002.5 A=0.168 P=2.54 MULT=1
MM1003 N_VPWR_M1003_d N_A_M1003_g N_A_83_260#_M1002_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75008
+ SB=75002 A=0.168 P=2.54 MULT=1
MM1015 N_VPWR_M1003_d N_A_M1015_g N_A_83_260#_M1015_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75008.4 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1019 N_VPWR_M1019_d N_A_M1019_g N_A_83_260#_M1015_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75008.9 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1029 N_VPWR_M1019_d N_A_M1029_g N_A_83_260#_M1029_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75009.3 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1035 N_VPWR_M1035_d N_A_M1035_g N_A_83_260#_M1029_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75009.8 SB=75000.2 A=0.168 P=2.54 MULT=1
DX44_noxref VNB VPB NWDIODE A=20.3484 P=25.6
c_97 VNB 0 3.07957e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_ls__buf_16.pxi.spice"
*
.ends
*
*
