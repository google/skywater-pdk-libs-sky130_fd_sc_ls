# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ls__sedfxtp_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ls__sedfxtp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  16.32000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 0.980000 0.805000 1.990000 ;
    END
  END D
  PIN DE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.515000 1.320000 1.845000 1.780000 ;
    END
  END DE
  PIN Q
    ANTENNADIFFAREA  0.560000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 15.375000 0.350000 15.705000 1.130000 ;
        RECT 15.460000 1.130000 15.705000 1.550000 ;
        RECT 15.460000 1.550000 16.195000 2.150000 ;
        RECT 15.460000 2.150000 15.705000 2.980000 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.955000 1.180000 5.410000 1.745000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.465000 1.180000 4.785000 1.510000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 6.395000 1.180000 6.725000 1.550000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 16.320000 0.085000 ;
        RECT  1.055000  0.085000  1.385000 0.810000 ;
        RECT  2.045000  0.085000  2.375000 1.005000 ;
        RECT  4.885000  0.085000  5.215000 1.010000 ;
        RECT  6.235000  0.085000  6.495000 0.680000 ;
        RECT  7.235000  0.085000  7.485000 1.130000 ;
        RECT 10.100000  0.085000 10.365000 0.680000 ;
        RECT 11.635000  0.085000 11.885000 0.680000 ;
        RECT 13.210000  0.085000 14.145000 0.680000 ;
        RECT 14.875000  0.085000 15.205000 0.950000 ;
        RECT 15.875000  0.085000 16.205000 1.130000 ;
      LAYER mcon ;
        RECT  0.155000 -0.085000  0.325000 0.085000 ;
        RECT  0.635000 -0.085000  0.805000 0.085000 ;
        RECT  1.115000 -0.085000  1.285000 0.085000 ;
        RECT  1.595000 -0.085000  1.765000 0.085000 ;
        RECT  2.075000 -0.085000  2.245000 0.085000 ;
        RECT  2.555000 -0.085000  2.725000 0.085000 ;
        RECT  3.035000 -0.085000  3.205000 0.085000 ;
        RECT  3.515000 -0.085000  3.685000 0.085000 ;
        RECT  3.995000 -0.085000  4.165000 0.085000 ;
        RECT  4.475000 -0.085000  4.645000 0.085000 ;
        RECT  4.955000 -0.085000  5.125000 0.085000 ;
        RECT  5.435000 -0.085000  5.605000 0.085000 ;
        RECT  5.915000 -0.085000  6.085000 0.085000 ;
        RECT  6.395000 -0.085000  6.565000 0.085000 ;
        RECT  6.875000 -0.085000  7.045000 0.085000 ;
        RECT  7.355000 -0.085000  7.525000 0.085000 ;
        RECT  7.835000 -0.085000  8.005000 0.085000 ;
        RECT  8.315000 -0.085000  8.485000 0.085000 ;
        RECT  8.795000 -0.085000  8.965000 0.085000 ;
        RECT  9.275000 -0.085000  9.445000 0.085000 ;
        RECT  9.755000 -0.085000  9.925000 0.085000 ;
        RECT 10.235000 -0.085000 10.405000 0.085000 ;
        RECT 10.715000 -0.085000 10.885000 0.085000 ;
        RECT 11.195000 -0.085000 11.365000 0.085000 ;
        RECT 11.675000 -0.085000 11.845000 0.085000 ;
        RECT 12.155000 -0.085000 12.325000 0.085000 ;
        RECT 12.635000 -0.085000 12.805000 0.085000 ;
        RECT 13.115000 -0.085000 13.285000 0.085000 ;
        RECT 13.595000 -0.085000 13.765000 0.085000 ;
        RECT 14.075000 -0.085000 14.245000 0.085000 ;
        RECT 14.555000 -0.085000 14.725000 0.085000 ;
        RECT 15.035000 -0.085000 15.205000 0.085000 ;
        RECT 15.515000 -0.085000 15.685000 0.085000 ;
        RECT 15.995000 -0.085000 16.165000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 16.320000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 3.245000 16.320000 3.415000 ;
        RECT  1.050000 2.630000  1.300000 3.245000 ;
        RECT  2.490000 2.630000  2.740000 3.245000 ;
        RECT  5.010000 2.595000  5.260000 3.245000 ;
        RECT  6.360000 2.710000  6.695000 3.245000 ;
        RECT  7.755000 2.710000  8.085000 3.245000 ;
        RECT 10.215000 2.730000 10.545000 3.245000 ;
        RECT 11.310000 2.730000 11.650000 3.245000 ;
        RECT 13.690000 2.650000 14.230000 3.245000 ;
        RECT 14.960000 1.950000 15.290000 3.245000 ;
        RECT 15.875000 2.320000 16.205000 3.245000 ;
      LAYER mcon ;
        RECT  0.155000 3.245000  0.325000 3.415000 ;
        RECT  0.635000 3.245000  0.805000 3.415000 ;
        RECT  1.115000 3.245000  1.285000 3.415000 ;
        RECT  1.595000 3.245000  1.765000 3.415000 ;
        RECT  2.075000 3.245000  2.245000 3.415000 ;
        RECT  2.555000 3.245000  2.725000 3.415000 ;
        RECT  3.035000 3.245000  3.205000 3.415000 ;
        RECT  3.515000 3.245000  3.685000 3.415000 ;
        RECT  3.995000 3.245000  4.165000 3.415000 ;
        RECT  4.475000 3.245000  4.645000 3.415000 ;
        RECT  4.955000 3.245000  5.125000 3.415000 ;
        RECT  5.435000 3.245000  5.605000 3.415000 ;
        RECT  5.915000 3.245000  6.085000 3.415000 ;
        RECT  6.395000 3.245000  6.565000 3.415000 ;
        RECT  6.875000 3.245000  7.045000 3.415000 ;
        RECT  7.355000 3.245000  7.525000 3.415000 ;
        RECT  7.835000 3.245000  8.005000 3.415000 ;
        RECT  8.315000 3.245000  8.485000 3.415000 ;
        RECT  8.795000 3.245000  8.965000 3.415000 ;
        RECT  9.275000 3.245000  9.445000 3.415000 ;
        RECT  9.755000 3.245000  9.925000 3.415000 ;
        RECT 10.235000 3.245000 10.405000 3.415000 ;
        RECT 10.715000 3.245000 10.885000 3.415000 ;
        RECT 11.195000 3.245000 11.365000 3.415000 ;
        RECT 11.675000 3.245000 11.845000 3.415000 ;
        RECT 12.155000 3.245000 12.325000 3.415000 ;
        RECT 12.635000 3.245000 12.805000 3.415000 ;
        RECT 13.115000 3.245000 13.285000 3.415000 ;
        RECT 13.595000 3.245000 13.765000 3.415000 ;
        RECT 14.075000 3.245000 14.245000 3.415000 ;
        RECT 14.555000 3.245000 14.725000 3.415000 ;
        RECT 15.035000 3.245000 15.205000 3.415000 ;
        RECT 15.515000 3.245000 15.685000 3.415000 ;
        RECT 15.995000 3.245000 16.165000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 16.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.085000 0.350000  0.565000 0.810000 ;
      RECT  0.085000 0.810000  0.255000 2.290000 ;
      RECT  0.085000 2.290000  1.640000 2.460000 ;
      RECT  0.085000 2.460000  0.510000 2.980000 ;
      RECT  0.975000 0.980000  1.865000 1.150000 ;
      RECT  0.975000 1.150000  1.305000 1.950000 ;
      RECT  0.975000 1.950000  2.385000 2.120000 ;
      RECT  1.470000 2.460000  1.640000 2.905000 ;
      RECT  1.470000 2.905000  2.320000 3.075000 ;
      RECT  1.615000 0.545000  1.865000 0.980000 ;
      RECT  1.810000 2.120000  1.980000 2.735000 ;
      RECT  2.055000 1.520000  2.385000 1.950000 ;
      RECT  2.150000 2.290000  3.500000 2.460000 ;
      RECT  2.150000 2.460000  2.320000 2.905000 ;
      RECT  2.555000 1.515000  3.070000 1.845000 ;
      RECT  2.865000 0.675000  3.340000 1.005000 ;
      RECT  3.170000 1.005000  3.340000 1.175000 ;
      RECT  3.170000 1.175000  3.500000 1.345000 ;
      RECT  3.250000 2.460000  3.500000 2.975000 ;
      RECT  3.330000 1.345000  3.500000 2.290000 ;
      RECT  3.510000 0.545000  3.840000 1.005000 ;
      RECT  3.670000 1.005000  3.840000 2.295000 ;
      RECT  3.670000 2.295000  3.950000 2.905000 ;
      RECT  3.670000 2.905000  4.840000 3.075000 ;
      RECT  4.010000 0.255000  4.295000 0.605000 ;
      RECT  4.010000 0.605000  4.715000 1.010000 ;
      RECT  4.010000 1.010000  4.295000 1.915000 ;
      RECT  4.010000 1.915000  5.885000 2.085000 ;
      RECT  4.125000 2.085000  4.295000 2.255000 ;
      RECT  4.125000 2.255000  4.500000 2.735000 ;
      RECT  4.670000 2.255000  6.225000 2.370000 ;
      RECT  4.670000 2.370000  8.425000 2.425000 ;
      RECT  4.670000 2.425000  4.840000 2.905000 ;
      RECT  5.620000 1.415000  5.885000 1.915000 ;
      RECT  5.675000 0.605000  6.005000 0.895000 ;
      RECT  5.675000 0.895000  6.225000 1.065000 ;
      RECT  5.800000 2.425000  8.425000 2.520000 ;
      RECT  5.800000 2.520000  9.015000 2.540000 ;
      RECT  5.800000 2.540000  6.130000 2.935000 ;
      RECT  6.055000 1.065000  6.225000 2.255000 ;
      RECT  6.675000 0.350000  7.065000 1.010000 ;
      RECT  6.895000 1.010000  7.065000 1.530000 ;
      RECT  6.895000 1.530000  7.615000 2.200000 ;
      RECT  7.665000 0.255000  9.495000 0.425000 ;
      RECT  7.665000 0.425000  7.995000 1.130000 ;
      RECT  7.865000 1.480000  8.475000 1.650000 ;
      RECT  7.865000 1.650000  8.035000 2.370000 ;
      RECT  8.205000 1.820000  8.815000 2.020000 ;
      RECT  8.205000 2.020000  9.005000 2.200000 ;
      RECT  8.225000 0.595000  8.475000 1.480000 ;
      RECT  8.255000 2.540000  9.015000 2.690000 ;
      RECT  8.645000 0.425000  8.815000 1.820000 ;
      RECT  8.645000 2.200000  9.005000 2.350000 ;
      RECT  8.765000 2.690000  9.015000 2.980000 ;
      RECT  8.985000 0.595000  9.155000 1.660000 ;
      RECT  8.985000 1.660000 10.785000 1.830000 ;
      RECT  9.185000 1.830000  9.355000 2.520000 ;
      RECT  9.185000 2.520000  9.545000 2.980000 ;
      RECT  9.325000 0.425000  9.495000 0.850000 ;
      RECT  9.325000 0.850000 10.705000 1.020000 ;
      RECT  9.325000 1.020000  9.655000 1.345000 ;
      RECT  9.525000 2.020000  9.885000 2.350000 ;
      RECT  9.715000 2.350000  9.885000 2.390000 ;
      RECT  9.715000 2.390000 12.730000 2.560000 ;
      RECT  9.915000 1.190000 11.800000 1.360000 ;
      RECT  9.915000 1.360000 10.245000 1.490000 ;
      RECT 10.455000 1.530000 10.785000 1.660000 ;
      RECT 10.535000 0.255000 11.465000 0.425000 ;
      RECT 10.535000 0.425000 10.705000 0.850000 ;
      RECT 10.750000 2.050000 11.125000 2.220000 ;
      RECT 10.875000 0.595000 11.125000 1.190000 ;
      RECT 10.955000 1.360000 11.800000 1.520000 ;
      RECT 10.955000 1.520000 11.125000 2.050000 ;
      RECT 11.295000 0.425000 11.465000 0.850000 ;
      RECT 11.295000 0.850000 12.210000 1.020000 ;
      RECT 12.040000 1.020000 12.210000 1.190000 ;
      RECT 12.040000 1.190000 13.450000 1.360000 ;
      RECT 12.040000 1.360000 12.370000 1.800000 ;
      RECT 12.390000 0.350000 12.720000 0.850000 ;
      RECT 12.390000 0.850000 13.790000 1.020000 ;
      RECT 12.560000 1.530000 12.910000 1.755000 ;
      RECT 12.560000 1.755000 12.730000 2.390000 ;
      RECT 12.900000 1.925000 13.250000 2.980000 ;
      RECT 13.080000 1.755000 14.410000 1.925000 ;
      RECT 13.120000 1.360000 13.450000 1.585000 ;
      RECT 13.510000 2.095000 13.840000 2.300000 ;
      RECT 13.510000 2.300000 14.750000 2.470000 ;
      RECT 13.620000 1.020000 13.790000 1.755000 ;
      RECT 14.080000 1.460000 14.410000 1.755000 ;
      RECT 14.080000 1.925000 14.410000 2.130000 ;
      RECT 14.315000 0.350000 14.645000 1.120000 ;
      RECT 14.315000 1.120000 14.750000 1.290000 ;
      RECT 14.400000 2.470000 14.750000 2.980000 ;
      RECT 14.580000 1.290000 14.750000 1.550000 ;
      RECT 14.580000 1.550000 15.235000 1.780000 ;
      RECT 14.580000 1.780000 14.750000 2.300000 ;
    LAYER mcon ;
      RECT  2.555000 1.580000  2.725000 1.750000 ;
      RECT 15.035000 1.580000 15.205000 1.750000 ;
    LAYER met1 ;
      RECT  2.495000 1.550000  2.785000 1.595000 ;
      RECT  2.495000 1.595000 15.265000 1.735000 ;
      RECT  2.495000 1.735000  2.785000 1.780000 ;
      RECT 14.975000 1.550000 15.265000 1.595000 ;
      RECT 14.975000 1.735000 15.265000 1.780000 ;
  END
END sky130_fd_sc_ls__sedfxtp_2
