* NGSPICE file created from sky130_fd_sc_ls__sdfsbp_1.ext - technology: sky130A

.subckt sky130_fd_sc_ls__sdfsbp_1 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q Q_N
M1000 a_1876_74# a_594_74# a_1762_74# VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=2.391e+11p ps=2.12e+06u
M1001 a_1954_74# a_1924_48# a_1876_74# VNB nshort w=420000u l=150000u
+  ad=1.638e+11p pd=1.62e+06u as=0p ps=0u
M1002 VGND a_1163_48# a_1115_74# VNB nshort w=420000u l=150000u
+  ad=2.17215e+12p pd=1.688e+07u as=1.008e+11p ps=1.32e+06u
M1003 a_1924_48# a_1762_74# VGND VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1004 a_1115_74# a_781_74# a_995_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.89e+11p ps=1.74e+06u
M1005 Q_N a_1762_74# VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1006 VPWR a_1924_48# a_1712_374# VPB phighvt w=420000u l=150000u
+  ad=2.1112e+12p pd=1.868e+07u as=3.744e+11p ps=4.45e+06u
M1007 VGND SET_B a_1954_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_1600_347# a_995_74# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=5.8e+11p pd=5.16e+06u as=0p ps=0u
M1009 a_1600_347# a_594_74# a_1762_74# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=4.393e+11p ps=4.2e+06u
M1010 VGND SET_B a_1411_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1011 a_392_74# SCE a_290_464# VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=3.0425e+11p ps=3.2e+06u
M1012 VGND SCD a_392_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR SET_B a_1163_48# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.848e+11p ps=1.72e+06u
M1014 a_290_464# D a_206_464# VPB phighvt w=640000u l=150000u
+  ad=4.269e+11p pd=3.65e+06u as=1.728e+11p ps=1.82e+06u
M1015 a_1762_74# SET_B VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND a_1762_74# a_2556_112# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1017 a_995_74# a_781_74# a_290_464# VPB phighvt w=420000u l=150000u
+  ad=2.11725e+11p pd=1.9e+06u as=0p ps=0u
M1018 a_1133_478# a_594_74# a_995_74# VPB phighvt w=420000u l=150000u
+  ad=1.674e+11p pd=1.73e+06u as=0p ps=0u
M1019 VPWR CLK a_594_74# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.248e+11p ps=2.82e+06u
M1020 a_781_74# a_594_74# VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1021 Q a_2556_112# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.248e+11p pd=2.82e+06u as=0p ps=0u
M1022 VGND CLK a_594_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1023 a_1684_74# a_995_74# VGND VNB nshort w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1024 a_1762_74# a_781_74# a_1684_74# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPWR a_1163_48# a_1133_478# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VPWR SCE a_27_74# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.888e+11p ps=1.87e+06u
M1027 a_206_464# SCE VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 Q a_2556_112# VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1029 a_781_74# a_594_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.192e+11p pd=2.81e+06u as=0p ps=0u
M1030 VPWR a_1762_74# a_2556_112# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=2.436e+11p ps=2.26e+06u
M1031 VPWR SCD a_416_464# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1032 VPWR a_1762_74# a_1924_48# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.218e+11p ps=1.42e+06u
M1033 VGND SCE a_27_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1034 a_995_74# a_594_74# a_290_464# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_1762_74# a_781_74# a_1712_374# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_228_74# a_27_74# VGND VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1037 a_290_464# D a_228_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 Q_N a_1762_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.248e+11p pd=2.82e+06u as=0p ps=0u
M1039 a_416_464# a_27_74# a_290_464# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1040 a_1163_48# a_995_74# VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1041 a_1411_74# a_995_74# a_1163_48# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
.ends

