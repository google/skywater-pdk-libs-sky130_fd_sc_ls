* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
M1000 VGND A2 a_52_123# VNB nshort w=640000u l=150000u
+  ad=4.426e+11p pd=4.38e+06u as=3.52e+11p ps=3.66e+06u
M1001 a_222_392# B2 a_132_392# VPB phighvt w=1e+06u l=150000u
+  ad=3.3e+11p pd=2.66e+06u as=6.9e+11p ps=5.38e+06u
M1002 VPWR A1 a_132_392# VPB phighvt w=1e+06u l=150000u
+  ad=8.88e+11p pd=5.95e+06u as=0p ps=0u
M1003 a_230_79# B2 VGND VNB nshort w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1004 a_132_392# A2 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_52_123# A1 a_222_392# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1006 X a_222_392# VGND VNB nshort w=740000u l=150000u
+  ad=1.961e+11p pd=2.01e+06u as=0p ps=0u
M1007 a_132_392# B1 a_222_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_222_392# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.08e+11p pd=2.79e+06u as=0p ps=0u
M1009 a_222_392# B1 a_230_79# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
