* File: sky130_fd_sc_ls__or2b_1.pex.spice
* Created: Fri Aug 28 13:57:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__OR2B_1%B_N 1 2 3 5 6 8 10 11
r34 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.29
+ $Y=1.385 $X2=0.29 $Y2=1.385
r35 13 15 12.2197 $w=3.55e-07 $l=9e-08 $layer=POLY_cond $X=0.36 $Y=1.295
+ $X2=0.36 $Y2=1.385
r36 11 16 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.29 $Y=1.295 $X2=0.29
+ $Y2=1.385
r37 8 10 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=0.88 $Y=1.22
+ $X2=0.88 $Y2=0.835
r38 7 13 22.9692 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=0.565 $Y=1.295
+ $X2=0.36 $Y2=1.295
r39 6 8 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.805 $Y=1.295
+ $X2=0.88 $Y2=1.22
r40 6 7 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=0.805 $Y=1.295
+ $X2=0.565 $Y2=1.295
r41 3 5 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.505 $Y=2.045
+ $X2=0.505 $Y2=2.54
r42 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.505 $Y=1.955 $X2=0.505
+ $Y2=2.045
r43 1 15 54.4585 $w=3.55e-07 $l=3.80657e-07 $layer=POLY_cond $X=0.505 $Y=1.7
+ $X2=0.36 $Y2=1.385
r44 1 2 99.121 $w=1.8e-07 $l=2.55e-07 $layer=POLY_cond $X=0.505 $Y=1.7 $X2=0.505
+ $Y2=1.955
.ends

.subckt PM_SKY130_FD_SC_LS__OR2B_1%A_27_112# 1 2 9 11 13 14 15 20 22 23 24 25 26
+ 28 32
c69 11 0 1.50793e-20 $X=1.69 $Y=1.765
r70 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.36
+ $Y=1.465 $X2=1.36 $Y2=1.465
r71 26 34 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=0.745 $Y=1.465
+ $X2=0.745 $Y2=1.845
r72 26 28 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=0.83 $Y=1.465
+ $X2=1.36 $Y2=1.465
r73 25 26 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=0.745 $Y=1.3
+ $X2=0.745 $Y2=1.465
r74 24 32 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.745 $Y=1.01
+ $X2=0.745 $Y2=0.845
r75 24 25 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.745 $Y=1.01
+ $X2=0.745 $Y2=1.3
r76 22 34 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.66 $Y=1.845
+ $X2=0.745 $Y2=1.845
r77 22 23 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=0.66 $Y=1.845
+ $X2=0.445 $Y2=1.845
r78 18 23 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=1.93
+ $X2=0.445 $Y2=1.845
r79 18 20 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.28 $Y=1.93
+ $X2=0.28 $Y2=2.265
r80 14 29 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=1.59 $Y=1.465
+ $X2=1.36 $Y2=1.465
r81 14 15 5.03009 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.59 $Y=1.465
+ $X2=1.59 $Y2=1.3
r82 11 15 37.0704 $w=1.5e-07 $l=5.12567e-07 $layer=POLY_cond $X=1.69 $Y=1.765
+ $X2=1.59 $Y2=1.3
r83 11 13 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.69 $Y=1.765
+ $X2=1.69 $Y2=2.34
r84 7 15 37.0704 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.665 $Y=1.3 $X2=1.59
+ $Y2=1.3
r85 7 9 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.665 $Y=1.3
+ $X2=1.665 $Y2=0.835
r86 2 20 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.12 $X2=0.28 $Y2=2.265
r87 1 32 91 $w=1.7e-07 $l=6.57229e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.56 $X2=0.665 $Y2=0.845
.ends

.subckt PM_SKY130_FD_SC_LS__OR2B_1%A 3 5 7 8 12
c32 12 0 1.50793e-20 $X=2.2 $Y=1.515
r33 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.2
+ $Y=1.515 $X2=2.2 $Y2=1.515
r34 8 12 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=2.2 $Y=1.665 $X2=2.2
+ $Y2=1.515
r35 5 11 51.7056 $w=3.11e-07 $l=2.88097e-07 $layer=POLY_cond $X=2.11 $Y=1.765
+ $X2=2.192 $Y2=1.515
r36 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.11 $Y=1.765
+ $X2=2.11 $Y2=2.34
r37 1 11 38.532 $w=3.11e-07 $l=2.07918e-07 $layer=POLY_cond $X=2.095 $Y=1.35
+ $X2=2.192 $Y2=1.515
r38 1 3 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=2.095 $Y=1.35
+ $X2=2.095 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_LS__OR2B_1%A_264_368# 1 2 7 9 12 16 20 23 24 29 31
r68 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.77
+ $Y=1.465 $X2=2.77 $Y2=1.465
r69 27 29 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.465 $Y=1.905
+ $X2=1.78 $Y2=1.905
r70 25 31 2.90867 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=2.045 $Y=1.095
+ $X2=1.87 $Y2=1.095
r71 24 34 15.4589 $w=2.92e-07 $l=4.59238e-07 $layer=LI1_cond $X=2.535 $Y=1.095
+ $X2=2.735 $Y2=1.465
r72 24 25 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=2.535 $Y=1.095
+ $X2=2.045 $Y2=1.095
r73 23 29 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.78 $Y=1.82
+ $X2=1.78 $Y2=1.905
r74 22 31 3.58051 $w=2.6e-07 $l=1.25499e-07 $layer=LI1_cond $X=1.78 $Y=1.18
+ $X2=1.87 $Y2=1.095
r75 22 23 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=1.78 $Y=1.18 $X2=1.78
+ $Y2=1.82
r76 18 31 3.58051 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.87 $Y=1.01 $X2=1.87
+ $Y2=1.095
r77 18 20 5.76222 $w=3.48e-07 $l=1.75e-07 $layer=LI1_cond $X=1.87 $Y=1.01
+ $X2=1.87 $Y2=0.835
r78 16 27 24.6204 $w=3.28e-07 $l=7.05e-07 $layer=LI1_cond $X=1.465 $Y=2.695
+ $X2=1.465 $Y2=1.99
r79 10 35 38.6549 $w=2.86e-07 $l=1.90526e-07 $layer=POLY_cond $X=2.825 $Y=1.3
+ $X2=2.77 $Y2=1.465
r80 10 12 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.825 $Y=1.3
+ $X2=2.825 $Y2=0.74
r81 7 35 61.4066 $w=2.86e-07 $l=3.3541e-07 $layer=POLY_cond $X=2.695 $Y=1.765
+ $X2=2.77 $Y2=1.465
r82 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.695 $Y=1.765
+ $X2=2.695 $Y2=2.4
r83 2 27 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.32
+ $Y=1.84 $X2=1.465 $Y2=1.985
r84 2 16 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.32
+ $Y=1.84 $X2=1.465 $Y2=2.695
r85 1 20 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=1.74
+ $Y=0.56 $X2=1.88 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_LS__OR2B_1%VPWR 1 2 9 13 18 19 20 22 35 36 39
r37 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r38 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r39 33 36 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r40 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r41 30 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r42 29 32 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r43 29 30 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r44 27 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=0.78 $Y2=3.33
r45 27 29 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=1.2 $Y2=3.33
r46 25 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r47 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r48 22 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.78 $Y2=3.33
r49 22 24 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.24 $Y2=3.33
r50 20 33 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r51 20 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r52 18 32 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=2.255 $Y=3.33
+ $X2=2.16 $Y2=3.33
r53 18 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.255 $Y=3.33
+ $X2=2.42 $Y2=3.33
r54 17 35 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=2.585 $Y=3.33
+ $X2=3.12 $Y2=3.33
r55 17 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.585 $Y=3.33
+ $X2=2.42 $Y2=3.33
r56 13 16 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=2.42 $Y=2.115 $X2=2.42
+ $Y2=2.815
r57 11 19 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.42 $Y=3.245
+ $X2=2.42 $Y2=3.33
r58 11 16 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.42 $Y=3.245
+ $X2=2.42 $Y2=2.815
r59 7 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=3.245 $X2=0.78
+ $Y2=3.33
r60 7 9 34.2241 $w=3.28e-07 $l=9.8e-07 $layer=LI1_cond $X=0.78 $Y=3.245 $X2=0.78
+ $Y2=2.265
r61 2 16 600 $w=1.7e-07 $l=1.08616e-06 $layer=licon1_PDIFF $count=1 $X=2.185
+ $Y=1.84 $X2=2.42 $Y2=2.815
r62 2 13 300 $w=1.7e-07 $l=3.745e-07 $layer=licon1_PDIFF $count=2 $X=2.185
+ $Y=1.84 $X2=2.42 $Y2=2.115
r63 1 9 300 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=2 $X=0.58
+ $Y=2.12 $X2=0.78 $Y2=2.265
.ends

.subckt PM_SKY130_FD_SC_LS__OR2B_1%X 1 2 9 13 14 15 16 31 32 35
r23 31 32 9.6413 $w=5.18e-07 $l=1.65e-07 $layer=LI1_cond $X=3.015 $Y=1.985
+ $X2=3.015 $Y2=1.82
r24 21 35 1.03507 $w=5.18e-07 $l=4.5e-08 $layer=LI1_cond $X=3.015 $Y=2.08
+ $X2=3.015 $Y2=2.035
r25 16 28 0.92006 $w=5.18e-07 $l=4e-08 $layer=LI1_cond $X=3.015 $Y=2.775
+ $X2=3.015 $Y2=2.815
r26 15 16 8.51056 $w=5.18e-07 $l=3.7e-07 $layer=LI1_cond $X=3.015 $Y=2.405
+ $X2=3.015 $Y2=2.775
r27 14 35 0.46003 $w=5.18e-07 $l=2e-08 $layer=LI1_cond $X=3.015 $Y=2.015
+ $X2=3.015 $Y2=2.035
r28 14 31 0.690045 $w=5.18e-07 $l=3e-08 $layer=LI1_cond $X=3.015 $Y=2.015
+ $X2=3.015 $Y2=1.985
r29 14 15 7.01546 $w=5.18e-07 $l=3.05e-07 $layer=LI1_cond $X=3.015 $Y=2.1
+ $X2=3.015 $Y2=2.405
r30 14 21 0.46003 $w=5.18e-07 $l=2e-08 $layer=LI1_cond $X=3.015 $Y=2.1 $X2=3.015
+ $Y2=2.08
r31 13 32 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.19 $Y=1.13 $X2=3.19
+ $Y2=1.82
r32 7 13 9.656 $w=3.98e-07 $l=2e-07 $layer=LI1_cond $X=3.075 $Y=0.93 $X2=3.075
+ $Y2=1.13
r33 7 9 11.9566 $w=3.98e-07 $l=4.15e-07 $layer=LI1_cond $X=3.075 $Y=0.93
+ $X2=3.075 $Y2=0.515
r34 2 31 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.77
+ $Y=1.84 $X2=2.92 $Y2=1.985
r35 2 28 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.77
+ $Y=1.84 $X2=2.92 $Y2=2.815
r36 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.9 $Y=0.37
+ $X2=3.04 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__OR2B_1%VGND 1 2 9 13 16 17 18 20 30 31 34
r38 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r39 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r40 28 31 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r41 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r42 25 34 11.6267 $w=1.7e-07 $l=2.63e-07 $layer=LI1_cond $X=1.525 $Y=0 $X2=1.262
+ $Y2=0
r43 25 27 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.525 $Y=0 $X2=2.16
+ $Y2=0
r44 23 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r45 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r46 20 34 11.6267 $w=1.7e-07 $l=2.62e-07 $layer=LI1_cond $X=1 $Y=0 $X2=1.262
+ $Y2=0
r47 20 22 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1 $Y=0 $X2=0.72
+ $Y2=0
r48 18 28 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r49 18 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r50 16 27 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=2.265 $Y=0 $X2=2.16
+ $Y2=0
r51 16 17 10.0494 $w=1.7e-07 $l=2.07e-07 $layer=LI1_cond $X=2.265 $Y=0 $X2=2.472
+ $Y2=0
r52 15 30 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=2.68 $Y=0 $X2=3.12
+ $Y2=0
r53 15 17 10.0494 $w=1.7e-07 $l=2.08e-07 $layer=LI1_cond $X=2.68 $Y=0 $X2=2.472
+ $Y2=0
r54 11 17 1.57254 $w=4.15e-07 $l=8.5e-08 $layer=LI1_cond $X=2.472 $Y=0.085
+ $X2=2.472 $Y2=0
r55 11 13 16.6618 $w=4.13e-07 $l=6e-07 $layer=LI1_cond $X=2.472 $Y=0.085
+ $X2=2.472 $Y2=0.685
r56 7 34 2.19831 $w=5.25e-07 $l=8.5e-08 $layer=LI1_cond $X=1.262 $Y=0.085
+ $X2=1.262 $Y2=0
r57 7 9 17.0868 $w=5.23e-07 $l=7.5e-07 $layer=LI1_cond $X=1.262 $Y=0.085
+ $X2=1.262 $Y2=0.835
r58 2 13 182 $w=1.7e-07 $l=3.51994e-07 $layer=licon1_NDIFF $count=1 $X=2.17
+ $Y=0.56 $X2=2.465 $Y2=0.685
r59 1 9 91 $w=1.7e-07 $l=6.01997e-07 $layer=licon1_NDIFF $count=2 $X=0.955
+ $Y=0.56 $X2=1.435 $Y2=0.835
.ends

