# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ls__xor3_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ls__xor3_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.56000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.910000 1.180000 1.285000 1.670000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.693000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.910000 1.180000 5.240000 1.550000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.381000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.810000 1.450000 7.070000 1.780000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  1.086400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.685000 1.820000 9.125000 2.980000 ;
        RECT 8.830000 0.350000 9.160000 1.085000 ;
        RECT 8.955000 1.085000 9.160000 1.300000 ;
        RECT 8.955000 1.300000 9.940000 1.470000 ;
        RECT 8.955000 1.470000 9.125000 1.820000 ;
        RECT 9.665000 1.470000 9.940000 1.550000 ;
        RECT 9.665000 1.550000 9.995000 2.980000 ;
        RECT 9.690000 0.350000 9.940000 1.300000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 10.560000 0.085000 ;
        RECT  0.625000  0.085000  1.035000 0.410000 ;
        RECT  5.250000  0.085000  5.500000 0.610000 ;
        RECT  8.330000  0.085000  8.660000 1.085000 ;
        RECT  9.340000  0.085000  9.510000 1.130000 ;
        RECT 10.120000  0.085000 10.450000 1.130000 ;
      LAYER mcon ;
        RECT  0.155000 -0.085000  0.325000 0.085000 ;
        RECT  0.635000 -0.085000  0.805000 0.085000 ;
        RECT  1.115000 -0.085000  1.285000 0.085000 ;
        RECT  1.595000 -0.085000  1.765000 0.085000 ;
        RECT  2.075000 -0.085000  2.245000 0.085000 ;
        RECT  2.555000 -0.085000  2.725000 0.085000 ;
        RECT  3.035000 -0.085000  3.205000 0.085000 ;
        RECT  3.515000 -0.085000  3.685000 0.085000 ;
        RECT  3.995000 -0.085000  4.165000 0.085000 ;
        RECT  4.475000 -0.085000  4.645000 0.085000 ;
        RECT  4.955000 -0.085000  5.125000 0.085000 ;
        RECT  5.435000 -0.085000  5.605000 0.085000 ;
        RECT  5.915000 -0.085000  6.085000 0.085000 ;
        RECT  6.395000 -0.085000  6.565000 0.085000 ;
        RECT  6.875000 -0.085000  7.045000 0.085000 ;
        RECT  7.355000 -0.085000  7.525000 0.085000 ;
        RECT  7.835000 -0.085000  8.005000 0.085000 ;
        RECT  8.315000 -0.085000  8.485000 0.085000 ;
        RECT  8.795000 -0.085000  8.965000 0.085000 ;
        RECT  9.275000 -0.085000  9.445000 0.085000 ;
        RECT  9.755000 -0.085000  9.925000 0.085000 ;
        RECT 10.235000 -0.085000 10.405000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.560000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 3.245000 10.560000 3.415000 ;
        RECT  0.565000 2.180000  0.895000 3.245000 ;
        RECT  4.905000 1.820000  5.235000 3.245000 ;
        RECT  7.945000 1.820000  8.115000 2.330000 ;
        RECT  7.945000 2.330000  8.500000 3.245000 ;
        RECT  9.295000 1.820000  9.465000 3.245000 ;
        RECT 10.195000 1.820000 10.445000 3.245000 ;
      LAYER mcon ;
        RECT  0.155000 3.245000  0.325000 3.415000 ;
        RECT  0.635000 3.245000  0.805000 3.415000 ;
        RECT  1.115000 3.245000  1.285000 3.415000 ;
        RECT  1.595000 3.245000  1.765000 3.415000 ;
        RECT  2.075000 3.245000  2.245000 3.415000 ;
        RECT  2.555000 3.245000  2.725000 3.415000 ;
        RECT  3.035000 3.245000  3.205000 3.415000 ;
        RECT  3.515000 3.245000  3.685000 3.415000 ;
        RECT  3.995000 3.245000  4.165000 3.415000 ;
        RECT  4.475000 3.245000  4.645000 3.415000 ;
        RECT  4.955000 3.245000  5.125000 3.415000 ;
        RECT  5.435000 3.245000  5.605000 3.415000 ;
        RECT  5.915000 3.245000  6.085000 3.415000 ;
        RECT  6.395000 3.245000  6.565000 3.415000 ;
        RECT  6.875000 3.245000  7.045000 3.415000 ;
        RECT  7.355000 3.245000  7.525000 3.415000 ;
        RECT  7.835000 3.245000  8.005000 3.415000 ;
        RECT  8.315000 3.245000  8.485000 3.415000 ;
        RECT  8.795000 3.245000  8.965000 3.415000 ;
        RECT  9.275000 3.245000  9.445000 3.415000 ;
        RECT  9.755000 3.245000  9.925000 3.415000 ;
        RECT 10.235000 3.245000 10.405000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 10.560000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085000 0.570000 0.445000 0.580000 ;
      RECT 0.085000 0.580000 1.965000 0.750000 ;
      RECT 0.085000 0.750000 0.445000 1.250000 ;
      RECT 0.085000 1.250000 0.255000 2.180000 ;
      RECT 0.085000 2.180000 0.365000 2.980000 ;
      RECT 0.425000 1.470000 0.700000 1.840000 ;
      RECT 0.425000 1.840000 1.625000 2.010000 ;
      RECT 1.065000 2.010000 1.395000 2.905000 ;
      RECT 1.065000 2.905000 3.825000 3.075000 ;
      RECT 1.455000 0.920000 1.625000 1.840000 ;
      RECT 1.600000 2.180000 1.930000 2.565000 ;
      RECT 1.600000 2.565000 3.485000 2.735000 ;
      RECT 1.795000 0.750000 1.965000 1.420000 ;
      RECT 1.795000 1.420000 2.805000 1.590000 ;
      RECT 2.135000 0.450000 3.145000 0.620000 ;
      RECT 2.135000 0.620000 2.385000 1.250000 ;
      RECT 2.135000 1.590000 2.385000 2.395000 ;
      RECT 2.555000 0.790000 2.805000 1.420000 ;
      RECT 2.555000 1.875000 3.145000 2.395000 ;
      RECT 2.975000 0.620000 3.145000 1.875000 ;
      RECT 3.315000 0.255000 5.080000 0.425000 ;
      RECT 3.315000 0.425000 3.485000 2.565000 ;
      RECT 3.655000 0.595000 4.740000 0.765000 ;
      RECT 3.655000 0.765000 3.825000 1.435000 ;
      RECT 3.655000 1.435000 3.985000 1.735000 ;
      RECT 3.655000 1.905000 4.325000 2.755000 ;
      RECT 3.655000 2.755000 3.825000 2.905000 ;
      RECT 3.995000 0.935000 4.325000 1.265000 ;
      RECT 4.155000 1.265000 4.325000 1.905000 ;
      RECT 4.535000 0.765000 4.740000 1.130000 ;
      RECT 4.535000 1.130000 4.705000 2.980000 ;
      RECT 4.910000 0.425000 5.080000 0.780000 ;
      RECT 4.910000 0.780000 5.960000 0.950000 ;
      RECT 5.405000 1.920000 5.795000 2.800000 ;
      RECT 5.435000 1.120000 6.300000 1.290000 ;
      RECT 5.435000 1.290000 5.605000 1.920000 ;
      RECT 5.710000 0.255000 7.410000 0.425000 ;
      RECT 5.710000 0.425000 5.960000 0.780000 ;
      RECT 5.775000 1.460000 6.135000 1.750000 ;
      RECT 5.965000 1.750000 6.135000 2.905000 ;
      RECT 5.965000 2.905000 7.500000 3.075000 ;
      RECT 6.130000 0.595000 7.070000 0.765000 ;
      RECT 6.130000 0.765000 6.300000 1.120000 ;
      RECT 6.305000 1.920000 6.640000 2.735000 ;
      RECT 6.470000 0.935000 6.640000 1.920000 ;
      RECT 6.820000 0.765000 7.070000 1.275000 ;
      RECT 6.835000 1.950000 7.410000 2.120000 ;
      RECT 6.835000 2.120000 7.085000 2.735000 ;
      RECT 7.240000 0.425000 7.410000 1.950000 ;
      RECT 7.330000 2.290000 7.750000 2.710000 ;
      RECT 7.330000 2.710000 7.500000 2.905000 ;
      RECT 7.580000 0.415000 8.150000 0.745000 ;
      RECT 7.580000 0.745000 7.750000 2.290000 ;
      RECT 7.920000 1.255000 8.785000 1.585000 ;
      RECT 8.285000 1.585000 8.515000 2.150000 ;
    LAYER mcon ;
      RECT 2.555000 1.950000 2.725000 2.120000 ;
      RECT 5.435000 1.950000 5.605000 2.120000 ;
      RECT 6.395000 1.950000 6.565000 2.120000 ;
      RECT 8.315000 1.950000 8.485000 2.120000 ;
    LAYER met1 ;
      RECT 2.495000 1.920000 2.785000 1.965000 ;
      RECT 2.495000 1.965000 5.665000 2.105000 ;
      RECT 2.495000 2.105000 2.785000 2.150000 ;
      RECT 5.375000 1.920000 5.665000 1.965000 ;
      RECT 5.375000 2.105000 5.665000 2.150000 ;
      RECT 6.335000 1.920000 6.625000 1.965000 ;
      RECT 6.335000 1.965000 8.545000 2.105000 ;
      RECT 6.335000 2.105000 6.625000 2.150000 ;
      RECT 8.255000 1.920000 8.545000 1.965000 ;
      RECT 8.255000 2.105000 8.545000 2.150000 ;
  END
END sky130_fd_sc_ls__xor3_4
