* File: sky130_fd_sc_ls__a21bo_1.spice
* Created: Fri Aug 28 12:50:07 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__a21bo_1.pex.spice"
.subckt sky130_fd_sc_ls__a21bo_1  VNB VPB A2 A1 B1_N VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B1_N	B1_N
* A1	A1
* A2	A2
* VPB	VPB
* VNB	VNB
MM1001 A_122_136# N_A2_M1001_g N_VGND_M1001_s VNB NSHORT L=0.15 W=0.64 AD=0.0672
+ AS=0.1696 PD=0.85 PS=1.81 NRD=9.372 NRS=0 M=1 R=4.26667 SA=75000.2 SB=75001.1
+ A=0.096 P=1.58 MULT=1
MM1007 N_A_194_136#_M1007_d N_A1_M1007_g A_122_136# VNB NSHORT L=0.15 W=0.64
+ AD=0.1248 AS=0.0672 PD=1.03 PS=0.85 NRD=3.744 NRS=9.372 M=1 R=4.26667
+ SA=75000.6 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1003 N_VGND_M1003_d N_A_272_110#_M1003_g N_A_194_136#_M1007_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.1696 AS=0.1248 PD=1.81 PS=1.03 NRD=0 NRS=16.872 M=1
+ R=4.26667 SA=75001.1 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1006 N_VGND_M1006_d N_B1_N_M1006_g N_A_272_110#_M1006_s VNB NSHORT L=0.15
+ W=0.55 AD=0.0964632 AS=0.15675 PD=0.90814 PS=1.67 NRD=4.356 NRS=0 M=1
+ R=3.66667 SA=75000.2 SB=75000.7 A=0.0825 P=1.4 MULT=1
MM1002 N_X_M1002_d N_A_194_136#_M1002_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.74
+ AD=0.1961 AS=0.129787 PD=2.01 PS=1.22186 NRD=0 NRS=4.044 M=1 R=4.93333
+ SA=75000.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1004 N_VPWR_M1004_d N_A2_M1004_g N_A_34_392#_M1004_s VPB PHIGHVT L=0.15 W=1
+ AD=0.165 AS=0.275 PD=1.33 PS=2.55 NRD=4.9053 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75001.1 A=0.15 P=2.3 MULT=1
MM1008 N_A_34_392#_M1008_d N_A1_M1008_g N_VPWR_M1004_d VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.165 PD=1.3 PS=1.33 NRD=1.9503 NRS=4.9053 M=1 R=6.66667 SA=75000.7
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1000 N_A_194_136#_M1000_d N_A_272_110#_M1000_g N_A_34_392#_M1008_d VPB PHIGHVT
+ L=0.15 W=1 AD=0.275 AS=0.15 PD=2.55 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75001.1 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1005 N_VPWR_M1005_d N_B1_N_M1005_g N_A_272_110#_M1005_s VPB PHIGHVT L=0.15
+ W=0.84 AD=0.174 AS=0.231 PD=1.29 PS=2.23 NRD=35.6767 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75000.7 A=0.126 P=1.98 MULT=1
MM1009 N_X_M1009_d N_A_194_136#_M1009_g N_VPWR_M1005_d VPB PHIGHVT L=0.15 W=1.12
+ AD=0.308 AS=0.232 PD=2.79 PS=1.72 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.6 SB=75000.2 A=0.168 P=2.54 MULT=1
DX10_noxref VNB VPB NWDIODE A=7.8492 P=12.16
c_42 VNB 0 9.10919e-20 $X=0 $Y=0
*
.include "sky130_fd_sc_ls__a21bo_1.pxi.spice"
*
.ends
*
*
