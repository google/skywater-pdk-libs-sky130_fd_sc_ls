* NGSPICE file created from sky130_fd_sc_ls__o221ai_2.ext - technology: sky130A

.subckt sky130_fd_sc_ls__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
M1000 a_376_368# B1 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=7.672e+11p pd=5.85e+06u as=1.904e+12p ps=1.236e+07u
M1001 Y A2 a_776_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=1.0248e+12p pd=8.55e+06u as=7.28e+11p ps=5.78e+06u
M1002 a_311_85# A2 VGND VNB nshort w=740000u l=150000u
+  ad=1.0841e+12p pd=1.033e+07u as=5.328e+11p ps=4.4e+06u
M1003 VGND A1 a_311_85# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_776_368# A2 Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_27_74# B2 a_311_85# VNB nshort w=740000u l=150000u
+  ad=9.287e+11p pd=8.43e+06u as=0p ps=0u
M1006 VPWR A1 a_776_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_376_368# B2 Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND A2 a_311_85# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y B2 a_376_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_27_74# B1 a_311_85# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_311_85# B1 a_27_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR B1 a_376_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 Y C1 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR C1 Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y C1 a_27_74# VNB nshort w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1016 a_27_74# C1 Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_311_85# A1 VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_776_368# A1 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_311_85# B2 a_27_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

