* NGSPICE file created from sky130_fd_sc_ls__o21a_2.ext - technology: sky130A

.subckt sky130_fd_sc_ls__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
M1000 a_244_368# A2 a_160_368# VPB phighvt w=1e+06u l=150000u
+  ad=4.2e+11p pd=2.84e+06u as=2.7e+11p ps=2.54e+06u
M1001 a_160_368# A1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=1.2676e+12p ps=8.84e+06u
M1002 X a_244_368# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=0p ps=0u
M1003 X a_244_368# VGND VNB nshort w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=8.14e+11p ps=6.64e+06u
M1004 a_54_74# A2 VGND VNB nshort w=740000u l=150000u
+  ad=5.032e+11p pd=4.32e+06u as=0p ps=0u
M1005 VPWR a_244_368# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND A1 a_54_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND a_244_368# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_244_368# B1 a_54_74# VNB nshort w=740000u l=150000u
+  ad=2.627e+11p pd=2.19e+06u as=0p ps=0u
M1009 VPWR B1 a_244_368# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

