* NGSPICE file created from sky130_fd_sc_ls__buf_8.ext - technology: sky130A

.subckt sky130_fd_sc_ls__buf_8 A VGND VNB VPB VPWR X
M1000 VPWR a_27_74# X VPB phighvt w=1.12e+06u l=150000u
+  ad=2.1616e+12p pd=1.73e+07u as=1.4168e+12p ps=1.149e+07u
M1001 a_27_74# A VGND VNB nshort w=740000u l=150000u
+  ad=4.181e+11p pd=4.09e+06u as=1.591e+12p ps=1.318e+07u
M1002 X a_27_74# VGND VNB nshort w=740000u l=150000u
+  ad=8.325e+11p pd=8.17e+06u as=0p ps=0u
M1003 VPWR a_27_74# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR a_27_74# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 X a_27_74# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 X a_27_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND a_27_74# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND A a_27_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND a_27_74# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR A a_27_74# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=6.664e+11p ps=5.67e+06u
M1011 a_27_74# A VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 X a_27_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR a_27_74# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND a_27_74# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR A a_27_74# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 X a_27_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND A a_27_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 X a_27_74# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND a_27_74# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 X a_27_74# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 X a_27_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

