* NGSPICE file created from sky130_fd_sc_ls__a41o_1.ext - technology: sky130A

.subckt sky130_fd_sc_ls__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
M1000 a_543_74# A2 a_449_74# VNB nshort w=740000u l=150000u
+  ad=3.108e+11p pd=2.32e+06u as=2.368e+11p ps=2.12e+06u
M1001 a_354_392# A2 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=9.45e+11p pd=7.89e+06u as=1.1804e+12p ps=8.53e+06u
M1002 a_354_392# A4 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_449_74# A1 a_83_244# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.072e+11p ps=2.04e+06u
M1004 VPWR A3 a_354_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_354_392# B1 a_83_244# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.95e+11p ps=2.59e+06u
M1006 VGND a_83_244# X VNB nshort w=740000u l=150000u
+  ad=5.217e+11p pd=4.37e+06u as=7.104e+11p ps=3.4e+06u
M1007 a_657_74# A3 a_543_74# VNB nshort w=740000u l=150000u
+  ad=3.108e+11p pd=2.32e+06u as=0p ps=0u
M1008 VPWR a_83_244# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.304e+11p ps=2.83e+06u
M1009 VPWR A1 a_354_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_83_244# B1 VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND A4 a_657_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

