* File: sky130_fd_sc_ls__and4_4.pex.spice
* Created: Fri Aug 28 13:05:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__AND4_4%A 3 5 7 10 12 14 15 22
c51 15 0 5.84547e-20 $X=1.2 $Y=1.665
c52 12 0 1.94138e-19 $X=1.405 $Y=1.885
r53 22 23 3.09769 $w=3.89e-07 $l=2.5e-08 $layer=POLY_cond $X=1.38 $Y=1.667
+ $X2=1.405 $Y2=1.667
r54 20 22 19.2057 $w=3.89e-07 $l=1.55e-07 $layer=POLY_cond $X=1.225 $Y=1.667
+ $X2=1.38 $Y2=1.667
r55 18 20 33.455 $w=3.89e-07 $l=2.7e-07 $layer=POLY_cond $X=0.955 $Y=1.667
+ $X2=1.225 $Y2=1.667
r56 17 18 0.619537 $w=3.89e-07 $l=5e-09 $layer=POLY_cond $X=0.95 $Y=1.667
+ $X2=0.955 $Y2=1.667
r57 15 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.225
+ $Y=1.615 $X2=1.225 $Y2=1.615
r58 12 23 25.1816 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=1.405 $Y=1.885
+ $X2=1.405 $Y2=1.667
r59 12 14 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.405 $Y=1.885
+ $X2=1.405 $Y2=2.46
r60 8 22 25.1816 $w=1.5e-07 $l=2.17e-07 $layer=POLY_cond $X=1.38 $Y=1.45
+ $X2=1.38 $Y2=1.667
r61 8 10 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=1.38 $Y=1.45 $X2=1.38
+ $Y2=0.915
r62 5 18 25.1816 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=0.955 $Y=1.885
+ $X2=0.955 $Y2=1.667
r63 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.955 $Y=1.885
+ $X2=0.955 $Y2=2.46
r64 1 17 25.1816 $w=1.5e-07 $l=2.17e-07 $layer=POLY_cond $X=0.95 $Y=1.45
+ $X2=0.95 $Y2=1.667
r65 1 3 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=0.95 $Y=1.45 $X2=0.95
+ $Y2=0.915
.ends

.subckt PM_SKY130_FD_SC_LS__AND4_4%B 1 3 7 8 9 13 16 18 20 21 22 26
c64 20 0 5.28639e-20 $X=1.832 $Y=1.46
c65 16 0 1.27581e-19 $X=1.87 $Y=1.885
r66 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.615 $X2=0.385 $Y2=1.615
r67 22 26 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=0.24 $Y=1.615
+ $X2=0.385 $Y2=1.615
r68 20 21 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=1.855 $Y=1.46
+ $X2=1.855 $Y2=1.7
r69 19 20 51.0119 $w=1.95e-07 $l=1.5e-07 $layer=POLY_cond $X=1.832 $Y=1.31
+ $X2=1.832 $Y2=1.46
r70 16 21 71.9113 $w=1.8e-07 $l=1.85e-07 $layer=POLY_cond $X=1.87 $Y=1.885
+ $X2=1.87 $Y2=1.7
r71 16 18 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.87 $Y=1.885
+ $X2=1.87 $Y2=2.46
r72 13 19 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.81 $Y=0.915
+ $X2=1.81 $Y2=1.31
r73 10 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.81 $Y=0.255
+ $X2=1.81 $Y2=0.915
r74 8 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.735 $Y=0.18
+ $X2=1.81 $Y2=0.255
r75 8 9 584.553 $w=1.5e-07 $l=1.14e-06 $layer=POLY_cond $X=1.735 $Y=0.18
+ $X2=0.595 $Y2=0.18
r76 5 25 38.5818 $w=3.27e-07 $l=2.14173e-07 $layer=POLY_cond $X=0.52 $Y=1.45
+ $X2=0.407 $Y2=1.615
r77 5 7 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=0.52 $Y=1.45 $X2=0.52
+ $Y2=0.915
r78 4 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.52 $Y=0.255
+ $X2=0.595 $Y2=0.18
r79 4 7 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.52 $Y=0.255 $X2=0.52
+ $Y2=0.915
r80 1 25 54.0589 $w=3.27e-07 $l=3.15214e-07 $layer=POLY_cond $X=0.505 $Y=1.885
+ $X2=0.407 $Y2=1.615
r81 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.505 $Y=1.885
+ $X2=0.505 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_LS__AND4_4%D 1 3 4 6 7 9 10 11 12 14 15 17
c61 17 0 4.10416e-20 $X=3.12 $Y=1.665
r62 22 24 18.9357 $w=4.2e-07 $l=1.65e-07 $layer=POLY_cond $X=3.095 $Y=1.615
+ $X2=3.26 $Y2=1.615
r63 20 22 31.5595 $w=4.2e-07 $l=2.75e-07 $layer=POLY_cond $X=2.82 $Y=1.615
+ $X2=3.095 $Y2=1.615
r64 17 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.095
+ $Y=1.635 $X2=3.095 $Y2=1.635
r65 12 15 64.3434 $w=1.8e-07 $l=1.6e-07 $layer=POLY_cond $X=3.705 $Y=1.885
+ $X2=3.705 $Y2=1.725
r66 12 14 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.705 $Y=1.885
+ $X2=3.705 $Y2=2.46
r67 11 24 29.6695 $w=4.2e-07 $l=1.42653e-07 $layer=POLY_cond $X=3.335 $Y=1.725
+ $X2=3.26 $Y2=1.615
r68 10 15 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.615 $Y=1.725
+ $X2=3.705 $Y2=1.725
r69 10 11 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.615 $Y=1.725
+ $X2=3.335 $Y2=1.725
r70 7 24 27.059 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=3.26 $Y=1.345 $X2=3.26
+ $Y2=1.615
r71 7 9 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.26 $Y=1.345 $X2=3.26
+ $Y2=0.915
r72 4 20 27.059 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.82 $Y=1.885 $X2=2.82
+ $Y2=1.615
r73 4 6 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.82 $Y=1.885
+ $X2=2.82 $Y2=2.46
r74 1 20 17.2143 $w=4.2e-07 $l=3.36749e-07 $layer=POLY_cond $X=2.67 $Y=1.345
+ $X2=2.82 $Y2=1.615
r75 1 3 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.67 $Y=1.345 $X2=2.67
+ $Y2=0.915
.ends

.subckt PM_SKY130_FD_SC_LS__AND4_4%C 4 9 10 11 14 16 19 20 22 24 25 26 27 28 32
c92 32 0 4.03165e-20 $X=4.2 $Y=1.51
c93 26 0 4.10416e-20 $X=2.347 $Y=1.885
r94 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.2
+ $Y=1.51 $X2=4.2 $Y2=1.51
r95 28 32 4.63971 $w=3.83e-07 $l=1.55e-07 $layer=LI1_cond $X=4.172 $Y=1.665
+ $X2=4.172 $Y2=1.51
r96 25 26 42.7811 $w=2.25e-07 $l=1.5e-07 $layer=POLY_cond $X=2.347 $Y=1.735
+ $X2=2.347 $Y2=1.885
r97 24 25 141.011 $w=1.5e-07 $l=2.75e-07 $layer=POLY_cond $X=2.31 $Y=1.46
+ $X2=2.31 $Y2=1.735
r98 23 24 43.7534 $w=2.2e-07 $l=1.5e-07 $layer=POLY_cond $X=2.275 $Y=1.31
+ $X2=2.275 $Y2=1.46
r99 20 31 76.233 $w=2.71e-07 $l=3.77492e-07 $layer=POLY_cond $X=4.205 $Y=1.885
+ $X2=4.2 $Y2=1.51
r100 20 22 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=4.205 $Y=1.885
+ $X2=4.205 $Y2=2.46
r101 19 31 38.8824 $w=2.71e-07 $l=1.65e-07 $layer=POLY_cond $X=4.2 $Y=1.345
+ $X2=4.2 $Y2=1.51
r102 18 19 558.915 $w=1.5e-07 $l=1.09e-06 $layer=POLY_cond $X=4.2 $Y=0.255
+ $X2=4.2 $Y2=1.345
r103 17 27 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.765 $Y=0.18
+ $X2=3.69 $Y2=0.18
r104 16 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.125 $Y=0.18
+ $X2=4.2 $Y2=0.255
r105 16 17 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=4.125 $Y=0.18
+ $X2=3.765 $Y2=0.18
r106 12 27 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.69 $Y=0.255
+ $X2=3.69 $Y2=0.18
r107 12 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.69 $Y=0.255
+ $X2=3.69 $Y2=0.915
r108 10 27 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.615 $Y=0.18
+ $X2=3.69 $Y2=0.18
r109 10 11 666.596 $w=1.5e-07 $l=1.3e-06 $layer=POLY_cond $X=3.615 $Y=0.18
+ $X2=2.315 $Y2=0.18
r110 9 26 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.37 $Y=2.46
+ $X2=2.37 $Y2=1.885
r111 4 23 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.24 $Y=0.915
+ $X2=2.24 $Y2=1.31
r112 1 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.24 $Y=0.255
+ $X2=2.315 $Y2=0.18
r113 1 4 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.24 $Y=0.255
+ $X2=2.24 $Y2=0.915
.ends

.subckt PM_SKY130_FD_SC_LS__AND4_4%A_116_392# 1 2 3 4 5 18 20 22 25 27 29 32 34
+ 36 39 41 43 45 46 48 50 53 56 58 59 61 64 66 70 72 75 76 81 87 89 91 100
c193 87 0 8.82342e-20 $X=1.645 $Y=2.105
c194 75 0 1.74227e-19 $X=4.62 $Y=1.95
c195 46 0 1.43623e-19 $X=0.89 $Y=1.13
c196 45 0 1.94138e-19 $X=0.805 $Y=1.95
c197 20 0 4.03165e-20 $X=4.765 $Y=1.765
c198 18 0 1.8401e-19 $X=4.75 $Y=0.74
r199 100 101 3.08184 $w=3.91e-07 $l=2.5e-08 $layer=POLY_cond $X=6.14 $Y=1.532
+ $X2=6.165 $Y2=1.532
r200 99 100 52.3913 $w=3.91e-07 $l=4.25e-07 $layer=POLY_cond $X=5.715 $Y=1.532
+ $X2=6.14 $Y2=1.532
r201 98 99 0.616368 $w=3.91e-07 $l=5e-09 $layer=POLY_cond $X=5.71 $Y=1.532
+ $X2=5.715 $Y2=1.532
r202 95 96 6.78005 $w=3.91e-07 $l=5.5e-08 $layer=POLY_cond $X=5.21 $Y=1.532
+ $X2=5.265 $Y2=1.532
r203 92 93 1.8491 $w=3.91e-07 $l=1.5e-08 $layer=POLY_cond $X=4.75 $Y=1.532
+ $X2=4.765 $Y2=1.532
r204 82 98 23.422 $w=3.91e-07 $l=1.9e-07 $layer=POLY_cond $X=5.52 $Y=1.532
+ $X2=5.71 $Y2=1.532
r205 82 96 31.4348 $w=3.91e-07 $l=2.55e-07 $layer=POLY_cond $X=5.52 $Y=1.532
+ $X2=5.265 $Y2=1.532
r206 81 82 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=5.52
+ $Y=1.465 $X2=5.52 $Y2=1.465
r207 79 95 45.6113 $w=3.91e-07 $l=3.7e-07 $layer=POLY_cond $X=4.84 $Y=1.532
+ $X2=5.21 $Y2=1.532
r208 79 93 9.24552 $w=3.91e-07 $l=7.5e-08 $layer=POLY_cond $X=4.84 $Y=1.532
+ $X2=4.765 $Y2=1.532
r209 78 81 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=4.84 $Y=1.465
+ $X2=5.52 $Y2=1.465
r210 78 79 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=4.84
+ $Y=1.465 $X2=4.84 $Y2=1.465
r211 76 78 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=4.705 $Y=1.465
+ $X2=4.84 $Y2=1.465
r212 74 76 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.62 $Y=1.63
+ $X2=4.705 $Y2=1.465
r213 74 75 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=4.62 $Y=1.63
+ $X2=4.62 $Y2=1.95
r214 73 91 8.61065 $w=1.7e-07 $l=1.69926e-07 $layer=LI1_cond $X=4.145 $Y=2.035
+ $X2=3.98 $Y2=2.045
r215 72 75 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.535 $Y=2.035
+ $X2=4.62 $Y2=1.95
r216 72 73 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=4.535 $Y=2.035
+ $X2=4.145 $Y2=2.035
r217 68 91 0.89609 $w=3.3e-07 $l=9.5e-08 $layer=LI1_cond $X=3.98 $Y=2.14
+ $X2=3.98 $Y2=2.045
r218 68 70 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=3.98 $Y=2.14
+ $X2=3.98 $Y2=2.815
r219 67 89 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.76 $Y=2.055
+ $X2=2.595 $Y2=2.055
r220 66 91 8.61065 $w=1.7e-07 $l=1.69926e-07 $layer=LI1_cond $X=3.815 $Y=2.055
+ $X2=3.98 $Y2=2.045
r221 66 67 68.8289 $w=1.68e-07 $l=1.055e-06 $layer=LI1_cond $X=3.815 $Y=2.055
+ $X2=2.76 $Y2=2.055
r222 62 89 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.595 $Y=2.14
+ $X2=2.595 $Y2=2.055
r223 62 64 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.595 $Y=2.14
+ $X2=2.595 $Y2=2.815
r224 61 89 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.595 $Y=1.97
+ $X2=2.595 $Y2=2.055
r225 60 61 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=2.595 $Y=1.77
+ $X2=2.595 $Y2=1.97
r226 58 60 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.43 $Y=1.685
+ $X2=2.595 $Y2=1.77
r227 58 59 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=2.43 $Y=1.685
+ $X2=1.73 $Y2=1.685
r228 54 87 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=1.645 $Y=2.24
+ $X2=1.645 $Y2=2.095
r229 54 56 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=1.645 $Y=2.24
+ $X2=1.645 $Y2=2.46
r230 53 87 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=1.645 $Y=1.95
+ $X2=1.645 $Y2=2.095
r231 52 59 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.645 $Y=1.77
+ $X2=1.73 $Y2=1.685
r232 52 53 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.645 $Y=1.77
+ $X2=1.645 $Y2=1.95
r233 51 85 3.14085 $w=2.9e-07 $l=1.63e-07 $layer=LI1_cond $X=0.89 $Y=2.095
+ $X2=0.727 $Y2=2.095
r234 50 87 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.56 $Y=2.095
+ $X2=1.645 $Y2=2.095
r235 50 51 26.6254 $w=2.88e-07 $l=6.7e-07 $layer=LI1_cond $X=1.56 $Y=2.095
+ $X2=0.89 $Y2=2.095
r236 46 48 12.6769 $w=2.48e-07 $l=2.75e-07 $layer=LI1_cond $X=0.89 $Y=1.13
+ $X2=1.165 $Y2=1.13
r237 45 85 4.29699 $w=1.7e-07 $l=1.79819e-07 $layer=LI1_cond $X=0.805 $Y=1.95
+ $X2=0.727 $Y2=2.095
r238 44 46 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.805 $Y=1.255
+ $X2=0.89 $Y2=1.13
r239 44 45 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=0.805 $Y=1.255
+ $X2=0.805 $Y2=1.95
r240 41 101 25.3065 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=6.165 $Y=1.765
+ $X2=6.165 $Y2=1.532
r241 41 43 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.165 $Y=1.765
+ $X2=6.165 $Y2=2.4
r242 37 100 25.3065 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=6.14 $Y=1.3
+ $X2=6.14 $Y2=1.532
r243 37 39 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=6.14 $Y=1.3
+ $X2=6.14 $Y2=0.74
r244 34 99 25.3065 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=5.715 $Y=1.765
+ $X2=5.715 $Y2=1.532
r245 34 36 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.715 $Y=1.765
+ $X2=5.715 $Y2=2.4
r246 30 98 25.3065 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=5.71 $Y=1.3
+ $X2=5.71 $Y2=1.532
r247 30 32 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=5.71 $Y=1.3
+ $X2=5.71 $Y2=0.74
r248 27 96 25.3065 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=5.265 $Y=1.765
+ $X2=5.265 $Y2=1.532
r249 27 29 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.265 $Y=1.765
+ $X2=5.265 $Y2=2.4
r250 23 95 25.3065 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=5.21 $Y=1.3
+ $X2=5.21 $Y2=1.532
r251 23 25 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=5.21 $Y=1.3
+ $X2=5.21 $Y2=0.74
r252 20 93 25.3065 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=4.765 $Y=1.765
+ $X2=4.765 $Y2=1.532
r253 20 22 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.765 $Y=1.765
+ $X2=4.765 $Y2=2.4
r254 16 92 25.3065 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=4.75 $Y=1.3
+ $X2=4.75 $Y2=1.532
r255 16 18 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.75 $Y=1.3
+ $X2=4.75 $Y2=0.74
r256 5 91 400 $w=1.7e-07 $l=2.66458e-07 $layer=licon1_PDIFF $count=1 $X=3.78
+ $Y=1.96 $X2=3.98 $Y2=2.115
r257 5 70 400 $w=1.7e-07 $l=9.4975e-07 $layer=licon1_PDIFF $count=1 $X=3.78
+ $Y=1.96 $X2=3.98 $Y2=2.815
r258 4 89 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.445
+ $Y=1.96 $X2=2.595 $Y2=2.105
r259 4 64 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=2.445
+ $Y=1.96 $X2=2.595 $Y2=2.815
r260 3 87 600 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_PDIFF $count=1 $X=1.48
+ $Y=1.96 $X2=1.645 $Y2=2.105
r261 3 56 300 $w=1.7e-07 $l=5.76628e-07 $layer=licon1_PDIFF $count=2 $X=1.48
+ $Y=1.96 $X2=1.645 $Y2=2.46
r262 2 85 600 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.96 $X2=0.73 $Y2=2.115
r263 1 48 182 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_NDIFF $count=1 $X=1.025
+ $Y=0.595 $X2=1.165 $Y2=1.09
.ends

.subckt PM_SKY130_FD_SC_LS__AND4_4%VPWR 1 2 3 4 5 6 7 22 24 30 34 40 44 48 50 52
+ 56 58 63 68 73 78 83 92 95 98 101 104 108
r100 107 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r101 104 105 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r102 101 102 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r103 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r104 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r105 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r106 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r107 87 108 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=6.48 $Y2=3.33
r108 87 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=5.52 $Y2=3.33
r109 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r110 84 104 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.655 $Y=3.33
+ $X2=5.53 $Y2=3.33
r111 84 86 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=5.655 $Y=3.33 $X2=6
+ $Y2=3.33
r112 83 107 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=6.275 $Y=3.33
+ $X2=6.497 $Y2=3.33
r113 83 86 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.275 $Y=3.33
+ $X2=6 $Y2=3.33
r114 82 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r115 82 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r116 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r117 79 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.645 $Y=3.33
+ $X2=4.48 $Y2=3.33
r118 79 81 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=4.645 $Y=3.33
+ $X2=5.04 $Y2=3.33
r119 78 104 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.405 $Y=3.33
+ $X2=5.53 $Y2=3.33
r120 78 81 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=5.405 $Y=3.33
+ $X2=5.04 $Y2=3.33
r121 77 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r122 76 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r123 74 98 13.8148 $w=1.7e-07 $l=3.58e-07 $layer=LI1_cond $X=3.645 $Y=3.33
+ $X2=3.287 $Y2=3.33
r124 74 76 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=3.645 $Y=3.33
+ $X2=4.08 $Y2=3.33
r125 73 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.315 $Y=3.33
+ $X2=4.48 $Y2=3.33
r126 73 76 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=4.315 $Y=3.33
+ $X2=4.08 $Y2=3.33
r127 72 99 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r128 72 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r129 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r130 69 95 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.26 $Y=3.33
+ $X2=2.095 $Y2=3.33
r131 69 71 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=2.26 $Y=3.33
+ $X2=2.64 $Y2=3.33
r132 68 98 13.8148 $w=1.7e-07 $l=3.57e-07 $layer=LI1_cond $X=2.93 $Y=3.33
+ $X2=3.287 $Y2=3.33
r133 68 71 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=2.93 $Y=3.33
+ $X2=2.64 $Y2=3.33
r134 67 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r135 67 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r136 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r137 64 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.345 $Y=3.33
+ $X2=1.18 $Y2=3.33
r138 64 66 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.345 $Y=3.33
+ $X2=1.68 $Y2=3.33
r139 63 95 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.93 $Y=3.33
+ $X2=2.095 $Y2=3.33
r140 63 66 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.93 $Y=3.33
+ $X2=1.68 $Y2=3.33
r141 62 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r142 62 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r143 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r144 59 89 4.27358 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=0.395 $Y=3.33
+ $X2=0.197 $Y2=3.33
r145 59 61 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.395 $Y=3.33
+ $X2=0.72 $Y2=3.33
r146 58 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.015 $Y=3.33
+ $X2=1.18 $Y2=3.33
r147 58 61 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.015 $Y=3.33
+ $X2=0.72 $Y2=3.33
r148 56 77 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=4.08 $Y2=3.33
r149 56 99 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=3.12 $Y2=3.33
r150 52 55 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=6.44 $Y=1.985
+ $X2=6.44 $Y2=2.815
r151 50 107 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=6.44 $Y=3.245
+ $X2=6.497 $Y2=3.33
r152 50 55 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=6.44 $Y=3.245
+ $X2=6.44 $Y2=2.815
r153 46 104 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.53 $Y=3.245
+ $X2=5.53 $Y2=3.33
r154 46 48 43.3319 $w=2.48e-07 $l=9.4e-07 $layer=LI1_cond $X=5.53 $Y=3.245
+ $X2=5.53 $Y2=2.305
r155 42 101 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.48 $Y=3.245
+ $X2=4.48 $Y2=3.33
r156 42 44 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=4.48 $Y=3.245
+ $X2=4.48 $Y2=2.455
r157 38 98 2.90666 $w=7.15e-07 $l=8.5e-08 $layer=LI1_cond $X=3.287 $Y=3.245
+ $X2=3.287 $Y2=3.33
r158 38 40 12.8808 $w=7.13e-07 $l=7.7e-07 $layer=LI1_cond $X=3.287 $Y=3.245
+ $X2=3.287 $Y2=2.475
r159 34 37 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=2.095 $Y=2.105
+ $X2=2.095 $Y2=2.815
r160 32 95 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.095 $Y=3.245
+ $X2=2.095 $Y2=3.33
r161 32 37 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.095 $Y=3.245
+ $X2=2.095 $Y2=2.815
r162 28 92 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.18 $Y=3.245
+ $X2=1.18 $Y2=3.33
r163 28 30 26.1919 $w=3.28e-07 $l=7.5e-07 $layer=LI1_cond $X=1.18 $Y=3.245
+ $X2=1.18 $Y2=2.495
r164 24 27 28.8111 $w=2.78e-07 $l=7e-07 $layer=LI1_cond $X=0.255 $Y=2.115
+ $X2=0.255 $Y2=2.815
r165 22 89 3.08647 $w=2.8e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.255 $Y=3.245
+ $X2=0.197 $Y2=3.33
r166 22 27 17.6982 $w=2.78e-07 $l=4.3e-07 $layer=LI1_cond $X=0.255 $Y=3.245
+ $X2=0.255 $Y2=2.815
r167 7 55 400 $w=1.7e-07 $l=1.07034e-06 $layer=licon1_PDIFF $count=1 $X=6.24
+ $Y=1.84 $X2=6.44 $Y2=2.815
r168 7 52 400 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=1 $X=6.24
+ $Y=1.84 $X2=6.44 $Y2=1.985
r169 6 48 300 $w=1.7e-07 $l=5.34766e-07 $layer=licon1_PDIFF $count=2 $X=5.34
+ $Y=1.84 $X2=5.49 $Y2=2.305
r170 5 44 300 $w=1.7e-07 $l=5.86536e-07 $layer=licon1_PDIFF $count=2 $X=4.28
+ $Y=1.96 $X2=4.48 $Y2=2.455
r171 4 40 150 $w=1.7e-07 $l=8.02185e-07 $layer=licon1_PDIFF $count=4 $X=2.895
+ $Y=1.96 $X2=3.48 $Y2=2.475
r172 3 37 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=1.945
+ $Y=1.96 $X2=2.095 $Y2=2.815
r173 3 34 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.945
+ $Y=1.96 $X2=2.095 $Y2=2.105
r174 2 30 300 $w=1.7e-07 $l=6.05372e-07 $layer=licon1_PDIFF $count=2 $X=1.03
+ $Y=1.96 $X2=1.18 $Y2=2.495
r175 1 27 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.28 $Y2=2.815
r176 1 24 400 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.28 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_LS__AND4_4%X 1 2 3 4 15 19 23 24 25 26 29 32 35 39 41 42
+ 43 44 47
c78 32 0 8.56004e-20 $X=5.98 $Y=1.8
c79 24 0 1.8401e-19 $X=5.08 $Y=1.045
r80 46 47 9.26965 $w=2.28e-07 $l=1.85e-07 $layer=LI1_cond $X=6.48 $Y=1.48
+ $X2=6.48 $Y2=1.295
r81 45 47 8.26753 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=6.48 $Y=1.13
+ $X2=6.48 $Y2=1.295
r82 41 46 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=6.365 $Y=1.565
+ $X2=6.48 $Y2=1.48
r83 41 42 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=6.365 $Y=1.565
+ $X2=6.105 $Y2=1.565
r84 40 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.09 $Y=1.045
+ $X2=5.925 $Y2=1.045
r85 39 45 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=6.365 $Y=1.045
+ $X2=6.48 $Y2=1.13
r86 39 40 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.365 $Y=1.045
+ $X2=6.09 $Y2=1.045
r87 35 37 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=5.98 $Y=1.985
+ $X2=5.98 $Y2=2.815
r88 33 44 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.98 $Y=1.97 $X2=5.98
+ $Y2=1.885
r89 33 35 0.691466 $w=2.48e-07 $l=1.5e-08 $layer=LI1_cond $X=5.98 $Y=1.97
+ $X2=5.98 $Y2=1.985
r90 32 44 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.98 $Y=1.8 $X2=5.98
+ $Y2=1.885
r91 31 42 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.98 $Y=1.65
+ $X2=6.105 $Y2=1.565
r92 31 32 6.91466 $w=2.48e-07 $l=1.5e-07 $layer=LI1_cond $X=5.98 $Y=1.65
+ $X2=5.98 $Y2=1.8
r93 27 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.925 $Y=0.96
+ $X2=5.925 $Y2=1.045
r94 27 29 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=5.925 $Y=0.96
+ $X2=5.925 $Y2=0.515
r95 25 44 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.855 $Y=1.885
+ $X2=5.98 $Y2=1.885
r96 25 26 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=5.855 $Y=1.885
+ $X2=5.205 $Y2=1.885
r97 23 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.76 $Y=1.045
+ $X2=5.925 $Y2=1.045
r98 23 24 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=5.76 $Y=1.045
+ $X2=5.08 $Y2=1.045
r99 19 21 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=5.04 $Y=1.985
+ $X2=5.04 $Y2=2.815
r100 17 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.04 $Y=1.97
+ $X2=5.205 $Y2=1.885
r101 17 19 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=5.04 $Y=1.97
+ $X2=5.04 $Y2=1.985
r102 13 24 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.955 $Y=0.96
+ $X2=5.08 $Y2=1.045
r103 13 15 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=4.955 $Y=0.96
+ $X2=4.955 $Y2=0.515
r104 4 37 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=5.79
+ $Y=1.84 $X2=5.94 $Y2=2.815
r105 4 35 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=5.79
+ $Y=1.84 $X2=5.94 $Y2=1.985
r106 3 21 400 $w=1.7e-07 $l=1.07034e-06 $layer=licon1_PDIFF $count=1 $X=4.84
+ $Y=1.84 $X2=5.04 $Y2=2.815
r107 3 19 400 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=1 $X=4.84
+ $Y=1.84 $X2=5.04 $Y2=1.985
r108 2 29 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.785
+ $Y=0.37 $X2=5.925 $Y2=0.515
r109 1 15 91 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_NDIFF $count=2 $X=4.825
+ $Y=0.37 $X2=4.995 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__AND4_4%A_32_119# 1 2 3 12 14 15 19 20 21
c49 21 0 1.2199e-19 $X=2.11 $Y=1.215
r50 20 23 14.9533 $w=2.29e-07 $l=2.97061e-07 $layer=LI1_cond $X=3.64 $Y=1.215
+ $X2=3.905 $Y2=1.147
r51 20 21 99.8182 $w=1.68e-07 $l=1.53e-06 $layer=LI1_cond $X=3.64 $Y=1.215
+ $X2=2.11 $Y2=1.215
r52 17 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.025 $Y=1.13
+ $X2=2.11 $Y2=1.215
r53 17 19 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=2.025 $Y=1.13
+ $X2=2.025 $Y2=0.74
r54 16 19 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.025 $Y=0.485
+ $X2=2.025 $Y2=0.74
r55 14 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.94 $Y=0.4
+ $X2=2.025 $Y2=0.485
r56 14 15 101.123 $w=1.68e-07 $l=1.55e-06 $layer=LI1_cond $X=1.94 $Y=0.4
+ $X2=0.39 $Y2=0.4
r57 10 15 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.265 $Y=0.485
+ $X2=0.39 $Y2=0.4
r58 10 12 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=0.265 $Y=0.485
+ $X2=0.265 $Y2=0.74
r59 3 23 182 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_NDIFF $count=1 $X=3.765
+ $Y=0.595 $X2=3.905 $Y2=1.085
r60 2 19 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.885
+ $Y=0.595 $X2=2.025 $Y2=0.74
r61 1 12 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.16
+ $Y=0.595 $X2=0.305 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__AND4_4%A_119_119# 1 2 11
r10 8 11 52.9899 $w=1.78e-07 $l=8.6e-07 $layer=LI1_cond $X=0.735 $Y=0.745
+ $X2=1.595 $Y2=0.745
r11 2 11 182 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=1 $X=1.455
+ $Y=0.595 $X2=1.595 $Y2=0.745
r12 1 8 182 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.595 $X2=0.735 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_LS__AND4_4%A_463_119# 1 2 7 10 15
r29 15 16 5.88214 $w=2.8e-07 $l=1.35e-07 $layer=LI1_cond $X=3.47 $Y=0.74
+ $X2=3.47 $Y2=0.875
r30 10 12 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=2.455 $Y=0.765
+ $X2=2.455 $Y2=0.875
r31 8 12 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.62 $Y=0.875
+ $X2=2.455 $Y2=0.875
r32 7 16 3.65648 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=3.3 $Y=0.875 $X2=3.47
+ $Y2=0.875
r33 7 8 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.3 $Y=0.875 $X2=2.62
+ $Y2=0.875
r34 2 15 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.335
+ $Y=0.595 $X2=3.475 $Y2=0.74
r35 1 10 182 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_NDIFF $count=1 $X=2.315
+ $Y=0.595 $X2=2.455 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LS__AND4_4%VGND 1 2 3 4 15 19 23 25 27 30 31 32 34 42 51
+ 56 59 63
r74 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r75 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r76 56 57 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r77 54 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r78 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6 $Y2=0
r79 51 62 3.99713 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=6.26 $Y=0 $X2=6.49
+ $Y2=0
r80 51 53 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=6.26 $Y=0 $X2=6
+ $Y2=0
r81 50 54 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=6
+ $Y2=0
r82 50 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.56
+ $Y2=0
r83 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r84 47 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.66 $Y=0 $X2=4.495
+ $Y2=0
r85 47 49 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=4.66 $Y=0 $X2=5.04
+ $Y2=0
r86 46 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r87 45 46 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r88 43 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.13 $Y=0 $X2=2.965
+ $Y2=0
r89 43 45 61.9786 $w=1.68e-07 $l=9.5e-07 $layer=LI1_cond $X=3.13 $Y=0 $X2=4.08
+ $Y2=0
r90 42 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.33 $Y=0 $X2=4.495
+ $Y2=0
r91 42 45 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=4.33 $Y=0 $X2=4.08
+ $Y2=0
r92 41 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r93 40 41 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r94 37 41 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=0.24 $Y=0 $X2=2.64
+ $Y2=0
r95 36 40 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=2.64
+ $Y2=0
r96 36 37 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r97 34 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.8 $Y=0 $X2=2.965
+ $Y2=0
r98 34 40 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=2.8 $Y=0 $X2=2.64
+ $Y2=0
r99 32 46 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.36 $Y=0 $X2=4.08
+ $Y2=0
r100 32 57 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.36 $Y=0
+ $X2=3.12 $Y2=0
r101 30 49 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=5.26 $Y=0 $X2=5.04
+ $Y2=0
r102 30 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.26 $Y=0 $X2=5.425
+ $Y2=0
r103 29 53 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=5.59 $Y=0 $X2=6
+ $Y2=0
r104 29 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.59 $Y=0 $X2=5.425
+ $Y2=0
r105 25 62 3.21509 $w=2.6e-07 $l=1.36015e-07 $layer=LI1_cond $X=6.39 $Y=0.085
+ $X2=6.49 $Y2=0
r106 25 27 19.0596 $w=2.58e-07 $l=4.3e-07 $layer=LI1_cond $X=6.39 $Y=0.085
+ $X2=6.39 $Y2=0.515
r107 21 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.425 $Y=0.085
+ $X2=5.425 $Y2=0
r108 21 23 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=5.425 $Y=0.085
+ $X2=5.425 $Y2=0.625
r109 17 59 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.495 $Y=0.085
+ $X2=4.495 $Y2=0
r110 17 19 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=4.495 $Y=0.085
+ $X2=4.495 $Y2=0.515
r111 13 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.965 $Y=0.085
+ $X2=2.965 $Y2=0
r112 13 15 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=2.965 $Y=0.085
+ $X2=2.965 $Y2=0.535
r113 4 27 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=6.215
+ $Y=0.37 $X2=6.355 $Y2=0.515
r114 3 23 182 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=1 $X=5.285
+ $Y=0.37 $X2=5.425 $Y2=0.625
r115 2 19 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=4.35
+ $Y=0.37 $X2=4.495 $Y2=0.515
r116 1 15 182 $w=1.7e-07 $l=2.48193e-07 $layer=licon1_NDIFF $count=1 $X=2.745
+ $Y=0.595 $X2=2.965 $Y2=0.535
.ends

