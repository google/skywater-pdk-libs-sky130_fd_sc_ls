* File: sky130_fd_sc_ls__sdfrtp_1.spice
* Created: Fri Aug 28 14:03:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__sdfrtp_1.pex.spice"
.subckt sky130_fd_sc_ls__sdfrtp_1  VNB VPB SCE D SCD CLK RESET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* RESET_B	RESET_B
* CLK	CLK
* SCD	SCD
* D	D
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1033 N_VGND_M1033_d N_SCE_M1033_g N_A_27_88#_M1033_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.1197 PD=1.41 PS=1.41 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1005 noxref_25 N_A_27_88#_M1005_g N_noxref_24_M1005_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.2 A=0.063 P=1.14 MULT=1
MM1006 N_A_300_464#_M1006_d N_D_M1006_g noxref_25 VNB NSHORT L=0.15 W=0.42
+ AD=0.13125 AS=0.0504 PD=1.045 PS=0.66 NRD=98.568 NRS=18.564 M=1 R=2.8
+ SA=75000.6 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1024 noxref_26 N_SCE_M1024_g N_A_300_464#_M1006_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.13125 PD=0.66 PS=1.045 NRD=18.564 NRS=0 M=1 R=2.8 SA=75001.4
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1012 N_noxref_24_M1012_d N_SCD_M1012_g noxref_26 VNB NSHORT L=0.15 W=0.42
+ AD=0.0651 AS=0.0504 PD=0.73 PS=0.66 NRD=2.856 NRS=18.564 M=1 R=2.8 SA=75001.8
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1037 N_VGND_M1037_d N_RESET_B_M1037_g N_noxref_24_M1012_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1197 AS=0.0651 PD=1.41 PS=0.73 NRD=0 NRS=5.712 M=1 R=2.8
+ SA=75002.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1028 N_VGND_M1028_d N_CLK_M1028_g N_A_835_98#_M1028_s VNB NSHORT L=0.15 W=0.74
+ AD=0.161125 AS=0.2619 PD=1.245 PS=2.38 NRD=10.536 NRS=10.536 M=1 R=4.93333
+ SA=75000.2 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1032 N_A_1034_392#_M1032_d N_A_835_98#_M1032_g N_VGND_M1028_d VNB NSHORT
+ L=0.15 W=0.74 AD=0.1961 AS=0.161125 PD=2.01 PS=1.245 NRD=0 NRS=10.536 M=1
+ R=4.93333 SA=75000.8 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1035 N_A_1234_119#_M1035_d N_A_835_98#_M1035_g N_A_300_464#_M1035_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75003.8 A=0.063 P=1.14 MULT=1
MM1000 A_1320_119# N_A_1034_392#_M1000_g N_A_1234_119#_M1035_d VNB NSHORT L=0.15
+ W=0.42 AD=0.04935 AS=0.0588 PD=0.655 PS=0.7 NRD=17.856 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75003.4 A=0.063 P=1.14 MULT=1
MM1019 A_1397_119# N_A_1367_93#_M1019_g A_1320_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.04935 PD=0.66 PS=0.655 NRD=18.564 NRS=17.856 M=1 R=2.8 SA=75001
+ SB=75003 A=0.063 P=1.14 MULT=1
MM1007 N_VGND_M1007_d N_RESET_B_M1007_g A_1397_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.211634 AS=0.0504 PD=1.27189 PS=0.66 NRD=128.244 NRS=18.564 M=1 R=2.8
+ SA=75001.4 SB=75002.6 A=0.063 P=1.14 MULT=1
MM1031 N_A_1367_93#_M1031_d N_A_1234_119#_M1031_g N_VGND_M1007_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.0896 AS=0.322491 PD=0.92 PS=1.93811 NRD=0 NRS=84.156 M=1
+ R=4.26667 SA=75001.7 SB=75002.1 A=0.096 P=1.58 MULT=1
MM1003 N_A_1745_74#_M1003_d N_A_1034_392#_M1003_g N_A_1367_93#_M1031_d VNB
+ NSHORT L=0.15 W=0.64 AD=0.282989 AS=0.0896 PD=1.96226 PS=0.92 NRD=132.18 NRS=0
+ M=1 R=4.26667 SA=75002.1 SB=75001.7 A=0.096 P=1.58 MULT=1
MM1002 A_1972_74# N_A_835_98#_M1002_g N_A_1745_74#_M1003_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.185711 PD=0.63 PS=1.28774 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75003 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_A_1997_272#_M1001_g A_1972_74# VNB NSHORT L=0.15 W=0.42
+ AD=0.06405 AS=0.0441 PD=0.725 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75003.3
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1036 A_2135_74# N_RESET_B_M1036_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.06405 PD=0.63 PS=0.725 NRD=14.28 NRS=7.14 M=1 R=2.8 SA=75003.8
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1021 N_A_1997_272#_M1021_d N_A_1745_74#_M1021_g A_2135_74# VNB NSHORT L=0.15
+ W=0.42 AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8
+ SA=75004.1 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1025 N_A_2399_424#_M1025_d N_A_1745_74#_M1025_g N_VGND_M1025_s VNB NSHORT
+ L=0.15 W=0.55 AD=0.15675 AS=0.1595 PD=1.67 PS=1.68 NRD=0 NRS=1.08 M=1
+ R=3.66667 SA=75000.2 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1004 N_Q_M1004_d N_A_2399_424#_M1004_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.2109 PD=2.05 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1020 N_VPWR_M1020_d N_SCE_M1020_g N_A_27_88#_M1020_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.112 AS=0.1888 PD=0.99 PS=1.87 NRD=18.4589 NRS=3.0732 M=1 R=4.26667
+ SA=75000.2 SB=75003.3 A=0.096 P=1.58 MULT=1
MM1017 A_216_464# N_SCE_M1017_g N_VPWR_M1020_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0864 AS=0.112 PD=0.91 PS=0.99 NRD=24.625 NRS=3.0732 M=1 R=4.26667
+ SA=75000.7 SB=75002.8 A=0.096 P=1.58 MULT=1
MM1011 N_A_300_464#_M1011_d N_D_M1011_g A_216_464# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.328 AS=0.0864 PD=1.665 PS=0.91 NRD=3.0732 NRS=24.625 M=1 R=4.26667
+ SA=75001.1 SB=75002.4 A=0.096 P=1.58 MULT=1
MM1022 A_535_464# N_A_27_88#_M1022_g N_A_300_464#_M1011_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0912 AS=0.328 PD=0.925 PS=1.665 NRD=26.9299 NRS=0 M=1 R=4.26667
+ SA=75002.3 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1026 N_VPWR_M1026_d N_SCD_M1026_g A_535_464# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1344 AS=0.0912 PD=1.06 PS=0.925 NRD=3.0732 NRS=26.9299 M=1 R=4.26667
+ SA=75002.8 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1038 N_A_300_464#_M1038_d N_RESET_B_M1038_g N_VPWR_M1026_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1888 AS=0.1344 PD=1.87 PS=1.06 NRD=3.0732 NRS=40.0107 M=1
+ R=4.26667 SA=75003.3 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1027 N_VPWR_M1027_d N_CLK_M1027_g N_A_835_98#_M1027_s VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.295 PD=1.3 PS=2.59 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75000.2
+ SB=75000.7 A=0.15 P=2.3 MULT=1
MM1030 N_A_1034_392#_M1030_d N_A_835_98#_M1030_g N_VPWR_M1027_d VPB PHIGHVT
+ L=0.15 W=1 AD=0.295 AS=0.15 PD=2.59 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75000.7 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1039 N_A_1234_119#_M1039_d N_A_1034_392#_M1039_g N_A_300_464#_M1039_s VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.0763 AS=0.1239 PD=0.795 PS=1.43 NRD=30.4759
+ NRS=4.6886 M=1 R=2.8 SA=75000.2 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1029 A_1343_461# N_A_835_98#_M1029_g N_A_1234_119#_M1039_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0567 AS=0.0763 PD=0.69 PS=0.795 NRD=37.5088 NRS=4.6886 M=1 R=2.8
+ SA=75000.7 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1008 N_VPWR_M1008_d N_A_1367_93#_M1008_g A_1343_461# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.135887 AS=0.0567 PD=1.14 PS=0.69 NRD=125.942 NRS=37.5088 M=1 R=2.8
+ SA=75001.1 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1009 N_A_1234_119#_M1009_d N_RESET_B_M1009_g N_VPWR_M1008_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1239 AS=0.135887 PD=1.43 PS=1.14 NRD=4.6886 NRS=125.942 M=1 R=2.8
+ SA=75001.7 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1013 N_A_1367_93#_M1013_d N_A_1234_119#_M1013_g N_VPWR_M1013_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.15 AS=0.295 PD=1.3 PS=2.59 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75001.2 A=0.15 P=2.3 MULT=1
MM1018 N_A_1745_74#_M1018_d N_A_835_98#_M1018_g N_A_1367_93#_M1013_d VPB PHIGHVT
+ L=0.15 W=1 AD=0.311954 AS=0.15 PD=2.56338 PS=1.3 NRD=40.3653 NRS=1.9503 M=1
+ R=6.66667 SA=75000.7 SB=75000.7 A=0.15 P=2.3 MULT=1
MM1014 A_1993_508# N_A_1034_392#_M1014_g N_A_1745_74#_M1018_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0567 AS=0.131021 PD=0.69 PS=1.07662 NRD=37.5088 NRS=53.9386 M=1
+ R=2.8 SA=75000.9 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1034 N_VPWR_M1034_d N_A_1997_272#_M1034_g A_1993_508# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.08925 AS=0.0567 PD=0.845 PS=0.69 NRD=21.0987 NRS=37.5088 M=1 R=2.8
+ SA=75001.3 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1016 N_A_1997_272#_M1016_d N_RESET_B_M1016_g N_VPWR_M1034_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.063 AS=0.08925 PD=0.72 PS=0.845 NRD=4.6886 NRS=46.886 M=1 R=2.8
+ SA=75001.9 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1023 N_VPWR_M1023_d N_A_1745_74#_M1023_g N_A_1997_272#_M1016_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.1092 AS=0.063 PD=0.85 PS=0.72 NRD=44.5417 NRS=4.6886 M=1
+ R=2.8 SA=75002.3 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1010 N_A_2399_424#_M1010_d N_A_1745_74#_M1010_g N_VPWR_M1023_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.2478 AS=0.2184 PD=2.27 PS=1.7 NRD=2.3443 NRS=14.0658 M=1
+ R=5.6 SA=75001.6 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1015 N_Q_M1015_d N_A_2399_424#_M1015_g N_VPWR_M1015_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.3304 AS=0.3304 PD=2.83 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.2 A=0.168 P=2.54 MULT=1
DX40_noxref VNB VPB NWDIODE A=25.8429 P=31.6
c_157 VNB 0 1.61901e-19 $X=0 $Y=0
c_2213 A_1343_461# 0 1.84284e-19 $X=6.715 $Y=2.305
c_2215 A_1993_508# 0 1.05093e-19 $X=9.965 $Y=2.54
*
.include "sky130_fd_sc_ls__sdfrtp_1.pxi.spice"
*
.ends
*
*
