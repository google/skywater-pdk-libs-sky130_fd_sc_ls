* File: sky130_fd_sc_ls__fa_1.pxi.spice
* Created: Wed Sep  2 11:07:31 2020
* 
x_PM_SKY130_FD_SC_LS__FA_1%A_69_260# N_A_69_260#_M1026_d N_A_69_260#_M1000_d
+ N_A_69_260#_M1024_g N_A_69_260#_c_158_n N_A_69_260#_M1021_g
+ N_A_69_260#_c_159_n N_A_69_260#_c_170_p N_A_69_260#_c_244_p
+ N_A_69_260#_c_163_n N_A_69_260#_c_172_p N_A_69_260#_c_164_n
+ N_A_69_260#_c_160_n N_A_69_260#_c_166_n N_A_69_260#_c_161_n
+ N_A_69_260#_c_182_p PM_SKY130_FD_SC_LS__FA_1%A_69_260#
x_PM_SKY130_FD_SC_LS__FA_1%A N_A_c_257_n N_A_M1011_g N_A_M1008_g N_A_c_259_n
+ N_A_M1015_g N_A_c_260_n N_A_M1003_g N_A_c_261_n N_A_M1009_g N_A_c_262_n
+ N_A_M1027_g N_A_c_263_n N_A_M1022_g N_A_c_264_n N_A_c_265_n N_A_M1018_g
+ N_A_c_266_n N_A_c_267_n N_A_c_268_n N_A_c_269_n N_A_c_270_n N_A_c_271_n
+ N_A_c_435_p N_A_c_310_p N_A_c_272_n A PM_SKY130_FD_SC_LS__FA_1%A
x_PM_SKY130_FD_SC_LS__FA_1%CIN N_CIN_M1026_g N_CIN_c_473_n N_CIN_M1000_g
+ N_CIN_M1002_g N_CIN_c_475_n N_CIN_M1007_g N_CIN_M1020_g N_CIN_c_477_n
+ N_CIN_M1014_g N_CIN_c_478_n N_CIN_c_479_n N_CIN_c_489_n N_CIN_c_490_n
+ N_CIN_c_491_n N_CIN_c_480_n N_CIN_c_481_n N_CIN_c_482_n CIN N_CIN_c_483_n
+ PM_SKY130_FD_SC_LS__FA_1%CIN
x_PM_SKY130_FD_SC_LS__FA_1%A_465_249# N_A_465_249#_M1016_d N_A_465_249#_M1010_d
+ N_A_465_249#_M1004_g N_A_465_249#_c_642_n N_A_465_249#_M1006_g
+ N_A_465_249#_c_651_n N_A_465_249#_M1023_g N_A_465_249#_M1017_g
+ N_A_465_249#_c_643_n N_A_465_249#_c_644_n N_A_465_249#_c_653_n
+ N_A_465_249#_c_668_n N_A_465_249#_c_654_n N_A_465_249#_c_661_n
+ N_A_465_249#_c_674_n N_A_465_249#_c_655_n N_A_465_249#_c_682_n
+ N_A_465_249#_c_645_n N_A_465_249#_c_646_n N_A_465_249#_c_647_n
+ N_A_465_249#_c_648_n N_A_465_249#_c_649_n N_A_465_249#_c_699_n
+ PM_SKY130_FD_SC_LS__FA_1%A_465_249#
x_PM_SKY130_FD_SC_LS__FA_1%B N_B_M1025_g N_B_M1005_g N_B_c_836_n N_B_c_837_n
+ N_B_M1012_g N_B_c_825_n N_B_c_826_n N_B_c_839_n N_B_c_840_n N_B_c_841_n
+ N_B_M1019_g N_B_c_843_n N_B_M1016_g N_B_c_827_n N_B_c_828_n N_B_c_845_n
+ N_B_c_846_n N_B_c_847_n N_B_M1010_g N_B_c_849_n N_B_M1001_g N_B_M1013_g
+ N_B_c_851_n N_B_c_830_n N_B_c_852_n N_B_c_831_n N_B_c_853_n N_B_c_854_n B
+ N_B_c_832_n N_B_c_833_n PM_SKY130_FD_SC_LS__FA_1%B
x_PM_SKY130_FD_SC_LS__FA_1%SUM N_SUM_M1024_s N_SUM_M1021_s N_SUM_c_1001_n
+ N_SUM_c_1002_n N_SUM_c_998_n SUM SUM SUM PM_SKY130_FD_SC_LS__FA_1%SUM
x_PM_SKY130_FD_SC_LS__FA_1%VPWR N_VPWR_M1021_d N_VPWR_M1019_d N_VPWR_M1007_d
+ N_VPWR_M1022_d N_VPWR_M1023_s N_VPWR_c_1019_n N_VPWR_c_1020_n N_VPWR_c_1021_n
+ N_VPWR_c_1022_n N_VPWR_c_1023_n N_VPWR_c_1024_n N_VPWR_c_1025_n VPWR
+ N_VPWR_c_1026_n N_VPWR_c_1027_n N_VPWR_c_1028_n N_VPWR_c_1029_n
+ N_VPWR_c_1030_n N_VPWR_c_1018_n N_VPWR_c_1032_n N_VPWR_c_1033_n
+ N_VPWR_c_1034_n N_VPWR_c_1035_n PM_SKY130_FD_SC_LS__FA_1%VPWR
x_PM_SKY130_FD_SC_LS__FA_1%A_509_347# N_A_509_347#_M1006_d N_A_509_347#_M1003_d
+ N_A_509_347#_c_1134_n N_A_509_347#_c_1132_n N_A_509_347#_c_1137_n
+ N_A_509_347#_c_1136_n N_A_509_347#_c_1133_n
+ PM_SKY130_FD_SC_LS__FA_1%A_509_347#
x_PM_SKY130_FD_SC_LS__FA_1%A_1107_347# N_A_1107_347#_M1014_d
+ N_A_1107_347#_M1001_d N_A_1107_347#_c_1179_n N_A_1107_347#_c_1174_n
+ N_A_1107_347#_c_1178_n N_A_1107_347#_c_1175_n N_A_1107_347#_c_1176_n
+ PM_SKY130_FD_SC_LS__FA_1%A_1107_347#
x_PM_SKY130_FD_SC_LS__FA_1%COUT N_COUT_M1017_d N_COUT_M1023_d COUT COUT COUT
+ COUT COUT COUT COUT COUT PM_SKY130_FD_SC_LS__FA_1%COUT
x_PM_SKY130_FD_SC_LS__FA_1%VGND N_VGND_M1024_d N_VGND_M1012_d N_VGND_M1002_d
+ N_VGND_M1018_d N_VGND_M1017_s N_VGND_c_1220_n N_VGND_c_1221_n N_VGND_c_1222_n
+ N_VGND_c_1223_n VGND N_VGND_c_1224_n N_VGND_c_1225_n N_VGND_c_1226_n
+ N_VGND_c_1227_n N_VGND_c_1228_n N_VGND_c_1229_n N_VGND_c_1230_n
+ N_VGND_c_1231_n N_VGND_c_1232_n N_VGND_c_1233_n PM_SKY130_FD_SC_LS__FA_1%VGND
x_PM_SKY130_FD_SC_LS__FA_1%A_501_75# N_A_501_75#_M1004_d N_A_501_75#_M1015_d
+ N_A_501_75#_c_1335_n N_A_501_75#_c_1332_n N_A_501_75#_c_1340_n
+ PM_SKY130_FD_SC_LS__FA_1%A_501_75#
x_PM_SKY130_FD_SC_LS__FA_1%A_1100_75# N_A_1100_75#_M1020_d N_A_1100_75#_M1013_d
+ N_A_1100_75#_c_1359_n N_A_1100_75#_c_1364_n N_A_1100_75#_c_1374_n
+ N_A_1100_75#_c_1365_n N_A_1100_75#_c_1360_n
+ PM_SKY130_FD_SC_LS__FA_1%A_1100_75#
cc_1 VNB N_A_69_260#_M1024_g 0.0264069f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_A_69_260#_c_158_n 0.0361844f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.765
cc_3 VNB N_A_69_260#_c_159_n 0.00139797f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.3
cc_4 VNB N_A_69_260#_c_160_n 0.00272515f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.465
cc_5 VNB N_A_69_260#_c_161_n 0.00289452f $X=-0.19 $Y=-0.245 $X2=2.105 $Y2=0.55
cc_6 VNB N_A_c_257_n 0.0341217f $X=-0.19 $Y=-0.245 $X2=1.965 $Y2=0.375
cc_7 VNB N_A_M1008_g 0.0233458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_c_259_n 0.0178818f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_9 VNB N_A_c_260_n 0.0386731f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.765
cc_10 VNB N_A_c_261_n 0.0382416f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=0.75
cc_11 VNB N_A_c_262_n 0.0170005f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=0.665
cc_12 VNB N_A_c_263_n 0.0375768f $X=-0.19 $Y=-0.245 $X2=2.08 $Y2=2.035
cc_13 VNB N_A_c_264_n 0.0254757f $X=-0.19 $Y=-0.245 $X2=2.245 $Y2=2.59
cc_14 VNB N_A_c_265_n 0.019979f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_c_266_n 0.0201195f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.465
cc_16 VNB N_A_c_267_n 0.00239261f $X=-0.19 $Y=-0.245 $X2=1.14 $Y2=2.035
cc_17 VNB N_A_c_268_n 0.00740945f $X=-0.19 $Y=-0.245 $X2=2.105 $Y2=0.55
cc_18 VNB N_A_c_269_n 0.00963516f $X=-0.19 $Y=-0.245 $X2=2.105 $Y2=0.665
cc_19 VNB N_A_c_270_n 0.00224455f $X=-0.19 $Y=-0.245 $X2=2.245 $Y2=1.91
cc_20 VNB N_A_c_271_n 0.00811052f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_c_272_n 0.00338796f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB A 0.00205822f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_CIN_M1026_g 0.0243526f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_CIN_c_473_n 0.0219431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_CIN_M1002_g 0.0252727f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_CIN_c_475_n 0.0239237f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_27 VNB N_CIN_M1020_g 0.025655f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=0.665
cc_28 VNB N_CIN_c_477_n 0.0223488f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=1.795
cc_29 VNB N_CIN_c_478_n 0.00103036f $X=-0.19 $Y=-0.245 $X2=2.245 $Y2=2.12
cc_30 VNB N_CIN_c_479_n 0.00370463f $X=-0.19 $Y=-0.245 $X2=2.245 $Y2=2.59
cc_31 VNB N_CIN_c_480_n 3.94034e-19 $X=-0.19 $Y=-0.245 $X2=1.14 $Y2=1.795
cc_32 VNB N_CIN_c_481_n 0.00392612f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_CIN_c_482_n 3.29665e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_CIN_c_483_n 0.00255009f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_465_249#_M1004_g 0.0261075f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_36 VNB N_A_465_249#_c_642_n 0.0217642f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.765
cc_37 VNB N_A_465_249#_c_643_n 0.0622009f $X=-0.19 $Y=-0.245 $X2=1.225 $Y2=2.035
cc_38 VNB N_A_465_249#_c_644_n 0.0221372f $X=-0.19 $Y=-0.245 $X2=2.245 $Y2=2.12
cc_39 VNB N_A_465_249#_c_645_n 0.0050609f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_465_249#_c_646_n 0.029447f $X=-0.19 $Y=-0.245 $X2=2.245 $Y2=1.91
cc_41 VNB N_A_465_249#_c_647_n 7.33795e-19 $X=-0.19 $Y=-0.245 $X2=2.245 $Y2=1.91
cc_42 VNB N_A_465_249#_c_648_n 0.00629526f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.465
cc_43 VNB N_A_465_249#_c_649_n 0.00566251f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_B_M1025_g 0.0387714f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_B_c_825_n 0.00627038f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=0.75
cc_46 VNB N_B_c_826_n 0.020951f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.3
cc_47 VNB N_B_c_827_n 0.00553036f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.465
cc_48 VNB N_B_c_828_n 0.0181796f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.465
cc_49 VNB N_B_M1013_g 0.0350093f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.465
cc_50 VNB N_B_c_830_n 0.0168615f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_B_c_831_n 0.014923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_B_c_832_n 0.0426944f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_B_c_833_n 0.00483187f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_SUM_c_998_n 0.0246106f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.3
cc_55 VNB SUM 0.0271795f $X=-0.19 $Y=-0.245 $X2=1.94 $Y2=0.665
cc_56 VNB SUM 0.0094822f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=0.665
cc_57 VNB N_VPWR_c_1018_n 0.362705f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB COUT 0.0263294f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.3
cc_59 VNB COUT 0.00845976f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_60 VNB COUT 0.0269902f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_61 VNB N_VGND_c_1220_n 0.018469f $X=-0.19 $Y=-0.245 $X2=1.94 $Y2=0.665
cc_62 VNB N_VGND_c_1221_n 0.00826643f $X=-0.19 $Y=-0.245 $X2=2.08 $Y2=2.035
cc_63 VNB N_VGND_c_1222_n 0.00547714f $X=-0.19 $Y=-0.245 $X2=2.245 $Y2=2.59
cc_64 VNB N_VGND_c_1223_n 0.0139843f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.465
cc_65 VNB N_VGND_c_1224_n 0.0343344f $X=-0.19 $Y=-0.245 $X2=1.14 $Y2=2.035
cc_66 VNB N_VGND_c_1225_n 0.0555224f $X=-0.19 $Y=-0.245 $X2=2.105 $Y2=0.665
cc_67 VNB N_VGND_c_1226_n 0.0578707f $X=-0.19 $Y=-0.245 $X2=2.245 $Y2=2.035
cc_68 VNB N_VGND_c_1227_n 0.019427f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_1228_n 0.0189924f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_1229_n 0.467822f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1230_n 0.0144116f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1231_n 0.00898487f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1232_n 0.00477762f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1233_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_1100_75#_c_1359_n 0.00362777f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.3
cc_76 VNB N_A_1100_75#_c_1360_n 0.00389169f $X=-0.19 $Y=-0.245 $X2=1.94
+ $Y2=0.665
cc_77 VPB N_A_69_260#_c_158_n 0.0273992f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.765
cc_78 VPB N_A_69_260#_c_163_n 0.00635828f $X=-0.19 $Y=1.66 $X2=1.055 $Y2=1.795
cc_79 VPB N_A_69_260#_c_164_n 0.0024405f $X=-0.19 $Y=1.66 $X2=2.245 $Y2=2.59
cc_80 VPB N_A_69_260#_c_160_n 4.96285e-19 $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.465
cc_81 VPB N_A_69_260#_c_166_n 0.00188689f $X=-0.19 $Y=1.66 $X2=1.14 $Y2=1.795
cc_82 VPB N_A_c_257_n 0.0220687f $X=-0.19 $Y=1.66 $X2=1.965 $Y2=0.375
cc_83 VPB N_A_c_260_n 0.021126f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.765
cc_84 VPB N_A_c_261_n 0.0192323f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=0.75
cc_85 VPB N_A_c_263_n 0.0279938f $X=-0.19 $Y=1.66 $X2=2.08 $Y2=2.035
cc_86 VPB N_A_c_272_n 9.06676e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_CIN_c_473_n 0.0242431f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_CIN_c_475_n 0.0230489f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_89 VPB N_CIN_c_477_n 0.0255466f $X=-0.19 $Y=1.66 $X2=0.705 $Y2=1.795
cc_90 VPB N_CIN_c_478_n 0.00300344f $X=-0.19 $Y=1.66 $X2=2.245 $Y2=2.12
cc_91 VPB N_CIN_c_479_n 0.00190949f $X=-0.19 $Y=1.66 $X2=2.245 $Y2=2.59
cc_92 VPB N_CIN_c_489_n 0.0102933f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.465
cc_93 VPB N_CIN_c_490_n 9.44822e-19 $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.465
cc_94 VPB N_CIN_c_491_n 0.00462727f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=1.795
cc_95 VPB N_CIN_c_480_n 6.01613e-19 $X=-0.19 $Y=1.66 $X2=1.14 $Y2=1.795
cc_96 VPB N_CIN_c_481_n 0.00371448f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_CIN_c_482_n 0.00316307f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_CIN_c_483_n 0.00392455f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB N_A_465_249#_c_642_n 0.0238795f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.765
cc_100 VPB N_A_465_249#_c_651_n 0.0218984f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=0.75
cc_101 VPB N_A_465_249#_c_643_n 0.00867073f $X=-0.19 $Y=1.66 $X2=1.225 $Y2=2.035
cc_102 VPB N_A_465_249#_c_653_n 0.00322579f $X=-0.19 $Y=1.66 $X2=2.245 $Y2=2.59
cc_103 VPB N_A_465_249#_c_654_n 0.00278199f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.465
cc_104 VPB N_A_465_249#_c_655_n 9.96124e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_105 VPB N_A_465_249#_c_645_n 0.00418629f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_A_465_249#_c_649_n 0.00348732f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB N_B_M1025_g 0.00521426f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_B_M1005_g 0.0110311f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_109 VPB N_B_c_836_n 0.100041f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_110 VPB N_B_c_837_n 0.0208605f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_B_c_826_n 8.27112e-19 $X=-0.19 $Y=1.66 $X2=0.62 $Y2=1.3
cc_112 VPB N_B_c_839_n 0.00742498f $X=-0.19 $Y=1.66 $X2=1.94 $Y2=0.665
cc_113 VPB N_B_c_840_n 0.0153402f $X=-0.19 $Y=1.66 $X2=0.705 $Y2=0.665
cc_114 VPB N_B_c_841_n 0.00574672f $X=-0.19 $Y=1.66 $X2=1.055 $Y2=1.795
cc_115 VPB N_B_M1019_g 0.00813881f $X=-0.19 $Y=1.66 $X2=1.225 $Y2=2.035
cc_116 VPB N_B_c_843_n 0.136579f $X=-0.19 $Y=1.66 $X2=2.245 $Y2=2.12
cc_117 VPB N_B_c_828_n 6.27797e-19 $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.465
cc_118 VPB N_B_c_845_n 0.00752662f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=1.795
cc_119 VPB N_B_c_846_n 0.016528f $X=-0.19 $Y=1.66 $X2=1.14 $Y2=1.795
cc_120 VPB N_B_c_847_n 0.00510734f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_B_M1010_g 0.00751154f $X=-0.19 $Y=1.66 $X2=2.105 $Y2=0.55
cc_122 VPB N_B_c_849_n 0.121778f $X=-0.19 $Y=1.66 $X2=2.105 $Y2=0.55
cc_123 VPB N_B_M1001_g 0.0117459f $X=-0.19 $Y=1.66 $X2=2.245 $Y2=1.91
cc_124 VPB N_B_c_851_n 0.0097805f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_B_c_852_n 0.0089864f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 VPB N_B_c_853_n 0.0089864f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_127 VPB N_B_c_854_n 0.0332515f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_B_c_832_n 0.0338556f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_129 VPB N_B_c_833_n 0.0118397f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_SUM_c_1001_n 0.00920368f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_131 VPB N_SUM_c_1002_n 0.0416756f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.765
cc_132 VPB N_SUM_c_998_n 0.00751766f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=1.3
cc_133 VPB N_VPWR_c_1019_n 0.00854695f $X=-0.19 $Y=1.66 $X2=1.055 $Y2=1.795
cc_134 VPB N_VPWR_c_1020_n 0.0132078f $X=-0.19 $Y=1.66 $X2=2.245 $Y2=2.59
cc_135 VPB N_VPWR_c_1021_n 0.0111988f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.465
cc_136 VPB N_VPWR_c_1022_n 0.0100542f $X=-0.19 $Y=1.66 $X2=1.14 $Y2=2.035
cc_137 VPB N_VPWR_c_1023_n 0.0352379f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_1024_n 0.0183142f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_1025_n 0.00436868f $X=-0.19 $Y=1.66 $X2=2.245 $Y2=2.035
cc_140 VPB N_VPWR_c_1026_n 0.0175529f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_1027_n 0.0658504f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_142 VPB N_VPWR_c_1028_n 0.0479018f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_143 VPB N_VPWR_c_1029_n 0.0266344f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_144 VPB N_VPWR_c_1030_n 0.0176701f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_145 VPB N_VPWR_c_1018_n 0.0941318f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_146 VPB N_VPWR_c_1032_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_147 VPB N_VPWR_c_1033_n 0.00436868f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_148 VPB N_VPWR_c_1034_n 0.00936252f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_149 VPB N_VPWR_c_1035_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_150 VPB N_A_509_347#_c_1132_n 0.00244184f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_151 VPB N_A_509_347#_c_1133_n 0.00274215f $X=-0.19 $Y=1.66 $X2=1.055
+ $Y2=1.795
cc_152 VPB N_A_1107_347#_c_1174_n 0.00272816f $X=-0.19 $Y=1.66 $X2=0.495
+ $Y2=0.74
cc_153 VPB N_A_1107_347#_c_1175_n 0.0045747f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_154 VPB N_A_1107_347#_c_1176_n 0.0120924f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=1.3
cc_155 VPB COUT 0.0548874f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_156 N_A_69_260#_M1024_g N_A_c_257_n 0.00308693f $X=0.495 $Y=0.74 $X2=-0.19
+ $Y2=-0.245
cc_157 N_A_69_260#_c_158_n N_A_c_257_n 0.042857f $X=0.495 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_158 N_A_69_260#_c_159_n N_A_c_257_n 2.60105e-19 $X=0.62 $Y=1.3 $X2=-0.19
+ $Y2=-0.245
cc_159 N_A_69_260#_c_170_p N_A_c_257_n 6.48432e-19 $X=1.94 $Y=0.665 $X2=-0.19
+ $Y2=-0.245
cc_160 N_A_69_260#_c_163_n N_A_c_257_n 0.0130079f $X=1.055 $Y=1.795 $X2=-0.19
+ $Y2=-0.245
cc_161 N_A_69_260#_c_172_p N_A_c_257_n 2.37377e-19 $X=2.08 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_162 N_A_69_260#_c_160_n N_A_c_257_n 0.00434044f $X=0.51 $Y=1.465 $X2=-0.19
+ $Y2=-0.245
cc_163 N_A_69_260#_c_166_n N_A_c_257_n 0.0138286f $X=1.14 $Y=1.795 $X2=-0.19
+ $Y2=-0.245
cc_164 N_A_69_260#_M1024_g N_A_M1008_g 0.0205774f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_165 N_A_69_260#_c_159_n N_A_M1008_g 0.00519091f $X=0.62 $Y=1.3 $X2=0 $Y2=0
cc_166 N_A_69_260#_c_170_p N_A_M1008_g 0.0119954f $X=1.94 $Y=0.665 $X2=0 $Y2=0
cc_167 N_A_69_260#_M1026_d N_A_c_266_n 0.00388826f $X=1.965 $Y=0.375 $X2=0 $Y2=0
cc_168 N_A_69_260#_c_170_p N_A_c_266_n 0.0369432f $X=1.94 $Y=0.665 $X2=0 $Y2=0
cc_169 N_A_69_260#_c_166_n N_A_c_266_n 2.80141e-19 $X=1.14 $Y=1.795 $X2=0 $Y2=0
cc_170 N_A_69_260#_c_161_n N_A_c_266_n 0.0209854f $X=2.105 $Y=0.55 $X2=0 $Y2=0
cc_171 N_A_69_260#_c_182_p N_A_c_266_n 0.00246004f $X=2.245 $Y=1.91 $X2=0 $Y2=0
cc_172 N_A_69_260#_M1024_g N_A_c_271_n 3.94697e-19 $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_173 N_A_69_260#_c_158_n N_A_c_271_n 2.83375e-19 $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_174 N_A_69_260#_c_159_n N_A_c_271_n 0.0190885f $X=0.62 $Y=1.3 $X2=0 $Y2=0
cc_175 N_A_69_260#_c_170_p N_A_c_271_n 0.0149495f $X=1.94 $Y=0.665 $X2=0 $Y2=0
cc_176 N_A_69_260#_c_163_n N_A_c_271_n 0.0123444f $X=1.055 $Y=1.795 $X2=0 $Y2=0
cc_177 N_A_69_260#_c_160_n N_A_c_271_n 0.0181292f $X=0.51 $Y=1.465 $X2=0 $Y2=0
cc_178 N_A_69_260#_c_166_n N_A_c_271_n 0.0133509f $X=1.14 $Y=1.795 $X2=0 $Y2=0
cc_179 N_A_69_260#_c_170_p N_CIN_M1026_g 0.00835085f $X=1.94 $Y=0.665 $X2=0
+ $Y2=0
cc_180 N_A_69_260#_c_161_n N_CIN_M1026_g 0.00569455f $X=2.105 $Y=0.55 $X2=0
+ $Y2=0
cc_181 N_A_69_260#_c_172_p N_CIN_c_473_n 0.0143532f $X=2.08 $Y=2.035 $X2=0 $Y2=0
cc_182 N_A_69_260#_c_164_n N_CIN_c_473_n 0.0122375f $X=2.245 $Y=2.59 $X2=0 $Y2=0
cc_183 N_A_69_260#_c_182_p N_CIN_c_473_n 0.00449716f $X=2.245 $Y=1.91 $X2=0
+ $Y2=0
cc_184 N_A_69_260#_M1000_d N_CIN_c_489_n 0.00212817f $X=2.095 $Y=1.735 $X2=0
+ $Y2=0
cc_185 N_A_69_260#_c_172_p N_CIN_c_489_n 0.00618871f $X=2.08 $Y=2.035 $X2=0
+ $Y2=0
cc_186 N_A_69_260#_c_182_p N_CIN_c_489_n 0.0124595f $X=2.245 $Y=1.91 $X2=0 $Y2=0
cc_187 N_A_69_260#_c_172_p N_CIN_c_490_n 0.00386746f $X=2.08 $Y=2.035 $X2=0
+ $Y2=0
cc_188 N_A_69_260#_c_166_n N_CIN_c_490_n 0.00166828f $X=1.14 $Y=1.795 $X2=0
+ $Y2=0
cc_189 N_A_69_260#_c_182_p N_CIN_c_490_n 9.59784e-19 $X=2.245 $Y=1.91 $X2=0
+ $Y2=0
cc_190 N_A_69_260#_c_172_p N_CIN_c_481_n 0.0185251f $X=2.08 $Y=2.035 $X2=0 $Y2=0
cc_191 N_A_69_260#_c_166_n N_CIN_c_481_n 0.0020521f $X=1.14 $Y=1.795 $X2=0 $Y2=0
cc_192 N_A_69_260#_c_182_p N_CIN_c_481_n 0.00272215f $X=2.245 $Y=1.91 $X2=0
+ $Y2=0
cc_193 N_A_69_260#_c_161_n N_A_465_249#_M1004_g 0.00476897f $X=2.105 $Y=0.55
+ $X2=0 $Y2=0
cc_194 N_A_69_260#_c_164_n N_A_465_249#_c_642_n 0.0068733f $X=2.245 $Y=2.59
+ $X2=0 $Y2=0
cc_195 N_A_69_260#_c_182_p N_A_465_249#_c_642_n 0.0056738f $X=2.245 $Y=1.91
+ $X2=0 $Y2=0
cc_196 N_A_69_260#_c_182_p N_A_465_249#_c_661_n 4.07793e-19 $X=2.245 $Y=1.91
+ $X2=0 $Y2=0
cc_197 N_A_69_260#_c_182_p N_A_465_249#_c_649_n 0.00334589f $X=2.245 $Y=1.91
+ $X2=0 $Y2=0
cc_198 N_A_69_260#_c_170_p N_B_M1025_g 0.0107797f $X=1.94 $Y=0.665 $X2=0 $Y2=0
cc_199 N_A_69_260#_c_166_n N_B_M1025_g 0.0023803f $X=1.14 $Y=1.795 $X2=0 $Y2=0
cc_200 N_A_69_260#_c_161_n N_B_M1025_g 0.00119451f $X=2.105 $Y=0.55 $X2=0 $Y2=0
cc_201 N_A_69_260#_c_172_p N_B_M1005_g 0.0181338f $X=2.08 $Y=2.035 $X2=0 $Y2=0
cc_202 N_A_69_260#_c_166_n N_B_M1005_g 0.0018123f $X=1.14 $Y=1.795 $X2=0 $Y2=0
cc_203 N_A_69_260#_c_182_p N_B_M1005_g 0.00302095f $X=2.245 $Y=1.91 $X2=0 $Y2=0
cc_204 N_A_69_260#_c_164_n N_B_c_836_n 0.00617372f $X=2.245 $Y=2.59 $X2=0 $Y2=0
cc_205 N_A_69_260#_c_182_p N_B_M1019_g 5.73377e-19 $X=2.245 $Y=1.91 $X2=0 $Y2=0
cc_206 N_A_69_260#_c_182_p N_B_c_851_n 8.23198e-19 $X=2.245 $Y=1.91 $X2=0 $Y2=0
cc_207 N_A_69_260#_c_158_n N_SUM_c_1001_n 0.00920527f $X=0.495 $Y=1.765 $X2=0
+ $Y2=0
cc_208 N_A_69_260#_c_160_n N_SUM_c_1001_n 0.00459508f $X=0.51 $Y=1.465 $X2=0
+ $Y2=0
cc_209 N_A_69_260#_M1024_g N_SUM_c_998_n 0.0034597f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_210 N_A_69_260#_c_158_n N_SUM_c_998_n 0.0121466f $X=0.495 $Y=1.765 $X2=0
+ $Y2=0
cc_211 N_A_69_260#_c_159_n N_SUM_c_998_n 0.00833638f $X=0.62 $Y=1.3 $X2=0 $Y2=0
cc_212 N_A_69_260#_c_160_n N_SUM_c_998_n 0.0344321f $X=0.51 $Y=1.465 $X2=0 $Y2=0
cc_213 N_A_69_260#_M1024_g SUM 0.00206152f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_214 N_A_69_260#_c_158_n SUM 8.44384e-19 $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_215 N_A_69_260#_c_159_n SUM 0.0136155f $X=0.62 $Y=1.3 $X2=0 $Y2=0
cc_216 N_A_69_260#_c_163_n N_VPWR_M1021_d 0.00182839f $X=1.055 $Y=1.795
+ $X2=-0.19 $Y2=-0.245
cc_217 N_A_69_260#_c_160_n N_VPWR_M1021_d 8.63167e-19 $X=0.51 $Y=1.465 $X2=-0.19
+ $Y2=-0.245
cc_218 N_A_69_260#_c_158_n N_VPWR_c_1019_n 0.0179282f $X=0.495 $Y=1.765 $X2=0
+ $Y2=0
cc_219 N_A_69_260#_c_163_n N_VPWR_c_1019_n 0.0140386f $X=1.055 $Y=1.795 $X2=0
+ $Y2=0
cc_220 N_A_69_260#_c_160_n N_VPWR_c_1019_n 0.0081754f $X=0.51 $Y=1.465 $X2=0
+ $Y2=0
cc_221 N_A_69_260#_c_158_n N_VPWR_c_1026_n 0.00413917f $X=0.495 $Y=1.765 $X2=0
+ $Y2=0
cc_222 N_A_69_260#_c_164_n N_VPWR_c_1027_n 0.00748518f $X=2.245 $Y=2.59 $X2=0
+ $Y2=0
cc_223 N_A_69_260#_c_158_n N_VPWR_c_1018_n 0.00821187f $X=0.495 $Y=1.765 $X2=0
+ $Y2=0
cc_224 N_A_69_260#_c_164_n N_VPWR_c_1018_n 0.00906792f $X=2.245 $Y=2.59 $X2=0
+ $Y2=0
cc_225 N_A_69_260#_c_172_p A_217_368# 0.0124597f $X=2.08 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_226 N_A_69_260#_c_166_n A_217_368# 0.0052193f $X=1.14 $Y=1.795 $X2=-0.19
+ $Y2=-0.245
cc_227 N_A_69_260#_c_172_p A_318_389# 0.0116474f $X=2.08 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_228 N_A_69_260#_c_182_p N_A_509_347#_c_1134_n 0.0217246f $X=2.245 $Y=1.91
+ $X2=0 $Y2=0
cc_229 N_A_69_260#_c_164_n N_A_509_347#_c_1132_n 0.0197755f $X=2.245 $Y=2.59
+ $X2=0 $Y2=0
cc_230 N_A_69_260#_c_164_n N_A_509_347#_c_1136_n 0.0123817f $X=2.245 $Y=2.59
+ $X2=0 $Y2=0
cc_231 N_A_69_260#_c_159_n N_VGND_M1024_d 0.00449182f $X=0.62 $Y=1.3 $X2=-0.19
+ $Y2=-0.245
cc_232 N_A_69_260#_c_170_p N_VGND_M1024_d 0.011913f $X=1.94 $Y=0.665 $X2=-0.19
+ $Y2=-0.245
cc_233 N_A_69_260#_c_244_p N_VGND_M1024_d 8.19949e-19 $X=0.705 $Y=0.665
+ $X2=-0.19 $Y2=-0.245
cc_234 N_A_69_260#_M1024_g N_VGND_c_1224_n 0.00806235f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_235 N_A_69_260#_c_170_p N_VGND_c_1224_n 0.0203993f $X=1.94 $Y=0.665 $X2=0
+ $Y2=0
cc_236 N_A_69_260#_c_244_p N_VGND_c_1224_n 0.00778467f $X=0.705 $Y=0.665 $X2=0
+ $Y2=0
cc_237 N_A_69_260#_c_170_p N_VGND_c_1225_n 0.0161153f $X=1.94 $Y=0.665 $X2=0
+ $Y2=0
cc_238 N_A_69_260#_c_161_n N_VGND_c_1225_n 0.0137352f $X=2.105 $Y=0.55 $X2=0
+ $Y2=0
cc_239 N_A_69_260#_M1024_g N_VGND_c_1229_n 0.00798259f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_240 N_A_69_260#_c_170_p N_VGND_c_1229_n 0.0279046f $X=1.94 $Y=0.665 $X2=0
+ $Y2=0
cc_241 N_A_69_260#_c_244_p N_VGND_c_1229_n 0.00315983f $X=0.705 $Y=0.665 $X2=0
+ $Y2=0
cc_242 N_A_69_260#_c_161_n N_VGND_c_1229_n 0.0117469f $X=2.105 $Y=0.55 $X2=0
+ $Y2=0
cc_243 N_A_69_260#_c_170_p A_237_75# 0.00339426f $X=1.94 $Y=0.665 $X2=-0.19
+ $Y2=-0.245
cc_244 N_A_69_260#_c_170_p A_315_75# 0.00339426f $X=1.94 $Y=0.665 $X2=-0.19
+ $Y2=-0.245
cc_245 N_A_69_260#_c_161_n N_A_501_75#_c_1332_n 0.0225265f $X=2.105 $Y=0.55
+ $X2=0 $Y2=0
cc_246 N_A_c_266_n N_CIN_M1026_g 0.010684f $X=3.3 $Y=1.005 $X2=0 $Y2=0
cc_247 N_A_c_266_n N_CIN_c_473_n 0.00464221f $X=3.3 $Y=1.005 $X2=0 $Y2=0
cc_248 N_A_c_259_n N_CIN_M1002_g 0.0222612f $X=3.53 $Y=1.125 $X2=0 $Y2=0
cc_249 N_A_c_260_n N_CIN_M1002_g 0.00627512f $X=3.54 $Y=1.66 $X2=0 $Y2=0
cc_250 N_A_c_261_n N_CIN_M1002_g 0.0045952f $X=4.505 $Y=1.66 $X2=0 $Y2=0
cc_251 N_A_c_262_n N_CIN_M1002_g 0.0180648f $X=4.605 $Y=1.125 $X2=0 $Y2=0
cc_252 N_A_c_267_n N_CIN_M1002_g 0.00149115f $X=3.465 $Y=1.29 $X2=0 $Y2=0
cc_253 N_A_c_268_n N_CIN_M1002_g 0.0150364f $X=4.38 $Y=1.005 $X2=0 $Y2=0
cc_254 N_A_c_310_p N_CIN_M1002_g 3.60835e-19 $X=4.545 $Y=1.012 $X2=0 $Y2=0
cc_255 A N_CIN_M1002_g 0.00111147f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_256 N_A_c_260_n N_CIN_c_475_n 0.0577557f $X=3.54 $Y=1.66 $X2=0 $Y2=0
cc_257 N_A_c_261_n N_CIN_c_475_n 0.0575503f $X=4.505 $Y=1.66 $X2=0 $Y2=0
cc_258 N_A_c_267_n N_CIN_c_475_n 7.86199e-19 $X=3.465 $Y=1.29 $X2=0 $Y2=0
cc_259 N_A_c_268_n N_CIN_c_475_n 0.00447738f $X=4.38 $Y=1.005 $X2=0 $Y2=0
cc_260 A N_CIN_c_475_n 3.40268e-19 $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_261 N_A_c_263_n N_CIN_M1020_g 0.00372458f $X=6.055 $Y=1.66 $X2=0 $Y2=0
cc_262 N_A_c_269_n N_CIN_M1020_g 0.01214f $X=5.81 $Y=1.02 $X2=0 $Y2=0
cc_263 N_A_c_270_n N_CIN_M1020_g 0.00259916f $X=5.895 $Y=1.32 $X2=0 $Y2=0
cc_264 N_A_c_263_n N_CIN_c_477_n 0.0410229f $X=6.055 $Y=1.66 $X2=0 $Y2=0
cc_265 N_A_c_269_n N_CIN_c_477_n 0.00433975f $X=5.81 $Y=1.02 $X2=0 $Y2=0
cc_266 N_A_c_270_n N_CIN_c_477_n 7.67886e-19 $X=5.895 $Y=1.32 $X2=0 $Y2=0
cc_267 N_A_c_272_n N_CIN_c_477_n 8.83241e-19 $X=6.045 $Y=1.41 $X2=0 $Y2=0
cc_268 N_A_c_261_n N_CIN_c_478_n 0.00353964f $X=4.505 $Y=1.66 $X2=0 $Y2=0
cc_269 N_A_c_269_n N_CIN_c_478_n 0.0167049f $X=5.81 $Y=1.02 $X2=0 $Y2=0
cc_270 A N_CIN_c_478_n 0.0108937f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_271 N_A_c_263_n N_CIN_c_479_n 3.27165e-19 $X=6.055 $Y=1.66 $X2=0 $Y2=0
cc_272 N_A_c_269_n N_CIN_c_479_n 0.0361598f $X=5.81 $Y=1.02 $X2=0 $Y2=0
cc_273 N_A_c_270_n N_CIN_c_479_n 0.00342339f $X=5.895 $Y=1.32 $X2=0 $Y2=0
cc_274 N_A_c_272_n N_CIN_c_479_n 0.0211108f $X=6.045 $Y=1.41 $X2=0 $Y2=0
cc_275 N_A_c_260_n N_CIN_c_489_n 0.00648335f $X=3.54 $Y=1.66 $X2=0 $Y2=0
cc_276 N_A_c_266_n N_CIN_c_489_n 0.0178463f $X=3.3 $Y=1.005 $X2=0 $Y2=0
cc_277 N_A_c_267_n N_CIN_c_489_n 0.00969257f $X=3.465 $Y=1.29 $X2=0 $Y2=0
cc_278 N_A_c_268_n N_CIN_c_489_n 0.00728431f $X=4.38 $Y=1.005 $X2=0 $Y2=0
cc_279 N_A_c_257_n N_CIN_c_490_n 7.71179e-19 $X=1.01 $Y=1.765 $X2=0 $Y2=0
cc_280 N_A_c_266_n N_CIN_c_490_n 0.00192258f $X=3.3 $Y=1.005 $X2=0 $Y2=0
cc_281 N_A_c_261_n N_CIN_c_491_n 0.00613522f $X=4.505 $Y=1.66 $X2=0 $Y2=0
cc_282 N_A_c_268_n N_CIN_c_491_n 0.00507703f $X=4.38 $Y=1.005 $X2=0 $Y2=0
cc_283 N_A_c_269_n N_CIN_c_491_n 0.00614904f $X=5.81 $Y=1.02 $X2=0 $Y2=0
cc_284 A N_CIN_c_491_n 0.00968886f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_285 N_A_c_261_n N_CIN_c_480_n 0.00135296f $X=4.505 $Y=1.66 $X2=0 $Y2=0
cc_286 N_A_c_268_n N_CIN_c_480_n 0.0021404f $X=4.38 $Y=1.005 $X2=0 $Y2=0
cc_287 N_A_c_257_n N_CIN_c_481_n 0.00169765f $X=1.01 $Y=1.765 $X2=0 $Y2=0
cc_288 N_A_c_266_n N_CIN_c_481_n 0.0408998f $X=3.3 $Y=1.005 $X2=0 $Y2=0
cc_289 N_A_c_271_n N_CIN_c_481_n 0.0123173f $X=1.05 $Y=1.005 $X2=0 $Y2=0
cc_290 N_A_c_261_n N_CIN_c_482_n 0.00128106f $X=4.505 $Y=1.66 $X2=0 $Y2=0
cc_291 N_A_c_269_n N_CIN_c_482_n 0.00210963f $X=5.81 $Y=1.02 $X2=0 $Y2=0
cc_292 N_A_c_260_n N_CIN_c_483_n 0.00383972f $X=3.54 $Y=1.66 $X2=0 $Y2=0
cc_293 N_A_c_261_n N_CIN_c_483_n 0.00695088f $X=4.505 $Y=1.66 $X2=0 $Y2=0
cc_294 N_A_c_267_n N_CIN_c_483_n 0.0124273f $X=3.465 $Y=1.29 $X2=0 $Y2=0
cc_295 N_A_c_268_n N_CIN_c_483_n 0.0261716f $X=4.38 $Y=1.005 $X2=0 $Y2=0
cc_296 A N_CIN_c_483_n 0.0145682f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_297 N_A_c_269_n N_A_465_249#_M1016_d 0.00176461f $X=5.81 $Y=1.02 $X2=-0.19
+ $Y2=-0.245
cc_298 N_A_c_266_n N_A_465_249#_M1004_g 0.0150305f $X=3.3 $Y=1.005 $X2=0 $Y2=0
cc_299 N_A_c_266_n N_A_465_249#_c_642_n 0.00428181f $X=3.3 $Y=1.005 $X2=0 $Y2=0
cc_300 N_A_c_260_n N_A_465_249#_c_653_n 0.00180782f $X=3.54 $Y=1.66 $X2=0 $Y2=0
cc_301 N_A_c_266_n N_A_465_249#_c_653_n 0.00808653f $X=3.3 $Y=1.005 $X2=0 $Y2=0
cc_302 N_A_c_260_n N_A_465_249#_c_668_n 0.00303197f $X=3.54 $Y=1.66 $X2=0 $Y2=0
cc_303 N_A_c_260_n N_A_465_249#_c_654_n 0.0135694f $X=3.54 $Y=1.66 $X2=0 $Y2=0
cc_304 N_A_c_261_n N_A_465_249#_c_654_n 0.0194312f $X=4.505 $Y=1.66 $X2=0 $Y2=0
cc_305 N_A_c_263_n N_A_465_249#_c_654_n 5.65261e-19 $X=6.055 $Y=1.66 $X2=0 $Y2=0
cc_306 N_A_c_267_n N_A_465_249#_c_654_n 0.00415742f $X=3.465 $Y=1.29 $X2=0 $Y2=0
cc_307 A N_A_465_249#_c_654_n 0.00389368f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_308 N_A_c_263_n N_A_465_249#_c_674_n 0.00461809f $X=6.055 $Y=1.66 $X2=0 $Y2=0
cc_309 N_A_c_265_n N_A_465_249#_c_674_n 0.0037443f $X=6.485 $Y=1.11 $X2=0 $Y2=0
cc_310 N_A_c_269_n N_A_465_249#_c_674_n 0.0400333f $X=5.81 $Y=1.02 $X2=0 $Y2=0
cc_311 N_A_c_272_n N_A_465_249#_c_674_n 0.00489085f $X=6.045 $Y=1.41 $X2=0 $Y2=0
cc_312 N_A_c_263_n N_A_465_249#_c_655_n 0.0157391f $X=6.055 $Y=1.66 $X2=0 $Y2=0
cc_313 N_A_c_264_n N_A_465_249#_c_655_n 0.00268633f $X=6.41 $Y=1.185 $X2=0 $Y2=0
cc_314 N_A_c_269_n N_A_465_249#_c_655_n 0.00480772f $X=5.81 $Y=1.02 $X2=0 $Y2=0
cc_315 N_A_c_272_n N_A_465_249#_c_655_n 0.0247281f $X=6.045 $Y=1.41 $X2=0 $Y2=0
cc_316 N_A_c_263_n N_A_465_249#_c_682_n 9.62124e-19 $X=6.055 $Y=1.66 $X2=0 $Y2=0
cc_317 N_A_c_265_n N_A_465_249#_c_682_n 0.00729181f $X=6.485 $Y=1.11 $X2=0 $Y2=0
cc_318 N_A_c_269_n N_A_465_249#_c_682_n 0.00366113f $X=5.81 $Y=1.02 $X2=0 $Y2=0
cc_319 N_A_c_263_n N_A_465_249#_c_645_n 0.00628146f $X=6.055 $Y=1.66 $X2=0 $Y2=0
cc_320 N_A_c_264_n N_A_465_249#_c_645_n 0.0104389f $X=6.41 $Y=1.185 $X2=0 $Y2=0
cc_321 N_A_c_270_n N_A_465_249#_c_645_n 0.00600815f $X=5.895 $Y=1.32 $X2=0 $Y2=0
cc_322 N_A_c_272_n N_A_465_249#_c_645_n 0.019392f $X=6.045 $Y=1.41 $X2=0 $Y2=0
cc_323 N_A_c_264_n N_A_465_249#_c_646_n 0.00113076f $X=6.41 $Y=1.185 $X2=0 $Y2=0
cc_324 N_A_c_265_n N_A_465_249#_c_646_n 0.00265319f $X=6.485 $Y=1.11 $X2=0 $Y2=0
cc_325 N_A_c_263_n N_A_465_249#_c_647_n 0.00258911f $X=6.055 $Y=1.66 $X2=0 $Y2=0
cc_326 N_A_c_264_n N_A_465_249#_c_647_n 0.00821163f $X=6.41 $Y=1.185 $X2=0 $Y2=0
cc_327 N_A_c_265_n N_A_465_249#_c_647_n 0.0070169f $X=6.485 $Y=1.11 $X2=0 $Y2=0
cc_328 N_A_c_269_n N_A_465_249#_c_647_n 0.0114981f $X=5.81 $Y=1.02 $X2=0 $Y2=0
cc_329 N_A_c_270_n N_A_465_249#_c_647_n 0.00335532f $X=5.895 $Y=1.32 $X2=0 $Y2=0
cc_330 N_A_c_272_n N_A_465_249#_c_647_n 0.00419754f $X=6.045 $Y=1.41 $X2=0 $Y2=0
cc_331 N_A_c_266_n N_A_465_249#_c_649_n 0.0313166f $X=3.3 $Y=1.005 $X2=0 $Y2=0
cc_332 N_A_c_267_n N_A_465_249#_c_649_n 0.00649172f $X=3.465 $Y=1.29 $X2=0 $Y2=0
cc_333 N_A_c_262_n N_A_465_249#_c_699_n 0.00105103f $X=4.605 $Y=1.125 $X2=0
+ $Y2=0
cc_334 N_A_c_269_n N_A_465_249#_c_699_n 0.0161182f $X=5.81 $Y=1.02 $X2=0 $Y2=0
cc_335 N_A_c_257_n N_B_M1025_g 0.0278764f $X=1.01 $Y=1.765 $X2=0 $Y2=0
cc_336 N_A_M1008_g N_B_M1025_g 0.0538361f $X=1.11 $Y=0.695 $X2=0 $Y2=0
cc_337 N_A_c_266_n N_B_M1025_g 0.0134851f $X=3.3 $Y=1.005 $X2=0 $Y2=0
cc_338 N_A_c_271_n N_B_M1025_g 0.00373251f $X=1.05 $Y=1.005 $X2=0 $Y2=0
cc_339 N_A_c_257_n N_B_M1005_g 0.0388508f $X=1.01 $Y=1.765 $X2=0 $Y2=0
cc_340 N_A_c_259_n N_B_c_825_n 8.46159e-19 $X=3.53 $Y=1.125 $X2=0 $Y2=0
cc_341 N_A_c_260_n N_B_c_825_n 0.0167155f $X=3.54 $Y=1.66 $X2=0 $Y2=0
cc_342 N_A_c_266_n N_B_c_825_n 0.00109957f $X=3.3 $Y=1.005 $X2=0 $Y2=0
cc_343 N_A_c_267_n N_B_c_825_n 0.00242117f $X=3.465 $Y=1.29 $X2=0 $Y2=0
cc_344 N_A_c_260_n N_B_c_826_n 0.00669739f $X=3.54 $Y=1.66 $X2=0 $Y2=0
cc_345 N_A_c_260_n N_B_c_839_n 0.00105762f $X=3.54 $Y=1.66 $X2=0 $Y2=0
cc_346 N_A_c_260_n N_B_M1019_g 0.0269033f $X=3.54 $Y=1.66 $X2=0 $Y2=0
cc_347 N_A_c_260_n N_B_c_843_n 0.0100467f $X=3.54 $Y=1.66 $X2=0 $Y2=0
cc_348 N_A_c_261_n N_B_c_843_n 0.0104018f $X=4.505 $Y=1.66 $X2=0 $Y2=0
cc_349 N_A_c_261_n N_B_c_827_n 0.0202139f $X=4.505 $Y=1.66 $X2=0 $Y2=0
cc_350 N_A_c_269_n N_B_c_827_n 0.00352699f $X=5.81 $Y=1.02 $X2=0 $Y2=0
cc_351 A N_B_c_827_n 0.00199957f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_352 N_A_c_261_n N_B_c_828_n 0.00818364f $X=4.505 $Y=1.66 $X2=0 $Y2=0
cc_353 N_A_c_261_n N_B_c_845_n 0.00209048f $X=4.505 $Y=1.66 $X2=0 $Y2=0
cc_354 N_A_c_261_n N_B_M1010_g 0.0390434f $X=4.505 $Y=1.66 $X2=0 $Y2=0
cc_355 N_A_c_263_n N_B_c_849_n 0.010379f $X=6.055 $Y=1.66 $X2=0 $Y2=0
cc_356 N_A_c_263_n N_B_M1001_g 0.0116289f $X=6.055 $Y=1.66 $X2=0 $Y2=0
cc_357 N_A_c_265_n N_B_M1013_g 0.0176832f $X=6.485 $Y=1.11 $X2=0 $Y2=0
cc_358 N_A_c_257_n N_B_c_851_n 0.0032909f $X=1.01 $Y=1.765 $X2=0 $Y2=0
cc_359 N_A_c_259_n N_B_c_830_n 0.0208927f $X=3.53 $Y=1.125 $X2=0 $Y2=0
cc_360 N_A_c_266_n N_B_c_830_n 0.0133079f $X=3.3 $Y=1.005 $X2=0 $Y2=0
cc_361 N_A_c_262_n N_B_c_831_n 0.0464607f $X=4.605 $Y=1.125 $X2=0 $Y2=0
cc_362 N_A_c_269_n N_B_c_831_n 0.011404f $X=5.81 $Y=1.02 $X2=0 $Y2=0
cc_363 N_A_c_263_n N_B_c_832_n 0.00542945f $X=6.055 $Y=1.66 $X2=0 $Y2=0
cc_364 N_A_c_257_n N_VPWR_c_1019_n 0.00788947f $X=1.01 $Y=1.765 $X2=0 $Y2=0
cc_365 N_A_c_260_n N_VPWR_c_1020_n 0.00401699f $X=3.54 $Y=1.66 $X2=0 $Y2=0
cc_366 N_A_c_260_n N_VPWR_c_1021_n 6.62299e-19 $X=3.54 $Y=1.66 $X2=0 $Y2=0
cc_367 N_A_c_261_n N_VPWR_c_1021_n 0.0126719f $X=4.505 $Y=1.66 $X2=0 $Y2=0
cc_368 N_A_c_263_n N_VPWR_c_1022_n 0.00760524f $X=6.055 $Y=1.66 $X2=0 $Y2=0
cc_369 N_A_c_257_n N_VPWR_c_1027_n 0.0049405f $X=1.01 $Y=1.765 $X2=0 $Y2=0
cc_370 N_A_c_257_n N_VPWR_c_1018_n 0.00508379f $X=1.01 $Y=1.765 $X2=0 $Y2=0
cc_371 N_A_c_260_n N_VPWR_c_1018_n 9.39239e-19 $X=3.54 $Y=1.66 $X2=0 $Y2=0
cc_372 N_A_c_261_n N_VPWR_c_1018_n 9.14192e-19 $X=4.505 $Y=1.66 $X2=0 $Y2=0
cc_373 N_A_c_263_n N_VPWR_c_1018_n 8.82885e-19 $X=6.055 $Y=1.66 $X2=0 $Y2=0
cc_374 N_A_c_260_n N_A_509_347#_c_1137_n 0.00978463f $X=3.54 $Y=1.66 $X2=0 $Y2=0
cc_375 N_A_c_260_n N_A_509_347#_c_1133_n 0.0070513f $X=3.54 $Y=1.66 $X2=0 $Y2=0
cc_376 N_A_c_263_n N_A_1107_347#_c_1174_n 3.90888e-19 $X=6.055 $Y=1.66 $X2=0
+ $Y2=0
cc_377 N_A_c_263_n N_A_1107_347#_c_1178_n 0.0139404f $X=6.055 $Y=1.66 $X2=0
+ $Y2=0
cc_378 N_A_c_266_n N_VGND_M1012_d 0.00252521f $X=3.3 $Y=1.005 $X2=0 $Y2=0
cc_379 N_A_c_435_p N_VGND_M1012_d 0.00106822f $X=3.465 $Y=1.005 $X2=0 $Y2=0
cc_380 N_A_c_268_n N_VGND_M1002_d 0.0035226f $X=4.38 $Y=1.005 $X2=0 $Y2=0
cc_381 N_A_c_310_p N_VGND_M1002_d 0.0011084f $X=4.545 $Y=1.012 $X2=0 $Y2=0
cc_382 N_A_c_259_n N_VGND_c_1220_n 0.00314919f $X=3.53 $Y=1.125 $X2=0 $Y2=0
cc_383 N_A_c_261_n N_VGND_c_1221_n 6.06391e-19 $X=4.505 $Y=1.66 $X2=0 $Y2=0
cc_384 N_A_c_262_n N_VGND_c_1221_n 0.016605f $X=4.605 $Y=1.125 $X2=0 $Y2=0
cc_385 N_A_c_268_n N_VGND_c_1221_n 0.0199906f $X=4.38 $Y=1.005 $X2=0 $Y2=0
cc_386 N_A_c_310_p N_VGND_c_1221_n 0.00871655f $X=4.545 $Y=1.012 $X2=0 $Y2=0
cc_387 N_A_c_265_n N_VGND_c_1222_n 9.17969e-19 $X=6.485 $Y=1.11 $X2=0 $Y2=0
cc_388 N_A_M1008_g N_VGND_c_1224_n 0.00407101f $X=1.11 $Y=0.695 $X2=0 $Y2=0
cc_389 N_A_M1008_g N_VGND_c_1225_n 0.00317047f $X=1.11 $Y=0.695 $X2=0 $Y2=0
cc_390 N_A_c_262_n N_VGND_c_1226_n 0.00379792f $X=4.605 $Y=1.125 $X2=0 $Y2=0
cc_391 N_A_c_265_n N_VGND_c_1226_n 0.0027564f $X=6.485 $Y=1.11 $X2=0 $Y2=0
cc_392 N_A_M1008_g N_VGND_c_1229_n 0.00544287f $X=1.11 $Y=0.695 $X2=0 $Y2=0
cc_393 N_A_c_259_n N_VGND_c_1229_n 0.00544287f $X=3.53 $Y=1.125 $X2=0 $Y2=0
cc_394 N_A_c_262_n N_VGND_c_1229_n 0.00457201f $X=4.605 $Y=1.125 $X2=0 $Y2=0
cc_395 N_A_c_265_n N_VGND_c_1229_n 0.00544287f $X=6.485 $Y=1.11 $X2=0 $Y2=0
cc_396 N_A_c_259_n N_VGND_c_1230_n 0.00397421f $X=3.53 $Y=1.125 $X2=0 $Y2=0
cc_397 N_A_c_266_n A_237_75# 0.00134267f $X=3.3 $Y=1.005 $X2=-0.19 $Y2=-0.245
cc_398 N_A_c_266_n A_315_75# 0.00134267f $X=3.3 $Y=1.005 $X2=-0.19 $Y2=-0.245
cc_399 N_A_c_266_n N_A_501_75#_M1004_d 0.0026214f $X=3.3 $Y=1.005 $X2=-0.19
+ $Y2=-0.245
cc_400 N_A_c_268_n N_A_501_75#_M1015_d 0.00176461f $X=4.38 $Y=1.005 $X2=0 $Y2=0
cc_401 N_A_c_259_n N_A_501_75#_c_1335_n 0.00936066f $X=3.53 $Y=1.125 $X2=0 $Y2=0
cc_402 N_A_c_260_n N_A_501_75#_c_1335_n 5.87191e-19 $X=3.54 $Y=1.66 $X2=0 $Y2=0
cc_403 N_A_c_435_p N_A_501_75#_c_1335_n 0.0171542f $X=3.465 $Y=1.005 $X2=0 $Y2=0
cc_404 N_A_c_259_n N_A_501_75#_c_1332_n 7.1726e-19 $X=3.53 $Y=1.125 $X2=0 $Y2=0
cc_405 N_A_c_266_n N_A_501_75#_c_1332_n 0.0472581f $X=3.3 $Y=1.005 $X2=0 $Y2=0
cc_406 N_A_c_259_n N_A_501_75#_c_1340_n 0.00483163f $X=3.53 $Y=1.125 $X2=0 $Y2=0
cc_407 N_A_c_262_n N_A_501_75#_c_1340_n 3.54619e-19 $X=4.605 $Y=1.125 $X2=0
+ $Y2=0
cc_408 N_A_c_268_n N_A_501_75#_c_1340_n 0.0144331f $X=4.38 $Y=1.005 $X2=0 $Y2=0
cc_409 N_A_c_435_p N_A_501_75#_c_1340_n 0.00185147f $X=3.465 $Y=1.005 $X2=0
+ $Y2=0
cc_410 N_A_c_269_n A_936_75# 0.0048076f $X=5.81 $Y=1.02 $X2=-0.19 $Y2=-0.245
cc_411 N_A_c_269_n N_A_1100_75#_M1020_d 0.00536422f $X=5.81 $Y=1.02 $X2=-0.19
+ $Y2=-0.245
cc_412 N_A_c_263_n N_A_1100_75#_c_1359_n 3.90359e-19 $X=6.055 $Y=1.66 $X2=0
+ $Y2=0
cc_413 N_A_c_265_n N_A_1100_75#_c_1359_n 0.0111244f $X=6.485 $Y=1.11 $X2=0 $Y2=0
cc_414 N_A_c_265_n N_A_1100_75#_c_1364_n 0.0104474f $X=6.485 $Y=1.11 $X2=0 $Y2=0
cc_415 N_A_c_265_n N_A_1100_75#_c_1365_n 0.00656693f $X=6.485 $Y=1.11 $X2=0
+ $Y2=0
cc_416 N_CIN_c_478_n N_A_465_249#_M1010_d 3.91994e-19 $X=5.155 $Y=1.425 $X2=0
+ $Y2=0
cc_417 N_CIN_c_482_n N_A_465_249#_M1010_d 8.14058e-19 $X=5.04 $Y=1.665 $X2=0
+ $Y2=0
cc_418 N_CIN_M1026_g N_A_465_249#_M1004_g 0.0258374f $X=1.89 $Y=0.695 $X2=0
+ $Y2=0
cc_419 N_CIN_c_473_n N_A_465_249#_c_642_n 0.0354191f $X=2.02 $Y=1.66 $X2=0 $Y2=0
cc_420 N_CIN_c_489_n N_A_465_249#_c_642_n 0.00982988f $X=3.935 $Y=1.665 $X2=0
+ $Y2=0
cc_421 N_CIN_c_481_n N_A_465_249#_c_642_n 3.95958e-19 $X=1.68 $Y=1.665 $X2=0
+ $Y2=0
cc_422 N_CIN_c_489_n N_A_465_249#_c_653_n 0.0201297f $X=3.935 $Y=1.665 $X2=0
+ $Y2=0
cc_423 N_CIN_c_483_n N_A_465_249#_c_653_n 0.00316748f $X=4.005 $Y=1.41 $X2=0
+ $Y2=0
cc_424 N_CIN_c_475_n N_A_465_249#_c_654_n 0.0154823f $X=4.045 $Y=1.66 $X2=0
+ $Y2=0
cc_425 N_CIN_c_477_n N_A_465_249#_c_654_n 0.0242973f $X=5.46 $Y=1.66 $X2=0 $Y2=0
cc_426 N_CIN_c_478_n N_A_465_249#_c_654_n 0.0137014f $X=5.155 $Y=1.425 $X2=0
+ $Y2=0
cc_427 N_CIN_c_479_n N_A_465_249#_c_654_n 0.0187439f $X=5.475 $Y=1.41 $X2=0
+ $Y2=0
cc_428 N_CIN_c_489_n N_A_465_249#_c_654_n 0.0227402f $X=3.935 $Y=1.665 $X2=0
+ $Y2=0
cc_429 N_CIN_c_491_n N_A_465_249#_c_654_n 0.0233361f $X=4.895 $Y=1.665 $X2=0
+ $Y2=0
cc_430 N_CIN_c_480_n N_A_465_249#_c_654_n 0.00339089f $X=4.225 $Y=1.665 $X2=0
+ $Y2=0
cc_431 N_CIN_c_482_n N_A_465_249#_c_654_n 0.00526688f $X=5.04 $Y=1.665 $X2=0
+ $Y2=0
cc_432 N_CIN_c_483_n N_A_465_249#_c_654_n 0.0171765f $X=4.005 $Y=1.41 $X2=0
+ $Y2=0
cc_433 N_CIN_M1020_g N_A_465_249#_c_674_n 0.0107451f $X=5.425 $Y=0.695 $X2=0
+ $Y2=0
cc_434 N_CIN_c_477_n N_A_465_249#_c_655_n 0.00750113f $X=5.46 $Y=1.66 $X2=0
+ $Y2=0
cc_435 N_CIN_c_479_n N_A_465_249#_c_655_n 0.00842675f $X=5.475 $Y=1.41 $X2=0
+ $Y2=0
cc_436 N_CIN_M1020_g N_A_465_249#_c_682_n 0.00366676f $X=5.425 $Y=0.695 $X2=0
+ $Y2=0
cc_437 N_CIN_M1020_g N_A_465_249#_c_647_n 3.99689e-19 $X=5.425 $Y=0.695 $X2=0
+ $Y2=0
cc_438 N_CIN_c_473_n N_A_465_249#_c_649_n 3.97232e-19 $X=2.02 $Y=1.66 $X2=0
+ $Y2=0
cc_439 N_CIN_c_489_n N_A_465_249#_c_649_n 0.0252619f $X=3.935 $Y=1.665 $X2=0
+ $Y2=0
cc_440 N_CIN_c_481_n N_A_465_249#_c_649_n 0.021248f $X=1.68 $Y=1.665 $X2=0 $Y2=0
cc_441 N_CIN_M1020_g N_A_465_249#_c_699_n 0.00851142f $X=5.425 $Y=0.695 $X2=0
+ $Y2=0
cc_442 N_CIN_M1026_g N_B_M1025_g 0.0555179f $X=1.89 $Y=0.695 $X2=0 $Y2=0
cc_443 N_CIN_c_473_n N_B_M1025_g 0.0261117f $X=2.02 $Y=1.66 $X2=0 $Y2=0
cc_444 N_CIN_c_490_n N_B_M1025_g 0.00332777f $X=1.825 $Y=1.665 $X2=0 $Y2=0
cc_445 N_CIN_c_481_n N_B_M1025_g 0.0115329f $X=1.68 $Y=1.665 $X2=0 $Y2=0
cc_446 N_CIN_c_473_n N_B_c_836_n 0.0103487f $X=2.02 $Y=1.66 $X2=0 $Y2=0
cc_447 N_CIN_c_489_n N_B_c_841_n 0.00282348f $X=3.935 $Y=1.665 $X2=0 $Y2=0
cc_448 N_CIN_c_475_n N_B_c_843_n 0.0103562f $X=4.045 $Y=1.66 $X2=0 $Y2=0
cc_449 N_CIN_M1020_g N_B_c_827_n 0.00833387f $X=5.425 $Y=0.695 $X2=0 $Y2=0
cc_450 N_CIN_c_477_n N_B_c_828_n 0.021431f $X=5.46 $Y=1.66 $X2=0 $Y2=0
cc_451 N_CIN_c_478_n N_B_c_828_n 0.0107765f $X=5.155 $Y=1.425 $X2=0 $Y2=0
cc_452 N_CIN_c_479_n N_B_c_828_n 4.59542e-19 $X=5.475 $Y=1.41 $X2=0 $Y2=0
cc_453 N_CIN_c_477_n N_B_c_845_n 0.00278823f $X=5.46 $Y=1.66 $X2=0 $Y2=0
cc_454 N_CIN_c_477_n N_B_c_847_n 0.00370009f $X=5.46 $Y=1.66 $X2=0 $Y2=0
cc_455 N_CIN_c_478_n N_B_c_847_n 0.00375646f $X=5.155 $Y=1.425 $X2=0 $Y2=0
cc_456 N_CIN_c_482_n N_B_c_847_n 5.45625e-19 $X=5.04 $Y=1.665 $X2=0 $Y2=0
cc_457 N_CIN_c_477_n N_B_M1010_g 0.0170667f $X=5.46 $Y=1.66 $X2=0 $Y2=0
cc_458 N_CIN_c_478_n N_B_M1010_g 0.00403934f $X=5.155 $Y=1.425 $X2=0 $Y2=0
cc_459 N_CIN_c_482_n N_B_M1010_g 0.00140427f $X=5.04 $Y=1.665 $X2=0 $Y2=0
cc_460 N_CIN_c_477_n N_B_c_849_n 0.00988928f $X=5.46 $Y=1.66 $X2=0 $Y2=0
cc_461 N_CIN_c_473_n N_B_c_851_n 0.040996f $X=2.02 $Y=1.66 $X2=0 $Y2=0
cc_462 N_CIN_c_490_n N_B_c_851_n 0.00115766f $X=1.825 $Y=1.665 $X2=0 $Y2=0
cc_463 N_CIN_c_481_n N_B_c_851_n 0.00186213f $X=1.68 $Y=1.665 $X2=0 $Y2=0
cc_464 N_CIN_M1020_g N_B_c_831_n 0.0214903f $X=5.425 $Y=0.695 $X2=0 $Y2=0
cc_465 N_CIN_c_489_n N_VPWR_M1019_d 0.00220021f $X=3.935 $Y=1.665 $X2=0 $Y2=0
cc_466 N_CIN_c_491_n N_VPWR_M1007_d 0.00169375f $X=4.895 $Y=1.665 $X2=0 $Y2=0
cc_467 N_CIN_c_480_n N_VPWR_M1007_d 0.00116927f $X=4.225 $Y=1.665 $X2=0 $Y2=0
cc_468 N_CIN_c_483_n N_VPWR_M1007_d 8.48983e-19 $X=4.005 $Y=1.41 $X2=0 $Y2=0
cc_469 N_CIN_c_475_n N_VPWR_c_1021_n 0.00927589f $X=4.045 $Y=1.66 $X2=0 $Y2=0
cc_470 N_CIN_c_477_n N_VPWR_c_1022_n 5.24658e-19 $X=5.46 $Y=1.66 $X2=0 $Y2=0
cc_471 N_CIN_c_473_n N_VPWR_c_1018_n 9.39239e-19 $X=2.02 $Y=1.66 $X2=0 $Y2=0
cc_472 N_CIN_c_475_n N_VPWR_c_1018_n 8.51577e-19 $X=4.045 $Y=1.66 $X2=0 $Y2=0
cc_473 N_CIN_c_477_n N_VPWR_c_1018_n 9.39239e-19 $X=5.46 $Y=1.66 $X2=0 $Y2=0
cc_474 N_CIN_c_489_n A_318_389# 9.88021e-19 $X=3.935 $Y=1.665 $X2=-0.19
+ $Y2=-0.245
cc_475 N_CIN_c_490_n A_318_389# 0.00169613f $X=1.825 $Y=1.665 $X2=-0.19
+ $Y2=-0.245
cc_476 N_CIN_c_481_n A_318_389# 0.00100152f $X=1.68 $Y=1.665 $X2=-0.19
+ $Y2=-0.245
cc_477 N_CIN_c_489_n N_A_509_347#_M1006_d 0.00129319f $X=3.935 $Y=1.665
+ $X2=-0.19 $Y2=-0.245
cc_478 N_CIN_c_489_n N_A_509_347#_M1003_d 0.00187641f $X=3.935 $Y=1.665 $X2=0
+ $Y2=0
cc_479 N_CIN_c_483_n N_A_509_347#_M1003_d 0.00147899f $X=4.005 $Y=1.41 $X2=0
+ $Y2=0
cc_480 N_CIN_c_489_n N_A_509_347#_c_1134_n 0.00184039f $X=3.935 $Y=1.665 $X2=0
+ $Y2=0
cc_481 N_CIN_c_489_n N_A_509_347#_c_1137_n 0.00149783f $X=3.935 $Y=1.665 $X2=0
+ $Y2=0
cc_482 N_CIN_c_475_n N_A_509_347#_c_1133_n 0.00254395f $X=4.045 $Y=1.66 $X2=0
+ $Y2=0
cc_483 N_CIN_c_491_n A_916_347# 0.00260705f $X=4.895 $Y=1.665 $X2=-0.19
+ $Y2=-0.245
cc_484 N_CIN_c_482_n A_916_347# 0.00103224f $X=5.04 $Y=1.665 $X2=-0.19
+ $Y2=-0.245
cc_485 N_CIN_c_477_n N_A_1107_347#_c_1179_n 0.00147836f $X=5.46 $Y=1.66 $X2=0
+ $Y2=0
cc_486 N_CIN_c_477_n N_A_1107_347#_c_1174_n 0.00402977f $X=5.46 $Y=1.66 $X2=0
+ $Y2=0
cc_487 N_CIN_M1002_g N_VGND_c_1220_n 0.00431894f $X=3.96 $Y=0.695 $X2=0 $Y2=0
cc_488 N_CIN_M1002_g N_VGND_c_1221_n 0.0064725f $X=3.96 $Y=0.695 $X2=0 $Y2=0
cc_489 N_CIN_M1026_g N_VGND_c_1225_n 0.00313567f $X=1.89 $Y=0.695 $X2=0 $Y2=0
cc_490 N_CIN_M1020_g N_VGND_c_1226_n 0.00316607f $X=5.425 $Y=0.695 $X2=0 $Y2=0
cc_491 N_CIN_M1026_g N_VGND_c_1229_n 0.00544287f $X=1.89 $Y=0.695 $X2=0 $Y2=0
cc_492 N_CIN_M1002_g N_VGND_c_1229_n 0.00544287f $X=3.96 $Y=0.695 $X2=0 $Y2=0
cc_493 N_CIN_M1020_g N_VGND_c_1229_n 0.00544287f $X=5.425 $Y=0.695 $X2=0 $Y2=0
cc_494 N_CIN_M1002_g N_A_501_75#_c_1340_n 0.00449722f $X=3.96 $Y=0.695 $X2=0
+ $Y2=0
cc_495 N_CIN_M1020_g N_A_1100_75#_c_1359_n 0.00645788f $X=5.425 $Y=0.695 $X2=0
+ $Y2=0
cc_496 N_A_465_249#_c_642_n N_B_c_836_n 0.0103487f $X=2.47 $Y=1.66 $X2=0 $Y2=0
cc_497 N_A_465_249#_c_642_n N_B_c_826_n 0.0197335f $X=2.47 $Y=1.66 $X2=0 $Y2=0
cc_498 N_A_465_249#_c_649_n N_B_c_826_n 0.00631568f $X=2.49 $Y=1.41 $X2=0 $Y2=0
cc_499 N_A_465_249#_c_642_n N_B_c_839_n 0.00226496f $X=2.47 $Y=1.66 $X2=0 $Y2=0
cc_500 N_A_465_249#_c_642_n N_B_c_841_n 0.00353516f $X=2.47 $Y=1.66 $X2=0 $Y2=0
cc_501 N_A_465_249#_c_653_n N_B_c_841_n 0.00516123f $X=3.03 $Y=1.71 $X2=0 $Y2=0
cc_502 N_A_465_249#_c_642_n N_B_M1019_g 0.0141617f $X=2.47 $Y=1.66 $X2=0 $Y2=0
cc_503 N_A_465_249#_c_653_n N_B_M1019_g 0.00854511f $X=3.03 $Y=1.71 $X2=0 $Y2=0
cc_504 N_A_465_249#_c_661_n N_B_M1019_g 0.0020345f $X=3.2 $Y=2.035 $X2=0 $Y2=0
cc_505 N_A_465_249#_c_654_n N_B_c_845_n 5.08057e-19 $X=5.07 $Y=2.035 $X2=0 $Y2=0
cc_506 N_A_465_249#_c_654_n N_B_M1010_g 0.0310668f $X=5.07 $Y=2.035 $X2=0 $Y2=0
cc_507 N_A_465_249#_c_654_n N_B_c_849_n 0.00427141f $X=5.07 $Y=2.035 $X2=0 $Y2=0
cc_508 N_A_465_249#_c_655_n N_B_M1001_g 0.00393101f $X=6.38 $Y=1.83 $X2=0 $Y2=0
cc_509 N_A_465_249#_c_643_n N_B_M1013_g 0.00323528f $X=8.055 $Y=1.385 $X2=0
+ $Y2=0
cc_510 N_A_465_249#_c_645_n N_B_M1013_g 0.00187649f $X=6.465 $Y=1.745 $X2=0
+ $Y2=0
cc_511 N_A_465_249#_c_646_n N_B_M1013_g 0.0136844f $X=7.71 $Y=1.065 $X2=0 $Y2=0
cc_512 N_A_465_249#_c_648_n N_B_M1013_g 0.00252947f $X=7.875 $Y=1.385 $X2=0
+ $Y2=0
cc_513 N_A_465_249#_M1004_g N_B_c_830_n 0.0225165f $X=2.43 $Y=0.695 $X2=0 $Y2=0
cc_514 N_A_465_249#_c_699_n N_B_c_831_n 0.00617071f $X=5.21 $Y=0.6 $X2=0 $Y2=0
cc_515 N_A_465_249#_c_643_n N_B_c_832_n 0.0154379f $X=8.055 $Y=1.385 $X2=0 $Y2=0
cc_516 N_A_465_249#_c_645_n N_B_c_832_n 0.00420628f $X=6.465 $Y=1.745 $X2=0
+ $Y2=0
cc_517 N_A_465_249#_c_646_n N_B_c_832_n 0.0036367f $X=7.71 $Y=1.065 $X2=0 $Y2=0
cc_518 N_A_465_249#_c_648_n N_B_c_832_n 9.69264e-19 $X=7.875 $Y=1.385 $X2=0
+ $Y2=0
cc_519 N_A_465_249#_c_651_n N_B_c_833_n 3.79438e-19 $X=8.145 $Y=1.765 $X2=0
+ $Y2=0
cc_520 N_A_465_249#_c_643_n N_B_c_833_n 0.00452614f $X=8.055 $Y=1.385 $X2=0
+ $Y2=0
cc_521 N_A_465_249#_c_655_n N_B_c_833_n 0.00248868f $X=6.38 $Y=1.83 $X2=0 $Y2=0
cc_522 N_A_465_249#_c_645_n N_B_c_833_n 0.0252993f $X=6.465 $Y=1.745 $X2=0 $Y2=0
cc_523 N_A_465_249#_c_646_n N_B_c_833_n 0.0511978f $X=7.71 $Y=1.065 $X2=0 $Y2=0
cc_524 N_A_465_249#_c_648_n N_B_c_833_n 0.0138522f $X=7.875 $Y=1.385 $X2=0 $Y2=0
cc_525 N_A_465_249#_c_653_n N_VPWR_M1019_d 9.32624e-19 $X=3.03 $Y=1.71 $X2=0
+ $Y2=0
cc_526 N_A_465_249#_c_668_n N_VPWR_M1019_d 0.00190874f $X=3.115 $Y=1.95 $X2=0
+ $Y2=0
cc_527 N_A_465_249#_c_654_n N_VPWR_M1019_d 0.00572787f $X=5.07 $Y=2.035 $X2=0
+ $Y2=0
cc_528 N_A_465_249#_c_661_n N_VPWR_M1019_d 0.00209835f $X=3.2 $Y=2.035 $X2=0
+ $Y2=0
cc_529 N_A_465_249#_c_654_n N_VPWR_M1007_d 0.00473314f $X=5.07 $Y=2.035 $X2=0
+ $Y2=0
cc_530 N_A_465_249#_c_655_n N_VPWR_M1022_d 0.00990454f $X=6.38 $Y=1.83 $X2=0
+ $Y2=0
cc_531 N_A_465_249#_c_654_n N_VPWR_c_1021_n 0.0270428f $X=5.07 $Y=2.035 $X2=0
+ $Y2=0
cc_532 N_A_465_249#_c_651_n N_VPWR_c_1023_n 0.0220569f $X=8.145 $Y=1.765 $X2=0
+ $Y2=0
cc_533 N_A_465_249#_c_643_n N_VPWR_c_1023_n 0.00353544f $X=8.055 $Y=1.385 $X2=0
+ $Y2=0
cc_534 N_A_465_249#_c_648_n N_VPWR_c_1023_n 0.017603f $X=7.875 $Y=1.385 $X2=0
+ $Y2=0
cc_535 N_A_465_249#_c_654_n N_VPWR_c_1028_n 0.00943889f $X=5.07 $Y=2.035 $X2=0
+ $Y2=0
cc_536 N_A_465_249#_c_651_n N_VPWR_c_1030_n 0.00413917f $X=8.145 $Y=1.765 $X2=0
+ $Y2=0
cc_537 N_A_465_249#_c_642_n N_VPWR_c_1018_n 9.39239e-19 $X=2.47 $Y=1.66 $X2=0
+ $Y2=0
cc_538 N_A_465_249#_c_651_n N_VPWR_c_1018_n 0.00821187f $X=8.145 $Y=1.765 $X2=0
+ $Y2=0
cc_539 N_A_465_249#_c_654_n N_VPWR_c_1018_n 0.0115663f $X=5.07 $Y=2.035 $X2=0
+ $Y2=0
cc_540 N_A_465_249#_c_653_n N_A_509_347#_M1006_d 7.65374e-19 $X=3.03 $Y=1.71
+ $X2=-0.19 $Y2=-0.245
cc_541 N_A_465_249#_c_649_n N_A_509_347#_M1006_d 0.00210526f $X=2.49 $Y=1.41
+ $X2=-0.19 $Y2=-0.245
cc_542 N_A_465_249#_c_654_n N_A_509_347#_M1003_d 0.0054536f $X=5.07 $Y=2.035
+ $X2=0 $Y2=0
cc_543 N_A_465_249#_c_642_n N_A_509_347#_c_1134_n 2.11228e-19 $X=2.47 $Y=1.66
+ $X2=0 $Y2=0
cc_544 N_A_465_249#_c_653_n N_A_509_347#_c_1134_n 0.00536428f $X=3.03 $Y=1.71
+ $X2=0 $Y2=0
cc_545 N_A_465_249#_c_649_n N_A_509_347#_c_1134_n 0.0112946f $X=2.49 $Y=1.41
+ $X2=0 $Y2=0
cc_546 N_A_465_249#_c_642_n N_A_509_347#_c_1132_n 0.00110996f $X=2.47 $Y=1.66
+ $X2=0 $Y2=0
cc_547 N_A_465_249#_c_653_n N_A_509_347#_c_1137_n 0.00343931f $X=3.03 $Y=1.71
+ $X2=0 $Y2=0
cc_548 N_A_465_249#_c_654_n N_A_509_347#_c_1137_n 0.0235205f $X=5.07 $Y=2.035
+ $X2=0 $Y2=0
cc_549 N_A_465_249#_c_661_n N_A_509_347#_c_1137_n 0.00872582f $X=3.2 $Y=2.035
+ $X2=0 $Y2=0
cc_550 N_A_465_249#_c_642_n N_A_509_347#_c_1136_n 0.00108366f $X=2.47 $Y=1.66
+ $X2=0 $Y2=0
cc_551 N_A_465_249#_c_654_n N_A_509_347#_c_1133_n 0.0193951f $X=5.07 $Y=2.035
+ $X2=0 $Y2=0
cc_552 N_A_465_249#_c_654_n A_916_347# 0.0124293f $X=5.07 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_553 N_A_465_249#_c_655_n N_A_1107_347#_M1014_d 0.0112797f $X=6.38 $Y=1.83
+ $X2=-0.19 $Y2=-0.245
cc_554 N_A_465_249#_c_654_n N_A_1107_347#_c_1179_n 0.0143691f $X=5.07 $Y=2.035
+ $X2=0 $Y2=0
cc_555 N_A_465_249#_c_655_n N_A_1107_347#_c_1179_n 0.0209652f $X=6.38 $Y=1.83
+ $X2=0 $Y2=0
cc_556 N_A_465_249#_c_654_n N_A_1107_347#_c_1174_n 0.0391091f $X=5.07 $Y=2.035
+ $X2=0 $Y2=0
cc_557 N_A_465_249#_c_655_n N_A_1107_347#_c_1178_n 0.0379011f $X=6.38 $Y=1.83
+ $X2=0 $Y2=0
cc_558 N_A_465_249#_c_644_n COUT 0.0139505f $X=8.145 $Y=1.22 $X2=0 $Y2=0
cc_559 N_A_465_249#_c_644_n COUT 0.00384336f $X=8.145 $Y=1.22 $X2=0 $Y2=0
cc_560 N_A_465_249#_c_646_n COUT 0.00654086f $X=7.71 $Y=1.065 $X2=0 $Y2=0
cc_561 N_A_465_249#_c_651_n COUT 0.00791945f $X=8.145 $Y=1.765 $X2=0 $Y2=0
cc_562 N_A_465_249#_c_644_n COUT 0.0209511f $X=8.145 $Y=1.22 $X2=0 $Y2=0
cc_563 N_A_465_249#_c_646_n COUT 0.00131142f $X=7.71 $Y=1.065 $X2=0 $Y2=0
cc_564 N_A_465_249#_c_648_n COUT 0.0238637f $X=7.875 $Y=1.385 $X2=0 $Y2=0
cc_565 N_A_465_249#_c_646_n N_VGND_M1018_d 0.00531596f $X=7.71 $Y=1.065 $X2=0
+ $Y2=0
cc_566 N_A_465_249#_c_646_n N_VGND_M1017_s 0.00320163f $X=7.71 $Y=1.065 $X2=0
+ $Y2=0
cc_567 N_A_465_249#_c_699_n N_VGND_c_1221_n 0.00896174f $X=5.21 $Y=0.6 $X2=0
+ $Y2=0
cc_568 N_A_465_249#_c_643_n N_VGND_c_1223_n 0.00116085f $X=8.055 $Y=1.385 $X2=0
+ $Y2=0
cc_569 N_A_465_249#_c_644_n N_VGND_c_1223_n 0.00564712f $X=8.145 $Y=1.22 $X2=0
+ $Y2=0
cc_570 N_A_465_249#_c_646_n N_VGND_c_1223_n 0.0189083f $X=7.71 $Y=1.065 $X2=0
+ $Y2=0
cc_571 N_A_465_249#_M1004_g N_VGND_c_1225_n 0.00430851f $X=2.43 $Y=0.695 $X2=0
+ $Y2=0
cc_572 N_A_465_249#_c_674_n N_VGND_c_1226_n 0.00284331f $X=6.15 $Y=0.68 $X2=0
+ $Y2=0
cc_573 N_A_465_249#_c_699_n N_VGND_c_1226_n 0.00841586f $X=5.21 $Y=0.6 $X2=0
+ $Y2=0
cc_574 N_A_465_249#_c_644_n N_VGND_c_1228_n 0.00434272f $X=8.145 $Y=1.22 $X2=0
+ $Y2=0
cc_575 N_A_465_249#_M1004_g N_VGND_c_1229_n 0.00544287f $X=2.43 $Y=0.695 $X2=0
+ $Y2=0
cc_576 N_A_465_249#_c_644_n N_VGND_c_1229_n 0.00828888f $X=8.145 $Y=1.22 $X2=0
+ $Y2=0
cc_577 N_A_465_249#_c_674_n N_VGND_c_1229_n 0.00593054f $X=6.15 $Y=0.68 $X2=0
+ $Y2=0
cc_578 N_A_465_249#_c_699_n N_VGND_c_1229_n 0.0109111f $X=5.21 $Y=0.6 $X2=0
+ $Y2=0
cc_579 N_A_465_249#_M1004_g N_A_501_75#_c_1332_n 0.00433986f $X=2.43 $Y=0.695
+ $X2=0 $Y2=0
cc_580 N_A_465_249#_c_674_n N_A_1100_75#_M1020_d 0.0217685f $X=6.15 $Y=0.68
+ $X2=-0.19 $Y2=-0.245
cc_581 N_A_465_249#_c_682_n N_A_1100_75#_M1020_d 0.00690281f $X=6.235 $Y=0.98
+ $X2=-0.19 $Y2=-0.245
cc_582 N_A_465_249#_c_647_n N_A_1100_75#_M1020_d 0.00149425f $X=6.55 $Y=1.065
+ $X2=-0.19 $Y2=-0.245
cc_583 N_A_465_249#_c_646_n N_A_1100_75#_M1013_d 0.00237104f $X=7.71 $Y=1.065
+ $X2=0 $Y2=0
cc_584 N_A_465_249#_c_674_n N_A_1100_75#_c_1359_n 0.0528994f $X=6.15 $Y=0.68
+ $X2=0 $Y2=0
cc_585 N_A_465_249#_c_647_n N_A_1100_75#_c_1359_n 0.00306218f $X=6.55 $Y=1.065
+ $X2=0 $Y2=0
cc_586 N_A_465_249#_c_674_n N_A_1100_75#_c_1364_n 0.0035178f $X=6.15 $Y=0.68
+ $X2=0 $Y2=0
cc_587 N_A_465_249#_c_646_n N_A_1100_75#_c_1374_n 0.0387969f $X=7.71 $Y=1.065
+ $X2=0 $Y2=0
cc_588 N_A_465_249#_c_674_n N_A_1100_75#_c_1365_n 0.0109254f $X=6.15 $Y=0.68
+ $X2=0 $Y2=0
cc_589 N_A_465_249#_c_682_n N_A_1100_75#_c_1365_n 0.00350045f $X=6.235 $Y=0.98
+ $X2=0 $Y2=0
cc_590 N_A_465_249#_c_647_n N_A_1100_75#_c_1365_n 0.00864961f $X=6.55 $Y=1.065
+ $X2=0 $Y2=0
cc_591 N_A_465_249#_c_644_n N_A_1100_75#_c_1360_n 7.49371e-19 $X=8.145 $Y=1.22
+ $X2=0 $Y2=0
cc_592 N_A_465_249#_c_646_n N_A_1100_75#_c_1360_n 0.020765f $X=7.71 $Y=1.065
+ $X2=0 $Y2=0
cc_593 N_B_M1005_g N_VPWR_c_1019_n 0.00299738f $X=1.515 $Y=2.445 $X2=0 $Y2=0
cc_594 N_B_c_837_n N_VPWR_c_1019_n 0.0039855f $X=1.605 $Y=3.15 $X2=0 $Y2=0
cc_595 N_B_c_839_n N_VPWR_c_1020_n 0.0108045f $X=2.955 $Y=2.9 $X2=0 $Y2=0
cc_596 N_B_M1019_g N_VPWR_c_1020_n 0.00245256f $X=2.955 $Y=2.235 $X2=0 $Y2=0
cc_597 N_B_c_843_n N_VPWR_c_1020_n 0.0242838f $X=4.92 $Y=3.15 $X2=0 $Y2=0
cc_598 N_B_c_843_n N_VPWR_c_1021_n 0.0257782f $X=4.92 $Y=3.15 $X2=0 $Y2=0
cc_599 N_B_c_845_n N_VPWR_c_1021_n 0.00593649f $X=5.01 $Y=2.9 $X2=0 $Y2=0
cc_600 N_B_M1010_g N_VPWR_c_1021_n 0.00159549f $X=5.01 $Y=2.235 $X2=0 $Y2=0
cc_601 N_B_c_849_n N_VPWR_c_1022_n 0.039246f $X=6.8 $Y=3.15 $X2=0 $Y2=0
cc_602 N_B_M1001_g N_VPWR_c_1022_n 0.00773265f $X=6.89 $Y=2.31 $X2=0 $Y2=0
cc_603 N_B_c_854_n N_VPWR_c_1022_n 0.0178816f $X=6.89 $Y=3.15 $X2=0 $Y2=0
cc_604 N_B_c_843_n N_VPWR_c_1024_n 0.0207894f $X=4.92 $Y=3.15 $X2=0 $Y2=0
cc_605 N_B_c_837_n N_VPWR_c_1027_n 0.0531734f $X=1.605 $Y=3.15 $X2=0 $Y2=0
cc_606 N_B_c_843_n N_VPWR_c_1028_n 0.0527197f $X=4.92 $Y=3.15 $X2=0 $Y2=0
cc_607 N_B_c_854_n N_VPWR_c_1029_n 0.00600312f $X=6.89 $Y=3.15 $X2=0 $Y2=0
cc_608 N_B_c_836_n N_VPWR_c_1018_n 0.0461871f $X=2.865 $Y=3.15 $X2=0 $Y2=0
cc_609 N_B_c_837_n N_VPWR_c_1018_n 0.0132496f $X=1.605 $Y=3.15 $X2=0 $Y2=0
cc_610 N_B_c_843_n N_VPWR_c_1018_n 0.0478036f $X=4.92 $Y=3.15 $X2=0 $Y2=0
cc_611 N_B_c_849_n N_VPWR_c_1018_n 0.0321787f $X=6.8 $Y=3.15 $X2=0 $Y2=0
cc_612 N_B_c_852_n N_VPWR_c_1018_n 0.0107686f $X=2.955 $Y=3.15 $X2=0 $Y2=0
cc_613 N_B_c_853_n N_VPWR_c_1018_n 0.0100229f $X=5.01 $Y=3.15 $X2=0 $Y2=0
cc_614 N_B_c_854_n N_VPWR_c_1018_n 0.0115945f $X=6.89 $Y=3.15 $X2=0 $Y2=0
cc_615 N_B_c_836_n N_A_509_347#_c_1132_n 0.00503771f $X=2.865 $Y=3.15 $X2=0
+ $Y2=0
cc_616 N_B_M1019_g N_A_509_347#_c_1137_n 0.0160572f $X=2.955 $Y=2.235 $X2=0
+ $Y2=0
cc_617 N_B_c_843_n N_A_509_347#_c_1137_n 0.0012079f $X=4.92 $Y=3.15 $X2=0 $Y2=0
cc_618 N_B_M1019_g N_A_509_347#_c_1133_n 8.63454e-19 $X=2.955 $Y=2.235 $X2=0
+ $Y2=0
cc_619 N_B_c_843_n N_A_509_347#_c_1133_n 0.00624256f $X=4.92 $Y=3.15 $X2=0 $Y2=0
cc_620 N_B_c_849_n N_A_1107_347#_c_1174_n 0.00572149f $X=6.8 $Y=3.15 $X2=0 $Y2=0
cc_621 N_B_M1001_g N_A_1107_347#_c_1178_n 0.0149337f $X=6.89 $Y=2.31 $X2=0 $Y2=0
cc_622 N_B_c_833_n N_A_1107_347#_c_1178_n 0.00803671f $X=7.305 $Y=1.485 $X2=0
+ $Y2=0
cc_623 N_B_c_832_n N_A_1107_347#_c_1175_n 0.00181486f $X=7.21 $Y=1.527 $X2=0
+ $Y2=0
cc_624 N_B_c_833_n N_A_1107_347#_c_1175_n 0.0280469f $X=7.305 $Y=1.485 $X2=0
+ $Y2=0
cc_625 N_B_M1001_g N_A_1107_347#_c_1176_n 0.00359019f $X=6.89 $Y=2.31 $X2=0
+ $Y2=0
cc_626 N_B_c_831_n N_VGND_c_1221_n 0.00171306f $X=5.01 $Y=1.09 $X2=0 $Y2=0
cc_627 N_B_M1013_g N_VGND_c_1222_n 0.00449178f $X=7.21 $Y=0.695 $X2=0 $Y2=0
cc_628 N_B_M1013_g N_VGND_c_1223_n 0.00562997f $X=7.21 $Y=0.695 $X2=0 $Y2=0
cc_629 N_B_M1025_g N_VGND_c_1225_n 0.00317047f $X=1.5 $Y=0.695 $X2=0 $Y2=0
cc_630 N_B_c_830_n N_VGND_c_1225_n 0.00313877f $X=2.955 $Y=1.09 $X2=0 $Y2=0
cc_631 N_B_c_831_n N_VGND_c_1226_n 0.00432196f $X=5.01 $Y=1.09 $X2=0 $Y2=0
cc_632 N_B_M1013_g N_VGND_c_1227_n 0.0032155f $X=7.21 $Y=0.695 $X2=0 $Y2=0
cc_633 N_B_M1025_g N_VGND_c_1229_n 0.00544287f $X=1.5 $Y=0.695 $X2=0 $Y2=0
cc_634 N_B_M1013_g N_VGND_c_1229_n 0.00544287f $X=7.21 $Y=0.695 $X2=0 $Y2=0
cc_635 N_B_c_830_n N_VGND_c_1229_n 0.00544287f $X=2.955 $Y=1.09 $X2=0 $Y2=0
cc_636 N_B_c_831_n N_VGND_c_1229_n 0.00544287f $X=5.01 $Y=1.09 $X2=0 $Y2=0
cc_637 N_B_c_830_n N_VGND_c_1230_n 0.00397421f $X=2.955 $Y=1.09 $X2=0 $Y2=0
cc_638 N_B_c_830_n N_A_501_75#_c_1335_n 0.0088188f $X=2.955 $Y=1.09 $X2=0 $Y2=0
cc_639 N_B_c_830_n N_A_501_75#_c_1332_n 0.00440744f $X=2.955 $Y=1.09 $X2=0 $Y2=0
cc_640 N_B_c_830_n N_A_501_75#_c_1340_n 8.04385e-19 $X=2.955 $Y=1.09 $X2=0 $Y2=0
cc_641 N_B_M1013_g N_A_1100_75#_c_1364_n 0.00140538f $X=7.21 $Y=0.695 $X2=0
+ $Y2=0
cc_642 N_B_M1013_g N_A_1100_75#_c_1374_n 0.0101012f $X=7.21 $Y=0.695 $X2=0 $Y2=0
cc_643 N_B_M1013_g N_A_1100_75#_c_1360_n 0.00493327f $X=7.21 $Y=0.695 $X2=0
+ $Y2=0
cc_644 N_SUM_c_1002_n N_VPWR_c_1019_n 0.0627545f $X=0.27 $Y=1.985 $X2=0 $Y2=0
cc_645 N_SUM_c_1002_n N_VPWR_c_1026_n 0.0119584f $X=0.27 $Y=1.985 $X2=0 $Y2=0
cc_646 N_SUM_c_1002_n N_VPWR_c_1018_n 0.00989813f $X=0.27 $Y=1.985 $X2=0 $Y2=0
cc_647 SUM N_VGND_c_1224_n 0.0135716f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_648 SUM N_VGND_c_1229_n 0.0102675f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_649 N_VPWR_c_1020_n N_A_509_347#_c_1132_n 0.00129215f $X=3.245 $Y=2.795 $X2=0
+ $Y2=0
cc_650 N_VPWR_c_1027_n N_A_509_347#_c_1132_n 0.00570949f $X=3.08 $Y=3.33 $X2=0
+ $Y2=0
cc_651 N_VPWR_c_1018_n N_A_509_347#_c_1132_n 0.00688066f $X=8.4 $Y=3.33 $X2=0
+ $Y2=0
cc_652 N_VPWR_M1019_d N_A_509_347#_c_1137_n 0.00723155f $X=3.03 $Y=1.735 $X2=0
+ $Y2=0
cc_653 N_VPWR_c_1020_n N_A_509_347#_c_1137_n 0.0261161f $X=3.245 $Y=2.795 $X2=0
+ $Y2=0
cc_654 N_VPWR_c_1020_n N_A_509_347#_c_1133_n 0.00502133f $X=3.245 $Y=2.795 $X2=0
+ $Y2=0
cc_655 N_VPWR_c_1021_n N_A_509_347#_c_1133_n 0.0172713f $X=4.27 $Y=2.47 $X2=0
+ $Y2=0
cc_656 N_VPWR_c_1024_n N_A_509_347#_c_1133_n 0.0073103f $X=4.105 $Y=3.33 $X2=0
+ $Y2=0
cc_657 N_VPWR_c_1018_n N_A_509_347#_c_1133_n 0.00891228f $X=8.4 $Y=3.33 $X2=0
+ $Y2=0
cc_658 N_VPWR_c_1022_n N_A_1107_347#_c_1174_n 0.0115183f $X=6.66 $Y=2.6 $X2=0
+ $Y2=0
cc_659 N_VPWR_c_1028_n N_A_1107_347#_c_1174_n 0.00650801f $X=6.12 $Y=3.33 $X2=0
+ $Y2=0
cc_660 N_VPWR_c_1018_n N_A_1107_347#_c_1174_n 0.00784572f $X=8.4 $Y=3.33 $X2=0
+ $Y2=0
cc_661 N_VPWR_M1022_d N_A_1107_347#_c_1178_n 0.021929f $X=6.13 $Y=1.735 $X2=0
+ $Y2=0
cc_662 N_VPWR_c_1022_n N_A_1107_347#_c_1178_n 0.0363925f $X=6.66 $Y=2.6 $X2=0
+ $Y2=0
cc_663 N_VPWR_c_1023_n N_A_1107_347#_c_1175_n 0.0137241f $X=7.92 $Y=1.985 $X2=0
+ $Y2=0
cc_664 N_VPWR_c_1022_n N_A_1107_347#_c_1176_n 0.0143566f $X=6.66 $Y=2.6 $X2=0
+ $Y2=0
cc_665 N_VPWR_c_1023_n N_A_1107_347#_c_1176_n 0.0249394f $X=7.92 $Y=1.985 $X2=0
+ $Y2=0
cc_666 N_VPWR_c_1029_n N_A_1107_347#_c_1176_n 0.0087946f $X=7.755 $Y=3.33 $X2=0
+ $Y2=0
cc_667 N_VPWR_c_1018_n N_A_1107_347#_c_1176_n 0.0106389f $X=8.4 $Y=3.33 $X2=0
+ $Y2=0
cc_668 N_VPWR_c_1023_n COUT 0.0779559f $X=7.92 $Y=1.985 $X2=0 $Y2=0
cc_669 N_VPWR_c_1030_n COUT 0.0112891f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_670 N_VPWR_c_1018_n COUT 0.00934413f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_671 COUT N_VGND_c_1223_n 0.0157813f $X=8.315 $Y=0.47 $X2=0 $Y2=0
cc_672 COUT N_VGND_c_1228_n 0.0145639f $X=8.315 $Y=0.47 $X2=0 $Y2=0
cc_673 COUT N_VGND_c_1229_n 0.0119984f $X=8.315 $Y=0.47 $X2=0 $Y2=0
cc_674 COUT N_A_1100_75#_c_1360_n 0.0011882f $X=8.315 $Y=0.47 $X2=0 $Y2=0
cc_675 N_VGND_M1012_d N_A_501_75#_c_1335_n 0.00734279f $X=3.015 $Y=0.375 $X2=0
+ $Y2=0
cc_676 N_VGND_c_1220_n N_A_501_75#_c_1335_n 0.0029521f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_677 N_VGND_c_1225_n N_A_501_75#_c_1335_n 0.00294479f $X=3.07 $Y=0 $X2=0 $Y2=0
cc_678 N_VGND_c_1229_n N_A_501_75#_c_1335_n 0.0111994f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_679 N_VGND_c_1230_n N_A_501_75#_c_1335_n 0.0243979f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_680 N_VGND_c_1225_n N_A_501_75#_c_1332_n 0.0114153f $X=3.07 $Y=0 $X2=0 $Y2=0
cc_681 N_VGND_c_1229_n N_A_501_75#_c_1332_n 0.01383f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_682 N_VGND_c_1220_n N_A_501_75#_c_1340_n 0.00882747f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_683 N_VGND_c_1229_n N_A_501_75#_c_1340_n 0.0110304f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_684 N_VGND_c_1229_n N_A_1100_75#_M1020_d 0.00738975f $X=8.4 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_685 N_VGND_M1018_d N_A_1100_75#_c_1359_n 4.88898e-19 $X=6.56 $Y=0.375 $X2=0
+ $Y2=0
cc_686 N_VGND_c_1222_n N_A_1100_75#_c_1359_n 0.014412f $X=6.915 $Y=0.305 $X2=0
+ $Y2=0
cc_687 N_VGND_c_1226_n N_A_1100_75#_c_1359_n 0.0709494f $X=6.83 $Y=0 $X2=0 $Y2=0
cc_688 N_VGND_c_1229_n N_A_1100_75#_c_1359_n 0.0410407f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_689 N_VGND_M1018_d N_A_1100_75#_c_1364_n 0.00300659f $X=6.56 $Y=0.375 $X2=0
+ $Y2=0
cc_690 N_VGND_c_1222_n N_A_1100_75#_c_1364_n 0.00332933f $X=6.915 $Y=0.305 $X2=0
+ $Y2=0
cc_691 N_VGND_M1018_d N_A_1100_75#_c_1374_n 0.0116084f $X=6.56 $Y=0.375 $X2=0
+ $Y2=0
cc_692 N_VGND_c_1222_n N_A_1100_75#_c_1374_n 0.0188598f $X=6.915 $Y=0.305 $X2=0
+ $Y2=0
cc_693 N_VGND_c_1226_n N_A_1100_75#_c_1374_n 0.00291923f $X=6.83 $Y=0 $X2=0
+ $Y2=0
cc_694 N_VGND_c_1227_n N_A_1100_75#_c_1374_n 0.0025393f $X=7.78 $Y=0 $X2=0 $Y2=0
cc_695 N_VGND_c_1229_n N_A_1100_75#_c_1374_n 0.0105139f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_696 N_VGND_M1018_d N_A_1100_75#_c_1365_n 4.74072e-19 $X=6.56 $Y=0.375 $X2=0
+ $Y2=0
cc_697 N_VGND_c_1223_n N_A_1100_75#_c_1360_n 0.0218711f $X=7.945 $Y=0.605 $X2=0
+ $Y2=0
cc_698 N_VGND_c_1227_n N_A_1100_75#_c_1360_n 0.00810949f $X=7.78 $Y=0 $X2=0
+ $Y2=0
cc_699 N_VGND_c_1229_n N_A_1100_75#_c_1360_n 0.0106855f $X=8.4 $Y=0 $X2=0 $Y2=0
