* File: sky130_fd_sc_ls__o31a_4.pex.spice
* Created: Fri Aug 28 13:53:00 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__O31A_4%A_86_260# 1 2 3 10 12 15 17 18 21 23 25 28 30
+ 32 35 37 39 42 49 53 56 58 60 64 68 70 72
c138 68 0 2.04502e-19 $X=2.465 $Y=1.3
c139 64 0 2.82748e-19 $X=3.105 $Y=0.77
c140 58 0 1.70893e-19 $X=2.94 $Y=1.215
c141 53 0 1.74626e-19 $X=2.63 $Y=2.105
c142 35 0 1.6164e-19 $X=1.83 $Y=0.74
r143 77 78 50.1574 $w=3.94e-07 $l=4.1e-07 $layer=POLY_cond $X=1.42 $Y=1.532
+ $X2=1.83 $Y2=1.532
r144 76 77 2.4467 $w=3.94e-07 $l=2e-08 $layer=POLY_cond $X=1.4 $Y=1.532 $X2=1.42
+ $Y2=1.532
r145 73 74 1.83503 $w=3.94e-07 $l=1.5e-08 $layer=POLY_cond $X=0.955 $Y=1.532
+ $X2=0.97 $Y2=1.532
r146 62 64 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=3.105 $Y=1.13
+ $X2=3.105 $Y2=0.77
r147 61 70 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.715 $Y=2.46
+ $X2=2.59 $Y2=2.46
r148 60 72 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.925 $Y=2.46
+ $X2=4.09 $Y2=2.46
r149 60 61 78.9412 $w=1.68e-07 $l=1.21e-06 $layer=LI1_cond $X=3.925 $Y=2.46
+ $X2=2.715 $Y2=2.46
r150 59 68 5.16603 $w=2.5e-07 $l=2.89396e-07 $layer=LI1_cond $X=2.715 $Y=1.215
+ $X2=2.465 $Y2=1.3
r151 58 62 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.94 $Y=1.215
+ $X2=3.105 $Y2=1.13
r152 58 59 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.94 $Y=1.215
+ $X2=2.715 $Y2=1.215
r153 54 70 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.59 $Y=2.545
+ $X2=2.59 $Y2=2.46
r154 54 56 12.4464 $w=2.48e-07 $l=2.7e-07 $layer=LI1_cond $X=2.59 $Y=2.545
+ $X2=2.59 $Y2=2.815
r155 51 70 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.59 $Y=2.375
+ $X2=2.59 $Y2=2.46
r156 51 53 12.4464 $w=2.48e-07 $l=2.7e-07 $layer=LI1_cond $X=2.59 $Y=2.375
+ $X2=2.59 $Y2=2.105
r157 50 68 1.34256 $w=2.5e-07 $l=3.87492e-07 $layer=LI1_cond $X=2.59 $Y=1.63
+ $X2=2.465 $Y2=1.3
r158 50 53 21.8964 $w=2.48e-07 $l=4.75e-07 $layer=LI1_cond $X=2.59 $Y=1.63
+ $X2=2.59 $Y2=2.105
r159 49 80 2.4467 $w=3.94e-07 $l=2e-08 $layer=POLY_cond $X=1.85 $Y=1.532
+ $X2=1.87 $Y2=1.532
r160 49 78 2.4467 $w=3.94e-07 $l=2e-08 $layer=POLY_cond $X=1.85 $Y=1.532
+ $X2=1.83 $Y2=1.532
r161 48 49 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.85
+ $Y=1.465 $X2=1.85 $Y2=1.465
r162 45 76 28.1371 $w=3.94e-07 $l=2.3e-07 $layer=POLY_cond $X=1.17 $Y=1.532
+ $X2=1.4 $Y2=1.532
r163 45 74 24.467 $w=3.94e-07 $l=2e-07 $layer=POLY_cond $X=1.17 $Y=1.532
+ $X2=0.97 $Y2=1.532
r164 44 48 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.17 $Y=1.465
+ $X2=1.85 $Y2=1.465
r165 44 45 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.17
+ $Y=1.465 $X2=1.17 $Y2=1.465
r166 42 68 5.16603 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=2.465 $Y=1.465
+ $X2=2.465 $Y2=1.3
r167 42 48 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=2.465 $Y=1.465
+ $X2=1.85 $Y2=1.465
r168 37 80 25.4929 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=1.87 $Y=1.765
+ $X2=1.87 $Y2=1.532
r169 37 39 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.87 $Y=1.765
+ $X2=1.87 $Y2=2.4
r170 33 78 25.4929 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=1.83 $Y=1.3
+ $X2=1.83 $Y2=1.532
r171 33 35 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.83 $Y=1.3
+ $X2=1.83 $Y2=0.74
r172 30 77 25.4929 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=1.42 $Y=1.765
+ $X2=1.42 $Y2=1.532
r173 30 32 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.42 $Y=1.765
+ $X2=1.42 $Y2=2.4
r174 26 76 25.4929 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=1.4 $Y=1.3 $X2=1.4
+ $Y2=1.532
r175 26 28 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.4 $Y=1.3 $X2=1.4
+ $Y2=0.74
r176 23 74 25.4929 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=0.97 $Y=1.765
+ $X2=0.97 $Y2=1.532
r177 23 25 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.97 $Y=1.765
+ $X2=0.97 $Y2=2.4
r178 19 73 25.4929 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=0.955 $Y=1.3
+ $X2=0.955 $Y2=1.532
r179 19 21 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.955 $Y=1.3
+ $X2=0.955 $Y2=0.74
r180 18 41 48.795 $w=1.8e-07 $l=1.2e-07 $layer=POLY_cond $X=0.52 $Y=1.42
+ $X2=0.52 $Y2=1.3
r181 17 73 16.4864 $w=3.94e-07 $l=1.4472e-07 $layer=POLY_cond $X=0.88 $Y=1.42
+ $X2=0.955 $Y2=1.532
r182 17 18 69.8776 $w=2.4e-07 $l=2.7e-07 $layer=POLY_cond $X=0.88 $Y=1.42
+ $X2=0.61 $Y2=1.42
r183 15 41 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.525 $Y=0.74
+ $X2=0.525 $Y2=1.3
r184 10 18 136.255 $w=1.8e-07 $l=3.45e-07 $layer=POLY_cond $X=0.52 $Y=1.765
+ $X2=0.52 $Y2=1.42
r185 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.52 $Y=1.765
+ $X2=0.52 $Y2=2.4
r186 3 72 300 $w=1.7e-07 $l=5.70088e-07 $layer=licon1_PDIFF $count=2 $X=3.94
+ $Y=1.96 $X2=4.09 $Y2=2.46
r187 2 70 600 $w=1.7e-07 $l=5.70088e-07 $layer=licon1_PDIFF $count=1 $X=2.48
+ $Y=1.96 $X2=2.63 $Y2=2.46
r188 2 56 600 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=2.48
+ $Y=1.96 $X2=2.63 $Y2=2.815
r189 2 53 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.48
+ $Y=1.96 $X2=2.63 $Y2=2.105
r190 1 64 91 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_NDIFF $count=2 $X=2.915
+ $Y=0.625 $X2=3.105 $Y2=0.77
.ends

.subckt PM_SKY130_FD_SC_LS__O31A_4%B1 2 3 5 6 7 10 12 14 17 19 20 26
c64 26 0 1.00449e-19 $X=3.07 $Y=1.635
c65 10 0 3.30533e-19 $X=2.84 $Y=0.945
c66 3 0 7.94108e-20 $X=2.405 $Y=1.885
c67 2 0 1.04054e-19 $X=2.405 $Y=1.795
r68 26 28 34.0395 $w=3.54e-07 $l=2.5e-07 $layer=POLY_cond $X=3.07 $Y=1.677
+ $X2=3.32 $Y2=1.677
r69 24 26 29.274 $w=3.54e-07 $l=2.15e-07 $layer=POLY_cond $X=2.855 $Y=1.677
+ $X2=3.07 $Y2=1.677
r70 23 24 2.04237 $w=3.54e-07 $l=1.5e-08 $layer=POLY_cond $X=2.84 $Y=1.677
+ $X2=2.855 $Y2=1.677
r71 19 20 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=3.07 $Y=1.635 $X2=3.07
+ $Y2=2.035
r72 19 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.07
+ $Y=1.635 $X2=3.07 $Y2=1.635
r73 15 28 22.9014 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.32 $Y=1.47
+ $X2=3.32 $Y2=1.677
r74 15 17 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=3.32 $Y=1.47
+ $X2=3.32 $Y2=0.945
r75 12 24 22.9014 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.855 $Y=1.885
+ $X2=2.855 $Y2=1.677
r76 12 14 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.855 $Y=1.885
+ $X2=2.855 $Y2=2.46
r77 8 23 22.9014 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.84 $Y=1.47
+ $X2=2.84 $Y2=1.677
r78 8 10 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=2.84 $Y=1.47
+ $X2=2.84 $Y2=0.945
r79 6 23 26.5778 $w=3.54e-07 $l=1.653e-07 $layer=POLY_cond $X=2.765 $Y=1.545
+ $X2=2.84 $Y2=1.677
r80 6 7 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.765 $Y=1.545
+ $X2=2.495 $Y2=1.545
r81 3 5 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.405 $Y=1.885
+ $X2=2.405 $Y2=2.46
r82 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.405 $Y=1.795 $X2=2.405
+ $Y2=1.885
r83 1 7 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=2.405 $Y=1.62
+ $X2=2.495 $Y2=1.545
r84 1 2 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=2.405 $Y=1.62
+ $X2=2.405 $Y2=1.795
.ends

.subckt PM_SKY130_FD_SC_LS__O31A_4%A3 1 3 6 8 10 13 15 16 17 18 28
c55 8 0 1.50942e-19 $X=4.315 $Y=1.885
c56 6 0 2.84737e-19 $X=3.91 $Y=0.945
r57 28 29 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=4.315 $Y=1.67
+ $X2=4.34 $Y2=1.67
r58 26 28 9.51316 $w=3.8e-07 $l=7.5e-08 $layer=POLY_cond $X=4.24 $Y=1.67
+ $X2=4.315 $Y2=1.67
r59 26 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.24
+ $Y=1.62 $X2=4.24 $Y2=1.62
r60 24 26 41.8579 $w=3.8e-07 $l=3.3e-07 $layer=POLY_cond $X=3.91 $Y=1.67
+ $X2=4.24 $Y2=1.67
r61 23 24 5.70789 $w=3.8e-07 $l=4.5e-08 $layer=POLY_cond $X=3.865 $Y=1.67
+ $X2=3.91 $Y2=1.67
r62 17 18 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=4.56 $Y=1.62
+ $X2=5.04 $Y2=1.62
r63 17 27 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=4.56 $Y=1.62
+ $X2=4.24 $Y2=1.62
r64 16 27 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=4.08 $Y=1.62 $X2=4.24
+ $Y2=1.62
r65 15 16 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=3.6 $Y=1.62 $X2=4.08
+ $Y2=1.62
r66 11 29 24.6126 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=4.34 $Y=1.455
+ $X2=4.34 $Y2=1.67
r67 11 13 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=4.34 $Y=1.455
+ $X2=4.34 $Y2=0.945
r68 8 28 24.6126 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=4.315 $Y=1.885
+ $X2=4.315 $Y2=1.67
r69 8 10 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=4.315 $Y=1.885
+ $X2=4.315 $Y2=2.46
r70 4 24 24.6126 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=3.91 $Y=1.455
+ $X2=3.91 $Y2=1.67
r71 4 6 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=3.91 $Y=1.455 $X2=3.91
+ $Y2=0.945
r72 1 23 24.6126 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=3.865 $Y=1.885
+ $X2=3.865 $Y2=1.67
r73 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.865 $Y=1.885
+ $X2=3.865 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_LS__O31A_4%A1 3 5 7 10 12 14 15 21 22
c52 22 0 1.91258e-19 $X=5.71 $Y=1.62
c53 10 0 1.6294e-19 $X=5.7 $Y=0.945
r54 21 23 0.637566 $w=3.78e-07 $l=5e-09 $layer=POLY_cond $X=5.71 $Y=1.67
+ $X2=5.715 $Y2=1.67
r55 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.71
+ $Y=1.62 $X2=5.71 $Y2=1.62
r56 19 21 1.27513 $w=3.78e-07 $l=1e-08 $layer=POLY_cond $X=5.7 $Y=1.67 $X2=5.71
+ $Y2=1.67
r57 18 19 61.8439 $w=3.78e-07 $l=4.85e-07 $layer=POLY_cond $X=5.215 $Y=1.67
+ $X2=5.7 $Y2=1.67
r58 17 18 1.9127 $w=3.78e-07 $l=1.5e-08 $layer=POLY_cond $X=5.2 $Y=1.67
+ $X2=5.215 $Y2=1.67
r59 15 22 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=5.52 $Y=1.62
+ $X2=5.71 $Y2=1.62
r60 12 23 24.4846 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=5.715 $Y=1.885
+ $X2=5.715 $Y2=1.67
r61 12 14 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.715 $Y=1.885
+ $X2=5.715 $Y2=2.46
r62 8 19 24.4846 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=5.7 $Y=1.455 $X2=5.7
+ $Y2=1.67
r63 8 10 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=5.7 $Y=1.455 $X2=5.7
+ $Y2=0.945
r64 5 18 24.4846 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=5.215 $Y=1.885
+ $X2=5.215 $Y2=1.67
r65 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.215 $Y=1.885
+ $X2=5.215 $Y2=2.46
r66 1 17 24.4846 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=5.2 $Y=1.455 $X2=5.2
+ $Y2=1.67
r67 1 3 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=5.2 $Y=1.455 $X2=5.2
+ $Y2=0.945
.ends

.subckt PM_SKY130_FD_SC_LS__O31A_4%A2 1 2 3 5 9 10 11 15 16 18 20
c61 9 0 1.44963e-19 $X=4.77 $Y=0.945
c62 3 0 1.50942e-19 $X=4.765 $Y=1.885
c63 2 0 1.91258e-19 $X=4.765 $Y=1.795
r64 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.28
+ $Y=1.62 $X2=6.28 $Y2=1.62
r65 20 24 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=6.48 $Y=1.62 $X2=6.28
+ $Y2=1.62
r66 16 23 54.9169 $w=2.95e-07 $l=3.00167e-07 $layer=POLY_cond $X=6.205 $Y=1.885
+ $X2=6.28 $Y2=1.62
r67 16 18 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.205 $Y=1.885
+ $X2=6.205 $Y2=2.46
r68 13 23 38.578 $w=2.95e-07 $l=2.0106e-07 $layer=POLY_cond $X=6.2 $Y=1.455
+ $X2=6.28 $Y2=1.62
r69 13 15 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=6.2 $Y=1.455 $X2=6.2
+ $Y2=0.945
r70 12 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.2 $Y=0.255 $X2=6.2
+ $Y2=0.945
r71 10 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.125 $Y=0.18
+ $X2=6.2 $Y2=0.255
r72 10 11 656.34 $w=1.5e-07 $l=1.28e-06 $layer=POLY_cond $X=6.125 $Y=0.18
+ $X2=4.845 $Y2=0.18
r73 9 19 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=4.77 $Y=0.945
+ $X2=4.77 $Y2=1.34
r74 6 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.77 $Y=0.255
+ $X2=4.845 $Y2=0.18
r75 6 9 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.77 $Y=0.255 $X2=4.77
+ $Y2=0.945
r76 3 5 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=4.765 $Y=1.885
+ $X2=4.765 $Y2=2.46
r77 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=4.765 $Y=1.795 $X2=4.765
+ $Y2=1.885
r78 1 19 36.2738 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=4.765 $Y=1.43 $X2=4.765
+ $Y2=1.34
r79 1 2 141.879 $w=1.8e-07 $l=3.65e-07 $layer=POLY_cond $X=4.765 $Y=1.43
+ $X2=4.765 $Y2=1.795
.ends

.subckt PM_SKY130_FD_SC_LS__O31A_4%VPWR 1 2 3 4 5 16 18 24 28 34 38 41 42 43 49
+ 53 58 68 69 75 78 81
r91 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r92 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r93 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r94 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r95 69 82 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=5.52 $Y2=3.33
r96 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r97 66 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.605 $Y=3.33
+ $X2=5.44 $Y2=3.33
r98 66 68 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=5.605 $Y=3.33
+ $X2=6.48 $Y2=3.33
r99 65 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r100 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r101 62 65 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=5.04 $Y2=3.33
r102 61 64 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=3.6 $Y=3.33
+ $X2=5.04 $Y2=3.33
r103 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r104 59 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.245 $Y=3.33
+ $X2=3.08 $Y2=3.33
r105 59 61 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=3.245 $Y=3.33
+ $X2=3.6 $Y2=3.33
r106 58 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.275 $Y=3.33
+ $X2=5.44 $Y2=3.33
r107 58 64 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=5.275 $Y=3.33
+ $X2=5.04 $Y2=3.33
r108 57 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r109 57 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r110 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r111 54 75 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.26 $Y=3.33
+ $X2=2.135 $Y2=3.33
r112 54 56 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=2.26 $Y=3.33
+ $X2=2.64 $Y2=3.33
r113 53 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.915 $Y=3.33
+ $X2=3.08 $Y2=3.33
r114 53 56 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.915 $Y=3.33
+ $X2=2.64 $Y2=3.33
r115 52 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r116 51 52 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r117 49 75 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.01 $Y=3.33
+ $X2=2.135 $Y2=3.33
r118 49 51 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.01 $Y=3.33
+ $X2=1.68 $Y2=3.33
r119 48 52 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r120 48 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r121 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r122 45 72 3.99177 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.38 $Y=3.33
+ $X2=0.19 $Y2=3.33
r123 45 47 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.38 $Y=3.33
+ $X2=0.72 $Y2=3.33
r124 43 62 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=3.6 $Y2=3.33
r125 43 79 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=3.12 $Y2=3.33
r126 41 47 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1.03 $Y=3.33
+ $X2=0.72 $Y2=3.33
r127 41 42 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.03 $Y=3.33
+ $X2=1.155 $Y2=3.33
r128 40 51 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=1.28 $Y=3.33 $X2=1.68
+ $Y2=3.33
r129 40 42 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.28 $Y=3.33
+ $X2=1.155 $Y2=3.33
r130 36 81 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.44 $Y=3.245
+ $X2=5.44 $Y2=3.33
r131 36 38 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=5.44 $Y=3.245
+ $X2=5.44 $Y2=2.8
r132 32 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.08 $Y=3.245
+ $X2=3.08 $Y2=3.33
r133 32 34 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=3.08 $Y=3.245
+ $X2=3.08 $Y2=2.805
r134 28 31 19.1306 $w=2.48e-07 $l=4.15e-07 $layer=LI1_cond $X=2.135 $Y=1.985
+ $X2=2.135 $Y2=2.4
r135 26 75 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.135 $Y=3.245
+ $X2=2.135 $Y2=3.33
r136 26 31 38.9526 $w=2.48e-07 $l=8.45e-07 $layer=LI1_cond $X=2.135 $Y=3.245
+ $X2=2.135 $Y2=2.4
r137 22 42 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.155 $Y=3.245
+ $X2=1.155 $Y2=3.33
r138 22 24 43.3319 $w=2.48e-07 $l=9.4e-07 $layer=LI1_cond $X=1.155 $Y=3.245
+ $X2=1.155 $Y2=2.305
r139 18 21 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=0.255 $Y=1.985
+ $X2=0.255 $Y2=2.815
r140 16 72 3.1514 $w=2.5e-07 $l=1.12916e-07 $layer=LI1_cond $X=0.255 $Y=3.245
+ $X2=0.19 $Y2=3.33
r141 16 21 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.255 $Y=3.245
+ $X2=0.255 $Y2=2.815
r142 5 38 600 $w=1.7e-07 $l=9.11921e-07 $layer=licon1_PDIFF $count=1 $X=5.29
+ $Y=1.96 $X2=5.44 $Y2=2.8
r143 4 34 600 $w=1.7e-07 $l=9.16938e-07 $layer=licon1_PDIFF $count=1 $X=2.93
+ $Y=1.96 $X2=3.08 $Y2=2.805
r144 3 31 300 $w=1.7e-07 $l=6.30555e-07 $layer=licon1_PDIFF $count=2 $X=1.945
+ $Y=1.84 $X2=2.095 $Y2=2.4
r145 3 28 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.945
+ $Y=1.84 $X2=2.095 $Y2=1.985
r146 2 24 300 $w=1.7e-07 $l=5.34766e-07 $layer=licon1_PDIFF $count=2 $X=1.045
+ $Y=1.84 $X2=1.195 $Y2=2.305
r147 1 21 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.15
+ $Y=1.84 $X2=0.295 $Y2=2.815
r148 1 18 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.15
+ $Y=1.84 $X2=0.295 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_LS__O31A_4%X 1 2 3 4 13 15 19 23 27 28 29 30 31 32 33 50
+ 60
c65 15 0 1.6164e-19 $X=1.45 $Y=1.045
c66 13 0 7.94108e-20 $X=1.48 $Y=1.885
r67 57 60 0.664871 $w=2.58e-07 $l=1.5e-08 $layer=LI1_cond $X=0.705 $Y=1.97
+ $X2=0.705 $Y2=1.985
r68 43 50 1.22229 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=0.74 $Y=0.96
+ $X2=0.74 $Y2=0.925
r69 32 33 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=0.705 $Y=2.405
+ $X2=0.705 $Y2=2.775
r70 31 52 3.58051 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=1.885
+ $X2=0.705 $Y2=1.8
r71 31 57 3.58051 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=1.885
+ $X2=0.705 $Y2=1.97
r72 31 32 15.9569 $w=2.58e-07 $l=3.6e-07 $layer=LI1_cond $X=0.705 $Y=2.045
+ $X2=0.705 $Y2=2.405
r73 31 60 2.65948 $w=2.58e-07 $l=6e-08 $layer=LI1_cond $X=0.705 $Y=2.045
+ $X2=0.705 $Y2=1.985
r74 30 52 5.98384 $w=2.58e-07 $l=1.35e-07 $layer=LI1_cond $X=0.705 $Y=1.665
+ $X2=0.705 $Y2=1.8
r75 29 30 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=0.705 $Y=1.295
+ $X2=0.705 $Y2=1.665
r76 29 51 7.31358 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=0.705 $Y=1.295
+ $X2=0.705 $Y2=1.13
r77 28 43 3.19717 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=0.74 $Y=1.045
+ $X2=0.74 $Y2=0.96
r78 28 51 3.19717 $w=2.95e-07 $l=1.00995e-07 $layer=LI1_cond $X=0.74 $Y=1.045
+ $X2=0.705 $Y2=1.13
r79 28 50 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=0.74 $Y=0.9
+ $X2=0.74 $Y2=0.925
r80 27 28 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=0.74 $Y=0.515
+ $X2=0.74 $Y2=0.9
r81 23 25 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=1.645 $Y=1.985
+ $X2=1.645 $Y2=2.815
r82 21 23 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=1.645 $Y=1.97
+ $X2=1.645 $Y2=1.985
r83 17 19 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=1.575 $Y=0.96
+ $X2=1.575 $Y2=0.515
r84 16 28 3.3845 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.905 $Y=1.045
+ $X2=0.74 $Y2=1.045
r85 15 17 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.45 $Y=1.045
+ $X2=1.575 $Y2=0.96
r86 15 16 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=1.45 $Y=1.045
+ $X2=0.905 $Y2=1.045
r87 14 31 2.90867 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.835 $Y=1.885
+ $X2=0.705 $Y2=1.885
r88 13 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.48 $Y=1.885
+ $X2=1.645 $Y2=1.97
r89 13 14 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=1.48 $Y=1.885
+ $X2=0.835 $Y2=1.885
r90 4 25 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.495
+ $Y=1.84 $X2=1.645 $Y2=2.815
r91 4 23 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.495
+ $Y=1.84 $X2=1.645 $Y2=1.985
r92 3 33 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.84 $X2=0.745 $Y2=2.815
r93 3 60 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.84 $X2=0.745 $Y2=1.985
r94 2 19 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.475
+ $Y=0.37 $X2=1.615 $Y2=0.515
r95 1 27 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.6
+ $Y=0.37 $X2=0.74 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__O31A_4%A_699_392# 1 2 3 10 16 18 20 22 25
c46 16 0 3.01885e-19 $X=4.54 $Y=2.475
r47 20 27 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.44 $Y=2.125 $X2=6.44
+ $Y2=2.04
r48 20 22 24.0965 $w=3.28e-07 $l=6.9e-07 $layer=LI1_cond $X=6.44 $Y=2.125
+ $X2=6.44 $Y2=2.815
r49 19 25 5.16603 $w=2.1e-07 $l=1.2339e-07 $layer=LI1_cond $X=4.645 $Y=2.04
+ $X2=4.54 $Y2=2.08
r50 18 27 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.275 $Y=2.04
+ $X2=6.44 $Y2=2.04
r51 18 19 106.342 $w=1.68e-07 $l=1.63e-06 $layer=LI1_cond $X=6.275 $Y=2.04
+ $X2=4.645 $Y2=2.04
r52 14 25 1.34256 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=4.54 $Y=2.205
+ $X2=4.54 $Y2=2.08
r53 14 16 14.2597 $w=2.08e-07 $l=2.7e-07 $layer=LI1_cond $X=4.54 $Y=2.205
+ $X2=4.54 $Y2=2.475
r54 10 25 5.16603 $w=2.1e-07 $l=1.05e-07 $layer=LI1_cond $X=4.435 $Y=2.08
+ $X2=4.54 $Y2=2.08
r55 10 12 36.6477 $w=2.48e-07 $l=7.95e-07 $layer=LI1_cond $X=4.435 $Y=2.08
+ $X2=3.64 $Y2=2.08
r56 3 27 400 $w=1.7e-07 $l=2.26274e-07 $layer=licon1_PDIFF $count=1 $X=6.28
+ $Y=1.96 $X2=6.44 $Y2=2.12
r57 3 22 400 $w=1.7e-07 $l=9.31571e-07 $layer=licon1_PDIFF $count=1 $X=6.28
+ $Y=1.96 $X2=6.44 $Y2=2.815
r58 2 25 600 $w=1.7e-07 $l=2.22711e-07 $layer=licon1_PDIFF $count=1 $X=4.39
+ $Y=1.96 $X2=4.54 $Y2=2.12
r59 2 16 300 $w=1.7e-07 $l=5.85214e-07 $layer=licon1_PDIFF $count=2 $X=4.39
+ $Y=1.96 $X2=4.54 $Y2=2.475
r60 1 12 600 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_PDIFF $count=1 $X=3.495
+ $Y=1.96 $X2=3.64 $Y2=2.12
.ends

.subckt PM_SKY130_FD_SC_LS__O31A_4%A_968_392# 1 2 7 9 11 18
r25 12 16 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.075 $Y=2.38
+ $X2=4.95 $Y2=2.38
r26 11 18 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.775 $Y=2.38
+ $X2=5.94 $Y2=2.38
r27 11 12 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=5.775 $Y=2.38
+ $X2=5.075 $Y2=2.38
r28 7 16 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.95 $Y=2.465 $X2=4.95
+ $Y2=2.38
r29 7 9 16.1342 $w=2.48e-07 $l=3.5e-07 $layer=LI1_cond $X=4.95 $Y=2.465 $X2=4.95
+ $Y2=2.815
r30 2 18 300 $w=1.7e-07 $l=4.89285e-07 $layer=licon1_PDIFF $count=2 $X=5.79
+ $Y=1.96 $X2=5.94 $Y2=2.38
r31 1 16 600 $w=1.7e-07 $l=4.89285e-07 $layer=licon1_PDIFF $count=1 $X=4.84
+ $Y=1.96 $X2=4.99 $Y2=2.38
r32 1 9 600 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=4.84
+ $Y=1.96 $X2=4.99 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_LS__O31A_4%VGND 1 2 3 4 5 6 19 21 25 29 33 37 41 44 45
+ 47 48 49 55 59 64 74 75 81 84 87
c96 59 0 1.61628e-19 $X=3.96 $Y=0
r97 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r98 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r99 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r100 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r101 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r102 72 75 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6.48
+ $Y2=0
r103 72 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r104 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r105 69 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.15 $Y=0 $X2=4.985
+ $Y2=0
r106 69 71 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=5.15 $Y=0 $X2=5.52
+ $Y2=0
r107 68 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r108 68 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r109 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r110 65 84 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.21 $Y=0 $X2=4.085
+ $Y2=0
r111 65 67 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=4.21 $Y=0 $X2=4.56
+ $Y2=0
r112 64 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.82 $Y=0 $X2=4.985
+ $Y2=0
r113 64 67 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=4.82 $Y=0 $X2=4.56
+ $Y2=0
r114 63 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r115 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r116 60 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.21 $Y=0 $X2=2.045
+ $Y2=0
r117 60 62 90.6845 $w=1.68e-07 $l=1.39e-06 $layer=LI1_cond $X=2.21 $Y=0 $X2=3.6
+ $Y2=0
r118 59 84 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.96 $Y=0 $X2=4.085
+ $Y2=0
r119 59 62 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=3.96 $Y=0 $X2=3.6
+ $Y2=0
r120 58 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r121 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r122 55 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.88 $Y=0 $X2=2.045
+ $Y2=0
r123 55 57 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=1.88 $Y=0 $X2=1.68
+ $Y2=0
r124 54 58 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r125 54 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r126 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r127 51 78 3.97288 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=0.395 $Y=0
+ $X2=0.197 $Y2=0
r128 51 53 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.395 $Y=0
+ $X2=0.72 $Y2=0
r129 49 63 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.36 $Y=0 $X2=3.6
+ $Y2=0
r130 49 82 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=3.36 $Y=0 $X2=2.16
+ $Y2=0
r131 47 71 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=5.75 $Y=0 $X2=5.52
+ $Y2=0
r132 47 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.75 $Y=0 $X2=5.915
+ $Y2=0
r133 46 74 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=6.08 $Y=0 $X2=6.48
+ $Y2=0
r134 46 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.08 $Y=0 $X2=5.915
+ $Y2=0
r135 44 53 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.085 $Y=0
+ $X2=0.72 $Y2=0
r136 44 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.085 $Y=0 $X2=1.17
+ $Y2=0
r137 43 57 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=1.255 $Y=0
+ $X2=1.68 $Y2=0
r138 43 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.255 $Y=0 $X2=1.17
+ $Y2=0
r139 39 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.915 $Y=0.085
+ $X2=5.915 $Y2=0
r140 39 41 24.0965 $w=3.28e-07 $l=6.9e-07 $layer=LI1_cond $X=5.915 $Y=0.085
+ $X2=5.915 $Y2=0.775
r141 35 87 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.985 $Y=0.085
+ $X2=4.985 $Y2=0
r142 35 37 24.0965 $w=3.28e-07 $l=6.9e-07 $layer=LI1_cond $X=4.985 $Y=0.085
+ $X2=4.985 $Y2=0.775
r143 31 84 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.085 $Y=0.085
+ $X2=4.085 $Y2=0
r144 31 33 31.8074 $w=2.48e-07 $l=6.9e-07 $layer=LI1_cond $X=4.085 $Y=0.085
+ $X2=4.085 $Y2=0.775
r145 27 81 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.045 $Y=0.085
+ $X2=2.045 $Y2=0
r146 27 29 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.045 $Y=0.085
+ $X2=2.045 $Y2=0.515
r147 23 45 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.17 $Y=0.085
+ $X2=1.17 $Y2=0
r148 23 25 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=1.17 $Y=0.085
+ $X2=1.17 $Y2=0.57
r149 19 78 3.17028 $w=2.5e-07 $l=1.15888e-07 $layer=LI1_cond $X=0.27 $Y=0.085
+ $X2=0.197 $Y2=0
r150 19 21 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.27 $Y=0.085
+ $X2=0.27 $Y2=0.515
r151 6 41 182 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=1 $X=5.775
+ $Y=0.625 $X2=5.915 $Y2=0.775
r152 5 37 182 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=1 $X=4.845
+ $Y=0.625 $X2=4.985 $Y2=0.775
r153 4 33 182 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=1 $X=3.985
+ $Y=0.625 $X2=4.125 $Y2=0.775
r154 3 29 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.905
+ $Y=0.37 $X2=2.045 $Y2=0.515
r155 2 25 182 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=1 $X=1.03
+ $Y=0.37 $X2=1.17 $Y2=0.57
r156 1 21 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.165
+ $Y=0.37 $X2=0.31 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__O31A_4%A_492_125# 1 2 3 4 5 18 20 21 25 26 27 30 32
+ 36 38 42 44 45
c86 36 0 1.6294e-19 $X=5.485 $Y=0.77
c87 30 0 1.44963e-19 $X=4.555 $Y=0.77
r88 40 42 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=6.415 $Y=1.115
+ $X2=6.415 $Y2=0.77
r89 39 45 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.57 $Y=1.2
+ $X2=5.445 $Y2=1.2
r90 38 40 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.25 $Y=1.2
+ $X2=6.415 $Y2=1.115
r91 38 39 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=6.25 $Y=1.2 $X2=5.57
+ $Y2=1.2
r92 34 45 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.445 $Y=1.115
+ $X2=5.445 $Y2=1.2
r93 34 36 15.9037 $w=2.48e-07 $l=3.45e-07 $layer=LI1_cond $X=5.445 $Y=1.115
+ $X2=5.445 $Y2=0.77
r94 33 44 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.64 $Y=1.2
+ $X2=4.515 $Y2=1.2
r95 32 45 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.32 $Y=1.2
+ $X2=5.445 $Y2=1.2
r96 32 33 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=5.32 $Y=1.2 $X2=4.64
+ $Y2=1.2
r97 28 44 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.515 $Y=1.115
+ $X2=4.515 $Y2=1.2
r98 28 30 15.9037 $w=2.48e-07 $l=3.45e-07 $layer=LI1_cond $X=4.515 $Y=1.115
+ $X2=4.515 $Y2=0.77
r99 26 44 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.39 $Y=1.2
+ $X2=4.515 $Y2=1.2
r100 26 27 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=4.39 $Y=1.2
+ $X2=3.78 $Y2=1.2
r101 23 27 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.615 $Y=1.115
+ $X2=3.78 $Y2=1.2
r102 23 25 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=3.615 $Y=1.115
+ $X2=3.615 $Y2=0.77
r103 22 25 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.615 $Y=0.435
+ $X2=3.615 $Y2=0.77
r104 20 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.45 $Y=0.35
+ $X2=3.615 $Y2=0.435
r105 20 21 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.45 $Y=0.35
+ $X2=2.77 $Y2=0.35
r106 16 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.605 $Y=0.435
+ $X2=2.77 $Y2=0.35
r107 16 18 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=2.605 $Y=0.435
+ $X2=2.605 $Y2=0.78
r108 5 42 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.275
+ $Y=0.625 $X2=6.415 $Y2=0.77
r109 4 36 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=5.275
+ $Y=0.625 $X2=5.485 $Y2=0.77
r110 3 30 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.415
+ $Y=0.625 $X2=4.555 $Y2=0.77
r111 2 25 91 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_NDIFF $count=2 $X=3.395
+ $Y=0.625 $X2=3.615 $Y2=0.77
r112 1 18 182 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=1 $X=2.46
+ $Y=0.625 $X2=2.605 $Y2=0.78
.ends

