* File: sky130_fd_sc_ls__a41o_1.spice
* Created: Fri Aug 28 13:01:10 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__a41o_1.pex.spice"
.subckt sky130_fd_sc_ls__a41o_1  VNB VPB B1 A1 A2 A3 A4 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A4	A4
* A3	A3
* A2	A2
* A1	A1
* B1	B1
* VPB	VPB
* VNB	VNB
MM1006 N_VGND_M1006_d N_A_83_244#_M1006_g N_X_M1006_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1554 AS=0.7104 PD=1.16 PS=3.4 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.9
+ SB=75002.8 A=0.111 P=1.78 MULT=1
MM1010 N_A_83_244#_M1010_d N_B1_M1010_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1554 PD=1.02 PS=1.16 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.5
+ SB=75002.2 A=0.111 P=1.78 MULT=1
MM1003 A_449_74# N_A1_M1003_g N_A_83_244#_M1010_d VNB NSHORT L=0.15 W=0.74
+ AD=0.1184 AS=0.1036 PD=1.06 PS=1.02 NRD=17.016 NRS=0 M=1 R=4.93333 SA=75001.9
+ SB=75001.8 A=0.111 P=1.78 MULT=1
MM1000 A_543_74# N_A2_M1000_g A_449_74# VNB NSHORT L=0.15 W=0.74 AD=0.1554
+ AS=0.1184 PD=1.16 PS=1.06 NRD=25.128 NRS=17.016 M=1 R=4.93333 SA=75002.4
+ SB=75001.4 A=0.111 P=1.78 MULT=1
MM1007 A_657_74# N_A3_M1007_g A_543_74# VNB NSHORT L=0.15 W=0.74 AD=0.1554
+ AS=0.1554 PD=1.16 PS=1.16 NRD=25.128 NRS=25.128 M=1 R=4.93333 SA=75002.9
+ SB=75000.8 A=0.111 P=1.78 MULT=1
MM1011 N_VGND_M1011_d N_A4_M1011_g A_657_74# VNB NSHORT L=0.15 W=0.74 AD=0.2109
+ AS=0.1554 PD=2.05 PS=1.16 NRD=0 NRS=25.128 M=1 R=4.93333 SA=75003.5 SB=75000.2
+ A=0.111 P=1.78 MULT=1
MM1008 N_VPWR_M1008_d N_A_83_244#_M1008_g N_X_M1008_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.3304 PD=2.83 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1005 N_A_354_392#_M1005_d N_B1_M1005_g N_A_83_244#_M1005_s VPB PHIGHVT L=0.15
+ W=1 AD=0.175 AS=0.295 PD=1.35 PS=2.59 NRD=11.8003 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75002.3 A=0.15 P=2.3 MULT=1
MM1009 N_VPWR_M1009_d N_A1_M1009_g N_A_354_392#_M1005_d VPB PHIGHVT L=0.15 W=1
+ AD=0.215 AS=0.175 PD=1.43 PS=1.35 NRD=11.8003 NRS=1.9503 M=1 R=6.66667
+ SA=75000.7 SB=75001.8 A=0.15 P=2.3 MULT=1
MM1001 N_A_354_392#_M1001_d N_A2_M1001_g N_VPWR_M1009_d VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.215 PD=1.3 PS=1.43 NRD=1.9503 NRS=17.73 M=1 R=6.66667 SA=75001.3
+ SB=75001.2 A=0.15 P=2.3 MULT=1
MM1004 N_VPWR_M1004_d N_A3_M1004_g N_A_354_392#_M1001_d VPB PHIGHVT L=0.15 W=1
+ AD=0.21 AS=0.15 PD=1.42 PS=1.3 NRD=11.8003 NRS=1.9503 M=1 R=6.66667 SA=75001.7
+ SB=75000.8 A=0.15 P=2.3 MULT=1
MM1002 N_A_354_392#_M1002_d N_A4_M1002_g N_VPWR_M1004_d VPB PHIGHVT L=0.15 W=1
+ AD=0.295 AS=0.21 PD=2.59 PS=1.42 NRD=1.9503 NRS=15.7403 M=1 R=6.66667
+ SA=75002.3 SB=75000.2 A=0.15 P=2.3 MULT=1
DX12_noxref VNB VPB NWDIODE A=8.742 P=13.12
*
.include "sky130_fd_sc_ls__a41o_1.pxi.spice"
*
.ends
*
*
