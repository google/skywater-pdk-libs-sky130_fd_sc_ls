* File: sky130_fd_sc_ls__clkinv_16.pex.spice
* Created: Fri Aug 28 13:10:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__CLKINV_16%A 3 5 7 10 12 14 17 19 21 24 26 28 31 33
+ 35 38 40 42 43 45 48 52 54 56 57 59 62 64 66 69 71 73 76 78 80 83 85 87 90 92
+ 94 97 99 101 104 108 110 112 113 115 116 118 119 121 122 124 125 127 128 130
+ 131 133 134 136 137 203 207 213 219 225 231 237 243 249 253
c417 203 0 1.31047e-19 $X=10.75 $Y=1.485
c418 83 0 1.88851e-19 $X=5.645 $Y=0.61
c419 48 0 1.6166e-19 $X=3.215 $Y=0.61
r420 250 253 1.84782 $w=2.3e-07 $l=2.88e-06 $layer=MET1_cond $X=7.83 $Y=1.295
+ $X2=10.71 $Y2=1.295
r421 249 253 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=10.71
+ $Y=1.295 $X2=10.71 $Y2=1.295
r422 249 250 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=7.83
+ $Y=1.295 $X2=7.83 $Y2=1.295
r423 244 250 0.718597 $w=2.3e-07 $l=1.12e-06 $layer=MET1_cond $X=6.71 $Y=1.295
+ $X2=7.83 $Y2=1.295
r424 243 244 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.71 $Y=1.295
+ $X2=6.71 $Y2=1.295
r425 237 238 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.76 $Y=1.295
+ $X2=5.76 $Y2=1.295
r426 232 238 0.538948 $w=2.3e-07 $l=8.4e-07 $layer=MET1_cond $X=4.92 $Y=1.295
+ $X2=5.76 $Y2=1.295
r427 231 232 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.92 $Y=1.295
+ $X2=4.92 $Y2=1.295
r428 226 232 0.635188 $w=2.3e-07 $l=9.9e-07 $layer=MET1_cond $X=3.93 $Y=1.295
+ $X2=4.92 $Y2=1.295
r429 225 226 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.93 $Y=1.295
+ $X2=3.93 $Y2=1.295
r430 220 226 0.596692 $w=2.3e-07 $l=9.3e-07 $layer=MET1_cond $X=3 $Y=1.295
+ $X2=3.93 $Y2=1.295
r431 219 220 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3 $Y=1.295 $X2=3
+ $Y2=1.295
r432 214 220 0.622356 $w=2.3e-07 $l=9.7e-07 $layer=MET1_cond $X=2.03 $Y=1.295
+ $X2=3 $Y2=1.295
r433 213 214 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.03 $Y=1.295
+ $X2=2.03 $Y2=1.295
r434 208 214 0.577444 $w=2.3e-07 $l=9e-07 $layer=MET1_cond $X=1.13 $Y=1.295
+ $X2=2.03 $Y2=1.295
r435 207 208 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.13 $Y=1.295
+ $X2=1.13 $Y2=1.295
r436 203 205 32.4188 $w=3.94e-07 $l=2.65e-07 $layer=POLY_cond $X=10.75 $Y=1.542
+ $X2=11.015 $Y2=1.542
r437 201 203 22.632 $w=3.94e-07 $l=1.85e-07 $layer=POLY_cond $X=10.565 $Y=1.542
+ $X2=10.75 $Y2=1.542
r438 200 201 55.0508 $w=3.94e-07 $l=4.5e-07 $layer=POLY_cond $X=10.115 $Y=1.542
+ $X2=10.565 $Y2=1.542
r439 199 200 55.0508 $w=3.94e-07 $l=4.5e-07 $layer=POLY_cond $X=9.665 $Y=1.542
+ $X2=10.115 $Y2=1.542
r440 198 199 55.0508 $w=3.94e-07 $l=4.5e-07 $layer=POLY_cond $X=9.215 $Y=1.542
+ $X2=9.665 $Y2=1.542
r441 197 198 55.0508 $w=3.94e-07 $l=4.5e-07 $layer=POLY_cond $X=8.765 $Y=1.542
+ $X2=9.215 $Y2=1.542
r442 196 197 55.0508 $w=3.94e-07 $l=4.5e-07 $layer=POLY_cond $X=8.315 $Y=1.542
+ $X2=8.765 $Y2=1.542
r443 195 196 55.0508 $w=3.94e-07 $l=4.5e-07 $layer=POLY_cond $X=7.865 $Y=1.542
+ $X2=8.315 $Y2=1.542
r444 194 249 0.683776 $w=3.388e-06 $l=1.9e-07 $layer=LI1_cond $X=9.22 $Y=1.485
+ $X2=9.22 $Y2=1.295
r445 194 203 29.056 $w=1.7e-07 $l=8.5e-07 $layer=licon1_POLY $count=5 $X=10.75
+ $Y=1.485 $X2=10.75 $Y2=1.485
r446 193 195 21.4086 $w=3.94e-07 $l=1.75e-07 $layer=POLY_cond $X=7.69 $Y=1.542
+ $X2=7.865 $Y2=1.542
r447 193 194 29.056 $w=1.7e-07 $l=8.5e-07 $layer=licon1_POLY $count=5 $X=7.69
+ $Y=1.485 $X2=7.69 $Y2=1.485
r448 191 193 33.6421 $w=3.94e-07 $l=2.75e-07 $layer=POLY_cond $X=7.415 $Y=1.542
+ $X2=7.69 $Y2=1.542
r449 190 191 6.11675 $w=3.94e-07 $l=5e-08 $layer=POLY_cond $X=7.365 $Y=1.542
+ $X2=7.415 $Y2=1.542
r450 189 190 52.6041 $w=3.94e-07 $l=4.3e-07 $layer=POLY_cond $X=6.935 $Y=1.542
+ $X2=7.365 $Y2=1.542
r451 188 189 3.67005 $w=3.94e-07 $l=3e-08 $layer=POLY_cond $X=6.905 $Y=1.542
+ $X2=6.935 $Y2=1.542
r452 187 243 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=6.71 $Y=1.485
+ $X2=6.71 $Y2=1.295
r453 186 188 23.8553 $w=3.94e-07 $l=1.95e-07 $layer=POLY_cond $X=6.71 $Y=1.542
+ $X2=6.905 $Y2=1.542
r454 186 187 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.71
+ $Y=1.485 $X2=6.71 $Y2=1.485
r455 184 186 25.0787 $w=3.94e-07 $l=2.05e-07 $layer=POLY_cond $X=6.505 $Y=1.542
+ $X2=6.71 $Y2=1.542
r456 183 184 12.2335 $w=3.94e-07 $l=1e-07 $layer=POLY_cond $X=6.405 $Y=1.542
+ $X2=6.505 $Y2=1.542
r457 182 183 40.3706 $w=3.94e-07 $l=3.3e-07 $layer=POLY_cond $X=6.075 $Y=1.542
+ $X2=6.405 $Y2=1.542
r458 181 182 14.6802 $w=3.94e-07 $l=1.2e-07 $layer=POLY_cond $X=5.955 $Y=1.542
+ $X2=6.075 $Y2=1.542
r459 180 237 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=5.76 $Y=1.485
+ $X2=5.76 $Y2=1.295
r460 179 181 23.8553 $w=3.94e-07 $l=1.95e-07 $layer=POLY_cond $X=5.76 $Y=1.542
+ $X2=5.955 $Y2=1.542
r461 179 180 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.76
+ $Y=1.485 $X2=5.76 $Y2=1.485
r462 177 179 14.0685 $w=3.94e-07 $l=1.15e-07 $layer=POLY_cond $X=5.645 $Y=1.542
+ $X2=5.76 $Y2=1.542
r463 176 177 23.2437 $w=3.94e-07 $l=1.9e-07 $layer=POLY_cond $X=5.455 $Y=1.542
+ $X2=5.645 $Y2=1.542
r464 175 176 29.3604 $w=3.94e-07 $l=2.4e-07 $layer=POLY_cond $X=5.215 $Y=1.542
+ $X2=5.455 $Y2=1.542
r465 174 175 25.6904 $w=3.94e-07 $l=2.1e-07 $layer=POLY_cond $X=5.005 $Y=1.542
+ $X2=5.215 $Y2=1.542
r466 173 231 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=4.92 $Y=1.485
+ $X2=4.92 $Y2=1.295
r467 172 174 10.3985 $w=3.94e-07 $l=8.5e-08 $layer=POLY_cond $X=4.92 $Y=1.542
+ $X2=5.005 $Y2=1.542
r468 172 173 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.92
+ $Y=1.485 $X2=4.92 $Y2=1.485
r469 170 172 33.6421 $w=3.94e-07 $l=2.75e-07 $layer=POLY_cond $X=4.645 $Y=1.542
+ $X2=4.92 $Y2=1.542
r470 169 170 11.0102 $w=3.94e-07 $l=9e-08 $layer=POLY_cond $X=4.555 $Y=1.542
+ $X2=4.645 $Y2=1.542
r471 168 169 41.5939 $w=3.94e-07 $l=3.4e-07 $layer=POLY_cond $X=4.215 $Y=1.542
+ $X2=4.555 $Y2=1.542
r472 167 168 13.4569 $w=3.94e-07 $l=1.1e-07 $layer=POLY_cond $X=4.105 $Y=1.542
+ $X2=4.215 $Y2=1.542
r473 166 225 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=3.93 $Y=1.485
+ $X2=3.93 $Y2=1.295
r474 165 167 21.4086 $w=3.94e-07 $l=1.75e-07 $layer=POLY_cond $X=3.93 $Y=1.542
+ $X2=4.105 $Y2=1.542
r475 165 166 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.93
+ $Y=1.485 $X2=3.93 $Y2=1.485
r476 163 165 33.6421 $w=3.94e-07 $l=2.75e-07 $layer=POLY_cond $X=3.655 $Y=1.542
+ $X2=3.93 $Y2=1.542
r477 162 163 1.22335 $w=3.94e-07 $l=1e-08 $layer=POLY_cond $X=3.645 $Y=1.542
+ $X2=3.655 $Y2=1.542
r478 161 162 52.6041 $w=3.94e-07 $l=4.3e-07 $layer=POLY_cond $X=3.215 $Y=1.542
+ $X2=3.645 $Y2=1.542
r479 160 161 1.22335 $w=3.94e-07 $l=1e-08 $layer=POLY_cond $X=3.205 $Y=1.542
+ $X2=3.215 $Y2=1.542
r480 159 219 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=3 $Y=1.485 $X2=3
+ $Y2=1.295
r481 158 160 25.0787 $w=3.94e-07 $l=2.05e-07 $layer=POLY_cond $X=3 $Y=1.542
+ $X2=3.205 $Y2=1.542
r482 158 159 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3
+ $Y=1.485 $X2=3 $Y2=1.485
r483 156 158 29.9721 $w=3.94e-07 $l=2.45e-07 $layer=POLY_cond $X=2.755 $Y=1.542
+ $X2=3 $Y2=1.542
r484 155 156 4.8934 $w=3.94e-07 $l=4e-08 $layer=POLY_cond $X=2.715 $Y=1.542
+ $X2=2.755 $Y2=1.542
r485 154 155 50.1574 $w=3.94e-07 $l=4.1e-07 $layer=POLY_cond $X=2.305 $Y=1.542
+ $X2=2.715 $Y2=1.542
r486 153 154 2.4467 $w=3.94e-07 $l=2e-08 $layer=POLY_cond $X=2.285 $Y=1.542
+ $X2=2.305 $Y2=1.542
r487 152 213 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=2.03 $Y=1.485
+ $X2=2.03 $Y2=1.295
r488 151 153 31.1954 $w=3.94e-07 $l=2.55e-07 $layer=POLY_cond $X=2.03 $Y=1.542
+ $X2=2.285 $Y2=1.542
r489 151 152 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.03
+ $Y=1.485 $X2=2.03 $Y2=1.485
r490 149 151 21.4086 $w=3.94e-07 $l=1.75e-07 $layer=POLY_cond $X=1.855 $Y=1.542
+ $X2=2.03 $Y2=1.542
r491 148 149 8.56345 $w=3.94e-07 $l=7e-08 $layer=POLY_cond $X=1.785 $Y=1.542
+ $X2=1.855 $Y2=1.542
r492 147 148 46.4873 $w=3.94e-07 $l=3.8e-07 $layer=POLY_cond $X=1.405 $Y=1.542
+ $X2=1.785 $Y2=1.542
r493 146 147 6.11675 $w=3.94e-07 $l=5e-08 $layer=POLY_cond $X=1.355 $Y=1.542
+ $X2=1.405 $Y2=1.542
r494 145 207 6.84263 $w=3.18e-07 $l=1.9e-07 $layer=LI1_cond $X=1.135 $Y=1.485
+ $X2=1.135 $Y2=1.295
r495 144 146 27.5254 $w=3.94e-07 $l=2.25e-07 $layer=POLY_cond $X=1.13 $Y=1.542
+ $X2=1.355 $Y2=1.542
r496 144 145 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.13
+ $Y=1.485 $X2=1.13 $Y2=1.485
r497 142 144 21.4086 $w=3.94e-07 $l=1.75e-07 $layer=POLY_cond $X=0.955 $Y=1.542
+ $X2=1.13 $Y2=1.542
r498 141 142 3.67005 $w=3.94e-07 $l=3e-08 $layer=POLY_cond $X=0.925 $Y=1.542
+ $X2=0.955 $Y2=1.542
r499 140 141 51.3807 $w=3.94e-07 $l=4.2e-07 $layer=POLY_cond $X=0.505 $Y=1.542
+ $X2=0.925 $Y2=1.542
r500 139 140 1.22335 $w=3.94e-07 $l=1e-08 $layer=POLY_cond $X=0.495 $Y=1.542
+ $X2=0.505 $Y2=1.542
r501 137 244 0.481203 $w=2.3e-07 $l=7.5e-07 $layer=MET1_cond $X=5.96 $Y=1.295
+ $X2=6.71 $Y2=1.295
r502 137 238 0.128321 $w=2.3e-07 $l=2e-07 $layer=MET1_cond $X=5.96 $Y=1.295
+ $X2=5.76 $Y2=1.295
r503 134 205 25.4929 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=11.015 $Y=1.765
+ $X2=11.015 $Y2=1.542
r504 134 136 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=11.015 $Y=1.765
+ $X2=11.015 $Y2=2.4
r505 131 201 25.4929 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=10.565 $Y=1.765
+ $X2=10.565 $Y2=1.542
r506 131 133 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=10.565 $Y=1.765
+ $X2=10.565 $Y2=2.4
r507 128 200 25.4929 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=10.115 $Y=1.765
+ $X2=10.115 $Y2=1.542
r508 128 130 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=10.115 $Y=1.765
+ $X2=10.115 $Y2=2.4
r509 125 199 25.4929 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=9.665 $Y=1.765
+ $X2=9.665 $Y2=1.542
r510 125 127 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=9.665 $Y=1.765
+ $X2=9.665 $Y2=2.4
r511 122 198 25.4929 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=9.215 $Y=1.765
+ $X2=9.215 $Y2=1.542
r512 122 124 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=9.215 $Y=1.765
+ $X2=9.215 $Y2=2.4
r513 119 197 25.4929 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=8.765 $Y=1.765
+ $X2=8.765 $Y2=1.542
r514 119 121 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.765 $Y=1.765
+ $X2=8.765 $Y2=2.4
r515 116 196 25.4929 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=8.315 $Y=1.765
+ $X2=8.315 $Y2=1.542
r516 116 118 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.315 $Y=1.765
+ $X2=8.315 $Y2=2.4
r517 113 195 25.4929 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=7.865 $Y=1.765
+ $X2=7.865 $Y2=1.542
r518 113 115 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.865 $Y=1.765
+ $X2=7.865 $Y2=2.4
r519 110 191 25.4929 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=7.415 $Y=1.765
+ $X2=7.415 $Y2=1.542
r520 110 112 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.415 $Y=1.765
+ $X2=7.415 $Y2=2.4
r521 106 190 25.4929 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=7.365 $Y=1.32
+ $X2=7.365 $Y2=1.542
r522 106 108 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=7.365 $Y=1.32
+ $X2=7.365 $Y2=0.61
r523 102 189 25.4929 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=6.935 $Y=1.32
+ $X2=6.935 $Y2=1.542
r524 102 104 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=6.935 $Y=1.32
+ $X2=6.935 $Y2=0.61
r525 99 188 25.4929 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=6.905 $Y=1.765
+ $X2=6.905 $Y2=1.542
r526 99 101 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.905 $Y=1.765
+ $X2=6.905 $Y2=2.4
r527 95 184 25.4929 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=6.505 $Y=1.32
+ $X2=6.505 $Y2=1.542
r528 95 97 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=6.505 $Y=1.32
+ $X2=6.505 $Y2=0.61
r529 92 183 25.4929 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=6.405 $Y=1.765
+ $X2=6.405 $Y2=1.542
r530 92 94 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.405 $Y=1.765
+ $X2=6.405 $Y2=2.4
r531 88 182 25.4929 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=6.075 $Y=1.32
+ $X2=6.075 $Y2=1.542
r532 88 90 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=6.075 $Y=1.32
+ $X2=6.075 $Y2=0.61
r533 85 181 25.4929 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=5.955 $Y=1.765
+ $X2=5.955 $Y2=1.542
r534 85 87 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.955 $Y=1.765
+ $X2=5.955 $Y2=2.4
r535 81 177 25.4929 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=5.645 $Y=1.32
+ $X2=5.645 $Y2=1.542
r536 81 83 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=5.645 $Y=1.32
+ $X2=5.645 $Y2=0.61
r537 78 176 25.4929 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=5.455 $Y=1.765
+ $X2=5.455 $Y2=1.542
r538 78 80 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.455 $Y=1.765
+ $X2=5.455 $Y2=2.4
r539 74 175 25.4929 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=5.215 $Y=1.32
+ $X2=5.215 $Y2=1.542
r540 74 76 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=5.215 $Y=1.32
+ $X2=5.215 $Y2=0.61
r541 71 174 25.4929 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=5.005 $Y=1.765
+ $X2=5.005 $Y2=1.542
r542 71 73 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.005 $Y=1.765
+ $X2=5.005 $Y2=2.4
r543 67 170 25.4929 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=4.645 $Y=1.32
+ $X2=4.645 $Y2=1.542
r544 67 69 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=4.645 $Y=1.32
+ $X2=4.645 $Y2=0.61
r545 64 169 25.4929 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=4.555 $Y=1.765
+ $X2=4.555 $Y2=1.542
r546 64 66 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.555 $Y=1.765
+ $X2=4.555 $Y2=2.4
r547 60 168 25.4929 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=4.215 $Y=1.32
+ $X2=4.215 $Y2=1.542
r548 60 62 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=4.215 $Y=1.32
+ $X2=4.215 $Y2=0.61
r549 57 167 25.4929 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=4.105 $Y=1.765
+ $X2=4.105 $Y2=1.542
r550 57 59 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.105 $Y=1.765
+ $X2=4.105 $Y2=2.4
r551 54 163 25.4929 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=3.655 $Y=1.765
+ $X2=3.655 $Y2=1.542
r552 54 56 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.655 $Y=1.765
+ $X2=3.655 $Y2=2.4
r553 50 162 25.4929 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=3.645 $Y=1.32
+ $X2=3.645 $Y2=1.542
r554 50 52 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=3.645 $Y=1.32
+ $X2=3.645 $Y2=0.61
r555 46 161 25.4929 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=3.215 $Y=1.32
+ $X2=3.215 $Y2=1.542
r556 46 48 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=3.215 $Y=1.32
+ $X2=3.215 $Y2=0.61
r557 43 160 25.4929 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=3.205 $Y=1.765
+ $X2=3.205 $Y2=1.542
r558 43 45 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.205 $Y=1.765
+ $X2=3.205 $Y2=2.4
r559 40 156 25.4929 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=2.755 $Y=1.765
+ $X2=2.755 $Y2=1.542
r560 40 42 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.755 $Y=1.765
+ $X2=2.755 $Y2=2.4
r561 36 155 25.4929 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=2.715 $Y=1.32
+ $X2=2.715 $Y2=1.542
r562 36 38 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=2.715 $Y=1.32
+ $X2=2.715 $Y2=0.61
r563 33 154 25.4929 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=2.305 $Y=1.765
+ $X2=2.305 $Y2=1.542
r564 33 35 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.305 $Y=1.765
+ $X2=2.305 $Y2=2.4
r565 29 153 25.4929 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=2.285 $Y=1.32
+ $X2=2.285 $Y2=1.542
r566 29 31 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=2.285 $Y=1.32
+ $X2=2.285 $Y2=0.61
r567 26 149 25.4929 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=1.855 $Y=1.765
+ $X2=1.855 $Y2=1.542
r568 26 28 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.855 $Y=1.765
+ $X2=1.855 $Y2=2.4
r569 22 148 25.4929 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=1.785 $Y=1.32
+ $X2=1.785 $Y2=1.542
r570 22 24 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.785 $Y=1.32
+ $X2=1.785 $Y2=0.61
r571 19 147 25.4929 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=1.405 $Y=1.765
+ $X2=1.405 $Y2=1.542
r572 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.405 $Y=1.765
+ $X2=1.405 $Y2=2.4
r573 15 146 25.4929 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=1.355 $Y=1.32
+ $X2=1.355 $Y2=1.542
r574 15 17 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.355 $Y=1.32
+ $X2=1.355 $Y2=0.61
r575 12 142 25.4929 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=0.955 $Y=1.765
+ $X2=0.955 $Y2=1.542
r576 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.955 $Y=1.765
+ $X2=0.955 $Y2=2.4
r577 8 141 25.4929 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=0.925 $Y=1.32
+ $X2=0.925 $Y2=1.542
r578 8 10 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=0.925 $Y=1.32
+ $X2=0.925 $Y2=0.61
r579 5 140 25.4929 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=1.542
r580 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.4
r581 1 139 25.4929 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=0.495 $Y=1.32
+ $X2=0.495 $Y2=1.542
r582 1 3 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=0.495 $Y=1.32
+ $X2=0.495 $Y2=0.61
.ends

.subckt PM_SKY130_FD_SC_LS__CLKINV_16%VPWR 1 2 3 4 5 6 7 8 9 10 11 12 13 40 42
+ 48 54 60 66 72 78 84 90 94 98 104 110 114 116 121 122 124 125 127 128 130 131
+ 133 134 136 137 139 140 141 142 143 170 175 180 189 192 195 199
r233 198 199 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r234 195 196 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r235 192 193 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r236 189 190 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r237 186 187 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r238 184 199 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=11.28 $Y2=3.33
r239 184 196 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=10.32 $Y2=3.33
r240 183 184 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r241 181 195 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.505 $Y=3.33
+ $X2=10.34 $Y2=3.33
r242 181 183 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=10.505 $Y=3.33
+ $X2=10.8 $Y2=3.33
r243 180 198 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=11.075 $Y=3.33
+ $X2=11.297 $Y2=3.33
r244 180 183 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=11.075 $Y=3.33
+ $X2=10.8 $Y2=3.33
r245 179 196 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=10.32 $Y2=3.33
r246 179 193 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=9.36 $Y2=3.33
r247 178 179 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r248 176 192 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.605 $Y=3.33
+ $X2=9.44 $Y2=3.33
r249 176 178 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=9.605 $Y=3.33
+ $X2=9.84 $Y2=3.33
r250 175 195 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.175 $Y=3.33
+ $X2=10.34 $Y2=3.33
r251 175 178 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=10.175 $Y=3.33
+ $X2=9.84 $Y2=3.33
r252 174 193 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=9.36 $Y2=3.33
r253 174 190 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=8.4 $Y2=3.33
r254 173 174 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r255 171 189 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.625 $Y=3.33
+ $X2=8.5 $Y2=3.33
r256 171 173 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=8.625 $Y=3.33
+ $X2=8.88 $Y2=3.33
r257 170 192 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.275 $Y=3.33
+ $X2=9.44 $Y2=3.33
r258 170 173 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=9.275 $Y=3.33
+ $X2=8.88 $Y2=3.33
r259 169 190 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=8.4 $Y2=3.33
r260 168 169 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r261 166 169 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=7.44 $Y2=3.33
r262 165 166 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r263 162 163 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r264 160 163 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r265 159 160 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r266 157 160 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r267 156 157 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r268 154 157 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r269 153 154 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r270 151 154 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r271 150 151 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r272 148 151 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r273 148 187 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r274 147 148 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r275 145 186 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.222 $Y2=3.33
r276 145 147 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.72 $Y2=3.33
r277 143 166 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=5.76 $Y=3.33
+ $X2=6.48 $Y2=3.33
r278 143 163 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=5.76 $Y=3.33
+ $X2=5.52 $Y2=3.33
r279 141 168 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=7.475 $Y=3.33
+ $X2=7.44 $Y2=3.33
r280 141 142 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.475 $Y=3.33
+ $X2=7.64 $Y2=3.33
r281 139 165 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=6.51 $Y=3.33
+ $X2=6.48 $Y2=3.33
r282 139 140 7.75133 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=6.51 $Y=3.33
+ $X2=6.652 $Y2=3.33
r283 138 168 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=6.795 $Y=3.33
+ $X2=7.44 $Y2=3.33
r284 138 140 7.75133 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=6.795 $Y=3.33
+ $X2=6.652 $Y2=3.33
r285 136 162 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=5.595 $Y=3.33
+ $X2=5.52 $Y2=3.33
r286 136 137 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.595 $Y=3.33
+ $X2=5.72 $Y2=3.33
r287 135 165 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=5.845 $Y=3.33
+ $X2=6.48 $Y2=3.33
r288 135 137 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.845 $Y=3.33
+ $X2=5.72 $Y2=3.33
r289 133 159 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=4.695 $Y=3.33
+ $X2=4.56 $Y2=3.33
r290 133 134 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.695 $Y=3.33
+ $X2=4.78 $Y2=3.33
r291 132 162 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=4.865 $Y=3.33
+ $X2=5.52 $Y2=3.33
r292 132 134 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.865 $Y=3.33
+ $X2=4.78 $Y2=3.33
r293 130 156 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=3.795 $Y=3.33
+ $X2=3.6 $Y2=3.33
r294 130 131 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.795 $Y=3.33
+ $X2=3.88 $Y2=3.33
r295 129 159 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=3.965 $Y=3.33
+ $X2=4.56 $Y2=3.33
r296 129 131 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.965 $Y=3.33
+ $X2=3.88 $Y2=3.33
r297 127 153 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.895 $Y=3.33
+ $X2=2.64 $Y2=3.33
r298 127 128 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.895 $Y=3.33
+ $X2=2.98 $Y2=3.33
r299 126 156 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=3.065 $Y=3.33
+ $X2=3.6 $Y2=3.33
r300 126 128 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.065 $Y=3.33
+ $X2=2.98 $Y2=3.33
r301 124 150 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.995 $Y=3.33
+ $X2=1.68 $Y2=3.33
r302 124 125 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.995 $Y=3.33
+ $X2=2.08 $Y2=3.33
r303 123 153 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=2.165 $Y=3.33
+ $X2=2.64 $Y2=3.33
r304 123 125 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.165 $Y=3.33
+ $X2=2.08 $Y2=3.33
r305 121 147 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.015 $Y=3.33
+ $X2=0.72 $Y2=3.33
r306 121 122 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.015 $Y=3.33
+ $X2=1.14 $Y2=3.33
r307 120 150 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=1.265 $Y=3.33
+ $X2=1.68 $Y2=3.33
r308 120 122 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.265 $Y=3.33
+ $X2=1.14 $Y2=3.33
r309 116 119 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=11.24 $Y=1.985
+ $X2=11.24 $Y2=2.815
r310 114 198 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=11.24 $Y=3.245
+ $X2=11.297 $Y2=3.33
r311 114 119 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=11.24 $Y=3.245
+ $X2=11.24 $Y2=2.815
r312 110 113 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=10.34 $Y=1.985
+ $X2=10.34 $Y2=2.815
r313 108 195 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.34 $Y=3.245
+ $X2=10.34 $Y2=3.33
r314 108 113 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=10.34 $Y=3.245
+ $X2=10.34 $Y2=2.815
r315 104 107 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=9.44 $Y=1.985
+ $X2=9.44 $Y2=2.815
r316 102 192 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.44 $Y=3.245
+ $X2=9.44 $Y2=3.33
r317 102 107 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=9.44 $Y=3.245
+ $X2=9.44 $Y2=2.815
r318 98 101 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=8.5 $Y=1.985
+ $X2=8.5 $Y2=2.815
r319 96 189 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.5 $Y=3.245
+ $X2=8.5 $Y2=3.33
r320 96 101 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=8.5 $Y=3.245
+ $X2=8.5 $Y2=2.815
r321 95 142 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.805 $Y=3.33
+ $X2=7.64 $Y2=3.33
r322 94 189 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.375 $Y=3.33
+ $X2=8.5 $Y2=3.33
r323 94 95 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=8.375 $Y=3.33
+ $X2=7.805 $Y2=3.33
r324 90 93 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=7.64 $Y=1.985
+ $X2=7.64 $Y2=2.815
r325 88 142 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.64 $Y=3.245
+ $X2=7.64 $Y2=3.33
r326 88 93 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=7.64 $Y=3.245
+ $X2=7.64 $Y2=2.815
r327 84 87 33.5624 $w=2.83e-07 $l=8.3e-07 $layer=LI1_cond $X=6.652 $Y=1.985
+ $X2=6.652 $Y2=2.815
r328 82 140 0.432977 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=6.652 $Y=3.245
+ $X2=6.652 $Y2=3.33
r329 82 87 17.3877 $w=2.83e-07 $l=4.3e-07 $layer=LI1_cond $X=6.652 $Y=3.245
+ $X2=6.652 $Y2=2.815
r330 78 81 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=5.72 $Y=1.985
+ $X2=5.72 $Y2=2.815
r331 76 137 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.72 $Y=3.245
+ $X2=5.72 $Y2=3.33
r332 76 81 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=5.72 $Y=3.245
+ $X2=5.72 $Y2=2.815
r333 72 75 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=4.78 $Y=1.985
+ $X2=4.78 $Y2=2.815
r334 70 134 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.78 $Y=3.245
+ $X2=4.78 $Y2=3.33
r335 70 75 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=4.78 $Y=3.245
+ $X2=4.78 $Y2=2.815
r336 66 69 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=3.88 $Y=1.985
+ $X2=3.88 $Y2=2.815
r337 64 131 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.88 $Y=3.245
+ $X2=3.88 $Y2=3.33
r338 64 69 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=3.88 $Y=3.245
+ $X2=3.88 $Y2=2.815
r339 60 63 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=2.98 $Y=1.985
+ $X2=2.98 $Y2=2.815
r340 58 128 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.98 $Y=3.245
+ $X2=2.98 $Y2=3.33
r341 58 63 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=2.98 $Y=3.245
+ $X2=2.98 $Y2=2.815
r342 54 57 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=2.08 $Y=1.985
+ $X2=2.08 $Y2=2.815
r343 52 125 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.08 $Y=3.245
+ $X2=2.08 $Y2=3.33
r344 52 57 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=2.08 $Y=3.245
+ $X2=2.08 $Y2=2.815
r345 48 51 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=1.14 $Y=1.985
+ $X2=1.14 $Y2=2.815
r346 46 122 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=3.245
+ $X2=1.14 $Y2=3.33
r347 46 51 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=1.14 $Y=3.245
+ $X2=1.14 $Y2=2.815
r348 42 45 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=0.28 $Y=1.985
+ $X2=0.28 $Y2=2.815
r349 40 186 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.222 $Y2=3.33
r350 40 45 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.28 $Y2=2.815
r351 13 119 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=11.09
+ $Y=1.84 $X2=11.24 $Y2=2.815
r352 13 116 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=11.09
+ $Y=1.84 $X2=11.24 $Y2=1.985
r353 12 113 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=10.19
+ $Y=1.84 $X2=10.34 $Y2=2.815
r354 12 110 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=10.19
+ $Y=1.84 $X2=10.34 $Y2=1.985
r355 11 107 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=9.29
+ $Y=1.84 $X2=9.44 $Y2=2.815
r356 11 104 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=9.29
+ $Y=1.84 $X2=9.44 $Y2=1.985
r357 10 101 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=8.39
+ $Y=1.84 $X2=8.54 $Y2=2.815
r358 10 98 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=8.39
+ $Y=1.84 $X2=8.54 $Y2=1.985
r359 9 93 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=7.49
+ $Y=1.84 $X2=7.64 $Y2=2.815
r360 9 90 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=7.49
+ $Y=1.84 $X2=7.64 $Y2=1.985
r361 8 87 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=6.48
+ $Y=1.84 $X2=6.63 $Y2=2.815
r362 8 84 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=6.48
+ $Y=1.84 $X2=6.63 $Y2=1.985
r363 7 81 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=5.53
+ $Y=1.84 $X2=5.68 $Y2=2.815
r364 7 78 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=5.53
+ $Y=1.84 $X2=5.68 $Y2=1.985
r365 6 75 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=4.63
+ $Y=1.84 $X2=4.78 $Y2=2.815
r366 6 72 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=4.63
+ $Y=1.84 $X2=4.78 $Y2=1.985
r367 5 69 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=3.73
+ $Y=1.84 $X2=3.88 $Y2=2.815
r368 5 66 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=3.73
+ $Y=1.84 $X2=3.88 $Y2=1.985
r369 4 63 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.83
+ $Y=1.84 $X2=2.98 $Y2=2.815
r370 4 60 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.83
+ $Y=1.84 $X2=2.98 $Y2=1.985
r371 3 57 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.93
+ $Y=1.84 $X2=2.08 $Y2=2.815
r372 3 54 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.93
+ $Y=1.84 $X2=2.08 $Y2=1.985
r373 2 51 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.03
+ $Y=1.84 $X2=1.18 $Y2=2.815
r374 2 48 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.03
+ $Y=1.84 $X2=1.18 $Y2=1.985
r375 1 45 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r376 1 42 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_LS__CLKINV_16%Y 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16
+ 17 18 19 20 63 71 77 81 85 86 89 94 95 97 101 106 111 114 115 120 123 124 125
+ 128 135 142 149 155 162 172 180 188 196 199 204 205 209 210
c325 210 0 1.6166e-19 $X=2.53 $Y=1.885
c326 86 0 1.88851e-19 $X=6.217 $Y=1.638
r327 209 212 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.035
+ $X2=2.53 $Y2=2.035
r328 209 210 3.61044 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=2.53 $Y=1.985
+ $X2=2.53 $Y2=1.885
r329 207 212 0.577444 $w=2.3e-07 $l=9e-07 $layer=MET1_cond $X=1.63 $Y=2.035
+ $X2=2.53 $Y2=2.035
r330 204 207 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.63 $Y=2.035
+ $X2=1.63 $Y2=2.035
r331 204 205 4.56265 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=1.63 $Y=1.985
+ $X2=1.63 $Y2=1.885
r332 196 201 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=10.79 $Y=1.985
+ $X2=10.79 $Y2=2.815
r333 196 199 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.79 $Y=2.035
+ $X2=10.79 $Y2=2.035
r334 191 199 0.577444 $w=2.3e-07 $l=9e-07 $layer=MET1_cond $X=9.89 $Y=2.035
+ $X2=10.79 $Y2=2.035
r335 188 193 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=9.89 $Y=1.985
+ $X2=9.89 $Y2=2.815
r336 188 191 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.89 $Y=2.035
+ $X2=9.89 $Y2=2.035
r337 183 191 0.577444 $w=2.3e-07 $l=9e-07 $layer=MET1_cond $X=8.99 $Y=2.035
+ $X2=9.89 $Y2=2.035
r338 180 185 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=8.99 $Y=1.985
+ $X2=8.99 $Y2=2.815
r339 180 183 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.99 $Y=2.035
+ $X2=8.99 $Y2=2.035
r340 175 183 0.577444 $w=2.3e-07 $l=9e-07 $layer=MET1_cond $X=8.09 $Y=2.035
+ $X2=8.99 $Y2=2.035
r341 172 177 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=8.09 $Y=1.985
+ $X2=8.09 $Y2=2.815
r342 172 175 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.09 $Y=2.035
+ $X2=8.09 $Y2=2.035
r343 167 175 0.596692 $w=2.3e-07 $l=9.3e-07 $layer=MET1_cond $X=7.16 $Y=2.035
+ $X2=8.09 $Y2=2.035
r344 165 169 39.0419 $w=2.43e-07 $l=8.3e-07 $layer=LI1_cond $X=7.167 $Y=1.985
+ $X2=7.167 $Y2=2.815
r345 165 167 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.16 $Y=2.035
+ $X2=7.16 $Y2=2.035
r346 162 165 64.6779 $w=2.43e-07 $l=1.375e-06 $layer=LI1_cond $X=7.167 $Y=0.61
+ $X2=7.167 $Y2=1.985
r347 157 167 0.628772 $w=2.3e-07 $l=9.8e-07 $layer=MET1_cond $X=6.18 $Y=2.035
+ $X2=7.16 $Y2=2.035
r348 155 159 30.366 $w=3.13e-07 $l=8.3e-07 $layer=LI1_cond $X=6.172 $Y=1.985
+ $X2=6.172 $Y2=2.815
r349 155 157 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.18 $Y=2.035
+ $X2=6.18 $Y2=2.035
r350 149 152 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=5.23 $Y=2.035
+ $X2=5.23 $Y2=2.815
r351 149 150 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.23 $Y=2.035
+ $X2=5.23 $Y2=2.035
r352 144 150 0.577444 $w=2.3e-07 $l=9e-07 $layer=MET1_cond $X=4.33 $Y=2.035
+ $X2=5.23 $Y2=2.035
r353 142 146 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=4.33 $Y=1.985
+ $X2=4.33 $Y2=2.815
r354 142 144 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.33 $Y=2.035
+ $X2=4.33 $Y2=2.035
r355 137 144 0.558196 $w=2.3e-07 $l=8.7e-07 $layer=MET1_cond $X=3.46 $Y=2.035
+ $X2=4.33 $Y2=2.035
r356 137 212 0.596692 $w=2.3e-07 $l=9.3e-07 $layer=MET1_cond $X=3.46 $Y=2.035
+ $X2=2.53 $Y2=2.035
r357 135 139 36.7895 $w=2.58e-07 $l=8.3e-07 $layer=LI1_cond $X=3.465 $Y=1.985
+ $X2=3.465 $Y2=2.815
r358 135 137 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.46 $Y=2.035
+ $X2=3.46 $Y2=2.035
r359 130 207 0.58386 $w=2.3e-07 $l=9.1e-07 $layer=MET1_cond $X=0.72 $Y=2.035
+ $X2=1.63 $Y2=2.035
r360 128 132 48.4498 $w=1.88e-07 $l=8.3e-07 $layer=LI1_cond $X=0.72 $Y=1.985
+ $X2=0.72 $Y2=2.815
r361 128 130 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=2.035
+ $X2=0.72 $Y2=2.035
r362 125 157 0.272682 $w=2.3e-07 $l=4.25e-07 $layer=MET1_cond $X=5.755 $Y=2.035
+ $X2=6.18 $Y2=2.035
r363 125 150 0.336842 $w=2.3e-07 $l=5.25e-07 $layer=MET1_cond $X=5.755 $Y=2.035
+ $X2=5.23 $Y2=2.035
r364 123 124 13.8636 $w=1.78e-07 $l=2.25e-07 $layer=LI1_cond $X=6.25 $Y=1.01
+ $X2=6.25 $Y2=0.785
r365 122 155 0.292684 $w=3.13e-07 $l=8e-09 $layer=LI1_cond $X=6.172 $Y=1.977
+ $X2=6.172 $Y2=1.985
r366 117 120 2.62582 $w=3.93e-07 $l=9e-08 $layer=LI1_cond $X=5.34 $Y=0.577
+ $X2=5.43 $Y2=0.577
r367 116 149 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=5.23 $Y=2.01
+ $X2=5.23 $Y2=2.035
r368 114 116 0.901327 $w=3.58e-07 $l=2.5e-08 $layer=LI1_cond $X=5.245 $Y=1.985
+ $X2=5.245 $Y2=2.01
r369 114 115 7.55066 $w=3.58e-07 $l=1.35e-07 $layer=LI1_cond $X=5.245 $Y=1.985
+ $X2=5.245 $Y2=1.85
r370 111 142 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=4.33 $Y=1.9
+ $X2=4.33 $Y2=1.985
r371 110 111 2.2967 $w=3.28e-07 $l=5e-08 $layer=LI1_cond $X=4.345 $Y=1.85
+ $X2=4.345 $Y2=1.9
r372 108 135 53.6329 $w=2.58e-07 $l=1.21e-06 $layer=LI1_cond $X=3.465 $Y=0.775
+ $X2=3.465 $Y2=1.985
r373 106 108 6.63702 $w=2.93e-07 $l=1.65e-07 $layer=LI1_cond $X=3.447 $Y=0.61
+ $X2=3.447 $Y2=0.775
r374 103 210 42.6404 $w=2.98e-07 $l=1.11e-06 $layer=LI1_cond $X=2.515 $Y=0.775
+ $X2=2.515 $Y2=1.885
r375 101 103 6.07341 $w=3.13e-07 $l=1.65e-07 $layer=LI1_cond $X=2.507 $Y=0.61
+ $X2=2.507 $Y2=0.775
r376 99 205 55.6179 $w=2.28e-07 $l=1.11e-06 $layer=LI1_cond $X=1.58 $Y=0.775
+ $X2=1.58 $Y2=1.885
r377 97 99 7.49534 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=1.57 $Y=0.61
+ $X2=1.57 $Y2=0.775
r378 94 128 4.08612 $w=1.88e-07 $l=7e-08 $layer=LI1_cond $X=0.72 $Y=1.915
+ $X2=0.72 $Y2=1.985
r379 94 95 5.58789 $w=1.88e-07 $l=9.5e-08 $layer=LI1_cond $X=0.72 $Y=1.915
+ $X2=0.72 $Y2=1.82
r380 93 95 64.3889 $w=1.78e-07 $l=1.045e-06 $layer=LI1_cond $X=0.715 $Y=0.775
+ $X2=0.715 $Y2=1.82
r381 87 124 6.23075 $w=2.23e-07 $l=1.12e-07 $layer=LI1_cond $X=6.272 $Y=0.673
+ $X2=6.272 $Y2=0.785
r382 87 89 3.22684 $w=2.23e-07 $l=6.3e-08 $layer=LI1_cond $X=6.272 $Y=0.673
+ $X2=6.272 $Y2=0.61
r383 86 122 15.0393 $w=2.75e-07 $l=3.60799e-07 $layer=LI1_cond $X=6.217 $Y=1.638
+ $X2=6.172 $Y2=1.977
r384 85 123 6.57226 $w=2.43e-07 $l=1.22e-07 $layer=LI1_cond $X=6.217 $Y=1.132
+ $X2=6.217 $Y2=1.01
r385 85 86 23.8015 $w=2.43e-07 $l=5.06e-07 $layer=LI1_cond $X=6.217 $Y=1.132
+ $X2=6.217 $Y2=1.638
r386 83 117 5.70203 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=5.34 $Y=0.775
+ $X2=5.34 $Y2=0.577
r387 83 115 70.1337 $w=1.68e-07 $l=1.075e-06 $layer=LI1_cond $X=5.34 $Y=0.775
+ $X2=5.34 $Y2=1.85
r388 81 110 54.9627 $w=2.58e-07 $l=1.24e-06 $layer=LI1_cond $X=4.395 $Y=0.61
+ $X2=4.395 $Y2=1.85
r389 75 209 2.26996 $w=3.28e-07 $l=6.5e-08 $layer=LI1_cond $X=2.53 $Y=2.05
+ $X2=2.53 $Y2=1.985
r390 75 77 26.7157 $w=3.28e-07 $l=7.65e-07 $layer=LI1_cond $X=2.53 $Y=2.05
+ $X2=2.53 $Y2=2.815
r391 69 204 2.26996 $w=3.28e-07 $l=6.5e-08 $layer=LI1_cond $X=1.63 $Y=2.05
+ $X2=1.63 $Y2=1.985
r392 69 71 26.7157 $w=3.28e-07 $l=7.65e-07 $layer=LI1_cond $X=1.63 $Y=2.05
+ $X2=1.63 $Y2=2.815
r393 61 93 5.58789 $w=1.88e-07 $l=9.5e-08 $layer=LI1_cond $X=0.71 $Y=0.68
+ $X2=0.71 $Y2=0.775
r394 61 63 4.08612 $w=1.88e-07 $l=7e-08 $layer=LI1_cond $X=0.71 $Y=0.68 $X2=0.71
+ $Y2=0.61
r395 20 201 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=10.64
+ $Y=1.84 $X2=10.79 $Y2=2.815
r396 20 196 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=10.64
+ $Y=1.84 $X2=10.79 $Y2=1.985
r397 19 193 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=9.74
+ $Y=1.84 $X2=9.89 $Y2=2.815
r398 19 188 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=9.74
+ $Y=1.84 $X2=9.89 $Y2=1.985
r399 18 185 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=8.84
+ $Y=1.84 $X2=8.99 $Y2=2.815
r400 18 180 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=8.84
+ $Y=1.84 $X2=8.99 $Y2=1.985
r401 17 177 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=7.94
+ $Y=1.84 $X2=8.09 $Y2=2.815
r402 17 172 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=7.94
+ $Y=1.84 $X2=8.09 $Y2=1.985
r403 16 169 400 $w=1.7e-07 $l=1.06119e-06 $layer=licon1_PDIFF $count=1 $X=6.98
+ $Y=1.84 $X2=7.16 $Y2=2.815
r404 16 165 400 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_PDIFF $count=1 $X=6.98
+ $Y=1.84 $X2=7.16 $Y2=1.985
r405 15 159 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=6.03
+ $Y=1.84 $X2=6.18 $Y2=2.815
r406 15 155 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=6.03
+ $Y=1.84 $X2=6.18 $Y2=1.985
r407 14 152 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=5.08
+ $Y=1.84 $X2=5.23 $Y2=2.815
r408 14 114 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=5.08
+ $Y=1.84 $X2=5.23 $Y2=1.985
r409 13 146 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=4.18
+ $Y=1.84 $X2=4.33 $Y2=2.815
r410 13 142 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=4.18
+ $Y=1.84 $X2=4.33 $Y2=1.985
r411 12 139 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=3.28
+ $Y=1.84 $X2=3.43 $Y2=2.815
r412 12 135 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=3.28
+ $Y=1.84 $X2=3.43 $Y2=1.985
r413 11 209 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.38
+ $Y=1.84 $X2=2.53 $Y2=1.985
r414 11 77 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.38
+ $Y=1.84 $X2=2.53 $Y2=2.815
r415 10 204 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.48
+ $Y=1.84 $X2=1.63 $Y2=1.985
r416 10 71 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.48
+ $Y=1.84 $X2=1.63 $Y2=2.815
r417 9 132 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.84 $X2=0.73 $Y2=2.815
r418 9 128 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.84 $X2=0.73 $Y2=1.985
r419 8 162 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=7.01
+ $Y=0.4 $X2=7.15 $Y2=0.61
r420 7 89 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=6.15
+ $Y=0.4 $X2=6.29 $Y2=0.61
r421 6 120 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=5.29
+ $Y=0.4 $X2=5.43 $Y2=0.61
r422 5 81 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.29
+ $Y=0.4 $X2=4.43 $Y2=0.61
r423 4 106 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.29
+ $Y=0.4 $X2=3.43 $Y2=0.61
r424 3 101 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.36
+ $Y=0.4 $X2=2.5 $Y2=0.61
r425 2 97 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.43
+ $Y=0.4 $X2=1.57 $Y2=0.61
r426 1 63 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.4 $X2=0.71 $Y2=0.61
.ends

.subckt PM_SKY130_FD_SC_LS__CLKINV_16%VGND 1 2 3 4 5 6 7 8 9 28 30 34 38 42 46
+ 50 54 58 61 62 64 65 67 68 70 71 73 74 76 77 79 80 82 85 86 114 122 123 130
c146 30 0 1.31047e-19 $X=0.28 $Y=0.61
r147 132 133 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r148 129 132 4.06215 $w=7.93e-07 $l=2.7e-07 $layer=LI1_cond $X=7.65 $Y=0.312
+ $X2=7.92 $Y2=0.312
r149 129 130 11.4033 $w=7.93e-07 $l=1.65e-07 $layer=LI1_cond $X=7.65 $Y=0.312
+ $X2=7.485 $Y2=0.312
r150 126 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r151 122 123 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r152 120 123 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=11.28 $Y2=0
r153 119 122 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=9.84 $Y=0
+ $X2=11.28 $Y2=0
r154 119 120 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.84 $Y=0
+ $X2=9.84 $Y2=0
r155 117 120 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=9.84 $Y2=0
r156 117 133 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=7.92 $Y2=0
r157 116 117 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r158 114 132 5.4162 $w=7.93e-07 $l=3.6e-07 $layer=LI1_cond $X=8.28 $Y=0.312
+ $X2=7.92 $Y2=0.312
r159 114 116 16.2486 $w=7.93e-07 $l=1.08e-06 $layer=LI1_cond $X=8.28 $Y=0.312
+ $X2=9.36 $Y2=0.312
r160 113 133 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=7.92 $Y2=0
r161 112 130 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=7.44 $Y=0
+ $X2=7.485 $Y2=0
r162 112 113 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r163 109 113 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=0
+ $X2=7.44 $Y2=0
r164 108 109 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r165 105 106 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r166 103 106 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=0
+ $X2=5.52 $Y2=0
r167 102 103 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r168 100 103 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0
+ $X2=4.56 $Y2=0
r169 99 100 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r170 97 100 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r171 96 97 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r172 94 97 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r173 93 94 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r174 91 94 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r175 91 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0
+ $X2=0.24 $Y2=0
r176 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r177 88 126 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=0
+ $X2=0.222 $Y2=0
r178 88 90 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=0
+ $X2=0.72 $Y2=0
r179 86 109 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=5.76 $Y=0
+ $X2=6.48 $Y2=0
r180 86 106 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=5.76 $Y=0
+ $X2=5.52 $Y2=0
r181 85 119 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=9.825 $Y=0
+ $X2=9.84 $Y2=0
r182 84 85 11.4033 $w=7.93e-07 $l=1.65e-07 $layer=LI1_cond $X=9.66 $Y=0.312
+ $X2=9.825 $Y2=0.312
r183 82 116 1.02306 $w=7.93e-07 $l=6.8e-08 $layer=LI1_cond $X=9.428 $Y=0.312
+ $X2=9.36 $Y2=0.312
r184 82 84 3.49044 $w=7.93e-07 $l=2.32e-07 $layer=LI1_cond $X=9.428 $Y=0.312
+ $X2=9.66 $Y2=0.312
r185 79 108 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=6.555 $Y=0
+ $X2=6.48 $Y2=0
r186 79 80 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=6.555 $Y=0 $X2=6.715
+ $Y2=0
r187 78 112 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=6.875 $Y=0
+ $X2=7.44 $Y2=0
r188 78 80 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=6.875 $Y=0 $X2=6.715
+ $Y2=0
r189 76 105 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=5.695 $Y=0
+ $X2=5.52 $Y2=0
r190 76 77 7.75133 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=5.695 $Y=0
+ $X2=5.837 $Y2=0
r191 75 108 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=5.98 $Y=0 $X2=6.48
+ $Y2=0
r192 75 77 7.75133 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=5.98 $Y=0 $X2=5.837
+ $Y2=0
r193 73 102 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=4.765 $Y=0
+ $X2=4.56 $Y2=0
r194 73 74 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=4.765 $Y=0 $X2=4.925
+ $Y2=0
r195 72 105 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=5.085 $Y=0
+ $X2=5.52 $Y2=0
r196 72 74 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=5.085 $Y=0 $X2=4.925
+ $Y2=0
r197 70 99 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.765 $Y=0 $X2=3.6
+ $Y2=0
r198 70 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.765 $Y=0 $X2=3.93
+ $Y2=0
r199 69 102 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=4.095 $Y=0
+ $X2=4.56 $Y2=0
r200 69 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.095 $Y=0 $X2=3.93
+ $Y2=0
r201 67 96 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=2.845 $Y=0
+ $X2=2.64 $Y2=0
r202 67 68 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.845 $Y=0 $X2=2.97
+ $Y2=0
r203 66 99 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=3.095 $Y=0 $X2=3.6
+ $Y2=0
r204 66 68 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.095 $Y=0 $X2=2.97
+ $Y2=0
r205 64 93 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.885 $Y=0
+ $X2=1.68 $Y2=0
r206 64 65 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=1.885 $Y=0 $X2=2.025
+ $Y2=0
r207 63 96 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=2.165 $Y=0
+ $X2=2.64 $Y2=0
r208 63 65 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.165 $Y=0 $X2=2.025
+ $Y2=0
r209 61 90 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.975 $Y=0
+ $X2=0.72 $Y2=0
r210 61 62 7.75133 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=0.975 $Y=0
+ $X2=1.117 $Y2=0
r211 60 93 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=1.26 $Y=0 $X2=1.68
+ $Y2=0
r212 60 62 7.75133 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=1.26 $Y=0 $X2=1.117
+ $Y2=0
r213 56 80 0.800721 $w=3.2e-07 $l=8.5e-08 $layer=LI1_cond $X=6.715 $Y=0.085
+ $X2=6.715 $Y2=0
r214 56 58 18.9073 $w=3.18e-07 $l=5.25e-07 $layer=LI1_cond $X=6.715 $Y=0.085
+ $X2=6.715 $Y2=0.61
r215 52 77 0.432977 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=5.837 $Y=0.085
+ $X2=5.837 $Y2=0
r216 52 54 21.2292 $w=2.83e-07 $l=5.25e-07 $layer=LI1_cond $X=5.837 $Y=0.085
+ $X2=5.837 $Y2=0.61
r217 48 74 0.800721 $w=3.2e-07 $l=8.5e-08 $layer=LI1_cond $X=4.925 $Y=0.085
+ $X2=4.925 $Y2=0
r218 48 50 18.9073 $w=3.18e-07 $l=5.25e-07 $layer=LI1_cond $X=4.925 $Y=0.085
+ $X2=4.925 $Y2=0.61
r219 44 71 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.93 $Y=0.085
+ $X2=3.93 $Y2=0
r220 44 46 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=3.93 $Y=0.085
+ $X2=3.93 $Y2=0.61
r221 40 68 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.97 $Y=0.085
+ $X2=2.97 $Y2=0
r222 40 42 24.2013 $w=2.48e-07 $l=5.25e-07 $layer=LI1_cond $X=2.97 $Y=0.085
+ $X2=2.97 $Y2=0.61
r223 36 65 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.025 $Y=0.085
+ $X2=2.025 $Y2=0
r224 36 38 21.6083 $w=2.78e-07 $l=5.25e-07 $layer=LI1_cond $X=2.025 $Y=0.085
+ $X2=2.025 $Y2=0.61
r225 32 62 0.432977 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=1.117 $Y=0.085
+ $X2=1.117 $Y2=0
r226 32 34 21.2292 $w=2.83e-07 $l=5.25e-07 $layer=LI1_cond $X=1.117 $Y=0.085
+ $X2=1.117 $Y2=0.61
r227 28 126 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.222 $Y2=0
r228 28 30 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.28 $Y2=0.61
r229 9 129 60.6667 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=3
+ $X=7.44 $Y=0.4 $X2=7.65 $Y2=0.545
r230 9 84 60.6667 $w=1.7e-07 $l=2.29135e-06 $layer=licon1_NDIFF $count=3 $X=7.44
+ $Y=0.4 $X2=9.66 $Y2=0.545
r231 8 58 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=6.58
+ $Y=0.4 $X2=6.72 $Y2=0.61
r232 7 54 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=5.72
+ $Y=0.4 $X2=5.86 $Y2=0.61
r233 6 50 182 $w=1.7e-07 $l=2.96985e-07 $layer=licon1_NDIFF $count=1 $X=4.72
+ $Y=0.4 $X2=4.93 $Y2=0.61
r234 5 46 182 $w=1.7e-07 $l=2.96985e-07 $layer=licon1_NDIFF $count=1 $X=3.72
+ $Y=0.4 $X2=3.93 $Y2=0.61
r235 4 42 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.79
+ $Y=0.4 $X2=2.93 $Y2=0.61
r236 3 38 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.86
+ $Y=0.4 $X2=2 $Y2=0.61
r237 2 34 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1 $Y=0.4
+ $X2=1.14 $Y2=0.61
r238 1 30 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.4 $X2=0.28 $Y2=0.61
.ends

