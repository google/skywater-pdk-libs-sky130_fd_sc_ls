* File: sky130_fd_sc_ls__nor2b_4.pxi.spice
* Created: Fri Aug 28 13:38:00 2020
* 
x_PM_SKY130_FD_SC_LS__NOR2B_4%A N_A_c_80_n N_A_c_91_n N_A_M1006_g N_A_c_81_n
+ N_A_c_93_n N_A_M1007_g N_A_c_82_n N_A_c_95_n N_A_M1011_g N_A_c_83_n
+ N_A_M1000_g N_A_c_96_n N_A_M1012_g N_A_c_84_n N_A_M1004_g N_A_c_85_n
+ N_A_c_86_n N_A_c_87_n N_A_c_88_n A A N_A_c_89_n PM_SKY130_FD_SC_LS__NOR2B_4%A
x_PM_SKY130_FD_SC_LS__NOR2B_4%A_353_323# N_A_353_323#_M1014_d
+ N_A_353_323#_M1010_d N_A_353_323#_c_197_n N_A_353_323#_M1001_g
+ N_A_353_323#_c_192_n N_A_353_323#_M1003_g N_A_353_323#_c_198_n
+ N_A_353_323#_M1002_g N_A_353_323#_c_193_n N_A_353_323#_M1008_g
+ N_A_353_323#_c_199_n N_A_353_323#_M1005_g N_A_353_323#_c_200_n
+ N_A_353_323#_M1009_g N_A_353_323#_c_201_n N_A_353_323#_c_202_n
+ N_A_353_323#_c_203_n N_A_353_323#_c_194_n N_A_353_323#_c_195_n
+ N_A_353_323#_c_196_n PM_SKY130_FD_SC_LS__NOR2B_4%A_353_323#
x_PM_SKY130_FD_SC_LS__NOR2B_4%B_N N_B_N_c_300_n N_B_N_M1010_g N_B_N_M1014_g
+ N_B_N_c_301_n N_B_N_M1013_g B_N B_N N_B_N_c_299_n
+ PM_SKY130_FD_SC_LS__NOR2B_4%B_N
x_PM_SKY130_FD_SC_LS__NOR2B_4%VPWR N_VPWR_M1006_s N_VPWR_M1007_s N_VPWR_M1012_s
+ N_VPWR_M1013_s N_VPWR_c_333_n N_VPWR_c_334_n N_VPWR_c_335_n N_VPWR_c_336_n
+ N_VPWR_c_337_n N_VPWR_c_338_n N_VPWR_c_339_n N_VPWR_c_340_n VPWR
+ N_VPWR_c_341_n N_VPWR_c_342_n N_VPWR_c_343_n N_VPWR_c_332_n
+ PM_SKY130_FD_SC_LS__NOR2B_4%VPWR
x_PM_SKY130_FD_SC_LS__NOR2B_4%A_116_368# N_A_116_368#_M1006_d
+ N_A_116_368#_M1011_d N_A_116_368#_M1002_s N_A_116_368#_M1009_s
+ N_A_116_368#_c_404_n N_A_116_368#_c_399_n N_A_116_368#_c_409_n
+ N_A_116_368#_c_411_n N_A_116_368#_c_412_n N_A_116_368#_c_400_n
+ N_A_116_368#_c_401_n N_A_116_368#_c_420_n N_A_116_368#_c_402_n
+ N_A_116_368#_c_416_n N_A_116_368#_c_403_n
+ PM_SKY130_FD_SC_LS__NOR2B_4%A_116_368#
x_PM_SKY130_FD_SC_LS__NOR2B_4%Y N_Y_M1003_d N_Y_M1000_d N_Y_M1001_d N_Y_M1005_d
+ N_Y_c_463_n N_Y_c_464_n N_Y_c_465_n N_Y_c_510_n N_Y_c_512_n N_Y_c_487_n
+ N_Y_c_517_n N_Y_c_520_n N_Y_c_466_n N_Y_c_467_n N_Y_c_468_n N_Y_c_523_n
+ N_Y_c_497_n Y Y Y PM_SKY130_FD_SC_LS__NOR2B_4%Y
x_PM_SKY130_FD_SC_LS__NOR2B_4%VGND N_VGND_M1003_s N_VGND_M1008_s N_VGND_M1004_s
+ N_VGND_c_559_n N_VGND_c_560_n VGND N_VGND_c_561_n N_VGND_c_562_n
+ N_VGND_c_563_n N_VGND_c_564_n N_VGND_c_565_n N_VGND_c_566_n N_VGND_c_567_n
+ N_VGND_c_568_n PM_SKY130_FD_SC_LS__NOR2B_4%VGND
cc_1 VNB N_A_c_80_n 0.0188384f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.675
cc_2 VNB N_A_c_81_n 0.0162349f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.675
cc_3 VNB N_A_c_82_n 0.0176514f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=1.675
cc_4 VNB N_A_c_83_n 0.0193643f $X=-0.19 $Y=-0.245 $X2=3.51 $Y2=1.22
cc_5 VNB N_A_c_84_n 0.016198f $X=-0.19 $Y=-0.245 $X2=3.94 $Y2=1.22
cc_6 VNB N_A_c_85_n 0.0136474f $X=-0.19 $Y=-0.245 $X2=3.645 $Y2=1.095
cc_7 VNB N_A_c_86_n 0.0161986f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=1.095
cc_8 VNB N_A_c_87_n 0.00205904f $X=-0.19 $Y=-0.245 $X2=3.81 $Y2=1.385
cc_9 VNB N_A_c_88_n 0.0521604f $X=-0.19 $Y=-0.245 $X2=3.81 $Y2=1.385
cc_10 VNB N_A_c_89_n 0.0863763f $X=-0.19 $Y=-0.245 $X2=1.295 $Y2=1.175
cc_11 VNB N_A_353_323#_c_192_n 0.0180618f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_12 VNB N_A_353_323#_c_193_n 0.0197816f $X=-0.19 $Y=-0.245 $X2=3.51 $Y2=1.22
cc_13 VNB N_A_353_323#_c_194_n 0.00529851f $X=-0.19 $Y=-0.245 $X2=0.955
+ $Y2=1.175
cc_14 VNB N_A_353_323#_c_195_n 0.107335f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=1.175
cc_15 VNB N_A_353_323#_c_196_n 0.0346171f $X=-0.19 $Y=-0.245 $X2=1.295 $Y2=1.21
cc_16 VNB N_B_N_M1014_g 0.0395613f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.34
cc_17 VNB B_N 0.0261981f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=1.34
cc_18 VNB N_B_N_c_299_n 0.0404365f $X=-0.19 $Y=-0.245 $X2=3.51 $Y2=0.74
cc_19 VNB N_VPWR_c_332_n 0.223389f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_Y_c_463_n 0.0115493f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=2.4
cc_21 VNB N_Y_c_464_n 0.00816012f $X=-0.19 $Y=-0.245 $X2=3.51 $Y2=0.74
cc_22 VNB N_Y_c_465_n 6.68229e-19 $X=-0.19 $Y=-0.245 $X2=3.705 $Y2=1.765
cc_23 VNB N_Y_c_466_n 8.97027e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_Y_c_467_n 0.00230198f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.21
cc_25 VNB N_Y_c_468_n 0.032652f $X=-0.19 $Y=-0.245 $X2=1.295 $Y2=1.175
cc_26 VNB Y 0.0283086f $X=-0.19 $Y=-0.245 $X2=1.295 $Y2=1.21
cc_27 VNB Y 0.0173879f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=1.21
cc_28 VNB N_VGND_c_559_n 0.0166025f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=1.675
cc_29 VNB N_VGND_c_560_n 0.00489167f $X=-0.19 $Y=-0.245 $X2=3.51 $Y2=0.74
cc_30 VNB N_VGND_c_561_n 0.0455645f $X=-0.19 $Y=-0.245 $X2=3.94 $Y2=1.22
cc_31 VNB N_VGND_c_562_n 0.0170209f $X=-0.19 $Y=-0.245 $X2=3.81 $Y2=1.385
cc_32 VNB N_VGND_c_563_n 0.0292937f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.175
cc_33 VNB N_VGND_c_564_n 0.303426f $X=-0.19 $Y=-0.245 $X2=1.295 $Y2=1.175
cc_34 VNB N_VGND_c_565_n 0.00631651f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=1.175
cc_35 VNB N_VGND_c_566_n 0.0186046f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.21
cc_36 VNB N_VGND_c_567_n 0.0247843f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_568_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VPB N_A_c_80_n 8.48304e-19 $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.675
cc_39 VPB N_A_c_91_n 0.0265442f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_40 VPB N_A_c_81_n 6.2759e-19 $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.675
cc_41 VPB N_A_c_93_n 0.0205685f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.765
cc_42 VPB N_A_c_82_n 6.28632e-19 $X=-0.19 $Y=1.66 $X2=1.405 $Y2=1.675
cc_43 VPB N_A_c_95_n 0.0203294f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=1.765
cc_44 VPB N_A_c_96_n 0.0158871f $X=-0.19 $Y=1.66 $X2=3.705 $Y2=1.765
cc_45 VPB N_A_c_88_n 0.00725861f $X=-0.19 $Y=1.66 $X2=3.81 $Y2=1.385
cc_46 VPB N_A_353_323#_c_197_n 0.0145915f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.675
cc_47 VPB N_A_353_323#_c_198_n 0.0147472f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=1.765
cc_48 VPB N_A_353_323#_c_199_n 0.0147503f $X=-0.19 $Y=1.66 $X2=3.705 $Y2=1.765
cc_49 VPB N_A_353_323#_c_200_n 0.0145086f $X=-0.19 $Y=1.66 $X2=3.94 $Y2=1.22
cc_50 VPB N_A_353_323#_c_201_n 7.49862e-19 $X=-0.19 $Y=1.66 $X2=3.645 $Y2=1.095
cc_51 VPB N_A_353_323#_c_202_n 0.017297f $X=-0.19 $Y=1.66 $X2=3.81 $Y2=1.385
cc_52 VPB N_A_353_323#_c_203_n 0.00704867f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_A_353_323#_c_195_n 0.0314269f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=1.175
cc_54 VPB N_B_N_c_300_n 0.0156104f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.34
cc_55 VPB N_B_N_c_301_n 0.0166598f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.765
cc_56 VPB B_N 0.00796315f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=1.34
cc_57 VPB N_B_N_c_299_n 0.0560576f $X=-0.19 $Y=1.66 $X2=3.51 $Y2=0.74
cc_58 VPB N_VPWR_c_333_n 0.0106521f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=1.765
cc_59 VPB N_VPWR_c_334_n 0.0535877f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=2.4
cc_60 VPB N_VPWR_c_335_n 0.00769929f $X=-0.19 $Y=1.66 $X2=3.705 $Y2=2.4
cc_61 VPB N_VPWR_c_336_n 0.013214f $X=-0.19 $Y=1.66 $X2=3.645 $Y2=1.095
cc_62 VPB N_VPWR_c_337_n 0.0117686f $X=-0.19 $Y=1.66 $X2=3.81 $Y2=1.385
cc_63 VPB N_VPWR_c_338_n 0.0541997f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_339_n 0.0597959f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_340_n 0.00631788f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_341_n 0.0206041f $X=-0.19 $Y=1.66 $X2=1.295 $Y2=1.175
cc_67 VPB N_VPWR_c_342_n 0.0212408f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_343_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_332_n 0.0824955f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_A_116_368#_c_399_n 0.00257348f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=2.4
cc_71 VPB N_A_116_368#_c_400_n 0.00259172f $X=-0.19 $Y=1.66 $X2=3.94 $Y2=0.74
cc_72 VPB N_A_116_368#_c_401_n 0.00171072f $X=-0.19 $Y=1.66 $X2=3.94 $Y2=0.74
cc_73 VPB N_A_116_368#_c_402_n 0.00467121f $X=-0.19 $Y=1.66 $X2=3.81 $Y2=1.385
cc_74 VPB N_A_116_368#_c_403_n 0.00218363f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=1.175
cc_75 VPB N_Y_c_464_n 0.00767295f $X=-0.19 $Y=1.66 $X2=3.51 $Y2=0.74
cc_76 VPB N_Y_c_465_n 7.22836e-19 $X=-0.19 $Y=1.66 $X2=3.705 $Y2=1.765
cc_77 VPB N_Y_c_466_n 0.00182538f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_Y_c_467_n 0.00101457f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.21
cc_79 VPB Y 0.00244476f $X=-0.19 $Y=1.66 $X2=1.68 $Y2=1.21
cc_80 N_A_c_95_n N_A_353_323#_c_197_n 0.0106506f $X=1.405 $Y=1.765 $X2=0 $Y2=0
cc_81 N_A_c_85_n N_A_353_323#_c_192_n 0.0125877f $X=3.645 $Y=1.095 $X2=0 $Y2=0
cc_82 N_A_c_86_n N_A_353_323#_c_192_n 0.00632392f $X=1.795 $Y=1.095 $X2=0 $Y2=0
cc_83 N_A_c_89_n N_A_353_323#_c_192_n 0.00840639f $X=1.295 $Y=1.175 $X2=0 $Y2=0
cc_84 N_A_c_85_n N_A_353_323#_c_193_n 0.0125331f $X=3.645 $Y=1.095 $X2=0 $Y2=0
cc_85 N_A_c_96_n N_A_353_323#_c_200_n 0.0248856f $X=3.705 $Y=1.765 $X2=0 $Y2=0
cc_86 N_A_c_85_n N_A_353_323#_c_201_n 0.0749937f $X=3.645 $Y=1.095 $X2=0 $Y2=0
cc_87 N_A_c_86_n N_A_353_323#_c_201_n 0.00262271f $X=1.795 $Y=1.095 $X2=0 $Y2=0
cc_88 N_A_c_87_n N_A_353_323#_c_201_n 0.00688023f $X=3.81 $Y=1.385 $X2=0 $Y2=0
cc_89 N_A_c_88_n N_A_353_323#_c_201_n 0.00187212f $X=3.81 $Y=1.385 $X2=0 $Y2=0
cc_90 N_A_c_96_n N_A_353_323#_c_202_n 0.0116494f $X=3.705 $Y=1.765 $X2=0 $Y2=0
cc_91 N_A_c_85_n N_A_353_323#_c_202_n 0.0132262f $X=3.645 $Y=1.095 $X2=0 $Y2=0
cc_92 N_A_c_87_n N_A_353_323#_c_202_n 0.0251788f $X=3.81 $Y=1.385 $X2=0 $Y2=0
cc_93 N_A_c_88_n N_A_353_323#_c_202_n 0.0127292f $X=3.81 $Y=1.385 $X2=0 $Y2=0
cc_94 N_A_c_96_n N_A_353_323#_c_203_n 7.76807e-19 $X=3.705 $Y=1.765 $X2=0 $Y2=0
cc_95 N_A_c_84_n N_A_353_323#_c_194_n 0.00177623f $X=3.94 $Y=1.22 $X2=0 $Y2=0
cc_96 N_A_c_85_n N_A_353_323#_c_194_n 0.00603876f $X=3.645 $Y=1.095 $X2=0 $Y2=0
cc_97 N_A_c_87_n N_A_353_323#_c_194_n 0.0123049f $X=3.81 $Y=1.385 $X2=0 $Y2=0
cc_98 N_A_c_88_n N_A_353_323#_c_194_n 7.7613e-19 $X=3.81 $Y=1.385 $X2=0 $Y2=0
cc_99 N_A_c_82_n N_A_353_323#_c_195_n 0.0156392f $X=1.405 $Y=1.675 $X2=0 $Y2=0
cc_100 N_A_c_85_n N_A_353_323#_c_195_n 0.027508f $X=3.645 $Y=1.095 $X2=0 $Y2=0
cc_101 N_A_c_86_n N_A_353_323#_c_195_n 2.05585e-19 $X=1.795 $Y=1.095 $X2=0 $Y2=0
cc_102 N_A_c_87_n N_A_353_323#_c_195_n 0.00151745f $X=3.81 $Y=1.385 $X2=0 $Y2=0
cc_103 N_A_c_88_n N_A_353_323#_c_195_n 0.0256104f $X=3.81 $Y=1.385 $X2=0 $Y2=0
cc_104 N_A_c_84_n N_A_353_323#_c_196_n 9.69162e-19 $X=3.94 $Y=1.22 $X2=0 $Y2=0
cc_105 N_A_c_96_n N_B_N_c_300_n 0.0200987f $X=3.705 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_106 N_A_c_84_n N_B_N_M1014_g 0.0194276f $X=3.94 $Y=1.22 $X2=0 $Y2=0
cc_107 N_A_c_85_n N_B_N_M1014_g 5.68631e-19 $X=3.645 $Y=1.095 $X2=0 $Y2=0
cc_108 N_A_c_87_n N_B_N_M1014_g 0.001297f $X=3.81 $Y=1.385 $X2=0 $Y2=0
cc_109 N_A_c_96_n N_B_N_c_299_n 0.00480143f $X=3.705 $Y=1.765 $X2=0 $Y2=0
cc_110 N_A_c_88_n N_B_N_c_299_n 0.0253143f $X=3.81 $Y=1.385 $X2=0 $Y2=0
cc_111 N_A_c_91_n N_VPWR_c_334_n 0.0102842f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_112 N_A_c_93_n N_VPWR_c_335_n 0.00496087f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_113 N_A_c_95_n N_VPWR_c_335_n 0.00341114f $X=1.405 $Y=1.765 $X2=0 $Y2=0
cc_114 N_A_c_96_n N_VPWR_c_336_n 0.00865448f $X=3.705 $Y=1.765 $X2=0 $Y2=0
cc_115 N_A_c_95_n N_VPWR_c_339_n 0.0044313f $X=1.405 $Y=1.765 $X2=0 $Y2=0
cc_116 N_A_c_96_n N_VPWR_c_339_n 0.0044313f $X=3.705 $Y=1.765 $X2=0 $Y2=0
cc_117 N_A_c_91_n N_VPWR_c_341_n 0.00445602f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_118 N_A_c_93_n N_VPWR_c_341_n 0.00445602f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_119 N_A_c_91_n N_VPWR_c_332_n 0.00861084f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_120 N_A_c_93_n N_VPWR_c_332_n 0.00857589f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_121 N_A_c_95_n N_VPWR_c_332_n 0.00853445f $X=1.405 $Y=1.765 $X2=0 $Y2=0
cc_122 N_A_c_96_n N_VPWR_c_332_n 0.00858005f $X=3.705 $Y=1.765 $X2=0 $Y2=0
cc_123 N_A_c_91_n N_A_116_368#_c_404_n 0.00203651f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_124 N_A_c_93_n N_A_116_368#_c_404_n 4.27055e-19 $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_125 N_A_c_91_n N_A_116_368#_c_399_n 0.00993054f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_126 N_A_c_93_n N_A_116_368#_c_399_n 0.0106476f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_127 N_A_c_95_n N_A_116_368#_c_399_n 6.54713e-19 $X=1.405 $Y=1.765 $X2=0 $Y2=0
cc_128 N_A_c_93_n N_A_116_368#_c_409_n 0.0119563f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_129 N_A_c_95_n N_A_116_368#_c_409_n 0.0120074f $X=1.405 $Y=1.765 $X2=0 $Y2=0
cc_130 N_A_c_95_n N_A_116_368#_c_411_n 4.27055e-19 $X=1.405 $Y=1.765 $X2=0 $Y2=0
cc_131 N_A_c_93_n N_A_116_368#_c_412_n 6.33901e-19 $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_132 N_A_c_95_n N_A_116_368#_c_412_n 0.00949598f $X=1.405 $Y=1.765 $X2=0 $Y2=0
cc_133 N_A_c_95_n N_A_116_368#_c_401_n 0.0032261f $X=1.405 $Y=1.765 $X2=0 $Y2=0
cc_134 N_A_c_96_n N_A_116_368#_c_402_n 0.00334791f $X=3.705 $Y=1.765 $X2=0 $Y2=0
cc_135 N_A_c_96_n N_A_116_368#_c_416_n 0.0083288f $X=3.705 $Y=1.765 $X2=0 $Y2=0
cc_136 N_A_c_85_n N_Y_M1003_d 0.00176891f $X=3.645 $Y=1.095 $X2=-0.19 $Y2=-0.245
cc_137 N_A_c_85_n N_Y_M1000_d 0.00178017f $X=3.645 $Y=1.095 $X2=0 $Y2=0
cc_138 N_A_c_81_n N_Y_c_464_n 0.00666041f $X=0.955 $Y=1.675 $X2=0 $Y2=0
cc_139 N_A_c_93_n N_Y_c_464_n 0.00517623f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_140 N_A_c_82_n N_Y_c_464_n 0.0063333f $X=1.405 $Y=1.675 $X2=0 $Y2=0
cc_141 N_A_c_95_n N_Y_c_464_n 0.00516033f $X=1.405 $Y=1.765 $X2=0 $Y2=0
cc_142 N_A_c_85_n N_Y_c_464_n 0.0037097f $X=3.645 $Y=1.095 $X2=0 $Y2=0
cc_143 N_A_c_86_n N_Y_c_464_n 0.0724897f $X=1.795 $Y=1.095 $X2=0 $Y2=0
cc_144 N_A_c_89_n N_Y_c_464_n 0.00294898f $X=1.295 $Y=1.175 $X2=0 $Y2=0
cc_145 N_A_c_95_n N_Y_c_465_n 7.85716e-19 $X=1.405 $Y=1.765 $X2=0 $Y2=0
cc_146 N_A_c_85_n N_Y_c_465_n 0.0101233f $X=3.645 $Y=1.095 $X2=0 $Y2=0
cc_147 N_A_c_83_n N_Y_c_487_n 0.0110659f $X=3.51 $Y=1.22 $X2=0 $Y2=0
cc_148 N_A_c_80_n N_Y_c_466_n 0.00793544f $X=0.505 $Y=1.675 $X2=0 $Y2=0
cc_149 N_A_c_91_n N_Y_c_466_n 0.00520862f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_150 N_A_c_80_n N_Y_c_467_n 0.00398727f $X=0.505 $Y=1.675 $X2=0 $Y2=0
cc_151 N_A_c_91_n N_Y_c_467_n 0.00602937f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_152 N_A_c_81_n N_Y_c_467_n 0.00180432f $X=0.955 $Y=1.675 $X2=0 $Y2=0
cc_153 N_A_c_89_n N_Y_c_467_n 5.58672e-19 $X=1.295 $Y=1.175 $X2=0 $Y2=0
cc_154 N_A_c_85_n N_Y_c_468_n 0.105987f $X=3.645 $Y=1.095 $X2=0 $Y2=0
cc_155 N_A_c_86_n N_Y_c_468_n 0.0773139f $X=1.795 $Y=1.095 $X2=0 $Y2=0
cc_156 N_A_c_89_n N_Y_c_468_n 0.0169587f $X=1.295 $Y=1.175 $X2=0 $Y2=0
cc_157 N_A_c_83_n N_Y_c_497_n 0.00837425f $X=3.51 $Y=1.22 $X2=0 $Y2=0
cc_158 N_A_c_85_n N_Y_c_497_n 0.0155098f $X=3.645 $Y=1.095 $X2=0 $Y2=0
cc_159 N_A_c_88_n N_Y_c_497_n 4.50695e-19 $X=3.81 $Y=1.385 $X2=0 $Y2=0
cc_160 N_A_c_86_n Y 0.0114186f $X=1.795 $Y=1.095 $X2=0 $Y2=0
cc_161 N_A_c_89_n Y 0.00943558f $X=1.295 $Y=1.175 $X2=0 $Y2=0
cc_162 N_A_c_86_n Y 0.00181037f $X=1.795 $Y=1.095 $X2=0 $Y2=0
cc_163 N_A_c_89_n Y 0.0083228f $X=1.295 $Y=1.175 $X2=0 $Y2=0
cc_164 N_A_c_85_n N_VGND_M1003_s 8.73801e-19 $X=3.645 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_165 N_A_c_86_n N_VGND_M1003_s 0.00289875f $X=1.795 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_166 N_A_c_85_n N_VGND_M1008_s 0.0116574f $X=3.645 $Y=1.095 $X2=0 $Y2=0
cc_167 N_A_c_83_n N_VGND_c_560_n 7.7967e-19 $X=3.51 $Y=1.22 $X2=0 $Y2=0
cc_168 N_A_c_84_n N_VGND_c_560_n 0.0122954f $X=3.94 $Y=1.22 $X2=0 $Y2=0
cc_169 N_A_c_83_n N_VGND_c_562_n 0.00327917f $X=3.51 $Y=1.22 $X2=0 $Y2=0
cc_170 N_A_c_84_n N_VGND_c_562_n 0.00383152f $X=3.94 $Y=1.22 $X2=0 $Y2=0
cc_171 N_A_c_83_n N_VGND_c_564_n 0.00418901f $X=3.51 $Y=1.22 $X2=0 $Y2=0
cc_172 N_A_c_84_n N_VGND_c_564_n 0.0075754f $X=3.94 $Y=1.22 $X2=0 $Y2=0
cc_173 N_A_c_83_n N_VGND_c_567_n 0.00641807f $X=3.51 $Y=1.22 $X2=0 $Y2=0
cc_174 N_A_353_323#_c_203_n N_B_N_c_300_n 0.014082f $X=4.515 $Y=2.16 $X2=-0.19
+ $Y2=-0.245
cc_175 N_A_353_323#_c_194_n N_B_N_M1014_g 0.0158316f $X=4.495 $Y=1.72 $X2=0
+ $Y2=0
cc_176 N_A_353_323#_c_196_n N_B_N_M1014_g 0.00981473f $X=5 $Y=0.505 $X2=0 $Y2=0
cc_177 N_A_353_323#_c_203_n N_B_N_c_301_n 0.0142331f $X=4.515 $Y=2.16 $X2=0
+ $Y2=0
cc_178 N_A_353_323#_c_203_n B_N 0.0085076f $X=4.515 $Y=2.16 $X2=0 $Y2=0
cc_179 N_A_353_323#_c_194_n B_N 0.0416881f $X=4.495 $Y=1.72 $X2=0 $Y2=0
cc_180 N_A_353_323#_c_196_n B_N 0.0366877f $X=5 $Y=0.505 $X2=0 $Y2=0
cc_181 N_A_353_323#_c_202_n N_B_N_c_299_n 0.01494f $X=4.35 $Y=1.805 $X2=0 $Y2=0
cc_182 N_A_353_323#_c_203_n N_B_N_c_299_n 0.0185926f $X=4.515 $Y=2.16 $X2=0
+ $Y2=0
cc_183 N_A_353_323#_c_194_n N_B_N_c_299_n 0.0132547f $X=4.495 $Y=1.72 $X2=0
+ $Y2=0
cc_184 N_A_353_323#_c_196_n N_B_N_c_299_n 0.00745827f $X=5 $Y=0.505 $X2=0 $Y2=0
cc_185 N_A_353_323#_c_202_n N_VPWR_M1012_s 0.00318354f $X=4.35 $Y=1.805 $X2=0
+ $Y2=0
cc_186 N_A_353_323#_c_202_n N_VPWR_c_336_n 0.0250024f $X=4.35 $Y=1.805 $X2=0
+ $Y2=0
cc_187 N_A_353_323#_c_203_n N_VPWR_c_336_n 0.0548038f $X=4.515 $Y=2.16 $X2=0
+ $Y2=0
cc_188 N_A_353_323#_c_203_n N_VPWR_c_338_n 0.0590788f $X=4.515 $Y=2.16 $X2=0
+ $Y2=0
cc_189 N_A_353_323#_c_197_n N_VPWR_c_339_n 0.00278271f $X=1.855 $Y=1.765 $X2=0
+ $Y2=0
cc_190 N_A_353_323#_c_198_n N_VPWR_c_339_n 0.00278257f $X=2.305 $Y=1.765 $X2=0
+ $Y2=0
cc_191 N_A_353_323#_c_199_n N_VPWR_c_339_n 0.00278257f $X=2.755 $Y=1.765 $X2=0
+ $Y2=0
cc_192 N_A_353_323#_c_200_n N_VPWR_c_339_n 0.00278271f $X=3.205 $Y=1.765 $X2=0
+ $Y2=0
cc_193 N_A_353_323#_c_203_n N_VPWR_c_342_n 0.0101887f $X=4.515 $Y=2.16 $X2=0
+ $Y2=0
cc_194 N_A_353_323#_c_197_n N_VPWR_c_332_n 0.00353907f $X=1.855 $Y=1.765 $X2=0
+ $Y2=0
cc_195 N_A_353_323#_c_198_n N_VPWR_c_332_n 0.00353822f $X=2.305 $Y=1.765 $X2=0
+ $Y2=0
cc_196 N_A_353_323#_c_199_n N_VPWR_c_332_n 0.00353822f $X=2.755 $Y=1.765 $X2=0
+ $Y2=0
cc_197 N_A_353_323#_c_200_n N_VPWR_c_332_n 0.00354337f $X=3.205 $Y=1.765 $X2=0
+ $Y2=0
cc_198 N_A_353_323#_c_203_n N_VPWR_c_332_n 0.0112927f $X=4.515 $Y=2.16 $X2=0
+ $Y2=0
cc_199 N_A_353_323#_c_202_n N_A_116_368#_M1009_s 0.00250873f $X=4.35 $Y=1.805
+ $X2=0 $Y2=0
cc_200 N_A_353_323#_c_197_n N_A_116_368#_c_400_n 0.0118389f $X=1.855 $Y=1.765
+ $X2=0 $Y2=0
cc_201 N_A_353_323#_c_198_n N_A_116_368#_c_400_n 0.00879888f $X=2.305 $Y=1.765
+ $X2=0 $Y2=0
cc_202 N_A_353_323#_c_197_n N_A_116_368#_c_420_n 4.50629e-19 $X=1.855 $Y=1.765
+ $X2=0 $Y2=0
cc_203 N_A_353_323#_c_198_n N_A_116_368#_c_420_n 0.00675073f $X=2.305 $Y=1.765
+ $X2=0 $Y2=0
cc_204 N_A_353_323#_c_199_n N_A_116_368#_c_420_n 0.00667767f $X=2.755 $Y=1.765
+ $X2=0 $Y2=0
cc_205 N_A_353_323#_c_200_n N_A_116_368#_c_420_n 4.45174e-19 $X=3.205 $Y=1.765
+ $X2=0 $Y2=0
cc_206 N_A_353_323#_c_199_n N_A_116_368#_c_402_n 0.00879888f $X=2.755 $Y=1.765
+ $X2=0 $Y2=0
cc_207 N_A_353_323#_c_200_n N_A_116_368#_c_402_n 0.0137438f $X=3.205 $Y=1.765
+ $X2=0 $Y2=0
cc_208 N_A_353_323#_c_202_n N_A_116_368#_c_416_n 0.0202249f $X=4.35 $Y=1.805
+ $X2=0 $Y2=0
cc_209 N_A_353_323#_c_198_n N_A_116_368#_c_403_n 0.00174703f $X=2.305 $Y=1.765
+ $X2=0 $Y2=0
cc_210 N_A_353_323#_c_199_n N_A_116_368#_c_403_n 0.00174703f $X=2.755 $Y=1.765
+ $X2=0 $Y2=0
cc_211 N_A_353_323#_c_201_n N_Y_M1005_d 7.90456e-19 $X=3.055 $Y=1.515 $X2=0
+ $Y2=0
cc_212 N_A_353_323#_c_195_n N_Y_c_464_n 0.00994398f $X=3.06 $Y=1.515 $X2=0 $Y2=0
cc_213 N_A_353_323#_c_197_n N_Y_c_465_n 0.00734514f $X=1.855 $Y=1.765 $X2=0
+ $Y2=0
cc_214 N_A_353_323#_c_198_n N_Y_c_465_n 0.00173224f $X=2.305 $Y=1.765 $X2=0
+ $Y2=0
cc_215 N_A_353_323#_c_201_n N_Y_c_465_n 0.00838044f $X=3.055 $Y=1.515 $X2=0
+ $Y2=0
cc_216 N_A_353_323#_c_195_n N_Y_c_465_n 0.0170298f $X=3.06 $Y=1.515 $X2=0 $Y2=0
cc_217 N_A_353_323#_c_197_n N_Y_c_510_n 0.00782087f $X=1.855 $Y=1.765 $X2=0
+ $Y2=0
cc_218 N_A_353_323#_c_198_n N_Y_c_510_n 0.0055062f $X=2.305 $Y=1.765 $X2=0 $Y2=0
cc_219 N_A_353_323#_c_198_n N_Y_c_512_n 0.0119989f $X=2.305 $Y=1.765 $X2=0 $Y2=0
cc_220 N_A_353_323#_c_199_n N_Y_c_512_n 0.0117277f $X=2.755 $Y=1.765 $X2=0 $Y2=0
cc_221 N_A_353_323#_c_201_n N_Y_c_512_n 0.0223329f $X=3.055 $Y=1.515 $X2=0 $Y2=0
cc_222 N_A_353_323#_c_195_n N_Y_c_512_n 0.00286417f $X=3.06 $Y=1.515 $X2=0 $Y2=0
cc_223 N_A_353_323#_c_193_n N_Y_c_487_n 0.0105158f $X=2.44 $Y=1.225 $X2=0 $Y2=0
cc_224 N_A_353_323#_c_200_n N_Y_c_517_n 0.00181586f $X=3.205 $Y=1.765 $X2=0
+ $Y2=0
cc_225 N_A_353_323#_c_201_n N_Y_c_517_n 0.00982093f $X=3.055 $Y=1.515 $X2=0
+ $Y2=0
cc_226 N_A_353_323#_c_195_n N_Y_c_517_n 0.00296562f $X=3.06 $Y=1.515 $X2=0 $Y2=0
cc_227 N_A_353_323#_c_199_n N_Y_c_520_n 0.00489913f $X=2.755 $Y=1.765 $X2=0
+ $Y2=0
cc_228 N_A_353_323#_c_200_n N_Y_c_520_n 0.00533243f $X=3.205 $Y=1.765 $X2=0
+ $Y2=0
cc_229 N_A_353_323#_c_192_n N_Y_c_468_n 0.0105158f $X=2.01 $Y=1.225 $X2=0 $Y2=0
cc_230 N_A_353_323#_c_192_n N_Y_c_523_n 0.00718488f $X=2.01 $Y=1.225 $X2=0 $Y2=0
cc_231 N_A_353_323#_c_193_n N_Y_c_523_n 0.00718488f $X=2.44 $Y=1.225 $X2=0 $Y2=0
cc_232 N_A_353_323#_c_192_n N_VGND_c_559_n 0.00789696f $X=2.01 $Y=1.225 $X2=0
+ $Y2=0
cc_233 N_A_353_323#_c_196_n N_VGND_c_560_n 0.0217307f $X=5 $Y=0.505 $X2=0 $Y2=0
cc_234 N_A_353_323#_c_196_n N_VGND_c_563_n 0.0340697f $X=5 $Y=0.505 $X2=0 $Y2=0
cc_235 N_A_353_323#_c_192_n N_VGND_c_564_n 0.00420785f $X=2.01 $Y=1.225 $X2=0
+ $Y2=0
cc_236 N_A_353_323#_c_193_n N_VGND_c_564_n 0.00420763f $X=2.44 $Y=1.225 $X2=0
+ $Y2=0
cc_237 N_A_353_323#_c_196_n N_VGND_c_564_n 0.027759f $X=5 $Y=0.505 $X2=0 $Y2=0
cc_238 N_A_353_323#_c_192_n N_VGND_c_566_n 0.00327334f $X=2.01 $Y=1.225 $X2=0
+ $Y2=0
cc_239 N_A_353_323#_c_193_n N_VGND_c_566_n 0.00327334f $X=2.44 $Y=1.225 $X2=0
+ $Y2=0
cc_240 N_A_353_323#_c_193_n N_VGND_c_567_n 0.00845421f $X=2.44 $Y=1.225 $X2=0
+ $Y2=0
cc_241 N_B_N_c_300_n N_VPWR_c_336_n 0.0110064f $X=4.29 $Y=1.94 $X2=0 $Y2=0
cc_242 N_B_N_c_301_n N_VPWR_c_338_n 0.0112416f $X=4.74 $Y=1.94 $X2=0 $Y2=0
cc_243 B_N N_VPWR_c_338_n 0.0223353f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_244 N_B_N_c_299_n N_VPWR_c_338_n 0.00508612f $X=4.74 $Y=1.717 $X2=0 $Y2=0
cc_245 N_B_N_c_300_n N_VPWR_c_342_n 0.00491343f $X=4.29 $Y=1.94 $X2=0 $Y2=0
cc_246 N_B_N_c_301_n N_VPWR_c_342_n 0.00491343f $X=4.74 $Y=1.94 $X2=0 $Y2=0
cc_247 N_B_N_c_300_n N_VPWR_c_332_n 0.00512916f $X=4.29 $Y=1.94 $X2=0 $Y2=0
cc_248 N_B_N_c_301_n N_VPWR_c_332_n 0.00512916f $X=4.74 $Y=1.94 $X2=0 $Y2=0
cc_249 N_B_N_M1014_g N_VGND_c_560_n 0.00333403f $X=4.37 $Y=0.74 $X2=0 $Y2=0
cc_250 N_B_N_M1014_g N_VGND_c_563_n 0.00421682f $X=4.37 $Y=0.74 $X2=0 $Y2=0
cc_251 N_B_N_M1014_g N_VGND_c_564_n 0.00784929f $X=4.37 $Y=0.74 $X2=0 $Y2=0
cc_252 N_VPWR_c_334_n N_A_116_368#_c_404_n 0.0121024f $X=0.28 $Y=2.015 $X2=0
+ $Y2=0
cc_253 N_VPWR_c_334_n N_A_116_368#_c_399_n 0.0596721f $X=0.28 $Y=2.015 $X2=0
+ $Y2=0
cc_254 N_VPWR_c_335_n N_A_116_368#_c_399_n 0.0469259f $X=1.18 $Y=2.425 $X2=0
+ $Y2=0
cc_255 N_VPWR_c_341_n N_A_116_368#_c_399_n 0.014552f $X=1.095 $Y=3.33 $X2=0
+ $Y2=0
cc_256 N_VPWR_c_332_n N_A_116_368#_c_399_n 0.0119791f $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_257 N_VPWR_M1007_s N_A_116_368#_c_409_n 0.00436806f $X=1.03 $Y=1.84 $X2=0
+ $Y2=0
cc_258 N_VPWR_c_335_n N_A_116_368#_c_409_n 0.0136682f $X=1.18 $Y=2.425 $X2=0
+ $Y2=0
cc_259 N_VPWR_c_335_n N_A_116_368#_c_412_n 0.0410966f $X=1.18 $Y=2.425 $X2=0
+ $Y2=0
cc_260 N_VPWR_c_339_n N_A_116_368#_c_400_n 0.0409869f $X=3.815 $Y=3.33 $X2=0
+ $Y2=0
cc_261 N_VPWR_c_332_n N_A_116_368#_c_400_n 0.0231342f $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_262 N_VPWR_c_335_n N_A_116_368#_c_401_n 0.0119328f $X=1.18 $Y=2.425 $X2=0
+ $Y2=0
cc_263 N_VPWR_c_339_n N_A_116_368#_c_401_n 0.017869f $X=3.815 $Y=3.33 $X2=0
+ $Y2=0
cc_264 N_VPWR_c_332_n N_A_116_368#_c_401_n 0.00965079f $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_265 N_VPWR_c_336_n N_A_116_368#_c_402_n 0.0119239f $X=3.98 $Y=2.145 $X2=0
+ $Y2=0
cc_266 N_VPWR_c_339_n N_A_116_368#_c_402_n 0.062632f $X=3.815 $Y=3.33 $X2=0
+ $Y2=0
cc_267 N_VPWR_c_332_n N_A_116_368#_c_402_n 0.0347638f $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_268 N_VPWR_c_339_n N_A_116_368#_c_403_n 0.0235381f $X=3.815 $Y=3.33 $X2=0
+ $Y2=0
cc_269 N_VPWR_c_332_n N_A_116_368#_c_403_n 0.0126899f $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_270 N_VPWR_c_334_n N_Y_c_466_n 7.06399e-19 $X=0.28 $Y=2.015 $X2=0 $Y2=0
cc_271 N_VPWR_c_334_n Y 0.0184311f $X=0.28 $Y=2.015 $X2=0 $Y2=0
cc_272 N_A_116_368#_c_400_n N_Y_M1001_d 0.00205104f $X=2.365 $Y=2.99 $X2=0 $Y2=0
cc_273 N_A_116_368#_c_402_n N_Y_M1005_d 0.00205104f $X=3.315 $Y=2.99 $X2=0 $Y2=0
cc_274 N_A_116_368#_c_409_n N_Y_c_464_n 0.0361701f $X=1.465 $Y=2.005 $X2=0 $Y2=0
cc_275 N_A_116_368#_c_411_n N_Y_c_464_n 0.017918f $X=1.59 $Y=2.09 $X2=0 $Y2=0
cc_276 N_A_116_368#_c_411_n N_Y_c_465_n 0.0141101f $X=1.59 $Y=2.09 $X2=0 $Y2=0
cc_277 N_A_116_368#_c_412_n N_Y_c_465_n 0.0112687f $X=1.63 $Y=2.815 $X2=0 $Y2=0
cc_278 N_A_116_368#_c_412_n N_Y_c_510_n 0.0378702f $X=1.63 $Y=2.815 $X2=0 $Y2=0
cc_279 N_A_116_368#_c_400_n N_Y_c_510_n 0.0165699f $X=2.365 $Y=2.99 $X2=0 $Y2=0
cc_280 N_A_116_368#_c_420_n N_Y_c_510_n 0.0226573f $X=2.53 $Y=2.485 $X2=0 $Y2=0
cc_281 N_A_116_368#_M1002_s N_Y_c_512_n 0.00448603f $X=2.38 $Y=1.84 $X2=0 $Y2=0
cc_282 N_A_116_368#_c_400_n N_Y_c_512_n 0.00306905f $X=2.365 $Y=2.99 $X2=0 $Y2=0
cc_283 N_A_116_368#_c_420_n N_Y_c_512_n 0.017171f $X=2.53 $Y=2.485 $X2=0 $Y2=0
cc_284 N_A_116_368#_c_402_n N_Y_c_512_n 0.00305835f $X=3.315 $Y=2.99 $X2=0 $Y2=0
cc_285 N_A_116_368#_c_420_n N_Y_c_520_n 0.0224621f $X=2.53 $Y=2.485 $X2=0 $Y2=0
cc_286 N_A_116_368#_c_402_n N_Y_c_520_n 0.0144241f $X=3.315 $Y=2.99 $X2=0 $Y2=0
cc_287 N_A_116_368#_c_404_n N_Y_c_467_n 0.0220201f $X=0.73 $Y=2.09 $X2=0 $Y2=0
cc_288 N_Y_c_468_n N_VGND_M1003_s 0.00811085f $X=2.06 $Y=0.685 $X2=-0.19
+ $Y2=-0.245
cc_289 N_Y_c_487_n N_VGND_M1008_s 0.0210657f $X=3.56 $Y=0.755 $X2=0 $Y2=0
cc_290 N_Y_c_468_n N_VGND_c_559_n 0.0252515f $X=2.06 $Y=0.685 $X2=0 $Y2=0
cc_291 N_Y_c_463_n N_VGND_c_561_n 0.00433932f $X=0.355 $Y=0.755 $X2=0 $Y2=0
cc_292 N_Y_c_468_n N_VGND_c_561_n 0.0202416f $X=2.06 $Y=0.685 $X2=0 $Y2=0
cc_293 N_Y_c_487_n N_VGND_c_562_n 0.0023667f $X=3.56 $Y=0.755 $X2=0 $Y2=0
cc_294 N_Y_c_497_n N_VGND_c_562_n 0.00544924f $X=3.725 $Y=0.675 $X2=0 $Y2=0
cc_295 N_Y_c_463_n N_VGND_c_564_n 0.00680159f $X=0.355 $Y=0.755 $X2=0 $Y2=0
cc_296 N_Y_c_487_n N_VGND_c_564_n 0.0121701f $X=3.56 $Y=0.755 $X2=0 $Y2=0
cc_297 N_Y_c_468_n N_VGND_c_564_n 0.0390596f $X=2.06 $Y=0.685 $X2=0 $Y2=0
cc_298 N_Y_c_523_n N_VGND_c_564_n 0.0101808f $X=2.39 $Y=0.685 $X2=0 $Y2=0
cc_299 N_Y_c_497_n N_VGND_c_564_n 0.00786294f $X=3.725 $Y=0.675 $X2=0 $Y2=0
cc_300 N_Y_c_487_n N_VGND_c_566_n 0.00236055f $X=3.56 $Y=0.755 $X2=0 $Y2=0
cc_301 N_Y_c_468_n N_VGND_c_566_n 0.00236055f $X=2.06 $Y=0.685 $X2=0 $Y2=0
cc_302 N_Y_c_523_n N_VGND_c_566_n 0.00642607f $X=2.39 $Y=0.685 $X2=0 $Y2=0
cc_303 N_Y_c_487_n N_VGND_c_567_n 0.061776f $X=3.56 $Y=0.755 $X2=0 $Y2=0
