# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ls__ebufn_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ls__ebufn_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.760000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 1.300000 0.805000 1.780000 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  0.951000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.975000 1.180000 1.285000 1.550000 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  1.101200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.970000 1.820000 5.205000 1.990000 ;
        RECT 3.970000 1.990000 4.300000 2.735000 ;
        RECT 4.015000 0.595000 4.345000 0.980000 ;
        RECT 4.015000 0.980000 5.205000 1.150000 ;
        RECT 4.870000 1.990000 5.205000 2.735000 ;
        RECT 4.875000 0.595000 5.205000 0.980000 ;
        RECT 5.035000 1.150000 5.205000 1.820000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.760000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.760000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.760000 0.085000 ;
      RECT 0.000000  3.245000 5.760000 3.415000 ;
      RECT 0.085000  0.350000 0.405000 1.130000 ;
      RECT 0.085000  1.130000 0.255000 1.950000 ;
      RECT 0.085000  1.950000 0.365000 2.390000 ;
      RECT 0.085000  2.390000 1.630000 2.560000 ;
      RECT 0.085000  2.560000 0.365000 2.980000 ;
      RECT 0.565000  2.730000 0.920000 3.245000 ;
      RECT 0.585000  0.085000 0.915000 1.010000 ;
      RECT 1.040000  1.720000 1.775000 1.890000 ;
      RECT 1.040000  1.890000 1.290000 2.220000 ;
      RECT 1.095000  0.300000 1.775000 1.010000 ;
      RECT 1.455000  1.010000 1.775000 1.720000 ;
      RECT 1.460000  2.060000 2.530000 2.230000 ;
      RECT 1.460000  2.230000 1.630000 2.390000 ;
      RECT 1.800000  2.400000 2.870000 2.570000 ;
      RECT 1.800000  2.570000 1.970000 2.820000 ;
      RECT 1.945000  0.350000 2.115000 1.140000 ;
      RECT 1.945000  1.140000 3.835000 1.150000 ;
      RECT 1.945000  1.150000 2.975000 1.310000 ;
      RECT 2.170000  2.740000 2.500000 3.245000 ;
      RECT 2.295000  0.085000 2.625000 0.970000 ;
      RECT 2.360000  1.480000 4.830000 1.650000 ;
      RECT 2.360000  1.650000 2.530000 2.060000 ;
      RECT 2.700000  1.820000 3.770000 1.990000 ;
      RECT 2.700000  1.990000 2.870000 2.400000 ;
      RECT 2.700000  2.570000 2.870000 2.980000 ;
      RECT 2.805000  0.350000 2.975000 0.980000 ;
      RECT 2.805000  0.980000 3.835000 1.140000 ;
      RECT 3.070000  2.160000 3.320000 3.245000 ;
      RECT 3.155000  0.085000 3.405000 0.810000 ;
      RECT 3.520000  1.990000 3.770000 2.905000 ;
      RECT 3.520000  2.905000 5.650000 3.075000 ;
      RECT 3.585000  0.255000 5.655000 0.425000 ;
      RECT 3.585000  0.425000 3.835000 0.980000 ;
      RECT 3.820000  1.320000 4.830000 1.480000 ;
      RECT 4.470000  2.160000 4.700000 2.905000 ;
      RECT 4.525000  0.425000 4.695000 0.810000 ;
      RECT 5.400000  1.820000 5.650000 2.905000 ;
      RECT 5.405000  0.425000 5.655000 1.130000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
  END
END sky130_fd_sc_ls__ebufn_4
