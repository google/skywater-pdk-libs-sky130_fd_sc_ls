* File: sky130_fd_sc_ls__a222oi_1.pex.spice
* Created: Fri Aug 28 12:54:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__A222OI_1%C1 2 3 5 8 9 12 13 14
r32 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.43 $Y=1.285
+ $X2=0.43 $Y2=1.45
r33 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.43 $Y=1.285
+ $X2=0.43 $Y2=1.12
r34 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.43
+ $Y=1.285 $X2=0.43 $Y2=1.285
r35 9 13 3.39186 $w=6.68e-07 $l=1.9e-07 $layer=LI1_cond $X=0.24 $Y=1.455
+ $X2=0.43 $Y2=1.455
r36 8 14 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=0.52 $Y=0.69 $X2=0.52
+ $Y2=1.12
r37 3 5 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.505 $Y=1.885
+ $X2=0.505 $Y2=2.46
r38 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.505 $Y=1.795 $X2=0.505
+ $Y2=1.885
r39 2 15 134.105 $w=1.8e-07 $l=3.45e-07 $layer=POLY_cond $X=0.505 $Y=1.795
+ $X2=0.505 $Y2=1.45
.ends

.subckt PM_SKY130_FD_SC_LS__A222OI_1%C2 1 3 4 6 7 8
r34 7 8 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=1.15 $Y=1.285 $X2=1.15
+ $Y2=1.665
r35 7 12 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.15
+ $Y=1.285 $X2=1.15 $Y2=1.285
r36 4 12 87.929 $w=4.42e-07 $l=6.34035e-07 $layer=POLY_cond $X=1.005 $Y=1.885
+ $X2=1.075 $Y2=1.285
r37 4 6 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.005 $Y=1.885
+ $X2=1.005 $Y2=2.46
r38 1 12 40.4924 $w=4.42e-07 $l=2.33345e-07 $layer=POLY_cond $X=0.91 $Y=1.12
+ $X2=1.075 $Y2=1.285
r39 1 3 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=0.91 $Y=1.12 $X2=0.91
+ $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_LS__A222OI_1%B2 1 3 6 8 9 10 11 15
r38 10 11 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=2.14 $Y=1.285
+ $X2=2.14 $Y2=1.665
r39 10 15 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.14
+ $Y=1.285 $X2=2.14 $Y2=1.285
r40 9 15 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.14 $Y=1.625
+ $X2=2.14 $Y2=1.285
r41 8 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.14 $Y=1.12
+ $X2=2.14 $Y2=1.285
r42 6 8 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.23 $Y=0.69 $X2=2.23
+ $Y2=1.12
r43 1 9 45.5709 $w=2.75e-07 $l=2.95127e-07 $layer=POLY_cond $X=2.215 $Y=1.885
+ $X2=2.14 $Y2=1.625
r44 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.215 $Y=1.885
+ $X2=2.215 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_LS__A222OI_1%B1 3 4 6 8 9 10 11 15
r38 10 11 12.5122 $w=3.48e-07 $l=3.8e-07 $layer=LI1_cond $X=2.7 $Y=1.285 $X2=2.7
+ $Y2=1.665
r39 10 15 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.71
+ $Y=1.285 $X2=2.71 $Y2=1.285
r40 9 15 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.71 $Y=1.625
+ $X2=2.71 $Y2=1.285
r41 8 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.71 $Y=1.12
+ $X2=2.71 $Y2=1.285
r42 4 9 45.5709 $w=2.75e-07 $l=2.62488e-07 $layer=POLY_cond $X=2.715 $Y=1.885
+ $X2=2.71 $Y2=1.625
r43 4 6 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.715 $Y=1.885
+ $X2=2.715 $Y2=2.46
r44 3 8 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.62 $Y=0.69 $X2=2.62
+ $Y2=1.12
.ends

.subckt PM_SKY130_FD_SC_LS__A222OI_1%A1 2 3 5 8 9 10 14 15 16
r37 14 16 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=3.305 $Y=1.285
+ $X2=3.305 $Y2=1.12
r38 14 15 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.32
+ $Y=1.285 $X2=3.32 $Y2=1.285
r39 9 10 7.90266 $w=5.58e-07 $l=3.7e-07 $layer=LI1_cond $X=3.435 $Y=1.295
+ $X2=3.435 $Y2=1.665
r40 9 15 0.213585 $w=5.58e-07 $l=1e-08 $layer=LI1_cond $X=3.435 $Y=1.295
+ $X2=3.435 $Y2=1.285
r41 8 16 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.41 $Y=0.69 $X2=3.41
+ $Y2=1.12
r42 3 5 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.215 $Y=1.885
+ $X2=3.215 $Y2=2.46
r43 2 3 44.6296 $w=2.97e-07 $l=3.1682e-07 $layer=POLY_cond $X=3.305 $Y=1.61
+ $X2=3.215 $Y2=1.885
r44 1 14 2.40434 $w=3.6e-07 $l=1.5e-08 $layer=POLY_cond $X=3.305 $Y=1.3
+ $X2=3.305 $Y2=1.285
r45 1 2 49.6898 $w=3.6e-07 $l=3.1e-07 $layer=POLY_cond $X=3.305 $Y=1.3 $X2=3.305
+ $Y2=1.61
.ends

.subckt PM_SKY130_FD_SC_LS__A222OI_1%A2 3 6 7 9 10 11 18
r29 16 18 41.0924 $w=3.3e-07 $l=2.35e-07 $layer=POLY_cond $X=3.815 $Y=1.345
+ $X2=4.05 $Y2=1.345
r30 14 16 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=3.8 $Y=1.345
+ $X2=3.815 $Y2=1.345
r31 10 11 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=4.05 $Y=1.295
+ $X2=4.05 $Y2=1.665
r32 10 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.05
+ $Y=1.345 $X2=4.05 $Y2=1.345
r33 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.815 $Y=1.885
+ $X2=3.815 $Y2=2.46
r34 6 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.815 $Y=1.795 $X2=3.815
+ $Y2=1.885
r35 5 16 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.815 $Y=1.51
+ $X2=3.815 $Y2=1.345
r36 5 6 110.782 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=3.815 $Y=1.51
+ $X2=3.815 $Y2=1.795
r37 1 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.8 $Y=1.18 $X2=3.8
+ $Y2=1.345
r38 1 3 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=3.8 $Y=1.18 $X2=3.8
+ $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_LS__A222OI_1%Y 1 2 3 4 13 15 19 21 23 24 28 34 36 37 39
+ 40 41 56
r80 48 56 1.48702 $w=3.08e-07 $l=4e-08 $layer=LI1_cond $X=1.64 $Y=1.625 $X2=1.64
+ $Y2=1.665
r81 41 58 5.79065 $w=3.08e-07 $l=9.3e-08 $layer=LI1_cond $X=1.64 $Y=1.687
+ $X2=1.64 $Y2=1.78
r82 41 56 0.817863 $w=3.08e-07 $l=2.2e-08 $layer=LI1_cond $X=1.64 $Y=1.687
+ $X2=1.64 $Y2=1.665
r83 41 48 0.855038 $w=3.08e-07 $l=2.3e-08 $layer=LI1_cond $X=1.64 $Y=1.602
+ $X2=1.64 $Y2=1.625
r84 40 41 11.4129 $w=3.08e-07 $l=3.07e-07 $layer=LI1_cond $X=1.64 $Y=1.295
+ $X2=1.64 $Y2=1.602
r85 39 47 0.701276 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.64 $Y=0.865
+ $X2=1.64 $Y2=0.95
r86 39 40 11.7103 $w=3.08e-07 $l=3.15e-07 $layer=LI1_cond $X=1.64 $Y=0.98
+ $X2=1.64 $Y2=1.295
r87 39 47 1.11527 $w=3.08e-07 $l=3e-08 $layer=LI1_cond $X=1.64 $Y=0.98 $X2=1.64
+ $Y2=0.95
r88 36 37 20.0288 $w=6.18e-07 $l=6.7e-07 $layer=LI1_cond $X=3.195 $Y=0.64
+ $X2=2.525 $Y2=0.64
r89 30 39 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=1.795 $Y=0.865
+ $X2=1.64 $Y2=0.865
r90 30 37 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.795 $Y=0.865
+ $X2=2.525 $Y2=0.865
r91 28 34 2.70057 $w=3.55e-07 $l=2.23495e-07 $layer=LI1_cond $X=1.57 $Y=1.96
+ $X2=1.385 $Y2=2.045
r92 28 58 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.57 $Y=1.96
+ $X2=1.57 $Y2=1.78
r93 23 39 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=1.485 $Y=0.865
+ $X2=1.64 $Y2=0.865
r94 23 24 66.2193 $w=1.68e-07 $l=1.015e-06 $layer=LI1_cond $X=1.485 $Y=0.865
+ $X2=0.47 $Y2=0.865
r95 22 32 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.445 $Y=2.045
+ $X2=0.28 $Y2=2.045
r96 21 34 4.08752 $w=1.7e-07 $l=2.7e-07 $layer=LI1_cond $X=1.115 $Y=2.045
+ $X2=1.385 $Y2=2.045
r97 21 22 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.115 $Y=2.045
+ $X2=0.445 $Y2=2.045
r98 17 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.305 $Y=0.78
+ $X2=0.47 $Y2=0.865
r99 17 19 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=0.305 $Y=0.78
+ $X2=0.305 $Y2=0.515
r100 13 32 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.28 $Y=2.13 $X2=0.28
+ $Y2=2.045
r101 13 15 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=0.28 $Y=2.13
+ $X2=0.28 $Y2=2.815
r102 4 34 300 $w=1.7e-07 $l=2.70185e-07 $layer=licon1_PDIFF $count=2 $X=1.08
+ $Y=1.96 $X2=1.28 $Y2=2.125
r103 3 32 400 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.28 $Y2=2.125
r104 3 15 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.28 $Y2=2.815
r105 2 36 45.5 $w=1.7e-07 $l=5.59017e-07 $layer=licon1_NDIFF $count=4 $X=2.695
+ $Y=0.37 $X2=3.195 $Y2=0.495
r106 1 19 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.16
+ $Y=0.37 $X2=0.305 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__A222OI_1%A_116_392# 1 2 9 11 12 15
r25 13 15 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=2.49 $Y=2.905
+ $X2=2.49 $Y2=2.465
r26 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.325 $Y=2.99
+ $X2=2.49 $Y2=2.905
r27 11 12 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.325 $Y=2.99
+ $X2=0.945 $Y2=2.99
r28 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.78 $Y=2.905
+ $X2=0.945 $Y2=2.99
r29 7 9 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=0.78 $Y=2.905 $X2=0.78
+ $Y2=2.465
r30 2 15 300 $w=1.7e-07 $l=5.96678e-07 $layer=licon1_PDIFF $count=2 $X=2.29
+ $Y=1.96 $X2=2.49 $Y2=2.465
r31 1 9 300 $w=1.7e-07 $l=5.96678e-07 $layer=licon1_PDIFF $count=2 $X=0.58
+ $Y=1.96 $X2=0.78 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LS__A222OI_1%A_369_392# 1 2 3 12 16 18 20 22 25 27
r43 20 29 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.04 $Y=2.13 $X2=4.04
+ $Y2=2.045
r44 20 22 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=4.04 $Y=2.13
+ $X2=4.04 $Y2=2.815
r45 19 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.155 $Y=2.045
+ $X2=2.99 $Y2=2.045
r46 18 29 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.875 $Y=2.045
+ $X2=4.04 $Y2=2.045
r47 18 19 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=3.875 $Y=2.045
+ $X2=3.155 $Y2=2.045
r48 14 27 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.99 $Y=2.13 $X2=2.99
+ $Y2=2.045
r49 14 16 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=2.99 $Y=2.13
+ $X2=2.99 $Y2=2.815
r50 13 25 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.155 $Y=2.045
+ $X2=1.99 $Y2=2.045
r51 12 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.825 $Y=2.045
+ $X2=2.99 $Y2=2.045
r52 12 13 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.825 $Y=2.045
+ $X2=2.155 $Y2=2.045
r53 3 29 400 $w=1.7e-07 $l=2.2798e-07 $layer=licon1_PDIFF $count=1 $X=3.89
+ $Y=1.96 $X2=4.04 $Y2=2.125
r54 3 22 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=3.89
+ $Y=1.96 $X2=4.04 $Y2=2.815
r55 2 27 400 $w=1.7e-07 $l=2.70185e-07 $layer=licon1_PDIFF $count=1 $X=2.79
+ $Y=1.96 $X2=2.99 $Y2=2.125
r56 2 16 400 $w=1.7e-07 $l=9.4975e-07 $layer=licon1_PDIFF $count=1 $X=2.79
+ $Y=1.96 $X2=2.99 $Y2=2.815
r57 1 25 300 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_PDIFF $count=2 $X=1.845
+ $Y=1.96 $X2=1.99 $Y2=2.125
.ends

.subckt PM_SKY130_FD_SC_LS__A222OI_1%VPWR 1 6 9 10 11 21 22
r35 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r36 19 22 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r37 18 19 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r38 14 18 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=3.12 $Y2=3.33
r39 14 15 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r40 11 19 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r41 11 15 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=0.24 $Y2=3.33
r42 9 18 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=3.325 $Y=3.33
+ $X2=3.12 $Y2=3.33
r43 9 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.325 $Y=3.33
+ $X2=3.49 $Y2=3.33
r44 8 21 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=3.655 $Y=3.33
+ $X2=4.08 $Y2=3.33
r45 8 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.655 $Y=3.33
+ $X2=3.49 $Y2=3.33
r46 4 10 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.49 $Y=3.245 $X2=3.49
+ $Y2=3.33
r47 4 6 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=3.49 $Y=3.245 $X2=3.49
+ $Y2=2.465
r48 1 6 300 $w=1.7e-07 $l=5.96678e-07 $layer=licon1_PDIFF $count=2 $X=3.29
+ $Y=1.96 $X2=3.49 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LS__A222OI_1%VGND 1 2 7 9 11 18 25 37 40
r42 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r43 35 37 8.17678 $w=6.83e-07 $l=2e-08 $layer=LI1_cond $X=2.16 $Y=0.257 $X2=2.18
+ $Y2=0.257
r44 33 35 2.53184 $w=6.83e-07 $l=1.45e-07 $layer=LI1_cond $X=2.015 $Y=0.257
+ $X2=2.16 $Y2=0.257
r45 30 33 5.84943 $w=6.83e-07 $l=3.35e-07 $layer=LI1_cond $X=1.68 $Y=0.257
+ $X2=2.015 $Y2=0.257
r46 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r47 28 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r48 27 30 8.38128 $w=6.83e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=0.257
+ $X2=1.68 $Y2=0.257
r49 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r50 24 27 1.30957 $w=6.83e-07 $l=7.5e-08 $layer=LI1_cond $X=1.125 $Y=0.257
+ $X2=1.2 $Y2=0.257
r51 24 25 10.7086 $w=6.83e-07 $l=1.65e-07 $layer=LI1_cond $X=1.125 $Y=0.257
+ $X2=0.96 $Y2=0.257
r52 22 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r53 21 37 92.6417 $w=1.68e-07 $l=1.42e-06 $layer=LI1_cond $X=3.6 $Y=0 $X2=2.18
+ $Y2=0
r54 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r55 18 39 4.67962 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=3.85 $Y=0 $X2=4.085
+ $Y2=0
r56 18 21 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.85 $Y=0 $X2=3.6
+ $Y2=0
r57 16 28 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r58 15 25 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=0.96
+ $Y2=0
r59 15 16 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r60 11 22 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.6
+ $Y2=0
r61 11 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r62 11 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r63 7 39 3.08656 $w=3.3e-07 $l=1.14782e-07 $layer=LI1_cond $X=4.015 $Y=0.085
+ $X2=4.085 $Y2=0
r64 7 9 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=4.015 $Y=0.085
+ $X2=4.015 $Y2=0.515
r65 2 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.875
+ $Y=0.37 $X2=4.015 $Y2=0.515
r66 1 33 121.333 $w=1.7e-07 $l=1.10011e-06 $layer=licon1_NDIFF $count=1 $X=0.985
+ $Y=0.37 $X2=2.015 $Y2=0.515
r67 1 24 121.333 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=0.985
+ $Y=0.37 $X2=1.125 $Y2=0.515
.ends

