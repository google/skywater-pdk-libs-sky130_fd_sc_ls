* File: sky130_fd_sc_ls__or3b_4.pex.spice
* Created: Wed Sep  2 11:25:20 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__OR3B_4%C_N 1 2 3 5 9 11 13 20 21
c37 3 0 1.15346e-19 $X=0.5 $Y=1.885
r38 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.61
+ $Y=0.405 $X2=0.61 $Y2=0.405
r39 18 20 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=0.515 $Y=0.405
+ $X2=0.61 $Y2=0.405
r40 16 21 10.1774 $w=3.83e-07 $l=3.4e-07 $layer=LI1_cond $X=0.27 $Y=0.447
+ $X2=0.61 $Y2=0.447
r41 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=0.405 $X2=0.27 $Y2=0.405
r42 13 18 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=0.44 $Y=0.405
+ $X2=0.515 $Y2=0.405
r43 13 15 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=0.44 $Y=0.405
+ $X2=0.27 $Y2=0.405
r44 11 16 0.898008 $w=3.83e-07 $l=3e-08 $layer=LI1_cond $X=0.24 $Y=0.447
+ $X2=0.27 $Y2=0.447
r45 9 10 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.515 $Y=1 $X2=0.515
+ $Y2=1.395
r46 6 18 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.515 $Y=0.57
+ $X2=0.515 $Y2=0.405
r47 6 9 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=0.515 $Y=0.57
+ $X2=0.515 $Y2=1
r48 3 5 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.5 $Y=1.885 $X2=0.5
+ $Y2=2.46
r49 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.5 $Y=1.795 $X2=0.5
+ $Y2=1.885
r50 1 10 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.5 $Y=1.485 $X2=0.5
+ $Y2=1.395
r51 1 2 120.5 $w=1.8e-07 $l=3.1e-07 $layer=POLY_cond $X=0.5 $Y=1.485 $X2=0.5
+ $Y2=1.795
.ends

.subckt PM_SKY130_FD_SC_LS__OR3B_4%A 1 3 6 8 9 11 14 17 18 19 23 25
c93 9 0 6.96018e-20 $X=3.405 $Y=1.885
r94 23 26 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.45 $Y=1.385
+ $X2=3.45 $Y2=1.55
r95 23 25 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.45 $Y=1.385
+ $X2=3.45 $Y2=1.22
r96 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.45
+ $Y=1.385 $X2=3.45 $Y2=1.385
r97 19 24 12.9453 $w=3.11e-07 $l=3.3e-07 $layer=LI1_cond $X=3.12 $Y=1.35
+ $X2=3.45 $Y2=1.35
r98 17 19 7.00102 $w=3.11e-07 $l=1.62635e-07 $layer=LI1_cond $X=3.005 $Y=1.235
+ $X2=3.12 $Y2=1.35
r99 17 18 122.326 $w=1.68e-07 $l=1.875e-06 $layer=LI1_cond $X=3.005 $Y=1.235
+ $X2=1.13 $Y2=1.235
r100 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.965
+ $Y=1.595 $X2=0.965 $Y2=1.595
r101 12 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.965 $Y=1.32
+ $X2=1.13 $Y2=1.235
r102 12 14 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=0.965 $Y=1.32
+ $X2=0.965 $Y2=1.595
r103 9 11 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.405 $Y=1.885
+ $X2=3.405 $Y2=2.46
r104 8 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.405 $Y=1.795
+ $X2=3.405 $Y2=1.885
r105 8 26 95.2339 $w=1.8e-07 $l=2.45e-07 $layer=POLY_cond $X=3.405 $Y=1.795
+ $X2=3.405 $Y2=1.55
r106 6 25 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.39 $Y=0.74 $X2=3.39
+ $Y2=1.22
r107 1 15 59.5544 $w=2.88e-07 $l=3.11689e-07 $layer=POLY_cond $X=1.01 $Y=1.885
+ $X2=0.965 $Y2=1.595
r108 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.01 $Y=1.885
+ $X2=1.01 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_LS__OR3B_4%B 1 3 4 6 9 11 12 13 23 26 37
c64 9 0 1.44963e-19 $X=2.96 $Y=0.74
r65 26 37 0.460977 $w=2.48e-07 $l=1e-08 $layer=LI1_cond $X=1.68 $Y=1.675
+ $X2=1.67 $Y2=1.675
r66 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.91
+ $Y=1.635 $X2=2.91 $Y2=1.635
r67 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.505
+ $Y=1.635 $X2=1.505 $Y2=1.635
r68 13 23 12.4464 $w=2.48e-07 $l=2.7e-07 $layer=LI1_cond $X=2.64 $Y=1.675
+ $X2=2.91 $Y2=1.675
r69 12 13 22.1269 $w=2.48e-07 $l=4.8e-07 $layer=LI1_cond $X=2.16 $Y=1.675
+ $X2=2.64 $Y2=1.675
r70 11 37 1.87799 $w=3.08e-07 $l=3.8e-08 $layer=LI1_cond $X=1.632 $Y=1.645
+ $X2=1.67 $Y2=1.645
r71 11 20 4.7213 $w=3.08e-07 $l=1.27e-07 $layer=LI1_cond $X=1.632 $Y=1.645
+ $X2=1.505 $Y2=1.645
r72 11 12 20.4213 $w=2.48e-07 $l=4.43e-07 $layer=LI1_cond $X=1.717 $Y=1.675
+ $X2=2.16 $Y2=1.675
r73 11 26 1.70562 $w=2.48e-07 $l=3.7e-08 $layer=LI1_cond $X=1.717 $Y=1.675
+ $X2=1.68 $Y2=1.675
r74 7 22 38.5562 $w=2.99e-07 $l=1.88348e-07 $layer=POLY_cond $X=2.96 $Y=1.47
+ $X2=2.91 $Y2=1.635
r75 7 9 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=2.96 $Y=1.47 $X2=2.96
+ $Y2=0.74
r76 4 22 52.2586 $w=2.99e-07 $l=2.57391e-07 $layer=POLY_cond $X=2.895 $Y=1.885
+ $X2=2.91 $Y2=1.635
r77 4 6 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.895 $Y=1.885
+ $X2=2.895 $Y2=2.46
r78 1 19 52.2586 $w=2.99e-07 $l=2.7157e-07 $layer=POLY_cond $X=1.46 $Y=1.885
+ $X2=1.505 $Y2=1.635
r79 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.46 $Y=1.885
+ $X2=1.46 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_LS__OR3B_4%A_27_392# 1 2 8 10 11 13 14 17 18 20 21 23 24
+ 25 29 32 36 37 40 41 43
r93 41 46 88.9594 $w=4.5e-07 $l=5.05e-07 $layer=POLY_cond $X=1.805 $Y=0.475
+ $X2=1.805 $Y2=0.98
r94 40 41 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.745
+ $Y=0.475 $X2=1.745 $Y2=0.475
r95 38 40 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.745 $Y=0.81
+ $X2=1.745 $Y2=0.475
r96 36 38 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.58 $Y=0.895
+ $X2=1.745 $Y2=0.81
r97 36 37 72.7433 $w=1.68e-07 $l=1.115e-06 $layer=LI1_cond $X=1.58 $Y=0.895
+ $X2=0.465 $Y2=0.895
r98 32 34 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=0.235 $Y=2.105
+ $X2=0.235 $Y2=2.815
r99 32 43 35.2648 $w=2.48e-07 $l=7.65e-07 $layer=LI1_cond $X=0.235 $Y=2.105
+ $X2=0.235 $Y2=1.34
r100 27 43 6.76842 $w=3.53e-07 $l=1.77e-07 $layer=LI1_cond $X=0.287 $Y=1.163
+ $X2=0.287 $Y2=1.34
r101 27 29 2.85676 $w=3.53e-07 $l=8.8e-08 $layer=LI1_cond $X=0.287 $Y=1.163
+ $X2=0.287 $Y2=1.075
r102 26 37 7.97992 $w=1.7e-07 $l=2.16365e-07 $layer=LI1_cond $X=0.287 $Y=0.98
+ $X2=0.465 $Y2=0.895
r103 26 29 3.084 $w=3.53e-07 $l=9.5e-08 $layer=LI1_cond $X=0.287 $Y=0.98
+ $X2=0.287 $Y2=1.075
r104 21 25 18.8402 $w=1.65e-07 $l=8.21584e-08 $layer=POLY_cond $X=2.46 $Y=1.185
+ $X2=2.445 $Y2=1.26
r105 21 23 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.46 $Y=1.185
+ $X2=2.46 $Y2=0.74
r106 18 20 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.445 $Y=1.885
+ $X2=2.445 $Y2=2.46
r107 17 18 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.445 $Y=1.795
+ $X2=2.445 $Y2=1.885
r108 16 25 18.8402 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=2.445 $Y=1.335
+ $X2=2.445 $Y2=1.26
r109 16 17 178.806 $w=1.8e-07 $l=4.6e-07 $layer=POLY_cond $X=2.445 $Y=1.335
+ $X2=2.445 $Y2=1.795
r110 15 24 6.66866 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.06 $Y=1.26 $X2=1.97
+ $Y2=1.26
r111 14 25 6.66866 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.355 $Y=1.26
+ $X2=2.445 $Y2=1.26
r112 14 15 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=2.355 $Y=1.26
+ $X2=2.06 $Y2=1.26
r113 11 13 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.97 $Y=1.885
+ $X2=1.97 $Y2=2.46
r114 10 11 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.97 $Y=1.795
+ $X2=1.97 $Y2=1.885
r115 9 24 18.8402 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=1.97 $Y=1.335
+ $X2=1.97 $Y2=1.26
r116 9 10 178.806 $w=1.8e-07 $l=4.6e-07 $layer=POLY_cond $X=1.97 $Y=1.335
+ $X2=1.97 $Y2=1.795
r117 8 24 18.8402 $w=1.65e-07 $l=8.21584e-08 $layer=POLY_cond $X=1.955 $Y=1.185
+ $X2=1.97 $Y2=1.26
r118 8 46 105.117 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=1.955 $Y=1.185
+ $X2=1.955 $Y2=0.98
r119 2 34 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.275 $Y2=2.815
r120 2 32 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.275 $Y2=2.105
r121 1 29 182 $w=1.7e-07 $l=4.61844e-07 $layer=licon1_NDIFF $count=1 $X=0.155
+ $Y=0.68 $X2=0.3 $Y2=1.075
.ends

.subckt PM_SKY130_FD_SC_LS__OR3B_4%A_409_392# 1 2 3 12 14 16 19 21 23 24 26 29
+ 33 35 37 40 42 44 45 48 50 53 55 61 67 69 70 79
c160 48 0 1.44963e-19 $X=3.175 $Y=0.515
r161 76 77 2.45293 $w=3.93e-07 $l=2e-08 $layer=POLY_cond $X=4.815 $Y=1.532
+ $X2=4.835 $Y2=1.532
r162 75 76 55.1908 $w=3.93e-07 $l=4.5e-07 $layer=POLY_cond $X=4.365 $Y=1.532
+ $X2=4.815 $Y2=1.532
r163 74 75 1.22646 $w=3.93e-07 $l=1e-08 $layer=POLY_cond $X=4.355 $Y=1.532
+ $X2=4.365 $Y2=1.532
r164 71 72 1.83969 $w=3.93e-07 $l=1.5e-08 $layer=POLY_cond $X=3.9 $Y=1.532
+ $X2=3.915 $Y2=1.532
r165 65 67 10.0544 $w=2.18e-07 $l=1.8e-07 $layer=LI1_cond $X=2.205 $Y=2.08
+ $X2=2.385 $Y2=2.08
r166 62 79 31.2748 $w=3.93e-07 $l=2.55e-07 $layer=POLY_cond $X=5.01 $Y=1.532
+ $X2=5.265 $Y2=1.532
r167 62 77 21.4631 $w=3.93e-07 $l=1.75e-07 $layer=POLY_cond $X=5.01 $Y=1.532
+ $X2=4.835 $Y2=1.532
r168 61 62 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.01
+ $Y=1.465 $X2=5.01 $Y2=1.465
r169 59 74 44.7659 $w=3.93e-07 $l=3.65e-07 $layer=POLY_cond $X=3.99 $Y=1.532
+ $X2=4.355 $Y2=1.532
r170 59 72 9.19847 $w=3.93e-07 $l=7.5e-08 $layer=POLY_cond $X=3.99 $Y=1.532
+ $X2=3.915 $Y2=1.532
r171 58 61 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=3.99 $Y=1.465
+ $X2=5.01 $Y2=1.465
r172 58 59 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.99
+ $Y=1.465 $X2=3.99 $Y2=1.465
r173 56 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.885 $Y=1.465
+ $X2=3.8 $Y2=1.465
r174 56 58 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=3.885 $Y=1.465
+ $X2=3.99 $Y2=1.465
r175 54 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.8 $Y=1.63 $X2=3.8
+ $Y2=1.465
r176 54 55 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=3.8 $Y=1.63 $X2=3.8
+ $Y2=1.97
r177 53 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.8 $Y=1.3 $X2=3.8
+ $Y2=1.465
r178 52 53 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=3.8 $Y=0.98 $X2=3.8
+ $Y2=1.3
r179 51 69 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.34 $Y=0.895
+ $X2=3.215 $Y2=0.895
r180 50 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.715 $Y=0.895
+ $X2=3.8 $Y2=0.98
r181 50 51 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=3.715 $Y=0.895
+ $X2=3.34 $Y2=0.895
r182 46 69 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.215 $Y=0.81
+ $X2=3.215 $Y2=0.895
r183 46 48 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=3.215 $Y=0.81
+ $X2=3.215 $Y2=0.515
r184 44 69 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.09 $Y=0.895
+ $X2=3.215 $Y2=0.895
r185 44 45 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.09 $Y=0.895
+ $X2=2.41 $Y2=0.895
r186 42 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.715 $Y=2.055
+ $X2=3.8 $Y2=1.97
r187 42 67 86.7701 $w=1.68e-07 $l=1.33e-06 $layer=LI1_cond $X=3.715 $Y=2.055
+ $X2=2.385 $Y2=2.055
r188 38 45 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.245 $Y=0.81
+ $X2=2.41 $Y2=0.895
r189 38 40 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.245 $Y=0.81
+ $X2=2.245 $Y2=0.515
r190 35 79 25.4309 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=5.265 $Y=1.765
+ $X2=5.265 $Y2=1.532
r191 35 37 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.265 $Y=1.765
+ $X2=5.265 $Y2=2.4
r192 31 79 25.4309 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=5.265 $Y=1.3
+ $X2=5.265 $Y2=1.532
r193 31 33 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=5.265 $Y=1.3
+ $X2=5.265 $Y2=0.74
r194 27 77 25.4309 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=4.835 $Y=1.3
+ $X2=4.835 $Y2=1.532
r195 27 29 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.835 $Y=1.3
+ $X2=4.835 $Y2=0.74
r196 24 76 25.4309 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=4.815 $Y=1.765
+ $X2=4.815 $Y2=1.532
r197 24 26 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.815 $Y=1.765
+ $X2=4.815 $Y2=2.4
r198 21 75 25.4309 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=4.365 $Y=1.765
+ $X2=4.365 $Y2=1.532
r199 21 23 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.365 $Y=1.765
+ $X2=4.365 $Y2=2.4
r200 17 74 25.4309 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=4.355 $Y=1.3
+ $X2=4.355 $Y2=1.532
r201 17 19 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.355 $Y=1.3
+ $X2=4.355 $Y2=0.74
r202 14 72 25.4309 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=3.915 $Y=1.765
+ $X2=3.915 $Y2=1.532
r203 14 16 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.915 $Y=1.765
+ $X2=3.915 $Y2=2.4
r204 10 71 25.4309 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=3.9 $Y=1.3 $X2=3.9
+ $Y2=1.532
r205 10 12 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.9 $Y=1.3 $X2=3.9
+ $Y2=0.74
r206 3 65 600 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_PDIFF $count=1 $X=2.045
+ $Y=1.96 $X2=2.205 $Y2=2.105
r207 2 69 182 $w=1.7e-07 $l=5.90868e-07 $layer=licon1_NDIFF $count=1 $X=3.035
+ $Y=0.37 $X2=3.175 $Y2=0.895
r208 2 48 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.035
+ $Y=0.37 $X2=3.175 $Y2=0.515
r209 1 40 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.105
+ $Y=0.37 $X2=2.245 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__OR3B_4%VPWR 1 2 3 4 15 21 25 27 29 31 33 38 46 51 57
+ 60 63 67
r72 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r73 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r74 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r75 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r76 55 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r77 55 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r78 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r79 52 63 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.675 $Y=3.33
+ $X2=4.55 $Y2=3.33
r80 52 54 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=4.675 $Y=3.33
+ $X2=5.04 $Y2=3.33
r81 51 66 4.02656 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=5.405 $Y=3.33
+ $X2=5.582 $Y2=3.33
r82 51 54 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=5.405 $Y=3.33
+ $X2=5.04 $Y2=3.33
r83 50 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r84 50 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r85 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r86 47 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.835 $Y=3.33
+ $X2=3.67 $Y2=3.33
r87 47 49 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=3.835 $Y=3.33
+ $X2=4.08 $Y2=3.33
r88 46 63 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.425 $Y=3.33
+ $X2=4.55 $Y2=3.33
r89 46 49 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=4.425 $Y=3.33
+ $X2=4.08 $Y2=3.33
r90 45 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r91 44 45 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r92 42 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r93 41 44 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=3.12 $Y2=3.33
r94 41 42 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r95 39 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.89 $Y=3.33
+ $X2=0.725 $Y2=3.33
r96 39 41 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.89 $Y=3.33 $X2=1.2
+ $Y2=3.33
r97 38 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.505 $Y=3.33
+ $X2=3.67 $Y2=3.33
r98 38 44 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=3.505 $Y=3.33
+ $X2=3.12 $Y2=3.33
r99 36 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r100 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r101 33 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.56 $Y=3.33
+ $X2=0.725 $Y2=3.33
r102 33 35 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.56 $Y=3.33
+ $X2=0.24 $Y2=3.33
r103 31 45 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=3.12 $Y2=3.33
r104 31 42 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=1.2 $Y2=3.33
r105 27 66 3.1166 $w=2.5e-07 $l=1.07912e-07 $layer=LI1_cond $X=5.53 $Y=3.245
+ $X2=5.582 $Y2=3.33
r106 27 29 43.3319 $w=2.48e-07 $l=9.4e-07 $layer=LI1_cond $X=5.53 $Y=3.245
+ $X2=5.53 $Y2=2.305
r107 23 63 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.55 $Y=3.245
+ $X2=4.55 $Y2=3.33
r108 23 25 43.3319 $w=2.48e-07 $l=9.4e-07 $layer=LI1_cond $X=4.55 $Y=3.245
+ $X2=4.55 $Y2=2.305
r109 19 60 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.67 $Y=3.245
+ $X2=3.67 $Y2=3.33
r110 19 21 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=3.67 $Y=3.245
+ $X2=3.67 $Y2=2.475
r111 15 18 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.725 $Y=2.105
+ $X2=0.725 $Y2=2.815
r112 13 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.725 $Y=3.245
+ $X2=0.725 $Y2=3.33
r113 13 18 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.725 $Y=3.245
+ $X2=0.725 $Y2=2.815
r114 4 29 300 $w=1.7e-07 $l=5.34766e-07 $layer=licon1_PDIFF $count=2 $X=5.34
+ $Y=1.84 $X2=5.49 $Y2=2.305
r115 3 25 300 $w=1.7e-07 $l=5.34766e-07 $layer=licon1_PDIFF $count=2 $X=4.44
+ $Y=1.84 $X2=4.59 $Y2=2.305
r116 2 21 300 $w=1.7e-07 $l=6.02557e-07 $layer=licon1_PDIFF $count=2 $X=3.48
+ $Y=1.96 $X2=3.67 $Y2=2.475
r117 1 18 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=0.575
+ $Y=1.96 $X2=0.725 $Y2=2.815
r118 1 15 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=0.575
+ $Y=1.96 $X2=0.725 $Y2=2.105
.ends

.subckt PM_SKY130_FD_SC_LS__OR3B_4%A_217_392# 1 2 9 13 15 19 21
c38 13 0 1.15346e-19 $X=1.235 $Y=2.815
r39 16 19 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.4 $Y=2.445
+ $X2=1.235 $Y2=2.445
r40 15 21 4.91858 $w=1.7e-07 $l=1.77059e-07 $layer=LI1_cond $X=3.005 $Y=2.445
+ $X2=3.17 $Y2=2.42
r41 15 16 104.711 $w=1.68e-07 $l=1.605e-06 $layer=LI1_cond $X=3.005 $Y=2.445
+ $X2=1.4 $Y2=2.445
r42 11 19 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.235 $Y=2.53
+ $X2=1.235 $Y2=2.445
r43 11 13 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=1.235 $Y=2.53
+ $X2=1.235 $Y2=2.815
r44 7 19 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.235 $Y=2.36
+ $X2=1.235 $Y2=2.445
r45 7 9 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=1.235 $Y=2.36
+ $X2=1.235 $Y2=2.135
r46 2 21 300 $w=1.7e-07 $l=6.06815e-07 $layer=licon1_PDIFF $count=2 $X=2.97
+ $Y=1.96 $X2=3.17 $Y2=2.475
r47 1 13 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=1.085
+ $Y=1.96 $X2=1.235 $Y2=2.815
r48 1 9 400 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=1 $X=1.085
+ $Y=1.96 $X2=1.235 $Y2=2.135
.ends

.subckt PM_SKY130_FD_SC_LS__OR3B_4%A_307_392# 1 2 11
c14 11 0 6.96018e-20 $X=2.67 $Y=2.8
r15 8 11 38.0718 $w=2.78e-07 $l=9.25e-07 $layer=LI1_cond $X=1.745 $Y=2.84
+ $X2=2.67 $Y2=2.84
r16 2 11 600 $w=1.7e-07 $l=9.11921e-07 $layer=licon1_PDIFF $count=1 $X=2.52
+ $Y=1.96 $X2=2.67 $Y2=2.8
r17 1 8 600 $w=1.7e-07 $l=9.39149e-07 $layer=licon1_PDIFF $count=1 $X=1.535
+ $Y=1.96 $X2=1.745 $Y2=2.8
.ends

.subckt PM_SKY130_FD_SC_LS__OR3B_4%X 1 2 3 4 15 19 23 24 25 26 29 35 37 39 41 42
+ 45 46
r83 45 46 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=5.52 $Y=1.295
+ $X2=5.52 $Y2=1.665
r84 44 46 6.76434 $w=2.28e-07 $l=1.35e-07 $layer=LI1_cond $X=5.52 $Y=1.8
+ $X2=5.52 $Y2=1.665
r85 43 45 8.26753 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=5.52 $Y=1.13
+ $X2=5.52 $Y2=1.295
r86 40 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.205 $Y=1.885
+ $X2=5.04 $Y2=1.885
r87 39 44 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=5.405 $Y=1.885
+ $X2=5.52 $Y2=1.8
r88 39 40 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=5.405 $Y=1.885
+ $X2=5.205 $Y2=1.885
r89 38 42 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.135 $Y=1.045
+ $X2=5.01 $Y2=1.045
r90 37 43 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=5.405 $Y=1.045
+ $X2=5.52 $Y2=1.13
r91 37 38 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=5.405 $Y=1.045
+ $X2=5.135 $Y2=1.045
r92 33 42 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.01 $Y=0.96
+ $X2=5.01 $Y2=1.045
r93 33 35 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=5.01 $Y=0.96
+ $X2=5.01 $Y2=0.515
r94 29 31 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=5.04 $Y=1.985
+ $X2=5.04 $Y2=2.815
r95 27 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.04 $Y=1.97 $X2=5.04
+ $Y2=1.885
r96 27 29 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=5.04 $Y=1.97
+ $X2=5.04 $Y2=1.985
r97 25 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.875 $Y=1.885
+ $X2=5.04 $Y2=1.885
r98 25 26 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=4.875 $Y=1.885
+ $X2=4.225 $Y2=1.885
r99 23 42 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.885 $Y=1.045
+ $X2=5.01 $Y2=1.045
r100 23 24 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=4.885 $Y=1.045
+ $X2=4.225 $Y2=1.045
r101 19 21 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=4.14 $Y=1.985
+ $X2=4.14 $Y2=2.815
r102 17 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.14 $Y=1.97
+ $X2=4.225 $Y2=1.885
r103 17 19 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=4.14 $Y=1.97
+ $X2=4.14 $Y2=1.985
r104 13 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.14 $Y=0.96
+ $X2=4.225 $Y2=1.045
r105 13 15 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=4.14 $Y=0.96
+ $X2=4.14 $Y2=0.515
r106 4 31 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=4.89
+ $Y=1.84 $X2=5.04 $Y2=2.815
r107 4 29 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=4.89
+ $Y=1.84 $X2=5.04 $Y2=1.985
r108 3 21 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=3.99
+ $Y=1.84 $X2=4.14 $Y2=2.815
r109 3 19 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=3.99
+ $Y=1.84 $X2=4.14 $Y2=1.985
r110 2 35 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.91
+ $Y=0.37 $X2=5.05 $Y2=0.515
r111 1 15 91 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=2 $X=3.975
+ $Y=0.37 $X2=4.14 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__OR3B_4%VGND 1 2 3 4 5 18 22 26 30 32 34 36 38 43 48
+ 53 58 64 67 70 73 77
r87 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r88 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r89 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r90 67 68 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r91 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r92 62 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r93 62 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.56
+ $Y2=0
r94 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r95 59 73 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.655 $Y=0 $X2=4.53
+ $Y2=0
r96 59 61 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=4.655 $Y=0 $X2=5.04
+ $Y2=0
r97 58 76 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=5.315 $Y=0 $X2=5.537
+ $Y2=0
r98 58 61 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=5.315 $Y=0 $X2=5.04
+ $Y2=0
r99 57 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r100 57 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r101 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r102 54 70 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=3.85 $Y=0 $X2=3.68
+ $Y2=0
r103 54 56 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=3.85 $Y=0 $X2=4.08
+ $Y2=0
r104 53 73 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.405 $Y=0 $X2=4.53
+ $Y2=0
r105 53 56 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=4.405 $Y=0
+ $X2=4.08 $Y2=0
r106 52 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r107 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r108 49 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.91 $Y=0 $X2=2.745
+ $Y2=0
r109 49 51 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=2.91 $Y=0 $X2=3.12
+ $Y2=0
r110 48 70 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=3.51 $Y=0 $X2=3.68
+ $Y2=0
r111 48 51 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=3.51 $Y=0 $X2=3.12
+ $Y2=0
r112 47 68 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r113 47 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r114 46 47 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r115 44 64 10.8012 $w=1.7e-07 $l=2.33e-07 $layer=LI1_cond $X=1.41 $Y=0 $X2=1.177
+ $Y2=0
r116 44 46 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=1.41 $Y=0 $X2=1.68
+ $Y2=0
r117 43 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.58 $Y=0 $X2=2.745
+ $Y2=0
r118 43 46 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=2.58 $Y=0 $X2=1.68
+ $Y2=0
r119 41 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r120 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r121 38 64 10.8012 $w=1.7e-07 $l=2.32e-07 $layer=LI1_cond $X=0.945 $Y=0
+ $X2=1.177 $Y2=0
r122 38 40 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.945 $Y=0
+ $X2=0.72 $Y2=0
r123 36 52 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=0
+ $X2=3.12 $Y2=0
r124 36 68 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=0
+ $X2=2.64 $Y2=0
r125 32 76 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=5.48 $Y=0.085
+ $X2=5.537 $Y2=0
r126 32 34 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=5.48 $Y=0.085
+ $X2=5.48 $Y2=0.625
r127 28 73 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.53 $Y=0.085
+ $X2=4.53 $Y2=0
r128 28 30 23.5098 $w=2.48e-07 $l=5.1e-07 $layer=LI1_cond $X=4.53 $Y=0.085
+ $X2=4.53 $Y2=0.595
r129 24 70 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=3.68 $Y=0.085
+ $X2=3.68 $Y2=0
r130 24 26 14.575 $w=3.38e-07 $l=4.3e-07 $layer=LI1_cond $X=3.68 $Y=0.085
+ $X2=3.68 $Y2=0.515
r131 20 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.745 $Y=0.085
+ $X2=2.745 $Y2=0
r132 20 22 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=2.745 $Y=0.085
+ $X2=2.745 $Y2=0.535
r133 16 64 1.88438 $w=4.65e-07 $l=8.5e-08 $layer=LI1_cond $X=1.177 $Y=0.085
+ $X2=1.177 $Y2=0
r134 16 18 10.0316 $w=4.63e-07 $l=3.9e-07 $layer=LI1_cond $X=1.177 $Y=0.085
+ $X2=1.177 $Y2=0.475
r135 5 34 182 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=1 $X=5.34
+ $Y=0.37 $X2=5.48 $Y2=0.625
r136 4 30 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=4.43
+ $Y=0.37 $X2=4.57 $Y2=0.595
r137 3 26 182 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_NDIFF $count=1 $X=3.465
+ $Y=0.37 $X2=3.68 $Y2=0.515
r138 2 22 182 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_NDIFF $count=1 $X=2.535
+ $Y=0.37 $X2=2.745 $Y2=0.535
r139 1 18 182 $w=1.7e-07 $l=6.79816e-07 $layer=licon1_NDIFF $count=1 $X=0.59
+ $Y=0.68 $X2=1.175 $Y2=0.475
.ends

