* File: sky130_fd_sc_ls__dlymetal6s6s_1.pxi.spice
* Created: Fri Aug 28 13:21:58 2020
* 
x_PM_SKY130_FD_SC_LS__DLYMETAL6S6S_1%A N_A_M1004_g N_A_c_88_n N_A_M1011_g A
+ N_A_c_89_n PM_SKY130_FD_SC_LS__DLYMETAL6S6S_1%A
x_PM_SKY130_FD_SC_LS__DLYMETAL6S6S_1%A_28_138# N_A_28_138#_M1004_s
+ N_A_28_138#_M1011_s N_A_28_138#_M1001_g N_A_28_138#_c_117_n
+ N_A_28_138#_M1009_g N_A_28_138#_c_118_n N_A_28_138#_c_132_n
+ N_A_28_138#_c_119_n N_A_28_138#_c_120_n N_A_28_138#_c_121_n
+ N_A_28_138#_c_124_n PM_SKY130_FD_SC_LS__DLYMETAL6S6S_1%A_28_138#
x_PM_SKY130_FD_SC_LS__DLYMETAL6S6S_1%A_209_74# N_A_209_74#_M1001_d
+ N_A_209_74#_M1009_d N_A_209_74#_M1006_g N_A_209_74#_c_179_n
+ N_A_209_74#_M1007_g N_A_209_74#_c_180_n N_A_209_74#_c_181_n
+ N_A_209_74#_c_182_n N_A_209_74#_c_187_n N_A_209_74#_c_183_n
+ N_A_209_74#_c_184_n N_A_209_74#_c_185_n N_A_209_74#_c_189_n
+ PM_SKY130_FD_SC_LS__DLYMETAL6S6S_1%A_209_74#
x_PM_SKY130_FD_SC_LS__DLYMETAL6S6S_1%A_316_138# N_A_316_138#_M1006_s
+ N_A_316_138#_M1007_s N_A_316_138#_M1010_g N_A_316_138#_c_244_n
+ N_A_316_138#_M1005_g N_A_316_138#_c_245_n N_A_316_138#_c_260_n
+ N_A_316_138#_c_246_n N_A_316_138#_c_247_n N_A_316_138#_c_248_n
+ N_A_316_138#_c_251_n PM_SKY130_FD_SC_LS__DLYMETAL6S6S_1%A_316_138#
x_PM_SKY130_FD_SC_LS__DLYMETAL6S6S_1%A_497_74# N_A_497_74#_M1010_d
+ N_A_497_74#_M1005_d N_A_497_74#_M1000_g N_A_497_74#_c_309_n
+ N_A_497_74#_M1008_g N_A_497_74#_c_310_n N_A_497_74#_c_317_n
+ N_A_497_74#_c_311_n N_A_497_74#_c_312_n N_A_497_74#_c_313_n
+ N_A_497_74#_c_314_n N_A_497_74#_c_318_n N_A_497_74#_c_315_n
+ PM_SKY130_FD_SC_LS__DLYMETAL6S6S_1%A_497_74#
x_PM_SKY130_FD_SC_LS__DLYMETAL6S6S_1%A_604_138# N_A_604_138#_M1000_s
+ N_A_604_138#_M1008_s N_A_604_138#_M1003_g N_A_604_138#_c_375_n
+ N_A_604_138#_M1002_g N_A_604_138#_c_387_n N_A_604_138#_c_376_n
+ N_A_604_138#_c_377_n N_A_604_138#_c_378_n N_A_604_138#_c_379_n
+ N_A_604_138#_c_382_n PM_SKY130_FD_SC_LS__DLYMETAL6S6S_1%A_604_138#
x_PM_SKY130_FD_SC_LS__DLYMETAL6S6S_1%VPWR N_VPWR_M1011_d N_VPWR_M1007_d
+ N_VPWR_M1008_d N_VPWR_c_435_n N_VPWR_c_436_n N_VPWR_c_437_n VPWR
+ N_VPWR_c_438_n N_VPWR_c_439_n N_VPWR_c_440_n N_VPWR_c_441_n N_VPWR_c_434_n
+ N_VPWR_c_443_n N_VPWR_c_444_n N_VPWR_c_445_n VPWR
+ PM_SKY130_FD_SC_LS__DLYMETAL6S6S_1%VPWR
x_PM_SKY130_FD_SC_LS__DLYMETAL6S6S_1%X N_X_M1003_d N_X_M1002_d N_X_c_485_n
+ N_X_c_488_n N_X_c_486_n X N_X_c_489_n N_X_c_487_n N_X_c_500_n N_X_c_491_n X
+ PM_SKY130_FD_SC_LS__DLYMETAL6S6S_1%X
x_PM_SKY130_FD_SC_LS__DLYMETAL6S6S_1%VGND N_VGND_M1004_d N_VGND_M1006_d
+ N_VGND_M1000_d N_VGND_c_536_n N_VGND_c_537_n N_VGND_c_538_n VGND
+ N_VGND_c_539_n N_VGND_c_540_n N_VGND_c_541_n N_VGND_c_542_n N_VGND_c_543_n
+ N_VGND_c_544_n N_VGND_c_545_n N_VGND_c_546_n VGND
+ PM_SKY130_FD_SC_LS__DLYMETAL6S6S_1%VGND
cc_1 VNB N_A_M1004_g 0.0286178f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=0.9
cc_2 VNB N_A_c_88_n 0.0428127f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.765
cc_3 VNB N_A_c_89_n 0.0129985f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.44
cc_4 VNB N_A_28_138#_M1001_g 0.0217641f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_5 VNB N_A_28_138#_c_117_n 0.0386283f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.44
cc_6 VNB N_A_28_138#_c_118_n 0.00533825f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_28_138#_c_119_n 0.00430876f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_28_138#_c_120_n 7.0366e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_28_138#_c_121_n 0.0201928f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_209_74#_M1006_g 0.0235592f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_209_74#_c_179_n 0.0423514f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.44
cc_12 VNB N_A_209_74#_c_180_n 0.0137727f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_209_74#_c_181_n 0.00523129f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_209_74#_c_182_n 0.0159058f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_209_74#_c_183_n 0.0013966f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_209_74#_c_184_n 0.00140045f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_209_74#_c_185_n 0.00344243f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_316_138#_M1010_g 0.0218556f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_316_138#_c_244_n 0.0384024f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.44
cc_20 VNB N_A_316_138#_c_245_n 0.00420983f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_316_138#_c_246_n 0.00578839f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_316_138#_c_247_n 9.03105e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_316_138#_c_248_n 0.00632352f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_497_74#_M1000_g 0.0234006f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_497_74#_c_309_n 0.0460635f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.44
cc_26 VNB N_A_497_74#_c_310_n 0.0147539f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_497_74#_c_311_n 0.00530393f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_497_74#_c_312_n 0.0160421f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_497_74#_c_313_n 0.00190862f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_497_74#_c_314_n 0.00344243f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_497_74#_c_315_n 0.00141674f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_604_138#_M1003_g 0.0223301f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_604_138#_c_375_n 0.0373543f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.44
cc_34 VNB N_A_604_138#_c_376_n 0.0029852f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_604_138#_c_377_n 0.00174446f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_604_138#_c_378_n 0.00547088f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_604_138#_c_379_n 9.14932e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VPWR_c_434_n 0.203486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_X_c_485_n 0.0318665f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_X_c_486_n 0.00832176f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_X_c_487_n 0.0274141f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_536_n 0.0187976f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.44
cc_43 VNB N_VGND_c_537_n 0.0125165f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_538_n 0.012298f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_539_n 0.0197723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_540_n 0.0312845f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_541_n 0.031135f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_542_n 0.0302512f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_543_n 0.314614f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_544_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_545_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_546_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VPB N_A_c_88_n 0.0336069f $X=-0.19 $Y=1.66 $X2=0.49 $Y2=1.765
cc_54 VPB N_A_c_89_n 0.00694124f $X=-0.19 $Y=1.66 $X2=0.39 $Y2=1.44
cc_55 VPB N_A_28_138#_c_117_n 0.0258859f $X=-0.19 $Y=1.66 $X2=0.39 $Y2=1.44
cc_56 VPB N_A_28_138#_c_120_n 0.00286642f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_A_28_138#_c_124_n 0.0138694f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_A_209_74#_c_179_n 0.0266515f $X=-0.19 $Y=1.66 $X2=0.39 $Y2=1.44
cc_59 VPB N_A_209_74#_c_187_n 0.00584205f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_A_209_74#_c_183_n 0.0042813f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_A_209_74#_c_189_n 0.0304457f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_A_316_138#_c_244_n 0.0247954f $X=-0.19 $Y=1.66 $X2=0.39 $Y2=1.44
cc_63 VPB N_A_316_138#_c_247_n 0.00320398f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_A_316_138#_c_251_n 0.0046748f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_A_497_74#_c_309_n 0.0266947f $X=-0.19 $Y=1.66 $X2=0.39 $Y2=1.44
cc_66 VPB N_A_497_74#_c_317_n 0.030369f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_A_497_74#_c_318_n 0.00734963f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_A_497_74#_c_315_n 0.00434639f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_A_604_138#_c_375_n 0.0269217f $X=-0.19 $Y=1.66 $X2=0.39 $Y2=1.44
cc_70 VPB N_A_604_138#_c_379_n 0.00329589f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_A_604_138#_c_382_n 0.00367379f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_435_n 0.0363206f $X=-0.19 $Y=1.66 $X2=0.39 $Y2=1.44
cc_73 VPB N_VPWR_c_436_n 0.0333726f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_437_n 0.0332872f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_438_n 0.0209183f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_439_n 0.035531f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_440_n 0.0349883f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_441_n 0.0284846f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_434_n 0.149501f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_443_n 0.00564836f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_444_n 0.00564836f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_445_n 0.00564503f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 VPB N_X_c_488_n 0.0368547f $X=-0.19 $Y=1.66 $X2=0.33 $Y2=1.44
cc_84 VPB N_X_c_489_n 0.0166148f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_X_c_487_n 0.00798828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_X_c_491_n 0.0730085f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 N_A_M1004_g N_A_28_138#_M1001_g 0.0165166f $X=0.48 $Y=0.9 $X2=0 $Y2=0
cc_88 N_A_M1004_g N_A_28_138#_c_117_n 7.45276e-19 $X=0.48 $Y=0.9 $X2=0 $Y2=0
cc_89 N_A_c_88_n N_A_28_138#_c_117_n 0.0406764f $X=0.49 $Y=1.765 $X2=0 $Y2=0
cc_90 N_A_c_89_n N_A_28_138#_c_117_n 2.61364e-19 $X=0.39 $Y=1.44 $X2=0 $Y2=0
cc_91 N_A_M1004_g N_A_28_138#_c_118_n 0.0142256f $X=0.48 $Y=0.9 $X2=0 $Y2=0
cc_92 N_A_c_88_n N_A_28_138#_c_118_n 0.00130174f $X=0.49 $Y=1.765 $X2=0 $Y2=0
cc_93 N_A_c_89_n N_A_28_138#_c_118_n 0.00983824f $X=0.39 $Y=1.44 $X2=0 $Y2=0
cc_94 N_A_c_88_n N_A_28_138#_c_132_n 0.0126821f $X=0.49 $Y=1.765 $X2=0 $Y2=0
cc_95 N_A_M1004_g N_A_28_138#_c_119_n 0.0027595f $X=0.48 $Y=0.9 $X2=0 $Y2=0
cc_96 N_A_c_88_n N_A_28_138#_c_119_n 0.00339828f $X=0.49 $Y=1.765 $X2=0 $Y2=0
cc_97 N_A_c_89_n N_A_28_138#_c_119_n 0.0202668f $X=0.39 $Y=1.44 $X2=0 $Y2=0
cc_98 N_A_c_88_n N_A_28_138#_c_120_n 0.0047408f $X=0.49 $Y=1.765 $X2=0 $Y2=0
cc_99 N_A_c_89_n N_A_28_138#_c_120_n 0.0122787f $X=0.39 $Y=1.44 $X2=0 $Y2=0
cc_100 N_A_M1004_g N_A_28_138#_c_121_n 0.00158922f $X=0.48 $Y=0.9 $X2=0 $Y2=0
cc_101 N_A_c_88_n N_A_28_138#_c_121_n 0.00417844f $X=0.49 $Y=1.765 $X2=0 $Y2=0
cc_102 N_A_c_89_n N_A_28_138#_c_121_n 0.0209233f $X=0.39 $Y=1.44 $X2=0 $Y2=0
cc_103 N_A_c_88_n N_A_28_138#_c_124_n 0.00342022f $X=0.49 $Y=1.765 $X2=0 $Y2=0
cc_104 N_A_c_89_n N_A_28_138#_c_124_n 0.0335534f $X=0.39 $Y=1.44 $X2=0 $Y2=0
cc_105 N_A_c_88_n N_A_209_74#_c_187_n 2.24143e-19 $X=0.49 $Y=1.765 $X2=0 $Y2=0
cc_106 N_A_c_88_n N_A_209_74#_c_189_n 7.0547e-19 $X=0.49 $Y=1.765 $X2=0 $Y2=0
cc_107 N_A_c_88_n N_VPWR_c_435_n 0.00229562f $X=0.49 $Y=1.765 $X2=0 $Y2=0
cc_108 N_A_M1004_g N_VGND_c_536_n 0.00429157f $X=0.48 $Y=0.9 $X2=0 $Y2=0
cc_109 N_A_M1004_g N_VGND_c_539_n 0.00382655f $X=0.48 $Y=0.9 $X2=0 $Y2=0
cc_110 N_A_M1004_g N_VGND_c_543_n 0.00451834f $X=0.48 $Y=0.9 $X2=0 $Y2=0
cc_111 N_A_28_138#_c_117_n N_A_209_74#_c_179_n 0.00507369f $X=1.005 $Y=1.765
+ $X2=0 $Y2=0
cc_112 N_A_28_138#_M1001_g N_A_209_74#_c_180_n 0.00268996f $X=0.97 $Y=0.74 $X2=0
+ $Y2=0
cc_113 N_A_28_138#_M1001_g N_A_209_74#_c_181_n 0.00332518f $X=0.97 $Y=0.74 $X2=0
+ $Y2=0
cc_114 N_A_28_138#_c_117_n N_A_209_74#_c_181_n 8.26384e-19 $X=1.005 $Y=1.765
+ $X2=0 $Y2=0
cc_115 N_A_28_138#_c_119_n N_A_209_74#_c_181_n 0.0122064f $X=0.81 $Y=1.605 $X2=0
+ $Y2=0
cc_116 N_A_28_138#_c_117_n N_A_209_74#_c_187_n 0.003773f $X=1.005 $Y=1.765 $X2=0
+ $Y2=0
cc_117 N_A_28_138#_c_120_n N_A_209_74#_c_187_n 0.00380646f $X=0.81 $Y=1.935
+ $X2=0 $Y2=0
cc_118 N_A_28_138#_c_117_n N_A_209_74#_c_183_n 0.00517269f $X=1.005 $Y=1.765
+ $X2=0 $Y2=0
cc_119 N_A_28_138#_c_120_n N_A_209_74#_c_183_n 0.0111914f $X=0.81 $Y=1.935 $X2=0
+ $Y2=0
cc_120 N_A_28_138#_c_117_n N_A_209_74#_c_184_n 0.00101945f $X=1.005 $Y=1.765
+ $X2=0 $Y2=0
cc_121 N_A_28_138#_c_117_n N_A_209_74#_c_185_n 0.00341845f $X=1.005 $Y=1.765
+ $X2=0 $Y2=0
cc_122 N_A_28_138#_c_119_n N_A_209_74#_c_185_n 0.0244957f $X=0.81 $Y=1.605 $X2=0
+ $Y2=0
cc_123 N_A_28_138#_c_117_n N_A_209_74#_c_189_n 0.0199377f $X=1.005 $Y=1.765
+ $X2=0 $Y2=0
cc_124 N_A_28_138#_c_132_n N_A_209_74#_c_189_n 0.00629937f $X=0.725 $Y=2.037
+ $X2=0 $Y2=0
cc_125 N_A_28_138#_c_119_n N_A_209_74#_c_189_n 0.00274452f $X=0.81 $Y=1.605
+ $X2=0 $Y2=0
cc_126 N_A_28_138#_c_120_n N_A_209_74#_c_189_n 4.40431e-19 $X=0.81 $Y=1.935
+ $X2=0 $Y2=0
cc_127 N_A_28_138#_c_124_n N_A_209_74#_c_189_n 0.00216674f $X=0.43 $Y=2.08 $X2=0
+ $Y2=0
cc_128 N_A_28_138#_c_117_n N_A_316_138#_c_251_n 6.18577e-19 $X=1.005 $Y=1.765
+ $X2=0 $Y2=0
cc_129 N_A_28_138#_c_132_n N_VPWR_M1011_d 0.00815077f $X=0.725 $Y=2.037
+ $X2=-0.19 $Y2=-0.245
cc_130 N_A_28_138#_c_120_n N_VPWR_M1011_d 0.00174917f $X=0.81 $Y=1.935 $X2=-0.19
+ $Y2=-0.245
cc_131 N_A_28_138#_c_117_n N_VPWR_c_435_n 0.00320844f $X=1.005 $Y=1.765 $X2=0
+ $Y2=0
cc_132 N_A_28_138#_c_132_n N_VPWR_c_435_n 0.0232529f $X=0.725 $Y=2.037 $X2=0
+ $Y2=0
cc_133 N_A_28_138#_c_117_n N_VPWR_c_439_n 0.00444353f $X=1.005 $Y=1.765 $X2=0
+ $Y2=0
cc_134 N_A_28_138#_c_117_n N_VPWR_c_434_n 0.00866222f $X=1.005 $Y=1.765 $X2=0
+ $Y2=0
cc_135 N_A_28_138#_c_117_n N_X_c_491_n 0.00653011f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_136 N_A_28_138#_c_118_n N_VGND_M1004_d 0.00119058f $X=0.725 $Y=1.06 $X2=-0.19
+ $Y2=-0.245
cc_137 N_A_28_138#_c_119_n N_VGND_M1004_d 0.00179209f $X=0.81 $Y=1.605 $X2=-0.19
+ $Y2=-0.245
cc_138 N_A_28_138#_M1001_g N_VGND_c_536_n 0.0132572f $X=0.97 $Y=0.74 $X2=0 $Y2=0
cc_139 N_A_28_138#_c_117_n N_VGND_c_536_n 3.45021e-19 $X=1.005 $Y=1.765 $X2=0
+ $Y2=0
cc_140 N_A_28_138#_c_118_n N_VGND_c_536_n 0.00915704f $X=0.725 $Y=1.06 $X2=0
+ $Y2=0
cc_141 N_A_28_138#_c_119_n N_VGND_c_536_n 0.0110081f $X=0.81 $Y=1.605 $X2=0
+ $Y2=0
cc_142 N_A_28_138#_c_121_n N_VGND_c_539_n 0.00444585f $X=0.265 $Y=0.865 $X2=0
+ $Y2=0
cc_143 N_A_28_138#_M1001_g N_VGND_c_540_n 0.00383152f $X=0.97 $Y=0.74 $X2=0
+ $Y2=0
cc_144 N_A_28_138#_M1001_g N_VGND_c_543_n 0.00762539f $X=0.97 $Y=0.74 $X2=0
+ $Y2=0
cc_145 N_A_28_138#_c_121_n N_VGND_c_543_n 0.00830526f $X=0.265 $Y=0.865 $X2=0
+ $Y2=0
cc_146 N_A_209_74#_M1006_g N_A_316_138#_M1010_g 0.0165204f $X=1.92 $Y=0.9 $X2=0
+ $Y2=0
cc_147 N_A_209_74#_M1006_g N_A_316_138#_c_244_n 5.933e-19 $X=1.92 $Y=0.9 $X2=0
+ $Y2=0
cc_148 N_A_209_74#_c_179_n N_A_316_138#_c_244_n 0.0429287f $X=1.975 $Y=1.765
+ $X2=0 $Y2=0
cc_149 N_A_209_74#_c_182_n N_A_316_138#_c_244_n 2.57095e-19 $X=1.83 $Y=1.44
+ $X2=0 $Y2=0
cc_150 N_A_209_74#_M1006_g N_A_316_138#_c_245_n 0.0140061f $X=1.92 $Y=0.9 $X2=0
+ $Y2=0
cc_151 N_A_209_74#_c_179_n N_A_316_138#_c_245_n 0.00323739f $X=1.975 $Y=1.765
+ $X2=0 $Y2=0
cc_152 N_A_209_74#_c_182_n N_A_316_138#_c_245_n 0.0113458f $X=1.83 $Y=1.44 $X2=0
+ $Y2=0
cc_153 N_A_209_74#_c_179_n N_A_316_138#_c_260_n 0.0126979f $X=1.975 $Y=1.765
+ $X2=0 $Y2=0
cc_154 N_A_209_74#_M1006_g N_A_316_138#_c_246_n 0.00276635f $X=1.92 $Y=0.9 $X2=0
+ $Y2=0
cc_155 N_A_209_74#_c_179_n N_A_316_138#_c_246_n 0.00302017f $X=1.975 $Y=1.765
+ $X2=0 $Y2=0
cc_156 N_A_209_74#_c_182_n N_A_316_138#_c_246_n 0.0244444f $X=1.83 $Y=1.44 $X2=0
+ $Y2=0
cc_157 N_A_209_74#_c_179_n N_A_316_138#_c_247_n 0.00670394f $X=1.975 $Y=1.765
+ $X2=0 $Y2=0
cc_158 N_A_209_74#_M1006_g N_A_316_138#_c_248_n 0.00158921f $X=1.92 $Y=0.9 $X2=0
+ $Y2=0
cc_159 N_A_209_74#_c_179_n N_A_316_138#_c_248_n 0.00407385f $X=1.975 $Y=1.765
+ $X2=0 $Y2=0
cc_160 N_A_209_74#_c_180_n N_A_316_138#_c_248_n 0.0359881f $X=1.185 $Y=0.57
+ $X2=0 $Y2=0
cc_161 N_A_209_74#_c_182_n N_A_316_138#_c_248_n 0.0233038f $X=1.83 $Y=1.44 $X2=0
+ $Y2=0
cc_162 N_A_209_74#_c_179_n N_A_316_138#_c_251_n 0.00464014f $X=1.975 $Y=1.765
+ $X2=0 $Y2=0
cc_163 N_A_209_74#_c_182_n N_A_316_138#_c_251_n 0.0214194f $X=1.83 $Y=1.44 $X2=0
+ $Y2=0
cc_164 N_A_209_74#_c_187_n N_A_316_138#_c_251_n 0.0265951f $X=1.222 $Y=1.992
+ $X2=0 $Y2=0
cc_165 N_A_209_74#_c_189_n N_A_316_138#_c_251_n 0.00174864f $X=1.23 $Y=2 $X2=0
+ $Y2=0
cc_166 N_A_209_74#_c_179_n N_A_497_74#_c_318_n 3.5276e-19 $X=1.975 $Y=1.765
+ $X2=0 $Y2=0
cc_167 N_A_209_74#_c_189_n N_VPWR_c_435_n 0.0308556f $X=1.23 $Y=2 $X2=0 $Y2=0
cc_168 N_A_209_74#_c_179_n N_VPWR_c_436_n 0.00186442f $X=1.975 $Y=1.765 $X2=0
+ $Y2=0
cc_169 N_A_209_74#_c_189_n N_VPWR_c_439_n 0.0223888f $X=1.23 $Y=2 $X2=0 $Y2=0
cc_170 N_A_209_74#_c_189_n N_VPWR_c_434_n 0.0121047f $X=1.23 $Y=2 $X2=0 $Y2=0
cc_171 N_A_209_74#_c_179_n N_X_c_491_n 0.00483253f $X=1.975 $Y=1.765 $X2=0 $Y2=0
cc_172 N_A_209_74#_c_189_n N_X_c_491_n 0.0681112f $X=1.23 $Y=2 $X2=0 $Y2=0
cc_173 N_A_209_74#_c_180_n N_VGND_c_536_n 0.0252885f $X=1.185 $Y=0.57 $X2=0
+ $Y2=0
cc_174 N_A_209_74#_M1006_g N_VGND_c_537_n 0.00261888f $X=1.92 $Y=0.9 $X2=0 $Y2=0
cc_175 N_A_209_74#_c_180_n N_VGND_c_537_n 0.0141693f $X=1.185 $Y=0.57 $X2=0
+ $Y2=0
cc_176 N_A_209_74#_M1006_g N_VGND_c_540_n 0.00382655f $X=1.92 $Y=0.9 $X2=0 $Y2=0
cc_177 N_A_209_74#_c_180_n N_VGND_c_540_n 0.0206458f $X=1.185 $Y=0.57 $X2=0
+ $Y2=0
cc_178 N_A_209_74#_M1006_g N_VGND_c_543_n 0.00451834f $X=1.92 $Y=0.9 $X2=0 $Y2=0
cc_179 N_A_209_74#_c_180_n N_VGND_c_543_n 0.0111968f $X=1.185 $Y=0.57 $X2=0
+ $Y2=0
cc_180 N_A_316_138#_c_244_n N_A_497_74#_c_309_n 0.00588998f $X=2.49 $Y=1.765
+ $X2=0 $Y2=0
cc_181 N_A_316_138#_c_246_n N_A_497_74#_c_309_n 2.02801e-19 $X=2.25 $Y=1.605
+ $X2=0 $Y2=0
cc_182 N_A_316_138#_M1010_g N_A_497_74#_c_310_n 0.00270228f $X=2.41 $Y=0.74
+ $X2=0 $Y2=0
cc_183 N_A_316_138#_c_244_n N_A_497_74#_c_317_n 0.00435535f $X=2.49 $Y=1.765
+ $X2=0 $Y2=0
cc_184 N_A_316_138#_M1010_g N_A_497_74#_c_311_n 0.00322309f $X=2.41 $Y=0.74
+ $X2=0 $Y2=0
cc_185 N_A_316_138#_c_244_n N_A_497_74#_c_311_n 6.2756e-19 $X=2.49 $Y=1.765
+ $X2=0 $Y2=0
cc_186 N_A_316_138#_c_246_n N_A_497_74#_c_311_n 0.0113527f $X=2.25 $Y=1.605
+ $X2=0 $Y2=0
cc_187 N_A_316_138#_c_244_n N_A_497_74#_c_313_n 0.00314148f $X=2.49 $Y=1.765
+ $X2=0 $Y2=0
cc_188 N_A_316_138#_c_244_n N_A_497_74#_c_314_n 0.00326086f $X=2.49 $Y=1.765
+ $X2=0 $Y2=0
cc_189 N_A_316_138#_c_246_n N_A_497_74#_c_314_n 0.0247198f $X=2.25 $Y=1.605
+ $X2=0 $Y2=0
cc_190 N_A_316_138#_c_244_n N_A_497_74#_c_318_n 0.0107864f $X=2.49 $Y=1.765
+ $X2=0 $Y2=0
cc_191 N_A_316_138#_c_260_n N_A_497_74#_c_318_n 0.024669f $X=2.165 $Y=2.017
+ $X2=0 $Y2=0
cc_192 N_A_316_138#_c_246_n N_A_497_74#_c_318_n 0.00484909f $X=2.25 $Y=1.605
+ $X2=0 $Y2=0
cc_193 N_A_316_138#_c_247_n N_A_497_74#_c_318_n 0.00443061f $X=2.25 $Y=1.895
+ $X2=0 $Y2=0
cc_194 N_A_316_138#_c_251_n N_A_497_74#_c_318_n 2.48727e-19 $X=1.87 $Y=2.06
+ $X2=0 $Y2=0
cc_195 N_A_316_138#_c_244_n N_A_497_74#_c_315_n 0.0052901f $X=2.49 $Y=1.765
+ $X2=0 $Y2=0
cc_196 N_A_316_138#_c_247_n N_A_497_74#_c_315_n 0.0102021f $X=2.25 $Y=1.895
+ $X2=0 $Y2=0
cc_197 N_A_316_138#_c_260_n N_VPWR_M1007_d 0.00769706f $X=2.165 $Y=2.017 $X2=0
+ $Y2=0
cc_198 N_A_316_138#_c_247_n N_VPWR_M1007_d 0.00133472f $X=2.25 $Y=1.895 $X2=0
+ $Y2=0
cc_199 N_A_316_138#_c_244_n N_VPWR_c_436_n 0.00352809f $X=2.49 $Y=1.765 $X2=0
+ $Y2=0
cc_200 N_A_316_138#_c_260_n N_VPWR_c_436_n 0.0185913f $X=2.165 $Y=2.017 $X2=0
+ $Y2=0
cc_201 N_A_316_138#_c_244_n N_VPWR_c_440_n 0.00461464f $X=2.49 $Y=1.765 $X2=0
+ $Y2=0
cc_202 N_A_316_138#_c_244_n N_VPWR_c_434_n 0.00917546f $X=2.49 $Y=1.765 $X2=0
+ $Y2=0
cc_203 N_A_316_138#_c_244_n N_X_c_491_n 0.00748895f $X=2.49 $Y=1.765 $X2=0 $Y2=0
cc_204 N_A_316_138#_c_260_n N_X_c_491_n 0.0116863f $X=2.165 $Y=2.017 $X2=0 $Y2=0
cc_205 N_A_316_138#_c_251_n N_X_c_491_n 0.0170914f $X=1.87 $Y=2.06 $X2=0 $Y2=0
cc_206 N_A_316_138#_c_245_n N_VGND_M1006_d 0.00119058f $X=2.165 $Y=1.06 $X2=0
+ $Y2=0
cc_207 N_A_316_138#_c_246_n N_VGND_M1006_d 0.00179209f $X=2.25 $Y=1.605 $X2=0
+ $Y2=0
cc_208 N_A_316_138#_M1010_g N_VGND_c_537_n 0.0132572f $X=2.41 $Y=0.74 $X2=0
+ $Y2=0
cc_209 N_A_316_138#_c_245_n N_VGND_c_537_n 0.00915704f $X=2.165 $Y=1.06 $X2=0
+ $Y2=0
cc_210 N_A_316_138#_c_246_n N_VGND_c_537_n 0.0110081f $X=2.25 $Y=1.605 $X2=0
+ $Y2=0
cc_211 N_A_316_138#_c_248_n N_VGND_c_540_n 0.00427375f $X=1.705 $Y=0.865 $X2=0
+ $Y2=0
cc_212 N_A_316_138#_M1010_g N_VGND_c_541_n 0.00383152f $X=2.41 $Y=0.74 $X2=0
+ $Y2=0
cc_213 N_A_316_138#_M1010_g N_VGND_c_543_n 0.00762539f $X=2.41 $Y=0.74 $X2=0
+ $Y2=0
cc_214 N_A_316_138#_c_248_n N_VGND_c_543_n 0.00802181f $X=1.705 $Y=0.865 $X2=0
+ $Y2=0
cc_215 N_A_497_74#_M1000_g N_A_604_138#_M1003_g 0.0165204f $X=3.36 $Y=0.9 $X2=0
+ $Y2=0
cc_216 N_A_497_74#_M1000_g N_A_604_138#_c_375_n 4.84716e-19 $X=3.36 $Y=0.9 $X2=0
+ $Y2=0
cc_217 N_A_497_74#_c_309_n N_A_604_138#_c_375_n 0.042757f $X=3.46 $Y=1.765 $X2=0
+ $Y2=0
cc_218 N_A_497_74#_c_312_n N_A_604_138#_c_375_n 2.23289e-19 $X=3.27 $Y=1.44
+ $X2=0 $Y2=0
cc_219 N_A_497_74#_c_310_n N_A_604_138#_c_387_n 0.0196927f $X=2.625 $Y=0.57
+ $X2=0 $Y2=0
cc_220 N_A_497_74#_M1000_g N_A_604_138#_c_376_n 0.0144149f $X=3.36 $Y=0.9 $X2=0
+ $Y2=0
cc_221 N_A_497_74#_c_309_n N_A_604_138#_c_376_n 0.00518557f $X=3.46 $Y=1.765
+ $X2=0 $Y2=0
cc_222 N_A_497_74#_c_312_n N_A_604_138#_c_376_n 0.0113081f $X=3.27 $Y=1.44 $X2=0
+ $Y2=0
cc_223 N_A_497_74#_c_309_n N_A_604_138#_c_377_n 0.0040983f $X=3.46 $Y=1.765
+ $X2=0 $Y2=0
cc_224 N_A_497_74#_c_312_n N_A_604_138#_c_377_n 0.0175411f $X=3.27 $Y=1.44 $X2=0
+ $Y2=0
cc_225 N_A_497_74#_c_313_n N_A_604_138#_c_377_n 0.013174f $X=2.697 $Y=1.075
+ $X2=0 $Y2=0
cc_226 N_A_497_74#_M1000_g N_A_604_138#_c_378_n 0.00277296f $X=3.36 $Y=0.9 $X2=0
+ $Y2=0
cc_227 N_A_497_74#_c_309_n N_A_604_138#_c_378_n 0.00335815f $X=3.46 $Y=1.765
+ $X2=0 $Y2=0
cc_228 N_A_497_74#_c_312_n N_A_604_138#_c_378_n 0.0246623f $X=3.27 $Y=1.44 $X2=0
+ $Y2=0
cc_229 N_A_497_74#_c_309_n N_A_604_138#_c_379_n 0.00733539f $X=3.46 $Y=1.765
+ $X2=0 $Y2=0
cc_230 N_A_497_74#_c_309_n N_A_604_138#_c_382_n 0.0211578f $X=3.46 $Y=1.765
+ $X2=0 $Y2=0
cc_231 N_A_497_74#_c_312_n N_A_604_138#_c_382_n 0.0171739f $X=3.27 $Y=1.44 $X2=0
+ $Y2=0
cc_232 N_A_497_74#_c_318_n N_A_604_138#_c_382_n 0.0250137f $X=2.715 $Y=2 $X2=0
+ $Y2=0
cc_233 N_A_497_74#_c_318_n N_VPWR_M1007_d 0.00207742f $X=2.715 $Y=2 $X2=0 $Y2=0
cc_234 N_A_497_74#_c_317_n N_VPWR_c_436_n 0.038177f $X=2.715 $Y=2.815 $X2=0
+ $Y2=0
cc_235 N_A_497_74#_c_309_n N_VPWR_c_437_n 0.00186878f $X=3.46 $Y=1.765 $X2=0
+ $Y2=0
cc_236 N_A_497_74#_c_317_n N_VPWR_c_440_n 0.0213627f $X=2.715 $Y=2.815 $X2=0
+ $Y2=0
cc_237 N_A_497_74#_c_317_n N_VPWR_c_434_n 0.0115856f $X=2.715 $Y=2.815 $X2=0
+ $Y2=0
cc_238 N_A_497_74#_c_309_n N_X_c_488_n 9.21606e-19 $X=3.46 $Y=1.765 $X2=0 $Y2=0
cc_239 N_A_497_74#_c_309_n N_X_c_489_n 3.56956e-19 $X=3.46 $Y=1.765 $X2=0 $Y2=0
cc_240 N_A_497_74#_c_309_n N_X_c_500_n 0.00261187f $X=3.46 $Y=1.765 $X2=0 $Y2=0
cc_241 N_A_497_74#_c_309_n N_X_c_491_n 0.00482652f $X=3.46 $Y=1.765 $X2=0 $Y2=0
cc_242 N_A_497_74#_c_317_n N_X_c_491_n 0.0369141f $X=2.715 $Y=2.815 $X2=0 $Y2=0
cc_243 N_A_497_74#_c_318_n N_X_c_491_n 0.03397f $X=2.715 $Y=2 $X2=0 $Y2=0
cc_244 N_A_497_74#_c_310_n N_VGND_c_537_n 0.0253911f $X=2.625 $Y=0.57 $X2=0
+ $Y2=0
cc_245 N_A_497_74#_M1000_g N_VGND_c_538_n 0.00254928f $X=3.36 $Y=0.9 $X2=0 $Y2=0
cc_246 N_A_497_74#_c_310_n N_VGND_c_538_n 0.0151085f $X=2.625 $Y=0.57 $X2=0
+ $Y2=0
cc_247 N_A_497_74#_M1000_g N_VGND_c_541_n 0.00382655f $X=3.36 $Y=0.9 $X2=0 $Y2=0
cc_248 N_A_497_74#_c_310_n N_VGND_c_541_n 0.0238717f $X=2.625 $Y=0.57 $X2=0
+ $Y2=0
cc_249 N_A_497_74#_M1000_g N_VGND_c_543_n 0.00451834f $X=3.36 $Y=0.9 $X2=0 $Y2=0
cc_250 N_A_497_74#_c_310_n N_VGND_c_543_n 0.0129463f $X=2.625 $Y=0.57 $X2=0
+ $Y2=0
cc_251 N_A_604_138#_c_379_n N_VPWR_M1008_d 0.00129487f $X=3.705 $Y=1.895 $X2=0
+ $Y2=0
cc_252 N_A_604_138#_c_382_n N_VPWR_M1008_d 0.00561191f $X=3.235 $Y=2.06 $X2=0
+ $Y2=0
cc_253 N_A_604_138#_c_375_n N_VPWR_c_437_n 0.00351639f $X=3.98 $Y=1.765 $X2=0
+ $Y2=0
cc_254 N_A_604_138#_c_382_n N_VPWR_c_437_n 0.0176897f $X=3.235 $Y=2.06 $X2=0
+ $Y2=0
cc_255 N_A_604_138#_c_375_n N_VPWR_c_441_n 0.00456575f $X=3.98 $Y=1.765 $X2=0
+ $Y2=0
cc_256 N_A_604_138#_c_375_n N_VPWR_c_434_n 0.00899198f $X=3.98 $Y=1.765 $X2=0
+ $Y2=0
cc_257 N_A_604_138#_M1003_g N_X_c_485_n 0.00271338f $X=3.85 $Y=0.74 $X2=0 $Y2=0
cc_258 N_A_604_138#_c_375_n N_X_c_488_n 0.0128767f $X=3.98 $Y=1.765 $X2=0 $Y2=0
cc_259 N_A_604_138#_c_382_n N_X_c_488_n 6.68901e-19 $X=3.235 $Y=2.06 $X2=0 $Y2=0
cc_260 N_A_604_138#_c_375_n N_X_c_486_n 0.00473153f $X=3.98 $Y=1.765 $X2=0 $Y2=0
cc_261 N_A_604_138#_c_378_n N_X_c_486_n 0.00241382f $X=3.705 $Y=1.605 $X2=0
+ $Y2=0
cc_262 N_A_604_138#_c_375_n X 0.00678614f $X=3.98 $Y=1.765 $X2=0 $Y2=0
cc_263 N_A_604_138#_c_375_n N_X_c_489_n 0.0097935f $X=3.98 $Y=1.765 $X2=0 $Y2=0
cc_264 N_A_604_138#_c_378_n N_X_c_489_n 0.00179568f $X=3.705 $Y=1.605 $X2=0
+ $Y2=0
cc_265 N_A_604_138#_c_379_n N_X_c_489_n 0.00449801f $X=3.705 $Y=1.895 $X2=0
+ $Y2=0
cc_266 N_A_604_138#_c_382_n N_X_c_489_n 0.017261f $X=3.235 $Y=2.06 $X2=0 $Y2=0
cc_267 N_A_604_138#_M1003_g N_X_c_487_n 0.00261251f $X=3.85 $Y=0.74 $X2=0 $Y2=0
cc_268 N_A_604_138#_c_375_n N_X_c_487_n 0.0127854f $X=3.98 $Y=1.765 $X2=0 $Y2=0
cc_269 N_A_604_138#_c_378_n N_X_c_487_n 0.0310126f $X=3.705 $Y=1.605 $X2=0 $Y2=0
cc_270 N_A_604_138#_c_379_n N_X_c_487_n 0.00788672f $X=3.705 $Y=1.895 $X2=0
+ $Y2=0
cc_271 N_A_604_138#_c_375_n N_X_c_500_n 0.0020164f $X=3.98 $Y=1.765 $X2=0 $Y2=0
cc_272 N_A_604_138#_c_378_n N_X_c_500_n 0.00573146f $X=3.705 $Y=1.605 $X2=0
+ $Y2=0
cc_273 N_A_604_138#_c_382_n N_X_c_500_n 0.0101289f $X=3.235 $Y=2.06 $X2=0 $Y2=0
cc_274 N_A_604_138#_c_382_n N_X_c_491_n 0.0271448f $X=3.235 $Y=2.06 $X2=0 $Y2=0
cc_275 N_A_604_138#_c_376_n N_VGND_M1000_d 0.00119058f $X=3.605 $Y=1.06 $X2=0
+ $Y2=0
cc_276 N_A_604_138#_c_378_n N_VGND_M1000_d 0.00179209f $X=3.705 $Y=1.605 $X2=0
+ $Y2=0
cc_277 N_A_604_138#_M1003_g N_VGND_c_538_n 0.0132572f $X=3.85 $Y=0.74 $X2=0
+ $Y2=0
cc_278 N_A_604_138#_c_376_n N_VGND_c_538_n 0.00915704f $X=3.605 $Y=1.06 $X2=0
+ $Y2=0
cc_279 N_A_604_138#_c_378_n N_VGND_c_538_n 0.0110542f $X=3.705 $Y=1.605 $X2=0
+ $Y2=0
cc_280 N_A_604_138#_c_387_n N_VGND_c_541_n 0.00310575f $X=3.145 $Y=0.865 $X2=0
+ $Y2=0
cc_281 N_A_604_138#_M1003_g N_VGND_c_542_n 0.00383152f $X=3.85 $Y=0.74 $X2=0
+ $Y2=0
cc_282 N_A_604_138#_M1003_g N_VGND_c_543_n 0.00762539f $X=3.85 $Y=0.74 $X2=0
+ $Y2=0
cc_283 N_A_604_138#_c_387_n N_VGND_c_543_n 0.00603761f $X=3.145 $Y=0.865 $X2=0
+ $Y2=0
cc_284 N_VPWR_c_437_n N_X_c_488_n 0.0353801f $X=3.75 $Y=2.475 $X2=0 $Y2=0
cc_285 N_VPWR_c_441_n N_X_c_488_n 0.0213486f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_286 N_VPWR_c_434_n N_X_c_488_n 0.0115672f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_287 N_VPWR_M1008_d X 9.9929e-19 $X=3.535 $Y=1.84 $X2=0 $Y2=0
cc_288 N_VPWR_c_437_n X 0.00438713f $X=3.75 $Y=2.475 $X2=0 $Y2=0
cc_289 N_VPWR_M1008_d N_X_c_500_n 0.00524614f $X=3.535 $Y=1.84 $X2=0 $Y2=0
cc_290 N_VPWR_c_437_n N_X_c_500_n 0.00133414f $X=3.75 $Y=2.475 $X2=0 $Y2=0
cc_291 N_VPWR_M1007_d N_X_c_491_n 8.55594e-19 $X=2.05 $Y=1.84 $X2=0 $Y2=0
cc_292 N_VPWR_c_435_n N_X_c_491_n 0.00566053f $X=0.78 $Y=2.475 $X2=0 $Y2=0
cc_293 N_VPWR_c_436_n N_X_c_491_n 0.0341338f $X=2.265 $Y=2.475 $X2=0 $Y2=0
cc_294 N_VPWR_c_437_n N_X_c_491_n 0.0288439f $X=3.75 $Y=2.475 $X2=0 $Y2=0
cc_295 N_X_c_485_n N_VGND_c_538_n 0.0254826f $X=4.065 $Y=0.57 $X2=0 $Y2=0
cc_296 N_X_c_485_n N_VGND_c_542_n 0.0270976f $X=4.065 $Y=0.57 $X2=0 $Y2=0
cc_297 N_X_c_485_n N_VGND_c_543_n 0.0146958f $X=4.065 $Y=0.57 $X2=0 $Y2=0
