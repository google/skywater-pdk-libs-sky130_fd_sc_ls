* File: sky130_fd_sc_ls__or3_1.spice
* Created: Fri Aug 28 13:58:13 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__or3_1.pex.spice"
.subckt sky130_fd_sc_ls__or3_1  VNB VPB C B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* C	C
* VPB	VPB
* VNB	VNB
MM1006 N_VGND_M1006_d N_C_M1006_g N_A_27_74#_M1006_s VNB NSHORT L=0.15 W=0.55
+ AD=0.09625 AS=0.15675 PD=0.9 PS=1.67 NRD=0 NRS=0 M=1 R=3.66667 SA=75000.2
+ SB=75002.1 A=0.0825 P=1.4 MULT=1
MM1002 N_A_27_74#_M1002_d N_B_M1002_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.55
+ AD=0.182875 AS=0.09625 PD=1.215 PS=0.9 NRD=0 NRS=15.264 M=1 R=3.66667
+ SA=75000.7 SB=75001.6 A=0.0825 P=1.4 MULT=1
MM1001 N_VGND_M1001_d N_A_M1001_g N_A_27_74#_M1002_d VNB NSHORT L=0.15 W=0.55
+ AD=0.11874 AS=0.182875 PD=0.989147 PS=1.215 NRD=15.264 NRS=0 M=1 R=3.66667
+ SA=75001.5 SB=75000.8 A=0.0825 P=1.4 MULT=1
MM1003 N_X_M1003_d N_A_27_74#_M1003_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.15976 PD=2.05 PS=1.33085 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75001.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1004 A_116_368# N_C_M1004_g N_A_27_74#_M1004_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.295 PD=1.27 PS=2.59 NRD=15.7403 NRS=1.9503 M=1 R=6.66667 SA=75000.2
+ SB=75002.1 A=0.15 P=2.3 MULT=1
MM1000 A_200_368# N_B_M1000_g A_116_368# VPB PHIGHVT L=0.15 W=1 AD=0.21 AS=0.135
+ PD=1.42 PS=1.27 NRD=30.5153 NRS=15.7403 M=1 R=6.66667 SA=75000.6 SB=75001.7
+ A=0.15 P=2.3 MULT=1
MM1007 N_VPWR_M1007_d N_A_M1007_g A_200_368# VPB PHIGHVT L=0.15 W=1 AD=0.35934
+ AS=0.21 PD=1.74528 PS=1.42 NRD=1.9503 NRS=30.5153 M=1 R=6.66667 SA=75001.2
+ SB=75001.1 A=0.15 P=2.3 MULT=1
MM1005 N_X_M1005_d N_A_27_74#_M1005_g N_VPWR_M1007_d VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.40246 PD=2.83 PS=1.95472 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.9 SB=75000.2 A=0.168 P=2.54 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.0636 P=10.24
*
.include "sky130_fd_sc_ls__or3_1.pxi.spice"
*
.ends
*
*
