* File: sky130_fd_sc_ls__a41o_2.pxi.spice
* Created: Wed Sep  2 10:53:32 2020
* 
x_PM_SKY130_FD_SC_LS__A41O_2%A4 N_A4_c_81_n N_A4_c_86_n N_A4_M1009_g N_A4_c_82_n
+ N_A4_M1005_g A4 N_A4_c_84_n PM_SKY130_FD_SC_LS__A41O_2%A4
x_PM_SKY130_FD_SC_LS__A41O_2%A3 N_A3_M1004_g N_A3_c_112_n N_A3_c_117_n
+ N_A3_M1008_g A3 A3 A3 N_A3_c_114_n N_A3_c_115_n PM_SKY130_FD_SC_LS__A41O_2%A3
x_PM_SKY130_FD_SC_LS__A41O_2%A2 N_A2_M1006_g N_A2_c_153_n N_A2_c_158_n
+ N_A2_M1013_g A2 A2 A2 N_A2_c_155_n N_A2_c_156_n PM_SKY130_FD_SC_LS__A41O_2%A2
x_PM_SKY130_FD_SC_LS__A41O_2%A1 N_A1_M1007_g N_A1_c_193_n N_A1_M1010_g A1
+ PM_SKY130_FD_SC_LS__A41O_2%A1
x_PM_SKY130_FD_SC_LS__A41O_2%B1 N_B1_M1002_g N_B1_c_229_n N_B1_M1000_g B1
+ N_B1_c_230_n PM_SKY130_FD_SC_LS__A41O_2%B1
x_PM_SKY130_FD_SC_LS__A41O_2%A_441_74# N_A_441_74#_M1007_d N_A_441_74#_M1000_d
+ N_A_441_74#_c_261_n N_A_441_74#_M1011_g N_A_441_74#_c_272_n
+ N_A_441_74#_M1001_g N_A_441_74#_c_262_n N_A_441_74#_M1012_g
+ N_A_441_74#_c_273_n N_A_441_74#_M1003_g N_A_441_74#_c_263_n
+ N_A_441_74#_c_264_n N_A_441_74#_c_265_n N_A_441_74#_c_266_n
+ N_A_441_74#_c_267_n N_A_441_74#_c_268_n N_A_441_74#_c_275_n
+ N_A_441_74#_c_269_n N_A_441_74#_c_276_n N_A_441_74#_c_270_n
+ N_A_441_74#_c_271_n PM_SKY130_FD_SC_LS__A41O_2%A_441_74#
x_PM_SKY130_FD_SC_LS__A41O_2%A_27_392# N_A_27_392#_M1009_s N_A_27_392#_M1008_d
+ N_A_27_392#_M1010_d N_A_27_392#_c_342_n N_A_27_392#_c_343_n
+ N_A_27_392#_c_344_n N_A_27_392#_c_345_n N_A_27_392#_c_346_n
+ N_A_27_392#_c_347_n N_A_27_392#_c_348_n N_A_27_392#_c_349_n
+ PM_SKY130_FD_SC_LS__A41O_2%A_27_392#
x_PM_SKY130_FD_SC_LS__A41O_2%VPWR N_VPWR_M1009_d N_VPWR_M1013_d N_VPWR_M1001_s
+ N_VPWR_M1003_s N_VPWR_c_403_n N_VPWR_c_404_n N_VPWR_c_405_n N_VPWR_c_406_n
+ N_VPWR_c_407_n N_VPWR_c_408_n VPWR N_VPWR_c_409_n N_VPWR_c_410_n
+ N_VPWR_c_411_n N_VPWR_c_412_n N_VPWR_c_413_n N_VPWR_c_414_n N_VPWR_c_402_n
+ PM_SKY130_FD_SC_LS__A41O_2%VPWR
x_PM_SKY130_FD_SC_LS__A41O_2%X N_X_M1011_d N_X_M1001_d N_X_c_462_n N_X_c_459_n
+ N_X_c_460_n N_X_c_472_n N_X_c_457_n X PM_SKY130_FD_SC_LS__A41O_2%X
x_PM_SKY130_FD_SC_LS__A41O_2%VGND N_VGND_M1005_s N_VGND_M1002_d N_VGND_M1012_s
+ N_VGND_c_493_n N_VGND_c_494_n N_VGND_c_495_n N_VGND_c_496_n N_VGND_c_497_n
+ VGND N_VGND_c_498_n N_VGND_c_499_n N_VGND_c_500_n
+ PM_SKY130_FD_SC_LS__A41O_2%VGND
cc_1 VNB N_A4_c_81_n 0.00976783f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.795
cc_2 VNB N_A4_c_82_n 0.0207173f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.22
cc_3 VNB A4 0.0082382f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_A4_c_84_n 0.058162f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.385
cc_5 VNB N_A3_c_112_n 0.00659705f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.46
cc_6 VNB A3 0.00532111f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_7 VNB N_A3_c_114_n 0.0306954f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.385
cc_8 VNB N_A3_c_115_n 0.0181058f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.295
cc_9 VNB N_A2_c_153_n 0.00678988f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.46
cc_10 VNB A2 0.0038768f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_11 VNB N_A2_c_155_n 0.0391048f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.385
cc_12 VNB N_A2_c_156_n 0.0200799f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.295
cc_13 VNB N_A1_M1007_g 0.0334159f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.885
cc_14 VNB N_A1_c_193_n 0.0205633f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.46
cc_15 VNB A1 0.00316184f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=0.74
cc_16 VNB N_B1_M1002_g 0.0325672f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.885
cc_17 VNB N_B1_c_229_n 0.018507f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.46
cc_18 VNB N_B1_c_230_n 0.00357093f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.385
cc_19 VNB N_A_441_74#_c_261_n 0.0187608f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=0.74
cc_20 VNB N_A_441_74#_c_262_n 0.0197849f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.385
cc_21 VNB N_A_441_74#_c_263_n 0.0165285f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_441_74#_c_264_n 0.0397326f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_441_74#_c_265_n 0.0722796f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_441_74#_c_266_n 0.0033626f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_441_74#_c_267_n 0.00990139f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_441_74#_c_268_n 0.0065138f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_441_74#_c_269_n 0.00557865f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_441_74#_c_270_n 0.00197732f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_441_74#_c_271_n 0.00285482f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VPWR_c_402_n 0.203486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_X_c_457_n 0.00545204f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB X 0.00329372f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.385
cc_33 VNB N_VGND_c_493_n 0.0131437f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_494_n 0.0344105f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.385
cc_35 VNB N_VGND_c_495_n 0.00985577f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.385
cc_36 VNB N_VGND_c_496_n 0.0655012f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_497_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_498_n 0.0217179f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_499_n 0.0492105f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_500_n 0.292499f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VPB N_A4_c_81_n 0.0101466f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.795
cc_42 VPB N_A4_c_86_n 0.0271866f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.885
cc_43 VPB N_A3_c_112_n 0.00724013f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.46
cc_44 VPB N_A3_c_117_n 0.0216084f $X=-0.19 $Y=1.66 $X2=0.53 $Y2=1.22
cc_45 VPB N_A2_c_153_n 0.00794645f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.46
cc_46 VPB N_A2_c_158_n 0.0235474f $X=-0.19 $Y=1.66 $X2=0.53 $Y2=1.22
cc_47 VPB N_A1_c_193_n 0.0389164f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.46
cc_48 VPB A1 0.00137218f $X=-0.19 $Y=1.66 $X2=0.53 $Y2=0.74
cc_49 VPB N_B1_c_229_n 0.0387086f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.46
cc_50 VPB N_B1_c_230_n 0.0024806f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.385
cc_51 VPB N_A_441_74#_c_272_n 0.0166815f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_A_441_74#_c_273_n 0.0174014f $X=-0.19 $Y=1.66 $X2=0.53 $Y2=1.385
cc_53 VPB N_A_441_74#_c_265_n 0.0174936f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_A_441_74#_c_275_n 0.0119461f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_A_441_74#_c_276_n 0.0120436f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_A_441_74#_c_270_n 0.00724087f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_A_27_392#_c_342_n 0.0443846f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.385
cc_58 VPB N_A_27_392#_c_343_n 0.0146284f $X=-0.19 $Y=1.66 $X2=0.53 $Y2=1.385
cc_59 VPB N_A_27_392#_c_344_n 0.00985309f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_A_27_392#_c_345_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_A_27_392#_c_346_n 0.0102508f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_A_27_392#_c_347_n 0.003977f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_A_27_392#_c_348_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_A_27_392#_c_349_n 0.00560004f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_403_n 0.00900305f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.385
cc_66 VPB N_VPWR_c_404_n 0.0186948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_405_n 0.0109589f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_406_n 0.0167107f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_407_n 0.0121909f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_408_n 0.0695592f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_409_n 0.0191515f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_410_n 0.0339528f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_411_n 0.0186948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_412_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_413_n 0.00978383f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_414_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_402_n 0.076804f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_X_c_459_n 0.00431889f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.385
cc_79 VPB N_X_c_460_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.385
cc_80 VPB N_X_c_457_n 0.00149334f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 N_A4_c_81_n N_A3_c_112_n 0.00598197f $X=0.505 $Y=1.795 $X2=0 $Y2=0
cc_82 N_A4_c_86_n N_A3_c_117_n 0.0317507f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_83 N_A4_c_82_n A3 0.00462195f $X=0.53 $Y=1.22 $X2=0 $Y2=0
cc_84 A4 A3 0.0147682f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_85 A4 N_A3_c_114_n 9.67587e-19 $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_86 N_A4_c_84_n N_A3_c_114_n 0.033243f $X=0.53 $Y=1.385 $X2=0 $Y2=0
cc_87 N_A4_c_82_n N_A3_c_115_n 0.033243f $X=0.53 $Y=1.22 $X2=0 $Y2=0
cc_88 N_A4_c_86_n N_A_27_392#_c_342_n 0.0140577f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_89 N_A4_c_81_n N_A_27_392#_c_343_n 0.00843106f $X=0.505 $Y=1.795 $X2=0 $Y2=0
cc_90 N_A4_c_86_n N_A_27_392#_c_343_n 0.00874324f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_91 A4 N_A_27_392#_c_343_n 6.17992e-19 $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_92 N_A4_c_84_n N_A_27_392#_c_343_n 4.15062e-19 $X=0.53 $Y=1.385 $X2=0 $Y2=0
cc_93 N_A4_c_81_n N_A_27_392#_c_344_n 0.00213197f $X=0.505 $Y=1.795 $X2=0 $Y2=0
cc_94 N_A4_c_86_n N_A_27_392#_c_344_n 0.00244188f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_95 A4 N_A_27_392#_c_344_n 0.0271109f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_96 N_A4_c_84_n N_A_27_392#_c_344_n 0.00228736f $X=0.53 $Y=1.385 $X2=0 $Y2=0
cc_97 N_A4_c_86_n N_A_27_392#_c_349_n 7.15392e-19 $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_98 N_A4_c_86_n N_VPWR_c_403_n 0.00874363f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_99 N_A4_c_86_n N_VPWR_c_409_n 0.00445602f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_100 N_A4_c_86_n N_VPWR_c_402_n 0.00861319f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_101 N_A4_c_82_n N_VGND_c_494_n 0.0159948f $X=0.53 $Y=1.22 $X2=0 $Y2=0
cc_102 A4 N_VGND_c_494_n 0.0241219f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_103 N_A4_c_84_n N_VGND_c_494_n 0.00199156f $X=0.53 $Y=1.385 $X2=0 $Y2=0
cc_104 N_A4_c_82_n N_VGND_c_496_n 0.00383152f $X=0.53 $Y=1.22 $X2=0 $Y2=0
cc_105 N_A4_c_82_n N_VGND_c_500_n 0.0075725f $X=0.53 $Y=1.22 $X2=0 $Y2=0
cc_106 N_A3_c_112_n N_A2_c_153_n 0.00843212f $X=1.055 $Y=1.795 $X2=0 $Y2=0
cc_107 N_A3_c_117_n N_A2_c_158_n 0.0165665f $X=1.055 $Y=1.885 $X2=0 $Y2=0
cc_108 A3 A2 0.0892488f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_109 N_A3_c_114_n A2 2.90162e-19 $X=1.01 $Y=1.385 $X2=0 $Y2=0
cc_110 N_A3_c_115_n A2 5.869e-19 $X=1.01 $Y=1.22 $X2=0 $Y2=0
cc_111 N_A3_c_114_n N_A2_c_155_n 0.0174537f $X=1.01 $Y=1.385 $X2=0 $Y2=0
cc_112 A3 N_A2_c_156_n 0.00916629f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_113 N_A3_c_115_n N_A2_c_156_n 0.0245047f $X=1.01 $Y=1.22 $X2=0 $Y2=0
cc_114 N_A3_c_117_n N_A_27_392#_c_342_n 7.1037e-19 $X=1.055 $Y=1.885 $X2=0 $Y2=0
cc_115 N_A3_c_112_n N_A_27_392#_c_343_n 0.0043556f $X=1.055 $Y=1.795 $X2=0 $Y2=0
cc_116 N_A3_c_117_n N_A_27_392#_c_343_n 0.00906272f $X=1.055 $Y=1.885 $X2=0
+ $Y2=0
cc_117 A3 N_A_27_392#_c_343_n 0.0209363f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_118 N_A3_c_114_n N_A_27_392#_c_343_n 8.27684e-19 $X=1.01 $Y=1.385 $X2=0 $Y2=0
cc_119 N_A3_c_117_n N_A_27_392#_c_345_n 0.00862222f $X=1.055 $Y=1.885 $X2=0
+ $Y2=0
cc_120 N_A3_c_112_n N_A_27_392#_c_349_n 0.00168439f $X=1.055 $Y=1.795 $X2=0
+ $Y2=0
cc_121 N_A3_c_117_n N_A_27_392#_c_349_n 0.00673667f $X=1.055 $Y=1.885 $X2=0
+ $Y2=0
cc_122 A3 N_A_27_392#_c_349_n 0.0181535f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_123 N_A3_c_114_n N_A_27_392#_c_349_n 2.37442e-19 $X=1.01 $Y=1.385 $X2=0 $Y2=0
cc_124 N_A3_c_117_n N_VPWR_c_403_n 0.00735548f $X=1.055 $Y=1.885 $X2=0 $Y2=0
cc_125 N_A3_c_117_n N_VPWR_c_404_n 0.00445602f $X=1.055 $Y=1.885 $X2=0 $Y2=0
cc_126 N_A3_c_117_n N_VPWR_c_402_n 0.00857909f $X=1.055 $Y=1.885 $X2=0 $Y2=0
cc_127 A3 N_VGND_c_494_n 0.0237984f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_128 N_A3_c_115_n N_VGND_c_494_n 0.00251629f $X=1.01 $Y=1.22 $X2=0 $Y2=0
cc_129 A3 N_VGND_c_496_n 0.0137277f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_130 N_A3_c_115_n N_VGND_c_496_n 0.00304348f $X=1.01 $Y=1.22 $X2=0 $Y2=0
cc_131 A3 N_VGND_c_500_n 0.0155751f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_132 N_A3_c_115_n N_VGND_c_500_n 0.00371612f $X=1.01 $Y=1.22 $X2=0 $Y2=0
cc_133 A3 A_199_74# 0.0136602f $X=1.115 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_134 A2 N_A1_M1007_g 0.00887723f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_135 N_A2_c_155_n N_A1_M1007_g 0.0127399f $X=1.65 $Y=1.385 $X2=0 $Y2=0
cc_136 N_A2_c_156_n N_A1_M1007_g 0.0197473f $X=1.615 $Y=1.22 $X2=0 $Y2=0
cc_137 N_A2_c_153_n N_A1_c_193_n 0.0097294f $X=1.505 $Y=1.795 $X2=0 $Y2=0
cc_138 N_A2_c_158_n N_A1_c_193_n 0.0175596f $X=1.505 $Y=1.885 $X2=0 $Y2=0
cc_139 A2 N_A1_c_193_n 3.48291e-19 $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_140 N_A2_c_155_n N_A1_c_193_n 0.006184f $X=1.65 $Y=1.385 $X2=0 $Y2=0
cc_141 N_A2_c_153_n A1 0.0012121f $X=1.505 $Y=1.795 $X2=0 $Y2=0
cc_142 A2 A1 0.00633735f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_143 N_A2_c_155_n A1 3.61063e-19 $X=1.65 $Y=1.385 $X2=0 $Y2=0
cc_144 A2 N_A_441_74#_c_268_n 0.00778382f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_145 N_A2_c_158_n N_A_27_392#_c_345_n 0.0144365f $X=1.505 $Y=1.885 $X2=0 $Y2=0
cc_146 N_A2_c_158_n N_A_27_392#_c_346_n 0.0161514f $X=1.505 $Y=1.885 $X2=0 $Y2=0
cc_147 A2 N_A_27_392#_c_346_n 0.0133989f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_148 N_A2_c_155_n N_A_27_392#_c_346_n 0.00127627f $X=1.65 $Y=1.385 $X2=0 $Y2=0
cc_149 N_A2_c_153_n N_A_27_392#_c_349_n 0.00416441f $X=1.505 $Y=1.795 $X2=0
+ $Y2=0
cc_150 N_A2_c_158_n N_A_27_392#_c_349_n 0.00978774f $X=1.505 $Y=1.885 $X2=0
+ $Y2=0
cc_151 N_A2_c_158_n N_VPWR_c_404_n 0.00445602f $X=1.505 $Y=1.885 $X2=0 $Y2=0
cc_152 N_A2_c_158_n N_VPWR_c_405_n 0.00775243f $X=1.505 $Y=1.885 $X2=0 $Y2=0
cc_153 N_A2_c_158_n N_VPWR_c_402_n 0.00859061f $X=1.505 $Y=1.885 $X2=0 $Y2=0
cc_154 A2 N_VGND_c_496_n 0.0094108f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_155 N_A2_c_156_n N_VGND_c_496_n 0.00378161f $X=1.615 $Y=1.22 $X2=0 $Y2=0
cc_156 A2 N_VGND_c_500_n 0.0110426f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_157 N_A2_c_156_n N_VGND_c_500_n 0.00629143f $X=1.615 $Y=1.22 $X2=0 $Y2=0
cc_158 A2 A_313_74# 0.0135149f $X=1.595 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_159 N_A1_M1007_g N_B1_M1002_g 0.0231835f $X=2.13 $Y=0.74 $X2=0 $Y2=0
cc_160 N_A1_c_193_n N_B1_c_229_n 0.0321211f $X=2.235 $Y=1.885 $X2=0 $Y2=0
cc_161 A1 N_B1_c_229_n 3.62235e-19 $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_162 N_A1_c_193_n N_B1_c_230_n 0.00201746f $X=2.235 $Y=1.885 $X2=0 $Y2=0
cc_163 A1 N_B1_c_230_n 0.0264884f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_164 N_A1_M1007_g N_A_441_74#_c_266_n 9.25648e-19 $X=2.13 $Y=0.74 $X2=0 $Y2=0
cc_165 N_A1_M1007_g N_A_441_74#_c_268_n 0.00253341f $X=2.13 $Y=0.74 $X2=0 $Y2=0
cc_166 N_A1_c_193_n N_A_441_74#_c_268_n 9.73364e-19 $X=2.235 $Y=1.885 $X2=0
+ $Y2=0
cc_167 A1 N_A_441_74#_c_268_n 0.0105084f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_168 N_A1_c_193_n N_A_27_392#_c_346_n 0.0143451f $X=2.235 $Y=1.885 $X2=0 $Y2=0
cc_169 A1 N_A_27_392#_c_346_n 0.0197776f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_170 N_A1_c_193_n N_A_27_392#_c_347_n 0.00120164f $X=2.235 $Y=1.885 $X2=0
+ $Y2=0
cc_171 A1 N_A_27_392#_c_347_n 0.00493222f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_172 N_A1_c_193_n N_A_27_392#_c_348_n 0.0144365f $X=2.235 $Y=1.885 $X2=0 $Y2=0
cc_173 N_A1_c_193_n N_A_27_392#_c_349_n 2.03256e-19 $X=2.235 $Y=1.885 $X2=0
+ $Y2=0
cc_174 A1 N_A_27_392#_c_349_n 0.00163617f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_175 N_A1_c_193_n N_VPWR_c_405_n 0.00928372f $X=2.235 $Y=1.885 $X2=0 $Y2=0
cc_176 N_A1_c_193_n N_VPWR_c_410_n 0.00445602f $X=2.235 $Y=1.885 $X2=0 $Y2=0
cc_177 N_A1_c_193_n N_VPWR_c_402_n 0.00859061f $X=2.235 $Y=1.885 $X2=0 $Y2=0
cc_178 N_A1_M1007_g N_VGND_c_496_n 0.00461464f $X=2.13 $Y=0.74 $X2=0 $Y2=0
cc_179 N_A1_M1007_g N_VGND_c_500_n 0.00912075f $X=2.13 $Y=0.74 $X2=0 $Y2=0
cc_180 N_B1_M1002_g N_A_441_74#_c_261_n 0.0260862f $X=2.67 $Y=0.74 $X2=0 $Y2=0
cc_181 N_B1_c_229_n N_A_441_74#_c_263_n 0.00525612f $X=2.685 $Y=1.885 $X2=0
+ $Y2=0
cc_182 N_B1_M1002_g N_A_441_74#_c_266_n 0.00451422f $X=2.67 $Y=0.74 $X2=0 $Y2=0
cc_183 N_B1_M1002_g N_A_441_74#_c_267_n 0.0160524f $X=2.67 $Y=0.74 $X2=0 $Y2=0
cc_184 N_B1_c_229_n N_A_441_74#_c_267_n 0.00411453f $X=2.685 $Y=1.885 $X2=0
+ $Y2=0
cc_185 N_B1_c_230_n N_A_441_74#_c_267_n 0.0269774f $X=2.76 $Y=1.615 $X2=0 $Y2=0
cc_186 N_B1_c_230_n N_A_441_74#_c_268_n 0.00309615f $X=2.76 $Y=1.615 $X2=0 $Y2=0
cc_187 N_B1_c_229_n N_A_441_74#_c_276_n 0.0232716f $X=2.685 $Y=1.885 $X2=0 $Y2=0
cc_188 N_B1_c_230_n N_A_441_74#_c_276_n 0.010879f $X=2.76 $Y=1.615 $X2=0 $Y2=0
cc_189 N_B1_c_229_n N_A_441_74#_c_270_n 0.00657778f $X=2.685 $Y=1.885 $X2=0
+ $Y2=0
cc_190 N_B1_c_230_n N_A_441_74#_c_270_n 0.0175146f $X=2.76 $Y=1.615 $X2=0 $Y2=0
cc_191 N_B1_M1002_g N_A_441_74#_c_271_n 0.00398645f $X=2.67 $Y=0.74 $X2=0 $Y2=0
cc_192 N_B1_c_229_n N_A_441_74#_c_271_n 3.86402e-19 $X=2.685 $Y=1.885 $X2=0
+ $Y2=0
cc_193 N_B1_c_230_n N_A_441_74#_c_271_n 0.00850124f $X=2.76 $Y=1.615 $X2=0 $Y2=0
cc_194 N_B1_c_229_n N_A_27_392#_c_347_n 0.00249431f $X=2.685 $Y=1.885 $X2=0
+ $Y2=0
cc_195 N_B1_c_230_n N_A_27_392#_c_347_n 0.0086545f $X=2.76 $Y=1.615 $X2=0 $Y2=0
cc_196 N_B1_c_229_n N_A_27_392#_c_348_n 0.00893311f $X=2.685 $Y=1.885 $X2=0
+ $Y2=0
cc_197 N_B1_c_229_n N_VPWR_c_406_n 0.00368752f $X=2.685 $Y=1.885 $X2=0 $Y2=0
cc_198 N_B1_c_229_n N_VPWR_c_410_n 0.00445602f $X=2.685 $Y=1.885 $X2=0 $Y2=0
cc_199 N_B1_c_229_n N_VPWR_c_402_n 0.00863237f $X=2.685 $Y=1.885 $X2=0 $Y2=0
cc_200 N_B1_M1002_g N_VGND_c_495_n 0.00693601f $X=2.67 $Y=0.74 $X2=0 $Y2=0
cc_201 N_B1_M1002_g N_VGND_c_496_n 0.00461464f $X=2.67 $Y=0.74 $X2=0 $Y2=0
cc_202 N_B1_M1002_g N_VGND_c_500_n 0.00910461f $X=2.67 $Y=0.74 $X2=0 $Y2=0
cc_203 N_A_441_74#_c_268_n N_A_27_392#_c_347_n 0.00610935f $X=2.56 $Y=1.195
+ $X2=0 $Y2=0
cc_204 N_A_441_74#_c_276_n N_A_27_392#_c_347_n 0.00755776f $X=2.96 $Y=2.115
+ $X2=0 $Y2=0
cc_205 N_A_441_74#_c_275_n N_A_27_392#_c_348_n 0.0330222f $X=2.96 $Y=2.815 $X2=0
+ $Y2=0
cc_206 N_A_441_74#_c_272_n N_VPWR_c_406_n 0.0172725f $X=3.795 $Y=1.765 $X2=0
+ $Y2=0
cc_207 N_A_441_74#_c_275_n N_VPWR_c_406_n 0.0478679f $X=2.96 $Y=2.815 $X2=0
+ $Y2=0
cc_208 N_A_441_74#_c_273_n N_VPWR_c_408_n 0.0261486f $X=4.245 $Y=1.765 $X2=0
+ $Y2=0
cc_209 N_A_441_74#_c_275_n N_VPWR_c_410_n 0.0146357f $X=2.96 $Y=2.815 $X2=0
+ $Y2=0
cc_210 N_A_441_74#_c_272_n N_VPWR_c_411_n 0.00445602f $X=3.795 $Y=1.765 $X2=0
+ $Y2=0
cc_211 N_A_441_74#_c_273_n N_VPWR_c_411_n 0.00445602f $X=4.245 $Y=1.765 $X2=0
+ $Y2=0
cc_212 N_A_441_74#_c_272_n N_VPWR_c_402_n 0.00861719f $X=3.795 $Y=1.765 $X2=0
+ $Y2=0
cc_213 N_A_441_74#_c_273_n N_VPWR_c_402_n 0.00860566f $X=4.245 $Y=1.765 $X2=0
+ $Y2=0
cc_214 N_A_441_74#_c_275_n N_VPWR_c_402_n 0.0121141f $X=2.96 $Y=2.815 $X2=0
+ $Y2=0
cc_215 N_A_441_74#_c_262_n N_X_c_462_n 0.0122008f $X=3.81 $Y=1.22 $X2=0 $Y2=0
cc_216 N_A_441_74#_c_265_n N_X_c_462_n 0.00376241f $X=3.81 $Y=1.492 $X2=0 $Y2=0
cc_217 N_A_441_74#_c_269_n N_X_c_462_n 0.0088769f $X=3.68 $Y=1.385 $X2=0 $Y2=0
cc_218 N_A_441_74#_c_272_n N_X_c_459_n 0.00427671f $X=3.795 $Y=1.765 $X2=0 $Y2=0
cc_219 N_A_441_74#_c_273_n N_X_c_459_n 0.00188635f $X=4.245 $Y=1.765 $X2=0 $Y2=0
cc_220 N_A_441_74#_c_265_n N_X_c_459_n 0.00241982f $X=3.81 $Y=1.492 $X2=0 $Y2=0
cc_221 N_A_441_74#_c_270_n N_X_c_459_n 0.00459661f $X=3.03 $Y=1.95 $X2=0 $Y2=0
cc_222 N_A_441_74#_c_272_n N_X_c_460_n 0.0171572f $X=3.795 $Y=1.765 $X2=0 $Y2=0
cc_223 N_A_441_74#_c_273_n N_X_c_460_n 0.0109216f $X=4.245 $Y=1.765 $X2=0 $Y2=0
cc_224 N_A_441_74#_c_276_n N_X_c_460_n 0.00459661f $X=2.96 $Y=2.115 $X2=0 $Y2=0
cc_225 N_A_441_74#_c_261_n N_X_c_472_n 0.00195381f $X=3.25 $Y=1.22 $X2=0 $Y2=0
cc_226 N_A_441_74#_c_264_n N_X_c_472_n 0.00136132f $X=3.705 $Y=1.385 $X2=0 $Y2=0
cc_227 N_A_441_74#_c_269_n N_X_c_472_n 0.0272424f $X=3.68 $Y=1.385 $X2=0 $Y2=0
cc_228 N_A_441_74#_c_272_n N_X_c_457_n 0.00116343f $X=3.795 $Y=1.765 $X2=0 $Y2=0
cc_229 N_A_441_74#_c_262_n N_X_c_457_n 0.00825937f $X=3.81 $Y=1.22 $X2=0 $Y2=0
cc_230 N_A_441_74#_c_273_n N_X_c_457_n 0.00251865f $X=4.245 $Y=1.765 $X2=0 $Y2=0
cc_231 N_A_441_74#_c_265_n N_X_c_457_n 0.0426768f $X=3.81 $Y=1.492 $X2=0 $Y2=0
cc_232 N_A_441_74#_c_269_n N_X_c_457_n 0.0337299f $X=3.68 $Y=1.385 $X2=0 $Y2=0
cc_233 N_A_441_74#_c_261_n X 0.0044265f $X=3.25 $Y=1.22 $X2=0 $Y2=0
cc_234 N_A_441_74#_c_271_n N_VGND_M1002_d 0.00279178f $X=3.18 $Y=1.33 $X2=0
+ $Y2=0
cc_235 N_A_441_74#_c_261_n N_VGND_c_495_n 0.00683054f $X=3.25 $Y=1.22 $X2=0
+ $Y2=0
cc_236 N_A_441_74#_c_266_n N_VGND_c_495_n 0.00127913f $X=2.395 $Y=0.515 $X2=0
+ $Y2=0
cc_237 N_A_441_74#_c_267_n N_VGND_c_495_n 0.0246062f $X=3.095 $Y=1.195 $X2=0
+ $Y2=0
cc_238 N_A_441_74#_c_271_n N_VGND_c_495_n 0.0021188f $X=3.18 $Y=1.33 $X2=0 $Y2=0
cc_239 N_A_441_74#_c_266_n N_VGND_c_496_n 0.0146357f $X=2.395 $Y=0.515 $X2=0
+ $Y2=0
cc_240 N_A_441_74#_c_261_n N_VGND_c_498_n 0.00461464f $X=3.25 $Y=1.22 $X2=0
+ $Y2=0
cc_241 N_A_441_74#_c_262_n N_VGND_c_498_n 0.00460063f $X=3.81 $Y=1.22 $X2=0
+ $Y2=0
cc_242 N_A_441_74#_c_261_n N_VGND_c_499_n 4.95096e-19 $X=3.25 $Y=1.22 $X2=0
+ $Y2=0
cc_243 N_A_441_74#_c_262_n N_VGND_c_499_n 0.00590656f $X=3.81 $Y=1.22 $X2=0
+ $Y2=0
cc_244 N_A_441_74#_c_265_n N_VGND_c_499_n 0.00517561f $X=3.81 $Y=1.492 $X2=0
+ $Y2=0
cc_245 N_A_441_74#_c_261_n N_VGND_c_500_n 0.00910813f $X=3.25 $Y=1.22 $X2=0
+ $Y2=0
cc_246 N_A_441_74#_c_262_n N_VGND_c_500_n 0.00442948f $X=3.81 $Y=1.22 $X2=0
+ $Y2=0
cc_247 N_A_441_74#_c_266_n N_VGND_c_500_n 0.0121141f $X=2.395 $Y=0.515 $X2=0
+ $Y2=0
cc_248 N_A_27_392#_c_346_n N_VPWR_M1013_d 0.00688982f $X=2.295 $Y=2.035 $X2=0
+ $Y2=0
cc_249 N_A_27_392#_c_342_n N_VPWR_c_403_n 0.0353111f $X=0.28 $Y=2.105 $X2=0
+ $Y2=0
cc_250 N_A_27_392#_c_343_n N_VPWR_c_403_n 0.0252372f $X=1.115 $Y=1.805 $X2=0
+ $Y2=0
cc_251 N_A_27_392#_c_349_n N_VPWR_c_403_n 0.0352735f $X=1.28 $Y=1.805 $X2=0
+ $Y2=0
cc_252 N_A_27_392#_c_345_n N_VPWR_c_404_n 0.014552f $X=1.28 $Y=2.815 $X2=0 $Y2=0
cc_253 N_A_27_392#_c_345_n N_VPWR_c_405_n 0.0267347f $X=1.28 $Y=2.815 $X2=0
+ $Y2=0
cc_254 N_A_27_392#_c_346_n N_VPWR_c_405_n 0.0379131f $X=2.295 $Y=2.035 $X2=0
+ $Y2=0
cc_255 N_A_27_392#_c_348_n N_VPWR_c_405_n 0.0267347f $X=2.46 $Y=2.815 $X2=0
+ $Y2=0
cc_256 N_A_27_392#_c_342_n N_VPWR_c_409_n 0.0145938f $X=0.28 $Y=2.105 $X2=0
+ $Y2=0
cc_257 N_A_27_392#_c_348_n N_VPWR_c_410_n 0.014552f $X=2.46 $Y=2.815 $X2=0 $Y2=0
cc_258 N_A_27_392#_c_342_n N_VPWR_c_402_n 0.0120466f $X=0.28 $Y=2.105 $X2=0
+ $Y2=0
cc_259 N_A_27_392#_c_345_n N_VPWR_c_402_n 0.0119791f $X=1.28 $Y=2.815 $X2=0
+ $Y2=0
cc_260 N_A_27_392#_c_348_n N_VPWR_c_402_n 0.0119791f $X=2.46 $Y=2.815 $X2=0
+ $Y2=0
cc_261 N_VPWR_c_408_n N_X_c_459_n 0.0450694f $X=4.52 $Y=1.985 $X2=0 $Y2=0
cc_262 N_VPWR_c_406_n N_X_c_460_n 0.0274314f $X=3.52 $Y=2.38 $X2=0 $Y2=0
cc_263 N_VPWR_c_411_n N_X_c_460_n 0.014552f $X=4.355 $Y=3.33 $X2=0 $Y2=0
cc_264 N_VPWR_c_402_n N_X_c_460_n 0.0119791f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_265 N_X_c_462_n N_VGND_M1012_s 0.0123021f $X=4.015 $Y=0.855 $X2=0 $Y2=0
cc_266 N_X_c_457_n N_VGND_M1012_s 0.00901369f $X=4.02 $Y=1.82 $X2=0 $Y2=0
cc_267 X N_VGND_c_495_n 0.0127255f $X=3.515 $Y=0.47 $X2=0 $Y2=0
cc_268 X N_VGND_c_498_n 0.0144853f $X=3.515 $Y=0.47 $X2=0 $Y2=0
cc_269 N_X_c_462_n N_VGND_c_499_n 0.0205938f $X=4.015 $Y=0.855 $X2=0 $Y2=0
cc_270 X N_VGND_c_499_n 0.0123663f $X=3.515 $Y=0.47 $X2=0 $Y2=0
cc_271 N_X_c_462_n N_VGND_c_500_n 0.00626145f $X=4.015 $Y=0.855 $X2=0 $Y2=0
cc_272 X N_VGND_c_500_n 0.0120561f $X=3.515 $Y=0.47 $X2=0 $Y2=0
