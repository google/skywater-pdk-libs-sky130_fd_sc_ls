* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
X0 a_309_390# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 VGND RESET_B a_1663_81# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 Q a_1921_409# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X3 a_30_78# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 VGND a_1271_74# a_1921_409# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X5 VPWR a_309_390# a_495_390# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 a_1525_212# a_1271_74# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 VGND a_309_390# a_495_390# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X8 VGND a_697_463# a_839_359# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X9 VPWR a_1921_409# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X10 a_30_78# a_495_390# a_697_463# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X11 a_309_390# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X12 a_839_359# a_309_390# a_1271_74# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 a_1271_74# a_495_390# a_1478_493# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X14 a_839_359# a_495_390# a_1271_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X15 a_30_78# a_309_390# a_697_463# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 VGND a_1921_409# Q VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X17 a_1478_493# a_1525_212# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X18 a_697_463# a_309_390# a_798_463# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X19 VPWR a_1271_74# a_1921_409# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X20 a_1663_81# a_1271_74# a_1525_212# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X21 a_697_463# a_495_390# a_823_138# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X22 VPWR D a_30_78# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X23 a_901_138# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X24 Q a_1921_409# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X25 a_1481_81# a_1525_212# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X26 a_117_78# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X27 VPWR RESET_B a_1525_212# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X28 VPWR a_697_463# a_839_359# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X29 a_30_78# D a_117_78# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X30 a_1271_74# a_309_390# a_1481_81# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X31 VPWR RESET_B a_697_463# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X32 a_798_463# a_839_359# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X33 a_823_138# a_839_359# a_901_138# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
