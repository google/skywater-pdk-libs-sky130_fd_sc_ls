* File: sky130_fd_sc_ls__sdfrbp_2.pex.spice
* Created: Wed Sep  2 11:27:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__SDFRBP_2%A_27_79# 1 2 9 11 13 14 17 20 23 27 30 34
+ 37 38
c83 30 0 1.3813e-19 $X=2.275 $Y=2.405
r84 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.44
+ $Y=1.995 $X2=2.44 $Y2=1.995
r85 32 34 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=2.44 $Y=2.32
+ $X2=2.44 $Y2=1.995
r86 31 38 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.445 $Y=2.405
+ $X2=0.28 $Y2=2.405
r87 30 32 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.275 $Y=2.405
+ $X2=2.44 $Y2=2.32
r88 30 31 119.39 $w=1.68e-07 $l=1.83e-06 $layer=LI1_cond $X=2.275 $Y=2.405
+ $X2=0.445 $Y2=2.405
r89 27 28 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.23
+ $Y=1.415 $X2=1.23 $Y2=1.415
r90 25 37 0.221902 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=0.365 $Y=1.415
+ $X2=0.24 $Y2=1.415
r91 25 27 30.208 $w=3.28e-07 $l=8.65e-07 $layer=LI1_cond $X=0.365 $Y=1.415
+ $X2=1.23 $Y2=1.415
r92 21 38 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.28 $Y=2.49 $X2=0.28
+ $Y2=2.405
r93 21 23 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=0.28 $Y=2.49 $X2=0.28
+ $Y2=2.65
r94 20 38 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=0.2 $Y=2.32
+ $X2=0.28 $Y2=2.405
r95 19 37 7.38875 $w=2.1e-07 $l=1.83916e-07 $layer=LI1_cond $X=0.2 $Y=1.58
+ $X2=0.24 $Y2=1.415
r96 19 20 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=0.2 $Y=1.58 $X2=0.2
+ $Y2=2.32
r97 15 37 7.38875 $w=2.1e-07 $l=1.65e-07 $layer=LI1_cond $X=0.24 $Y=1.25
+ $X2=0.24 $Y2=1.415
r98 15 17 29.733 $w=2.48e-07 $l=6.45e-07 $layer=LI1_cond $X=0.24 $Y=1.25
+ $X2=0.24 $Y2=0.605
r99 14 28 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=1.4 $Y=1.415
+ $X2=1.23 $Y2=1.415
r100 11 35 50.023 $w=3.78e-07 $l=3.06186e-07 $layer=POLY_cond $X=2.615 $Y=2.245
+ $X2=2.49 $Y2=1.995
r101 11 13 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.615 $Y=2.245
+ $X2=2.615 $Y2=2.64
r102 7 14 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=1.475 $Y=1.25
+ $X2=1.4 $Y2=1.415
r103 7 9 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=1.475 $Y=1.25
+ $X2=1.475 $Y2=0.605
r104 2 23 600 $w=1.7e-07 $l=3.95917e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.32 $X2=0.28 $Y2=2.65
r105 1 17 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.395 $X2=0.28 $Y2=0.605
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRBP_2%SCE 2 3 5 6 8 9 11 14 18 23 24 26 27 29 30
+ 31 36 46
r86 41 42 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.385
+ $Y=1.985 $X2=1.385 $Y2=1.985
r87 36 41 12.5952 $w=3.3e-07 $l=1.11041e-07 $layer=POLY_cond $X=1.37 $Y=1.985
+ $X2=1.46 $Y2=2.032
r88 36 38 116.283 $w=3.3e-07 $l=6.65e-07 $layer=POLY_cond $X=1.37 $Y=1.985
+ $X2=0.705 $Y2=1.985
r89 31 46 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.71 $Y=1.985
+ $X2=1.625 $Y2=1.985
r90 31 46 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=1.61 $Y=1.985
+ $X2=1.625 $Y2=1.985
r91 31 42 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=1.61 $Y=1.985
+ $X2=1.385 $Y2=1.985
r92 30 42 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=1.2 $Y=1.985
+ $X2=1.385 $Y2=1.985
r93 29 30 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=0.705 $Y=1.985
+ $X2=1.2 $Y2=1.985
r94 29 38 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.705
+ $Y=1.985 $X2=0.705 $Y2=1.985
r95 27 44 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.57 $Y=1.455
+ $X2=2.57 $Y2=1.29
r96 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.57
+ $Y=1.455 $X2=2.57 $Y2=1.455
r97 24 26 34.3517 $w=2.58e-07 $l=7.75e-07 $layer=LI1_cond $X=1.795 $Y=1.49
+ $X2=2.57 $Y2=1.49
r98 23 31 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.71 $Y=1.82
+ $X2=1.71 $Y2=1.985
r99 22 24 7.21222 $w=2.6e-07 $l=1.67183e-07 $layer=LI1_cond $X=1.71 $Y=1.62
+ $X2=1.795 $Y2=1.49
r100 22 23 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=1.71 $Y=1.62 $X2=1.71
+ $Y2=1.82
r101 21 38 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=0.595 $Y=1.985
+ $X2=0.705 $Y2=1.985
r102 16 18 43.5851 $w=1.5e-07 $l=8.5e-08 $layer=POLY_cond $X=0.41 $Y=0.965
+ $X2=0.495 $Y2=0.965
r103 14 44 351.245 $w=1.5e-07 $l=6.85e-07 $layer=POLY_cond $X=2.66 $Y=0.605
+ $X2=2.66 $Y2=1.29
r104 9 41 19.5823 $w=1.5e-07 $l=2.13e-07 $layer=POLY_cond $X=1.46 $Y=2.245
+ $X2=1.46 $Y2=2.032
r105 9 11 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.46 $Y=2.245
+ $X2=1.46 $Y2=2.64
r106 6 21 64.077 $w=2.08e-07 $l=2.79285e-07 $layer=POLY_cond $X=0.505 $Y=2.245
+ $X2=0.465 $Y2=1.985
r107 6 8 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.505 $Y=2.245
+ $X2=0.505 $Y2=2.64
r108 3 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.495 $Y=0.89
+ $X2=0.495 $Y2=0.965
r109 3 5 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.495 $Y=0.89
+ $X2=0.495 $Y2=0.605
r110 2 21 42.0626 $w=2.08e-07 $l=1.90526e-07 $layer=POLY_cond $X=0.41 $Y=1.82
+ $X2=0.465 $Y2=1.985
r111 1 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.41 $Y=1.04
+ $X2=0.41 $Y2=0.965
r112 1 2 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=0.41 $Y=1.04 $X2=0.41
+ $Y2=1.82
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRBP_2%D 3 5 6 8 9 12 13 14
r47 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.925 $Y=1.09
+ $X2=1.925 $Y2=1.255
r48 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.925 $Y=1.09
+ $X2=1.925 $Y2=0.925
r49 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.925
+ $Y=1.09 $X2=1.925 $Y2=1.09
r50 9 13 7.43022 $w=3.78e-07 $l=2.45e-07 $layer=LI1_cond $X=1.68 $Y=1 $X2=1.925
+ $Y2=1
r51 6 8 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.88 $Y=2.245
+ $X2=1.88 $Y2=2.64
r52 5 6 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.88 $Y=2.155 $X2=1.88
+ $Y2=2.245
r53 5 15 349.839 $w=1.8e-07 $l=9e-07 $layer=POLY_cond $X=1.88 $Y=2.155 $X2=1.88
+ $Y2=1.255
r54 3 14 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.865 $Y=0.605
+ $X2=1.865 $Y2=0.925
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRBP_2%SCD 1 3 6 10 11 12 16
c44 11 0 1.32376e-19 $X=3.12 $Y=1.665
c45 1 0 1.3813e-19 $X=3.035 $Y=2.245
r46 11 12 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.11 $Y=1.605
+ $X2=3.11 $Y2=2.035
r47 11 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.11
+ $Y=1.605 $X2=3.11 $Y2=1.605
r48 10 16 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.11 $Y=1.945
+ $X2=3.11 $Y2=1.605
r49 9 16 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.11 $Y=1.44
+ $X2=3.11 $Y2=1.605
r50 6 9 428.16 $w=1.5e-07 $l=8.35e-07 $layer=POLY_cond $X=3.05 $Y=0.605 $X2=3.05
+ $Y2=1.44
r51 1 10 55.1908 $w=2.62e-07 $l=3.3541e-07 $layer=POLY_cond $X=3.035 $Y=2.245
+ $X2=3.11 $Y2=1.945
r52 1 3 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.035 $Y=2.245
+ $X2=3.035 $Y2=2.64
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRBP_2%CLK 1 3 6 8
c41 6 0 6.36774e-20 $X=4.645 $Y=2.46
c42 1 0 9.8593e-20 $X=4.62 $Y=1.445
r43 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.02
+ $Y=1.385 $X2=4.02 $Y2=1.385
r44 8 12 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=4.07 $Y=1.295 $X2=4.07
+ $Y2=1.385
r45 4 14 20.933 $w=1.5e-07 $l=2.78e-07 $layer=POLY_cond $X=4.645 $Y=1.775
+ $X2=4.645 $Y2=1.497
r46 4 6 351.245 $w=1.5e-07 $l=6.85e-07 $layer=POLY_cond $X=4.645 $Y=1.775
+ $X2=4.645 $Y2=2.46
r47 1 14 3.69632 $w=3.26e-07 $l=2.5e-08 $layer=POLY_cond $X=4.62 $Y=1.497
+ $X2=4.645 $Y2=1.497
r48 1 11 88.7117 $w=3.26e-07 $l=6e-07 $layer=POLY_cond $X=4.62 $Y=1.497 $X2=4.02
+ $Y2=1.497
r49 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.62 $Y=1.445 $X2=4.62
+ $Y2=0.965
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRBP_2%A_1025_119# 1 2 8 9 11 12 16 18 20 21 22 23
+ 25 29 30 31 33 34 37 38 39 41 46 50 54 61 62 65 67 69
c194 69 0 1.10669e-19 $X=6.045 $Y=1.575
c195 62 0 3.21364e-19 $X=9.475 $Y=1.07
c196 34 0 1.50504e-19 $X=8.155 $Y=0.665
c197 16 0 6.36741e-20 $X=6.54 $Y=0.805
r198 65 67 5.06676 $w=4.43e-07 $l=1.65e-07 $layer=LI1_cond $X=9.532 $Y=2.03
+ $X2=9.532 $Y2=1.865
r199 65 66 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.615
+ $Y=2.03 $X2=9.615 $Y2=2.03
r200 62 75 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=9.475 $Y=1.07
+ $X2=9.475 $Y2=1.165
r201 61 62 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.475
+ $Y=1.07 $X2=9.475 $Y2=1.07
r202 58 61 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=9.185 $Y=1.07
+ $X2=9.475 $Y2=1.07
r203 54 56 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=7.085 $Y=0.395
+ $X2=7.085 $Y2=0.665
r204 53 72 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.045 $Y=1.665
+ $X2=6.045 $Y2=1.83
r205 53 69 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=6.045 $Y=1.665
+ $X2=6.045 $Y2=1.575
r206 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.045
+ $Y=1.665 $X2=6.045 $Y2=1.665
r207 50 52 12.6702 $w=4.67e-07 $l=4.85e-07 $layer=LI1_cond $X=5.56 $Y=1.87
+ $X2=6.045 $Y2=1.87
r208 49 50 6.26981 $w=4.67e-07 $l=3.86814e-07 $layer=LI1_cond $X=5.32 $Y=2.155
+ $X2=5.56 $Y2=1.87
r209 42 61 0.716491 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=9.475 $Y=1.235
+ $X2=9.475 $Y2=1.07
r210 42 67 22.0012 $w=3.28e-07 $l=6.3e-07 $layer=LI1_cond $X=9.475 $Y=1.235
+ $X2=9.475 $Y2=1.865
r211 41 58 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.185 $Y=0.905
+ $X2=9.185 $Y2=1.07
r212 40 41 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=9.185 $Y=0.425
+ $X2=9.185 $Y2=0.905
r213 38 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.1 $Y=0.34
+ $X2=9.185 $Y2=0.425
r214 38 39 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=9.1 $Y=0.34
+ $X2=8.325 $Y2=0.34
r215 36 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.24 $Y=0.425
+ $X2=8.325 $Y2=0.34
r216 36 37 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=8.24 $Y=0.425
+ $X2=8.24 $Y2=0.58
r217 35 56 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.17 $Y=0.665
+ $X2=7.085 $Y2=0.665
r218 34 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.155 $Y=0.665
+ $X2=8.24 $Y2=0.58
r219 34 35 64.262 $w=1.68e-07 $l=9.85e-07 $layer=LI1_cond $X=8.155 $Y=0.665
+ $X2=7.17 $Y2=0.665
r220 33 50 6.73017 $w=1.7e-07 $l=3.7e-07 $layer=LI1_cond $X=5.56 $Y=1.5 $X2=5.56
+ $Y2=1.87
r221 32 46 3.76007 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=5.56 $Y=1.275
+ $X2=5.56 $Y2=1.132
r222 32 33 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=5.56 $Y=1.275
+ $X2=5.56 $Y2=1.5
r223 30 54 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7 $Y=0.395
+ $X2=7.085 $Y2=0.395
r224 30 31 102.428 $w=1.68e-07 $l=1.57e-06 $layer=LI1_cond $X=7 $Y=0.395
+ $X2=5.43 $Y2=0.395
r225 27 46 11.9288 $w=2.83e-07 $l=2.95e-07 $layer=LI1_cond $X=5.265 $Y=1.132
+ $X2=5.56 $Y2=1.132
r226 27 29 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=5.265 $Y=0.99
+ $X2=5.265 $Y2=0.74
r227 26 31 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.265 $Y=0.48
+ $X2=5.43 $Y2=0.395
r228 26 29 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=5.265 $Y=0.48
+ $X2=5.265 $Y2=0.74
r229 23 66 51.8789 $w=3.07e-07 $l=2.87228e-07 $layer=POLY_cond $X=9.7 $Y=2.28
+ $X2=9.62 $Y2=2.03
r230 23 25 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=9.7 $Y=2.28 $X2=9.7
+ $Y2=2.565
r231 21 75 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.31 $Y=1.165
+ $X2=9.475 $Y2=1.165
r232 21 22 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=9.31 $Y=1.165
+ $X2=8.95 $Y2=1.165
r233 18 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.875 $Y=1.09
+ $X2=8.95 $Y2=1.165
r234 18 20 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=8.875 $Y=1.09
+ $X2=8.875 $Y2=0.695
r235 14 16 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=6.54 $Y=1.5
+ $X2=6.54 $Y2=0.805
r236 13 69 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.21 $Y=1.575
+ $X2=6.045 $Y2=1.575
r237 12 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.465 $Y=1.575
+ $X2=6.54 $Y2=1.5
r238 12 13 130.755 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=6.465 $Y=1.575
+ $X2=6.21 $Y2=1.575
r239 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.1 $Y=2.21 $X2=6.1
+ $Y2=2.495
r240 8 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.1 $Y=2.12 $X2=6.1
+ $Y2=2.21
r241 8 72 112.726 $w=1.8e-07 $l=2.9e-07 $layer=POLY_cond $X=6.1 $Y=2.12 $X2=6.1
+ $Y2=1.83
r242 2 49 600 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=5.17
+ $Y=1.96 $X2=5.32 $Y2=2.155
r243 1 29 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.125
+ $Y=0.595 $X2=5.265 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRBP_2%A_1370_290# 1 2 8 11 13 15 18 19 22 23 25
+ 33 34 36
c95 34 0 1.91015e-19 $X=8.845 $Y=0.842
c96 22 0 6.53341e-20 $X=7.21 $Y=1.005
c97 13 0 1.69775e-19 $X=6.94 $Y=2.21
c98 11 0 1.56765e-19 $X=6.93 $Y=0.805
r99 37 39 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=6.93 $Y=1.615 $X2=6.94
+ $Y2=1.615
r100 32 34 4.47019 $w=4.93e-07 $l=1.85e-07 $layer=LI1_cond $X=8.66 $Y=0.842
+ $X2=8.845 $Y2=0.842
r101 32 33 9.48656 $w=4.93e-07 $l=1.65e-07 $layer=LI1_cond $X=8.66 $Y=0.842
+ $X2=8.495 $Y2=0.842
r102 29 34 7.09362 $w=1.7e-07 $l=2.48e-07 $layer=LI1_cond $X=8.845 $Y=1.09
+ $X2=8.845 $Y2=0.842
r103 29 36 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=8.845 $Y=1.09
+ $X2=8.845 $Y2=1.745
r104 25 27 27.0228 $w=2.88e-07 $l=6.8e-07 $layer=LI1_cond $X=8.785 $Y=1.91
+ $X2=8.785 $Y2=2.59
r105 23 36 7.71909 $w=2.88e-07 $l=1.45e-07 $layer=LI1_cond $X=8.785 $Y=1.89
+ $X2=8.785 $Y2=1.745
r106 23 25 0.794788 $w=2.88e-07 $l=2e-08 $layer=LI1_cond $X=8.785 $Y=1.89
+ $X2=8.785 $Y2=1.91
r107 22 33 83.8342 $w=1.68e-07 $l=1.285e-06 $layer=LI1_cond $X=7.21 $Y=1.005
+ $X2=8.495 $Y2=1.005
r108 19 39 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.105 $Y=1.615
+ $X2=6.94 $Y2=1.615
r109 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.105
+ $Y=1.615 $X2=7.105 $Y2=1.615
r110 16 22 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=7.105 $Y=1.09
+ $X2=7.21 $Y2=1.005
r111 16 18 27.7273 $w=2.08e-07 $l=5.25e-07 $layer=LI1_cond $X=7.105 $Y=1.09
+ $X2=7.105 $Y2=1.615
r112 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.94 $Y=2.21
+ $X2=6.94 $Y2=2.495
r113 9 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.93 $Y=1.45
+ $X2=6.93 $Y2=1.615
r114 9 11 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=6.93 $Y=1.45
+ $X2=6.93 $Y2=0.805
r115 8 13 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.94 $Y=2.12 $X2=6.94
+ $Y2=2.21
r116 7 39 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.94 $Y=1.78
+ $X2=6.94 $Y2=1.615
r117 7 8 132.161 $w=1.8e-07 $l=3.4e-07 $layer=POLY_cond $X=6.94 $Y=1.78 $X2=6.94
+ $Y2=2.12
r118 2 27 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=8.575
+ $Y=1.735 $X2=8.725 $Y2=2.59
r119 2 25 400 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=1 $X=8.575
+ $Y=1.735 $X2=8.725 $Y2=1.91
r120 1 32 182 $w=1.7e-07 $l=5.00125e-07 $layer=licon1_NDIFF $count=1 $X=8.52
+ $Y=0.375 $X2=8.66 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRBP_2%RESET_B 4 5 7 8 9 13 14 15 16 18 20 23 26
+ 27 29 32 34 35 36 37 45 48 51 53 56 67
c203 67 0 1.25229e-19 $X=10.8 $Y=2.035
c204 48 0 1.32376e-19 $X=3.605 $Y=2.032
c205 8 0 1.66e-21 $X=7.245 $Y=0.18
c206 5 0 9.37604e-20 $X=3.605 $Y=2.245
r207 58 67 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.945
+ $Y=1.985 $X2=10.945 $Y2=1.985
r208 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.825
+ $Y=1.96 $X2=7.825 $Y2=1.96
r209 53 55 14.7051 $w=2.95e-07 $l=9e-08 $layer=POLY_cond $X=7.735 $Y=2.002
+ $X2=7.825 $Y2=2.002
r210 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.95
+ $Y=1.985 $X2=3.95 $Y2=1.985
r211 48 50 46.1917 $w=3.6e-07 $l=3.45e-07 $layer=POLY_cond $X=3.605 $Y=2.032
+ $X2=3.95 $Y2=2.032
r212 47 48 4.68611 $w=3.6e-07 $l=3.5e-08 $layer=POLY_cond $X=3.57 $Y=2.032
+ $X2=3.605 $Y2=2.032
r213 45 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=2.035
+ $X2=10.8 $Y2=2.035
r214 43 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=2.035
+ $X2=7.92 $Y2=2.035
r215 39 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=2.035
+ $X2=4.08 $Y2=2.035
r216 37 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.065 $Y=2.035
+ $X2=7.92 $Y2=2.035
r217 36 45 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=10.655 $Y=2.035
+ $X2=10.8 $Y2=2.035
r218 36 37 3.20544 $w=1.4e-07 $l=2.59e-06 $layer=MET1_cond $X=10.655 $Y=2.035
+ $X2=8.065 $Y2=2.035
r219 35 39 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.225 $Y=2.035
+ $X2=4.08 $Y2=2.035
r220 34 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.775 $Y=2.035
+ $X2=7.92 $Y2=2.035
r221 34 35 4.39356 $w=1.4e-07 $l=3.55e-06 $layer=MET1_cond $X=7.775 $Y=2.035
+ $X2=4.225 $Y2=2.035
r222 30 32 71.7872 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=10.715 $Y=1.55
+ $X2=10.855 $Y2=1.55
r223 27 58 60.4771 $w=2.87e-07 $l=3.23612e-07 $layer=POLY_cond $X=11.005 $Y=2.28
+ $X2=10.945 $Y2=1.985
r224 27 29 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=11.005 $Y=2.28
+ $X2=11.005 $Y2=2.565
r225 26 58 38.6443 $w=2.87e-07 $l=2.05122e-07 $layer=POLY_cond $X=10.855 $Y=1.82
+ $X2=10.945 $Y2=1.985
r226 25 32 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.855 $Y=1.625
+ $X2=10.855 $Y2=1.55
r227 25 26 99.9894 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=10.855 $Y=1.625
+ $X2=10.855 $Y2=1.82
r228 21 30 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.715 $Y=1.475
+ $X2=10.715 $Y2=1.55
r229 21 23 458.926 $w=1.5e-07 $l=8.95e-07 $layer=POLY_cond $X=10.715 $Y=1.475
+ $X2=10.715 $Y2=0.58
r230 20 53 18.5736 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.735 $Y=1.795
+ $X2=7.735 $Y2=2.002
r231 19 20 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=7.735 $Y=1.24
+ $X2=7.735 $Y2=1.795
r232 16 53 34.3119 $w=2.95e-07 $l=2.96277e-07 $layer=POLY_cond $X=7.525 $Y=2.21
+ $X2=7.735 $Y2=2.002
r233 16 18 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.525 $Y=2.21
+ $X2=7.525 $Y2=2.495
r234 14 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.66 $Y=1.165
+ $X2=7.735 $Y2=1.24
r235 14 15 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=7.66 $Y=1.165
+ $X2=7.395 $Y2=1.165
r236 11 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.32 $Y=1.09
+ $X2=7.395 $Y2=1.165
r237 11 13 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.32 $Y=1.09
+ $X2=7.32 $Y2=0.805
r238 10 13 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=7.32 $Y=0.255
+ $X2=7.32 $Y2=0.805
r239 8 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.245 $Y=0.18
+ $X2=7.32 $Y2=0.255
r240 8 9 1845.96 $w=1.5e-07 $l=3.6e-06 $layer=POLY_cond $X=7.245 $Y=0.18
+ $X2=3.645 $Y2=0.18
r241 5 48 23.3057 $w=1.5e-07 $l=2.13e-07 $layer=POLY_cond $X=3.605 $Y=2.245
+ $X2=3.605 $Y2=2.032
r242 5 7 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.605 $Y=2.245
+ $X2=3.605 $Y2=2.64
r243 2 47 23.3057 $w=1.5e-07 $l=2.12e-07 $layer=POLY_cond $X=3.57 $Y=1.82
+ $X2=3.57 $Y2=2.032
r244 2 4 623.011 $w=1.5e-07 $l=1.215e-06 $layer=POLY_cond $X=3.57 $Y=1.82
+ $X2=3.57 $Y2=0.605
r245 1 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.57 $Y=0.255
+ $X2=3.645 $Y2=0.18
r246 1 4 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=3.57 $Y=0.255
+ $X2=3.57 $Y2=0.605
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRBP_2%A_1223_119# 1 2 3 12 14 16 17 21 27 30 31
+ 33 36 37
c108 36 0 3.02968e-20 $X=6.78 $Y=2.425
c109 33 0 1.03439e-19 $X=8.425 $Y=1.41
c110 21 0 2.62023e-19 $X=6.66 $Y=2.61
r111 36 38 8.88342 $w=2.38e-07 $l=1.85e-07 $layer=LI1_cond $X=6.78 $Y=2.425
+ $X2=6.78 $Y2=2.61
r112 36 37 5.07737 $w=2.38e-07 $l=8.5e-08 $layer=LI1_cond $X=6.78 $Y=2.425
+ $X2=6.78 $Y2=2.34
r113 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.425
+ $Y=1.41 $X2=8.425 $Y2=1.41
r114 31 33 32.0123 $w=3.13e-07 $l=8.75e-07 $layer=LI1_cond $X=7.55 $Y=1.417
+ $X2=8.425 $Y2=1.417
r115 30 42 10.3482 $w=3.36e-07 $l=3.72552e-07 $layer=LI1_cond $X=7.465 $Y=2.32
+ $X2=7.75 $Y2=2.522
r116 29 31 7.64049 $w=3.15e-07 $l=1.95944e-07 $layer=LI1_cond $X=7.465 $Y=1.575
+ $X2=7.55 $Y2=1.417
r117 29 30 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=7.465 $Y=1.575
+ $X2=7.465 $Y2=2.32
r118 28 36 2.75731 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=6.9 $Y=2.425
+ $X2=6.78 $Y2=2.425
r119 27 30 6.05874 $w=3.36e-07 $l=1.41244e-07 $layer=LI1_cond $X=7.38 $Y=2.425
+ $X2=7.465 $Y2=2.32
r120 27 28 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=7.38 $Y=2.425
+ $X2=6.9 $Y2=2.425
r121 25 37 90.6845 $w=1.68e-07 $l=1.39e-06 $layer=LI1_cond $X=6.745 $Y=0.95
+ $X2=6.745 $Y2=2.34
r122 21 38 0.974673 $w=2.3e-07 $l=1.2e-07 $layer=LI1_cond $X=6.66 $Y=2.61
+ $X2=6.78 $Y2=2.61
r123 21 23 16.7856 $w=2.28e-07 $l=3.35e-07 $layer=LI1_cond $X=6.66 $Y=2.61
+ $X2=6.325 $Y2=2.61
r124 17 25 7.51767 $w=3e-07 $l=1.8775e-07 $layer=LI1_cond $X=6.66 $Y=0.8
+ $X2=6.745 $Y2=0.95
r125 17 19 12.8689 $w=2.98e-07 $l=3.35e-07 $layer=LI1_cond $X=6.66 $Y=0.8
+ $X2=6.325 $Y2=0.8
r126 14 34 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=8.5 $Y=1.66
+ $X2=8.425 $Y2=1.41
r127 14 16 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=8.5 $Y=1.66
+ $X2=8.5 $Y2=2.235
r128 10 34 38.5562 $w=2.99e-07 $l=1.74714e-07 $layer=POLY_cond $X=8.445 $Y=1.245
+ $X2=8.425 $Y2=1.41
r129 10 12 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=8.445 $Y=1.245
+ $X2=8.445 $Y2=0.695
r130 3 42 600 $w=1.7e-07 $l=3.00791e-07 $layer=licon1_PDIFF $count=1 $X=7.6
+ $Y=2.285 $X2=7.75 $Y2=2.52
r131 2 23 600 $w=1.7e-07 $l=3.62319e-07 $layer=licon1_PDIFF $count=1 $X=6.175
+ $Y=2.285 $X2=6.325 $Y2=2.58
r132 1 19 182 $w=1.7e-07 $l=2.95212e-07 $layer=licon1_NDIFF $count=1 $X=6.115
+ $Y=0.595 $X2=6.325 $Y2=0.8
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRBP_2%A_852_119# 1 2 7 9 12 15 17 18 19 20 21 22
+ 24 25 26 27 29 30 32 33 37 38 39 42 44 46 50 54 63
c170 63 0 5.1675e-20 $X=5.595 $Y=1.61
c171 54 0 2.0443e-19 $X=4.49 $Y=1.847
c172 39 0 1.30843e-19 $X=9.04 $Y=1.55
c173 38 0 1.34905e-19 $X=9.85 $Y=1.55
c174 17 0 1.55925e-19 $X=5.595 $Y=3.075
c175 12 0 1.11043e-19 $X=5.095 $Y=2.46
r176 62 63 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=5.58 $Y=1.61
+ $X2=5.595 $Y2=1.61
r177 58 60 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=5.05 $Y=1.61
+ $X2=5.095 $Y2=1.61
r178 57 62 76.939 $w=3.3e-07 $l=4.4e-07 $layer=POLY_cond $X=5.14 $Y=1.61
+ $X2=5.58 $Y2=1.61
r179 57 60 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=5.14 $Y=1.61
+ $X2=5.095 $Y2=1.61
r180 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.14
+ $Y=1.61 $X2=5.14 $Y2=1.61
r181 54 56 16.1179 $w=4.92e-07 $l=7.59309e-07 $layer=LI1_cond $X=4.49 $Y=1.847
+ $X2=5.14 $Y2=1.61
r182 53 54 1.73577 $w=4.92e-07 $l=7e-08 $layer=LI1_cond $X=4.42 $Y=1.847
+ $X2=4.49 $Y2=1.847
r183 48 50 2.36043 $w=4.13e-07 $l=8.5e-08 $layer=LI1_cond $X=4.405 $Y=0.802
+ $X2=4.49 $Y2=0.802
r184 46 54 7.05553 $w=1.7e-07 $l=4.02e-07 $layer=LI1_cond $X=4.49 $Y=1.445
+ $X2=4.49 $Y2=1.847
r185 45 50 6.00275 $w=1.7e-07 $l=2.08e-07 $layer=LI1_cond $X=4.49 $Y=1.01
+ $X2=4.49 $Y2=0.802
r186 45 46 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=4.49 $Y=1.01
+ $X2=4.49 $Y2=1.445
r187 40 42 458.926 $w=1.5e-07 $l=8.95e-07 $layer=POLY_cond $X=9.925 $Y=1.475
+ $X2=9.925 $Y2=0.58
r188 38 40 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.85 $Y=1.55
+ $X2=9.925 $Y2=1.475
r189 38 39 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=9.85 $Y=1.55
+ $X2=9.04 $Y2=1.55
r190 35 37 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=8.95 $Y=2.81
+ $X2=8.95 $Y2=2.235
r191 34 39 26.9307 $w=1.5e-07 $l=1.48324e-07 $layer=POLY_cond $X=8.95 $Y=1.66
+ $X2=9.04 $Y2=1.55
r192 34 37 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=8.95 $Y=1.66
+ $X2=8.95 $Y2=2.235
r193 32 35 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=8.95 $Y=2.9 $X2=8.95
+ $Y2=2.81
r194 32 33 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=8.95 $Y=2.9
+ $X2=8.95 $Y2=3.075
r195 31 44 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=6.64 $Y=3.15 $X2=6.55
+ $Y2=3.15
r196 30 33 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=8.86 $Y=3.15
+ $X2=8.95 $Y2=3.075
r197 30 31 1138.34 $w=1.5e-07 $l=2.22e-06 $layer=POLY_cond $X=8.86 $Y=3.15
+ $X2=6.64 $Y2=3.15
r198 27 29 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.55 $Y=2.78
+ $X2=6.55 $Y2=2.495
r199 26 44 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=6.55 $Y=3.075
+ $X2=6.55 $Y2=3.15
r200 25 27 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.55 $Y=2.87 $X2=6.55
+ $Y2=2.78
r201 25 26 79.6855 $w=1.8e-07 $l=2.05e-07 $layer=POLY_cond $X=6.55 $Y=2.87
+ $X2=6.55 $Y2=3.075
r202 22 24 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.04 $Y=1.09
+ $X2=6.04 $Y2=0.805
r203 20 44 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=6.46 $Y=3.15 $X2=6.55
+ $Y2=3.15
r204 20 21 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=6.46 $Y=3.15
+ $X2=5.67 $Y2=3.15
r205 18 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.965 $Y=1.165
+ $X2=6.04 $Y2=1.09
r206 18 19 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=5.965 $Y=1.165
+ $X2=5.67 $Y2=1.165
r207 17 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.595 $Y=3.075
+ $X2=5.67 $Y2=3.15
r208 16 63 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.595 $Y=1.775
+ $X2=5.595 $Y2=1.61
r209 16 17 666.596 $w=1.5e-07 $l=1.3e-06 $layer=POLY_cond $X=5.595 $Y=1.775
+ $X2=5.595 $Y2=3.075
r210 15 62 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.58 $Y=1.445
+ $X2=5.58 $Y2=1.61
r211 14 19 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=5.58 $Y=1.24
+ $X2=5.67 $Y2=1.165
r212 14 15 79.6855 $w=1.8e-07 $l=2.05e-07 $layer=POLY_cond $X=5.58 $Y=1.24
+ $X2=5.58 $Y2=1.445
r213 10 60 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.095 $Y=1.775
+ $X2=5.095 $Y2=1.61
r214 10 12 351.245 $w=1.5e-07 $l=6.85e-07 $layer=POLY_cond $X=5.095 $Y=1.775
+ $X2=5.095 $Y2=2.46
r215 7 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.05 $Y=1.445
+ $X2=5.05 $Y2=1.61
r216 7 9 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.05 $Y=1.445 $X2=5.05
+ $Y2=0.965
r217 2 53 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=4.275
+ $Y=1.96 $X2=4.42 $Y2=2.085
r218 1 48 182 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_NDIFF $count=1 $X=4.26
+ $Y=0.595 $X2=4.405 $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRBP_2%A_2006_373# 1 2 7 9 12 17 19 20 21 22 25 27
+ 28 30 31 37
c110 21 0 3.10546e-20 $X=11.065 $Y=2.405
c111 20 0 1.34905e-19 $X=10.545 $Y=1.565
c112 12 0 1.25229e-19 $X=10.285 $Y=0.58
r113 36 37 22.2151 $w=3.58e-07 $l=1.65e-07 $layer=POLY_cond $X=10.12 $Y=2.072
+ $X2=10.285 $Y2=2.072
r114 31 34 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=11.23 $Y=2.405
+ $X2=11.23 $Y2=2.565
r115 29 30 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=11.775 $Y=0.875
+ $X2=11.775 $Y2=1.48
r116 27 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.69 $Y=0.79
+ $X2=11.775 $Y2=0.875
r117 27 28 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=11.69 $Y=0.79
+ $X2=11.455 $Y2=0.79
r118 23 28 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=11.29 $Y=0.705
+ $X2=11.455 $Y2=0.79
r119 23 25 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=11.29 $Y=0.705
+ $X2=11.29 $Y2=0.58
r120 21 31 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.065 $Y=2.405
+ $X2=11.23 $Y2=2.405
r121 21 22 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=11.065 $Y=2.405
+ $X2=10.545 $Y2=2.405
r122 19 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.69 $Y=1.565
+ $X2=11.775 $Y2=1.48
r123 19 20 74.7005 $w=1.68e-07 $l=1.145e-06 $layer=LI1_cond $X=11.69 $Y=1.565
+ $X2=10.545 $Y2=1.565
r124 18 37 16.1564 $w=3.58e-07 $l=1.2e-07 $layer=POLY_cond $X=10.405 $Y=2.072
+ $X2=10.285 $Y2=2.072
r125 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.405
+ $Y=2.03 $X2=10.405 $Y2=2.03
r126 15 22 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=10.405 $Y=2.32
+ $X2=10.545 $Y2=2.405
r127 15 17 11.936 $w=2.78e-07 $l=2.9e-07 $layer=LI1_cond $X=10.405 $Y=2.32
+ $X2=10.405 $Y2=2.03
r128 14 20 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=10.405 $Y=1.65
+ $X2=10.545 $Y2=1.565
r129 14 17 15.6403 $w=2.78e-07 $l=3.8e-07 $layer=LI1_cond $X=10.405 $Y=1.65
+ $X2=10.405 $Y2=2.03
r130 10 37 23.1716 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=10.285 $Y=1.865
+ $X2=10.285 $Y2=2.072
r131 10 12 658.904 $w=1.5e-07 $l=1.285e-06 $layer=POLY_cond $X=10.285 $Y=1.865
+ $X2=10.285 $Y2=0.58
r132 7 36 23.1716 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=10.12 $Y=2.28
+ $X2=10.12 $Y2=2.072
r133 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=10.12 $Y=2.28
+ $X2=10.12 $Y2=2.565
r134 2 34 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=11.08
+ $Y=2.355 $X2=11.23 $Y2=2.565
r135 1 25 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=11.15
+ $Y=0.37 $X2=11.29 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRBP_2%A_1790_75# 1 2 9 11 12 13 15 16 18 20 23 25
+ 27 30 32 33 34 36 39 47 51 56 58 61 64
c151 58 0 1.03069e-19 $X=10.01 $Y=2.365
c152 56 0 1.57754e-19 $X=10.01 $Y=1.045
c153 13 0 3.10546e-20 $X=11.455 $Y=2.28
c154 12 0 7.64129e-20 $X=11.455 $Y=2.19
r155 61 62 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.355
+ $Y=1.175 $X2=11.355 $Y2=1.175
r156 59 64 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=10.095 $Y=1.177
+ $X2=10.01 $Y2=1.177
r157 59 61 54.7954 $w=2.63e-07 $l=1.26e-06 $layer=LI1_cond $X=10.095 $Y=1.177
+ $X2=11.355 $Y2=1.177
r158 57 64 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=10.01 $Y=1.31
+ $X2=10.01 $Y2=1.177
r159 57 58 68.8289 $w=1.68e-07 $l=1.055e-06 $layer=LI1_cond $X=10.01 $Y=1.31
+ $X2=10.01 $Y2=2.365
r160 56 64 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=10.01 $Y=1.045
+ $X2=10.01 $Y2=1.177
r161 55 56 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=10.01 $Y=0.735
+ $X2=10.01 $Y2=1.045
r162 51 55 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.925 $Y=0.57
+ $X2=10.01 $Y2=0.735
r163 51 53 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=9.925 $Y=0.57
+ $X2=9.655 $Y2=0.57
r164 47 58 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.925 $Y=2.53
+ $X2=10.01 $Y2=2.365
r165 47 49 19.382 $w=3.28e-07 $l=5.55e-07 $layer=LI1_cond $X=9.925 $Y=2.53
+ $X2=9.37 $Y2=2.53
r166 43 44 9.38961 $w=3.85e-07 $l=7.5e-08 $layer=POLY_cond $X=12.44 $Y=1.51
+ $X2=12.515 $Y2=1.51
r167 42 43 44.4442 $w=3.85e-07 $l=3.55e-07 $layer=POLY_cond $X=12.085 $Y=1.51
+ $X2=12.44 $Y2=1.51
r168 41 42 11.8935 $w=3.85e-07 $l=9.5e-08 $layer=POLY_cond $X=11.99 $Y=1.51
+ $X2=12.085 $Y2=1.51
r169 37 46 24.9301 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=12.99 $Y=1.255
+ $X2=12.99 $Y2=1.51
r170 37 39 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=12.99 $Y=1.255
+ $X2=12.99 $Y2=0.69
r171 34 36 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=12.945 $Y=1.885
+ $X2=12.945 $Y2=2.46
r172 33 34 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=12.945 $Y=1.795
+ $X2=12.945 $Y2=1.885
r173 32 46 5.63377 $w=3.85e-07 $l=4.5e-08 $layer=POLY_cond $X=12.945 $Y=1.51
+ $X2=12.99 $Y2=1.51
r174 32 44 53.8338 $w=3.85e-07 $l=4.3e-07 $layer=POLY_cond $X=12.945 $Y=1.51
+ $X2=12.515 $Y2=1.51
r175 32 33 81.629 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=12.945 $Y=1.585
+ $X2=12.945 $Y2=1.795
r176 28 44 24.9301 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=12.515 $Y=1.255
+ $X2=12.515 $Y2=1.51
r177 28 30 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=12.515 $Y=1.255
+ $X2=12.515 $Y2=0.74
r178 25 43 24.9301 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=12.44 $Y=1.765
+ $X2=12.44 $Y2=1.51
r179 25 27 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=12.44 $Y=1.765
+ $X2=12.44 $Y2=2.4
r180 21 42 24.9301 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=12.085 $Y=1.255
+ $X2=12.085 $Y2=1.51
r181 21 23 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=12.085 $Y=1.255
+ $X2=12.085 $Y2=0.74
r182 18 41 24.9301 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=11.99 $Y=1.765
+ $X2=11.99 $Y2=1.51
r183 18 20 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=11.99 $Y=1.765
+ $X2=11.99 $Y2=2.4
r184 17 62 36.297 $w=3.28e-07 $l=3.76776e-07 $layer=POLY_cond $X=11.545 $Y=1.422
+ $X2=11.272 $Y2=1.175
r185 16 41 12.2091 $w=3.85e-07 $l=1.2657e-07 $layer=POLY_cond $X=11.9 $Y=1.422
+ $X2=11.99 $Y2=1.51
r186 16 17 61.1493 $w=3.35e-07 $l=3.55e-07 $layer=POLY_cond $X=11.9 $Y=1.422
+ $X2=11.545 $Y2=1.422
r187 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=11.455 $Y=2.28
+ $X2=11.455 $Y2=2.565
r188 12 13 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=11.455 $Y=2.19
+ $X2=11.455 $Y2=2.28
r189 11 17 34.4294 $w=3.28e-07 $l=2.08192e-07 $layer=POLY_cond $X=11.455 $Y=1.59
+ $X2=11.545 $Y2=1.422
r190 11 12 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=11.455 $Y=1.59
+ $X2=11.455 $Y2=2.19
r191 7 62 38.5876 $w=3.28e-07 $l=2.67047e-07 $layer=POLY_cond $X=11.075 $Y=1.01
+ $X2=11.272 $Y2=1.175
r192 7 9 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=11.075 $Y=1.01
+ $X2=11.075 $Y2=0.58
r193 2 49 600 $w=1.7e-07 $l=9.51998e-07 $layer=licon1_PDIFF $count=1 $X=9.025
+ $Y=1.735 $X2=9.37 $Y2=2.53
r194 1 53 182 $w=1.7e-07 $l=7.96555e-07 $layer=licon1_NDIFF $count=1 $X=8.95
+ $Y=0.375 $X2=9.655 $Y2=0.57
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRBP_2%A_2604_392# 1 2 7 9 12 14 16 19 21 24 28 32
+ 38 41
r51 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=13.8
+ $Y=1.465 $X2=13.8 $Y2=1.465
r52 36 41 0.499868 $w=3.3e-07 $l=1.3e-07 $layer=LI1_cond $X=13.325 $Y=1.465
+ $X2=13.195 $Y2=1.465
r53 36 38 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=13.325 $Y=1.465
+ $X2=13.8 $Y2=1.465
r54 32 34 31.4706 $w=2.58e-07 $l=7.1e-07 $layer=LI1_cond $X=13.195 $Y=2.105
+ $X2=13.195 $Y2=2.815
r55 30 41 6.26932 $w=2.6e-07 $l=1.65e-07 $layer=LI1_cond $X=13.195 $Y=1.63
+ $X2=13.195 $Y2=1.465
r56 30 32 21.0542 $w=2.58e-07 $l=4.75e-07 $layer=LI1_cond $X=13.195 $Y=1.63
+ $X2=13.195 $Y2=2.105
r57 26 41 6.26932 $w=2.6e-07 $l=1.65e-07 $layer=LI1_cond $X=13.195 $Y=1.3
+ $X2=13.195 $Y2=1.465
r58 26 28 34.7949 $w=2.58e-07 $l=7.85e-07 $layer=LI1_cond $X=13.195 $Y=1.3
+ $X2=13.195 $Y2=0.515
r59 24 25 1.77641 $w=4.07e-07 $l=1.5e-08 $layer=POLY_cond $X=14.385 $Y=1.532
+ $X2=14.4 $Y2=1.532
r60 23 24 49.1474 $w=4.07e-07 $l=4.15e-07 $layer=POLY_cond $X=13.97 $Y=1.532
+ $X2=14.385 $Y2=1.532
r61 22 23 4.14496 $w=4.07e-07 $l=3.5e-08 $layer=POLY_cond $X=13.935 $Y=1.532
+ $X2=13.97 $Y2=1.532
r62 21 39 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=13.845 $Y=1.465
+ $X2=13.8 $Y2=1.465
r63 21 22 12.5251 $w=4.07e-07 $l=1.1887e-07 $layer=POLY_cond $X=13.845 $Y=1.465
+ $X2=13.935 $Y2=1.532
r64 17 25 26.2866 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=14.4 $Y=1.3
+ $X2=14.4 $Y2=1.532
r65 17 19 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=14.4 $Y=1.3 $X2=14.4
+ $Y2=0.74
r66 14 24 26.2866 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=14.385 $Y=1.765
+ $X2=14.385 $Y2=1.532
r67 14 16 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=14.385 $Y=1.765
+ $X2=14.385 $Y2=2.4
r68 10 23 26.2866 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=13.97 $Y=1.3
+ $X2=13.97 $Y2=1.532
r69 10 12 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=13.97 $Y=1.3
+ $X2=13.97 $Y2=0.74
r70 7 22 26.2866 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=13.935 $Y=1.765
+ $X2=13.935 $Y2=1.532
r71 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=13.935 $Y=1.765
+ $X2=13.935 $Y2=2.4
r72 2 34 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=13.02
+ $Y=1.96 $X2=13.17 $Y2=2.815
r73 2 32 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=13.02
+ $Y=1.96 $X2=13.17 $Y2=2.105
r74 1 28 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=13.065
+ $Y=0.37 $X2=13.205 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRBP_2%VPWR 1 2 3 4 5 6 7 8 9 10 33 37 41 45 49 53
+ 59 65 69 71 76 77 79 80 81 88 106 110 115 120 125 133 136 138 141 144 151 154
+ 157 161
r188 160 161 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.64 $Y=3.33
+ $X2=14.64 $Y2=3.33
r189 157 158 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=3.33
+ $X2=13.68 $Y2=3.33
r190 154 155 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r191 151 152 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r192 142 148 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=10.32 $Y2=3.33
r193 141 142 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r194 138 139 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r195 135 136 10.7086 $w=6.83e-07 $l=1.65e-07 $layer=LI1_cond $X=1.235 $Y=3.072
+ $X2=1.4 $Y2=3.072
r196 131 135 0.611135 $w=6.83e-07 $l=3.5e-08 $layer=LI1_cond $X=1.2 $Y=3.072
+ $X2=1.235 $Y2=3.072
r197 131 133 18.0422 $w=6.83e-07 $l=5.85e-07 $layer=LI1_cond $X=1.2 $Y=3.072
+ $X2=0.615 $Y2=3.072
r198 131 132 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r199 129 161 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.16 $Y=3.33
+ $X2=14.64 $Y2=3.33
r200 129 158 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.16 $Y=3.33
+ $X2=13.68 $Y2=3.33
r201 128 129 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.16 $Y=3.33
+ $X2=14.16 $Y2=3.33
r202 126 157 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.875 $Y=3.33
+ $X2=13.71 $Y2=3.33
r203 126 128 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=13.875 $Y=3.33
+ $X2=14.16 $Y2=3.33
r204 125 160 4.29523 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=14.495 $Y=3.33
+ $X2=14.687 $Y2=3.33
r205 125 128 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=14.495 $Y=3.33
+ $X2=14.16 $Y2=3.33
r206 124 158 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=3.33
+ $X2=13.68 $Y2=3.33
r207 124 155 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=3.33
+ $X2=12.72 $Y2=3.33
r208 123 124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=3.33
+ $X2=13.2 $Y2=3.33
r209 121 154 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=12.83 $Y=3.33
+ $X2=12.685 $Y2=3.33
r210 121 123 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=12.83 $Y=3.33
+ $X2=13.2 $Y2=3.33
r211 120 157 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.545 $Y=3.33
+ $X2=13.71 $Y2=3.33
r212 120 123 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=13.545 $Y=3.33
+ $X2=13.2 $Y2=3.33
r213 119 155 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=12.72 $Y2=3.33
r214 119 152 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=11.76 $Y2=3.33
r215 118 119 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r216 116 151 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.85 $Y=3.33
+ $X2=11.725 $Y2=3.33
r217 116 118 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=11.85 $Y=3.33
+ $X2=12.24 $Y2=3.33
r218 115 154 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=12.54 $Y=3.33
+ $X2=12.685 $Y2=3.33
r219 115 118 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=12.54 $Y=3.33
+ $X2=12.24 $Y2=3.33
r220 114 152 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=11.76 $Y2=3.33
r221 114 148 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=10.32 $Y2=3.33
r222 113 114 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r223 111 113 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=10.86 $Y=3.33
+ $X2=11.28 $Y2=3.33
r224 110 151 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.6 $Y=3.33
+ $X2=11.725 $Y2=3.33
r225 110 113 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=11.6 $Y=3.33
+ $X2=11.28 $Y2=3.33
r226 109 142 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r227 108 109 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r228 106 141 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.19 $Y=3.33
+ $X2=8.315 $Y2=3.33
r229 106 108 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=8.19 $Y=3.33
+ $X2=7.92 $Y2=3.33
r230 104 105 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r231 102 105 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=6.96 $Y2=3.33
r232 101 104 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=5.04 $Y=3.33
+ $X2=6.96 $Y2=3.33
r233 101 102 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r234 99 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r235 98 99 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r236 96 99 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r237 96 139 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r238 95 98 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.6 $Y=3.33 $X2=4.56
+ $Y2=3.33
r239 95 96 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r240 93 138 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.445 $Y=3.33
+ $X2=3.28 $Y2=3.33
r241 93 95 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=3.445 $Y=3.33
+ $X2=3.6 $Y2=3.33
r242 92 139 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=3.12 $Y2=3.33
r243 92 132 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r244 91 136 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1.68 $Y=3.33
+ $X2=1.4 $Y2=3.33
r245 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r246 88 138 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.115 $Y=3.33
+ $X2=3.28 $Y2=3.33
r247 88 91 93.6203 $w=1.68e-07 $l=1.435e-06 $layer=LI1_cond $X=3.115 $Y=3.33
+ $X2=1.68 $Y2=3.33
r248 86 132 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r249 85 133 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=0.615 $Y2=3.33
r250 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r251 81 109 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r252 81 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6.96 $Y2=3.33
r253 79 104 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=7.07 $Y=3.33
+ $X2=6.96 $Y2=3.33
r254 79 80 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.07 $Y=3.33
+ $X2=7.195 $Y2=3.33
r255 78 108 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=7.32 $Y=3.33
+ $X2=7.92 $Y2=3.33
r256 78 80 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.32 $Y=3.33
+ $X2=7.195 $Y2=3.33
r257 76 98 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=4.705 $Y=3.33
+ $X2=4.56 $Y2=3.33
r258 76 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.705 $Y=3.33
+ $X2=4.87 $Y2=3.33
r259 75 101 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=5.035 $Y=3.33
+ $X2=5.04 $Y2=3.33
r260 75 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.035 $Y=3.33
+ $X2=4.87 $Y2=3.33
r261 71 74 34.1617 $w=2.78e-07 $l=8.3e-07 $layer=LI1_cond $X=14.635 $Y=1.985
+ $X2=14.635 $Y2=2.815
r262 69 160 3.06482 $w=2.8e-07 $l=1.07912e-07 $layer=LI1_cond $X=14.635 $Y=3.245
+ $X2=14.687 $Y2=3.33
r263 69 74 17.6982 $w=2.78e-07 $l=4.3e-07 $layer=LI1_cond $X=14.635 $Y=3.245
+ $X2=14.635 $Y2=2.815
r264 65 68 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=13.71 $Y=1.985
+ $X2=13.71 $Y2=2.815
r265 63 157 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.71 $Y=3.245
+ $X2=13.71 $Y2=3.33
r266 63 68 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=13.71 $Y=3.245
+ $X2=13.71 $Y2=2.815
r267 59 62 29.0098 $w=2.88e-07 $l=7.3e-07 $layer=LI1_cond $X=12.685 $Y=2.085
+ $X2=12.685 $Y2=2.815
r268 57 154 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=12.685 $Y=3.245
+ $X2=12.685 $Y2=3.33
r269 57 62 17.0879 $w=2.88e-07 $l=4.3e-07 $layer=LI1_cond $X=12.685 $Y=3.245
+ $X2=12.685 $Y2=2.815
r270 53 56 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=11.725 $Y=1.985
+ $X2=11.725 $Y2=2.815
r271 51 151 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=11.725 $Y=3.245
+ $X2=11.725 $Y2=3.33
r272 51 56 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=11.725 $Y=3.245
+ $X2=11.725 $Y2=2.815
r273 50 141 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.44 $Y=3.33
+ $X2=8.315 $Y2=3.33
r274 49 111 8.26286 $w=1.7e-07 $l=2.98e-07 $layer=LI1_cond $X=10.562 $Y=3.33
+ $X2=10.86 $Y2=3.33
r275 49 148 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r276 49 144 10.1516 $w=5.93e-07 $l=5.05e-07 $layer=LI1_cond $X=10.562 $Y=3.33
+ $X2=10.562 $Y2=2.825
r277 49 50 119.064 $w=1.68e-07 $l=1.825e-06 $layer=LI1_cond $X=10.265 $Y=3.33
+ $X2=8.44 $Y2=3.33
r278 45 48 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=8.315 $Y=1.91
+ $X2=8.315 $Y2=2.59
r279 43 141 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.315 $Y=3.245
+ $X2=8.315 $Y2=3.33
r280 43 48 30.194 $w=2.48e-07 $l=6.55e-07 $layer=LI1_cond $X=8.315 $Y=3.245
+ $X2=8.315 $Y2=2.59
r281 39 80 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.195 $Y=3.245
+ $X2=7.195 $Y2=3.33
r282 39 41 18.4391 $w=2.48e-07 $l=4e-07 $layer=LI1_cond $X=7.195 $Y=3.245
+ $X2=7.195 $Y2=2.845
r283 35 77 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.87 $Y=3.245
+ $X2=4.87 $Y2=3.33
r284 35 37 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=4.87 $Y=3.245
+ $X2=4.87 $Y2=2.835
r285 31 138 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.28 $Y=3.245
+ $X2=3.28 $Y2=3.33
r286 31 33 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=3.28 $Y=3.245
+ $X2=3.28 $Y2=2.78
r287 10 74 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=14.46
+ $Y=1.84 $X2=14.61 $Y2=2.815
r288 10 71 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=14.46
+ $Y=1.84 $X2=14.61 $Y2=1.985
r289 9 68 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=13.565
+ $Y=1.84 $X2=13.71 $Y2=2.815
r290 9 65 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=13.565
+ $Y=1.84 $X2=13.71 $Y2=1.985
r291 8 62 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=12.515
+ $Y=1.84 $X2=12.665 $Y2=2.815
r292 8 59 400 $w=1.7e-07 $l=3.11087e-07 $layer=licon1_PDIFF $count=1 $X=12.515
+ $Y=1.84 $X2=12.665 $Y2=2.085
r293 7 56 600 $w=1.7e-07 $l=5.6542e-07 $layer=licon1_PDIFF $count=1 $X=11.53
+ $Y=2.355 $X2=11.765 $Y2=2.815
r294 7 53 300 $w=1.7e-07 $l=4.73128e-07 $layer=licon1_PDIFF $count=2 $X=11.53
+ $Y=2.355 $X2=11.765 $Y2=1.985
r295 6 144 600 $w=1.7e-07 $l=6.26458e-07 $layer=licon1_PDIFF $count=1 $X=10.195
+ $Y=2.355 $X2=10.56 $Y2=2.825
r296 5 48 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=8.15
+ $Y=1.735 $X2=8.275 $Y2=2.59
r297 5 45 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=8.15
+ $Y=1.735 $X2=8.275 $Y2=1.91
r298 4 41 600 $w=1.7e-07 $l=6.60908e-07 $layer=licon1_PDIFF $count=1 $X=7.015
+ $Y=2.285 $X2=7.235 $Y2=2.845
r299 3 37 600 $w=1.7e-07 $l=9.47035e-07 $layer=licon1_PDIFF $count=1 $X=4.72
+ $Y=1.96 $X2=4.87 $Y2=2.835
r300 2 33 600 $w=1.7e-07 $l=5.38331e-07 $layer=licon1_PDIFF $count=1 $X=3.11
+ $Y=2.32 $X2=3.28 $Y2=2.78
r301 1 135 300 $w=1.7e-07 $l=8.679e-07 $layer=licon1_PDIFF $count=2 $X=0.58
+ $Y=2.32 $X2=1.235 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRBP_2%A_388_79# 1 2 3 4 5 16 22 24 25 27 28 29 31
+ 32 37 40 41 43 44 46 49 50 52 56
c156 56 0 3.02968e-20 $X=5.847 $Y=2.495
c157 50 0 4.7366e-20 $X=4.645 $Y=2.5
c158 46 0 5.1675e-20 $X=6.405 $Y=2.155
r159 56 58 1.5641 $w=2.34e-07 $l=3e-08 $layer=LI1_cond $X=5.847 $Y=2.495
+ $X2=5.847 $Y2=2.525
r160 55 56 13.2949 $w=2.34e-07 $l=2.55e-07 $layer=LI1_cond $X=5.847 $Y=2.24
+ $X2=5.847 $Y2=2.495
r161 49 50 4.62121 $w=1.78e-07 $l=7.5e-08 $layer=LI1_cond $X=4.57 $Y=2.5
+ $X2=4.645 $Y2=2.5
r162 47 48 2.50513 $w=4.87e-07 $l=1e-07 $layer=LI1_cond $X=3.72 $Y=2.405
+ $X2=3.72 $Y2=2.505
r163 45 46 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=6.405 $Y=1.29
+ $X2=6.405 $Y2=2.155
r164 43 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.32 $Y=1.205
+ $X2=6.405 $Y2=1.29
r165 43 44 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=6.32 $Y=1.205
+ $X2=5.99 $Y2=1.205
r166 42 55 2.60974 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=5.985 $Y=2.24
+ $X2=5.847 $Y2=2.24
r167 41 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.32 $Y=2.24
+ $X2=6.405 $Y2=2.155
r168 41 42 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=6.32 $Y=2.24
+ $X2=5.985 $Y2=2.24
r169 40 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.905 $Y=1.12
+ $X2=5.99 $Y2=1.205
r170 39 52 0.716491 $w=1.7e-07 $l=1.18427e-07 $layer=LI1_cond $X=5.905 $Y=0.82
+ $X2=5.825 $Y2=0.735
r171 39 40 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=5.905 $Y=0.82
+ $X2=5.905 $Y2=1.12
r172 37 56 2.60974 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=5.71 $Y=2.495
+ $X2=5.847 $Y2=2.495
r173 37 50 69.4813 $w=1.68e-07 $l=1.065e-06 $layer=LI1_cond $X=5.71 $Y=2.495
+ $X2=4.645 $Y2=2.495
r174 36 48 6.9916 $w=1.7e-07 $l=2.75e-07 $layer=LI1_cond $X=3.995 $Y=2.505
+ $X2=3.72 $Y2=2.505
r175 36 49 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=3.995 $Y=2.505
+ $X2=4.57 $Y2=2.505
r176 32 48 2.75122 $w=4.87e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.805 $Y=2.59
+ $X2=3.72 $Y2=2.505
r177 32 34 1.92632 $w=3.8e-07 $l=6e-08 $layer=LI1_cond $X=3.805 $Y=2.59
+ $X2=3.805 $Y2=2.65
r178 31 47 7.62281 $w=4.87e-07 $l=2.28583e-07 $layer=LI1_cond $X=3.53 $Y=2.32
+ $X2=3.72 $Y2=2.405
r179 30 31 74.7005 $w=1.68e-07 $l=1.145e-06 $layer=LI1_cond $X=3.53 $Y=1.175
+ $X2=3.53 $Y2=2.32
r180 28 47 6.9916 $w=1.7e-07 $l=2.75e-07 $layer=LI1_cond $X=3.445 $Y=2.405
+ $X2=3.72 $Y2=2.405
r181 28 29 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=3.445 $Y=2.405
+ $X2=2.945 $Y2=2.405
r182 26 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.86 $Y=2.49
+ $X2=2.945 $Y2=2.405
r183 26 27 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.86 $Y=2.49
+ $X2=2.86 $Y2=2.66
r184 24 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.445 $Y=1.09
+ $X2=3.53 $Y2=1.175
r185 24 25 54.4759 $w=1.68e-07 $l=8.35e-07 $layer=LI1_cond $X=3.445 $Y=1.09
+ $X2=2.61 $Y2=1.09
r186 20 25 7.93686 $w=1.7e-07 $l=2.13307e-07 $layer=LI1_cond $X=2.435 $Y=1.005
+ $X2=2.61 $Y2=1.09
r187 20 22 10.7013 $w=3.48e-07 $l=3.25e-07 $layer=LI1_cond $X=2.435 $Y=1.005
+ $X2=2.435 $Y2=0.68
r188 16 27 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.775 $Y=2.785
+ $X2=2.86 $Y2=2.66
r189 16 18 24.4318 $w=2.48e-07 $l=5.3e-07 $layer=LI1_cond $X=2.775 $Y=2.785
+ $X2=2.245 $Y2=2.785
r190 5 58 600 $w=1.7e-07 $l=3.01993e-07 $layer=licon1_PDIFF $count=1 $X=5.745
+ $Y=2.285 $X2=5.885 $Y2=2.525
r191 4 34 600 $w=1.7e-07 $l=3.97995e-07 $layer=licon1_PDIFF $count=1 $X=3.68
+ $Y=2.32 $X2=3.83 $Y2=2.65
r192 3 18 600 $w=1.7e-07 $l=5.51249e-07 $layer=licon1_PDIFF $count=1 $X=1.955
+ $Y=2.32 $X2=2.245 $Y2=2.745
r193 2 52 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=5.68
+ $Y=0.595 $X2=5.825 $Y2=0.735
r194 1 22 182 $w=1.7e-07 $l=6.21369e-07 $layer=licon1_NDIFF $count=1 $X=1.94
+ $Y=0.395 $X2=2.435 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRBP_2%Q_N 1 2 7 8 9 16 30
r28 30 31 0.96397 $w=4.33e-07 $l=1e-08 $layer=LI1_cond $X=12.247 $Y=0.925
+ $X2=12.247 $Y2=0.915
r29 25 27 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=12.195 $Y=1.985
+ $X2=12.195 $Y2=2.815
r30 9 25 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=12.195 $Y=1.665
+ $X2=12.195 $Y2=1.985
r31 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=12.195 $Y=1.295
+ $X2=12.195 $Y2=1.665
r32 8 33 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=12.195 $Y=1.295
+ $X2=12.195 $Y2=1.085
r33 7 33 3.95767 $w=4.33e-07 $l=1.23e-07 $layer=LI1_cond $X=12.247 $Y=0.962
+ $X2=12.247 $Y2=1.085
r34 7 30 0.980239 $w=4.33e-07 $l=3.7e-08 $layer=LI1_cond $X=12.247 $Y=0.962
+ $X2=12.247 $Y2=0.925
r35 7 31 1.32706 $w=3.28e-07 $l=3.8e-08 $layer=LI1_cond $X=12.3 $Y=0.877
+ $X2=12.3 $Y2=0.915
r36 7 16 12.642 $w=3.28e-07 $l=3.62e-07 $layer=LI1_cond $X=12.3 $Y=0.877
+ $X2=12.3 $Y2=0.515
r37 2 27 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=12.065
+ $Y=1.84 $X2=12.215 $Y2=2.815
r38 2 25 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=12.065
+ $Y=1.84 $X2=12.215 $Y2=1.985
r39 1 16 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=12.16
+ $Y=0.37 $X2=12.3 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRBP_2%Q 1 2 7 10
r16 7 16 35.427 $w=2.68e-07 $l=8.3e-07 $layer=LI1_cond $X=14.19 $Y=1.985
+ $X2=14.19 $Y2=2.815
r17 7 10 62.7441 $w=2.68e-07 $l=1.47e-06 $layer=LI1_cond $X=14.19 $Y=1.985
+ $X2=14.19 $Y2=0.515
r18 2 16 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=14.01
+ $Y=1.84 $X2=14.16 $Y2=2.815
r19 2 7 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=14.01
+ $Y=1.84 $X2=14.16 $Y2=1.985
r20 1 10 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=14.045
+ $Y=0.37 $X2=14.185 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRBP_2%VGND 1 2 3 4 5 6 7 8 9 30 34 38 42 46 50 52
+ 56 58 60 63 64 66 67 69 70 71 73 99 103 108 114 118 122 124 127 130 134
c155 134 0 6.26159e-21 $X=14.64 $Y=0
c156 38 0 9.8593e-20 $X=4.835 $Y=0.965
r157 133 134 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.64 $Y=0
+ $X2=14.64 $Y2=0
r158 130 131 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.68 $Y=0
+ $X2=13.68 $Y2=0
r159 128 131 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=12.72 $Y=0
+ $X2=13.68 $Y2=0
r160 127 128 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r161 124 125 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r162 120 122 7.07024 $w=4.93e-07 $l=6.5e-08 $layer=LI1_cond $X=7.92 $Y=0.162
+ $X2=7.985 $Y2=0.162
r163 120 121 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r164 117 120 4.95346 $w=4.93e-07 $l=2.05e-07 $layer=LI1_cond $X=7.715 $Y=0.162
+ $X2=7.92 $Y2=0.162
r165 117 118 11.9029 $w=4.93e-07 $l=2.65e-07 $layer=LI1_cond $X=7.715 $Y=0.162
+ $X2=7.45 $Y2=0.162
r166 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0
+ $X2=0.72 $Y2=0
r167 112 134 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.16 $Y=0
+ $X2=14.64 $Y2=0
r168 112 131 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.16 $Y=0
+ $X2=13.68 $Y2=0
r169 111 112 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.16 $Y=0
+ $X2=14.16 $Y2=0
r170 109 130 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.84 $Y=0
+ $X2=13.755 $Y2=0
r171 109 111 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=13.84 $Y=0
+ $X2=14.16 $Y2=0
r172 108 133 4.34417 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=14.495 $Y=0
+ $X2=14.687 $Y2=0
r173 108 111 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=14.495 $Y=0
+ $X2=14.16 $Y2=0
r174 107 128 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=12.72 $Y2=0
r175 107 125 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=11.76 $Y2=0
r176 106 107 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r177 104 124 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.895 $Y=0
+ $X2=11.77 $Y2=0
r178 104 106 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=11.895 $Y=0
+ $X2=12.24 $Y2=0
r179 103 127 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=12.635 $Y=0
+ $X2=12.765 $Y2=0
r180 103 106 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=12.635 $Y=0
+ $X2=12.24 $Y2=0
r181 102 125 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=11.76 $Y2=0
r182 101 102 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r183 99 124 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.645 $Y=0
+ $X2=11.77 $Y2=0
r184 99 101 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=11.645 $Y=0
+ $X2=11.28 $Y2=0
r185 98 102 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=11.28 $Y2=0
r186 98 121 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=7.92 $Y2=0
r187 97 122 152.337 $w=1.68e-07 $l=2.335e-06 $layer=LI1_cond $X=10.32 $Y=0
+ $X2=7.985 $Y2=0
r188 97 98 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r189 93 118 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=7.44 $Y=0 $X2=7.45
+ $Y2=0
r190 90 93 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=5.04 $Y=0 $X2=7.44
+ $Y2=0
r191 90 91 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r192 87 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r193 86 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r194 84 87 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r195 83 84 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r196 81 84 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=3.6
+ $Y2=0
r197 81 115 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r198 80 83 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=3.6
+ $Y2=0
r199 80 81 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r200 78 114 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.875 $Y=0
+ $X2=0.71 $Y2=0
r201 78 80 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=1.2
+ $Y2=0
r202 76 115 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0
+ $X2=0.72 $Y2=0
r203 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r204 73 114 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.545 $Y=0
+ $X2=0.71 $Y2=0
r205 73 75 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0
+ $X2=0.24 $Y2=0
r206 71 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=7.92 $Y2=0
r207 71 91 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=7.44 $Y=0 $X2=5.04
+ $Y2=0
r208 71 93 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r209 69 97 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=10.335 $Y=0
+ $X2=10.32 $Y2=0
r210 69 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.335 $Y=0
+ $X2=10.5 $Y2=0
r211 68 101 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=10.665 $Y=0
+ $X2=11.28 $Y2=0
r212 68 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.665 $Y=0
+ $X2=10.5 $Y2=0
r213 66 86 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=4.75 $Y=0 $X2=4.56
+ $Y2=0
r214 66 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.75 $Y=0 $X2=4.835
+ $Y2=0
r215 65 90 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=4.92 $Y=0 $X2=5.04
+ $Y2=0
r216 65 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.92 $Y=0 $X2=4.835
+ $Y2=0
r217 63 83 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=3.64 $Y=0 $X2=3.6
+ $Y2=0
r218 63 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.64 $Y=0 $X2=3.805
+ $Y2=0
r219 62 86 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=3.97 $Y=0 $X2=4.56
+ $Y2=0
r220 62 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.97 $Y=0 $X2=3.805
+ $Y2=0
r221 58 133 3.0545 $w=2.85e-07 $l=1.07121e-07 $layer=LI1_cond $X=14.637 $Y=0.085
+ $X2=14.687 $Y2=0
r222 58 60 17.3877 $w=2.83e-07 $l=4.3e-07 $layer=LI1_cond $X=14.637 $Y=0.085
+ $X2=14.637 $Y2=0.515
r223 54 130 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.755 $Y=0.085
+ $X2=13.755 $Y2=0
r224 54 56 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=13.755 $Y=0.085
+ $X2=13.755 $Y2=0.515
r225 53 127 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=12.895 $Y=0
+ $X2=12.765 $Y2=0
r226 52 130 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.67 $Y=0
+ $X2=13.755 $Y2=0
r227 52 53 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=13.67 $Y=0
+ $X2=12.895 $Y2=0
r228 48 127 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=12.765 $Y=0.085
+ $X2=12.765 $Y2=0
r229 48 50 20.3894 $w=2.58e-07 $l=4.6e-07 $layer=LI1_cond $X=12.765 $Y=0.085
+ $X2=12.765 $Y2=0.545
r230 44 124 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=11.77 $Y=0.085
+ $X2=11.77 $Y2=0
r231 44 46 13.1378 $w=2.48e-07 $l=2.85e-07 $layer=LI1_cond $X=11.77 $Y=0.085
+ $X2=11.77 $Y2=0.37
r232 40 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.5 $Y=0.085
+ $X2=10.5 $Y2=0
r233 40 42 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=10.5 $Y=0.085
+ $X2=10.5 $Y2=0.58
r234 36 67 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.835 $Y=0.085
+ $X2=4.835 $Y2=0
r235 36 38 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=4.835 $Y=0.085
+ $X2=4.835 $Y2=0.965
r236 32 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.805 $Y=0.085
+ $X2=3.805 $Y2=0
r237 32 34 18.1597 $w=3.28e-07 $l=5.2e-07 $layer=LI1_cond $X=3.805 $Y=0.085
+ $X2=3.805 $Y2=0.605
r238 28 114 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0
r239 28 30 18.1597 $w=3.28e-07 $l=5.2e-07 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0.605
r240 9 60 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=14.475
+ $Y=0.37 $X2=14.615 $Y2=0.515
r241 8 56 91 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=2 $X=13.6
+ $Y=0.37 $X2=13.755 $Y2=0.515
r242 7 50 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=12.59
+ $Y=0.37 $X2=12.73 $Y2=0.545
r243 6 46 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=11.685
+ $Y=0.225 $X2=11.81 $Y2=0.37
r244 5 42 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=10.36
+ $Y=0.37 $X2=10.5 $Y2=0.58
r245 4 117 182 $w=1.7e-07 $l=4.34511e-07 $layer=licon1_NDIFF $count=1 $X=7.395
+ $Y=0.595 $X2=7.715 $Y2=0.325
r246 3 38 182 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_NDIFF $count=1 $X=4.695
+ $Y=0.595 $X2=4.835 $Y2=0.965
r247 2 34 182 $w=1.7e-07 $l=2.78747e-07 $layer=licon1_NDIFF $count=1 $X=3.645
+ $Y=0.395 $X2=3.805 $Y2=0.605
r248 1 30 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.395 $X2=0.71 $Y2=0.605
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRBP_2%noxref_25 1 2 9 11 12 15
r35 13 15 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=3.265 $Y=0.425
+ $X2=3.265 $Y2=0.605
r36 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.1 $Y=0.34
+ $X2=3.265 $Y2=0.425
r37 11 12 114.497 $w=1.68e-07 $l=1.755e-06 $layer=LI1_cond $X=3.1 $Y=0.34
+ $X2=1.345 $Y2=0.34
r38 7 12 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.22 $Y=0.425
+ $X2=1.345 $Y2=0.34
r39 7 9 8.29759 $w=2.48e-07 $l=1.8e-07 $layer=LI1_cond $X=1.22 $Y=0.425 $X2=1.22
+ $Y2=0.605
r40 2 15 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.125
+ $Y=0.395 $X2=3.265 $Y2=0.605
r41 1 9 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=1.115
+ $Y=0.395 $X2=1.26 $Y2=0.605
.ends

