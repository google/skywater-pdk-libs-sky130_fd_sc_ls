* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_ls__sedfxtp_4 CLK D DE SCD SCE VGND VNB VPB VPWR Q
*.PININFO CLK:I D:I DE:I SCD:I SCE:I VGND:I VNB:I VPB:I VPWR:I Q:O
MI14 net146 M1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=1.12 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI13 S0 clkneg net146 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S0 VPWR VPB pfet_01v8_hvt m=4 w=1.12 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net114 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=1.12 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net118 q1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net118 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net114 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 q1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net107 deneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 net98 sceneg db VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 VPWR SCD net98 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 net95 D net107 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 net95 SCE db VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 net87 q1 net95 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI36 deneg DE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 VPWR DE net87 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 sceneg SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.74 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.74 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net222 q1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net222 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S0 VGND VNB nfet_01v8 m=4 w=0.74 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net211 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 M0 clkpos net211 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 net95 sceneg db VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 q1 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 sceneg SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net95 D net167 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 net187 M1 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI15 S0 clkpos net187 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI41 net174 q1 net95 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 VGND deneg net174 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 deneg DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net167 DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI49 net163 SCE db VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI48 VGND SCD net163 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_sc_ls__sedfxtp_4
