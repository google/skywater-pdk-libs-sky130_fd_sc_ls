* NGSPICE file created from sky130_fd_sc_ls__a21bo_1.ext - technology: sky130A

.subckt sky130_fd_sc_ls__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
M1000 a_194_136# a_272_110# a_34_392# VPB phighvt w=1e+06u l=150000u
+  ad=2.75e+11p pd=2.55e+06u as=5.75e+11p ps=5.15e+06u
M1001 a_122_136# A2 VGND VNB nshort w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=5.6545e+11p ps=5.75e+06u
M1002 X a_194_136# VGND VNB nshort w=740000u l=150000u
+  ad=1.961e+11p pd=2.01e+06u as=0p ps=0u
M1003 VGND a_272_110# a_194_136# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=2.496e+11p ps=2.06e+06u
M1004 VPWR A2 a_34_392# VPB phighvt w=1e+06u l=150000u
+  ad=7.36e+11p pd=5.67e+06u as=0p ps=0u
M1005 VPWR B1_N a_272_110# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=2.31e+11p ps=2.23e+06u
M1006 VGND B1_N a_272_110# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1007 a_194_136# A1 a_122_136# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_34_392# A1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 X a_194_136# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.08e+11p pd=2.79e+06u as=0p ps=0u
.ends

