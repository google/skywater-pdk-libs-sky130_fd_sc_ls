* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__dfsbp_2 CLK D SET_B VGND VNB VPB VPWR Q Q_N
X0 a_2221_74# a_1339_74# VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X1 a_1521_508# a_1501_92# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 a_225_74# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X3 VGND a_2221_74# Q VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X4 a_595_97# a_225_74# a_706_463# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 VPWR a_2221_74# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X6 a_1339_74# a_398_74# a_1521_508# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 a_595_97# a_398_74# a_731_97# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_225_74# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X9 VPWR a_595_97# a_1258_341# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_706_463# a_757_401# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X11 a_731_97# a_757_401# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 a_757_401# a_595_97# a_1001_74# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 VGND a_1339_74# Q_N VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X14 VGND a_225_74# a_398_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X15 Q a_2221_74# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X16 VPWR a_595_97# a_757_401# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X17 VPWR SET_B a_1339_74# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X18 a_757_401# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X19 a_27_74# a_225_74# a_595_97# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 VPWR a_1339_74# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X21 a_1001_74# SET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X22 a_1261_74# a_398_74# a_1339_74# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X23 a_1339_74# a_225_74# a_1453_118# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X24 Q a_2221_74# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X25 a_2221_74# a_1339_74# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X26 a_27_74# a_398_74# a_595_97# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X27 VGND a_595_97# a_1261_74# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X28 a_1258_341# a_225_74# a_1339_74# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X29 VPWR a_225_74# a_398_74# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X30 a_1453_118# a_1501_92# a_1531_118# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X31 VGND a_1339_74# a_1501_92# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X32 a_27_74# D VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X33 Q_N a_1339_74# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X34 a_27_74# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X35 Q_N a_1339_74# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X36 a_1501_92# a_1339_74# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X37 a_1531_118# SET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
