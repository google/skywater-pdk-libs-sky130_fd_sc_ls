* File: sky130_fd_sc_ls__dfstp_4.spice
* Created: Wed Sep  2 11:01:56 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__dfstp_4.pex.spice"
.subckt sky130_fd_sc_ls__dfstp_4  VNB VPB D CLK SET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* SET_B	SET_B
* CLK	CLK
* D	D
* VPB	VPB
* VNB	VNB
MM1035 N_VGND_M1035_d N_D_M1035_g N_A_27_74#_M1035_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.1197 PD=1.41 PS=1.41 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1037 N_VGND_M1037_d N_CLK_M1037_g N_A_225_74#_M1037_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1022 N_A_398_74#_M1022_d N_A_225_74#_M1022_g N_VGND_M1037_d VNB NSHORT L=0.15
+ W=0.74 AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1027 N_A_612_74#_M1027_d N_A_225_74#_M1027_g N_A_27_74#_M1027_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0945 AS=0.18665 PD=0.87 PS=1.8 NRD=48.564 NRS=24.276 M=1
+ R=2.8 SA=75000.3 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1017 A_732_74# N_A_398_74#_M1017_g N_A_612_74#_M1027_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.0945 PD=0.66 PS=0.87 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75000.9 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_A_767_402#_M1001_g A_732_74# VNB NSHORT L=0.15 W=0.42
+ AD=0.147 AS=0.0504 PD=1.54 PS=0.66 NRD=8.568 NRS=18.564 M=1 R=2.8 SA=75001.3
+ SB=75000.3 A=0.063 P=1.14 MULT=1
MM1029 A_1035_118# N_A_612_74#_M1029_g N_A_767_402#_M1029_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.1491 PD=0.66 PS=1.55 NRD=18.564 NRS=9.996 M=1 R=2.8
+ SA=75000.3 SB=75003.3 A=0.063 P=1.14 MULT=1
MM1020 N_VGND_M1020_d N_SET_B_M1020_g A_1035_118# VNB NSHORT L=0.15 W=0.42
+ AD=0.0930736 AS=0.0504 PD=0.832075 PS=0.66 NRD=37.848 NRS=18.564 M=1 R=2.8
+ SA=75000.7 SB=75002.9 A=0.063 P=1.14 MULT=1
MM1031 A_1225_74# N_A_612_74#_M1031_g N_VGND_M1020_d VNB NSHORT L=0.15 W=0.64
+ AD=0.1264 AS=0.141826 PD=1.035 PS=1.26792 NRD=26.712 NRS=0 M=1 R=4.26667
+ SA=75000.9 SB=75002.4 A=0.096 P=1.58 MULT=1
MM1003 N_A_1321_392#_M1003_d N_A_398_74#_M1003_g A_1225_74# VNB NSHORT L=0.15
+ W=0.64 AD=0.127668 AS=0.1264 PD=1.20755 PS=1.035 NRD=0 NRS=26.712 M=1
+ R=4.26667 SA=75001.4 SB=75001.8 A=0.096 P=1.58 MULT=1
MM1018 A_1436_88# N_A_225_74#_M1018_g N_A_1321_392#_M1003_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.0837821 PD=0.66 PS=0.792453 NRD=18.564 NRS=22.848 M=1
+ R=2.8 SA=75001.9 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1004 A_1514_88# N_A_1484_62#_M1004_g A_1436_88# VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0504 PD=0.66 PS=0.66 NRD=18.564 NRS=18.564 M=1 R=2.8 SA=75002.3
+ SB=75001.8 A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1005_d N_SET_B_M1005_g A_1514_88# VNB NSHORT L=0.15 W=0.42
+ AD=0.21735 AS=0.0504 PD=1.455 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75002.7
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1002 N_A_1484_62#_M1002_d N_A_1321_392#_M1002_g N_VGND_M1005_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.1197 AS=0.21735 PD=1.41 PS=1.455 NRD=0 NRS=19.992 M=1 R=2.8
+ SA=75003.9 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1038 N_VGND_M1038_d N_A_1321_392#_M1038_g N_A_1940_74#_M1038_s VNB NSHORT
+ L=0.15 W=0.74 AD=0.1295 AS=0.2627 PD=1.09 PS=2.19 NRD=0 NRS=11.34 M=1
+ R=4.93333 SA=75000.3 SB=75002.5 A=0.111 P=1.78 MULT=1
MM1006 N_Q_M1006_d N_A_1940_74#_M1006_g N_VGND_M1038_d VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75000.8
+ SB=75002 A=0.111 P=1.78 MULT=1
MM1009 N_Q_M1006_d N_A_1940_74#_M1009_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.2627 PD=1.02 PS=1.45 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.2
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1021 N_Q_M1021_d N_A_1940_74#_M1021_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.74
+ AD=0.12025 AS=0.2627 PD=1.065 PS=1.45 NRD=7.296 NRS=0 M=1 R=4.93333 SA=75002.1
+ SB=75000.8 A=0.111 P=1.78 MULT=1
MM1036 N_Q_M1021_d N_A_1940_74#_M1036_g N_VGND_M1036_s VNB NSHORT L=0.15 W=0.74
+ AD=0.12025 AS=0.2627 PD=1.065 PS=2.19 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75002.5
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1033 N_VPWR_M1033_d N_D_M1033_g N_A_27_74#_M1033_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1239 AS=0.1239 PD=1.43 PS=1.43 NRD=4.6886 NRS=4.6886 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1026 N_VPWR_M1026_d N_CLK_M1026_g N_A_225_74#_M1026_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1034 N_A_398_74#_M1034_d N_A_225_74#_M1034_g N_VPWR_M1026_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1010 N_A_612_74#_M1010_d N_A_398_74#_M1010_g N_A_27_74#_M1010_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0735 AS=0.1239 PD=0.77 PS=1.43 NRD=28.1316 NRS=4.6886 M=1
+ R=2.8 SA=75000.2 SB=75004.5 A=0.063 P=1.14 MULT=1
MM1019 A_716_463# N_A_225_74#_M1019_g N_A_612_74#_M1010_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0567 AS=0.0735 PD=0.69 PS=0.77 NRD=37.5088 NRS=4.6886 M=1 R=2.8
+ SA=75000.7 SB=75004 A=0.063 P=1.14 MULT=1
MM1011 N_VPWR_M1011_d N_A_767_402#_M1011_g A_716_463# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.16485 AS=0.0567 PD=1.205 PS=0.69 NRD=11.7215 NRS=37.5088 M=1 R=2.8
+ SA=75001.1 SB=75003.6 A=0.063 P=1.14 MULT=1
MM1000 N_A_767_402#_M1000_d N_A_612_74#_M1000_g N_VPWR_M1011_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.063 AS=0.16485 PD=0.72 PS=1.205 NRD=4.6886 NRS=225.132 M=1
+ R=2.8 SA=75002.1 SB=75002.6 A=0.063 P=1.14 MULT=1
MM1007 N_VPWR_M1007_d N_SET_B_M1007_g N_A_767_402#_M1000_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.115648 AS=0.063 PD=0.925775 PS=0.72 NRD=114.91 NRS=4.6886 M=1
+ R=2.8 SA=75002.5 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1014 A_1220_347# N_A_612_74#_M1014_g N_VPWR_M1007_d VPB PHIGHVT L=0.15 W=1
+ AD=0.197187 AS=0.275352 PD=1.58 PS=2.20423 NRD=27.9937 NRS=7.8603 M=1
+ R=6.66667 SA=75001.5 SB=75000.9 A=0.15 P=2.3 MULT=1
MM1013 N_A_1321_392#_M1013_d N_A_225_74#_M1013_g A_1220_347# VPB PHIGHVT L=0.15
+ W=1 AD=0.305141 AS=0.197187 PD=2.3169 PS=1.58 NRD=1.9503 NRS=27.9937 M=1
+ R=6.66667 SA=75001.9 SB=75000.9 A=0.15 P=2.3 MULT=1
MM1028 A_1480_508# N_A_398_74#_M1028_g N_A_1321_392#_M1013_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0567 AS=0.128159 PD=0.69 PS=0.973099 NRD=37.5088 NRS=86.7588 M=1
+ R=2.8 SA=75002.6 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1024 N_VPWR_M1024_d N_A_1484_62#_M1024_g A_1480_508# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.063 AS=0.0567 PD=0.72 PS=0.69 NRD=4.6886 NRS=37.5088 M=1 R=2.8 SA=75003.1
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1032 N_A_1321_392#_M1032_d N_SET_B_M1032_g N_VPWR_M1024_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1155 AS=0.063 PD=1.39 PS=0.72 NRD=4.6886 NRS=4.6886 M=1 R=2.8
+ SA=75003.5 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1030 N_A_1484_62#_M1030_d N_A_1321_392#_M1030_g N_VPWR_M1030_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.1155 AS=0.1176 PD=1.39 PS=1.4 NRD=4.6886 NRS=4.6886 M=1
+ R=2.8 SA=75000.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1012 N_A_1940_74#_M1012_d N_A_1321_392#_M1012_g N_VPWR_M1012_s VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.126 AS=0.2352 PD=1.14 PS=2.24 NRD=2.3443 NRS=2.3443 M=1
+ R=5.6 SA=75000.2 SB=75002.5 A=0.126 P=1.98 MULT=1
MM1023 N_A_1940_74#_M1012_d N_A_1321_392#_M1023_g N_VPWR_M1023_s VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.126 AS=0.1668 PD=1.14 PS=1.27714 NRD=2.3443 NRS=18.7544 M=1
+ R=5.6 SA=75000.7 SB=75002.1 A=0.126 P=1.98 MULT=1
MM1008 N_VPWR_M1023_s N_A_1940_74#_M1008_g N_Q_M1008_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.2224 AS=0.168 PD=1.70286 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.9 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1015 N_VPWR_M1015_d N_A_1940_74#_M1015_g N_Q_M1008_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.4 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1016 N_VPWR_M1015_d N_A_1940_74#_M1016_g N_Q_M1016_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.8 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1025 N_VPWR_M1025_d N_A_1940_74#_M1025_g N_Q_M1016_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3192 AS=0.168 PD=2.81 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.3 SB=75000.2 A=0.168 P=2.54 MULT=1
DX39_noxref VNB VPB NWDIODE A=24.9216 P=30.61
c_136 VNB 0 7.64129e-20 $X=0 $Y=0
c_1752 A_716_463# 0 1.99261e-20 $X=3.58 $Y=2.315
*
.include "sky130_fd_sc_ls__dfstp_4.pxi.spice"
*
.ends
*
*
