* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__xnor3_4 A B C VGND VNB VPB VPWR X
X0 X a_1057_74# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X1 a_324_373# a_386_23# a_75_227# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X2 X a_1057_74# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X3 VGND A a_75_227# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X4 a_27_373# a_75_227# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_75_227# B a_324_373# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X6 VPWR a_1057_74# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X7 a_27_373# a_75_227# VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X8 a_1024_300# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X9 VPWR A a_75_227# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 VPWR a_1057_74# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X11 a_386_23# B VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X12 a_27_373# B a_321_77# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X13 a_321_77# a_386_23# a_27_373# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 a_386_23# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X15 a_75_227# B a_321_77# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X16 X a_1057_74# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X17 a_1024_300# C VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 VGND a_1057_74# X VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X19 a_321_77# a_386_23# a_75_227# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X20 a_321_77# a_1024_300# a_1057_74# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X21 X a_1057_74# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X22 a_1057_74# C a_321_77# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X23 a_324_373# a_1024_300# a_1057_74# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X24 a_1057_74# C a_324_373# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X25 a_324_373# a_386_23# a_27_373# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X26 a_27_373# B a_324_373# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X27 VGND a_1057_74# X VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
.ends
