* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__sdfxtp_2 CLK D SCD SCE VGND VNB VPB VPWR Q
M1000 VGND SCD a_442_74# VNB nshort w=420000u l=150000u
+  ad=1.84785e+12p pd=1.542e+07u as=1.008e+11p ps=1.32e+06u
M1001 VGND a_1829_398# Q VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.405e+11p ps=2.13e+06u
M1002 a_1219_100# a_846_74# a_1044_100# VNB nshort w=420000u l=150000u
+  ad=1.764e+11p pd=1.68e+06u as=3.045e+11p ps=2.29e+06u
M1003 a_1287_320# a_1044_100# VGND VNB nshort w=550000u l=150000u
+  ad=3.795e+11p pd=2.48e+06u as=0p ps=0u
M1004 a_634_74# CLK VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=2.86313e+12p ps=2.094e+07u
M1005 VPWR a_1287_320# a_1210_508# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.68e+11p ps=1.64e+06u
M1006 a_439_453# a_27_74# a_300_453# VPB phighvt w=640000u l=150000u
+  ad=1.728e+11p pd=1.82e+06u as=4.727e+11p ps=3.8e+06u
M1007 a_1287_320# a_1044_100# VPWR VPB phighvt w=840000u l=150000u
+  ad=4.452e+11p pd=2.74e+06u as=0p ps=0u
M1008 VGND a_1287_320# a_1219_100# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Q a_1829_398# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=0p ps=0u
M1010 a_1592_424# a_846_74# a_1287_320# VNB nshort w=550000u l=150000u
+  ad=1.8825e+11p pd=1.82e+06u as=0p ps=0u
M1011 a_1704_496# a_846_74# a_1592_424# VPB phighvt w=420000u l=150000u
+  ad=2.688e+11p pd=2.12e+06u as=2.943e+11p ps=2.5e+06u
M1012 a_442_74# SCE a_300_453# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=3.528e+11p ps=3.36e+06u
M1013 a_300_453# D a_216_453# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1014 a_223_74# a_27_74# VGND VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1015 a_300_453# D a_223_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_1829_398# a_1592_424# VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1017 VPWR SCD a_439_453# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_1829_398# a_1592_424# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.95e+11p pd=2.59e+06u as=0p ps=0u
M1019 VPWR a_1829_398# Q VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_1787_74# a_634_74# a_1592_424# VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1021 VGND a_1829_398# a_1787_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_216_453# SCE VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 Q a_1829_398# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VPWR SCE a_27_74# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.888e+11p ps=1.87e+06u
M1025 a_1592_424# a_634_74# a_1287_320# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_1044_100# a_846_74# a_300_453# VPB phighvt w=420000u l=150000u
+  ad=1.26e+11p pd=1.44e+06u as=0p ps=0u
M1027 a_846_74# a_634_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=0p ps=0u
M1028 a_846_74# a_634_74# VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1029 a_634_74# CLK VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1030 VGND SCE a_27_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.386e+11p ps=1.5e+06u
M1031 a_1210_508# a_634_74# a_1044_100# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 VPWR a_1829_398# a_1704_496# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_1044_100# a_634_74# a_300_453# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
