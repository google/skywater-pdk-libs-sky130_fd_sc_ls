# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_ls__nand2b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_ls__nand2b_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A_N
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.350000 0.570000 1.780000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445000 1.350000 2.775000 1.780000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  0.879200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.645000 1.820000 2.275000 1.950000 ;
        RECT 1.645000 1.950000 2.795000 2.200000 ;
        RECT 1.700000 0.630000 1.870000 1.220000 ;
        RECT 1.700000 1.220000 2.275000 1.390000 ;
        RECT 2.045000 1.390000 2.275000 1.820000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000000 0.000000 3.360000 0.245000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.660000 3.550000 3.520000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.115000  0.350000 0.445000 1.010000 ;
      RECT 0.115000  1.010000 0.975000 1.140000 ;
      RECT 0.115000  1.140000 1.135000 1.180000 ;
      RECT 0.115000  1.950000 0.975000 2.120000 ;
      RECT 0.115000  2.120000 0.445000 2.860000 ;
      RECT 0.615000  0.085000 0.875000 0.840000 ;
      RECT 0.725000  2.290000 1.095000 3.245000 ;
      RECT 0.805000  1.180000 1.135000 1.470000 ;
      RECT 0.805000  1.470000 0.975000 1.950000 ;
      RECT 1.190000  0.255000 2.380000 0.425000 ;
      RECT 1.190000  0.425000 1.520000 0.970000 ;
      RECT 1.305000  0.970000 1.475000 2.370000 ;
      RECT 1.305000  2.370000 3.245000 2.540000 ;
      RECT 2.015000  2.710000 2.345000 3.245000 ;
      RECT 2.050000  0.425000 2.380000 1.050000 ;
      RECT 2.560000  0.085000 2.730000 1.130000 ;
      RECT 2.915000  0.350000 3.245000 1.130000 ;
      RECT 2.915000  2.710000 3.245000 3.245000 ;
      RECT 3.075000  1.130000 3.245000 2.370000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_ls__nand2b_2
END LIBRARY
