* File: sky130_fd_sc_ls__bufbuf_8.pxi.spice
* Created: Fri Aug 28 13:07:45 2020
* 
x_PM_SKY130_FD_SC_LS__BUFBUF_8%A N_A_M1015_g N_A_c_126_n N_A_M1018_g A
+ N_A_c_127_n PM_SKY130_FD_SC_LS__BUFBUF_8%A
x_PM_SKY130_FD_SC_LS__BUFBUF_8%A_27_112# N_A_27_112#_M1015_s N_A_27_112#_M1018_s
+ N_A_27_112#_c_159_n N_A_27_112#_M1000_g N_A_27_112#_M1012_g
+ N_A_27_112#_c_161_n N_A_27_112#_c_167_n N_A_27_112#_c_168_n
+ N_A_27_112#_c_178_n N_A_27_112#_c_162_n N_A_27_112#_c_163_n
+ N_A_27_112#_c_164_n N_A_27_112#_c_165_n PM_SKY130_FD_SC_LS__BUFBUF_8%A_27_112#
x_PM_SKY130_FD_SC_LS__BUFBUF_8%A_221_368# N_A_221_368#_M1012_d
+ N_A_221_368#_M1000_d N_A_221_368#_c_241_n N_A_221_368#_M1007_g
+ N_A_221_368#_M1004_g N_A_221_368#_c_242_n N_A_221_368#_M1014_g
+ N_A_221_368#_M1013_g N_A_221_368#_M1022_g N_A_221_368#_c_243_n
+ N_A_221_368#_M1020_g N_A_221_368#_c_244_n N_A_221_368#_c_233_n
+ N_A_221_368#_c_234_n N_A_221_368#_c_235_n N_A_221_368#_c_245_n
+ N_A_221_368#_c_236_n N_A_221_368#_c_237_n N_A_221_368#_c_238_n
+ N_A_221_368#_c_239_n N_A_221_368#_c_240_n
+ PM_SKY130_FD_SC_LS__BUFBUF_8%A_221_368#
x_PM_SKY130_FD_SC_LS__BUFBUF_8%A_334_368# N_A_334_368#_M1004_d
+ N_A_334_368#_M1013_d N_A_334_368#_M1007_s N_A_334_368#_M1014_s
+ N_A_334_368#_M1002_g N_A_334_368#_c_343_n N_A_334_368#_M1001_g
+ N_A_334_368#_M1005_g N_A_334_368#_c_344_n N_A_334_368#_M1003_g
+ N_A_334_368#_M1006_g N_A_334_368#_c_345_n N_A_334_368#_M1008_g
+ N_A_334_368#_M1010_g N_A_334_368#_c_346_n N_A_334_368#_M1009_g
+ N_A_334_368#_M1011_g N_A_334_368#_c_347_n N_A_334_368#_M1016_g
+ N_A_334_368#_M1019_g N_A_334_368#_c_348_n N_A_334_368#_M1017_g
+ N_A_334_368#_c_349_n N_A_334_368#_M1021_g N_A_334_368#_M1023_g
+ N_A_334_368#_M1025_g N_A_334_368#_c_350_n N_A_334_368#_M1024_g
+ N_A_334_368#_c_351_n N_A_334_368#_c_352_n N_A_334_368#_c_337_n
+ N_A_334_368#_c_338_n N_A_334_368#_c_353_n N_A_334_368#_c_354_n
+ N_A_334_368#_c_339_n N_A_334_368#_c_340_n N_A_334_368#_c_356_n
+ N_A_334_368#_c_341_n N_A_334_368#_c_342_n
+ PM_SKY130_FD_SC_LS__BUFBUF_8%A_334_368#
x_PM_SKY130_FD_SC_LS__BUFBUF_8%VPWR N_VPWR_M1018_d N_VPWR_M1007_d N_VPWR_M1020_d
+ N_VPWR_M1003_s N_VPWR_M1009_s N_VPWR_M1017_s N_VPWR_M1024_s N_VPWR_c_526_n
+ N_VPWR_c_527_n N_VPWR_c_528_n N_VPWR_c_529_n N_VPWR_c_530_n N_VPWR_c_531_n
+ N_VPWR_c_532_n N_VPWR_c_533_n N_VPWR_c_534_n N_VPWR_c_535_n VPWR
+ N_VPWR_c_536_n N_VPWR_c_537_n N_VPWR_c_538_n N_VPWR_c_539_n N_VPWR_c_540_n
+ N_VPWR_c_541_n N_VPWR_c_542_n N_VPWR_c_543_n N_VPWR_c_544_n N_VPWR_c_545_n
+ N_VPWR_c_546_n N_VPWR_c_525_n PM_SKY130_FD_SC_LS__BUFBUF_8%VPWR
x_PM_SKY130_FD_SC_LS__BUFBUF_8%X N_X_M1002_d N_X_M1006_d N_X_M1011_d N_X_M1023_d
+ N_X_M1001_d N_X_M1008_d N_X_M1016_d N_X_M1021_d N_X_c_634_n N_X_c_639_n
+ N_X_c_635_n N_X_c_636_n N_X_c_640_n N_X_c_641_n N_X_c_642_n N_X_c_643_n
+ N_X_c_644_n N_X_c_645_n N_X_c_637_n N_X_c_638_n N_X_c_647_n N_X_c_648_n
+ N_X_c_649_n X X PM_SKY130_FD_SC_LS__BUFBUF_8%X
x_PM_SKY130_FD_SC_LS__BUFBUF_8%VGND N_VGND_M1015_d N_VGND_M1004_s N_VGND_M1022_s
+ N_VGND_M1005_s N_VGND_M1010_s N_VGND_M1019_s N_VGND_M1025_s N_VGND_c_744_n
+ N_VGND_c_745_n N_VGND_c_746_n N_VGND_c_747_n N_VGND_c_748_n N_VGND_c_749_n
+ N_VGND_c_750_n N_VGND_c_751_n VGND N_VGND_c_752_n N_VGND_c_753_n
+ N_VGND_c_754_n N_VGND_c_755_n N_VGND_c_756_n N_VGND_c_757_n N_VGND_c_758_n
+ N_VGND_c_759_n N_VGND_c_760_n N_VGND_c_761_n N_VGND_c_762_n N_VGND_c_763_n
+ N_VGND_c_764_n N_VGND_c_765_n PM_SKY130_FD_SC_LS__BUFBUF_8%VGND
cc_1 VNB N_A_M1015_g 0.0339682f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.835
cc_2 VNB N_A_c_126_n 0.027776f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_3 VNB N_A_c_127_n 0.0150187f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.515
cc_4 VNB N_A_27_112#_c_159_n 0.0350459f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.26
cc_5 VNB N_A_27_112#_M1012_g 0.0274055f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.515
cc_6 VNB N_A_27_112#_c_161_n 0.0214174f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.565
cc_7 VNB N_A_27_112#_c_162_n 0.00593404f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_27_112#_c_163_n 0.00982632f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_27_112#_c_164_n 0.00808778f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_27_112#_c_165_n 4.00537e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_221_368#_M1004_g 0.0258021f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.515
cc_12 VNB N_A_221_368#_M1013_g 0.0203202f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_221_368#_M1022_g 0.0198048f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_221_368#_c_233_n 0.00853307f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_221_368#_c_234_n 0.00360834f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_221_368#_c_235_n 0.00327963f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_221_368#_c_236_n 6.23805e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_221_368#_c_237_n 0.00819829f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_221_368#_c_238_n 0.00231516f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_221_368#_c_239_n 0.0485727f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_221_368#_c_240_n 0.069295f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_334_368#_M1002_g 0.0223012f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_334_368#_M1005_g 0.0217877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_334_368#_M1006_g 0.0212331f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_334_368#_M1010_g 0.0203701f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_334_368#_M1011_g 0.0211262f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_334_368#_M1019_g 0.021979f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_334_368#_M1023_g 0.0210832f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_334_368#_M1025_g 0.0260098f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_334_368#_c_337_n 0.00373398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_334_368#_c_338_n 0.00690186f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_334_368#_c_339_n 2.73442e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_334_368#_c_340_n 0.00736042f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_334_368#_c_341_n 0.0120893f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_334_368#_c_342_n 0.219745f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VPWR_c_525_n 0.302998f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_X_c_634_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_X_c_635_n 0.0131511f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_X_c_636_n 0.00230427f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_X_c_637_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_X_c_638_n 0.0229756f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_744_n 0.0168478f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_745_n 0.00323505f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_746_n 0.00498656f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_747_n 0.00498656f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_748_n 0.00258815f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_749_n 0.00506929f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_750_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_751_n 0.041823f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_752_n 0.0202692f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_753_n 0.0319969f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_754_n 0.016486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_755_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_756_n 0.016486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_757_n 0.0183953f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_758_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_759_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_760_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_761_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_762_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_763_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_764_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_765_n 0.421461f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VPB N_A_c_126_n 0.0335881f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_65 VPB N_A_c_127_n 0.00758331f $X=-0.19 $Y=1.66 $X2=0.405 $Y2=1.515
cc_66 VPB N_A_27_112#_c_159_n 0.0280835f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.26
cc_67 VPB N_A_27_112#_c_167_n 0.010868f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_A_27_112#_c_168_n 0.0222078f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_A_27_112#_c_165_n 0.00281858f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_A_221_368#_c_241_n 0.0195927f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.26
cc_71 VPB N_A_221_368#_c_242_n 0.0153937f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_A_221_368#_c_243_n 0.0159418f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_A_221_368#_c_244_n 0.0130657f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_A_221_368#_c_245_n 0.00891107f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_A_221_368#_c_236_n 0.00348542f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_A_221_368#_c_240_n 0.0205477f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_A_334_368#_c_343_n 0.0158416f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_A_334_368#_c_344_n 0.0157265f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 VPB N_A_334_368#_c_345_n 0.0153396f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 VPB N_A_334_368#_c_346_n 0.0153788f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_A_334_368#_c_347_n 0.0153784f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 VPB N_A_334_368#_c_348_n 0.0153394f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 VPB N_A_334_368#_c_349_n 0.015193f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_84 VPB N_A_334_368#_c_350_n 0.0180049f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_A_334_368#_c_351_n 0.00349831f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_A_334_368#_c_352_n 0.0107973f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_A_334_368#_c_353_n 0.00187314f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_A_334_368#_c_354_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_A_334_368#_c_339_n 0.00150252f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB N_A_334_368#_c_356_n 0.00119925f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB N_A_334_368#_c_342_n 0.0524541f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_526_n 0.0190202f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_527_n 0.00790074f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_528_n 0.0186948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_529_n 0.00845326f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_530_n 0.0185672f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_531_n 0.00755981f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_532_n 0.00771277f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_533_n 0.00764f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_534_n 0.0131454f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_535_n 0.0513568f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_102 VPB N_VPWR_c_536_n 0.0189402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 VPB N_VPWR_c_537_n 0.0334841f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB N_VPWR_c_538_n 0.0183651f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_105 VPB N_VPWR_c_539_n 0.0178906f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_VPWR_c_540_n 0.0178906f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB N_VPWR_c_541_n 0.00680245f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_VPWR_c_542_n 0.0043981f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_109 VPB N_VPWR_c_543_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_110 VPB N_VPWR_c_544_n 0.00487897f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_VPWR_c_545_n 0.00526366f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_546_n 0.00516749f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_VPWR_c_525_n 0.0966136f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_X_c_639_n 0.00268029f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_X_c_640_n 0.00216667f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_X_c_641_n 0.00209466f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_X_c_642_n 0.00253854f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_X_c_643_n 0.00199268f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_X_c_644_n 0.00271871f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_X_c_645_n 0.00216921f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_X_c_638_n 0.0117101f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_X_c_647_n 0.00271871f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_X_c_648_n 0.00153495f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_X_c_649_n 0.00165774f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 N_A_M1015_g N_A_27_112#_c_159_n 0.0178757f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_126 N_A_c_126_n N_A_27_112#_c_159_n 0.0258689f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_127 N_A_c_127_n N_A_27_112#_c_159_n 3.14462e-19 $X=0.405 $Y=1.515 $X2=0 $Y2=0
cc_128 N_A_M1015_g N_A_27_112#_M1012_g 0.0175574f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_129 N_A_M1015_g N_A_27_112#_c_161_n 0.00900949f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_130 N_A_c_126_n N_A_27_112#_c_167_n 8.45428e-19 $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_131 N_A_c_127_n N_A_27_112#_c_167_n 0.0222448f $X=0.405 $Y=1.515 $X2=0 $Y2=0
cc_132 N_A_c_126_n N_A_27_112#_c_168_n 0.00208622f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_133 N_A_c_126_n N_A_27_112#_c_178_n 0.0151929f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_134 N_A_c_127_n N_A_27_112#_c_178_n 0.0126353f $X=0.405 $Y=1.515 $X2=0 $Y2=0
cc_135 N_A_M1015_g N_A_27_112#_c_162_n 0.0112899f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_136 N_A_c_126_n N_A_27_112#_c_162_n 2.93656e-19 $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_137 N_A_c_127_n N_A_27_112#_c_162_n 0.00908651f $X=0.405 $Y=1.515 $X2=0 $Y2=0
cc_138 N_A_M1015_g N_A_27_112#_c_163_n 0.00377582f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_139 N_A_c_126_n N_A_27_112#_c_163_n 0.00418411f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_140 N_A_c_127_n N_A_27_112#_c_163_n 0.0277302f $X=0.405 $Y=1.515 $X2=0 $Y2=0
cc_141 N_A_M1015_g N_A_27_112#_c_164_n 0.00384276f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_142 N_A_c_126_n N_A_27_112#_c_164_n 9.84981e-19 $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_143 N_A_c_127_n N_A_27_112#_c_164_n 0.0221059f $X=0.405 $Y=1.515 $X2=0 $Y2=0
cc_144 N_A_c_126_n N_A_27_112#_c_165_n 0.00450098f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_145 N_A_c_127_n N_A_27_112#_c_165_n 0.0109521f $X=0.405 $Y=1.515 $X2=0 $Y2=0
cc_146 N_A_c_126_n N_A_221_368#_c_244_n 8.64489e-19 $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_147 N_A_M1015_g N_A_221_368#_c_233_n 8.51156e-19 $X=0.495 $Y=0.835 $X2=0
+ $Y2=0
cc_148 N_A_c_126_n N_VPWR_c_526_n 0.010189f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_149 N_A_c_126_n N_VPWR_c_536_n 0.00361294f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_150 N_A_c_126_n N_VPWR_c_525_n 0.00419404f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_151 N_A_M1015_g N_VGND_c_744_n 0.00507175f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_152 N_A_M1015_g N_VGND_c_752_n 0.0043356f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_153 N_A_M1015_g N_VGND_c_765_n 0.00487769f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_154 N_A_27_112#_c_159_n N_A_221_368#_c_244_n 0.012536f $X=1.03 $Y=1.765 $X2=0
+ $Y2=0
cc_155 N_A_27_112#_M1012_g N_A_221_368#_c_233_n 0.00926861f $X=1.075 $Y=0.74
+ $X2=0 $Y2=0
cc_156 N_A_27_112#_M1012_g N_A_221_368#_c_234_n 0.00367276f $X=1.075 $Y=0.74
+ $X2=0 $Y2=0
cc_157 N_A_27_112#_c_164_n N_A_221_368#_c_234_n 0.0074024f $X=0.835 $Y=1.63
+ $X2=0 $Y2=0
cc_158 N_A_27_112#_c_159_n N_A_221_368#_c_245_n 0.00357744f $X=1.03 $Y=1.765
+ $X2=0 $Y2=0
cc_159 N_A_27_112#_c_164_n N_A_221_368#_c_245_n 0.00375309f $X=0.835 $Y=1.63
+ $X2=0 $Y2=0
cc_160 N_A_27_112#_c_165_n N_A_221_368#_c_245_n 0.00571905f $X=0.835 $Y=1.95
+ $X2=0 $Y2=0
cc_161 N_A_27_112#_c_159_n N_A_221_368#_c_236_n 0.00403171f $X=1.03 $Y=1.765
+ $X2=0 $Y2=0
cc_162 N_A_27_112#_c_165_n N_A_221_368#_c_236_n 0.00796192f $X=0.835 $Y=1.95
+ $X2=0 $Y2=0
cc_163 N_A_27_112#_M1012_g N_A_221_368#_c_237_n 0.00358918f $X=1.075 $Y=0.74
+ $X2=0 $Y2=0
cc_164 N_A_27_112#_c_164_n N_A_221_368#_c_237_n 0.00977888f $X=0.835 $Y=1.63
+ $X2=0 $Y2=0
cc_165 N_A_27_112#_c_159_n N_A_221_368#_c_238_n 0.0027735f $X=1.03 $Y=1.765
+ $X2=0 $Y2=0
cc_166 N_A_27_112#_c_164_n N_A_221_368#_c_238_n 0.0282875f $X=0.835 $Y=1.63
+ $X2=0 $Y2=0
cc_167 N_A_27_112#_c_159_n N_A_221_368#_c_239_n 0.00950058f $X=1.03 $Y=1.765
+ $X2=0 $Y2=0
cc_168 N_A_27_112#_c_164_n N_A_221_368#_c_239_n 2.93865e-19 $X=0.835 $Y=1.63
+ $X2=0 $Y2=0
cc_169 N_A_27_112#_c_159_n N_A_334_368#_c_351_n 3.03895e-19 $X=1.03 $Y=1.765
+ $X2=0 $Y2=0
cc_170 N_A_27_112#_c_159_n N_A_334_368#_c_352_n 0.00142359f $X=1.03 $Y=1.765
+ $X2=0 $Y2=0
cc_171 N_A_27_112#_M1012_g N_A_334_368#_c_337_n 5.09056e-19 $X=1.075 $Y=0.74
+ $X2=0 $Y2=0
cc_172 N_A_27_112#_M1012_g N_A_334_368#_c_338_n 9.49225e-19 $X=1.075 $Y=0.74
+ $X2=0 $Y2=0
cc_173 N_A_27_112#_c_178_n N_VPWR_M1018_d 0.00921861f $X=0.75 $Y=2.075 $X2=-0.19
+ $Y2=-0.245
cc_174 N_A_27_112#_c_165_n N_VPWR_M1018_d 0.0020968f $X=0.835 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_175 N_A_27_112#_c_159_n N_VPWR_c_526_n 0.0106117f $X=1.03 $Y=1.765 $X2=0
+ $Y2=0
cc_176 N_A_27_112#_c_168_n N_VPWR_c_526_n 0.0124215f $X=0.28 $Y=2.535 $X2=0
+ $Y2=0
cc_177 N_A_27_112#_c_178_n N_VPWR_c_526_n 0.0237523f $X=0.75 $Y=2.075 $X2=0
+ $Y2=0
cc_178 N_A_27_112#_c_168_n N_VPWR_c_536_n 0.00538193f $X=0.28 $Y=2.535 $X2=0
+ $Y2=0
cc_179 N_A_27_112#_c_159_n N_VPWR_c_537_n 0.00445602f $X=1.03 $Y=1.765 $X2=0
+ $Y2=0
cc_180 N_A_27_112#_c_159_n N_VPWR_c_525_n 0.00866521f $X=1.03 $Y=1.765 $X2=0
+ $Y2=0
cc_181 N_A_27_112#_c_168_n N_VPWR_c_525_n 0.00801054f $X=0.28 $Y=2.535 $X2=0
+ $Y2=0
cc_182 N_A_27_112#_c_162_n N_VGND_M1015_d 0.00129688f $X=0.75 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_183 N_A_27_112#_c_164_n N_VGND_M1015_d 0.00373674f $X=0.835 $Y=1.63 $X2=-0.19
+ $Y2=-0.245
cc_184 N_A_27_112#_c_159_n N_VGND_c_744_n 6.47755e-19 $X=1.03 $Y=1.765 $X2=0
+ $Y2=0
cc_185 N_A_27_112#_M1012_g N_VGND_c_744_n 0.00879154f $X=1.075 $Y=0.74 $X2=0
+ $Y2=0
cc_186 N_A_27_112#_c_161_n N_VGND_c_744_n 0.0115116f $X=0.28 $Y=0.835 $X2=0
+ $Y2=0
cc_187 N_A_27_112#_c_162_n N_VGND_c_744_n 0.00997062f $X=0.75 $Y=1.095 $X2=0
+ $Y2=0
cc_188 N_A_27_112#_c_164_n N_VGND_c_744_n 0.0163934f $X=0.835 $Y=1.63 $X2=0
+ $Y2=0
cc_189 N_A_27_112#_c_161_n N_VGND_c_752_n 0.00811255f $X=0.28 $Y=0.835 $X2=0
+ $Y2=0
cc_190 N_A_27_112#_M1012_g N_VGND_c_753_n 0.00434272f $X=1.075 $Y=0.74 $X2=0
+ $Y2=0
cc_191 N_A_27_112#_M1012_g N_VGND_c_765_n 0.00830058f $X=1.075 $Y=0.74 $X2=0
+ $Y2=0
cc_192 N_A_27_112#_c_161_n N_VGND_c_765_n 0.0106114f $X=0.28 $Y=0.835 $X2=0
+ $Y2=0
cc_193 N_A_221_368#_M1022_g N_A_334_368#_M1002_g 0.0264864f $X=2.925 $Y=0.74
+ $X2=0 $Y2=0
cc_194 N_A_221_368#_c_243_n N_A_334_368#_c_343_n 0.0211957f $X=2.94 $Y=1.765
+ $X2=0 $Y2=0
cc_195 N_A_221_368#_c_241_n N_A_334_368#_c_351_n 8.43177e-19 $X=2.04 $Y=1.765
+ $X2=0 $Y2=0
cc_196 N_A_221_368#_c_235_n N_A_334_368#_c_351_n 0.0254944f $X=2.37 $Y=1.465
+ $X2=0 $Y2=0
cc_197 N_A_221_368#_c_245_n N_A_334_368#_c_351_n 0.0152201f $X=1.255 $Y=1.985
+ $X2=0 $Y2=0
cc_198 N_A_221_368#_c_239_n N_A_334_368#_c_351_n 0.00689902f $X=1.95 $Y=1.465
+ $X2=0 $Y2=0
cc_199 N_A_221_368#_c_240_n N_A_334_368#_c_351_n 4.36456e-19 $X=2.925 $Y=1.532
+ $X2=0 $Y2=0
cc_200 N_A_221_368#_c_241_n N_A_334_368#_c_352_n 0.0122589f $X=2.04 $Y=1.765
+ $X2=0 $Y2=0
cc_201 N_A_221_368#_c_242_n N_A_334_368#_c_352_n 6.50051e-19 $X=2.49 $Y=1.765
+ $X2=0 $Y2=0
cc_202 N_A_221_368#_c_245_n N_A_334_368#_c_352_n 0.0834061f $X=1.255 $Y=1.985
+ $X2=0 $Y2=0
cc_203 N_A_221_368#_c_233_n N_A_334_368#_c_337_n 0.0194438f $X=1.29 $Y=0.515
+ $X2=0 $Y2=0
cc_204 N_A_221_368#_c_235_n N_A_334_368#_c_337_n 0.0210833f $X=2.37 $Y=1.465
+ $X2=0 $Y2=0
cc_205 N_A_221_368#_c_239_n N_A_334_368#_c_337_n 0.00582391f $X=1.95 $Y=1.465
+ $X2=0 $Y2=0
cc_206 N_A_221_368#_M1004_g N_A_334_368#_c_338_n 0.00159319f $X=2.065 $Y=0.74
+ $X2=0 $Y2=0
cc_207 N_A_221_368#_c_233_n N_A_334_368#_c_338_n 0.0380854f $X=1.29 $Y=0.515
+ $X2=0 $Y2=0
cc_208 N_A_221_368#_c_241_n N_A_334_368#_c_353_n 0.0121163f $X=2.04 $Y=1.765
+ $X2=0 $Y2=0
cc_209 N_A_221_368#_c_242_n N_A_334_368#_c_353_n 0.013573f $X=2.49 $Y=1.765
+ $X2=0 $Y2=0
cc_210 N_A_221_368#_c_235_n N_A_334_368#_c_353_n 0.0350772f $X=2.37 $Y=1.465
+ $X2=0 $Y2=0
cc_211 N_A_221_368#_c_240_n N_A_334_368#_c_353_n 0.00754501f $X=2.925 $Y=1.532
+ $X2=0 $Y2=0
cc_212 N_A_221_368#_c_241_n N_A_334_368#_c_354_n 6.50051e-19 $X=2.04 $Y=1.765
+ $X2=0 $Y2=0
cc_213 N_A_221_368#_c_242_n N_A_334_368#_c_354_n 0.0117289f $X=2.49 $Y=1.765
+ $X2=0 $Y2=0
cc_214 N_A_221_368#_c_243_n N_A_334_368#_c_354_n 0.0104444f $X=2.94 $Y=1.765
+ $X2=0 $Y2=0
cc_215 N_A_221_368#_c_242_n N_A_334_368#_c_339_n 0.00127309f $X=2.49 $Y=1.765
+ $X2=0 $Y2=0
cc_216 N_A_221_368#_c_243_n N_A_334_368#_c_339_n 0.00141301f $X=2.94 $Y=1.765
+ $X2=0 $Y2=0
cc_217 N_A_221_368#_c_240_n N_A_334_368#_c_339_n 0.00717782f $X=2.925 $Y=1.532
+ $X2=0 $Y2=0
cc_218 N_A_221_368#_c_240_n N_A_334_368#_c_340_n 5.22192e-19 $X=2.925 $Y=1.532
+ $X2=0 $Y2=0
cc_219 N_A_221_368#_c_242_n N_A_334_368#_c_356_n 0.00124523f $X=2.49 $Y=1.765
+ $X2=0 $Y2=0
cc_220 N_A_221_368#_c_243_n N_A_334_368#_c_356_n 0.00187043f $X=2.94 $Y=1.765
+ $X2=0 $Y2=0
cc_221 N_A_221_368#_c_240_n N_A_334_368#_c_356_n 0.00504592f $X=2.925 $Y=1.532
+ $X2=0 $Y2=0
cc_222 N_A_221_368#_M1004_g N_A_334_368#_c_341_n 0.0147157f $X=2.065 $Y=0.74
+ $X2=0 $Y2=0
cc_223 N_A_221_368#_M1013_g N_A_334_368#_c_341_n 0.0214947f $X=2.495 $Y=0.74
+ $X2=0 $Y2=0
cc_224 N_A_221_368#_M1022_g N_A_334_368#_c_341_n 0.0174616f $X=2.925 $Y=0.74
+ $X2=0 $Y2=0
cc_225 N_A_221_368#_c_235_n N_A_334_368#_c_341_n 0.0695695f $X=2.37 $Y=1.465
+ $X2=0 $Y2=0
cc_226 N_A_221_368#_c_239_n N_A_334_368#_c_341_n 0.0013449f $X=1.95 $Y=1.465
+ $X2=0 $Y2=0
cc_227 N_A_221_368#_c_240_n N_A_334_368#_c_341_n 0.0354411f $X=2.925 $Y=1.532
+ $X2=0 $Y2=0
cc_228 N_A_221_368#_c_240_n N_A_334_368#_c_342_n 0.018262f $X=2.925 $Y=1.532
+ $X2=0 $Y2=0
cc_229 N_A_221_368#_c_244_n N_VPWR_c_526_n 0.0242806f $X=1.255 $Y=2.815 $X2=0
+ $Y2=0
cc_230 N_A_221_368#_c_241_n N_VPWR_c_527_n 0.00348001f $X=2.04 $Y=1.765 $X2=0
+ $Y2=0
cc_231 N_A_221_368#_c_242_n N_VPWR_c_527_n 0.00220054f $X=2.49 $Y=1.765 $X2=0
+ $Y2=0
cc_232 N_A_221_368#_c_242_n N_VPWR_c_528_n 0.00445602f $X=2.49 $Y=1.765 $X2=0
+ $Y2=0
cc_233 N_A_221_368#_c_243_n N_VPWR_c_528_n 0.00445602f $X=2.94 $Y=1.765 $X2=0
+ $Y2=0
cc_234 N_A_221_368#_c_243_n N_VPWR_c_529_n 0.00804627f $X=2.94 $Y=1.765 $X2=0
+ $Y2=0
cc_235 N_A_221_368#_c_241_n N_VPWR_c_537_n 0.00445602f $X=2.04 $Y=1.765 $X2=0
+ $Y2=0
cc_236 N_A_221_368#_c_244_n N_VPWR_c_537_n 0.0172711f $X=1.255 $Y=2.815 $X2=0
+ $Y2=0
cc_237 N_A_221_368#_c_241_n N_VPWR_c_525_n 0.00861719f $X=2.04 $Y=1.765 $X2=0
+ $Y2=0
cc_238 N_A_221_368#_c_242_n N_VPWR_c_525_n 0.00856917f $X=2.49 $Y=1.765 $X2=0
+ $Y2=0
cc_239 N_A_221_368#_c_243_n N_VPWR_c_525_n 0.00857432f $X=2.94 $Y=1.765 $X2=0
+ $Y2=0
cc_240 N_A_221_368#_c_244_n N_VPWR_c_525_n 0.0142626f $X=1.255 $Y=2.815 $X2=0
+ $Y2=0
cc_241 N_A_221_368#_M1022_g N_X_c_634_n 8.24855e-19 $X=2.925 $Y=0.74 $X2=0 $Y2=0
cc_242 N_A_221_368#_M1022_g N_X_c_636_n 2.28512e-19 $X=2.925 $Y=0.74 $X2=0 $Y2=0
cc_243 N_A_221_368#_c_233_n N_VGND_c_744_n 0.0193831f $X=1.29 $Y=0.515 $X2=0
+ $Y2=0
cc_244 N_A_221_368#_M1004_g N_VGND_c_745_n 0.0109645f $X=2.065 $Y=0.74 $X2=0
+ $Y2=0
cc_245 N_A_221_368#_M1013_g N_VGND_c_745_n 0.0105568f $X=2.495 $Y=0.74 $X2=0
+ $Y2=0
cc_246 N_A_221_368#_M1022_g N_VGND_c_745_n 0.00138519f $X=2.925 $Y=0.74 $X2=0
+ $Y2=0
cc_247 N_A_221_368#_M1013_g N_VGND_c_746_n 0.00138519f $X=2.495 $Y=0.74 $X2=0
+ $Y2=0
cc_248 N_A_221_368#_M1022_g N_VGND_c_746_n 0.0105635f $X=2.925 $Y=0.74 $X2=0
+ $Y2=0
cc_249 N_A_221_368#_M1004_g N_VGND_c_753_n 0.00383152f $X=2.065 $Y=0.74 $X2=0
+ $Y2=0
cc_250 N_A_221_368#_c_233_n N_VGND_c_753_n 0.0156794f $X=1.29 $Y=0.515 $X2=0
+ $Y2=0
cc_251 N_A_221_368#_M1013_g N_VGND_c_754_n 0.00383152f $X=2.495 $Y=0.74 $X2=0
+ $Y2=0
cc_252 N_A_221_368#_M1022_g N_VGND_c_754_n 0.00383152f $X=2.925 $Y=0.74 $X2=0
+ $Y2=0
cc_253 N_A_221_368#_M1004_g N_VGND_c_765_n 0.00762539f $X=2.065 $Y=0.74 $X2=0
+ $Y2=0
cc_254 N_A_221_368#_M1013_g N_VGND_c_765_n 0.0075754f $X=2.495 $Y=0.74 $X2=0
+ $Y2=0
cc_255 N_A_221_368#_M1022_g N_VGND_c_765_n 0.0075754f $X=2.925 $Y=0.74 $X2=0
+ $Y2=0
cc_256 N_A_221_368#_c_233_n N_VGND_c_765_n 0.0129217f $X=1.29 $Y=0.515 $X2=0
+ $Y2=0
cc_257 N_A_334_368#_c_353_n N_VPWR_M1007_d 0.00197722f $X=2.55 $Y=1.905 $X2=0
+ $Y2=0
cc_258 N_A_334_368#_c_352_n N_VPWR_c_527_n 0.0315168f $X=1.815 $Y=2.815 $X2=0
+ $Y2=0
cc_259 N_A_334_368#_c_353_n N_VPWR_c_527_n 0.0151327f $X=2.55 $Y=1.905 $X2=0
+ $Y2=0
cc_260 N_A_334_368#_c_354_n N_VPWR_c_527_n 0.0315168f $X=2.715 $Y=2.815 $X2=0
+ $Y2=0
cc_261 N_A_334_368#_c_354_n N_VPWR_c_528_n 0.014552f $X=2.715 $Y=2.815 $X2=0
+ $Y2=0
cc_262 N_A_334_368#_c_343_n N_VPWR_c_529_n 0.0164564f $X=3.44 $Y=1.765 $X2=0
+ $Y2=0
cc_263 N_A_334_368#_c_344_n N_VPWR_c_529_n 6.35908e-19 $X=3.94 $Y=1.765 $X2=0
+ $Y2=0
cc_264 N_A_334_368#_c_354_n N_VPWR_c_529_n 0.0379001f $X=2.715 $Y=2.815 $X2=0
+ $Y2=0
cc_265 N_A_334_368#_c_340_n N_VPWR_c_529_n 0.0205825f $X=5.895 $Y=1.465 $X2=0
+ $Y2=0
cc_266 N_A_334_368#_c_356_n N_VPWR_c_529_n 0.00795491f $X=2.715 $Y=1.985 $X2=0
+ $Y2=0
cc_267 N_A_334_368#_c_341_n N_VPWR_c_529_n 0.00631924f $X=2.71 $Y=0.965 $X2=0
+ $Y2=0
cc_268 N_A_334_368#_c_342_n N_VPWR_c_529_n 4.75507e-19 $X=6.635 $Y=1.532 $X2=0
+ $Y2=0
cc_269 N_A_334_368#_c_343_n N_VPWR_c_530_n 0.00413917f $X=3.44 $Y=1.765 $X2=0
+ $Y2=0
cc_270 N_A_334_368#_c_344_n N_VPWR_c_530_n 0.00461464f $X=3.94 $Y=1.765 $X2=0
+ $Y2=0
cc_271 N_A_334_368#_c_344_n N_VPWR_c_531_n 0.00238553f $X=3.94 $Y=1.765 $X2=0
+ $Y2=0
cc_272 N_A_334_368#_c_345_n N_VPWR_c_531_n 0.00234284f $X=4.39 $Y=1.765 $X2=0
+ $Y2=0
cc_273 N_A_334_368#_c_346_n N_VPWR_c_532_n 0.00242236f $X=4.84 $Y=1.765 $X2=0
+ $Y2=0
cc_274 N_A_334_368#_c_347_n N_VPWR_c_532_n 0.00240779f $X=5.295 $Y=1.765 $X2=0
+ $Y2=0
cc_275 N_A_334_368#_c_348_n N_VPWR_c_533_n 0.00219104f $X=5.745 $Y=1.765 $X2=0
+ $Y2=0
cc_276 N_A_334_368#_c_349_n N_VPWR_c_533_n 0.00219104f $X=6.195 $Y=1.765 $X2=0
+ $Y2=0
cc_277 N_A_334_368#_c_350_n N_VPWR_c_535_n 0.00379697f $X=6.645 $Y=1.765 $X2=0
+ $Y2=0
cc_278 N_A_334_368#_c_352_n N_VPWR_c_537_n 0.0145938f $X=1.815 $Y=2.815 $X2=0
+ $Y2=0
cc_279 N_A_334_368#_c_345_n N_VPWR_c_538_n 0.00461464f $X=4.39 $Y=1.765 $X2=0
+ $Y2=0
cc_280 N_A_334_368#_c_346_n N_VPWR_c_538_n 0.00461464f $X=4.84 $Y=1.765 $X2=0
+ $Y2=0
cc_281 N_A_334_368#_c_347_n N_VPWR_c_539_n 0.00461464f $X=5.295 $Y=1.765 $X2=0
+ $Y2=0
cc_282 N_A_334_368#_c_348_n N_VPWR_c_539_n 0.00461464f $X=5.745 $Y=1.765 $X2=0
+ $Y2=0
cc_283 N_A_334_368#_c_349_n N_VPWR_c_540_n 0.00461464f $X=6.195 $Y=1.765 $X2=0
+ $Y2=0
cc_284 N_A_334_368#_c_350_n N_VPWR_c_540_n 0.00461464f $X=6.645 $Y=1.765 $X2=0
+ $Y2=0
cc_285 N_A_334_368#_c_343_n N_VPWR_c_525_n 0.00818187f $X=3.44 $Y=1.765 $X2=0
+ $Y2=0
cc_286 N_A_334_368#_c_344_n N_VPWR_c_525_n 0.00908404f $X=3.94 $Y=1.765 $X2=0
+ $Y2=0
cc_287 N_A_334_368#_c_345_n N_VPWR_c_525_n 0.00908055f $X=4.39 $Y=1.765 $X2=0
+ $Y2=0
cc_288 N_A_334_368#_c_346_n N_VPWR_c_525_n 0.00907879f $X=4.84 $Y=1.765 $X2=0
+ $Y2=0
cc_289 N_A_334_368#_c_347_n N_VPWR_c_525_n 0.00907879f $X=5.295 $Y=1.765 $X2=0
+ $Y2=0
cc_290 N_A_334_368#_c_348_n N_VPWR_c_525_n 0.00907831f $X=5.745 $Y=1.765 $X2=0
+ $Y2=0
cc_291 N_A_334_368#_c_349_n N_VPWR_c_525_n 0.00907831f $X=6.195 $Y=1.765 $X2=0
+ $Y2=0
cc_292 N_A_334_368#_c_350_n N_VPWR_c_525_n 0.0091148f $X=6.645 $Y=1.765 $X2=0
+ $Y2=0
cc_293 N_A_334_368#_c_352_n N_VPWR_c_525_n 0.0120466f $X=1.815 $Y=2.815 $X2=0
+ $Y2=0
cc_294 N_A_334_368#_c_354_n N_VPWR_c_525_n 0.0119791f $X=2.715 $Y=2.815 $X2=0
+ $Y2=0
cc_295 N_A_334_368#_M1002_g N_X_c_634_n 0.00812804f $X=3.425 $Y=0.74 $X2=0 $Y2=0
cc_296 N_A_334_368#_M1005_g N_X_c_634_n 0.00812804f $X=3.855 $Y=0.74 $X2=0 $Y2=0
cc_297 N_A_334_368#_M1006_g N_X_c_634_n 8.24855e-19 $X=4.355 $Y=0.74 $X2=0 $Y2=0
cc_298 N_A_334_368#_c_343_n N_X_c_639_n 0.00527536f $X=3.44 $Y=1.765 $X2=0 $Y2=0
cc_299 N_A_334_368#_c_344_n N_X_c_639_n 4.44808e-19 $X=3.94 $Y=1.765 $X2=0 $Y2=0
cc_300 N_A_334_368#_M1005_g N_X_c_635_n 0.01369f $X=3.855 $Y=0.74 $X2=0 $Y2=0
cc_301 N_A_334_368#_M1006_g N_X_c_635_n 0.0151745f $X=4.355 $Y=0.74 $X2=0 $Y2=0
cc_302 N_A_334_368#_M1010_g N_X_c_635_n 0.0146497f $X=4.785 $Y=0.74 $X2=0 $Y2=0
cc_303 N_A_334_368#_M1011_g N_X_c_635_n 0.0146863f $X=5.215 $Y=0.74 $X2=0 $Y2=0
cc_304 N_A_334_368#_M1019_g N_X_c_635_n 0.0152668f $X=5.705 $Y=0.74 $X2=0 $Y2=0
cc_305 N_A_334_368#_M1023_g N_X_c_635_n 0.0154892f $X=6.205 $Y=0.74 $X2=0 $Y2=0
cc_306 N_A_334_368#_c_340_n N_X_c_635_n 0.168617f $X=5.895 $Y=1.465 $X2=0 $Y2=0
cc_307 N_A_334_368#_c_342_n N_X_c_635_n 0.0159694f $X=6.635 $Y=1.532 $X2=0 $Y2=0
cc_308 N_A_334_368#_M1002_g N_X_c_636_n 0.00418335f $X=3.425 $Y=0.74 $X2=0 $Y2=0
cc_309 N_A_334_368#_M1005_g N_X_c_636_n 0.00115621f $X=3.855 $Y=0.74 $X2=0 $Y2=0
cc_310 N_A_334_368#_c_340_n N_X_c_636_n 0.0276081f $X=5.895 $Y=1.465 $X2=0 $Y2=0
cc_311 N_A_334_368#_c_341_n N_X_c_636_n 0.0121173f $X=2.71 $Y=0.965 $X2=0 $Y2=0
cc_312 N_A_334_368#_c_342_n N_X_c_636_n 0.00232957f $X=6.635 $Y=1.532 $X2=0
+ $Y2=0
cc_313 N_A_334_368#_c_344_n N_X_c_640_n 0.0135845f $X=3.94 $Y=1.765 $X2=0 $Y2=0
cc_314 N_A_334_368#_c_345_n N_X_c_640_n 0.0136118f $X=4.39 $Y=1.765 $X2=0 $Y2=0
cc_315 N_A_334_368#_c_340_n N_X_c_640_n 0.04878f $X=5.895 $Y=1.465 $X2=0 $Y2=0
cc_316 N_A_334_368#_c_342_n N_X_c_640_n 0.00923296f $X=6.635 $Y=1.532 $X2=0
+ $Y2=0
cc_317 N_A_334_368#_c_343_n N_X_c_641_n 0.00151063f $X=3.44 $Y=1.765 $X2=0 $Y2=0
cc_318 N_A_334_368#_c_340_n N_X_c_641_n 0.0223483f $X=5.895 $Y=1.465 $X2=0 $Y2=0
cc_319 N_A_334_368#_c_342_n N_X_c_641_n 0.00682414f $X=6.635 $Y=1.532 $X2=0
+ $Y2=0
cc_320 N_A_334_368#_c_345_n N_X_c_642_n 4.0177e-19 $X=4.39 $Y=1.765 $X2=0 $Y2=0
cc_321 N_A_334_368#_c_346_n N_X_c_642_n 4.03786e-19 $X=4.84 $Y=1.765 $X2=0 $Y2=0
cc_322 N_A_334_368#_c_346_n N_X_c_643_n 0.0136408f $X=4.84 $Y=1.765 $X2=0 $Y2=0
cc_323 N_A_334_368#_c_347_n N_X_c_643_n 0.0136408f $X=5.295 $Y=1.765 $X2=0 $Y2=0
cc_324 N_A_334_368#_c_340_n N_X_c_643_n 0.0469011f $X=5.895 $Y=1.465 $X2=0 $Y2=0
cc_325 N_A_334_368#_c_342_n N_X_c_643_n 0.00882293f $X=6.635 $Y=1.532 $X2=0
+ $Y2=0
cc_326 N_A_334_368#_c_347_n N_X_c_644_n 4.07589e-19 $X=5.295 $Y=1.765 $X2=0
+ $Y2=0
cc_327 N_A_334_368#_c_348_n N_X_c_644_n 4.07589e-19 $X=5.745 $Y=1.765 $X2=0
+ $Y2=0
cc_328 N_A_334_368#_c_348_n N_X_c_645_n 0.0136118f $X=5.745 $Y=1.765 $X2=0 $Y2=0
cc_329 N_A_334_368#_c_349_n N_X_c_645_n 0.0139827f $X=6.195 $Y=1.765 $X2=0 $Y2=0
cc_330 N_A_334_368#_c_340_n N_X_c_645_n 0.0268326f $X=5.895 $Y=1.465 $X2=0 $Y2=0
cc_331 N_A_334_368#_c_342_n N_X_c_645_n 0.00834795f $X=6.635 $Y=1.532 $X2=0
+ $Y2=0
cc_332 N_A_334_368#_M1019_g N_X_c_637_n 8.24855e-19 $X=5.705 $Y=0.74 $X2=0 $Y2=0
cc_333 N_A_334_368#_M1023_g N_X_c_637_n 0.00812804f $X=6.205 $Y=0.74 $X2=0 $Y2=0
cc_334 N_A_334_368#_M1025_g N_X_c_637_n 0.00682285f $X=6.635 $Y=0.74 $X2=0 $Y2=0
cc_335 N_A_334_368#_M1019_g N_X_c_638_n 5.6669e-19 $X=5.705 $Y=0.74 $X2=0 $Y2=0
cc_336 N_A_334_368#_c_349_n N_X_c_638_n 0.00180659f $X=6.195 $Y=1.765 $X2=0
+ $Y2=0
cc_337 N_A_334_368#_M1023_g N_X_c_638_n 0.00530912f $X=6.205 $Y=0.74 $X2=0 $Y2=0
cc_338 N_A_334_368#_M1025_g N_X_c_638_n 0.0195857f $X=6.635 $Y=0.74 $X2=0 $Y2=0
cc_339 N_A_334_368#_c_350_n N_X_c_638_n 0.0102113f $X=6.645 $Y=1.765 $X2=0 $Y2=0
cc_340 N_A_334_368#_c_340_n N_X_c_638_n 0.0213782f $X=5.895 $Y=1.465 $X2=0 $Y2=0
cc_341 N_A_334_368#_c_342_n N_X_c_638_n 0.0489768f $X=6.635 $Y=1.532 $X2=0 $Y2=0
cc_342 N_A_334_368#_c_349_n N_X_c_647_n 4.07589e-19 $X=6.195 $Y=1.765 $X2=0
+ $Y2=0
cc_343 N_A_334_368#_c_350_n N_X_c_647_n 4.07589e-19 $X=6.645 $Y=1.765 $X2=0
+ $Y2=0
cc_344 N_A_334_368#_c_340_n N_X_c_648_n 0.0210833f $X=5.895 $Y=1.465 $X2=0 $Y2=0
cc_345 N_A_334_368#_c_342_n N_X_c_648_n 0.00641554f $X=6.635 $Y=1.532 $X2=0
+ $Y2=0
cc_346 N_A_334_368#_c_340_n N_X_c_649_n 0.02277f $X=5.895 $Y=1.465 $X2=0 $Y2=0
cc_347 N_A_334_368#_c_342_n N_X_c_649_n 0.00674341f $X=6.635 $Y=1.532 $X2=0
+ $Y2=0
cc_348 N_A_334_368#_c_341_n N_VGND_M1004_s 0.00178571f $X=2.71 $Y=0.965 $X2=0
+ $Y2=0
cc_349 N_A_334_368#_c_341_n N_VGND_M1022_s 0.00347359f $X=2.71 $Y=0.965 $X2=0
+ $Y2=0
cc_350 N_A_334_368#_c_338_n N_VGND_c_745_n 0.0136308f $X=1.85 $Y=0.515 $X2=0
+ $Y2=0
cc_351 N_A_334_368#_c_341_n N_VGND_c_745_n 0.0175375f $X=2.71 $Y=0.965 $X2=0
+ $Y2=0
cc_352 N_A_334_368#_M1002_g N_VGND_c_746_n 0.00365073f $X=3.425 $Y=0.74 $X2=0
+ $Y2=0
cc_353 N_A_334_368#_c_340_n N_VGND_c_746_n 0.00611161f $X=5.895 $Y=1.465 $X2=0
+ $Y2=0
cc_354 N_A_334_368#_c_341_n N_VGND_c_746_n 0.00803013f $X=2.71 $Y=0.965 $X2=0
+ $Y2=0
cc_355 N_A_334_368#_M1005_g N_VGND_c_747_n 0.00365073f $X=3.855 $Y=0.74 $X2=0
+ $Y2=0
cc_356 N_A_334_368#_M1006_g N_VGND_c_747_n 0.0105645f $X=4.355 $Y=0.74 $X2=0
+ $Y2=0
cc_357 N_A_334_368#_M1010_g N_VGND_c_747_n 0.00138519f $X=4.785 $Y=0.74 $X2=0
+ $Y2=0
cc_358 N_A_334_368#_M1006_g N_VGND_c_748_n 0.00138519f $X=4.355 $Y=0.74 $X2=0
+ $Y2=0
cc_359 N_A_334_368#_M1010_g N_VGND_c_748_n 0.0105568f $X=4.785 $Y=0.74 $X2=0
+ $Y2=0
cc_360 N_A_334_368#_M1011_g N_VGND_c_748_n 0.0111547f $X=5.215 $Y=0.74 $X2=0
+ $Y2=0
cc_361 N_A_334_368#_M1019_g N_VGND_c_748_n 0.00143792f $X=5.705 $Y=0.74 $X2=0
+ $Y2=0
cc_362 N_A_334_368#_M1011_g N_VGND_c_749_n 0.00143792f $X=5.215 $Y=0.74 $X2=0
+ $Y2=0
cc_363 N_A_334_368#_M1019_g N_VGND_c_749_n 0.0111624f $X=5.705 $Y=0.74 $X2=0
+ $Y2=0
cc_364 N_A_334_368#_M1023_g N_VGND_c_749_n 0.00365073f $X=6.205 $Y=0.74 $X2=0
+ $Y2=0
cc_365 N_A_334_368#_M1025_g N_VGND_c_751_n 0.0178469f $X=6.635 $Y=0.74 $X2=0
+ $Y2=0
cc_366 N_A_334_368#_c_338_n N_VGND_c_753_n 0.011066f $X=1.85 $Y=0.515 $X2=0
+ $Y2=0
cc_367 N_A_334_368#_M1002_g N_VGND_c_755_n 0.00434272f $X=3.425 $Y=0.74 $X2=0
+ $Y2=0
cc_368 N_A_334_368#_M1005_g N_VGND_c_755_n 0.00434272f $X=3.855 $Y=0.74 $X2=0
+ $Y2=0
cc_369 N_A_334_368#_M1006_g N_VGND_c_756_n 0.00383152f $X=4.355 $Y=0.74 $X2=0
+ $Y2=0
cc_370 N_A_334_368#_M1010_g N_VGND_c_756_n 0.00383152f $X=4.785 $Y=0.74 $X2=0
+ $Y2=0
cc_371 N_A_334_368#_M1011_g N_VGND_c_757_n 0.00383152f $X=5.215 $Y=0.74 $X2=0
+ $Y2=0
cc_372 N_A_334_368#_M1019_g N_VGND_c_757_n 0.00383152f $X=5.705 $Y=0.74 $X2=0
+ $Y2=0
cc_373 N_A_334_368#_M1023_g N_VGND_c_758_n 0.00434272f $X=6.205 $Y=0.74 $X2=0
+ $Y2=0
cc_374 N_A_334_368#_M1025_g N_VGND_c_758_n 0.00434272f $X=6.635 $Y=0.74 $X2=0
+ $Y2=0
cc_375 N_A_334_368#_M1002_g N_VGND_c_765_n 0.00820772f $X=3.425 $Y=0.74 $X2=0
+ $Y2=0
cc_376 N_A_334_368#_M1005_g N_VGND_c_765_n 0.00820718f $X=3.855 $Y=0.74 $X2=0
+ $Y2=0
cc_377 N_A_334_368#_M1006_g N_VGND_c_765_n 0.0075754f $X=4.355 $Y=0.74 $X2=0
+ $Y2=0
cc_378 N_A_334_368#_M1010_g N_VGND_c_765_n 0.0075754f $X=4.785 $Y=0.74 $X2=0
+ $Y2=0
cc_379 N_A_334_368#_M1011_g N_VGND_c_765_n 0.00758109f $X=5.215 $Y=0.74 $X2=0
+ $Y2=0
cc_380 N_A_334_368#_M1019_g N_VGND_c_765_n 0.00758109f $X=5.705 $Y=0.74 $X2=0
+ $Y2=0
cc_381 N_A_334_368#_M1023_g N_VGND_c_765_n 0.00820718f $X=6.205 $Y=0.74 $X2=0
+ $Y2=0
cc_382 N_A_334_368#_M1025_g N_VGND_c_765_n 0.00823934f $X=6.635 $Y=0.74 $X2=0
+ $Y2=0
cc_383 N_A_334_368#_c_338_n N_VGND_c_765_n 0.00915947f $X=1.85 $Y=0.515 $X2=0
+ $Y2=0
cc_384 N_VPWR_c_529_n N_X_c_639_n 0.0361347f $X=3.215 $Y=1.985 $X2=0 $Y2=0
cc_385 N_VPWR_c_530_n N_X_c_639_n 0.0117353f $X=4.035 $Y=3.33 $X2=0 $Y2=0
cc_386 N_VPWR_c_531_n N_X_c_639_n 0.00133675f $X=4.165 $Y=2.305 $X2=0 $Y2=0
cc_387 N_VPWR_c_525_n N_X_c_639_n 0.00971347f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_388 N_VPWR_M1003_s N_X_c_640_n 0.00197722f $X=4.015 $Y=1.84 $X2=0 $Y2=0
cc_389 N_VPWR_c_531_n N_X_c_640_n 0.0151327f $X=4.165 $Y=2.305 $X2=0 $Y2=0
cc_390 N_VPWR_c_529_n N_X_c_641_n 0.00611657f $X=3.215 $Y=1.985 $X2=0 $Y2=0
cc_391 N_VPWR_c_531_n N_X_c_642_n 0.00133086f $X=4.165 $Y=2.305 $X2=0 $Y2=0
cc_392 N_VPWR_c_532_n N_X_c_642_n 0.00143844f $X=5.065 $Y=2.305 $X2=0 $Y2=0
cc_393 N_VPWR_c_538_n N_X_c_642_n 0.011066f $X=4.93 $Y=3.33 $X2=0 $Y2=0
cc_394 N_VPWR_c_525_n N_X_c_642_n 0.00915947f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_395 N_VPWR_M1009_s N_X_c_643_n 0.00203037f $X=4.915 $Y=1.84 $X2=0 $Y2=0
cc_396 N_VPWR_c_532_n N_X_c_643_n 0.0155395f $X=5.065 $Y=2.305 $X2=0 $Y2=0
cc_397 N_VPWR_c_532_n N_X_c_644_n 0.001475f $X=5.065 $Y=2.305 $X2=0 $Y2=0
cc_398 N_VPWR_c_533_n N_X_c_644_n 0.00147295f $X=5.97 $Y=2.305 $X2=0 $Y2=0
cc_399 N_VPWR_c_539_n N_X_c_644_n 0.0119584f $X=5.835 $Y=3.33 $X2=0 $Y2=0
cc_400 N_VPWR_c_525_n N_X_c_644_n 0.00989813f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_401 N_VPWR_M1017_s N_X_c_645_n 0.00197722f $X=5.82 $Y=1.84 $X2=0 $Y2=0
cc_402 N_VPWR_c_533_n N_X_c_645_n 0.0151327f $X=5.97 $Y=2.305 $X2=0 $Y2=0
cc_403 N_VPWR_c_535_n N_X_c_638_n 0.0254744f $X=6.875 $Y=2.115 $X2=0 $Y2=0
cc_404 N_VPWR_c_533_n N_X_c_647_n 0.00147295f $X=5.97 $Y=2.305 $X2=0 $Y2=0
cc_405 N_VPWR_c_535_n N_X_c_647_n 0.00148667f $X=6.875 $Y=2.115 $X2=0 $Y2=0
cc_406 N_VPWR_c_540_n N_X_c_647_n 0.0119584f $X=6.735 $Y=3.33 $X2=0 $Y2=0
cc_407 N_VPWR_c_525_n N_X_c_647_n 0.00989813f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_408 N_X_c_635_n N_VGND_M1005_s 0.00253871f $X=6.255 $Y=1.005 $X2=0 $Y2=0
cc_409 N_X_c_635_n N_VGND_M1010_s 0.00178571f $X=6.255 $Y=1.005 $X2=0 $Y2=0
cc_410 N_X_c_635_n N_VGND_M1019_s 0.00253871f $X=6.255 $Y=1.005 $X2=0 $Y2=0
cc_411 N_X_c_634_n N_VGND_c_746_n 0.0142986f $X=3.64 $Y=0.515 $X2=0 $Y2=0
cc_412 N_X_c_634_n N_VGND_c_747_n 0.0142986f $X=3.64 $Y=0.515 $X2=0 $Y2=0
cc_413 N_X_c_635_n N_VGND_c_747_n 0.0215485f $X=6.255 $Y=1.005 $X2=0 $Y2=0
cc_414 N_X_c_635_n N_VGND_c_748_n 0.0175375f $X=6.255 $Y=1.005 $X2=0 $Y2=0
cc_415 N_X_c_635_n N_VGND_c_749_n 0.0215485f $X=6.255 $Y=1.005 $X2=0 $Y2=0
cc_416 N_X_c_637_n N_VGND_c_749_n 0.0142986f $X=6.42 $Y=0.515 $X2=0 $Y2=0
cc_417 N_X_c_637_n N_VGND_c_751_n 0.0206398f $X=6.42 $Y=0.515 $X2=0 $Y2=0
cc_418 N_X_c_638_n N_VGND_c_751_n 0.0284003f $X=6.42 $Y=1.97 $X2=0 $Y2=0
cc_419 N_X_c_634_n N_VGND_c_755_n 0.0144922f $X=3.64 $Y=0.515 $X2=0 $Y2=0
cc_420 N_X_c_637_n N_VGND_c_758_n 0.0144922f $X=6.42 $Y=0.515 $X2=0 $Y2=0
cc_421 N_X_c_634_n N_VGND_c_765_n 0.0118826f $X=3.64 $Y=0.515 $X2=0 $Y2=0
cc_422 N_X_c_637_n N_VGND_c_765_n 0.0118826f $X=6.42 $Y=0.515 $X2=0 $Y2=0
