* NGSPICE file created from sky130_fd_sc_ls__dlxtn_1.ext - technology: sky130A

.subckt sky130_fd_sc_ls__dlxtn_1 D GATE_N VGND VNB VPB VPWR Q
M1000 a_812_508# a_217_419# a_669_392# VPB phighvt w=420000u l=150000u
+  ad=1.134e+11p pd=1.38e+06u as=5.128e+11p ps=3.13e+06u
M1001 Q a_863_441# VGND VNB nshort w=740000u l=150000u
+  ad=2.146e+11p pd=2.06e+06u as=1.31878e+12p ps=1.016e+07u
M1002 VGND a_217_419# a_369_392# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1003 VPWR a_217_419# a_369_392# VPB phighvt w=840000u l=150000u
+  ad=1.57875e+12p pd=1.174e+07u as=2.478e+11p ps=2.27e+06u
M1004 VGND D a_27_115# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1005 a_871_139# a_369_392# a_669_392# VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=2.786e+11p ps=2.52e+06u
M1006 a_217_419# GATE_N VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1007 a_863_441# a_669_392# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.95e+11p pd=2.59e+06u as=0p ps=0u
M1008 a_669_392# a_369_392# a_585_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1009 Q a_863_441# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=0p ps=0u
M1010 VPWR D a_27_115# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=2.478e+11p ps=2.27e+06u
M1011 a_217_419# GATE_N VPWR VPB phighvt w=840000u l=150000u
+  ad=3.192e+11p pd=2.44e+06u as=0p ps=0u
M1012 a_585_392# a_27_115# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND a_863_441# a_871_139# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_863_441# a_669_392# VGND VNB nshort w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=0p ps=0u
M1015 a_655_79# a_27_115# VGND VNB nshort w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1016 a_669_392# a_217_419# a_655_79# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR a_863_441# a_812_508# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

