* File: sky130_fd_sc_ls__sdfxtp_1.pex.spice
* Created: Wed Sep  2 11:28:27 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__SDFXTP_1%A_35_74# 1 2 9 11 13 14 16 19 21 25 26 31
+ 38 39
c96 39 0 1.8681e-19 $X=0.825 $Y=1.825
c97 38 0 1.35641e-19 $X=0.66 $Y=1.69
r98 37 39 10.1561 $w=5.98e-07 $l=1.65e-07 $layer=LI1_cond $X=0.66 $Y=1.825
+ $X2=0.825 $Y2=1.825
r99 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.66
+ $Y=1.69 $X2=0.66 $Y2=1.69
r100 35 37 6.77778 $w=5.98e-07 $l=3.4e-07 $layer=LI1_cond $X=0.32 $Y=1.825
+ $X2=0.66 $Y2=1.825
r101 33 35 2.9902 $w=5.98e-07 $l=1.5e-07 $layer=LI1_cond $X=0.17 $Y=1.825
+ $X2=0.32 $Y2=1.825
r102 28 31 3.97394 $w=4.33e-07 $l=1.5e-07 $layer=LI1_cond $X=0.17 $Y=0.567
+ $X2=0.32 $Y2=0.567
r103 25 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.03
+ $Y=1.635 $X2=2.03 $Y2=1.635
r104 23 25 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=2.03 $Y=1.955
+ $X2=2.03 $Y2=1.635
r105 21 23 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.865 $Y=2.04
+ $X2=2.03 $Y2=1.955
r106 21 39 67.8503 $w=1.68e-07 $l=1.04e-06 $layer=LI1_cond $X=1.865 $Y=2.04
+ $X2=0.825 $Y2=2.04
r107 17 35 2.16985 $w=4.7e-07 $l=3e-07 $layer=LI1_cond $X=0.32 $Y=2.125 $X2=0.32
+ $Y2=1.825
r108 17 19 8.65248 $w=4.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.32 $Y=2.125
+ $X2=0.32 $Y2=2.465
r109 16 33 8.31678 $w=1.7e-07 $l=3e-07 $layer=LI1_cond $X=0.17 $Y=1.525 $X2=0.17
+ $Y2=1.825
r110 15 28 6.29128 $w=1.7e-07 $l=2.18e-07 $layer=LI1_cond $X=0.17 $Y=0.785
+ $X2=0.17 $Y2=0.567
r111 15 16 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=0.17 $Y=0.785
+ $X2=0.17 $Y2=1.525
r112 14 26 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.03 $Y=1.975
+ $X2=2.03 $Y2=1.635
r113 11 14 48.0221 $w=2.71e-07 $l=2.91633e-07 $layer=POLY_cond $X=1.985 $Y=2.245
+ $X2=2.03 $Y2=1.975
r114 11 13 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.985 $Y=2.245
+ $X2=1.985 $Y2=2.64
r115 7 38 74.7592 $w=2.45e-07 $l=4.55082e-07 $layer=POLY_cond $X=1.04 $Y=1.525
+ $X2=0.66 $Y2=1.69
r116 7 9 484.564 $w=1.5e-07 $l=9.45e-07 $layer=POLY_cond $X=1.04 $Y=1.525
+ $X2=1.04 $Y2=0.58
r117 2 19 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.245
+ $Y=2.32 $X2=0.39 $Y2=2.465
r118 1 31 182 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_NDIFF $count=1 $X=0.175
+ $Y=0.37 $X2=0.32 $Y2=0.565
.ends

.subckt PM_SKY130_FD_SC_LS__SDFXTP_1%SCE 2 3 4 5 6 9 11 13 14 16 18 21 22 26 30
+ 31 33 40 43 45
r88 33 45 3.36024 $w=4.73e-07 $l=1.15e-07 $layer=LI1_cond $X=1.2 $Y=1.047
+ $X2=1.315 $Y2=1.047
r89 33 43 4.02225 $w=4.73e-07 $l=1.15e-07 $layer=LI1_cond $X=1.2 $Y=1.047
+ $X2=1.085 $Y2=1.047
r90 31 40 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.085 $Y=1.065
+ $X2=2.085 $Y2=0.9
r91 30 45 23.0489 $w=3.83e-07 $l=7.7e-07 $layer=LI1_cond $X=2.085 $Y=1.092
+ $X2=1.315 $Y2=1.092
r92 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.085
+ $Y=1.065 $X2=2.085 $Y2=1.065
r93 26 37 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.59 $Y=1.12 $X2=0.59
+ $Y2=1.21
r94 26 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.59 $Y=1.12
+ $X2=0.59 $Y2=0.955
r95 25 43 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=0.59 $Y=1.12
+ $X2=1.085 $Y2=1.12
r96 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.59
+ $Y=1.12 $X2=0.59 $Y2=1.12
r97 21 40 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.175 $Y=0.58
+ $X2=2.175 $Y2=0.9
r98 16 18 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.115 $Y=2.245
+ $X2=1.115 $Y2=2.64
r99 15 22 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.69 $Y=2.17
+ $X2=0.615 $Y2=2.17
r100 14 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.04 $Y=2.17
+ $X2=1.115 $Y2=2.245
r101 14 15 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=1.04 $Y=2.17
+ $X2=0.69 $Y2=2.17
r102 11 22 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.615 $Y=2.245
+ $X2=0.615 $Y2=2.17
r103 11 13 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.615 $Y=2.245
+ $X2=0.615 $Y2=2.64
r104 9 36 192.287 $w=1.5e-07 $l=3.75e-07 $layer=POLY_cond $X=0.535 $Y=0.58
+ $X2=0.535 $Y2=0.955
r105 5 22 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.54 $Y=2.17
+ $X2=0.615 $Y2=2.17
r106 5 6 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.54 $Y=2.17
+ $X2=0.255 $Y2=2.17
r107 3 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.425 $Y=1.21
+ $X2=0.59 $Y2=1.21
r108 3 4 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=0.425 $Y=1.21
+ $X2=0.255 $Y2=1.21
r109 2 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.18 $Y=2.095
+ $X2=0.255 $Y2=2.17
r110 1 4 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.18 $Y=1.285
+ $X2=0.255 $Y2=1.21
r111 1 2 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=0.18 $Y=1.285 $X2=0.18
+ $Y2=2.095
.ends

.subckt PM_SKY130_FD_SC_LS__SDFXTP_1%D 3 6 7 9 10 13 14
c42 13 0 1.8681e-19 $X=1.49 $Y=1.62
r43 13 16 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.49 $Y=1.62
+ $X2=1.49 $Y2=1.785
r44 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.49 $Y=1.62
+ $X2=1.49 $Y2=1.455
r45 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.49
+ $Y=1.62 $X2=1.49 $Y2=1.62
r46 10 14 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=1.2 $Y=1.62 $X2=1.49
+ $Y2=1.62
r47 7 9 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.535 $Y=2.245
+ $X2=1.535 $Y2=2.64
r48 6 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.535 $Y=2.155 $X2=1.535
+ $Y2=2.245
r49 6 16 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=1.535 $Y=2.155
+ $X2=1.535 $Y2=1.785
r50 3 15 448.67 $w=1.5e-07 $l=8.75e-07 $layer=POLY_cond $X=1.43 $Y=0.58 $X2=1.43
+ $Y2=1.455
.ends

.subckt PM_SKY130_FD_SC_LS__SDFXTP_1%SCD 1 3 6 10 11 14
c46 6 0 7.17504e-20 $X=2.565 $Y=0.58
r47 11 14 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.57
+ $Y=1.635 $X2=2.57 $Y2=1.635
r48 10 14 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.57 $Y=1.975
+ $X2=2.57 $Y2=1.635
r49 9 14 37.7798 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.57 $Y=1.47
+ $X2=2.57 $Y2=1.635
r50 6 9 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=2.565 $Y=0.58
+ $X2=2.565 $Y2=1.47
r51 1 10 48.0221 $w=2.71e-07 $l=2.91633e-07 $layer=POLY_cond $X=2.525 $Y=2.245
+ $X2=2.57 $Y2=1.975
r52 1 3 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.525 $Y=2.245
+ $X2=2.525 $Y2=2.64
.ends

.subckt PM_SKY130_FD_SC_LS__SDFXTP_1%CLK 1 3 4 6 7
c40 7 0 7.17504e-20 $X=3.6 $Y=1.295
r41 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.415
+ $Y=1.385 $X2=3.415 $Y2=1.385
r42 7 11 5.76222 $w=3.68e-07 $l=1.85e-07 $layer=LI1_cond $X=3.6 $Y=1.365
+ $X2=3.415 $Y2=1.365
r43 4 10 66.8274 $w=3.74e-07 $l=4.06571e-07 $layer=POLY_cond $X=3.235 $Y=1.765
+ $X2=3.29 $Y2=1.385
r44 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.235 $Y=1.765
+ $X2=3.235 $Y2=2.4
r45 1 10 39.1188 $w=3.74e-07 $l=2.85832e-07 $layer=POLY_cond $X=3.075 $Y=1.22
+ $X2=3.29 $Y2=1.385
r46 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.075 $Y=1.22 $X2=3.075
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__SDFXTP_1%A_828_74# 1 2 7 9 10 12 15 17 18 20 21 24
+ 26 27 29 30 33 36 37 39 42 43 44 47 51 52 57 58 60 61 63 64 65 78
c203 64 0 7.65965e-20 $X=7.57 $Y=1.195
c204 57 0 4.42023e-21 $X=5.12 $Y=2.215
c205 51 0 1.06419e-19 $X=8.47 $Y=1.57
c206 47 0 7.308e-20 $X=8.07 $Y=1.275
c207 33 0 1.68607e-19 $X=5.82 $Y=0.69
c208 29 0 1.77768e-19 $X=5.14 $Y=2.05
c209 18 0 1.30629e-20 $X=8.365 $Y=2.465
c210 17 0 1.24984e-19 $X=8.365 $Y=2.375
r211 64 78 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.57 $Y=1.195
+ $X2=7.57 $Y2=1.03
r212 63 66 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=7.65 $Y=1.195 $X2=7.65
+ $Y2=1.275
r213 63 65 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.65 $Y=1.195
+ $X2=7.65 $Y2=1.03
r214 63 64 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.57
+ $Y=1.195 $X2=7.57 $Y2=1.195
r215 58 72 54.032 $w=2.81e-07 $l=3.15e-07 $layer=POLY_cond $X=5.12 $Y=2.257
+ $X2=5.435 $Y2=2.257
r216 57 58 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.12
+ $Y=2.215 $X2=5.12 $Y2=2.215
r217 55 57 17.8075 $w=3.22e-07 $l=4.7e-07 $layer=LI1_cond $X=4.65 $Y=2.1
+ $X2=5.12 $Y2=2.1
r218 51 52 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.47
+ $Y=1.57 $X2=8.47 $Y2=1.57
r219 49 51 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=8.43 $Y=1.49 $X2=8.43
+ $Y2=1.57
r220 48 66 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.815 $Y=1.275
+ $X2=7.65 $Y2=1.275
r221 47 49 20.9966 $w=2.15e-07 $l=3.91152e-07 $layer=LI1_cond $X=8.07 $Y=1.275
+ $X2=8.43 $Y2=1.34
r222 47 48 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=8.07 $Y=1.275
+ $X2=7.815 $Y2=1.275
r223 45 65 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=7.73 $Y=0.425
+ $X2=7.73 $Y2=1.03
r224 43 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.645 $Y=0.34
+ $X2=7.73 $Y2=0.425
r225 43 44 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.645 $Y=0.34
+ $X2=6.975 $Y2=0.34
r226 41 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.89 $Y=0.425
+ $X2=6.975 $Y2=0.34
r227 41 42 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=6.89 $Y=0.425
+ $X2=6.89 $Y2=0.69
r228 40 61 2.11342 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.985 $Y=0.775
+ $X2=5.86 $Y2=0.775
r229 39 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.805 $Y=0.775
+ $X2=6.89 $Y2=0.69
r230 39 40 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=6.805 $Y=0.775
+ $X2=5.985 $Y2=0.775
r231 37 73 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=5.82 $Y=1.195
+ $X2=5.695 $Y2=1.195
r232 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.82
+ $Y=1.195 $X2=5.82 $Y2=1.195
r233 34 61 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=5.86 $Y=0.86 $X2=5.86
+ $Y2=0.775
r234 34 36 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=5.86 $Y=0.86
+ $X2=5.86 $Y2=1.195
r235 33 61 4.3182 $w=2.1e-07 $l=1.03078e-07 $layer=LI1_cond $X=5.82 $Y=0.69
+ $X2=5.86 $Y2=0.775
r236 32 33 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=5.82 $Y=0.425
+ $X2=5.82 $Y2=0.69
r237 31 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.225 $Y=0.34
+ $X2=5.14 $Y2=0.34
r238 30 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.735 $Y=0.34
+ $X2=5.82 $Y2=0.425
r239 30 31 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=5.735 $Y=0.34
+ $X2=5.225 $Y2=0.34
r240 29 57 0.757764 $w=3.22e-07 $l=2e-08 $layer=LI1_cond $X=5.14 $Y=2.1 $X2=5.12
+ $Y2=2.1
r241 28 60 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.14 $Y=0.425
+ $X2=5.14 $Y2=0.34
r242 28 29 106.016 $w=1.68e-07 $l=1.625e-06 $layer=LI1_cond $X=5.14 $Y=0.425
+ $X2=5.14 $Y2=2.05
r243 26 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.055 $Y=0.34
+ $X2=5.14 $Y2=0.34
r244 26 27 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=5.055 $Y=0.34
+ $X2=4.445 $Y2=0.34
r245 22 27 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.32 $Y=0.425
+ $X2=4.445 $Y2=0.34
r246 22 24 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=4.32 $Y=0.425
+ $X2=4.32 $Y2=0.515
r247 21 52 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=8.47 $Y=1.91
+ $X2=8.47 $Y2=1.57
r248 18 20 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=8.365 $Y=2.465
+ $X2=8.365 $Y2=2.75
r249 17 18 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=8.365 $Y=2.375
+ $X2=8.365 $Y2=2.465
r250 16 21 44.3718 $w=2.77e-07 $l=3.02985e-07 $layer=POLY_cond $X=8.365 $Y=2.165
+ $X2=8.47 $Y2=1.91
r251 16 17 81.629 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=8.365 $Y=2.165
+ $X2=8.365 $Y2=2.375
r252 15 78 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=7.525 $Y=0.645
+ $X2=7.525 $Y2=1.03
r253 10 73 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.695 $Y=1.03
+ $X2=5.695 $Y2=1.195
r254 10 12 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=5.695 $Y=1.03
+ $X2=5.695 $Y2=0.71
r255 7 72 17.4353 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=5.435 $Y=2.465
+ $X2=5.435 $Y2=2.257
r256 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=5.435 $Y=2.465
+ $X2=5.435 $Y2=2.75
r257 2 55 600 $w=1.7e-07 $l=2.43721e-07 $layer=licon1_PDIFF $count=1 $X=4.5
+ $Y=1.84 $X2=4.65 $Y2=2.02
r258 1 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.14
+ $Y=0.37 $X2=4.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__SDFXTP_1%A_630_74# 1 2 9 11 13 15 16 20 22 27 28 30
+ 31 33 35 36 37 38 40 41 43 48 50 54 55 58 61 62 64 65 66 68 69 72 74 79 80 87
c212 68 0 1.7275e-19 $X=7.63 $Y=2.52
c213 66 0 1.30859e-19 $X=6.215 $Y=2.605
c214 43 0 1.89404e-19 $X=5.015 $Y=1.555
c215 36 0 1.41929e-19 $X=8.29 $Y=1.09
c216 31 0 3.01141e-19 $X=7.66 $Y=2.045
c217 28 0 7.56861e-20 $X=5.935 $Y=2.465
c218 27 0 4.42023e-21 $X=5.935 $Y=2.375
c219 20 0 1.68607e-19 $X=5.015 $Y=0.71
c220 13 0 1.77768e-19 $X=4.425 $Y=1.765
r221 80 88 11.9702 $w=3.02e-07 $l=7.5e-08 $layer=POLY_cond $X=7.735 $Y=1.822
+ $X2=7.66 $Y2=1.822
r222 79 80 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.735
+ $Y=1.765 $X2=7.735 $Y2=1.765
r223 76 79 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=7.63 $Y=1.765
+ $X2=7.735 $Y2=1.765
r224 72 87 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.9 $Y=2.035
+ $X2=5.9 $Y2=2.2
r225 71 74 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=5.9 $Y=2.035
+ $X2=6.13 $Y2=2.035
r226 71 72 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.9
+ $Y=2.035 $X2=5.9 $Y2=2.035
r227 67 76 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.63 $Y=1.93
+ $X2=7.63 $Y2=1.765
r228 67 68 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=7.63 $Y=1.93
+ $X2=7.63 $Y2=2.52
r229 65 68 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.545 $Y=2.605
+ $X2=7.63 $Y2=2.52
r230 65 66 86.7701 $w=1.68e-07 $l=1.33e-06 $layer=LI1_cond $X=7.545 $Y=2.605
+ $X2=6.215 $Y2=2.605
r231 64 66 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.13 $Y=2.52
+ $X2=6.215 $Y2=2.605
r232 63 74 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.13 $Y=2.2
+ $X2=6.13 $Y2=2.035
r233 63 64 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=6.13 $Y=2.2 $X2=6.13
+ $Y2=2.52
r234 62 84 14.8382 $w=3.5e-07 $l=9e-08 $layer=POLY_cond $X=3.965 $Y=1.465
+ $X2=3.965 $Y2=1.555
r235 62 83 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.965 $Y=1.465
+ $X2=3.965 $Y2=1.3
r236 61 62 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.955
+ $Y=1.465 $X2=3.955 $Y2=1.465
r237 59 61 19.6864 $w=1.98e-07 $l=3.55e-07 $layer=LI1_cond $X=3.955 $Y=1.82
+ $X2=3.955 $Y2=1.465
r238 58 69 5.8268 $w=1.98e-07 $l=1e-07 $layer=LI1_cond $X=3.955 $Y=1.4 $X2=3.955
+ $Y2=1.3
r239 58 61 3.60455 $w=1.98e-07 $l=6.5e-08 $layer=LI1_cond $X=3.955 $Y=1.4
+ $X2=3.955 $Y2=1.465
r240 56 69 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=3.94 $Y=0.96
+ $X2=3.94 $Y2=1.3
r241 54 56 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.855 $Y=0.875
+ $X2=3.94 $Y2=0.96
r242 54 55 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=3.855 $Y=0.875
+ $X2=3.455 $Y2=0.875
r243 50 59 7.29955 $w=3.2e-07 $l=2.03961e-07 $layer=LI1_cond $X=3.855 $Y=1.98
+ $X2=3.955 $Y2=1.82
r244 50 52 14.2255 $w=3.18e-07 $l=3.95e-07 $layer=LI1_cond $X=3.855 $Y=1.98
+ $X2=3.46 $Y2=1.98
r245 46 55 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.29 $Y=0.79
+ $X2=3.455 $Y2=0.875
r246 46 48 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.29 $Y=0.79
+ $X2=3.29 $Y2=0.515
r247 43 44 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=5.015 $Y=1.555
+ $X2=5.015 $Y2=1.765
r248 38 40 98.0067 $w=1.5e-07 $l=3.05e-07 $layer=POLY_cond $X=8.365 $Y=1.015
+ $X2=8.365 $Y2=0.71
r249 36 38 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.29 $Y=1.09
+ $X2=8.365 $Y2=1.015
r250 36 37 99.9894 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=8.29 $Y=1.09
+ $X2=8.095 $Y2=1.09
r251 35 80 45.4868 $w=3.02e-07 $l=3.80125e-07 $layer=POLY_cond $X=8.02 $Y=1.6
+ $X2=7.735 $Y2=1.822
r252 34 37 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.02 $Y=1.165
+ $X2=8.095 $Y2=1.09
r253 34 35 223.053 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.02 $Y=1.165
+ $X2=8.02 $Y2=1.6
r254 31 88 19.1248 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=7.66 $Y=2.045
+ $X2=7.66 $Y2=1.822
r255 31 33 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=7.66 $Y=2.045
+ $X2=7.66 $Y2=2.54
r256 28 30 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=5.935 $Y=2.465
+ $X2=5.935 $Y2=2.75
r257 27 28 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.935 $Y=2.375
+ $X2=5.935 $Y2=2.465
r258 27 87 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=5.935 $Y=2.375
+ $X2=5.935 $Y2=2.2
r259 24 72 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=5.9 $Y=1.84
+ $X2=5.9 $Y2=2.035
r260 23 44 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.09 $Y=1.765
+ $X2=5.015 $Y2=1.765
r261 22 24 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=5.735 $Y=1.765
+ $X2=5.9 $Y2=1.84
r262 22 23 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=5.735 $Y=1.765
+ $X2=5.09 $Y2=1.765
r263 18 43 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.015 $Y=1.48
+ $X2=5.015 $Y2=1.555
r264 18 20 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=5.015 $Y=1.48
+ $X2=5.015 $Y2=0.71
r265 17 41 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.515 $Y=1.555
+ $X2=4.425 $Y2=1.555
r266 16 43 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.94 $Y=1.555
+ $X2=5.015 $Y2=1.555
r267 16 17 217.926 $w=1.5e-07 $l=4.25e-07 $layer=POLY_cond $X=4.94 $Y=1.555
+ $X2=4.515 $Y2=1.555
r268 13 41 83.7788 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=4.425 $Y=1.765
+ $X2=4.425 $Y2=1.555
r269 13 15 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.425 $Y=1.765
+ $X2=4.425 $Y2=2.4
r270 12 84 22.6286 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=4.14 $Y=1.555
+ $X2=3.965 $Y2=1.555
r271 11 41 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.335 $Y=1.555
+ $X2=4.425 $Y2=1.555
r272 11 12 99.9894 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=4.335 $Y=1.555
+ $X2=4.14 $Y2=1.555
r273 9 83 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.065 $Y=0.74
+ $X2=4.065 $Y2=1.3
r274 2 52 600 $w=1.7e-07 $l=2.43721e-07 $layer=licon1_PDIFF $count=1 $X=3.31
+ $Y=1.84 $X2=3.46 $Y2=2.02
r275 1 48 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.15
+ $Y=0.37 $X2=3.29 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__SDFXTP_1%A_1239_74# 1 2 9 10 12 15 16 19 22 26 27 30
+ 33 35
c74 27 0 1.94723e-19 $X=7.195 $Y=2.1
c75 10 0 1.40468e-19 $X=6.335 $Y=2.465
r76 30 32 8.8114 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=7.31 $Y=0.685
+ $X2=7.31 $Y2=0.86
r77 26 27 8.51103 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=7.195 $Y=2.265
+ $X2=7.195 $Y2=2.1
r78 23 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.23 $Y=1.36
+ $X2=7.23 $Y2=1.195
r79 23 27 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=7.23 $Y=1.36
+ $X2=7.23 $Y2=2.1
r80 22 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.23 $Y=1.03
+ $X2=7.23 $Y2=1.195
r81 22 32 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=7.23 $Y=1.03
+ $X2=7.23 $Y2=0.86
r82 19 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.36 $Y=1.195
+ $X2=6.36 $Y2=1.36
r83 19 35 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.36 $Y=1.195
+ $X2=6.36 $Y2=1.03
r84 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.36
+ $Y=1.195 $X2=6.36 $Y2=1.195
r85 16 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.145 $Y=1.195
+ $X2=7.23 $Y2=1.195
r86 16 18 27.4142 $w=3.28e-07 $l=7.85e-07 $layer=LI1_cond $X=7.145 $Y=1.195
+ $X2=6.36 $Y2=1.195
r87 15 36 489.691 $w=1.5e-07 $l=9.55e-07 $layer=POLY_cond $X=6.35 $Y=2.315
+ $X2=6.35 $Y2=1.36
r88 10 15 58.3064 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=6.335 $Y=2.465
+ $X2=6.335 $Y2=2.315
r89 10 12 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.335 $Y=2.465
+ $X2=6.335 $Y2=2.75
r90 9 35 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.27 $Y=0.71 $X2=6.27
+ $Y2=1.03
r91 2 26 600 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_PDIFF $count=1 $X=7.03
+ $Y=2.12 $X2=7.195 $Y2=2.265
r92 1 30 182 $w=1.7e-07 $l=3.80657e-07 $layer=licon1_NDIFF $count=1 $X=7.165
+ $Y=0.37 $X2=7.31 $Y2=0.685
.ends

.subckt PM_SKY130_FD_SC_LS__SDFXTP_1%A_1018_100# 1 2 7 9 12 16 22 24 26 27 28 29
c87 28 0 1.40468e-19 $X=5.635 $Y=2.54
c88 26 0 1.97671e-19 $X=5.48 $Y=1.615
c89 7 0 3.4703e-20 $X=6.955 $Y=2.045
r90 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.81
+ $Y=1.765 $X2=6.81 $Y2=1.765
r91 29 32 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=6.81 $Y=1.615
+ $X2=6.81 $Y2=1.765
r92 27 28 8.63679 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=5.635 $Y=2.37
+ $X2=5.635 $Y2=2.54
r93 25 26 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.565 $Y=1.615
+ $X2=5.48 $Y2=1.615
r94 24 29 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.645 $Y=1.615
+ $X2=6.81 $Y2=1.615
r95 24 25 70.4599 $w=1.68e-07 $l=1.08e-06 $layer=LI1_cond $X=6.645 $Y=1.615
+ $X2=5.565 $Y2=1.615
r96 22 28 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=5.71 $Y=2.75
+ $X2=5.71 $Y2=2.54
r97 18 26 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.48 $Y=1.7 $X2=5.48
+ $Y2=1.615
r98 18 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.48 $Y=1.7 $X2=5.48
+ $Y2=2.37
r99 14 26 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.48 $Y=1.53 $X2=5.48
+ $Y2=1.615
r100 14 16 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=5.48 $Y=1.53
+ $X2=5.48 $Y2=0.765
r101 10 33 40.2632 $w=4.32e-07 $l=2.5446e-07 $layer=POLY_cond $X=7.09 $Y=1.6
+ $X2=6.905 $Y2=1.765
r102 10 12 489.691 $w=1.5e-07 $l=9.55e-07 $layer=POLY_cond $X=7.09 $Y=1.6
+ $X2=7.09 $Y2=0.645
r103 7 33 53.0942 $w=4.32e-07 $l=3.03974e-07 $layer=POLY_cond $X=6.955 $Y=2.045
+ $X2=6.905 $Y2=1.765
r104 7 9 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=6.955 $Y=2.045
+ $X2=6.955 $Y2=2.54
r105 2 22 600 $w=1.7e-07 $l=2.93428e-07 $layer=licon1_PDIFF $count=1 $X=5.51
+ $Y=2.54 $X2=5.71 $Y2=2.75
r106 1 16 182 $w=1.7e-07 $l=5.05421e-07 $layer=licon1_NDIFF $count=1 $X=5.09
+ $Y=0.5 $X2=5.48 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LS__SDFXTP_1%A_1736_74# 1 2 7 9 10 12 14 15 17 20 24 26
+ 27 28 37 39 42 43 51
c85 43 0 1.61732e-19 $X=9.762 $Y=2.1
c86 28 0 4.59464e-20 $X=9.65 $Y=1.195
c87 26 0 4.09155e-20 $X=10.45 $Y=1.485
c88 14 0 7.308e-20 $X=8.95 $Y=2.315
r89 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.08
+ $Y=1.485 $X2=10.08 $Y2=1.485
r90 44 46 8.48441 $w=4.17e-07 $l=2.9e-07 $layer=LI1_cond $X=9.947 $Y=1.195
+ $X2=9.947 $Y2=1.485
r91 42 43 8.4794 $w=3.43e-07 $l=1.65e-07 $layer=LI1_cond $X=9.762 $Y=2.265
+ $X2=9.762 $Y2=2.1
r92 39 46 9.23389 $w=4.17e-07 $l=2.07918e-07 $layer=LI1_cond $X=9.85 $Y=1.65
+ $X2=9.947 $Y2=1.485
r93 39 43 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=9.85 $Y=1.65
+ $X2=9.85 $Y2=2.1
r94 35 44 5.39268 $w=4.17e-07 $l=2.21371e-07 $layer=LI1_cond $X=9.815 $Y=1.03
+ $X2=9.947 $Y2=1.195
r95 35 37 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=9.815 $Y=1.03
+ $X2=9.815 $Y2=0.645
r96 31 51 33.8246 $w=2.85e-07 $l=2e-07 $layer=POLY_cond $X=9.15 $Y=1.187
+ $X2=8.95 $Y2=1.187
r97 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.15
+ $Y=1.195 $X2=9.15 $Y2=1.195
r98 28 44 2.11011 $w=3.3e-07 $l=2.97e-07 $layer=LI1_cond $X=9.65 $Y=1.195
+ $X2=9.947 $Y2=1.195
r99 28 30 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=9.65 $Y=1.195 $X2=9.15
+ $Y2=1.195
r100 26 47 64.6987 $w=3.3e-07 $l=3.7e-07 $layer=POLY_cond $X=10.45 $Y=1.485
+ $X2=10.08 $Y2=1.485
r101 26 27 5.03009 $w=3.3e-07 $l=1.15022e-07 $layer=POLY_cond $X=10.45 $Y=1.485
+ $X2=10.54 $Y2=1.542
r102 22 24 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.785 $Y=2.39
+ $X2=8.95 $Y2=2.39
r103 18 27 37.0704 $w=1.5e-07 $l=2.29377e-07 $layer=POLY_cond $X=10.555 $Y=1.32
+ $X2=10.54 $Y2=1.542
r104 18 20 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=10.555 $Y=1.32
+ $X2=10.555 $Y2=0.76
r105 15 27 37.0704 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=10.54 $Y=1.765
+ $X2=10.54 $Y2=1.542
r106 15 17 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=10.54 $Y=1.765
+ $X2=10.54 $Y2=2.4
r107 14 24 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.95 $Y=2.315
+ $X2=8.95 $Y2=2.39
r108 13 51 17.7656 $w=1.5e-07 $l=1.73e-07 $layer=POLY_cond $X=8.95 $Y=1.36
+ $X2=8.95 $Y2=1.187
r109 13 14 489.691 $w=1.5e-07 $l=9.55e-07 $layer=POLY_cond $X=8.95 $Y=1.36
+ $X2=8.95 $Y2=2.315
r110 10 22 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.785 $Y=2.465
+ $X2=8.785 $Y2=2.39
r111 10 12 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=8.785 $Y=2.465
+ $X2=8.785 $Y2=2.75
r112 7 51 32.9789 $w=2.85e-07 $l=2.67516e-07 $layer=POLY_cond $X=8.755 $Y=1.015
+ $X2=8.95 $Y2=1.187
r113 7 9 98.0067 $w=1.5e-07 $l=3.05e-07 $layer=POLY_cond $X=8.755 $Y=1.015
+ $X2=8.755 $Y2=0.71
r114 2 42 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=9.605
+ $Y=2.12 $X2=9.755 $Y2=2.265
r115 1 37 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=9.675
+ $Y=0.37 $X2=9.815 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_LS__SDFXTP_1%A_1520_74# 1 2 7 9 12 14 16 18 21 23 26 32
+ 34
c86 32 0 7.65965e-20 $X=8.15 $Y=0.71
c87 26 0 4.09155e-20 $X=9.43 $Y=1.765
c88 21 0 9.5983e-20 $X=8.81 $Y=1.6
r89 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.43
+ $Y=1.765 $X2=9.43 $Y2=1.765
r90 24 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.895 $Y=1.765
+ $X2=8.81 $Y2=1.765
r91 24 26 18.6835 $w=3.28e-07 $l=5.35e-07 $layer=LI1_cond $X=8.895 $Y=1.765
+ $X2=9.43 $Y2=1.765
r92 22 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.81 $Y=1.93
+ $X2=8.81 $Y2=1.765
r93 22 23 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=8.81 $Y=1.93
+ $X2=8.81 $Y2=2.245
r94 21 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.81 $Y=1.6 $X2=8.81
+ $Y2=1.765
r95 20 32 25.6433 $w=3.14e-07 $l=8.1037e-07 $layer=LI1_cond $X=8.81 $Y=1.15
+ $X2=8.15 $Y2=0.815
r96 20 21 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=8.81 $Y=1.15
+ $X2=8.81 $Y2=1.6
r97 19 30 3.97288 $w=1.7e-07 $l=1.57321e-07 $layer=LI1_cond $X=8.135 $Y=2.33
+ $X2=8.01 $Y2=2.257
r98 18 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.725 $Y=2.33
+ $X2=8.81 $Y2=2.245
r99 18 19 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=8.725 $Y=2.33
+ $X2=8.135 $Y2=2.33
r100 14 30 3.17028 $w=2.5e-07 $l=1.58e-07 $layer=LI1_cond $X=8.01 $Y=2.415
+ $X2=8.01 $Y2=2.257
r101 14 16 18.4391 $w=2.48e-07 $l=4e-07 $layer=LI1_cond $X=8.01 $Y=2.415
+ $X2=8.01 $Y2=2.815
r102 10 27 38.7839 $w=3.5e-07 $l=2.20624e-07 $layer=POLY_cond $X=9.6 $Y=1.6
+ $X2=9.47 $Y2=1.765
r103 10 12 489.691 $w=1.5e-07 $l=9.55e-07 $layer=POLY_cond $X=9.6 $Y=1.6 $X2=9.6
+ $Y2=0.645
r104 7 27 54.6211 $w=3.5e-07 $l=3.08545e-07 $layer=POLY_cond $X=9.53 $Y=2.045
+ $X2=9.47 $Y2=1.765
r105 7 9 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=9.53 $Y=2.045
+ $X2=9.53 $Y2=2.54
r106 2 30 600 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=1 $X=7.735
+ $Y=2.12 $X2=7.97 $Y2=2.265
r107 2 16 600 $w=1.7e-07 $l=8.03959e-07 $layer=licon1_PDIFF $count=1 $X=7.735
+ $Y=2.12 $X2=7.97 $Y2=2.815
r108 1 32 182 $w=1.7e-07 $l=6.99643e-07 $layer=licon1_NDIFF $count=1 $X=7.6
+ $Y=0.37 $X2=8.15 $Y2=0.71
.ends

.subckt PM_SKY130_FD_SC_LS__SDFXTP_1%VPWR 1 2 3 4 5 6 21 25 29 33 37 41 46 47 49
+ 50 52 53 54 66 70 75 85 86 89 92 95
c121 21 0 1.35641e-19 $X=0.89 $Y=2.465
r122 95 96 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r123 92 93 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r124 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r125 85 86 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r126 83 86 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=10.8 $Y2=3.33
r127 83 96 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=8.88 $Y2=3.33
r128 82 83 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r129 80 95 12.2593 $w=1.7e-07 $l=2.88e-07 $layer=LI1_cond $X=9.42 $Y=3.33
+ $X2=9.132 $Y2=3.33
r130 80 82 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=9.42 $Y=3.33
+ $X2=9.84 $Y2=3.33
r131 79 96 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=8.88 $Y2=3.33
r132 79 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6.48 $Y2=3.33
r133 78 79 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r134 76 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.81 $Y=3.33
+ $X2=6.645 $Y2=3.33
r135 76 78 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=6.81 $Y=3.33
+ $X2=6.96 $Y2=3.33
r136 75 95 12.2593 $w=1.7e-07 $l=2.87e-07 $layer=LI1_cond $X=8.845 $Y=3.33
+ $X2=9.132 $Y2=3.33
r137 75 78 122.979 $w=1.68e-07 $l=1.885e-06 $layer=LI1_cond $X=8.845 $Y=3.33
+ $X2=6.96 $Y2=3.33
r138 74 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r139 73 74 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r140 71 89 11.4275 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=4.365 $Y=3.33
+ $X2=4.11 $Y2=3.33
r141 71 73 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=4.365 $Y=3.33
+ $X2=4.56 $Y2=3.33
r142 70 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.48 $Y=3.33
+ $X2=6.645 $Y2=3.33
r143 70 73 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=6.48 $Y=3.33
+ $X2=4.56 $Y2=3.33
r144 69 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r145 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r146 66 89 11.4275 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=3.855 $Y=3.33
+ $X2=4.11 $Y2=3.33
r147 66 68 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=3.855 $Y=3.33
+ $X2=3.6 $Y2=3.33
r148 65 69 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r149 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r150 62 65 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r151 61 64 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r152 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r153 58 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r154 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r155 54 93 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6.48 $Y2=3.33
r156 54 74 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=4.56 $Y2=3.33
r157 52 82 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=10.15 $Y=3.33
+ $X2=9.84 $Y2=3.33
r158 52 53 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.15 $Y=3.33
+ $X2=10.275 $Y2=3.33
r159 51 85 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=10.4 $Y=3.33 $X2=10.8
+ $Y2=3.33
r160 51 53 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.4 $Y=3.33
+ $X2=10.275 $Y2=3.33
r161 49 64 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=2.67 $Y=3.33 $X2=2.64
+ $Y2=3.33
r162 49 50 11.3601 $w=1.7e-07 $l=2.52e-07 $layer=LI1_cond $X=2.67 $Y=3.33
+ $X2=2.922 $Y2=3.33
r163 48 68 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=3.175 $Y=3.33
+ $X2=3.6 $Y2=3.33
r164 48 50 11.3601 $w=1.7e-07 $l=2.53e-07 $layer=LI1_cond $X=3.175 $Y=3.33
+ $X2=2.922 $Y2=3.33
r165 46 57 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=0.725 $Y=3.33
+ $X2=0.72 $Y2=3.33
r166 46 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.725 $Y=3.33
+ $X2=0.89 $Y2=3.33
r167 45 61 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=1.055 $Y=3.33
+ $X2=1.2 $Y2=3.33
r168 45 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.055 $Y=3.33
+ $X2=0.89 $Y2=3.33
r169 41 44 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=10.275 $Y=1.985
+ $X2=10.275 $Y2=2.815
r170 39 53 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=10.275 $Y=3.245
+ $X2=10.275 $Y2=3.33
r171 39 44 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=10.275 $Y=3.245
+ $X2=10.275 $Y2=2.815
r172 35 95 2.42056 $w=5.75e-07 $l=8.5e-08 $layer=LI1_cond $X=9.132 $Y=3.245
+ $X2=9.132 $Y2=3.33
r173 35 37 8.94459 $w=5.73e-07 $l=4.3e-07 $layer=LI1_cond $X=9.132 $Y=3.245
+ $X2=9.132 $Y2=2.815
r174 31 92 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.645 $Y=3.245
+ $X2=6.645 $Y2=3.33
r175 31 33 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=6.645 $Y=3.245
+ $X2=6.645 $Y2=3.025
r176 27 89 2.12513 $w=5.1e-07 $l=8.5e-08 $layer=LI1_cond $X=4.11 $Y=3.245
+ $X2=4.11 $Y2=3.33
r177 27 29 10.0846 $w=5.08e-07 $l=4.3e-07 $layer=LI1_cond $X=4.11 $Y=3.245
+ $X2=4.11 $Y2=2.815
r178 23 50 2.09999 $w=5.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.922 $Y=3.245
+ $X2=2.922 $Y2=3.33
r179 23 25 10.1844 $w=5.03e-07 $l=4.3e-07 $layer=LI1_cond $X=2.922 $Y=3.245
+ $X2=2.922 $Y2=2.815
r180 19 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.89 $Y=3.245
+ $X2=0.89 $Y2=3.33
r181 19 21 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=0.89 $Y=3.245
+ $X2=0.89 $Y2=2.465
r182 6 44 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=10.17
+ $Y=1.84 $X2=10.315 $Y2=2.815
r183 6 41 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=10.17
+ $Y=1.84 $X2=10.315 $Y2=1.985
r184 5 37 600 $w=1.7e-07 $l=3.87137e-07 $layer=licon1_PDIFF $count=1 $X=8.86
+ $Y=2.54 $X2=9.13 $Y2=2.815
r185 4 33 600 $w=1.7e-07 $l=5.90931e-07 $layer=licon1_PDIFF $count=1 $X=6.41
+ $Y=2.54 $X2=6.645 $Y2=3.025
r186 3 29 600 $w=1.7e-07 $l=1.08616e-06 $layer=licon1_PDIFF $count=1 $X=3.875
+ $Y=1.84 $X2=4.11 $Y2=2.815
r187 2 25 600 $w=1.7e-07 $l=6.35157e-07 $layer=licon1_PDIFF $count=1 $X=2.6
+ $Y=2.32 $X2=2.92 $Y2=2.815
r188 1 21 300 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=2 $X=0.69
+ $Y=2.32 $X2=0.89 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LS__SDFXTP_1%A_301_74# 1 2 3 4 13 19 22 23 24 26 27 30
+ 31 32 34 36 37 39 42 43 44 49
c135 39 0 7.56861e-20 $X=5.21 $Y=2.805
c136 31 0 1.89404e-19 $X=4.615 $Y=1.565
c137 30 0 8.2679e-20 $X=4.31 $Y=2.31
r138 46 49 3.34041 $w=3.43e-07 $l=1e-07 $layer=LI1_cond $X=4.7 $Y=0.767 $X2=4.8
+ $Y2=0.767
r139 44 45 16.3723 $w=2.31e-07 $l=3.1e-07 $layer=LI1_cond $X=4.31 $Y=2.435
+ $X2=4.62 $Y2=2.435
r140 37 39 21.555 $w=2.68e-07 $l=5.05e-07 $layer=LI1_cond $X=4.705 $Y=2.845
+ $X2=5.21 $Y2=2.845
r141 35 46 4.88813 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=4.7 $Y=0.94 $X2=4.7
+ $Y2=0.767
r142 35 36 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=4.7 $Y=0.94 $X2=4.7
+ $Y2=1.48
r143 34 37 7.28469 $w=2.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=4.62 $Y=2.71
+ $X2=4.705 $Y2=2.845
r144 33 45 2.5345 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.62 $Y=2.56
+ $X2=4.62 $Y2=2.435
r145 33 34 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=4.62 $Y=2.56
+ $X2=4.62 $Y2=2.71
r146 31 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.615 $Y=1.565
+ $X2=4.7 $Y2=1.48
r147 31 32 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=4.615 $Y=1.565
+ $X2=4.395 $Y2=1.565
r148 30 44 2.5345 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.31 $Y=2.31
+ $X2=4.31 $Y2=2.435
r149 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.31 $Y=1.65
+ $X2=4.395 $Y2=1.565
r150 29 30 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=4.31 $Y=1.65
+ $X2=4.31 $Y2=2.31
r151 28 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.08 $Y=2.395
+ $X2=2.995 $Y2=2.395
r152 27 44 51.8401 $w=2.31e-07 $l=9.84797e-07 $layer=LI1_cond $X=3.345 $Y=2.395
+ $X2=4.31 $Y2=2.435
r153 27 28 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.345 $Y=2.395
+ $X2=3.08 $Y2=2.395
r154 26 43 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.995 $Y=2.31
+ $X2=2.995 $Y2=2.395
r155 25 26 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=2.995 $Y=1.3
+ $X2=2.995 $Y2=2.31
r156 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.91 $Y=1.215
+ $X2=2.995 $Y2=1.3
r157 23 24 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2.91 $Y=1.215
+ $X2=2.59 $Y2=1.215
r158 22 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.505 $Y=1.13
+ $X2=2.59 $Y2=1.215
r159 21 22 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=2.505 $Y=0.73
+ $X2=2.505 $Y2=1.13
r160 20 42 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.925 $Y=2.395
+ $X2=1.76 $Y2=2.395
r161 19 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.91 $Y=2.395
+ $X2=2.995 $Y2=2.395
r162 19 20 64.262 $w=1.68e-07 $l=9.85e-07 $layer=LI1_cond $X=2.91 $Y=2.395
+ $X2=1.925 $Y2=2.395
r163 13 21 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.42 $Y=0.565
+ $X2=2.505 $Y2=0.73
r164 13 15 21.1281 $w=3.28e-07 $l=6.05e-07 $layer=LI1_cond $X=2.42 $Y=0.565
+ $X2=1.815 $Y2=0.565
r165 4 39 600 $w=1.7e-07 $l=3.29621e-07 $layer=licon1_PDIFF $count=1 $X=5.065
+ $Y=2.54 $X2=5.21 $Y2=2.805
r166 3 42 300 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=2 $X=1.61
+ $Y=2.32 $X2=1.76 $Y2=2.475
r167 2 49 182 $w=1.7e-07 $l=3.21481e-07 $layer=licon1_NDIFF $count=1 $X=4.675
+ $Y=0.5 $X2=4.8 $Y2=0.765
r168 1 15 182 $w=1.7e-07 $l=3.95664e-07 $layer=licon1_NDIFF $count=1 $X=1.505
+ $Y=0.37 $X2=1.815 $Y2=0.565
.ends

.subckt PM_SKY130_FD_SC_LS__SDFXTP_1%Q 1 2 7 8 9 10 11 12 13
r13 12 13 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=10.767 $Y=2.405
+ $X2=10.767 $Y2=2.775
r14 11 12 14.4485 $w=3.33e-07 $l=4.2e-07 $layer=LI1_cond $X=10.767 $Y=1.985
+ $X2=10.767 $Y2=2.405
r15 10 11 11.0084 $w=3.33e-07 $l=3.2e-07 $layer=LI1_cond $X=10.767 $Y=1.665
+ $X2=10.767 $Y2=1.985
r16 9 10 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=10.767 $Y=1.295
+ $X2=10.767 $Y2=1.665
r17 8 9 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=10.767 $Y=0.925
+ $X2=10.767 $Y2=1.295
r18 7 8 13.4165 $w=3.33e-07 $l=3.9e-07 $layer=LI1_cond $X=10.767 $Y=0.535
+ $X2=10.767 $Y2=0.925
r19 2 13 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=10.615
+ $Y=1.84 $X2=10.765 $Y2=2.815
r20 2 11 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=10.615
+ $Y=1.84 $X2=10.765 $Y2=1.985
r21 1 7 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.63
+ $Y=0.39 $X2=10.77 $Y2=0.535
.ends

.subckt PM_SKY130_FD_SC_LS__SDFXTP_1%VGND 1 2 3 4 5 6 21 25 29 33 37 41 44 45 47
+ 48 49 51 66 73 78 85 86 89 92 95 100
r124 100 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r125 96 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0 $X2=8.88
+ $Y2=0
r126 95 98 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r127 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r128 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r129 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r130 86 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=10.32 $Y2=0
r131 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=0 $X2=10.8
+ $Y2=0
r132 83 100 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.425 $Y=0
+ $X2=10.3 $Y2=0
r133 83 85 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=10.425 $Y=0
+ $X2=10.8 $Y2=0
r134 82 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=10.32 $Y2=0
r135 82 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0 $X2=9.36
+ $Y2=0
r136 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r137 79 95 13.399 $w=1.7e-07 $l=3.38e-07 $layer=LI1_cond $X=9.48 $Y=0 $X2=9.142
+ $Y2=0
r138 79 81 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=9.48 $Y=0 $X2=9.84
+ $Y2=0
r139 78 100 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.175 $Y=0
+ $X2=10.3 $Y2=0
r140 78 81 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=10.175 $Y=0
+ $X2=9.84 $Y2=0
r141 77 98 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6.96 $Y=0
+ $X2=8.88 $Y2=0
r142 77 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=6.48
+ $Y2=0
r143 76 77 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r144 74 92 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.635 $Y=0 $X2=6.51
+ $Y2=0
r145 74 76 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=6.635 $Y=0
+ $X2=6.96 $Y2=0
r146 73 95 13.399 $w=1.7e-07 $l=3.37e-07 $layer=LI1_cond $X=8.805 $Y=0 $X2=9.142
+ $Y2=0
r147 73 76 120.369 $w=1.68e-07 $l=1.845e-06 $layer=LI1_cond $X=8.805 $Y=0
+ $X2=6.96 $Y2=0
r148 72 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r149 71 72 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6
+ $Y2=0
r150 68 71 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.08 $Y=0 $X2=6
+ $Y2=0
r151 68 69 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r152 66 92 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.385 $Y=0 $X2=6.51
+ $Y2=0
r153 66 71 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=6.385 $Y=0 $X2=6
+ $Y2=0
r154 65 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r155 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r156 62 65 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r157 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r158 59 62 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r159 59 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r160 58 61 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r161 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r162 56 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.915 $Y=0 $X2=0.75
+ $Y2=0
r163 56 58 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.915 $Y=0 $X2=1.2
+ $Y2=0
r164 54 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r165 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r166 51 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.585 $Y=0 $X2=0.75
+ $Y2=0
r167 51 53 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.585 $Y=0 $X2=0.24
+ $Y2=0
r168 49 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r169 49 69 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=5.52 $Y=0
+ $X2=4.08 $Y2=0
r170 47 64 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.685 $Y=0 $X2=3.6
+ $Y2=0
r171 47 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.685 $Y=0 $X2=3.85
+ $Y2=0
r172 46 68 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=4.015 $Y=0 $X2=4.08
+ $Y2=0
r173 46 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.015 $Y=0 $X2=3.85
+ $Y2=0
r174 44 61 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=2.775 $Y=0
+ $X2=2.64 $Y2=0
r175 44 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.775 $Y=0 $X2=2.86
+ $Y2=0
r176 43 64 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=2.945 $Y=0 $X2=3.6
+ $Y2=0
r177 43 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.945 $Y=0 $X2=2.86
+ $Y2=0
r178 39 100 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=10.3 $Y=0.085
+ $X2=10.3 $Y2=0
r179 39 41 20.744 $w=2.48e-07 $l=4.5e-07 $layer=LI1_cond $X=10.3 $Y=0.085
+ $X2=10.3 $Y2=0.535
r180 35 95 2.78459 $w=6.75e-07 $l=8.5e-08 $layer=LI1_cond $X=9.142 $Y=0.085
+ $X2=9.142 $Y2=0
r181 35 37 9.92302 $w=6.73e-07 $l=5.6e-07 $layer=LI1_cond $X=9.142 $Y=0.085
+ $X2=9.142 $Y2=0.645
r182 31 92 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.51 $Y=0.085
+ $X2=6.51 $Y2=0
r183 31 33 12.4464 $w=2.48e-07 $l=2.7e-07 $layer=LI1_cond $X=6.51 $Y=0.085
+ $X2=6.51 $Y2=0.355
r184 27 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.85 $Y=0.085
+ $X2=3.85 $Y2=0
r185 27 29 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=3.85 $Y=0.085
+ $X2=3.85 $Y2=0.525
r186 23 45 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.86 $Y=0.085
+ $X2=2.86 $Y2=0
r187 23 25 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=2.86 $Y=0.085
+ $X2=2.86 $Y2=0.625
r188 19 89 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=0.085
+ $X2=0.75 $Y2=0
r189 19 21 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.75 $Y=0.085
+ $X2=0.75 $Y2=0.565
r190 6 41 91 $w=1.7e-07 $l=1.99687e-07 $layer=licon1_NDIFF $count=2 $X=10.21
+ $Y=0.39 $X2=10.34 $Y2=0.535
r191 5 37 91 $w=1.7e-07 $l=5.52766e-07 $layer=licon1_NDIFF $count=2 $X=8.83
+ $Y=0.5 $X2=9.315 $Y2=0.645
r192 4 33 182 $w=1.7e-07 $l=2.67862e-07 $layer=licon1_NDIFF $count=1 $X=6.345
+ $Y=0.5 $X2=6.55 $Y2=0.355
r193 3 29 182 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=1 $X=3.705
+ $Y=0.37 $X2=3.85 $Y2=0.525
r194 2 25 182 $w=1.7e-07 $l=3.4803e-07 $layer=licon1_NDIFF $count=1 $X=2.64
+ $Y=0.37 $X2=2.86 $Y2=0.625
r195 1 21 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=0.61
+ $Y=0.37 $X2=0.75 $Y2=0.565
.ends

