# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ls__tapvpwrvgnd_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ls__tapvpwrvgnd_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  0.480000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 0.480000 0.085000 ;
        RECT 0.090000  0.085000 0.390000 1.105000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 0.480000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 0.480000 3.415000 ;
        RECT 0.090000 2.205000 0.390000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 0.480000 3.575000 ;
    END
  END VPWR
END sky130_fd_sc_ls__tapvpwrvgnd_1
