* File: sky130_fd_sc_ls__or2b_1.spice
* Created: Fri Aug 28 13:57:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__or2b_1.pex.spice"
.subckt sky130_fd_sc_ls__or2b_1  VNB VPB B_N A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B_N	B_N
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_B_N_M1003_g N_A_27_112#_M1003_s VNB NSHORT L=0.15 W=0.55
+ AD=0.174625 AS=0.3685 PD=1.185 PS=2.44 NRD=0 NRS=0 M=1 R=3.66667 SA=75000.6
+ SB=75002.2 A=0.0825 P=1.4 MULT=1
MM1000 N_A_264_368#_M1000_d N_A_27_112#_M1000_g N_VGND_M1003_d VNB NSHORT L=0.15
+ W=0.55 AD=0.077 AS=0.174625 PD=0.83 PS=1.185 NRD=0 NRS=3.264 M=1 R=3.66667
+ SA=75001.4 SB=75001.4 A=0.0825 P=1.4 MULT=1
MM1001 N_VGND_M1001_d N_A_M1001_g N_A_264_368#_M1000_d VNB NSHORT L=0.15 W=0.55
+ AD=0.164766 AS=0.077 PD=1.12558 PS=0.83 NRD=33.816 NRS=0 M=1 R=3.66667
+ SA=75001.8 SB=75000.9 A=0.0825 P=1.4 MULT=1
MM1007 N_X_M1007_d N_A_264_368#_M1007_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.221684 PD=2.05 PS=1.51442 NRD=0 NRS=23.508 M=1 R=4.93333
+ SA=75002 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1005 N_VPWR_M1005_d N_B_N_M1005_g N_A_27_112#_M1005_s VPB PHIGHVT L=0.15
+ W=0.84 AD=0.2898 AS=0.2478 PD=2.37 PS=2.27 NRD=14.0658 NRS=2.3443 M=1 R=5.6
+ SA=75000.2 SB=75000.3 A=0.126 P=1.98 MULT=1
MM1004 A_353_368# N_A_27_112#_M1004_g N_A_264_368#_M1004_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.295 PD=1.27 PS=2.59 NRD=15.7403 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75001.2 A=0.15 P=2.3 MULT=1
MM1002 N_VPWR_M1002_d N_A_M1002_g A_353_368# VPB PHIGHVT L=0.15 W=1 AD=0.224717
+ AS=0.135 PD=1.46698 PS=1.27 NRD=19.0302 NRS=15.7403 M=1 R=6.66667 SA=75000.6
+ SB=75000.8 A=0.15 P=2.3 MULT=1
MM1006 N_X_M1006_d N_A_264_368#_M1006_g N_VPWR_M1002_d VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.251683 PD=2.83 PS=1.64302 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75001.1 SB=75000.2 A=0.168 P=2.54 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.9564 P=11.2
*
.include "sky130_fd_sc_ls__or2b_1.pxi.spice"
*
.ends
*
*
