* File: sky130_fd_sc_ls__dlrtn_4.pex.spice
* Created: Wed Sep  2 11:03:51 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__DLRTN_4%D 3 5 7 8
r29 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.59
+ $Y=1.615 $X2=0.59 $Y2=1.615
r30 8 12 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=0.72 $Y=1.615
+ $X2=0.59 $Y2=1.615
r31 5 11 57.4383 $w=2.94e-07 $l=3.04893e-07 $layer=POLY_cond $X=0.535 $Y=1.895
+ $X2=0.587 $Y2=1.615
r32 5 7 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.535 $Y=1.895
+ $X2=0.535 $Y2=2.39
r33 1 11 38.5845 $w=2.94e-07 $l=2.05925e-07 $layer=POLY_cond $X=0.495 $Y=1.45
+ $X2=0.587 $Y2=1.615
r34 1 3 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.495 $Y=1.45
+ $X2=0.495 $Y2=0.955
.ends

.subckt PM_SKY130_FD_SC_LS__DLRTN_4%GATE_N 3 5 7 8
r33 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.13
+ $Y=1.615 $X2=1.13 $Y2=1.615
r34 5 11 57.6553 $w=2.91e-07 $l=3.01662e-07 $layer=POLY_cond $X=1.085 $Y=1.895
+ $X2=1.13 $Y2=1.615
r35 5 7 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.085 $Y=1.895
+ $X2=1.085 $Y2=2.39
r36 1 11 38.6072 $w=2.91e-07 $l=1.86145e-07 $layer=POLY_cond $X=1.085 $Y=1.45
+ $X2=1.13 $Y2=1.615
r37 1 3 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=1.085 $Y=1.45
+ $X2=1.085 $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_LS__DLRTN_4%A_232_98# 1 2 7 9 12 16 18 20 22 24 25 30 35
+ 36 39 40 43 44 46 48
c114 7 0 1.26581e-19 $X=2.11 $Y=1.885
r115 46 49 8.6688 $w=4.03e-07 $l=1.65e-07 $layer=LI1_cond $X=1.662 $Y=1.585
+ $X2=1.662 $Y2=1.75
r116 46 48 8.6688 $w=4.03e-07 $l=1.65e-07 $layer=LI1_cond $X=1.662 $Y=1.585
+ $X2=1.662 $Y2=1.42
r117 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.7
+ $Y=1.585 $X2=1.7 $Y2=1.585
r118 44 49 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=1.545 $Y=1.95
+ $X2=1.545 $Y2=1.75
r119 43 44 9.42615 $w=4.83e-07 $l=1.65e-07 $layer=LI1_cond $X=1.387 $Y=2.115
+ $X2=1.387 $Y2=1.95
r120 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.035
+ $Y=2.195 $X2=4.035 $Y2=2.195
r121 37 39 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=4.035 $Y=2.6
+ $X2=4.035 $Y2=2.195
r122 35 37 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.87 $Y=2.685
+ $X2=4.035 $Y2=2.6
r123 35 36 146.139 $w=1.68e-07 $l=2.24e-06 $layer=LI1_cond $X=3.87 $Y=2.685
+ $X2=1.63 $Y2=2.685
r124 31 48 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.545 $Y=1.25
+ $X2=1.545 $Y2=1.42
r125 30 36 9.10402 $w=1.7e-07 $l=2.82319e-07 $layer=LI1_cond $X=1.387 $Y=2.6
+ $X2=1.63 $Y2=2.685
r126 29 43 1.89893 $w=4.83e-07 $l=7.7e-08 $layer=LI1_cond $X=1.387 $Y=2.192
+ $X2=1.387 $Y2=2.115
r127 29 30 10.0619 $w=4.83e-07 $l=4.08e-07 $layer=LI1_cond $X=1.387 $Y=2.192
+ $X2=1.387 $Y2=2.6
r128 25 31 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.46 $Y=1.125
+ $X2=1.545 $Y2=1.25
r129 25 27 5.07075 $w=2.48e-07 $l=1.1e-07 $layer=LI1_cond $X=1.46 $Y=1.125
+ $X2=1.35 $Y2=1.125
r130 23 40 49.8355 $w=3.3e-07 $l=2.85e-07 $layer=POLY_cond $X=3.75 $Y=2.195
+ $X2=4.035 $Y2=2.195
r131 23 24 5.03009 $w=3.3e-07 $l=1.08995e-07 $layer=POLY_cond $X=3.75 $Y=2.195
+ $X2=3.66 $Y2=2.237
r132 22 47 55.9556 $w=3.3e-07 $l=3.2e-07 $layer=POLY_cond $X=2.02 $Y=1.585
+ $X2=1.7 $Y2=1.585
r133 18 24 37.0704 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.66 $Y=2.445
+ $X2=3.66 $Y2=2.237
r134 18 20 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.66 $Y=2.445
+ $X2=3.66 $Y2=2.73
r135 14 24 37.0704 $w=1.5e-07 $l=2.14369e-07 $layer=POLY_cond $X=3.645 $Y=2.03
+ $X2=3.66 $Y2=2.237
r136 14 16 687.106 $w=1.5e-07 $l=1.34e-06 $layer=POLY_cond $X=3.645 $Y=2.03
+ $X2=3.645 $Y2=0.69
r137 10 22 43.2316 $w=1.97e-07 $l=1.85257e-07 $layer=POLY_cond $X=2.18 $Y=1.42
+ $X2=2.137 $Y2=1.585
r138 10 12 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.18 $Y=1.42
+ $X2=2.18 $Y2=0.86
r139 7 22 76.2621 $w=1.97e-07 $l=3.13209e-07 $layer=POLY_cond $X=2.11 $Y=1.885
+ $X2=2.137 $Y2=1.585
r140 7 9 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.11 $Y=1.885
+ $X2=2.11 $Y2=2.38
r141 2 43 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=1.16
+ $Y=1.97 $X2=1.31 $Y2=2.115
r142 1 27 182 $w=1.7e-07 $l=6.83429e-07 $layer=licon1_NDIFF $count=1 $X=1.16
+ $Y=0.49 $X2=1.35 $Y2=1.085
.ends

.subckt PM_SKY130_FD_SC_LS__DLRTN_4%A_27_136# 1 2 7 9 10 12 14 18 23 24 27 30 32
+ 33
c75 27 0 1.26581e-19 $X=2.655 $Y=1.505
c76 7 0 1.51556e-19 $X=2.73 $Y=1.885
r77 32 33 8.60763 $w=3.88e-07 $l=1.65e-07 $layer=LI1_cond $X=0.28 $Y=2.115
+ $X2=0.28 $Y2=1.95
r78 30 33 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=0.17 $Y=1.25 $X2=0.17
+ $Y2=1.95
r79 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.655
+ $Y=1.505 $X2=2.655 $Y2=1.505
r80 25 27 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.655 $Y=0.83
+ $X2=2.655 $Y2=1.505
r81 23 25 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.49 $Y=0.745
+ $X2=2.655 $Y2=0.83
r82 23 24 133.417 $w=1.68e-07 $l=2.045e-06 $layer=LI1_cond $X=2.49 $Y=0.745
+ $X2=0.445 $Y2=0.745
r83 16 30 8.99121 $w=3.58e-07 $l=1.8e-07 $layer=LI1_cond $X=0.265 $Y=1.07
+ $X2=0.265 $Y2=1.25
r84 16 18 3.68142 $w=3.58e-07 $l=1.15e-07 $layer=LI1_cond $X=0.265 $Y=1.07
+ $X2=0.265 $Y2=0.955
r85 15 24 8.02311 $w=1.7e-07 $l=2.18403e-07 $layer=LI1_cond $X=0.265 $Y=0.83
+ $X2=0.445 $Y2=0.745
r86 15 18 4.00154 $w=3.58e-07 $l=1.25e-07 $layer=LI1_cond $X=0.265 $Y=0.83
+ $X2=0.265 $Y2=0.955
r87 12 14 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.255 $Y=1.085
+ $X2=3.255 $Y2=0.69
r88 11 28 71.6767 $w=2.32e-07 $l=4.19464e-07 $layer=POLY_cond $X=2.82 $Y=1.16
+ $X2=2.655 $Y2=1.505
r89 10 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.18 $Y=1.16
+ $X2=3.255 $Y2=1.085
r90 10 11 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=3.18 $Y=1.16
+ $X2=2.82 $Y2=1.16
r91 7 28 84.9572 $w=2.32e-07 $l=4.15812e-07 $layer=POLY_cond $X=2.73 $Y=1.885
+ $X2=2.655 $Y2=1.505
r92 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.73 $Y=1.885
+ $X2=2.73 $Y2=2.46
r93 2 32 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.165
+ $Y=1.97 $X2=0.31 $Y2=2.115
r94 1 18 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.68 $X2=0.28 $Y2=0.955
.ends

.subckt PM_SKY130_FD_SC_LS__DLRTN_4%A_348_392# 1 2 7 9 12 15 16 21 23 25 26 31
+ 37
c87 31 0 1.51556e-19 $X=2.12 $Y=1.125
r88 36 37 7.70264 $w=5.08e-07 $l=8.5e-08 $layer=LI1_cond $X=2.12 $Y=2.175
+ $X2=2.205 $Y2=2.175
r89 34 36 5.51134 $w=5.08e-07 $l=2.35e-07 $layer=LI1_cond $X=1.885 $Y=2.175
+ $X2=2.12 $Y2=2.175
r90 29 31 7.14515 $w=2.48e-07 $l=1.55e-07 $layer=LI1_cond $X=1.965 $Y=1.125
+ $X2=2.12 $Y2=1.125
r91 26 40 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.095 $Y=1.355
+ $X2=4.095 $Y2=1.19
r92 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.095
+ $Y=1.355 $X2=4.095 $Y2=1.355
r93 23 25 25.668 $w=3.28e-07 $l=7.35e-07 $layer=LI1_cond $X=3.36 $Y=1.355
+ $X2=4.095 $Y2=1.355
r94 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.195
+ $Y=1.61 $X2=3.195 $Y2=1.61
r95 19 21 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=3.195 $Y=1.92
+ $X2=3.195 $Y2=1.61
r96 18 23 6.81649 $w=3.3e-07 $l=2.33345e-07 $layer=LI1_cond $X=3.195 $Y=1.52
+ $X2=3.36 $Y2=1.355
r97 18 21 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=3.195 $Y=1.52
+ $X2=3.195 $Y2=1.61
r98 16 19 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.03 $Y=2.005
+ $X2=3.195 $Y2=1.92
r99 16 37 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=3.03 $Y=2.005
+ $X2=2.205 $Y2=2.005
r100 15 36 7.28118 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=2.12 $Y=1.92
+ $X2=2.12 $Y2=2.175
r101 14 31 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.12 $Y=1.25
+ $X2=2.12 $Y2=1.125
r102 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.12 $Y=1.25
+ $X2=2.12 $Y2=1.92
r103 12 40 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.12 $Y=0.58
+ $X2=4.12 $Y2=1.19
r104 7 22 56.7567 $w=2.92e-07 $l=3.10242e-07 $layer=POLY_cond $X=3.12 $Y=1.885
+ $X2=3.195 $Y2=1.61
r105 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.12 $Y=1.885
+ $X2=3.12 $Y2=2.46
r106 2 34 600 $w=1.7e-07 $l=2.88531e-07 $layer=licon1_PDIFF $count=1 $X=1.74
+ $Y=1.96 $X2=1.885 $Y2=2.185
r107 1 29 182 $w=1.7e-07 $l=6.63551e-07 $layer=licon1_NDIFF $count=1 $X=1.82
+ $Y=0.49 $X2=1.965 $Y2=1.085
.ends

.subckt PM_SKY130_FD_SC_LS__DLRTN_4%A_888_406# 1 2 3 10 12 15 17 18 19 21 22 26
+ 28 30 33 35 37 40 42 44 47 50 52 58 63 65 69 78 81 83 84 85 86 95
c189 58 0 1.15495e-20 $X=5.655 $Y=2.03
r190 92 93 31.5204 $w=3.67e-07 $l=2.4e-07 $layer=POLY_cond $X=8.435 $Y=1.532
+ $X2=8.675 $Y2=1.532
r191 91 92 24.9537 $w=3.67e-07 $l=1.9e-07 $layer=POLY_cond $X=8.245 $Y=1.532
+ $X2=8.435 $Y2=1.532
r192 88 89 15.7602 $w=3.67e-07 $l=1.2e-07 $layer=POLY_cond $X=7.815 $Y=1.532
+ $X2=7.935 $Y2=1.532
r193 85 86 8.63679 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=7.725 $Y=1.545
+ $X2=7.895 $Y2=1.545
r194 79 95 9.85014 $w=3.67e-07 $l=7.5e-08 $layer=POLY_cond $X=8.91 $Y=1.532
+ $X2=8.985 $Y2=1.532
r195 79 93 30.8638 $w=3.67e-07 $l=2.35e-07 $layer=POLY_cond $X=8.91 $Y=1.532
+ $X2=8.675 $Y2=1.532
r196 78 79 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=8.91
+ $Y=1.465 $X2=8.91 $Y2=1.465
r197 76 91 1.97003 $w=3.67e-07 $l=1.5e-08 $layer=POLY_cond $X=8.23 $Y=1.532
+ $X2=8.245 $Y2=1.532
r198 76 89 38.7439 $w=3.67e-07 $l=2.95e-07 $layer=POLY_cond $X=8.23 $Y=1.532
+ $X2=7.935 $Y2=1.532
r199 75 78 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=8.23 $Y=1.465
+ $X2=8.91 $Y2=1.465
r200 75 86 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=8.23 $Y=1.465
+ $X2=7.895 $Y2=1.465
r201 75 76 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=8.23
+ $Y=1.465 $X2=8.23 $Y2=1.465
r202 72 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.82 $Y=1.705
+ $X2=6.655 $Y2=1.705
r203 72 85 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=6.82 $Y=1.705
+ $X2=7.725 $Y2=1.705
r204 67 84 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.655 $Y=1.79
+ $X2=6.655 $Y2=1.705
r205 67 69 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=6.655 $Y=1.79
+ $X2=6.655 $Y2=2.245
r206 66 81 2.76166 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=5.835 $Y=1.705
+ $X2=5.662 $Y2=1.705
r207 65 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.49 $Y=1.705
+ $X2=6.655 $Y2=1.705
r208 65 66 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=6.49 $Y=1.705
+ $X2=5.835 $Y2=1.705
r209 61 81 3.70735 $w=2.5e-07 $l=1.23386e-07 $layer=LI1_cond $X=5.75 $Y=1.62
+ $X2=5.662 $Y2=1.705
r210 61 63 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=5.75 $Y=1.62
+ $X2=5.75 $Y2=0.81
r211 58 83 5.16603 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=5.655 $Y=2.03
+ $X2=5.655 $Y2=2.195
r212 57 81 3.70735 $w=2.5e-07 $l=8.84308e-08 $layer=LI1_cond $X=5.655 $Y=1.79
+ $X2=5.662 $Y2=1.705
r213 57 58 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=5.655 $Y=1.79
+ $X2=5.655 $Y2=2.03
r214 54 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.605
+ $Y=2.195 $X2=4.605 $Y2=2.195
r215 52 83 1.34256 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=5.49 $Y=2.195
+ $X2=5.655 $Y2=2.195
r216 52 54 30.9064 $w=3.28e-07 $l=8.85e-07 $layer=LI1_cond $X=5.49 $Y=2.195
+ $X2=4.605 $Y2=2.195
r217 45 95 15.7602 $w=3.67e-07 $l=2.85769e-07 $layer=POLY_cond $X=9.105 $Y=1.3
+ $X2=8.985 $Y2=1.532
r218 45 47 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=9.105 $Y=1.3
+ $X2=9.105 $Y2=0.74
r219 42 95 23.77 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=8.985 $Y=1.765
+ $X2=8.985 $Y2=1.532
r220 42 44 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.985 $Y=1.765
+ $X2=8.985 $Y2=2.4
r221 38 93 23.77 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=8.675 $Y=1.3
+ $X2=8.675 $Y2=1.532
r222 38 40 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=8.675 $Y=1.3
+ $X2=8.675 $Y2=0.74
r223 35 92 23.77 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=8.435 $Y=1.765
+ $X2=8.435 $Y2=1.532
r224 35 37 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.435 $Y=1.765
+ $X2=8.435 $Y2=2.4
r225 31 91 23.77 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=8.245 $Y=1.3
+ $X2=8.245 $Y2=1.532
r226 31 33 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=8.245 $Y=1.3
+ $X2=8.245 $Y2=0.74
r227 28 89 23.77 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=7.935 $Y=1.765
+ $X2=7.935 $Y2=1.532
r228 28 30 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.935 $Y=1.765
+ $X2=7.935 $Y2=2.4
r229 24 88 23.77 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=7.815 $Y=1.3
+ $X2=7.815 $Y2=1.532
r230 24 26 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=7.815 $Y=1.3
+ $X2=7.815 $Y2=0.74
r231 23 50 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=7.575 $Y=1.555
+ $X2=7.485 $Y2=1.555
r232 22 88 27.1901 $w=3.67e-07 $l=8.57321e-08 $layer=POLY_cond $X=7.74 $Y=1.555
+ $X2=7.815 $Y2=1.532
r233 22 23 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.74 $Y=1.555
+ $X2=7.575 $Y2=1.555
r234 19 50 83.7788 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=7.485 $Y=1.765
+ $X2=7.485 $Y2=1.555
r235 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.485 $Y=1.765
+ $X2=7.485 $Y2=2.4
r236 18 55 34.1752 $w=2.99e-07 $l=1.86145e-07 $layer=POLY_cond $X=4.56 $Y=2.03
+ $X2=4.605 $Y2=2.195
r237 17 49 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=4.56 $Y=1.825
+ $X2=4.56 $Y2=1.735
r238 17 18 79.6855 $w=1.8e-07 $l=2.05e-07 $layer=POLY_cond $X=4.56 $Y=1.825
+ $X2=4.56 $Y2=2.03
r239 15 49 592.245 $w=1.5e-07 $l=1.155e-06 $layer=POLY_cond $X=4.545 $Y=0.58
+ $X2=4.545 $Y2=1.735
r240 10 55 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=4.53 $Y=2.445
+ $X2=4.605 $Y2=2.195
r241 10 12 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.53 $Y=2.445
+ $X2=4.53 $Y2=2.73
r242 3 69 300 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=2 $X=6.455
+ $Y=2.1 $X2=6.655 $Y2=2.245
r243 2 83 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=5.505
+ $Y=2.1 $X2=5.655 $Y2=2.245
r244 1 63 182 $w=1.7e-07 $l=5.05173e-07 $layer=licon1_NDIFF $count=1 $X=5.61
+ $Y=0.37 $X2=5.75 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_LS__DLRTN_4%A_639_392# 1 2 8 9 11 12 14 16 17 19 20 22
+ 23 28 29 30 33 35 36 37 38 46
c118 46 0 1.47145e-19 $X=5.88 $Y=1.455
r119 46 47 6.42163 $w=6.38e-07 $l=8.5e-08 $layer=POLY_cond $X=5.88 $Y=1.455
+ $X2=5.965 $Y2=1.455
r120 45 46 26.0643 $w=6.38e-07 $l=3.45e-07 $layer=POLY_cond $X=5.535 $Y=1.455
+ $X2=5.88 $Y2=1.455
r121 44 45 7.9326 $w=6.38e-07 $l=1.05e-07 $layer=POLY_cond $X=5.43 $Y=1.455
+ $X2=5.535 $Y2=1.455
r122 42 44 28.3307 $w=6.38e-07 $l=3.75e-07 $layer=POLY_cond $X=5.055 $Y=1.455
+ $X2=5.43 $Y2=1.455
r123 41 42 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.055
+ $Y=1.285 $X2=5.055 $Y2=1.285
r124 39 41 15.8148 $w=2.7e-07 $l=3.5e-07 $layer=LI1_cond $X=4.985 $Y=0.935
+ $X2=4.985 $Y2=1.285
r125 37 41 2.4733 $w=4.05e-07 $l=5.05272e-08 $layer=LI1_cond $X=5.017 $Y=1.322
+ $X2=4.985 $Y2=1.285
r126 37 38 10.4716 $w=4.03e-07 $l=3.68e-07 $layer=LI1_cond $X=5.017 $Y=1.322
+ $X2=5.017 $Y2=1.69
r127 35 39 3.44395 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=4.815 $Y=0.935
+ $X2=4.985 $Y2=0.935
r128 35 36 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=4.815 $Y=0.935
+ $X2=4.07 $Y2=0.935
r129 31 36 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.905 $Y=0.85
+ $X2=4.07 $Y2=0.935
r130 31 33 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=3.905 $Y=0.85
+ $X2=3.905 $Y2=0.565
r131 29 38 8.41448 $w=1.7e-07 $l=2.40778e-07 $layer=LI1_cond $X=4.815 $Y=1.775
+ $X2=5.017 $Y2=1.69
r132 29 30 72.7433 $w=1.68e-07 $l=1.115e-06 $layer=LI1_cond $X=4.815 $Y=1.775
+ $X2=3.7 $Y2=1.775
r133 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.615 $Y=1.86
+ $X2=3.7 $Y2=1.775
r134 27 28 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=3.615 $Y=1.86
+ $X2=3.615 $Y2=2.26
r135 23 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.53 $Y=2.345
+ $X2=3.615 $Y2=2.26
r136 23 25 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=3.53 $Y=2.345
+ $X2=3.345 $Y2=2.345
r137 20 47 37.6732 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=5.965 $Y=1.12
+ $X2=5.965 $Y2=1.455
r138 20 22 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=5.965 $Y=1.12
+ $X2=5.965 $Y2=0.69
r139 17 19 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=5.88 $Y=2.025
+ $X2=5.88 $Y2=2.52
r140 16 17 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.88 $Y=1.935
+ $X2=5.88 $Y2=2.025
r141 15 46 32.9664 $w=1.8e-07 $l=3.35e-07 $layer=POLY_cond $X=5.88 $Y=1.79
+ $X2=5.88 $Y2=1.455
r142 15 16 56.3629 $w=1.8e-07 $l=1.45e-07 $layer=POLY_cond $X=5.88 $Y=1.79
+ $X2=5.88 $Y2=1.935
r143 12 45 37.6732 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=5.535 $Y=1.12
+ $X2=5.535 $Y2=1.455
r144 12 14 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=5.535 $Y=1.12
+ $X2=5.535 $Y2=0.69
r145 9 11 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=5.43 $Y=2.025
+ $X2=5.43 $Y2=2.52
r146 8 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.43 $Y=1.935 $X2=5.43
+ $Y2=2.025
r147 7 44 32.9664 $w=1.8e-07 $l=3.35e-07 $layer=POLY_cond $X=5.43 $Y=1.79
+ $X2=5.43 $Y2=1.455
r148 7 8 56.3629 $w=1.8e-07 $l=1.45e-07 $layer=POLY_cond $X=5.43 $Y=1.79
+ $X2=5.43 $Y2=1.935
r149 2 25 600 $w=1.7e-07 $l=4.53845e-07 $layer=licon1_PDIFF $count=1 $X=3.195
+ $Y=1.96 $X2=3.345 $Y2=2.345
r150 1 33 182 $w=1.7e-07 $l=2.72213e-07 $layer=licon1_NDIFF $count=1 $X=3.72
+ $Y=0.37 $X2=3.905 $Y2=0.565
.ends

.subckt PM_SKY130_FD_SC_LS__DLRTN_4%RESET_B 2 3 5 6 8 9 11 13 14 16 17 18 19 26
c62 3 0 1.15495e-20 $X=6.38 $Y=2.025
r63 26 28 7.94506 $w=4.55e-07 $l=7.5e-08 $layer=POLY_cond $X=6.825 $Y=1.355
+ $X2=6.9 $Y2=1.355
r64 26 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.825
+ $Y=1.285 $X2=6.825 $Y2=1.285
r65 24 26 45.5516 $w=4.55e-07 $l=4.3e-07 $layer=POLY_cond $X=6.395 $Y=1.355
+ $X2=6.825 $Y2=1.355
r66 23 24 1.58901 $w=4.55e-07 $l=1.5e-08 $layer=POLY_cond $X=6.38 $Y=1.355
+ $X2=6.395 $Y2=1.355
r67 18 19 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=6.96 $Y=1.285
+ $X2=7.44 $Y2=1.285
r68 18 27 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=6.96 $Y=1.285
+ $X2=6.825 $Y2=1.285
r69 17 27 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=6.48 $Y=1.285
+ $X2=6.825 $Y2=1.285
r70 14 16 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=6.9 $Y=2.025 $X2=6.9
+ $Y2=2.52
r71 13 14 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.9 $Y=1.935 $X2=6.9
+ $Y2=2.025
r72 12 28 24.5593 $w=1.8e-07 $l=2.35e-07 $layer=POLY_cond $X=6.9 $Y=1.59 $X2=6.9
+ $Y2=1.355
r73 12 13 134.105 $w=1.8e-07 $l=3.45e-07 $layer=POLY_cond $X=6.9 $Y=1.59 $X2=6.9
+ $Y2=1.935
r74 9 26 29.0417 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=6.825 $Y=1.12
+ $X2=6.825 $Y2=1.355
r75 9 11 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=6.825 $Y=1.12
+ $X2=6.825 $Y2=0.69
r76 6 24 29.0417 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=6.395 $Y=1.12
+ $X2=6.395 $Y2=1.355
r77 6 8 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=6.395 $Y=1.12
+ $X2=6.395 $Y2=0.69
r78 3 5 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=6.38 $Y=2.025 $X2=6.38
+ $Y2=2.52
r79 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.38 $Y=1.935 $X2=6.38
+ $Y2=2.025
r80 1 23 24.5593 $w=1.8e-07 $l=2.35e-07 $layer=POLY_cond $X=6.38 $Y=1.59
+ $X2=6.38 $Y2=1.355
r81 1 2 134.105 $w=1.8e-07 $l=3.45e-07 $layer=POLY_cond $X=6.38 $Y=1.59 $X2=6.38
+ $Y2=1.935
.ends

.subckt PM_SKY130_FD_SC_LS__DLRTN_4%VPWR 1 2 3 4 5 6 7 26 28 32 36 40 42 44 47
+ 50 54 55 57 58 59 82 87 92 95 97 101
r104 100 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r105 97 98 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r106 94 95 11.3415 $w=7.83e-07 $l=1.65e-07 $layer=LI1_cond $X=5.155 $Y=3.022
+ $X2=5.32 $Y2=3.022
r107 91 98 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33 $X2=6
+ $Y2=3.33
r108 90 94 1.75222 $w=7.83e-07 $l=1.15e-07 $layer=LI1_cond $X=5.04 $Y=3.022
+ $X2=5.155 $Y2=3.022
r109 90 92 15.6839 $w=7.83e-07 $l=4.5e-07 $layer=LI1_cond $X=5.04 $Y=3.022
+ $X2=4.59 $Y2=3.022
r110 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r111 87 88 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r112 85 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=9.36 $Y2=3.33
r113 84 85 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r114 82 100 4.53846 $w=1.7e-07 $l=2.77e-07 $layer=LI1_cond $X=9.045 $Y=3.33
+ $X2=9.322 $Y2=3.33
r115 82 84 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=9.045 $Y=3.33
+ $X2=8.88 $Y2=3.33
r116 81 85 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.88 $Y2=3.33
r117 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r118 78 81 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.92 $Y2=3.33
r119 78 98 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=3.33 $X2=6
+ $Y2=3.33
r120 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r121 75 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.32 $Y=3.33
+ $X2=6.155 $Y2=3.33
r122 75 77 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=6.32 $Y=3.33
+ $X2=6.96 $Y2=3.33
r123 73 92 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=4.56 $Y=3.33 $X2=4.59
+ $Y2=3.33
r124 73 74 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r125 71 74 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=4.56 $Y2=3.33
r126 70 73 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=2.64 $Y=3.33
+ $X2=4.56 $Y2=3.33
r127 70 71 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r128 67 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r129 66 67 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r130 64 67 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r131 64 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r132 63 66 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r133 63 64 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r134 61 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.975 $Y=3.33
+ $X2=0.81 $Y2=3.33
r135 61 63 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.975 $Y=3.33
+ $X2=1.2 $Y2=3.33
r136 59 91 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.8 $Y=3.33
+ $X2=5.04 $Y2=3.33
r137 59 74 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.8 $Y=3.33
+ $X2=4.56 $Y2=3.33
r138 57 80 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=8.045 $Y=3.33
+ $X2=7.92 $Y2=3.33
r139 57 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.045 $Y=3.33
+ $X2=8.21 $Y2=3.33
r140 56 84 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=8.375 $Y=3.33
+ $X2=8.88 $Y2=3.33
r141 56 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.375 $Y=3.33
+ $X2=8.21 $Y2=3.33
r142 54 77 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=7.045 $Y=3.33
+ $X2=6.96 $Y2=3.33
r143 54 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.045 $Y=3.33
+ $X2=7.21 $Y2=3.33
r144 53 80 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=7.375 $Y=3.33
+ $X2=7.92 $Y2=3.33
r145 53 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.375 $Y=3.33
+ $X2=7.21 $Y2=3.33
r146 51 70 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=2.585 $Y=3.33
+ $X2=2.64 $Y2=3.33
r147 50 66 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=2.255 $Y=3.33
+ $X2=2.16 $Y2=3.33
r148 49 51 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.42 $Y=3.33
+ $X2=2.585 $Y2=3.33
r149 49 50 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.42 $Y=3.33
+ $X2=2.255 $Y2=3.33
r150 47 49 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=2.42 $Y=3.025
+ $X2=2.42 $Y2=3.33
r151 42 100 3.22771 $w=3.3e-07 $l=1.4854e-07 $layer=LI1_cond $X=9.21 $Y=3.245
+ $X2=9.322 $Y2=3.33
r152 42 44 32.8272 $w=3.28e-07 $l=9.4e-07 $layer=LI1_cond $X=9.21 $Y=3.245
+ $X2=9.21 $Y2=2.305
r153 38 58 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.21 $Y=3.245
+ $X2=8.21 $Y2=3.33
r154 38 40 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=8.21 $Y=3.245
+ $X2=8.21 $Y2=2.465
r155 34 55 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.21 $Y=3.245
+ $X2=7.21 $Y2=3.33
r156 34 36 34.9225 $w=3.28e-07 $l=1e-06 $layer=LI1_cond $X=7.21 $Y=3.245
+ $X2=7.21 $Y2=2.245
r157 30 97 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.155 $Y=3.245
+ $X2=6.155 $Y2=3.33
r158 30 32 34.9225 $w=3.28e-07 $l=1e-06 $layer=LI1_cond $X=6.155 $Y=3.245
+ $X2=6.155 $Y2=2.245
r159 28 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.99 $Y=3.33
+ $X2=6.155 $Y2=3.33
r160 28 95 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.99 $Y=3.33
+ $X2=5.32 $Y2=3.33
r161 24 87 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.81 $Y=3.245
+ $X2=0.81 $Y2=3.33
r162 24 26 39.4624 $w=3.28e-07 $l=1.13e-06 $layer=LI1_cond $X=0.81 $Y=3.245
+ $X2=0.81 $Y2=2.115
r163 7 44 300 $w=1.7e-07 $l=5.34766e-07 $layer=licon1_PDIFF $count=2 $X=9.06
+ $Y=1.84 $X2=9.21 $Y2=2.305
r164 6 40 300 $w=1.7e-07 $l=7.1807e-07 $layer=licon1_PDIFF $count=2 $X=8.01
+ $Y=1.84 $X2=8.21 $Y2=2.465
r165 5 36 300 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=2 $X=6.975
+ $Y=2.1 $X2=7.21 $Y2=2.245
r166 4 32 300 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=2 $X=5.955
+ $Y=2.1 $X2=6.155 $Y2=2.245
r167 3 94 300 $w=1.7e-07 $l=6.7361e-07 $layer=licon1_PDIFF $count=2 $X=4.605
+ $Y=2.52 $X2=5.155 $Y2=2.795
r168 2 47 600 $w=1.7e-07 $l=1.17665e-06 $layer=licon1_PDIFF $count=1 $X=2.185
+ $Y=1.96 $X2=2.42 $Y2=3.025
r169 1 26 300 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=2 $X=0.61
+ $Y=1.97 $X2=0.81 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_LS__DLRTN_4%Q 1 2 3 4 13 15 17 21 24 27 31 33 37 43 44
+ 45 55
r76 55 56 6.0176 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=8.795 $Y=0.965
+ $X2=8.89 $Y2=0.965
r77 44 45 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=9.36 $Y=1.295
+ $X2=9.36 $Y2=1.665
r78 44 49 8.26753 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=9.36 $Y=1.295
+ $X2=9.36 $Y2=1.13
r79 43 49 2.85155 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=9.36 $Y=0.965
+ $X2=9.36 $Y2=1.13
r80 43 56 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=9.36 $Y=0.965
+ $X2=8.89 $Y2=0.965
r81 42 45 6.76434 $w=2.28e-07 $l=1.35e-07 $layer=LI1_cond $X=9.36 $Y=1.8
+ $X2=9.36 $Y2=1.665
r82 40 41 2.09535 $w=3.28e-07 $l=6e-08 $layer=LI1_cond $X=8.71 $Y=1.985 $X2=8.71
+ $Y2=2.045
r83 37 40 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=8.71 $Y=1.885 $X2=8.71
+ $Y2=1.985
r84 34 37 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.875 $Y=1.885
+ $X2=8.71 $Y2=1.885
r85 33 42 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=9.245 $Y=1.885
+ $X2=9.36 $Y2=1.8
r86 33 34 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=9.245 $Y=1.885
+ $X2=8.875 $Y2=1.885
r87 29 56 3.96751 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=8.89 $Y=0.8 $X2=8.89
+ $Y2=0.965
r88 29 31 16.0526 $w=1.88e-07 $l=2.75e-07 $layer=LI1_cond $X=8.89 $Y=0.8
+ $X2=8.89 $Y2=0.525
r89 25 41 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=8.71 $Y=2.13
+ $X2=8.71 $Y2=2.045
r90 25 27 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=8.71 $Y=2.13
+ $X2=8.71 $Y2=2.4
r91 24 55 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.125 $Y=1.045
+ $X2=8.795 $Y2=1.045
r92 19 24 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=8.03 $Y=0.96
+ $X2=8.125 $Y2=1.045
r93 19 21 25.3923 $w=1.88e-07 $l=4.35e-07 $layer=LI1_cond $X=8.03 $Y=0.96
+ $X2=8.03 $Y2=0.525
r94 18 36 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.875 $Y=2.045
+ $X2=7.71 $Y2=2.045
r95 17 41 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.545 $Y=2.045
+ $X2=8.71 $Y2=2.045
r96 17 18 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.545 $Y=2.045
+ $X2=7.875 $Y2=2.045
r97 13 36 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.71 $Y=2.13 $X2=7.71
+ $Y2=2.045
r98 13 15 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=7.71 $Y=2.13
+ $X2=7.71 $Y2=2.815
r99 4 40 600 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=1 $X=8.51
+ $Y=1.84 $X2=8.71 $Y2=1.985
r100 4 27 300 $w=1.7e-07 $l=6.5238e-07 $layer=licon1_PDIFF $count=2 $X=8.51
+ $Y=1.84 $X2=8.71 $Y2=2.4
r101 3 36 400 $w=1.7e-07 $l=3.52101e-07 $layer=licon1_PDIFF $count=1 $X=7.56
+ $Y=1.84 $X2=7.71 $Y2=2.125
r102 3 15 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=7.56
+ $Y=1.84 $X2=7.71 $Y2=2.815
r103 2 56 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=8.75
+ $Y=0.37 $X2=8.89 $Y2=0.965
r104 2 31 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=8.75
+ $Y=0.37 $X2=8.89 $Y2=0.525
r105 1 21 91 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=2 $X=7.89
+ $Y=0.37 $X2=8.03 $Y2=0.525
.ends

.subckt PM_SKY130_FD_SC_LS__DLRTN_4%VGND 1 2 3 4 5 6 7 24 28 32 34 38 42 44 46
+ 49 50 51 53 70 74 79 85 90 96 98 101 104 108
c119 28 0 1.47145e-19 $X=4.76 $Y=0.515
r120 107 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r121 104 105 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r122 101 102 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r123 99 102 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=0
+ $X2=7.44 $Y2=0
r124 98 99 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r125 94 96 6.66521 $w=5.73e-07 $l=5e-09 $layer=LI1_cond $X=3.12 $Y=0.202
+ $X2=3.125 $Y2=0.202
r126 94 95 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r127 92 94 3.32822 $w=5.73e-07 $l=1.6e-07 $layer=LI1_cond $X=2.96 $Y=0.202
+ $X2=3.12 $Y2=0.202
r128 89 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r129 88 92 6.65644 $w=5.73e-07 $l=3.2e-07 $layer=LI1_cond $X=2.64 $Y=0.202
+ $X2=2.96 $Y2=0.202
r130 88 90 13.4257 $w=5.73e-07 $l=3.3e-07 $layer=LI1_cond $X=2.64 $Y=0.202
+ $X2=2.31 $Y2=0.202
r131 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r132 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r133 83 108 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0
+ $X2=9.36 $Y2=0
r134 83 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=8.4
+ $Y2=0
r135 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r136 80 104 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.625 $Y=0
+ $X2=8.46 $Y2=0
r137 80 82 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=8.625 $Y=0
+ $X2=8.88 $Y2=0
r138 79 107 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=9.155 $Y=0
+ $X2=9.377 $Y2=0
r139 79 82 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=9.155 $Y=0
+ $X2=8.88 $Y2=0
r140 78 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.4
+ $Y2=0
r141 78 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0
+ $X2=7.44 $Y2=0
r142 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r143 75 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.765 $Y=0 $X2=7.6
+ $Y2=0
r144 75 77 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=7.765 $Y=0
+ $X2=7.92 $Y2=0
r145 74 104 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.295 $Y=0
+ $X2=8.46 $Y2=0
r146 74 77 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=8.295 $Y=0
+ $X2=7.92 $Y2=0
r147 73 99 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=6.48 $Y2=0
r148 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r149 70 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.445 $Y=0 $X2=6.61
+ $Y2=0
r150 70 72 91.6631 $w=1.68e-07 $l=1.405e-06 $layer=LI1_cond $X=6.445 $Y=0
+ $X2=5.04 $Y2=0
r151 69 95 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.56 $Y=0
+ $X2=3.12 $Y2=0
r152 68 96 93.6203 $w=1.68e-07 $l=1.435e-06 $layer=LI1_cond $X=4.56 $Y=0
+ $X2=3.125 $Y2=0
r153 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r154 65 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r155 64 90 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=2.16 $Y=0 $X2=2.31
+ $Y2=0
r156 64 65 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r157 62 65 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r158 62 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r159 61 64 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r160 61 62 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r161 59 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=0.79
+ $Y2=0
r162 59 61 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=1.2
+ $Y2=0
r163 56 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r164 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r165 53 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.625 $Y=0 $X2=0.79
+ $Y2=0
r166 53 55 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.625 $Y=0
+ $X2=0.24 $Y2=0
r167 51 73 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.8 $Y=0 $X2=5.04
+ $Y2=0
r168 51 69 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.8 $Y=0 $X2=4.56
+ $Y2=0
r169 49 68 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=4.595 $Y=0 $X2=4.56
+ $Y2=0
r170 49 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.595 $Y=0 $X2=4.76
+ $Y2=0
r171 48 72 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=4.925 $Y=0
+ $X2=5.04 $Y2=0
r172 48 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.925 $Y=0 $X2=4.76
+ $Y2=0
r173 44 107 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=9.32 $Y=0.085
+ $X2=9.377 $Y2=0
r174 44 46 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=9.32 $Y=0.085
+ $X2=9.32 $Y2=0.53
r175 40 104 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.46 $Y=0.085
+ $X2=8.46 $Y2=0
r176 40 42 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=8.46 $Y=0.085
+ $X2=8.46 $Y2=0.625
r177 36 101 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.6 $Y=0.085
+ $X2=7.6 $Y2=0
r178 36 38 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=7.6 $Y=0.085
+ $X2=7.6 $Y2=0.525
r179 35 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.775 $Y=0 $X2=6.61
+ $Y2=0
r180 34 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.435 $Y=0 $X2=7.6
+ $Y2=0
r181 34 35 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=7.435 $Y=0
+ $X2=6.775 $Y2=0
r182 30 98 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.61 $Y=0.085
+ $X2=6.61 $Y2=0
r183 30 32 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=6.61 $Y=0.085
+ $X2=6.61 $Y2=0.515
r184 26 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.76 $Y=0.085
+ $X2=4.76 $Y2=0
r185 26 28 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=4.76 $Y=0.085
+ $X2=4.76 $Y2=0.515
r186 22 85 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.79 $Y=0.085
+ $X2=0.79 $Y2=0
r187 22 24 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=0.79 $Y=0.085
+ $X2=0.79 $Y2=0.325
r188 7 46 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=9.18
+ $Y=0.37 $X2=9.32 $Y2=0.53
r189 6 42 182 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=1 $X=8.32
+ $Y=0.37 $X2=8.46 $Y2=0.625
r190 5 38 91 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=2 $X=7.455
+ $Y=0.37 $X2=7.6 $Y2=0.525
r191 4 32 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=6.47
+ $Y=0.37 $X2=6.61 $Y2=0.515
r192 3 28 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=4.62
+ $Y=0.37 $X2=4.76 $Y2=0.515
r193 2 92 91 $w=1.7e-07 $l=7.83167e-07 $layer=licon1_NDIFF $count=2 $X=2.255
+ $Y=0.49 $X2=2.96 $Y2=0.325
r194 1 24 182 $w=1.7e-07 $l=4.51802e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.68 $X2=0.79 $Y2=0.325
.ends

.subckt PM_SKY130_FD_SC_LS__DLRTN_4%A_1035_74# 1 2 3 12 14 15 17 19 20 22 24
r45 22 29 2.91016 $w=2.6e-07 $l=9e-08 $layer=LI1_cond $X=7.075 $Y=0.77 $X2=7.075
+ $Y2=0.86
r46 22 24 11.0812 $w=2.58e-07 $l=2.5e-07 $layer=LI1_cond $X=7.075 $Y=0.77
+ $X2=7.075 $Y2=0.52
r47 21 27 4.10122 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=6.265 $Y=0.86
+ $X2=6.14 $Y2=0.86
r48 20 29 4.20357 $w=1.8e-07 $l=1.3e-07 $layer=LI1_cond $X=6.945 $Y=0.86
+ $X2=7.075 $Y2=0.86
r49 20 21 41.899 $w=1.78e-07 $l=6.8e-07 $layer=LI1_cond $X=6.945 $Y=0.86
+ $X2=6.265 $Y2=0.86
r50 17 27 2.95288 $w=2.5e-07 $l=9e-08 $layer=LI1_cond $X=6.14 $Y=0.77 $X2=6.14
+ $Y2=0.86
r51 17 19 12.6769 $w=2.48e-07 $l=2.75e-07 $layer=LI1_cond $X=6.14 $Y=0.77
+ $X2=6.14 $Y2=0.495
r52 16 19 3.22684 $w=2.48e-07 $l=7e-08 $layer=LI1_cond $X=6.14 $Y=0.425 $X2=6.14
+ $Y2=0.495
r53 14 16 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.015 $Y=0.34
+ $X2=6.14 $Y2=0.425
r54 14 15 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=6.015 $Y=0.34
+ $X2=5.485 $Y2=0.34
r55 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.32 $Y=0.425
+ $X2=5.485 $Y2=0.34
r56 10 12 2.44458 $w=3.28e-07 $l=7e-08 $layer=LI1_cond $X=5.32 $Y=0.425 $X2=5.32
+ $Y2=0.495
r57 3 29 182 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_NDIFF $count=1 $X=6.9
+ $Y=0.37 $X2=7.04 $Y2=0.86
r58 3 24 182 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=1 $X=6.9
+ $Y=0.37 $X2=7.04 $Y2=0.52
r59 2 27 182 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_NDIFF $count=1 $X=6.04
+ $Y=0.37 $X2=6.18 $Y2=0.865
r60 2 19 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=6.04
+ $Y=0.37 $X2=6.18 $Y2=0.495
r61 1 12 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=5.175
+ $Y=0.37 $X2=5.32 $Y2=0.495
.ends

