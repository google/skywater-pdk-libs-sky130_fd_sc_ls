* NGSPICE file created from sky130_fd_sc_ls__a211o_4.ext - technology: sky130A

.subckt sky130_fd_sc_ls__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
M1000 a_1064_123# A2 VGND VNB nshort w=640000u l=150000u
+  ad=3.584e+11p pd=3.68e+06u as=1.50765e+12p ps=1.284e+07u
M1001 X a_105_280# VGND VNB nshort w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=0p ps=0u
M1002 a_105_280# A1 a_1064_123# VNB nshort w=640000u l=150000u
+  ad=5.79525e+11p pd=5.76e+06u as=0p ps=0u
M1003 a_517_392# B1 a_602_392# VPB phighvt w=1e+06u l=150000u
+  ad=1.155e+12p pd=1.031e+07u as=6.75e+11p ps=5.35e+06u
M1004 a_105_280# C1 a_602_392# VPB phighvt w=1e+06u l=150000u
+  ad=3e+11p pd=2.6e+06u as=0p ps=0u
M1005 a_105_280# B1 VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR A2 a_517_392# VPB phighvt w=1e+06u l=150000u
+  ad=1.907e+12p pd=1.433e+07u as=0p ps=0u
M1007 VPWR A1 a_517_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR a_105_280# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=6.72e+11p ps=5.68e+06u
M1009 a_602_392# C1 a_105_280# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND a_105_280# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 X a_105_280# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_517_392# A1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 X a_105_280# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_517_392# A2 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND B1 a_105_280# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 X a_105_280# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_1064_123# A1 a_105_280# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND a_105_280# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR a_105_280# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND C1 a_105_280# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_105_280# C1 VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND A2 a_1064_123# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_602_392# B1 a_517_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

