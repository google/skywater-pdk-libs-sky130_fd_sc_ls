* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
M1000 a_841_368# A3 Y VPB phighvt w=1.12e+06u l=150000u
+  ad=1.8592e+12p pd=1.452e+07u as=1.8536e+12p ps=1.227e+07u
M1001 VGND A2 a_459_74# VNB nshort w=740000u l=150000u
+  ad=2.19225e+12p pd=1.657e+07u as=1.7316e+12p ps=1.652e+07u
M1002 a_459_74# B1 a_27_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=1.02765e+12p ps=1.022e+07u
M1003 Y C1 a_27_74# VNB nshort w=740000u l=150000u
+  ad=4.181e+11p pd=4.09e+06u as=0p ps=0u
M1004 a_459_74# A2 VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND A1 a_459_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_841_368# A2 a_1350_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=1.4e+12p ps=1.146e+07u
M1007 VPWR A1 a_1350_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=3.6176e+12p pd=1.99e+07u as=0p ps=0u
M1008 VGND A3 a_459_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_841_368# A3 Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_459_74# A3 VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR C1 Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_459_74# A1 VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_1350_368# A1 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_27_74# B1 a_459_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_27_74# B1 a_459_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_459_74# A2 VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_1350_368# A1 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_27_74# C1 Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_27_74# C1 Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 Y B1 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_1350_368# A2 a_841_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 Y C1 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VPWR A1 a_1350_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND A3 a_459_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VGND A2 a_459_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_841_368# A2 a_1350_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_459_74# B1 a_27_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VPWR B1 Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 Y C1 a_27_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 Y A3 a_841_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_459_74# A3 VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 Y A3 a_841_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_1350_368# A2 a_841_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 VGND A1 a_459_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_459_74# A1 VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
