* File: sky130_fd_sc_ls__and3b_2.spice
* Created: Wed Sep  2 10:55:11 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__and3b_2.pex.spice"
.subckt sky130_fd_sc_ls__and3b_2  VNB VPB A_N B C VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* C	C
* B	B
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1010 N_VGND_M1010_d N_A_N_M1010_g N_A_27_88#_M1010_s VNB NSHORT L=0.15 W=0.55
+ AD=0.16225 AS=0.15675 PD=1.69 PS=1.67 NRD=0 NRS=0 M=1 R=3.66667 SA=75000.2
+ SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1006 A_376_74# N_A_27_88#_M1006_g N_A_284_368#_M1006_s VNB NSHORT L=0.15
+ W=0.74 AD=0.0888 AS=0.2109 PD=0.98 PS=2.05 NRD=10.536 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75002.2 A=0.111 P=1.78 MULT=1
MM1005 A_454_74# N_B_M1005_g A_376_74# VNB NSHORT L=0.15 W=0.74 AD=0.1554
+ AS=0.0888 PD=1.16 PS=0.98 NRD=25.128 NRS=10.536 M=1 R=4.93333 SA=75000.6
+ SB=75001.8 A=0.111 P=1.78 MULT=1
MM1000 N_VGND_M1000_d N_C_M1000_g A_454_74# VNB NSHORT L=0.15 W=0.74 AD=0.1554
+ AS=0.1554 PD=1.16 PS=1.16 NRD=0 NRS=25.128 M=1 R=4.93333 SA=75001.2 SB=75001.2
+ A=0.111 P=1.78 MULT=1
MM1002 N_X_M1002_d N_A_284_368#_M1002_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1554 PD=1.02 PS=1.16 NRD=0 NRS=22.692 M=1 R=4.93333 SA=75001.7
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1011 N_X_M1002_d N_A_284_368#_M1011_g N_VGND_M1011_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1007 N_VPWR_M1007_d N_A_N_M1007_g N_A_27_88#_M1007_s VPB PHIGHVT L=0.15 W=0.84
+ AD=0.2562 AS=0.2478 PD=2.29 PS=2.27 NRD=3.5066 NRS=2.3443 M=1 R=5.6 SA=75000.2
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1003 N_VPWR_M1003_d N_A_27_88#_M1003_g N_A_284_368#_M1003_s VPB PHIGHVT L=0.15
+ W=1 AD=0.21 AS=0.295 PD=1.42 PS=2.59 NRD=11.8003 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75002.2 A=0.15 P=2.3 MULT=1
MM1001 N_A_284_368#_M1001_d N_B_M1001_g N_VPWR_M1003_d VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.21 PD=1.3 PS=1.42 NRD=1.9503 NRS=15.7403 M=1 R=6.66667 SA=75000.8
+ SB=75001.7 A=0.15 P=2.3 MULT=1
MM1004 N_VPWR_M1004_d N_C_M1004_g N_A_284_368#_M1001_d VPB PHIGHVT L=0.15 W=1
+ AD=0.20066 AS=0.15 PD=1.42453 PS=1.3 NRD=19.7 NRS=1.9503 M=1 R=6.66667
+ SA=75001.2 SB=75001.2 A=0.15 P=2.3 MULT=1
MM1008 N_VPWR_M1004_d N_A_284_368#_M1008_g N_X_M1008_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.22474 AS=0.1764 PD=1.59547 PS=1.435 NRD=1.7533 NRS=2.6201 M=1 R=7.46667
+ SA=75001.6 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1009 N_VPWR_M1009_d N_A_284_368#_M1009_g N_X_M1008_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.1764 PD=2.83 PS=1.435 NRD=1.7533 NRS=3.5066 M=1 R=7.46667
+ SA=75002.1 SB=75000.2 A=0.168 P=2.54 MULT=1
DX12_noxref VNB VPB NWDIODE A=8.742 P=13.12
*
.include "sky130_fd_sc_ls__and3b_2.pxi.spice"
*
.ends
*
*
