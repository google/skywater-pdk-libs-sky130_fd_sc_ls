* File: sky130_fd_sc_ls__dlrbp_1.pxi.spice
* Created: Wed Sep  2 11:03:24 2020
* 
x_PM_SKY130_FD_SC_LS__DLRBP_1%D N_D_M1001_g N_D_c_159_n N_D_M1021_g D
+ PM_SKY130_FD_SC_LS__DLRBP_1%D
x_PM_SKY130_FD_SC_LS__DLRBP_1%GATE N_GATE_M1016_g N_GATE_c_191_n N_GATE_M1018_g
+ GATE PM_SKY130_FD_SC_LS__DLRBP_1%GATE
x_PM_SKY130_FD_SC_LS__DLRBP_1%A_226_104# N_A_226_104#_M1016_d
+ N_A_226_104#_M1018_d N_A_226_104#_c_224_n N_A_226_104#_M1002_g
+ N_A_226_104#_c_226_n N_A_226_104#_M1014_g N_A_226_104#_c_239_n
+ N_A_226_104#_M1010_g N_A_226_104#_c_240_n N_A_226_104#_c_241_n
+ N_A_226_104#_M1015_g N_A_226_104#_c_228_n N_A_226_104#_c_229_n
+ N_A_226_104#_c_243_n N_A_226_104#_c_244_n N_A_226_104#_c_230_n
+ N_A_226_104#_c_231_n N_A_226_104#_c_232_n N_A_226_104#_c_233_n
+ N_A_226_104#_c_234_n N_A_226_104#_c_235_n N_A_226_104#_c_236_n
+ N_A_226_104#_c_237_n PM_SKY130_FD_SC_LS__DLRBP_1%A_226_104#
x_PM_SKY130_FD_SC_LS__DLRBP_1%A_27_142# N_A_27_142#_M1001_s N_A_27_142#_M1021_s
+ N_A_27_142#_c_370_n N_A_27_142#_M1022_g N_A_27_142#_c_371_n
+ N_A_27_142#_M1007_g N_A_27_142#_c_372_n N_A_27_142#_c_373_n
+ N_A_27_142#_c_374_n N_A_27_142#_c_379_n N_A_27_142#_c_380_n
+ N_A_27_142#_c_381_n N_A_27_142#_c_382_n N_A_27_142#_c_375_n
+ N_A_27_142#_c_383_n N_A_27_142#_c_376_n N_A_27_142#_c_377_n
+ PM_SKY130_FD_SC_LS__DLRBP_1%A_27_142#
x_PM_SKY130_FD_SC_LS__DLRBP_1%A_353_98# N_A_353_98#_M1002_s N_A_353_98#_M1014_s
+ N_A_353_98#_M1008_g N_A_353_98#_c_465_n N_A_353_98#_M1004_g
+ N_A_353_98#_c_458_n N_A_353_98#_c_459_n N_A_353_98#_c_460_n
+ N_A_353_98#_c_570_p N_A_353_98#_c_461_n N_A_353_98#_c_468_n
+ N_A_353_98#_c_469_n N_A_353_98#_c_470_n N_A_353_98#_c_471_n
+ N_A_353_98#_c_506_n N_A_353_98#_c_462_n N_A_353_98#_c_463_n
+ N_A_353_98#_c_464_n PM_SKY130_FD_SC_LS__DLRBP_1%A_353_98#
x_PM_SKY130_FD_SC_LS__DLRBP_1%A_823_98# N_A_823_98#_M1019_s N_A_823_98#_M1009_d
+ N_A_823_98#_c_576_n N_A_823_98#_M1005_g N_A_823_98#_c_577_n
+ N_A_823_98#_c_590_n N_A_823_98#_M1006_g N_A_823_98#_M1000_g
+ N_A_823_98#_c_579_n N_A_823_98#_M1003_g N_A_823_98#_c_580_n
+ N_A_823_98#_M1012_g N_A_823_98#_c_582_n N_A_823_98#_c_593_n
+ N_A_823_98#_M1011_g N_A_823_98#_c_583_n N_A_823_98#_c_584_n
+ N_A_823_98#_c_594_n N_A_823_98#_c_595_n N_A_823_98#_c_585_n
+ N_A_823_98#_c_596_n N_A_823_98#_c_597_n N_A_823_98#_c_586_n
+ N_A_823_98#_c_587_n N_A_823_98#_c_599_n N_A_823_98#_c_588_n
+ PM_SKY130_FD_SC_LS__DLRBP_1%A_823_98#
x_PM_SKY130_FD_SC_LS__DLRBP_1%A_642_392# N_A_642_392#_M1008_d
+ N_A_642_392#_M1010_d N_A_642_392#_c_729_n N_A_642_392#_M1009_g
+ N_A_642_392#_M1019_g N_A_642_392#_c_723_n N_A_642_392#_c_724_n
+ N_A_642_392#_c_737_n N_A_642_392#_c_725_n N_A_642_392#_c_726_n
+ N_A_642_392#_c_727_n N_A_642_392#_c_747_n N_A_642_392#_c_734_n
+ N_A_642_392#_c_728_n PM_SKY130_FD_SC_LS__DLRBP_1%A_642_392#
x_PM_SKY130_FD_SC_LS__DLRBP_1%RESET_B N_RESET_B_c_811_n N_RESET_B_M1017_g
+ N_RESET_B_c_812_n N_RESET_B_M1023_g RESET_B N_RESET_B_c_813_n
+ PM_SKY130_FD_SC_LS__DLRBP_1%RESET_B
x_PM_SKY130_FD_SC_LS__DLRBP_1%A_1342_74# N_A_1342_74#_M1012_s
+ N_A_1342_74#_M1011_s N_A_1342_74#_M1020_g N_A_1342_74#_c_844_n
+ N_A_1342_74#_M1013_g N_A_1342_74#_c_845_n N_A_1342_74#_c_850_n
+ N_A_1342_74#_c_846_n N_A_1342_74#_c_847_n N_A_1342_74#_c_848_n
+ PM_SKY130_FD_SC_LS__DLRBP_1%A_1342_74#
x_PM_SKY130_FD_SC_LS__DLRBP_1%VPWR N_VPWR_M1021_d N_VPWR_M1014_d N_VPWR_M1006_d
+ N_VPWR_M1023_d N_VPWR_M1011_d N_VPWR_c_902_n N_VPWR_c_903_n N_VPWR_c_904_n
+ N_VPWR_c_905_n VPWR N_VPWR_c_906_n N_VPWR_c_907_n N_VPWR_c_908_n
+ N_VPWR_c_909_n N_VPWR_c_910_n N_VPWR_c_901_n N_VPWR_c_912_n N_VPWR_c_913_n
+ N_VPWR_c_914_n N_VPWR_c_915_n N_VPWR_c_916_n PM_SKY130_FD_SC_LS__DLRBP_1%VPWR
x_PM_SKY130_FD_SC_LS__DLRBP_1%Q N_Q_M1000_d N_Q_M1003_d N_Q_c_992_n N_Q_c_993_n
+ N_Q_c_995_n N_Q_c_994_n Q Q PM_SKY130_FD_SC_LS__DLRBP_1%Q
x_PM_SKY130_FD_SC_LS__DLRBP_1%Q_N N_Q_N_M1020_d N_Q_N_M1013_d N_Q_N_c_1033_n
+ N_Q_N_c_1034_n N_Q_N_c_1030_n Q_N Q_N Q_N PM_SKY130_FD_SC_LS__DLRBP_1%Q_N
x_PM_SKY130_FD_SC_LS__DLRBP_1%VGND N_VGND_M1001_d N_VGND_M1002_d N_VGND_M1005_d
+ N_VGND_M1017_d N_VGND_M1012_d N_VGND_c_1052_n N_VGND_c_1053_n N_VGND_c_1054_n
+ N_VGND_c_1055_n N_VGND_c_1056_n N_VGND_c_1057_n VGND N_VGND_c_1058_n
+ N_VGND_c_1059_n N_VGND_c_1060_n N_VGND_c_1061_n N_VGND_c_1062_n
+ N_VGND_c_1063_n N_VGND_c_1064_n N_VGND_c_1065_n N_VGND_c_1066_n
+ N_VGND_c_1067_n PM_SKY130_FD_SC_LS__DLRBP_1%VGND
cc_1 VNB N_D_M1001_g 0.0287436f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.985
cc_2 VNB N_D_c_159_n 0.0213869f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.915
cc_3 VNB D 0.00163867f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_4 VNB N_GATE_M1016_g 0.0268455f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.985
cc_5 VNB N_GATE_c_191_n 0.018171f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.915
cc_6 VNB GATE 0.00260178f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_7 VNB N_A_226_104#_c_224_n 0.015812f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.41
cc_8 VNB N_A_226_104#_M1002_g 0.0280298f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.615
cc_9 VNB N_A_226_104#_c_226_n 0.0105025f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.615
cc_10 VNB N_A_226_104#_M1015_g 0.04132f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_226_104#_c_228_n 0.00790686f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_226_104#_c_229_n 0.00496729f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_226_104#_c_230_n 0.00358065f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_226_104#_c_231_n 0.00163151f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_226_104#_c_232_n 0.00858829f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_226_104#_c_233_n 0.0444271f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_226_104#_c_234_n 0.0106508f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_226_104#_c_235_n 0.00483006f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_226_104#_c_236_n 0.00286045f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_226_104#_c_237_n 0.0221744f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_27_142#_c_370_n 0.0195808f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.41
cc_22 VNB N_A_27_142#_c_371_n 0.0111327f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.615
cc_23 VNB N_A_27_142#_c_372_n 0.0144876f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.615
cc_24 VNB N_A_27_142#_c_373_n 0.0083007f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_27_142#_c_374_n 0.0207946f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_27_142#_c_375_n 0.0129596f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_27_142#_c_376_n 0.0178451f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_27_142#_c_377_n 0.00167974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_353_98#_c_458_n 0.00208878f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_353_98#_c_459_n 0.0161497f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.615
cc_31 VNB N_A_353_98#_c_460_n 0.00294809f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_353_98#_c_461_n 0.0028445f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_353_98#_c_462_n 0.00711509f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_353_98#_c_463_n 0.0305419f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_353_98#_c_464_n 0.0159056f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_823_98#_c_576_n 0.0171346f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.41
cc_37 VNB N_A_823_98#_c_577_n 0.0236589f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.615
cc_38 VNB N_A_823_98#_M1000_g 0.0301114f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_823_98#_c_579_n 0.0234118f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_823_98#_c_580_n 0.0481818f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_823_98#_M1012_g 0.0437361f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_823_98#_c_582_n 0.00816122f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_823_98#_c_583_n 0.0200553f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_823_98#_c_584_n 0.00412378f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_823_98#_c_585_n 0.00790788f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_823_98#_c_586_n 7.85697e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_823_98#_c_587_n 0.00533523f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_823_98#_c_588_n 0.00752343f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_642_392#_M1019_g 0.027719f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.615
cc_50 VNB N_A_642_392#_c_723_n 0.0346804f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_642_392#_c_724_n 0.012237f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.615
cc_52 VNB N_A_642_392#_c_725_n 0.00569027f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_642_392#_c_726_n 0.0131155f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_642_392#_c_727_n 0.00719536f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_642_392#_c_728_n 0.00952616f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_RESET_B_c_811_n 0.0169211f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.45
cc_57 VNB N_RESET_B_c_812_n 0.0334739f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_RESET_B_c_813_n 0.00980122f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.615
cc_59 VNB N_A_1342_74#_M1020_g 0.0274092f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_1342_74#_c_844_n 0.0384415f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.615
cc_61 VNB N_A_1342_74#_c_845_n 0.00331897f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.615
cc_62 VNB N_A_1342_74#_c_846_n 0.00745708f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_1342_74#_c_847_n 0.00729284f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_1342_74#_c_848_n 0.00133875f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VPWR_c_901_n 0.342803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_Q_c_992_n 0.00885771f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_Q_c_993_n 0.013309f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.615
cc_68 VNB N_Q_c_994_n 0.00547807f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_Q_N_c_1030_n 0.029039f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.615
cc_70 VNB Q_N 0.0232158f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB Q_N 0.00662967f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1052_n 0.037441f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1053_n 0.0221825f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1054_n 0.00647919f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1055_n 0.00712978f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1056_n 0.0296399f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1057_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1058_n 0.0206435f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1059_n 0.0373847f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1060_n 0.0393212f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1061_n 0.0345892f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1062_n 0.0193536f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1063_n 0.478218f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1064_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1065_n 0.0180279f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1066_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1067_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VPB N_D_c_159_n 0.0451535f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.915
cc_89 VPB D 0.00137225f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_90 VPB N_GATE_c_191_n 0.0421514f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.915
cc_91 VPB GATE 0.0015683f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_92 VPB N_A_226_104#_c_226_n 0.0345729f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.615
cc_93 VPB N_A_226_104#_c_239_n 0.0147131f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB N_A_226_104#_c_240_n 0.0416418f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_95 VPB N_A_226_104#_c_241_n 0.010091f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB N_A_226_104#_M1015_g 0.00175587f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_A_226_104#_c_243_n 0.0101573f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_A_226_104#_c_244_n 0.00437403f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB N_A_226_104#_c_235_n 0.00394788f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 VPB N_A_226_104#_c_237_n 0.0149765f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB N_A_27_142#_c_370_n 0.0363578f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.41
cc_102 VPB N_A_27_142#_c_379_n 0.00947227f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 VPB N_A_27_142#_c_380_n 0.0089607f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB N_A_27_142#_c_381_n 0.0221307f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_105 VPB N_A_27_142#_c_382_n 0.00116019f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_A_27_142#_c_383_n 0.0131772f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB N_A_27_142#_c_376_n 0.0147556f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_A_353_98#_c_465_n 0.0644066f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.615
cc_109 VPB N_A_353_98#_c_458_n 0.00325226f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_110 VPB N_A_353_98#_c_461_n 0.00226155f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_A_353_98#_c_468_n 0.00642419f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_A_353_98#_c_469_n 0.00197776f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_A_353_98#_c_470_n 0.00452839f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_A_353_98#_c_471_n 0.00519173f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_A_823_98#_c_577_n 0.0241914f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.615
cc_116 VPB N_A_823_98#_c_590_n 0.0624523f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.615
cc_117 VPB N_A_823_98#_c_579_n 0.0320213f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_A_823_98#_c_582_n 0.0156586f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_A_823_98#_c_593_n 0.0189233f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_A_823_98#_c_594_n 0.0186498f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_A_823_98#_c_595_n 0.0103861f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_A_823_98#_c_596_n 0.00290171f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_A_823_98#_c_597_n 0.00851415f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_A_823_98#_c_586_n 7.43912e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_A_823_98#_c_599_n 0.00907059f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 VPB N_A_642_392#_c_729_n 0.0175575f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.41
cc_127 VPB N_A_642_392#_c_723_n 0.0148713f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_A_642_392#_c_724_n 0.00704601f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.615
cc_129 VPB N_A_642_392#_c_726_n 0.00986883f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_A_642_392#_c_727_n 2.20751e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_A_642_392#_c_734_n 0.00483148f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_A_642_392#_c_728_n 0.00417831f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_RESET_B_c_812_n 0.0224068f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_A_1342_74#_c_844_n 0.0295319f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.615
cc_135 VPB N_A_1342_74#_c_850_n 0.00598072f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_VPWR_c_902_n 0.0186796f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_VPWR_c_903_n 0.012678f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_904_n 0.00886117f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_905_n 0.00774436f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_140 VPB N_VPWR_c_906_n 0.0435325f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_907_n 0.0431663f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_142 VPB N_VPWR_c_908_n 0.0196813f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_143 VPB N_VPWR_c_909_n 0.0323599f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_144 VPB N_VPWR_c_910_n 0.0192325f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_145 VPB N_VPWR_c_901_n 0.113085f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_146 VPB N_VPWR_c_912_n 0.027025f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_147 VPB N_VPWR_c_913_n 0.00623769f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_148 VPB N_VPWR_c_914_n 0.0231504f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_149 VPB N_VPWR_c_915_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_150 VPB N_VPWR_c_916_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_151 VPB N_Q_c_995_n 0.00301309f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_152 VPB N_Q_c_994_n 0.00597653f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_153 VPB Q 0.0127496f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_154 VPB N_Q_N_c_1033_n 0.0409189f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_155 VPB N_Q_N_c_1034_n 0.0124896f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_156 VPB N_Q_N_c_1030_n 0.00765777f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.615
cc_157 N_D_M1001_g N_GATE_M1016_g 0.0137684f $X=0.495 $Y=0.985 $X2=0 $Y2=0
cc_158 N_D_c_159_n N_GATE_c_191_n 0.0498165f $X=0.505 $Y=1.915 $X2=0 $Y2=0
cc_159 D N_GATE_c_191_n 0.00109805f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_160 N_D_c_159_n GATE 3.77615e-19 $X=0.505 $Y=1.915 $X2=0 $Y2=0
cc_161 D GATE 0.0264532f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_162 N_D_c_159_n N_A_226_104#_c_243_n 0.00108177f $X=0.505 $Y=1.915 $X2=0
+ $Y2=0
cc_163 N_D_M1001_g N_A_27_142#_c_374_n 0.00684784f $X=0.495 $Y=0.985 $X2=0 $Y2=0
cc_164 N_D_c_159_n N_A_27_142#_c_379_n 0.00620811f $X=0.505 $Y=1.915 $X2=0 $Y2=0
cc_165 N_D_c_159_n N_A_27_142#_c_380_n 0.0140459f $X=0.505 $Y=1.915 $X2=0 $Y2=0
cc_166 D N_A_27_142#_c_380_n 0.0087727f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_167 N_D_c_159_n N_A_27_142#_c_381_n 0.00765878f $X=0.505 $Y=1.915 $X2=0 $Y2=0
cc_168 N_D_M1001_g N_A_27_142#_c_375_n 0.00477757f $X=0.495 $Y=0.985 $X2=0 $Y2=0
cc_169 N_D_c_159_n N_A_27_142#_c_375_n 2.25073e-19 $X=0.505 $Y=1.915 $X2=0 $Y2=0
cc_170 D N_A_27_142#_c_375_n 7.1032e-19 $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_171 N_D_c_159_n N_A_27_142#_c_383_n 0.00519173f $X=0.505 $Y=1.915 $X2=0 $Y2=0
cc_172 D N_A_27_142#_c_383_n 6.56837e-19 $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_173 N_D_M1001_g N_A_27_142#_c_376_n 0.00415844f $X=0.495 $Y=0.985 $X2=0 $Y2=0
cc_174 N_D_c_159_n N_A_27_142#_c_376_n 0.0126706f $X=0.505 $Y=1.915 $X2=0 $Y2=0
cc_175 D N_A_27_142#_c_376_n 0.0249896f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_176 N_D_c_159_n N_VPWR_c_902_n 0.0043785f $X=0.505 $Y=1.915 $X2=0 $Y2=0
cc_177 N_D_c_159_n N_VPWR_c_901_n 0.00505379f $X=0.505 $Y=1.915 $X2=0 $Y2=0
cc_178 N_D_c_159_n N_VPWR_c_912_n 0.00475032f $X=0.505 $Y=1.915 $X2=0 $Y2=0
cc_179 N_D_M1001_g N_VGND_c_1052_n 0.00673272f $X=0.495 $Y=0.985 $X2=0 $Y2=0
cc_180 N_D_c_159_n N_VGND_c_1052_n 0.0032381f $X=0.505 $Y=1.915 $X2=0 $Y2=0
cc_181 D N_VGND_c_1052_n 0.0152608f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_182 N_D_M1001_g N_VGND_c_1058_n 0.00360349f $X=0.495 $Y=0.985 $X2=0 $Y2=0
cc_183 N_D_M1001_g N_VGND_c_1063_n 0.00446563f $X=0.495 $Y=0.985 $X2=0 $Y2=0
cc_184 N_GATE_M1016_g N_A_226_104#_c_228_n 0.0048812f $X=1.055 $Y=0.89 $X2=0
+ $Y2=0
cc_185 N_GATE_c_191_n N_A_226_104#_c_243_n 0.0085111f $X=1.125 $Y=1.915 $X2=0
+ $Y2=0
cc_186 GATE N_A_226_104#_c_243_n 0.0084864f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_187 N_GATE_c_191_n N_A_226_104#_c_244_n 0.00593692f $X=1.125 $Y=1.915 $X2=0
+ $Y2=0
cc_188 N_GATE_M1016_g N_A_226_104#_c_234_n 0.0102394f $X=1.055 $Y=0.89 $X2=0
+ $Y2=0
cc_189 N_GATE_c_191_n N_A_226_104#_c_234_n 0.00285212f $X=1.125 $Y=1.915 $X2=0
+ $Y2=0
cc_190 GATE N_A_226_104#_c_234_n 0.0100357f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_191 N_GATE_c_191_n N_A_226_104#_c_235_n 0.00124686f $X=1.125 $Y=1.915 $X2=0
+ $Y2=0
cc_192 GATE N_A_226_104#_c_235_n 0.0262997f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_193 N_GATE_M1016_g N_A_226_104#_c_236_n 0.00457461f $X=1.055 $Y=0.89 $X2=0
+ $Y2=0
cc_194 N_GATE_M1016_g N_A_226_104#_c_237_n 7.24666e-19 $X=1.055 $Y=0.89 $X2=0
+ $Y2=0
cc_195 N_GATE_c_191_n N_A_226_104#_c_237_n 0.0165331f $X=1.125 $Y=1.915 $X2=0
+ $Y2=0
cc_196 GATE N_A_226_104#_c_237_n 3.29883e-19 $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_197 N_GATE_c_191_n N_A_27_142#_c_380_n 0.0172965f $X=1.125 $Y=1.915 $X2=0
+ $Y2=0
cc_198 GATE N_A_27_142#_c_380_n 0.00457372f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_199 N_GATE_c_191_n N_A_27_142#_c_381_n 7.68435e-19 $X=1.125 $Y=1.915 $X2=0
+ $Y2=0
cc_200 N_GATE_c_191_n N_A_27_142#_c_383_n 0.00183087f $X=1.125 $Y=1.915 $X2=0
+ $Y2=0
cc_201 N_GATE_c_191_n N_A_353_98#_c_471_n 3.77523e-19 $X=1.125 $Y=1.915 $X2=0
+ $Y2=0
cc_202 N_GATE_c_191_n N_VPWR_c_902_n 0.00663705f $X=1.125 $Y=1.915 $X2=0 $Y2=0
cc_203 N_GATE_c_191_n N_VPWR_c_906_n 0.00487664f $X=1.125 $Y=1.915 $X2=0 $Y2=0
cc_204 N_GATE_c_191_n N_VPWR_c_901_n 0.00505379f $X=1.125 $Y=1.915 $X2=0 $Y2=0
cc_205 N_GATE_M1016_g N_VGND_c_1052_n 0.00584542f $X=1.055 $Y=0.89 $X2=0 $Y2=0
cc_206 N_GATE_M1016_g N_VGND_c_1059_n 0.00475172f $X=1.055 $Y=0.89 $X2=0 $Y2=0
cc_207 N_GATE_M1016_g N_VGND_c_1063_n 0.00499434f $X=1.055 $Y=0.89 $X2=0 $Y2=0
cc_208 N_A_226_104#_c_226_n N_A_27_142#_c_370_n 0.0452168f $X=2.205 $Y=1.885
+ $X2=0 $Y2=0
cc_209 N_A_226_104#_c_239_n N_A_27_142#_c_370_n 0.0547763f $X=3.135 $Y=1.885
+ $X2=0 $Y2=0
cc_210 N_A_226_104#_c_241_n N_A_27_142#_c_370_n 0.0119964f $X=3.225 $Y=1.765
+ $X2=0 $Y2=0
cc_211 N_A_226_104#_c_226_n N_A_27_142#_c_371_n 0.00502555f $X=2.205 $Y=1.885
+ $X2=0 $Y2=0
cc_212 N_A_226_104#_M1002_g N_A_27_142#_c_372_n 0.0210344f $X=2.19 $Y=0.86 $X2=0
+ $Y2=0
cc_213 N_A_226_104#_c_230_n N_A_27_142#_c_372_n 0.00969944f $X=2.82 $Y=0.665
+ $X2=0 $Y2=0
cc_214 N_A_226_104#_c_231_n N_A_27_142#_c_372_n 0.00983971f $X=2.99 $Y=0.382
+ $X2=0 $Y2=0
cc_215 N_A_226_104#_c_232_n N_A_27_142#_c_372_n 2.18501e-19 $X=3.74 $Y=0.345
+ $X2=0 $Y2=0
cc_216 N_A_226_104#_M1002_g N_A_27_142#_c_373_n 0.00502555f $X=2.19 $Y=0.86
+ $X2=0 $Y2=0
cc_217 N_A_226_104#_M1018_d N_A_27_142#_c_380_n 0.0107584f $X=1.2 $Y=1.99 $X2=0
+ $Y2=0
cc_218 N_A_226_104#_c_226_n N_A_27_142#_c_380_n 0.0160955f $X=2.205 $Y=1.885
+ $X2=0 $Y2=0
cc_219 N_A_226_104#_c_243_n N_A_27_142#_c_380_n 0.0313572f $X=1.475 $Y=2.095
+ $X2=0 $Y2=0
cc_220 N_A_226_104#_c_235_n N_A_27_142#_c_380_n 0.0046631f $X=1.71 $Y=1.585
+ $X2=0 $Y2=0
cc_221 N_A_226_104#_c_237_n N_A_27_142#_c_380_n 0.00116795f $X=1.71 $Y=1.495
+ $X2=0 $Y2=0
cc_222 N_A_226_104#_c_226_n N_A_27_142#_c_382_n 0.00650368f $X=2.205 $Y=1.885
+ $X2=0 $Y2=0
cc_223 N_A_226_104#_c_239_n N_A_27_142#_c_382_n 2.88046e-19 $X=3.135 $Y=1.885
+ $X2=0 $Y2=0
cc_224 N_A_226_104#_c_226_n N_A_27_142#_c_377_n 0.00120511f $X=2.205 $Y=1.885
+ $X2=0 $Y2=0
cc_225 N_A_226_104#_c_230_n N_A_353_98#_M1002_s 0.00970401f $X=2.82 $Y=0.665
+ $X2=-0.19 $Y2=-0.245
cc_226 N_A_226_104#_c_239_n N_A_353_98#_c_465_n 0.0205927f $X=3.135 $Y=1.885
+ $X2=0 $Y2=0
cc_227 N_A_226_104#_c_240_n N_A_353_98#_c_465_n 0.018086f $X=3.725 $Y=1.765
+ $X2=0 $Y2=0
cc_228 N_A_226_104#_c_224_n N_A_353_98#_c_458_n 0.00598126f $X=2.115 $Y=1.495
+ $X2=0 $Y2=0
cc_229 N_A_226_104#_M1002_g N_A_353_98#_c_458_n 0.00474446f $X=2.19 $Y=0.86
+ $X2=0 $Y2=0
cc_230 N_A_226_104#_c_226_n N_A_353_98#_c_458_n 0.0140246f $X=2.205 $Y=1.885
+ $X2=0 $Y2=0
cc_231 N_A_226_104#_c_244_n N_A_353_98#_c_458_n 0.00789954f $X=1.56 $Y=1.97
+ $X2=0 $Y2=0
cc_232 N_A_226_104#_c_235_n N_A_353_98#_c_458_n 0.02461f $X=1.71 $Y=1.585 $X2=0
+ $Y2=0
cc_233 N_A_226_104#_c_236_n N_A_353_98#_c_458_n 0.00496061f $X=1.675 $Y=1.42
+ $X2=0 $Y2=0
cc_234 N_A_226_104#_c_237_n N_A_353_98#_c_458_n 0.00102115f $X=1.71 $Y=1.495
+ $X2=0 $Y2=0
cc_235 N_A_226_104#_M1002_g N_A_353_98#_c_459_n 0.0066394f $X=2.19 $Y=0.86 $X2=0
+ $Y2=0
cc_236 N_A_226_104#_c_226_n N_A_353_98#_c_459_n 0.00106272f $X=2.205 $Y=1.885
+ $X2=0 $Y2=0
cc_237 N_A_226_104#_c_230_n N_A_353_98#_c_459_n 0.0202971f $X=2.82 $Y=0.665
+ $X2=0 $Y2=0
cc_238 N_A_226_104#_c_231_n N_A_353_98#_c_459_n 0.0060371f $X=2.99 $Y=0.382
+ $X2=0 $Y2=0
cc_239 N_A_226_104#_c_232_n N_A_353_98#_c_459_n 4.49052e-19 $X=3.74 $Y=0.345
+ $X2=0 $Y2=0
cc_240 N_A_226_104#_M1002_g N_A_353_98#_c_460_n 0.00975883f $X=2.19 $Y=0.86
+ $X2=0 $Y2=0
cc_241 N_A_226_104#_c_229_n N_A_353_98#_c_460_n 0.0274006f $X=1.415 $Y=1.05
+ $X2=0 $Y2=0
cc_242 N_A_226_104#_c_230_n N_A_353_98#_c_460_n 0.0255279f $X=2.82 $Y=0.665
+ $X2=0 $Y2=0
cc_243 N_A_226_104#_c_234_n N_A_353_98#_c_460_n 0.00241323f $X=1.415 $Y=1.28
+ $X2=0 $Y2=0
cc_244 N_A_226_104#_c_235_n N_A_353_98#_c_460_n 0.00391614f $X=1.71 $Y=1.585
+ $X2=0 $Y2=0
cc_245 N_A_226_104#_c_237_n N_A_353_98#_c_460_n 0.00670506f $X=1.71 $Y=1.495
+ $X2=0 $Y2=0
cc_246 N_A_226_104#_c_239_n N_A_353_98#_c_461_n 0.00207212f $X=3.135 $Y=1.885
+ $X2=0 $Y2=0
cc_247 N_A_226_104#_c_241_n N_A_353_98#_c_461_n 0.0068682f $X=3.225 $Y=1.765
+ $X2=0 $Y2=0
cc_248 N_A_226_104#_M1015_g N_A_353_98#_c_461_n 8.96735e-19 $X=3.8 $Y=0.83 $X2=0
+ $Y2=0
cc_249 N_A_226_104#_c_239_n N_A_353_98#_c_468_n 0.0132105f $X=3.135 $Y=1.885
+ $X2=0 $Y2=0
cc_250 N_A_226_104#_c_239_n N_A_353_98#_c_470_n 5.066e-19 $X=3.135 $Y=1.885
+ $X2=0 $Y2=0
cc_251 N_A_226_104#_c_240_n N_A_353_98#_c_470_n 7.29778e-19 $X=3.725 $Y=1.765
+ $X2=0 $Y2=0
cc_252 N_A_226_104#_c_224_n N_A_353_98#_c_471_n 0.00521549f $X=2.115 $Y=1.495
+ $X2=0 $Y2=0
cc_253 N_A_226_104#_c_226_n N_A_353_98#_c_471_n 0.00667592f $X=2.205 $Y=1.885
+ $X2=0 $Y2=0
cc_254 N_A_226_104#_c_243_n N_A_353_98#_c_471_n 0.0217728f $X=1.475 $Y=2.095
+ $X2=0 $Y2=0
cc_255 N_A_226_104#_c_244_n N_A_353_98#_c_471_n 0.00230777f $X=1.56 $Y=1.97
+ $X2=0 $Y2=0
cc_256 N_A_226_104#_c_235_n N_A_353_98#_c_471_n 0.00425849f $X=1.71 $Y=1.585
+ $X2=0 $Y2=0
cc_257 N_A_226_104#_c_237_n N_A_353_98#_c_471_n 4.22751e-19 $X=1.71 $Y=1.495
+ $X2=0 $Y2=0
cc_258 N_A_226_104#_c_239_n N_A_353_98#_c_506_n 0.00945501f $X=3.135 $Y=1.885
+ $X2=0 $Y2=0
cc_259 N_A_226_104#_c_241_n N_A_353_98#_c_462_n 0.00117082f $X=3.225 $Y=1.765
+ $X2=0 $Y2=0
cc_260 N_A_226_104#_M1015_g N_A_353_98#_c_462_n 4.00213e-19 $X=3.8 $Y=0.83 $X2=0
+ $Y2=0
cc_261 N_A_226_104#_c_232_n N_A_353_98#_c_462_n 0.00446145f $X=3.74 $Y=0.345
+ $X2=0 $Y2=0
cc_262 N_A_226_104#_c_241_n N_A_353_98#_c_463_n 0.0208047f $X=3.225 $Y=1.765
+ $X2=0 $Y2=0
cc_263 N_A_226_104#_M1015_g N_A_353_98#_c_463_n 0.0113395f $X=3.8 $Y=0.83 $X2=0
+ $Y2=0
cc_264 N_A_226_104#_M1015_g N_A_353_98#_c_464_n 0.0138701f $X=3.8 $Y=0.83 $X2=0
+ $Y2=0
cc_265 N_A_226_104#_c_231_n N_A_353_98#_c_464_n 0.00506575f $X=2.99 $Y=0.382
+ $X2=0 $Y2=0
cc_266 N_A_226_104#_c_232_n N_A_353_98#_c_464_n 0.013663f $X=3.74 $Y=0.345 $X2=0
+ $Y2=0
cc_267 N_A_226_104#_c_233_n N_A_353_98#_c_464_n 0.00778027f $X=3.74 $Y=0.345
+ $X2=0 $Y2=0
cc_268 N_A_226_104#_M1015_g N_A_823_98#_c_576_n 0.0388657f $X=3.8 $Y=0.83 $X2=0
+ $Y2=0
cc_269 N_A_226_104#_c_233_n N_A_823_98#_c_576_n 0.00120024f $X=3.74 $Y=0.345
+ $X2=0 $Y2=0
cc_270 N_A_226_104#_M1015_g N_A_823_98#_c_577_n 0.0206399f $X=3.8 $Y=0.83 $X2=0
+ $Y2=0
cc_271 N_A_226_104#_c_232_n N_A_642_392#_M1008_d 0.00211965f $X=3.74 $Y=0.345
+ $X2=-0.19 $Y2=-0.245
cc_272 N_A_226_104#_M1015_g N_A_642_392#_c_737_n 0.00898495f $X=3.8 $Y=0.83
+ $X2=0 $Y2=0
cc_273 N_A_226_104#_c_231_n N_A_642_392#_c_737_n 0.00265955f $X=2.99 $Y=0.382
+ $X2=0 $Y2=0
cc_274 N_A_226_104#_c_232_n N_A_642_392#_c_737_n 0.0307459f $X=3.74 $Y=0.345
+ $X2=0 $Y2=0
cc_275 N_A_226_104#_c_233_n N_A_642_392#_c_737_n 0.00324473f $X=3.74 $Y=0.345
+ $X2=0 $Y2=0
cc_276 N_A_226_104#_c_240_n N_A_642_392#_c_725_n 0.00150476f $X=3.725 $Y=1.765
+ $X2=0 $Y2=0
cc_277 N_A_226_104#_M1015_g N_A_642_392#_c_725_n 0.0200584f $X=3.8 $Y=0.83 $X2=0
+ $Y2=0
cc_278 N_A_226_104#_c_240_n N_A_642_392#_c_726_n 0.00411388f $X=3.725 $Y=1.765
+ $X2=0 $Y2=0
cc_279 N_A_226_104#_M1015_g N_A_642_392#_c_726_n 0.00645726f $X=3.8 $Y=0.83
+ $X2=0 $Y2=0
cc_280 N_A_226_104#_c_240_n N_A_642_392#_c_727_n 0.0168023f $X=3.725 $Y=1.765
+ $X2=0 $Y2=0
cc_281 N_A_226_104#_M1015_g N_A_642_392#_c_727_n 9.72505e-19 $X=3.8 $Y=0.83
+ $X2=0 $Y2=0
cc_282 N_A_226_104#_c_239_n N_A_642_392#_c_747_n 0.0038846f $X=3.135 $Y=1.885
+ $X2=0 $Y2=0
cc_283 N_A_226_104#_c_240_n N_A_642_392#_c_747_n 0.00238029f $X=3.725 $Y=1.765
+ $X2=0 $Y2=0
cc_284 N_A_226_104#_c_239_n N_A_642_392#_c_734_n 0.00613548f $X=3.135 $Y=1.885
+ $X2=0 $Y2=0
cc_285 N_A_226_104#_c_240_n N_A_642_392#_c_734_n 0.00595874f $X=3.725 $Y=1.765
+ $X2=0 $Y2=0
cc_286 N_A_226_104#_c_241_n N_A_642_392#_c_734_n 9.46059e-19 $X=3.225 $Y=1.765
+ $X2=0 $Y2=0
cc_287 N_A_226_104#_c_226_n N_VPWR_c_903_n 0.00560625f $X=2.205 $Y=1.885 $X2=0
+ $Y2=0
cc_288 N_A_226_104#_c_239_n N_VPWR_c_903_n 2.70003e-19 $X=3.135 $Y=1.885 $X2=0
+ $Y2=0
cc_289 N_A_226_104#_c_226_n N_VPWR_c_906_n 0.00469064f $X=2.205 $Y=1.885 $X2=0
+ $Y2=0
cc_290 N_A_226_104#_c_239_n N_VPWR_c_907_n 0.00278271f $X=3.135 $Y=1.885 $X2=0
+ $Y2=0
cc_291 N_A_226_104#_c_226_n N_VPWR_c_901_n 0.0049649f $X=2.205 $Y=1.885 $X2=0
+ $Y2=0
cc_292 N_A_226_104#_c_239_n N_VPWR_c_901_n 0.0035428f $X=3.135 $Y=1.885 $X2=0
+ $Y2=0
cc_293 N_A_226_104#_c_230_n N_VGND_M1002_d 0.00912757f $X=2.82 $Y=0.665 $X2=0
+ $Y2=0
cc_294 N_A_226_104#_c_228_n N_VGND_c_1052_n 0.00131648f $X=1.415 $Y=0.75 $X2=0
+ $Y2=0
cc_295 N_A_226_104#_c_234_n N_VGND_c_1052_n 0.00131206f $X=1.415 $Y=1.28 $X2=0
+ $Y2=0
cc_296 N_A_226_104#_M1015_g N_VGND_c_1053_n 0.0019797f $X=3.8 $Y=0.83 $X2=0
+ $Y2=0
cc_297 N_A_226_104#_c_232_n N_VGND_c_1053_n 0.01269f $X=3.74 $Y=0.345 $X2=0
+ $Y2=0
cc_298 N_A_226_104#_c_233_n N_VGND_c_1053_n 0.00337434f $X=3.74 $Y=0.345 $X2=0
+ $Y2=0
cc_299 N_A_226_104#_M1002_g N_VGND_c_1059_n 0.00374721f $X=2.19 $Y=0.86 $X2=0
+ $Y2=0
cc_300 N_A_226_104#_c_228_n N_VGND_c_1059_n 0.0127217f $X=1.415 $Y=0.75 $X2=0
+ $Y2=0
cc_301 N_A_226_104#_c_230_n N_VGND_c_1059_n 0.0123272f $X=2.82 $Y=0.665 $X2=0
+ $Y2=0
cc_302 N_A_226_104#_c_230_n N_VGND_c_1060_n 0.00276577f $X=2.82 $Y=0.665 $X2=0
+ $Y2=0
cc_303 N_A_226_104#_c_231_n N_VGND_c_1060_n 0.0117598f $X=2.99 $Y=0.382 $X2=0
+ $Y2=0
cc_304 N_A_226_104#_c_232_n N_VGND_c_1060_n 0.0596213f $X=3.74 $Y=0.345 $X2=0
+ $Y2=0
cc_305 N_A_226_104#_c_233_n N_VGND_c_1060_n 0.00653686f $X=3.74 $Y=0.345 $X2=0
+ $Y2=0
cc_306 N_A_226_104#_M1002_g N_VGND_c_1063_n 0.00508379f $X=2.19 $Y=0.86 $X2=0
+ $Y2=0
cc_307 N_A_226_104#_c_228_n N_VGND_c_1063_n 0.0153896f $X=1.415 $Y=0.75 $X2=0
+ $Y2=0
cc_308 N_A_226_104#_c_230_n N_VGND_c_1063_n 0.0266335f $X=2.82 $Y=0.665 $X2=0
+ $Y2=0
cc_309 N_A_226_104#_c_231_n N_VGND_c_1063_n 0.00647831f $X=2.99 $Y=0.382 $X2=0
+ $Y2=0
cc_310 N_A_226_104#_c_232_n N_VGND_c_1063_n 0.0332028f $X=3.74 $Y=0.345 $X2=0
+ $Y2=0
cc_311 N_A_226_104#_c_233_n N_VGND_c_1063_n 0.0102677f $X=3.74 $Y=0.345 $X2=0
+ $Y2=0
cc_312 N_A_226_104#_M1002_g N_VGND_c_1065_n 0.0014541f $X=2.19 $Y=0.86 $X2=0
+ $Y2=0
cc_313 N_A_226_104#_c_230_n N_VGND_c_1065_n 0.0244722f $X=2.82 $Y=0.665 $X2=0
+ $Y2=0
cc_314 N_A_226_104#_c_231_n N_VGND_c_1065_n 0.0113011f $X=2.99 $Y=0.382 $X2=0
+ $Y2=0
cc_315 N_A_226_104#_c_231_n A_571_80# 0.00407179f $X=2.99 $Y=0.382 $X2=-0.19
+ $Y2=-0.245
cc_316 N_A_226_104#_c_232_n A_571_80# 5.69087e-19 $X=3.74 $Y=0.345 $X2=-0.19
+ $Y2=-0.245
cc_317 N_A_27_142#_c_380_n N_A_353_98#_M1014_s 0.0080688f $X=2.505 $Y=2.475
+ $X2=0 $Y2=0
cc_318 N_A_27_142#_c_370_n N_A_353_98#_c_458_n 0.00118939f $X=2.745 $Y=1.885
+ $X2=0 $Y2=0
cc_319 N_A_27_142#_c_371_n N_A_353_98#_c_458_n 8.80243e-19 $X=2.76 $Y=1.47 $X2=0
+ $Y2=0
cc_320 N_A_27_142#_c_377_n N_A_353_98#_c_458_n 0.0220582f $X=2.67 $Y=1.635 $X2=0
+ $Y2=0
cc_321 N_A_27_142#_c_370_n N_A_353_98#_c_459_n 0.00126003f $X=2.745 $Y=1.885
+ $X2=0 $Y2=0
cc_322 N_A_27_142#_c_371_n N_A_353_98#_c_459_n 0.00324086f $X=2.76 $Y=1.47 $X2=0
+ $Y2=0
cc_323 N_A_27_142#_c_373_n N_A_353_98#_c_459_n 0.00869943f $X=2.77 $Y=1.265
+ $X2=0 $Y2=0
cc_324 N_A_27_142#_c_377_n N_A_353_98#_c_459_n 0.0249573f $X=2.67 $Y=1.635 $X2=0
+ $Y2=0
cc_325 N_A_27_142#_c_372_n N_A_353_98#_c_460_n 9.94999e-19 $X=2.77 $Y=1.115
+ $X2=0 $Y2=0
cc_326 N_A_27_142#_c_370_n N_A_353_98#_c_461_n 0.00551206f $X=2.745 $Y=1.885
+ $X2=0 $Y2=0
cc_327 N_A_27_142#_c_382_n N_A_353_98#_c_461_n 0.00712086f $X=2.59 $Y=2.39 $X2=0
+ $Y2=0
cc_328 N_A_27_142#_c_370_n N_A_353_98#_c_469_n 0.00111115f $X=2.745 $Y=1.885
+ $X2=0 $Y2=0
cc_329 N_A_27_142#_c_370_n N_A_353_98#_c_471_n 2.62068e-19 $X=2.745 $Y=1.885
+ $X2=0 $Y2=0
cc_330 N_A_27_142#_c_380_n N_A_353_98#_c_471_n 0.02544f $X=2.505 $Y=2.475 $X2=0
+ $Y2=0
cc_331 N_A_27_142#_c_382_n N_A_353_98#_c_471_n 0.0138942f $X=2.59 $Y=2.39 $X2=0
+ $Y2=0
cc_332 N_A_27_142#_c_371_n N_A_353_98#_c_462_n 0.0050162f $X=2.76 $Y=1.47 $X2=0
+ $Y2=0
cc_333 N_A_27_142#_c_377_n N_A_353_98#_c_462_n 0.0248145f $X=2.67 $Y=1.635 $X2=0
+ $Y2=0
cc_334 N_A_27_142#_c_371_n N_A_353_98#_c_463_n 0.0114717f $X=2.76 $Y=1.47 $X2=0
+ $Y2=0
cc_335 N_A_27_142#_c_373_n N_A_353_98#_c_463_n 0.0310886f $X=2.77 $Y=1.265 $X2=0
+ $Y2=0
cc_336 N_A_27_142#_c_372_n N_A_353_98#_c_464_n 0.0310886f $X=2.77 $Y=1.115 $X2=0
+ $Y2=0
cc_337 N_A_27_142#_c_372_n N_A_642_392#_c_737_n 0.00107367f $X=2.77 $Y=1.115
+ $X2=0 $Y2=0
cc_338 N_A_27_142#_c_380_n N_VPWR_M1021_d 0.0147931f $X=2.505 $Y=2.475 $X2=-0.19
+ $Y2=-0.245
cc_339 N_A_27_142#_c_380_n N_VPWR_M1014_d 0.00967039f $X=2.505 $Y=2.475 $X2=0
+ $Y2=0
cc_340 N_A_27_142#_c_382_n N_VPWR_M1014_d 0.00479677f $X=2.59 $Y=2.39 $X2=0
+ $Y2=0
cc_341 N_A_27_142#_c_380_n N_VPWR_c_902_n 0.0259408f $X=2.505 $Y=2.475 $X2=0
+ $Y2=0
cc_342 N_A_27_142#_c_381_n N_VPWR_c_902_n 0.00816548f $X=0.445 $Y=2.475 $X2=0
+ $Y2=0
cc_343 N_A_27_142#_c_370_n N_VPWR_c_903_n 0.00687706f $X=2.745 $Y=1.885 $X2=0
+ $Y2=0
cc_344 N_A_27_142#_c_380_n N_VPWR_c_903_n 0.0218683f $X=2.505 $Y=2.475 $X2=0
+ $Y2=0
cc_345 N_A_27_142#_c_370_n N_VPWR_c_907_n 0.00413917f $X=2.745 $Y=1.885 $X2=0
+ $Y2=0
cc_346 N_A_27_142#_c_370_n N_VPWR_c_901_n 0.00817239f $X=2.745 $Y=1.885 $X2=0
+ $Y2=0
cc_347 N_A_27_142#_c_380_n N_VPWR_c_901_n 0.0589062f $X=2.505 $Y=2.475 $X2=0
+ $Y2=0
cc_348 N_A_27_142#_c_381_n N_VPWR_c_901_n 0.0118514f $X=0.445 $Y=2.475 $X2=0
+ $Y2=0
cc_349 N_A_27_142#_c_381_n N_VPWR_c_912_n 0.0101564f $X=0.445 $Y=2.475 $X2=0
+ $Y2=0
cc_350 N_A_27_142#_c_374_n N_VGND_c_1052_n 0.02282f $X=0.27 $Y=1.105 $X2=0 $Y2=0
cc_351 N_A_27_142#_c_374_n N_VGND_c_1058_n 0.00622364f $X=0.27 $Y=1.105 $X2=0
+ $Y2=0
cc_352 N_A_27_142#_c_372_n N_VGND_c_1060_n 0.00347067f $X=2.77 $Y=1.115 $X2=0
+ $Y2=0
cc_353 N_A_27_142#_c_372_n N_VGND_c_1063_n 0.00414706f $X=2.77 $Y=1.115 $X2=0
+ $Y2=0
cc_354 N_A_27_142#_c_374_n N_VGND_c_1063_n 0.0100744f $X=0.27 $Y=1.105 $X2=0
+ $Y2=0
cc_355 N_A_27_142#_c_372_n N_VGND_c_1065_n 0.00245071f $X=2.77 $Y=1.115 $X2=0
+ $Y2=0
cc_356 N_A_353_98#_c_465_n N_A_823_98#_c_590_n 0.0332545f $X=3.69 $Y=2.465 $X2=0
+ $Y2=0
cc_357 N_A_353_98#_c_468_n N_A_823_98#_c_590_n 0.00173515f $X=3.685 $Y=2.99
+ $X2=0 $Y2=0
cc_358 N_A_353_98#_c_470_n N_A_823_98#_c_590_n 0.00938739f $X=3.85 $Y=2.215
+ $X2=0 $Y2=0
cc_359 N_A_353_98#_c_465_n N_A_823_98#_c_595_n 9.76153e-19 $X=3.69 $Y=2.465
+ $X2=0 $Y2=0
cc_360 N_A_353_98#_c_470_n N_A_823_98#_c_595_n 0.0181165f $X=3.85 $Y=2.215 $X2=0
+ $Y2=0
cc_361 N_A_353_98#_c_468_n N_A_642_392#_M1010_d 0.004439f $X=3.685 $Y=2.99 $X2=0
+ $Y2=0
cc_362 N_A_353_98#_c_462_n N_A_642_392#_c_737_n 0.0141269f $X=3.2 $Y=1.215 $X2=0
+ $Y2=0
cc_363 N_A_353_98#_c_463_n N_A_642_392#_c_737_n 0.0010954f $X=3.23 $Y=1.315
+ $X2=0 $Y2=0
cc_364 N_A_353_98#_c_464_n N_A_642_392#_c_737_n 0.00939294f $X=3.23 $Y=1.15
+ $X2=0 $Y2=0
cc_365 N_A_353_98#_c_461_n N_A_642_392#_c_725_n 0.00700637f $X=3.09 $Y=1.97
+ $X2=0 $Y2=0
cc_366 N_A_353_98#_c_462_n N_A_642_392#_c_725_n 0.0250855f $X=3.2 $Y=1.215 $X2=0
+ $Y2=0
cc_367 N_A_353_98#_c_463_n N_A_642_392#_c_725_n 0.00224196f $X=3.23 $Y=1.315
+ $X2=0 $Y2=0
cc_368 N_A_353_98#_c_464_n N_A_642_392#_c_725_n 0.00309916f $X=3.23 $Y=1.15
+ $X2=0 $Y2=0
cc_369 N_A_353_98#_c_465_n N_A_642_392#_c_726_n 9.19261e-19 $X=3.69 $Y=2.465
+ $X2=0 $Y2=0
cc_370 N_A_353_98#_c_465_n N_A_642_392#_c_727_n 8.6097e-19 $X=3.69 $Y=2.465
+ $X2=0 $Y2=0
cc_371 N_A_353_98#_c_461_n N_A_642_392#_c_727_n 0.0131205f $X=3.09 $Y=1.97 $X2=0
+ $Y2=0
cc_372 N_A_353_98#_c_470_n N_A_642_392#_c_727_n 0.0200797f $X=3.85 $Y=2.215
+ $X2=0 $Y2=0
cc_373 N_A_353_98#_c_462_n N_A_642_392#_c_727_n 0.00371746f $X=3.2 $Y=1.215
+ $X2=0 $Y2=0
cc_374 N_A_353_98#_c_465_n N_A_642_392#_c_747_n 0.00221007f $X=3.69 $Y=2.465
+ $X2=0 $Y2=0
cc_375 N_A_353_98#_c_468_n N_A_642_392#_c_747_n 0.0193955f $X=3.685 $Y=2.99
+ $X2=0 $Y2=0
cc_376 N_A_353_98#_c_465_n N_A_642_392#_c_734_n 0.00376484f $X=3.69 $Y=2.465
+ $X2=0 $Y2=0
cc_377 N_A_353_98#_c_461_n N_A_642_392#_c_734_n 0.0106062f $X=3.09 $Y=1.97 $X2=0
+ $Y2=0
cc_378 N_A_353_98#_c_470_n N_A_642_392#_c_734_n 0.0516937f $X=3.85 $Y=2.215
+ $X2=0 $Y2=0
cc_379 N_A_353_98#_c_506_n N_A_642_392#_c_734_n 0.0124377f $X=3.09 $Y=2.055
+ $X2=0 $Y2=0
cc_380 N_A_353_98#_c_469_n N_VPWR_c_903_n 0.0117385f $X=3.025 $Y=2.99 $X2=0
+ $Y2=0
cc_381 N_A_353_98#_c_465_n N_VPWR_c_907_n 0.00278193f $X=3.69 $Y=2.465 $X2=0
+ $Y2=0
cc_382 N_A_353_98#_c_468_n N_VPWR_c_907_n 0.0651631f $X=3.685 $Y=2.99 $X2=0
+ $Y2=0
cc_383 N_A_353_98#_c_469_n N_VPWR_c_907_n 0.0121867f $X=3.025 $Y=2.99 $X2=0
+ $Y2=0
cc_384 N_A_353_98#_c_465_n N_VPWR_c_901_n 0.00356387f $X=3.69 $Y=2.465 $X2=0
+ $Y2=0
cc_385 N_A_353_98#_c_468_n N_VPWR_c_901_n 0.0362648f $X=3.685 $Y=2.99 $X2=0
+ $Y2=0
cc_386 N_A_353_98#_c_469_n N_VPWR_c_901_n 0.00660921f $X=3.025 $Y=2.99 $X2=0
+ $Y2=0
cc_387 N_A_353_98#_c_465_n N_VPWR_c_914_n 4.0437e-19 $X=3.69 $Y=2.465 $X2=0
+ $Y2=0
cc_388 N_A_353_98#_c_468_n N_VPWR_c_914_n 0.00799935f $X=3.685 $Y=2.99 $X2=0
+ $Y2=0
cc_389 N_A_353_98#_c_470_n N_VPWR_c_914_n 0.0109969f $X=3.85 $Y=2.215 $X2=0
+ $Y2=0
cc_390 N_A_353_98#_c_570_p A_564_392# 0.00327032f $X=2.94 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_391 N_A_353_98#_c_506_n A_564_392# 0.00289737f $X=3.09 $Y=2.055 $X2=-0.19
+ $Y2=-0.245
cc_392 N_A_353_98#_c_468_n A_753_508# 9.16612e-19 $X=3.685 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_393 N_A_353_98#_c_470_n A_753_508# 0.00589473f $X=3.85 $Y=2.215 $X2=-0.19
+ $Y2=-0.245
cc_394 N_A_353_98#_c_459_n N_VGND_M1002_d 0.00334301f $X=3.005 $Y=1.215 $X2=0
+ $Y2=0
cc_395 N_A_353_98#_c_464_n N_VGND_c_1060_n 9.29978e-19 $X=3.23 $Y=1.15 $X2=0
+ $Y2=0
cc_396 N_A_823_98#_c_577_n N_A_642_392#_c_729_n 0.00307848f $X=4.3 $Y=1.99 $X2=0
+ $Y2=0
cc_397 N_A_823_98#_c_590_n N_A_642_392#_c_729_n 0.0138232f $X=4.345 $Y=2.465
+ $X2=0 $Y2=0
cc_398 N_A_823_98#_c_596_n N_A_642_392#_c_729_n 3.04524e-19 $X=5.415 $Y=2.4
+ $X2=0 $Y2=0
cc_399 N_A_823_98#_c_599_n N_A_642_392#_c_729_n 0.0215216f $X=5.332 $Y=1.805
+ $X2=0 $Y2=0
cc_400 N_A_823_98#_c_585_n N_A_642_392#_M1019_g 0.0154535f $X=4.965 $Y=0.515
+ $X2=0 $Y2=0
cc_401 N_A_823_98#_c_587_n N_A_642_392#_M1019_g 0.00612197f $X=5.027 $Y=1.13
+ $X2=0 $Y2=0
cc_402 N_A_823_98#_c_588_n N_A_642_392#_M1019_g 0.00748864f $X=5.332 $Y=1.72
+ $X2=0 $Y2=0
cc_403 N_A_823_98#_c_577_n N_A_642_392#_c_723_n 0.0224688f $X=4.3 $Y=1.99 $X2=0
+ $Y2=0
cc_404 N_A_823_98#_c_595_n N_A_642_392#_c_723_n 0.00658112f $X=5.085 $Y=2.155
+ $X2=0 $Y2=0
cc_405 N_A_823_98#_c_587_n N_A_642_392#_c_723_n 0.00805879f $X=5.027 $Y=1.13
+ $X2=0 $Y2=0
cc_406 N_A_823_98#_c_577_n N_A_642_392#_c_724_n 7.78544e-19 $X=4.3 $Y=1.99 $X2=0
+ $Y2=0
cc_407 N_A_823_98#_c_599_n N_A_642_392#_c_724_n 0.00183897f $X=5.332 $Y=1.805
+ $X2=0 $Y2=0
cc_408 N_A_823_98#_c_588_n N_A_642_392#_c_724_n 0.0139553f $X=5.332 $Y=1.72
+ $X2=0 $Y2=0
cc_409 N_A_823_98#_c_576_n N_A_642_392#_c_737_n 7.06024e-19 $X=4.19 $Y=1.115
+ $X2=0 $Y2=0
cc_410 N_A_823_98#_c_576_n N_A_642_392#_c_725_n 0.00134833f $X=4.19 $Y=1.115
+ $X2=0 $Y2=0
cc_411 N_A_823_98#_c_577_n N_A_642_392#_c_725_n 0.00183254f $X=4.3 $Y=1.99 $X2=0
+ $Y2=0
cc_412 N_A_823_98#_c_577_n N_A_642_392#_c_726_n 0.0132396f $X=4.3 $Y=1.99 $X2=0
+ $Y2=0
cc_413 N_A_823_98#_c_590_n N_A_642_392#_c_726_n 0.00423928f $X=4.345 $Y=2.465
+ $X2=0 $Y2=0
cc_414 N_A_823_98#_c_583_n N_A_642_392#_c_726_n 0.00363508f $X=4.3 $Y=1.19 $X2=0
+ $Y2=0
cc_415 N_A_823_98#_c_595_n N_A_642_392#_c_726_n 0.0266186f $X=5.085 $Y=2.155
+ $X2=0 $Y2=0
cc_416 N_A_823_98#_c_577_n N_A_642_392#_c_728_n 0.00227906f $X=4.3 $Y=1.99 $X2=0
+ $Y2=0
cc_417 N_A_823_98#_c_595_n N_A_642_392#_c_728_n 0.0280515f $X=5.085 $Y=2.155
+ $X2=0 $Y2=0
cc_418 N_A_823_98#_c_587_n N_A_642_392#_c_728_n 0.0080797f $X=5.027 $Y=1.13
+ $X2=0 $Y2=0
cc_419 N_A_823_98#_c_588_n N_A_642_392#_c_728_n 0.0349453f $X=5.332 $Y=1.72
+ $X2=0 $Y2=0
cc_420 N_A_823_98#_M1000_g N_RESET_B_c_811_n 0.0175421f $X=6.08 $Y=0.74
+ $X2=-0.19 $Y2=-0.245
cc_421 N_A_823_98#_c_585_n N_RESET_B_c_811_n 0.00338875f $X=4.965 $Y=0.515
+ $X2=-0.19 $Y2=-0.245
cc_422 N_A_823_98#_M1000_g N_RESET_B_c_812_n 0.0208694f $X=6.08 $Y=0.74 $X2=0
+ $Y2=0
cc_423 N_A_823_98#_c_579_n N_RESET_B_c_812_n 0.0363792f $X=6.14 $Y=1.765 $X2=0
+ $Y2=0
cc_424 N_A_823_98#_c_596_n N_RESET_B_c_812_n 0.00740145f $X=5.415 $Y=2.4 $X2=0
+ $Y2=0
cc_425 N_A_823_98#_c_597_n N_RESET_B_c_812_n 0.014703f $X=6.005 $Y=1.805 $X2=0
+ $Y2=0
cc_426 N_A_823_98#_c_586_n N_RESET_B_c_812_n 0.00191442f $X=6.17 $Y=1.515 $X2=0
+ $Y2=0
cc_427 N_A_823_98#_c_599_n N_RESET_B_c_812_n 0.0115893f $X=5.332 $Y=1.805 $X2=0
+ $Y2=0
cc_428 N_A_823_98#_c_588_n N_RESET_B_c_812_n 0.00146036f $X=5.332 $Y=1.72 $X2=0
+ $Y2=0
cc_429 N_A_823_98#_M1000_g N_RESET_B_c_813_n 0.0025692f $X=6.08 $Y=0.74 $X2=0
+ $Y2=0
cc_430 N_A_823_98#_c_597_n N_RESET_B_c_813_n 0.0157396f $X=6.005 $Y=1.805 $X2=0
+ $Y2=0
cc_431 N_A_823_98#_c_586_n N_RESET_B_c_813_n 0.0127618f $X=6.17 $Y=1.515 $X2=0
+ $Y2=0
cc_432 N_A_823_98#_c_599_n N_RESET_B_c_813_n 0.0131268f $X=5.332 $Y=1.805 $X2=0
+ $Y2=0
cc_433 N_A_823_98#_c_588_n N_RESET_B_c_813_n 0.028157f $X=5.332 $Y=1.72 $X2=0
+ $Y2=0
cc_434 N_A_823_98#_M1012_g N_A_1342_74#_M1020_g 0.0218445f $X=7.07 $Y=0.645
+ $X2=0 $Y2=0
cc_435 N_A_823_98#_M1012_g N_A_1342_74#_c_844_n 0.0181135f $X=7.07 $Y=0.645
+ $X2=0 $Y2=0
cc_436 N_A_823_98#_c_582_n N_A_1342_74#_c_844_n 0.00678052f $X=7.07 $Y=1.89
+ $X2=0 $Y2=0
cc_437 N_A_823_98#_c_593_n N_A_1342_74#_c_844_n 0.0190055f $X=7.15 $Y=2.045
+ $X2=0 $Y2=0
cc_438 N_A_823_98#_c_594_n N_A_1342_74#_c_844_n 0.00531731f $X=7.07 $Y=1.967
+ $X2=0 $Y2=0
cc_439 N_A_823_98#_M1000_g N_A_1342_74#_c_845_n 4.11576e-19 $X=6.08 $Y=0.74
+ $X2=0 $Y2=0
cc_440 N_A_823_98#_M1012_g N_A_1342_74#_c_845_n 0.0163105f $X=7.07 $Y=0.645
+ $X2=0 $Y2=0
cc_441 N_A_823_98#_c_579_n N_A_1342_74#_c_850_n 0.001306f $X=6.14 $Y=1.765 $X2=0
+ $Y2=0
cc_442 N_A_823_98#_c_582_n N_A_1342_74#_c_850_n 0.00843693f $X=7.07 $Y=1.89
+ $X2=0 $Y2=0
cc_443 N_A_823_98#_c_593_n N_A_1342_74#_c_850_n 0.00865733f $X=7.15 $Y=2.045
+ $X2=0 $Y2=0
cc_444 N_A_823_98#_c_594_n N_A_1342_74#_c_850_n 0.00602621f $X=7.07 $Y=1.967
+ $X2=0 $Y2=0
cc_445 N_A_823_98#_M1012_g N_A_1342_74#_c_846_n 0.00653346f $X=7.07 $Y=0.645
+ $X2=0 $Y2=0
cc_446 N_A_823_98#_c_582_n N_A_1342_74#_c_846_n 0.00895789f $X=7.07 $Y=1.89
+ $X2=0 $Y2=0
cc_447 N_A_823_98#_c_584_n N_A_1342_74#_c_846_n 0.00331626f $X=7.07 $Y=1.425
+ $X2=0 $Y2=0
cc_448 N_A_823_98#_c_594_n N_A_1342_74#_c_846_n 0.00342021f $X=7.07 $Y=1.967
+ $X2=0 $Y2=0
cc_449 N_A_823_98#_M1000_g N_A_1342_74#_c_847_n 0.00102563f $X=6.08 $Y=0.74
+ $X2=0 $Y2=0
cc_450 N_A_823_98#_c_580_n N_A_1342_74#_c_847_n 0.00407734f $X=6.995 $Y=1.425
+ $X2=0 $Y2=0
cc_451 N_A_823_98#_M1012_g N_A_1342_74#_c_847_n 0.00739433f $X=7.07 $Y=0.645
+ $X2=0 $Y2=0
cc_452 N_A_823_98#_c_580_n N_A_1342_74#_c_848_n 0.00971855f $X=6.995 $Y=1.425
+ $X2=0 $Y2=0
cc_453 N_A_823_98#_M1012_g N_A_1342_74#_c_848_n 5.74881e-19 $X=7.07 $Y=0.645
+ $X2=0 $Y2=0
cc_454 N_A_823_98#_c_582_n N_A_1342_74#_c_848_n 0.00287486f $X=7.07 $Y=1.89
+ $X2=0 $Y2=0
cc_455 N_A_823_98#_c_584_n N_A_1342_74#_c_848_n 3.53117e-19 $X=7.07 $Y=1.425
+ $X2=0 $Y2=0
cc_456 N_A_823_98#_c_595_n N_VPWR_M1006_d 0.00709733f $X=5.085 $Y=2.155 $X2=0
+ $Y2=0
cc_457 N_A_823_98#_c_597_n N_VPWR_M1023_d 0.00271393f $X=6.005 $Y=1.805 $X2=0
+ $Y2=0
cc_458 N_A_823_98#_c_579_n N_VPWR_c_904_n 0.00800305f $X=6.14 $Y=1.765 $X2=0
+ $Y2=0
cc_459 N_A_823_98#_c_597_n N_VPWR_c_904_n 0.0184553f $X=6.005 $Y=1.805 $X2=0
+ $Y2=0
cc_460 N_A_823_98#_c_599_n N_VPWR_c_904_n 0.0622316f $X=5.332 $Y=1.805 $X2=0
+ $Y2=0
cc_461 N_A_823_98#_c_593_n N_VPWR_c_905_n 0.0183582f $X=7.15 $Y=2.045 $X2=0
+ $Y2=0
cc_462 N_A_823_98#_c_594_n N_VPWR_c_905_n 4.25443e-19 $X=7.07 $Y=1.967 $X2=0
+ $Y2=0
cc_463 N_A_823_98#_c_590_n N_VPWR_c_907_n 0.00415318f $X=4.345 $Y=2.465 $X2=0
+ $Y2=0
cc_464 N_A_823_98#_c_596_n N_VPWR_c_908_n 0.0145938f $X=5.415 $Y=2.4 $X2=0 $Y2=0
cc_465 N_A_823_98#_c_579_n N_VPWR_c_909_n 0.00445602f $X=6.14 $Y=1.765 $X2=0
+ $Y2=0
cc_466 N_A_823_98#_c_593_n N_VPWR_c_909_n 0.00413917f $X=7.15 $Y=2.045 $X2=0
+ $Y2=0
cc_467 N_A_823_98#_c_590_n N_VPWR_c_901_n 0.0085718f $X=4.345 $Y=2.465 $X2=0
+ $Y2=0
cc_468 N_A_823_98#_c_579_n N_VPWR_c_901_n 0.00862233f $X=6.14 $Y=1.765 $X2=0
+ $Y2=0
cc_469 N_A_823_98#_c_593_n N_VPWR_c_901_n 0.00822528f $X=7.15 $Y=2.045 $X2=0
+ $Y2=0
cc_470 N_A_823_98#_c_596_n N_VPWR_c_901_n 0.0120466f $X=5.415 $Y=2.4 $X2=0 $Y2=0
cc_471 N_A_823_98#_c_590_n N_VPWR_c_914_n 0.0121988f $X=4.345 $Y=2.465 $X2=0
+ $Y2=0
cc_472 N_A_823_98#_c_595_n N_VPWR_c_914_n 0.0311617f $X=5.085 $Y=2.155 $X2=0
+ $Y2=0
cc_473 N_A_823_98#_c_596_n N_VPWR_c_914_n 0.00167116f $X=5.415 $Y=2.4 $X2=0
+ $Y2=0
cc_474 N_A_823_98#_c_597_n N_Q_M1003_d 0.00114126f $X=6.005 $Y=1.805 $X2=0 $Y2=0
cc_475 N_A_823_98#_M1000_g N_Q_c_992_n 0.00882067f $X=6.08 $Y=0.74 $X2=0 $Y2=0
cc_476 N_A_823_98#_M1012_g N_Q_c_992_n 0.0019166f $X=7.07 $Y=0.645 $X2=0 $Y2=0
cc_477 N_A_823_98#_M1000_g N_Q_c_993_n 0.00541399f $X=6.08 $Y=0.74 $X2=0 $Y2=0
cc_478 N_A_823_98#_c_579_n N_Q_c_993_n 0.00648394f $X=6.14 $Y=1.765 $X2=0 $Y2=0
cc_479 N_A_823_98#_c_580_n N_Q_c_993_n 8.36337e-19 $X=6.995 $Y=1.425 $X2=0 $Y2=0
cc_480 N_A_823_98#_M1012_g N_Q_c_993_n 9.06455e-19 $X=7.07 $Y=0.645 $X2=0 $Y2=0
cc_481 N_A_823_98#_c_586_n N_Q_c_993_n 0.0155222f $X=6.17 $Y=1.515 $X2=0 $Y2=0
cc_482 N_A_823_98#_c_579_n N_Q_c_995_n 0.00302201f $X=6.14 $Y=1.765 $X2=0 $Y2=0
cc_483 N_A_823_98#_c_580_n N_Q_c_995_n 0.00450563f $X=6.995 $Y=1.425 $X2=0 $Y2=0
cc_484 N_A_823_98#_c_597_n N_Q_c_995_n 0.00626536f $X=6.005 $Y=1.805 $X2=0 $Y2=0
cc_485 N_A_823_98#_M1000_g N_Q_c_994_n 0.00481732f $X=6.08 $Y=0.74 $X2=0 $Y2=0
cc_486 N_A_823_98#_c_579_n N_Q_c_994_n 0.00771233f $X=6.14 $Y=1.765 $X2=0 $Y2=0
cc_487 N_A_823_98#_c_580_n N_Q_c_994_n 0.0135079f $X=6.995 $Y=1.425 $X2=0 $Y2=0
cc_488 N_A_823_98#_M1012_g N_Q_c_994_n 8.40314e-19 $X=7.07 $Y=0.645 $X2=0 $Y2=0
cc_489 N_A_823_98#_c_582_n N_Q_c_994_n 0.00226262f $X=7.07 $Y=1.89 $X2=0 $Y2=0
cc_490 N_A_823_98#_c_597_n N_Q_c_994_n 0.0142023f $X=6.005 $Y=1.805 $X2=0 $Y2=0
cc_491 N_A_823_98#_c_586_n N_Q_c_994_n 0.0273368f $X=6.17 $Y=1.515 $X2=0 $Y2=0
cc_492 N_A_823_98#_c_579_n Q 0.0115149f $X=6.14 $Y=1.765 $X2=0 $Y2=0
cc_493 N_A_823_98#_c_593_n N_Q_N_c_1033_n 5.4831e-19 $X=7.15 $Y=2.045 $X2=0
+ $Y2=0
cc_494 N_A_823_98#_c_582_n N_Q_N_c_1034_n 3.0923e-19 $X=7.07 $Y=1.89 $X2=0 $Y2=0
cc_495 N_A_823_98#_c_594_n N_Q_N_c_1034_n 7.61515e-19 $X=7.07 $Y=1.967 $X2=0
+ $Y2=0
cc_496 N_A_823_98#_c_576_n N_VGND_c_1053_n 0.014495f $X=4.19 $Y=1.115 $X2=0
+ $Y2=0
cc_497 N_A_823_98#_c_583_n N_VGND_c_1053_n 0.00424774f $X=4.3 $Y=1.19 $X2=0
+ $Y2=0
cc_498 N_A_823_98#_c_585_n N_VGND_c_1053_n 0.0490224f $X=4.965 $Y=0.515 $X2=0
+ $Y2=0
cc_499 N_A_823_98#_M1000_g N_VGND_c_1054_n 0.00658431f $X=6.08 $Y=0.74 $X2=0
+ $Y2=0
cc_500 N_A_823_98#_c_585_n N_VGND_c_1054_n 0.0274648f $X=4.965 $Y=0.515 $X2=0
+ $Y2=0
cc_501 N_A_823_98#_M1012_g N_VGND_c_1055_n 0.00628291f $X=7.07 $Y=0.645 $X2=0
+ $Y2=0
cc_502 N_A_823_98#_c_585_n N_VGND_c_1056_n 0.0197679f $X=4.965 $Y=0.515 $X2=0
+ $Y2=0
cc_503 N_A_823_98#_c_576_n N_VGND_c_1060_n 0.00347405f $X=4.19 $Y=1.115 $X2=0
+ $Y2=0
cc_504 N_A_823_98#_M1000_g N_VGND_c_1061_n 0.00434272f $X=6.08 $Y=0.74 $X2=0
+ $Y2=0
cc_505 N_A_823_98#_M1012_g N_VGND_c_1061_n 0.00434272f $X=7.07 $Y=0.645 $X2=0
+ $Y2=0
cc_506 N_A_823_98#_c_576_n N_VGND_c_1063_n 0.00395485f $X=4.19 $Y=1.115 $X2=0
+ $Y2=0
cc_507 N_A_823_98#_M1000_g N_VGND_c_1063_n 0.00826076f $X=6.08 $Y=0.74 $X2=0
+ $Y2=0
cc_508 N_A_823_98#_M1012_g N_VGND_c_1063_n 0.00826076f $X=7.07 $Y=0.645 $X2=0
+ $Y2=0
cc_509 N_A_823_98#_c_585_n N_VGND_c_1063_n 0.0160121f $X=4.965 $Y=0.515 $X2=0
+ $Y2=0
cc_510 N_A_642_392#_M1019_g N_RESET_B_c_811_n 0.047894f $X=5.18 $Y=0.74
+ $X2=-0.19 $Y2=-0.245
cc_511 N_A_642_392#_c_729_n N_RESET_B_c_812_n 0.0090227f $X=5.165 $Y=1.765 $X2=0
+ $Y2=0
cc_512 N_A_642_392#_M1019_g N_RESET_B_c_812_n 0.0208526f $X=5.18 $Y=0.74 $X2=0
+ $Y2=0
cc_513 N_A_642_392#_c_724_n N_RESET_B_c_812_n 0.00996096f $X=5.165 $Y=1.557
+ $X2=0 $Y2=0
cc_514 N_A_642_392#_M1019_g N_RESET_B_c_813_n 0.00213108f $X=5.18 $Y=0.74 $X2=0
+ $Y2=0
cc_515 N_A_642_392#_c_729_n N_VPWR_c_908_n 0.00461464f $X=5.165 $Y=1.765 $X2=0
+ $Y2=0
cc_516 N_A_642_392#_c_729_n N_VPWR_c_901_n 0.00910532f $X=5.165 $Y=1.765 $X2=0
+ $Y2=0
cc_517 N_A_642_392#_c_729_n N_VPWR_c_914_n 0.00437435f $X=5.165 $Y=1.765 $X2=0
+ $Y2=0
cc_518 N_A_642_392#_M1019_g N_VGND_c_1053_n 0.00414178f $X=5.18 $Y=0.74 $X2=0
+ $Y2=0
cc_519 N_A_642_392#_c_737_n N_VGND_c_1053_n 0.00827174f $X=3.58 $Y=0.835 $X2=0
+ $Y2=0
cc_520 N_A_642_392#_c_725_n N_VGND_c_1053_n 0.00300042f $X=3.665 $Y=1.65 $X2=0
+ $Y2=0
cc_521 N_A_642_392#_c_726_n N_VGND_c_1053_n 0.0109917f $X=4.585 $Y=1.735 $X2=0
+ $Y2=0
cc_522 N_A_642_392#_M1019_g N_VGND_c_1054_n 0.00230844f $X=5.18 $Y=0.74 $X2=0
+ $Y2=0
cc_523 N_A_642_392#_M1019_g N_VGND_c_1056_n 0.00292646f $X=5.18 $Y=0.74 $X2=0
+ $Y2=0
cc_524 N_A_642_392#_M1019_g N_VGND_c_1063_n 0.00362778f $X=5.18 $Y=0.74 $X2=0
+ $Y2=0
cc_525 N_RESET_B_c_812_n N_VPWR_c_904_n 0.00713672f $X=5.64 $Y=1.765 $X2=0 $Y2=0
cc_526 N_RESET_B_c_812_n N_VPWR_c_908_n 0.00445602f $X=5.64 $Y=1.765 $X2=0 $Y2=0
cc_527 N_RESET_B_c_812_n N_VPWR_c_901_n 0.00858408f $X=5.64 $Y=1.765 $X2=0 $Y2=0
cc_528 N_RESET_B_c_811_n N_Q_c_993_n 5.64132e-19 $X=5.57 $Y=1.22 $X2=0 $Y2=0
cc_529 N_RESET_B_c_811_n N_VGND_c_1054_n 0.0141029f $X=5.57 $Y=1.22 $X2=0 $Y2=0
cc_530 N_RESET_B_c_812_n N_VGND_c_1054_n 9.00286e-19 $X=5.64 $Y=1.765 $X2=0
+ $Y2=0
cc_531 N_RESET_B_c_813_n N_VGND_c_1054_n 0.0124443f $X=5.63 $Y=1.385 $X2=0 $Y2=0
cc_532 N_RESET_B_c_811_n N_VGND_c_1056_n 0.00383152f $X=5.57 $Y=1.22 $X2=0 $Y2=0
cc_533 N_RESET_B_c_811_n N_VGND_c_1063_n 0.0075725f $X=5.57 $Y=1.22 $X2=0 $Y2=0
cc_534 N_A_1342_74#_c_844_n N_VPWR_c_905_n 0.0109024f $X=7.655 $Y=1.765 $X2=0
+ $Y2=0
cc_535 N_A_1342_74#_c_850_n N_VPWR_c_905_n 0.0573751f $X=6.925 $Y=2.265 $X2=0
+ $Y2=0
cc_536 N_A_1342_74#_c_846_n N_VPWR_c_905_n 0.0132717f $X=7.55 $Y=1.485 $X2=0
+ $Y2=0
cc_537 N_A_1342_74#_c_850_n N_VPWR_c_909_n 0.00749631f $X=6.925 $Y=2.265 $X2=0
+ $Y2=0
cc_538 N_A_1342_74#_c_844_n N_VPWR_c_910_n 0.00445602f $X=7.655 $Y=1.765 $X2=0
+ $Y2=0
cc_539 N_A_1342_74#_c_844_n N_VPWR_c_901_n 0.00861079f $X=7.655 $Y=1.765 $X2=0
+ $Y2=0
cc_540 N_A_1342_74#_c_850_n N_VPWR_c_901_n 0.0062048f $X=6.925 $Y=2.265 $X2=0
+ $Y2=0
cc_541 N_A_1342_74#_c_845_n N_Q_c_992_n 0.00762129f $X=6.93 $Y=1.32 $X2=0 $Y2=0
cc_542 N_A_1342_74#_c_847_n N_Q_c_992_n 0.033035f $X=6.855 $Y=0.625 $X2=0 $Y2=0
cc_543 N_A_1342_74#_c_845_n N_Q_c_993_n 0.0139769f $X=6.93 $Y=1.32 $X2=0 $Y2=0
cc_544 N_A_1342_74#_c_845_n N_Q_c_994_n 0.0105495f $X=6.93 $Y=1.32 $X2=0 $Y2=0
cc_545 N_A_1342_74#_c_850_n N_Q_c_994_n 0.104675f $X=6.925 $Y=2.265 $X2=0 $Y2=0
cc_546 N_A_1342_74#_c_848_n N_Q_c_994_n 0.0266283f $X=6.93 $Y=1.485 $X2=0 $Y2=0
cc_547 N_A_1342_74#_c_844_n N_Q_N_c_1033_n 0.0120819f $X=7.655 $Y=1.765 $X2=0
+ $Y2=0
cc_548 N_A_1342_74#_c_844_n N_Q_N_c_1034_n 0.00509602f $X=7.655 $Y=1.765 $X2=0
+ $Y2=0
cc_549 N_A_1342_74#_M1020_g N_Q_N_c_1030_n 0.00736672f $X=7.58 $Y=0.74 $X2=0
+ $Y2=0
cc_550 N_A_1342_74#_c_844_n N_Q_N_c_1030_n 0.0121388f $X=7.655 $Y=1.765 $X2=0
+ $Y2=0
cc_551 N_A_1342_74#_c_846_n N_Q_N_c_1030_n 0.0262114f $X=7.55 $Y=1.485 $X2=0
+ $Y2=0
cc_552 N_A_1342_74#_M1020_g Q_N 0.0132824f $X=7.58 $Y=0.74 $X2=0 $Y2=0
cc_553 N_A_1342_74#_c_844_n Q_N 0.00140046f $X=7.655 $Y=1.765 $X2=0 $Y2=0
cc_554 N_A_1342_74#_M1020_g N_VGND_c_1055_n 0.0136941f $X=7.58 $Y=0.74 $X2=0
+ $Y2=0
cc_555 N_A_1342_74#_c_844_n N_VGND_c_1055_n 0.00221326f $X=7.655 $Y=1.765 $X2=0
+ $Y2=0
cc_556 N_A_1342_74#_c_846_n N_VGND_c_1055_n 0.0139393f $X=7.55 $Y=1.485 $X2=0
+ $Y2=0
cc_557 N_A_1342_74#_c_847_n N_VGND_c_1055_n 0.0223138f $X=6.855 $Y=0.625 $X2=0
+ $Y2=0
cc_558 N_A_1342_74#_c_847_n N_VGND_c_1061_n 0.0144085f $X=6.855 $Y=0.625 $X2=0
+ $Y2=0
cc_559 N_A_1342_74#_M1020_g N_VGND_c_1062_n 0.00383152f $X=7.58 $Y=0.74 $X2=0
+ $Y2=0
cc_560 N_A_1342_74#_M1020_g N_VGND_c_1063_n 0.00761455f $X=7.58 $Y=0.74 $X2=0
+ $Y2=0
cc_561 N_A_1342_74#_c_847_n N_VGND_c_1063_n 0.0119386f $X=6.855 $Y=0.625 $X2=0
+ $Y2=0
cc_562 N_VPWR_c_904_n N_Q_c_995_n 0.0371576f $X=5.865 $Y=2.225 $X2=0 $Y2=0
cc_563 N_VPWR_c_909_n Q 0.0208407f $X=7.21 $Y=3.33 $X2=0 $Y2=0
cc_564 N_VPWR_c_901_n Q 0.0172173f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_565 N_VPWR_c_905_n N_Q_N_c_1033_n 0.0331828f $X=7.375 $Y=2.265 $X2=0 $Y2=0
cc_566 N_VPWR_c_910_n N_Q_N_c_1033_n 0.01504f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_567 N_VPWR_c_901_n N_Q_N_c_1033_n 0.0124159f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_568 N_Q_c_992_n N_VGND_c_1054_n 0.0244145f $X=6.295 $Y=0.515 $X2=0 $Y2=0
cc_569 N_Q_c_992_n N_VGND_c_1061_n 0.0145323f $X=6.295 $Y=0.515 $X2=0 $Y2=0
cc_570 N_Q_c_992_n N_VGND_c_1063_n 0.0119861f $X=6.295 $Y=0.515 $X2=0 $Y2=0
cc_571 Q_N N_VGND_c_1055_n 0.0219107f $X=7.835 $Y=0.47 $X2=0 $Y2=0
cc_572 Q_N N_VGND_c_1062_n 0.0153133f $X=7.835 $Y=0.47 $X2=0 $Y2=0
cc_573 Q_N N_VGND_c_1063_n 0.0126713f $X=7.835 $Y=0.47 $X2=0 $Y2=0
