# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ls__nand2_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_ls__nand2_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.160000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  1.560000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.185000 1.220000 7.555000 1.550000 ;
        RECT 5.965000 1.550000 7.555000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.560000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.350000 4.195000 1.780000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  2.284800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.140000 1.950000 4.710000 2.120000 ;
        RECT 2.140000 2.120000 2.470000 2.980000 ;
        RECT 4.335000 0.770000 7.895000 1.050000 ;
        RECT 4.335000 1.050000 4.710000 1.130000 ;
        RECT 4.380000 1.130000 4.710000 1.950000 ;
        RECT 4.380000 2.120000 4.710000 2.980000 ;
        RECT 5.940000 1.950000 7.895000 2.120000 ;
        RECT 5.940000 2.120000 6.270000 2.980000 ;
        RECT 7.320000 2.120000 7.550000 2.980000 ;
        RECT 7.725000 1.050000 7.895000 1.950000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.160000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.160000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.160000 0.085000 ;
      RECT 0.000000  3.245000 8.160000 3.415000 ;
      RECT 0.105000  0.350000 0.355000 1.165000 ;
      RECT 0.105000  1.165000 4.155000 1.180000 ;
      RECT 0.105000  1.180000 1.860000 1.355000 ;
      RECT 0.535000  0.085000 0.865000 0.995000 ;
      RECT 0.660000  1.950000 1.970000 3.245000 ;
      RECT 1.035000  0.350000 1.225000 1.010000 ;
      RECT 1.035000  1.010000 4.155000 1.165000 ;
      RECT 1.395000  0.085000 1.725000 0.840000 ;
      RECT 1.895000  0.350000 2.155000 1.010000 ;
      RECT 2.325000  0.085000 2.905000 0.840000 ;
      RECT 2.640000  2.290000 4.210000 3.245000 ;
      RECT 3.075000  0.350000 3.305000 1.010000 ;
      RECT 3.475000  0.085000 3.805000 0.840000 ;
      RECT 3.985000  0.350000 8.045000 0.600000 ;
      RECT 3.985000  0.600000 4.155000 1.010000 ;
      RECT 4.880000  1.820000 5.210000 3.245000 ;
      RECT 5.440000  1.820000 5.770000 3.245000 ;
      RECT 6.440000  2.290000 7.150000 3.245000 ;
      RECT 7.720000  2.290000 8.050000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
  END
END sky130_fd_sc_ls__nand2_8
END LIBRARY
