* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__clkdlyinv5sd2_1 A VGND VNB VPB VPWR Y
M1000 a_549_74# a_288_74# VGND VNB nshort w=420000u l=180000u
+  ad=1.113e+11p pd=1.37e+06u as=7.371e+11p ps=6.03e+06u
M1001 a_549_74# a_288_74# VPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.65e+11p pd=2.53e+06u as=1.6848e+12p ps=9.72e+06u
M1002 Y a_682_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1003 VGND a_549_74# a_682_74# VNB nshort w=420000u l=180000u
+  ad=0p pd=0u as=2.457e+11p ps=2.01e+06u
M1004 VPWR a_549_74# a_682_74# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=5.1e+11p ps=3.02e+06u
M1005 Y a_682_74# VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1006 a_288_74# a_28_74# VGND VNB nshort w=420000u l=180000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1007 VGND A a_28_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1008 VPWR A a_28_74# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1009 a_288_74# a_28_74# VPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.6e+11p pd=2.52e+06u as=0p ps=0u
.ends
