* NGSPICE file created from sky130_fd_sc_ls__dlxbn_1.ext - technology: sky130A

.subckt sky130_fd_sc_ls__dlxbn_1 D GATE_N VGND VNB VPB VPWR Q Q_N
M1000 a_805_392# a_232_82# a_653_79# VPB phighvt w=420000u l=150000u
+  ad=1.407e+11p pd=1.51e+06u as=4.057e+11p ps=3.2e+06u
M1001 a_232_82# GATE_N VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=1.4754e+12p ps=1.217e+07u
M1002 a_863_294# a_653_79# VGND VNB nshort w=740000u l=150000u
+  ad=2.183e+11p pd=2.07e+06u as=0p ps=0u
M1003 a_571_392# a_27_120# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.7e+11p pd=2.54e+06u as=1.8056e+12p ps=1.431e+07u
M1004 VGND a_863_294# a_852_123# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1005 Q_N a_1347_424# VGND VNB nshort w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1006 VPWR D a_27_120# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=2.94e+11p ps=2.38e+06u
M1007 VGND a_232_82# a_343_80# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=3.182e+11p ps=2.34e+06u
M1008 VGND a_863_294# Q VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1009 Q_N a_1347_424# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=0p ps=0u
M1010 a_852_123# a_343_80# a_653_79# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=4.099e+11p ps=2.97e+06u
M1011 a_232_82# GATE_N VPWR VPB phighvt w=840000u l=150000u
+  ad=2.478e+11p pd=2.27e+06u as=0p ps=0u
M1012 a_653_79# a_232_82# a_575_79# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=1.536e+11p ps=1.76e+06u
M1013 a_575_79# a_27_120# VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_863_294# a_653_79# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1015 VPWR a_863_294# a_805_392# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_1347_424# a_863_294# VGND VNB nshort w=550000u l=150000u
+  ad=1.5675e+11p pd=1.67e+06u as=0p ps=0u
M1017 VGND D a_27_120# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1018 VPWR a_232_82# a_343_80# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=2.478e+11p ps=2.27e+06u
M1019 VPWR a_863_294# Q VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1020 a_1347_424# a_863_294# VPWR VPB phighvt w=840000u l=150000u
+  ad=2.478e+11p pd=2.27e+06u as=0p ps=0u
M1021 a_653_79# a_343_80# a_571_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

