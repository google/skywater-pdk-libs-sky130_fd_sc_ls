* File: sky130_fd_sc_ls__sdfrbp_2.pxi.spice
* Created: Wed Sep  2 11:27:01 2020
* 
x_PM_SKY130_FD_SC_LS__SDFRBP_2%A_27_79# N_A_27_79#_M1027_s N_A_27_79#_M1026_s
+ N_A_27_79#_M1007_g N_A_27_79#_c_281_n N_A_27_79#_M1014_g N_A_27_79#_c_276_n
+ N_A_27_79#_c_277_n N_A_27_79#_c_278_n N_A_27_79#_c_283_n N_A_27_79#_c_279_n
+ N_A_27_79#_c_295_p N_A_27_79#_c_284_n N_A_27_79#_c_280_n N_A_27_79#_c_285_n
+ PM_SKY130_FD_SC_LS__SDFRBP_2%A_27_79#
x_PM_SKY130_FD_SC_LS__SDFRBP_2%SCE N_SCE_c_358_n N_SCE_c_359_n N_SCE_M1027_g
+ N_SCE_c_367_n N_SCE_M1026_g N_SCE_c_368_n N_SCE_M1030_g N_SCE_M1028_g
+ N_SCE_c_361_n N_SCE_c_362_n N_SCE_c_363_n N_SCE_c_364_n N_SCE_c_365_n SCE SCE
+ SCE N_SCE_c_370_n N_SCE_c_371_n PM_SKY130_FD_SC_LS__SDFRBP_2%SCE
x_PM_SKY130_FD_SC_LS__SDFRBP_2%D N_D_M1023_g N_D_c_444_n N_D_c_449_n N_D_M1018_g
+ D N_D_c_445_n N_D_c_446_n N_D_c_447_n PM_SKY130_FD_SC_LS__SDFRBP_2%D
x_PM_SKY130_FD_SC_LS__SDFRBP_2%SCD N_SCD_c_495_n N_SCD_M1031_g N_SCD_M1008_g
+ N_SCD_c_492_n SCD SCD N_SCD_c_494_n PM_SKY130_FD_SC_LS__SDFRBP_2%SCD
x_PM_SKY130_FD_SC_LS__SDFRBP_2%CLK N_CLK_c_535_n N_CLK_M1019_g N_CLK_M1032_g CLK
+ PM_SKY130_FD_SC_LS__SDFRBP_2%CLK
x_PM_SKY130_FD_SC_LS__SDFRBP_2%A_1025_119# N_A_1025_119#_M1029_d
+ N_A_1025_119#_M1035_d N_A_1025_119#_c_596_n N_A_1025_119#_c_597_n
+ N_A_1025_119#_M1033_g N_A_1025_119#_c_576_n N_A_1025_119#_M1011_g
+ N_A_1025_119#_c_578_n N_A_1025_119#_M1016_g N_A_1025_119#_c_579_n
+ N_A_1025_119#_c_580_n N_A_1025_119#_c_598_n N_A_1025_119#_M1024_g
+ N_A_1025_119#_c_581_n N_A_1025_119#_c_582_n N_A_1025_119#_c_583_n
+ N_A_1025_119#_c_584_n N_A_1025_119#_c_585_n N_A_1025_119#_c_746_p
+ N_A_1025_119#_c_586_n N_A_1025_119#_c_587_n N_A_1025_119#_c_588_n
+ N_A_1025_119#_c_589_n N_A_1025_119#_c_590_n N_A_1025_119#_c_591_n
+ N_A_1025_119#_c_592_n N_A_1025_119#_c_593_n N_A_1025_119#_c_600_n
+ N_A_1025_119#_c_594_n N_A_1025_119#_c_595_n
+ PM_SKY130_FD_SC_LS__SDFRBP_2%A_1025_119#
x_PM_SKY130_FD_SC_LS__SDFRBP_2%A_1370_290# N_A_1370_290#_M1002_d
+ N_A_1370_290#_M1039_d N_A_1370_290#_c_776_n N_A_1370_290#_M1040_g
+ N_A_1370_290#_c_777_n N_A_1370_290#_M1042_g N_A_1370_290#_c_771_n
+ N_A_1370_290#_c_772_n N_A_1370_290#_c_791_n N_A_1370_290#_c_793_n
+ N_A_1370_290#_c_780_n N_A_1370_290#_c_773_n N_A_1370_290#_c_774_n
+ N_A_1370_290#_c_775_n PM_SKY130_FD_SC_LS__SDFRBP_2%A_1370_290#
x_PM_SKY130_FD_SC_LS__SDFRBP_2%RESET_B N_RESET_B_M1000_g N_RESET_B_c_875_n
+ N_RESET_B_M1044_g N_RESET_B_c_866_n N_RESET_B_c_867_n N_RESET_B_M1006_g
+ N_RESET_B_c_869_n N_RESET_B_c_870_n N_RESET_B_c_876_n N_RESET_B_M1015_g
+ N_RESET_B_c_871_n N_RESET_B_M1020_g N_RESET_B_c_878_n N_RESET_B_c_879_n
+ N_RESET_B_M1009_g N_RESET_B_c_873_n N_RESET_B_c_881_n N_RESET_B_c_882_n
+ N_RESET_B_c_883_n N_RESET_B_c_884_n RESET_B N_RESET_B_c_886_n
+ N_RESET_B_c_887_n N_RESET_B_c_888_n N_RESET_B_c_889_n N_RESET_B_c_890_n
+ PM_SKY130_FD_SC_LS__SDFRBP_2%RESET_B
x_PM_SKY130_FD_SC_LS__SDFRBP_2%A_1223_119# N_A_1223_119#_M1010_d
+ N_A_1223_119#_M1033_d N_A_1223_119#_M1015_d N_A_1223_119#_M1002_g
+ N_A_1223_119#_c_1069_n N_A_1223_119#_M1039_g N_A_1223_119#_c_1082_n
+ N_A_1223_119#_c_1075_n N_A_1223_119#_c_1095_n N_A_1223_119#_c_1070_n
+ N_A_1223_119#_c_1071_n N_A_1223_119#_c_1072_n N_A_1223_119#_c_1078_n
+ N_A_1223_119#_c_1073_n PM_SKY130_FD_SC_LS__SDFRBP_2%A_1223_119#
x_PM_SKY130_FD_SC_LS__SDFRBP_2%A_852_119# N_A_852_119#_M1019_s
+ N_A_852_119#_M1032_s N_A_852_119#_c_1176_n N_A_852_119#_M1029_g
+ N_A_852_119#_M1035_g N_A_852_119#_c_1177_n N_A_852_119#_c_1189_n
+ N_A_852_119#_c_1178_n N_A_852_119#_c_1179_n N_A_852_119#_c_1190_n
+ N_A_852_119#_c_1191_n N_A_852_119#_c_1180_n N_A_852_119#_M1010_g
+ N_A_852_119#_c_1192_n N_A_852_119#_c_1193_n N_A_852_119#_c_1194_n
+ N_A_852_119#_M1022_g N_A_852_119#_c_1195_n N_A_852_119#_c_1196_n
+ N_A_852_119#_c_1197_n N_A_852_119#_M1004_g N_A_852_119#_c_1181_n
+ N_A_852_119#_c_1182_n N_A_852_119#_M1045_g N_A_852_119#_c_1201_n
+ N_A_852_119#_c_1184_n N_A_852_119#_c_1185_n N_A_852_119#_c_1186_n
+ N_A_852_119#_c_1187_n PM_SKY130_FD_SC_LS__SDFRBP_2%A_852_119#
x_PM_SKY130_FD_SC_LS__SDFRBP_2%A_2006_373# N_A_2006_373#_M1013_d
+ N_A_2006_373#_M1009_d N_A_2006_373#_c_1353_n N_A_2006_373#_M1001_g
+ N_A_2006_373#_M1041_g N_A_2006_373#_c_1355_n N_A_2006_373#_c_1347_n
+ N_A_2006_373#_c_1348_n N_A_2006_373#_c_1357_n N_A_2006_373#_c_1358_n
+ N_A_2006_373#_c_1349_n N_A_2006_373#_c_1350_n N_A_2006_373#_c_1351_n
+ N_A_2006_373#_c_1352_n N_A_2006_373#_c_1359_n N_A_2006_373#_c_1360_n
+ PM_SKY130_FD_SC_LS__SDFRBP_2%A_2006_373#
x_PM_SKY130_FD_SC_LS__SDFRBP_2%A_1790_75# N_A_1790_75#_M1016_d
+ N_A_1790_75#_M1004_d N_A_1790_75#_M1013_g N_A_1790_75#_c_1457_n
+ N_A_1790_75#_c_1467_n N_A_1790_75#_c_1468_n N_A_1790_75#_M1025_g
+ N_A_1790_75#_c_1458_n N_A_1790_75#_c_1469_n N_A_1790_75#_M1003_g
+ N_A_1790_75#_M1021_g N_A_1790_75#_c_1470_n N_A_1790_75#_M1036_g
+ N_A_1790_75#_M1037_g N_A_1790_75#_c_1461_n N_A_1790_75#_c_1462_n
+ N_A_1790_75#_c_1473_n N_A_1790_75#_M1012_g N_A_1790_75#_M1005_g
+ N_A_1790_75#_c_1478_n N_A_1790_75#_c_1480_n N_A_1790_75#_c_1464_n
+ N_A_1790_75#_c_1465_n N_A_1790_75#_c_1466_n N_A_1790_75#_c_1490_n
+ PM_SKY130_FD_SC_LS__SDFRBP_2%A_1790_75#
x_PM_SKY130_FD_SC_LS__SDFRBP_2%A_2604_392# N_A_2604_392#_M1005_d
+ N_A_2604_392#_M1012_d N_A_2604_392#_c_1614_n N_A_2604_392#_M1034_g
+ N_A_2604_392#_M1017_g N_A_2604_392#_c_1615_n N_A_2604_392#_M1043_g
+ N_A_2604_392#_M1038_g N_A_2604_392#_c_1609_n N_A_2604_392#_c_1610_n
+ N_A_2604_392#_c_1611_n N_A_2604_392#_c_1612_n N_A_2604_392#_c_1631_p
+ N_A_2604_392#_c_1613_n PM_SKY130_FD_SC_LS__SDFRBP_2%A_2604_392#
x_PM_SKY130_FD_SC_LS__SDFRBP_2%VPWR N_VPWR_M1026_d N_VPWR_M1031_d N_VPWR_M1032_d
+ N_VPWR_M1042_d N_VPWR_M1039_s N_VPWR_M1001_d N_VPWR_M1025_d N_VPWR_M1036_d
+ N_VPWR_M1034_s N_VPWR_M1043_s N_VPWR_c_1659_n N_VPWR_c_1660_n N_VPWR_c_1661_n
+ N_VPWR_c_1662_n N_VPWR_c_1663_n N_VPWR_c_1664_n N_VPWR_c_1665_n
+ N_VPWR_c_1666_n N_VPWR_c_1667_n N_VPWR_c_1668_n N_VPWR_c_1669_n
+ N_VPWR_c_1670_n N_VPWR_c_1671_n N_VPWR_c_1672_n VPWR N_VPWR_c_1673_n
+ N_VPWR_c_1674_n N_VPWR_c_1675_n N_VPWR_c_1676_n N_VPWR_c_1677_n
+ N_VPWR_c_1678_n N_VPWR_c_1679_n N_VPWR_c_1680_n N_VPWR_c_1681_n
+ N_VPWR_c_1682_n N_VPWR_c_1683_n N_VPWR_c_1684_n N_VPWR_c_1685_n
+ N_VPWR_c_1686_n N_VPWR_c_1658_n PM_SKY130_FD_SC_LS__SDFRBP_2%VPWR
x_PM_SKY130_FD_SC_LS__SDFRBP_2%A_388_79# N_A_388_79#_M1023_d N_A_388_79#_M1010_s
+ N_A_388_79#_M1018_d N_A_388_79#_M1044_d N_A_388_79#_M1033_s
+ N_A_388_79#_c_1865_n N_A_388_79#_c_1847_n N_A_388_79#_c_1848_n
+ N_A_388_79#_c_1849_n N_A_388_79#_c_1867_n N_A_388_79#_c_1888_n
+ N_A_388_79#_c_1856_n N_A_388_79#_c_1850_n N_A_388_79#_c_1858_n
+ N_A_388_79#_c_1859_n N_A_388_79#_c_1851_n N_A_388_79#_c_1860_n
+ N_A_388_79#_c_1852_n N_A_388_79#_c_1853_n N_A_388_79#_c_1854_n
+ N_A_388_79#_c_1862_n N_A_388_79#_c_1902_n N_A_388_79#_c_1855_n
+ N_A_388_79#_c_1863_n PM_SKY130_FD_SC_LS__SDFRBP_2%A_388_79#
x_PM_SKY130_FD_SC_LS__SDFRBP_2%Q_N N_Q_N_M1021_d N_Q_N_M1003_s Q_N Q_N Q_N
+ N_Q_N_c_2009_n Q_N PM_SKY130_FD_SC_LS__SDFRBP_2%Q_N
x_PM_SKY130_FD_SC_LS__SDFRBP_2%Q N_Q_M1017_d N_Q_M1034_d Q N_Q_c_2036_n
+ PM_SKY130_FD_SC_LS__SDFRBP_2%Q
x_PM_SKY130_FD_SC_LS__SDFRBP_2%VGND N_VGND_M1027_d N_VGND_M1000_d N_VGND_M1019_d
+ N_VGND_M1006_d N_VGND_M1041_d N_VGND_M1021_s N_VGND_M1037_s N_VGND_M1017_s
+ N_VGND_M1038_s N_VGND_c_2052_n N_VGND_c_2053_n N_VGND_c_2054_n N_VGND_c_2055_n
+ N_VGND_c_2056_n N_VGND_c_2057_n N_VGND_c_2058_n N_VGND_c_2059_n
+ N_VGND_c_2060_n N_VGND_c_2061_n N_VGND_c_2062_n N_VGND_c_2063_n
+ N_VGND_c_2064_n N_VGND_c_2065_n N_VGND_c_2066_n N_VGND_c_2067_n VGND
+ N_VGND_c_2068_n N_VGND_c_2069_n N_VGND_c_2070_n N_VGND_c_2071_n
+ N_VGND_c_2072_n N_VGND_c_2073_n N_VGND_c_2074_n N_VGND_c_2075_n
+ N_VGND_c_2076_n N_VGND_c_2077_n N_VGND_c_2078_n
+ PM_SKY130_FD_SC_LS__SDFRBP_2%VGND
x_PM_SKY130_FD_SC_LS__SDFRBP_2%noxref_25 N_noxref_25_M1007_s N_noxref_25_M1008_d
+ N_noxref_25_c_2207_n N_noxref_25_c_2208_n N_noxref_25_c_2209_n
+ N_noxref_25_c_2210_n PM_SKY130_FD_SC_LS__SDFRBP_2%noxref_25
cc_1 VNB N_A_27_79#_M1007_g 0.0455097f $X=-0.19 $Y=-0.245 $X2=1.475 $Y2=0.605
cc_2 VNB N_A_27_79#_c_276_n 0.0789787f $X=-0.19 $Y=-0.245 $X2=1.4 $Y2=1.415
cc_3 VNB N_A_27_79#_c_277_n 0.0355558f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=0.605
cc_4 VNB N_A_27_79#_c_278_n 0.00354448f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=2.32
cc_5 VNB N_A_27_79#_c_279_n 0.00484068f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=1.415
cc_6 VNB N_A_27_79#_c_280_n 0.0159647f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.415
cc_7 VNB N_SCE_c_358_n 0.0443833f $X=-0.19 $Y=-0.245 $X2=0.135 $Y2=2.32
cc_8 VNB N_SCE_c_359_n 0.0211781f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_SCE_M1028_g 0.0363026f $X=-0.19 $Y=-0.245 $X2=1.4 $Y2=1.415
cc_10 VNB N_SCE_c_361_n 0.0216296f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_SCE_c_362_n 0.00133979f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.65
cc_12 VNB N_SCE_c_363_n 0.00450757f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_SCE_c_364_n 0.0230028f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=1.415
cc_14 VNB N_SCE_c_365_n 0.0330707f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=1.415
cc_15 VNB N_D_c_444_n 0.0238331f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_D_c_445_n 0.0310845f $X=-0.19 $Y=-0.245 $X2=2.615 $Y2=2.64
cc_17 VNB N_D_c_446_n 0.00902418f $X=-0.19 $Y=-0.245 $X2=2.615 $Y2=2.64
cc_18 VNB N_D_c_447_n 0.0162587f $X=-0.19 $Y=-0.245 $X2=1.4 $Y2=1.415
cc_19 VNB N_SCD_M1008_g 0.042619f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_SCD_c_492_n 0.00499797f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB SCD 0.00197778f $X=-0.19 $Y=-0.245 $X2=2.615 $Y2=2.245
cc_22 VNB N_SCD_c_494_n 0.0164016f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.605
cc_23 VNB N_CLK_c_535_n 0.103954f $X=-0.19 $Y=-0.245 $X2=0.135 $Y2=0.395
cc_24 VNB CLK 0.0128351f $X=-0.19 $Y=-0.245 $X2=1.475 $Y2=0.605
cc_25 VNB N_A_1025_119#_c_576_n 0.0269582f $X=-0.19 $Y=-0.245 $X2=2.615 $Y2=2.64
cc_26 VNB N_A_1025_119#_M1011_g 0.0361986f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.605
cc_27 VNB N_A_1025_119#_c_578_n 0.0167906f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_1025_119#_c_579_n 0.0173598f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.49
cc_29 VNB N_A_1025_119#_c_580_n 0.00726011f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.65
cc_30 VNB N_A_1025_119#_c_581_n 0.0063026f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_1025_119#_c_582_n 0.0213285f $X=-0.19 $Y=-0.245 $X2=2.275
+ $Y2=2.405
cc_32 VNB N_A_1025_119#_c_583_n 0.00390562f $X=-0.19 $Y=-0.245 $X2=0.445
+ $Y2=2.405
cc_33 VNB N_A_1025_119#_c_584_n 0.00193797f $X=-0.19 $Y=-0.245 $X2=2.44
+ $Y2=1.995
cc_34 VNB N_A_1025_119#_c_585_n 0.00174335f $X=-0.19 $Y=-0.245 $X2=2.44
+ $Y2=1.995
cc_35 VNB N_A_1025_119#_c_586_n 0.00716745f $X=-0.19 $Y=-0.245 $X2=0.28
+ $Y2=2.405
cc_36 VNB N_A_1025_119#_c_587_n 0.00251082f $X=-0.19 $Y=-0.245 $X2=1.23
+ $Y2=1.415
cc_37 VNB N_A_1025_119#_c_588_n 0.00159202f $X=-0.19 $Y=-0.245 $X2=2.49
+ $Y2=1.995
cc_38 VNB N_A_1025_119#_c_589_n 0.00445673f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_1025_119#_c_590_n 0.00416989f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_1025_119#_c_591_n 0.00358753f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_1025_119#_c_592_n 0.00459644f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_1025_119#_c_593_n 0.0333667f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_1025_119#_c_594_n 0.00474639f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_1025_119#_c_595_n 0.0130177f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_1370_290#_M1040_g 0.0295995f $X=-0.19 $Y=-0.245 $X2=2.615
+ $Y2=2.245
cc_46 VNB N_A_1370_290#_c_771_n 0.00357226f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_1370_290#_c_772_n 0.0255382f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=1.58
cc_48 VNB N_A_1370_290#_c_773_n 0.00909034f $X=-0.19 $Y=-0.245 $X2=2.44
+ $Y2=1.995
cc_49 VNB N_A_1370_290#_c_774_n 0.00431592f $X=-0.19 $Y=-0.245 $X2=2.44
+ $Y2=1.995
cc_50 VNB N_A_1370_290#_c_775_n 0.00658141f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_RESET_B_M1000_g 0.0567158f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_RESET_B_c_866_n 0.271622f $X=-0.19 $Y=-0.245 $X2=1.475 $Y2=0.605
cc_53 VNB N_RESET_B_c_867_n 0.0126359f $X=-0.19 $Y=-0.245 $X2=1.475 $Y2=0.605
cc_54 VNB N_RESET_B_M1006_g 0.0292065f $X=-0.19 $Y=-0.245 $X2=2.615 $Y2=2.64
cc_55 VNB N_RESET_B_c_869_n 0.0258223f $X=-0.19 $Y=-0.245 $X2=1.4 $Y2=1.415
cc_56 VNB N_RESET_B_c_870_n 0.0119677f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.25
cc_57 VNB N_RESET_B_c_871_n 0.0223419f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=2.32
cc_58 VNB N_RESET_B_M1020_g 0.0456332f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.65
cc_59 VNB N_RESET_B_c_873_n 0.0112292f $X=-0.19 $Y=-0.245 $X2=2.44 $Y2=2.32
cc_60 VNB N_A_1223_119#_M1002_g 0.0268009f $X=-0.19 $Y=-0.245 $X2=2.615 $Y2=2.64
cc_61 VNB N_A_1223_119#_c_1069_n 0.0288104f $X=-0.19 $Y=-0.245 $X2=1.4 $Y2=1.415
cc_62 VNB N_A_1223_119#_c_1070_n 0.00155425f $X=-0.19 $Y=-0.245 $X2=2.275
+ $Y2=2.405
cc_63 VNB N_A_1223_119#_c_1071_n 0.00408417f $X=-0.19 $Y=-0.245 $X2=0.445
+ $Y2=2.405
cc_64 VNB N_A_1223_119#_c_1072_n 0.00984593f $X=-0.19 $Y=-0.245 $X2=2.44
+ $Y2=1.995
cc_65 VNB N_A_1223_119#_c_1073_n 0.0108902f $X=-0.19 $Y=-0.245 $X2=0.24
+ $Y2=1.415
cc_66 VNB N_A_852_119#_c_1176_n 0.0166255f $X=-0.19 $Y=-0.245 $X2=1.475 $Y2=1.25
cc_67 VNB N_A_852_119#_c_1177_n 0.0108198f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.25
cc_68 VNB N_A_852_119#_c_1178_n 0.025462f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_852_119#_c_1179_n 0.0105739f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=1.58
cc_70 VNB N_A_852_119#_c_1180_n 0.0149335f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.65
cc_71 VNB N_A_852_119#_c_1181_n 0.0298264f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.405
cc_72 VNB N_A_852_119#_c_1182_n 0.00535099f $X=-0.19 $Y=-0.245 $X2=1.23
+ $Y2=1.415
cc_73 VNB N_A_852_119#_M1045_g 0.045335f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_852_119#_c_1184_n 6.70936e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_852_119#_c_1185_n 0.00599319f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_852_119#_c_1186_n 0.00828774f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_852_119#_c_1187_n 0.0430016f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_2006_373#_M1041_g 0.0481405f $X=-0.19 $Y=-0.245 $X2=2.615 $Y2=2.64
cc_79 VNB N_A_2006_373#_c_1347_n 0.00410394f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=1.58
cc_80 VNB N_A_2006_373#_c_1348_n 0.00173724f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=2.32
cc_81 VNB N_A_2006_373#_c_1349_n 0.0070639f $X=-0.19 $Y=-0.245 $X2=0.365
+ $Y2=1.415
cc_82 VNB N_A_2006_373#_c_1350_n 0.00667447f $X=-0.19 $Y=-0.245 $X2=1.23
+ $Y2=1.415
cc_83 VNB N_A_2006_373#_c_1351_n 0.00230863f $X=-0.19 $Y=-0.245 $X2=1.23
+ $Y2=1.415
cc_84 VNB N_A_2006_373#_c_1352_n 0.00172407f $X=-0.19 $Y=-0.245 $X2=2.275
+ $Y2=2.405
cc_85 VNB N_A_1790_75#_M1013_g 0.0262898f $X=-0.19 $Y=-0.245 $X2=1.475 $Y2=0.605
cc_86 VNB N_A_1790_75#_c_1457_n 0.0559917f $X=-0.19 $Y=-0.245 $X2=2.615
+ $Y2=2.245
cc_87 VNB N_A_1790_75#_c_1458_n 0.0318785f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.605
cc_88 VNB N_A_1790_75#_M1021_g 0.0197591f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.65
cc_89 VNB N_A_1790_75#_M1037_g 0.0192815f $X=-0.19 $Y=-0.245 $X2=2.275 $Y2=2.405
cc_90 VNB N_A_1790_75#_c_1461_n 0.0729414f $X=-0.19 $Y=-0.245 $X2=2.44 $Y2=2.32
cc_91 VNB N_A_1790_75#_c_1462_n 0.00428291f $X=-0.19 $Y=-0.245 $X2=2.44
+ $Y2=1.995
cc_92 VNB N_A_1790_75#_M1005_g 0.027051f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=1.415
cc_93 VNB N_A_1790_75#_c_1464_n 0.00230536f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_1790_75#_c_1465_n 0.00223918f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_1790_75#_c_1466_n 0.021329f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_2604_392#_M1017_g 0.023917f $X=-0.19 $Y=-0.245 $X2=2.615 $Y2=2.64
cc_97 VNB N_A_2604_392#_M1038_g 0.0268211f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=1.58
cc_98 VNB N_A_2604_392#_c_1609_n 0.0652038f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.49
cc_99 VNB N_A_2604_392#_c_1610_n 0.0587782f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_A_2604_392#_c_1611_n 0.0102396f $X=-0.19 $Y=-0.245 $X2=1.23
+ $Y2=1.415
cc_101 VNB N_A_2604_392#_c_1612_n 7.2775e-19 $X=-0.19 $Y=-0.245 $X2=2.44
+ $Y2=2.32
cc_102 VNB N_A_2604_392#_c_1613_n 0.00109231f $X=-0.19 $Y=-0.245 $X2=2.49
+ $Y2=1.995
cc_103 VNB N_VPWR_c_1658_n 0.621437f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_A_388_79#_c_1847_n 0.00214649f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.65
cc_105 VNB N_A_388_79#_c_1848_n 0.0235335f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_A_388_79#_c_1849_n 0.00417762f $X=-0.19 $Y=-0.245 $X2=0.365
+ $Y2=1.415
cc_107 VNB N_A_388_79#_c_1850_n 0.0041886f $X=-0.19 $Y=-0.245 $X2=0.445
+ $Y2=2.405
cc_108 VNB N_A_388_79#_c_1851_n 5.87737e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_A_388_79#_c_1852_n 0.00626889f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_A_388_79#_c_1853_n 0.00170831f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_A_388_79#_c_1854_n 0.00300845f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_A_388_79#_c_1855_n 0.00181996f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB Q_N 0.00143966f $X=-0.19 $Y=-0.245 $X2=1.475 $Y2=0.605
cc_114 VNB N_Q_N_c_2009_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.605
cc_115 VNB N_Q_c_2036_n 0.0065793f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_VGND_c_2052_n 0.0153683f $X=-0.19 $Y=-0.245 $X2=2.275 $Y2=2.405
cc_117 VNB N_VGND_c_2053_n 0.0225435f $X=-0.19 $Y=-0.245 $X2=2.44 $Y2=1.995
cc_118 VNB N_VGND_c_2054_n 0.0139405f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.405
cc_119 VNB N_VGND_c_2055_n 0.00692506f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_VGND_c_2056_n 0.00869988f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_VGND_c_2057_n 0.0114612f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_VGND_c_2058_n 0.0225701f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB N_VGND_c_2059_n 0.00935384f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_VGND_c_2060_n 0.0108727f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_2061_n 0.0526431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_2062_n 0.0649427f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_VGND_c_2063_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_2064_n 0.0210525f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_2065_n 0.00226387f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_2066_n 0.0583825f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_2067_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_VGND_c_2068_n 0.0176416f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_VGND_c_2069_n 0.0276584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_VGND_c_2070_n 0.0209223f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_VGND_c_2071_n 0.0186734f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_VGND_c_2072_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_VGND_c_2073_n 0.0605454f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB N_VGND_c_2074_n 0.0190429f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VNB N_VGND_c_2075_n 0.00478044f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_VGND_c_2076_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_141 VNB N_VGND_c_2077_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_142 VNB N_VGND_c_2078_n 0.772554f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_143 VNB N_noxref_25_c_2207_n 0.00622698f $X=-0.19 $Y=-0.245 $X2=1.475
+ $Y2=0.605
cc_144 VNB N_noxref_25_c_2208_n 0.017862f $X=-0.19 $Y=-0.245 $X2=2.615 $Y2=2.245
cc_145 VNB N_noxref_25_c_2209_n 0.00386383f $X=-0.19 $Y=-0.245 $X2=2.615
+ $Y2=2.64
cc_146 VNB N_noxref_25_c_2210_n 0.00276768f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.25
cc_147 VPB N_A_27_79#_c_281_n 0.0656313f $X=-0.19 $Y=1.66 $X2=2.615 $Y2=2.245
cc_148 VPB N_A_27_79#_c_278_n 0.031275f $X=-0.19 $Y=1.66 $X2=0.2 $Y2=2.32
cc_149 VPB N_A_27_79#_c_283_n 0.0213374f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.65
cc_150 VPB N_A_27_79#_c_284_n 0.00449549f $X=-0.19 $Y=1.66 $X2=2.44 $Y2=1.995
cc_151 VPB N_A_27_79#_c_285_n 0.00957909f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.405
cc_152 VPB N_SCE_c_358_n 0.013397f $X=-0.19 $Y=1.66 $X2=0.135 $Y2=2.32
cc_153 VPB N_SCE_c_367_n 0.052364f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_154 VPB N_SCE_c_368_n 0.0413346f $X=-0.19 $Y=1.66 $X2=1.475 $Y2=0.605
cc_155 VPB N_SCE_c_362_n 0.00700226f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.65
cc_156 VPB N_SCE_c_370_n 0.0605067f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_157 VPB N_SCE_c_371_n 0.00222208f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_158 VPB N_D_c_444_n 0.0324711f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_159 VPB N_D_c_449_n 0.0243702f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_160 VPB N_SCD_c_495_n 0.0168486f $X=-0.19 $Y=1.66 $X2=0.135 $Y2=0.395
cc_161 VPB N_SCD_c_492_n 0.0497542f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_162 VPB SCD 0.00164304f $X=-0.19 $Y=1.66 $X2=2.615 $Y2=2.245
cc_163 VPB N_CLK_M1032_g 0.023763f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_164 VPB N_A_1025_119#_c_596_n 0.0178704f $X=-0.19 $Y=1.66 $X2=1.475 $Y2=0.605
cc_165 VPB N_A_1025_119#_c_597_n 0.0194025f $X=-0.19 $Y=1.66 $X2=1.475 $Y2=0.605
cc_166 VPB N_A_1025_119#_c_598_n 0.0554159f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.65
cc_167 VPB N_A_1025_119#_c_590_n 0.00720545f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_168 VPB N_A_1025_119#_c_600_n 0.00662341f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_169 VPB N_A_1025_119#_c_594_n 0.0041865f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_170 VPB N_A_1025_119#_c_595_n 0.0168953f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_171 VPB N_A_1370_290#_c_776_n 0.024486f $X=-0.19 $Y=1.66 $X2=1.475 $Y2=0.605
cc_172 VPB N_A_1370_290#_c_777_n 0.0207961f $X=-0.19 $Y=1.66 $X2=2.615 $Y2=2.64
cc_173 VPB N_A_1370_290#_c_771_n 0.00212444f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_174 VPB N_A_1370_290#_c_772_n 0.0186985f $X=-0.19 $Y=1.66 $X2=0.2 $Y2=1.58
cc_175 VPB N_A_1370_290#_c_780_n 0.0024203f $X=-0.19 $Y=1.66 $X2=0.365 $Y2=1.415
cc_176 VPB N_A_1370_290#_c_775_n 0.00166674f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_177 VPB N_RESET_B_M1000_g 0.00640222f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_178 VPB N_RESET_B_c_875_n 0.0215686f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_179 VPB N_RESET_B_c_876_n 0.0164974f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=0.605
cc_180 VPB N_RESET_B_c_871_n 0.00915309f $X=-0.19 $Y=1.66 $X2=0.2 $Y2=2.32
cc_181 VPB N_RESET_B_c_878_n 0.0120728f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=1.415
cc_182 VPB N_RESET_B_c_879_n 0.0547375f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=1.415
cc_183 VPB N_RESET_B_c_873_n 0.00587573f $X=-0.19 $Y=1.66 $X2=2.44 $Y2=2.32
cc_184 VPB N_RESET_B_c_881_n 0.02191f $X=-0.19 $Y=1.66 $X2=2.44 $Y2=1.995
cc_185 VPB N_RESET_B_c_882_n 0.00347238f $X=-0.19 $Y=1.66 $X2=2.44 $Y2=1.995
cc_186 VPB N_RESET_B_c_883_n 0.00850003f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_187 VPB N_RESET_B_c_884_n 0.00382672f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.415
cc_188 VPB RESET_B 0.00298374f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_189 VPB N_RESET_B_c_886_n 0.0668095f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_190 VPB N_RESET_B_c_887_n 0.00207352f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_191 VPB N_RESET_B_c_888_n 0.0565102f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_192 VPB N_RESET_B_c_889_n 0.00232432f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_193 VPB N_RESET_B_c_890_n 0.0062794f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_194 VPB N_A_1223_119#_c_1069_n 0.0272296f $X=-0.19 $Y=1.66 $X2=1.4 $Y2=1.415
cc_195 VPB N_A_1223_119#_c_1075_n 0.0032604f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.49
cc_196 VPB N_A_1223_119#_c_1070_n 0.01535f $X=-0.19 $Y=1.66 $X2=2.275 $Y2=2.405
cc_197 VPB N_A_1223_119#_c_1072_n 0.00370269f $X=-0.19 $Y=1.66 $X2=2.44
+ $Y2=1.995
cc_198 VPB N_A_1223_119#_c_1078_n 0.0020586f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_199 VPB N_A_1223_119#_c_1073_n 0.0113579f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.415
cc_200 VPB N_A_852_119#_M1035_g 0.0213965f $X=-0.19 $Y=1.66 $X2=2.615 $Y2=2.64
cc_201 VPB N_A_852_119#_c_1189_n 0.0706807f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=0.605
cc_202 VPB N_A_852_119#_c_1190_n 0.0543441f $X=-0.19 $Y=1.66 $X2=0.2 $Y2=2.32
cc_203 VPB N_A_852_119#_c_1191_n 0.0123654f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.49
cc_204 VPB N_A_852_119#_c_1192_n 0.00707596f $X=-0.19 $Y=1.66 $X2=0.365
+ $Y2=1.415
cc_205 VPB N_A_852_119#_c_1193_n 0.0191676f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=1.415
cc_206 VPB N_A_852_119#_c_1194_n 0.013948f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=1.415
cc_207 VPB N_A_852_119#_c_1195_n 0.179501f $X=-0.19 $Y=1.66 $X2=2.275 $Y2=2.405
cc_208 VPB N_A_852_119#_c_1196_n 0.00747951f $X=-0.19 $Y=1.66 $X2=2.44 $Y2=2.32
cc_209 VPB N_A_852_119#_c_1197_n 0.0161081f $X=-0.19 $Y=1.66 $X2=2.44 $Y2=1.995
cc_210 VPB N_A_852_119#_M1004_g 0.00865924f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.415
cc_211 VPB N_A_852_119#_c_1181_n 0.0303876f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.405
cc_212 VPB N_A_852_119#_c_1182_n 0.00515977f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=1.415
cc_213 VPB N_A_852_119#_c_1201_n 0.0089867f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_214 VPB N_A_852_119#_c_1186_n 0.00464413f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_215 VPB N_A_2006_373#_c_1353_n 0.0154015f $X=-0.19 $Y=1.66 $X2=1.475 $Y2=1.25
cc_216 VPB N_A_2006_373#_M1041_g 0.0146783f $X=-0.19 $Y=1.66 $X2=2.615 $Y2=2.64
cc_217 VPB N_A_2006_373#_c_1355_n 0.0043277f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=0.605
cc_218 VPB N_A_2006_373#_c_1347_n 0.010942f $X=-0.19 $Y=1.66 $X2=0.2 $Y2=1.58
cc_219 VPB N_A_2006_373#_c_1357_n 0.00277764f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.49
cc_220 VPB N_A_2006_373#_c_1358_n 2.07695e-19 $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.65
cc_221 VPB N_A_2006_373#_c_1359_n 0.00608544f $X=-0.19 $Y=1.66 $X2=0.445
+ $Y2=2.405
cc_222 VPB N_A_2006_373#_c_1360_n 0.0572791f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.415
cc_223 VPB N_A_1790_75#_c_1467_n 0.0332504f $X=-0.19 $Y=1.66 $X2=2.615 $Y2=2.64
cc_224 VPB N_A_1790_75#_c_1468_n 0.0220882f $X=-0.19 $Y=1.66 $X2=2.615 $Y2=2.64
cc_225 VPB N_A_1790_75#_c_1469_n 0.0159809f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_226 VPB N_A_1790_75#_c_1470_n 0.0160546f $X=-0.19 $Y=1.66 $X2=0.365 $Y2=1.415
cc_227 VPB N_A_1790_75#_c_1461_n 0.0202262f $X=-0.19 $Y=1.66 $X2=2.44 $Y2=2.32
cc_228 VPB N_A_1790_75#_c_1462_n 0.00804325f $X=-0.19 $Y=1.66 $X2=2.44 $Y2=1.995
cc_229 VPB N_A_1790_75#_c_1473_n 0.0246892f $X=-0.19 $Y=1.66 $X2=2.44 $Y2=1.995
cc_230 VPB N_A_1790_75#_c_1465_n 0.00737395f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_231 VPB N_A_2604_392#_c_1614_n 0.0177068f $X=-0.19 $Y=1.66 $X2=1.475 $Y2=1.25
cc_232 VPB N_A_2604_392#_c_1615_n 0.0174134f $X=-0.19 $Y=1.66 $X2=1.4 $Y2=1.415
cc_233 VPB N_A_2604_392#_c_1610_n 0.0176653f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_234 VPB N_A_2604_392#_c_1612_n 0.0195039f $X=-0.19 $Y=1.66 $X2=2.44 $Y2=2.32
cc_235 VPB N_VPWR_c_1659_n 0.00985307f $X=-0.19 $Y=1.66 $X2=2.44 $Y2=1.995
cc_236 VPB N_VPWR_c_1660_n 0.00396467f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.415
cc_237 VPB N_VPWR_c_1661_n 0.0079126f $X=-0.19 $Y=1.66 $X2=2.49 $Y2=1.995
cc_238 VPB N_VPWR_c_1662_n 0.0135327f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_239 VPB N_VPWR_c_1663_n 0.0511217f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_240 VPB N_VPWR_c_1664_n 0.0221602f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_241 VPB N_VPWR_c_1665_n 0.0103382f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_242 VPB N_VPWR_c_1666_n 0.0184711f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_243 VPB N_VPWR_c_1667_n 0.0109102f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_244 VPB N_VPWR_c_1668_n 0.0663373f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_245 VPB N_VPWR_c_1669_n 0.0343579f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_246 VPB N_VPWR_c_1670_n 0.00601569f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_247 VPB N_VPWR_c_1671_n 0.0563142f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_248 VPB N_VPWR_c_1672_n 0.00330333f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_249 VPB N_VPWR_c_1673_n 0.0474691f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_250 VPB N_VPWR_c_1674_n 0.0237904f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_251 VPB N_VPWR_c_1675_n 0.0217361f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_252 VPB N_VPWR_c_1676_n 0.0193312f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_253 VPB N_VPWR_c_1677_n 0.0206736f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_254 VPB N_VPWR_c_1678_n 0.0174144f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_255 VPB N_VPWR_c_1679_n 0.0191515f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_256 VPB N_VPWR_c_1680_n 0.0263586f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_257 VPB N_VPWR_c_1681_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_258 VPB N_VPWR_c_1682_n 0.00330333f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_259 VPB N_VPWR_c_1683_n 0.0389406f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_260 VPB N_VPWR_c_1684_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_261 VPB N_VPWR_c_1685_n 0.00555219f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_262 VPB N_VPWR_c_1686_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_263 VPB N_VPWR_c_1658_n 0.130753f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_264 VPB N_A_388_79#_c_1856_n 0.0051238f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_265 VPB N_A_388_79#_c_1850_n 0.00481007f $X=-0.19 $Y=1.66 $X2=0.445 $Y2=2.405
cc_266 VPB N_A_388_79#_c_1858_n 0.0124567f $X=-0.19 $Y=1.66 $X2=2.44 $Y2=2.32
cc_267 VPB N_A_388_79#_c_1859_n 0.00269448f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.415
cc_268 VPB N_A_388_79#_c_1860_n 5.99802e-19 $X=-0.19 $Y=1.66 $X2=2.49 $Y2=1.995
cc_269 VPB N_A_388_79#_c_1854_n 0.00737551f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_270 VPB N_A_388_79#_c_1862_n 0.00834887f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_271 VPB N_A_388_79#_c_1863_n 0.00668435f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_272 VPB Q_N 0.00344098f $X=-0.19 $Y=1.66 $X2=1.475 $Y2=0.605
cc_273 VPB N_Q_c_2036_n 0.00405531f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_274 N_A_27_79#_c_276_n N_SCE_c_358_n 0.0181735f $X=1.4 $Y=1.415 $X2=0 $Y2=0
cc_275 N_A_27_79#_c_277_n N_SCE_c_358_n 0.0127444f $X=0.28 $Y=0.605 $X2=0 $Y2=0
cc_276 N_A_27_79#_c_278_n N_SCE_c_358_n 0.0140797f $X=0.2 $Y=2.32 $X2=0 $Y2=0
cc_277 N_A_27_79#_c_279_n N_SCE_c_358_n 0.0179605f $X=1.23 $Y=1.415 $X2=0 $Y2=0
cc_278 N_A_27_79#_c_280_n N_SCE_c_358_n 0.00851213f $X=0.24 $Y=1.415 $X2=0 $Y2=0
cc_279 N_A_27_79#_c_277_n N_SCE_c_359_n 0.00367837f $X=0.28 $Y=0.605 $X2=0 $Y2=0
cc_280 N_A_27_79#_c_278_n N_SCE_c_367_n 0.0112444f $X=0.2 $Y=2.32 $X2=0 $Y2=0
cc_281 N_A_27_79#_c_283_n N_SCE_c_367_n 0.0155777f $X=0.28 $Y=2.65 $X2=0 $Y2=0
cc_282 N_A_27_79#_c_279_n N_SCE_c_367_n 0.00644399f $X=1.23 $Y=1.415 $X2=0 $Y2=0
cc_283 N_A_27_79#_c_295_p N_SCE_c_367_n 0.0138322f $X=2.275 $Y=2.405 $X2=0 $Y2=0
cc_284 N_A_27_79#_c_285_n N_SCE_c_367_n 0.00605135f $X=0.28 $Y=2.405 $X2=0 $Y2=0
cc_285 N_A_27_79#_c_295_p N_SCE_c_368_n 0.0137373f $X=2.275 $Y=2.405 $X2=0 $Y2=0
cc_286 N_A_27_79#_c_277_n N_SCE_c_361_n 0.0100023f $X=0.28 $Y=0.605 $X2=0 $Y2=0
cc_287 N_A_27_79#_c_279_n N_SCE_c_361_n 0.00327315f $X=1.23 $Y=1.415 $X2=0 $Y2=0
cc_288 N_A_27_79#_c_281_n N_SCE_c_362_n 0.00102331f $X=2.615 $Y=2.245 $X2=0
+ $Y2=0
cc_289 N_A_27_79#_c_295_p N_SCE_c_362_n 0.0123483f $X=2.275 $Y=2.405 $X2=0 $Y2=0
cc_290 N_A_27_79#_c_284_n N_SCE_c_362_n 0.0109466f $X=2.44 $Y=1.995 $X2=0 $Y2=0
cc_291 N_A_27_79#_c_276_n N_SCE_c_363_n 0.00219996f $X=1.4 $Y=1.415 $X2=0 $Y2=0
cc_292 N_A_27_79#_c_279_n N_SCE_c_363_n 0.0155382f $X=1.23 $Y=1.415 $X2=0 $Y2=0
cc_293 N_A_27_79#_c_281_n N_SCE_c_364_n 0.00192643f $X=2.615 $Y=2.245 $X2=0
+ $Y2=0
cc_294 N_A_27_79#_c_284_n N_SCE_c_364_n 0.0221869f $X=2.44 $Y=1.995 $X2=0 $Y2=0
cc_295 N_A_27_79#_c_281_n N_SCE_c_365_n 0.0202521f $X=2.615 $Y=2.245 $X2=0 $Y2=0
cc_296 N_A_27_79#_c_284_n N_SCE_c_365_n 7.02495e-19 $X=2.44 $Y=1.995 $X2=0 $Y2=0
cc_297 N_A_27_79#_c_276_n N_SCE_c_370_n 0.0448734f $X=1.4 $Y=1.415 $X2=0 $Y2=0
cc_298 N_A_27_79#_c_279_n N_SCE_c_370_n 0.00247218f $X=1.23 $Y=1.415 $X2=0 $Y2=0
cc_299 N_A_27_79#_c_295_p N_SCE_c_370_n 0.0171512f $X=2.275 $Y=2.405 $X2=0 $Y2=0
cc_300 N_A_27_79#_c_276_n N_SCE_c_371_n 0.00363355f $X=1.4 $Y=1.415 $X2=0 $Y2=0
cc_301 N_A_27_79#_c_278_n N_SCE_c_371_n 0.0192999f $X=0.2 $Y=2.32 $X2=0 $Y2=0
cc_302 N_A_27_79#_c_279_n N_SCE_c_371_n 0.0494351f $X=1.23 $Y=1.415 $X2=0 $Y2=0
cc_303 N_A_27_79#_c_295_p N_SCE_c_371_n 0.0736349f $X=2.275 $Y=2.405 $X2=0 $Y2=0
cc_304 N_A_27_79#_c_281_n N_D_c_444_n 0.0130861f $X=2.615 $Y=2.245 $X2=0 $Y2=0
cc_305 N_A_27_79#_c_276_n N_D_c_444_n 0.0185925f $X=1.4 $Y=1.415 $X2=0 $Y2=0
cc_306 N_A_27_79#_c_279_n N_D_c_444_n 6.63701e-19 $X=1.23 $Y=1.415 $X2=0 $Y2=0
cc_307 N_A_27_79#_c_284_n N_D_c_444_n 0.00129661f $X=2.44 $Y=1.995 $X2=0 $Y2=0
cc_308 N_A_27_79#_c_281_n N_D_c_449_n 0.0173318f $X=2.615 $Y=2.245 $X2=0 $Y2=0
cc_309 N_A_27_79#_c_295_p N_D_c_449_n 0.0174363f $X=2.275 $Y=2.405 $X2=0 $Y2=0
cc_310 N_A_27_79#_c_284_n N_D_c_449_n 0.00352705f $X=2.44 $Y=1.995 $X2=0 $Y2=0
cc_311 N_A_27_79#_M1007_g N_D_c_445_n 0.0200462f $X=1.475 $Y=0.605 $X2=0 $Y2=0
cc_312 N_A_27_79#_M1007_g N_D_c_446_n 0.0109288f $X=1.475 $Y=0.605 $X2=0 $Y2=0
cc_313 N_A_27_79#_M1007_g N_D_c_447_n 0.03521f $X=1.475 $Y=0.605 $X2=0 $Y2=0
cc_314 N_A_27_79#_c_281_n N_SCD_c_495_n 0.0359696f $X=2.615 $Y=2.245 $X2=-0.19
+ $Y2=-0.245
cc_315 N_A_27_79#_c_284_n N_SCD_c_495_n 3.88432e-19 $X=2.44 $Y=1.995 $X2=-0.19
+ $Y2=-0.245
cc_316 N_A_27_79#_c_281_n N_SCD_c_492_n 0.0223785f $X=2.615 $Y=2.245 $X2=0 $Y2=0
cc_317 N_A_27_79#_c_284_n N_SCD_c_492_n 0.00149955f $X=2.44 $Y=1.995 $X2=0 $Y2=0
cc_318 N_A_27_79#_c_281_n SCD 0.00131261f $X=2.615 $Y=2.245 $X2=0 $Y2=0
cc_319 N_A_27_79#_c_284_n SCD 0.0137554f $X=2.44 $Y=1.995 $X2=0 $Y2=0
cc_320 N_A_27_79#_c_295_p N_VPWR_M1026_d 0.0181551f $X=2.275 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_321 N_A_27_79#_c_281_n N_VPWR_c_1673_n 0.00300876f $X=2.615 $Y=2.245 $X2=0
+ $Y2=0
cc_322 N_A_27_79#_c_283_n N_VPWR_c_1679_n 0.0145785f $X=0.28 $Y=2.65 $X2=0 $Y2=0
cc_323 N_A_27_79#_c_283_n N_VPWR_c_1680_n 0.0102732f $X=0.28 $Y=2.65 $X2=0 $Y2=0
cc_324 N_A_27_79#_c_295_p N_VPWR_c_1680_n 0.0418977f $X=2.275 $Y=2.405 $X2=0
+ $Y2=0
cc_325 N_A_27_79#_c_281_n N_VPWR_c_1658_n 0.00370805f $X=2.615 $Y=2.245 $X2=0
+ $Y2=0
cc_326 N_A_27_79#_c_283_n N_VPWR_c_1658_n 0.0120406f $X=0.28 $Y=2.65 $X2=0 $Y2=0
cc_327 N_A_27_79#_c_295_p N_VPWR_c_1658_n 0.0250254f $X=2.275 $Y=2.405 $X2=0
+ $Y2=0
cc_328 N_A_27_79#_c_295_p A_307_464# 0.00479553f $X=2.275 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_329 N_A_27_79#_c_295_p N_A_388_79#_M1018_d 0.0167952f $X=2.275 $Y=2.405 $X2=0
+ $Y2=0
cc_330 N_A_27_79#_c_281_n N_A_388_79#_c_1865_n 0.0181967f $X=2.615 $Y=2.245
+ $X2=0 $Y2=0
cc_331 N_A_27_79#_c_295_p N_A_388_79#_c_1865_n 0.0419607f $X=2.275 $Y=2.405
+ $X2=0 $Y2=0
cc_332 N_A_27_79#_c_281_n N_A_388_79#_c_1867_n 0.00384668f $X=2.615 $Y=2.245
+ $X2=0 $Y2=0
cc_333 N_A_27_79#_c_281_n N_A_388_79#_c_1856_n 0.0012654f $X=2.615 $Y=2.245
+ $X2=0 $Y2=0
cc_334 N_A_27_79#_c_295_p N_A_388_79#_c_1856_n 0.0148585f $X=2.275 $Y=2.405
+ $X2=0 $Y2=0
cc_335 N_A_27_79#_M1007_g N_VGND_c_2052_n 5.90987e-19 $X=1.475 $Y=0.605 $X2=0
+ $Y2=0
cc_336 N_A_27_79#_c_276_n N_VGND_c_2052_n 0.00297438f $X=1.4 $Y=1.415 $X2=0
+ $Y2=0
cc_337 N_A_27_79#_c_277_n N_VGND_c_2052_n 0.0179429f $X=0.28 $Y=0.605 $X2=0
+ $Y2=0
cc_338 N_A_27_79#_c_279_n N_VGND_c_2052_n 0.0148785f $X=1.23 $Y=1.415 $X2=0
+ $Y2=0
cc_339 N_A_27_79#_M1007_g N_VGND_c_2062_n 9.44495e-19 $X=1.475 $Y=0.605 $X2=0
+ $Y2=0
cc_340 N_A_27_79#_c_277_n N_VGND_c_2068_n 0.0100552f $X=0.28 $Y=0.605 $X2=0
+ $Y2=0
cc_341 N_A_27_79#_c_277_n N_VGND_c_2078_n 0.00902019f $X=0.28 $Y=0.605 $X2=0
+ $Y2=0
cc_342 N_A_27_79#_M1007_g N_noxref_25_c_2207_n 7.43016e-19 $X=1.475 $Y=0.605
+ $X2=0 $Y2=0
cc_343 N_A_27_79#_c_276_n N_noxref_25_c_2207_n 0.0048989f $X=1.4 $Y=1.415 $X2=0
+ $Y2=0
cc_344 N_A_27_79#_c_279_n N_noxref_25_c_2207_n 0.0106151f $X=1.23 $Y=1.415 $X2=0
+ $Y2=0
cc_345 N_A_27_79#_M1007_g N_noxref_25_c_2208_n 0.0154771f $X=1.475 $Y=0.605
+ $X2=0 $Y2=0
cc_346 N_SCE_c_368_n N_D_c_444_n 0.0238606f $X=1.46 $Y=2.245 $X2=0 $Y2=0
cc_347 N_SCE_M1028_g N_D_c_444_n 8.48778e-19 $X=2.66 $Y=0.605 $X2=0 $Y2=0
cc_348 N_SCE_c_362_n N_D_c_444_n 0.0202953f $X=1.71 $Y=1.82 $X2=0 $Y2=0
cc_349 N_SCE_c_363_n N_D_c_444_n 0.00239218f $X=1.795 $Y=1.49 $X2=0 $Y2=0
cc_350 N_SCE_c_364_n N_D_c_444_n 0.0188764f $X=2.57 $Y=1.455 $X2=0 $Y2=0
cc_351 N_SCE_c_365_n N_D_c_444_n 0.00894005f $X=2.57 $Y=1.455 $X2=0 $Y2=0
cc_352 N_SCE_c_368_n N_D_c_449_n 0.0403591f $X=1.46 $Y=2.245 $X2=0 $Y2=0
cc_353 N_SCE_M1028_g N_D_c_445_n 0.00730331f $X=2.66 $Y=0.605 $X2=0 $Y2=0
cc_354 N_SCE_c_363_n N_D_c_445_n 7.56204e-19 $X=1.795 $Y=1.49 $X2=0 $Y2=0
cc_355 N_SCE_c_364_n N_D_c_445_n 0.002936f $X=2.57 $Y=1.455 $X2=0 $Y2=0
cc_356 N_SCE_M1028_g N_D_c_446_n 5.42624e-19 $X=2.66 $Y=0.605 $X2=0 $Y2=0
cc_357 N_SCE_c_363_n N_D_c_446_n 0.0150217f $X=1.795 $Y=1.49 $X2=0 $Y2=0
cc_358 N_SCE_c_364_n N_D_c_446_n 0.0224216f $X=2.57 $Y=1.455 $X2=0 $Y2=0
cc_359 N_SCE_c_371_n N_D_c_446_n 0.0020111f $X=1.625 $Y=1.985 $X2=0 $Y2=0
cc_360 N_SCE_M1028_g N_D_c_447_n 0.00705002f $X=2.66 $Y=0.605 $X2=0 $Y2=0
cc_361 N_SCE_M1028_g N_SCD_M1008_g 0.0628756f $X=2.66 $Y=0.605 $X2=0 $Y2=0
cc_362 N_SCE_c_364_n N_SCD_M1008_g 5.04484e-19 $X=2.57 $Y=1.455 $X2=0 $Y2=0
cc_363 N_SCE_c_364_n SCD 0.0120234f $X=2.57 $Y=1.455 $X2=0 $Y2=0
cc_364 N_SCE_c_365_n SCD 2.2546e-19 $X=2.57 $Y=1.455 $X2=0 $Y2=0
cc_365 N_SCE_c_364_n N_SCD_c_494_n 6.19299e-19 $X=2.57 $Y=1.455 $X2=0 $Y2=0
cc_366 N_SCE_c_365_n N_SCD_c_494_n 0.0113035f $X=2.57 $Y=1.455 $X2=0 $Y2=0
cc_367 N_SCE_c_368_n N_VPWR_c_1673_n 0.00413917f $X=1.46 $Y=2.245 $X2=0 $Y2=0
cc_368 N_SCE_c_367_n N_VPWR_c_1679_n 0.00445602f $X=0.505 $Y=2.245 $X2=0 $Y2=0
cc_369 N_SCE_c_367_n N_VPWR_c_1680_n 0.0101493f $X=0.505 $Y=2.245 $X2=0 $Y2=0
cc_370 N_SCE_c_368_n N_VPWR_c_1680_n 0.0101104f $X=1.46 $Y=2.245 $X2=0 $Y2=0
cc_371 N_SCE_c_367_n N_VPWR_c_1658_n 0.00460319f $X=0.505 $Y=2.245 $X2=0 $Y2=0
cc_372 N_SCE_c_368_n N_VPWR_c_1658_n 0.00412661f $X=1.46 $Y=2.245 $X2=0 $Y2=0
cc_373 N_SCE_c_368_n N_A_388_79#_c_1865_n 8.44751e-19 $X=1.46 $Y=2.245 $X2=0
+ $Y2=0
cc_374 N_SCE_M1028_g N_A_388_79#_c_1847_n 0.0103246f $X=2.66 $Y=0.605 $X2=0
+ $Y2=0
cc_375 N_SCE_M1028_g N_A_388_79#_c_1848_n 0.0087327f $X=2.66 $Y=0.605 $X2=0
+ $Y2=0
cc_376 N_SCE_c_364_n N_A_388_79#_c_1848_n 0.00815275f $X=2.57 $Y=1.455 $X2=0
+ $Y2=0
cc_377 N_SCE_M1028_g N_A_388_79#_c_1849_n 0.00327429f $X=2.66 $Y=0.605 $X2=0
+ $Y2=0
cc_378 N_SCE_c_364_n N_A_388_79#_c_1849_n 0.0273677f $X=2.57 $Y=1.455 $X2=0
+ $Y2=0
cc_379 N_SCE_c_365_n N_A_388_79#_c_1849_n 0.00449985f $X=2.57 $Y=1.455 $X2=0
+ $Y2=0
cc_380 N_SCE_c_359_n N_VGND_c_2052_n 0.0143331f $X=0.495 $Y=0.89 $X2=0 $Y2=0
cc_381 N_SCE_M1028_g N_VGND_c_2062_n 9.44495e-19 $X=2.66 $Y=0.605 $X2=0 $Y2=0
cc_382 N_SCE_c_359_n N_VGND_c_2068_n 0.00465077f $X=0.495 $Y=0.89 $X2=0 $Y2=0
cc_383 N_SCE_c_359_n N_VGND_c_2078_n 0.00451796f $X=0.495 $Y=0.89 $X2=0 $Y2=0
cc_384 N_SCE_c_359_n N_noxref_25_c_2207_n 7.27954e-19 $X=0.495 $Y=0.89 $X2=0
+ $Y2=0
cc_385 N_SCE_M1028_g N_noxref_25_c_2208_n 0.0128121f $X=2.66 $Y=0.605 $X2=0
+ $Y2=0
cc_386 N_SCE_c_359_n N_noxref_25_c_2209_n 6.46792e-19 $X=0.495 $Y=0.89 $X2=0
+ $Y2=0
cc_387 N_SCE_M1028_g N_noxref_25_c_2210_n 0.00151906f $X=2.66 $Y=0.605 $X2=0
+ $Y2=0
cc_388 N_D_c_449_n N_VPWR_c_1673_n 0.00445405f $X=1.88 $Y=2.245 $X2=0 $Y2=0
cc_389 N_D_c_449_n N_VPWR_c_1680_n 0.00139022f $X=1.88 $Y=2.245 $X2=0 $Y2=0
cc_390 N_D_c_449_n N_VPWR_c_1658_n 0.00457269f $X=1.88 $Y=2.245 $X2=0 $Y2=0
cc_391 N_D_c_446_n N_A_388_79#_M1023_d 0.00145733f $X=1.925 $Y=1.09 $X2=-0.19
+ $Y2=-0.245
cc_392 N_D_c_449_n N_A_388_79#_c_1865_n 0.00949498f $X=1.88 $Y=2.245 $X2=0 $Y2=0
cc_393 N_D_c_445_n N_A_388_79#_c_1847_n 3.29098e-19 $X=1.925 $Y=1.09 $X2=0 $Y2=0
cc_394 N_D_c_446_n N_A_388_79#_c_1847_n 0.0164816f $X=1.925 $Y=1.09 $X2=0 $Y2=0
cc_395 N_D_c_447_n N_A_388_79#_c_1847_n 0.00523412f $X=1.925 $Y=0.925 $X2=0
+ $Y2=0
cc_396 N_D_c_445_n N_A_388_79#_c_1849_n 7.8315e-19 $X=1.925 $Y=1.09 $X2=0 $Y2=0
cc_397 N_D_c_446_n N_A_388_79#_c_1849_n 0.0148785f $X=1.925 $Y=1.09 $X2=0 $Y2=0
cc_398 N_D_c_447_n N_VGND_c_2062_n 9.44495e-19 $X=1.925 $Y=0.925 $X2=0 $Y2=0
cc_399 N_D_c_446_n N_noxref_25_c_2207_n 0.00134475f $X=1.925 $Y=1.09 $X2=0 $Y2=0
cc_400 N_D_c_445_n N_noxref_25_c_2208_n 5.75063e-19 $X=1.925 $Y=1.09 $X2=0 $Y2=0
cc_401 N_D_c_446_n N_noxref_25_c_2208_n 0.0127007f $X=1.925 $Y=1.09 $X2=0 $Y2=0
cc_402 N_D_c_447_n N_noxref_25_c_2208_n 0.0123465f $X=1.925 $Y=0.925 $X2=0 $Y2=0
cc_403 N_D_c_446_n noxref_26 0.00197445f $X=1.925 $Y=1.09 $X2=-0.19 $Y2=-0.245
cc_404 N_SCD_M1008_g N_RESET_B_M1000_g 0.0292104f $X=3.05 $Y=0.605 $X2=0 $Y2=0
cc_405 SCD N_RESET_B_M1000_g 7.60177e-19 $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_406 N_SCD_c_494_n N_RESET_B_M1000_g 0.0196966f $X=3.11 $Y=1.605 $X2=0 $Y2=0
cc_407 N_SCD_c_495_n N_RESET_B_c_875_n 0.0148826f $X=3.035 $Y=2.245 $X2=0 $Y2=0
cc_408 N_SCD_c_492_n N_RESET_B_c_886_n 0.0237049f $X=3.11 $Y=1.945 $X2=0 $Y2=0
cc_409 N_SCD_c_495_n N_VPWR_c_1659_n 0.00395262f $X=3.035 $Y=2.245 $X2=0 $Y2=0
cc_410 N_SCD_c_495_n N_VPWR_c_1673_n 0.00461464f $X=3.035 $Y=2.245 $X2=0 $Y2=0
cc_411 N_SCD_c_495_n N_VPWR_c_1658_n 0.00463738f $X=3.035 $Y=2.245 $X2=0 $Y2=0
cc_412 N_SCD_M1008_g N_A_388_79#_c_1847_n 0.00151803f $X=3.05 $Y=0.605 $X2=0
+ $Y2=0
cc_413 N_SCD_M1008_g N_A_388_79#_c_1848_n 0.0127975f $X=3.05 $Y=0.605 $X2=0
+ $Y2=0
cc_414 SCD N_A_388_79#_c_1848_n 0.0182456f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_415 N_SCD_c_494_n N_A_388_79#_c_1848_n 0.00113125f $X=3.11 $Y=1.605 $X2=0
+ $Y2=0
cc_416 N_SCD_c_495_n N_A_388_79#_c_1888_n 0.011884f $X=3.035 $Y=2.245 $X2=0
+ $Y2=0
cc_417 N_SCD_c_492_n N_A_388_79#_c_1888_n 8.43385e-19 $X=3.11 $Y=1.945 $X2=0
+ $Y2=0
cc_418 SCD N_A_388_79#_c_1888_n 0.023597f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_419 N_SCD_c_495_n N_A_388_79#_c_1850_n 0.00133602f $X=3.035 $Y=2.245 $X2=0
+ $Y2=0
cc_420 N_SCD_M1008_g N_A_388_79#_c_1850_n 0.00475298f $X=3.05 $Y=0.605 $X2=0
+ $Y2=0
cc_421 N_SCD_c_492_n N_A_388_79#_c_1850_n 0.00181866f $X=3.11 $Y=1.945 $X2=0
+ $Y2=0
cc_422 SCD N_A_388_79#_c_1850_n 0.0534506f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_423 N_SCD_c_494_n N_A_388_79#_c_1850_n 0.00361663f $X=3.11 $Y=1.605 $X2=0
+ $Y2=0
cc_424 N_SCD_c_495_n N_A_388_79#_c_1858_n 3.22195e-19 $X=3.035 $Y=2.245 $X2=0
+ $Y2=0
cc_425 N_SCD_M1008_g N_VGND_c_2053_n 2.27924e-19 $X=3.05 $Y=0.605 $X2=0 $Y2=0
cc_426 N_SCD_M1008_g N_VGND_c_2062_n 9.63557e-19 $X=3.05 $Y=0.605 $X2=0 $Y2=0
cc_427 N_SCD_M1008_g N_noxref_25_c_2208_n 0.0110567f $X=3.05 $Y=0.605 $X2=0
+ $Y2=0
cc_428 N_SCD_M1008_g N_noxref_25_c_2210_n 0.00775324f $X=3.05 $Y=0.605 $X2=0
+ $Y2=0
cc_429 N_CLK_c_535_n N_A_1025_119#_c_589_n 3.98191e-19 $X=4.62 $Y=1.445 $X2=0
+ $Y2=0
cc_430 N_CLK_M1032_g N_A_1025_119#_c_590_n 8.53953e-19 $X=4.645 $Y=2.46 $X2=0
+ $Y2=0
cc_431 N_CLK_c_535_n N_RESET_B_M1000_g 0.0266275f $X=4.62 $Y=1.445 $X2=0 $Y2=0
cc_432 CLK N_RESET_B_M1000_g 0.00170133f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_433 N_CLK_c_535_n N_RESET_B_c_866_n 0.0102778f $X=4.62 $Y=1.445 $X2=0 $Y2=0
cc_434 N_CLK_c_535_n N_RESET_B_c_881_n 0.00244269f $X=4.62 $Y=1.445 $X2=0 $Y2=0
cc_435 N_CLK_M1032_g N_RESET_B_c_881_n 0.00240281f $X=4.645 $Y=2.46 $X2=0 $Y2=0
cc_436 CLK N_RESET_B_c_881_n 2.97792e-19 $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_437 N_CLK_c_535_n N_RESET_B_c_882_n 0.00157986f $X=4.62 $Y=1.445 $X2=0 $Y2=0
cc_438 CLK N_RESET_B_c_882_n 0.00364034f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_439 N_CLK_c_535_n N_RESET_B_c_886_n 0.0165248f $X=4.62 $Y=1.445 $X2=0 $Y2=0
cc_440 N_CLK_M1032_g N_RESET_B_c_886_n 0.00537889f $X=4.645 $Y=2.46 $X2=0 $Y2=0
cc_441 CLK N_RESET_B_c_886_n 6.66082e-19 $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_442 N_CLK_c_535_n N_RESET_B_c_887_n 0.00233965f $X=4.62 $Y=1.445 $X2=0 $Y2=0
cc_443 N_CLK_M1032_g N_RESET_B_c_887_n 3.35987e-19 $X=4.645 $Y=2.46 $X2=0 $Y2=0
cc_444 CLK N_RESET_B_c_887_n 0.012296f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_445 N_CLK_c_535_n N_A_852_119#_c_1176_n 0.0230093f $X=4.62 $Y=1.445 $X2=0
+ $Y2=0
cc_446 N_CLK_M1032_g N_A_852_119#_M1035_g 0.0417462f $X=4.645 $Y=2.46 $X2=0
+ $Y2=0
cc_447 N_CLK_c_535_n N_A_852_119#_c_1184_n 0.0123834f $X=4.62 $Y=1.445 $X2=0
+ $Y2=0
cc_448 CLK N_A_852_119#_c_1184_n 0.0207634f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_449 N_CLK_c_535_n N_A_852_119#_c_1185_n 0.0104784f $X=4.62 $Y=1.445 $X2=0
+ $Y2=0
cc_450 N_CLK_c_535_n N_A_852_119#_c_1186_n 0.0415927f $X=4.62 $Y=1.445 $X2=0
+ $Y2=0
cc_451 N_CLK_M1032_g N_A_852_119#_c_1186_n 0.00994609f $X=4.645 $Y=2.46 $X2=0
+ $Y2=0
cc_452 CLK N_A_852_119#_c_1186_n 0.00838159f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_453 N_CLK_c_535_n N_A_852_119#_c_1187_n 0.0215538f $X=4.62 $Y=1.445 $X2=0
+ $Y2=0
cc_454 N_CLK_M1032_g N_VPWR_c_1660_n 0.0164315f $X=4.645 $Y=2.46 $X2=0 $Y2=0
cc_455 N_CLK_M1032_g N_VPWR_c_1669_n 0.00303184f $X=4.645 $Y=2.46 $X2=0 $Y2=0
cc_456 N_CLK_M1032_g N_VPWR_c_1658_n 0.00397656f $X=4.645 $Y=2.46 $X2=0 $Y2=0
cc_457 N_CLK_c_535_n N_A_388_79#_c_1850_n 0.00163069f $X=4.62 $Y=1.445 $X2=0
+ $Y2=0
cc_458 CLK N_A_388_79#_c_1850_n 0.0174094f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_459 N_CLK_M1032_g N_A_388_79#_c_1858_n 0.01216f $X=4.645 $Y=2.46 $X2=0 $Y2=0
cc_460 N_CLK_M1032_g N_A_388_79#_c_1859_n 0.00649693f $X=4.645 $Y=2.46 $X2=0
+ $Y2=0
cc_461 N_CLK_c_535_n N_A_388_79#_c_1862_n 6.9817e-19 $X=4.62 $Y=1.445 $X2=0
+ $Y2=0
cc_462 N_CLK_M1032_g N_A_388_79#_c_1902_n 0.00900509f $X=4.645 $Y=2.46 $X2=0
+ $Y2=0
cc_463 N_CLK_c_535_n N_VGND_c_2053_n 0.00604615f $X=4.62 $Y=1.445 $X2=0 $Y2=0
cc_464 CLK N_VGND_c_2053_n 0.00344374f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_465 N_CLK_c_535_n N_VGND_c_2054_n 0.00381935f $X=4.62 $Y=1.445 $X2=0 $Y2=0
cc_466 N_CLK_c_535_n N_VGND_c_2078_n 9.39239e-19 $X=4.62 $Y=1.445 $X2=0 $Y2=0
cc_467 N_A_1025_119#_c_586_n N_A_1370_290#_M1002_d 0.00176891f $X=9.1 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_468 N_A_1025_119#_c_596_n N_A_1370_290#_c_776_n 0.00201631f $X=6.1 $Y=2.12
+ $X2=0 $Y2=0
cc_469 N_A_1025_119#_M1011_g N_A_1370_290#_M1040_g 0.0462355f $X=6.54 $Y=0.805
+ $X2=0 $Y2=0
cc_470 N_A_1025_119#_c_582_n N_A_1370_290#_M1040_g 0.00762221f $X=7 $Y=0.395
+ $X2=0 $Y2=0
cc_471 N_A_1025_119#_c_591_n N_A_1370_290#_M1040_g 0.00542036f $X=7.085 $Y=0.395
+ $X2=0 $Y2=0
cc_472 N_A_1025_119#_c_597_n N_A_1370_290#_c_777_n 0.00201631f $X=6.1 $Y=2.21
+ $X2=0 $Y2=0
cc_473 N_A_1025_119#_M1011_g N_A_1370_290#_c_772_n 0.0105382f $X=6.54 $Y=0.805
+ $X2=0 $Y2=0
cc_474 N_A_1025_119#_c_591_n N_A_1370_290#_c_772_n 3.83611e-19 $X=7.085 $Y=0.395
+ $X2=0 $Y2=0
cc_475 N_A_1025_119#_c_595_n N_A_1370_290#_c_772_n 0.00192784f $X=6.045 $Y=1.575
+ $X2=0 $Y2=0
cc_476 N_A_1025_119#_c_585_n N_A_1370_290#_c_791_n 0.00146445f $X=8.155 $Y=0.665
+ $X2=0 $Y2=0
cc_477 N_A_1025_119#_c_591_n N_A_1370_290#_c_791_n 0.00967347f $X=7.085 $Y=0.395
+ $X2=0 $Y2=0
cc_478 N_A_1025_119#_c_598_n N_A_1370_290#_c_793_n 3.85264e-19 $X=9.7 $Y=2.28
+ $X2=0 $Y2=0
cc_479 N_A_1025_119#_c_600_n N_A_1370_290#_c_793_n 0.0194716f $X=9.615 $Y=2.03
+ $X2=0 $Y2=0
cc_480 N_A_1025_119#_c_598_n N_A_1370_290#_c_780_n 0.00120571f $X=9.7 $Y=2.28
+ $X2=0 $Y2=0
cc_481 N_A_1025_119#_c_585_n N_A_1370_290#_c_773_n 0.0737203f $X=8.155 $Y=0.665
+ $X2=0 $Y2=0
cc_482 N_A_1025_119#_c_586_n N_A_1370_290#_c_773_n 0.00353238f $X=9.1 $Y=0.34
+ $X2=0 $Y2=0
cc_483 N_A_1025_119#_c_578_n N_A_1370_290#_c_774_n 0.0120063f $X=8.875 $Y=1.09
+ $X2=0 $Y2=0
cc_484 N_A_1025_119#_c_586_n N_A_1370_290#_c_774_n 0.0229775f $X=9.1 $Y=0.34
+ $X2=0 $Y2=0
cc_485 N_A_1025_119#_c_588_n N_A_1370_290#_c_774_n 0.0234316f $X=9.185 $Y=0.905
+ $X2=0 $Y2=0
cc_486 N_A_1025_119#_c_592_n N_A_1370_290#_c_774_n 0.0158022f $X=9.475 $Y=1.07
+ $X2=0 $Y2=0
cc_487 N_A_1025_119#_c_580_n N_A_1370_290#_c_775_n 0.00714514f $X=8.95 $Y=1.165
+ $X2=0 $Y2=0
cc_488 N_A_1025_119#_c_592_n N_A_1370_290#_c_775_n 0.0107601f $X=9.475 $Y=1.07
+ $X2=0 $Y2=0
cc_489 N_A_1025_119#_c_594_n N_A_1370_290#_c_775_n 0.0194716f $X=9.532 $Y=1.865
+ $X2=0 $Y2=0
cc_490 N_A_1025_119#_M1011_g N_RESET_B_c_866_n 0.00880557f $X=6.54 $Y=0.805
+ $X2=0 $Y2=0
cc_491 N_A_1025_119#_c_582_n N_RESET_B_c_866_n 0.0286159f $X=7 $Y=0.395 $X2=0
+ $Y2=0
cc_492 N_A_1025_119#_c_583_n N_RESET_B_c_866_n 0.00755311f $X=5.43 $Y=0.395
+ $X2=0 $Y2=0
cc_493 N_A_1025_119#_c_591_n N_RESET_B_c_866_n 0.00357516f $X=7.085 $Y=0.395
+ $X2=0 $Y2=0
cc_494 N_A_1025_119#_c_585_n N_RESET_B_M1006_g 0.0123884f $X=8.155 $Y=0.665
+ $X2=0 $Y2=0
cc_495 N_A_1025_119#_c_591_n N_RESET_B_M1006_g 0.00727728f $X=7.085 $Y=0.395
+ $X2=0 $Y2=0
cc_496 N_A_1025_119#_c_596_n N_RESET_B_c_881_n 0.00557922f $X=6.1 $Y=2.12 $X2=0
+ $Y2=0
cc_497 N_A_1025_119#_c_576_n N_RESET_B_c_881_n 0.00395271f $X=6.465 $Y=1.575
+ $X2=0 $Y2=0
cc_498 N_A_1025_119#_c_590_n N_RESET_B_c_881_n 0.0617736f $X=5.56 $Y=1.87 $X2=0
+ $Y2=0
cc_499 N_A_1025_119#_c_595_n N_RESET_B_c_881_n 4.9282e-19 $X=6.045 $Y=1.575
+ $X2=0 $Y2=0
cc_500 N_A_1025_119#_c_598_n N_RESET_B_c_883_n 0.00170256f $X=9.7 $Y=2.28 $X2=0
+ $Y2=0
cc_501 N_A_1025_119#_c_600_n N_RESET_B_c_883_n 0.0277328f $X=9.615 $Y=2.03 $X2=0
+ $Y2=0
cc_502 N_A_1025_119#_c_578_n N_A_1223_119#_M1002_g 0.026603f $X=8.875 $Y=1.09
+ $X2=0 $Y2=0
cc_503 N_A_1025_119#_c_586_n N_A_1223_119#_M1002_g 0.0116384f $X=9.1 $Y=0.34
+ $X2=0 $Y2=0
cc_504 N_A_1025_119#_c_576_n N_A_1223_119#_c_1082_n 6.10614e-19 $X=6.465
+ $Y=1.575 $X2=0 $Y2=0
cc_505 N_A_1025_119#_M1011_g N_A_1223_119#_c_1082_n 0.0146944f $X=6.54 $Y=0.805
+ $X2=0 $Y2=0
cc_506 N_A_1025_119#_c_582_n N_A_1223_119#_c_1082_n 0.0431682f $X=7 $Y=0.395
+ $X2=0 $Y2=0
cc_507 N_A_1025_119#_c_597_n N_A_1223_119#_c_1075_n 0.00283015f $X=6.1 $Y=2.21
+ $X2=0 $Y2=0
cc_508 N_A_1025_119#_c_597_n N_A_1223_119#_c_1073_n 3.46279e-19 $X=6.1 $Y=2.21
+ $X2=0 $Y2=0
cc_509 N_A_1025_119#_M1011_g N_A_1223_119#_c_1073_n 0.00527914f $X=6.54 $Y=0.805
+ $X2=0 $Y2=0
cc_510 N_A_1025_119#_c_581_n N_A_852_119#_c_1176_n 0.00874347f $X=5.265 $Y=0.74
+ $X2=0 $Y2=0
cc_511 N_A_1025_119#_c_583_n N_A_852_119#_c_1176_n 6.62904e-19 $X=5.43 $Y=0.395
+ $X2=0 $Y2=0
cc_512 N_A_1025_119#_c_584_n N_A_852_119#_c_1176_n 0.00276356f $X=5.56 $Y=1.5
+ $X2=0 $Y2=0
cc_513 N_A_1025_119#_c_589_n N_A_852_119#_c_1176_n 0.00435367f $X=5.56 $Y=1.132
+ $X2=0 $Y2=0
cc_514 N_A_1025_119#_c_590_n N_A_852_119#_M1035_g 0.00666545f $X=5.56 $Y=1.87
+ $X2=0 $Y2=0
cc_515 N_A_1025_119#_c_584_n N_A_852_119#_c_1177_n 0.00718429f $X=5.56 $Y=1.5
+ $X2=0 $Y2=0
cc_516 N_A_1025_119#_c_589_n N_A_852_119#_c_1177_n 0.00193283f $X=5.56 $Y=1.132
+ $X2=0 $Y2=0
cc_517 N_A_1025_119#_c_596_n N_A_852_119#_c_1189_n 0.0134932f $X=6.1 $Y=2.12
+ $X2=0 $Y2=0
cc_518 N_A_1025_119#_c_597_n N_A_852_119#_c_1189_n 0.0137907f $X=6.1 $Y=2.21
+ $X2=0 $Y2=0
cc_519 N_A_1025_119#_c_590_n N_A_852_119#_c_1189_n 0.0185474f $X=5.56 $Y=1.87
+ $X2=0 $Y2=0
cc_520 N_A_1025_119#_c_590_n N_A_852_119#_c_1178_n 0.00597693f $X=5.56 $Y=1.87
+ $X2=0 $Y2=0
cc_521 N_A_1025_119#_c_595_n N_A_852_119#_c_1178_n 0.0117155f $X=6.045 $Y=1.575
+ $X2=0 $Y2=0
cc_522 N_A_1025_119#_c_582_n N_A_852_119#_c_1179_n 0.00126052f $X=7 $Y=0.395
+ $X2=0 $Y2=0
cc_523 N_A_1025_119#_c_589_n N_A_852_119#_c_1179_n 0.00907962f $X=5.56 $Y=1.132
+ $X2=0 $Y2=0
cc_524 N_A_1025_119#_c_597_n N_A_852_119#_c_1190_n 0.00899647f $X=6.1 $Y=2.21
+ $X2=0 $Y2=0
cc_525 N_A_1025_119#_M1011_g N_A_852_119#_c_1180_n 0.0192564f $X=6.54 $Y=0.805
+ $X2=0 $Y2=0
cc_526 N_A_1025_119#_c_581_n N_A_852_119#_c_1180_n 0.00427994f $X=5.265 $Y=0.74
+ $X2=0 $Y2=0
cc_527 N_A_1025_119#_c_582_n N_A_852_119#_c_1180_n 0.00544855f $X=7 $Y=0.395
+ $X2=0 $Y2=0
cc_528 N_A_1025_119#_c_589_n N_A_852_119#_c_1180_n 5.42723e-19 $X=5.56 $Y=1.132
+ $X2=0 $Y2=0
cc_529 N_A_1025_119#_c_597_n N_A_852_119#_c_1192_n 0.00278823f $X=6.1 $Y=2.21
+ $X2=0 $Y2=0
cc_530 N_A_1025_119#_c_597_n N_A_852_119#_c_1194_n 0.0128753f $X=6.1 $Y=2.21
+ $X2=0 $Y2=0
cc_531 N_A_1025_119#_c_576_n N_A_852_119#_c_1194_n 0.00375991f $X=6.465 $Y=1.575
+ $X2=0 $Y2=0
cc_532 N_A_1025_119#_c_598_n N_A_852_119#_c_1196_n 0.00247489f $X=9.7 $Y=2.28
+ $X2=0 $Y2=0
cc_533 N_A_1025_119#_c_598_n N_A_852_119#_M1004_g 0.0185475f $X=9.7 $Y=2.28
+ $X2=0 $Y2=0
cc_534 N_A_1025_119#_c_594_n N_A_852_119#_M1004_g 0.00632245f $X=9.532 $Y=1.865
+ $X2=0 $Y2=0
cc_535 N_A_1025_119#_c_579_n N_A_852_119#_c_1181_n 0.0230767f $X=9.31 $Y=1.165
+ $X2=0 $Y2=0
cc_536 N_A_1025_119#_c_598_n N_A_852_119#_c_1181_n 0.0184752f $X=9.7 $Y=2.28
+ $X2=0 $Y2=0
cc_537 N_A_1025_119#_c_592_n N_A_852_119#_c_1181_n 0.00156342f $X=9.475 $Y=1.07
+ $X2=0 $Y2=0
cc_538 N_A_1025_119#_c_600_n N_A_852_119#_c_1181_n 7.40372e-19 $X=9.615 $Y=2.03
+ $X2=0 $Y2=0
cc_539 N_A_1025_119#_c_594_n N_A_852_119#_c_1181_n 0.0189852f $X=9.532 $Y=1.865
+ $X2=0 $Y2=0
cc_540 N_A_1025_119#_c_580_n N_A_852_119#_c_1182_n 0.0230767f $X=8.95 $Y=1.165
+ $X2=0 $Y2=0
cc_541 N_A_1025_119#_c_594_n N_A_852_119#_c_1182_n 7.05953e-19 $X=9.532 $Y=1.865
+ $X2=0 $Y2=0
cc_542 N_A_1025_119#_c_586_n N_A_852_119#_M1045_g 0.00370958f $X=9.1 $Y=0.34
+ $X2=0 $Y2=0
cc_543 N_A_1025_119#_c_588_n N_A_852_119#_M1045_g 0.00214927f $X=9.185 $Y=0.905
+ $X2=0 $Y2=0
cc_544 N_A_1025_119#_c_592_n N_A_852_119#_M1045_g 0.00105258f $X=9.475 $Y=1.07
+ $X2=0 $Y2=0
cc_545 N_A_1025_119#_c_593_n N_A_852_119#_M1045_g 0.0199966f $X=9.475 $Y=1.07
+ $X2=0 $Y2=0
cc_546 N_A_1025_119#_c_594_n N_A_852_119#_M1045_g 0.00469019f $X=9.532 $Y=1.865
+ $X2=0 $Y2=0
cc_547 N_A_1025_119#_c_589_n N_A_852_119#_c_1184_n 0.00426584f $X=5.56 $Y=1.132
+ $X2=0 $Y2=0
cc_548 N_A_1025_119#_c_584_n N_A_852_119#_c_1186_n 0.00415559f $X=5.56 $Y=1.5
+ $X2=0 $Y2=0
cc_549 N_A_1025_119#_c_589_n N_A_852_119#_c_1186_n 0.0134677f $X=5.56 $Y=1.132
+ $X2=0 $Y2=0
cc_550 N_A_1025_119#_c_590_n N_A_852_119#_c_1186_n 0.0493185f $X=5.56 $Y=1.87
+ $X2=0 $Y2=0
cc_551 N_A_1025_119#_c_584_n N_A_852_119#_c_1187_n 0.00254352f $X=5.56 $Y=1.5
+ $X2=0 $Y2=0
cc_552 N_A_1025_119#_c_589_n N_A_852_119#_c_1187_n 0.00333735f $X=5.56 $Y=1.132
+ $X2=0 $Y2=0
cc_553 N_A_1025_119#_c_590_n N_A_852_119#_c_1187_n 0.0167058f $X=5.56 $Y=1.87
+ $X2=0 $Y2=0
cc_554 N_A_1025_119#_c_595_n N_A_852_119#_c_1187_n 0.0214737f $X=6.045 $Y=1.575
+ $X2=0 $Y2=0
cc_555 N_A_1025_119#_c_598_n N_A_2006_373#_c_1353_n 0.0292474f $X=9.7 $Y=2.28
+ $X2=0 $Y2=0
cc_556 N_A_1025_119#_c_598_n N_A_2006_373#_c_1360_n 0.0224077f $X=9.7 $Y=2.28
+ $X2=0 $Y2=0
cc_557 N_A_1025_119#_c_600_n N_A_2006_373#_c_1360_n 3.95315e-19 $X=9.615 $Y=2.03
+ $X2=0 $Y2=0
cc_558 N_A_1025_119#_c_586_n N_A_1790_75#_M1016_d 0.00348304f $X=9.1 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_559 N_A_1025_119#_c_588_n N_A_1790_75#_M1016_d 0.0113451f $X=9.185 $Y=0.905
+ $X2=-0.19 $Y2=-0.245
cc_560 N_A_1025_119#_c_592_n N_A_1790_75#_M1016_d 0.00122753f $X=9.475 $Y=1.07
+ $X2=-0.19 $Y2=-0.245
cc_561 N_A_1025_119#_c_598_n N_A_1790_75#_c_1478_n 0.0204256f $X=9.7 $Y=2.28
+ $X2=0 $Y2=0
cc_562 N_A_1025_119#_c_600_n N_A_1790_75#_c_1478_n 0.0316971f $X=9.615 $Y=2.03
+ $X2=0 $Y2=0
cc_563 N_A_1025_119#_c_578_n N_A_1790_75#_c_1480_n 5.95394e-19 $X=8.875 $Y=1.09
+ $X2=0 $Y2=0
cc_564 N_A_1025_119#_c_586_n N_A_1790_75#_c_1480_n 0.00170833f $X=9.1 $Y=0.34
+ $X2=0 $Y2=0
cc_565 N_A_1025_119#_c_588_n N_A_1790_75#_c_1480_n 0.0250265f $X=9.185 $Y=0.905
+ $X2=0 $Y2=0
cc_566 N_A_1025_119#_c_592_n N_A_1790_75#_c_1480_n 0.0155252f $X=9.475 $Y=1.07
+ $X2=0 $Y2=0
cc_567 N_A_1025_119#_c_593_n N_A_1790_75#_c_1480_n 0.00457036f $X=9.475 $Y=1.07
+ $X2=0 $Y2=0
cc_568 N_A_1025_119#_c_588_n N_A_1790_75#_c_1464_n 0.00427034f $X=9.185 $Y=0.905
+ $X2=0 $Y2=0
cc_569 N_A_1025_119#_c_592_n N_A_1790_75#_c_1464_n 0.00683662f $X=9.475 $Y=1.07
+ $X2=0 $Y2=0
cc_570 N_A_1025_119#_c_598_n N_A_1790_75#_c_1465_n 0.00539734f $X=9.7 $Y=2.28
+ $X2=0 $Y2=0
cc_571 N_A_1025_119#_c_600_n N_A_1790_75#_c_1465_n 0.0241297f $X=9.615 $Y=2.03
+ $X2=0 $Y2=0
cc_572 N_A_1025_119#_c_594_n N_A_1790_75#_c_1465_n 0.0288004f $X=9.532 $Y=1.865
+ $X2=0 $Y2=0
cc_573 N_A_1025_119#_c_592_n N_A_1790_75#_c_1490_n 0.0103633f $X=9.475 $Y=1.07
+ $X2=0 $Y2=0
cc_574 N_A_1025_119#_c_593_n N_A_1790_75#_c_1490_n 2.34254e-19 $X=9.475 $Y=1.07
+ $X2=0 $Y2=0
cc_575 N_A_1025_119#_c_594_n N_A_1790_75#_c_1490_n 0.00424934f $X=9.532 $Y=1.865
+ $X2=0 $Y2=0
cc_576 N_A_1025_119#_c_598_n N_VPWR_c_1663_n 0.00349642f $X=9.7 $Y=2.28 $X2=0
+ $Y2=0
cc_577 N_A_1025_119#_c_597_n N_VPWR_c_1658_n 9.49986e-19 $X=6.1 $Y=2.21 $X2=0
+ $Y2=0
cc_578 N_A_1025_119#_c_598_n N_VPWR_c_1658_n 0.00489211f $X=9.7 $Y=2.28 $X2=0
+ $Y2=0
cc_579 N_A_1025_119#_M1035_d N_A_388_79#_c_1859_n 0.00633458f $X=5.17 $Y=1.96
+ $X2=0 $Y2=0
cc_580 N_A_1025_119#_c_590_n N_A_388_79#_c_1859_n 0.0321431f $X=5.56 $Y=1.87
+ $X2=0 $Y2=0
cc_581 N_A_1025_119#_M1011_g N_A_388_79#_c_1851_n 4.31453e-19 $X=6.54 $Y=0.805
+ $X2=0 $Y2=0
cc_582 N_A_1025_119#_c_581_n N_A_388_79#_c_1851_n 0.00733866f $X=5.265 $Y=0.74
+ $X2=0 $Y2=0
cc_583 N_A_1025_119#_c_589_n N_A_388_79#_c_1851_n 0.0101686f $X=5.56 $Y=1.132
+ $X2=0 $Y2=0
cc_584 N_A_1025_119#_c_597_n N_A_388_79#_c_1860_n 0.015022f $X=6.1 $Y=2.21 $X2=0
+ $Y2=0
cc_585 N_A_1025_119#_c_576_n N_A_388_79#_c_1860_n 0.00262689f $X=6.465 $Y=1.575
+ $X2=0 $Y2=0
cc_586 N_A_1025_119#_c_590_n N_A_388_79#_c_1860_n 0.00995354f $X=5.56 $Y=1.87
+ $X2=0 $Y2=0
cc_587 N_A_1025_119#_c_595_n N_A_388_79#_c_1860_n 7.55924e-19 $X=6.045 $Y=1.575
+ $X2=0 $Y2=0
cc_588 N_A_1025_119#_M1011_g N_A_388_79#_c_1852_n 0.00493912f $X=6.54 $Y=0.805
+ $X2=0 $Y2=0
cc_589 N_A_1025_119#_c_582_n N_A_388_79#_c_1852_n 0.00414539f $X=7 $Y=0.395
+ $X2=0 $Y2=0
cc_590 N_A_1025_119#_c_590_n N_A_388_79#_c_1852_n 0.0105782f $X=5.56 $Y=1.87
+ $X2=0 $Y2=0
cc_591 N_A_1025_119#_c_595_n N_A_388_79#_c_1852_n 0.00651441f $X=6.045 $Y=1.575
+ $X2=0 $Y2=0
cc_592 N_A_1025_119#_c_584_n N_A_388_79#_c_1853_n 0.00118296f $X=5.56 $Y=1.5
+ $X2=0 $Y2=0
cc_593 N_A_1025_119#_c_589_n N_A_388_79#_c_1853_n 0.0126221f $X=5.56 $Y=1.132
+ $X2=0 $Y2=0
cc_594 N_A_1025_119#_c_590_n N_A_388_79#_c_1853_n 0.012515f $X=5.56 $Y=1.87
+ $X2=0 $Y2=0
cc_595 N_A_1025_119#_c_595_n N_A_388_79#_c_1853_n 4.25051e-19 $X=6.045 $Y=1.575
+ $X2=0 $Y2=0
cc_596 N_A_1025_119#_c_596_n N_A_388_79#_c_1854_n 0.0048812f $X=6.1 $Y=2.12
+ $X2=0 $Y2=0
cc_597 N_A_1025_119#_c_576_n N_A_388_79#_c_1854_n 0.0124449f $X=6.465 $Y=1.575
+ $X2=0 $Y2=0
cc_598 N_A_1025_119#_M1011_g N_A_388_79#_c_1854_n 0.00569051f $X=6.54 $Y=0.805
+ $X2=0 $Y2=0
cc_599 N_A_1025_119#_c_584_n N_A_388_79#_c_1854_n 0.00522378f $X=5.56 $Y=1.5
+ $X2=0 $Y2=0
cc_600 N_A_1025_119#_c_590_n N_A_388_79#_c_1854_n 0.0386275f $X=5.56 $Y=1.87
+ $X2=0 $Y2=0
cc_601 N_A_1025_119#_c_595_n N_A_388_79#_c_1854_n 0.00205284f $X=6.045 $Y=1.575
+ $X2=0 $Y2=0
cc_602 N_A_1025_119#_c_581_n N_A_388_79#_c_1855_n 0.0113657f $X=5.265 $Y=0.74
+ $X2=0 $Y2=0
cc_603 N_A_1025_119#_c_582_n N_A_388_79#_c_1855_n 0.0212057f $X=7 $Y=0.395 $X2=0
+ $Y2=0
cc_604 N_A_1025_119#_c_597_n N_A_388_79#_c_1863_n 2.02597e-19 $X=6.1 $Y=2.21
+ $X2=0 $Y2=0
cc_605 N_A_1025_119#_c_590_n N_A_388_79#_c_1863_n 0.0231507f $X=5.56 $Y=1.87
+ $X2=0 $Y2=0
cc_606 N_A_1025_119#_c_595_n N_A_388_79#_c_1863_n 5.61328e-19 $X=6.045 $Y=1.575
+ $X2=0 $Y2=0
cc_607 N_A_1025_119#_c_585_n N_VGND_M1006_d 0.0231466f $X=8.155 $Y=0.665 $X2=0
+ $Y2=0
cc_608 N_A_1025_119#_c_746_p N_VGND_M1006_d 0.00612573f $X=8.24 $Y=0.58 $X2=0
+ $Y2=0
cc_609 N_A_1025_119#_c_587_n N_VGND_M1006_d 0.00119488f $X=8.325 $Y=0.34 $X2=0
+ $Y2=0
cc_610 N_A_1025_119#_c_581_n N_VGND_c_2054_n 0.0223626f $X=5.265 $Y=0.74 $X2=0
+ $Y2=0
cc_611 N_A_1025_119#_c_583_n N_VGND_c_2054_n 0.0137189f $X=5.43 $Y=0.395 $X2=0
+ $Y2=0
cc_612 N_A_1025_119#_c_578_n N_VGND_c_2066_n 0.00278271f $X=8.875 $Y=1.09 $X2=0
+ $Y2=0
cc_613 N_A_1025_119#_c_585_n N_VGND_c_2066_n 0.003347f $X=8.155 $Y=0.665 $X2=0
+ $Y2=0
cc_614 N_A_1025_119#_c_586_n N_VGND_c_2066_n 0.0611382f $X=9.1 $Y=0.34 $X2=0
+ $Y2=0
cc_615 N_A_1025_119#_c_587_n N_VGND_c_2066_n 0.0118998f $X=8.325 $Y=0.34 $X2=0
+ $Y2=0
cc_616 N_A_1025_119#_c_582_n N_VGND_c_2073_n 0.0751677f $X=7 $Y=0.395 $X2=0
+ $Y2=0
cc_617 N_A_1025_119#_c_583_n N_VGND_c_2073_n 0.0175158f $X=5.43 $Y=0.395 $X2=0
+ $Y2=0
cc_618 N_A_1025_119#_c_585_n N_VGND_c_2073_n 0.00545957f $X=8.155 $Y=0.665 $X2=0
+ $Y2=0
cc_619 N_A_1025_119#_c_591_n N_VGND_c_2073_n 0.00863901f $X=7.085 $Y=0.395 $X2=0
+ $Y2=0
cc_620 N_A_1025_119#_c_585_n N_VGND_c_2074_n 0.0398776f $X=8.155 $Y=0.665 $X2=0
+ $Y2=0
cc_621 N_A_1025_119#_c_587_n N_VGND_c_2074_n 0.0140562f $X=8.325 $Y=0.34 $X2=0
+ $Y2=0
cc_622 N_A_1025_119#_c_591_n N_VGND_c_2074_n 0.00577425f $X=7.085 $Y=0.395 $X2=0
+ $Y2=0
cc_623 N_A_1025_119#_c_578_n N_VGND_c_2078_n 0.00358525f $X=8.875 $Y=1.09 $X2=0
+ $Y2=0
cc_624 N_A_1025_119#_c_582_n N_VGND_c_2078_n 0.0507418f $X=7 $Y=0.395 $X2=0
+ $Y2=0
cc_625 N_A_1025_119#_c_583_n N_VGND_c_2078_n 0.0111521f $X=5.43 $Y=0.395 $X2=0
+ $Y2=0
cc_626 N_A_1025_119#_c_585_n N_VGND_c_2078_n 0.015012f $X=8.155 $Y=0.665 $X2=0
+ $Y2=0
cc_627 N_A_1025_119#_c_586_n N_VGND_c_2078_n 0.0343665f $X=9.1 $Y=0.34 $X2=0
+ $Y2=0
cc_628 N_A_1025_119#_c_587_n N_VGND_c_2078_n 0.00655543f $X=8.325 $Y=0.34 $X2=0
+ $Y2=0
cc_629 N_A_1025_119#_c_591_n N_VGND_c_2078_n 0.0055945f $X=7.085 $Y=0.395 $X2=0
+ $Y2=0
cc_630 N_A_1025_119#_c_585_n A_1401_119# 5.60515e-19 $X=8.155 $Y=0.665 $X2=-0.19
+ $Y2=-0.245
cc_631 N_A_1025_119#_c_591_n A_1401_119# 0.00145656f $X=7.085 $Y=0.395 $X2=-0.19
+ $Y2=-0.245
cc_632 N_A_1370_290#_M1040_g N_RESET_B_c_866_n 0.00881802f $X=6.93 $Y=0.805
+ $X2=0 $Y2=0
cc_633 N_A_1370_290#_M1040_g N_RESET_B_M1006_g 0.0413828f $X=6.93 $Y=0.805 $X2=0
+ $Y2=0
cc_634 N_A_1370_290#_c_773_n N_RESET_B_M1006_g 0.0149052f $X=8.495 $Y=0.842
+ $X2=0 $Y2=0
cc_635 N_A_1370_290#_c_773_n N_RESET_B_c_869_n 0.0110159f $X=8.495 $Y=0.842
+ $X2=0 $Y2=0
cc_636 N_A_1370_290#_c_771_n N_RESET_B_c_870_n 0.00392043f $X=7.105 $Y=1.615
+ $X2=0 $Y2=0
cc_637 N_A_1370_290#_c_772_n N_RESET_B_c_870_n 0.00184962f $X=7.105 $Y=1.615
+ $X2=0 $Y2=0
cc_638 N_A_1370_290#_c_777_n N_RESET_B_c_876_n 0.013937f $X=6.94 $Y=2.21 $X2=0
+ $Y2=0
cc_639 N_A_1370_290#_c_776_n N_RESET_B_c_871_n 0.00165672f $X=6.94 $Y=2.12 $X2=0
+ $Y2=0
cc_640 N_A_1370_290#_M1040_g N_RESET_B_c_871_n 0.00134145f $X=6.93 $Y=0.805
+ $X2=0 $Y2=0
cc_641 N_A_1370_290#_c_771_n N_RESET_B_c_871_n 4.1836e-19 $X=7.105 $Y=1.615
+ $X2=0 $Y2=0
cc_642 N_A_1370_290#_c_772_n N_RESET_B_c_871_n 0.00818789f $X=7.105 $Y=1.615
+ $X2=0 $Y2=0
cc_643 N_A_1370_290#_c_776_n N_RESET_B_c_881_n 0.0118824f $X=6.94 $Y=2.12 $X2=0
+ $Y2=0
cc_644 N_A_1370_290#_c_771_n N_RESET_B_c_881_n 0.00636364f $X=7.105 $Y=1.615
+ $X2=0 $Y2=0
cc_645 N_A_1370_290#_c_772_n N_RESET_B_c_881_n 0.00145933f $X=7.105 $Y=1.615
+ $X2=0 $Y2=0
cc_646 N_A_1370_290#_M1039_d N_RESET_B_c_883_n 0.00455663f $X=8.575 $Y=1.735
+ $X2=0 $Y2=0
cc_647 N_A_1370_290#_c_780_n N_RESET_B_c_883_n 0.0380147f $X=8.725 $Y=1.91 $X2=0
+ $Y2=0
cc_648 N_A_1370_290#_c_776_n N_RESET_B_c_888_n 0.00541842f $X=6.94 $Y=2.12 $X2=0
+ $Y2=0
cc_649 N_A_1370_290#_c_773_n N_A_1223_119#_M1002_g 0.01076f $X=8.495 $Y=0.842
+ $X2=0 $Y2=0
cc_650 N_A_1370_290#_c_774_n N_A_1223_119#_M1002_g 0.0115634f $X=8.845 $Y=0.842
+ $X2=0 $Y2=0
cc_651 N_A_1370_290#_c_775_n N_A_1223_119#_M1002_g 0.00299356f $X=8.785 $Y=1.745
+ $X2=0 $Y2=0
cc_652 N_A_1370_290#_c_793_n N_A_1223_119#_c_1069_n 0.00358587f $X=8.785 $Y=1.89
+ $X2=0 $Y2=0
cc_653 N_A_1370_290#_c_773_n N_A_1223_119#_c_1069_n 0.00251001f $X=8.495
+ $Y=0.842 $X2=0 $Y2=0
cc_654 N_A_1370_290#_c_774_n N_A_1223_119#_c_1069_n 0.00187812f $X=8.845
+ $Y=0.842 $X2=0 $Y2=0
cc_655 N_A_1370_290#_c_775_n N_A_1223_119#_c_1069_n 0.00588778f $X=8.785
+ $Y=1.745 $X2=0 $Y2=0
cc_656 N_A_1370_290#_c_777_n N_A_1223_119#_c_1095_n 0.0081651f $X=6.94 $Y=2.21
+ $X2=0 $Y2=0
cc_657 N_A_1370_290#_c_771_n N_A_1223_119#_c_1095_n 0.00227639f $X=7.105
+ $Y=1.615 $X2=0 $Y2=0
cc_658 N_A_1370_290#_c_772_n N_A_1223_119#_c_1095_n 0.0023271f $X=7.105 $Y=1.615
+ $X2=0 $Y2=0
cc_659 N_A_1370_290#_c_776_n N_A_1223_119#_c_1070_n 0.00408734f $X=6.94 $Y=2.12
+ $X2=0 $Y2=0
cc_660 N_A_1370_290#_c_777_n N_A_1223_119#_c_1070_n 0.00158906f $X=6.94 $Y=2.21
+ $X2=0 $Y2=0
cc_661 N_A_1370_290#_c_771_n N_A_1223_119#_c_1070_n 0.0148532f $X=7.105 $Y=1.615
+ $X2=0 $Y2=0
cc_662 N_A_1370_290#_c_772_n N_A_1223_119#_c_1070_n 0.00180559f $X=7.105
+ $Y=1.615 $X2=0 $Y2=0
cc_663 N_A_1370_290#_M1040_g N_A_1223_119#_c_1071_n 7.20903e-19 $X=6.93 $Y=0.805
+ $X2=0 $Y2=0
cc_664 N_A_1370_290#_c_771_n N_A_1223_119#_c_1071_n 0.0265063f $X=7.105 $Y=1.615
+ $X2=0 $Y2=0
cc_665 N_A_1370_290#_c_772_n N_A_1223_119#_c_1071_n 0.00122451f $X=7.105
+ $Y=1.615 $X2=0 $Y2=0
cc_666 N_A_1370_290#_c_773_n N_A_1223_119#_c_1071_n 0.0142918f $X=8.495 $Y=0.842
+ $X2=0 $Y2=0
cc_667 N_A_1370_290#_c_773_n N_A_1223_119#_c_1072_n 0.080152f $X=8.495 $Y=0.842
+ $X2=0 $Y2=0
cc_668 N_A_1370_290#_c_775_n N_A_1223_119#_c_1072_n 0.0250137f $X=8.785 $Y=1.745
+ $X2=0 $Y2=0
cc_669 N_A_1370_290#_c_777_n N_A_1223_119#_c_1078_n 0.00914809f $X=6.94 $Y=2.21
+ $X2=0 $Y2=0
cc_670 N_A_1370_290#_M1040_g N_A_1223_119#_c_1073_n 0.00323506f $X=6.93 $Y=0.805
+ $X2=0 $Y2=0
cc_671 N_A_1370_290#_c_777_n N_A_1223_119#_c_1073_n 0.00107886f $X=6.94 $Y=2.21
+ $X2=0 $Y2=0
cc_672 N_A_1370_290#_c_771_n N_A_1223_119#_c_1073_n 0.0500464f $X=7.105 $Y=1.615
+ $X2=0 $Y2=0
cc_673 N_A_1370_290#_c_772_n N_A_1223_119#_c_1073_n 0.0103325f $X=7.105 $Y=1.615
+ $X2=0 $Y2=0
cc_674 N_A_1370_290#_c_791_n N_A_1223_119#_c_1073_n 0.00869313f $X=7.21 $Y=1.005
+ $X2=0 $Y2=0
cc_675 N_A_1370_290#_c_777_n N_A_852_119#_c_1192_n 0.00322542f $X=6.94 $Y=2.21
+ $X2=0 $Y2=0
cc_676 N_A_1370_290#_c_777_n N_A_852_119#_c_1194_n 0.0313261f $X=6.94 $Y=2.21
+ $X2=0 $Y2=0
cc_677 N_A_1370_290#_c_777_n N_A_852_119#_c_1195_n 0.00853677f $X=6.94 $Y=2.21
+ $X2=0 $Y2=0
cc_678 N_A_1370_290#_c_780_n N_A_852_119#_c_1195_n 0.00262042f $X=8.725 $Y=1.91
+ $X2=0 $Y2=0
cc_679 N_A_1370_290#_c_780_n N_A_852_119#_c_1196_n 5.08057e-19 $X=8.725 $Y=1.91
+ $X2=0 $Y2=0
cc_680 N_A_1370_290#_c_793_n N_A_852_119#_M1004_g 0.00259852f $X=8.785 $Y=1.89
+ $X2=0 $Y2=0
cc_681 N_A_1370_290#_c_780_n N_A_852_119#_M1004_g 0.0157448f $X=8.725 $Y=1.91
+ $X2=0 $Y2=0
cc_682 N_A_1370_290#_c_775_n N_A_852_119#_M1004_g 0.00201426f $X=8.785 $Y=1.745
+ $X2=0 $Y2=0
cc_683 N_A_1370_290#_c_775_n N_A_852_119#_c_1182_n 0.00700961f $X=8.785 $Y=1.745
+ $X2=0 $Y2=0
cc_684 N_A_1370_290#_c_780_n N_A_1790_75#_c_1478_n 0.0268437f $X=8.725 $Y=1.91
+ $X2=0 $Y2=0
cc_685 N_A_1370_290#_c_777_n N_VPWR_c_1661_n 0.00337046f $X=6.94 $Y=2.21 $X2=0
+ $Y2=0
cc_686 N_A_1370_290#_c_793_n N_VPWR_c_1662_n 0.0654619f $X=8.785 $Y=1.89 $X2=0
+ $Y2=0
cc_687 N_A_1370_290#_c_780_n N_VPWR_c_1663_n 0.00650548f $X=8.725 $Y=1.91 $X2=0
+ $Y2=0
cc_688 N_A_1370_290#_c_777_n N_VPWR_c_1658_n 9.49986e-19 $X=6.94 $Y=2.21 $X2=0
+ $Y2=0
cc_689 N_A_1370_290#_c_780_n N_VPWR_c_1658_n 0.00790777f $X=8.725 $Y=1.91 $X2=0
+ $Y2=0
cc_690 N_A_1370_290#_c_773_n N_VGND_M1006_d 0.0123706f $X=8.495 $Y=0.842 $X2=0
+ $Y2=0
cc_691 N_A_1370_290#_c_791_n A_1401_119# 0.00131009f $X=7.21 $Y=1.005 $X2=-0.19
+ $Y2=-0.245
cc_692 N_RESET_B_c_869_n N_A_1223_119#_M1002_g 0.00460948f $X=7.66 $Y=1.165
+ $X2=0 $Y2=0
cc_693 N_RESET_B_c_871_n N_A_1223_119#_c_1069_n 0.0123417f $X=7.735 $Y=1.795
+ $X2=0 $Y2=0
cc_694 N_RESET_B_c_883_n N_A_1223_119#_c_1069_n 0.00747349f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_695 N_RESET_B_c_881_n N_A_1223_119#_c_1075_n 0.00709547f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_696 N_RESET_B_c_881_n N_A_1223_119#_c_1095_n 0.0165692f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_697 N_RESET_B_c_876_n N_A_1223_119#_c_1070_n 0.0168337f $X=7.525 $Y=2.21
+ $X2=0 $Y2=0
cc_698 N_RESET_B_c_871_n N_A_1223_119#_c_1070_n 0.00611723f $X=7.735 $Y=1.795
+ $X2=0 $Y2=0
cc_699 N_RESET_B_c_881_n N_A_1223_119#_c_1070_n 0.0319772f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_700 N_RESET_B_c_884_n N_A_1223_119#_c_1070_n 0.00394987f $X=8.065 $Y=2.035
+ $X2=0 $Y2=0
cc_701 N_RESET_B_c_888_n N_A_1223_119#_c_1070_n 0.0177116f $X=7.735 $Y=2.002
+ $X2=0 $Y2=0
cc_702 N_RESET_B_c_889_n N_A_1223_119#_c_1070_n 0.0379481f $X=7.825 $Y=1.96
+ $X2=0 $Y2=0
cc_703 N_RESET_B_c_870_n N_A_1223_119#_c_1071_n 0.00420432f $X=7.395 $Y=1.165
+ $X2=0 $Y2=0
cc_704 N_RESET_B_c_869_n N_A_1223_119#_c_1072_n 0.00254634f $X=7.66 $Y=1.165
+ $X2=0 $Y2=0
cc_705 N_RESET_B_c_871_n N_A_1223_119#_c_1072_n 0.0171699f $X=7.735 $Y=1.795
+ $X2=0 $Y2=0
cc_706 N_RESET_B_c_881_n N_A_1223_119#_c_1072_n 0.00645679f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_707 N_RESET_B_c_883_n N_A_1223_119#_c_1072_n 0.0108792f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_708 N_RESET_B_c_884_n N_A_1223_119#_c_1072_n 0.00336108f $X=8.065 $Y=2.035
+ $X2=0 $Y2=0
cc_709 N_RESET_B_c_888_n N_A_1223_119#_c_1072_n 0.00671537f $X=7.735 $Y=2.002
+ $X2=0 $Y2=0
cc_710 N_RESET_B_c_889_n N_A_1223_119#_c_1072_n 0.0174718f $X=7.825 $Y=1.96
+ $X2=0 $Y2=0
cc_711 N_RESET_B_c_876_n N_A_1223_119#_c_1078_n 6.31808e-19 $X=7.525 $Y=2.21
+ $X2=0 $Y2=0
cc_712 N_RESET_B_c_881_n N_A_1223_119#_c_1078_n 0.00286392f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_713 N_RESET_B_c_881_n N_A_1223_119#_c_1073_n 0.0252869f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_714 N_RESET_B_c_881_n N_A_852_119#_M1032_s 0.00215597f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_715 N_RESET_B_c_866_n N_A_852_119#_c_1176_n 0.0101478f $X=7.245 $Y=0.18 $X2=0
+ $Y2=0
cc_716 N_RESET_B_c_881_n N_A_852_119#_M1035_g 0.00360778f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_717 N_RESET_B_c_881_n N_A_852_119#_c_1189_n 9.73062e-19 $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_718 N_RESET_B_c_866_n N_A_852_119#_c_1180_n 0.00880557f $X=7.245 $Y=0.18
+ $X2=0 $Y2=0
cc_719 N_RESET_B_c_881_n N_A_852_119#_c_1194_n 0.00256252f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_720 N_RESET_B_c_876_n N_A_852_119#_c_1195_n 0.00850098f $X=7.525 $Y=2.21
+ $X2=0 $Y2=0
cc_721 N_RESET_B_c_883_n N_A_852_119#_M1004_g 0.00873993f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_722 N_RESET_B_c_883_n N_A_852_119#_c_1181_n 0.00840564f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_723 N_RESET_B_c_883_n N_A_852_119#_c_1182_n 3.03408e-19 $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_724 N_RESET_B_M1000_g N_A_852_119#_c_1185_n 0.00467265f $X=3.57 $Y=0.605
+ $X2=0 $Y2=0
cc_725 N_RESET_B_c_866_n N_A_852_119#_c_1185_n 0.00566977f $X=7.245 $Y=0.18
+ $X2=0 $Y2=0
cc_726 N_RESET_B_c_881_n N_A_852_119#_c_1186_n 0.0464929f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_727 N_RESET_B_c_882_n N_A_852_119#_c_1186_n 0.00281985f $X=4.225 $Y=2.035
+ $X2=0 $Y2=0
cc_728 N_RESET_B_c_886_n N_A_852_119#_c_1186_n 0.00315294f $X=3.605 $Y=2.032
+ $X2=0 $Y2=0
cc_729 N_RESET_B_c_887_n N_A_852_119#_c_1186_n 0.0250832f $X=3.95 $Y=1.985 $X2=0
+ $Y2=0
cc_730 N_RESET_B_M1020_g N_A_2006_373#_M1041_g 0.0455699f $X=10.715 $Y=0.58
+ $X2=0 $Y2=0
cc_731 N_RESET_B_c_878_n N_A_2006_373#_M1041_g 0.00569933f $X=10.855 $Y=1.82
+ $X2=0 $Y2=0
cc_732 N_RESET_B_c_878_n N_A_2006_373#_c_1355_n 0.00379957f $X=10.855 $Y=1.82
+ $X2=0 $Y2=0
cc_733 N_RESET_B_c_879_n N_A_2006_373#_c_1355_n 0.00369134f $X=11.005 $Y=2.28
+ $X2=0 $Y2=0
cc_734 N_RESET_B_c_883_n N_A_2006_373#_c_1355_n 0.0257703f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_735 RESET_B N_A_2006_373#_c_1355_n 0.00275621f $X=10.715 $Y=1.95 $X2=0 $Y2=0
cc_736 N_RESET_B_c_890_n N_A_2006_373#_c_1355_n 0.0241058f $X=10.8 $Y=2.035
+ $X2=0 $Y2=0
cc_737 N_RESET_B_c_878_n N_A_2006_373#_c_1347_n 0.00306368f $X=10.855 $Y=1.82
+ $X2=0 $Y2=0
cc_738 N_RESET_B_c_879_n N_A_2006_373#_c_1347_n 0.0031248f $X=11.005 $Y=2.28
+ $X2=0 $Y2=0
cc_739 N_RESET_B_c_873_n N_A_2006_373#_c_1347_n 0.012737f $X=10.855 $Y=1.55
+ $X2=0 $Y2=0
cc_740 N_RESET_B_c_883_n N_A_2006_373#_c_1347_n 0.00282721f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_741 RESET_B N_A_2006_373#_c_1347_n 0.00310808f $X=10.715 $Y=1.95 $X2=0 $Y2=0
cc_742 N_RESET_B_c_890_n N_A_2006_373#_c_1347_n 0.0505438f $X=10.8 $Y=2.035
+ $X2=0 $Y2=0
cc_743 N_RESET_B_c_879_n N_A_2006_373#_c_1357_n 0.0144067f $X=11.005 $Y=2.28
+ $X2=0 $Y2=0
cc_744 N_RESET_B_c_873_n N_A_2006_373#_c_1357_n 4.02079e-19 $X=10.855 $Y=1.55
+ $X2=0 $Y2=0
cc_745 N_RESET_B_c_883_n N_A_2006_373#_c_1357_n 0.00318931f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_746 RESET_B N_A_2006_373#_c_1357_n 0.0077273f $X=10.715 $Y=1.95 $X2=0 $Y2=0
cc_747 N_RESET_B_c_890_n N_A_2006_373#_c_1357_n 0.0232665f $X=10.8 $Y=2.035
+ $X2=0 $Y2=0
cc_748 N_RESET_B_M1020_g N_A_2006_373#_c_1349_n 9.65407e-19 $X=10.715 $Y=0.58
+ $X2=0 $Y2=0
cc_749 N_RESET_B_M1020_g N_A_2006_373#_c_1351_n 6.07222e-19 $X=10.715 $Y=0.58
+ $X2=0 $Y2=0
cc_750 N_RESET_B_c_879_n N_A_2006_373#_c_1359_n 0.0117118f $X=11.005 $Y=2.28
+ $X2=0 $Y2=0
cc_751 N_RESET_B_c_890_n N_A_2006_373#_c_1359_n 0.0277898f $X=10.8 $Y=2.035
+ $X2=0 $Y2=0
cc_752 N_RESET_B_c_879_n N_A_2006_373#_c_1360_n 0.0215739f $X=11.005 $Y=2.28
+ $X2=0 $Y2=0
cc_753 N_RESET_B_c_883_n N_A_2006_373#_c_1360_n 0.0142613f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_754 RESET_B N_A_2006_373#_c_1360_n 0.00149024f $X=10.715 $Y=1.95 $X2=0 $Y2=0
cc_755 N_RESET_B_c_890_n N_A_2006_373#_c_1360_n 0.00155699f $X=10.8 $Y=2.035
+ $X2=0 $Y2=0
cc_756 N_RESET_B_c_883_n N_A_1790_75#_M1004_d 0.00975786f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_757 N_RESET_B_M1020_g N_A_1790_75#_M1013_g 0.0556926f $X=10.715 $Y=0.58 $X2=0
+ $Y2=0
cc_758 N_RESET_B_M1020_g N_A_1790_75#_c_1457_n 0.0094439f $X=10.715 $Y=0.58
+ $X2=0 $Y2=0
cc_759 N_RESET_B_c_879_n N_A_1790_75#_c_1457_n 0.00125789f $X=11.005 $Y=2.28
+ $X2=0 $Y2=0
cc_760 N_RESET_B_c_873_n N_A_1790_75#_c_1457_n 0.00511143f $X=10.855 $Y=1.55
+ $X2=0 $Y2=0
cc_761 N_RESET_B_c_878_n N_A_1790_75#_c_1467_n 0.00511143f $X=10.855 $Y=1.82
+ $X2=0 $Y2=0
cc_762 N_RESET_B_c_879_n N_A_1790_75#_c_1467_n 0.0232392f $X=11.005 $Y=2.28
+ $X2=0 $Y2=0
cc_763 N_RESET_B_c_890_n N_A_1790_75#_c_1467_n 0.0083262f $X=10.8 $Y=2.035 $X2=0
+ $Y2=0
cc_764 N_RESET_B_c_879_n N_A_1790_75#_c_1468_n 0.00947913f $X=11.005 $Y=2.28
+ $X2=0 $Y2=0
cc_765 N_RESET_B_c_883_n N_A_1790_75#_c_1478_n 0.0195683f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_766 N_RESET_B_c_883_n N_A_1790_75#_c_1465_n 0.0213448f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_767 N_RESET_B_M1020_g N_A_1790_75#_c_1466_n 0.0184362f $X=10.715 $Y=0.58
+ $X2=0 $Y2=0
cc_768 N_RESET_B_c_873_n N_A_1790_75#_c_1466_n 0.00370089f $X=10.855 $Y=1.55
+ $X2=0 $Y2=0
cc_769 N_RESET_B_c_881_n N_VPWR_M1032_d 0.00305774f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_770 N_RESET_B_c_883_n N_VPWR_M1039_s 0.00198285f $X=10.655 $Y=2.035 $X2=0
+ $Y2=0
cc_771 N_RESET_B_c_875_n N_VPWR_c_1659_n 0.00579128f $X=3.605 $Y=2.245 $X2=0
+ $Y2=0
cc_772 N_RESET_B_c_876_n N_VPWR_c_1661_n 0.00314968f $X=7.525 $Y=2.21 $X2=0
+ $Y2=0
cc_773 N_RESET_B_c_876_n N_VPWR_c_1662_n 0.00490213f $X=7.525 $Y=2.21 $X2=0
+ $Y2=0
cc_774 N_RESET_B_c_871_n N_VPWR_c_1662_n 4.78591e-19 $X=7.735 $Y=1.795 $X2=0
+ $Y2=0
cc_775 N_RESET_B_c_883_n N_VPWR_c_1662_n 0.0236795f $X=10.655 $Y=2.035 $X2=0
+ $Y2=0
cc_776 N_RESET_B_c_884_n N_VPWR_c_1662_n 0.0027362f $X=8.065 $Y=2.035 $X2=0
+ $Y2=0
cc_777 N_RESET_B_c_888_n N_VPWR_c_1662_n 0.0020516f $X=7.735 $Y=2.002 $X2=0
+ $Y2=0
cc_778 N_RESET_B_c_889_n N_VPWR_c_1662_n 0.0258087f $X=7.825 $Y=1.96 $X2=0 $Y2=0
cc_779 N_RESET_B_c_890_n N_VPWR_c_1664_n 0.0233946f $X=10.8 $Y=2.035 $X2=0 $Y2=0
cc_780 N_RESET_B_c_875_n N_VPWR_c_1669_n 0.00388952f $X=3.605 $Y=2.245 $X2=0
+ $Y2=0
cc_781 N_RESET_B_c_879_n N_VPWR_c_1675_n 0.00443738f $X=11.005 $Y=2.28 $X2=0
+ $Y2=0
cc_782 N_RESET_B_c_879_n N_VPWR_c_1683_n 0.00802674f $X=11.005 $Y=2.28 $X2=0
+ $Y2=0
cc_783 N_RESET_B_c_883_n N_VPWR_c_1683_n 0.00135379f $X=10.655 $Y=2.035 $X2=0
+ $Y2=0
cc_784 N_RESET_B_c_875_n N_VPWR_c_1658_n 0.00423691f $X=3.605 $Y=2.245 $X2=0
+ $Y2=0
cc_785 N_RESET_B_c_876_n N_VPWR_c_1658_n 9.49986e-19 $X=7.525 $Y=2.21 $X2=0
+ $Y2=0
cc_786 N_RESET_B_c_879_n N_VPWR_c_1658_n 0.00489211f $X=11.005 $Y=2.28 $X2=0
+ $Y2=0
cc_787 N_RESET_B_M1000_g N_A_388_79#_c_1848_n 0.0179961f $X=3.57 $Y=0.605 $X2=0
+ $Y2=0
cc_788 N_RESET_B_M1000_g N_A_388_79#_c_1850_n 0.022108f $X=3.57 $Y=0.605 $X2=0
+ $Y2=0
cc_789 N_RESET_B_c_875_n N_A_388_79#_c_1850_n 0.00392187f $X=3.605 $Y=2.245
+ $X2=0 $Y2=0
cc_790 N_RESET_B_c_882_n N_A_388_79#_c_1850_n 0.00108246f $X=4.225 $Y=2.035
+ $X2=0 $Y2=0
cc_791 N_RESET_B_c_886_n N_A_388_79#_c_1850_n 0.0151779f $X=3.605 $Y=2.032 $X2=0
+ $Y2=0
cc_792 N_RESET_B_c_887_n N_A_388_79#_c_1850_n 0.0228178f $X=3.95 $Y=1.985 $X2=0
+ $Y2=0
cc_793 N_RESET_B_c_875_n N_A_388_79#_c_1858_n 0.0248771f $X=3.605 $Y=2.245 $X2=0
+ $Y2=0
cc_794 N_RESET_B_c_882_n N_A_388_79#_c_1858_n 0.001474f $X=4.225 $Y=2.035 $X2=0
+ $Y2=0
cc_795 N_RESET_B_c_886_n N_A_388_79#_c_1858_n 0.00751654f $X=3.605 $Y=2.032
+ $X2=0 $Y2=0
cc_796 N_RESET_B_c_887_n N_A_388_79#_c_1858_n 0.0165337f $X=3.95 $Y=1.985 $X2=0
+ $Y2=0
cc_797 N_RESET_B_c_881_n N_A_388_79#_c_1859_n 0.00436641f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_798 N_RESET_B_c_881_n N_A_388_79#_c_1860_n 0.0125677f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_799 N_RESET_B_c_881_n N_A_388_79#_c_1854_n 0.0149539f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_800 N_RESET_B_c_881_n N_A_388_79#_c_1862_n 0.00680456f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_801 N_RESET_B_c_882_n N_A_388_79#_c_1862_n 0.00654599f $X=4.225 $Y=2.035
+ $X2=0 $Y2=0
cc_802 N_RESET_B_c_886_n N_A_388_79#_c_1862_n 0.00181987f $X=3.605 $Y=2.032
+ $X2=0 $Y2=0
cc_803 N_RESET_B_c_887_n N_A_388_79#_c_1862_n 0.00668852f $X=3.95 $Y=1.985 $X2=0
+ $Y2=0
cc_804 N_RESET_B_c_881_n N_A_388_79#_c_1902_n 0.0134265f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_805 N_RESET_B_c_881_n N_A_388_79#_c_1863_n 0.00782023f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_806 N_RESET_B_M1000_g N_VGND_c_2053_n 0.00775196f $X=3.57 $Y=0.605 $X2=0
+ $Y2=0
cc_807 N_RESET_B_c_866_n N_VGND_c_2053_n 0.0196811f $X=7.245 $Y=0.18 $X2=0 $Y2=0
cc_808 N_RESET_B_c_867_n N_VGND_c_2053_n 0.00321798f $X=3.645 $Y=0.18 $X2=0
+ $Y2=0
cc_809 N_RESET_B_c_866_n N_VGND_c_2054_n 0.0170937f $X=7.245 $Y=0.18 $X2=0 $Y2=0
cc_810 N_RESET_B_M1020_g N_VGND_c_2055_n 0.0122664f $X=10.715 $Y=0.58 $X2=0
+ $Y2=0
cc_811 N_RESET_B_c_867_n N_VGND_c_2062_n 0.00564095f $X=3.645 $Y=0.18 $X2=0
+ $Y2=0
cc_812 N_RESET_B_c_866_n N_VGND_c_2064_n 0.0237832f $X=7.245 $Y=0.18 $X2=0 $Y2=0
cc_813 N_RESET_B_M1020_g N_VGND_c_2069_n 0.00383152f $X=10.715 $Y=0.58 $X2=0
+ $Y2=0
cc_814 N_RESET_B_c_866_n N_VGND_c_2073_n 0.0558684f $X=7.245 $Y=0.18 $X2=0 $Y2=0
cc_815 N_RESET_B_c_866_n N_VGND_c_2074_n 0.0109384f $X=7.245 $Y=0.18 $X2=0 $Y2=0
cc_816 N_RESET_B_c_866_n N_VGND_c_2078_n 0.0937386f $X=7.245 $Y=0.18 $X2=0 $Y2=0
cc_817 N_RESET_B_c_867_n N_VGND_c_2078_n 0.0110707f $X=3.645 $Y=0.18 $X2=0 $Y2=0
cc_818 N_RESET_B_M1020_g N_VGND_c_2078_n 0.0075694f $X=10.715 $Y=0.58 $X2=0
+ $Y2=0
cc_819 N_RESET_B_M1000_g N_noxref_25_c_2208_n 0.00204561f $X=3.57 $Y=0.605 $X2=0
+ $Y2=0
cc_820 N_RESET_B_M1000_g N_noxref_25_c_2210_n 0.0037218f $X=3.57 $Y=0.605 $X2=0
+ $Y2=0
cc_821 N_A_1223_119#_c_1075_n N_A_852_119#_c_1190_n 0.0036476f $X=6.66 $Y=2.61
+ $X2=0 $Y2=0
cc_822 N_A_1223_119#_c_1075_n N_A_852_119#_c_1192_n 9.70565e-19 $X=6.66 $Y=2.61
+ $X2=0 $Y2=0
cc_823 N_A_1223_119#_c_1075_n N_A_852_119#_c_1194_n 0.0101282f $X=6.66 $Y=2.61
+ $X2=0 $Y2=0
cc_824 N_A_1223_119#_c_1078_n N_A_852_119#_c_1194_n 4.9181e-19 $X=6.78 $Y=2.425
+ $X2=0 $Y2=0
cc_825 N_A_1223_119#_c_1073_n N_A_852_119#_c_1194_n 0.00166513f $X=6.78 $Y=2.34
+ $X2=0 $Y2=0
cc_826 N_A_1223_119#_c_1069_n N_A_852_119#_c_1195_n 0.0103562f $X=8.5 $Y=1.66
+ $X2=0 $Y2=0
cc_827 N_A_1223_119#_c_1095_n N_A_852_119#_c_1195_n 0.00255374f $X=7.38 $Y=2.425
+ $X2=0 $Y2=0
cc_828 N_A_1223_119#_c_1070_n N_A_852_119#_c_1195_n 0.00749106f $X=7.465 $Y=2.32
+ $X2=0 $Y2=0
cc_829 N_A_1223_119#_c_1078_n N_A_852_119#_c_1195_n 0.00275309f $X=6.78 $Y=2.425
+ $X2=0 $Y2=0
cc_830 N_A_1223_119#_c_1069_n N_A_852_119#_c_1196_n 0.00249951f $X=8.5 $Y=1.66
+ $X2=0 $Y2=0
cc_831 N_A_1223_119#_c_1069_n N_A_852_119#_M1004_g 0.00579836f $X=8.5 $Y=1.66
+ $X2=0 $Y2=0
cc_832 N_A_1223_119#_c_1069_n N_A_852_119#_c_1182_n 0.00845345f $X=8.5 $Y=1.66
+ $X2=0 $Y2=0
cc_833 N_A_1223_119#_c_1095_n N_VPWR_M1042_d 0.00730901f $X=7.38 $Y=2.425 $X2=0
+ $Y2=0
cc_834 N_A_1223_119#_c_1070_n N_VPWR_M1042_d 8.72177e-19 $X=7.465 $Y=2.32 $X2=0
+ $Y2=0
cc_835 N_A_1223_119#_c_1095_n N_VPWR_c_1661_n 0.0190336f $X=7.38 $Y=2.425 $X2=0
+ $Y2=0
cc_836 N_A_1223_119#_c_1070_n N_VPWR_c_1661_n 0.00274183f $X=7.465 $Y=2.32 $X2=0
+ $Y2=0
cc_837 N_A_1223_119#_c_1078_n N_VPWR_c_1661_n 0.00236604f $X=6.78 $Y=2.425 $X2=0
+ $Y2=0
cc_838 N_A_1223_119#_c_1069_n N_VPWR_c_1662_n 0.0179689f $X=8.5 $Y=1.66 $X2=0
+ $Y2=0
cc_839 N_A_1223_119#_c_1070_n N_VPWR_c_1662_n 0.0295999f $X=7.465 $Y=2.32 $X2=0
+ $Y2=0
cc_840 N_A_1223_119#_c_1072_n N_VPWR_c_1662_n 0.0170777f $X=8.425 $Y=1.41 $X2=0
+ $Y2=0
cc_841 N_A_1223_119#_c_1075_n N_VPWR_c_1671_n 0.009596f $X=6.66 $Y=2.61 $X2=0
+ $Y2=0
cc_842 N_A_1223_119#_c_1078_n N_VPWR_c_1671_n 0.00499509f $X=6.78 $Y=2.425 $X2=0
+ $Y2=0
cc_843 N_A_1223_119#_c_1070_n N_VPWR_c_1674_n 0.00745648f $X=7.465 $Y=2.32 $X2=0
+ $Y2=0
cc_844 N_A_1223_119#_c_1069_n N_VPWR_c_1658_n 8.51577e-19 $X=8.5 $Y=1.66 $X2=0
+ $Y2=0
cc_845 N_A_1223_119#_c_1075_n N_VPWR_c_1658_n 0.012602f $X=6.66 $Y=2.61 $X2=0
+ $Y2=0
cc_846 N_A_1223_119#_c_1095_n N_VPWR_c_1658_n 0.00768901f $X=7.38 $Y=2.425 $X2=0
+ $Y2=0
cc_847 N_A_1223_119#_c_1070_n N_VPWR_c_1658_n 0.0153115f $X=7.465 $Y=2.32 $X2=0
+ $Y2=0
cc_848 N_A_1223_119#_c_1078_n N_VPWR_c_1658_n 0.00635167f $X=6.78 $Y=2.425 $X2=0
+ $Y2=0
cc_849 N_A_1223_119#_c_1073_n N_A_388_79#_c_1851_n 0.00327725f $X=6.78 $Y=2.34
+ $X2=0 $Y2=0
cc_850 N_A_1223_119#_M1033_d N_A_388_79#_c_1860_n 0.00201424f $X=6.175 $Y=2.285
+ $X2=0 $Y2=0
cc_851 N_A_1223_119#_c_1075_n N_A_388_79#_c_1860_n 0.0159467f $X=6.66 $Y=2.61
+ $X2=0 $Y2=0
cc_852 N_A_1223_119#_c_1073_n N_A_388_79#_c_1860_n 0.0120507f $X=6.78 $Y=2.34
+ $X2=0 $Y2=0
cc_853 N_A_1223_119#_c_1082_n N_A_388_79#_c_1852_n 0.0240423f $X=6.66 $Y=0.8
+ $X2=0 $Y2=0
cc_854 N_A_1223_119#_c_1073_n N_A_388_79#_c_1852_n 0.0135678f $X=6.78 $Y=2.34
+ $X2=0 $Y2=0
cc_855 N_A_1223_119#_c_1073_n N_A_388_79#_c_1854_n 0.0629989f $X=6.78 $Y=2.34
+ $X2=0 $Y2=0
cc_856 N_A_1223_119#_c_1075_n N_A_388_79#_c_1863_n 0.00971511f $X=6.66 $Y=2.61
+ $X2=0 $Y2=0
cc_857 N_A_1223_119#_M1002_g N_VGND_c_2066_n 0.00278271f $X=8.445 $Y=0.695 $X2=0
+ $Y2=0
cc_858 N_A_1223_119#_M1002_g N_VGND_c_2074_n 0.00116012f $X=8.445 $Y=0.695 $X2=0
+ $Y2=0
cc_859 N_A_1223_119#_M1002_g N_VGND_c_2078_n 0.00358525f $X=8.445 $Y=0.695 $X2=0
+ $Y2=0
cc_860 N_A_1223_119#_c_1082_n A_1323_119# 0.0012023f $X=6.66 $Y=0.8 $X2=-0.19
+ $Y2=-0.245
cc_861 N_A_852_119#_M1045_g N_A_2006_373#_M1041_g 0.0830829f $X=9.925 $Y=0.58
+ $X2=0 $Y2=0
cc_862 N_A_852_119#_M1004_g N_A_1790_75#_c_1478_n 0.00371138f $X=8.95 $Y=2.235
+ $X2=0 $Y2=0
cc_863 N_A_852_119#_M1045_g N_A_1790_75#_c_1480_n 0.0113037f $X=9.925 $Y=0.58
+ $X2=0 $Y2=0
cc_864 N_A_852_119#_M1045_g N_A_1790_75#_c_1464_n 0.00782202f $X=9.925 $Y=0.58
+ $X2=0 $Y2=0
cc_865 N_A_852_119#_c_1181_n N_A_1790_75#_c_1465_n 0.00624492f $X=9.85 $Y=1.55
+ $X2=0 $Y2=0
cc_866 N_A_852_119#_M1045_g N_A_1790_75#_c_1465_n 0.0034675f $X=9.925 $Y=0.58
+ $X2=0 $Y2=0
cc_867 N_A_852_119#_M1045_g N_A_1790_75#_c_1490_n 0.00668381f $X=9.925 $Y=0.58
+ $X2=0 $Y2=0
cc_868 N_A_852_119#_c_1186_n N_VPWR_M1032_d 0.00199165f $X=4.49 $Y=1.847 $X2=0
+ $Y2=0
cc_869 N_A_852_119#_M1035_g N_VPWR_c_1660_n 0.00840339f $X=5.095 $Y=2.46 $X2=0
+ $Y2=0
cc_870 N_A_852_119#_c_1189_n N_VPWR_c_1660_n 0.00168763f $X=5.595 $Y=3.075 $X2=0
+ $Y2=0
cc_871 N_A_852_119#_c_1191_n N_VPWR_c_1660_n 0.00241263f $X=5.67 $Y=3.15 $X2=0
+ $Y2=0
cc_872 N_A_852_119#_c_1192_n N_VPWR_c_1661_n 0.00673937f $X=6.55 $Y=2.87 $X2=0
+ $Y2=0
cc_873 N_A_852_119#_c_1195_n N_VPWR_c_1661_n 0.0209699f $X=8.86 $Y=3.15 $X2=0
+ $Y2=0
cc_874 N_A_852_119#_c_1195_n N_VPWR_c_1662_n 0.0213056f $X=8.86 $Y=3.15 $X2=0
+ $Y2=0
cc_875 N_A_852_119#_c_1196_n N_VPWR_c_1662_n 0.00613773f $X=8.95 $Y=2.9 $X2=0
+ $Y2=0
cc_876 N_A_852_119#_M1004_g N_VPWR_c_1662_n 6.31058e-19 $X=8.95 $Y=2.235 $X2=0
+ $Y2=0
cc_877 N_A_852_119#_c_1195_n N_VPWR_c_1663_n 0.0188492f $X=8.86 $Y=3.15 $X2=0
+ $Y2=0
cc_878 N_A_852_119#_M1035_g N_VPWR_c_1671_n 0.00303678f $X=5.095 $Y=2.46 $X2=0
+ $Y2=0
cc_879 N_A_852_119#_c_1191_n N_VPWR_c_1671_n 0.0438713f $X=5.67 $Y=3.15 $X2=0
+ $Y2=0
cc_880 N_A_852_119#_c_1195_n N_VPWR_c_1674_n 0.0266609f $X=8.86 $Y=3.15 $X2=0
+ $Y2=0
cc_881 N_A_852_119#_M1035_g N_VPWR_c_1658_n 0.00394565f $X=5.095 $Y=2.46 $X2=0
+ $Y2=0
cc_882 N_A_852_119#_c_1190_n N_VPWR_c_1658_n 0.0231728f $X=6.46 $Y=3.15 $X2=0
+ $Y2=0
cc_883 N_A_852_119#_c_1191_n N_VPWR_c_1658_n 0.00688548f $X=5.67 $Y=3.15 $X2=0
+ $Y2=0
cc_884 N_A_852_119#_c_1195_n N_VPWR_c_1658_n 0.0670958f $X=8.86 $Y=3.15 $X2=0
+ $Y2=0
cc_885 N_A_852_119#_c_1201_n N_VPWR_c_1658_n 0.00504011f $X=6.55 $Y=3.15 $X2=0
+ $Y2=0
cc_886 N_A_852_119#_M1035_g N_A_388_79#_c_1859_n 0.0141206f $X=5.095 $Y=2.46
+ $X2=0 $Y2=0
cc_887 N_A_852_119#_c_1189_n N_A_388_79#_c_1859_n 0.013013f $X=5.595 $Y=3.075
+ $X2=0 $Y2=0
cc_888 N_A_852_119#_c_1186_n N_A_388_79#_c_1859_n 0.0014292f $X=4.49 $Y=1.847
+ $X2=0 $Y2=0
cc_889 N_A_852_119#_c_1176_n N_A_388_79#_c_1851_n 5.04404e-19 $X=5.05 $Y=1.445
+ $X2=0 $Y2=0
cc_890 N_A_852_119#_c_1178_n N_A_388_79#_c_1851_n 0.00417422f $X=5.965 $Y=1.165
+ $X2=0 $Y2=0
cc_891 N_A_852_119#_c_1180_n N_A_388_79#_c_1851_n 0.00690249f $X=6.04 $Y=1.09
+ $X2=0 $Y2=0
cc_892 N_A_852_119#_c_1194_n N_A_388_79#_c_1860_n 0.00417216f $X=6.55 $Y=2.78
+ $X2=0 $Y2=0
cc_893 N_A_852_119#_c_1178_n N_A_388_79#_c_1852_n 0.00708724f $X=5.965 $Y=1.165
+ $X2=0 $Y2=0
cc_894 N_A_852_119#_c_1178_n N_A_388_79#_c_1853_n 0.00497709f $X=5.965 $Y=1.165
+ $X2=0 $Y2=0
cc_895 N_A_852_119#_c_1177_n N_A_388_79#_c_1854_n 0.00257235f $X=5.58 $Y=1.445
+ $X2=0 $Y2=0
cc_896 N_A_852_119#_M1032_s N_A_388_79#_c_1862_n 0.00821428f $X=4.275 $Y=1.96
+ $X2=0 $Y2=0
cc_897 N_A_852_119#_c_1186_n N_A_388_79#_c_1862_n 0.0134136f $X=4.49 $Y=1.847
+ $X2=0 $Y2=0
cc_898 N_A_852_119#_c_1186_n N_A_388_79#_c_1902_n 0.00787817f $X=4.49 $Y=1.847
+ $X2=0 $Y2=0
cc_899 N_A_852_119#_c_1178_n N_A_388_79#_c_1855_n 5.32864e-19 $X=5.965 $Y=1.165
+ $X2=0 $Y2=0
cc_900 N_A_852_119#_c_1179_n N_A_388_79#_c_1855_n 0.00500227f $X=5.67 $Y=1.165
+ $X2=0 $Y2=0
cc_901 N_A_852_119#_c_1180_n N_A_388_79#_c_1855_n 0.00209515f $X=6.04 $Y=1.09
+ $X2=0 $Y2=0
cc_902 N_A_852_119#_c_1189_n N_A_388_79#_c_1863_n 0.00912689f $X=5.595 $Y=3.075
+ $X2=0 $Y2=0
cc_903 N_A_852_119#_c_1190_n N_A_388_79#_c_1863_n 0.0043692f $X=6.46 $Y=3.15
+ $X2=0 $Y2=0
cc_904 N_A_852_119#_c_1185_n N_VGND_c_2053_n 0.0144881f $X=4.49 $Y=0.802 $X2=0
+ $Y2=0
cc_905 N_A_852_119#_c_1176_n N_VGND_c_2054_n 0.00166106f $X=5.05 $Y=1.445 $X2=0
+ $Y2=0
cc_906 N_A_852_119#_c_1186_n N_VGND_c_2054_n 0.00961843f $X=4.49 $Y=1.847 $X2=0
+ $Y2=0
cc_907 N_A_852_119#_M1045_g N_VGND_c_2055_n 0.00120934f $X=9.925 $Y=0.58 $X2=0
+ $Y2=0
cc_908 N_A_852_119#_c_1185_n N_VGND_c_2064_n 0.00623819f $X=4.49 $Y=0.802 $X2=0
+ $Y2=0
cc_909 N_A_852_119#_M1045_g N_VGND_c_2066_n 0.00298877f $X=9.925 $Y=0.58 $X2=0
+ $Y2=0
cc_910 N_A_852_119#_c_1176_n N_VGND_c_2078_n 7.82699e-19 $X=5.05 $Y=1.445 $X2=0
+ $Y2=0
cc_911 N_A_852_119#_M1045_g N_VGND_c_2078_n 0.00370514f $X=9.925 $Y=0.58 $X2=0
+ $Y2=0
cc_912 N_A_852_119#_c_1185_n N_VGND_c_2078_n 0.00887442f $X=4.49 $Y=0.802 $X2=0
+ $Y2=0
cc_913 N_A_2006_373#_c_1349_n N_A_1790_75#_M1013_g 0.00658176f $X=11.29 $Y=0.58
+ $X2=0 $Y2=0
cc_914 N_A_2006_373#_c_1351_n N_A_1790_75#_M1013_g 0.00562994f $X=11.455 $Y=0.79
+ $X2=0 $Y2=0
cc_915 N_A_2006_373#_c_1352_n N_A_1790_75#_M1013_g 0.00311727f $X=11.775 $Y=1.48
+ $X2=0 $Y2=0
cc_916 N_A_2006_373#_c_1347_n N_A_1790_75#_c_1457_n 0.0111503f $X=11.69 $Y=1.565
+ $X2=0 $Y2=0
cc_917 N_A_2006_373#_c_1350_n N_A_1790_75#_c_1457_n 0.00258531f $X=11.69 $Y=0.79
+ $X2=0 $Y2=0
cc_918 N_A_2006_373#_c_1351_n N_A_1790_75#_c_1457_n 0.0075729f $X=11.455 $Y=0.79
+ $X2=0 $Y2=0
cc_919 N_A_2006_373#_c_1352_n N_A_1790_75#_c_1457_n 0.00284108f $X=11.775
+ $Y=1.48 $X2=0 $Y2=0
cc_920 N_A_2006_373#_c_1347_n N_A_1790_75#_c_1467_n 0.00952908f $X=11.69
+ $Y=1.565 $X2=0 $Y2=0
cc_921 N_A_2006_373#_c_1359_n N_A_1790_75#_c_1468_n 0.00686533f $X=11.23
+ $Y=2.405 $X2=0 $Y2=0
cc_922 N_A_2006_373#_c_1347_n N_A_1790_75#_c_1458_n 0.0131208f $X=11.69 $Y=1.565
+ $X2=0 $Y2=0
cc_923 N_A_2006_373#_c_1350_n N_A_1790_75#_c_1458_n 0.00113849f $X=11.69 $Y=0.79
+ $X2=0 $Y2=0
cc_924 N_A_2006_373#_c_1352_n N_A_1790_75#_c_1458_n 0.0180935f $X=11.775 $Y=1.48
+ $X2=0 $Y2=0
cc_925 N_A_2006_373#_c_1349_n N_A_1790_75#_M1021_g 0.00446735f $X=11.29 $Y=0.58
+ $X2=0 $Y2=0
cc_926 N_A_2006_373#_c_1350_n N_A_1790_75#_M1021_g 0.00377396f $X=11.69 $Y=0.79
+ $X2=0 $Y2=0
cc_927 N_A_2006_373#_c_1352_n N_A_1790_75#_M1021_g 0.00455681f $X=11.775 $Y=1.48
+ $X2=0 $Y2=0
cc_928 N_A_2006_373#_c_1347_n N_A_1790_75#_c_1461_n 5.76097e-19 $X=11.69
+ $Y=1.565 $X2=0 $Y2=0
cc_929 N_A_2006_373#_c_1353_n N_A_1790_75#_c_1478_n 0.0150017f $X=10.12 $Y=2.28
+ $X2=0 $Y2=0
cc_930 N_A_2006_373#_c_1358_n N_A_1790_75#_c_1478_n 0.0109254f $X=10.545
+ $Y=2.405 $X2=0 $Y2=0
cc_931 N_A_2006_373#_M1041_g N_A_1790_75#_c_1480_n 0.00245703f $X=10.285 $Y=0.58
+ $X2=0 $Y2=0
cc_932 N_A_2006_373#_M1041_g N_A_1790_75#_c_1464_n 0.00544577f $X=10.285 $Y=0.58
+ $X2=0 $Y2=0
cc_933 N_A_2006_373#_c_1353_n N_A_1790_75#_c_1465_n 0.00156196f $X=10.12 $Y=2.28
+ $X2=0 $Y2=0
cc_934 N_A_2006_373#_M1041_g N_A_1790_75#_c_1465_n 0.0092441f $X=10.285 $Y=0.58
+ $X2=0 $Y2=0
cc_935 N_A_2006_373#_c_1355_n N_A_1790_75#_c_1465_n 0.0474407f $X=10.405 $Y=2.03
+ $X2=0 $Y2=0
cc_936 N_A_2006_373#_c_1348_n N_A_1790_75#_c_1465_n 0.0135848f $X=10.545
+ $Y=1.565 $X2=0 $Y2=0
cc_937 N_A_2006_373#_c_1358_n N_A_1790_75#_c_1465_n 0.00357879f $X=10.545
+ $Y=2.405 $X2=0 $Y2=0
cc_938 N_A_2006_373#_c_1360_n N_A_1790_75#_c_1465_n 0.0108982f $X=10.285
+ $Y=2.072 $X2=0 $Y2=0
cc_939 N_A_2006_373#_M1041_g N_A_1790_75#_c_1466_n 0.0192761f $X=10.285 $Y=0.58
+ $X2=0 $Y2=0
cc_940 N_A_2006_373#_c_1347_n N_A_1790_75#_c_1466_n 0.0718198f $X=11.69 $Y=1.565
+ $X2=0 $Y2=0
cc_941 N_A_2006_373#_c_1348_n N_A_1790_75#_c_1466_n 0.0235777f $X=10.545
+ $Y=1.565 $X2=0 $Y2=0
cc_942 N_A_2006_373#_c_1350_n N_A_1790_75#_c_1466_n 0.00476671f $X=11.69 $Y=0.79
+ $X2=0 $Y2=0
cc_943 N_A_2006_373#_c_1351_n N_A_1790_75#_c_1466_n 0.026725f $X=11.455 $Y=0.79
+ $X2=0 $Y2=0
cc_944 N_A_2006_373#_c_1352_n N_A_1790_75#_c_1466_n 0.0207312f $X=11.775 $Y=1.48
+ $X2=0 $Y2=0
cc_945 N_A_2006_373#_c_1360_n N_A_1790_75#_c_1466_n 0.00394383f $X=10.285
+ $Y=2.072 $X2=0 $Y2=0
cc_946 N_A_2006_373#_c_1357_n N_VPWR_M1001_d 0.00487963f $X=11.065 $Y=2.405
+ $X2=0 $Y2=0
cc_947 N_A_2006_373#_c_1358_n N_VPWR_M1001_d 0.00589954f $X=10.545 $Y=2.405
+ $X2=0 $Y2=0
cc_948 N_A_2006_373#_c_1353_n N_VPWR_c_1663_n 0.00419312f $X=10.12 $Y=2.28 $X2=0
+ $Y2=0
cc_949 N_A_2006_373#_c_1347_n N_VPWR_c_1664_n 0.0223739f $X=11.69 $Y=1.565 $X2=0
+ $Y2=0
cc_950 N_A_2006_373#_c_1359_n N_VPWR_c_1664_n 0.031333f $X=11.23 $Y=2.405 $X2=0
+ $Y2=0
cc_951 N_A_2006_373#_c_1359_n N_VPWR_c_1675_n 0.00802713f $X=11.23 $Y=2.405
+ $X2=0 $Y2=0
cc_952 N_A_2006_373#_c_1353_n N_VPWR_c_1683_n 0.0101552f $X=10.12 $Y=2.28 $X2=0
+ $Y2=0
cc_953 N_A_2006_373#_c_1357_n N_VPWR_c_1683_n 0.0240529f $X=11.065 $Y=2.405
+ $X2=0 $Y2=0
cc_954 N_A_2006_373#_c_1358_n N_VPWR_c_1683_n 0.0238431f $X=10.545 $Y=2.405
+ $X2=0 $Y2=0
cc_955 N_A_2006_373#_c_1359_n N_VPWR_c_1683_n 0.0095412f $X=11.23 $Y=2.405 $X2=0
+ $Y2=0
cc_956 N_A_2006_373#_c_1360_n N_VPWR_c_1683_n 0.00121809f $X=10.285 $Y=2.072
+ $X2=0 $Y2=0
cc_957 N_A_2006_373#_c_1353_n N_VPWR_c_1658_n 0.00489211f $X=10.12 $Y=2.28 $X2=0
+ $Y2=0
cc_958 N_A_2006_373#_c_1357_n N_VPWR_c_1658_n 0.00766785f $X=11.065 $Y=2.405
+ $X2=0 $Y2=0
cc_959 N_A_2006_373#_c_1358_n N_VPWR_c_1658_n 0.00101543f $X=10.545 $Y=2.405
+ $X2=0 $Y2=0
cc_960 N_A_2006_373#_c_1359_n N_VPWR_c_1658_n 0.010512f $X=11.23 $Y=2.405 $X2=0
+ $Y2=0
cc_961 N_A_2006_373#_c_1347_n Q_N 0.0138399f $X=11.69 $Y=1.565 $X2=0 $Y2=0
cc_962 N_A_2006_373#_c_1350_n N_Q_N_c_2009_n 0.00970057f $X=11.69 $Y=0.79 $X2=0
+ $Y2=0
cc_963 N_A_2006_373#_c_1352_n N_Q_N_c_2009_n 0.00199024f $X=11.775 $Y=1.48 $X2=0
+ $Y2=0
cc_964 N_A_2006_373#_c_1352_n Q_N 0.0415299f $X=11.775 $Y=1.48 $X2=0 $Y2=0
cc_965 N_A_2006_373#_c_1350_n N_VGND_M1021_s 0.00517852f $X=11.69 $Y=0.79 $X2=0
+ $Y2=0
cc_966 N_A_2006_373#_c_1352_n N_VGND_M1021_s 0.00675628f $X=11.775 $Y=1.48 $X2=0
+ $Y2=0
cc_967 N_A_2006_373#_M1041_g N_VGND_c_2055_n 0.0105628f $X=10.285 $Y=0.58 $X2=0
+ $Y2=0
cc_968 N_A_2006_373#_c_1349_n N_VGND_c_2055_n 0.0118606f $X=11.29 $Y=0.58 $X2=0
+ $Y2=0
cc_969 N_A_2006_373#_c_1351_n N_VGND_c_2055_n 0.00372607f $X=11.455 $Y=0.79
+ $X2=0 $Y2=0
cc_970 N_A_2006_373#_c_1349_n N_VGND_c_2056_n 0.0139523f $X=11.29 $Y=0.58 $X2=0
+ $Y2=0
cc_971 N_A_2006_373#_c_1350_n N_VGND_c_2056_n 0.0181192f $X=11.69 $Y=0.79 $X2=0
+ $Y2=0
cc_972 N_A_2006_373#_M1041_g N_VGND_c_2066_n 0.00383152f $X=10.285 $Y=0.58 $X2=0
+ $Y2=0
cc_973 N_A_2006_373#_c_1349_n N_VGND_c_2069_n 0.0142949f $X=11.29 $Y=0.58 $X2=0
+ $Y2=0
cc_974 N_A_2006_373#_c_1350_n N_VGND_c_2069_n 0.00298753f $X=11.69 $Y=0.79 $X2=0
+ $Y2=0
cc_975 N_A_2006_373#_M1041_g N_VGND_c_2078_n 0.0075694f $X=10.285 $Y=0.58 $X2=0
+ $Y2=0
cc_976 N_A_2006_373#_c_1349_n N_VGND_c_2078_n 0.011894f $X=11.29 $Y=0.58 $X2=0
+ $Y2=0
cc_977 N_A_2006_373#_c_1350_n N_VGND_c_2078_n 0.00611276f $X=11.69 $Y=0.79 $X2=0
+ $Y2=0
cc_978 N_A_1790_75#_c_1461_n N_A_2604_392#_c_1609_n 0.0166552f $X=12.945
+ $Y=1.585 $X2=0 $Y2=0
cc_979 N_A_1790_75#_c_1462_n N_A_2604_392#_c_1609_n 0.00200517f $X=12.945
+ $Y=1.795 $X2=0 $Y2=0
cc_980 N_A_1790_75#_M1005_g N_A_2604_392#_c_1611_n 0.0121223f $X=12.99 $Y=0.69
+ $X2=0 $Y2=0
cc_981 N_A_1790_75#_c_1462_n N_A_2604_392#_c_1612_n 0.0108738f $X=12.945
+ $Y=1.795 $X2=0 $Y2=0
cc_982 N_A_1790_75#_c_1473_n N_A_2604_392#_c_1612_n 0.00283082f $X=12.945
+ $Y=1.885 $X2=0 $Y2=0
cc_983 N_A_1790_75#_c_1461_n N_A_2604_392#_c_1613_n 0.0099279f $X=12.945
+ $Y=1.585 $X2=0 $Y2=0
cc_984 N_A_1790_75#_c_1462_n N_A_2604_392#_c_1613_n 0.00145958f $X=12.945
+ $Y=1.795 $X2=0 $Y2=0
cc_985 N_A_1790_75#_c_1478_n N_VPWR_c_1663_n 0.0165613f $X=9.925 $Y=2.53 $X2=0
+ $Y2=0
cc_986 N_A_1790_75#_c_1467_n N_VPWR_c_1664_n 0.00657334f $X=11.455 $Y=2.19 $X2=0
+ $Y2=0
cc_987 N_A_1790_75#_c_1468_n N_VPWR_c_1664_n 0.00817866f $X=11.455 $Y=2.28 $X2=0
+ $Y2=0
cc_988 N_A_1790_75#_c_1458_n N_VPWR_c_1664_n 0.00168841f $X=11.9 $Y=1.422 $X2=0
+ $Y2=0
cc_989 N_A_1790_75#_c_1469_n N_VPWR_c_1664_n 0.00877379f $X=11.99 $Y=1.765 $X2=0
+ $Y2=0
cc_990 N_A_1790_75#_c_1470_n N_VPWR_c_1665_n 0.00328506f $X=12.44 $Y=1.765 $X2=0
+ $Y2=0
cc_991 N_A_1790_75#_c_1461_n N_VPWR_c_1665_n 0.0105801f $X=12.945 $Y=1.585 $X2=0
+ $Y2=0
cc_992 N_A_1790_75#_c_1473_n N_VPWR_c_1665_n 0.00894992f $X=12.945 $Y=1.885
+ $X2=0 $Y2=0
cc_993 N_A_1790_75#_c_1473_n N_VPWR_c_1666_n 0.00461748f $X=12.945 $Y=1.885
+ $X2=0 $Y2=0
cc_994 N_A_1790_75#_c_1468_n N_VPWR_c_1675_n 0.00443738f $X=11.455 $Y=2.28 $X2=0
+ $Y2=0
cc_995 N_A_1790_75#_c_1469_n N_VPWR_c_1676_n 0.00422942f $X=11.99 $Y=1.765 $X2=0
+ $Y2=0
cc_996 N_A_1790_75#_c_1470_n N_VPWR_c_1676_n 0.00461464f $X=12.44 $Y=1.765 $X2=0
+ $Y2=0
cc_997 N_A_1790_75#_c_1473_n N_VPWR_c_1677_n 0.00461464f $X=12.945 $Y=1.885
+ $X2=0 $Y2=0
cc_998 N_A_1790_75#_c_1478_n N_VPWR_c_1683_n 0.00301353f $X=9.925 $Y=2.53 $X2=0
+ $Y2=0
cc_999 N_A_1790_75#_c_1468_n N_VPWR_c_1658_n 0.00489211f $X=11.455 $Y=2.28 $X2=0
+ $Y2=0
cc_1000 N_A_1790_75#_c_1469_n N_VPWR_c_1658_n 0.00789017f $X=11.99 $Y=1.765
+ $X2=0 $Y2=0
cc_1001 N_A_1790_75#_c_1470_n N_VPWR_c_1658_n 0.0090856f $X=12.44 $Y=1.765 $X2=0
+ $Y2=0
cc_1002 N_A_1790_75#_c_1473_n N_VPWR_c_1658_n 0.00913697f $X=12.945 $Y=1.885
+ $X2=0 $Y2=0
cc_1003 N_A_1790_75#_c_1478_n N_VPWR_c_1658_n 0.0291224f $X=9.925 $Y=2.53 $X2=0
+ $Y2=0
cc_1004 N_A_1790_75#_c_1478_n A_1955_471# 0.00419128f $X=9.925 $Y=2.53 $X2=-0.19
+ $Y2=-0.245
cc_1005 N_A_1790_75#_c_1467_n Q_N 9.68335e-19 $X=11.455 $Y=2.19 $X2=0 $Y2=0
cc_1006 N_A_1790_75#_c_1469_n Q_N 0.0159647f $X=11.99 $Y=1.765 $X2=0 $Y2=0
cc_1007 N_A_1790_75#_M1021_g Q_N 0.00434424f $X=12.085 $Y=0.74 $X2=0 $Y2=0
cc_1008 N_A_1790_75#_c_1470_n Q_N 0.00257754f $X=12.44 $Y=1.765 $X2=0 $Y2=0
cc_1009 N_A_1790_75#_M1037_g Q_N 0.00444052f $X=12.515 $Y=0.74 $X2=0 $Y2=0
cc_1010 N_A_1790_75#_c_1461_n Q_N 0.0512546f $X=12.945 $Y=1.585 $X2=0 $Y2=0
cc_1011 N_A_1790_75#_c_1462_n Q_N 8.09244e-19 $X=12.945 $Y=1.795 $X2=0 $Y2=0
cc_1012 N_A_1790_75#_M1021_g N_Q_N_c_2009_n 0.0129348f $X=12.085 $Y=0.74 $X2=0
+ $Y2=0
cc_1013 N_A_1790_75#_M1037_g N_Q_N_c_2009_n 0.0062067f $X=12.515 $Y=0.74 $X2=0
+ $Y2=0
cc_1014 N_A_1790_75#_M1005_g N_Q_N_c_2009_n 2.82358e-19 $X=12.99 $Y=0.69 $X2=0
+ $Y2=0
cc_1015 N_A_1790_75#_M1021_g Q_N 0.00845569f $X=12.085 $Y=0.74 $X2=0 $Y2=0
cc_1016 N_A_1790_75#_M1037_g Q_N 0.00357919f $X=12.515 $Y=0.74 $X2=0 $Y2=0
cc_1017 N_A_1790_75#_M1013_g N_VGND_c_2055_n 0.00182072f $X=11.075 $Y=0.58 $X2=0
+ $Y2=0
cc_1018 N_A_1790_75#_c_1480_n N_VGND_c_2055_n 0.0208351f $X=9.925 $Y=0.57 $X2=0
+ $Y2=0
cc_1019 N_A_1790_75#_c_1464_n N_VGND_c_2055_n 0.00424796f $X=10.01 $Y=1.045
+ $X2=0 $Y2=0
cc_1020 N_A_1790_75#_c_1466_n N_VGND_c_2055_n 0.0223381f $X=11.355 $Y=1.175
+ $X2=0 $Y2=0
cc_1021 N_A_1790_75#_M1013_g N_VGND_c_2056_n 0.00310691f $X=11.075 $Y=0.58 $X2=0
+ $Y2=0
cc_1022 N_A_1790_75#_M1021_g N_VGND_c_2056_n 0.00814486f $X=12.085 $Y=0.74 $X2=0
+ $Y2=0
cc_1023 N_A_1790_75#_M1037_g N_VGND_c_2057_n 0.0030832f $X=12.515 $Y=0.74 $X2=0
+ $Y2=0
cc_1024 N_A_1790_75#_c_1461_n N_VGND_c_2057_n 0.00620549f $X=12.945 $Y=1.585
+ $X2=0 $Y2=0
cc_1025 N_A_1790_75#_M1005_g N_VGND_c_2057_n 0.00352391f $X=12.99 $Y=0.69 $X2=0
+ $Y2=0
cc_1026 N_A_1790_75#_M1005_g N_VGND_c_2058_n 0.00461464f $X=12.99 $Y=0.69 $X2=0
+ $Y2=0
cc_1027 N_A_1790_75#_M1005_g N_VGND_c_2059_n 0.00385314f $X=12.99 $Y=0.69 $X2=0
+ $Y2=0
cc_1028 N_A_1790_75#_c_1480_n N_VGND_c_2066_n 0.0202724f $X=9.925 $Y=0.57 $X2=0
+ $Y2=0
cc_1029 N_A_1790_75#_M1013_g N_VGND_c_2069_n 0.00434272f $X=11.075 $Y=0.58 $X2=0
+ $Y2=0
cc_1030 N_A_1790_75#_M1021_g N_VGND_c_2070_n 0.00434272f $X=12.085 $Y=0.74 $X2=0
+ $Y2=0
cc_1031 N_A_1790_75#_M1037_g N_VGND_c_2070_n 0.00434272f $X=12.515 $Y=0.74 $X2=0
+ $Y2=0
cc_1032 N_A_1790_75#_M1013_g N_VGND_c_2078_n 0.00825669f $X=11.075 $Y=0.58 $X2=0
+ $Y2=0
cc_1033 N_A_1790_75#_M1021_g N_VGND_c_2078_n 0.00826269f $X=12.085 $Y=0.74 $X2=0
+ $Y2=0
cc_1034 N_A_1790_75#_M1037_g N_VGND_c_2078_n 0.00820493f $X=12.515 $Y=0.74 $X2=0
+ $Y2=0
cc_1035 N_A_1790_75#_M1005_g N_VGND_c_2078_n 0.00912981f $X=12.99 $Y=0.69 $X2=0
+ $Y2=0
cc_1036 N_A_1790_75#_c_1480_n N_VGND_c_2078_n 0.0221648f $X=9.925 $Y=0.57 $X2=0
+ $Y2=0
cc_1037 N_A_1790_75#_c_1480_n A_2000_74# 0.00371855f $X=9.925 $Y=0.57 $X2=-0.19
+ $Y2=-0.245
cc_1038 N_A_1790_75#_c_1464_n A_2000_74# 5.09211e-19 $X=10.01 $Y=1.045 $X2=-0.19
+ $Y2=-0.245
cc_1039 N_A_2604_392#_c_1612_n N_VPWR_c_1665_n 0.00374141f $X=13.17 $Y=2.105
+ $X2=0 $Y2=0
cc_1040 N_A_2604_392#_c_1614_n N_VPWR_c_1666_n 0.0177685f $X=13.935 $Y=1.765
+ $X2=0 $Y2=0
cc_1041 N_A_2604_392#_c_1615_n N_VPWR_c_1666_n 6.92538e-19 $X=14.385 $Y=1.765
+ $X2=0 $Y2=0
cc_1042 N_A_2604_392#_c_1609_n N_VPWR_c_1666_n 0.00687596f $X=13.845 $Y=1.465
+ $X2=0 $Y2=0
cc_1043 N_A_2604_392#_c_1610_n N_VPWR_c_1666_n 4.36456e-19 $X=14.385 $Y=1.532
+ $X2=0 $Y2=0
cc_1044 N_A_2604_392#_c_1612_n N_VPWR_c_1666_n 0.0792204f $X=13.17 $Y=2.105
+ $X2=0 $Y2=0
cc_1045 N_A_2604_392#_c_1631_p N_VPWR_c_1666_n 0.0253438f $X=13.8 $Y=1.465 $X2=0
+ $Y2=0
cc_1046 N_A_2604_392#_c_1615_n N_VPWR_c_1668_n 0.00508676f $X=14.385 $Y=1.765
+ $X2=0 $Y2=0
cc_1047 N_A_2604_392#_c_1612_n N_VPWR_c_1677_n 0.0115122f $X=13.17 $Y=2.105
+ $X2=0 $Y2=0
cc_1048 N_A_2604_392#_c_1614_n N_VPWR_c_1678_n 0.00413917f $X=13.935 $Y=1.765
+ $X2=0 $Y2=0
cc_1049 N_A_2604_392#_c_1615_n N_VPWR_c_1678_n 0.00445602f $X=14.385 $Y=1.765
+ $X2=0 $Y2=0
cc_1050 N_A_2604_392#_c_1614_n N_VPWR_c_1658_n 0.00817726f $X=13.935 $Y=1.765
+ $X2=0 $Y2=0
cc_1051 N_A_2604_392#_c_1615_n N_VPWR_c_1658_n 0.00860378f $X=14.385 $Y=1.765
+ $X2=0 $Y2=0
cc_1052 N_A_2604_392#_c_1612_n N_VPWR_c_1658_n 0.0095288f $X=13.17 $Y=2.105
+ $X2=0 $Y2=0
cc_1053 N_A_2604_392#_c_1611_n Q_N 0.00105746f $X=13.205 $Y=0.515 $X2=0 $Y2=0
cc_1054 N_A_2604_392#_c_1614_n N_Q_c_2036_n 0.00199967f $X=13.935 $Y=1.765 $X2=0
+ $Y2=0
cc_1055 N_A_2604_392#_M1017_g N_Q_c_2036_n 0.00531072f $X=13.97 $Y=0.74 $X2=0
+ $Y2=0
cc_1056 N_A_2604_392#_c_1615_n N_Q_c_2036_n 0.0153858f $X=14.385 $Y=1.765 $X2=0
+ $Y2=0
cc_1057 N_A_2604_392#_M1038_g N_Q_c_2036_n 0.00534388f $X=14.4 $Y=0.74 $X2=0
+ $Y2=0
cc_1058 N_A_2604_392#_c_1610_n N_Q_c_2036_n 0.045774f $X=14.385 $Y=1.532 $X2=0
+ $Y2=0
cc_1059 N_A_2604_392#_c_1631_p N_Q_c_2036_n 0.0258081f $X=13.8 $Y=1.465 $X2=0
+ $Y2=0
cc_1060 N_A_2604_392#_c_1611_n N_VGND_c_2057_n 0.0303376f $X=13.205 $Y=0.515
+ $X2=0 $Y2=0
cc_1061 N_A_2604_392#_c_1611_n N_VGND_c_2058_n 0.0115122f $X=13.205 $Y=0.515
+ $X2=0 $Y2=0
cc_1062 N_A_2604_392#_M1017_g N_VGND_c_2059_n 0.00508752f $X=13.97 $Y=0.74 $X2=0
+ $Y2=0
cc_1063 N_A_2604_392#_c_1609_n N_VGND_c_2059_n 0.00391367f $X=13.845 $Y=1.465
+ $X2=0 $Y2=0
cc_1064 N_A_2604_392#_c_1611_n N_VGND_c_2059_n 0.0350664f $X=13.205 $Y=0.515
+ $X2=0 $Y2=0
cc_1065 N_A_2604_392#_c_1631_p N_VGND_c_2059_n 0.014168f $X=13.8 $Y=1.465 $X2=0
+ $Y2=0
cc_1066 N_A_2604_392#_M1038_g N_VGND_c_2061_n 0.00543765f $X=14.4 $Y=0.74 $X2=0
+ $Y2=0
cc_1067 N_A_2604_392#_M1017_g N_VGND_c_2071_n 0.00461464f $X=13.97 $Y=0.74 $X2=0
+ $Y2=0
cc_1068 N_A_2604_392#_M1038_g N_VGND_c_2071_n 0.00461464f $X=14.4 $Y=0.74 $X2=0
+ $Y2=0
cc_1069 N_A_2604_392#_M1017_g N_VGND_c_2078_n 0.00913331f $X=13.97 $Y=0.74 $X2=0
+ $Y2=0
cc_1070 N_A_2604_392#_M1038_g N_VGND_c_2078_n 0.00911154f $X=14.4 $Y=0.74 $X2=0
+ $Y2=0
cc_1071 N_A_2604_392#_c_1611_n N_VGND_c_2078_n 0.0095288f $X=13.205 $Y=0.515
+ $X2=0 $Y2=0
cc_1072 N_VPWR_c_1673_n N_A_388_79#_c_1865_n 0.0287061f $X=3.115 $Y=3.33 $X2=0
+ $Y2=0
cc_1073 N_VPWR_c_1680_n N_A_388_79#_c_1865_n 0.00580289f $X=1.4 $Y=3.072 $X2=0
+ $Y2=0
cc_1074 N_VPWR_c_1658_n N_A_388_79#_c_1865_n 0.0336043f $X=14.64 $Y=3.33 $X2=0
+ $Y2=0
cc_1075 N_VPWR_M1031_d N_A_388_79#_c_1888_n 0.0106464f $X=3.11 $Y=2.32 $X2=0
+ $Y2=0
cc_1076 N_VPWR_c_1659_n N_A_388_79#_c_1888_n 0.0220425f $X=3.28 $Y=2.78 $X2=0
+ $Y2=0
cc_1077 N_VPWR_c_1658_n N_A_388_79#_c_1888_n 0.00587028f $X=14.64 $Y=3.33 $X2=0
+ $Y2=0
cc_1078 N_VPWR_M1031_d N_A_388_79#_c_1858_n 6.64982e-19 $X=3.11 $Y=2.32 $X2=0
+ $Y2=0
cc_1079 N_VPWR_c_1659_n N_A_388_79#_c_1858_n 0.0251321f $X=3.28 $Y=2.78 $X2=0
+ $Y2=0
cc_1080 N_VPWR_c_1669_n N_A_388_79#_c_1858_n 0.0166395f $X=4.705 $Y=3.33 $X2=0
+ $Y2=0
cc_1081 N_VPWR_c_1658_n N_A_388_79#_c_1858_n 0.0196698f $X=14.64 $Y=3.33 $X2=0
+ $Y2=0
cc_1082 N_VPWR_M1032_d N_A_388_79#_c_1859_n 0.0047096f $X=4.72 $Y=1.96 $X2=0
+ $Y2=0
cc_1083 N_VPWR_c_1660_n N_A_388_79#_c_1859_n 0.0166205f $X=4.87 $Y=2.835 $X2=0
+ $Y2=0
cc_1084 N_VPWR_c_1669_n N_A_388_79#_c_1859_n 7.47605e-19 $X=4.705 $Y=3.33 $X2=0
+ $Y2=0
cc_1085 N_VPWR_c_1671_n N_A_388_79#_c_1859_n 0.00867576f $X=7.07 $Y=3.33 $X2=0
+ $Y2=0
cc_1086 N_VPWR_c_1658_n N_A_388_79#_c_1859_n 0.0185655f $X=14.64 $Y=3.33 $X2=0
+ $Y2=0
cc_1087 N_VPWR_c_1669_n N_A_388_79#_c_1862_n 0.00886663f $X=4.705 $Y=3.33 $X2=0
+ $Y2=0
cc_1088 N_VPWR_c_1658_n N_A_388_79#_c_1862_n 0.0167388f $X=14.64 $Y=3.33 $X2=0
+ $Y2=0
cc_1089 N_VPWR_c_1671_n N_A_388_79#_c_1863_n 0.00576571f $X=7.07 $Y=3.33 $X2=0
+ $Y2=0
cc_1090 N_VPWR_c_1658_n N_A_388_79#_c_1863_n 0.00730692f $X=14.64 $Y=3.33 $X2=0
+ $Y2=0
cc_1091 N_VPWR_c_1664_n Q_N 0.0844051f $X=11.765 $Y=1.985 $X2=0 $Y2=0
cc_1092 N_VPWR_c_1665_n Q_N 0.00150368f $X=12.665 $Y=2.085 $X2=0 $Y2=0
cc_1093 N_VPWR_c_1676_n Q_N 0.014534f $X=12.54 $Y=3.33 $X2=0 $Y2=0
cc_1094 N_VPWR_c_1658_n Q_N 0.0119501f $X=14.64 $Y=3.33 $X2=0 $Y2=0
cc_1095 N_VPWR_c_1666_n N_Q_c_2036_n 0.0430489f $X=13.71 $Y=1.985 $X2=0 $Y2=0
cc_1096 N_VPWR_c_1668_n N_Q_c_2036_n 0.0437503f $X=14.61 $Y=1.985 $X2=0 $Y2=0
cc_1097 N_VPWR_c_1678_n N_Q_c_2036_n 0.0119166f $X=14.495 $Y=3.33 $X2=0 $Y2=0
cc_1098 N_VPWR_c_1658_n N_Q_c_2036_n 0.00983061f $X=14.64 $Y=3.33 $X2=0 $Y2=0
cc_1099 N_A_388_79#_c_1865_n A_538_464# 0.00358318f $X=2.775 $Y=2.785 $X2=-0.19
+ $Y2=-0.245
cc_1100 N_A_388_79#_c_1867_n A_538_464# 0.00186299f $X=2.86 $Y=2.66 $X2=-0.19
+ $Y2=-0.245
cc_1101 N_A_388_79#_c_1856_n A_538_464# 0.00712083f $X=2.945 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_1102 N_A_388_79#_M1023_d N_noxref_25_c_2208_n 0.011077f $X=1.94 $Y=0.395
+ $X2=0 $Y2=0
cc_1103 N_A_388_79#_c_1847_n N_noxref_25_c_2208_n 0.0217278f $X=2.435 $Y=0.68
+ $X2=0 $Y2=0
cc_1104 N_A_388_79#_c_1848_n N_noxref_25_c_2208_n 0.0118204f $X=3.445 $Y=1.09
+ $X2=0 $Y2=0
cc_1105 N_A_388_79#_c_1847_n N_noxref_25_c_2210_n 0.00763776f $X=2.435 $Y=0.68
+ $X2=0 $Y2=0
cc_1106 N_A_388_79#_c_1848_n N_noxref_25_c_2210_n 0.0271448f $X=3.445 $Y=1.09
+ $X2=0 $Y2=0
cc_1107 N_Q_N_c_2009_n N_VGND_c_2056_n 0.010788f $X=12.3 $Y=0.515 $X2=0 $Y2=0
cc_1108 N_Q_N_c_2009_n N_VGND_c_2057_n 0.0272093f $X=12.3 $Y=0.515 $X2=0 $Y2=0
cc_1109 N_Q_N_c_2009_n N_VGND_c_2070_n 0.0144922f $X=12.3 $Y=0.515 $X2=0 $Y2=0
cc_1110 N_Q_N_c_2009_n N_VGND_c_2078_n 0.0118826f $X=12.3 $Y=0.515 $X2=0 $Y2=0
cc_1111 N_Q_c_2036_n N_VGND_c_2059_n 0.00251281f $X=14.185 $Y=0.515 $X2=0 $Y2=0
cc_1112 N_Q_c_2036_n N_VGND_c_2061_n 0.0305242f $X=14.185 $Y=0.515 $X2=0 $Y2=0
cc_1113 N_Q_c_2036_n N_VGND_c_2071_n 0.0119584f $X=14.185 $Y=0.515 $X2=0 $Y2=0
cc_1114 N_Q_c_2036_n N_VGND_c_2078_n 0.00989813f $X=14.185 $Y=0.515 $X2=0 $Y2=0
cc_1115 N_VGND_c_2052_n N_noxref_25_c_2207_n 0.0278855f $X=0.71 $Y=0.605 $X2=0
+ $Y2=0
cc_1116 N_VGND_c_2053_n N_noxref_25_c_2208_n 0.0121474f $X=3.805 $Y=0.605 $X2=0
+ $Y2=0
cc_1117 N_VGND_c_2062_n N_noxref_25_c_2208_n 0.136372f $X=3.64 $Y=0 $X2=0 $Y2=0
cc_1118 N_VGND_c_2078_n N_noxref_25_c_2208_n 0.078753f $X=14.64 $Y=0 $X2=0 $Y2=0
cc_1119 N_VGND_c_2052_n N_noxref_25_c_2209_n 0.0125436f $X=0.71 $Y=0.605 $X2=0
+ $Y2=0
cc_1120 N_VGND_c_2062_n N_noxref_25_c_2209_n 0.0177095f $X=3.64 $Y=0 $X2=0 $Y2=0
cc_1121 N_VGND_c_2078_n N_noxref_25_c_2209_n 0.00967952f $X=14.64 $Y=0 $X2=0
+ $Y2=0
cc_1122 N_VGND_c_2053_n N_noxref_25_c_2210_n 0.0270493f $X=3.805 $Y=0.605 $X2=0
+ $Y2=0
cc_1123 N_noxref_25_c_2208_n noxref_26 0.00198134f $X=3.1 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_1124 N_noxref_25_c_2208_n noxref_27 0.00246354f $X=3.1 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
