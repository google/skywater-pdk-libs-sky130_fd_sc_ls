* File: sky130_fd_sc_ls__o21a_1.pxi.spice
* Created: Wed Sep  2 11:17:52 2020
* 
x_PM_SKY130_FD_SC_LS__O21A_1%A_83_244# N_A_83_244#_M1002_s N_A_83_244#_M1003_d
+ N_A_83_244#_c_50_n N_A_83_244#_M1006_g N_A_83_244#_c_51_n N_A_83_244#_M1005_g
+ N_A_83_244#_c_52_n N_A_83_244#_c_53_n N_A_83_244#_c_65_p N_A_83_244#_c_84_p
+ N_A_83_244#_c_54_n N_A_83_244#_c_55_n N_A_83_244#_c_58_n
+ PM_SKY130_FD_SC_LS__O21A_1%A_83_244#
x_PM_SKY130_FD_SC_LS__O21A_1%B1 N_B1_c_109_n N_B1_c_110_n N_B1_M1003_g
+ N_B1_M1002_g N_B1_c_111_n N_B1_c_112_n B1 PM_SKY130_FD_SC_LS__O21A_1%B1
x_PM_SKY130_FD_SC_LS__O21A_1%A2 N_A2_c_151_n N_A2_M1004_g N_A2_M1007_g A2
+ PM_SKY130_FD_SC_LS__O21A_1%A2
x_PM_SKY130_FD_SC_LS__O21A_1%A1 N_A1_c_182_n N_A1_M1000_g N_A1_M1001_g A1
+ N_A1_c_184_n PM_SKY130_FD_SC_LS__O21A_1%A1
x_PM_SKY130_FD_SC_LS__O21A_1%X N_X_M1006_s N_X_M1005_s X X X X X X X X
+ PM_SKY130_FD_SC_LS__O21A_1%X
x_PM_SKY130_FD_SC_LS__O21A_1%VPWR N_VPWR_M1005_d N_VPWR_M1000_d N_VPWR_c_221_n
+ N_VPWR_c_222_n N_VPWR_c_223_n VPWR N_VPWR_c_224_n N_VPWR_c_225_n
+ N_VPWR_c_226_n N_VPWR_c_220_n PM_SKY130_FD_SC_LS__O21A_1%VPWR
x_PM_SKY130_FD_SC_LS__O21A_1%VGND N_VGND_M1006_d N_VGND_M1007_d N_VGND_c_253_n
+ N_VGND_c_254_n VGND N_VGND_c_255_n N_VGND_c_256_n N_VGND_c_257_n
+ N_VGND_c_258_n N_VGND_c_259_n N_VGND_c_260_n PM_SKY130_FD_SC_LS__O21A_1%VGND
x_PM_SKY130_FD_SC_LS__O21A_1%A_320_74# N_A_320_74#_M1002_d N_A_320_74#_M1001_d
+ N_A_320_74#_c_292_n N_A_320_74#_c_293_n N_A_320_74#_c_294_n
+ N_A_320_74#_c_295_n PM_SKY130_FD_SC_LS__O21A_1%A_320_74#
cc_1 VNB N_A_83_244#_c_50_n 0.0225546f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.22
cc_2 VNB N_A_83_244#_c_51_n 0.0528845f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_3 VNB N_A_83_244#_c_52_n 0.00153256f $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=1.95
cc_4 VNB N_A_83_244#_c_53_n 0.0117976f $X=-0.19 $Y=-0.245 $X2=1.145 $Y2=1.19
cc_5 VNB N_A_83_244#_c_54_n 0.0105126f $X=-0.19 $Y=-0.245 $X2=1.31 $Y2=0.515
cc_6 VNB N_A_83_244#_c_55_n 0.00418063f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.19
cc_7 VNB N_B1_c_109_n 0.0264753f $X=-0.19 $Y=-0.245 $X2=1.375 $Y2=1.935
cc_8 VNB N_B1_c_110_n 0.00343846f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_B1_c_111_n 0.0169352f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_10 VNB N_B1_c_112_n 0.0349012f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_11 VNB B1 0.00336589f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_12 VNB N_A2_c_151_n 0.0182098f $X=-0.19 $Y=-0.245 $X2=1.165 $Y2=0.37
cc_13 VNB N_A2_M1007_g 0.0344726f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB A2 0.00593863f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_15 VNB N_A1_c_182_n 0.0606108f $X=-0.19 $Y=-0.245 $X2=1.165 $Y2=0.37
cc_16 VNB N_A1_M1001_g 0.03507f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A1_c_184_n 0.00431187f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_18 VNB X 0.0582938f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.22
cc_19 VNB N_VPWR_c_220_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_253_n 0.012579f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_21 VNB N_VGND_c_254_n 0.00396467f $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=1.55
cc_22 VNB N_VGND_c_255_n 0.0173909f $X=-0.19 $Y=-0.245 $X2=1.36 $Y2=2.035
cc_23 VNB N_VGND_c_256_n 0.0318625f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_257_n 0.0173909f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.385
cc_25 VNB N_VGND_c_258_n 0.197018f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.55
cc_26 VNB N_VGND_c_259_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.385
cc_27 VNB N_VGND_c_260_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_320_74#_c_292_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_29 VNB N_A_320_74#_c_293_n 0.013225f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_30 VNB N_A_320_74#_c_294_n 0.00558639f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_31 VNB N_A_320_74#_c_295_n 0.0247745f $X=-0.19 $Y=-0.245 $X2=1.145 $Y2=1.19
cc_32 VPB N_A_83_244#_c_51_n 0.0286454f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_33 VPB N_A_83_244#_c_52_n 0.00457714f $X=-0.19 $Y=1.66 $X2=0.78 $Y2=1.95
cc_34 VPB N_A_83_244#_c_58_n 0.0010391f $X=-0.19 $Y=1.66 $X2=1.525 $Y2=2.115
cc_35 VPB N_B1_c_110_n 0.0365124f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_36 VPB B1 0.00338512f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_37 VPB N_A2_c_151_n 0.0355028f $X=-0.19 $Y=1.66 $X2=1.165 $Y2=0.37
cc_38 VPB A2 0.015944f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_39 VPB N_A1_c_182_n 0.0353772f $X=-0.19 $Y=1.66 $X2=1.165 $Y2=0.37
cc_40 VPB N_A1_c_184_n 0.00764817f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_41 VPB X 0.00767567f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.22
cc_42 VPB X 0.0490703f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_43 VPB N_VPWR_c_221_n 0.0160289f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_44 VPB N_VPWR_c_222_n 0.0121909f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_45 VPB N_VPWR_c_223_n 0.0494883f $X=-0.19 $Y=1.66 $X2=0.78 $Y2=1.55
cc_46 VPB N_VPWR_c_224_n 0.0191515f $X=-0.19 $Y=1.66 $X2=1.27 $Y2=1.105
cc_47 VPB N_VPWR_c_225_n 0.0380926f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_226_n 0.0108417f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.385
cc_49 VPB N_VPWR_c_220_n 0.0806326f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 N_A_83_244#_c_51_n N_B1_c_109_n 0.00355615f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_51 N_A_83_244#_c_52_n N_B1_c_109_n 8.17514e-19 $X=0.78 $Y=1.95 $X2=0 $Y2=0
cc_52 N_A_83_244#_c_53_n N_B1_c_109_n 0.0062815f $X=1.145 $Y=1.19 $X2=0 $Y2=0
cc_53 N_A_83_244#_c_55_n N_B1_c_109_n 0.00132844f $X=0.7 $Y=1.19 $X2=0 $Y2=0
cc_54 N_A_83_244#_c_51_n N_B1_c_110_n 0.00829673f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_55 N_A_83_244#_c_52_n N_B1_c_110_n 0.00326333f $X=0.78 $Y=1.95 $X2=0 $Y2=0
cc_56 N_A_83_244#_c_65_p N_B1_c_110_n 0.0137036f $X=1.36 $Y=2.035 $X2=0 $Y2=0
cc_57 N_A_83_244#_c_58_n N_B1_c_110_n 0.0149767f $X=1.525 $Y=2.115 $X2=0 $Y2=0
cc_58 N_A_83_244#_c_54_n N_B1_c_111_n 0.00209693f $X=1.31 $Y=0.515 $X2=0 $Y2=0
cc_59 N_A_83_244#_c_50_n N_B1_c_112_n 0.00248076f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_60 N_A_83_244#_c_51_n N_B1_c_112_n 0.0189893f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_61 N_A_83_244#_c_53_n N_B1_c_112_n 0.00899946f $X=1.145 $Y=1.19 $X2=0 $Y2=0
cc_62 N_A_83_244#_c_54_n N_B1_c_112_n 0.00716644f $X=1.31 $Y=0.515 $X2=0 $Y2=0
cc_63 N_A_83_244#_c_51_n B1 6.62181e-19 $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_64 N_A_83_244#_c_53_n B1 0.0243916f $X=1.145 $Y=1.19 $X2=0 $Y2=0
cc_65 N_A_83_244#_c_65_p B1 0.018413f $X=1.36 $Y=2.035 $X2=0 $Y2=0
cc_66 N_A_83_244#_c_55_n B1 0.0220981f $X=0.7 $Y=1.19 $X2=0 $Y2=0
cc_67 N_A_83_244#_c_58_n B1 0.00374369f $X=1.525 $Y=2.115 $X2=0 $Y2=0
cc_68 N_A_83_244#_c_53_n N_A2_M1007_g 6.62318e-19 $X=1.145 $Y=1.19 $X2=0 $Y2=0
cc_69 N_A_83_244#_c_50_n X 0.0040121f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_70 N_A_83_244#_c_51_n X 0.0159981f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_71 N_A_83_244#_c_52_n X 0.0131415f $X=0.78 $Y=1.95 $X2=0 $Y2=0
cc_72 N_A_83_244#_c_55_n X 0.0341729f $X=0.7 $Y=1.19 $X2=0 $Y2=0
cc_73 N_A_83_244#_c_51_n X 0.0211799f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_74 N_A_83_244#_c_52_n X 0.00713749f $X=0.78 $Y=1.95 $X2=0 $Y2=0
cc_75 N_A_83_244#_c_84_p X 0.0104069f $X=0.865 $Y=2.035 $X2=0 $Y2=0
cc_76 N_A_83_244#_c_52_n N_VPWR_M1005_d 0.00214909f $X=0.78 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_77 N_A_83_244#_c_65_p N_VPWR_M1005_d 0.00999462f $X=1.36 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_78 N_A_83_244#_c_84_p N_VPWR_M1005_d 0.00515892f $X=0.865 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_79 N_A_83_244#_c_51_n N_VPWR_c_221_n 0.00548634f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_80 N_A_83_244#_c_65_p N_VPWR_c_221_n 0.0246152f $X=1.36 $Y=2.035 $X2=0 $Y2=0
cc_81 N_A_83_244#_c_84_p N_VPWR_c_221_n 0.0152373f $X=0.865 $Y=2.035 $X2=0 $Y2=0
cc_82 N_A_83_244#_c_58_n N_VPWR_c_221_n 0.0189233f $X=1.525 $Y=2.115 $X2=0 $Y2=0
cc_83 N_A_83_244#_c_51_n N_VPWR_c_224_n 0.00445602f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_84 N_A_83_244#_c_58_n N_VPWR_c_225_n 0.00786289f $X=1.525 $Y=2.115 $X2=0
+ $Y2=0
cc_85 N_A_83_244#_c_51_n N_VPWR_c_220_n 0.00865213f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_86 N_A_83_244#_c_58_n N_VPWR_c_220_n 0.010689f $X=1.525 $Y=2.115 $X2=0 $Y2=0
cc_87 N_A_83_244#_c_55_n N_VGND_M1006_d 0.00251343f $X=0.7 $Y=1.19 $X2=-0.19
+ $Y2=-0.245
cc_88 N_A_83_244#_c_50_n N_VGND_c_253_n 0.014482f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_89 N_A_83_244#_c_51_n N_VGND_c_253_n 0.00160934f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_90 N_A_83_244#_c_53_n N_VGND_c_253_n 7.60144e-19 $X=1.145 $Y=1.19 $X2=0 $Y2=0
cc_91 N_A_83_244#_c_54_n N_VGND_c_253_n 0.0345891f $X=1.31 $Y=0.515 $X2=0 $Y2=0
cc_92 N_A_83_244#_c_55_n N_VGND_c_253_n 0.0231389f $X=0.7 $Y=1.19 $X2=0 $Y2=0
cc_93 N_A_83_244#_c_50_n N_VGND_c_255_n 0.00383152f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_94 N_A_83_244#_c_54_n N_VGND_c_256_n 0.011066f $X=1.31 $Y=0.515 $X2=0 $Y2=0
cc_95 N_A_83_244#_c_50_n N_VGND_c_258_n 0.00761198f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_96 N_A_83_244#_c_54_n N_VGND_c_258_n 0.00915947f $X=1.31 $Y=0.515 $X2=0 $Y2=0
cc_97 N_A_83_244#_c_54_n N_A_320_74#_c_292_n 0.0216462f $X=1.31 $Y=0.515 $X2=0
+ $Y2=0
cc_98 N_A_83_244#_c_53_n N_A_320_74#_c_294_n 0.00198425f $X=1.145 $Y=1.19 $X2=0
+ $Y2=0
cc_99 N_A_83_244#_c_54_n N_A_320_74#_c_294_n 0.00929448f $X=1.31 $Y=0.515 $X2=0
+ $Y2=0
cc_100 N_B1_c_109_n N_A2_c_151_n 0.014966f $X=1.27 $Y=1.61 $X2=-0.19 $Y2=-0.245
cc_101 N_B1_c_110_n N_A2_c_151_n 0.0239503f $X=1.3 $Y=1.86 $X2=-0.19 $Y2=-0.245
cc_102 B1 N_A2_c_151_n 4.22595e-19 $X=1.115 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_103 N_B1_c_109_n N_A2_M1007_g 0.00719084f $X=1.27 $Y=1.61 $X2=0 $Y2=0
cc_104 N_B1_c_111_n N_A2_M1007_g 0.016626f $X=1.352 $Y=1.085 $X2=0 $Y2=0
cc_105 N_B1_c_109_n A2 4.2012e-19 $X=1.27 $Y=1.61 $X2=0 $Y2=0
cc_106 B1 A2 0.0176587f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_107 N_B1_c_110_n N_VPWR_c_221_n 0.00512313f $X=1.3 $Y=1.86 $X2=0 $Y2=0
cc_108 N_B1_c_110_n N_VPWR_c_225_n 0.00443738f $X=1.3 $Y=1.86 $X2=0 $Y2=0
cc_109 N_B1_c_110_n N_VPWR_c_220_n 0.00489211f $X=1.3 $Y=1.86 $X2=0 $Y2=0
cc_110 N_B1_c_111_n N_VGND_c_253_n 0.00372626f $X=1.352 $Y=1.085 $X2=0 $Y2=0
cc_111 N_B1_c_111_n N_VGND_c_254_n 6.90953e-19 $X=1.352 $Y=1.085 $X2=0 $Y2=0
cc_112 N_B1_c_111_n N_VGND_c_256_n 0.00434272f $X=1.352 $Y=1.085 $X2=0 $Y2=0
cc_113 N_B1_c_111_n N_VGND_c_258_n 0.00826366f $X=1.352 $Y=1.085 $X2=0 $Y2=0
cc_114 N_B1_c_111_n N_A_320_74#_c_292_n 0.00705529f $X=1.352 $Y=1.085 $X2=0
+ $Y2=0
cc_115 N_B1_c_111_n N_A_320_74#_c_294_n 0.00221692f $X=1.352 $Y=1.085 $X2=0
+ $Y2=0
cc_116 N_B1_c_112_n N_A_320_74#_c_294_n 0.00241027f $X=1.352 $Y=1.235 $X2=0
+ $Y2=0
cc_117 N_A2_c_151_n N_A1_c_182_n 0.0519818f $X=1.805 $Y=1.86 $X2=-0.19
+ $Y2=-0.245
cc_118 A2 N_A1_c_182_n 0.00293271f $X=2.075 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_119 N_A2_M1007_g N_A1_M1001_g 0.037899f $X=1.955 $Y=0.69 $X2=0 $Y2=0
cc_120 N_A2_c_151_n N_A1_c_184_n 2.29563e-19 $X=1.805 $Y=1.86 $X2=0 $Y2=0
cc_121 N_A2_M1007_g N_A1_c_184_n 6.91913e-19 $X=1.955 $Y=0.69 $X2=0 $Y2=0
cc_122 A2 N_A1_c_184_n 0.0276317f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_123 N_A2_c_151_n N_VPWR_c_221_n 0.0045081f $X=1.805 $Y=1.86 $X2=0 $Y2=0
cc_124 N_A2_c_151_n N_VPWR_c_223_n 0.00500475f $X=1.805 $Y=1.86 $X2=0 $Y2=0
cc_125 N_A2_c_151_n N_VPWR_c_225_n 0.00559701f $X=1.805 $Y=1.86 $X2=0 $Y2=0
cc_126 N_A2_c_151_n N_VPWR_c_220_n 0.00537853f $X=1.805 $Y=1.86 $X2=0 $Y2=0
cc_127 N_A2_M1007_g N_VGND_c_254_n 0.00929444f $X=1.955 $Y=0.69 $X2=0 $Y2=0
cc_128 N_A2_M1007_g N_VGND_c_256_n 0.00383152f $X=1.955 $Y=0.69 $X2=0 $Y2=0
cc_129 N_A2_M1007_g N_VGND_c_258_n 0.00757637f $X=1.955 $Y=0.69 $X2=0 $Y2=0
cc_130 N_A2_c_151_n N_A_320_74#_c_293_n 0.00159962f $X=1.805 $Y=1.86 $X2=0 $Y2=0
cc_131 N_A2_M1007_g N_A_320_74#_c_293_n 0.0144314f $X=1.955 $Y=0.69 $X2=0 $Y2=0
cc_132 A2 N_A_320_74#_c_293_n 0.0217572f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_133 N_A2_c_151_n N_A_320_74#_c_294_n 0.00268926f $X=1.805 $Y=1.86 $X2=0 $Y2=0
cc_134 A2 N_A_320_74#_c_294_n 0.00587011f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_135 N_A1_c_182_n N_VPWR_c_223_n 0.0268832f $X=2.375 $Y=1.86 $X2=0 $Y2=0
cc_136 N_A1_c_184_n N_VPWR_c_223_n 0.0258019f $X=2.61 $Y=1.465 $X2=0 $Y2=0
cc_137 N_A1_c_182_n N_VPWR_c_225_n 0.00502391f $X=2.375 $Y=1.86 $X2=0 $Y2=0
cc_138 N_A1_c_182_n N_VPWR_c_220_n 0.00487653f $X=2.375 $Y=1.86 $X2=0 $Y2=0
cc_139 N_A1_M1001_g N_VGND_c_254_n 0.0121806f $X=2.385 $Y=0.69 $X2=0 $Y2=0
cc_140 N_A1_M1001_g N_VGND_c_257_n 0.00383152f $X=2.385 $Y=0.69 $X2=0 $Y2=0
cc_141 N_A1_M1001_g N_VGND_c_258_n 0.00761198f $X=2.385 $Y=0.69 $X2=0 $Y2=0
cc_142 N_A1_c_182_n N_A_320_74#_c_293_n 0.00303926f $X=2.375 $Y=1.86 $X2=0 $Y2=0
cc_143 N_A1_M1001_g N_A_320_74#_c_293_n 0.0187748f $X=2.385 $Y=0.69 $X2=0 $Y2=0
cc_144 N_A1_c_184_n N_A_320_74#_c_293_n 0.0270164f $X=2.61 $Y=1.465 $X2=0 $Y2=0
cc_145 N_A1_M1001_g N_A_320_74#_c_295_n 4.43891e-19 $X=2.385 $Y=0.69 $X2=0 $Y2=0
cc_146 X N_VPWR_c_221_n 0.0267478f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_147 X N_VPWR_c_224_n 0.0145938f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_148 X N_VPWR_c_220_n 0.0120466f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_149 X N_VGND_c_253_n 0.0216951f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_150 X N_VGND_c_255_n 0.011066f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_151 X N_VGND_c_258_n 0.00915947f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_152 N_VGND_c_254_n N_A_320_74#_c_292_n 0.0164981f $X=2.17 $Y=0.57 $X2=0 $Y2=0
cc_153 N_VGND_c_256_n N_A_320_74#_c_292_n 0.0109942f $X=2.005 $Y=0 $X2=0 $Y2=0
cc_154 N_VGND_c_258_n N_A_320_74#_c_292_n 0.00904371f $X=2.64 $Y=0 $X2=0 $Y2=0
cc_155 N_VGND_M1007_d N_A_320_74#_c_293_n 0.00176461f $X=2.03 $Y=0.37 $X2=0
+ $Y2=0
cc_156 N_VGND_c_254_n N_A_320_74#_c_293_n 0.0171619f $X=2.17 $Y=0.57 $X2=0 $Y2=0
cc_157 N_VGND_c_254_n N_A_320_74#_c_295_n 0.0164982f $X=2.17 $Y=0.57 $X2=0 $Y2=0
cc_158 N_VGND_c_257_n N_A_320_74#_c_295_n 0.011066f $X=2.64 $Y=0 $X2=0 $Y2=0
cc_159 N_VGND_c_258_n N_A_320_74#_c_295_n 0.00915947f $X=2.64 $Y=0 $X2=0 $Y2=0
