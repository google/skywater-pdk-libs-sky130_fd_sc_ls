* File: sky130_fd_sc_ls__o2bb2a_2.pxi.spice
* Created: Fri Aug 28 13:50:12 2020
* 
x_PM_SKY130_FD_SC_LS__O2BB2A_2%B1 N_B1_M1011_g N_B1_c_84_n N_B1_M1007_g B1
+ N_B1_c_85_n PM_SKY130_FD_SC_LS__O2BB2A_2%B1
x_PM_SKY130_FD_SC_LS__O2BB2A_2%B2 N_B2_M1012_g N_B2_c_107_n N_B2_M1001_g B2
+ PM_SKY130_FD_SC_LS__O2BB2A_2%B2
x_PM_SKY130_FD_SC_LS__O2BB2A_2%A_270_48# N_A_270_48#_M1006_s N_A_270_48#_M1000_d
+ N_A_270_48#_M1009_g N_A_270_48#_c_136_n N_A_270_48#_M1002_g
+ N_A_270_48#_c_143_n N_A_270_48#_c_137_n N_A_270_48#_c_138_n
+ N_A_270_48#_c_171_p N_A_270_48#_c_153_p N_A_270_48#_c_139_n
+ N_A_270_48#_c_140_n N_A_270_48#_c_141_n PM_SKY130_FD_SC_LS__O2BB2A_2%A_270_48#
x_PM_SKY130_FD_SC_LS__O2BB2A_2%A2_N N_A2_N_c_203_n N_A2_N_M1000_g N_A2_N_c_204_n
+ N_A2_N_c_205_n N_A2_N_M1006_g N_A2_N_c_206_n A2_N
+ PM_SKY130_FD_SC_LS__O2BB2A_2%A2_N
x_PM_SKY130_FD_SC_LS__O2BB2A_2%A1_N N_A1_N_c_247_n N_A1_N_M1004_g N_A1_N_M1010_g
+ A1_N PM_SKY130_FD_SC_LS__O2BB2A_2%A1_N
x_PM_SKY130_FD_SC_LS__O2BB2A_2%A_201_392# N_A_201_392#_M1009_d
+ N_A_201_392#_M1001_d N_A_201_392#_c_296_n N_A_201_392#_M1005_g
+ N_A_201_392#_M1003_g N_A_201_392#_M1013_g N_A_201_392#_c_297_n
+ N_A_201_392#_M1008_g N_A_201_392#_c_298_n N_A_201_392#_c_299_n
+ N_A_201_392#_c_310_n N_A_201_392#_c_287_n N_A_201_392#_c_288_n
+ N_A_201_392#_c_289_n N_A_201_392#_c_290_n N_A_201_392#_c_291_n
+ N_A_201_392#_c_292_n N_A_201_392#_c_293_n N_A_201_392#_c_294_n
+ N_A_201_392#_c_327_n N_A_201_392#_c_295_n
+ PM_SKY130_FD_SC_LS__O2BB2A_2%A_201_392#
x_PM_SKY130_FD_SC_LS__O2BB2A_2%VPWR N_VPWR_M1007_s N_VPWR_M1002_d N_VPWR_M1004_d
+ N_VPWR_M1008_s N_VPWR_c_407_n N_VPWR_c_408_n N_VPWR_c_409_n N_VPWR_c_410_n
+ N_VPWR_c_411_n N_VPWR_c_412_n VPWR N_VPWR_c_413_n N_VPWR_c_414_n
+ N_VPWR_c_415_n N_VPWR_c_416_n N_VPWR_c_417_n N_VPWR_c_406_n
+ PM_SKY130_FD_SC_LS__O2BB2A_2%VPWR
x_PM_SKY130_FD_SC_LS__O2BB2A_2%X N_X_M1003_d N_X_M1005_d N_X_c_459_n N_X_c_460_n
+ X X X X N_X_c_461_n PM_SKY130_FD_SC_LS__O2BB2A_2%X
x_PM_SKY130_FD_SC_LS__O2BB2A_2%A_27_74# N_A_27_74#_M1011_s N_A_27_74#_M1012_d
+ N_A_27_74#_c_491_n N_A_27_74#_c_492_n N_A_27_74#_c_493_n N_A_27_74#_c_494_n
+ PM_SKY130_FD_SC_LS__O2BB2A_2%A_27_74#
x_PM_SKY130_FD_SC_LS__O2BB2A_2%VGND N_VGND_M1011_d N_VGND_M1010_d N_VGND_M1013_s
+ N_VGND_c_517_n N_VGND_c_518_n N_VGND_c_519_n N_VGND_c_520_n VGND
+ N_VGND_c_521_n N_VGND_c_522_n N_VGND_c_523_n N_VGND_c_524_n N_VGND_c_525_n
+ N_VGND_c_526_n PM_SKY130_FD_SC_LS__O2BB2A_2%VGND
cc_1 VNB N_B1_M1011_g 0.0379819f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_B1_c_84_n 0.0211941f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.885
cc_3 VNB N_B1_c_85_n 0.0104121f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.615
cc_4 VNB N_B2_M1012_g 0.0287799f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_5 VNB N_B2_c_107_n 0.0162389f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.885
cc_6 VNB B2 0.00404778f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_7 VNB N_A_270_48#_M1009_g 0.0364177f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_270_48#_c_136_n 0.0249562f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.615
cc_9 VNB N_A_270_48#_c_137_n 0.0149601f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_270_48#_c_138_n 0.00375376f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_270_48#_c_139_n 0.00589746f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_270_48#_c_140_n 0.00166222f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_270_48#_c_141_n 0.00298596f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A2_N_c_203_n 0.0177131f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.45
cc_15 VNB N_A2_N_c_204_n 0.0156143f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.885
cc_16 VNB N_A2_N_c_205_n 0.0171957f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.46
cc_17 VNB N_A2_N_c_206_n 0.0246559f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.615
cc_18 VNB A2_N 0.00165787f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.615
cc_19 VNB N_A1_N_c_247_n 0.0176223f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.45
cc_20 VNB N_A1_N_M1010_g 0.0363411f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.46
cc_21 VNB A1_N 0.00156355f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_22 VNB N_A_201_392#_M1003_g 0.0231615f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.615
cc_23 VNB N_A_201_392#_M1013_g 0.0263481f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.615
cc_24 VNB N_A_201_392#_c_287_n 0.00607937f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_201_392#_c_288_n 0.0166771f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_201_392#_c_289_n 0.00278702f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_201_392#_c_290_n 0.00184446f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_201_392#_c_291_n 0.00941197f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_201_392#_c_292_n 0.00210357f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_201_392#_c_293_n 0.00980048f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_201_392#_c_294_n 3.33931e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_201_392#_c_295_n 0.0750155f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VPWR_c_406_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_X_c_459_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_X_c_460_n 0.004293f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.615
cc_36 VNB N_X_c_461_n 0.00113445f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_27_74#_c_491_n 0.0302831f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_27_74#_c_492_n 0.0189843f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.615
cc_39 VNB N_A_27_74#_c_493_n 0.00975977f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.615
cc_40 VNB N_A_27_74#_c_494_n 0.00252706f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_517_n 0.00396467f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.615
cc_42 VNB N_VGND_c_518_n 0.00671515f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.615
cc_43 VNB N_VGND_c_519_n 0.0111565f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_520_n 0.0505285f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_521_n 0.0173909f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_522_n 0.0497142f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_523_n 0.0203669f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_524_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_525_n 0.00617641f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_526_n 0.256918f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VPB N_B1_c_84_n 0.0433409f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.885
cc_52 VPB N_B1_c_85_n 0.00566928f $X=-0.19 $Y=1.66 $X2=0.405 $Y2=1.615
cc_53 VPB N_B2_c_107_n 0.0361519f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.885
cc_54 VPB B2 0.00287247f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_55 VPB N_A_270_48#_c_136_n 0.0416577f $X=-0.19 $Y=1.66 $X2=0.405 $Y2=1.615
cc_56 VPB N_A_270_48#_c_143_n 0.0033648f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_A_270_48#_c_140_n 0.00138703f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_A2_N_c_203_n 0.0381399f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.45
cc_59 VPB A2_N 0.00138199f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.615
cc_60 VPB N_A1_N_c_247_n 0.0410346f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.45
cc_61 VPB A1_N 0.00102491f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_62 VPB N_A_201_392#_c_296_n 0.016431f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=2.46
cc_63 VPB N_A_201_392#_c_297_n 0.0173613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_A_201_392#_c_298_n 0.004308f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_A_201_392#_c_299_n 0.00296785f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_A_201_392#_c_294_n 0.00286179f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_A_201_392#_c_295_n 0.0169003f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_407_n 0.0121183f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.615
cc_69 VPB N_VPWR_c_408_n 0.0507181f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_409_n 0.0150337f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_410_n 0.0159763f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_411_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_412_n 0.0645697f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_413_n 0.033334f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_414_n 0.0263486f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_415_n 0.020646f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_416_n 0.00680245f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_417_n 0.00862975f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_406_n 0.0787592f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 VPB X 0.00182746f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB X 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 VPB N_X_c_461_n 8.32938e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 N_B1_M1011_g N_B2_M1012_g 0.0246174f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_84 N_B1_c_84_n N_B2_c_107_n 0.0785742f $X=0.51 $Y=1.885 $X2=0 $Y2=0
cc_85 N_B1_c_85_n N_B2_c_107_n 4.07543e-19 $X=0.405 $Y=1.615 $X2=0 $Y2=0
cc_86 N_B1_c_84_n B2 7.67374e-19 $X=0.51 $Y=1.885 $X2=0 $Y2=0
cc_87 N_B1_c_85_n B2 0.0198037f $X=0.405 $Y=1.615 $X2=0 $Y2=0
cc_88 N_B1_c_84_n N_VPWR_c_408_n 0.0282388f $X=0.51 $Y=1.885 $X2=0 $Y2=0
cc_89 N_B1_c_85_n N_VPWR_c_408_n 0.0277354f $X=0.405 $Y=1.615 $X2=0 $Y2=0
cc_90 N_B1_c_84_n N_VPWR_c_413_n 0.00413917f $X=0.51 $Y=1.885 $X2=0 $Y2=0
cc_91 N_B1_c_84_n N_VPWR_c_406_n 0.00817532f $X=0.51 $Y=1.885 $X2=0 $Y2=0
cc_92 N_B1_M1011_g N_A_27_74#_c_491_n 0.00159319f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_93 N_B1_M1011_g N_A_27_74#_c_492_n 0.0156808f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_94 N_B1_c_84_n N_A_27_74#_c_492_n 0.00219605f $X=0.51 $Y=1.885 $X2=0 $Y2=0
cc_95 N_B1_c_85_n N_A_27_74#_c_492_n 0.0148079f $X=0.405 $Y=1.615 $X2=0 $Y2=0
cc_96 N_B1_c_84_n N_A_27_74#_c_493_n 0.00291196f $X=0.51 $Y=1.885 $X2=0 $Y2=0
cc_97 N_B1_c_85_n N_A_27_74#_c_493_n 0.0207147f $X=0.405 $Y=1.615 $X2=0 $Y2=0
cc_98 N_B1_M1011_g N_VGND_c_517_n 0.0134383f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_99 N_B1_M1011_g N_VGND_c_521_n 0.00383152f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_100 N_B1_M1011_g N_VGND_c_526_n 0.00761198f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_101 N_B2_M1012_g N_A_270_48#_M1009_g 0.0253735f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_102 N_B2_c_107_n N_A_270_48#_c_136_n 0.0442787f $X=0.93 $Y=1.885 $X2=0 $Y2=0
cc_103 B2 N_A_270_48#_c_136_n 0.00246192f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_104 N_B2_c_107_n N_A_270_48#_c_140_n 2.64325e-19 $X=0.93 $Y=1.885 $X2=0 $Y2=0
cc_105 B2 N_A_270_48#_c_140_n 0.0268544f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_106 N_B2_c_107_n N_A_201_392#_c_298_n 0.00453614f $X=0.93 $Y=1.885 $X2=0
+ $Y2=0
cc_107 B2 N_A_201_392#_c_298_n 0.0203326f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_108 N_B2_c_107_n N_A_201_392#_c_299_n 0.00239916f $X=0.93 $Y=1.885 $X2=0
+ $Y2=0
cc_109 N_B2_M1012_g N_A_201_392#_c_289_n 3.08164e-19 $X=0.925 $Y=0.74 $X2=0
+ $Y2=0
cc_110 N_B2_c_107_n N_VPWR_c_408_n 0.00358919f $X=0.93 $Y=1.885 $X2=0 $Y2=0
cc_111 N_B2_c_107_n N_VPWR_c_413_n 0.00461464f $X=0.93 $Y=1.885 $X2=0 $Y2=0
cc_112 N_B2_c_107_n N_VPWR_c_406_n 0.00910115f $X=0.93 $Y=1.885 $X2=0 $Y2=0
cc_113 N_B2_M1012_g N_A_27_74#_c_492_n 0.0143059f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_114 N_B2_c_107_n N_A_27_74#_c_492_n 0.00416048f $X=0.93 $Y=1.885 $X2=0 $Y2=0
cc_115 B2 N_A_27_74#_c_492_n 0.0378094f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_116 N_B2_M1012_g N_A_27_74#_c_494_n 4.69391e-19 $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_117 N_B2_M1012_g N_VGND_c_517_n 0.0106075f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_118 N_B2_M1012_g N_VGND_c_522_n 0.00383152f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_119 N_B2_M1012_g N_VGND_c_526_n 0.00758251f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_120 N_A_270_48#_c_136_n N_A2_N_c_203_n 0.0414162f $X=1.44 $Y=1.885 $X2=-0.19
+ $Y2=-0.245
cc_121 N_A_270_48#_c_143_n N_A2_N_c_203_n 0.00382678f $X=1.7 $Y=1.975 $X2=-0.19
+ $Y2=-0.245
cc_122 N_A_270_48#_c_137_n N_A2_N_c_203_n 0.00135594f $X=2.045 $Y=1.22 $X2=-0.19
+ $Y2=-0.245
cc_123 N_A_270_48#_c_153_p N_A2_N_c_203_n 0.0125037f $X=2.355 $Y=2.14 $X2=-0.19
+ $Y2=-0.245
cc_124 N_A_270_48#_c_140_n N_A2_N_c_203_n 0.00106229f $X=1.62 $Y=1.615 $X2=-0.19
+ $Y2=-0.245
cc_125 N_A_270_48#_c_136_n N_A2_N_c_204_n 8.57091e-19 $X=1.44 $Y=1.885 $X2=0
+ $Y2=0
cc_126 N_A_270_48#_c_137_n N_A2_N_c_204_n 0.00498608f $X=2.045 $Y=1.22 $X2=0
+ $Y2=0
cc_127 N_A_270_48#_c_141_n N_A2_N_c_204_n 0.00265089f $X=1.62 $Y=1.45 $X2=0
+ $Y2=0
cc_128 N_A_270_48#_c_139_n N_A2_N_c_205_n 0.00725711f $X=2.21 $Y=0.81 $X2=0
+ $Y2=0
cc_129 N_A_270_48#_M1009_g N_A2_N_c_206_n 0.00362293f $X=1.425 $Y=0.74 $X2=0
+ $Y2=0
cc_130 N_A_270_48#_c_137_n N_A2_N_c_206_n 0.00538493f $X=2.045 $Y=1.22 $X2=0
+ $Y2=0
cc_131 N_A_270_48#_c_139_n N_A2_N_c_206_n 0.00587895f $X=2.21 $Y=0.81 $X2=0
+ $Y2=0
cc_132 N_A_270_48#_c_136_n A2_N 0.00111877f $X=1.44 $Y=1.885 $X2=0 $Y2=0
cc_133 N_A_270_48#_c_137_n A2_N 0.0267167f $X=2.045 $Y=1.22 $X2=0 $Y2=0
cc_134 N_A_270_48#_c_153_p A2_N 0.0218955f $X=2.355 $Y=2.14 $X2=0 $Y2=0
cc_135 N_A_270_48#_c_140_n A2_N 0.0208999f $X=1.62 $Y=1.615 $X2=0 $Y2=0
cc_136 N_A_270_48#_c_153_p N_A1_N_c_247_n 0.00500523f $X=2.355 $Y=2.14 $X2=-0.19
+ $Y2=-0.245
cc_137 N_A_270_48#_c_137_n N_A1_N_M1010_g 2.68167e-19 $X=2.045 $Y=1.22 $X2=0
+ $Y2=0
cc_138 N_A_270_48#_c_153_p A1_N 0.00204545f $X=2.355 $Y=2.14 $X2=0 $Y2=0
cc_139 N_A_270_48#_c_136_n N_A_201_392#_c_298_n 0.00824224f $X=1.44 $Y=1.885
+ $X2=0 $Y2=0
cc_140 N_A_270_48#_c_143_n N_A_201_392#_c_298_n 0.00142443f $X=1.7 $Y=1.975
+ $X2=0 $Y2=0
cc_141 N_A_270_48#_c_171_p N_A_201_392#_c_298_n 0.0160892f $X=1.785 $Y=2.1 $X2=0
+ $Y2=0
cc_142 N_A_270_48#_c_136_n N_A_201_392#_c_299_n 0.00648576f $X=1.44 $Y=1.885
+ $X2=0 $Y2=0
cc_143 N_A_270_48#_M1000_d N_A_201_392#_c_310_n 0.00830827f $X=2.16 $Y=1.965
+ $X2=0 $Y2=0
cc_144 N_A_270_48#_c_136_n N_A_201_392#_c_310_n 0.013643f $X=1.44 $Y=1.885 $X2=0
+ $Y2=0
cc_145 N_A_270_48#_c_171_p N_A_201_392#_c_310_n 0.0137412f $X=1.785 $Y=2.1 $X2=0
+ $Y2=0
cc_146 N_A_270_48#_c_153_p N_A_201_392#_c_310_n 0.0446228f $X=2.355 $Y=2.14
+ $X2=0 $Y2=0
cc_147 N_A_270_48#_c_140_n N_A_201_392#_c_310_n 0.00334664f $X=1.62 $Y=1.615
+ $X2=0 $Y2=0
cc_148 N_A_270_48#_M1009_g N_A_201_392#_c_287_n 0.00610421f $X=1.425 $Y=0.74
+ $X2=0 $Y2=0
cc_149 N_A_270_48#_c_136_n N_A_201_392#_c_287_n 0.00120384f $X=1.44 $Y=1.885
+ $X2=0 $Y2=0
cc_150 N_A_270_48#_c_137_n N_A_201_392#_c_287_n 0.00157271f $X=2.045 $Y=1.22
+ $X2=0 $Y2=0
cc_151 N_A_270_48#_c_138_n N_A_201_392#_c_287_n 0.0156773f $X=1.785 $Y=1.22
+ $X2=0 $Y2=0
cc_152 N_A_270_48#_c_139_n N_A_201_392#_c_287_n 0.0242222f $X=2.21 $Y=0.81 $X2=0
+ $Y2=0
cc_153 N_A_270_48#_c_140_n N_A_201_392#_c_287_n 0.00385199f $X=1.62 $Y=1.615
+ $X2=0 $Y2=0
cc_154 N_A_270_48#_M1006_s N_A_201_392#_c_288_n 0.00264658f $X=2.065 $Y=0.37
+ $X2=0 $Y2=0
cc_155 N_A_270_48#_c_139_n N_A_201_392#_c_288_n 0.020634f $X=2.21 $Y=0.81 $X2=0
+ $Y2=0
cc_156 N_A_270_48#_M1009_g N_A_201_392#_c_289_n 0.00544881f $X=1.425 $Y=0.74
+ $X2=0 $Y2=0
cc_157 N_A_270_48#_c_139_n N_A_201_392#_c_290_n 0.0248147f $X=2.21 $Y=0.81 $X2=0
+ $Y2=0
cc_158 N_A_270_48#_c_137_n N_A_201_392#_c_292_n 0.0155236f $X=2.045 $Y=1.22
+ $X2=0 $Y2=0
cc_159 N_A_270_48#_c_153_p N_A_201_392#_c_294_n 0.0081071f $X=2.355 $Y=2.14
+ $X2=0 $Y2=0
cc_160 N_A_270_48#_c_136_n N_A_201_392#_c_327_n 2.24111e-19 $X=1.44 $Y=1.885
+ $X2=0 $Y2=0
cc_161 N_A_270_48#_c_143_n N_VPWR_M1002_d 3.68124e-19 $X=1.7 $Y=1.975 $X2=0
+ $Y2=0
cc_162 N_A_270_48#_c_171_p N_VPWR_M1002_d 0.00655923f $X=1.785 $Y=2.1 $X2=0
+ $Y2=0
cc_163 N_A_270_48#_c_153_p N_VPWR_M1002_d 0.00574422f $X=2.355 $Y=2.14 $X2=0
+ $Y2=0
cc_164 N_A_270_48#_c_136_n N_VPWR_c_409_n 0.00764758f $X=1.44 $Y=1.885 $X2=0
+ $Y2=0
cc_165 N_A_270_48#_c_136_n N_VPWR_c_413_n 0.00445602f $X=1.44 $Y=1.885 $X2=0
+ $Y2=0
cc_166 N_A_270_48#_c_136_n N_VPWR_c_406_n 0.00441354f $X=1.44 $Y=1.885 $X2=0
+ $Y2=0
cc_167 N_A_270_48#_M1009_g N_A_27_74#_c_492_n 0.00252956f $X=1.425 $Y=0.74 $X2=0
+ $Y2=0
cc_168 N_A_270_48#_c_138_n N_A_27_74#_c_492_n 0.00890055f $X=1.785 $Y=1.22 $X2=0
+ $Y2=0
cc_169 N_A_270_48#_M1009_g N_A_27_74#_c_494_n 0.00402051f $X=1.425 $Y=0.74 $X2=0
+ $Y2=0
cc_170 N_A_270_48#_M1009_g N_VGND_c_517_n 5.20809e-19 $X=1.425 $Y=0.74 $X2=0
+ $Y2=0
cc_171 N_A_270_48#_M1009_g N_VGND_c_522_n 0.00430908f $X=1.425 $Y=0.74 $X2=0
+ $Y2=0
cc_172 N_A_270_48#_M1009_g N_VGND_c_526_n 0.00822378f $X=1.425 $Y=0.74 $X2=0
+ $Y2=0
cc_173 N_A2_N_c_203_n N_A1_N_c_247_n 0.046381f $X=2.085 $Y=1.89 $X2=-0.19
+ $Y2=-0.245
cc_174 A2_N N_A1_N_c_247_n 4.04807e-19 $X=2.075 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_175 N_A2_N_c_204_n N_A1_N_M1010_g 0.0078326f $X=2.25 $Y=1.475 $X2=0 $Y2=0
cc_176 N_A2_N_c_205_n N_A1_N_M1010_g 0.0451706f $X=2.425 $Y=1.085 $X2=0 $Y2=0
cc_177 N_A2_N_c_203_n A1_N 0.00187659f $X=2.085 $Y=1.89 $X2=0 $Y2=0
cc_178 A2_N A1_N 0.0231358f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_179 N_A2_N_c_203_n N_A_201_392#_c_298_n 9.06284e-19 $X=2.085 $Y=1.89 $X2=0
+ $Y2=0
cc_180 N_A2_N_c_203_n N_A_201_392#_c_299_n 7.70097e-19 $X=2.085 $Y=1.89 $X2=0
+ $Y2=0
cc_181 N_A2_N_c_203_n N_A_201_392#_c_310_n 0.0129975f $X=2.085 $Y=1.89 $X2=0
+ $Y2=0
cc_182 N_A2_N_c_205_n N_A_201_392#_c_287_n 0.00494986f $X=2.425 $Y=1.085 $X2=0
+ $Y2=0
cc_183 N_A2_N_c_205_n N_A_201_392#_c_288_n 0.0143941f $X=2.425 $Y=1.085 $X2=0
+ $Y2=0
cc_184 N_A2_N_c_206_n N_A_201_392#_c_288_n 4.10115e-19 $X=2.425 $Y=1.16 $X2=0
+ $Y2=0
cc_185 N_A2_N_c_205_n N_A_201_392#_c_290_n 0.00304192f $X=2.425 $Y=1.085 $X2=0
+ $Y2=0
cc_186 N_A2_N_c_204_n N_A_201_392#_c_292_n 2.70295e-19 $X=2.25 $Y=1.475 $X2=0
+ $Y2=0
cc_187 N_A2_N_c_206_n N_A_201_392#_c_292_n 8.38832e-19 $X=2.425 $Y=1.16 $X2=0
+ $Y2=0
cc_188 N_A2_N_c_203_n N_VPWR_c_409_n 0.00590139f $X=2.085 $Y=1.89 $X2=0 $Y2=0
cc_189 N_A2_N_c_203_n N_VPWR_c_414_n 0.00472107f $X=2.085 $Y=1.89 $X2=0 $Y2=0
cc_190 N_A2_N_c_203_n N_VPWR_c_406_n 0.0049796f $X=2.085 $Y=1.89 $X2=0 $Y2=0
cc_191 N_A2_N_c_205_n N_VGND_c_518_n 3.72445e-19 $X=2.425 $Y=1.085 $X2=0 $Y2=0
cc_192 N_A2_N_c_205_n N_VGND_c_522_n 0.00278271f $X=2.425 $Y=1.085 $X2=0 $Y2=0
cc_193 N_A2_N_c_205_n N_VGND_c_526_n 0.00358137f $X=2.425 $Y=1.085 $X2=0 $Y2=0
cc_194 N_A1_N_c_247_n N_A_201_392#_c_296_n 0.0167426f $X=2.625 $Y=1.89 $X2=0
+ $Y2=0
cc_195 N_A1_N_M1010_g N_A_201_392#_M1003_g 0.0165087f $X=2.815 $Y=0.69 $X2=0
+ $Y2=0
cc_196 N_A1_N_c_247_n N_A_201_392#_c_310_n 0.0182845f $X=2.625 $Y=1.89 $X2=0
+ $Y2=0
cc_197 A1_N N_A_201_392#_c_310_n 0.00721403f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_198 N_A1_N_M1010_g N_A_201_392#_c_288_n 0.0011351f $X=2.815 $Y=0.69 $X2=0
+ $Y2=0
cc_199 N_A1_N_M1010_g N_A_201_392#_c_290_n 0.0052743f $X=2.815 $Y=0.69 $X2=0
+ $Y2=0
cc_200 N_A1_N_c_247_n N_A_201_392#_c_291_n 5.5832e-19 $X=2.625 $Y=1.89 $X2=0
+ $Y2=0
cc_201 N_A1_N_M1010_g N_A_201_392#_c_291_n 0.0153044f $X=2.815 $Y=0.69 $X2=0
+ $Y2=0
cc_202 A1_N N_A_201_392#_c_291_n 0.0107679f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_203 N_A1_N_c_247_n N_A_201_392#_c_292_n 0.00457362f $X=2.625 $Y=1.89 $X2=0
+ $Y2=0
cc_204 A1_N N_A_201_392#_c_292_n 0.0143367f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_205 N_A1_N_M1010_g N_A_201_392#_c_293_n 0.00478972f $X=2.815 $Y=0.69 $X2=0
+ $Y2=0
cc_206 A1_N N_A_201_392#_c_293_n 0.0105181f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_207 N_A1_N_c_247_n N_A_201_392#_c_294_n 0.00958751f $X=2.625 $Y=1.89 $X2=0
+ $Y2=0
cc_208 A1_N N_A_201_392#_c_294_n 0.0105017f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_209 N_A1_N_c_247_n N_A_201_392#_c_295_n 0.0031468f $X=2.625 $Y=1.89 $X2=0
+ $Y2=0
cc_210 N_A1_N_M1010_g N_A_201_392#_c_295_n 0.020241f $X=2.815 $Y=0.69 $X2=0
+ $Y2=0
cc_211 N_A1_N_c_247_n N_VPWR_c_410_n 0.00635186f $X=2.625 $Y=1.89 $X2=0 $Y2=0
cc_212 N_A1_N_c_247_n N_VPWR_c_414_n 0.00472107f $X=2.625 $Y=1.89 $X2=0 $Y2=0
cc_213 N_A1_N_c_247_n N_VPWR_c_406_n 0.0049796f $X=2.625 $Y=1.89 $X2=0 $Y2=0
cc_214 N_A1_N_M1010_g N_X_c_460_n 6.44522e-19 $X=2.815 $Y=0.69 $X2=0 $Y2=0
cc_215 N_A1_N_M1010_g N_VGND_c_518_n 0.00814171f $X=2.815 $Y=0.69 $X2=0 $Y2=0
cc_216 N_A1_N_M1010_g N_VGND_c_522_n 0.00444681f $X=2.815 $Y=0.69 $X2=0 $Y2=0
cc_217 N_A1_N_M1010_g N_VGND_c_526_n 0.00877228f $X=2.815 $Y=0.69 $X2=0 $Y2=0
cc_218 N_A_201_392#_c_310_n N_VPWR_M1002_d 0.00955667f $X=3.085 $Y=2.48 $X2=0
+ $Y2=0
cc_219 N_A_201_392#_c_310_n N_VPWR_M1004_d 0.0182171f $X=3.085 $Y=2.48 $X2=0
+ $Y2=0
cc_220 N_A_201_392#_c_294_n N_VPWR_M1004_d 0.012403f $X=3.17 $Y=2.395 $X2=0
+ $Y2=0
cc_221 N_A_201_392#_c_298_n N_VPWR_c_408_n 0.00603256f $X=1.215 $Y=2.115 $X2=0
+ $Y2=0
cc_222 N_A_201_392#_c_299_n N_VPWR_c_408_n 0.00580658f $X=1.215 $Y=2.815 $X2=0
+ $Y2=0
cc_223 N_A_201_392#_c_299_n N_VPWR_c_409_n 0.016592f $X=1.215 $Y=2.815 $X2=0
+ $Y2=0
cc_224 N_A_201_392#_c_310_n N_VPWR_c_409_n 0.0278856f $X=3.085 $Y=2.48 $X2=0
+ $Y2=0
cc_225 N_A_201_392#_c_296_n N_VPWR_c_410_n 0.00803088f $X=3.365 $Y=1.765 $X2=0
+ $Y2=0
cc_226 N_A_201_392#_c_310_n N_VPWR_c_410_n 0.0364237f $X=3.085 $Y=2.48 $X2=0
+ $Y2=0
cc_227 N_A_201_392#_c_297_n N_VPWR_c_412_n 0.00981831f $X=3.815 $Y=1.765 $X2=0
+ $Y2=0
cc_228 N_A_201_392#_c_299_n N_VPWR_c_413_n 0.0145938f $X=1.215 $Y=2.815 $X2=0
+ $Y2=0
cc_229 N_A_201_392#_c_296_n N_VPWR_c_415_n 0.00445602f $X=3.365 $Y=1.765 $X2=0
+ $Y2=0
cc_230 N_A_201_392#_c_297_n N_VPWR_c_415_n 0.00428607f $X=3.815 $Y=1.765 $X2=0
+ $Y2=0
cc_231 N_A_201_392#_c_296_n N_VPWR_c_406_n 0.00862503f $X=3.365 $Y=1.765 $X2=0
+ $Y2=0
cc_232 N_A_201_392#_c_297_n N_VPWR_c_406_n 0.00806054f $X=3.815 $Y=1.765 $X2=0
+ $Y2=0
cc_233 N_A_201_392#_c_299_n N_VPWR_c_406_n 0.0120466f $X=1.215 $Y=2.815 $X2=0
+ $Y2=0
cc_234 N_A_201_392#_c_310_n N_VPWR_c_406_n 0.040738f $X=3.085 $Y=2.48 $X2=0
+ $Y2=0
cc_235 N_A_201_392#_M1003_g N_X_c_459_n 0.00812178f $X=3.38 $Y=0.74 $X2=0 $Y2=0
cc_236 N_A_201_392#_M1013_g N_X_c_459_n 0.0081896f $X=3.81 $Y=0.74 $X2=0 $Y2=0
cc_237 N_A_201_392#_M1003_g N_X_c_460_n 0.00485634f $X=3.38 $Y=0.74 $X2=0 $Y2=0
cc_238 N_A_201_392#_M1013_g N_X_c_460_n 0.00215589f $X=3.81 $Y=0.74 $X2=0 $Y2=0
cc_239 N_A_201_392#_c_295_n N_X_c_460_n 0.0024311f $X=3.81 $Y=1.535 $X2=0 $Y2=0
cc_240 N_A_201_392#_c_296_n X 0.0026829f $X=3.365 $Y=1.765 $X2=0 $Y2=0
cc_241 N_A_201_392#_c_297_n X 0.0022003f $X=3.815 $Y=1.765 $X2=0 $Y2=0
cc_242 N_A_201_392#_c_294_n X 0.0223997f $X=3.17 $Y=2.395 $X2=0 $Y2=0
cc_243 N_A_201_392#_c_295_n X 0.00751256f $X=3.81 $Y=1.535 $X2=0 $Y2=0
cc_244 N_A_201_392#_c_296_n X 0.0166429f $X=3.365 $Y=1.765 $X2=0 $Y2=0
cc_245 N_A_201_392#_c_297_n X 0.012401f $X=3.815 $Y=1.765 $X2=0 $Y2=0
cc_246 N_A_201_392#_M1003_g N_X_c_461_n 9.7705e-19 $X=3.38 $Y=0.74 $X2=0 $Y2=0
cc_247 N_A_201_392#_M1013_g N_X_c_461_n 0.00886097f $X=3.81 $Y=0.74 $X2=0 $Y2=0
cc_248 N_A_201_392#_c_297_n N_X_c_461_n 0.00295823f $X=3.815 $Y=1.765 $X2=0
+ $Y2=0
cc_249 N_A_201_392#_c_293_n N_X_c_461_n 0.0302315f $X=3.17 $Y=1.635 $X2=0 $Y2=0
cc_250 N_A_201_392#_c_294_n N_X_c_461_n 0.00618574f $X=3.17 $Y=2.395 $X2=0 $Y2=0
cc_251 N_A_201_392#_c_295_n N_X_c_461_n 0.0342738f $X=3.81 $Y=1.535 $X2=0 $Y2=0
cc_252 N_A_201_392#_c_298_n N_A_27_74#_c_492_n 7.14544e-19 $X=1.215 $Y=2.115
+ $X2=0 $Y2=0
cc_253 N_A_201_392#_c_289_n N_A_27_74#_c_494_n 0.00392044f $X=1.805 $Y=0.34
+ $X2=0 $Y2=0
cc_254 N_A_201_392#_c_289_n N_VGND_c_517_n 0.00266256f $X=1.805 $Y=0.34 $X2=0
+ $Y2=0
cc_255 N_A_201_392#_M1003_g N_VGND_c_518_n 0.00866971f $X=3.38 $Y=0.74 $X2=0
+ $Y2=0
cc_256 N_A_201_392#_c_288_n N_VGND_c_518_n 0.0117236f $X=2.545 $Y=0.34 $X2=0
+ $Y2=0
cc_257 N_A_201_392#_c_291_n N_VGND_c_518_n 0.013791f $X=3.085 $Y=1.22 $X2=0
+ $Y2=0
cc_258 N_A_201_392#_c_293_n N_VGND_c_518_n 0.0118589f $X=3.17 $Y=1.635 $X2=0
+ $Y2=0
cc_259 N_A_201_392#_c_295_n N_VGND_c_518_n 6.03907e-19 $X=3.81 $Y=1.535 $X2=0
+ $Y2=0
cc_260 N_A_201_392#_M1013_g N_VGND_c_520_n 0.00646793f $X=3.81 $Y=0.74 $X2=0
+ $Y2=0
cc_261 N_A_201_392#_c_288_n N_VGND_c_522_n 0.0593614f $X=2.545 $Y=0.34 $X2=0
+ $Y2=0
cc_262 N_A_201_392#_c_289_n N_VGND_c_522_n 0.0236456f $X=1.805 $Y=0.34 $X2=0
+ $Y2=0
cc_263 N_A_201_392#_M1003_g N_VGND_c_523_n 0.00434272f $X=3.38 $Y=0.74 $X2=0
+ $Y2=0
cc_264 N_A_201_392#_M1013_g N_VGND_c_523_n 0.00422942f $X=3.81 $Y=0.74 $X2=0
+ $Y2=0
cc_265 N_A_201_392#_M1003_g N_VGND_c_526_n 0.00822284f $X=3.38 $Y=0.74 $X2=0
+ $Y2=0
cc_266 N_A_201_392#_M1013_g N_VGND_c_526_n 0.00787305f $X=3.81 $Y=0.74 $X2=0
+ $Y2=0
cc_267 N_A_201_392#_c_288_n N_VGND_c_526_n 0.0337409f $X=2.545 $Y=0.34 $X2=0
+ $Y2=0
cc_268 N_A_201_392#_c_289_n N_VGND_c_526_n 0.0127298f $X=1.805 $Y=0.34 $X2=0
+ $Y2=0
cc_269 N_A_201_392#_c_290_n A_500_74# 0.00249342f $X=2.63 $Y=1.135 $X2=-0.19
+ $Y2=-0.245
cc_270 N_VPWR_c_412_n X 0.0828853f $X=4.04 $Y=1.985 $X2=0 $Y2=0
cc_271 N_VPWR_c_410_n X 0.0169587f $X=2.995 $Y=2.9 $X2=0 $Y2=0
cc_272 N_VPWR_c_415_n X 0.0151764f $X=3.955 $Y=3.33 $X2=0 $Y2=0
cc_273 N_VPWR_c_406_n X 0.0124607f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_274 N_X_c_459_n N_VGND_c_518_n 0.0399419f $X=3.595 $Y=0.515 $X2=0 $Y2=0
cc_275 N_X_c_459_n N_VGND_c_520_n 0.0308798f $X=3.595 $Y=0.515 $X2=0 $Y2=0
cc_276 N_X_c_459_n N_VGND_c_523_n 0.0149085f $X=3.595 $Y=0.515 $X2=0 $Y2=0
cc_277 N_X_c_459_n N_VGND_c_526_n 0.0122037f $X=3.595 $Y=0.515 $X2=0 $Y2=0
cc_278 N_A_27_74#_c_491_n N_VGND_c_517_n 0.0218743f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_279 N_A_27_74#_c_492_n N_VGND_c_517_n 0.0216087f $X=1.055 $Y=1.195 $X2=0
+ $Y2=0
cc_280 N_A_27_74#_c_494_n N_VGND_c_517_n 0.0218743f $X=1.14 $Y=0.515 $X2=0 $Y2=0
cc_281 N_A_27_74#_c_491_n N_VGND_c_521_n 0.011066f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_282 N_A_27_74#_c_494_n N_VGND_c_522_n 0.011066f $X=1.14 $Y=0.515 $X2=0 $Y2=0
cc_283 N_A_27_74#_c_491_n N_VGND_c_526_n 0.00915947f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_284 N_A_27_74#_c_494_n N_VGND_c_526_n 0.00915947f $X=1.14 $Y=0.515 $X2=0
+ $Y2=0
