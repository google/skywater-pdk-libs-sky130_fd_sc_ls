* File: sky130_fd_sc_ls__nor2_8.pex.spice
* Created: Fri Aug 28 13:37:18 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__NOR2_8%A 1 3 4 5 6 8 9 11 13 14 18 20 22 25 27 29 30
+ 32 35 37 39 42 44 46 47 48 49 50 51 52 53 72
r139 70 72 37.2747 $w=3.75e-07 $l=2.9e-07 $layer=POLY_cond $X=3.42 $Y=1.557
+ $X2=3.71 $Y2=1.557
r140 70 71 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=3.42
+ $Y=1.515 $X2=3.42 $Y2=1.515
r141 68 70 14.7813 $w=3.75e-07 $l=1.15e-07 $layer=POLY_cond $X=3.305 $Y=1.557
+ $X2=3.42 $Y2=1.557
r142 67 68 12.2107 $w=3.75e-07 $l=9.5e-08 $layer=POLY_cond $X=3.21 $Y=1.557
+ $X2=3.305 $Y2=1.557
r143 66 67 45.6293 $w=3.75e-07 $l=3.55e-07 $layer=POLY_cond $X=2.855 $Y=1.557
+ $X2=3.21 $Y2=1.557
r144 65 66 64.2667 $w=3.75e-07 $l=5e-07 $layer=POLY_cond $X=2.355 $Y=1.557
+ $X2=2.855 $Y2=1.557
r145 64 65 5.784 $w=3.75e-07 $l=4.5e-08 $layer=POLY_cond $X=2.31 $Y=1.557
+ $X2=2.355 $Y2=1.557
r146 62 64 32.1333 $w=3.75e-07 $l=2.5e-07 $layer=POLY_cond $X=2.06 $Y=1.557
+ $X2=2.31 $Y2=1.557
r147 62 63 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=2.06
+ $Y=1.515 $X2=2.06 $Y2=1.515
r148 60 62 19.9227 $w=3.75e-07 $l=1.55e-07 $layer=POLY_cond $X=1.905 $Y=1.557
+ $X2=2.06 $Y2=1.557
r149 59 60 12.2107 $w=3.75e-07 $l=9.5e-08 $layer=POLY_cond $X=1.81 $Y=1.557
+ $X2=1.905 $Y2=1.557
r150 53 71 4.82418 $w=4.28e-07 $l=1.8e-07 $layer=LI1_cond $X=3.6 $Y=1.565
+ $X2=3.42 $Y2=1.565
r151 52 71 8.0403 $w=4.28e-07 $l=3e-07 $layer=LI1_cond $X=3.12 $Y=1.565 $X2=3.42
+ $Y2=1.565
r152 51 52 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=2.64 $Y=1.565
+ $X2=3.12 $Y2=1.565
r153 50 51 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=2.16 $Y=1.565
+ $X2=2.64 $Y2=1.565
r154 50 63 2.6801 $w=4.28e-07 $l=1e-07 $layer=LI1_cond $X=2.16 $Y=1.565 $X2=2.06
+ $Y2=1.565
r155 49 63 10.1844 $w=4.28e-07 $l=3.8e-07 $layer=LI1_cond $X=1.68 $Y=1.565
+ $X2=2.06 $Y2=1.565
r156 44 72 18.6373 $w=3.75e-07 $l=2.70969e-07 $layer=POLY_cond $X=3.855 $Y=1.765
+ $X2=3.71 $Y2=1.557
r157 44 46 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.855 $Y=1.765
+ $X2=3.855 $Y2=2.4
r158 40 72 24.2915 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.71 $Y=1.35
+ $X2=3.71 $Y2=1.557
r159 40 42 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.71 $Y=1.35
+ $X2=3.71 $Y2=0.74
r160 37 68 24.2915 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.305 $Y=1.765
+ $X2=3.305 $Y2=1.557
r161 37 39 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.305 $Y=1.765
+ $X2=3.305 $Y2=2.4
r162 33 67 24.2915 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.21 $Y=1.35
+ $X2=3.21 $Y2=1.557
r163 33 35 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.21 $Y=1.35
+ $X2=3.21 $Y2=0.74
r164 30 66 24.2915 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.855 $Y=1.765
+ $X2=2.855 $Y2=1.557
r165 30 32 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.855 $Y=1.765
+ $X2=2.855 $Y2=2.4
r166 27 65 24.2915 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.355 $Y=1.765
+ $X2=2.355 $Y2=1.557
r167 27 29 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.355 $Y=1.765
+ $X2=2.355 $Y2=2.4
r168 23 64 24.2915 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.31 $Y=1.35
+ $X2=2.31 $Y2=1.557
r169 23 25 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.31 $Y=1.35
+ $X2=2.31 $Y2=0.74
r170 20 60 24.2915 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.905 $Y=1.765
+ $X2=1.905 $Y2=1.557
r171 20 22 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.905 $Y=1.765
+ $X2=1.905 $Y2=2.4
r172 16 59 24.2915 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.81 $Y=1.35
+ $X2=1.81 $Y2=1.557
r173 16 18 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.81 $Y=1.35
+ $X2=1.81 $Y2=0.74
r174 15 48 20.4101 $w=1.5e-07 $l=9.94987e-08 $layer=POLY_cond $X=1.545 $Y=1.65
+ $X2=1.455 $Y2=1.67
r175 14 59 27.567 $w=3.75e-07 $l=1.24996e-07 $layer=POLY_cond $X=1.735 $Y=1.65
+ $X2=1.81 $Y2=1.557
r176 14 15 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=1.735 $Y=1.65
+ $X2=1.545 $Y2=1.65
r177 11 48 5.30422 $w=1.5e-07 $l=9.5e-08 $layer=POLY_cond $X=1.455 $Y=1.765
+ $X2=1.455 $Y2=1.67
r178 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.455 $Y=1.765
+ $X2=1.455 $Y2=2.4
r179 10 47 20.4101 $w=1.5e-07 $l=9.94987e-08 $layer=POLY_cond $X=1.095 $Y=1.65
+ $X2=1.005 $Y2=1.67
r180 9 48 20.4101 $w=1.5e-07 $l=9.94987e-08 $layer=POLY_cond $X=1.365 $Y=1.65
+ $X2=1.455 $Y2=1.67
r181 9 10 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=1.365 $Y=1.65
+ $X2=1.095 $Y2=1.65
r182 6 47 5.30422 $w=1.5e-07 $l=9.5e-08 $layer=POLY_cond $X=1.005 $Y=1.765
+ $X2=1.005 $Y2=1.67
r183 6 8 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.005 $Y=1.765
+ $X2=1.005 $Y2=2.4
r184 4 47 20.4101 $w=1.5e-07 $l=9.94987e-08 $layer=POLY_cond $X=0.915 $Y=1.65
+ $X2=1.005 $Y2=1.67
r185 4 5 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.915 $Y=1.65
+ $X2=0.595 $Y2=1.65
r186 1 5 26.9307 $w=1.5e-07 $l=1.53542e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.595 $Y2=1.65
r187 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__NOR2_8%B 1 3 5 6 8 9 12 13 15 16 19 20 22 23 25 26
+ 29 30 32 33 35 37 38 40 41 43 44 45 47 48 50 51 54 55 57 59 60 62 63 64 65 70
+ 72 74 75 79 80
c154 38 0 4.12053e-20 $X=6.205 $Y=1.765
r155 83 84 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=7.39
+ $Y=1.145 $X2=7.39 $Y2=1.145
r156 79 83 57.7492 $w=6.3e-07 $l=6.8e-07 $layer=POLY_cond $X=7.38 $Y=0.465
+ $X2=7.38 $Y2=1.145
r157 79 80 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=7.39
+ $Y=0.465 $X2=7.39 $Y2=0.465
r158 75 84 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=7.39 $Y=0.925
+ $X2=7.39 $Y2=1.145
r159 74 75 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=7.39 $Y=0.555
+ $X2=7.39 $Y2=0.925
r160 74 80 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=7.39 $Y=0.555
+ $X2=7.39 $Y2=0.465
r161 71 83 3.39701 $w=6.3e-07 $l=4e-08 $layer=POLY_cond $X=7.38 $Y=1.185
+ $X2=7.38 $Y2=1.145
r162 71 72 6.3694 $w=6.3e-07 $l=7.5e-08 $layer=POLY_cond $X=7.38 $Y=1.185
+ $X2=7.38 $Y2=1.26
r163 60 62 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.605 $Y=1.765
+ $X2=7.605 $Y2=2.4
r164 59 60 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=7.605 $Y=1.675
+ $X2=7.605 $Y2=1.765
r165 55 57 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.155 $Y=1.765
+ $X2=7.155 $Y2=2.4
r166 54 55 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=7.155 $Y=1.675
+ $X2=7.155 $Y2=1.765
r167 53 72 36.8168 $w=6.3e-07 $l=7.5e-08 $layer=POLY_cond $X=7.38 $Y=1.335
+ $X2=7.38 $Y2=1.26
r168 53 59 132.161 $w=1.8e-07 $l=3.4e-07 $layer=POLY_cond $X=7.605 $Y=1.335
+ $X2=7.605 $Y2=1.675
r169 53 54 132.161 $w=1.8e-07 $l=3.4e-07 $layer=POLY_cond $X=7.155 $Y=1.335
+ $X2=7.155 $Y2=1.675
r170 52 70 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=6.745 $Y=1.26
+ $X2=6.655 $Y2=1.26
r171 51 72 37.3437 $w=1.5e-07 $l=3.15e-07 $layer=POLY_cond $X=7.065 $Y=1.26
+ $X2=7.38 $Y2=1.26
r172 51 52 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=7.065 $Y=1.26
+ $X2=6.745 $Y2=1.26
r173 48 50 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.655 $Y=1.765
+ $X2=6.655 $Y2=2.4
r174 47 48 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.655 $Y=1.675
+ $X2=6.655 $Y2=1.765
r175 46 70 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=6.655 $Y=1.335
+ $X2=6.655 $Y2=1.26
r176 46 47 132.161 $w=1.8e-07 $l=3.4e-07 $layer=POLY_cond $X=6.655 $Y=1.335
+ $X2=6.655 $Y2=1.675
r177 45 69 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.4 $Y=1.26
+ $X2=6.325 $Y2=1.26
r178 44 70 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=6.565 $Y=1.26
+ $X2=6.655 $Y2=1.26
r179 44 45 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.565 $Y=1.26
+ $X2=6.4 $Y2=1.26
r180 41 69 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.325 $Y=1.185
+ $X2=6.325 $Y2=1.26
r181 41 43 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=6.325 $Y=1.185
+ $X2=6.325 $Y2=0.74
r182 38 40 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.205 $Y=1.765
+ $X2=6.205 $Y2=2.4
r183 37 38 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.205 $Y=1.675
+ $X2=6.205 $Y2=1.765
r184 36 69 61.5319 $w=1.5e-07 $l=1.2e-07 $layer=POLY_cond $X=6.205 $Y=1.26
+ $X2=6.325 $Y2=1.26
r185 36 67 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=6.205 $Y=1.26
+ $X2=5.895 $Y2=1.26
r186 36 37 132.161 $w=1.8e-07 $l=3.4e-07 $layer=POLY_cond $X=6.205 $Y=1.335
+ $X2=6.205 $Y2=1.675
r187 33 67 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.895 $Y=1.185
+ $X2=5.895 $Y2=1.26
r188 33 35 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=5.895 $Y=1.185
+ $X2=5.895 $Y2=0.74
r189 30 32 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.755 $Y=1.765
+ $X2=5.755 $Y2=2.4
r190 29 30 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.755 $Y=1.675
+ $X2=5.755 $Y2=1.765
r191 28 67 71.7872 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=5.755 $Y=1.26
+ $X2=5.895 $Y2=1.26
r192 28 29 132.161 $w=1.8e-07 $l=3.4e-07 $layer=POLY_cond $X=5.755 $Y=1.335
+ $X2=5.755 $Y2=1.675
r193 27 65 13.2179 $w=1.5e-07 $l=9.3e-08 $layer=POLY_cond $X=5.4 $Y=1.26
+ $X2=5.307 $Y2=1.26
r194 26 28 46.1489 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=5.665 $Y=1.26
+ $X2=5.755 $Y2=1.26
r195 26 27 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=5.665 $Y=1.26
+ $X2=5.4 $Y2=1.26
r196 23 65 10.9219 $w=1.5e-07 $l=8.35165e-08 $layer=POLY_cond $X=5.325 $Y=1.185
+ $X2=5.307 $Y2=1.26
r197 23 25 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=5.325 $Y=1.185
+ $X2=5.325 $Y2=0.74
r198 20 22 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.305 $Y=1.765
+ $X2=5.305 $Y2=2.4
r199 19 20 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.305 $Y=1.675
+ $X2=5.305 $Y2=1.765
r200 18 65 10.9219 $w=1.8e-07 $l=7.59934e-08 $layer=POLY_cond $X=5.305 $Y=1.335
+ $X2=5.307 $Y2=1.26
r201 18 19 132.161 $w=1.8e-07 $l=3.4e-07 $layer=POLY_cond $X=5.305 $Y=1.335
+ $X2=5.305 $Y2=1.675
r202 17 64 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.895 $Y=1.26
+ $X2=4.805 $Y2=1.26
r203 16 65 13.2179 $w=1.5e-07 $l=9.2e-08 $layer=POLY_cond $X=5.215 $Y=1.26
+ $X2=5.307 $Y2=1.26
r204 16 17 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=5.215 $Y=1.26
+ $X2=4.895 $Y2=1.26
r205 13 15 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.805 $Y=1.765
+ $X2=4.805 $Y2=2.4
r206 12 13 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=4.805 $Y=1.675
+ $X2=4.805 $Y2=1.765
r207 11 64 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=4.805 $Y=1.335
+ $X2=4.805 $Y2=1.26
r208 11 12 132.161 $w=1.8e-07 $l=3.4e-07 $layer=POLY_cond $X=4.805 $Y=1.335
+ $X2=4.805 $Y2=1.675
r209 10 63 6.66866 $w=1.5e-07 $l=1.3e-07 $layer=POLY_cond $X=4.395 $Y=1.26
+ $X2=4.265 $Y2=1.26
r210 9 64 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.715 $Y=1.26
+ $X2=4.805 $Y2=1.26
r211 9 10 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.715 $Y=1.26
+ $X2=4.395 $Y2=1.26
r212 6 8 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.305 $Y=1.765
+ $X2=4.305 $Y2=2.4
r213 5 6 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=4.305 $Y=1.675
+ $X2=4.305 $Y2=1.765
r214 4 63 18.8402 $w=1.65e-07 $l=9.28709e-08 $layer=POLY_cond $X=4.305 $Y=1.335
+ $X2=4.265 $Y2=1.26
r215 4 5 132.161 $w=1.8e-07 $l=3.4e-07 $layer=POLY_cond $X=4.305 $Y=1.335
+ $X2=4.305 $Y2=1.675
r216 1 63 18.8402 $w=1.65e-07 $l=9.87421e-08 $layer=POLY_cond $X=4.21 $Y=1.185
+ $X2=4.265 $Y2=1.26
r217 1 3 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=4.21 $Y=1.185
+ $X2=4.21 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__NOR2_8%A_27_368# 1 2 3 4 5 6 7 8 9 30 34 35 38 40 44
+ 46 50 52 54 57 58 59 62 66 70 74 78 82 86 90 95 97 100 101 102
r139 90 93 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.23 $Y=1.865
+ $X2=1.23 $Y2=2.035
r140 86 89 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=7.88 $Y=1.985
+ $X2=7.88 $Y2=2.815
r141 84 89 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=7.88 $Y=2.905
+ $X2=7.88 $Y2=2.815
r142 83 102 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=7.035 $Y=2.99
+ $X2=6.905 $Y2=2.99
r143 82 84 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.715 $Y=2.99
+ $X2=7.88 $Y2=2.905
r144 82 83 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=7.715 $Y=2.99
+ $X2=7.035 $Y2=2.99
r145 78 81 36.7895 $w=2.58e-07 $l=8.3e-07 $layer=LI1_cond $X=6.905 $Y=1.985
+ $X2=6.905 $Y2=2.815
r146 76 102 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=6.905 $Y=2.905
+ $X2=6.905 $Y2=2.99
r147 76 81 3.98923 $w=2.58e-07 $l=9e-08 $layer=LI1_cond $X=6.905 $Y=2.905
+ $X2=6.905 $Y2=2.815
r148 75 101 6.01921 $w=1.7e-07 $l=1.03e-07 $layer=LI1_cond $X=6.08 $Y=2.99
+ $X2=5.977 $Y2=2.99
r149 74 102 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.775 $Y=2.99
+ $X2=6.905 $Y2=2.99
r150 74 75 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=6.775 $Y=2.99
+ $X2=6.08 $Y2=2.99
r151 70 73 44.9047 $w=2.03e-07 $l=8.3e-07 $layer=LI1_cond $X=5.977 $Y=1.985
+ $X2=5.977 $Y2=2.815
r152 68 101 0.677923 $w=2.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.977 $Y=2.905
+ $X2=5.977 $Y2=2.99
r153 68 73 4.86918 $w=2.03e-07 $l=9e-08 $layer=LI1_cond $X=5.977 $Y=2.905
+ $X2=5.977 $Y2=2.815
r154 67 100 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.185 $Y=2.99
+ $X2=5.055 $Y2=2.99
r155 66 101 6.01921 $w=1.7e-07 $l=1.02e-07 $layer=LI1_cond $X=5.875 $Y=2.99
+ $X2=5.977 $Y2=2.99
r156 66 67 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.875 $Y=2.99
+ $X2=5.185 $Y2=2.99
r157 62 65 31.0273 $w=2.58e-07 $l=7e-07 $layer=LI1_cond $X=5.055 $Y=2.115
+ $X2=5.055 $Y2=2.815
r158 60 100 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=5.055 $Y=2.905
+ $X2=5.055 $Y2=2.99
r159 60 65 3.98923 $w=2.58e-07 $l=9e-08 $layer=LI1_cond $X=5.055 $Y=2.905
+ $X2=5.055 $Y2=2.815
r160 58 100 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.925 $Y=2.99
+ $X2=5.055 $Y2=2.99
r161 58 59 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.925 $Y=2.99
+ $X2=4.245 $Y2=2.99
r162 55 59 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.08 $Y=2.905
+ $X2=4.245 $Y2=2.99
r163 55 57 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=4.08 $Y=2.905
+ $X2=4.08 $Y2=2.815
r164 54 99 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.08 $Y=2.12 $X2=4.08
+ $Y2=2.035
r165 54 57 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=4.08 $Y=2.12
+ $X2=4.08 $Y2=2.815
r166 53 97 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.245 $Y=2.035
+ $X2=3.12 $Y2=2.035
r167 52 99 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.915 $Y=2.035
+ $X2=4.08 $Y2=2.035
r168 52 53 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.915 $Y=2.035
+ $X2=3.245 $Y2=2.035
r169 48 97 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.12 $Y=2.12
+ $X2=3.12 $Y2=2.035
r170 48 50 14.5208 $w=2.48e-07 $l=3.15e-07 $layer=LI1_cond $X=3.12 $Y=2.12
+ $X2=3.12 $Y2=2.435
r171 47 95 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.295 $Y=2.035
+ $X2=2.17 $Y2=2.035
r172 46 97 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.995 $Y=2.035
+ $X2=3.12 $Y2=2.035
r173 46 47 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=2.995 $Y=2.035
+ $X2=2.295 $Y2=2.035
r174 42 95 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.17 $Y=2.12
+ $X2=2.17 $Y2=2.035
r175 42 44 14.5208 $w=2.48e-07 $l=3.15e-07 $layer=LI1_cond $X=2.17 $Y=2.12
+ $X2=2.17 $Y2=2.435
r176 41 93 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.315 $Y=2.035
+ $X2=1.23 $Y2=2.035
r177 40 95 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.045 $Y=2.035
+ $X2=2.17 $Y2=2.035
r178 40 41 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=2.045 $Y=2.035
+ $X2=1.315 $Y2=2.035
r179 36 93 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.23 $Y=2.12
+ $X2=1.23 $Y2=2.035
r180 36 38 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.23 $Y=2.12
+ $X2=1.23 $Y2=2.435
r181 34 90 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.145 $Y=1.865
+ $X2=1.23 $Y2=1.865
r182 34 35 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.145 $Y=1.865
+ $X2=0.445 $Y2=1.865
r183 30 32 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=0.28 $Y=1.985
+ $X2=0.28 $Y2=2.815
r184 28 35 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=1.95
+ $X2=0.445 $Y2=1.865
r185 28 30 1.22229 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=0.28 $Y=1.95
+ $X2=0.28 $Y2=1.985
r186 9 89 400 $w=1.7e-07 $l=1.07034e-06 $layer=licon1_PDIFF $count=1 $X=7.68
+ $Y=1.84 $X2=7.88 $Y2=2.815
r187 9 86 400 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=1 $X=7.68
+ $Y=1.84 $X2=7.88 $Y2=1.985
r188 8 81 400 $w=1.7e-07 $l=1.07034e-06 $layer=licon1_PDIFF $count=1 $X=6.73
+ $Y=1.84 $X2=6.93 $Y2=2.815
r189 8 78 400 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=1 $X=6.73
+ $Y=1.84 $X2=6.93 $Y2=1.985
r190 7 73 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=5.83
+ $Y=1.84 $X2=5.98 $Y2=2.815
r191 7 70 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=5.83
+ $Y=1.84 $X2=5.98 $Y2=1.985
r192 6 65 400 $w=1.7e-07 $l=1.07034e-06 $layer=licon1_PDIFF $count=1 $X=4.88
+ $Y=1.84 $X2=5.08 $Y2=2.815
r193 6 62 400 $w=1.7e-07 $l=3.61421e-07 $layer=licon1_PDIFF $count=1 $X=4.88
+ $Y=1.84 $X2=5.08 $Y2=2.115
r194 5 99 400 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=3.93
+ $Y=1.84 $X2=4.08 $Y2=2.035
r195 5 57 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=3.93
+ $Y=1.84 $X2=4.08 $Y2=2.815
r196 4 97 600 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=2.93
+ $Y=1.84 $X2=3.08 $Y2=2.035
r197 4 50 300 $w=1.7e-07 $l=6.65789e-07 $layer=licon1_PDIFF $count=2 $X=2.93
+ $Y=1.84 $X2=3.08 $Y2=2.435
r198 3 95 600 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=1.98
+ $Y=1.84 $X2=2.13 $Y2=2.035
r199 3 44 300 $w=1.7e-07 $l=6.65789e-07 $layer=licon1_PDIFF $count=2 $X=1.98
+ $Y=1.84 $X2=2.13 $Y2=2.435
r200 2 93 600 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=1.08
+ $Y=1.84 $X2=1.23 $Y2=2.035
r201 2 38 300 $w=1.7e-07 $l=6.65789e-07 $layer=licon1_PDIFF $count=2 $X=1.08
+ $Y=1.84 $X2=1.23 $Y2=2.435
r202 1 32 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r203 1 30 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_LS__NOR2_8%VPWR 1 2 3 4 15 19 23 27 29 31 36 41 46 56 57
+ 60 63 66 69
r99 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r100 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r101 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r102 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r103 56 57 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r104 53 56 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=4.08 $Y=3.33
+ $X2=7.92 $Y2=3.33
r105 51 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.745 $Y=3.33
+ $X2=3.58 $Y2=3.33
r106 51 53 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=3.745 $Y=3.33
+ $X2=4.08 $Y2=3.33
r107 50 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r108 50 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r109 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r110 47 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.795 $Y=3.33
+ $X2=2.63 $Y2=3.33
r111 47 49 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.795 $Y=3.33
+ $X2=3.12 $Y2=3.33
r112 46 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.415 $Y=3.33
+ $X2=3.58 $Y2=3.33
r113 46 49 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.415 $Y=3.33
+ $X2=3.12 $Y2=3.33
r114 45 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r115 45 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r116 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r117 42 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.845 $Y=3.33
+ $X2=1.68 $Y2=3.33
r118 42 44 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.845 $Y=3.33
+ $X2=2.16 $Y2=3.33
r119 41 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.465 $Y=3.33
+ $X2=2.63 $Y2=3.33
r120 41 44 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.465 $Y=3.33
+ $X2=2.16 $Y2=3.33
r121 40 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r122 40 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r123 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r124 37 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=0.78 $Y2=3.33
r125 37 39 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=1.2 $Y2=3.33
r126 36 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.515 $Y=3.33
+ $X2=1.68 $Y2=3.33
r127 36 39 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.515 $Y=3.33
+ $X2=1.2 $Y2=3.33
r128 34 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r129 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r130 31 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.78 $Y2=3.33
r131 31 33 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.24 $Y2=3.33
r132 29 57 1.07034 $w=4.9e-07 $l=3.84e-06 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=7.92 $Y2=3.33
r133 29 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r134 29 53 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r135 25 69 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.58 $Y=3.245
+ $X2=3.58 $Y2=3.33
r136 25 27 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=3.58 $Y=3.245
+ $X2=3.58 $Y2=2.455
r137 21 66 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.63 $Y=3.245
+ $X2=2.63 $Y2=3.33
r138 21 23 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=2.63 $Y=3.245
+ $X2=2.63 $Y2=2.455
r139 17 63 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.68 $Y=3.245
+ $X2=1.68 $Y2=3.33
r140 17 19 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=1.68 $Y=3.245
+ $X2=1.68 $Y2=2.455
r141 13 60 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=3.245
+ $X2=0.78 $Y2=3.33
r142 13 15 33.5256 $w=3.28e-07 $l=9.6e-07 $layer=LI1_cond $X=0.78 $Y=3.245
+ $X2=0.78 $Y2=2.285
r143 4 27 300 $w=1.7e-07 $l=7.07972e-07 $layer=licon1_PDIFF $count=2 $X=3.38
+ $Y=1.84 $X2=3.58 $Y2=2.455
r144 3 23 300 $w=1.7e-07 $l=7.07972e-07 $layer=licon1_PDIFF $count=2 $X=2.43
+ $Y=1.84 $X2=2.63 $Y2=2.455
r145 2 19 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=1.53
+ $Y=1.84 $X2=1.68 $Y2=2.455
r146 1 15 300 $w=1.7e-07 $l=5.35747e-07 $layer=licon1_PDIFF $count=2 $X=0.58
+ $Y=1.84 $X2=0.78 $Y2=2.285
.ends

.subckt PM_SKY130_FD_SC_LS__NOR2_8%Y 1 2 3 4 5 6 7 8 27 29 30 33 35 39 45 51 55
+ 59 60 63 67 68 73
c120 60 0 4.12053e-20 $X=6.595 $Y=1.565
r121 76 77 5.99298 $w=8.55e-07 $l=4.2e-07 $layer=LI1_cond $X=5.11 $Y=1.14
+ $X2=5.53 $Y2=1.14
r122 74 76 7.56257 $w=8.55e-07 $l=5.3e-07 $layer=LI1_cond $X=4.58 $Y=1.14
+ $X2=5.11 $Y2=1.14
r123 73 74 0.28538 $w=8.55e-07 $l=2e-08 $layer=LI1_cond $X=4.56 $Y=1.14 $X2=4.58
+ $Y2=1.14
r124 71 73 1.92632 $w=8.55e-07 $l=1.35e-07 $layer=LI1_cond $X=4.425 $Y=1.14
+ $X2=4.56 $Y2=1.14
r125 68 73 10.6563 $w=1.7e-07 $l=5.25e-07 $layer=LI1_cond $X=4.56 $Y=1.665
+ $X2=4.56 $Y2=1.14
r126 63 65 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=7.38 $Y=1.97
+ $X2=7.38 $Y2=2.65
r127 61 63 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=7.38 $Y=1.65
+ $X2=7.38 $Y2=1.97
r128 59 61 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.215 $Y=1.565
+ $X2=7.38 $Y2=1.65
r129 59 60 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=7.215 $Y=1.565
+ $X2=6.595 $Y2=1.565
r130 55 57 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=6.43 $Y=1.97
+ $X2=6.43 $Y2=2.65
r131 53 60 12.0026 $w=8.55e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.43 $Y=1.65
+ $X2=6.595 $Y2=1.565
r132 53 55 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=6.43 $Y=1.65
+ $X2=6.43 $Y2=1.97
r133 49 53 4.56608 $w=8.55e-07 $l=6.50615e-07 $layer=LI1_cond $X=6.11 $Y=1.14
+ $X2=6.43 $Y2=1.65
r134 49 77 8.27602 $w=8.55e-07 $l=5.8e-07 $layer=LI1_cond $X=6.11 $Y=1.14
+ $X2=5.53 $Y2=1.14
r135 49 51 21.8266 $w=3.28e-07 $l=6.25e-07 $layer=LI1_cond $X=6.11 $Y=1.14
+ $X2=6.11 $Y2=0.515
r136 45 47 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=5.53 $Y=1.97
+ $X2=5.53 $Y2=2.65
r137 43 77 6.368 $w=3.3e-07 $l=6.4e-07 $layer=LI1_cond $X=5.53 $Y=1.78 $X2=5.53
+ $Y2=1.14
r138 43 45 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=5.53 $Y=1.78
+ $X2=5.53 $Y2=1.97
r139 39 41 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=4.58 $Y=1.97
+ $X2=4.58 $Y2=2.65
r140 37 74 6.368 $w=3.3e-07 $l=6.4e-07 $layer=LI1_cond $X=4.58 $Y=1.78 $X2=4.58
+ $Y2=1.14
r141 37 39 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=4.58 $Y=1.78
+ $X2=4.58 $Y2=1.97
r142 36 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.59 $Y=1.095
+ $X2=3.425 $Y2=1.095
r143 35 71 12.0026 $w=8.55e-07 $l=1.86145e-07 $layer=LI1_cond $X=4.26 $Y=1.095
+ $X2=4.425 $Y2=1.14
r144 35 36 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.26 $Y=1.095
+ $X2=3.59 $Y2=1.095
r145 31 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.425 $Y=1.01
+ $X2=3.425 $Y2=1.095
r146 31 33 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=3.425 $Y=1.01
+ $X2=3.425 $Y2=0.515
r147 29 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.26 $Y=1.095
+ $X2=3.425 $Y2=1.095
r148 29 30 69.8075 $w=1.68e-07 $l=1.07e-06 $layer=LI1_cond $X=3.26 $Y=1.095
+ $X2=2.19 $Y2=1.095
r149 25 30 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.025 $Y=1.01
+ $X2=2.19 $Y2=1.095
r150 25 27 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=2.025 $Y=1.01
+ $X2=2.025 $Y2=0.515
r151 8 65 400 $w=1.7e-07 $l=8.81816e-07 $layer=licon1_PDIFF $count=1 $X=7.23
+ $Y=1.84 $X2=7.38 $Y2=2.65
r152 8 63 400 $w=1.7e-07 $l=2.04939e-07 $layer=licon1_PDIFF $count=1 $X=7.23
+ $Y=1.84 $X2=7.38 $Y2=1.97
r153 7 57 400 $w=1.7e-07 $l=8.81816e-07 $layer=licon1_PDIFF $count=1 $X=6.28
+ $Y=1.84 $X2=6.43 $Y2=2.65
r154 7 55 400 $w=1.7e-07 $l=2.04939e-07 $layer=licon1_PDIFF $count=1 $X=6.28
+ $Y=1.84 $X2=6.43 $Y2=1.97
r155 6 47 400 $w=1.7e-07 $l=8.81816e-07 $layer=licon1_PDIFF $count=1 $X=5.38
+ $Y=1.84 $X2=5.53 $Y2=2.65
r156 6 45 400 $w=1.7e-07 $l=2.04939e-07 $layer=licon1_PDIFF $count=1 $X=5.38
+ $Y=1.84 $X2=5.53 $Y2=1.97
r157 5 41 400 $w=1.7e-07 $l=9.04489e-07 $layer=licon1_PDIFF $count=1 $X=4.38
+ $Y=1.84 $X2=4.58 $Y2=2.65
r158 5 39 400 $w=1.7e-07 $l=2.56905e-07 $layer=licon1_PDIFF $count=1 $X=4.38
+ $Y=1.84 $X2=4.58 $Y2=1.97
r159 4 51 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.97
+ $Y=0.37 $X2=6.11 $Y2=0.515
r160 3 76 60.6667 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_NDIFF $count=3
+ $X=4.285 $Y=0.37 $X2=5.11 $Y2=0.515
r161 3 71 60.6667 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=3
+ $X=4.285 $Y=0.37 $X2=4.425 $Y2=0.515
r162 2 33 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.285
+ $Y=0.37 $X2=3.425 $Y2=0.515
r163 1 27 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.885
+ $Y=0.37 $X2=2.025 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__NOR2_8%VGND 1 2 3 4 5 20 25 29 31 35 37 41 43 45 50
+ 60 61 64 69 72 75 78
r78 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r79 76 79 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6.48
+ $Y2=0
r80 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r81 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r82 65 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r83 64 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r84 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r85 60 61 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r86 58 61 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.92
+ $Y2=0
r87 58 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=6.48
+ $Y2=0
r88 57 60 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=6.96 $Y=0 $X2=7.92
+ $Y2=0
r89 57 58 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r90 55 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.775 $Y=0 $X2=6.61
+ $Y2=0
r91 55 57 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=6.775 $Y=0 $X2=6.96
+ $Y2=0
r92 54 70 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=2.64
+ $Y2=0
r93 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r94 51 69 13.9655 $w=1.7e-07 $l=3.65e-07 $layer=LI1_cond $X=3.09 $Y=0 $X2=2.725
+ $Y2=0
r95 51 53 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=3.09 $Y=0 $X2=3.6
+ $Y2=0
r96 50 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.76 $Y=0 $X2=3.925
+ $Y2=0
r97 50 53 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=3.76 $Y=0 $X2=3.6
+ $Y2=0
r98 49 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r99 49 65 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.2
+ $Y2=0
r100 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r101 46 64 16.5844 $w=1.7e-07 $l=5.2e-07 $layer=LI1_cond $X=1.69 $Y=0 $X2=1.17
+ $Y2=0
r102 46 48 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=1.69 $Y=0 $X2=2.16
+ $Y2=0
r103 45 69 13.9655 $w=1.7e-07 $l=3.65e-07 $layer=LI1_cond $X=2.36 $Y=0 $X2=2.725
+ $Y2=0
r104 45 48 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=2.36 $Y=0 $X2=2.16
+ $Y2=0
r105 43 76 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.08 $Y=0
+ $X2=5.52 $Y2=0
r106 43 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r107 43 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r108 39 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.61 $Y=0.085
+ $X2=6.61 $Y2=0
r109 39 41 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=6.61 $Y=0.085
+ $X2=6.61 $Y2=0.515
r110 38 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.775 $Y=0 $X2=5.61
+ $Y2=0
r111 37 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.445 $Y=0 $X2=6.61
+ $Y2=0
r112 37 38 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.445 $Y=0
+ $X2=5.775 $Y2=0
r113 33 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.61 $Y=0.085
+ $X2=5.61 $Y2=0
r114 33 35 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=5.61 $Y=0.085
+ $X2=5.61 $Y2=0.515
r115 32 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.09 $Y=0 $X2=3.925
+ $Y2=0
r116 31 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.445 $Y=0 $X2=5.61
+ $Y2=0
r117 31 32 88.4011 $w=1.68e-07 $l=1.355e-06 $layer=LI1_cond $X=5.445 $Y=0
+ $X2=4.09 $Y2=0
r118 27 72 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.925 $Y=0.085
+ $X2=3.925 $Y2=0
r119 27 29 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=3.925 $Y=0.085
+ $X2=3.925 $Y2=0.675
r120 23 69 2.94957 $w=7.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.725 $Y=0.085
+ $X2=2.725 $Y2=0
r121 23 25 9.66693 $w=7.28e-07 $l=5.9e-07 $layer=LI1_cond $X=2.725 $Y=0.085
+ $X2=2.725 $Y2=0.675
r122 18 64 3.59326 $w=1.04e-06 $l=8.5e-08 $layer=LI1_cond $X=1.17 $Y=0.085
+ $X2=1.17 $Y2=0
r123 18 20 5.04423 $w=1.038e-06 $l=4.3e-07 $layer=LI1_cond $X=1.17 $Y=0.085
+ $X2=1.17 $Y2=0.515
r124 5 41 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=6.4
+ $Y=0.37 $X2=6.61 $Y2=0.515
r125 4 35 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=5.4
+ $Y=0.37 $X2=5.61 $Y2=0.515
r126 3 29 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=3.785
+ $Y=0.37 $X2=3.925 $Y2=0.675
r127 2 25 91 $w=1.7e-07 $l=7.47094e-07 $layer=licon1_NDIFF $count=2 $X=2.385
+ $Y=0.37 $X2=2.995 $Y2=0.675
r128 1 20 60.6667 $w=1.7e-07 $l=9.94862e-07 $layer=licon1_NDIFF $count=3 $X=0.67
+ $Y=0.37 $X2=1.595 $Y2=0.515
r129 1 20 60.6667 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_NDIFF $count=3 $X=0.67
+ $Y=0.37 $X2=0.885 $Y2=0.515
.ends

