# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ls__o41a_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ls__o41a_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.160000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.528000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.330000 1.420000 7.075000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.528000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.305000 0.255000 7.635000 0.335000 ;
        RECT 7.305000 0.335000 8.035000 0.505000 ;
        RECT 7.805000 0.505000 8.035000 0.670000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.528000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.875000 0.255000 4.205000 0.670000 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.528000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445000 1.425000 5.180000 1.780000 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.444000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.280000 1.440000 4.195000 1.780000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  1.086400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.930000 1.855000 1.100000 ;
        RECT 0.125000 1.100000 0.295000 1.770000 ;
        RECT 0.125000 1.770000 2.125000 1.940000 ;
        RECT 0.125000 1.940000 0.355000 2.890000 ;
        RECT 0.675000 0.350000 0.925000 0.930000 ;
        RECT 0.895000 1.940000 1.225000 2.980000 ;
        RECT 1.605000 0.350000 1.855000 0.930000 ;
        RECT 1.795000 1.940000 2.125000 2.980000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.160000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.160000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.160000 0.085000 ;
      RECT 0.000000  3.245000 8.160000 3.415000 ;
      RECT 0.175000  0.085000 0.505000 0.760000 ;
      RECT 0.525000  2.110000 0.695000 3.245000 ;
      RECT 0.585000  1.270000 3.110000 1.600000 ;
      RECT 1.105000  0.085000 1.435000 0.760000 ;
      RECT 1.425000  2.110000 1.595000 3.245000 ;
      RECT 2.035000  0.085000 2.365000 1.100000 ;
      RECT 2.325000  1.910000 2.575000 3.245000 ;
      RECT 2.595000  0.260000 3.705000 0.430000 ;
      RECT 2.595000  0.430000 2.925000 0.930000 ;
      RECT 2.780000  1.600000 3.110000 1.950000 ;
      RECT 2.780000  1.950000 5.030000 2.120000 ;
      RECT 2.780000  2.120000 3.110000 2.790000 ;
      RECT 2.940000  1.100000 3.275000 1.270000 ;
      RECT 3.105000  0.600000 3.275000 1.100000 ;
      RECT 3.310000  2.290000 3.560000 3.245000 ;
      RECT 3.455000  0.430000 3.705000 1.085000 ;
      RECT 3.455000  1.085000 7.635000 1.250000 ;
      RECT 3.455000  1.250000 5.845000 1.255000 ;
      RECT 3.455000  1.255000 3.705000 1.270000 ;
      RECT 3.790000  2.290000 5.850000 2.460000 ;
      RECT 3.790000  2.460000 4.040000 2.980000 ;
      RECT 4.240000  2.630000 5.480000 2.980000 ;
      RECT 4.375000  0.085000 4.545000 0.915000 ;
      RECT 4.725000  0.580000 4.975000 1.085000 ;
      RECT 5.155000  0.085000 5.485000 0.915000 ;
      RECT 5.665000  0.580000 5.845000 1.080000 ;
      RECT 5.665000  1.080000 7.635000 1.085000 ;
      RECT 5.680000  1.820000 5.850000 1.950000 ;
      RECT 5.680000  1.950000 7.870000 2.120000 ;
      RECT 5.680000  2.120000 5.850000 2.290000 ;
      RECT 5.680000  2.460000 5.850000 2.980000 ;
      RECT 6.025000  0.085000 6.275000 0.910000 ;
      RECT 6.050000  2.290000 7.370000 2.460000 ;
      RECT 6.050000  2.460000 6.380000 2.980000 ;
      RECT 6.455000  0.580000 6.705000 1.080000 ;
      RECT 6.580000  2.650000 6.870000 3.245000 ;
      RECT 6.885000  0.085000 7.135000 0.910000 ;
      RECT 7.040000  2.460000 7.370000 2.980000 ;
      RECT 7.385000  0.675000 7.635000 1.080000 ;
      RECT 7.385000  1.250000 7.635000 1.275000 ;
      RECT 7.540000  1.820000 7.870000 1.950000 ;
      RECT 7.540000  2.120000 7.870000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
  END
END sky130_fd_sc_ls__o41a_4
