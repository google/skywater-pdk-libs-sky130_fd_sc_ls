* File: sky130_fd_sc_ls__clkdlyinv5sd1_1.spice
* Created: Wed Sep  2 10:58:15 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__clkdlyinv5sd1_1.pex.spice"
.subckt sky130_fd_sc_ls__clkdlyinv5sd1_1  VNB VPB A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1006 N_VGND_M1006_d N_A_M1006_g N_A_28_74#_M1006_s VNB NSHORT L=0.15 W=0.42
+ AD=0.15435 AS=0.1113 PD=1.155 PS=1.37 NRD=15.708 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1009 N_A_288_74#_M1009_d N_A_28_74#_M1009_g N_VGND_M1006_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.15435 PD=1.37 PS=1.155 NRD=0 NRS=114.276 M=1 R=2.8
+ SA=75001.1 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1001 N_A_549_74#_M1001_d N_A_288_74#_M1001_g N_VGND_M1001_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.2604 PD=1.37 PS=2.08 NRD=0 NRS=99.996 M=1 R=2.8
+ SA=75000.5 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_A_549_74#_M1003_g N_A_682_74#_M1003_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0966 AS=0.2583 PD=0.88 PS=2.07 NRD=51.42 NRS=99.996 M=1 R=2.8
+ SA=75000.5 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1002 N_Y_M1002_d N_A_682_74#_M1002_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0966 PD=1.37 PS=0.88 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1007 N_VPWR_M1007_d N_A_M1007_g N_A_28_74#_M1007_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.397177 AS=0.3136 PD=1.94415 PS=2.8 NRD=5.2599 NRS=2.6201 M=1 R=7.46667
+ SA=75000.2 SB=75001 A=0.168 P=2.54 MULT=1
MM1008 N_A_288_74#_M1008_d N_A_28_74#_M1008_g N_VPWR_M1007_d VPB PHIGHVT L=0.15
+ W=1 AD=0.265 AS=0.354623 PD=2.53 PS=1.73585 NRD=0 NRS=80.77 M=1 R=6.66667
+ SA=75001.1 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1004 N_A_549_74#_M1004_d N_A_288_74#_M1004_g N_VPWR_M1004_s VPB PHIGHVT L=0.15
+ W=1 AD=0.265 AS=0.62 PD=2.53 PS=3.24 NRD=0 NRS=69.9153 M=1 R=6.66667
+ SA=75000.5 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1005 N_VPWR_M1005_d N_A_549_74#_M1005_g N_A_682_74#_M1005_s VPB PHIGHVT L=0.15
+ W=1 AD=0.239623 AS=0.61 PD=1.50472 PS=3.22 NRD=36.7602 NRS=67.9453 M=1
+ R=6.66667 SA=75000.5 SB=75000.8 A=0.15 P=2.3 MULT=1
MM1000 N_Y_M1000_d N_A_682_74#_M1000_g N_VPWR_M1005_d VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3136 AS=0.268377 PD=2.8 PS=1.68528 NRD=2.6201 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75000.2 A=0.168 P=2.54 MULT=1
DX10_noxref VNB VPB NWDIODE A=10.5276 P=15.04
*
.include "sky130_fd_sc_ls__clkdlyinv5sd1_1.pxi.spice"
*
.ends
*
*
