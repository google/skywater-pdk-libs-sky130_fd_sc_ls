* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__dfrbp_1 CLK D RESET_B VGND VNB VPB VPWR Q Q_N
X0 VPWR RESET_B a_1482_48# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_38_78# a_500_392# a_705_463# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 a_705_463# a_500_392# a_832_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 VGND a_705_463# a_841_401# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X4 a_796_463# a_841_401# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 VGND a_2026_424# Q VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X6 a_38_78# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 a_125_78# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_841_401# a_319_392# a_1224_74# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 a_1624_74# a_1224_74# a_1482_48# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_38_78# D a_125_78# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 VPWR a_705_463# a_841_401# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 VGND a_1224_74# Q_N VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X13 VPWR a_319_392# a_500_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 a_319_392# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X15 a_1465_471# a_1482_48# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X16 a_1482_48# a_1224_74# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X17 a_910_119# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 a_2026_424# a_1224_74# VGND VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X19 a_319_392# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X20 a_705_463# a_319_392# a_796_463# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X21 VPWR RESET_B a_705_463# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X22 a_1224_74# a_500_392# a_1465_471# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X23 VPWR a_1224_74# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X24 a_1224_74# a_319_392# a_1434_74# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X25 VGND RESET_B a_1624_74# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X26 a_2026_424# a_1224_74# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X27 VGND a_319_392# a_500_392# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X28 a_1434_74# a_1482_48# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X29 VPWR a_2026_424# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X30 a_832_119# a_841_401# a_910_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X31 a_38_78# a_319_392# a_705_463# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X32 VPWR D a_38_78# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X33 a_841_401# a_500_392# a_1224_74# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
.ends
