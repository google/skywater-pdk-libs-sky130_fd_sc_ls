* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
M1000 a_303_84# B1 a_30_84# VNB nshort w=740000u l=150000u
+  ad=7.067e+11p pd=6.35e+06u as=6.882e+11p ps=6.3e+06u
M1001 VPWR A1 a_505_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=1.3888e+12p pd=1.144e+07u as=9.968e+11p ps=8.5e+06u
M1002 Y C1 a_30_84# VNB nshort w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1003 a_30_84# C1 Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND A2 a_303_84# VNB nshort w=740000u l=150000u
+  ad=6.512e+11p pd=6.2e+06u as=0p ps=0u
M1005 Y B1 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=1.008e+12p pd=8.52e+06u as=0p ps=0u
M1006 a_303_84# A1 VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_505_368# A1 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR B1 Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_303_84# A2 VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND A1 a_303_84# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Y A2 a_505_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_505_368# A2 Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_30_84# B1 a_303_84# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Y C1 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR C1 Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
