# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ls__dlxbp_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ls__dlxbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.160000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.208500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.435000 1.220000 0.835000 1.890000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.537600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.765000 1.820000 6.125000 2.980000 ;
        RECT 5.795000 0.370000 6.125000 1.150000 ;
        RECT 5.955000 1.150000 6.125000 1.820000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.535700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.715000 0.350000 8.050000 2.980000 ;
    END
  END Q_N
  PIN GATE
    ANTENNAGATEAREA  0.237000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.005000 1.180000 1.335000 1.550000 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 8.160000 0.085000 ;
        RECT 0.630000  0.085000 0.960000 1.010000 ;
        RECT 2.355000  0.085000 2.740000 0.410000 ;
        RECT 4.520000  0.085000 4.850000 1.060000 ;
        RECT 6.295000  0.085000 6.545000 1.150000 ;
        RECT 7.285000  0.085000 7.535000 1.130000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
        RECT 6.395000 -0.085000 6.565000 0.085000 ;
        RECT 6.875000 -0.085000 7.045000 0.085000 ;
        RECT 7.355000 -0.085000 7.525000 0.085000 ;
        RECT 7.835000 -0.085000 8.005000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.160000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 8.160000 3.415000 ;
        RECT 0.640000 2.885000 0.970000 3.245000 ;
        RECT 2.380000 2.780000 2.710000 3.245000 ;
        RECT 4.490000 2.545000 5.035000 3.245000 ;
        RECT 6.295000 2.100000 6.545000 3.245000 ;
        RECT 7.270000 1.820000 7.520000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
        RECT 6.395000 3.245000 6.565000 3.415000 ;
        RECT 6.875000 3.245000 7.045000 3.415000 ;
        RECT 7.355000 3.245000 7.525000 3.415000 ;
        RECT 7.835000 3.245000 8.005000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 8.160000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.095000 0.540000 0.450000 1.050000 ;
      RECT 0.095000 1.050000 0.265000 2.060000 ;
      RECT 0.095000 2.060000 0.440000 2.545000 ;
      RECT 0.095000 2.545000 1.760000 2.715000 ;
      RECT 0.095000 2.715000 0.440000 2.925000 ;
      RECT 1.130000 0.350000 1.675000 0.580000 ;
      RECT 1.130000 0.580000 3.080000 0.750000 ;
      RECT 1.130000 0.750000 1.675000 1.010000 ;
      RECT 1.170000 1.720000 2.330000 1.890000 ;
      RECT 1.170000 1.890000 1.420000 2.375000 ;
      RECT 1.505000 1.010000 1.675000 1.470000 ;
      RECT 1.505000 1.470000 2.330000 1.720000 ;
      RECT 1.590000 2.060000 2.875000 2.230000 ;
      RECT 1.590000 2.230000 1.760000 2.545000 ;
      RECT 1.845000 0.920000 2.175000 1.020000 ;
      RECT 1.845000 1.020000 3.515000 1.190000 ;
      RECT 1.930000 2.400000 2.180000 2.440000 ;
      RECT 1.930000 2.440000 4.100000 2.610000 ;
      RECT 1.930000 2.610000 2.180000 2.820000 ;
      RECT 2.545000 1.470000 2.875000 2.060000 ;
      RECT 2.910000 0.255000 4.075000 0.510000 ;
      RECT 2.910000 0.510000 3.080000 0.580000 ;
      RECT 3.045000 1.190000 3.515000 1.480000 ;
      RECT 3.045000 1.480000 3.215000 2.440000 ;
      RECT 3.310000 0.680000 3.950000 0.850000 ;
      RECT 3.385000 1.650000 5.035000 1.820000 ;
      RECT 3.385000 1.820000 3.555000 2.270000 ;
      RECT 3.770000 2.050000 4.100000 2.440000 ;
      RECT 3.780000 0.850000 3.950000 1.650000 ;
      RECT 4.315000 1.990000 5.535000 2.320000 ;
      RECT 4.705000 1.240000 5.035000 1.650000 ;
      RECT 5.020000 0.350000 5.375000 1.070000 ;
      RECT 5.205000 1.070000 5.375000 1.320000 ;
      RECT 5.205000 1.320000 5.775000 1.650000 ;
      RECT 5.205000 1.650000 5.535000 1.990000 ;
      RECT 5.205000 2.320000 5.535000 2.980000 ;
      RECT 6.720000 0.560000 7.055000 1.320000 ;
      RECT 6.720000 1.320000 7.320000 1.650000 ;
      RECT 6.720000 1.650000 7.050000 2.980000 ;
  END
END sky130_fd_sc_ls__dlxbp_1
