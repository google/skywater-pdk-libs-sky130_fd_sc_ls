* File: sky130_fd_sc_ls__and4bb_1.pex.spice
* Created: Fri Aug 28 13:06:06 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__AND4BB_1%A_N 3 5 7 8 12
c26 3 0 1.61433e-19 $X=0.495 $Y=0.645
r27 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.465 $X2=0.27 $Y2=1.465
r28 8 12 7.81317 $w=2.93e-07 $l=2e-07 $layer=LI1_cond $X=0.252 $Y=1.665
+ $X2=0.252 $Y2=1.465
r29 5 11 55.8528 $w=4e-07 $l=3.69459e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.35 $Y2=1.465
r30 5 7 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.26
r31 1 11 39.5853 $w=4e-07 $l=2.26164e-07 $layer=POLY_cond $X=0.495 $Y=1.3
+ $X2=0.35 $Y2=1.465
r32 1 3 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.495 $Y=1.3
+ $X2=0.495 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_LS__AND4BB_1%A_179_48# 1 2 3 12 14 16 20 21 22 24 27 29
+ 33 37 39 42 46
c105 21 0 6.72583e-20 $X=1.82 $Y=0.945
c106 20 0 1.23538e-19 $X=1.525 $Y=1.3
c107 12 0 9.12013e-20 $X=0.97 $Y=0.74
r108 36 39 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=1.38 $Y=1.465
+ $X2=1.525 $Y2=1.465
r109 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.38
+ $Y=1.465 $X2=1.38 $Y2=1.465
r110 31 33 2.26996 $w=3.28e-07 $l=6.5e-08 $layer=LI1_cond $X=3.46 $Y=2.2
+ $X2=3.46 $Y2=2.265
r111 30 46 2.76166 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=2.625 $Y=2.115
+ $X2=2.42 $Y2=2.115
r112 29 31 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.295 $Y=2.115
+ $X2=3.46 $Y2=2.2
r113 29 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.295 $Y=2.115
+ $X2=2.625 $Y2=2.115
r114 25 46 3.70735 $w=2.5e-07 $l=1.03078e-07 $layer=LI1_cond $X=2.46 $Y=2.2
+ $X2=2.42 $Y2=2.115
r115 25 27 2.26996 $w=3.28e-07 $l=6.5e-08 $layer=LI1_cond $X=2.46 $Y=2.2
+ $X2=2.46 $Y2=2.265
r116 24 46 3.70735 $w=2.5e-07 $l=1.56844e-07 $layer=LI1_cond $X=2.3 $Y=2.03
+ $X2=2.42 $Y2=2.115
r117 24 45 65.2406 $w=1.68e-07 $l=1e-06 $layer=LI1_cond $X=2.3 $Y=2.03 $X2=2.3
+ $Y2=1.03
r118 21 45 8.23509 $w=5.63e-07 $l=8.5e-08 $layer=LI1_cond $X=2.102 $Y=0.945
+ $X2=2.102 $Y2=1.03
r119 21 42 9.1029 $w=5.63e-07 $l=4.3e-07 $layer=LI1_cond $X=2.102 $Y=0.945
+ $X2=2.102 $Y2=0.515
r120 21 22 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=1.82 $Y=0.945
+ $X2=1.61 $Y2=0.945
r121 20 39 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.525 $Y=1.3
+ $X2=1.525 $Y2=1.465
r122 19 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.525 $Y=1.03
+ $X2=1.61 $Y2=0.945
r123 19 20 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=1.525 $Y=1.03
+ $X2=1.525 $Y2=1.3
r124 18 37 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=1.13 $Y=1.465
+ $X2=1.38 $Y2=1.465
r125 14 18 76.2621 $w=1.97e-07 $l=3.13688e-07 $layer=POLY_cond $X=1.04 $Y=1.765
+ $X2=1.012 $Y2=1.465
r126 14 16 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.04 $Y=1.765
+ $X2=1.04 $Y2=2.4
r127 10 18 43.2316 $w=1.97e-07 $l=1.84811e-07 $layer=POLY_cond $X=0.97 $Y=1.3
+ $X2=1.012 $Y2=1.465
r128 10 12 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.97 $Y=1.3
+ $X2=0.97 $Y2=0.74
r129 3 33 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=3.31
+ $Y=2.12 $X2=3.46 $Y2=2.265
r130 2 27 300 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=2 $X=2.26
+ $Y=2.12 $X2=2.46 $Y2=2.265
r131 1 42 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=1.84
+ $Y=0.37 $X2=1.985 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__AND4BB_1%A_27_74# 1 2 7 9 12 16 18 19 21 22 26 30
c82 12 0 2.32305e-19 $X=2.2 $Y=0.69
c83 7 0 2.14739e-19 $X=2.185 $Y=2.045
r84 30 31 6.52768 $w=5.42e-07 $l=2.9e-07 $layer=LI1_cond $X=0.427 $Y=2.115
+ $X2=0.427 $Y2=2.405
r85 26 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.92
+ $Y=1.455 $X2=1.92 $Y2=1.455
r86 24 26 37.6175 $w=2.63e-07 $l=8.65e-07 $layer=LI1_cond $X=1.912 $Y=2.32
+ $X2=1.912 $Y2=1.455
r87 23 31 7.66608 $w=1.7e-07 $l=3.13e-07 $layer=LI1_cond $X=0.74 $Y=2.405
+ $X2=0.427 $Y2=2.405
r88 22 24 7.24806 $w=1.7e-07 $l=1.69245e-07 $layer=LI1_cond $X=1.78 $Y=2.405
+ $X2=1.912 $Y2=2.32
r89 22 23 67.8503 $w=1.68e-07 $l=1.04e-06 $layer=LI1_cond $X=1.78 $Y=2.405
+ $X2=0.74 $Y2=2.405
r90 21 30 9.97635 $w=5.42e-07 $l=2.99339e-07 $layer=LI1_cond $X=0.655 $Y=1.95
+ $X2=0.427 $Y2=2.115
r91 20 21 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=0.655 $Y=1.13
+ $X2=0.655 $Y2=1.95
r92 18 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.57 $Y=1.045
+ $X2=0.655 $Y2=1.13
r93 18 19 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=0.57 $Y=1.045
+ $X2=0.365 $Y2=1.045
r94 14 19 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.24 $Y=0.96
+ $X2=0.365 $Y2=1.045
r95 14 16 14.5208 $w=2.48e-07 $l=3.15e-07 $layer=LI1_cond $X=0.24 $Y=0.96
+ $X2=0.24 $Y2=0.645
r96 10 27 41.4407 $w=4.81e-07 $l=2.5446e-07 $layer=POLY_cond $X=2.2 $Y=1.29
+ $X2=2.015 $Y2=1.455
r97 10 12 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=2.2 $Y=1.29 $X2=2.2
+ $Y2=0.69
r98 7 27 84.0291 $w=4.81e-07 $l=6.69627e-07 $layer=POLY_cond $X=2.185 $Y=2.045
+ $X2=2.015 $Y2=1.455
r99 7 9 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.185 $Y=2.045
+ $X2=2.185 $Y2=2.54
r100 2 30 300 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.115
r101 1 16 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_LS__AND4BB_1%A_503_48# 1 2 9 11 12 14 16 17 18 21 22 25
+ 27 28 30 32 36
c92 25 0 1.65047e-19 $X=2.845 $Y=0.935
r93 35 36 5.28416 $w=1.78e-07 $l=8.5e-08 $layer=LI1_cond $X=4.145 $Y=0.94
+ $X2=4.06 $Y2=0.94
r94 32 35 23.1061 $w=1.78e-07 $l=3.75e-07 $layer=LI1_cond $X=4.52 $Y=0.94
+ $X2=4.145 $Y2=0.94
r95 32 34 4.25152 $w=3.3e-07 $l=1.15e-07 $layer=LI1_cond $X=4.52 $Y=0.85
+ $X2=4.52 $Y2=0.735
r96 28 39 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=4.48 $Y=2.035
+ $X2=4.145 $Y2=2.035
r97 28 30 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=4.48 $Y=2.12
+ $X2=4.48 $Y2=2.265
r98 27 39 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.145 $Y=1.95
+ $X2=4.145 $Y2=2.035
r99 26 35 1.06262 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=4.145 $Y=1.03 $X2=4.145
+ $Y2=0.94
r100 26 27 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=4.145 $Y=1.03
+ $X2=4.145 $Y2=1.95
r101 25 36 79.2674 $w=1.68e-07 $l=1.215e-06 $layer=LI1_cond $X=2.845 $Y=0.935
+ $X2=4.06 $Y2=0.935
r102 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.68
+ $Y=1.285 $X2=2.68 $Y2=1.285
r103 19 25 7.43784 $w=1.7e-07 $l=1.8262e-07 $layer=LI1_cond $X=2.7 $Y=1.02
+ $X2=2.845 $Y2=0.935
r104 19 21 10.5309 $w=2.88e-07 $l=2.65e-07 $layer=LI1_cond $X=2.7 $Y=1.02
+ $X2=2.7 $Y2=1.285
r105 17 22 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.68 $Y=1.625
+ $X2=2.68 $Y2=1.285
r106 17 18 34.9753 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.68 $Y=1.625
+ $X2=2.68 $Y2=1.79
r107 16 22 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.68 $Y=1.12
+ $X2=2.68 $Y2=1.285
r108 12 14 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.685 $Y=2.045
+ $X2=2.685 $Y2=2.54
r109 11 12 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.685 $Y=1.955
+ $X2=2.685 $Y2=2.045
r110 11 18 64.1371 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.685 $Y=1.955
+ $X2=2.685 $Y2=1.79
r111 9 16 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.59 $Y=0.69
+ $X2=2.59 $Y2=1.12
r112 2 30 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=4.33
+ $Y=2.12 $X2=4.48 $Y2=2.265
r113 1 34 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=4.38
+ $Y=0.46 $X2=4.52 $Y2=0.735
.ends

.subckt PM_SKY130_FD_SC_LS__AND4BB_1%C 3 5 7 10 11 14 15
r40 14 15 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.22
+ $Y=1.355 $X2=3.22 $Y2=1.355
r41 11 15 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=3.18 $Y=1.665
+ $X2=3.18 $Y2=1.355
r42 10 14 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.22 $Y=1.695
+ $X2=3.22 $Y2=1.355
r43 9 14 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.22 $Y=1.19
+ $X2=3.22 $Y2=1.355
r44 5 10 67.48 $w=2.5e-07 $l=3.57421e-07 $layer=POLY_cond $X=3.235 $Y=2.045
+ $X2=3.22 $Y2=1.695
r45 5 7 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=3.235 $Y=2.045
+ $X2=3.235 $Y2=2.54
r46 3 9 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=3.16 $Y=0.69 $X2=3.16
+ $Y2=1.19
.ends

.subckt PM_SKY130_FD_SC_LS__AND4BB_1%D 3 5 7 10 11 14 15
r43 14 15 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.76
+ $Y=1.355 $X2=3.76 $Y2=1.355
r44 11 15 2.85631 $w=6.68e-07 $l=1.6e-07 $layer=LI1_cond $X=3.6 $Y=1.525
+ $X2=3.76 $Y2=1.525
r45 10 14 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.76 $Y=1.695
+ $X2=3.76 $Y2=1.355
r46 9 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.76 $Y=1.19
+ $X2=3.76 $Y2=1.355
r47 5 10 67.48 $w=2.5e-07 $l=3.85681e-07 $layer=POLY_cond $X=3.685 $Y=2.045
+ $X2=3.76 $Y2=1.695
r48 5 7 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=3.685 $Y=2.045
+ $X2=3.685 $Y2=2.54
r49 3 9 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=3.67 $Y=0.69 $X2=3.67
+ $Y2=1.19
.ends

.subckt PM_SKY130_FD_SC_LS__AND4BB_1%B_N 2 3 5 8 10 16 17
r33 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.53
+ $Y=1.465 $X2=4.53 $Y2=1.465
r34 14 16 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=4.305 $Y=1.465
+ $X2=4.53 $Y2=1.465
r35 12 14 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=4.255 $Y=1.465
+ $X2=4.305 $Y2=1.465
r36 10 17 7.81317 $w=2.93e-07 $l=2e-07 $layer=LI1_cond $X=4.547 $Y=1.665
+ $X2=4.547 $Y2=1.465
r37 6 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.305 $Y=1.3
+ $X2=4.305 $Y2=1.465
r38 6 8 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=4.305 $Y=1.3
+ $X2=4.305 $Y2=0.735
r39 3 5 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=4.255 $Y=2.045
+ $X2=4.255 $Y2=2.54
r40 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=4.255 $Y=1.955 $X2=4.255
+ $Y2=2.045
r41 1 12 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.255 $Y=1.63
+ $X2=4.255 $Y2=1.465
r42 1 2 126.331 $w=1.8e-07 $l=3.25e-07 $layer=POLY_cond $X=4.255 $Y=1.63
+ $X2=4.255 $Y2=1.955
.ends

.subckt PM_SKY130_FD_SC_LS__AND4BB_1%VPWR 1 2 3 4 17 21 25 29 32 33 35 36 38 39
+ 40 53 54 57
r64 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r65 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r66 51 54 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r67 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r68 48 51 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r69 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r70 45 58 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r71 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r72 42 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.98 $Y=3.33
+ $X2=0.815 $Y2=3.33
r73 42 44 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=0.98 $Y=3.33 $X2=1.68
+ $Y2=3.33
r74 40 48 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=2.64 $Y2=3.33
r75 40 45 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=1.68 $Y2=3.33
r76 38 50 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=3.815 $Y=3.33
+ $X2=3.6 $Y2=3.33
r77 38 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.815 $Y=3.33
+ $X2=3.98 $Y2=3.33
r78 37 53 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=4.145 $Y=3.33
+ $X2=4.56 $Y2=3.33
r79 37 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.145 $Y=3.33
+ $X2=3.98 $Y2=3.33
r80 35 47 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=2.795 $Y=3.33
+ $X2=2.64 $Y2=3.33
r81 35 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.795 $Y=3.33
+ $X2=2.96 $Y2=3.33
r82 34 50 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=3.125 $Y=3.33
+ $X2=3.6 $Y2=3.33
r83 34 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.125 $Y=3.33
+ $X2=2.96 $Y2=3.33
r84 32 44 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=1.795 $Y=3.33
+ $X2=1.68 $Y2=3.33
r85 32 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.795 $Y=3.33
+ $X2=1.96 $Y2=3.33
r86 31 47 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=2.125 $Y=3.33
+ $X2=2.64 $Y2=3.33
r87 31 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.125 $Y=3.33
+ $X2=1.96 $Y2=3.33
r88 27 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.98 $Y=3.245
+ $X2=3.98 $Y2=3.33
r89 27 29 29.8588 $w=3.28e-07 $l=8.55e-07 $layer=LI1_cond $X=3.98 $Y=3.245
+ $X2=3.98 $Y2=2.39
r90 23 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.96 $Y=3.245
+ $X2=2.96 $Y2=3.33
r91 23 25 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=2.96 $Y=3.245
+ $X2=2.96 $Y2=2.455
r92 19 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.96 $Y=3.245
+ $X2=1.96 $Y2=3.33
r93 19 21 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=1.96 $Y=3.245
+ $X2=1.96 $Y2=2.78
r94 15 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=3.245
+ $X2=0.815 $Y2=3.33
r95 15 17 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=0.815 $Y=3.245
+ $X2=0.815 $Y2=2.78
r96 4 29 300 $w=1.7e-07 $l=3.63731e-07 $layer=licon1_PDIFF $count=2 $X=3.76
+ $Y=2.12 $X2=3.98 $Y2=2.39
r97 3 25 300 $w=1.7e-07 $l=4.2335e-07 $layer=licon1_PDIFF $count=2 $X=2.76
+ $Y=2.12 $X2=2.96 $Y2=2.455
r98 2 21 600 $w=1.7e-07 $l=7.28903e-07 $layer=licon1_PDIFF $count=1 $X=1.815
+ $Y=2.12 $X2=1.96 $Y2=2.78
r99 1 17 600 $w=1.7e-07 $l=1.05095e-06 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.84 $X2=0.815 $Y2=2.78
.ends

.subckt PM_SKY130_FD_SC_LS__AND4BB_1%X 1 2 8 11 15 17 18 23
c35 17 0 1.20215e-19 $X=1.08 $Y=1.985
c36 15 0 1.61433e-19 $X=1.175 $Y=1.045
r37 18 23 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=1.2 $Y=1.985
+ $X2=1.33 $Y2=1.985
r38 17 18 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=1.08 $Y=1.985 $X2=1.2
+ $Y2=1.985
r39 13 15 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.995 $Y=1.045
+ $X2=1.175 $Y2=1.045
r40 9 15 0.0262452 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.175 $Y=0.96
+ $X2=1.175 $Y2=1.045
r41 9 11 25.9761 $w=1.88e-07 $l=4.45e-07 $layer=LI1_cond $X=1.175 $Y=0.96
+ $X2=1.175 $Y2=0.515
r42 8 17 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.995 $Y=1.82
+ $X2=1.08 $Y2=1.985
r43 7 13 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.995 $Y=1.13
+ $X2=0.995 $Y2=1.045
r44 7 8 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=0.995 $Y=1.13 $X2=0.995
+ $Y2=1.82
r45 2 23 600 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_PDIFF $count=1 $X=1.115
+ $Y=1.84 $X2=1.33 $Y2=1.985
r46 1 11 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.045
+ $Y=0.37 $X2=1.185 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__AND4BB_1%VGND 1 2 9 13 16 17 18 20 33 34 37
r47 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r48 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r49 31 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r50 30 31 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r51 28 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r52 27 30 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=3.6
+ $Y2=0
r53 27 28 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r54 25 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=0.71
+ $Y2=0
r55 25 27 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=1.2
+ $Y2=0
r56 23 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r57 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r58 20 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.71
+ $Y2=0
r59 20 22 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.24
+ $Y2=0
r60 18 31 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=2.4 $Y=0 $X2=3.6
+ $Y2=0
r61 18 28 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=2.4 $Y=0 $X2=1.2
+ $Y2=0
r62 16 30 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=3.72 $Y=0 $X2=3.6
+ $Y2=0
r63 16 17 9.6488 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=3.72 $Y=0 $X2=3.915
+ $Y2=0
r64 15 33 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=4.11 $Y=0 $X2=4.56
+ $Y2=0
r65 15 17 9.6488 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=4.11 $Y=0 $X2=3.915
+ $Y2=0
r66 11 17 1.39532 $w=3.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.915 $Y=0.085
+ $X2=3.915 $Y2=0
r67 11 13 12.7064 $w=3.88e-07 $l=4.3e-07 $layer=LI1_cond $X=3.915 $Y=0.085
+ $X2=3.915 $Y2=0.515
r68 7 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=0.085 $X2=0.71
+ $Y2=0
r69 7 9 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=0.71 $Y=0.085 $X2=0.71
+ $Y2=0.625
r70 2 13 182 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_NDIFF $count=1 $X=3.745
+ $Y=0.37 $X2=3.945 $Y2=0.515
r71 1 9 182 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.625
.ends

