* File: sky130_fd_sc_ls__nor3b_1.pex.spice
* Created: Fri Aug 28 13:38:58 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__NOR3B_1%C_N 1 3 4 6 7
r27 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.61
+ $Y=1.385 $X2=0.61 $Y2=1.385
r28 7 11 3.42618 $w=3.68e-07 $l=1.1e-07 $layer=LI1_cond $X=0.72 $Y=1.365
+ $X2=0.61 $Y2=1.365
r29 4 10 38.9026 $w=2.7e-07 $l=2.05122e-07 $layer=POLY_cond $X=0.7 $Y=1.22
+ $X2=0.61 $Y2=1.385
r30 4 6 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=0.7 $Y=1.22 $X2=0.7
+ $Y2=0.835
r31 1 10 77.2841 $w=2.7e-07 $l=4.01871e-07 $layer=POLY_cond $X=0.655 $Y=1.765
+ $X2=0.61 $Y2=1.385
r32 1 3 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.655 $Y=1.765
+ $X2=0.655 $Y2=2.26
.ends

.subckt PM_SKY130_FD_SC_LS__NOR3B_1%A 1 3 6 8 12
r29 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.15
+ $Y=1.515 $X2=1.15 $Y2=1.515
r30 8 12 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.15 $Y=1.665
+ $X2=1.15 $Y2=1.515
r31 4 11 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=1.24 $Y=1.35
+ $X2=1.15 $Y2=1.515
r32 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.24 $Y=1.35 $X2=1.24
+ $Y2=0.74
r33 1 11 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=1.225 $Y=1.765
+ $X2=1.15 $Y2=1.515
r34 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.225 $Y=1.765
+ $X2=1.225 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__NOR3B_1%B 1 3 6 8 12
r33 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.72
+ $Y=1.515 $X2=1.72 $Y2=1.515
r34 8 12 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.72 $Y=1.665
+ $X2=1.72 $Y2=1.515
r35 4 11 38.5562 $w=2.99e-07 $l=1.69926e-07 $layer=POLY_cond $X=1.71 $Y=1.35
+ $X2=1.72 $Y2=1.515
r36 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.71 $Y=1.35 $X2=1.71
+ $Y2=0.74
r37 1 11 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=1.645 $Y=1.765
+ $X2=1.72 $Y2=1.515
r38 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.645 $Y=1.765
+ $X2=1.645 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__NOR3B_1%A_27_112# 1 2 7 9 12 18 21 25 28 29 30 32
r62 32 35 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.29 $Y=1.515
+ $X2=2.29 $Y2=1.68
r63 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.29
+ $Y=1.515 $X2=2.29 $Y2=1.515
r64 28 30 1.22049 $w=4.88e-07 $l=5e-08 $layer=LI1_cond $X=0.35 $Y=1.985 $X2=0.35
+ $Y2=2.035
r65 28 29 9.45624 $w=4.88e-07 $l=1.65e-07 $layer=LI1_cond $X=0.35 $Y=1.985
+ $X2=0.35 $Y2=1.82
r66 22 25 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.19 $Y=0.845
+ $X2=0.485 $Y2=0.845
r67 21 35 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=2.21 $Y=1.95 $X2=2.21
+ $Y2=1.68
r68 19 30 7.03003 $w=1.7e-07 $l=2.45e-07 $layer=LI1_cond $X=0.595 $Y=2.035
+ $X2=0.35 $Y2=2.035
r69 18 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.125 $Y=2.035
+ $X2=2.21 $Y2=1.95
r70 18 19 99.8182 $w=1.68e-07 $l=1.53e-06 $layer=LI1_cond $X=2.125 $Y=2.035
+ $X2=0.595 $Y2=2.035
r71 14 22 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.19 $Y=1.01
+ $X2=0.19 $Y2=0.845
r72 14 29 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=0.19 $Y=1.01
+ $X2=0.19 $Y2=1.82
r73 10 33 38.5562 $w=2.99e-07 $l=1.69926e-07 $layer=POLY_cond $X=2.28 $Y=1.35
+ $X2=2.29 $Y2=1.515
r74 10 12 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.28 $Y=1.35
+ $X2=2.28 $Y2=0.74
r75 7 33 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=2.215 $Y=1.765
+ $X2=2.29 $Y2=1.515
r76 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.215 $Y=1.765
+ $X2=2.215 $Y2=2.4
r77 2 28 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.285
+ $Y=1.84 $X2=0.43 $Y2=1.985
r78 1 25 182 $w=1.7e-07 $l=4.71434e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.56 $X2=0.485 $Y2=0.845
.ends

.subckt PM_SKY130_FD_SC_LS__NOR3B_1%VPWR 1 6 9 10 11 21 22
r24 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r25 18 21 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r26 18 19 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r27 15 19 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r28 14 15 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r29 11 22 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=2.64 $Y2=3.33
r30 11 19 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.2 $Y2=3.33
r31 9 14 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=0.835 $Y=3.33
+ $X2=0.72 $Y2=3.33
r32 9 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.835 $Y=3.33 $X2=1
+ $Y2=3.33
r33 8 18 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=1.165 $Y=3.33 $X2=1.2
+ $Y2=3.33
r34 8 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.165 $Y=3.33 $X2=1
+ $Y2=3.33
r35 4 10 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1 $Y=3.245 $X2=1
+ $Y2=3.33
r36 4 6 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=1 $Y=3.245 $X2=1
+ $Y2=2.455
r37 1 6 300 $w=1.7e-07 $l=7.3775e-07 $layer=licon1_PDIFF $count=2 $X=0.73
+ $Y=1.84 $X2=1 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_LS__NOR3B_1%Y 1 2 3 12 14 15 19 20 22 23 29 35
r45 23 35 2.40447 $w=4.02e-07 $l=1.17707e-07 $layer=LI1_cond $X=2.64 $Y=1.01
+ $X2=2.562 $Y2=1.095
r46 22 23 9.51718 $w=4.63e-07 $l=3.7e-07 $layer=LI1_cond $X=2.562 $Y=0.555
+ $X2=2.562 $Y2=0.925
r47 22 29 1.02888 $w=4.63e-07 $l=4e-08 $layer=LI1_cond $X=2.562 $Y=0.555
+ $X2=2.562 $Y2=0.515
r48 19 20 9.6413 $w=5.18e-07 $l=1.65e-07 $layer=LI1_cond $X=2.535 $Y=2.455
+ $X2=2.535 $Y2=2.29
r49 16 35 2.40447 $w=4.02e-07 $l=1.85699e-07 $layer=LI1_cond $X=2.71 $Y=1.18
+ $X2=2.562 $Y2=1.095
r50 16 20 72.4171 $w=1.68e-07 $l=1.11e-06 $layer=LI1_cond $X=2.71 $Y=1.18
+ $X2=2.71 $Y2=2.29
r51 14 35 4.56719 $w=1.7e-07 $l=2.32e-07 $layer=LI1_cond $X=2.33 $Y=1.095
+ $X2=2.562 $Y2=1.095
r52 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.33 $Y=1.095
+ $X2=1.66 $Y2=1.095
r53 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.495 $Y=1.01
+ $X2=1.66 $Y2=1.095
r54 10 12 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=1.495 $Y=1.01
+ $X2=1.495 $Y2=0.515
r55 3 19 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=2.29
+ $Y=1.84 $X2=2.44 $Y2=2.455
r56 2 29 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.355
+ $Y=0.37 $X2=2.495 $Y2=0.515
r57 1 12 91 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_NDIFF $count=2 $X=1.315
+ $Y=0.37 $X2=1.495 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__NOR3B_1%VGND 1 2 9 13 16 17 19 20 21 31 32
r33 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r34 29 32 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r35 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r36 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r37 21 29 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.68
+ $Y2=0
r38 21 25 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=0.72
+ $Y2=0
r39 19 28 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=1.83 $Y=0 $X2=1.68
+ $Y2=0
r40 19 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.83 $Y=0 $X2=1.995
+ $Y2=0
r41 18 31 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r42 18 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.16 $Y=0 $X2=1.995
+ $Y2=0
r43 16 24 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=0.83 $Y=0 $X2=0.72
+ $Y2=0
r44 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.83 $Y=0 $X2=0.995
+ $Y2=0
r45 15 28 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.16 $Y=0 $X2=1.68
+ $Y2=0
r46 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.16 $Y=0 $X2=0.995
+ $Y2=0
r47 11 20 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.995 $Y=0.085
+ $X2=1.995 $Y2=0
r48 11 13 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=1.995 $Y=0.085
+ $X2=1.995 $Y2=0.675
r49 7 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.995 $Y=0.085
+ $X2=0.995 $Y2=0
r50 7 9 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.995 $Y=0.085
+ $X2=0.995 $Y2=0.515
r51 2 13 182 $w=1.7e-07 $l=3.96327e-07 $layer=licon1_NDIFF $count=1 $X=1.785
+ $Y=0.37 $X2=1.995 $Y2=0.675
r52 1 9 91 $w=1.7e-07 $l=2.41454e-07 $layer=licon1_NDIFF $count=2 $X=0.775
+ $Y=0.56 $X2=0.995 $Y2=0.515
.ends

