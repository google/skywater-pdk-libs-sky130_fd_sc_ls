* File: sky130_fd_sc_ls__nor4_1.spice
* Created: Fri Aug 28 13:39:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__nor4_1.pex.spice"
.subckt sky130_fd_sc_ls__nor4_1  VNB VPB A B C D VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* D	D
* C	C
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1000 N_Y_M1000_d N_A_M1000_g N_VGND_M1000_s VNB NSHORT L=0.15 W=0.74 AD=0.1036
+ AS=0.2627 PD=1.02 PS=2.19 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.3 SB=75001.8
+ A=0.111 P=1.78 MULT=1
MM1004 N_VGND_M1004_d N_B_M1004_g N_Y_M1000_d VNB NSHORT L=0.15 W=0.74 AD=0.1924
+ AS=0.1036 PD=1.26 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.7 SB=75001.3
+ A=0.111 P=1.78 MULT=1
MM1005 N_Y_M1005_d N_C_M1005_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.74 AD=0.1036
+ AS=0.1924 PD=1.02 PS=1.26 NRD=0 NRS=27.564 M=1 R=4.93333 SA=75001.4 SB=75000.7
+ A=0.111 P=1.78 MULT=1
MM1006 N_VGND_M1006_d N_D_M1006_g N_Y_M1005_d VNB NSHORT L=0.15 W=0.74
+ AD=0.23225 AS=0.1036 PD=2.19 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.8
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1007 A_144_368# N_A_M1007_g N_VPWR_M1007_s VPB PHIGHVT L=0.15 W=1.12 AD=0.1512
+ AS=0.3304 PD=1.39 PS=2.83 NRD=14.0658 NRS=1.7533 M=1 R=7.46667 SA=75000.2
+ SB=75001.8 A=0.168 P=2.54 MULT=1
MM1002 A_228_368# N_B_M1002_g A_144_368# VPB PHIGHVT L=0.15 W=1.12 AD=0.2352
+ AS=0.1512 PD=1.54 PS=1.39 NRD=27.2451 NRS=14.0658 M=1 R=7.46667 SA=75000.6
+ SB=75001.4 A=0.168 P=2.54 MULT=1
MM1003 A_342_368# N_C_M1003_g A_228_368# VPB PHIGHVT L=0.15 W=1.12 AD=0.2352
+ AS=0.2352 PD=1.54 PS=1.54 NRD=27.2451 NRS=27.2451 M=1 R=7.46667 SA=75001.2
+ SB=75000.8 A=0.168 P=2.54 MULT=1
MM1001 N_Y_M1001_d N_D_M1001_g A_342_368# VPB PHIGHVT L=0.15 W=1.12 AD=0.3304
+ AS=0.2352 PD=2.83 PS=1.54 NRD=1.7533 NRS=27.2451 M=1 R=7.46667 SA=75001.8
+ SB=75000.2 A=0.168 P=2.54 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.0636 P=10.24
*
.include "sky130_fd_sc_ls__nor4_1.pxi.spice"
*
.ends
*
*
