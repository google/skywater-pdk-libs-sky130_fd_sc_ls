* File: sky130_fd_sc_ls__inv_16.spice
* Created: Fri Aug 28 13:27:55 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__inv_16.pex.spice"
.subckt sky130_fd_sc_ls__inv_16  VNB VPB A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1002 N_Y_M1002_d N_A_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.74 AD=0.1036
+ AS=0.1961 PD=1.02 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2 SB=75007.2
+ A=0.111 P=1.78 MULT=1
MM1003 N_Y_M1002_d N_A_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.74 AD=0.1036
+ AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75000.6 SB=75006.8
+ A=0.111 P=1.78 MULT=1
MM1005 N_Y_M1005_d N_A_M1005_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.74 AD=0.1036
+ AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1 SB=75006.3
+ A=0.111 P=1.78 MULT=1
MM1008 N_Y_M1005_d N_A_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.74 AD=0.1036
+ AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.6 SB=75005.9
+ A=0.111 P=1.78 MULT=1
MM1009 N_Y_M1009_d N_A_M1009_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.74 AD=0.1036
+ AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75002.1 SB=75005.4
+ A=0.111 P=1.78 MULT=1
MM1011 N_Y_M1009_d N_A_M1011_g N_VGND_M1011_s VNB NSHORT L=0.15 W=0.74 AD=0.1036
+ AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=8.1 M=1 R=4.93333 SA=75002.5 SB=75004.9
+ A=0.111 P=1.78 MULT=1
MM1012 N_Y_M1012_d N_A_M1012_g N_VGND_M1011_s VNB NSHORT L=0.15 W=0.74 AD=0.1036
+ AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=3.24 M=1 R=4.93333 SA=75003 SB=75004.4
+ A=0.111 P=1.78 MULT=1
MM1013 N_Y_M1012_d N_A_M1013_g N_VGND_M1013_s VNB NSHORT L=0.15 W=0.74 AD=0.1036
+ AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75003.4 SB=75004
+ A=0.111 P=1.78 MULT=1
MM1014 N_Y_M1014_d N_A_M1014_g N_VGND_M1013_s VNB NSHORT L=0.15 W=0.74 AD=0.1036
+ AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75003.8 SB=75003.6
+ A=0.111 P=1.78 MULT=1
MM1015 N_Y_M1014_d N_A_M1015_g N_VGND_M1015_s VNB NSHORT L=0.15 W=0.74 AD=0.1036
+ AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=5.664 M=1 R=4.93333 SA=75004.3 SB=75003.1
+ A=0.111 P=1.78 MULT=1
MM1018 N_Y_M1018_d N_A_M1018_g N_VGND_M1015_s VNB NSHORT L=0.15 W=0.74 AD=0.1036
+ AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=5.664 M=1 R=4.93333 SA=75004.8 SB=75002.6
+ A=0.111 P=1.78 MULT=1
MM1019 N_Y_M1018_d N_A_M1019_g N_VGND_M1019_s VNB NSHORT L=0.15 W=0.74 AD=0.1036
+ AS=0.1554 PD=1.02 PS=1.16 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75005.2 SB=75002.2
+ A=0.111 P=1.78 MULT=1
MM1023 N_Y_M1023_d N_A_M1023_g N_VGND_M1019_s VNB NSHORT L=0.15 W=0.74 AD=0.1036
+ AS=0.1554 PD=1.02 PS=1.16 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75005.8 SB=75001.6
+ A=0.111 P=1.78 MULT=1
MM1027 N_Y_M1023_d N_A_M1027_g N_VGND_M1027_s VNB NSHORT L=0.15 W=0.74 AD=0.1036
+ AS=0.1628 PD=1.02 PS=1.18 NRD=0 NRS=12.972 M=1 R=4.93333 SA=75006.2 SB=75001.2
+ A=0.111 P=1.78 MULT=1
MM1029 N_Y_M1029_d N_A_M1029_g N_VGND_M1027_s VNB NSHORT L=0.15 W=0.74 AD=0.1036
+ AS=0.1628 PD=1.02 PS=1.18 NRD=0 NRS=12.972 M=1 R=4.93333 SA=75006.8 SB=75000.6
+ A=0.111 P=1.78 MULT=1
MM1031 N_Y_M1029_d N_A_M1031_g N_VGND_M1031_s VNB NSHORT L=0.15 W=0.74 AD=0.1036
+ AS=0.1961 PD=1.02 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333 SA=75007.2 SB=75000.2
+ A=0.111 P=1.78 MULT=1
MM1000 N_VPWR_M1000_d N_A_M1000_g N_Y_M1000_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75007.4 A=0.168 P=2.54 MULT=1
MM1001 N_VPWR_M1001_d N_A_M1001_g N_Y_M1000_s VPB PHIGHVT L=0.15 W=1.12 AD=0.196
+ AS=0.168 PD=1.47 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75000.7
+ SB=75006.9 A=0.168 P=2.54 MULT=1
MM1004 N_VPWR_M1001_d N_A_M1004_g N_Y_M1004_s VPB PHIGHVT L=0.15 W=1.12 AD=0.196
+ AS=0.168 PD=1.47 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667 SA=75001.2
+ SB=75006.4 A=0.168 P=2.54 MULT=1
MM1006 N_VPWR_M1006_d N_A_M1006_g N_Y_M1004_s VPB PHIGHVT L=0.15 W=1.12 AD=0.196
+ AS=0.168 PD=1.47 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75001.6
+ SB=75006 A=0.168 P=2.54 MULT=1
MM1007 N_VPWR_M1006_d N_A_M1007_g N_Y_M1007_s VPB PHIGHVT L=0.15 W=1.12 AD=0.196
+ AS=0.168 PD=1.47 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667 SA=75002.1
+ SB=75005.5 A=0.168 P=2.54 MULT=1
MM1010 N_VPWR_M1010_d N_A_M1010_g N_Y_M1007_s VPB PHIGHVT L=0.15 W=1.12 AD=0.196
+ AS=0.168 PD=1.47 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75002.6
+ SB=75005 A=0.168 P=2.54 MULT=1
MM1016 N_VPWR_M1010_d N_A_M1016_g N_Y_M1016_s VPB PHIGHVT L=0.15 W=1.12 AD=0.196
+ AS=0.168 PD=1.47 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667 SA=75003.1
+ SB=75004.5 A=0.168 P=2.54 MULT=1
MM1017 N_VPWR_M1017_d N_A_M1017_g N_Y_M1016_s VPB PHIGHVT L=0.15 W=1.12 AD=0.168
+ AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75003.5
+ SB=75004.1 A=0.168 P=2.54 MULT=1
MM1020 N_VPWR_M1017_d N_A_M1020_g N_Y_M1020_s VPB PHIGHVT L=0.15 W=1.12 AD=0.168
+ AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75004
+ SB=75003.6 A=0.168 P=2.54 MULT=1
MM1021 N_VPWR_M1021_d N_A_M1021_g N_Y_M1020_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.1792 AS=0.168 PD=1.44 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75004.4 SB=75003.2 A=0.168 P=2.54 MULT=1
MM1022 N_VPWR_M1021_d N_A_M1022_g N_Y_M1022_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.1792 AS=0.1848 PD=1.44 PS=1.45 NRD=5.2599 NRS=7.0329 M=1 R=7.46667
+ SA=75004.9 SB=75002.7 A=0.168 P=2.54 MULT=1
MM1024 N_VPWR_M1024_d N_A_M1024_g N_Y_M1022_s VPB PHIGHVT L=0.15 W=1.12 AD=0.224
+ AS=0.1848 PD=1.52 PS=1.45 NRD=10.5395 NRS=1.7533 M=1 R=7.46667 SA=75005.4
+ SB=75002.2 A=0.168 P=2.54 MULT=1
MM1025 N_VPWR_M1024_d N_A_M1025_g N_Y_M1025_s VPB PHIGHVT L=0.15 W=1.12 AD=0.224
+ AS=0.168 PD=1.52 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667 SA=75005.9
+ SB=75001.7 A=0.168 P=2.54 MULT=1
MM1026 N_VPWR_M1026_d N_A_M1026_g N_Y_M1025_s VPB PHIGHVT L=0.15 W=1.12 AD=0.224
+ AS=0.168 PD=1.52 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667 SA=75006.4
+ SB=75001.2 A=0.168 P=2.54 MULT=1
MM1028 N_VPWR_M1026_d N_A_M1028_g N_Y_M1028_s VPB PHIGHVT L=0.15 W=1.12 AD=0.224
+ AS=0.168 PD=1.52 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667 SA=75006.9
+ SB=75000.7 A=0.168 P=2.54 MULT=1
MM1030 N_VPWR_M1030_d N_A_M1030_g N_Y_M1028_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75007.4 SB=75000.2 A=0.168 P=2.54 MULT=1
DX32_noxref VNB VPB NWDIODE A=15.8844 P=20.8
c_69 VNB 0 1.71499e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_ls__inv_16.pxi.spice"
*
.ends
*
*
