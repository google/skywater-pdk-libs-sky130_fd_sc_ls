* File: sky130_fd_sc_ls__maj3_2.pxi.spice
* Created: Fri Aug 28 13:29:08 2020
* 
x_PM_SKY130_FD_SC_LS__MAJ3_2%A_87_264# N_A_87_264#_M1009_d N_A_87_264#_M1012_d
+ N_A_87_264#_M1014_d N_A_87_264#_M1005_d N_A_87_264#_M1010_g N_A_87_264#_c_85_n
+ N_A_87_264#_M1002_g N_A_87_264#_M1013_g N_A_87_264#_c_86_n N_A_87_264#_M1003_g
+ N_A_87_264#_c_87_n N_A_87_264#_c_79_n N_A_87_264#_c_80_n N_A_87_264#_c_100_p
+ N_A_87_264#_c_81_n N_A_87_264#_c_89_n N_A_87_264#_c_90_n N_A_87_264#_c_82_n
+ N_A_87_264#_c_83_n N_A_87_264#_c_92_n N_A_87_264#_c_84_n
+ PM_SKY130_FD_SC_LS__MAJ3_2%A_87_264#
x_PM_SKY130_FD_SC_LS__MAJ3_2%B N_B_M1009_g N_B_c_214_n N_B_M1014_g N_B_M1001_g
+ N_B_c_215_n N_B_M1015_g B N_B_c_212_n N_B_c_213_n PM_SKY130_FD_SC_LS__MAJ3_2%B
x_PM_SKY130_FD_SC_LS__MAJ3_2%C N_C_M1004_g N_C_c_256_n N_C_M1000_g N_C_M1012_g
+ N_C_c_258_n N_C_M1005_g N_C_c_259_n C N_C_c_260_n PM_SKY130_FD_SC_LS__MAJ3_2%C
x_PM_SKY130_FD_SC_LS__MAJ3_2%A N_A_c_314_n N_A_M1006_g N_A_c_315_n N_A_M1008_g
+ N_A_c_322_n N_A_c_316_n N_A_M1007_g N_A_M1011_g N_A_c_318_n N_A_c_326_n
+ N_A_c_327_n A PM_SKY130_FD_SC_LS__MAJ3_2%A
x_PM_SKY130_FD_SC_LS__MAJ3_2%VPWR N_VPWR_M1002_s N_VPWR_M1003_s N_VPWR_M1000_d
+ N_VPWR_c_393_n N_VPWR_c_394_n N_VPWR_c_395_n N_VPWR_c_396_n VPWR
+ N_VPWR_c_397_n N_VPWR_c_398_n N_VPWR_c_399_n N_VPWR_c_392_n N_VPWR_c_401_n
+ N_VPWR_c_402_n PM_SKY130_FD_SC_LS__MAJ3_2%VPWR
x_PM_SKY130_FD_SC_LS__MAJ3_2%X N_X_M1010_s N_X_M1002_d N_X_c_443_n N_X_c_444_n X
+ X X X N_X_c_445_n PM_SKY130_FD_SC_LS__MAJ3_2%X
x_PM_SKY130_FD_SC_LS__MAJ3_2%VGND N_VGND_M1010_d N_VGND_M1013_d N_VGND_M1004_d
+ N_VGND_c_477_n N_VGND_c_478_n N_VGND_c_479_n N_VGND_c_480_n VGND
+ N_VGND_c_481_n N_VGND_c_482_n N_VGND_c_483_n N_VGND_c_484_n N_VGND_c_485_n
+ N_VGND_c_486_n PM_SKY130_FD_SC_LS__MAJ3_2%VGND
cc_1 VNB N_A_87_264#_M1010_g 0.0275446f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=0.74
cc_2 VNB N_A_87_264#_M1013_g 0.0258102f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=0.74
cc_3 VNB N_A_87_264#_c_79_n 0.00315813f $X=-0.19 $Y=-0.245 $X2=2.05 $Y2=1.78
cc_4 VNB N_A_87_264#_c_80_n 0.0153736f $X=-0.19 $Y=-0.245 $X2=4.33 $Y2=0.99
cc_5 VNB N_A_87_264#_c_81_n 0.0237216f $X=-0.19 $Y=-0.245 $X2=4.495 $Y2=0.515
cc_6 VNB N_A_87_264#_c_82_n 0.00814668f $X=-0.19 $Y=-0.245 $X2=1.06 $Y2=1.485
cc_7 VNB N_A_87_264#_c_83_n 0.00446828f $X=-0.19 $Y=-0.245 $X2=2.76 $Y2=0.712
cc_8 VNB N_A_87_264#_c_84_n 0.072573f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.542
cc_9 VNB N_B_M1009_g 0.0182529f $X=-0.19 $Y=-0.245 $X2=2.47 $Y2=1.735
cc_10 VNB N_B_M1001_g 0.0193109f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_B_c_212_n 0.0387344f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=1.32
cc_12 VNB N_B_c_213_n 0.00176754f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=0.74
cc_13 VNB N_C_M1004_g 0.020459f $X=-0.19 $Y=-0.245 $X2=2.47 $Y2=1.735
cc_14 VNB N_C_c_256_n 0.0255382f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_C_M1012_g 0.0299104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_C_c_258_n 0.0353374f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_C_c_259_n 0.0202004f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.765
cc_18 VNB N_C_c_260_n 0.00433354f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.765
cc_19 VNB N_A_c_314_n 0.0260089f $X=-0.19 $Y=-0.245 $X2=2.455 $Y2=0.37
cc_20 VNB N_A_c_315_n 0.0193072f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_c_316_n 0.00137966f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_M1011_g 0.0343707f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_c_318_n 0.0375928f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=2.4
cc_24 VNB A 0.0072112f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=2.4
cc_25 VNB N_VPWR_c_392_n 0.203486f $X=-0.19 $Y=-0.245 $X2=1.06 $Y2=1.485
cc_26 VNB N_X_c_443_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_X_c_444_n 0.00429968f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.32
cc_28 VNB N_X_c_445_n 0.00139976f $X=-0.19 $Y=-0.245 $X2=2.76 $Y2=0.99
cc_29 VNB N_VGND_c_477_n 0.011316f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_478_n 0.0505285f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_479_n 0.0141402f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_480_n 0.00492322f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=1.32
cc_33 VNB N_VGND_c_481_n 0.0192531f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.765
cc_34 VNB N_VGND_c_482_n 0.042745f $X=-0.19 $Y=-0.245 $X2=2.05 $Y2=1.075
cc_35 VNB N_VGND_c_483_n 0.0299721f $X=-0.19 $Y=-0.245 $X2=4.52 $Y2=2.12
cc_36 VNB N_VGND_c_484_n 0.29124f $X=-0.19 $Y=-0.245 $X2=4.52 $Y2=2.695
cc_37 VNB N_VGND_c_485_n 0.013849f $X=-0.19 $Y=-0.245 $X2=1.255 $Y2=1.865
cc_38 VNB N_VGND_c_486_n 0.00923827f $X=-0.19 $Y=-0.245 $X2=2.76 $Y2=0.712
cc_39 VPB N_A_87_264#_c_85_n 0.017357f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=1.765
cc_40 VPB N_A_87_264#_c_86_n 0.016171f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.765
cc_41 VPB N_A_87_264#_c_87_n 0.0101982f $X=-0.19 $Y=1.66 $X2=1.965 $Y2=1.865
cc_42 VPB N_A_87_264#_c_79_n 0.00121077f $X=-0.19 $Y=1.66 $X2=2.05 $Y2=1.78
cc_43 VPB N_A_87_264#_c_89_n 0.0192421f $X=-0.19 $Y=1.66 $X2=4.52 $Y2=2.12
cc_44 VPB N_A_87_264#_c_90_n 0.0314293f $X=-0.19 $Y=1.66 $X2=4.52 $Y2=2.695
cc_45 VPB N_A_87_264#_c_82_n 0.00311528f $X=-0.19 $Y=1.66 $X2=1.06 $Y2=1.485
cc_46 VPB N_A_87_264#_c_92_n 0.00317265f $X=-0.19 $Y=1.66 $X2=2.375 $Y2=2.035
cc_47 VPB N_A_87_264#_c_84_n 0.0168368f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.542
cc_48 VPB N_B_c_214_n 0.0129339f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 VPB N_B_c_215_n 0.0127923f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_B_c_212_n 0.0210434f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=1.32
cc_51 VPB N_B_c_213_n 0.00163146f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=0.74
cc_52 VPB N_C_c_256_n 0.0249986f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_C_c_258_n 0.0297039f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_C_c_259_n 9.84389e-19 $X=-0.19 $Y=1.66 $X2=0.525 $Y2=1.765
cc_55 VPB N_C_c_260_n 0.00289875f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.765
cc_56 VPB N_A_c_314_n 0.0102776f $X=-0.19 $Y=1.66 $X2=2.455 $Y2=0.37
cc_57 VPB N_A_M1006_g 0.0100721f $X=-0.19 $Y=1.66 $X2=4.37 $Y2=1.84
cc_58 VPB N_A_c_322_n 0.139308f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_A_c_316_n 0.00900129f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_A_M1007_g 0.00874122f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=1.32
cc_61 VPB N_A_M1011_g 0.00103027f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_A_c_326_n 0.0292965f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=1.32
cc_63 VPB N_A_c_327_n 0.0289797f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_393_n 0.0112901f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_394_n 0.0644986f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_395_n 0.0169003f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=2.4
cc_67 VPB N_VPWR_c_396_n 0.00880841f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.765
cc_68 VPB N_VPWR_c_397_n 0.0194151f $X=-0.19 $Y=1.66 $X2=1.255 $Y2=1.865
cc_69 VPB N_VPWR_c_398_n 0.049034f $X=-0.19 $Y=1.66 $X2=4.355 $Y2=2.035
cc_70 VPB N_VPWR_c_399_n 0.0304171f $X=-0.19 $Y=1.66 $X2=1.075 $Y2=1.485
cc_71 VPB N_VPWR_c_392_n 0.0693167f $X=-0.19 $Y=1.66 $X2=1.06 $Y2=1.485
cc_72 VPB N_VPWR_c_401_n 0.0133423f $X=-0.19 $Y=1.66 $X2=2.595 $Y2=0.515
cc_73 VPB N_VPWR_c_402_n 0.00435574f $X=-0.19 $Y=1.66 $X2=2.375 $Y2=2.035
cc_74 VPB X 0.00195651f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=0.74
cc_75 VPB X 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_X_c_445_n 8.51199e-19 $X=-0.19 $Y=1.66 $X2=2.76 $Y2=0.99
cc_77 N_A_87_264#_c_79_n N_B_M1009_g 0.00606835f $X=2.05 $Y=1.78 $X2=0 $Y2=0
cc_78 N_A_87_264#_c_83_n N_B_M1009_g 0.0214115f $X=2.76 $Y=0.712 $X2=0 $Y2=0
cc_79 N_A_87_264#_c_79_n N_B_c_214_n 3.8425e-19 $X=2.05 $Y=1.78 $X2=0 $Y2=0
cc_80 N_A_87_264#_c_92_n N_B_c_214_n 0.0327982f $X=2.375 $Y=2.035 $X2=0 $Y2=0
cc_81 N_A_87_264#_c_80_n N_B_M1001_g 0.0112064f $X=4.33 $Y=0.99 $X2=0 $Y2=0
cc_82 N_A_87_264#_c_83_n N_B_M1001_g 0.0119906f $X=2.76 $Y=0.712 $X2=0 $Y2=0
cc_83 N_A_87_264#_c_100_p N_B_c_215_n 0.0120063f $X=4.355 $Y=2.035 $X2=0 $Y2=0
cc_84 N_A_87_264#_c_92_n N_B_c_215_n 0.0143462f $X=2.375 $Y=2.035 $X2=0 $Y2=0
cc_85 N_A_87_264#_c_80_n N_B_c_212_n 4.99319e-19 $X=4.33 $Y=0.99 $X2=0 $Y2=0
cc_86 N_A_87_264#_c_83_n N_B_c_212_n 7.90856e-19 $X=2.76 $Y=0.712 $X2=0 $Y2=0
cc_87 N_A_87_264#_c_92_n N_B_c_212_n 0.0011523f $X=2.375 $Y=2.035 $X2=0 $Y2=0
cc_88 N_A_87_264#_M1014_d N_B_c_213_n 0.00204332f $X=2.47 $Y=1.735 $X2=0 $Y2=0
cc_89 N_A_87_264#_c_79_n N_B_c_213_n 0.0408189f $X=2.05 $Y=1.78 $X2=0 $Y2=0
cc_90 N_A_87_264#_c_100_p N_B_c_213_n 0.0100458f $X=4.355 $Y=2.035 $X2=0 $Y2=0
cc_91 N_A_87_264#_c_83_n N_B_c_213_n 0.0472156f $X=2.76 $Y=0.712 $X2=0 $Y2=0
cc_92 N_A_87_264#_c_92_n N_B_c_213_n 0.0301095f $X=2.375 $Y=2.035 $X2=0 $Y2=0
cc_93 N_A_87_264#_c_80_n N_C_M1004_g 0.0151982f $X=4.33 $Y=0.99 $X2=0 $Y2=0
cc_94 N_A_87_264#_c_83_n N_C_M1004_g 0.0020622f $X=2.76 $Y=0.712 $X2=0 $Y2=0
cc_95 N_A_87_264#_c_80_n N_C_c_256_n 0.0011427f $X=4.33 $Y=0.99 $X2=0 $Y2=0
cc_96 N_A_87_264#_c_100_p N_C_c_256_n 0.0164325f $X=4.355 $Y=2.035 $X2=0 $Y2=0
cc_97 N_A_87_264#_c_92_n N_C_c_256_n 0.00297601f $X=2.375 $Y=2.035 $X2=0 $Y2=0
cc_98 N_A_87_264#_c_80_n N_C_M1012_g 0.0130655f $X=4.33 $Y=0.99 $X2=0 $Y2=0
cc_99 N_A_87_264#_c_81_n N_C_M1012_g 0.0112749f $X=4.495 $Y=0.515 $X2=0 $Y2=0
cc_100 N_A_87_264#_c_80_n N_C_c_258_n 0.0042771f $X=4.33 $Y=0.99 $X2=0 $Y2=0
cc_101 N_A_87_264#_c_100_p N_C_c_258_n 0.0125334f $X=4.355 $Y=2.035 $X2=0 $Y2=0
cc_102 N_A_87_264#_c_89_n N_C_c_258_n 0.0070094f $X=4.52 $Y=2.12 $X2=0 $Y2=0
cc_103 N_A_87_264#_c_90_n N_C_c_258_n 0.0131256f $X=4.52 $Y=2.695 $X2=0 $Y2=0
cc_104 N_A_87_264#_c_80_n N_C_c_259_n 0.0494717f $X=4.33 $Y=0.99 $X2=0 $Y2=0
cc_105 N_A_87_264#_c_100_p N_C_c_259_n 0.0257911f $X=4.355 $Y=2.035 $X2=0 $Y2=0
cc_106 N_A_87_264#_c_89_n N_C_c_259_n 0.0138934f $X=4.52 $Y=2.12 $X2=0 $Y2=0
cc_107 N_A_87_264#_c_80_n N_C_c_260_n 0.0366919f $X=4.33 $Y=0.99 $X2=0 $Y2=0
cc_108 N_A_87_264#_c_100_p N_C_c_260_n 0.0334181f $X=4.355 $Y=2.035 $X2=0 $Y2=0
cc_109 N_A_87_264#_c_87_n N_A_c_314_n 7.11218e-19 $X=1.965 $Y=1.865 $X2=-0.19
+ $Y2=-0.245
cc_110 N_A_87_264#_c_79_n N_A_c_314_n 0.0219162f $X=2.05 $Y=1.78 $X2=-0.19
+ $Y2=-0.245
cc_111 N_A_87_264#_c_82_n N_A_c_314_n 0.00445641f $X=1.06 $Y=1.485 $X2=-0.19
+ $Y2=-0.245
cc_112 N_A_87_264#_c_84_n N_A_c_314_n 0.00155618f $X=0.975 $Y=1.542 $X2=-0.19
+ $Y2=-0.245
cc_113 N_A_87_264#_c_87_n N_A_M1006_g 0.0193817f $X=1.965 $Y=1.865 $X2=0 $Y2=0
cc_114 N_A_87_264#_c_79_n N_A_M1006_g 3.73525e-19 $X=2.05 $Y=1.78 $X2=0 $Y2=0
cc_115 N_A_87_264#_c_82_n N_A_M1006_g 3.31563e-19 $X=1.06 $Y=1.485 $X2=0 $Y2=0
cc_116 N_A_87_264#_c_92_n N_A_M1006_g 0.0266137f $X=2.375 $Y=2.035 $X2=0 $Y2=0
cc_117 N_A_87_264#_c_79_n N_A_c_315_n 0.00640847f $X=2.05 $Y=1.78 $X2=0 $Y2=0
cc_118 N_A_87_264#_c_83_n N_A_c_315_n 0.0224413f $X=2.76 $Y=0.712 $X2=0 $Y2=0
cc_119 N_A_87_264#_c_92_n N_A_c_322_n 0.0132081f $X=2.375 $Y=2.035 $X2=0 $Y2=0
cc_120 N_A_87_264#_c_100_p N_A_M1007_g 0.0160299f $X=4.355 $Y=2.035 $X2=0 $Y2=0
cc_121 N_A_87_264#_c_89_n N_A_M1007_g 6.25842e-19 $X=4.52 $Y=2.12 $X2=0 $Y2=0
cc_122 N_A_87_264#_c_90_n N_A_M1007_g 0.00245895f $X=4.52 $Y=2.695 $X2=0 $Y2=0
cc_123 N_A_87_264#_c_80_n N_A_M1011_g 0.0152913f $X=4.33 $Y=0.99 $X2=0 $Y2=0
cc_124 N_A_87_264#_c_81_n N_A_M1011_g 0.00204644f $X=4.495 $Y=0.515 $X2=0 $Y2=0
cc_125 N_A_87_264#_M1013_g N_A_c_318_n 0.00312895f $X=0.945 $Y=0.74 $X2=0 $Y2=0
cc_126 N_A_87_264#_c_87_n N_A_c_318_n 0.00236155f $X=1.965 $Y=1.865 $X2=0 $Y2=0
cc_127 N_A_87_264#_c_82_n N_A_c_318_n 0.00152219f $X=1.06 $Y=1.485 $X2=0 $Y2=0
cc_128 N_A_87_264#_c_84_n N_A_c_318_n 0.0128112f $X=0.975 $Y=1.542 $X2=0 $Y2=0
cc_129 N_A_87_264#_M1013_g A 0.00166385f $X=0.945 $Y=0.74 $X2=0 $Y2=0
cc_130 N_A_87_264#_c_87_n A 0.0199019f $X=1.965 $Y=1.865 $X2=0 $Y2=0
cc_131 N_A_87_264#_c_79_n A 0.0265523f $X=2.05 $Y=1.78 $X2=0 $Y2=0
cc_132 N_A_87_264#_c_82_n A 0.0157135f $X=1.06 $Y=1.485 $X2=0 $Y2=0
cc_133 N_A_87_264#_c_84_n A 2.7436e-19 $X=0.975 $Y=1.542 $X2=0 $Y2=0
cc_134 N_A_87_264#_c_87_n N_VPWR_M1003_s 0.00762293f $X=1.965 $Y=1.865 $X2=0
+ $Y2=0
cc_135 N_A_87_264#_c_82_n N_VPWR_M1003_s 0.0025351f $X=1.06 $Y=1.485 $X2=0 $Y2=0
cc_136 N_A_87_264#_c_100_p N_VPWR_M1000_d 0.00829456f $X=4.355 $Y=2.035 $X2=0
+ $Y2=0
cc_137 N_A_87_264#_c_85_n N_VPWR_c_394_n 0.00954146f $X=0.525 $Y=1.765 $X2=0
+ $Y2=0
cc_138 N_A_87_264#_c_86_n N_VPWR_c_395_n 0.00827096f $X=0.975 $Y=1.765 $X2=0
+ $Y2=0
cc_139 N_A_87_264#_c_87_n N_VPWR_c_395_n 0.0408869f $X=1.965 $Y=1.865 $X2=0
+ $Y2=0
cc_140 N_A_87_264#_c_82_n N_VPWR_c_395_n 0.0132688f $X=1.06 $Y=1.485 $X2=0 $Y2=0
cc_141 N_A_87_264#_c_84_n N_VPWR_c_395_n 5.39386e-19 $X=0.975 $Y=1.542 $X2=0
+ $Y2=0
cc_142 N_A_87_264#_c_100_p N_VPWR_c_396_n 0.0219335f $X=4.355 $Y=2.035 $X2=0
+ $Y2=0
cc_143 N_A_87_264#_c_90_n N_VPWR_c_396_n 0.0165759f $X=4.52 $Y=2.695 $X2=0 $Y2=0
cc_144 N_A_87_264#_c_85_n N_VPWR_c_397_n 0.00411612f $X=0.525 $Y=1.765 $X2=0
+ $Y2=0
cc_145 N_A_87_264#_c_86_n N_VPWR_c_397_n 0.00445602f $X=0.975 $Y=1.765 $X2=0
+ $Y2=0
cc_146 N_A_87_264#_c_92_n N_VPWR_c_398_n 0.0176311f $X=2.375 $Y=2.035 $X2=0
+ $Y2=0
cc_147 N_A_87_264#_c_90_n N_VPWR_c_399_n 0.0097982f $X=4.52 $Y=2.695 $X2=0 $Y2=0
cc_148 N_A_87_264#_c_85_n N_VPWR_c_392_n 0.00751088f $X=0.525 $Y=1.765 $X2=0
+ $Y2=0
cc_149 N_A_87_264#_c_86_n N_VPWR_c_392_n 0.00861719f $X=0.975 $Y=1.765 $X2=0
+ $Y2=0
cc_150 N_A_87_264#_c_90_n N_VPWR_c_392_n 0.0111907f $X=4.52 $Y=2.695 $X2=0 $Y2=0
cc_151 N_A_87_264#_c_92_n N_VPWR_c_392_n 0.0225398f $X=2.375 $Y=2.035 $X2=0
+ $Y2=0
cc_152 N_A_87_264#_M1010_g N_X_c_443_n 0.0081896f $X=0.515 $Y=0.74 $X2=0 $Y2=0
cc_153 N_A_87_264#_M1013_g N_X_c_443_n 0.00783249f $X=0.945 $Y=0.74 $X2=0 $Y2=0
cc_154 N_A_87_264#_M1010_g N_X_c_444_n 0.00215589f $X=0.515 $Y=0.74 $X2=0 $Y2=0
cc_155 N_A_87_264#_M1013_g N_X_c_444_n 0.00717489f $X=0.945 $Y=0.74 $X2=0 $Y2=0
cc_156 N_A_87_264#_c_84_n N_X_c_444_n 0.00239209f $X=0.975 $Y=1.542 $X2=0 $Y2=0
cc_157 N_A_87_264#_c_85_n X 0.00240464f $X=0.525 $Y=1.765 $X2=0 $Y2=0
cc_158 N_A_87_264#_c_86_n X 0.0038841f $X=0.975 $Y=1.765 $X2=0 $Y2=0
cc_159 N_A_87_264#_c_82_n X 0.00739958f $X=1.06 $Y=1.485 $X2=0 $Y2=0
cc_160 N_A_87_264#_c_84_n X 0.00822959f $X=0.975 $Y=1.542 $X2=0 $Y2=0
cc_161 N_A_87_264#_c_85_n X 0.0130738f $X=0.525 $Y=1.765 $X2=0 $Y2=0
cc_162 N_A_87_264#_c_86_n X 0.0146975f $X=0.975 $Y=1.765 $X2=0 $Y2=0
cc_163 N_A_87_264#_M1010_g N_X_c_445_n 0.00963174f $X=0.515 $Y=0.74 $X2=0 $Y2=0
cc_164 N_A_87_264#_c_85_n N_X_c_445_n 0.0030228f $X=0.525 $Y=1.765 $X2=0 $Y2=0
cc_165 N_A_87_264#_M1013_g N_X_c_445_n 0.00298176f $X=0.945 $Y=0.74 $X2=0 $Y2=0
cc_166 N_A_87_264#_c_82_n N_X_c_445_n 0.0292292f $X=1.06 $Y=1.485 $X2=0 $Y2=0
cc_167 N_A_87_264#_c_84_n N_X_c_445_n 0.033069f $X=0.975 $Y=1.542 $X2=0 $Y2=0
cc_168 N_A_87_264#_c_79_n A_393_368# 3.70148e-19 $X=2.05 $Y=1.78 $X2=-0.19
+ $Y2=-0.245
cc_169 N_A_87_264#_c_92_n A_393_368# 0.0149642f $X=2.375 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_170 N_A_87_264#_c_100_p A_584_347# 0.014957f $X=4.355 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_171 N_A_87_264#_c_100_p A_790_368# 0.00818206f $X=4.355 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_172 N_A_87_264#_c_80_n N_VGND_M1004_d 0.00817304f $X=4.33 $Y=0.99 $X2=0 $Y2=0
cc_173 N_A_87_264#_M1010_g N_VGND_c_478_n 0.00646793f $X=0.515 $Y=0.74 $X2=0
+ $Y2=0
cc_174 N_A_87_264#_M1013_g N_VGND_c_479_n 0.00552888f $X=0.945 $Y=0.74 $X2=0
+ $Y2=0
cc_175 N_A_87_264#_c_82_n N_VGND_c_479_n 0.00986737f $X=1.06 $Y=1.485 $X2=0
+ $Y2=0
cc_176 N_A_87_264#_c_83_n N_VGND_c_479_n 0.0576083f $X=2.76 $Y=0.712 $X2=0 $Y2=0
cc_177 N_A_87_264#_c_84_n N_VGND_c_479_n 0.00109081f $X=0.975 $Y=1.542 $X2=0
+ $Y2=0
cc_178 N_A_87_264#_c_80_n N_VGND_c_480_n 0.0251177f $X=4.33 $Y=0.99 $X2=0 $Y2=0
cc_179 N_A_87_264#_c_81_n N_VGND_c_480_n 0.0107976f $X=4.495 $Y=0.515 $X2=0
+ $Y2=0
cc_180 N_A_87_264#_c_83_n N_VGND_c_480_n 0.00980679f $X=2.76 $Y=0.712 $X2=0
+ $Y2=0
cc_181 N_A_87_264#_M1010_g N_VGND_c_481_n 0.00422942f $X=0.515 $Y=0.74 $X2=0
+ $Y2=0
cc_182 N_A_87_264#_M1013_g N_VGND_c_481_n 0.00434272f $X=0.945 $Y=0.74 $X2=0
+ $Y2=0
cc_183 N_A_87_264#_c_83_n N_VGND_c_482_n 0.0345112f $X=2.76 $Y=0.712 $X2=0 $Y2=0
cc_184 N_A_87_264#_c_81_n N_VGND_c_483_n 0.0145639f $X=4.495 $Y=0.515 $X2=0
+ $Y2=0
cc_185 N_A_87_264#_M1010_g N_VGND_c_484_n 0.00787322f $X=0.515 $Y=0.74 $X2=0
+ $Y2=0
cc_186 N_A_87_264#_M1013_g N_VGND_c_484_n 0.00825283f $X=0.945 $Y=0.74 $X2=0
+ $Y2=0
cc_187 N_A_87_264#_c_81_n N_VGND_c_484_n 0.0119984f $X=4.495 $Y=0.515 $X2=0
+ $Y2=0
cc_188 N_A_87_264#_c_83_n N_VGND_c_484_n 0.0280173f $X=2.76 $Y=0.712 $X2=0 $Y2=0
cc_189 N_A_87_264#_c_79_n A_413_74# 4.41425e-19 $X=2.05 $Y=1.78 $X2=-0.19
+ $Y2=-0.245
cc_190 N_A_87_264#_c_83_n A_413_74# 0.00517808f $X=2.76 $Y=0.712 $X2=-0.19
+ $Y2=-0.245
cc_191 N_A_87_264#_c_80_n A_577_74# 0.0155294f $X=4.33 $Y=0.99 $X2=-0.19
+ $Y2=-0.245
cc_192 N_A_87_264#_c_80_n A_793_74# 0.00632546f $X=4.33 $Y=0.99 $X2=-0.19
+ $Y2=-0.245
cc_193 N_B_M1001_g N_C_M1004_g 0.0375136f $X=2.81 $Y=0.74 $X2=0 $Y2=0
cc_194 N_B_c_215_n N_C_c_256_n 0.0481751f $X=2.845 $Y=1.66 $X2=0 $Y2=0
cc_195 N_B_c_212_n N_C_c_256_n 0.0215943f $X=2.81 $Y=1.41 $X2=0 $Y2=0
cc_196 N_B_c_213_n N_C_c_256_n 0.00212676f $X=2.81 $Y=1.41 $X2=0 $Y2=0
cc_197 N_B_c_215_n N_C_c_260_n 3.05774e-19 $X=2.845 $Y=1.66 $X2=0 $Y2=0
cc_198 N_B_c_212_n N_C_c_260_n 0.00149111f $X=2.81 $Y=1.41 $X2=0 $Y2=0
cc_199 N_B_c_213_n N_C_c_260_n 0.0314385f $X=2.81 $Y=1.41 $X2=0 $Y2=0
cc_200 N_B_c_214_n N_A_c_314_n 0.0036509f $X=2.395 $Y=1.66 $X2=-0.19 $Y2=-0.245
cc_201 N_B_c_212_n N_A_c_314_n 0.0392774f $X=2.81 $Y=1.41 $X2=-0.19 $Y2=-0.245
cc_202 N_B_c_213_n N_A_c_314_n 6.77874e-19 $X=2.81 $Y=1.41 $X2=-0.19 $Y2=-0.245
cc_203 N_B_c_214_n N_A_M1006_g 0.0358626f $X=2.395 $Y=1.66 $X2=0 $Y2=0
cc_204 N_B_M1009_g N_A_c_315_n 0.0355006f $X=2.38 $Y=0.74 $X2=0 $Y2=0
cc_205 N_B_c_214_n N_A_c_322_n 0.00969102f $X=2.395 $Y=1.66 $X2=0 $Y2=0
cc_206 N_B_c_215_n N_A_c_322_n 0.0103438f $X=2.845 $Y=1.66 $X2=0 $Y2=0
cc_207 N_B_c_214_n N_VPWR_c_392_n 9.39239e-19 $X=2.395 $Y=1.66 $X2=0 $Y2=0
cc_208 N_B_c_215_n N_VPWR_c_392_n 9.39239e-19 $X=2.845 $Y=1.66 $X2=0 $Y2=0
cc_209 N_B_M1001_g N_VGND_c_480_n 0.00153831f $X=2.81 $Y=0.74 $X2=0 $Y2=0
cc_210 N_B_M1009_g N_VGND_c_482_n 0.00291649f $X=2.38 $Y=0.74 $X2=0 $Y2=0
cc_211 N_B_M1001_g N_VGND_c_482_n 0.00433162f $X=2.81 $Y=0.74 $X2=0 $Y2=0
cc_212 N_B_M1009_g N_VGND_c_484_n 0.00358831f $X=2.38 $Y=0.74 $X2=0 $Y2=0
cc_213 N_B_M1001_g N_VGND_c_484_n 0.00818163f $X=2.81 $Y=0.74 $X2=0 $Y2=0
cc_214 N_C_c_256_n N_A_c_322_n 0.0104164f $X=3.305 $Y=1.66 $X2=0 $Y2=0
cc_215 N_C_c_256_n N_A_c_316_n 0.00369026f $X=3.305 $Y=1.66 $X2=0 $Y2=0
cc_216 N_C_c_258_n N_A_c_316_n 0.0407404f $X=4.295 $Y=1.765 $X2=0 $Y2=0
cc_217 N_C_c_259_n N_A_c_316_n 0.0044568f $X=4.37 $Y=1.465 $X2=0 $Y2=0
cc_218 N_C_c_260_n N_A_c_316_n 0.00419048f $X=3.38 $Y=1.41 $X2=0 $Y2=0
cc_219 N_C_c_256_n N_A_M1007_g 0.0205934f $X=3.305 $Y=1.66 $X2=0 $Y2=0
cc_220 N_C_c_258_n N_A_M1007_g 0.0517799f $X=4.295 $Y=1.765 $X2=0 $Y2=0
cc_221 N_C_c_260_n N_A_M1007_g 4.44044e-19 $X=3.38 $Y=1.41 $X2=0 $Y2=0
cc_222 N_C_M1004_g N_A_M1011_g 0.027073f $X=3.29 $Y=0.74 $X2=0 $Y2=0
cc_223 N_C_c_256_n N_A_M1011_g 0.0163516f $X=3.305 $Y=1.66 $X2=0 $Y2=0
cc_224 N_C_M1012_g N_A_M1011_g 0.0407404f $X=4.28 $Y=0.74 $X2=0 $Y2=0
cc_225 N_C_c_259_n N_A_M1011_g 0.0120146f $X=4.37 $Y=1.465 $X2=0 $Y2=0
cc_226 N_C_c_260_n N_A_M1011_g 0.00200531f $X=3.38 $Y=1.41 $X2=0 $Y2=0
cc_227 N_C_c_258_n N_A_c_327_n 0.00281763f $X=4.295 $Y=1.765 $X2=0 $Y2=0
cc_228 N_C_c_260_n N_VPWR_M1000_d 0.00233213f $X=3.38 $Y=1.41 $X2=0 $Y2=0
cc_229 N_C_c_256_n N_VPWR_c_396_n 0.0155631f $X=3.305 $Y=1.66 $X2=0 $Y2=0
cc_230 N_C_c_258_n N_VPWR_c_396_n 0.00216473f $X=4.295 $Y=1.765 $X2=0 $Y2=0
cc_231 N_C_c_258_n N_VPWR_c_399_n 0.00481995f $X=4.295 $Y=1.765 $X2=0 $Y2=0
cc_232 N_C_c_256_n N_VPWR_c_392_n 9.39239e-19 $X=3.305 $Y=1.66 $X2=0 $Y2=0
cc_233 N_C_c_258_n N_VPWR_c_392_n 0.00508379f $X=4.295 $Y=1.765 $X2=0 $Y2=0
cc_234 N_C_M1004_g N_VGND_c_480_n 0.0164979f $X=3.29 $Y=0.74 $X2=0 $Y2=0
cc_235 N_C_M1012_g N_VGND_c_480_n 0.00149046f $X=4.28 $Y=0.74 $X2=0 $Y2=0
cc_236 N_C_M1004_g N_VGND_c_482_n 0.00383152f $X=3.29 $Y=0.74 $X2=0 $Y2=0
cc_237 N_C_M1012_g N_VGND_c_483_n 0.00434272f $X=4.28 $Y=0.74 $X2=0 $Y2=0
cc_238 N_C_M1004_g N_VGND_c_484_n 0.00758084f $X=3.29 $Y=0.74 $X2=0 $Y2=0
cc_239 N_C_M1012_g N_VGND_c_484_n 0.0082472f $X=4.28 $Y=0.74 $X2=0 $Y2=0
cc_240 N_A_M1006_g N_VPWR_c_395_n 0.00428685f $X=1.89 $Y=2.34 $X2=0 $Y2=0
cc_241 N_A_c_326_n N_VPWR_c_395_n 0.0143412f $X=1.89 $Y=3.15 $X2=0 $Y2=0
cc_242 N_A_c_322_n N_VPWR_c_396_n 0.0206374f $X=3.785 $Y=3.15 $X2=0 $Y2=0
cc_243 N_A_M1007_g N_VPWR_c_396_n 0.0120759f $X=3.875 $Y=2.34 $X2=0 $Y2=0
cc_244 N_A_c_327_n N_VPWR_c_396_n 0.0133659f $X=3.875 $Y=3.15 $X2=0 $Y2=0
cc_245 N_A_c_326_n N_VPWR_c_398_n 0.0507819f $X=1.89 $Y=3.15 $X2=0 $Y2=0
cc_246 N_A_c_327_n N_VPWR_c_399_n 0.00580471f $X=3.875 $Y=3.15 $X2=0 $Y2=0
cc_247 N_A_c_322_n N_VPWR_c_392_n 0.0525554f $X=3.785 $Y=3.15 $X2=0 $Y2=0
cc_248 N_A_c_326_n N_VPWR_c_392_n 0.0126101f $X=1.89 $Y=3.15 $X2=0 $Y2=0
cc_249 N_A_c_327_n N_VPWR_c_392_n 0.0112834f $X=3.875 $Y=3.15 $X2=0 $Y2=0
cc_250 N_A_c_315_n N_VGND_c_479_n 0.0187277f $X=1.99 $Y=1.22 $X2=0 $Y2=0
cc_251 N_A_c_318_n N_VGND_c_479_n 0.00232901f $X=1.8 $Y=1.385 $X2=0 $Y2=0
cc_252 A N_VGND_c_479_n 0.0288088f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_253 N_A_M1011_g N_VGND_c_480_n 0.0157197f $X=3.89 $Y=0.74 $X2=0 $Y2=0
cc_254 N_A_c_315_n N_VGND_c_482_n 0.00348254f $X=1.99 $Y=1.22 $X2=0 $Y2=0
cc_255 N_A_M1011_g N_VGND_c_483_n 0.00383152f $X=3.89 $Y=0.74 $X2=0 $Y2=0
cc_256 N_A_c_315_n N_VGND_c_484_n 0.00547229f $X=1.99 $Y=1.22 $X2=0 $Y2=0
cc_257 N_A_M1011_g N_VGND_c_484_n 0.0075725f $X=3.89 $Y=0.74 $X2=0 $Y2=0
cc_258 N_VPWR_c_394_n X 0.0887573f $X=0.3 $Y=1.985 $X2=0 $Y2=0
cc_259 N_VPWR_c_395_n X 0.0335865f $X=1.205 $Y=2.285 $X2=0 $Y2=0
cc_260 N_VPWR_c_397_n X 0.0158009f $X=1.085 $Y=3.33 $X2=0 $Y2=0
cc_261 N_VPWR_c_392_n X 0.0129424f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_262 N_X_c_443_n N_VGND_c_478_n 0.0308798f $X=0.73 $Y=0.515 $X2=0 $Y2=0
cc_263 N_X_c_443_n N_VGND_c_479_n 0.0245818f $X=0.73 $Y=0.515 $X2=0 $Y2=0
cc_264 N_X_c_443_n N_VGND_c_481_n 0.0149085f $X=0.73 $Y=0.515 $X2=0 $Y2=0
cc_265 N_X_c_443_n N_VGND_c_484_n 0.0122037f $X=0.73 $Y=0.515 $X2=0 $Y2=0
