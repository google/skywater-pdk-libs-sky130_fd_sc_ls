* NGSPICE file created from sky130_fd_sc_ls__dlrbp_1.ext - technology: sky130A

.subckt sky130_fd_sc_ls__dlrbp_1 D GATE RESET_B VGND VNB VPB VPWR Q Q_N
M1000 Q a_823_98# VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=1.30975e+12p ps=1.109e+07u
M1001 VGND D a_27_142# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1002 VGND a_226_104# a_353_98# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.59e+11p ps=2.18e+06u
M1003 Q a_823_98# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=2.0626e+12p ps=1.529e+07u
M1004 a_753_508# a_353_98# a_642_392# VPB phighvt w=420000u l=150000u
+  ad=2.121e+11p pd=1.85e+06u as=3.528e+11p ps=2.81e+06u
M1005 VGND a_823_98# a_775_124# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1006 VPWR a_823_98# a_753_508# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_571_80# a_27_142# VGND VNB nshort w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1008 a_642_392# a_353_98# a_571_80# VNB nshort w=640000u l=150000u
+  ad=2.692e+11p pd=2.3e+06u as=0p ps=0u
M1009 a_823_98# a_642_392# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.64e+11p pd=2.89e+06u as=0p ps=0u
M1010 a_642_392# a_226_104# a_564_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.4e+11p ps=2.48e+06u
M1011 VPWR a_823_98# a_1342_74# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=2.478e+11p ps=2.27e+06u
M1012 VGND a_823_98# a_1342_74# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1013 Q_N a_1342_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=0p ps=0u
M1014 VPWR a_226_104# a_353_98# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=2.478e+11p ps=2.27e+06u
M1015 a_775_124# a_226_104# a_642_392# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_226_104# GATE VGND VNB nshort w=740000u l=150000u
+  ad=2.701e+11p pd=2.21e+06u as=0p ps=0u
M1017 VGND RESET_B a_1051_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=1.776e+11p ps=1.96e+06u
M1018 a_226_104# GATE VPWR VPB phighvt w=840000u l=150000u
+  ad=3.066e+11p pd=2.41e+06u as=0p ps=0u
M1019 a_1051_74# a_642_392# a_823_98# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1020 Q_N a_1342_74# VGND VNB nshort w=740000u l=150000u
+  ad=2.738e+11p pd=2.22e+06u as=0p ps=0u
M1021 VPWR D a_27_142# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=2.478e+11p ps=2.27e+06u
M1022 a_564_392# a_27_142# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VPWR RESET_B a_823_98# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

