* File: sky130_fd_sc_ls__decap_4.pex.spice
* Created: Fri Aug 28 13:11:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__DECAP_4%VGND 1 9 12 13 16 17 19 21 24 26 30 40
r28 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r29 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r30 34 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r31 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r32 31 36 6.87129 $w=1.7e-07 $l=4.28e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=0.427
+ $Y2=0
r33 31 33 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=1.2
+ $Y2=0
r34 30 39 3.92207 $w=1.7e-07 $l=2.47e-07 $layer=LI1_cond $X=1.425 $Y=0 $X2=1.672
+ $Y2=0
r35 30 33 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=1.425 $Y=0 $X2=1.2
+ $Y2=0
r36 26 34 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=1.2
+ $Y2=0
r37 26 37 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=0.72
+ $Y2=0
r38 24 25 7.54852 $w=6.13e-07 $l=1.65e-07 $layer=LI1_cond $X=0.547 $Y=0.55
+ $X2=0.547 $Y2=0.715
r39 19 39 3.25516 $w=2.55e-07 $l=1.56844e-07 $layer=LI1_cond $X=1.552 $Y=0.085
+ $X2=1.672 $Y2=0
r40 19 21 21.0151 $w=2.53e-07 $l=4.65e-07 $layer=LI1_cond $X=1.552 $Y=0.085
+ $X2=1.552 $Y2=0.55
r41 16 25 32.4989 $w=2.48e-07 $l=7.05e-07 $layer=LI1_cond $X=0.73 $Y=1.42
+ $X2=0.73 $Y2=0.715
r42 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.69
+ $Y=1.42 $X2=0.69 $Y2=1.42
r43 13 24 2.76168 $w=6.13e-07 $l=1.42e-07 $layer=LI1_cond $X=0.547 $Y=0.408
+ $X2=0.547 $Y2=0.55
r44 12 36 3.29116 $w=6.15e-07 $l=1.56844e-07 $layer=LI1_cond $X=0.547 $Y=0.085
+ $X2=0.427 $Y2=0
r45 12 13 6.28184 $w=6.13e-07 $l=3.23e-07 $layer=LI1_cond $X=0.547 $Y=0.085
+ $X2=0.547 $Y2=0.408
r46 10 17 57.7274 $w=3.95e-07 $l=4.1e-07 $layer=POLY_cond $X=0.657 $Y=1.83
+ $X2=0.657 $Y2=1.42
r47 9 10 51.8833 $w=1e-06 $l=6.3e-07 $layer=POLY_cond $X=0.96 $Y=2.46 $X2=0.96
+ $Y2=1.83
r48 1 24 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.46
+ $Y=0.425 $X2=0.325 $Y2=0.55
r49 1 21 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=1.46
+ $Y=0.425 $X2=1.595 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_LS__DECAP_4%VPWR 1 8 10 13 15 19 20 22 26 37 40
r27 38 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r28 37 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r29 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r30 35 37 9.02691 $w=6.69e-07 $l=4.95e-07 $layer=LI1_cond $X=1.492 $Y=2.835
+ $X2=1.492 $Y2=3.33
r31 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r32 30 33 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r33 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r34 27 32 3.88906 $w=1.7e-07 $l=2.45e-07 $layer=LI1_cond $X=0.49 $Y=3.33
+ $X2=0.245 $Y2=3.33
r35 27 29 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=0.49 $Y=3.33
+ $X2=0.72 $Y2=3.33
r36 26 37 9.02406 $w=1.7e-07 $l=4.27e-07 $layer=LI1_cond $X=1.065 $Y=3.33
+ $X2=1.492 $Y2=3.33
r37 26 29 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.065 $Y=3.33
+ $X2=0.72 $Y2=3.33
r38 22 38 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=1.2 $Y2=3.33
r39 22 30 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=0.72 $Y2=3.33
r40 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.23
+ $Y=1.415 $X2=1.23 $Y2=1.415
r41 17 35 8.02051 $w=6.69e-07 $l=3.75545e-07 $layer=LI1_cond $X=1.19 $Y=2.67
+ $X2=1.492 $Y2=2.835
r42 17 19 57.8526 $w=2.48e-07 $l=1.255e-06 $layer=LI1_cond $X=1.19 $Y=2.67
+ $X2=1.19 $Y2=1.415
r43 13 32 3.25411 $w=2.5e-07 $l=1.56844e-07 $layer=LI1_cond $X=0.365 $Y=3.245
+ $X2=0.245 $Y2=3.33
r44 13 15 18.9001 $w=2.48e-07 $l=4.1e-07 $layer=LI1_cond $X=0.365 $Y=3.245
+ $X2=0.365 $Y2=2.835
r45 11 20 52.0954 $w=3.95e-07 $l=3.7e-07 $layer=POLY_cond $X=1.262 $Y=1.045
+ $X2=1.262 $Y2=1.415
r46 10 11 19.5871 $w=3.95e-07 $l=4.05e-07 $layer=POLY_cond $X=1.262 $Y=0.64
+ $X2=1.262 $Y2=1.045
r47 8 10 19.1703 $w=8.1e-07 $l=3.02e-07 $layer=POLY_cond $X=0.96 $Y=0.64
+ $X2=1.262 $Y2=0.64
r48 1 35 600 $w=1.7e-07 $l=9.4008e-07 $layer=licon1_PDIFF $count=1 $X=1.46
+ $Y=1.96 $X2=1.595 $Y2=2.835
r49 1 15 600 $w=1.7e-07 $l=9.44722e-07 $layer=licon1_PDIFF $count=1 $X=1.46
+ $Y=1.96 $X2=0.325 $Y2=2.835
.ends

