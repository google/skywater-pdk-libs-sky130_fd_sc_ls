* File: sky130_fd_sc_ls__xor3_2.spice
* Created: Wed Sep  2 11:31:22 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__xor3_2.pex.spice"
.subckt sky130_fd_sc_ls__xor3_2  VNB VPB A B C VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* C	C
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1017 N_VGND_M1017_d N_A_83_289#_M1017_g N_A_27_134#_M1017_s VNB NSHORT L=0.15
+ W=0.64 AD=0.34745 AS=0.1824 PD=1.81 PS=1.85 NRD=91.476 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75002.9 A=0.096 P=1.58 MULT=1
MM1022 N_A_83_289#_M1022_d N_A_M1022_g N_VGND_M1017_d VNB NSHORT L=0.15 W=0.64
+ AD=0.169862 AS=0.34745 PD=1.275 PS=1.81 NRD=0 NRS=91.476 M=1 R=4.26667
+ SA=75001 SB=75002 A=0.096 P=1.58 MULT=1
MM1019 N_A_416_113#_M1019_d N_B_M1019_g N_A_83_289#_M1022_d VNB NSHORT L=0.15
+ W=0.64 AD=0.125283 AS=0.169862 PD=1.19547 PS=1.275 NRD=0 NRS=47.808 M=1
+ R=4.26667 SA=75001.5 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1008 N_A_27_134#_M1008_d N_A_440_315#_M1008_g N_A_416_113#_M1019_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.125326 AS=0.082217 PD=0.919245 PS=0.784528 NRD=19.992
+ NRS=20.712 M=1 R=2.8 SA=75002.2 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1016 N_A_372_419#_M1016_d N_B_M1016_g N_A_27_134#_M1008_d VNB NSHORT L=0.15
+ W=0.64 AD=0.1495 AS=0.190974 PD=1.14 PS=1.40075 NRD=15.468 NRS=31.872 M=1
+ R=4.26667 SA=75002 SB=75000.9 A=0.096 P=1.58 MULT=1
MM1020 N_A_83_289#_M1020_d N_A_440_315#_M1020_g N_A_372_419#_M1016_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.2848 AS=0.1495 PD=2.17 PS=1.14 NRD=31.872 NRS=15.468 M=1
+ R=4.26667 SA=75002.6 SB=75000.4 A=0.096 P=1.58 MULT=1
MM1009 N_VGND_M1009_d N_B_M1009_g N_A_440_315#_M1009_s VNB NSHORT L=0.15 W=0.74
+ AD=0.46725 AS=0.2035 PD=2.88 PS=2.03 NRD=93.468 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.4 A=0.111 P=1.78 MULT=1
MM1004 N_A_1195_424#_M1004_d N_A_1162_379#_M1004_g N_A_372_419#_M1004_s VNB
+ NSHORT L=0.15 W=0.64 AD=0.169775 AS=0.176 PD=1.24 PS=1.83 NRD=47.808 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75000.9 A=0.096 P=1.58 MULT=1
MM1007 N_A_416_113#_M1007_d N_C_M1007_g N_A_1195_424#_M1004_d VNB NSHORT L=0.15
+ W=0.64 AD=0.2144 AS=0.169775 PD=1.95 PS=1.24 NRD=4.68 NRS=0 M=1 R=4.26667
+ SA=75000.8 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1018 N_VGND_M1018_d N_C_M1018_g N_A_1162_379#_M1018_s VNB NSHORT L=0.15 W=0.42
+ AD=0.106521 AS=0.1197 PD=0.847241 PS=1.41 NRD=22.848 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1018_d N_A_1195_424#_M1002_g N_X_M1002_s VNB NSHORT L=0.15 W=0.74
+ AD=0.187679 AS=0.1036 PD=1.49276 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1014 N_VGND_M1014_d N_A_1195_424#_M1014_g N_X_M1002_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1000 N_VPWR_M1000_d N_A_83_289#_M1000_g N_A_27_134#_M1000_s VPB PHIGHVT L=0.15
+ W=1 AD=0.2225 AS=0.295 PD=1.445 PS=2.59 NRD=11.8003 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75002.4 A=0.15 P=2.3 MULT=1
MM1006 N_A_83_289#_M1006_d N_A_M1006_g N_VPWR_M1000_d VPB PHIGHVT L=0.15 W=1
+ AD=0.201413 AS=0.2225 PD=1.50543 PS=1.445 NRD=1.9503 NRS=20.685 M=1 R=6.66667
+ SA=75000.8 SB=75001.9 A=0.15 P=2.3 MULT=1
MM1012 N_A_372_419#_M1012_d N_B_M1012_g N_A_83_289#_M1006_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.159032 AS=0.169187 PD=1.35649 PS=1.26457 NRD=3.5066 NRS=22.261 M=1
+ R=5.6 SA=75001.3 SB=75001.6 A=0.126 P=1.98 MULT=1
MM1015 N_A_27_134#_M1015_d N_A_440_315#_M1015_g N_A_372_419#_M1012_d VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.096 AS=0.121168 PD=0.94 PS=1.03351 NRD=3.0732 NRS=18.4589
+ M=1 R=4.26667 SA=75001.9 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1021 N_A_416_113#_M1021_d N_B_M1021_g N_A_27_134#_M1015_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.132065 AS=0.096 PD=1.05946 PS=0.94 NRD=30.7714 NRS=3.0732 M=1
+ R=4.26667 SA=75002.3 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1003 N_A_83_289#_M1003_d N_A_440_315#_M1003_g N_A_416_113#_M1021_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.5544 AS=0.173335 PD=3 PS=1.39054 NRD=75.0373 NRS=2.3443 M=1
+ R=5.6 SA=75002.2 SB=75000.6 A=0.126 P=1.98 MULT=1
MM1011 N_VPWR_M1011_d N_B_M1011_g N_A_440_315#_M1011_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.3304 PD=2.83 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1013 N_A_1195_424#_M1013_d N_A_1162_379#_M1013_g N_A_416_113#_M1013_s VPB
+ PHIGHVT L=0.15 W=0.84 AD=0.2562 AS=0.2478 PD=1.45 PS=2.27 NRD=75.0373
+ NRS=2.3443 M=1 R=5.6 SA=75000.2 SB=75001 A=0.126 P=1.98 MULT=1
MM1023 N_A_372_419#_M1023_d N_C_M1023_g N_A_1195_424#_M1013_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.2478 AS=0.2562 PD=2.27 PS=1.45 NRD=2.3443 NRS=2.3443 M=1 R=5.6
+ SA=75001 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1010 N_VPWR_M1010_d N_C_M1010_g N_A_1162_379#_M1010_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.287709 AS=0.24 PD=1.35636 PS=2.03 NRD=30.0031 NRS=27.6982 M=1
+ R=4.26667 SA=75000.3 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1001 N_X_M1001_d N_A_1195_424#_M1001_g N_VPWR_M1010_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.503491 PD=1.42 PS=2.37364 NRD=1.7533 NRS=65.0691 M=1
+ R=7.46667 SA=75000.9 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1005 N_X_M1001_d N_A_1195_424#_M1005_g N_VPWR_M1005_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.4 SB=75000.2 A=0.168 P=2.54 MULT=1
DX24_noxref VNB VPB NWDIODE A=18.5628 P=23.68
c_106 VNB 0 1.49322e-19 $X=0 $Y=0
c_195 VPB 0 3.36481e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_ls__xor3_2.pxi.spice"
*
.ends
*
*
