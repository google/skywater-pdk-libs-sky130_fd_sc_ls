* NGSPICE file created from sky130_fd_sc_ls__a211oi_1.ext - technology: sky130A

.subckt sky130_fd_sc_ls__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
M1000 a_71_368# A1 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=6.44e+11p pd=5.63e+06u as=4.368e+11p ps=3.02e+06u
M1001 Y A1 a_159_74# VNB nshort w=740000u l=150000u
+  ad=4.847e+11p pd=4.27e+06u as=1.554e+11p ps=1.9e+06u
M1002 a_354_368# B1 a_71_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=3.696e+11p pd=2.9e+06u as=0p ps=0u
M1003 a_159_74# A2 VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=4.847e+11p ps=4.27e+06u
M1004 VGND B1 Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR A2 a_71_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y C1 a_354_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=3.08e+11p pd=2.79e+06u as=0p ps=0u
M1007 Y C1 VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

