* File: sky130_fd_sc_ls__nor3_1.spice
* Created: Wed Sep  2 11:14:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__nor3_1.pex.spice"
.subckt sky130_fd_sc_ls__nor3_1  VNB VPB A B C VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* C	C
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1004 N_Y_M1004_d N_A_M1004_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.74 AD=0.1036
+ AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0.396 M=1 R=4.93333 SA=75000.2 SB=75001.1
+ A=0.111 P=1.78 MULT=1
MM1005 N_VGND_M1005_d N_B_M1005_g N_Y_M1004_d VNB NSHORT L=0.15 W=0.74 AD=0.1295
+ AS=0.1036 PD=1.09 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6 SB=75000.7
+ A=0.111 P=1.78 MULT=1
MM1002 N_Y_M1002_d N_C_M1002_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.74 AD=0.2109
+ AS=0.1295 PD=2.05 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.1 SB=75000.2
+ A=0.111 P=1.78 MULT=1
MM1003 A_114_368# N_A_M1003_g N_VPWR_M1003_s VPB PHIGHVT L=0.15 W=1.12 AD=0.1512
+ AS=0.3192 PD=1.39 PS=2.81 NRD=14.0658 NRS=1.7533 M=1 R=7.46667 SA=75000.2
+ SB=75001.1 A=0.168 P=2.54 MULT=1
MM1001 A_198_368# N_B_M1001_g A_114_368# VPB PHIGHVT L=0.15 W=1.12 AD=0.2016
+ AS=0.1512 PD=1.48 PS=1.39 NRD=21.9852 NRS=14.0658 M=1 R=7.46667 SA=75000.6
+ SB=75000.7 A=0.168 P=2.54 MULT=1
MM1000 N_Y_M1000_d N_C_M1000_g A_198_368# VPB PHIGHVT L=0.15 W=1.12 AD=0.3192
+ AS=0.2016 PD=2.81 PS=1.48 NRD=1.7533 NRS=21.9852 M=1 R=7.46667 SA=75001.1
+ SB=75000.2 A=0.168 P=2.54 MULT=1
DX6_noxref VNB VPB NWDIODE A=4.278 P=8.32
*
.include "sky130_fd_sc_ls__nor3_1.pxi.spice"
*
.ends
*
*
