* File: sky130_fd_sc_ls__a21boi_4.pxi.spice
* Created: Fri Aug 28 12:51:10 2020
* 
x_PM_SKY130_FD_SC_LS__A21BOI_4%A1 N_A1_c_125_n N_A1_M1002_g N_A1_M1000_g
+ N_A1_c_126_n N_A1_M1016_g N_A1_M1003_g N_A1_c_127_n N_A1_M1017_g N_A1_M1004_g
+ N_A1_c_128_n N_A1_M1022_g N_A1_M1013_g A1 A1 A1 A1 N_A1_c_124_n
+ PM_SKY130_FD_SC_LS__A21BOI_4%A1
x_PM_SKY130_FD_SC_LS__A21BOI_4%A2 N_A2_M1010_g N_A2_c_206_n N_A2_M1008_g
+ N_A2_M1011_g N_A2_c_207_n N_A2_M1015_g N_A2_M1019_g N_A2_c_208_n N_A2_M1021_g
+ N_A2_M1026_g N_A2_c_209_n N_A2_M1024_g A2 A2 A2 N_A2_c_205_n
+ PM_SKY130_FD_SC_LS__A21BOI_4%A2
x_PM_SKY130_FD_SC_LS__A21BOI_4%A_803_323# N_A_803_323#_M1001_d
+ N_A_803_323#_M1007_d N_A_803_323#_c_299_n N_A_803_323#_M1005_g
+ N_A_803_323#_c_286_n N_A_803_323#_c_287_n N_A_803_323#_c_288_n
+ N_A_803_323#_M1006_g N_A_803_323#_M1012_g N_A_803_323#_c_290_n
+ N_A_803_323#_M1018_g N_A_803_323#_c_303_n N_A_803_323#_M1009_g
+ N_A_803_323#_M1020_g N_A_803_323#_c_304_n N_A_803_323#_M1025_g
+ N_A_803_323#_M1023_g N_A_803_323#_c_294_n N_A_803_323#_c_295_n
+ N_A_803_323#_c_306_n N_A_803_323#_c_296_n N_A_803_323#_c_307_n
+ N_A_803_323#_c_308_n N_A_803_323#_c_297_n N_A_803_323#_c_309_n
+ N_A_803_323#_c_298_n PM_SKY130_FD_SC_LS__A21BOI_4%A_803_323#
x_PM_SKY130_FD_SC_LS__A21BOI_4%B1_N N_B1_N_M1001_g N_B1_N_c_413_n N_B1_N_M1007_g
+ N_B1_N_c_414_n N_B1_N_M1014_g B1_N B1_N B1_N N_B1_N_c_412_n
+ PM_SKY130_FD_SC_LS__A21BOI_4%B1_N
x_PM_SKY130_FD_SC_LS__A21BOI_4%A_31_368# N_A_31_368#_M1002_d N_A_31_368#_M1016_d
+ N_A_31_368#_M1022_d N_A_31_368#_M1015_s N_A_31_368#_M1024_s
+ N_A_31_368#_M1006_s N_A_31_368#_M1025_s N_A_31_368#_c_447_n
+ N_A_31_368#_c_448_n N_A_31_368#_c_460_n N_A_31_368#_c_449_n
+ N_A_31_368#_c_466_n N_A_31_368#_c_450_n N_A_31_368#_c_475_n
+ N_A_31_368#_c_451_n N_A_31_368#_c_483_n N_A_31_368#_c_487_n
+ N_A_31_368#_c_488_n N_A_31_368#_c_452_n N_A_31_368#_c_453_n
+ N_A_31_368#_c_498_n N_A_31_368#_c_454_n N_A_31_368#_c_455_n
+ N_A_31_368#_c_471_n N_A_31_368#_c_456_n N_A_31_368#_c_492_n
+ N_A_31_368#_c_457_n PM_SKY130_FD_SC_LS__A21BOI_4%A_31_368#
x_PM_SKY130_FD_SC_LS__A21BOI_4%VPWR N_VPWR_M1002_s N_VPWR_M1017_s N_VPWR_M1008_d
+ N_VPWR_M1021_d N_VPWR_M1007_s N_VPWR_M1014_s N_VPWR_c_556_n N_VPWR_c_557_n
+ N_VPWR_c_558_n N_VPWR_c_559_n N_VPWR_c_560_n N_VPWR_c_561_n N_VPWR_c_562_n
+ N_VPWR_c_563_n N_VPWR_c_564_n N_VPWR_c_565_n N_VPWR_c_566_n N_VPWR_c_567_n
+ N_VPWR_c_568_n N_VPWR_c_569_n VPWR N_VPWR_c_570_n N_VPWR_c_571_n
+ N_VPWR_c_572_n N_VPWR_c_555_n N_VPWR_c_574_n N_VPWR_c_575_n
+ PM_SKY130_FD_SC_LS__A21BOI_4%VPWR
x_PM_SKY130_FD_SC_LS__A21BOI_4%Y N_Y_M1000_s N_Y_M1004_s N_Y_M1012_d N_Y_M1020_d
+ N_Y_M1005_d N_Y_M1009_d N_Y_c_675_n N_Y_c_665_n N_Y_c_666_n N_Y_c_710_n
+ N_Y_c_667_n N_Y_c_673_n N_Y_c_668_n N_Y_c_674_n N_Y_c_728_n N_Y_c_669_n
+ N_Y_c_670_n N_Y_c_671_n Y Y PM_SKY130_FD_SC_LS__A21BOI_4%Y
x_PM_SKY130_FD_SC_LS__A21BOI_4%A_46_74# N_A_46_74#_M1000_d N_A_46_74#_M1003_d
+ N_A_46_74#_M1013_d N_A_46_74#_M1011_s N_A_46_74#_M1026_s N_A_46_74#_c_776_n
+ N_A_46_74#_c_788_n N_A_46_74#_c_804_n N_A_46_74#_c_790_n N_A_46_74#_c_777_n
+ N_A_46_74#_c_807_n N_A_46_74#_c_778_n PM_SKY130_FD_SC_LS__A21BOI_4%A_46_74#
x_PM_SKY130_FD_SC_LS__A21BOI_4%VGND N_VGND_M1010_d N_VGND_M1019_d N_VGND_M1012_s
+ N_VGND_M1018_s N_VGND_M1023_s N_VGND_c_830_n N_VGND_c_831_n N_VGND_c_832_n
+ N_VGND_c_833_n N_VGND_c_834_n N_VGND_c_835_n N_VGND_c_836_n N_VGND_c_837_n
+ N_VGND_c_838_n N_VGND_c_839_n N_VGND_c_840_n N_VGND_c_841_n VGND
+ N_VGND_c_842_n N_VGND_c_843_n N_VGND_c_844_n N_VGND_c_845_n N_VGND_c_846_n
+ PM_SKY130_FD_SC_LS__A21BOI_4%VGND
cc_1 VNB N_A1_M1000_g 0.0337982f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=0.74
cc_2 VNB N_A1_M1003_g 0.0235163f $X=-0.19 $Y=-0.245 $X2=1 $Y2=0.74
cc_3 VNB N_A1_M1004_g 0.022969f $X=-0.19 $Y=-0.245 $X2=1.43 $Y2=0.74
cc_4 VNB N_A1_M1013_g 0.0226731f $X=-0.19 $Y=-0.245 $X2=1.86 $Y2=0.74
cc_5 VNB A1 0.0153254f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_6 VNB N_A1_c_124_n 0.0774836f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=1.557
cc_7 VNB N_A2_M1010_g 0.0222064f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_8 VNB N_A2_M1011_g 0.0218258f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_9 VNB N_A2_M1019_g 0.0218258f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=2.4
cc_10 VNB N_A2_M1026_g 0.0262254f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=2.4
cc_11 VNB A2 0.00232653f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_12 VNB N_A2_c_205_n 0.0720397f $X=-0.19 $Y=-0.245 $X2=1.86 $Y2=1.557
cc_13 VNB N_A_803_323#_c_286_n 0.00993983f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_14 VNB N_A_803_323#_c_287_n 0.00613301f $X=-0.19 $Y=-0.245 $X2=1 $Y2=1.35
cc_15 VNB N_A_803_323#_c_288_n 0.00629408f $X=-0.19 $Y=-0.245 $X2=1 $Y2=0.74
cc_16 VNB N_A_803_323#_M1012_g 0.0345749f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=2.4
cc_17 VNB N_A_803_323#_c_290_n 0.0138f $X=-0.19 $Y=-0.245 $X2=1.43 $Y2=0.74
cc_18 VNB N_A_803_323#_M1018_g 0.0211895f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=2.4
cc_19 VNB N_A_803_323#_M1020_g 0.0217754f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_20 VNB N_A_803_323#_M1023_g 0.0218825f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.557
cc_21 VNB N_A_803_323#_c_294_n 0.00605926f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=1.515
cc_22 VNB N_A_803_323#_c_295_n 0.0677327f $X=-0.19 $Y=-0.245 $X2=1.43 $Y2=1.557
cc_23 VNB N_A_803_323#_c_296_n 0.0112317f $X=-0.19 $Y=-0.245 $X2=1.6 $Y2=1.515
cc_24 VNB N_A_803_323#_c_297_n 0.0330377f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.605
cc_25 VNB N_A_803_323#_c_298_n 0.00664811f $X=-0.19 $Y=-0.245 $X2=1.6 $Y2=1.605
cc_26 VNB N_B1_N_M1001_g 0.0401523f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_27 VNB B1_N 0.0314342f $X=-0.19 $Y=-0.245 $X2=1 $Y2=0.74
cc_28 VNB N_B1_N_c_412_n 0.0500872f $X=-0.19 $Y=-0.245 $X2=1.43 $Y2=0.74
cc_29 VNB N_VPWR_c_555_n 0.322901f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_Y_c_665_n 0.022664f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_Y_c_666_n 0.0211712f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=2.4
cc_32 VNB N_Y_c_667_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_33 VNB N_Y_c_668_n 0.00533449f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_Y_c_669_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=1.515
cc_35 VNB N_Y_c_670_n 0.0023338f $X=-0.19 $Y=-0.245 $X2=1 $Y2=1.557
cc_36 VNB N_Y_c_671_n 0.00227381f $X=-0.19 $Y=-0.245 $X2=1.43 $Y2=1.557
cc_37 VNB N_A_46_74#_c_776_n 0.00914219f $X=-0.19 $Y=-0.245 $X2=1.43 $Y2=1.35
cc_38 VNB N_A_46_74#_c_777_n 0.0370051f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_39 VNB N_A_46_74#_c_778_n 0.00481051f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.557
cc_40 VNB N_VGND_c_830_n 0.00323505f $X=-0.19 $Y=-0.245 $X2=1.43 $Y2=1.35
cc_41 VNB N_VGND_c_831_n 0.00266156f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=1.765
cc_42 VNB N_VGND_c_832_n 0.0133983f $X=-0.19 $Y=-0.245 $X2=1.86 $Y2=0.74
cc_43 VNB N_VGND_c_833_n 0.0172524f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_834_n 0.00420208f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_45 VNB N_VGND_c_835_n 0.00334323f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_836_n 0.0604496f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=1.557
cc_47 VNB N_VGND_c_837_n 0.00601569f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=1.515
cc_48 VNB N_VGND_c_838_n 0.014238f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.557
cc_49 VNB N_VGND_c_839_n 0.00601569f $X=-0.19 $Y=-0.245 $X2=1 $Y2=1.557
cc_50 VNB N_VGND_c_840_n 0.0184034f $X=-0.19 $Y=-0.245 $X2=1.26 $Y2=1.557
cc_51 VNB N_VGND_c_841_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=1.26 $Y2=1.515
cc_52 VNB N_VGND_c_842_n 0.0172524f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_843_n 0.0461117f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_844_n 0.451501f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_845_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_846_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VPB N_A1_c_125_n 0.0201401f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_58 VPB N_A1_c_126_n 0.0149968f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.765
cc_59 VPB N_A1_c_127_n 0.014996f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=1.765
cc_60 VPB N_A1_c_128_n 0.015369f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=1.765
cc_61 VPB A1 0.0165319f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.58
cc_62 VPB N_A1_c_124_n 0.0478075f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=1.557
cc_63 VPB N_A2_c_206_n 0.015369f $X=-0.19 $Y=1.66 $X2=0.57 $Y2=0.74
cc_64 VPB N_A2_c_207_n 0.0155119f $X=-0.19 $Y=1.66 $X2=1 $Y2=0.74
cc_65 VPB N_A2_c_208_n 0.0155127f $X=-0.19 $Y=1.66 $X2=1.43 $Y2=0.74
cc_66 VPB N_A2_c_209_n 0.0153123f $X=-0.19 $Y=1.66 $X2=1.86 $Y2=0.74
cc_67 VPB A2 0.00851521f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_68 VPB N_A2_c_205_n 0.0465732f $X=-0.19 $Y=1.66 $X2=1.86 $Y2=1.557
cc_69 VPB N_A_803_323#_c_299_n 0.0144998f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_A_803_323#_c_286_n 0.00675749f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_71 VPB N_A_803_323#_c_287_n 0.00369877f $X=-0.19 $Y=1.66 $X2=1 $Y2=1.35
cc_72 VPB N_A_803_323#_c_288_n 0.0177271f $X=-0.19 $Y=1.66 $X2=1 $Y2=0.74
cc_73 VPB N_A_803_323#_c_303_n 0.0145642f $X=-0.19 $Y=1.66 $X2=1.86 $Y2=1.35
cc_74 VPB N_A_803_323#_c_304_n 0.0171142f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.58
cc_75 VPB N_A_803_323#_c_295_n 0.0142886f $X=-0.19 $Y=1.66 $X2=1.43 $Y2=1.557
cc_76 VPB N_A_803_323#_c_306_n 0.00703151f $X=-0.19 $Y=1.66 $X2=1.6 $Y2=1.515
cc_77 VPB N_A_803_323#_c_307_n 0.00366357f $X=-0.19 $Y=1.66 $X2=1.86 $Y2=1.557
cc_78 VPB N_A_803_323#_c_308_n 0.00273598f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.605
cc_79 VPB N_A_803_323#_c_309_n 0.00243101f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 VPB N_B1_N_c_413_n 0.0173817f $X=-0.19 $Y=1.66 $X2=0.57 $Y2=0.74
cc_81 VPB N_B1_N_c_414_n 0.0174317f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.765
cc_82 VPB B1_N 0.0244129f $X=-0.19 $Y=1.66 $X2=1 $Y2=0.74
cc_83 VPB N_B1_N_c_412_n 0.0555178f $X=-0.19 $Y=1.66 $X2=1.43 $Y2=0.74
cc_84 VPB N_A_31_368#_c_447_n 0.00786417f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=1.765
cc_85 VPB N_A_31_368#_c_448_n 0.0345863f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=2.4
cc_86 VPB N_A_31_368#_c_449_n 0.00180921f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_87 VPB N_A_31_368#_c_450_n 0.00180921f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_A_31_368#_c_451_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.557
cc_89 VPB N_A_31_368#_c_452_n 0.0026202f $X=-0.19 $Y=1.66 $X2=1.6 $Y2=1.515
cc_90 VPB N_A_31_368#_c_453_n 0.00192911f $X=-0.19 $Y=1.66 $X2=1.6 $Y2=1.515
cc_91 VPB N_A_31_368#_c_454_n 0.00660678f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_92 VPB N_A_31_368#_c_455_n 0.0125757f $X=-0.19 $Y=1.66 $X2=1.2 $Y2=1.605
cc_93 VPB N_A_31_368#_c_456_n 0.0030519f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB N_A_31_368#_c_457_n 0.00167433f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_556_n 0.00329129f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_557_n 0.00261791f $X=-0.19 $Y=1.66 $X2=1.86 $Y2=1.35
cc_97 VPB N_VPWR_c_558_n 0.00504372f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_98 VPB N_VPWR_c_559_n 0.00769929f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_560_n 0.011866f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.557
cc_100 VPB N_VPWR_c_561_n 0.0469329f $X=-0.19 $Y=1.66 $X2=0.92 $Y2=1.515
cc_101 VPB N_VPWR_c_562_n 0.0164465f $X=-0.19 $Y=1.66 $X2=1.26 $Y2=1.557
cc_102 VPB N_VPWR_c_563_n 0.00460249f $X=-0.19 $Y=1.66 $X2=1.26 $Y2=1.515
cc_103 VPB N_VPWR_c_564_n 0.0206041f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=1.557
cc_104 VPB N_VPWR_c_565_n 0.00324402f $X=-0.19 $Y=1.66 $X2=1.43 $Y2=1.557
cc_105 VPB N_VPWR_c_566_n 0.0594566f $X=-0.19 $Y=1.66 $X2=1.6 $Y2=1.515
cc_106 VPB N_VPWR_c_567_n 0.00614127f $X=-0.19 $Y=1.66 $X2=1.6 $Y2=1.515
cc_107 VPB N_VPWR_c_568_n 0.0182909f $X=-0.19 $Y=1.66 $X2=1.86 $Y2=1.557
cc_108 VPB N_VPWR_c_569_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.605
cc_109 VPB N_VPWR_c_570_n 0.0180274f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.605
cc_110 VPB N_VPWR_c_571_n 0.0164465f $X=-0.19 $Y=1.66 $X2=1.26 $Y2=1.605
cc_111 VPB N_VPWR_c_572_n 0.0153494f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_555_n 0.110805f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_VPWR_c_574_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_VPWR_c_575_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_Y_c_666_n 0.00382854f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=2.4
cc_116 VPB N_Y_c_673_n 0.00160061f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_117 VPB N_Y_c_674_n 0.00183525f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 N_A1_M1013_g N_A2_M1010_g 0.032151f $X=1.86 $Y=0.74 $X2=0 $Y2=0
cc_119 N_A1_c_128_n N_A2_c_206_n 0.00946162f $X=1.855 $Y=1.765 $X2=0 $Y2=0
cc_120 A1 A2 0.0107734f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_121 N_A1_c_124_n A2 0.00116888f $X=1.855 $Y=1.557 $X2=0 $Y2=0
cc_122 A1 N_A2_c_205_n 0.00116888f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_123 N_A1_c_124_n N_A2_c_205_n 0.022585f $X=1.855 $Y=1.557 $X2=0 $Y2=0
cc_124 A1 N_A_31_368#_c_447_n 0.0209486f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_125 N_A1_c_125_n N_A_31_368#_c_448_n 0.00634858f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_126 N_A1_c_125_n N_A_31_368#_c_460_n 0.0126853f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_127 N_A1_c_126_n N_A_31_368#_c_460_n 0.0126853f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_128 A1 N_A_31_368#_c_460_n 0.0467841f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_129 N_A1_c_124_n N_A_31_368#_c_460_n 0.00150005f $X=1.855 $Y=1.557 $X2=0
+ $Y2=0
cc_130 N_A1_c_126_n N_A_31_368#_c_449_n 0.00554978f $X=0.955 $Y=1.765 $X2=0
+ $Y2=0
cc_131 N_A1_c_127_n N_A_31_368#_c_449_n 0.00554978f $X=1.405 $Y=1.765 $X2=0
+ $Y2=0
cc_132 N_A1_c_127_n N_A_31_368#_c_466_n 0.0126853f $X=1.405 $Y=1.765 $X2=0 $Y2=0
cc_133 N_A1_c_128_n N_A_31_368#_c_466_n 0.0167336f $X=1.855 $Y=1.765 $X2=0 $Y2=0
cc_134 A1 N_A_31_368#_c_466_n 0.0341468f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_135 N_A1_c_124_n N_A_31_368#_c_466_n 0.00150005f $X=1.855 $Y=1.557 $X2=0
+ $Y2=0
cc_136 N_A1_c_128_n N_A_31_368#_c_450_n 0.00576879f $X=1.855 $Y=1.765 $X2=0
+ $Y2=0
cc_137 A1 N_A_31_368#_c_471_n 0.0148009f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_138 N_A1_c_124_n N_A_31_368#_c_471_n 0.00104296f $X=1.855 $Y=1.557 $X2=0
+ $Y2=0
cc_139 N_A1_c_128_n N_A_31_368#_c_456_n 0.00262483f $X=1.855 $Y=1.765 $X2=0
+ $Y2=0
cc_140 N_A1_c_125_n N_VPWR_c_556_n 0.0141019f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_141 N_A1_c_126_n N_VPWR_c_556_n 0.0110266f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_142 N_A1_c_127_n N_VPWR_c_556_n 5.35985e-19 $X=1.405 $Y=1.765 $X2=0 $Y2=0
cc_143 N_A1_c_126_n N_VPWR_c_557_n 5.35985e-19 $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_144 N_A1_c_127_n N_VPWR_c_557_n 0.0110266f $X=1.405 $Y=1.765 $X2=0 $Y2=0
cc_145 N_A1_c_128_n N_VPWR_c_557_n 0.0110266f $X=1.855 $Y=1.765 $X2=0 $Y2=0
cc_146 N_A1_c_128_n N_VPWR_c_558_n 5.37805e-19 $X=1.855 $Y=1.765 $X2=0 $Y2=0
cc_147 N_A1_c_128_n N_VPWR_c_562_n 0.00413917f $X=1.855 $Y=1.765 $X2=0 $Y2=0
cc_148 N_A1_c_125_n N_VPWR_c_570_n 0.00413917f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_149 N_A1_c_126_n N_VPWR_c_571_n 0.00413917f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_150 N_A1_c_127_n N_VPWR_c_571_n 0.00413917f $X=1.405 $Y=1.765 $X2=0 $Y2=0
cc_151 N_A1_c_125_n N_VPWR_c_555_n 0.00821221f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_152 N_A1_c_126_n N_VPWR_c_555_n 0.00817726f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_153 N_A1_c_127_n N_VPWR_c_555_n 0.00817726f $X=1.405 $Y=1.765 $X2=0 $Y2=0
cc_154 N_A1_c_128_n N_VPWR_c_555_n 0.0081781f $X=1.855 $Y=1.765 $X2=0 $Y2=0
cc_155 N_A1_M1003_g N_Y_c_675_n 0.00924655f $X=1 $Y=0.74 $X2=0 $Y2=0
cc_156 N_A1_M1004_g N_Y_c_675_n 0.00971392f $X=1.43 $Y=0.74 $X2=0 $Y2=0
cc_157 A1 N_Y_c_675_n 0.0148057f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_158 N_A1_c_124_n N_Y_c_675_n 0.00193117f $X=1.855 $Y=1.557 $X2=0 $Y2=0
cc_159 N_A1_M1013_g N_Y_c_665_n 0.0134911f $X=1.86 $Y=0.74 $X2=0 $Y2=0
cc_160 N_A1_c_124_n N_Y_c_665_n 4.21656e-19 $X=1.855 $Y=1.557 $X2=0 $Y2=0
cc_161 N_A1_M1003_g N_Y_c_670_n 0.00516369f $X=1 $Y=0.74 $X2=0 $Y2=0
cc_162 N_A1_M1004_g N_Y_c_670_n 6.39903e-19 $X=1.43 $Y=0.74 $X2=0 $Y2=0
cc_163 A1 N_Y_c_670_n 0.0129494f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_164 N_A1_c_124_n N_Y_c_670_n 0.00231456f $X=1.855 $Y=1.557 $X2=0 $Y2=0
cc_165 N_A1_M1003_g N_Y_c_671_n 0.00127276f $X=1 $Y=0.74 $X2=0 $Y2=0
cc_166 N_A1_M1004_g N_Y_c_671_n 0.00903278f $X=1.43 $Y=0.74 $X2=0 $Y2=0
cc_167 N_A1_M1013_g N_Y_c_671_n 0.00849971f $X=1.86 $Y=0.74 $X2=0 $Y2=0
cc_168 A1 N_Y_c_671_n 0.0257396f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_169 N_A1_c_124_n N_Y_c_671_n 0.00253745f $X=1.855 $Y=1.557 $X2=0 $Y2=0
cc_170 N_A1_M1000_g N_A_46_74#_c_776_n 0.0128206f $X=0.57 $Y=0.74 $X2=0 $Y2=0
cc_171 N_A1_M1003_g N_A_46_74#_c_776_n 0.010203f $X=1 $Y=0.74 $X2=0 $Y2=0
cc_172 N_A1_M1004_g N_A_46_74#_c_776_n 0.0101343f $X=1.43 $Y=0.74 $X2=0 $Y2=0
cc_173 N_A1_M1013_g N_A_46_74#_c_776_n 0.0129923f $X=1.86 $Y=0.74 $X2=0 $Y2=0
cc_174 N_A1_M1000_g N_A_46_74#_c_777_n 0.0100735f $X=0.57 $Y=0.74 $X2=0 $Y2=0
cc_175 N_A1_M1003_g N_A_46_74#_c_777_n 9.10353e-19 $X=1 $Y=0.74 $X2=0 $Y2=0
cc_176 A1 N_A_46_74#_c_777_n 0.0190532f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_177 N_A1_c_124_n N_A_46_74#_c_777_n 0.00216428f $X=1.855 $Y=1.557 $X2=0 $Y2=0
cc_178 N_A1_M1013_g N_VGND_c_830_n 7.0229e-19 $X=1.86 $Y=0.74 $X2=0 $Y2=0
cc_179 N_A1_M1000_g N_VGND_c_836_n 0.00291626f $X=0.57 $Y=0.74 $X2=0 $Y2=0
cc_180 N_A1_M1003_g N_VGND_c_836_n 0.00291649f $X=1 $Y=0.74 $X2=0 $Y2=0
cc_181 N_A1_M1004_g N_VGND_c_836_n 0.00291649f $X=1.43 $Y=0.74 $X2=0 $Y2=0
cc_182 N_A1_M1013_g N_VGND_c_836_n 0.00291649f $X=1.86 $Y=0.74 $X2=0 $Y2=0
cc_183 N_A1_M1000_g N_VGND_c_844_n 0.00362992f $X=0.57 $Y=0.74 $X2=0 $Y2=0
cc_184 N_A1_M1003_g N_VGND_c_844_n 0.00358174f $X=1 $Y=0.74 $X2=0 $Y2=0
cc_185 N_A1_M1004_g N_VGND_c_844_n 0.00358174f $X=1.43 $Y=0.74 $X2=0 $Y2=0
cc_186 N_A1_M1013_g N_VGND_c_844_n 0.00359219f $X=1.86 $Y=0.74 $X2=0 $Y2=0
cc_187 N_A2_c_209_n N_A_803_323#_c_299_n 0.0118912f $X=3.655 $Y=1.765 $X2=0
+ $Y2=0
cc_188 N_A2_c_205_n N_A_803_323#_c_287_n 0.00618447f $X=3.58 $Y=1.557 $X2=0
+ $Y2=0
cc_189 N_A2_c_206_n N_A_31_368#_c_450_n 0.0039133f $X=2.305 $Y=1.765 $X2=0 $Y2=0
cc_190 N_A2_c_206_n N_A_31_368#_c_475_n 0.0167336f $X=2.305 $Y=1.765 $X2=0 $Y2=0
cc_191 N_A2_c_207_n N_A_31_368#_c_475_n 0.0120074f $X=2.755 $Y=1.765 $X2=0 $Y2=0
cc_192 A2 N_A_31_368#_c_475_n 0.0300859f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_193 N_A2_c_205_n N_A_31_368#_c_475_n 0.00130859f $X=3.58 $Y=1.557 $X2=0 $Y2=0
cc_194 N_A2_c_206_n N_A_31_368#_c_451_n 6.69308e-19 $X=2.305 $Y=1.765 $X2=0
+ $Y2=0
cc_195 N_A2_c_207_n N_A_31_368#_c_451_n 0.0105452f $X=2.755 $Y=1.765 $X2=0 $Y2=0
cc_196 N_A2_c_208_n N_A_31_368#_c_451_n 0.0103431f $X=3.205 $Y=1.765 $X2=0 $Y2=0
cc_197 N_A2_c_209_n N_A_31_368#_c_451_n 6.45594e-19 $X=3.655 $Y=1.765 $X2=0
+ $Y2=0
cc_198 N_A2_c_208_n N_A_31_368#_c_483_n 0.0119563f $X=3.205 $Y=1.765 $X2=0 $Y2=0
cc_199 N_A2_c_209_n N_A_31_368#_c_483_n 0.0120074f $X=3.655 $Y=1.765 $X2=0 $Y2=0
cc_200 A2 N_A_31_368#_c_483_n 0.0386622f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_201 N_A2_c_205_n N_A_31_368#_c_483_n 0.00130859f $X=3.58 $Y=1.557 $X2=0 $Y2=0
cc_202 N_A2_c_209_n N_A_31_368#_c_487_n 8.76854e-19 $X=3.655 $Y=1.765 $X2=0
+ $Y2=0
cc_203 N_A2_c_208_n N_A_31_368#_c_488_n 6.23807e-19 $X=3.205 $Y=1.765 $X2=0
+ $Y2=0
cc_204 N_A2_c_209_n N_A_31_368#_c_488_n 0.00919154f $X=3.655 $Y=1.765 $X2=0
+ $Y2=0
cc_205 N_A2_c_209_n N_A_31_368#_c_453_n 0.0032261f $X=3.655 $Y=1.765 $X2=0 $Y2=0
cc_206 N_A2_c_206_n N_A_31_368#_c_456_n 0.00262483f $X=2.305 $Y=1.765 $X2=0
+ $Y2=0
cc_207 N_A2_c_207_n N_A_31_368#_c_492_n 4.27055e-19 $X=2.755 $Y=1.765 $X2=0
+ $Y2=0
cc_208 N_A2_c_208_n N_A_31_368#_c_492_n 4.27055e-19 $X=3.205 $Y=1.765 $X2=0
+ $Y2=0
cc_209 A2 N_A_31_368#_c_492_n 0.0233234f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_210 N_A2_c_205_n N_A_31_368#_c_492_n 0.00144162f $X=3.58 $Y=1.557 $X2=0 $Y2=0
cc_211 N_A2_c_206_n N_VPWR_c_557_n 5.35985e-19 $X=2.305 $Y=1.765 $X2=0 $Y2=0
cc_212 N_A2_c_206_n N_VPWR_c_558_n 0.0106464f $X=2.305 $Y=1.765 $X2=0 $Y2=0
cc_213 N_A2_c_207_n N_VPWR_c_558_n 0.00526215f $X=2.755 $Y=1.765 $X2=0 $Y2=0
cc_214 N_A2_c_208_n N_VPWR_c_559_n 0.00486623f $X=3.205 $Y=1.765 $X2=0 $Y2=0
cc_215 N_A2_c_209_n N_VPWR_c_559_n 0.00331651f $X=3.655 $Y=1.765 $X2=0 $Y2=0
cc_216 N_A2_c_206_n N_VPWR_c_562_n 0.00413917f $X=2.305 $Y=1.765 $X2=0 $Y2=0
cc_217 N_A2_c_207_n N_VPWR_c_564_n 0.00445602f $X=2.755 $Y=1.765 $X2=0 $Y2=0
cc_218 N_A2_c_208_n N_VPWR_c_564_n 0.00445602f $X=3.205 $Y=1.765 $X2=0 $Y2=0
cc_219 N_A2_c_209_n N_VPWR_c_566_n 0.0044313f $X=3.655 $Y=1.765 $X2=0 $Y2=0
cc_220 N_A2_c_206_n N_VPWR_c_555_n 0.0081781f $X=2.305 $Y=1.765 $X2=0 $Y2=0
cc_221 N_A2_c_207_n N_VPWR_c_555_n 0.00857589f $X=2.755 $Y=1.765 $X2=0 $Y2=0
cc_222 N_A2_c_208_n N_VPWR_c_555_n 0.00857589f $X=3.205 $Y=1.765 $X2=0 $Y2=0
cc_223 N_A2_c_209_n N_VPWR_c_555_n 0.00853445f $X=3.655 $Y=1.765 $X2=0 $Y2=0
cc_224 N_A2_M1010_g N_Y_c_665_n 0.0149909f $X=2.29 $Y=0.74 $X2=0 $Y2=0
cc_225 N_A2_M1011_g N_Y_c_665_n 0.0104926f $X=2.72 $Y=0.74 $X2=0 $Y2=0
cc_226 N_A2_M1019_g N_Y_c_665_n 0.0104926f $X=3.15 $Y=0.74 $X2=0 $Y2=0
cc_227 N_A2_M1026_g N_Y_c_665_n 0.0125331f $X=3.58 $Y=0.74 $X2=0 $Y2=0
cc_228 A2 N_Y_c_665_n 0.100241f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_229 N_A2_c_205_n N_Y_c_665_n 0.00960894f $X=3.58 $Y=1.557 $X2=0 $Y2=0
cc_230 N_A2_M1026_g N_Y_c_666_n 0.0031715f $X=3.58 $Y=0.74 $X2=0 $Y2=0
cc_231 N_A2_c_209_n N_Y_c_666_n 7.34383e-19 $X=3.655 $Y=1.765 $X2=0 $Y2=0
cc_232 A2 N_Y_c_666_n 0.0231776f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_233 N_A2_c_205_n N_Y_c_666_n 0.00596607f $X=3.58 $Y=1.557 $X2=0 $Y2=0
cc_234 N_A2_M1010_g N_Y_c_671_n 9.08556e-19 $X=2.29 $Y=0.74 $X2=0 $Y2=0
cc_235 N_A2_M1010_g N_A_46_74#_c_776_n 8.36418e-19 $X=2.29 $Y=0.74 $X2=0 $Y2=0
cc_236 N_A2_M1010_g N_A_46_74#_c_788_n 0.0097843f $X=2.29 $Y=0.74 $X2=0 $Y2=0
cc_237 N_A2_M1011_g N_A_46_74#_c_788_n 0.0097843f $X=2.72 $Y=0.74 $X2=0 $Y2=0
cc_238 N_A2_M1019_g N_A_46_74#_c_790_n 0.0097843f $X=3.15 $Y=0.74 $X2=0 $Y2=0
cc_239 N_A2_M1026_g N_A_46_74#_c_790_n 0.0097843f $X=3.58 $Y=0.74 $X2=0 $Y2=0
cc_240 N_A2_M1010_g N_VGND_c_830_n 0.00676719f $X=2.29 $Y=0.74 $X2=0 $Y2=0
cc_241 N_A2_M1011_g N_VGND_c_830_n 0.00779025f $X=2.72 $Y=0.74 $X2=0 $Y2=0
cc_242 N_A2_M1019_g N_VGND_c_830_n 8.17314e-19 $X=3.15 $Y=0.74 $X2=0 $Y2=0
cc_243 N_A2_M1011_g N_VGND_c_831_n 8.17314e-19 $X=2.72 $Y=0.74 $X2=0 $Y2=0
cc_244 N_A2_M1019_g N_VGND_c_831_n 0.00779025f $X=3.15 $Y=0.74 $X2=0 $Y2=0
cc_245 N_A2_M1026_g N_VGND_c_831_n 0.00903439f $X=3.58 $Y=0.74 $X2=0 $Y2=0
cc_246 N_A2_M1026_g N_VGND_c_832_n 0.00461687f $X=3.58 $Y=0.74 $X2=0 $Y2=0
cc_247 N_A2_M1010_g N_VGND_c_836_n 0.00281141f $X=2.29 $Y=0.74 $X2=0 $Y2=0
cc_248 N_A2_M1011_g N_VGND_c_838_n 0.00281141f $X=2.72 $Y=0.74 $X2=0 $Y2=0
cc_249 N_A2_M1019_g N_VGND_c_838_n 0.00281141f $X=3.15 $Y=0.74 $X2=0 $Y2=0
cc_250 N_A2_M1026_g N_VGND_c_840_n 0.00281141f $X=3.58 $Y=0.74 $X2=0 $Y2=0
cc_251 N_A2_M1010_g N_VGND_c_844_n 0.00365164f $X=2.29 $Y=0.74 $X2=0 $Y2=0
cc_252 N_A2_M1011_g N_VGND_c_844_n 0.00365066f $X=2.72 $Y=0.74 $X2=0 $Y2=0
cc_253 N_A2_M1019_g N_VGND_c_844_n 0.00365066f $X=3.15 $Y=0.74 $X2=0 $Y2=0
cc_254 N_A2_M1026_g N_VGND_c_844_n 0.00370065f $X=3.58 $Y=0.74 $X2=0 $Y2=0
cc_255 N_A_803_323#_M1023_g N_B1_N_M1001_g 0.0148997f $X=5.85 $Y=0.74 $X2=0
+ $Y2=0
cc_256 N_A_803_323#_c_296_n N_B1_N_M1001_g 0.0166978f $X=6.4 $Y=1.235 $X2=0
+ $Y2=0
cc_257 N_A_803_323#_c_297_n N_B1_N_M1001_g 0.00321641f $X=6.495 $Y=0.515 $X2=0
+ $Y2=0
cc_258 N_A_803_323#_c_298_n N_B1_N_M1001_g 0.00733653f $X=6.11 $Y=1.4 $X2=0
+ $Y2=0
cc_259 N_A_803_323#_c_307_n N_B1_N_c_413_n 0.0109952f $X=6.535 $Y=2.075 $X2=0
+ $Y2=0
cc_260 N_A_803_323#_c_309_n N_B1_N_c_413_n 9.00673e-19 $X=6.65 $Y=2.265 $X2=0
+ $Y2=0
cc_261 N_A_803_323#_c_307_n N_B1_N_c_414_n 0.00407678f $X=6.535 $Y=2.075 $X2=0
+ $Y2=0
cc_262 N_A_803_323#_c_309_n N_B1_N_c_414_n 0.0107901f $X=6.65 $Y=2.265 $X2=0
+ $Y2=0
cc_263 N_A_803_323#_c_306_n B1_N 0.0134675f $X=6.11 $Y=1.99 $X2=0 $Y2=0
cc_264 N_A_803_323#_c_296_n B1_N 0.0245195f $X=6.4 $Y=1.235 $X2=0 $Y2=0
cc_265 N_A_803_323#_c_307_n B1_N 0.0356589f $X=6.535 $Y=2.075 $X2=0 $Y2=0
cc_266 N_A_803_323#_c_298_n B1_N 0.0141734f $X=6.11 $Y=1.4 $X2=0 $Y2=0
cc_267 N_A_803_323#_c_295_n N_B1_N_c_412_n 0.0151702f $X=5.76 $Y=1.485 $X2=0
+ $Y2=0
cc_268 N_A_803_323#_c_306_n N_B1_N_c_412_n 0.0106445f $X=6.11 $Y=1.99 $X2=0
+ $Y2=0
cc_269 N_A_803_323#_c_296_n N_B1_N_c_412_n 0.00807778f $X=6.4 $Y=1.235 $X2=0
+ $Y2=0
cc_270 N_A_803_323#_c_307_n N_B1_N_c_412_n 0.0154625f $X=6.535 $Y=2.075 $X2=0
+ $Y2=0
cc_271 N_A_803_323#_c_299_n N_A_31_368#_c_452_n 0.0128006f $X=4.105 $Y=1.765
+ $X2=0 $Y2=0
cc_272 N_A_803_323#_c_288_n N_A_31_368#_c_452_n 0.0128349f $X=4.555 $Y=1.765
+ $X2=0 $Y2=0
cc_273 N_A_803_323#_c_290_n N_A_31_368#_c_498_n 2.69463e-19 $X=4.915 $Y=1.575
+ $X2=0 $Y2=0
cc_274 N_A_803_323#_c_303_n N_A_31_368#_c_454_n 0.0127907f $X=5.005 $Y=1.765
+ $X2=0 $Y2=0
cc_275 N_A_803_323#_c_304_n N_A_31_368#_c_454_n 0.0137046f $X=5.455 $Y=1.765
+ $X2=0 $Y2=0
cc_276 N_A_803_323#_c_304_n N_A_31_368#_c_455_n 0.00143221f $X=5.455 $Y=1.765
+ $X2=0 $Y2=0
cc_277 N_A_803_323#_c_294_n N_A_31_368#_c_455_n 0.0234447f $X=6.025 $Y=1.485
+ $X2=0 $Y2=0
cc_278 N_A_803_323#_c_295_n N_A_31_368#_c_455_n 0.00717826f $X=5.76 $Y=1.485
+ $X2=0 $Y2=0
cc_279 N_A_803_323#_c_306_n N_A_31_368#_c_455_n 0.0127429f $X=6.11 $Y=1.99 $X2=0
+ $Y2=0
cc_280 N_A_803_323#_c_308_n N_A_31_368#_c_455_n 0.0142731f $X=6.195 $Y=2.075
+ $X2=0 $Y2=0
cc_281 N_A_803_323#_c_307_n N_VPWR_M1007_s 0.00103113f $X=6.535 $Y=2.075 $X2=0
+ $Y2=0
cc_282 N_A_803_323#_c_308_n N_VPWR_M1007_s 0.00150507f $X=6.195 $Y=2.075 $X2=0
+ $Y2=0
cc_283 N_A_803_323#_c_304_n N_VPWR_c_560_n 8.71134e-19 $X=5.455 $Y=1.765 $X2=0
+ $Y2=0
cc_284 N_A_803_323#_c_307_n N_VPWR_c_560_n 0.00896099f $X=6.535 $Y=2.075 $X2=0
+ $Y2=0
cc_285 N_A_803_323#_c_308_n N_VPWR_c_560_n 0.0144736f $X=6.195 $Y=2.075 $X2=0
+ $Y2=0
cc_286 N_A_803_323#_c_309_n N_VPWR_c_560_n 0.0251606f $X=6.65 $Y=2.265 $X2=0
+ $Y2=0
cc_287 N_A_803_323#_c_307_n N_VPWR_c_561_n 0.00430094f $X=6.535 $Y=2.075 $X2=0
+ $Y2=0
cc_288 N_A_803_323#_c_309_n N_VPWR_c_561_n 0.0543079f $X=6.65 $Y=2.265 $X2=0
+ $Y2=0
cc_289 N_A_803_323#_c_299_n N_VPWR_c_566_n 0.00278271f $X=4.105 $Y=1.765 $X2=0
+ $Y2=0
cc_290 N_A_803_323#_c_288_n N_VPWR_c_566_n 0.00278271f $X=4.555 $Y=1.765 $X2=0
+ $Y2=0
cc_291 N_A_803_323#_c_303_n N_VPWR_c_566_n 0.00278271f $X=5.005 $Y=1.765 $X2=0
+ $Y2=0
cc_292 N_A_803_323#_c_304_n N_VPWR_c_566_n 0.00278271f $X=5.455 $Y=1.765 $X2=0
+ $Y2=0
cc_293 N_A_803_323#_c_309_n N_VPWR_c_568_n 0.0123628f $X=6.65 $Y=2.265 $X2=0
+ $Y2=0
cc_294 N_A_803_323#_c_299_n N_VPWR_c_555_n 0.00353907f $X=4.105 $Y=1.765 $X2=0
+ $Y2=0
cc_295 N_A_803_323#_c_288_n N_VPWR_c_555_n 0.00353823f $X=4.555 $Y=1.765 $X2=0
+ $Y2=0
cc_296 N_A_803_323#_c_303_n N_VPWR_c_555_n 0.00353823f $X=5.005 $Y=1.765 $X2=0
+ $Y2=0
cc_297 N_A_803_323#_c_304_n N_VPWR_c_555_n 0.00358624f $X=5.455 $Y=1.765 $X2=0
+ $Y2=0
cc_298 N_A_803_323#_c_309_n N_VPWR_c_555_n 0.0101999f $X=6.65 $Y=2.265 $X2=0
+ $Y2=0
cc_299 N_A_803_323#_c_299_n N_Y_c_666_n 0.0118882f $X=4.105 $Y=1.765 $X2=0 $Y2=0
cc_300 N_A_803_323#_c_286_n N_Y_c_666_n 0.0138742f $X=4.48 $Y=1.69 $X2=0 $Y2=0
cc_301 N_A_803_323#_c_287_n N_Y_c_666_n 0.00701865f $X=4.18 $Y=1.69 $X2=0 $Y2=0
cc_302 N_A_803_323#_c_288_n N_Y_c_666_n 0.0216289f $X=4.555 $Y=1.765 $X2=0 $Y2=0
cc_303 N_A_803_323#_M1012_g N_Y_c_666_n 0.030234f $X=4.56 $Y=0.74 $X2=0 $Y2=0
cc_304 N_A_803_323#_c_290_n N_Y_c_666_n 0.00778004f $X=4.915 $Y=1.575 $X2=0
+ $Y2=0
cc_305 N_A_803_323#_M1018_g N_Y_c_666_n 0.00333031f $X=4.99 $Y=0.74 $X2=0 $Y2=0
cc_306 N_A_803_323#_c_294_n N_Y_c_666_n 0.0285716f $X=6.025 $Y=1.485 $X2=0 $Y2=0
cc_307 N_A_803_323#_c_295_n N_Y_c_666_n 0.00388253f $X=5.76 $Y=1.485 $X2=0 $Y2=0
cc_308 N_A_803_323#_c_299_n N_Y_c_710_n 0.00721451f $X=4.105 $Y=1.765 $X2=0
+ $Y2=0
cc_309 N_A_803_323#_c_288_n N_Y_c_710_n 0.0085809f $X=4.555 $Y=1.765 $X2=0 $Y2=0
cc_310 N_A_803_323#_c_303_n N_Y_c_710_n 5.86053e-19 $X=5.005 $Y=1.765 $X2=0
+ $Y2=0
cc_311 N_A_803_323#_M1012_g N_Y_c_667_n 0.0101f $X=4.56 $Y=0.74 $X2=0 $Y2=0
cc_312 N_A_803_323#_M1018_g N_Y_c_667_n 3.97481e-19 $X=4.99 $Y=0.74 $X2=0 $Y2=0
cc_313 N_A_803_323#_c_290_n N_Y_c_673_n 0.00470466f $X=4.915 $Y=1.575 $X2=0
+ $Y2=0
cc_314 N_A_803_323#_c_303_n N_Y_c_673_n 0.0120074f $X=5.005 $Y=1.765 $X2=0 $Y2=0
cc_315 N_A_803_323#_c_294_n N_Y_c_673_n 0.010734f $X=6.025 $Y=1.485 $X2=0 $Y2=0
cc_316 N_A_803_323#_c_295_n N_Y_c_673_n 4.52619e-19 $X=5.76 $Y=1.485 $X2=0 $Y2=0
cc_317 N_A_803_323#_M1018_g N_Y_c_668_n 0.0126841f $X=4.99 $Y=0.74 $X2=0 $Y2=0
cc_318 N_A_803_323#_M1020_g N_Y_c_668_n 0.0122543f $X=5.42 $Y=0.74 $X2=0 $Y2=0
cc_319 N_A_803_323#_M1023_g N_Y_c_668_n 0.00123832f $X=5.85 $Y=0.74 $X2=0 $Y2=0
cc_320 N_A_803_323#_c_294_n N_Y_c_668_n 0.0616244f $X=6.025 $Y=1.485 $X2=0 $Y2=0
cc_321 N_A_803_323#_c_295_n N_Y_c_668_n 0.00457162f $X=5.76 $Y=1.485 $X2=0 $Y2=0
cc_322 N_A_803_323#_c_303_n N_Y_c_674_n 6.83942e-19 $X=5.005 $Y=1.765 $X2=0
+ $Y2=0
cc_323 N_A_803_323#_c_304_n N_Y_c_674_n 0.00216099f $X=5.455 $Y=1.765 $X2=0
+ $Y2=0
cc_324 N_A_803_323#_c_294_n N_Y_c_674_n 0.0276944f $X=6.025 $Y=1.485 $X2=0 $Y2=0
cc_325 N_A_803_323#_c_295_n N_Y_c_674_n 0.00789892f $X=5.76 $Y=1.485 $X2=0 $Y2=0
cc_326 N_A_803_323#_c_288_n N_Y_c_728_n 5.86053e-19 $X=4.555 $Y=1.765 $X2=0
+ $Y2=0
cc_327 N_A_803_323#_c_303_n N_Y_c_728_n 0.0085809f $X=5.005 $Y=1.765 $X2=0 $Y2=0
cc_328 N_A_803_323#_c_304_n N_Y_c_728_n 0.00759832f $X=5.455 $Y=1.765 $X2=0
+ $Y2=0
cc_329 N_A_803_323#_M1018_g N_Y_c_669_n 6.3583e-19 $X=4.99 $Y=0.74 $X2=0 $Y2=0
cc_330 N_A_803_323#_M1020_g N_Y_c_669_n 0.00887299f $X=5.42 $Y=0.74 $X2=0 $Y2=0
cc_331 N_A_803_323#_M1023_g N_Y_c_669_n 3.97481e-19 $X=5.85 $Y=0.74 $X2=0 $Y2=0
cc_332 N_A_803_323#_M1012_g N_A_46_74#_c_778_n 8.70183e-19 $X=4.56 $Y=0.74 $X2=0
+ $Y2=0
cc_333 N_A_803_323#_M1012_g N_VGND_c_832_n 0.00639168f $X=4.56 $Y=0.74 $X2=0
+ $Y2=0
cc_334 N_A_803_323#_M1012_g N_VGND_c_833_n 0.00434272f $X=4.56 $Y=0.74 $X2=0
+ $Y2=0
cc_335 N_A_803_323#_M1018_g N_VGND_c_833_n 0.00383152f $X=4.99 $Y=0.74 $X2=0
+ $Y2=0
cc_336 N_A_803_323#_M1012_g N_VGND_c_834_n 5.11602e-19 $X=4.56 $Y=0.74 $X2=0
+ $Y2=0
cc_337 N_A_803_323#_M1018_g N_VGND_c_834_n 0.00953461f $X=4.99 $Y=0.74 $X2=0
+ $Y2=0
cc_338 N_A_803_323#_M1020_g N_VGND_c_834_n 0.00192252f $X=5.42 $Y=0.74 $X2=0
+ $Y2=0
cc_339 N_A_803_323#_M1020_g N_VGND_c_835_n 5.60973e-19 $X=5.42 $Y=0.74 $X2=0
+ $Y2=0
cc_340 N_A_803_323#_M1023_g N_VGND_c_835_n 0.0110422f $X=5.85 $Y=0.74 $X2=0
+ $Y2=0
cc_341 N_A_803_323#_c_294_n N_VGND_c_835_n 0.00478652f $X=6.025 $Y=1.485 $X2=0
+ $Y2=0
cc_342 N_A_803_323#_c_296_n N_VGND_c_835_n 0.00212635f $X=6.4 $Y=1.235 $X2=0
+ $Y2=0
cc_343 N_A_803_323#_c_297_n N_VGND_c_835_n 0.0244016f $X=6.495 $Y=0.515 $X2=0
+ $Y2=0
cc_344 N_A_803_323#_c_298_n N_VGND_c_835_n 0.0135092f $X=6.11 $Y=1.4 $X2=0 $Y2=0
cc_345 N_A_803_323#_M1020_g N_VGND_c_842_n 0.00434272f $X=5.42 $Y=0.74 $X2=0
+ $Y2=0
cc_346 N_A_803_323#_M1023_g N_VGND_c_842_n 0.00383152f $X=5.85 $Y=0.74 $X2=0
+ $Y2=0
cc_347 N_A_803_323#_c_297_n N_VGND_c_843_n 0.0115122f $X=6.495 $Y=0.515 $X2=0
+ $Y2=0
cc_348 N_A_803_323#_M1012_g N_VGND_c_844_n 0.00825283f $X=4.56 $Y=0.74 $X2=0
+ $Y2=0
cc_349 N_A_803_323#_M1018_g N_VGND_c_844_n 0.0075754f $X=4.99 $Y=0.74 $X2=0
+ $Y2=0
cc_350 N_A_803_323#_M1020_g N_VGND_c_844_n 0.00820284f $X=5.42 $Y=0.74 $X2=0
+ $Y2=0
cc_351 N_A_803_323#_M1023_g N_VGND_c_844_n 0.0075754f $X=5.85 $Y=0.74 $X2=0
+ $Y2=0
cc_352 N_A_803_323#_c_297_n N_VGND_c_844_n 0.0095288f $X=6.495 $Y=0.515 $X2=0
+ $Y2=0
cc_353 N_B1_N_c_413_n N_A_31_368#_c_454_n 5.75404e-19 $X=6.425 $Y=2.045 $X2=0
+ $Y2=0
cc_354 N_B1_N_c_413_n N_A_31_368#_c_455_n 0.00383047f $X=6.425 $Y=2.045 $X2=0
+ $Y2=0
cc_355 N_B1_N_c_412_n N_A_31_368#_c_455_n 4.62469e-19 $X=6.53 $Y=1.655 $X2=0
+ $Y2=0
cc_356 N_B1_N_c_413_n N_VPWR_c_560_n 0.0112901f $X=6.425 $Y=2.045 $X2=0 $Y2=0
cc_357 N_B1_N_c_414_n N_VPWR_c_560_n 5.8666e-19 $X=6.875 $Y=2.045 $X2=0 $Y2=0
cc_358 N_B1_N_c_414_n N_VPWR_c_561_n 0.00990078f $X=6.875 $Y=2.045 $X2=0 $Y2=0
cc_359 B1_N N_VPWR_c_561_n 0.0154871f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_360 N_B1_N_c_413_n N_VPWR_c_568_n 0.00413917f $X=6.425 $Y=2.045 $X2=0 $Y2=0
cc_361 N_B1_N_c_414_n N_VPWR_c_568_n 0.00445602f $X=6.875 $Y=2.045 $X2=0 $Y2=0
cc_362 N_B1_N_c_413_n N_VPWR_c_555_n 0.00817726f $X=6.425 $Y=2.045 $X2=0 $Y2=0
cc_363 N_B1_N_c_414_n N_VPWR_c_555_n 0.00862391f $X=6.875 $Y=2.045 $X2=0 $Y2=0
cc_364 N_B1_N_M1001_g N_VGND_c_835_n 0.0137119f $X=6.28 $Y=0.74 $X2=0 $Y2=0
cc_365 N_B1_N_M1001_g N_VGND_c_843_n 0.00383152f $X=6.28 $Y=0.74 $X2=0 $Y2=0
cc_366 N_B1_N_M1001_g N_VGND_c_844_n 0.00762539f $X=6.28 $Y=0.74 $X2=0 $Y2=0
cc_367 N_A_31_368#_c_460_n N_VPWR_M1002_s 0.00359365f $X=1.095 $Y=2.035
+ $X2=-0.19 $Y2=1.66
cc_368 N_A_31_368#_c_466_n N_VPWR_M1017_s 0.00359365f $X=1.995 $Y=2.035 $X2=0
+ $Y2=0
cc_369 N_A_31_368#_c_475_n N_VPWR_M1008_d 0.00384138f $X=2.815 $Y=2.035 $X2=0
+ $Y2=0
cc_370 N_A_31_368#_c_483_n N_VPWR_M1021_d 0.00408911f $X=3.715 $Y=2.035 $X2=0
+ $Y2=0
cc_371 N_A_31_368#_c_448_n N_VPWR_c_556_n 0.0462948f $X=0.28 $Y=2.815 $X2=0
+ $Y2=0
cc_372 N_A_31_368#_c_460_n N_VPWR_c_556_n 0.0171813f $X=1.095 $Y=2.035 $X2=0
+ $Y2=0
cc_373 N_A_31_368#_c_449_n N_VPWR_c_556_n 0.0449718f $X=1.18 $Y=2.815 $X2=0
+ $Y2=0
cc_374 N_A_31_368#_c_449_n N_VPWR_c_557_n 0.0449718f $X=1.18 $Y=2.815 $X2=0
+ $Y2=0
cc_375 N_A_31_368#_c_466_n N_VPWR_c_557_n 0.0171813f $X=1.995 $Y=2.035 $X2=0
+ $Y2=0
cc_376 N_A_31_368#_c_450_n N_VPWR_c_557_n 0.0449718f $X=2.08 $Y=2.4 $X2=0 $Y2=0
cc_377 N_A_31_368#_c_450_n N_VPWR_c_558_n 0.0440249f $X=2.08 $Y=2.4 $X2=0 $Y2=0
cc_378 N_A_31_368#_c_475_n N_VPWR_c_558_n 0.0154248f $X=2.815 $Y=2.035 $X2=0
+ $Y2=0
cc_379 N_A_31_368#_c_451_n N_VPWR_c_558_n 0.0462948f $X=2.98 $Y=2.815 $X2=0
+ $Y2=0
cc_380 N_A_31_368#_c_451_n N_VPWR_c_559_n 0.0449718f $X=2.98 $Y=2.815 $X2=0
+ $Y2=0
cc_381 N_A_31_368#_c_483_n N_VPWR_c_559_n 0.0136682f $X=3.715 $Y=2.035 $X2=0
+ $Y2=0
cc_382 N_A_31_368#_c_488_n N_VPWR_c_559_n 0.0395235f $X=3.88 $Y=2.815 $X2=0
+ $Y2=0
cc_383 N_A_31_368#_c_453_n N_VPWR_c_559_n 0.0119328f $X=3.995 $Y=2.99 $X2=0
+ $Y2=0
cc_384 N_A_31_368#_c_454_n N_VPWR_c_560_n 0.0139f $X=5.565 $Y=2.99 $X2=0 $Y2=0
cc_385 N_A_31_368#_c_455_n N_VPWR_c_560_n 0.0436952f $X=5.68 $Y=1.985 $X2=0
+ $Y2=0
cc_386 N_A_31_368#_c_450_n N_VPWR_c_562_n 0.00749631f $X=2.08 $Y=2.4 $X2=0 $Y2=0
cc_387 N_A_31_368#_c_451_n N_VPWR_c_564_n 0.014552f $X=2.98 $Y=2.815 $X2=0 $Y2=0
cc_388 N_A_31_368#_c_452_n N_VPWR_c_566_n 0.0422287f $X=4.665 $Y=2.99 $X2=0
+ $Y2=0
cc_389 N_A_31_368#_c_453_n N_VPWR_c_566_n 0.0200196f $X=3.995 $Y=2.99 $X2=0
+ $Y2=0
cc_390 N_A_31_368#_c_454_n N_VPWR_c_566_n 0.062301f $X=5.565 $Y=2.99 $X2=0 $Y2=0
cc_391 N_A_31_368#_c_457_n N_VPWR_c_566_n 0.016488f $X=4.78 $Y=2.99 $X2=0 $Y2=0
cc_392 N_A_31_368#_c_448_n N_VPWR_c_570_n 0.011066f $X=0.28 $Y=2.815 $X2=0 $Y2=0
cc_393 N_A_31_368#_c_449_n N_VPWR_c_571_n 0.00749631f $X=1.18 $Y=2.815 $X2=0
+ $Y2=0
cc_394 N_A_31_368#_c_448_n N_VPWR_c_555_n 0.00915947f $X=0.28 $Y=2.815 $X2=0
+ $Y2=0
cc_395 N_A_31_368#_c_449_n N_VPWR_c_555_n 0.0062048f $X=1.18 $Y=2.815 $X2=0
+ $Y2=0
cc_396 N_A_31_368#_c_450_n N_VPWR_c_555_n 0.0062048f $X=2.08 $Y=2.4 $X2=0 $Y2=0
cc_397 N_A_31_368#_c_451_n N_VPWR_c_555_n 0.0119791f $X=2.98 $Y=2.815 $X2=0
+ $Y2=0
cc_398 N_A_31_368#_c_452_n N_VPWR_c_555_n 0.0238173f $X=4.665 $Y=2.99 $X2=0
+ $Y2=0
cc_399 N_A_31_368#_c_453_n N_VPWR_c_555_n 0.0108171f $X=3.995 $Y=2.99 $X2=0
+ $Y2=0
cc_400 N_A_31_368#_c_454_n N_VPWR_c_555_n 0.0347031f $X=5.565 $Y=2.99 $X2=0
+ $Y2=0
cc_401 N_A_31_368#_c_457_n N_VPWR_c_555_n 0.00894187f $X=4.78 $Y=2.99 $X2=0
+ $Y2=0
cc_402 N_A_31_368#_c_452_n N_Y_M1005_d 0.00197722f $X=4.665 $Y=2.99 $X2=0 $Y2=0
cc_403 N_A_31_368#_c_454_n N_Y_M1009_d 0.00197722f $X=5.565 $Y=2.99 $X2=0 $Y2=0
cc_404 N_A_31_368#_c_456_n N_Y_c_665_n 0.00626207f $X=2.08 $Y=1.985 $X2=0 $Y2=0
cc_405 N_A_31_368#_M1006_s N_Y_c_666_n 6.41842e-19 $X=4.63 $Y=1.84 $X2=0 $Y2=0
cc_406 N_A_31_368#_c_487_n N_Y_c_666_n 0.0017692f $X=3.855 $Y=2.12 $X2=0 $Y2=0
cc_407 N_A_31_368#_c_498_n N_Y_c_666_n 0.00522938f $X=4.78 $Y=2.325 $X2=0 $Y2=0
cc_408 N_A_31_368#_c_452_n N_Y_c_710_n 0.0160777f $X=4.665 $Y=2.99 $X2=0 $Y2=0
cc_409 N_A_31_368#_M1006_s N_Y_c_673_n 0.00135003f $X=4.63 $Y=1.84 $X2=0 $Y2=0
cc_410 N_A_31_368#_c_498_n N_Y_c_673_n 0.0103774f $X=4.78 $Y=2.325 $X2=0 $Y2=0
cc_411 N_A_31_368#_c_455_n N_Y_c_674_n 0.00793541f $X=5.68 $Y=1.985 $X2=0 $Y2=0
cc_412 N_A_31_368#_c_454_n N_Y_c_728_n 0.0160777f $X=5.565 $Y=2.99 $X2=0 $Y2=0
cc_413 N_Y_c_675_n N_A_46_74#_M1003_d 0.00436671f $X=1.48 $Y=0.855 $X2=0 $Y2=0
cc_414 N_Y_c_665_n N_A_46_74#_M1013_d 0.00176461f $X=3.965 $Y=1.175 $X2=0 $Y2=0
cc_415 N_Y_c_665_n N_A_46_74#_M1011_s 0.00176461f $X=3.965 $Y=1.175 $X2=0 $Y2=0
cc_416 N_Y_c_665_n N_A_46_74#_M1026_s 0.00230047f $X=3.965 $Y=1.175 $X2=0 $Y2=0
cc_417 N_Y_M1000_s N_A_46_74#_c_776_n 0.00178571f $X=0.645 $Y=0.37 $X2=0 $Y2=0
cc_418 N_Y_M1004_s N_A_46_74#_c_776_n 0.00178571f $X=1.505 $Y=0.37 $X2=0 $Y2=0
cc_419 N_Y_c_675_n N_A_46_74#_c_776_n 0.0288691f $X=1.48 $Y=0.855 $X2=0 $Y2=0
cc_420 N_Y_c_665_n N_A_46_74#_c_776_n 0.00367211f $X=3.965 $Y=1.175 $X2=0 $Y2=0
cc_421 N_Y_c_670_n N_A_46_74#_c_776_n 0.0144527f $X=0.825 $Y=0.855 $X2=0 $Y2=0
cc_422 N_Y_c_671_n N_A_46_74#_c_776_n 0.0165193f $X=1.645 $Y=0.855 $X2=0 $Y2=0
cc_423 N_Y_c_665_n N_A_46_74#_c_788_n 0.0323235f $X=3.965 $Y=1.175 $X2=0 $Y2=0
cc_424 N_Y_c_665_n N_A_46_74#_c_804_n 0.0133131f $X=3.965 $Y=1.175 $X2=0 $Y2=0
cc_425 N_Y_c_665_n N_A_46_74#_c_790_n 0.0323235f $X=3.965 $Y=1.175 $X2=0 $Y2=0
cc_426 N_Y_c_670_n N_A_46_74#_c_777_n 0.0136308f $X=0.825 $Y=0.855 $X2=0 $Y2=0
cc_427 N_Y_c_665_n N_A_46_74#_c_807_n 0.0129669f $X=3.965 $Y=1.175 $X2=0 $Y2=0
cc_428 N_Y_c_665_n N_A_46_74#_c_778_n 0.0194084f $X=3.965 $Y=1.175 $X2=0 $Y2=0
cc_429 N_Y_c_667_n N_A_46_74#_c_778_n 0.00109563f $X=4.775 $Y=0.515 $X2=0 $Y2=0
cc_430 N_Y_c_665_n N_VGND_M1010_d 0.00176891f $X=3.965 $Y=1.175 $X2=-0.19
+ $Y2=-0.245
cc_431 N_Y_c_665_n N_VGND_M1019_d 0.00176891f $X=3.965 $Y=1.175 $X2=0 $Y2=0
cc_432 N_Y_c_666_n N_VGND_M1012_s 0.00261869f $X=4.33 $Y=1.99 $X2=0 $Y2=0
cc_433 N_Y_c_668_n N_VGND_M1018_s 0.00176461f $X=5.47 $Y=1.065 $X2=0 $Y2=0
cc_434 N_Y_c_666_n N_VGND_c_832_n 0.0191564f $X=4.33 $Y=1.99 $X2=0 $Y2=0
cc_435 N_Y_c_667_n N_VGND_c_832_n 0.0189326f $X=4.775 $Y=0.515 $X2=0 $Y2=0
cc_436 N_Y_c_667_n N_VGND_c_833_n 0.0109942f $X=4.775 $Y=0.515 $X2=0 $Y2=0
cc_437 N_Y_c_667_n N_VGND_c_834_n 0.0165282f $X=4.775 $Y=0.515 $X2=0 $Y2=0
cc_438 N_Y_c_668_n N_VGND_c_834_n 0.0152916f $X=5.47 $Y=1.065 $X2=0 $Y2=0
cc_439 N_Y_c_669_n N_VGND_c_834_n 0.0165282f $X=5.635 $Y=0.515 $X2=0 $Y2=0
cc_440 N_Y_c_669_n N_VGND_c_835_n 0.023308f $X=5.635 $Y=0.515 $X2=0 $Y2=0
cc_441 N_Y_c_669_n N_VGND_c_842_n 0.0109942f $X=5.635 $Y=0.515 $X2=0 $Y2=0
cc_442 N_Y_c_667_n N_VGND_c_844_n 0.00904371f $X=4.775 $Y=0.515 $X2=0 $Y2=0
cc_443 N_Y_c_669_n N_VGND_c_844_n 0.00904371f $X=5.635 $Y=0.515 $X2=0 $Y2=0
cc_444 N_A_46_74#_c_788_n N_VGND_M1010_d 0.0033542f $X=2.85 $Y=0.835 $X2=-0.19
+ $Y2=-0.245
cc_445 N_A_46_74#_c_790_n N_VGND_M1019_d 0.0033542f $X=3.71 $Y=0.835 $X2=0 $Y2=0
cc_446 N_A_46_74#_c_776_n N_VGND_c_830_n 0.00913089f $X=1.99 $Y=0.475 $X2=0
+ $Y2=0
cc_447 N_A_46_74#_c_788_n N_VGND_c_830_n 0.0165203f $X=2.85 $Y=0.835 $X2=0 $Y2=0
cc_448 N_A_46_74#_c_790_n N_VGND_c_831_n 0.0165203f $X=3.71 $Y=0.835 $X2=0 $Y2=0
cc_449 N_A_46_74#_c_778_n N_VGND_c_832_n 0.0246655f $X=3.795 $Y=0.725 $X2=0
+ $Y2=0
cc_450 N_A_46_74#_c_776_n N_VGND_c_836_n 0.0668236f $X=1.99 $Y=0.475 $X2=0 $Y2=0
cc_451 N_A_46_74#_c_788_n N_VGND_c_836_n 0.00197156f $X=2.85 $Y=0.835 $X2=0
+ $Y2=0
cc_452 N_A_46_74#_c_777_n N_VGND_c_836_n 0.0146502f $X=0.355 $Y=0.515 $X2=0
+ $Y2=0
cc_453 N_A_46_74#_c_788_n N_VGND_c_838_n 0.00197156f $X=2.85 $Y=0.835 $X2=0
+ $Y2=0
cc_454 N_A_46_74#_c_790_n N_VGND_c_838_n 0.00197156f $X=3.71 $Y=0.835 $X2=0
+ $Y2=0
cc_455 N_A_46_74#_c_807_n N_VGND_c_838_n 0.00418578f $X=2.935 $Y=0.725 $X2=0
+ $Y2=0
cc_456 N_A_46_74#_c_790_n N_VGND_c_840_n 0.00197156f $X=3.71 $Y=0.835 $X2=0
+ $Y2=0
cc_457 N_A_46_74#_c_778_n N_VGND_c_840_n 0.00623759f $X=3.795 $Y=0.725 $X2=0
+ $Y2=0
cc_458 N_A_46_74#_c_776_n N_VGND_c_844_n 0.0560338f $X=1.99 $Y=0.475 $X2=0 $Y2=0
cc_459 N_A_46_74#_c_788_n N_VGND_c_844_n 0.00938768f $X=2.85 $Y=0.835 $X2=0
+ $Y2=0
cc_460 N_A_46_74#_c_790_n N_VGND_c_844_n 0.00939316f $X=3.71 $Y=0.835 $X2=0
+ $Y2=0
cc_461 N_A_46_74#_c_777_n N_VGND_c_844_n 0.0120674f $X=0.355 $Y=0.515 $X2=0
+ $Y2=0
cc_462 N_A_46_74#_c_807_n N_VGND_c_844_n 0.00545294f $X=2.935 $Y=0.725 $X2=0
+ $Y2=0
cc_463 N_A_46_74#_c_778_n N_VGND_c_844_n 0.0080625f $X=3.795 $Y=0.725 $X2=0
+ $Y2=0
