* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__nor2b_2 A B_N VGND VNB VPB VPWR Y
M1000 VPWR A a_228_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=6.31e+11p pd=5.43e+06u as=9.912e+11p ps=8.49e+06u
M1001 Y a_27_392# VGND VNB nshort w=740000u l=150000u
+  ad=4.884e+11p pd=4.28e+06u as=7.744e+11p ps=6.56e+06u
M1002 VGND B_N a_27_392# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1003 a_228_368# A VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND a_27_392# Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y A VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y a_27_392# a_228_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=0p ps=0u
M1007 VGND A Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR B_N a_27_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1009 a_228_368# a_27_392# Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
