* File: sky130_fd_sc_ls__dfbbp_1.pex.spice
* Created: Fri Aug 28 13:13:41 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__DFBBP_1%CLK 1 3 4 6 7
r32 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.52
+ $Y=1.385 $X2=0.52 $Y2=1.385
r33 7 11 6.22942 $w=3.68e-07 $l=2e-07 $layer=LI1_cond $X=0.72 $Y=1.365 $X2=0.52
+ $Y2=1.365
r34 4 10 77.2841 $w=2.7e-07 $l=4.15812e-07 $layer=POLY_cond $X=0.595 $Y=1.765
+ $X2=0.52 $Y2=1.385
r35 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.595 $Y=1.765
+ $X2=0.595 $Y2=2.4
r36 1 10 38.9026 $w=2.7e-07 $l=1.77059e-07 $layer=POLY_cond $X=0.495 $Y=1.22
+ $X2=0.52 $Y2=1.385
r37 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.495 $Y=1.22 $X2=0.495
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__DFBBP_1%D 3 5 7 8 12
r38 12 14 72.1174 $w=2.64e-07 $l=3.95e-07 $layer=POLY_cond $X=2.125 $Y=2.032
+ $X2=2.52 $Y2=2.032
r39 10 12 16.4318 $w=2.64e-07 $l=9e-08 $layer=POLY_cond $X=2.035 $Y=2.032
+ $X2=2.125 $Y2=2.032
r40 8 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.125
+ $Y=1.99 $X2=2.125 $Y2=1.99
r41 5 14 15.9823 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.52 $Y=2.24
+ $X2=2.52 $Y2=2.032
r42 5 7 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.52 $Y=2.24 $X2=2.52
+ $Y2=2.525
r43 1 10 15.9823 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.035 $Y=1.825
+ $X2=2.035 $Y2=2.032
r44 1 3 507.638 $w=1.5e-07 $l=9.9e-07 $layer=POLY_cond $X=2.035 $Y=1.825
+ $X2=2.035 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_LS__DFBBP_1%A_671_93# 1 2 7 9 11 12 14 16 17 19 20 22 24
+ 27 28 30 31 34 36 37 38 39 43 47 49 54
c164 43 0 6.96239e-20 $X=5.935 $Y=1.825
c165 39 0 9.97901e-20 $X=5.335 $Y=0.925
c166 31 0 5.24889e-20 $X=3.72 $Y=0.815
c167 27 0 9.83523e-20 $X=3.59 $Y=1.29
c168 17 0 1.41852e-19 $X=5.94 $Y=1.82
c169 7 0 1.68855e-19 $X=3.43 $Y=1.125
r170 48 57 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.015 $Y=1.42
+ $X2=6.015 $Y2=1.585
r171 48 54 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=6.015 $Y=1.42
+ $X2=6.015 $Y2=1.295
r172 47 50 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=6.015 $Y=1.42
+ $X2=6.015 $Y2=1.585
r173 47 49 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=6.015 $Y=1.42
+ $X2=6.015 $Y2=1.255
r174 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.015
+ $Y=1.42 $X2=6.015 $Y2=1.42
r175 43 50 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=5.935 $Y=1.825
+ $X2=5.935 $Y2=1.585
r176 40 49 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=5.935 $Y=1.01
+ $X2=5.935 $Y2=1.255
r177 39 45 9.11221 $w=3.9e-07 $l=2.17991e-07 $layer=LI1_cond $X=5.335 $Y=0.925
+ $X2=5.17 $Y2=0.802
r178 38 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.85 $Y=0.925
+ $X2=5.935 $Y2=1.01
r179 38 39 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=5.85 $Y=0.925
+ $X2=5.335 $Y2=0.925
r180 36 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.85 $Y=1.91
+ $X2=5.935 $Y2=1.825
r181 36 37 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=5.85 $Y=1.91 $X2=4.95
+ $Y2=1.91
r182 32 37 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.825 $Y=1.995
+ $X2=4.95 $Y2=1.91
r183 32 34 2.0744 $w=2.48e-07 $l=4.5e-08 $layer=LI1_cond $X=4.825 $Y=1.995
+ $X2=4.825 $Y2=2.04
r184 30 45 8.79939 $w=3.9e-07 $l=1.61369e-07 $layer=LI1_cond $X=5.015 $Y=0.815
+ $X2=5.17 $Y2=0.802
r185 30 31 84.4866 $w=1.68e-07 $l=1.295e-06 $layer=LI1_cond $X=5.015 $Y=0.815
+ $X2=3.72 $Y2=0.815
r186 28 51 28.8839 $w=2.67e-07 $l=1.6e-07 $layer=POLY_cond $X=3.59 $Y=1.29
+ $X2=3.43 $Y2=1.29
r187 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.59
+ $Y=1.29 $X2=3.59 $Y2=1.29
r188 25 31 7.17723 $w=1.7e-07 $l=1.65118e-07 $layer=LI1_cond $X=3.592 $Y=0.9
+ $X2=3.72 $Y2=0.815
r189 25 27 17.6256 $w=2.53e-07 $l=3.9e-07 $layer=LI1_cond $X=3.592 $Y=0.9
+ $X2=3.592 $Y2=1.29
r190 22 24 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=6.515 $Y=1.22
+ $X2=6.515 $Y2=0.87
r191 21 54 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.18 $Y=1.295
+ $X2=6.015 $Y2=1.295
r192 20 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.44 $Y=1.295
+ $X2=6.515 $Y2=1.22
r193 20 21 133.319 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=6.44 $Y=1.295
+ $X2=6.18 $Y2=1.295
r194 17 19 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=5.94 $Y=1.82
+ $X2=5.94 $Y2=2.315
r195 16 17 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.94 $Y=1.73 $X2=5.94
+ $Y2=1.82
r196 16 57 56.3629 $w=1.8e-07 $l=1.45e-07 $layer=POLY_cond $X=5.94 $Y=1.73
+ $X2=5.94 $Y2=1.585
r197 12 14 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.88 $Y=1.82
+ $X2=3.88 $Y2=2.105
r198 11 12 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.88 $Y=1.73 $X2=3.88
+ $Y2=1.82
r199 10 28 52.3521 $w=2.67e-07 $l=3.63249e-07 $layer=POLY_cond $X=3.88 $Y=1.455
+ $X2=3.59 $Y2=1.29
r200 10 11 106.895 $w=1.8e-07 $l=2.75e-07 $layer=POLY_cond $X=3.88 $Y=1.455
+ $X2=3.88 $Y2=1.73
r201 7 51 16.2448 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.43 $Y=1.125
+ $X2=3.43 $Y2=1.29
r202 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.43 $Y=1.125
+ $X2=3.43 $Y2=0.805
r203 2 34 300 $w=1.7e-07 $l=3.03974e-07 $layer=licon1_PDIFF $count=2 $X=4.545
+ $Y=1.895 $X2=4.785 $Y2=2.04
r204 1 45 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=5.03
+ $Y=0.595 $X2=5.17 $Y2=0.8
.ends

.subckt PM_SKY130_FD_SC_LS__DFBBP_1%SET_B 3 5 7 10 12 14 16 17 18 20 21 22 24 25
+ 26 28 29 30 35 37
c164 12 0 1.01328e-19 $X=8.48 $Y=1.885
r165 37 45 7.33544 $w=3.16e-07 $l=1.9e-07 $layer=LI1_cond $X=8.405 $Y=1.635
+ $X2=8.405 $Y2=1.825
r166 37 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.405
+ $Y=1.635 $X2=8.405 $Y2=1.635
r167 32 35 2.35192 $w=2.43e-07 $l=5e-08 $layer=LI1_cond $X=4.395 $Y=1.532
+ $X2=4.445 $Y2=1.532
r168 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.395
+ $Y=1.53 $X2=4.395 $Y2=1.53
r169 29 45 4.36715 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.24 $Y=1.825
+ $X2=8.405 $Y2=1.825
r170 29 30 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=8.24 $Y=1.825
+ $X2=7.45 $Y2=1.825
r171 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.365 $Y=1.91
+ $X2=7.45 $Y2=1.825
r172 27 28 64.9144 $w=1.68e-07 $l=9.95e-07 $layer=LI1_cond $X=7.365 $Y=1.91
+ $X2=7.365 $Y2=2.905
r173 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.28 $Y=2.99
+ $X2=7.365 $Y2=2.905
r174 25 26 69.8075 $w=1.68e-07 $l=1.07e-06 $layer=LI1_cond $X=7.28 $Y=2.99
+ $X2=6.21 $Y2=2.99
r175 24 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.125 $Y=2.905
+ $X2=6.21 $Y2=2.99
r176 23 24 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=6.125 $Y=2.335
+ $X2=6.125 $Y2=2.905
r177 21 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.04 $Y=2.25
+ $X2=6.125 $Y2=2.335
r178 21 22 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=6.04 $Y=2.25
+ $X2=5.33 $Y2=2.25
r179 19 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.245 $Y=2.335
+ $X2=5.33 $Y2=2.25
r180 19 20 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=5.245 $Y=2.335
+ $X2=5.245 $Y2=2.905
r181 17 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.16 $Y=2.99
+ $X2=5.245 $Y2=2.905
r182 17 18 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=5.16 $Y=2.99
+ $X2=4.53 $Y2=2.99
r183 16 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.445 $Y=2.905
+ $X2=4.53 $Y2=2.99
r184 15 35 2.87745 $w=1.7e-07 $l=1.23e-07 $layer=LI1_cond $X=4.445 $Y=1.655
+ $X2=4.445 $Y2=1.532
r185 15 16 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=4.445 $Y=1.655
+ $X2=4.445 $Y2=2.905
r186 12 41 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=8.48 $Y=1.885
+ $X2=8.405 $Y2=1.635
r187 12 14 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=8.48 $Y=1.885
+ $X2=8.48 $Y2=2.46
r188 8 41 38.5562 $w=2.99e-07 $l=1.92678e-07 $layer=POLY_cond $X=8.465 $Y=1.47
+ $X2=8.405 $Y2=1.635
r189 8 10 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=8.465 $Y=1.47
+ $X2=8.465 $Y2=0.74
r190 5 33 58.4261 $w=3.03e-07 $l=3.29773e-07 $layer=POLY_cond $X=4.47 $Y=1.82
+ $X2=4.385 $Y2=1.53
r191 5 7 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=4.47 $Y=1.82 $X2=4.47
+ $Y2=2.315
r192 1 33 38.5416 $w=3.03e-07 $l=2.09105e-07 $layer=POLY_cond $X=4.285 $Y=1.365
+ $X2=4.385 $Y2=1.53
r193 1 3 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=4.285 $Y=1.365
+ $X2=4.285 $Y2=0.87
.ends

.subckt PM_SKY130_FD_SC_LS__DFBBP_1%A_520_87# 1 2 9 11 12 14 15 20 23 25 28 29
+ 30 31 35 37
c109 35 0 9.97901e-20 $X=4.935 $Y=1.42
c110 30 0 1.68855e-19 $X=4.06 $Y=1.155
r111 35 38 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.935 $Y=1.42
+ $X2=4.935 $Y2=1.585
r112 35 37 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.935 $Y=1.42
+ $X2=4.935 $Y2=1.255
r113 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.935
+ $Y=1.42 $X2=4.935 $Y2=1.42
r114 29 34 11.2257 $w=2.88e-07 $l=3.42243e-07 $layer=LI1_cond $X=4.745 $Y=1.155
+ $X2=4.922 $Y2=1.42
r115 29 30 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=4.745 $Y=1.155
+ $X2=4.06 $Y2=1.155
r116 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.975 $Y=1.24
+ $X2=4.06 $Y2=1.155
r117 27 28 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=3.975 $Y=1.24
+ $X2=3.975 $Y2=1.625
r118 26 31 2.57001 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=3.43 $Y=1.71
+ $X2=3.277 $Y2=1.71
r119 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.89 $Y=1.71
+ $X2=3.975 $Y2=1.625
r120 25 26 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=3.89 $Y=1.71
+ $X2=3.43 $Y2=1.71
r121 21 31 3.87901 $w=2.37e-07 $l=8.5e-08 $layer=LI1_cond $X=3.277 $Y=1.795
+ $X2=3.277 $Y2=1.71
r122 21 23 14.1694 $w=3.03e-07 $l=3.75e-07 $layer=LI1_cond $X=3.277 $Y=1.795
+ $X2=3.277 $Y2=2.17
r123 20 31 3.87901 $w=2.37e-07 $l=1.13666e-07 $layer=LI1_cond $X=3.21 $Y=1.625
+ $X2=3.277 $Y2=1.71
r124 19 20 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=3.21 $Y=0.745
+ $X2=3.21 $Y2=1.625
r125 15 19 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.125 $Y=0.58
+ $X2=3.21 $Y2=0.745
r126 15 17 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=3.125 $Y=0.58
+ $X2=2.74 $Y2=0.58
r127 12 14 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=5.01 $Y=1.82
+ $X2=5.01 $Y2=2.315
r128 11 12 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.01 $Y=1.73 $X2=5.01
+ $Y2=1.82
r129 11 38 56.3629 $w=1.8e-07 $l=1.45e-07 $layer=POLY_cond $X=5.01 $Y=1.73
+ $X2=5.01 $Y2=1.585
r130 9 37 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=4.955 $Y=0.87
+ $X2=4.955 $Y2=1.255
r131 2 23 600 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_PDIFF $count=1 $X=3.045
+ $Y=2.315 $X2=3.265 $Y2=2.17
r132 1 17 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.6
+ $Y=0.435 $X2=2.74 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_LS__DFBBP_1%A_1062_93# 1 2 9 11 12 14 16 17 19 20 22 23
+ 25 29 33 35 40 42 43 46 49 50 53 55 57 65
c151 57 0 9.47353e-20 $X=9.875 $Y=1.295
c152 12 0 6.96239e-20 $X=5.43 $Y=1.82
r153 53 56 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.475 $Y=1.42
+ $X2=5.475 $Y2=1.585
r154 53 55 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.475 $Y=1.42
+ $X2=5.475 $Y2=1.255
r155 50 65 6.55126 $w=3.53e-07 $l=1.05e-07 $layer=LI1_cond $X=9.887 $Y=1.295
+ $X2=9.887 $Y2=1.19
r156 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=1.295
+ $X2=9.84 $Y2=1.295
r157 46 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.475
+ $Y=1.42 $X2=5.475 $Y2=1.42
r158 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=1.295
+ $X2=5.52 $Y2=1.295
r159 43 45 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.665 $Y=1.295
+ $X2=5.52 $Y2=1.295
r160 42 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.695 $Y=1.295
+ $X2=9.84 $Y2=1.295
r161 42 43 4.98761 $w=1.4e-07 $l=4.03e-06 $layer=MET1_cond $X=9.695 $Y=1.295
+ $X2=5.665 $Y2=1.295
r162 37 40 6.24041 $w=4.58e-07 $l=2.4e-07 $layer=LI1_cond $X=9.98 $Y=0.58
+ $X2=10.22 $Y2=0.58
r163 33 35 8.0671 $w=2.48e-07 $l=1.75e-07 $layer=LI1_cond $X=10.065 $Y=1.945
+ $X2=10.24 $Y2=1.945
r164 31 37 6.6364 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=9.98 $Y=0.81 $X2=9.98
+ $Y2=0.58
r165 31 65 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=9.98 $Y=0.81
+ $X2=9.98 $Y2=1.19
r166 30 57 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=9.875 $Y=1.385
+ $X2=9.875 $Y2=1.295
r167 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.875
+ $Y=1.385 $X2=9.875 $Y2=1.385
r168 27 33 7.08698 $w=2.5e-07 $l=2.32237e-07 $layer=LI1_cond $X=9.887 $Y=1.82
+ $X2=10.065 $Y2=1.945
r169 27 29 14.1215 $w=3.53e-07 $l=4.35e-07 $layer=LI1_cond $X=9.887 $Y=1.82
+ $X2=9.887 $Y2=1.385
r170 26 50 2.33735 $w=3.53e-07 $l=7.2e-08 $layer=LI1_cond $X=9.887 $Y=1.367
+ $X2=9.887 $Y2=1.295
r171 26 29 0.584337 $w=3.53e-07 $l=1.8e-08 $layer=LI1_cond $X=9.887 $Y=1.367
+ $X2=9.887 $Y2=1.385
r172 24 25 6.66866 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=9.5 $Y=1.295 $X2=9.41
+ $Y2=1.295
r173 23 57 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.71 $Y=1.295
+ $X2=9.875 $Y2=1.295
r174 23 24 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=9.71 $Y=1.295
+ $X2=9.5 $Y2=1.295
r175 20 22 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=9.41 $Y=1.885
+ $X2=9.41 $Y2=2.46
r176 17 25 18.8402 $w=1.65e-07 $l=7.98436e-08 $layer=POLY_cond $X=9.4 $Y=1.22
+ $X2=9.41 $Y2=1.295
r177 17 19 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=9.4 $Y=1.22 $X2=9.4
+ $Y2=0.74
r178 16 20 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=9.41 $Y=1.795
+ $X2=9.41 $Y2=1.885
r179 15 25 18.8402 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=9.41 $Y=1.37
+ $X2=9.41 $Y2=1.295
r180 15 16 165.202 $w=1.8e-07 $l=4.25e-07 $layer=POLY_cond $X=9.41 $Y=1.37
+ $X2=9.41 $Y2=1.795
r181 12 14 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=5.43 $Y=1.82
+ $X2=5.43 $Y2=2.315
r182 11 12 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.43 $Y=1.73 $X2=5.43
+ $Y2=1.82
r183 11 56 56.3629 $w=1.8e-07 $l=1.45e-07 $layer=POLY_cond $X=5.43 $Y=1.73
+ $X2=5.43 $Y2=1.585
r184 9 55 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=5.385 $Y=0.87
+ $X2=5.385 $Y2=1.255
r185 2 35 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=10.115
+ $Y=1.84 $X2=10.24 $Y2=1.985
r186 1 40 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=10.075
+ $Y=0.37 $X2=10.22 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_LS__DFBBP_1%A_27_74# 1 2 9 11 13 14 17 18 19 21 22 23 26
+ 28 29 30 32 33 35 38 41 43 45 48 51 54 58 62 67 68 71 72 74 75 77 79 85
c224 77 0 1.41852e-19 $X=6.605 $Y=1.775
c225 71 0 1.41865e-20 $X=7.505 $Y=1.065
c226 30 0 9.83523e-20 $X=3.49 $Y=2.39
c227 26 0 1.57784e-19 $X=2.525 $Y=0.645
c228 17 0 9.68576e-20 $X=1.525 $Y=1.3
c229 11 0 7.24936e-20 $X=1.175 $Y=1.765
c230 9 0 6.93165e-20 $X=0.995 $Y=0.74
r231 77 79 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=6.605 $Y=1.775
+ $X2=6.605 $Y2=1.61
r232 77 78 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.605
+ $Y=1.775 $X2=6.605 $Y2=1.775
r233 72 85 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.505 $Y=1.065
+ $X2=7.505 $Y2=0.9
r234 71 72 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.505
+ $Y=1.065 $X2=7.505 $Y2=1.065
r235 69 71 22.6943 $w=3.23e-07 $l=6.4e-07 $layer=LI1_cond $X=7.507 $Y=0.425
+ $X2=7.507 $Y2=1.065
r236 67 69 7.72402 $w=1.7e-07 $l=2.00035e-07 $layer=LI1_cond $X=7.345 $Y=0.34
+ $X2=7.507 $Y2=0.425
r237 67 68 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=7.345 $Y=0.34
+ $X2=6.77 $Y2=0.34
r238 65 68 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.685 $Y=0.425
+ $X2=6.77 $Y2=0.34
r239 65 79 77.3102 $w=1.68e-07 $l=1.185e-06 $layer=LI1_cond $X=6.685 $Y=0.425
+ $X2=6.685 $Y2=1.61
r240 63 81 13.8153 $w=3.14e-07 $l=9e-08 $layer=POLY_cond $X=1.08 $Y=1.465
+ $X2=1.08 $Y2=1.375
r241 62 63 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.06
+ $Y=1.465 $X2=1.06 $Y2=1.465
r242 60 62 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.06 $Y=1.72
+ $X2=1.06 $Y2=1.465
r243 59 75 3.57226 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=0.535 $Y=1.805
+ $X2=0.31 $Y2=1.805
r244 58 60 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.975 $Y=1.805
+ $X2=1.06 $Y2=1.72
r245 58 59 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=0.975 $Y=1.805
+ $X2=0.535 $Y2=1.805
r246 54 56 22.061 $w=4.48e-07 $l=8.3e-07 $layer=LI1_cond $X=0.31 $Y=1.985
+ $X2=0.31 $Y2=2.815
r247 52 75 3.05675 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.31 $Y=1.89
+ $X2=0.31 $Y2=1.805
r248 52 54 2.52505 $w=4.48e-07 $l=9.5e-08 $layer=LI1_cond $X=0.31 $Y=1.89
+ $X2=0.31 $Y2=1.985
r249 51 75 3.05675 $w=3.1e-07 $l=1.77482e-07 $layer=LI1_cond $X=0.17 $Y=1.72
+ $X2=0.31 $Y2=1.805
r250 51 74 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=0.17 $Y=1.72
+ $X2=0.17 $Y2=1.01
r251 46 74 8.99121 $w=3.58e-07 $l=1.8e-07 $layer=LI1_cond $X=0.265 $Y=0.83
+ $X2=0.265 $Y2=1.01
r252 46 48 10.0839 $w=3.58e-07 $l=3.15e-07 $layer=LI1_cond $X=0.265 $Y=0.83
+ $X2=0.265 $Y2=0.515
r253 42 43 76.9149 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=1.525 $Y=1.375
+ $X2=1.675 $Y2=1.375
r254 41 85 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=7.415 $Y=0.58
+ $X2=7.415 $Y2=0.9
r255 36 38 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=6.48 $Y=3.035
+ $X2=6.48 $Y2=2.54
r256 35 78 53.8969 $w=3.31e-07 $l=3.1607e-07 $layer=POLY_cond $X=6.48 $Y=2.045
+ $X2=6.58 $Y2=1.775
r257 35 38 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=6.48 $Y=2.045
+ $X2=6.48 $Y2=2.54
r258 34 45 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.58 $Y=3.15 $X2=3.49
+ $Y2=3.15
r259 33 36 26.9307 $w=1.5e-07 $l=1.53542e-07 $layer=POLY_cond $X=6.39 $Y=3.15
+ $X2=6.48 $Y2=3.035
r260 33 34 1440.87 $w=1.5e-07 $l=2.81e-06 $layer=POLY_cond $X=6.39 $Y=3.15
+ $X2=3.58 $Y2=3.15
r261 30 32 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.49 $Y=2.39
+ $X2=3.49 $Y2=2.105
r262 29 45 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=3.49 $Y=3.075
+ $X2=3.49 $Y2=3.15
r263 28 30 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.49 $Y=2.48 $X2=3.49
+ $Y2=2.39
r264 28 29 231.282 $w=1.8e-07 $l=5.95e-07 $layer=POLY_cond $X=3.49 $Y=2.48
+ $X2=3.49 $Y2=3.075
r265 24 26 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=2.525 $Y=0.255
+ $X2=2.525 $Y2=0.645
r266 22 45 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.4 $Y=3.15 $X2=3.49
+ $Y2=3.15
r267 22 23 846.064 $w=1.5e-07 $l=1.65e-06 $layer=POLY_cond $X=3.4 $Y=3.15
+ $X2=1.75 $Y2=3.15
r268 21 23 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.675 $Y=3.075
+ $X2=1.75 $Y2=3.15
r269 20 43 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.675 $Y=1.45
+ $X2=1.675 $Y2=1.375
r270 20 21 833.245 $w=1.5e-07 $l=1.625e-06 $layer=POLY_cond $X=1.675 $Y=1.45
+ $X2=1.675 $Y2=3.075
r271 18 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.45 $Y=0.18
+ $X2=2.525 $Y2=0.255
r272 18 19 435.851 $w=1.5e-07 $l=8.5e-07 $layer=POLY_cond $X=2.45 $Y=0.18
+ $X2=1.6 $Y2=0.18
r273 17 42 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.525 $Y=1.3
+ $X2=1.525 $Y2=1.375
r274 16 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.525 $Y=0.255
+ $X2=1.6 $Y2=0.18
r275 16 17 535.84 $w=1.5e-07 $l=1.045e-06 $layer=POLY_cond $X=1.525 $Y=0.255
+ $X2=1.525 $Y2=1.3
r276 15 81 20.044 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=1.265 $Y=1.375
+ $X2=1.08 $Y2=1.375
r277 14 42 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.45 $Y=1.375
+ $X2=1.525 $Y2=1.375
r278 14 15 94.8617 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=1.45 $Y=1.375
+ $X2=1.265 $Y2=1.375
r279 11 63 59.2576 $w=3.14e-07 $l=3.44238e-07 $layer=POLY_cond $X=1.175 $Y=1.765
+ $X2=1.08 $Y2=1.465
r280 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.175 $Y=1.765
+ $X2=1.175 $Y2=2.4
r281 7 81 24.7194 $w=3.14e-07 $l=1.16619e-07 $layer=POLY_cond $X=0.995 $Y=1.3
+ $X2=1.08 $Y2=1.375
r282 7 9 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.995 $Y=1.3
+ $X2=0.995 $Y2=0.74
r283 2 56 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.225
+ $Y=1.84 $X2=0.37 $Y2=2.815
r284 2 54 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.225
+ $Y=1.84 $X2=0.37 $Y2=1.985
r285 1 48 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__DFBBP_1%A_214_74# 1 2 7 12 14 15 17 18 19 23 24 26
+ 28 29 32 36 38 40 46 50
c140 46 0 1.57784e-19 $X=2.485 $Y=1.42
c141 32 0 1.41865e-20 $X=7.055 $Y=1.295
c142 12 0 5.24889e-20 $X=2.955 $Y=0.645
r143 47 50 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.485 $Y=1.42
+ $X2=2.485 $Y2=1.33
r144 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.485
+ $Y=1.42 $X2=2.485 $Y2=1.42
r145 44 46 32.1287 $w=3.28e-07 $l=9.2e-07 $layer=LI1_cond $X=1.565 $Y=1.42
+ $X2=2.485 $Y2=1.42
r146 40 42 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=1.44 $Y=1.985
+ $X2=1.44 $Y2=2.815
r147 38 44 7.64946 $w=2.65e-07 $l=2.07123e-07 $layer=LI1_cond $X=1.44 $Y=1.585
+ $X2=1.345 $Y2=1.42
r148 38 40 18.4391 $w=2.48e-07 $l=4e-07 $layer=LI1_cond $X=1.44 $Y=1.585
+ $X2=1.44 $Y2=1.985
r149 34 44 16.8014 $w=3.6e-07 $l=4.89592e-07 $layer=LI1_cond $X=1.305 $Y=0.95
+ $X2=1.345 $Y2=1.42
r150 34 36 13.9254 $w=3.58e-07 $l=4.35e-07 $layer=LI1_cond $X=1.305 $Y=0.95
+ $X2=1.305 $Y2=0.515
r151 30 32 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=6.875 $Y=1.295
+ $X2=7.055 $Y2=1.295
r152 27 32 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.055 $Y=1.37
+ $X2=7.055 $Y2=1.295
r153 27 28 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=7.055 $Y=1.37
+ $X2=7.055 $Y2=2.18
r154 24 28 71.1762 $w=1.93e-07 $l=3.04344e-07 $layer=POLY_cond $X=7.015 $Y=2.465
+ $X2=7.055 $Y2=2.18
r155 24 26 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.015 $Y=2.465
+ $X2=7.015 $Y2=2.75
r156 21 30 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.875 $Y=1.22
+ $X2=6.875 $Y2=1.295
r157 21 23 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=6.875 $Y=1.22
+ $X2=6.875 $Y2=0.87
r158 20 23 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=6.875 $Y=0.255
+ $X2=6.875 $Y2=0.87
r159 18 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.8 $Y=0.18
+ $X2=6.875 $Y2=0.255
r160 18 19 1933.13 $w=1.5e-07 $l=3.77e-06 $layer=POLY_cond $X=6.8 $Y=0.18
+ $X2=3.03 $Y2=0.18
r161 15 17 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.97 $Y=2.24
+ $X2=2.97 $Y2=2.525
r162 14 15 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.97 $Y=2.15 $X2=2.97
+ $Y2=2.24
r163 13 29 18.8402 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=2.97 $Y=1.405
+ $X2=2.97 $Y2=1.33
r164 13 14 289.589 $w=1.8e-07 $l=7.45e-07 $layer=POLY_cond $X=2.97 $Y=1.405
+ $X2=2.97 $Y2=2.15
r165 10 29 18.8402 $w=1.65e-07 $l=8.21584e-08 $layer=POLY_cond $X=2.955 $Y=1.255
+ $X2=2.97 $Y2=1.33
r166 10 12 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.955 $Y=1.255
+ $X2=2.955 $Y2=0.645
r167 9 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.955 $Y=0.255
+ $X2=3.03 $Y2=0.18
r168 9 12 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=2.955 $Y=0.255
+ $X2=2.955 $Y2=0.645
r169 8 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.65 $Y=1.33
+ $X2=2.485 $Y2=1.33
r170 7 29 6.66866 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.88 $Y=1.33 $X2=2.97
+ $Y2=1.33
r171 7 8 117.936 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=2.88 $Y=1.33 $X2=2.65
+ $Y2=1.33
r172 2 42 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.25
+ $Y=1.84 $X2=1.4 $Y2=2.815
r173 2 40 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.25
+ $Y=1.84 $X2=1.4 $Y2=1.985
r174 1 36 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.07
+ $Y=0.37 $X2=1.21 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__DFBBP_1%A_1474_446# 1 2 7 9 11 14 16 18 21 23 24 26
+ 28 29 31 32 34 37 41 43 46 51 55 58 59 62 65 68 72 77
c187 62 0 1.25678e-19 $X=10.865 $Y=2.24
c188 51 0 4.99671e-20 $X=7.785 $Y=2.215
c189 37 0 1.35822e-19 $X=7.955 $Y=1.81
c190 16 0 2.32792e-19 $X=10.98 $Y=1.765
c191 11 0 2.35385e-20 $X=7.875 $Y=2.05
r192 84 85 4.22807 $w=3.99e-07 $l=3.5e-08 $layer=POLY_cond $X=10.98 $Y=1.542
+ $X2=11.015 $Y2=1.542
r193 78 84 3.02005 $w=3.99e-07 $l=2.5e-08 $layer=POLY_cond $X=10.955 $Y=1.542
+ $X2=10.98 $Y2=1.542
r194 77 78 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.955
+ $Y=1.485 $X2=10.955 $Y2=1.485
r195 74 77 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=10.865 $Y=1.485
+ $X2=10.955 $Y2=1.485
r196 70 72 3.63098 $w=3.63e-07 $l=1.15e-07 $layer=LI1_cond $X=9.185 $Y=0.777
+ $X2=9.3 $Y2=0.777
r197 67 68 6.73996 $w=4.38e-07 $l=8.5e-08 $layer=LI1_cond $X=9.3 $Y=2.19
+ $X2=9.385 $Y2=2.19
r198 66 67 12.834 $w=4.38e-07 $l=4.9e-07 $layer=LI1_cond $X=8.81 $Y=2.19 $X2=9.3
+ $Y2=2.19
r199 64 66 1.04768 $w=4.38e-07 $l=4e-08 $layer=LI1_cond $X=8.77 $Y=2.19 $X2=8.81
+ $Y2=2.19
r200 64 65 3.40064 $w=4.38e-07 $l=8.5e-08 $layer=LI1_cond $X=8.77 $Y=2.19
+ $X2=8.685 $Y2=2.19
r201 61 74 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.865 $Y=1.65
+ $X2=10.865 $Y2=1.485
r202 61 62 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=10.865 $Y=1.65
+ $X2=10.865 $Y2=2.24
r203 59 62 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.78 $Y=2.325
+ $X2=10.865 $Y2=2.24
r204 59 68 91.0107 $w=1.68e-07 $l=1.395e-06 $layer=LI1_cond $X=10.78 $Y=2.325
+ $X2=9.385 $Y2=2.325
r205 58 67 6.36164 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=9.3 $Y=1.97 $X2=9.3
+ $Y2=2.19
r206 57 72 5.2253 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=9.3 $Y=0.96 $X2=9.3
+ $Y2=0.777
r207 57 58 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=9.3 $Y=0.96
+ $X2=9.3 $Y2=1.97
r208 53 66 4.04531 $w=2.5e-07 $l=2.2e-07 $layer=LI1_cond $X=8.81 $Y=2.41
+ $X2=8.81 $Y2=2.19
r209 53 55 2.99635 $w=2.48e-07 $l=6.5e-08 $layer=LI1_cond $X=8.81 $Y=2.41
+ $X2=8.81 $Y2=2.475
r210 51 82 15.6043 $w=2.78e-07 $l=9e-08 $layer=POLY_cond $X=7.785 $Y=2.257
+ $X2=7.875 $Y2=2.257
r211 51 80 56.3489 $w=2.78e-07 $l=3.25e-07 $layer=POLY_cond $X=7.785 $Y=2.257
+ $X2=7.46 $Y2=2.257
r212 50 65 34.5733 $w=2.98e-07 $l=9e-07 $layer=LI1_cond $X=7.785 $Y=2.23
+ $X2=8.685 $Y2=2.23
r213 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.785
+ $Y=2.215 $X2=7.785 $Y2=2.215
r214 44 46 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=11.71 $Y=1.9
+ $X2=11.95 $Y2=1.9
r215 39 41 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=11.71 $Y=0.94
+ $X2=12.005 $Y2=0.94
r216 35 37 41.0213 $w=1.5e-07 $l=8e-08 $layer=POLY_cond $X=7.875 $Y=1.81
+ $X2=7.955 $Y2=1.81
r217 32 41 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.005 $Y=0.865
+ $X2=12.005 $Y2=0.94
r218 32 34 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=12.005 $Y=0.865
+ $X2=12.005 $Y2=0.58
r219 29 46 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.95 $Y=1.975
+ $X2=11.95 $Y2=1.9
r220 29 31 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=11.95 $Y=1.975
+ $X2=11.95 $Y2=2.47
r221 28 44 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.71 $Y=1.825
+ $X2=11.71 $Y2=1.9
r222 27 43 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.71 $Y=1.65
+ $X2=11.71 $Y2=1.485
r223 27 28 89.734 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=11.71 $Y=1.65
+ $X2=11.71 $Y2=1.825
r224 26 43 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.71 $Y=1.32
+ $X2=11.71 $Y2=1.485
r225 25 39 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.71 $Y=1.015
+ $X2=11.71 $Y2=0.94
r226 25 26 156.394 $w=1.5e-07 $l=3.05e-07 $layer=POLY_cond $X=11.71 $Y=1.015
+ $X2=11.71 $Y2=1.32
r227 24 85 10.6442 $w=3.99e-07 $l=9.94987e-08 $layer=POLY_cond $X=11.09 $Y=1.485
+ $X2=11.015 $Y2=1.542
r228 23 43 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=11.635 $Y=1.485
+ $X2=11.71 $Y2=1.485
r229 23 24 95.2994 $w=3.3e-07 $l=5.45e-07 $layer=POLY_cond $X=11.635 $Y=1.485
+ $X2=11.09 $Y2=1.485
r230 19 85 25.8008 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=11.015 $Y=1.32
+ $X2=11.015 $Y2=1.542
r231 19 21 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=11.015 $Y=1.32
+ $X2=11.015 $Y2=0.74
r232 16 84 25.8008 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=10.98 $Y=1.765
+ $X2=10.98 $Y2=1.542
r233 16 18 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=10.98 $Y=1.765
+ $X2=10.98 $Y2=2.4
r234 12 37 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.955 $Y=1.735
+ $X2=7.955 $Y2=1.81
r235 12 14 592.245 $w=1.5e-07 $l=1.155e-06 $layer=POLY_cond $X=7.955 $Y=1.735
+ $X2=7.955 $Y2=0.58
r236 11 82 17.1848 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.875 $Y=2.05
+ $X2=7.875 $Y2=2.257
r237 10 35 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.875 $Y=1.885
+ $X2=7.875 $Y2=1.81
r238 10 11 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.875 $Y=1.885
+ $X2=7.875 $Y2=2.05
r239 7 80 17.1848 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=7.46 $Y=2.465
+ $X2=7.46 $Y2=2.257
r240 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.46 $Y=2.465 $X2=7.46
+ $Y2=2.75
r241 2 64 600 $w=1.7e-07 $l=2.89569e-07 $layer=licon1_PDIFF $count=1 $X=8.555
+ $Y=1.96 $X2=8.77 $Y2=2.135
r242 2 55 300 $w=1.7e-07 $l=6.13148e-07 $layer=licon1_PDIFF $count=2 $X=8.555
+ $Y=1.96 $X2=8.77 $Y2=2.475
r243 1 70 182 $w=1.7e-07 $l=4.71964e-07 $layer=licon1_NDIFF $count=1 $X=9.04
+ $Y=0.37 $X2=9.185 $Y2=0.775
.ends

.subckt PM_SKY130_FD_SC_LS__DFBBP_1%A_1311_424# 1 2 9 11 12 14 17 21 24 25 27 32
+ 34 35 43 46
c108 32 0 4.99671e-20 $X=7.025 $Y=2.195
c109 27 0 1.01328e-19 $X=8.78 $Y=1.215
c110 24 0 1.59361e-19 $X=7.025 $Y=2.11
r111 43 47 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.945 $Y=1.385
+ $X2=8.945 $Y2=1.55
r112 43 46 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.945 $Y=1.385
+ $X2=8.945 $Y2=1.22
r113 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.945
+ $Y=1.385 $X2=8.945 $Y2=1.385
r114 35 37 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=7.985 $Y=1.215
+ $X2=7.985 $Y2=1.485
r115 30 32 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=6.705 $Y=2.195
+ $X2=7.025 $Y2=2.195
r116 28 35 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.07 $Y=1.215
+ $X2=7.985 $Y2=1.215
r117 27 42 7.39303 $w=2.63e-07 $l=1.7e-07 $layer=LI1_cond $X=8.912 $Y=1.215
+ $X2=8.912 $Y2=1.385
r118 27 28 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=8.78 $Y=1.215
+ $X2=8.07 $Y2=1.215
r119 26 34 1.97946 $w=1.7e-07 $l=1.18e-07 $layer=LI1_cond $X=7.175 $Y=1.485
+ $X2=7.057 $Y2=1.485
r120 25 37 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.9 $Y=1.485
+ $X2=7.985 $Y2=1.485
r121 25 26 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=7.9 $Y=1.485
+ $X2=7.175 $Y2=1.485
r122 24 32 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.025 $Y=2.11
+ $X2=7.025 $Y2=2.195
r123 23 34 4.45556 $w=2.02e-07 $l=9.97246e-08 $layer=LI1_cond $X=7.025 $Y=1.57
+ $X2=7.057 $Y2=1.485
r124 23 24 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=7.025 $Y=1.57
+ $X2=7.025 $Y2=2.11
r125 19 34 4.45556 $w=2.02e-07 $l=8.5e-08 $layer=LI1_cond $X=7.057 $Y=1.4
+ $X2=7.057 $Y2=1.485
r126 19 21 31.3857 $w=2.33e-07 $l=6.4e-07 $layer=LI1_cond $X=7.057 $Y=1.4
+ $X2=7.057 $Y2=0.76
r127 17 30 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=6.705 $Y=2.65
+ $X2=6.705 $Y2=2.28
r128 12 14 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=8.995 $Y=1.885
+ $X2=8.995 $Y2=2.46
r129 11 12 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=8.995 $Y=1.795
+ $X2=8.995 $Y2=1.885
r130 11 47 95.2339 $w=1.8e-07 $l=2.45e-07 $layer=POLY_cond $X=8.995 $Y=1.795
+ $X2=8.995 $Y2=1.55
r131 9 46 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=8.965 $Y=0.74
+ $X2=8.965 $Y2=1.22
r132 2 30 600 $w=1.7e-07 $l=2.12132e-07 $layer=licon1_PDIFF $count=1 $X=6.555
+ $Y=2.12 $X2=6.705 $Y2=2.27
r133 2 17 600 $w=1.7e-07 $l=6.00333e-07 $layer=licon1_PDIFF $count=1 $X=6.555
+ $Y=2.12 $X2=6.705 $Y2=2.65
r134 1 21 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=6.95
+ $Y=0.595 $X2=7.09 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_LS__DFBBP_1%RESET_B 3 5 7 10 11 14 15
c46 14 0 1.55842e-19 $X=10.415 $Y=1.145
r47 14 15 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=10.415
+ $Y=1.145 $X2=10.415 $Y2=1.145
r48 11 15 1.69593 $w=6.68e-07 $l=9.5e-08 $layer=LI1_cond $X=10.32 $Y=1.315
+ $X2=10.415 $Y2=1.315
r49 10 14 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=10.415 $Y=1.485
+ $X2=10.415 $Y2=1.145
r50 9 14 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.415 $Y=0.98
+ $X2=10.415 $Y2=1.145
r51 5 10 50.3582 $w=2.68e-07 $l=3.03974e-07 $layer=POLY_cond $X=10.465 $Y=1.765
+ $X2=10.415 $Y2=1.485
r52 5 7 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=10.465 $Y=1.765
+ $X2=10.465 $Y2=2.16
r53 3 9 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=10.435 $Y=0.58
+ $X2=10.435 $Y2=0.98
.ends

.subckt PM_SKY130_FD_SC_LS__DFBBP_1%A_2320_410# 1 2 7 9 12 15 19 23 25 29 32 33
c62 33 0 1.92742e-19 $X=11.765 $Y=2.03
c63 15 0 1.21275e-19 $X=12.375 $Y=1.42
r64 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.19
+ $Y=1.42 $X2=12.19 $Y2=1.42
r65 27 32 0.341012 $w=3.3e-07 $l=1.18e-07 $layer=LI1_cond $X=11.875 $Y=1.42
+ $X2=11.757 $Y2=1.42
r66 27 29 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=11.875 $Y=1.42
+ $X2=12.19 $Y2=1.42
r67 23 33 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=11.765 $Y=2.155
+ $X2=11.765 $Y2=2.03
r68 23 25 1.84391 $w=2.48e-07 $l=4e-08 $layer=LI1_cond $X=11.765 $Y=2.155
+ $X2=11.765 $Y2=2.195
r69 21 32 7.59124 $w=2.02e-07 $l=1.80291e-07 $layer=LI1_cond $X=11.725 $Y=1.585
+ $X2=11.757 $Y2=1.42
r70 21 33 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=11.725 $Y=1.585
+ $X2=11.725 $Y2=2.03
r71 17 32 7.59124 $w=2.02e-07 $l=1.65e-07 $layer=LI1_cond $X=11.757 $Y=1.255
+ $X2=11.757 $Y2=1.42
r72 17 19 33.1021 $w=2.33e-07 $l=6.75e-07 $layer=LI1_cond $X=11.757 $Y=1.255
+ $X2=11.757 $Y2=0.58
r73 15 30 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=12.375 $Y=1.42
+ $X2=12.19 $Y2=1.42
r74 15 16 66.2869 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=12.465 $Y=1.42
+ $X2=12.465 $Y2=1.255
r75 12 16 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=12.48 $Y=0.74
+ $X2=12.48 $Y2=1.255
r76 7 15 136.255 $w=1.8e-07 $l=3.45e-07 $layer=POLY_cond $X=12.465 $Y=1.765
+ $X2=12.465 $Y2=1.42
r77 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=12.465 $Y=1.765
+ $X2=12.465 $Y2=2.4
r78 2 25 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=11.6
+ $Y=2.05 $X2=11.725 $Y2=2.195
r79 1 19 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=11.645
+ $Y=0.37 $X2=11.79 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_LS__DFBBP_1%VPWR 1 2 3 4 5 6 7 8 29 35 39 43 47 51 55 60
+ 61 62 64 69 77 94 98 105 106 109 112 115 118 123 129 131 134
c148 35 0 7.24936e-20 $X=2.29 $Y=2.59
r149 134 135 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r150 131 132 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r151 127 129 8.95 $w=7.63e-07 $l=2e-08 $layer=LI1_cond $X=8.4 $Y=3.032 $X2=8.42
+ $Y2=3.032
r152 127 128 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r153 125 127 2.26708 $w=7.63e-07 $l=1.45e-07 $layer=LI1_cond $X=8.255 $Y=3.032
+ $X2=8.4 $Y2=3.032
r154 122 128 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r155 121 125 5.23773 $w=7.63e-07 $l=3.35e-07 $layer=LI1_cond $X=7.92 $Y=3.032
+ $X2=8.255 $Y2=3.032
r156 121 123 13.3278 $w=7.63e-07 $l=3e-07 $layer=LI1_cond $X=7.92 $Y=3.032
+ $X2=7.62 $Y2=3.032
r157 121 122 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r158 118 119 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r159 115 116 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r160 112 113 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r161 109 110 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r162 106 135 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=12.24 $Y2=3.33
r163 105 106 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r164 103 134 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.325 $Y=3.33
+ $X2=12.2 $Y2=3.33
r165 103 105 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=12.325 $Y=3.33
+ $X2=12.72 $Y2=3.33
r166 102 135 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=12.24 $Y2=3.33
r167 102 132 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=10.8 $Y2=3.33
r168 101 102 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r169 99 131 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.92 $Y=3.33
+ $X2=10.755 $Y2=3.33
r170 99 101 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=10.92 $Y=3.33
+ $X2=11.76 $Y2=3.33
r171 98 134 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.075 $Y=3.33
+ $X2=12.2 $Y2=3.33
r172 98 101 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=12.075 $Y=3.33
+ $X2=11.76 $Y2=3.33
r173 97 132 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=10.8 $Y2=3.33
r174 96 97 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r175 94 131 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.59 $Y=3.33
+ $X2=10.755 $Y2=3.33
r176 94 96 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=10.59 $Y=3.33
+ $X2=10.32 $Y2=3.33
r177 93 97 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=10.32 $Y2=3.33
r178 93 128 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=8.4 $Y2=3.33
r179 92 129 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=9.36 $Y=3.33
+ $X2=8.42 $Y2=3.33
r180 92 93 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r181 89 122 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r182 88 123 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=7.44 $Y=3.33
+ $X2=7.62 $Y2=3.33
r183 88 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r184 86 119 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=5.52 $Y2=3.33
r185 85 88 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=6 $Y=3.33 $X2=7.44
+ $Y2=3.33
r186 85 86 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r187 83 118 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=5.87 $Y=3.33
+ $X2=5.685 $Y2=3.33
r188 83 85 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=5.87 $Y=3.33 $X2=6
+ $Y2=3.33
r189 81 119 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r190 81 116 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r191 80 81 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r192 78 115 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.19 $Y=3.33
+ $X2=4.065 $Y2=3.33
r193 78 80 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=4.19 $Y=3.33
+ $X2=4.56 $Y2=3.33
r194 77 118 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=5.5 $Y=3.33
+ $X2=5.685 $Y2=3.33
r195 77 80 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=5.5 $Y=3.33
+ $X2=4.56 $Y2=3.33
r196 76 116 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r197 75 76 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r198 73 76 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r199 73 113 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r200 72 75 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.64 $Y=3.33 $X2=3.6
+ $Y2=3.33
r201 72 73 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r202 70 112 12.6176 $w=1.7e-07 $l=3.03e-07 $layer=LI1_cond $X=2.41 $Y=3.33
+ $X2=2.107 $Y2=3.33
r203 70 72 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=2.41 $Y=3.33
+ $X2=2.64 $Y2=3.33
r204 69 115 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.94 $Y=3.33
+ $X2=4.065 $Y2=3.33
r205 69 75 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=3.94 $Y=3.33
+ $X2=3.6 $Y2=3.33
r206 68 113 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r207 68 110 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r208 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r209 65 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.035 $Y=3.33
+ $X2=0.87 $Y2=3.33
r210 65 67 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=1.035 $Y=3.33
+ $X2=1.68 $Y2=3.33
r211 64 112 12.6176 $w=1.7e-07 $l=3.02e-07 $layer=LI1_cond $X=1.805 $Y=3.33
+ $X2=2.107 $Y2=3.33
r212 64 67 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=1.805 $Y=3.33
+ $X2=1.68 $Y2=3.33
r213 62 89 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=7.44 $Y2=3.33
r214 62 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33 $X2=6
+ $Y2=3.33
r215 60 92 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=9.47 $Y=3.33
+ $X2=9.36 $Y2=3.33
r216 60 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.47 $Y=3.33
+ $X2=9.635 $Y2=3.33
r217 59 96 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=9.8 $Y=3.33
+ $X2=10.32 $Y2=3.33
r218 59 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.8 $Y=3.33
+ $X2=9.635 $Y2=3.33
r219 55 58 19.1306 $w=2.48e-07 $l=4.15e-07 $layer=LI1_cond $X=12.2 $Y=1.985
+ $X2=12.2 $Y2=2.4
r220 53 134 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=12.2 $Y=3.245
+ $X2=12.2 $Y2=3.33
r221 53 58 38.9526 $w=2.48e-07 $l=8.45e-07 $layer=LI1_cond $X=12.2 $Y=3.245
+ $X2=12.2 $Y2=2.4
r222 49 131 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.755 $Y=3.245
+ $X2=10.755 $Y2=3.33
r223 49 51 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=10.755 $Y=3.245
+ $X2=10.755 $Y2=2.745
r224 45 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.635 $Y=3.245
+ $X2=9.635 $Y2=3.33
r225 45 47 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=9.635 $Y=3.245
+ $X2=9.635 $Y2=2.78
r226 41 118 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.685 $Y=3.245
+ $X2=5.685 $Y2=3.33
r227 41 43 20.4014 $w=3.68e-07 $l=6.55e-07 $layer=LI1_cond $X=5.685 $Y=3.245
+ $X2=5.685 $Y2=2.59
r228 37 115 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.065 $Y=3.245
+ $X2=4.065 $Y2=3.33
r229 37 39 50.477 $w=2.48e-07 $l=1.095e-06 $layer=LI1_cond $X=4.065 $Y=3.245
+ $X2=4.065 $Y2=2.15
r230 33 112 2.53987 $w=6.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.107 $Y=3.245
+ $X2=2.107 $Y2=3.33
r231 33 35 12.9493 $w=6.03e-07 $l=6.55e-07 $layer=LI1_cond $X=2.107 $Y=3.245
+ $X2=2.107 $Y2=2.59
r232 29 32 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.87 $Y=2.145
+ $X2=0.87 $Y2=2.825
r233 27 109 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.87 $Y=3.245
+ $X2=0.87 $Y2=3.33
r234 27 32 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=0.87 $Y=3.245
+ $X2=0.87 $Y2=2.825
r235 8 58 300 $w=1.7e-07 $l=4.44691e-07 $layer=licon1_PDIFF $count=2 $X=12.025
+ $Y=2.05 $X2=12.24 $Y2=2.4
r236 8 55 600 $w=1.7e-07 $l=2.45357e-07 $layer=licon1_PDIFF $count=1 $X=12.025
+ $Y=2.05 $X2=12.24 $Y2=1.985
r237 7 51 600 $w=1.7e-07 $l=1.00678e-06 $layer=licon1_PDIFF $count=1 $X=10.54
+ $Y=1.84 $X2=10.755 $Y2=2.745
r238 6 47 600 $w=1.7e-07 $l=8.91852e-07 $layer=licon1_PDIFF $count=1 $X=9.485
+ $Y=1.96 $X2=9.635 $Y2=2.78
r239 5 125 300 $w=1.7e-07 $l=8.46404e-07 $layer=licon1_PDIFF $count=2 $X=7.535
+ $Y=2.54 $X2=8.255 $Y2=2.815
r240 4 43 600 $w=1.7e-07 $l=7.79824e-07 $layer=licon1_PDIFF $count=1 $X=5.505
+ $Y=1.895 $X2=5.685 $Y2=2.59
r241 3 39 600 $w=1.7e-07 $l=3.21364e-07 $layer=licon1_PDIFF $count=1 $X=3.955
+ $Y=1.895 $X2=4.105 $Y2=2.15
r242 2 35 300 $w=1.7e-07 $l=5.866e-07 $layer=licon1_PDIFF $count=2 $X=1.825
+ $Y=2.315 $X2=2.29 $Y2=2.59
r243 1 32 400 $w=1.7e-07 $l=1.08038e-06 $layer=licon1_PDIFF $count=1 $X=0.67
+ $Y=1.84 $X2=0.87 $Y2=2.825
r244 1 29 400 $w=1.7e-07 $l=3.9246e-07 $layer=licon1_PDIFF $count=1 $X=0.67
+ $Y=1.84 $X2=0.87 $Y2=2.145
.ends

.subckt PM_SKY130_FD_SC_LS__DFBBP_1%A_422_125# 1 2 9 11 12 16 17
c49 12 0 9.68576e-20 $X=2.335 $Y=1
r50 16 17 10.552 $w=3.73e-07 $l=2.3e-07 $layer=LI1_cond $X=2.767 $Y=2.525
+ $X2=2.767 $Y2=2.295
r51 13 17 78.9412 $w=1.68e-07 $l=1.21e-06 $layer=LI1_cond $X=2.87 $Y=1.085
+ $X2=2.87 $Y2=2.295
r52 11 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.785 $Y=1
+ $X2=2.87 $Y2=1.085
r53 11 12 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=2.785 $Y=1 $X2=2.335
+ $Y2=1
r54 7 12 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.21 $Y=0.915
+ $X2=2.335 $Y2=1
r55 7 9 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=2.21 $Y=0.915 $X2=2.21
+ $Y2=0.835
r56 2 16 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=2.595
+ $Y=2.315 $X2=2.745 $Y2=2.525
r57 1 9 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.11
+ $Y=0.625 $X2=2.25 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_LS__DFBBP_1%Q_N 1 2 9 13 14 15 16 23 32
c38 32 0 1.61325e-19 $X=11.29 $Y=1.82
c39 13 0 1.55842e-19 $X=11.262 $Y=1.13
r40 21 23 1.52529 $w=3.38e-07 $l=4.5e-08 $layer=LI1_cond $X=11.29 $Y=1.99
+ $X2=11.29 $Y2=2.035
r41 15 16 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=11.29 $Y=2.405
+ $X2=11.29 $Y2=2.775
r42 14 21 0.677908 $w=3.38e-07 $l=2e-08 $layer=LI1_cond $X=11.29 $Y=1.97
+ $X2=11.29 $Y2=1.99
r43 14 32 7.96349 $w=3.38e-07 $l=1.5e-07 $layer=LI1_cond $X=11.29 $Y=1.97
+ $X2=11.29 $Y2=1.82
r44 14 15 11.8634 $w=3.38e-07 $l=3.5e-07 $layer=LI1_cond $X=11.29 $Y=2.055
+ $X2=11.29 $Y2=2.405
r45 14 23 0.677908 $w=3.38e-07 $l=2e-08 $layer=LI1_cond $X=11.29 $Y=2.055
+ $X2=11.29 $Y2=2.035
r46 13 32 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=11.375 $Y=1.13
+ $X2=11.375 $Y2=1.82
r47 7 13 9.56083 $w=3.93e-07 $l=1.97e-07 $layer=LI1_cond $X=11.262 $Y=0.933
+ $X2=11.262 $Y2=1.13
r48 7 9 12.1955 $w=3.93e-07 $l=4.18e-07 $layer=LI1_cond $X=11.262 $Y=0.933
+ $X2=11.262 $Y2=0.515
r49 2 14 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=11.055
+ $Y=1.84 $X2=11.205 $Y2=1.985
r50 2 16 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=11.055
+ $Y=1.84 $X2=11.205 $Y2=2.815
r51 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=11.09
+ $Y=0.37 $X2=11.23 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__DFBBP_1%Q 1 2 7 8 9 10 11 12 13
r14 12 13 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=12.692 $Y=2.405
+ $X2=12.692 $Y2=2.775
r15 11 12 14.4485 $w=3.33e-07 $l=4.2e-07 $layer=LI1_cond $X=12.692 $Y=1.985
+ $X2=12.692 $Y2=2.405
r16 10 11 11.0084 $w=3.33e-07 $l=3.2e-07 $layer=LI1_cond $X=12.692 $Y=1.665
+ $X2=12.692 $Y2=1.985
r17 9 10 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=12.692 $Y=1.295
+ $X2=12.692 $Y2=1.665
r18 8 9 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=12.692 $Y=0.925
+ $X2=12.692 $Y2=1.295
r19 7 8 14.1045 $w=3.33e-07 $l=4.1e-07 $layer=LI1_cond $X=12.692 $Y=0.515
+ $X2=12.692 $Y2=0.925
r20 2 13 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=12.54
+ $Y=1.84 $X2=12.69 $Y2=2.815
r21 2 11 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=12.54
+ $Y=1.84 $X2=12.69 $Y2=1.985
r22 1 7 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=12.555
+ $Y=0.37 $X2=12.695 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__DFBBP_1%VGND 1 2 3 4 5 6 7 24 26 30 33 36 40 44 48
+ 51 52 54 57 58 59 61 66 75 82 92 93 96 99 111 114
c159 30 0 6.93165e-20 $X=1.82 $Y=0.835
r160 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=0
+ $X2=10.8 $Y2=0
r161 111 112 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.4 $Y=0
+ $X2=8.4 $Y2=0
r162 104 106 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0
+ $X2=4.08 $Y2=0
r163 99 100 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0
+ $X2=1.68 $Y2=0
r164 97 100 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0
+ $X2=1.68 $Y2=0
r165 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r166 92 93 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r167 90 93 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=12.72 $Y2=0
r168 90 115 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=10.8 $Y2=0
r169 89 90 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r170 87 114 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.895 $Y=0
+ $X2=10.73 $Y2=0
r171 87 89 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=10.895 $Y=0
+ $X2=11.76 $Y2=0
r172 86 115 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=10.8 $Y2=0
r173 86 112 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=8.4 $Y2=0
r174 85 86 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r175 83 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.415 $Y=0
+ $X2=8.25 $Y2=0
r176 83 85 124.283 $w=1.68e-07 $l=1.905e-06 $layer=LI1_cond $X=8.415 $Y=0
+ $X2=10.32 $Y2=0
r177 82 114 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.565 $Y=0
+ $X2=10.73 $Y2=0
r178 82 85 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=10.565 $Y=0
+ $X2=10.32 $Y2=0
r179 81 112 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.4
+ $Y2=0
r180 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r181 77 80 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=6.48 $Y=0 $X2=7.92
+ $Y2=0
r182 75 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.085 $Y=0
+ $X2=8.25 $Y2=0
r183 75 80 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=8.085 $Y=0
+ $X2=7.92 $Y2=0
r184 74 106 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6 $Y=0 $X2=4.08
+ $Y2=0
r185 73 74 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6
+ $Y2=0
r186 71 73 120.369 $w=1.68e-07 $l=1.845e-06 $layer=LI1_cond $X=4.155 $Y=0 $X2=6
+ $Y2=0
r187 70 104 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=3.6 $Y2=0
r188 70 100 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=1.68 $Y2=0
r189 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r190 67 99 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.905 $Y=0 $X2=1.78
+ $Y2=0
r191 67 69 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.905 $Y=0
+ $X2=2.16 $Y2=0
r192 66 108 9.54852 $w=5.93e-07 $l=4.75e-07 $layer=LI1_cond $X=3.857 $Y=0
+ $X2=3.857 $Y2=0.475
r193 66 71 8.26286 $w=1.7e-07 $l=2.98e-07 $layer=LI1_cond $X=3.857 $Y=0
+ $X2=4.155 $Y2=0
r194 66 106 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r195 66 104 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r196 66 69 91.3369 $w=1.68e-07 $l=1.4e-06 $layer=LI1_cond $X=3.56 $Y=0 $X2=2.16
+ $Y2=0
r197 64 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r198 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r199 61 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.78
+ $Y2=0
r200 61 63 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=0
+ $X2=0.24 $Y2=0
r201 59 81 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=6.48 $Y=0
+ $X2=7.92 $Y2=0
r202 59 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r203 59 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r204 57 89 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=12.055 $Y=0
+ $X2=11.76 $Y2=0
r205 57 58 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.055 $Y=0
+ $X2=12.18 $Y2=0
r206 56 92 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=12.305 $Y=0
+ $X2=12.72 $Y2=0
r207 56 58 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.305 $Y=0
+ $X2=12.18 $Y2=0
r208 54 55 6.55957 $w=3.68e-07 $l=1.65e-07 $layer=LI1_cond $X=6.245 $Y=0.505
+ $X2=6.245 $Y2=0.67
r209 51 73 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=6.06 $Y=0 $X2=6 $Y2=0
r210 51 52 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=6.06 $Y=0 $X2=6.245
+ $Y2=0
r211 50 77 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=6.43 $Y=0 $X2=6.48
+ $Y2=0
r212 50 52 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=6.43 $Y=0 $X2=6.245
+ $Y2=0
r213 46 58 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=12.18 $Y=0.085
+ $X2=12.18 $Y2=0
r214 46 48 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=12.18 $Y=0.085
+ $X2=12.18 $Y2=0.58
r215 42 114 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.73 $Y=0.085
+ $X2=10.73 $Y2=0
r216 42 44 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=10.73 $Y=0.085
+ $X2=10.73 $Y2=0.58
r217 38 111 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.25 $Y=0.085
+ $X2=8.25 $Y2=0
r218 38 40 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=8.25 $Y=0.085
+ $X2=8.25 $Y2=0.495
r219 36 55 12.0046 $w=2.38e-07 $l=2.5e-07 $layer=LI1_cond $X=6.31 $Y=0.92
+ $X2=6.31 $Y2=0.67
r220 33 54 0.622942 $w=3.68e-07 $l=2e-08 $layer=LI1_cond $X=6.245 $Y=0.485
+ $X2=6.245 $Y2=0.505
r221 32 52 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.245 $Y=0.085
+ $X2=6.245 $Y2=0
r222 32 33 12.4588 $w=3.68e-07 $l=4e-07 $layer=LI1_cond $X=6.245 $Y=0.085
+ $X2=6.245 $Y2=0.485
r223 28 99 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.78 $Y=0.085
+ $X2=1.78 $Y2=0
r224 28 30 34.5733 $w=2.48e-07 $l=7.5e-07 $layer=LI1_cond $X=1.78 $Y=0.085
+ $X2=1.78 $Y2=0.835
r225 27 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=0.78
+ $Y2=0
r226 26 99 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.655 $Y=0 $X2=1.78
+ $Y2=0
r227 26 27 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=1.655 $Y=0
+ $X2=0.945 $Y2=0
r228 22 96 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=0.085
+ $X2=0.78 $Y2=0
r229 22 24 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.78 $Y=0.085
+ $X2=0.78 $Y2=0.515
r230 7 48 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=12.08
+ $Y=0.37 $X2=12.22 $Y2=0.58
r231 6 44 182 $w=1.7e-07 $l=3.07571e-07 $layer=licon1_NDIFF $count=1 $X=10.51
+ $Y=0.37 $X2=10.73 $Y2=0.58
r232 5 40 91 $w=1.7e-07 $l=2.755e-07 $layer=licon1_NDIFF $count=2 $X=8.03
+ $Y=0.37 $X2=8.25 $Y2=0.495
r233 4 54 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=6.085
+ $Y=0.36 $X2=6.225 $Y2=0.505
r234 4 36 182 $w=1.7e-07 $l=6.58787e-07 $layer=licon1_NDIFF $count=1 $X=6.085
+ $Y=0.36 $X2=6.3 $Y2=0.92
r235 3 108 182 $w=1.7e-07 $l=4.05586e-07 $layer=licon1_NDIFF $count=1 $X=3.505
+ $Y=0.595 $X2=3.855 $Y2=0.475
r236 2 30 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=1.675
+ $Y=0.625 $X2=1.82 $Y2=0.835
r237 1 24 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=0.57
+ $Y=0.37 $X2=0.78 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__DFBBP_1%A_872_119# 1 2 7 9 14
r27 14 17 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=5.675 $Y=0.34
+ $X2=5.675 $Y2=0.5
r28 9 12 3.79463 $w=4.08e-07 $l=1.35e-07 $layer=LI1_cond $X=4.62 $Y=0.34
+ $X2=4.62 $Y2=0.475
r29 8 9 5.92876 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=4.825 $Y=0.34 $X2=4.62
+ $Y2=0.34
r30 7 14 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.51 $Y=0.34
+ $X2=5.675 $Y2=0.34
r31 7 8 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=5.51 $Y=0.34
+ $X2=4.825 $Y2=0.34
r32 2 17 182 $w=1.7e-07 $l=2.58167e-07 $layer=licon1_NDIFF $count=1 $X=5.46
+ $Y=0.595 $X2=5.675 $Y2=0.5
r33 1 12 182 $w=1.7e-07 $l=3.14325e-07 $layer=licon1_NDIFF $count=1 $X=4.36
+ $Y=0.595 $X2=4.62 $Y2=0.475
.ends

.subckt PM_SKY130_FD_SC_LS__DFBBP_1%A_1708_74# 1 2 9 11 12 15
c29 15 0 9.47353e-20 $X=9.64 $Y=0.515
r30 13 15 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=9.64 $Y=0.425 $X2=9.64
+ $Y2=0.515
r31 11 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.555 $Y=0.34
+ $X2=9.64 $Y2=0.425
r32 11 12 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=9.555 $Y=0.34
+ $X2=8.915 $Y2=0.34
r33 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.75 $Y=0.425
+ $X2=8.915 $Y2=0.34
r34 7 9 2.44458 $w=3.28e-07 $l=7e-08 $layer=LI1_cond $X=8.75 $Y=0.425 $X2=8.75
+ $Y2=0.495
r35 2 15 91 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=2 $X=9.475
+ $Y=0.37 $X2=9.64 $Y2=0.515
r36 1 9 91 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=2 $X=8.54
+ $Y=0.37 $X2=8.75 $Y2=0.495
.ends

