* File: sky130_fd_sc_ls__a311o_2.spice
* Created: Fri Aug 28 12:57:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__a311o_2.pex.spice"
.subckt sky130_fd_sc_ls__a311o_2  VNB VPB A3 A2 A1 B1 C1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* C1	C1
* B1	B1
* A1	A1
* A2	A2
* A3	A3
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_A_21_270#_M1003_g N_X_M1003_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1961 AS=0.1036 PD=2.01 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75003.2 A=0.111 P=1.78 MULT=1
MM1009 N_VGND_M1009_d N_A_21_270#_M1009_g N_X_M1003_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1554 AS=0.1036 PD=1.16 PS=1.02 NRD=17.016 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75002.7 A=0.111 P=1.78 MULT=1
MM1006 A_351_74# N_A3_M1006_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.74 AD=0.0777
+ AS=0.1554 PD=0.95 PS=1.16 NRD=8.1 NRS=5.664 M=1 R=4.93333 SA=75001.2
+ SB=75002.2 A=0.111 P=1.78 MULT=1
MM1001 A_423_74# N_A2_M1001_g A_351_74# VNB NSHORT L=0.15 W=0.74 AD=0.1443
+ AS=0.0777 PD=1.13 PS=0.95 NRD=22.692 NRS=8.1 M=1 R=4.93333 SA=75001.6
+ SB=75001.8 A=0.111 P=1.78 MULT=1
MM1012 N_A_21_270#_M1012_d N_A1_M1012_g A_423_74# VNB NSHORT L=0.15 W=0.74
+ AD=0.1443 AS=0.1443 PD=1.13 PS=1.13 NRD=3.24 NRS=22.692 M=1 R=4.93333
+ SA=75002.1 SB=75001.3 A=0.111 P=1.78 MULT=1
MM1004 N_VGND_M1004_d N_B1_M1004_g N_A_21_270#_M1012_d VNB NSHORT L=0.15 W=0.74
+ AD=0.1443 AS=0.1443 PD=1.13 PS=1.13 NRD=3.24 NRS=14.592 M=1 R=4.93333
+ SA=75002.6 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1008 N_A_21_270#_M1008_d N_C1_M1008_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.74
+ AD=0.1961 AS=0.1443 PD=2.01 PS=1.13 NRD=0 NRS=14.592 M=1 R=4.93333 SA=75003.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1007 N_VPWR_M1007_d N_A_21_270#_M1007_g N_X_M1007_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.308 AS=0.168 PD=2.79 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75003 A=0.168 P=2.54 MULT=1
MM1010 N_VPWR_M1010_d N_A_21_270#_M1010_g N_X_M1007_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.212906 AS=0.168 PD=1.57434 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.6 SB=75002.5 A=0.168 P=2.54 MULT=1
MM1013 N_A_330_392#_M1013_d N_A3_M1013_g N_VPWR_M1010_d VPB PHIGHVT L=0.15 W=1
+ AD=0.165 AS=0.190094 PD=1.33 PS=1.40566 NRD=1.9503 NRS=15.7403 M=1 R=6.66667
+ SA=75001.2 SB=75002.3 A=0.15 P=2.3 MULT=1
MM1000 N_VPWR_M1000_d N_A2_M1000_g N_A_330_392#_M1013_d VPB PHIGHVT L=0.15 W=1
+ AD=0.27 AS=0.165 PD=1.54 PS=1.33 NRD=25.5903 NRS=7.8603 M=1 R=6.66667
+ SA=75001.6 SB=75001.8 A=0.15 P=2.3 MULT=1
MM1011 N_A_330_392#_M1011_d N_A1_M1011_g N_VPWR_M1000_d VPB PHIGHVT L=0.15 W=1
+ AD=0.165 AS=0.27 PD=1.33 PS=1.54 NRD=7.8603 NRS=25.5903 M=1 R=6.66667
+ SA=75002.3 SB=75001.1 A=0.15 P=2.3 MULT=1
MM1005 A_660_392# N_B1_M1005_g N_A_330_392#_M1011_d VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.165 PD=1.27 PS=1.33 NRD=15.7403 NRS=1.9503 M=1 R=6.66667
+ SA=75002.8 SB=75000.6 A=0.15 P=2.3 MULT=1
MM1002 N_A_21_270#_M1002_d N_C1_M1002_g A_660_392# VPB PHIGHVT L=0.15 W=1
+ AD=0.275 AS=0.135 PD=2.55 PS=1.27 NRD=1.9503 NRS=15.7403 M=1 R=6.66667
+ SA=75003.2 SB=75000.2 A=0.15 P=2.3 MULT=1
DX14_noxref VNB VPB NWDIODE A=8.742 P=13.12
*
.include "sky130_fd_sc_ls__a311o_2.pxi.spice"
*
.ends
*
*
