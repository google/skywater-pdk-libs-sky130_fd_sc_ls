* File: sky130_fd_sc_ls__and2b_2.pex.spice
* Created: Fri Aug 28 13:03:20 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__AND2B_2%A_N 3 5 7 8 12
c27 5 0 1.61228e-19 $X=0.505 $Y=1.765
c28 3 0 1.67496e-19 $X=0.495 $Y=0.645
r29 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.515 $X2=0.385 $Y2=1.515
r30 8 12 4.06745 $w=4.23e-07 $l=1.5e-07 $layer=LI1_cond $X=0.337 $Y=1.665
+ $X2=0.337 $Y2=1.515
r31 5 11 50.8664 $w=3.35e-07 $l=2.94958e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.407 $Y2=1.515
r32 5 7 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.26
r33 1 11 38.6365 $w=3.35e-07 $l=2.04316e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.407 $Y2=1.515
r34 1 3 361.5 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=0.495 $Y=1.35 $X2=0.495
+ $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_LS__AND2B_2%A_198_48# 1 2 9 11 13 16 18 20 24 25 26 27
+ 29 33 36 38 43
c98 18 0 3.46076e-20 $X=1.575 $Y=1.765
r99 42 43 10.1474 $w=3.8e-07 $l=8e-08 $layer=POLY_cond $X=1.495 $Y=1.532
+ $X2=1.575 $Y2=1.532
r100 41 42 46.9316 $w=3.8e-07 $l=3.7e-07 $layer=POLY_cond $X=1.125 $Y=1.532
+ $X2=1.495 $Y2=1.532
r101 40 41 7.61053 $w=3.8e-07 $l=6e-08 $layer=POLY_cond $X=1.065 $Y=1.532
+ $X2=1.125 $Y2=1.532
r102 37 43 5.70789 $w=3.8e-07 $l=4.5e-08 $layer=POLY_cond $X=1.62 $Y=1.532
+ $X2=1.575 $Y2=1.532
r103 36 39 8.64761 $w=3.98e-07 $l=1.65e-07 $layer=LI1_cond $X=1.655 $Y=1.465
+ $X2=1.655 $Y2=1.63
r104 36 38 8.64761 $w=3.98e-07 $l=1.65e-07 $layer=LI1_cond $X=1.655 $Y=1.465
+ $X2=1.655 $Y2=1.3
r105 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.62
+ $Y=1.465 $X2=1.62 $Y2=1.465
r106 31 33 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=3.055 $Y=0.84
+ $X2=3.055 $Y2=0.515
r107 27 29 31.898 $w=2.78e-07 $l=7.75e-07 $layer=LI1_cond $X=1.855 $Y=2.01
+ $X2=2.63 $Y2=2.01
r108 25 31 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.89 $Y=0.925
+ $X2=3.055 $Y2=0.84
r109 25 26 67.5241 $w=1.68e-07 $l=1.035e-06 $layer=LI1_cond $X=2.89 $Y=0.925
+ $X2=1.855 $Y2=0.925
r110 24 27 7.36005 $w=2.8e-07 $l=1.77482e-07 $layer=LI1_cond $X=1.77 $Y=1.87
+ $X2=1.855 $Y2=2.01
r111 24 39 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=1.77 $Y=1.87
+ $X2=1.77 $Y2=1.63
r112 21 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.77 $Y=1.01
+ $X2=1.855 $Y2=0.925
r113 21 38 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.77 $Y=1.01
+ $X2=1.77 $Y2=1.3
r114 18 43 24.6126 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=1.575 $Y=1.765
+ $X2=1.575 $Y2=1.532
r115 18 20 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.575 $Y=1.765
+ $X2=1.575 $Y2=2.4
r116 14 42 24.6126 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=1.495 $Y=1.3
+ $X2=1.495 $Y2=1.532
r117 14 16 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.495 $Y=1.3
+ $X2=1.495 $Y2=0.74
r118 11 41 24.6126 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=1.125 $Y=1.765
+ $X2=1.125 $Y2=1.532
r119 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.125 $Y=1.765
+ $X2=1.125 $Y2=2.4
r120 7 40 24.6126 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=1.065 $Y=1.3
+ $X2=1.065 $Y2=1.532
r121 7 9 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.065 $Y=1.3
+ $X2=1.065 $Y2=0.74
r122 2 29 600 $w=1.7e-07 $l=2.22711e-07 $layer=licon1_PDIFF $count=1 $X=2.48
+ $Y=1.89 $X2=2.63 $Y2=2.05
r123 1 33 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.915
+ $Y=0.37 $X2=3.055 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__AND2B_2%B 2 3 5 8 9 12 13 14
r40 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.36 $Y=1.385
+ $X2=2.36 $Y2=1.55
r41 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.36 $Y=1.385
+ $X2=2.36 $Y2=1.22
r42 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.36
+ $Y=1.385 $X2=2.36 $Y2=1.385
r43 9 13 6.22942 $w=3.68e-07 $l=2e-07 $layer=LI1_cond $X=2.16 $Y=1.365 $X2=2.36
+ $Y2=1.365
r44 8 14 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.45 $Y=0.74 $X2=2.45
+ $Y2=1.22
r45 3 5 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.405 $Y=1.815
+ $X2=2.405 $Y2=2.39
r46 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.405 $Y=1.725 $X2=2.405
+ $Y2=1.815
r47 2 15 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=2.405 $Y=1.725
+ $X2=2.405 $Y2=1.55
.ends

.subckt PM_SKY130_FD_SC_LS__AND2B_2%A_27_74# 1 2 9 11 13 16 18 19 21 22 23 25 33
r84 30 33 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=2.93 $Y=1.465
+ $X2=3.05 $Y2=1.465
r85 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.93
+ $Y=1.465 $X2=2.93 $Y2=1.465
r86 27 28 10.1828 $w=6.29e-07 $l=5.25e-07 $layer=LI1_cond $X=0.28 $Y=2.325
+ $X2=0.805 $Y2=2.325
r87 24 33 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.05 $Y=1.63
+ $X2=3.05 $Y2=1.465
r88 24 25 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.05 $Y=1.63 $X2=3.05
+ $Y2=2.32
r89 23 28 9.00042 $w=6.29e-07 $l=1.18427e-07 $layer=LI1_cond $X=0.89 $Y=2.405
+ $X2=0.805 $Y2=2.325
r90 22 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.965 $Y=2.405
+ $X2=3.05 $Y2=2.32
r91 22 23 135.374 $w=1.68e-07 $l=2.075e-06 $layer=LI1_cond $X=2.965 $Y=2.405
+ $X2=0.89 $Y2=2.405
r92 21 28 8.62214 $w=1.7e-07 $l=3.75e-07 $layer=LI1_cond $X=0.805 $Y=1.95
+ $X2=0.805 $Y2=2.325
r93 20 21 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=0.805 $Y=1.18
+ $X2=0.805 $Y2=1.95
r94 18 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.72 $Y=1.095
+ $X2=0.805 $Y2=1.18
r95 18 19 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.72 $Y=1.095
+ $X2=0.445 $Y2=1.095
r96 14 19 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=1.01
+ $X2=0.445 $Y2=1.095
r97 14 16 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=0.28 $Y=1.01
+ $X2=0.28 $Y2=0.645
r98 11 31 71.0994 $w=2.76e-07 $l=3.85681e-07 $layer=POLY_cond $X=2.855 $Y=1.815
+ $X2=2.93 $Y2=1.465
r99 11 13 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.855 $Y=1.815
+ $X2=2.855 $Y2=2.39
r100 7 31 38.7914 $w=2.76e-07 $l=2.05122e-07 $layer=POLY_cond $X=2.84 $Y=1.3
+ $X2=2.93 $Y2=1.465
r101 7 9 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.84 $Y=1.3 $X2=2.84
+ $Y2=0.74
r102 2 27 300 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.115
r103 1 16 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_LS__AND2B_2%VPWR 1 2 3 14 16 18 20 22 24 30 33 43
r42 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r43 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r44 28 43 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r45 28 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r46 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r47 25 27 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=2.26 $Y=3.33
+ $X2=2.64 $Y2=3.33
r48 24 42 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=2.915 $Y=3.33
+ $X2=3.137 $Y2=3.33
r49 24 27 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.915 $Y=3.33
+ $X2=2.64 $Y2=3.33
r50 22 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r51 22 31 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r52 18 42 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=3.08 $Y=3.245
+ $X2=3.137 $Y2=3.33
r53 18 20 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=3.08 $Y=3.245 $X2=3.08
+ $Y2=2.745
r54 17 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.98 $Y=3.33
+ $X2=0.815 $Y2=3.33
r55 16 25 8.58075 $w=1.7e-07 $l=3.13e-07 $layer=LI1_cond $X=1.947 $Y=3.33
+ $X2=2.26 $Y2=3.33
r56 16 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r57 16 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r58 16 33 11.1953 $w=6.23e-07 $l=5.85e-07 $layer=LI1_cond $X=1.947 $Y=3.33
+ $X2=1.947 $Y2=2.745
r59 16 17 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=1.635 $Y=3.33
+ $X2=0.98 $Y2=3.33
r60 12 30 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=3.245
+ $X2=0.815 $Y2=3.33
r61 12 14 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=0.815 $Y=3.245
+ $X2=0.815 $Y2=2.825
r62 3 20 600 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=2.93
+ $Y=1.89 $X2=3.08 $Y2=2.745
r63 2 33 600 $w=1.7e-07 $l=1.04211e-06 $layer=licon1_PDIFF $count=1 $X=1.65
+ $Y=1.84 $X2=1.945 $Y2=2.745
r64 1 14 600 $w=1.7e-07 $l=1.09622e-06 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.84 $X2=0.815 $Y2=2.825
.ends

.subckt PM_SKY130_FD_SC_LS__AND2B_2%X 1 2 9 13 14 17 18
c36 18 0 8.17288e-20 $X=1.3 $Y=1.82
c37 17 0 1.61228e-19 $X=1.35 $Y=1.985
c38 13 0 1.20374e-19 $X=1.28 $Y=1.13
r39 17 18 8.78489 $w=4.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.3 $Y=1.985
+ $X2=1.3 $Y2=1.82
r40 14 17 1.34005 $w=4.28e-07 $l=5e-08 $layer=LI1_cond $X=1.3 $Y=2.035 $X2=1.3
+ $Y2=1.985
r41 13 18 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.2 $Y=1.13 $X2=1.2
+ $Y2=1.82
r42 7 13 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.28 $Y=0.965
+ $X2=1.28 $Y2=1.13
r43 7 9 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=1.28 $Y=0.965 $X2=1.28
+ $Y2=0.515
r44 2 17 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.2
+ $Y=1.84 $X2=1.35 $Y2=1.985
r45 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.14
+ $Y=0.37 $X2=1.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__AND2B_2%VGND 1 2 9 13 15 22 23 26 31 37
r41 36 37 10.7086 $w=6.83e-07 $l=1.65e-07 $layer=LI1_cond $X=2.235 $Y=0.257
+ $X2=2.4 $Y2=0.257
r42 33 36 1.30957 $w=6.83e-07 $l=7.5e-08 $layer=LI1_cond $X=2.16 $Y=0.257
+ $X2=2.235 $Y2=0.257
r43 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r44 29 33 8.38128 $w=6.83e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=0.257
+ $X2=2.16 $Y2=0.257
r45 29 31 8.96253 $w=6.83e-07 $l=6.5e-08 $layer=LI1_cond $X=1.68 $Y=0.257
+ $X2=1.615 $Y2=0.257
r46 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r47 23 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.16
+ $Y2=0
r48 22 37 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=3.12 $Y=0 $X2=2.4
+ $Y2=0
r49 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r50 18 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r51 17 18 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r52 15 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.78
+ $Y2=0
r53 15 17 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.24
+ $Y2=0
r54 13 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r55 13 27 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r56 13 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r57 12 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=0.78
+ $Y2=0
r58 12 31 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=1.615
+ $Y2=0
r59 7 26 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=0.085 $X2=0.78
+ $Y2=0
r60 7 9 19.2074 $w=3.28e-07 $l=5.5e-07 $layer=LI1_cond $X=0.78 $Y=0.085 $X2=0.78
+ $Y2=0.635
r61 2 36 91 $w=1.7e-07 $l=7.33928e-07 $layer=licon1_NDIFF $count=2 $X=1.57
+ $Y=0.37 $X2=2.235 $Y2=0.515
r62 1 9 182 $w=1.7e-07 $l=3.54789e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.78 $Y2=0.635
.ends

