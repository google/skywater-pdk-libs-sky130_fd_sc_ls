* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__dfbbn_1 CLK_N D RESET_B SET_B VGND VNB VPB VPWR Q Q_N
M1000 VGND a_1534_446# a_2412_410# VNB nshort w=420000u l=150000u
+  ad=1.55002e+12p pd=1.351e+07u as=1.134e+11p ps=1.38e+06u
M1001 a_595_119# a_27_74# a_523_119# VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=8.82e+10p ps=1.26e+06u
M1002 VPWR a_1534_446# a_2412_410# VPB phighvt w=840000u l=150000u
+  ad=2.57262e+12p pd=2.063e+07u as=2.394e+11p ps=2.25e+06u
M1003 a_1349_114# a_200_74# a_1297_424# VPB phighvt w=840000u l=150000u
+  ad=2.877e+11p pd=2.46e+06u as=2.016e+11p ps=2.16e+06u
M1004 a_311_119# a_200_74# a_595_119# VNB nshort w=420000u l=150000u
+  ad=5.1975e+11p pd=3.99e+06u as=0p ps=0u
M1005 VPWR RESET_B a_978_357# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1006 Q a_2412_410# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.192e+11p pd=2.81e+06u as=0p ps=0u
M1007 VPWR SET_B a_1534_446# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=5.75e+11p ps=5.15e+06u
M1008 VGND RESET_B a_978_357# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1009 Q a_2412_410# VGND VNB nshort w=740000u l=150000u
+  ad=1.998e+11p pd=2.02e+06u as=0p ps=0u
M1010 VPWR a_1534_446# a_1483_508# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1011 a_523_119# a_474_405# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_1483_508# a_27_74# a_1349_114# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND D a_311_119# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_1818_76# SET_B VGND VNB nshort w=740000u l=150000u
+  ad=5.032e+11p pd=4.56e+06u as=0p ps=0u
M1015 a_537_503# a_474_405# VPWR VPB phighvt w=420000u l=150000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1016 a_474_405# a_595_119# a_867_119# VNB nshort w=550000u l=150000u
+  ad=1.925e+11p pd=1.8e+06u as=3.4925e+11p ps=3.47e+06u
M1017 a_1297_424# a_474_405# VPWR VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_1611_140# a_200_74# a_1349_114# VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=6.2825e+11p ps=3.42e+06u
M1019 a_933_424# a_595_119# a_474_405# VPB phighvt w=840000u l=150000u
+  ad=2.016e+11p pd=2.16e+06u as=4.704e+11p ps=4.48e+06u
M1020 VPWR a_978_357# a_933_424# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_1254_119# a_474_405# VGND VNB nshort w=550000u l=150000u
+  ad=1.83125e+11p pd=1.8e+06u as=0p ps=0u
M1022 VGND SET_B a_867_119# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 Q_N a_1534_446# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1024 a_1349_114# a_27_74# a_1254_119# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 Q_N a_1534_446# VGND VNB nshort w=740000u l=150000u
+  ad=1.998e+11p pd=2.02e+06u as=0p ps=0u
M1026 a_867_119# a_978_357# a_474_405# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_474_405# SET_B VPWR VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_1534_446# a_1349_114# a_1917_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1029 a_1818_76# a_1349_114# a_1534_446# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.368e+11p ps=2.12e+06u
M1030 VPWR CLK_N a_27_74# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.192e+11p ps=2.81e+06u
M1031 a_200_74# a_27_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1032 a_1534_446# a_978_357# a_1818_76# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VGND CLK_N a_27_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1034 a_200_74# a_27_74# VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1035 a_595_119# a_200_74# a_537_503# VPB phighvt w=420000u l=150000u
+  ad=1.512e+11p pd=1.56e+06u as=0p ps=0u
M1036 a_311_119# a_27_74# a_595_119# VPB phighvt w=420000u l=150000u
+  ad=3.4845e+11p pd=3.47e+06u as=0p ps=0u
M1037 VPWR D a_311_119# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 VGND a_1534_446# a_1611_140# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_1917_392# a_978_357# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
