* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__or3_4 A B C VGND VNB VPB VPWR X
M1000 a_116_388# B a_206_388# VPB phighvt w=1e+06u l=150000u
+  ad=6.5e+11p pd=5.3e+06u as=6.85e+11p ps=5.37e+06u
M1001 X a_302_388# VGND VNB nshort w=740000u l=150000u
+  ad=4.181e+11p pd=4.09e+06u as=9.879e+11p ps=8.59e+06u
M1002 a_116_388# A VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=1.3788e+12p ps=1.127e+07u
M1003 a_206_388# B a_116_388# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND A a_302_388# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=4.625e+11p ps=4.21e+06u
M1005 X a_302_388# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=6.72e+11p pd=5.68e+06u as=0p ps=0u
M1006 VPWR A a_116_388# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND a_302_388# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND C a_302_388# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND a_302_388# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR a_302_388# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 X a_302_388# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_302_388# B VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_302_388# C a_206_388# VPB phighvt w=1e+06u l=150000u
+  ad=3e+11p pd=2.6e+06u as=0p ps=0u
M1014 VPWR a_302_388# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 X a_302_388# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_206_388# C a_302_388# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
