# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ls__dfbbn_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ls__dfbbn_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  14.40000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.955000 1.180000 2.755000 1.510000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.515000 1.770000 14.035000 1.940000 ;
        RECT 13.515000 1.940000 13.845000 2.980000 ;
        RECT 13.540000 0.350000 13.800000 0.850000 ;
        RECT 13.540000 0.850000 14.035000 1.100000 ;
        RECT 13.865000 1.100000 14.035000 1.770000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.630000 0.440000 11.985000 1.180000 ;
        RECT 11.645000 1.850000 11.985000 2.020000 ;
        RECT 11.645000 2.020000 11.815000 2.980000 ;
        RECT 11.815000 1.180000 11.985000 1.850000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.715000 1.350000 11.115000 1.780000 ;
    END
  END RESET_B
  PIN SET_B
    ANTENNAGATEAREA  0.469500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.415000 1.630000 5.745000 2.150000 ;
        RECT 8.765000 1.450000 9.160000 1.780000 ;
        RECT 8.765000 1.780000 8.995000 2.120000 ;
      LAYER mcon ;
        RECT 5.435000 1.950000 5.605000 2.120000 ;
        RECT 8.795000 1.950000 8.965000 2.120000 ;
      LAYER met1 ;
        RECT 5.375000 1.920000 5.665000 1.965000 ;
        RECT 5.375000 1.965000 9.025000 2.105000 ;
        RECT 5.375000 2.105000 5.665000 2.150000 ;
        RECT 8.735000 1.920000 9.025000 1.965000 ;
        RECT 8.735000 2.105000 9.025000 2.150000 ;
    END
  END SET_B
  PIN CLK_N
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.300000 0.495000 1.780000 ;
    END
  END CLK_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 14.400000 0.085000 ;
        RECT  0.545000  0.085000  0.875000 0.790000 ;
        RECT  2.045000  0.085000  2.440000 0.670000 ;
        RECT  5.745000  0.085000  6.075000 1.025000 ;
        RECT  8.785000  0.085000  8.955000 0.840000 ;
        RECT 10.665000  0.085000 11.450000 0.500000 ;
        RECT 12.155000  0.085000 12.405000 1.260000 ;
        RECT 13.095000  0.085000 13.370000 1.050000 ;
        RECT 13.970000  0.085000 14.300000 0.680000 ;
      LAYER mcon ;
        RECT  0.155000 -0.085000  0.325000 0.085000 ;
        RECT  0.635000 -0.085000  0.805000 0.085000 ;
        RECT  1.115000 -0.085000  1.285000 0.085000 ;
        RECT  1.595000 -0.085000  1.765000 0.085000 ;
        RECT  2.075000 -0.085000  2.245000 0.085000 ;
        RECT  2.555000 -0.085000  2.725000 0.085000 ;
        RECT  3.035000 -0.085000  3.205000 0.085000 ;
        RECT  3.515000 -0.085000  3.685000 0.085000 ;
        RECT  3.995000 -0.085000  4.165000 0.085000 ;
        RECT  4.475000 -0.085000  4.645000 0.085000 ;
        RECT  4.955000 -0.085000  5.125000 0.085000 ;
        RECT  5.435000 -0.085000  5.605000 0.085000 ;
        RECT  5.915000 -0.085000  6.085000 0.085000 ;
        RECT  6.395000 -0.085000  6.565000 0.085000 ;
        RECT  6.875000 -0.085000  7.045000 0.085000 ;
        RECT  7.355000 -0.085000  7.525000 0.085000 ;
        RECT  7.835000 -0.085000  8.005000 0.085000 ;
        RECT  8.315000 -0.085000  8.485000 0.085000 ;
        RECT  8.795000 -0.085000  8.965000 0.085000 ;
        RECT  9.275000 -0.085000  9.445000 0.085000 ;
        RECT  9.755000 -0.085000  9.925000 0.085000 ;
        RECT 10.235000 -0.085000 10.405000 0.085000 ;
        RECT 10.715000 -0.085000 10.885000 0.085000 ;
        RECT 11.195000 -0.085000 11.365000 0.085000 ;
        RECT 11.675000 -0.085000 11.845000 0.085000 ;
        RECT 12.155000 -0.085000 12.325000 0.085000 ;
        RECT 12.635000 -0.085000 12.805000 0.085000 ;
        RECT 13.115000 -0.085000 13.285000 0.085000 ;
        RECT 13.595000 -0.085000 13.765000 0.085000 ;
        RECT 14.075000 -0.085000 14.245000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 14.400000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 3.245000 14.400000 3.415000 ;
        RECT  0.635000 2.290000  0.805000 3.245000 ;
        RECT  2.295000 2.525000  2.465000 3.245000 ;
        RECT  5.055000 2.660000  5.385000 3.245000 ;
        RECT  6.095000 2.660000  6.425000 3.245000 ;
        RECT  8.010000 2.970000  8.340000 3.245000 ;
        RECT  9.105000 2.970000  9.435000 3.245000 ;
        RECT 11.115000 2.630000 11.445000 3.245000 ;
        RECT 12.015000 2.190000 12.345000 3.245000 ;
        RECT 13.065000 1.820000 13.315000 3.245000 ;
        RECT 14.045000 2.110000 14.295000 3.245000 ;
      LAYER mcon ;
        RECT  0.155000 3.245000  0.325000 3.415000 ;
        RECT  0.635000 3.245000  0.805000 3.415000 ;
        RECT  1.115000 3.245000  1.285000 3.415000 ;
        RECT  1.595000 3.245000  1.765000 3.415000 ;
        RECT  2.075000 3.245000  2.245000 3.415000 ;
        RECT  2.555000 3.245000  2.725000 3.415000 ;
        RECT  3.035000 3.245000  3.205000 3.415000 ;
        RECT  3.515000 3.245000  3.685000 3.415000 ;
        RECT  3.995000 3.245000  4.165000 3.415000 ;
        RECT  4.475000 3.245000  4.645000 3.415000 ;
        RECT  4.955000 3.245000  5.125000 3.415000 ;
        RECT  5.435000 3.245000  5.605000 3.415000 ;
        RECT  5.915000 3.245000  6.085000 3.415000 ;
        RECT  6.395000 3.245000  6.565000 3.415000 ;
        RECT  6.875000 3.245000  7.045000 3.415000 ;
        RECT  7.355000 3.245000  7.525000 3.415000 ;
        RECT  7.835000 3.245000  8.005000 3.415000 ;
        RECT  8.315000 3.245000  8.485000 3.415000 ;
        RECT  8.795000 3.245000  8.965000 3.415000 ;
        RECT  9.275000 3.245000  9.445000 3.415000 ;
        RECT  9.755000 3.245000  9.925000 3.415000 ;
        RECT 10.235000 3.245000 10.405000 3.415000 ;
        RECT 10.715000 3.245000 10.885000 3.415000 ;
        RECT 11.195000 3.245000 11.365000 3.415000 ;
        RECT 11.675000 3.245000 11.845000 3.415000 ;
        RECT 12.155000 3.245000 12.325000 3.415000 ;
        RECT 12.635000 3.245000 12.805000 3.415000 ;
        RECT 13.115000 3.245000 13.285000 3.415000 ;
        RECT 13.595000 3.245000 13.765000 3.415000 ;
        RECT 14.075000 3.245000 14.245000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 14.400000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.105000 1.950000  0.835000 2.120000 ;
      RECT  0.105000 2.120000  0.435000 2.980000 ;
      RECT  0.115000 0.350000  0.365000 0.960000 ;
      RECT  0.115000 0.960000  0.835000 1.130000 ;
      RECT  0.665000 1.130000  0.835000 1.300000 ;
      RECT  0.665000 1.300000  1.105000 1.630000 ;
      RECT  0.665000 1.630000  0.835000 1.950000 ;
      RECT  1.005000 1.820000  1.445000 2.905000 ;
      RECT  1.005000 2.905000  2.125000 3.075000 ;
      RECT  1.055000 0.350000  1.445000 1.130000 ;
      RECT  1.275000 1.130000  1.445000 1.820000 ;
      RECT  1.615000 0.575000  1.865000 0.840000 ;
      RECT  1.615000 0.840000  2.780000 1.010000 ;
      RECT  1.615000 1.010000  1.785000 2.735000 ;
      RECT  1.955000 1.685000  3.230000 1.855000 ;
      RECT  1.955000 1.855000  2.125000 2.905000 ;
      RECT  2.365000 2.025000  2.805000 2.355000 ;
      RECT  2.610000 0.255000  4.225000 0.425000 ;
      RECT  2.610000 0.425000  2.780000 0.840000 ;
      RECT  2.635000 2.355000  2.805000 2.905000 ;
      RECT  2.635000 2.905000  4.605000 3.075000 ;
      RECT  2.975000 1.855000  3.230000 2.355000 ;
      RECT  2.980000 0.595000  3.310000 0.785000 ;
      RECT  2.980000 0.785000  3.885000 0.955000 ;
      RECT  3.005000 1.125000  3.545000 1.455000 ;
      RECT  3.005000 1.455000  3.230000 1.685000 ;
      RECT  3.085000 2.565000  3.570000 2.735000 ;
      RECT  3.400000 1.625000  4.095000 1.795000 ;
      RECT  3.400000 1.795000  3.570000 2.565000 ;
      RECT  3.490000 0.425000  4.225000 0.615000 ;
      RECT  3.715000 0.955000  3.885000 1.465000 ;
      RECT  3.715000 1.465000  4.095000 1.625000 ;
      RECT  3.740000 1.965000  4.435000 2.135000 ;
      RECT  3.740000 2.135000  3.990000 2.735000 ;
      RECT  4.055000 0.615000  4.225000 1.125000 ;
      RECT  4.055000 1.125000  4.435000 1.295000 ;
      RECT  4.185000 2.305000  4.775000 2.320000 ;
      RECT  4.185000 2.320000  6.380000 2.490000 ;
      RECT  4.185000 2.490000  4.605000 2.905000 ;
      RECT  4.265000 1.295000  4.435000 1.965000 ;
      RECT  4.395000 0.265000  5.575000 0.435000 ;
      RECT  4.395000 0.435000  4.565000 0.955000 ;
      RECT  4.605000 1.125000  4.905000 1.295000 ;
      RECT  4.605000 1.295000  4.775000 2.305000 ;
      RECT  4.735000 0.605000  5.075000 1.120000 ;
      RECT  4.735000 1.120000  4.905000 1.125000 ;
      RECT  4.945000 1.610000  5.245000 1.940000 ;
      RECT  5.075000 1.290000  6.415000 1.460000 ;
      RECT  5.075000 1.460000  5.245000 1.610000 ;
      RECT  5.245000 0.435000  5.575000 1.025000 ;
      RECT  5.565000 2.490000  5.895000 2.980000 ;
      RECT  6.050000 1.630000  6.380000 2.320000 ;
      RECT  6.245000 0.340000  8.615000 0.510000 ;
      RECT  6.245000 0.510000  6.415000 1.290000 ;
      RECT  6.650000 0.680000  8.275000 1.010000 ;
      RECT  6.785000 1.180000  7.935000 1.410000 ;
      RECT  6.785000 1.410000  7.115000 1.910000 ;
      RECT  6.965000 2.100000  7.455000 2.980000 ;
      RECT  7.285000 1.720000  8.595000 1.890000 ;
      RECT  7.285000 1.890000  7.455000 2.100000 ;
      RECT  7.685000 1.410000  7.935000 1.550000 ;
      RECT  7.925000 2.060000  8.255000 2.630000 ;
      RECT  7.925000 2.630000 10.390000 2.800000 ;
      RECT  8.105000 1.010000  8.275000 1.720000 ;
      RECT  8.425000 1.890000  8.595000 2.290000 ;
      RECT  8.425000 2.290000  9.890000 2.460000 ;
      RECT  8.445000 0.510000  8.615000 1.010000 ;
      RECT  8.445000 1.010000 10.990000 1.180000 ;
      RECT  8.570000 2.800000  8.900000 2.980000 ;
      RECT  9.135000 0.255000 10.440000 0.425000 ;
      RECT  9.135000 0.425000  9.385000 0.840000 ;
      RECT  9.370000 1.180000  9.700000 1.550000 ;
      RECT  9.605000 0.595000  9.935000 0.670000 ;
      RECT  9.605000 0.670000 11.460000 0.840000 ;
      RECT  9.720000 1.720000 10.205000 1.890000 ;
      RECT  9.720000 1.890000  9.890000 2.290000 ;
      RECT  9.910000 1.470000 10.205000 1.720000 ;
      RECT 10.060000 2.290000 11.460000 2.460000 ;
      RECT 10.060000 2.460000 10.390000 2.630000 ;
      RECT 10.060000 2.800000 10.390000 2.980000 ;
      RECT 10.110000 0.425000 10.440000 0.500000 ;
      RECT 10.375000 1.180000 10.545000 1.950000 ;
      RECT 10.375000 1.950000 10.920000 2.120000 ;
      RECT 11.290000 0.840000 11.460000 1.350000 ;
      RECT 11.290000 1.350000 11.645000 1.680000 ;
      RECT 11.290000 1.680000 11.460000 2.290000 ;
      RECT 12.545000 1.820000 12.875000 2.860000 ;
      RECT 12.635000 0.350000 12.885000 1.270000 ;
      RECT 12.635000 1.270000 13.695000 1.600000 ;
      RECT 12.635000 1.600000 12.875000 1.820000 ;
    LAYER mcon ;
      RECT 3.035000 1.210000 3.205000 1.380000 ;
      RECT 6.875000 1.210000 7.045000 1.380000 ;
    LAYER met1 ;
      RECT 2.975000 1.180000 3.265000 1.225000 ;
      RECT 2.975000 1.225000 7.105000 1.365000 ;
      RECT 2.975000 1.365000 3.265000 1.410000 ;
      RECT 6.815000 1.180000 7.105000 1.225000 ;
      RECT 6.815000 1.365000 7.105000 1.410000 ;
  END
END sky130_fd_sc_ls__dfbbn_2
