* File: sky130_fd_sc_ls__o211ai_2.pex.spice
* Created: Fri Aug 28 13:43:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__O211AI_2%C1 3 5 7 10 12 14 15 19 22
c47 12 0 1.27308e-19 $X=0.985 $Y=1.765
r48 22 23 6.19714 $w=3.5e-07 $l=4.5e-08 $layer=POLY_cond $X=0.94 $Y=1.557
+ $X2=0.985 $Y2=1.557
r49 21 22 55.7743 $w=3.5e-07 $l=4.05e-07 $layer=POLY_cond $X=0.535 $Y=1.557
+ $X2=0.94 $Y2=1.557
r50 20 21 3.44286 $w=3.5e-07 $l=2.5e-08 $layer=POLY_cond $X=0.51 $Y=1.557
+ $X2=0.535 $Y2=1.557
r51 18 20 17.2143 $w=3.5e-07 $l=1.25e-07 $layer=POLY_cond $X=0.385 $Y=1.557
+ $X2=0.51 $Y2=1.557
r52 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.515 $X2=0.385 $Y2=1.515
r53 15 19 4.06745 $w=4.23e-07 $l=1.5e-07 $layer=LI1_cond $X=0.337 $Y=1.665
+ $X2=0.337 $Y2=1.515
r54 12 23 22.6286 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.985 $Y=1.765
+ $X2=0.985 $Y2=1.557
r55 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.985 $Y=1.765
+ $X2=0.985 $Y2=2.4
r56 8 22 22.6286 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.94 $Y=1.35
+ $X2=0.94 $Y2=1.557
r57 8 10 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.94 $Y=1.35 $X2=0.94
+ $Y2=0.79
r58 5 21 22.6286 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.535 $Y=1.765
+ $X2=0.535 $Y2=1.557
r59 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.535 $Y=1.765
+ $X2=0.535 $Y2=2.4
r60 1 20 22.6286 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.51 $Y=1.35
+ $X2=0.51 $Y2=1.557
r61 1 3 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.51 $Y=1.35 $X2=0.51
+ $Y2=0.79
.ends

.subckt PM_SKY130_FD_SC_LS__O211AI_2%B1 1 3 6 8 10 13 15 16 23 24
c51 24 0 1.83227e-19 $X=1.885 $Y=1.557
c52 23 0 1.27308e-19 $X=1.85 $Y=1.515
c53 13 0 1.66856e-19 $X=1.94 $Y=0.79
c54 8 0 8.69002e-20 $X=1.885 $Y=1.765
c55 6 0 1.74665e-19 $X=1.44 $Y=0.79
r56 24 25 7.06933 $w=3.75e-07 $l=5.5e-08 $layer=POLY_cond $X=1.885 $Y=1.557
+ $X2=1.94 $Y2=1.557
r57 22 24 4.49867 $w=3.75e-07 $l=3.5e-08 $layer=POLY_cond $X=1.85 $Y=1.557
+ $X2=1.885 $Y2=1.557
r58 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.85
+ $Y=1.515 $X2=1.85 $Y2=1.515
r59 20 22 52.6987 $w=3.75e-07 $l=4.1e-07 $layer=POLY_cond $X=1.44 $Y=1.557
+ $X2=1.85 $Y2=1.557
r60 19 20 0.642667 $w=3.75e-07 $l=5e-09 $layer=POLY_cond $X=1.435 $Y=1.557
+ $X2=1.44 $Y2=1.557
r61 16 23 4.55617 $w=4.28e-07 $l=1.7e-07 $layer=LI1_cond $X=1.68 $Y=1.565
+ $X2=1.85 $Y2=1.565
r62 15 16 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.565
+ $X2=1.68 $Y2=1.565
r63 11 25 24.2915 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.94 $Y=1.35
+ $X2=1.94 $Y2=1.557
r64 11 13 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.94 $Y=1.35
+ $X2=1.94 $Y2=0.79
r65 8 24 24.2915 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.885 $Y=1.765
+ $X2=1.885 $Y2=1.557
r66 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.885 $Y=1.765
+ $X2=1.885 $Y2=2.4
r67 4 20 24.2915 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.44 $Y=1.35
+ $X2=1.44 $Y2=1.557
r68 4 6 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.44 $Y=1.35 $X2=1.44
+ $Y2=0.79
r69 1 19 24.2915 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.435 $Y=1.765
+ $X2=1.435 $Y2=1.557
r70 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.435 $Y=1.765
+ $X2=1.435 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__O211AI_2%A2 1 3 6 8 10 13 15 16 19 29 31
c58 31 0 2.53756e-19 $X=3.005 $Y=1.55
c59 8 0 1.88567e-19 $X=3.345 $Y=1.765
r60 29 30 3.05838 $w=3.94e-07 $l=2.5e-08 $layer=POLY_cond $X=3.345 $Y=1.542
+ $X2=3.37 $Y2=1.542
r61 27 29 7.95178 $w=3.94e-07 $l=6.5e-08 $layer=POLY_cond $X=3.28 $Y=1.542
+ $X2=3.345 $Y2=1.542
r62 27 28 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.28
+ $Y=1.485 $X2=3.28 $Y2=1.485
r63 25 27 41.5939 $w=3.94e-07 $l=3.4e-07 $layer=POLY_cond $X=2.94 $Y=1.542
+ $X2=3.28 $Y2=1.542
r64 24 25 5.50508 $w=3.94e-07 $l=4.5e-08 $layer=POLY_cond $X=2.895 $Y=1.542
+ $X2=2.94 $Y2=1.542
r65 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.6
+ $Y=1.485 $X2=2.6 $Y2=1.485
r66 19 24 12.4234 $w=3.94e-07 $l=1.15022e-07 $layer=POLY_cond $X=2.805 $Y=1.485
+ $X2=2.895 $Y2=1.542
r67 19 21 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=2.805 $Y=1.485
+ $X2=2.6 $Y2=1.485
r68 16 28 4.91688 $w=3.97e-07 $l=1.6e-07 $layer=LI1_cond $X=3.12 $Y=1.55
+ $X2=3.28 $Y2=1.55
r69 16 31 3.3124 $w=4.6e-07 $l=1.15e-07 $layer=LI1_cond $X=3.12 $Y=1.55
+ $X2=3.005 $Y2=1.55
r70 15 31 9.49062 $w=4.58e-07 $l=3.65e-07 $layer=LI1_cond $X=2.64 $Y=1.55
+ $X2=3.005 $Y2=1.55
r71 15 22 1.04007 $w=4.58e-07 $l=4e-08 $layer=LI1_cond $X=2.64 $Y=1.55 $X2=2.6
+ $Y2=1.55
r72 11 30 25.4929 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=3.37 $Y=1.32
+ $X2=3.37 $Y2=1.542
r73 11 13 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.37 $Y=1.32
+ $X2=3.37 $Y2=0.74
r74 8 29 25.4929 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=3.345 $Y=1.765
+ $X2=3.345 $Y2=1.542
r75 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.345 $Y=1.765
+ $X2=3.345 $Y2=2.4
r76 4 25 25.4929 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=2.94 $Y=1.32
+ $X2=2.94 $Y2=1.542
r77 4 6 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.94 $Y=1.32 $X2=2.94
+ $Y2=0.74
r78 1 24 25.4929 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=2.895 $Y=1.765
+ $X2=2.895 $Y2=1.542
r79 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.895 $Y=1.765
+ $X2=2.895 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__O211AI_2%A1 1 3 6 10 12 14 20 26 31
r49 29 31 5.27442 $w=4.68e-07 $l=1.65e-07 $layer=LI1_cond $X=4.53 $Y=1.415
+ $X2=4.365 $Y2=1.415
r50 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.53
+ $Y=1.465 $X2=4.53 $Y2=1.465
r51 26 28 29.4974 $w=3.84e-07 $l=2.35e-07 $layer=POLY_cond $X=4.295 $Y=1.532
+ $X2=4.53 $Y2=1.532
r52 25 26 1.88281 $w=3.84e-07 $l=1.5e-08 $layer=POLY_cond $X=4.28 $Y=1.532
+ $X2=4.295 $Y2=1.532
r53 22 23 1.25521 $w=3.84e-07 $l=1e-08 $layer=POLY_cond $X=3.795 $Y=1.532
+ $X2=3.805 $Y2=1.532
r54 20 29 0.763454 $w=4.68e-07 $l=3e-08 $layer=LI1_cond $X=4.56 $Y=1.415
+ $X2=4.53 $Y2=1.415
r55 18 25 11.2969 $w=3.84e-07 $l=9e-08 $layer=POLY_cond $X=4.19 $Y=1.532
+ $X2=4.28 $Y2=1.532
r56 18 23 48.3255 $w=3.84e-07 $l=3.85e-07 $layer=POLY_cond $X=4.19 $Y=1.532
+ $X2=3.805 $Y2=1.532
r57 17 31 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=4.19 $Y=1.485
+ $X2=4.365 $Y2=1.485
r58 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.19
+ $Y=1.485 $X2=4.19 $Y2=1.485
r59 12 26 24.8669 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=4.295 $Y=1.765
+ $X2=4.295 $Y2=1.532
r60 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.295 $Y=1.765
+ $X2=4.295 $Y2=2.4
r61 8 25 24.8669 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=4.28 $Y=1.3 $X2=4.28
+ $Y2=1.532
r62 8 10 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.28 $Y=1.3 $X2=4.28
+ $Y2=0.74
r63 4 23 24.8669 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=3.805 $Y=1.3
+ $X2=3.805 $Y2=1.532
r64 4 6 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.805 $Y=1.3 $X2=3.805
+ $Y2=0.74
r65 1 22 24.8669 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=3.795 $Y=1.765
+ $X2=3.795 $Y2=1.532
r66 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.795 $Y=1.765
+ $X2=3.795 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__O211AI_2%VPWR 1 2 3 4 13 15 19 23 27 31 33 35 40 50
+ 51 57 60 63
c65 31 0 1.88567e-19 $X=4.02 $Y=2.325
r66 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r67 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r68 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r69 55 58 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r70 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r71 51 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r72 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r73 48 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.185 $Y=3.33
+ $X2=4.02 $Y2=3.33
r74 48 50 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=4.185 $Y=3.33
+ $X2=4.56 $Y2=3.33
r75 47 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r76 46 47 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r77 44 47 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r78 43 46 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.64 $Y=3.33 $X2=3.6
+ $Y2=3.33
r79 43 44 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r80 41 60 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.275 $Y=3.33
+ $X2=2.15 $Y2=3.33
r81 41 43 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.275 $Y=3.33
+ $X2=2.64 $Y2=3.33
r82 40 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.855 $Y=3.33
+ $X2=4.02 $Y2=3.33
r83 40 46 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=3.855 $Y=3.33
+ $X2=3.6 $Y2=3.33
r84 39 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r85 39 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r86 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r87 36 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.295 $Y=3.33
+ $X2=1.21 $Y2=3.33
r88 36 38 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=1.295 $Y=3.33
+ $X2=1.68 $Y2=3.33
r89 35 60 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.025 $Y=3.33
+ $X2=2.15 $Y2=3.33
r90 35 38 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.025 $Y=3.33
+ $X2=1.68 $Y2=3.33
r91 33 44 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=2.64 $Y2=3.33
r92 33 61 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=2.16 $Y2=3.33
r93 29 63 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.02 $Y=3.245
+ $X2=4.02 $Y2=3.33
r94 29 31 32.1287 $w=3.28e-07 $l=9.2e-07 $layer=LI1_cond $X=4.02 $Y=3.245
+ $X2=4.02 $Y2=2.325
r95 25 60 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.15 $Y=3.245
+ $X2=2.15 $Y2=3.33
r96 25 27 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=2.15 $Y=3.245
+ $X2=2.15 $Y2=2.455
r97 21 57 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.21 $Y=3.245
+ $X2=1.21 $Y2=3.33
r98 21 23 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=1.21 $Y=3.245
+ $X2=1.21 $Y2=2.455
r99 20 54 3.97288 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=0.395 $Y=3.33
+ $X2=0.197 $Y2=3.33
r100 19 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.125 $Y=3.33
+ $X2=1.21 $Y2=3.33
r101 19 20 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.125 $Y=3.33
+ $X2=0.395 $Y2=3.33
r102 15 18 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=0.27 $Y=2.115
+ $X2=0.27 $Y2=2.815
r103 13 54 3.17028 $w=2.5e-07 $l=1.15888e-07 $layer=LI1_cond $X=0.27 $Y=3.245
+ $X2=0.197 $Y2=3.33
r104 13 18 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.27 $Y=3.245
+ $X2=0.27 $Y2=2.815
r105 4 31 300 $w=1.7e-07 $l=5.54955e-07 $layer=licon1_PDIFF $count=2 $X=3.87
+ $Y=1.84 $X2=4.02 $Y2=2.325
r106 3 27 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=1.96
+ $Y=1.84 $X2=2.11 $Y2=2.455
r107 2 23 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=1.06
+ $Y=1.84 $X2=1.21 $Y2=2.455
r108 1 18 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.165
+ $Y=1.84 $X2=0.31 $Y2=2.815
r109 1 15 400 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.165
+ $Y=1.84 $X2=0.31 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_LS__O211AI_2%Y 1 2 3 4 15 18 19 23 25 29 32 34 36 37 38
c69 18 0 1.83227e-19 $X=0.805 $Y=1.95
c70 15 0 1.74665e-19 $X=0.725 $Y=0.68
r71 37 38 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.76 $Y=2.405
+ $X2=0.76 $Y2=2.775
r72 30 37 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=0.76 $Y=2.12
+ $X2=0.76 $Y2=2.405
r73 30 32 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.76 $Y=2.12 $X2=0.76
+ $Y2=2.035
r74 26 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.825 $Y=2.035
+ $X2=1.66 $Y2=2.035
r75 25 36 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.955 $Y=2.035
+ $X2=3.12 $Y2=2.035
r76 25 26 73.7219 $w=1.68e-07 $l=1.13e-06 $layer=LI1_cond $X=2.955 $Y=2.035
+ $X2=1.825 $Y2=2.035
r77 21 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.66 $Y=2.12 $X2=1.66
+ $Y2=2.035
r78 21 23 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=1.66 $Y=2.12
+ $X2=1.66 $Y2=2.815
r79 20 32 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.925 $Y=2.035
+ $X2=0.76 $Y2=2.035
r80 19 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.495 $Y=2.035
+ $X2=1.66 $Y2=2.035
r81 19 20 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.495 $Y=2.035
+ $X2=0.925 $Y2=2.035
r82 18 32 3.70735 $w=2.5e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.805 $Y=1.95
+ $X2=0.76 $Y2=2.035
r83 18 29 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=0.805 $Y=1.95
+ $X2=0.805 $Y2=1.18
r84 13 29 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.725 $Y=1.015
+ $X2=0.725 $Y2=1.18
r85 13 15 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.725 $Y=1.015
+ $X2=0.725 $Y2=0.68
r86 4 36 300 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=2 $X=2.97
+ $Y=1.84 $X2=3.12 $Y2=2.115
r87 3 34 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=1.51
+ $Y=1.84 $X2=1.66 $Y2=2.115
r88 3 23 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.51
+ $Y=1.84 $X2=1.66 $Y2=2.815
r89 2 38 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=0.61
+ $Y=1.84 $X2=0.76 $Y2=2.815
r90 2 32 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=0.61
+ $Y=1.84 $X2=0.76 $Y2=2.115
r91 1 15 91 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_NDIFF $count=2 $X=0.585
+ $Y=0.42 $X2=0.725 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_LS__O211AI_2%A_505_368# 1 2 3 12 14 15 16 19 20 22 24
r44 22 29 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.52 $Y=1.99 $X2=4.52
+ $Y2=1.905
r45 22 24 28.8111 $w=3.28e-07 $l=8.25e-07 $layer=LI1_cond $X=4.52 $Y=1.99
+ $X2=4.52 $Y2=2.815
r46 21 27 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.655 $Y=1.905
+ $X2=3.57 $Y2=1.905
r47 20 29 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.355 $Y=1.905
+ $X2=4.52 $Y2=1.905
r48 20 21 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=4.355 $Y=1.905
+ $X2=3.655 $Y2=1.905
r49 17 19 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=3.57 $Y=2.905 $X2=3.57
+ $Y2=2.815
r50 16 27 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.57 $Y=1.99 $X2=3.57
+ $Y2=1.905
r51 16 19 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=3.57 $Y=1.99
+ $X2=3.57 $Y2=2.815
r52 14 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.485 $Y=2.99
+ $X2=3.57 $Y2=2.905
r53 14 15 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=3.485 $Y=2.99
+ $X2=2.755 $Y2=2.99
r54 10 15 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.63 $Y=2.905
+ $X2=2.755 $Y2=2.99
r55 10 12 20.744 $w=2.48e-07 $l=4.5e-07 $layer=LI1_cond $X=2.63 $Y=2.905
+ $X2=2.63 $Y2=2.455
r56 3 29 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=4.37
+ $Y=1.84 $X2=4.52 $Y2=1.985
r57 3 24 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=4.37
+ $Y=1.84 $X2=4.52 $Y2=2.815
r58 2 27 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=3.42
+ $Y=1.84 $X2=3.57 $Y2=1.985
r59 2 19 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=3.42
+ $Y=1.84 $X2=3.57 $Y2=2.815
r60 1 12 300 $w=1.7e-07 $l=6.83667e-07 $layer=licon1_PDIFF $count=2 $X=2.525
+ $Y=1.84 $X2=2.67 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_LS__O211AI_2%A_30_84# 1 2 3 12 14 15 20 23
r38 18 23 5.2656 $w=3.22e-07 $l=1.65e-07 $layer=LI1_cond $X=1.39 $Y=0.492
+ $X2=1.225 $Y2=0.492
r39 18 20 19.3891 $w=4.73e-07 $l=7.7e-07 $layer=LI1_cond $X=1.39 $Y=0.492
+ $X2=2.16 $Y2=0.492
r40 14 23 5.2656 $w=3.22e-07 $l=2.28703e-07 $layer=LI1_cond $X=1.06 $Y=0.34
+ $X2=1.225 $Y2=0.492
r41 14 15 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.06 $Y=0.34
+ $X2=0.38 $Y2=0.34
r42 10 15 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.255 $Y=0.425
+ $X2=0.38 $Y2=0.34
r43 10 12 6.45368 $w=2.48e-07 $l=1.4e-07 $layer=LI1_cond $X=0.255 $Y=0.425
+ $X2=0.255 $Y2=0.565
r44 3 20 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=2.015
+ $Y=0.42 $X2=2.16 $Y2=0.565
r45 2 23 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=1.015
+ $Y=0.42 $X2=1.225 $Y2=0.565
r46 1 12 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.15
+ $Y=0.42 $X2=0.295 $Y2=0.565
.ends

.subckt PM_SKY130_FD_SC_LS__O211AI_2%A_303_84# 1 2 3 10 14 16 20 25 26
r47 23 25 8.55689 $w=2.78e-07 $l=1.65e-07 $layer=LI1_cond $X=1.725 $Y=1.04
+ $X2=1.89 $Y2=1.04
r48 18 20 23.8172 $w=2.23e-07 $l=4.65e-07 $layer=LI1_cond $X=4.047 $Y=0.98
+ $X2=4.047 $Y2=0.515
r49 17 26 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.24 $Y=1.065
+ $X2=3.155 $Y2=1.065
r50 16 18 6.9898 $w=1.7e-07 $l=1.4854e-07 $layer=LI1_cond $X=3.935 $Y=1.065
+ $X2=4.047 $Y2=0.98
r51 16 17 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=3.935 $Y=1.065
+ $X2=3.24 $Y2=1.065
r52 12 26 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.155 $Y=0.98
+ $X2=3.155 $Y2=1.065
r53 12 14 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=3.155 $Y=0.98
+ $X2=3.155 $Y2=0.515
r54 10 26 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.07 $Y=1.065
+ $X2=3.155 $Y2=1.065
r55 10 25 76.984 $w=1.68e-07 $l=1.18e-06 $layer=LI1_cond $X=3.07 $Y=1.065
+ $X2=1.89 $Y2=1.065
r56 3 20 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.88
+ $Y=0.37 $X2=4.02 $Y2=0.515
r57 2 14 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.015
+ $Y=0.37 $X2=3.155 $Y2=0.515
r58 1 23 182 $w=1.7e-07 $l=6.76905e-07 $layer=licon1_NDIFF $count=1 $X=1.515
+ $Y=0.42 $X2=1.725 $Y2=1
.ends

.subckt PM_SKY130_FD_SC_LS__O211AI_2%VGND 1 2 3 12 16 18 20 22 24 29 34 40 43 47
r55 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r56 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r57 40 41 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r58 38 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r59 38 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r60 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r61 35 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.75 $Y=0 $X2=3.585
+ $Y2=0
r62 35 37 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=3.75 $Y=0 $X2=4.08
+ $Y2=0
r63 34 46 4.96106 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=4.33 $Y=0 $X2=4.565
+ $Y2=0
r64 34 37 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=4.33 $Y=0 $X2=4.08
+ $Y2=0
r65 33 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r66 33 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r67 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r68 30 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.89 $Y=0 $X2=2.725
+ $Y2=0
r69 30 32 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=2.89 $Y=0 $X2=3.12
+ $Y2=0
r70 29 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.42 $Y=0 $X2=3.585
+ $Y2=0
r71 29 32 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=3.42 $Y=0 $X2=3.12
+ $Y2=0
r72 26 27 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r73 24 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.56 $Y=0 $X2=2.725
+ $Y2=0
r74 24 26 151.358 $w=1.68e-07 $l=2.32e-06 $layer=LI1_cond $X=2.56 $Y=0 $X2=0.24
+ $Y2=0
r75 22 41 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=2.64
+ $Y2=0
r76 22 27 0.602067 $w=4.9e-07 $l=2.16e-06 $layer=MET1_cond $X=2.4 $Y=0 $X2=0.24
+ $Y2=0
r77 18 46 3.01886 $w=3.55e-07 $l=1.1025e-07 $layer=LI1_cond $X=4.507 $Y=0.085
+ $X2=4.565 $Y2=0
r78 18 20 13.9592 $w=3.53e-07 $l=4.3e-07 $layer=LI1_cond $X=4.507 $Y=0.085
+ $X2=4.507 $Y2=0.515
r79 14 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.585 $Y=0.085
+ $X2=3.585 $Y2=0
r80 14 16 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=3.585 $Y=0.085
+ $X2=3.585 $Y2=0.63
r81 10 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.725 $Y=0.085
+ $X2=2.725 $Y2=0
r82 10 12 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=2.725 $Y=0.085
+ $X2=2.725 $Y2=0.63
r83 3 20 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.355
+ $Y=0.37 $X2=4.495 $Y2=0.515
r84 2 16 182 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_NDIFF $count=1 $X=3.445
+ $Y=0.37 $X2=3.585 $Y2=0.63
r85 1 12 182 $w=1.7e-07 $l=3.245e-07 $layer=licon1_NDIFF $count=1 $X=2.58
+ $Y=0.37 $X2=2.725 $Y2=0.63
.ends

