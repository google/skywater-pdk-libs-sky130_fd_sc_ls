* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__a41oi_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
X0 a_277_74# A3 a_355_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X1 a_116_368# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X2 VPWR A1 a_116_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X3 a_355_74# A2 a_469_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X4 VGND A4 a_277_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X5 a_469_74# A1 Y VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X6 Y B1 a_116_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X7 a_116_368# A4 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X8 VPWR A3 a_116_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X9 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
.ends
