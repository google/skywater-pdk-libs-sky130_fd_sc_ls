* File: sky130_fd_sc_ls__dlclkp_2.pex.spice
* Created: Wed Sep  2 11:02:54 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__DLCLKP_2%A_83_244# 1 2 7 9 10 12 14 15 17 18 20 22
+ 23 25 27 29 31
c85 17 0 5.18245e-20 $X=1.535 $Y=2.035
c86 10 0 1.23149e-19 $X=0.505 $Y=1.765
r87 34 36 8.48848 $w=3.48e-07 $l=1.65e-07 $layer=LI1_cond $X=0.61 $Y=1.385
+ $X2=0.61 $Y2=1.55
r88 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.6
+ $Y=1.385 $X2=0.6 $Y2=1.385
r89 31 34 6.25612 $w=3.48e-07 $l=1.9e-07 $layer=LI1_cond $X=0.61 $Y=1.195
+ $X2=0.61 $Y2=1.385
r90 27 29 18.6835 $w=3.28e-07 $l=5.35e-07 $layer=LI1_cond $X=1.705 $Y=2.715
+ $X2=2.24 $Y2=2.715
r91 23 25 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=1.56 $Y=0.785
+ $X2=1.985 $Y2=0.785
r92 22 27 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.62 $Y=2.55
+ $X2=1.705 $Y2=2.715
r93 21 22 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=1.62 $Y=2.12
+ $X2=1.62 $Y2=2.55
r94 19 23 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.475 $Y=0.95
+ $X2=1.56 $Y2=0.785
r95 19 20 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=1.475 $Y=0.95
+ $X2=1.475 $Y2=1.11
r96 17 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.535 $Y=2.035
+ $X2=1.62 $Y2=2.12
r97 17 18 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=1.535 $Y=2.035
+ $X2=0.785 $Y2=2.035
r98 16 31 4.974 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=0.785 $Y=1.195
+ $X2=0.61 $Y2=1.195
r99 15 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.39 $Y=1.195
+ $X2=1.475 $Y2=1.11
r100 15 16 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=1.39 $Y=1.195
+ $X2=0.785 $Y2=1.195
r101 14 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.7 $Y=1.95
+ $X2=0.785 $Y2=2.035
r102 14 36 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=0.7 $Y=1.95 $X2=0.7
+ $Y2=1.55
r103 10 35 75.4509 $w=2.82e-07 $l=4.20357e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.59 $Y2=1.385
r104 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.4
r105 7 35 38.7026 $w=2.82e-07 $l=2.07123e-07 $layer=POLY_cond $X=0.495 $Y=1.22
+ $X2=0.59 $Y2=1.385
r106 7 9 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.495 $Y=1.22
+ $X2=0.495 $Y2=0.74
r107 2 29 300 $w=1.7e-07 $l=9.73409e-07 $layer=licon1_PDIFF $count=2 $X=1.74
+ $Y=1.96 $X2=2.24 $Y2=2.715
r108 1 25 182 $w=1.7e-07 $l=5.29268e-07 $layer=licon1_NDIFF $count=1 $X=1.725
+ $Y=0.37 $X2=1.985 $Y2=0.785
.ends

.subckt PM_SKY130_FD_SC_LS__DLCLKP_2%GATE 1 3 6 8
c35 8 0 1.23149e-19 $X=1.2 $Y=1.665
r36 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.17
+ $Y=1.615 $X2=1.17 $Y2=1.615
r37 4 11 38.5916 $w=2.93e-07 $l=2.05122e-07 $layer=POLY_cond $X=1.26 $Y=1.45
+ $X2=1.17 $Y2=1.615
r38 4 6 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=1.26 $Y=1.45 $X2=1.26
+ $Y2=0.69
r39 1 11 55.8646 $w=2.93e-07 $l=3.05205e-07 $layer=POLY_cond $X=1.245 $Y=1.885
+ $X2=1.17 $Y2=1.615
r40 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.245 $Y=1.885
+ $X2=1.245 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_LS__DLCLKP_2%A_315_48# 1 2 7 9 10 12 13 15 18 20 24 26
+ 28 29 32 35 44 45 51 52 54 59 61 63 65 66 74
c146 35 0 1.73462e-19 $X=4.43 $Y=0.74
c147 29 0 1.92985e-19 $X=3.155 $Y=2.135
c148 10 0 5.18245e-20 $X=2.465 $Y=2.465
c149 7 0 1.30966e-19 $X=1.65 $Y=1.12
r150 65 66 8.46614 $w=3.33e-07 $l=1.65e-07 $layer=LI1_cond $X=4.377 $Y=2.24
+ $X2=4.377 $Y2=2.075
r151 62 66 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=4.295 $Y=1.885
+ $X2=4.295 $Y2=2.075
r152 61 63 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=4.295 $Y=1.555
+ $X2=4.295 $Y2=1.275
r153 60 74 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.16 $Y=1.72 $X2=4.16
+ $Y2=1.63
r154 59 62 8.58894 $w=3.83e-07 $l=1.65e-07 $layer=LI1_cond $X=4.187 $Y=1.72
+ $X2=4.187 $Y2=1.885
r155 59 61 8.58894 $w=3.83e-07 $l=1.65e-07 $layer=LI1_cond $X=4.187 $Y=1.72
+ $X2=4.187 $Y2=1.555
r156 59 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.16
+ $Y=1.72 $X2=4.16 $Y2=1.72
r157 54 57 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.32 $Y=1.72
+ $X2=3.32 $Y2=1.885
r158 54 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.32
+ $Y=1.72 $X2=3.32 $Y2=1.72
r159 49 52 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.39 $Y=2.215
+ $X2=2.555 $Y2=2.215
r160 49 51 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.39 $Y=2.215
+ $X2=2.225 $Y2=2.215
r161 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.39
+ $Y=2.215 $X2=2.39 $Y2=2.215
r162 45 69 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=1.88 $Y=1.285
+ $X2=1.65 $Y2=1.285
r163 44 47 8.46257 $w=3.13e-07 $l=1.65e-07 $layer=LI1_cond $X=1.887 $Y=1.285
+ $X2=1.887 $Y2=1.45
r164 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.88
+ $Y=1.285 $X2=1.88 $Y2=1.285
r165 33 63 9.39714 $w=3.83e-07 $l=1.92e-07 $layer=LI1_cond $X=4.402 $Y=1.083
+ $X2=4.402 $Y2=1.275
r166 33 35 10.2672 $w=3.83e-07 $l=3.43e-07 $layer=LI1_cond $X=4.402 $Y=1.083
+ $X2=4.402 $Y2=0.74
r167 32 57 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.24 $Y=2.05
+ $X2=3.24 $Y2=1.885
r168 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.155 $Y=2.135
+ $X2=3.24 $Y2=2.05
r169 29 52 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=3.155 $Y=2.135
+ $X2=2.555 $Y2=2.135
r170 28 51 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.045 $Y=2.135
+ $X2=2.225 $Y2=2.135
r171 26 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.96 $Y=2.05
+ $X2=2.045 $Y2=2.135
r172 26 47 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=1.96 $Y=2.05 $X2=1.96
+ $Y2=1.45
r173 24 55 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=3.505 $Y=1.72
+ $X2=3.32 $Y2=1.72
r174 22 24 24.6477 $w=1.76e-07 $l=9e-08 $layer=POLY_cond $X=3.617 $Y=1.63
+ $X2=3.617 $Y2=1.72
r175 21 22 6.61437 $w=1.5e-07 $l=1.13e-07 $layer=POLY_cond $X=3.73 $Y=1.63
+ $X2=3.617 $Y2=1.63
r176 20 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.995 $Y=1.63
+ $X2=4.16 $Y2=1.63
r177 20 21 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=3.995 $Y=1.63
+ $X2=3.73 $Y2=1.63
r178 16 22 21.729 $w=1.76e-07 $l=9.20598e-08 $layer=POLY_cond $X=3.655 $Y=1.555
+ $X2=3.617 $Y2=1.63
r179 16 18 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.655 $Y=1.555
+ $X2=3.655 $Y2=0.995
r180 13 24 90.195 $w=1.76e-07 $l=3.3582e-07 $layer=POLY_cond $X=3.595 $Y=2.045
+ $X2=3.617 $Y2=1.72
r181 13 15 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=3.595 $Y=2.045
+ $X2=3.595 $Y2=2.54
r182 10 50 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=2.465 $Y=2.465
+ $X2=2.39 $Y2=2.215
r183 10 12 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.465 $Y=2.465
+ $X2=2.465 $Y2=2.75
r184 7 69 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.65 $Y=1.12
+ $X2=1.65 $Y2=1.285
r185 7 9 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.65 $Y=1.12 $X2=1.65
+ $Y2=0.69
r186 2 65 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=4.235
+ $Y=2.095 $X2=4.38 $Y2=2.24
r187 1 35 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=4.285
+ $Y=0.595 $X2=4.43 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__DLCLKP_2%A_315_338# 1 2 7 9 10 11 14 18 19 21 22 27
+ 31 33 34
c98 27 0 6.54874e-20 $X=3.82 $Y=2.265
c99 19 0 1.92985e-19 $X=2.42 $Y=1.675
r100 29 33 3.70735 $w=2.5e-07 $l=9.66954e-08 $layer=LI1_cond $X=3.87 $Y=1.215
+ $X2=3.845 $Y2=1.3
r101 29 31 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=3.87 $Y=1.215
+ $X2=3.87 $Y2=0.77
r102 27 34 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.82 $Y=2.265
+ $X2=3.82 $Y2=2.1
r103 23 33 3.70735 $w=2.5e-07 $l=1.41244e-07 $layer=LI1_cond $X=3.74 $Y=1.385
+ $X2=3.845 $Y2=1.3
r104 23 34 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=3.74 $Y=1.385
+ $X2=3.74 $Y2=2.1
r105 21 33 2.76166 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.655 $Y=1.3
+ $X2=3.845 $Y2=1.3
r106 21 22 69.8075 $w=1.68e-07 $l=1.07e-06 $layer=LI1_cond $X=3.655 $Y=1.3
+ $X2=2.585 $Y2=1.3
r107 19 37 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.42 $Y=1.675
+ $X2=2.42 $Y2=1.765
r108 19 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.42 $Y=1.675
+ $X2=2.42 $Y2=1.51
r109 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.42
+ $Y=1.675 $X2=2.42 $Y2=1.675
r110 16 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.42 $Y=1.385
+ $X2=2.585 $Y2=1.3
r111 16 18 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=2.42 $Y=1.385
+ $X2=2.42 $Y2=1.675
r112 14 36 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=2.395 $Y=0.8
+ $X2=2.395 $Y2=1.51
r113 10 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.255 $Y=1.765
+ $X2=2.42 $Y2=1.765
r114 10 11 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=2.255 $Y=1.765
+ $X2=1.755 $Y2=1.765
r115 7 11 26.9307 $w=1.5e-07 $l=1.58745e-07 $layer=POLY_cond $X=1.665 $Y=1.885
+ $X2=1.755 $Y2=1.765
r116 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.665 $Y=1.885
+ $X2=1.665 $Y2=2.46
r117 2 27 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=3.67
+ $Y=2.12 $X2=3.82 $Y2=2.265
r118 1 31 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.73
+ $Y=0.625 $X2=3.87 $Y2=0.77
.ends

.subckt PM_SKY130_FD_SC_LS__DLCLKP_2%CLK 2 3 5 6 8 9 11 12 14 15 22
c50 15 0 1.30706e-19 $X=5.04 $Y=1.665
c51 12 0 1.73462e-19 $X=5.145 $Y=1.445
c52 9 0 1.73671e-19 $X=5.13 $Y=1.86
r53 22 23 2.05398 $w=3.52e-07 $l=1.5e-08 $layer=POLY_cond $X=5.13 $Y=1.652
+ $X2=5.145 $Y2=1.652
r54 20 22 10.2699 $w=3.52e-07 $l=7.5e-08 $layer=POLY_cond $X=5.055 $Y=1.652
+ $X2=5.13 $Y2=1.652
r55 18 20 56.142 $w=3.52e-07 $l=4.1e-07 $layer=POLY_cond $X=4.645 $Y=1.652
+ $X2=5.055 $Y2=1.652
r56 15 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.055
+ $Y=1.61 $X2=5.055 $Y2=1.61
r57 12 23 22.7654 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.145 $Y=1.445
+ $X2=5.145 $Y2=1.652
r58 12 14 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.145 $Y=1.445
+ $X2=5.145 $Y2=0.965
r59 9 22 22.7654 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=5.13 $Y=1.86
+ $X2=5.13 $Y2=1.652
r60 9 11 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.13 $Y=1.86
+ $X2=5.13 $Y2=2.435
r61 6 18 22.7654 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.645 $Y=1.445
+ $X2=4.645 $Y2=1.652
r62 6 8 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.645 $Y=1.445
+ $X2=4.645 $Y2=0.965
r63 3 5 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=4.625 $Y=2.02
+ $X2=4.625 $Y2=2.515
r64 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=4.625 $Y=1.93 $X2=4.625
+ $Y2=2.02
r65 1 18 2.73864 $w=3.52e-07 $l=2e-08 $layer=POLY_cond $X=4.625 $Y=1.652
+ $X2=4.645 $Y2=1.652
r66 1 2 60.25 $w=1.8e-07 $l=1.55e-07 $layer=POLY_cond $X=4.625 $Y=1.775
+ $X2=4.625 $Y2=1.93
.ends

.subckt PM_SKY130_FD_SC_LS__DLCLKP_2%A_27_74# 1 2 10 11 12 13 15 16 21 23 24 26
+ 29 32 38 40 43 44 45 46 48 49 50 56
c132 40 0 1.30966e-19 $X=1.05 $Y=0.855
c133 29 0 1.30706e-19 $X=5.562 $Y=1.56
c134 11 0 6.54874e-20 $X=2.885 $Y=2.215
r135 54 59 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=2.977 $Y=0.42
+ $X2=2.977 $Y2=0.585
r136 54 56 37.9425 $w=3.65e-07 $l=2.4e-07 $layer=POLY_cond $X=2.977 $Y=0.42
+ $X2=2.977 $Y2=0.18
r137 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.995
+ $Y=0.42 $X2=2.995 $Y2=0.42
r138 50 53 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=2.995 $Y=0.34
+ $X2=2.995 $Y2=0.42
r139 48 49 8.48848 $w=3.48e-07 $l=1.65e-07 $layer=LI1_cond $X=0.27 $Y=1.985
+ $X2=0.27 $Y2=1.82
r140 44 50 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.83 $Y=0.34
+ $X2=2.995 $Y2=0.34
r141 44 45 105.037 $w=1.68e-07 $l=1.61e-06 $layer=LI1_cond $X=2.83 $Y=0.34
+ $X2=1.22 $Y2=0.34
r142 42 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.135 $Y=0.425
+ $X2=1.22 $Y2=0.34
r143 42 43 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.135 $Y=0.425
+ $X2=1.135 $Y2=0.77
r144 41 46 2.28545 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.365 $Y=0.855
+ $X2=0.23 $Y2=0.855
r145 40 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.05 $Y=0.855
+ $X2=1.135 $Y2=0.77
r146 40 41 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=1.05 $Y=0.855
+ $X2=0.365 $Y2=0.855
r147 36 48 0.329269 $w=3.48e-07 $l=1e-08 $layer=LI1_cond $X=0.27 $Y=1.995
+ $X2=0.27 $Y2=1.985
r148 36 38 27.0001 $w=3.48e-07 $l=8.2e-07 $layer=LI1_cond $X=0.27 $Y=1.995
+ $X2=0.27 $Y2=2.815
r149 34 46 4.14756 $w=2.2e-07 $l=1.07121e-07 $layer=LI1_cond $X=0.18 $Y=0.94
+ $X2=0.23 $Y2=0.855
r150 34 49 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=0.18 $Y=0.94
+ $X2=0.18 $Y2=1.82
r151 30 46 4.14756 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=0.23 $Y=0.77
+ $X2=0.23 $Y2=0.855
r152 30 32 5.33538 $w=2.68e-07 $l=1.25e-07 $layer=LI1_cond $X=0.23 $Y=0.77
+ $X2=0.23 $Y2=0.645
r153 28 29 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=5.562 $Y=1.41
+ $X2=5.562 $Y2=1.56
r154 24 26 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.605 $Y=1.86
+ $X2=5.605 $Y2=2.435
r155 23 24 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.605 $Y=1.77
+ $X2=5.605 $Y2=1.86
r156 23 29 81.629 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=5.605 $Y=1.77
+ $X2=5.605 $Y2=1.56
r157 21 28 228.181 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=5.505 $Y=0.965
+ $X2=5.505 $Y2=1.41
r158 18 21 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=5.505 $Y=0.255
+ $X2=5.505 $Y2=0.965
r159 17 56 23.6381 $w=1.5e-07 $l=1.83e-07 $layer=POLY_cond $X=3.16 $Y=0.18
+ $X2=2.977 $Y2=0.18
r160 16 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.43 $Y=0.18
+ $X2=5.505 $Y2=0.255
r161 16 17 1163.98 $w=1.5e-07 $l=2.27e-06 $layer=POLY_cond $X=5.43 $Y=0.18
+ $X2=3.16 $Y2=0.18
r162 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.885 $Y=2.465
+ $X2=2.885 $Y2=2.75
r163 12 13 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.885 $Y=2.375
+ $X2=2.885 $Y2=2.465
r164 11 27 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.885 $Y=2.215
+ $X2=2.885 $Y2=2.125
r165 11 12 62.1936 $w=1.8e-07 $l=1.6e-07 $layer=POLY_cond $X=2.885 $Y=2.215
+ $X2=2.885 $Y2=2.375
r166 10 27 625.574 $w=1.5e-07 $l=1.22e-06 $layer=POLY_cond $X=2.87 $Y=0.905
+ $X2=2.87 $Y2=2.125
r167 10 59 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.87 $Y=0.905
+ $X2=2.87 $Y2=0.585
r168 2 48 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
r169 2 38 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r170 1 32 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_LS__DLCLKP_2%A_1041_387# 1 2 7 8 9 11 14 16 18 20 21 23
+ 29 35 38 39 44 45
c64 29 0 1.73671e-19 $X=5.38 $Y=2.81
r65 44 45 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.14
+ $Y=1.105 $X2=6.14 $Y2=1.105
r66 42 44 7.49781 $w=6.68e-07 $l=4.2e-07 $layer=LI1_cond $X=5.72 $Y=1.275
+ $X2=6.14 $Y2=1.275
r67 40 42 4.37372 $w=6.68e-07 $l=2.45e-07 $layer=LI1_cond $X=5.475 $Y=1.275
+ $X2=5.72 $Y2=1.275
r68 38 39 7.81132 $w=3.43e-07 $l=1.45e-07 $layer=LI1_cond $X=5.387 $Y=2.095
+ $X2=5.387 $Y2=1.95
r69 33 42 4.89075 $w=3.3e-07 $l=3.35e-07 $layer=LI1_cond $X=5.72 $Y=0.94
+ $X2=5.72 $Y2=1.275
r70 33 35 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=5.72 $Y=0.94 $X2=5.72
+ $Y2=0.74
r71 31 40 9.03384 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=5.475 $Y=1.61
+ $X2=5.475 $Y2=1.275
r72 31 39 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=5.475 $Y=1.61
+ $X2=5.475 $Y2=1.95
r73 27 38 0.901912 $w=3.43e-07 $l=2.7e-08 $layer=LI1_cond $X=5.387 $Y=2.122
+ $X2=5.387 $Y2=2.095
r74 27 29 22.9821 $w=3.43e-07 $l=6.88e-07 $layer=LI1_cond $X=5.387 $Y=2.122
+ $X2=5.387 $Y2=2.81
r75 24 45 46.3382 $w=3.3e-07 $l=2.65e-07 $layer=POLY_cond $X=6.14 $Y=1.37
+ $X2=6.14 $Y2=1.105
r76 21 23 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=7.185 $Y=1.31
+ $X2=7.185 $Y2=0.83
r77 18 20 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.175 $Y=1.765
+ $X2=7.175 $Y2=2.4
r78 16 18 76.5018 $w=1.76e-07 $l=2.75e-07 $layer=POLY_cond $X=7.175 $Y=1.49
+ $X2=7.175 $Y2=1.765
r79 16 21 50.4847 $w=1.76e-07 $l=1.84932e-07 $layer=POLY_cond $X=7.175 $Y=1.49
+ $X2=7.185 $Y2=1.31
r80 12 14 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=6.755 $Y=1.37
+ $X2=6.755 $Y2=0.83
r81 9 11 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.725 $Y=1.765
+ $X2=6.725 $Y2=2.4
r82 8 24 27.8133 $w=2.4e-07 $l=2.16852e-07 $layer=POLY_cond $X=6.305 $Y=1.49
+ $X2=6.14 $Y2=1.37
r83 7 9 72.3211 $w=1.89e-07 $l=2.78478e-07 $layer=POLY_cond $X=6.732 $Y=1.49
+ $X2=6.725 $Y2=1.765
r84 7 12 32.792 $w=1.89e-07 $l=1.30996e-07 $layer=POLY_cond $X=6.732 $Y=1.49
+ $X2=6.755 $Y2=1.37
r85 7 16 65.9955 $w=2.4e-07 $l=2.55e-07 $layer=POLY_cond $X=6.83 $Y=1.49
+ $X2=7.085 $Y2=1.49
r86 7 8 85.4059 $w=2.4e-07 $l=3.3e-07 $layer=POLY_cond $X=6.635 $Y=1.49
+ $X2=6.305 $Y2=1.49
r87 2 38 400 $w=1.7e-07 $l=2.42126e-07 $layer=licon1_PDIFF $count=1 $X=5.205
+ $Y=1.935 $X2=5.38 $Y2=2.095
r88 2 29 400 $w=1.7e-07 $l=9.58514e-07 $layer=licon1_PDIFF $count=1 $X=5.205
+ $Y=1.935 $X2=5.38 $Y2=2.81
r89 1 35 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.58
+ $Y=0.595 $X2=5.72 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__DLCLKP_2%VPWR 1 2 3 4 5 20 24 28 32 36 38 43 44 45
+ 47 62 66 72 75 78 82
r82 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r83 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r84 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r85 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r86 70 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.44 $Y2=3.33
r87 70 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6.48 $Y2=3.33
r88 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r89 67 78 15.5458 $w=1.7e-07 $l=4.53e-07 $layer=LI1_cond $X=6.635 $Y=3.33
+ $X2=6.182 $Y2=3.33
r90 67 69 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=6.635 $Y=3.33
+ $X2=6.96 $Y2=3.33
r91 66 81 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=7.315 $Y=3.33
+ $X2=7.497 $Y2=3.33
r92 66 69 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=7.315 $Y=3.33
+ $X2=6.96 $Y2=3.33
r93 65 79 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6.48 $Y2=3.33
r94 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r95 62 78 15.5458 $w=1.7e-07 $l=4.52e-07 $layer=LI1_cond $X=5.73 $Y=3.33
+ $X2=6.182 $Y2=3.33
r96 62 64 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=5.73 $Y=3.33
+ $X2=5.52 $Y2=3.33
r97 61 65 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r98 60 61 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r99 58 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r100 57 60 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.6 $Y=3.33 $X2=4.56
+ $Y2=3.33
r101 57 58 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r102 55 75 11.8214 $w=1.7e-07 $l=2.7e-07 $layer=LI1_cond $X=3.485 $Y=3.33
+ $X2=3.215 $Y2=3.33
r103 55 57 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=3.485 $Y=3.33
+ $X2=3.6 $Y2=3.33
r104 54 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r105 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r106 51 54 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r107 51 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r108 50 53 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r109 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r110 48 72 9.6488 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=1.075 $Y=3.33
+ $X2=0.88 $Y2=3.33
r111 48 50 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=1.075 $Y=3.33
+ $X2=1.2 $Y2=3.33
r112 47 75 11.8214 $w=1.7e-07 $l=2.7e-07 $layer=LI1_cond $X=2.945 $Y=3.33
+ $X2=3.215 $Y2=3.33
r113 47 53 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.945 $Y=3.33
+ $X2=2.64 $Y2=3.33
r114 45 61 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=4.56 $Y2=3.33
r115 45 58 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=3.6 $Y2=3.33
r116 43 60 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=4.715 $Y=3.33
+ $X2=4.56 $Y2=3.33
r117 43 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.715 $Y=3.33
+ $X2=4.88 $Y2=3.33
r118 42 64 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=5.045 $Y=3.33
+ $X2=5.52 $Y2=3.33
r119 42 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.045 $Y=3.33
+ $X2=4.88 $Y2=3.33
r120 38 41 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=7.44 $Y=1.985
+ $X2=7.44 $Y2=2.815
r121 36 81 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=7.44 $Y=3.245
+ $X2=7.497 $Y2=3.33
r122 36 41 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=7.44 $Y=3.245
+ $X2=7.44 $Y2=2.815
r123 32 35 9.36906 $w=9.03e-07 $l=6.95e-07 $layer=LI1_cond $X=6.182 $Y=2.115
+ $X2=6.182 $Y2=2.81
r124 30 78 3.35974 $w=9.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.182 $Y=3.245
+ $X2=6.182 $Y2=3.33
r125 30 35 5.86409 $w=9.03e-07 $l=4.35e-07 $layer=LI1_cond $X=6.182 $Y=3.245
+ $X2=6.182 $Y2=2.81
r126 26 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.88 $Y=3.245
+ $X2=4.88 $Y2=3.33
r127 26 28 35.0971 $w=3.28e-07 $l=1.005e-06 $layer=LI1_cond $X=4.88 $Y=3.245
+ $X2=4.88 $Y2=2.24
r128 22 75 2.26835 $w=5.4e-07 $l=8.5e-08 $layer=LI1_cond $X=3.215 $Y=3.245
+ $X2=3.215 $Y2=3.33
r129 22 24 9.52433 $w=5.38e-07 $l=4.3e-07 $layer=LI1_cond $X=3.215 $Y=3.245
+ $X2=3.215 $Y2=2.815
r130 18 72 1.39532 $w=3.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.88 $Y=3.245
+ $X2=0.88 $Y2=3.33
r131 18 20 25.4128 $w=3.88e-07 $l=8.6e-07 $layer=LI1_cond $X=0.88 $Y=3.245
+ $X2=0.88 $Y2=2.385
r132 5 41 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=7.25
+ $Y=1.84 $X2=7.4 $Y2=2.815
r133 5 38 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=7.25
+ $Y=1.84 $X2=7.4 $Y2=1.985
r134 4 35 200 $w=1.7e-07 $l=9.49342e-07 $layer=licon1_PDIFF $count=3 $X=5.68
+ $Y=1.935 $X2=5.835 $Y2=2.81
r135 4 32 200 $w=1.7e-07 $l=2.45561e-07 $layer=licon1_PDIFF $count=3 $X=5.68
+ $Y=1.935 $X2=5.835 $Y2=2.115
r136 3 28 300 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_PDIFF $count=2 $X=4.7
+ $Y=2.095 $X2=4.88 $Y2=2.24
r137 2 24 600 $w=1.7e-07 $l=3.81772e-07 $layer=licon1_PDIFF $count=1 $X=2.96
+ $Y=2.54 $X2=3.215 $Y2=2.815
r138 1 20 300 $w=1.7e-07 $l=6.7862e-07 $layer=licon1_PDIFF $count=2 $X=0.58
+ $Y=1.84 $X2=0.88 $Y2=2.385
.ends

.subckt PM_SKY130_FD_SC_LS__DLCLKP_2%GCLK 1 2 7 8 9 10 11 12 13
r17 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=6.97 $Y=2.405
+ $X2=6.97 $Y2=2.775
r18 11 12 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=6.97 $Y=1.985
+ $X2=6.97 $Y2=2.405
r19 10 11 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=6.97 $Y=1.665
+ $X2=6.97 $Y2=1.985
r20 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=6.97 $Y=1.295
+ $X2=6.97 $Y2=1.665
r21 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=6.97 $Y=0.925 $X2=6.97
+ $Y2=1.295
r22 7 8 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=6.97 $Y=0.555 $X2=6.97
+ $Y2=0.925
r23 2 13 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=6.8
+ $Y=1.84 $X2=6.95 $Y2=2.815
r24 2 11 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=6.8
+ $Y=1.84 $X2=6.95 $Y2=1.985
r25 1 7 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.83
+ $Y=0.46 $X2=6.97 $Y2=0.605
.ends

.subckt PM_SKY130_FD_SC_LS__DLCLKP_2%VGND 1 2 3 4 5 18 20 25 28 32 34 36 39 40
+ 43 45 57 64 69 75 78 81 85
r92 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r93 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r94 78 79 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r95 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r96 73 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r97 73 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=6.48
+ $Y2=0
r98 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r99 70 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.635 $Y=0 $X2=6.47
+ $Y2=0
r100 70 72 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=6.635 $Y=0
+ $X2=6.96 $Y2=0
r101 69 84 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=7.315 $Y=0
+ $X2=7.497 $Y2=0
r102 69 72 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=7.315 $Y=0
+ $X2=6.96 $Y2=0
r103 68 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r104 68 79 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.04
+ $Y2=0
r105 67 68 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r106 65 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.095 $Y=0 $X2=4.93
+ $Y2=0
r107 65 67 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=5.095 $Y=0 $X2=6
+ $Y2=0
r108 64 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.305 $Y=0 $X2=6.47
+ $Y2=0
r109 64 67 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=6.305 $Y=0 $X2=6
+ $Y2=0
r110 63 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r111 62 63 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r112 59 62 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r113 59 60 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r114 57 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.765 $Y=0 $X2=4.93
+ $Y2=0
r115 57 62 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=4.765 $Y=0
+ $X2=4.56 $Y2=0
r116 56 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r117 55 56 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r118 53 56 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r119 53 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r120 52 55 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r121 52 53 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r122 50 75 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=0.88 $Y=0 $X2=0.712
+ $Y2=0
r123 50 52 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.88 $Y=0 $X2=1.2
+ $Y2=0
r124 48 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r125 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r126 45 75 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=0.545 $Y=0
+ $X2=0.712 $Y2=0
r127 45 47 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0
+ $X2=0.24 $Y2=0
r128 43 63 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.84 $Y=0 $X2=4.56
+ $Y2=0
r129 43 60 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=0 $X2=3.6
+ $Y2=0
r130 39 55 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=3.34 $Y=0 $X2=3.12
+ $Y2=0
r131 39 40 5.78184 $w=1.7e-07 $l=9.7e-08 $layer=LI1_cond $X=3.34 $Y=0 $X2=3.437
+ $Y2=0
r132 38 59 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=3.535 $Y=0 $X2=3.6
+ $Y2=0
r133 38 40 5.78184 $w=1.7e-07 $l=9.8e-08 $layer=LI1_cond $X=3.535 $Y=0 $X2=3.437
+ $Y2=0
r134 34 84 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=7.44 $Y=0.085
+ $X2=7.497 $Y2=0
r135 34 36 23.9708 $w=2.48e-07 $l=5.2e-07 $layer=LI1_cond $X=7.44 $Y=0.085
+ $X2=7.44 $Y2=0.605
r136 30 81 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.47 $Y=0.085
+ $X2=6.47 $Y2=0
r137 30 32 18.1597 $w=3.28e-07 $l=5.2e-07 $layer=LI1_cond $X=6.47 $Y=0.085
+ $X2=6.47 $Y2=0.605
r138 26 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.93 $Y=0.085
+ $X2=4.93 $Y2=0
r139 26 28 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=4.93 $Y=0.085
+ $X2=4.93 $Y2=0.74
r140 25 42 3.91487 $w=1.95e-07 $l=1.25e-07 $layer=LI1_cond $X=3.437 $Y=0.755
+ $X2=3.437 $Y2=0.88
r141 24 40 0.85348 $w=1.95e-07 $l=8.5e-08 $layer=LI1_cond $X=3.437 $Y=0.085
+ $X2=3.437 $Y2=0
r142 24 25 38.1072 $w=1.93e-07 $l=6.7e-07 $layer=LI1_cond $X=3.437 $Y=0.085
+ $X2=3.437 $Y2=0.755
r143 20 42 3.03794 $w=2.5e-07 $l=9.7e-08 $layer=LI1_cond $X=3.34 $Y=0.88
+ $X2=3.437 $Y2=0.88
r144 20 22 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=3.34 $Y=0.88
+ $X2=3.085 $Y2=0.88
r145 16 75 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=0.712 $Y=0.085
+ $X2=0.712 $Y2=0
r146 16 18 14.7926 $w=3.33e-07 $l=4.3e-07 $layer=LI1_cond $X=0.712 $Y=0.085
+ $X2=0.712 $Y2=0.515
r147 5 36 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.26
+ $Y=0.46 $X2=7.4 $Y2=0.605
r148 4 32 182 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=1 $X=6.315
+ $Y=0.46 $X2=6.47 $Y2=0.605
r149 3 28 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=4.72
+ $Y=0.595 $X2=4.93 $Y2=0.74
r150 2 42 182 $w=1.7e-07 $l=5.6285e-07 $layer=licon1_NDIFF $count=1 $X=2.945
+ $Y=0.695 $X2=3.44 $Y2=0.84
r151 2 22 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.945
+ $Y=0.695 $X2=3.085 $Y2=0.84
r152 1 18 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.515
.ends

