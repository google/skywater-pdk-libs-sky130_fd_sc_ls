* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
X0 VPWR a_83_256# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X1 VGND a_83_256# X VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X2 a_564_74# A3 VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X3 a_1234_392# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 VGND A2 a_564_74# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X5 a_564_74# B2 a_83_256# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X6 a_534_388# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 a_83_256# A3 a_961_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 a_564_74# B1 a_83_256# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X9 a_534_388# B2 a_83_256# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_1234_392# A2 a_961_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 X a_83_256# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X12 a_564_74# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X13 X a_83_256# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X14 VPWR a_83_256# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X15 a_83_256# B1 a_564_74# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X16 X a_83_256# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X17 VGND A3 a_564_74# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X18 VPWR B1 a_534_388# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 a_961_392# A3 a_83_256# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X20 a_564_74# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X21 a_961_392# A2 a_1234_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X22 a_83_256# B2 a_534_388# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X23 VGND a_83_256# X VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X24 VPWR A1 a_1234_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X25 X a_83_256# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X26 a_83_256# B2 a_564_74# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X27 VGND A1 a_564_74# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
.ends
