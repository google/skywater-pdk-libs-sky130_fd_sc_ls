* File: sky130_fd_sc_ls__sedfxtp_4.spice
* Created: Fri Aug 28 14:07:44 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__sedfxtp_4.pex.spice"
.subckt sky130_fd_sc_ls__sedfxtp_4  VNB VPB D DE SCD SCE CLK VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* CLK	CLK
* SCE	SCE
* SCD	SCD
* DE	DE
* D	D
* VPB	VPB
* VNB	VNB
MM1000 A_135_74# N_D_M1000_g N_A_37_464#_M1000_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1029 N_VGND_M1029_d N_DE_M1029_g A_135_74# VNB NSHORT L=0.15 W=0.42 AD=0.1197
+ AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.6 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_DE_M1004_g N_A_177_290#_M1004_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75001.7
+ A=0.063 P=1.14 MULT=1
MM1035 A_497_113# N_A_177_290#_M1035_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0588 PD=0.66 PS=0.7 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1020 N_A_37_464#_M1020_d N_A_545_87#_M1020_g A_497_113# VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.0504 PD=0.7 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001
+ SB=75000.9 A=0.063 P=1.14 MULT=1
MM1021 N_A_661_113#_M1021_d N_A_631_87#_M1021_g N_A_37_464#_M1020_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.21 AS=0.0588 PD=1.84 PS=0.7 NRD=39.996 NRS=0 M=1 R=2.8
+ SA=75001.5 SB=75000.4 A=0.063 P=1.14 MULT=1
MM1042 N_VGND_M1042_d N_SCE_M1042_g N_A_631_87#_M1042_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75001
+ A=0.063 P=1.14 MULT=1
MM1007 A_1044_125# N_SCD_M1007_g N_VGND_M1042_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1001 N_A_661_113#_M1001_d N_SCE_M1001_g A_1044_125# VNB NSHORT L=0.15 W=0.42
+ AD=0.1176 AS=0.0441 PD=1.4 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1022 N_A_1313_74#_M1022_d N_CLK_M1022_g N_VGND_M1022_s VNB NSHORT L=0.15
+ W=0.74 AD=0.2072 AS=0.2109 PD=2.04 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1011 N_A_1510_74#_M1011_d N_A_1313_74#_M1011_g N_VGND_M1011_s VNB NSHORT
+ L=0.15 W=0.74 AD=0.2072 AS=0.2109 PD=2.04 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1037 N_A_1756_97#_M1037_d N_A_1313_74#_M1037_g N_A_661_113#_M1037_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.083475 AS=0.2226 PD=0.87 PS=1.9 NRD=0 NRS=71.424 M=1 R=2.8
+ SA=75000.5 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1032 A_1858_79# N_A_1510_74#_M1032_g N_A_1756_97#_M1037_d VNB NSHORT L=0.15
+ W=0.42 AD=0.08925 AS=0.083475 PD=0.845 PS=0.87 NRD=45 NRS=24.276 M=1 R=2.8
+ SA=75000.8 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1027 N_VGND_M1027_d N_A_1943_53#_M1027_g A_1858_79# VNB NSHORT L=0.15 W=0.42
+ AD=0.109992 AS=0.08925 PD=0.92717 PS=0.845 NRD=0 NRS=45 M=1 R=2.8 SA=75001.4
+ SB=75000.9 A=0.063 P=1.14 MULT=1
MM1046 N_A_1943_53#_M1046_d N_A_1756_97#_M1046_g N_VGND_M1027_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.1824 AS=0.167608 PD=1.85 PS=1.41283 NRD=0 NRS=46.872 M=1
+ R=4.26667 SA=75001.4 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1047 A_2331_74# N_A_1943_53#_M1047_g N_VGND_M1047_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0672 AS=0.1824 PD=0.85 PS=1.85 NRD=9.372 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75001.9 A=0.096 P=1.58 MULT=1
MM1026 N_A_2403_74#_M1026_d N_A_1510_74#_M1026_g A_2331_74# VNB NSHORT L=0.15
+ W=0.64 AD=0.115623 AS=0.0672 PD=1.16528 PS=0.85 NRD=8.436 NRS=9.372 M=1
+ R=4.26667 SA=75000.6 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1013 A_2498_74# N_A_1313_74#_M1013_g N_A_2403_74#_M1026_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.0758774 PD=0.66 PS=0.764717 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75001 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1014 N_VGND_M1014_d N_A_545_87#_M1014_g A_2498_74# VNB NSHORT L=0.15 W=0.42
+ AD=0.21 AS=0.0504 PD=1.42 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.4
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1016 N_A_545_87#_M1016_d N_A_2403_74#_M1016_g N_VGND_M1014_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1197 AS=0.21 PD=1.41 PS=1.42 NRD=0 NRS=19.992 M=1 R=2.8 SA=75002.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1019 N_Q_M1019_d N_A_2403_74#_M1019_g N_VGND_M1019_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1036 N_Q_M1019_d N_A_2403_74#_M1036_g N_VGND_M1036_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75000.6
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1039 N_Q_M1039_d N_A_2403_74#_M1039_g N_VGND_M1036_s VNB NSHORT L=0.15 W=0.74
+ AD=0.10915 AS=0.1295 PD=1.035 PS=1.09 NRD=0.804 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1040 N_Q_M1039_d N_A_2403_74#_M1040_g N_VGND_M1040_s VNB NSHORT L=0.15 W=0.74
+ AD=0.10915 AS=0.1998 PD=1.035 PS=2.02 NRD=1.62 NRS=0 M=1 R=4.93333 SA=75001.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1023 A_126_464# N_D_M1023_g N_A_37_464#_M1023_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0864 AS=0.1888 PD=0.91 PS=1.87 NRD=24.625 NRS=3.0732 M=1 R=4.26667
+ SA=75000.2 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1005 N_VPWR_M1005_d N_A_177_290#_M1005_g A_126_464# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1888 AS=0.0864 PD=1.87 PS=0.91 NRD=3.0732 NRS=24.625 M=1 R=4.26667
+ SA=75000.6 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1010 N_VPWR_M1010_d N_DE_M1010_g N_A_177_290#_M1010_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1696 AS=0.1888 PD=1.17 PS=1.87 NRD=73.8553 NRS=3.0732 M=1
+ R=4.26667 SA=75000.2 SB=75001.7 A=0.096 P=1.58 MULT=1
MM1028 A_572_463# N_DE_M1028_g N_VPWR_M1010_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0768 AS=0.1696 PD=0.88 PS=1.17 NRD=19.9955 NRS=3.0732 M=1 R=4.26667
+ SA=75000.9 SB=75001 A=0.096 P=1.58 MULT=1
MM1006 N_A_37_464#_M1006_d N_A_545_87#_M1006_g A_572_463# VPB PHIGHVT L=0.15
+ W=0.64 AD=0.096 AS=0.0768 PD=0.94 PS=0.88 NRD=3.0732 NRS=19.9955 M=1 R=4.26667
+ SA=75001.3 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1015 N_A_661_113#_M1015_d N_SCE_M1015_g N_A_37_464#_M1006_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.176 AS=0.096 PD=1.83 PS=0.94 NRD=3.0732 NRS=3.0732 M=1 R=4.26667
+ SA=75001.7 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1044 N_VPWR_M1044_d N_SCE_M1044_g N_A_631_87#_M1044_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1696 AS=0.1792 PD=1.17 PS=1.84 NRD=73.8553 NRS=3.0732 M=1
+ R=4.26667 SA=75000.2 SB=75001.3 A=0.096 P=1.58 MULT=1
MM1012 A_1071_455# N_SCD_M1012_g N_VPWR_M1044_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0768 AS=0.1696 PD=0.88 PS=1.17 NRD=19.9955 NRS=3.0732 M=1 R=4.26667
+ SA=75000.9 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1034 N_A_661_113#_M1034_d N_A_631_87#_M1034_g A_1071_455# VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1792 AS=0.0768 PD=1.84 PS=0.88 NRD=3.0732 NRS=19.9955 M=1
+ R=4.26667 SA=75001.3 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1041 N_A_1313_74#_M1041_d N_CLK_M1041_g N_VPWR_M1041_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.308 AS=0.3136 PD=2.79 PS=2.8 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1017 N_A_1510_74#_M1017_d N_A_1313_74#_M1017_g N_VPWR_M1017_s VPB PHIGHVT
+ L=0.15 W=1.12 AD=0.308 AS=0.308 PD=2.79 PS=2.79 NRD=1.7533 NRS=1.7533 M=1
+ R=7.46667 SA=75000.2 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1018 N_A_1756_97#_M1018_d N_A_1510_74#_M1018_g N_A_661_113#_M1018_s VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.063 AS=0.1155 PD=0.72 PS=1.39 NRD=4.6886 NRS=4.6886
+ M=1 R=2.8 SA=75000.2 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1025 A_1899_508# N_A_1313_74#_M1025_g N_A_1756_97#_M1018_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0693 AS=0.063 PD=0.75 PS=0.72 NRD=51.5943 NRS=4.6886 M=1 R=2.8
+ SA=75000.6 SB=75001 A=0.063 P=1.14 MULT=1
MM1009 N_VPWR_M1009_d N_A_1943_53#_M1009_g A_1899_508# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0957833 AS=0.0693 PD=0.89 PS=0.75 NRD=4.6886 NRS=51.5943 M=1 R=2.8
+ SA=75001.1 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1002 N_A_1943_53#_M1002_d N_A_1756_97#_M1002_g N_VPWR_M1009_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.231 AS=0.191567 PD=2.23 PS=1.78 NRD=2.3443 NRS=18.7544 M=1
+ R=5.6 SA=75000.7 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1043 A_2292_392# N_A_1943_53#_M1043_g N_VPWR_M1043_s VPB PHIGHVT L=0.15 W=1
+ AD=0.405 AS=0.275 PD=1.81 PS=2.55 NRD=68.9303 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75001.8 A=0.15 P=2.3 MULT=1
MM1008 N_A_2403_74#_M1008_d N_A_1313_74#_M1008_g A_2292_392# VPB PHIGHVT L=0.15
+ W=1 AD=0.214718 AS=0.405 PD=1.91549 PS=1.81 NRD=13.7703 NRS=68.9303 M=1
+ R=6.66667 SA=75001.2 SB=75000.9 A=0.15 P=2.3 MULT=1
MM1045 A_2586_508# N_A_1510_74#_M1045_g N_A_2403_74#_M1008_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0567 AS=0.0901817 PD=0.69 PS=0.804507 NRD=37.5088 NRS=4.6886 M=1
+ R=2.8 SA=75001.7 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1030 N_VPWR_M1030_d N_A_545_87#_M1030_g A_2586_508# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.116292 AS=0.0567 PD=0.950943 PS=0.69 NRD=53.9386 NRS=37.5088 M=1 R=2.8
+ SA=75002.1 SB=75000.9 A=0.063 P=1.14 MULT=1
MM1031 N_A_545_87#_M1031_d N_A_2403_74#_M1031_g N_VPWR_M1030_d VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.176 AS=0.177208 PD=1.83 PS=1.44906 NRD=3.0732 NRS=50.7866
+ M=1 R=4.26667 SA=75001.9 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1003 N_VPWR_M1003_d N_A_2403_74#_M1003_g N_Q_M1003_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.308 AS=0.168 PD=2.79 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1024 N_VPWR_M1024_d N_A_2403_74#_M1024_g N_Q_M1003_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.6 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1033 N_VPWR_M1024_d N_A_2403_74#_M1033_g N_Q_M1033_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1038 N_VPWR_M1038_d N_A_2403_74#_M1038_g N_Q_M1033_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3192 AS=0.168 PD=2.81 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.5 SB=75000.2 A=0.168 P=2.54 MULT=1
DX48_noxref VNB VPB NWDIODE A=31.9921 P=38.15
c_177 VNB 0 1.36415e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_ls__sedfxtp_4.pxi.spice"
*
.ends
*
*
