* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__mux2i_4 A0 A1 S VGND VNB VPB VPWR Y
M1000 Y A1 a_116_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=1.792e+12p pd=1.44e+07u as=1.4336e+12p ps=1.152e+07u
M1001 a_478_368# A0 Y VPB phighvt w=1.12e+06u l=150000u
+  ad=1.4448e+12p pd=1.154e+07u as=0p ps=0u
M1002 a_116_368# a_1030_268# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=2.5466e+12p ps=1.762e+07u
M1003 VPWR S a_478_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_475_85# A0 Y VNB nshort w=740000u l=150000u
+  ad=8.806e+11p pd=8.3e+06u as=1.0767e+12p ps=1.031e+07u
M1005 a_114_85# S VGND VNB nshort w=740000u l=150000u
+  ad=8.917e+11p pd=8.33e+06u as=1.795e+12p ps=1.331e+07u
M1006 a_475_85# a_1030_268# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND a_1030_268# a_475_85# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_478_368# S VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_114_85# S VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 Y A0 a_478_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_114_85# A1 Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Y A1 a_114_85# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_1030_268# S VGND VNB nshort w=740000u l=150000u
+  ad=2.627e+11p pd=2.19e+06u as=0p ps=0u
M1014 a_116_368# A1 Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y A1 a_116_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR S a_478_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_1030_268# S VPWR VPB phighvt w=840000u l=150000u
+  ad=2.52e+11p pd=2.28e+06u as=0p ps=0u
M1018 a_116_368# a_1030_268# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND S a_114_85# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_478_368# A0 Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND a_1030_268# a_475_85# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND S a_114_85# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VPWR a_1030_268# a_116_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_475_85# a_1030_268# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_116_368# A1 Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VPWR S a_1030_268# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 Y A0 a_475_85# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 Y A0 a_475_85# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 Y A0 a_478_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VPWR a_1030_268# a_116_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_475_85# A0 Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 Y A1 a_114_85# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_478_368# S VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_114_85# A1 Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
