# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_ls__dlrtn_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_ls__dlrtn_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.200000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.208500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.435000 1.450000 0.835000 1.780000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.600500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.730000 0.350000 7.115000 1.130000 ;
        RECT 6.755000 1.820000 7.115000 2.980000 ;
        RECT 6.945000 1.130000 7.115000 1.820000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.885000 1.180000 6.235000 1.550000 ;
    END
  END RESET_B
  PIN VNB
    PORT
      LAYER pwell ;
        RECT 0.000000 0.000000 7.200000 0.245000 ;
    END
  END VNB
  PIN VPB
    PORT
      LAYER nwell ;
        RECT -0.190000 1.660000 7.390000 3.520000 ;
    END
  END VPB
  PIN GATE_N
    ANTENNAGATEAREA  0.237000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.005000 1.450000 1.335000 1.780000 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.200000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 7.200000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.200000 0.085000 ;
      RECT 0.000000  3.245000 7.200000 3.415000 ;
      RECT 0.095000  0.580000 2.865000 0.750000 ;
      RECT 0.095000  0.750000 0.445000 1.250000 ;
      RECT 0.095000  1.250000 0.265000 1.950000 ;
      RECT 0.095000  1.950000 0.450000 2.830000 ;
      RECT 0.625000  0.085000 0.955000 0.410000 ;
      RECT 0.655000  1.950000 0.985000 3.245000 ;
      RECT 1.065000  0.920000 1.675000 1.250000 ;
      RECT 1.190000  1.950000 1.675000 2.520000 ;
      RECT 1.190000  2.520000 4.245000 2.690000 ;
      RECT 1.190000  2.690000 1.675000 2.830000 ;
      RECT 1.505000  1.250000 1.675000 1.340000 ;
      RECT 1.505000  1.340000 1.905000 1.670000 ;
      RECT 1.505000  1.670000 1.675000 1.950000 ;
      RECT 1.845000  0.920000 2.245000 1.170000 ;
      RECT 1.845000  1.840000 3.405000 2.010000 ;
      RECT 1.845000  2.010000 2.245000 2.350000 ;
      RECT 2.075000  1.170000 2.245000 1.840000 ;
      RECT 2.300000  2.860000 2.630000 3.245000 ;
      RECT 2.355000  0.085000 3.200000 0.410000 ;
      RECT 2.535000  0.750000 2.865000 1.590000 ;
      RECT 3.075000  1.190000 4.335000 1.520000 ;
      RECT 3.075000  1.520000 3.405000 1.840000 ;
      RECT 3.255000  2.180000 3.745000 2.350000 ;
      RECT 3.575000  1.690000 5.070000 1.860000 ;
      RECT 3.575000  1.860000 3.745000 2.180000 ;
      RECT 3.815000  0.350000 4.145000 0.850000 ;
      RECT 3.815000  0.850000 5.070000 1.020000 ;
      RECT 3.915000  2.030000 4.245000 2.520000 ;
      RECT 4.485000  2.030000 5.965000 2.360000 ;
      RECT 4.635000  2.530000 5.430000 3.245000 ;
      RECT 4.670000  0.085000 5.010000 0.680000 ;
      RECT 4.900000  1.020000 5.070000 1.300000 ;
      RECT 4.900000  1.300000 5.295000 1.630000 ;
      RECT 4.900000  1.630000 5.070000 1.690000 ;
      RECT 5.240000  0.350000 5.635000 1.130000 ;
      RECT 5.465000  1.130000 5.635000 1.720000 ;
      RECT 5.465000  1.720000 6.585000 1.890000 ;
      RECT 5.465000  1.890000 5.965000 2.030000 ;
      RECT 5.635000  2.360000 5.965000 2.860000 ;
      RECT 6.140000  0.085000 6.470000 1.010000 ;
      RECT 6.255000  2.060000 6.585000 3.245000 ;
      RECT 6.415000  1.320000 6.775000 1.650000 ;
      RECT 6.415000  1.650000 6.585000 1.720000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
  END
END sky130_fd_sc_ls__dlrtn_1
END LIBRARY
