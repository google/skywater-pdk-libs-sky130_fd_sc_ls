* File: sky130_fd_sc_ls__bufbuf_16.pex.spice
* Created: Fri Aug 28 13:07:31 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__BUFBUF_16%A 1 3 6 8 12
c32 1 0 5.40859e-20 $X=0.505 $Y=1.765
r33 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.34
+ $Y=1.465 $X2=0.34 $Y2=1.465
r34 8 12 6.06549 $w=3.78e-07 $l=2e-07 $layer=LI1_cond $X=0.315 $Y=1.665
+ $X2=0.315 $Y2=1.465
r35 4 11 38.7839 $w=3.5e-07 $l=2.18746e-07 $layer=POLY_cond $X=0.51 $Y=1.3
+ $X2=0.385 $Y2=1.465
r36 4 6 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.51 $Y=1.3 $X2=0.51
+ $Y2=0.74
r37 1 11 57.3754 $w=3.5e-07 $l=3.54965e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.385 $Y2=1.465
r38 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__BUFBUF_16%A_27_368# 1 2 9 11 13 16 18 20 23 25 27 28
+ 30 34 36 37 38 41 43 49 54 61
c110 9 0 1.78628e-19 $X=0.94 $Y=0.74
r111 61 62 6.07053 $w=3.97e-07 $l=5e-08 $layer=POLY_cond $X=1.805 $Y=1.532
+ $X2=1.855 $Y2=1.532
r112 58 59 4.24937 $w=3.97e-07 $l=3.5e-08 $layer=POLY_cond $X=1.37 $Y=1.532
+ $X2=1.405 $Y2=1.532
r113 55 56 1.82116 $w=3.97e-07 $l=1.5e-08 $layer=POLY_cond $X=0.94 $Y=1.532
+ $X2=0.955 $Y2=1.532
r114 50 61 11.534 $w=3.97e-07 $l=9.5e-08 $layer=POLY_cond $X=1.71 $Y=1.532
+ $X2=1.805 $Y2=1.532
r115 50 59 37.0302 $w=3.97e-07 $l=3.05e-07 $layer=POLY_cond $X=1.71 $Y=1.532
+ $X2=1.405 $Y2=1.532
r116 49 50 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.71
+ $Y=1.465 $X2=1.71 $Y2=1.465
r117 47 58 41.2796 $w=3.97e-07 $l=3.4e-07 $layer=POLY_cond $X=1.03 $Y=1.532
+ $X2=1.37 $Y2=1.532
r118 47 56 9.10579 $w=3.97e-07 $l=7.5e-08 $layer=POLY_cond $X=1.03 $Y=1.532
+ $X2=0.955 $Y2=1.532
r119 46 49 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.03 $Y=1.465
+ $X2=1.71 $Y2=1.465
r120 46 47 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.03
+ $Y=1.465 $X2=1.03 $Y2=1.465
r121 44 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.845 $Y=1.465
+ $X2=0.76 $Y2=1.465
r122 44 46 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=0.845 $Y=1.465
+ $X2=1.03 $Y2=1.465
r123 42 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.76 $Y=1.63
+ $X2=0.76 $Y2=1.465
r124 42 43 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.76 $Y=1.63
+ $X2=0.76 $Y2=1.95
r125 41 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.76 $Y=1.3
+ $X2=0.76 $Y2=1.465
r126 40 41 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.76 $Y=1.13
+ $X2=0.76 $Y2=1.3
r127 39 53 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.445 $Y=2.035
+ $X2=0.28 $Y2=2.035
r128 38 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.675 $Y=2.035
+ $X2=0.76 $Y2=1.95
r129 38 39 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=0.675 $Y=2.035
+ $X2=0.445 $Y2=2.035
r130 36 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.675 $Y=1.045
+ $X2=0.76 $Y2=1.13
r131 36 37 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.675 $Y=1.045
+ $X2=0.38 $Y2=1.045
r132 32 37 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.255 $Y=0.96
+ $X2=0.38 $Y2=1.045
r133 32 34 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=0.255 $Y=0.96
+ $X2=0.255 $Y2=0.515
r134 28 53 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.28 $Y=2.12 $X2=0.28
+ $Y2=2.035
r135 28 30 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=0.28 $Y=2.12
+ $X2=0.28 $Y2=2.815
r136 25 62 25.678 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=1.855 $Y=1.765
+ $X2=1.855 $Y2=1.532
r137 25 27 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.855 $Y=1.765
+ $X2=1.855 $Y2=2.4
r138 21 61 25.678 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=1.805 $Y=1.3
+ $X2=1.805 $Y2=1.532
r139 21 23 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.805 $Y=1.3
+ $X2=1.805 $Y2=0.74
r140 18 59 25.678 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=1.405 $Y=1.765
+ $X2=1.405 $Y2=1.532
r141 18 20 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.405 $Y=1.765
+ $X2=1.405 $Y2=2.4
r142 14 58 25.678 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=1.37 $Y=1.3
+ $X2=1.37 $Y2=1.532
r143 14 16 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.37 $Y=1.3
+ $X2=1.37 $Y2=0.74
r144 11 56 25.678 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=0.955 $Y=1.765
+ $X2=0.955 $Y2=1.532
r145 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.955 $Y=1.765
+ $X2=0.955 $Y2=2.4
r146 7 55 25.678 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=0.94 $Y=1.3 $X2=0.94
+ $Y2=1.532
r147 7 9 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.94 $Y=1.3 $X2=0.94
+ $Y2=0.74
r148 2 53 400 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.115
r149 2 30 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r150 1 34 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.15
+ $Y=0.37 $X2=0.295 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__BUFBUF_16%A_203_74# 1 2 3 4 15 17 19 22 24 26 27 29
+ 32 36 38 40 41 43 46 48 50 53 57 63 65 66 67 68 71 75 80 82 88 91 92 93 106
c194 68 0 5.40859e-20 $X=1.345 $Y=1.885
c195 66 0 1.78628e-19 $X=1.24 $Y=1.045
c196 48 0 3.06714e-20 $X=5.14 $Y=1.765
r197 106 107 1.90263 $w=3.8e-07 $l=1.5e-08 $layer=POLY_cond $X=5.14 $Y=1.542
+ $X2=5.155 $Y2=1.542
r198 105 106 52.6395 $w=3.8e-07 $l=4.15e-07 $layer=POLY_cond $X=4.725 $Y=1.542
+ $X2=5.14 $Y2=1.542
r199 104 105 4.43947 $w=3.8e-07 $l=3.5e-08 $layer=POLY_cond $X=4.69 $Y=1.542
+ $X2=4.725 $Y2=1.542
r200 101 102 0.634211 $w=3.8e-07 $l=5e-09 $layer=POLY_cond $X=4.225 $Y=1.542
+ $X2=4.23 $Y2=1.542
r201 100 101 54.5421 $w=3.8e-07 $l=4.3e-07 $layer=POLY_cond $X=3.795 $Y=1.542
+ $X2=4.225 $Y2=1.542
r202 99 100 1.90263 $w=3.8e-07 $l=1.5e-08 $layer=POLY_cond $X=3.78 $Y=1.542
+ $X2=3.795 $Y2=1.542
r203 98 99 57.0789 $w=3.8e-07 $l=4.5e-07 $layer=POLY_cond $X=3.33 $Y=1.542
+ $X2=3.78 $Y2=1.542
r204 97 98 4.43947 $w=3.8e-07 $l=3.5e-08 $layer=POLY_cond $X=3.295 $Y=1.542
+ $X2=3.33 $Y2=1.542
r205 94 95 1.90263 $w=3.8e-07 $l=1.5e-08 $layer=POLY_cond $X=2.865 $Y=1.542
+ $X2=2.88 $Y2=1.542
r206 89 104 47.5658 $w=3.8e-07 $l=3.75e-07 $layer=POLY_cond $X=4.315 $Y=1.542
+ $X2=4.69 $Y2=1.542
r207 89 102 10.7816 $w=3.8e-07 $l=8.5e-08 $layer=POLY_cond $X=4.315 $Y=1.542
+ $X2=4.23 $Y2=1.542
r208 88 89 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=4.315
+ $Y=1.485 $X2=4.315 $Y2=1.485
r209 86 97 43.1263 $w=3.8e-07 $l=3.4e-07 $layer=POLY_cond $X=2.955 $Y=1.542
+ $X2=3.295 $Y2=1.542
r210 86 95 9.51316 $w=3.8e-07 $l=7.5e-08 $layer=POLY_cond $X=2.955 $Y=1.542
+ $X2=2.88 $Y2=1.542
r211 85 88 47.4946 $w=3.28e-07 $l=1.36e-06 $layer=LI1_cond $X=2.955 $Y=1.485
+ $X2=4.315 $Y2=1.485
r212 85 86 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=2.955
+ $Y=1.485 $X2=2.955 $Y2=1.485
r213 83 93 0.63164 $w=3.3e-07 $l=1e-07 $layer=LI1_cond $X=2.245 $Y=1.485
+ $X2=2.145 $Y2=1.485
r214 83 85 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=2.245 $Y=1.485
+ $X2=2.955 $Y2=1.485
r215 82 92 3.52026 $w=2.65e-07 $l=1.12916e-07 $layer=LI1_cond $X=2.145 $Y=1.8
+ $X2=2.08 $Y2=1.885
r216 81 93 8.10876 $w=1.85e-07 $l=1.65e-07 $layer=LI1_cond $X=2.145 $Y=1.65
+ $X2=2.145 $Y2=1.485
r217 81 82 8.31818 $w=1.98e-07 $l=1.5e-07 $layer=LI1_cond $X=2.145 $Y=1.65
+ $X2=2.145 $Y2=1.8
r218 80 93 8.10876 $w=1.85e-07 $l=1.72337e-07 $layer=LI1_cond $X=2.13 $Y=1.32
+ $X2=2.145 $Y2=1.485
r219 79 91 3.52026 $w=2.65e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.13 $Y=1.13
+ $X2=2.035 $Y2=1.045
r220 79 80 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=2.13 $Y=1.13
+ $X2=2.13 $Y2=1.32
r221 75 77 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=2.08 $Y=1.985
+ $X2=2.08 $Y2=2.815
r222 73 92 3.52026 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=2.08 $Y=1.97
+ $X2=2.08 $Y2=1.885
r223 73 75 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=2.08 $Y=1.97
+ $X2=2.08 $Y2=1.985
r224 69 91 3.52026 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=2.035 $Y=0.96
+ $X2=2.035 $Y2=1.045
r225 69 71 14.2455 $w=3.58e-07 $l=4.45e-07 $layer=LI1_cond $X=2.035 $Y=0.96
+ $X2=2.035 $Y2=0.515
r226 67 92 2.98021 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.915 $Y=1.885
+ $X2=2.08 $Y2=1.885
r227 67 68 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.915 $Y=1.885
+ $X2=1.345 $Y2=1.885
r228 65 91 2.98021 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=1.855 $Y=1.045
+ $X2=2.035 $Y2=1.045
r229 65 66 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=1.855 $Y=1.045
+ $X2=1.24 $Y2=1.045
r230 61 66 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.155 $Y=0.96
+ $X2=1.24 $Y2=1.045
r231 61 63 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=1.155 $Y=0.96
+ $X2=1.155 $Y2=0.515
r232 57 59 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=1.18 $Y=1.985
+ $X2=1.18 $Y2=2.815
r233 55 68 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.18 $Y=1.97
+ $X2=1.345 $Y2=1.885
r234 55 57 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=1.18 $Y=1.97
+ $X2=1.18 $Y2=1.985
r235 51 107 24.6126 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=5.155 $Y=1.32
+ $X2=5.155 $Y2=1.542
r236 51 53 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=5.155 $Y=1.32
+ $X2=5.155 $Y2=0.74
r237 48 106 24.6126 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=5.14 $Y=1.765
+ $X2=5.14 $Y2=1.542
r238 48 50 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.14 $Y=1.765
+ $X2=5.14 $Y2=2.4
r239 44 105 24.6126 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=4.725 $Y=1.32
+ $X2=4.725 $Y2=1.542
r240 44 46 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=4.725 $Y=1.32
+ $X2=4.725 $Y2=0.74
r241 41 104 24.6126 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=4.69 $Y=1.765
+ $X2=4.69 $Y2=1.542
r242 41 43 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.69 $Y=1.765
+ $X2=4.69 $Y2=2.4
r243 38 102 24.6126 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=4.23 $Y=1.765
+ $X2=4.23 $Y2=1.542
r244 38 40 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.23 $Y=1.765
+ $X2=4.23 $Y2=2.4
r245 34 101 24.6126 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=4.225 $Y=1.32
+ $X2=4.225 $Y2=1.542
r246 34 36 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=4.225 $Y=1.32
+ $X2=4.225 $Y2=0.74
r247 30 100 24.6126 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=3.795 $Y=1.32
+ $X2=3.795 $Y2=1.542
r248 30 32 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.795 $Y=1.32
+ $X2=3.795 $Y2=0.74
r249 27 99 24.6126 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=3.78 $Y=1.765
+ $X2=3.78 $Y2=1.542
r250 27 29 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.78 $Y=1.765
+ $X2=3.78 $Y2=2.4
r251 24 98 24.6126 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=3.33 $Y=1.765
+ $X2=3.33 $Y2=1.542
r252 24 26 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.33 $Y=1.765
+ $X2=3.33 $Y2=2.4
r253 20 97 24.6126 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=3.295 $Y=1.32
+ $X2=3.295 $Y2=1.542
r254 20 22 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.295 $Y=1.32
+ $X2=3.295 $Y2=0.74
r255 17 95 24.6126 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=2.88 $Y=1.765
+ $X2=2.88 $Y2=1.542
r256 17 19 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.88 $Y=1.765
+ $X2=2.88 $Y2=2.4
r257 13 94 24.6126 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=2.865 $Y=1.32
+ $X2=2.865 $Y2=1.542
r258 13 15 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.865 $Y=1.32
+ $X2=2.865 $Y2=0.74
r259 4 77 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.93
+ $Y=1.84 $X2=2.08 $Y2=2.815
r260 4 75 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.93
+ $Y=1.84 $X2=2.08 $Y2=1.985
r261 3 59 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.03
+ $Y=1.84 $X2=1.18 $Y2=2.815
r262 3 57 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.03
+ $Y=1.84 $X2=1.18 $Y2=1.985
r263 2 71 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.88
+ $Y=0.37 $X2=2.02 $Y2=0.515
r264 1 63 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.015
+ $Y=0.37 $X2=1.155 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__BUFBUF_16%A_588_74# 1 2 3 4 5 6 21 23 25 28 30 32 35
+ 37 39 42 44 46 49 51 53 56 58 60 63 65 67 70 72 74 77 79 81 84 86 88 91 93 95
+ 98 100 102 105 107 109 112 114 116 117 119 122 126 128 130 133 135 137 139 140
+ 141 145 149 151 153 155 157 161 164 168 169 170 194 203 210 217 224 231 238
+ 245 248
c482 155 0 1.38532e-19 $X=4.915 $Y=1.99
c483 112 0 9.40629e-20 $X=11.455 $Y=0.74
c484 37 0 1.0086e-19 $X=6.55 $Y=1.765
c485 30 0 1.79811e-19 $X=6.05 $Y=1.765
c486 23 0 1.89809e-19 $X=5.6 $Y=1.765
r487 279 281 2.0766 $w=4.7e-07 $l=8e-08 $layer=LI1_cond $X=5.077 $Y=1.905
+ $X2=5.077 $Y2=1.985
r488 248 249 7.03183 $w=3.77e-07 $l=5.5e-08 $layer=POLY_cond $X=12.395 $Y=1.542
+ $X2=12.45 $Y2=1.542
r489 247 248 54.9761 $w=3.77e-07 $l=4.3e-07 $layer=POLY_cond $X=11.965 $Y=1.542
+ $X2=12.395 $Y2=1.542
r490 246 247 1.91777 $w=3.77e-07 $l=1.5e-08 $layer=POLY_cond $X=11.95 $Y=1.542
+ $X2=11.965 $Y2=1.542
r491 244 246 33.8806 $w=3.77e-07 $l=2.65e-07 $layer=POLY_cond $X=11.685 $Y=1.542
+ $X2=11.95 $Y2=1.542
r492 244 245 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.685
+ $Y=1.485 $X2=11.685 $Y2=1.485
r493 242 244 23.6525 $w=3.77e-07 $l=1.85e-07 $layer=POLY_cond $X=11.5 $Y=1.542
+ $X2=11.685 $Y2=1.542
r494 241 242 5.75332 $w=3.77e-07 $l=4.5e-08 $layer=POLY_cond $X=11.455 $Y=1.542
+ $X2=11.5 $Y2=1.542
r495 240 241 51.7798 $w=3.77e-07 $l=4.05e-07 $layer=POLY_cond $X=11.05 $Y=1.542
+ $X2=11.455 $Y2=1.542
r496 239 240 3.19629 $w=3.77e-07 $l=2.5e-08 $layer=POLY_cond $X=11.025 $Y=1.542
+ $X2=11.05 $Y2=1.542
r497 237 239 33.8806 $w=3.77e-07 $l=2.65e-07 $layer=POLY_cond $X=10.76 $Y=1.542
+ $X2=11.025 $Y2=1.542
r498 237 238 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.76
+ $Y=1.485 $X2=10.76 $Y2=1.485
r499 235 237 20.4562 $w=3.77e-07 $l=1.6e-07 $layer=POLY_cond $X=10.6 $Y=1.542
+ $X2=10.76 $Y2=1.542
r500 234 235 9.58886 $w=3.77e-07 $l=7.5e-08 $layer=POLY_cond $X=10.525 $Y=1.542
+ $X2=10.6 $Y2=1.542
r501 233 234 47.9443 $w=3.77e-07 $l=3.75e-07 $layer=POLY_cond $X=10.15 $Y=1.542
+ $X2=10.525 $Y2=1.542
r502 232 233 7.03183 $w=3.77e-07 $l=5.5e-08 $layer=POLY_cond $X=10.095 $Y=1.542
+ $X2=10.15 $Y2=1.542
r503 230 232 35.7984 $w=3.77e-07 $l=2.8e-07 $layer=POLY_cond $X=9.815 $Y=1.542
+ $X2=10.095 $Y2=1.542
r504 230 231 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.815
+ $Y=1.485 $X2=9.815 $Y2=1.485
r505 228 230 14.7029 $w=3.77e-07 $l=1.15e-07 $layer=POLY_cond $X=9.7 $Y=1.542
+ $X2=9.815 $Y2=1.542
r506 227 228 13.4244 $w=3.77e-07 $l=1.05e-07 $layer=POLY_cond $X=9.595 $Y=1.542
+ $X2=9.7 $Y2=1.542
r507 226 227 44.1088 $w=3.77e-07 $l=3.45e-07 $layer=POLY_cond $X=9.25 $Y=1.542
+ $X2=9.595 $Y2=1.542
r508 225 226 10.8674 $w=3.77e-07 $l=8.5e-08 $layer=POLY_cond $X=9.165 $Y=1.542
+ $X2=9.25 $Y2=1.542
r509 223 225 33.2414 $w=3.77e-07 $l=2.6e-07 $layer=POLY_cond $X=8.905 $Y=1.542
+ $X2=9.165 $Y2=1.542
r510 223 224 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.905
+ $Y=1.485 $X2=8.905 $Y2=1.485
r511 221 223 13.4244 $w=3.77e-07 $l=1.05e-07 $layer=POLY_cond $X=8.8 $Y=1.542
+ $X2=8.905 $Y2=1.542
r512 220 221 17.2599 $w=3.77e-07 $l=1.35e-07 $layer=POLY_cond $X=8.665 $Y=1.542
+ $X2=8.8 $Y2=1.542
r513 219 220 40.2732 $w=3.77e-07 $l=3.15e-07 $layer=POLY_cond $X=8.35 $Y=1.542
+ $X2=8.665 $Y2=1.542
r514 218 219 14.7029 $w=3.77e-07 $l=1.15e-07 $layer=POLY_cond $X=8.235 $Y=1.542
+ $X2=8.35 $Y2=1.542
r515 216 218 31.9629 $w=3.77e-07 $l=2.5e-07 $layer=POLY_cond $X=7.985 $Y=1.542
+ $X2=8.235 $Y2=1.542
r516 216 217 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.985
+ $Y=1.485 $X2=7.985 $Y2=1.485
r517 214 216 10.8674 $w=3.77e-07 $l=8.5e-08 $layer=POLY_cond $X=7.9 $Y=1.542
+ $X2=7.985 $Y2=1.542
r518 213 214 21.0955 $w=3.77e-07 $l=1.65e-07 $layer=POLY_cond $X=7.735 $Y=1.542
+ $X2=7.9 $Y2=1.542
r519 212 213 36.4377 $w=3.77e-07 $l=2.85e-07 $layer=POLY_cond $X=7.45 $Y=1.542
+ $X2=7.735 $Y2=1.542
r520 211 212 18.5385 $w=3.77e-07 $l=1.45e-07 $layer=POLY_cond $X=7.305 $Y=1.542
+ $X2=7.45 $Y2=1.542
r521 209 211 28.1273 $w=3.77e-07 $l=2.2e-07 $layer=POLY_cond $X=7.085 $Y=1.542
+ $X2=7.305 $Y2=1.542
r522 209 210 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.085
+ $Y=1.485 $X2=7.085 $Y2=1.485
r523 207 209 10.8674 $w=3.77e-07 $l=8.5e-08 $layer=POLY_cond $X=7 $Y=1.542
+ $X2=7.085 $Y2=1.542
r524 206 207 15.9814 $w=3.77e-07 $l=1.25e-07 $layer=POLY_cond $X=6.875 $Y=1.542
+ $X2=7 $Y2=1.542
r525 205 206 41.5517 $w=3.77e-07 $l=3.25e-07 $layer=POLY_cond $X=6.55 $Y=1.542
+ $X2=6.875 $Y2=1.542
r526 204 205 13.4244 $w=3.77e-07 $l=1.05e-07 $layer=POLY_cond $X=6.445 $Y=1.542
+ $X2=6.55 $Y2=1.542
r527 202 204 30.0451 $w=3.77e-07 $l=2.35e-07 $layer=POLY_cond $X=6.21 $Y=1.542
+ $X2=6.445 $Y2=1.542
r528 202 203 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.21
+ $Y=1.485 $X2=6.21 $Y2=1.485
r529 200 202 20.4562 $w=3.77e-07 $l=1.6e-07 $layer=POLY_cond $X=6.05 $Y=1.542
+ $X2=6.21 $Y2=1.542
r530 199 200 4.4748 $w=3.77e-07 $l=3.5e-08 $layer=POLY_cond $X=6.015 $Y=1.542
+ $X2=6.05 $Y2=1.542
r531 198 199 53.0584 $w=3.77e-07 $l=4.15e-07 $layer=POLY_cond $X=5.6 $Y=1.542
+ $X2=6.015 $Y2=1.542
r532 197 198 1.91777 $w=3.77e-07 $l=1.5e-08 $layer=POLY_cond $X=5.585 $Y=1.542
+ $X2=5.6 $Y2=1.542
r533 195 245 5.25164 $w=3.93e-07 $l=1.8e-07 $layer=LI1_cond $X=11.692 $Y=1.665
+ $X2=11.692 $Y2=1.485
r534 194 195 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.685 $Y=1.665
+ $X2=11.685 $Y2=1.665
r535 192 238 5.53173 $w=3.73e-07 $l=1.8e-07 $layer=LI1_cond $X=10.752 $Y=1.665
+ $X2=10.752 $Y2=1.485
r536 191 194 0.593484 $w=2.3e-07 $l=9.25e-07 $layer=MET1_cond $X=10.76 $Y=1.665
+ $X2=11.685 $Y2=1.665
r537 191 192 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.76 $Y=1.665
+ $X2=10.76 $Y2=1.665
r538 189 231 6.38276 $w=3.23e-07 $l=1.8e-07 $layer=LI1_cond $X=9.812 $Y=1.665
+ $X2=9.812 $Y2=1.485
r539 188 191 0.606316 $w=2.3e-07 $l=9.45e-07 $layer=MET1_cond $X=9.815 $Y=1.665
+ $X2=10.76 $Y2=1.665
r540 188 189 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.815 $Y=1.665
+ $X2=9.815 $Y2=1.665
r541 186 224 7.03186 $w=2.93e-07 $l=1.8e-07 $layer=LI1_cond $X=8.897 $Y=1.665
+ $X2=8.897 $Y2=1.485
r542 185 188 0.58386 $w=2.3e-07 $l=9.1e-07 $layer=MET1_cond $X=8.905 $Y=1.665
+ $X2=9.815 $Y2=1.665
r543 185 186 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.905 $Y=1.665
+ $X2=8.905 $Y2=1.665
r544 183 217 7.82791 $w=2.63e-07 $l=1.8e-07 $layer=LI1_cond $X=7.982 $Y=1.665
+ $X2=7.982 $Y2=1.485
r545 182 185 0.590276 $w=2.3e-07 $l=9.2e-07 $layer=MET1_cond $X=7.985 $Y=1.665
+ $X2=8.905 $Y2=1.665
r546 182 183 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.985 $Y=1.665
+ $X2=7.985 $Y2=1.665
r547 180 210 7.82791 $w=2.63e-07 $l=1.8e-07 $layer=LI1_cond $X=7.082 $Y=1.665
+ $X2=7.082 $Y2=1.485
r548 179 182 0.577444 $w=2.3e-07 $l=9e-07 $layer=MET1_cond $X=7.085 $Y=1.665
+ $X2=7.985 $Y2=1.665
r549 179 180 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.085 $Y=1.665
+ $X2=7.085 $Y2=1.665
r550 177 203 6.6916 $w=3.08e-07 $l=1.8e-07 $layer=LI1_cond $X=6.21 $Y=1.665
+ $X2=6.21 $Y2=1.485
r551 176 179 0.561404 $w=2.3e-07 $l=8.75e-07 $layer=MET1_cond $X=6.21 $Y=1.665
+ $X2=7.085 $Y2=1.665
r552 176 177 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=1.665
+ $X2=6.21 $Y2=1.665
r553 173 279 6.22979 $w=4.7e-07 $l=2.4e-07 $layer=LI1_cond $X=5.077 $Y=1.665
+ $X2=5.077 $Y2=1.905
r554 172 176 0.606316 $w=2.3e-07 $l=9.45e-07 $layer=MET1_cond $X=5.265 $Y=1.665
+ $X2=6.21 $Y2=1.665
r555 172 173 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.265 $Y=1.665
+ $X2=5.265 $Y2=1.665
r556 164 173 11.3723 $w=4.7e-07 $l=3.92702e-07 $layer=LI1_cond $X=4.975 $Y=1.32
+ $X2=5.077 $Y2=1.665
r557 163 170 3.64284 $w=2.55e-07 $l=1.00995e-07 $layer=LI1_cond $X=4.975 $Y=1.15
+ $X2=4.94 $Y2=1.065
r558 163 164 7.5352 $w=2.58e-07 $l=1.7e-07 $layer=LI1_cond $X=4.975 $Y=1.15
+ $X2=4.975 $Y2=1.32
r559 159 170 3.64284 $w=2.55e-07 $l=1.03078e-07 $layer=LI1_cond $X=4.9 $Y=0.98
+ $X2=4.94 $Y2=1.065
r560 159 161 21.4354 $w=2.48e-07 $l=4.65e-07 $layer=LI1_cond $X=4.9 $Y=0.98
+ $X2=4.9 $Y2=0.515
r561 155 281 1.22671 $w=4.7e-07 $l=1.64481e-07 $layer=LI1_cond $X=4.915 $Y=1.99
+ $X2=5.077 $Y2=1.985
r562 155 157 28.8111 $w=3.28e-07 $l=8.25e-07 $layer=LI1_cond $X=4.915 $Y=1.99
+ $X2=4.915 $Y2=2.815
r563 154 168 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.17 $Y=1.905
+ $X2=4.005 $Y2=1.905
r564 153 279 6.76998 $w=1.7e-07 $l=3.27e-07 $layer=LI1_cond $X=4.75 $Y=1.905
+ $X2=5.077 $Y2=1.905
r565 153 154 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=4.75 $Y=1.905
+ $X2=4.17 $Y2=1.905
r566 152 169 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.095 $Y=1.065
+ $X2=3.97 $Y2=1.065
r567 151 170 2.83584 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.775 $Y=1.065
+ $X2=4.94 $Y2=1.065
r568 151 152 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.775 $Y=1.065
+ $X2=4.095 $Y2=1.065
r569 147 169 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.97 $Y=0.98
+ $X2=3.97 $Y2=1.065
r570 147 149 21.4354 $w=2.48e-07 $l=4.65e-07 $layer=LI1_cond $X=3.97 $Y=0.98
+ $X2=3.97 $Y2=0.515
r571 143 168 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.005 $Y=1.99
+ $X2=4.005 $Y2=1.905
r572 143 145 28.8111 $w=3.28e-07 $l=8.25e-07 $layer=LI1_cond $X=4.005 $Y=1.99
+ $X2=4.005 $Y2=2.815
r573 142 166 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.27 $Y=1.905
+ $X2=3.105 $Y2=1.905
r574 141 168 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.84 $Y=1.905
+ $X2=4.005 $Y2=1.905
r575 141 142 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=3.84 $Y=1.905
+ $X2=3.27 $Y2=1.905
r576 139 169 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.845 $Y=1.065
+ $X2=3.97 $Y2=1.065
r577 139 140 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.845 $Y=1.065
+ $X2=3.165 $Y2=1.065
r578 135 166 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.105 $Y=1.99
+ $X2=3.105 $Y2=1.905
r579 135 137 28.8111 $w=3.28e-07 $l=8.25e-07 $layer=LI1_cond $X=3.105 $Y=1.99
+ $X2=3.105 $Y2=2.815
r580 131 140 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.04 $Y=0.98
+ $X2=3.165 $Y2=1.065
r581 131 133 21.4354 $w=2.48e-07 $l=4.65e-07 $layer=LI1_cond $X=3.04 $Y=0.98
+ $X2=3.04 $Y2=0.515
r582 128 249 24.4204 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=12.45 $Y=1.765
+ $X2=12.45 $Y2=1.542
r583 128 130 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=12.45 $Y=1.765
+ $X2=12.45 $Y2=2.4
r584 124 248 24.4204 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=12.395 $Y=1.32
+ $X2=12.395 $Y2=1.542
r585 124 126 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=12.395 $Y=1.32
+ $X2=12.395 $Y2=0.74
r586 120 247 24.4204 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=11.965 $Y=1.32
+ $X2=11.965 $Y2=1.542
r587 120 122 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=11.965 $Y=1.32
+ $X2=11.965 $Y2=0.74
r588 117 246 24.4204 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=11.95 $Y=1.765
+ $X2=11.95 $Y2=1.542
r589 117 119 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=11.95 $Y=1.765
+ $X2=11.95 $Y2=2.4
r590 114 242 24.4204 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=11.5 $Y=1.765
+ $X2=11.5 $Y2=1.542
r591 114 116 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=11.5 $Y=1.765
+ $X2=11.5 $Y2=2.4
r592 110 241 24.4204 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=11.455 $Y=1.32
+ $X2=11.455 $Y2=1.542
r593 110 112 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=11.455 $Y=1.32
+ $X2=11.455 $Y2=0.74
r594 107 240 24.4204 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=11.05 $Y=1.765
+ $X2=11.05 $Y2=1.542
r595 107 109 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=11.05 $Y=1.765
+ $X2=11.05 $Y2=2.4
r596 103 239 24.4204 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=11.025 $Y=1.32
+ $X2=11.025 $Y2=1.542
r597 103 105 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=11.025 $Y=1.32
+ $X2=11.025 $Y2=0.74
r598 100 235 24.4204 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=10.6 $Y=1.765
+ $X2=10.6 $Y2=1.542
r599 100 102 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=10.6 $Y=1.765
+ $X2=10.6 $Y2=2.4
r600 96 234 24.4204 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=10.525 $Y=1.32
+ $X2=10.525 $Y2=1.542
r601 96 98 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=10.525 $Y=1.32
+ $X2=10.525 $Y2=0.74
r602 93 233 24.4204 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=10.15 $Y=1.765
+ $X2=10.15 $Y2=1.542
r603 93 95 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=10.15 $Y=1.765
+ $X2=10.15 $Y2=2.4
r604 89 232 24.4204 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=10.095 $Y=1.32
+ $X2=10.095 $Y2=1.542
r605 89 91 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=10.095 $Y=1.32
+ $X2=10.095 $Y2=0.74
r606 86 228 24.4204 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=9.7 $Y=1.765
+ $X2=9.7 $Y2=1.542
r607 86 88 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=9.7 $Y=1.765
+ $X2=9.7 $Y2=2.4
r608 82 227 24.4204 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=9.595 $Y=1.32
+ $X2=9.595 $Y2=1.542
r609 82 84 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=9.595 $Y=1.32
+ $X2=9.595 $Y2=0.74
r610 79 226 24.4204 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=9.25 $Y=1.765
+ $X2=9.25 $Y2=1.542
r611 79 81 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=9.25 $Y=1.765
+ $X2=9.25 $Y2=2.4
r612 75 225 24.4204 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=9.165 $Y=1.32
+ $X2=9.165 $Y2=1.542
r613 75 77 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=9.165 $Y=1.32
+ $X2=9.165 $Y2=0.74
r614 72 221 24.4204 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=8.8 $Y=1.765
+ $X2=8.8 $Y2=1.542
r615 72 74 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.8 $Y=1.765
+ $X2=8.8 $Y2=2.4
r616 68 220 24.4204 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=8.665 $Y=1.32
+ $X2=8.665 $Y2=1.542
r617 68 70 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=8.665 $Y=1.32
+ $X2=8.665 $Y2=0.74
r618 65 219 24.4204 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=8.35 $Y=1.765
+ $X2=8.35 $Y2=1.542
r619 65 67 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.35 $Y=1.765
+ $X2=8.35 $Y2=2.4
r620 61 218 24.4204 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=8.235 $Y=1.32
+ $X2=8.235 $Y2=1.542
r621 61 63 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=8.235 $Y=1.32
+ $X2=8.235 $Y2=0.74
r622 58 214 24.4204 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=7.9 $Y=1.765
+ $X2=7.9 $Y2=1.542
r623 58 60 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.9 $Y=1.765
+ $X2=7.9 $Y2=2.4
r624 54 213 24.4204 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=7.735 $Y=1.32
+ $X2=7.735 $Y2=1.542
r625 54 56 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=7.735 $Y=1.32
+ $X2=7.735 $Y2=0.74
r626 51 212 24.4204 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=7.45 $Y=1.765
+ $X2=7.45 $Y2=1.542
r627 51 53 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.45 $Y=1.765
+ $X2=7.45 $Y2=2.4
r628 47 211 24.4204 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=7.305 $Y=1.32
+ $X2=7.305 $Y2=1.542
r629 47 49 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=7.305 $Y=1.32
+ $X2=7.305 $Y2=0.74
r630 44 207 24.4204 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=7 $Y=1.765 $X2=7
+ $Y2=1.542
r631 44 46 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7 $Y=1.765 $X2=7
+ $Y2=2.4
r632 40 206 24.4204 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=6.875 $Y=1.32
+ $X2=6.875 $Y2=1.542
r633 40 42 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.875 $Y=1.32
+ $X2=6.875 $Y2=0.74
r634 37 205 24.4204 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=6.55 $Y=1.765
+ $X2=6.55 $Y2=1.542
r635 37 39 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.55 $Y=1.765
+ $X2=6.55 $Y2=2.4
r636 33 204 24.4204 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=6.445 $Y=1.32
+ $X2=6.445 $Y2=1.542
r637 33 35 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.445 $Y=1.32
+ $X2=6.445 $Y2=0.74
r638 30 200 24.4204 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=6.05 $Y=1.765
+ $X2=6.05 $Y2=1.542
r639 30 32 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.05 $Y=1.765
+ $X2=6.05 $Y2=2.4
r640 26 199 24.4204 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=6.015 $Y=1.32
+ $X2=6.015 $Y2=1.542
r641 26 28 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.015 $Y=1.32
+ $X2=6.015 $Y2=0.74
r642 23 198 24.4204 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=5.6 $Y=1.765
+ $X2=5.6 $Y2=1.542
r643 23 25 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.6 $Y=1.765
+ $X2=5.6 $Y2=2.4
r644 19 197 24.4204 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=5.585 $Y=1.32
+ $X2=5.585 $Y2=1.542
r645 19 21 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=5.585 $Y=1.32
+ $X2=5.585 $Y2=0.74
r646 6 281 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=4.765
+ $Y=1.84 $X2=4.915 $Y2=1.985
r647 6 157 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=4.765
+ $Y=1.84 $X2=4.915 $Y2=2.815
r648 5 168 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=3.855
+ $Y=1.84 $X2=4.005 $Y2=1.985
r649 5 145 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=3.855
+ $Y=1.84 $X2=4.005 $Y2=2.815
r650 4 166 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.955
+ $Y=1.84 $X2=3.105 $Y2=1.985
r651 4 137 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.955
+ $Y=1.84 $X2=3.105 $Y2=2.815
r652 3 161 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.8
+ $Y=0.37 $X2=4.94 $Y2=0.515
r653 2 149 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.87
+ $Y=0.37 $X2=4.01 $Y2=0.515
r654 1 133 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.94
+ $Y=0.37 $X2=3.08 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__BUFBUF_16%VPWR 1 2 3 4 5 6 7 8 9 10 11 12 13 14 47
+ 51 55 61 65 69 75 79 83 89 93 97 101 105 111 115 117 122 123 125 126 128 129
+ 131 132 134 135 137 138 140 141 142 143 144 150 176 181 187 190 193 196 199
+ 203
r232 202 203 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r233 199 200 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r234 196 197 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r235 194 197 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=10.8 $Y2=3.33
r236 193 194 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r237 190 191 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r238 187 188 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r239 185 203 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=12.72 $Y2=3.33
r240 185 200 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=11.76 $Y2=3.33
r241 184 185 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r242 182 199 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.89 $Y=3.33
+ $X2=11.765 $Y2=3.33
r243 182 184 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=11.89 $Y=3.33
+ $X2=12.24 $Y2=3.33
r244 181 202 4.0045 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=12.59 $Y=3.33
+ $X2=12.775 $Y2=3.33
r245 181 184 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=12.59 $Y=3.33
+ $X2=12.24 $Y2=3.33
r246 180 200 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=11.76 $Y2=3.33
r247 180 197 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=10.8 $Y2=3.33
r248 179 180 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r249 177 196 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.91 $Y=3.33
+ $X2=10.825 $Y2=3.33
r250 177 179 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=10.91 $Y=3.33
+ $X2=11.28 $Y2=3.33
r251 176 199 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.64 $Y=3.33
+ $X2=11.765 $Y2=3.33
r252 176 179 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=11.64 $Y=3.33
+ $X2=11.28 $Y2=3.33
r253 175 194 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=9.84 $Y2=3.33
r254 174 175 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r255 172 175 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.88 $Y2=3.33
r256 171 172 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r257 169 172 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.92 $Y2=3.33
r258 168 169 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r259 165 166 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r260 163 166 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=6 $Y2=3.33
r261 162 163 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r262 160 163 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r263 159 160 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r264 157 160 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r265 157 191 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r266 156 157 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r267 154 190 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.74 $Y=3.33
+ $X2=2.615 $Y2=3.33
r268 154 156 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=2.74 $Y=3.33
+ $X2=3.12 $Y2=3.33
r269 153 191 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r270 152 153 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r271 150 190 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.49 $Y=3.33
+ $X2=2.615 $Y2=3.33
r272 150 152 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.49 $Y=3.33
+ $X2=2.16 $Y2=3.33
r273 149 153 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r274 149 188 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r275 148 149 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r276 146 187 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=3.33
+ $X2=0.73 $Y2=3.33
r277 146 148 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.815 $Y=3.33
+ $X2=1.2 $Y2=3.33
r278 144 169 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6.96 $Y2=3.33
r279 144 166 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6 $Y2=3.33
r280 142 174 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=8.94 $Y=3.33
+ $X2=8.88 $Y2=3.33
r281 142 143 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.94 $Y=3.33
+ $X2=9.025 $Y2=3.33
r282 140 171 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=8.04 $Y=3.33
+ $X2=7.92 $Y2=3.33
r283 140 141 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.04 $Y=3.33
+ $X2=8.125 $Y2=3.33
r284 139 174 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.21 $Y=3.33
+ $X2=8.88 $Y2=3.33
r285 139 141 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.21 $Y=3.33
+ $X2=8.125 $Y2=3.33
r286 137 168 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=7.14 $Y=3.33
+ $X2=6.96 $Y2=3.33
r287 137 138 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.14 $Y=3.33
+ $X2=7.225 $Y2=3.33
r288 136 171 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=7.31 $Y=3.33
+ $X2=7.92 $Y2=3.33
r289 136 138 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.31 $Y=3.33
+ $X2=7.225 $Y2=3.33
r290 134 165 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=6.16 $Y=3.33
+ $X2=6 $Y2=3.33
r291 134 135 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.16 $Y=3.33
+ $X2=6.285 $Y2=3.33
r292 133 168 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=6.41 $Y=3.33
+ $X2=6.96 $Y2=3.33
r293 133 135 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.41 $Y=3.33
+ $X2=6.285 $Y2=3.33
r294 131 162 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=5.28 $Y=3.33
+ $X2=5.04 $Y2=3.33
r295 131 132 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.28 $Y=3.33
+ $X2=5.365 $Y2=3.33
r296 130 165 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=5.45 $Y=3.33
+ $X2=6 $Y2=3.33
r297 130 132 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.45 $Y=3.33
+ $X2=5.365 $Y2=3.33
r298 128 159 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=4.37 $Y=3.33
+ $X2=4.08 $Y2=3.33
r299 128 129 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.37 $Y=3.33
+ $X2=4.455 $Y2=3.33
r300 127 162 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=4.54 $Y=3.33
+ $X2=5.04 $Y2=3.33
r301 127 129 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.54 $Y=3.33
+ $X2=4.455 $Y2=3.33
r302 125 156 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=3.47 $Y=3.33
+ $X2=3.12 $Y2=3.33
r303 125 126 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.47 $Y=3.33
+ $X2=3.555 $Y2=3.33
r304 124 159 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=3.64 $Y=3.33
+ $X2=4.08 $Y2=3.33
r305 124 126 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.64 $Y=3.33
+ $X2=3.555 $Y2=3.33
r306 122 148 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.545 $Y=3.33
+ $X2=1.2 $Y2=3.33
r307 122 123 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.545 $Y=3.33
+ $X2=1.63 $Y2=3.33
r308 121 152 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=1.715 $Y=3.33
+ $X2=2.16 $Y2=3.33
r309 121 123 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.715 $Y=3.33
+ $X2=1.63 $Y2=3.33
r310 117 120 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=12.715 $Y=1.985
+ $X2=12.715 $Y2=2.815
r311 115 202 3.13866 $w=2.5e-07 $l=1.11018e-07 $layer=LI1_cond $X=12.715
+ $Y=3.245 $X2=12.775 $Y2=3.33
r312 115 120 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=12.715 $Y=3.245
+ $X2=12.715 $Y2=2.815
r313 111 114 33.4208 $w=2.48e-07 $l=7.25e-07 $layer=LI1_cond $X=11.765 $Y=2.09
+ $X2=11.765 $Y2=2.815
r314 109 199 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=11.765 $Y=3.245
+ $X2=11.765 $Y2=3.33
r315 109 114 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=11.765 $Y=3.245
+ $X2=11.765 $Y2=2.815
r316 105 108 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=10.825 $Y=2.09
+ $X2=10.825 $Y2=2.815
r317 103 196 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.825 $Y=3.245
+ $X2=10.825 $Y2=3.33
r318 103 108 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=10.825 $Y=3.245
+ $X2=10.825 $Y2=2.815
r319 102 193 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.01 $Y=3.33
+ $X2=9.925 $Y2=3.33
r320 101 196 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.74 $Y=3.33
+ $X2=10.825 $Y2=3.33
r321 101 102 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=10.74 $Y=3.33
+ $X2=10.01 $Y2=3.33
r322 97 100 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=9.925 $Y=2.09
+ $X2=9.925 $Y2=2.815
r323 95 193 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.925 $Y=3.245
+ $X2=9.925 $Y2=3.33
r324 95 100 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=9.925 $Y=3.245
+ $X2=9.925 $Y2=2.815
r325 94 143 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.11 $Y=3.33
+ $X2=9.025 $Y2=3.33
r326 93 193 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.84 $Y=3.33
+ $X2=9.925 $Y2=3.33
r327 93 94 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=9.84 $Y=3.33
+ $X2=9.11 $Y2=3.33
r328 89 92 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=9.025 $Y=2.09
+ $X2=9.025 $Y2=2.815
r329 87 143 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.025 $Y=3.245
+ $X2=9.025 $Y2=3.33
r330 87 92 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=9.025 $Y=3.245
+ $X2=9.025 $Y2=2.815
r331 83 86 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=8.125 $Y=2.09
+ $X2=8.125 $Y2=2.815
r332 81 141 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.125 $Y=3.245
+ $X2=8.125 $Y2=3.33
r333 81 86 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=8.125 $Y=3.245
+ $X2=8.125 $Y2=2.815
r334 77 138 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.225 $Y=3.245
+ $X2=7.225 $Y2=3.33
r335 77 79 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=7.225 $Y=3.245
+ $X2=7.225 $Y2=2.325
r336 73 135 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.285 $Y=3.245
+ $X2=6.285 $Y2=3.33
r337 73 75 42.4099 $w=2.48e-07 $l=9.2e-07 $layer=LI1_cond $X=6.285 $Y=3.245
+ $X2=6.285 $Y2=2.325
r338 69 72 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=5.365 $Y=2.09
+ $X2=5.365 $Y2=2.815
r339 67 132 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.365 $Y=3.245
+ $X2=5.365 $Y2=3.33
r340 67 72 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=5.365 $Y=3.245
+ $X2=5.365 $Y2=2.815
r341 63 129 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.455 $Y=3.245
+ $X2=4.455 $Y2=3.33
r342 63 65 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=4.455 $Y=3.245
+ $X2=4.455 $Y2=2.325
r343 59 126 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.555 $Y=3.245
+ $X2=3.555 $Y2=3.33
r344 59 61 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=3.555 $Y=3.245
+ $X2=3.555 $Y2=2.325
r345 55 58 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=2.615 $Y=1.985
+ $X2=2.615 $Y2=2.815
r346 53 190 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.615 $Y=3.245
+ $X2=2.615 $Y2=3.33
r347 53 58 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=2.615 $Y=3.245
+ $X2=2.615 $Y2=2.815
r348 49 123 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.63 $Y=3.245
+ $X2=1.63 $Y2=3.33
r349 49 51 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=1.63 $Y=3.245
+ $X2=1.63 $Y2=2.305
r350 45 187 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=3.33
r351 45 47 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=2.455
r352 14 120 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=12.525
+ $Y=1.84 $X2=12.675 $Y2=2.815
r353 14 117 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=12.525
+ $Y=1.84 $X2=12.675 $Y2=1.985
r354 13 114 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=11.575
+ $Y=1.84 $X2=11.725 $Y2=2.815
r355 13 111 400 $w=1.7e-07 $l=3.16228e-07 $layer=licon1_PDIFF $count=1 $X=11.575
+ $Y=1.84 $X2=11.725 $Y2=2.09
r356 12 108 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=10.675
+ $Y=1.84 $X2=10.825 $Y2=2.815
r357 12 105 400 $w=1.7e-07 $l=3.16228e-07 $layer=licon1_PDIFF $count=1 $X=10.675
+ $Y=1.84 $X2=10.825 $Y2=2.09
r358 11 100 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=9.775
+ $Y=1.84 $X2=9.925 $Y2=2.815
r359 11 97 400 $w=1.7e-07 $l=3.16228e-07 $layer=licon1_PDIFF $count=1 $X=9.775
+ $Y=1.84 $X2=9.925 $Y2=2.09
r360 10 92 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=8.875
+ $Y=1.84 $X2=9.025 $Y2=2.815
r361 10 89 400 $w=1.7e-07 $l=3.16228e-07 $layer=licon1_PDIFF $count=1 $X=8.875
+ $Y=1.84 $X2=9.025 $Y2=2.09
r362 9 86 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=7.975
+ $Y=1.84 $X2=8.125 $Y2=2.815
r363 9 83 400 $w=1.7e-07 $l=3.16228e-07 $layer=licon1_PDIFF $count=1 $X=7.975
+ $Y=1.84 $X2=8.125 $Y2=2.09
r364 8 79 300 $w=1.7e-07 $l=5.54955e-07 $layer=licon1_PDIFF $count=2 $X=7.075
+ $Y=1.84 $X2=7.225 $Y2=2.325
r365 7 75 300 $w=1.7e-07 $l=5.7639e-07 $layer=licon1_PDIFF $count=2 $X=6.125
+ $Y=1.84 $X2=6.325 $Y2=2.325
r366 6 72 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=5.215
+ $Y=1.84 $X2=5.365 $Y2=2.815
r367 6 69 400 $w=1.7e-07 $l=3.16228e-07 $layer=licon1_PDIFF $count=1 $X=5.215
+ $Y=1.84 $X2=5.365 $Y2=2.09
r368 5 65 300 $w=1.7e-07 $l=5.54955e-07 $layer=licon1_PDIFF $count=2 $X=4.305
+ $Y=1.84 $X2=4.455 $Y2=2.325
r369 4 61 300 $w=1.7e-07 $l=5.54955e-07 $layer=licon1_PDIFF $count=2 $X=3.405
+ $Y=1.84 $X2=3.555 $Y2=2.325
r370 3 58 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=2.51
+ $Y=1.84 $X2=2.655 $Y2=2.815
r371 3 55 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=2.51
+ $Y=1.84 $X2=2.655 $Y2=1.985
r372 2 51 300 $w=1.7e-07 $l=5.34766e-07 $layer=licon1_PDIFF $count=2 $X=1.48
+ $Y=1.84 $X2=1.63 $Y2=2.305
r373 1 47 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=0.58
+ $Y=1.84 $X2=0.73 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_LS__BUFBUF_16%X 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16
+ 51 53 55 59 65 69 75 79 85 89 95 99 105 109 113 117 122 125 127 128 129 130
+ 131 132 133 140 141 145 146 150 151 155 156 160 161 165 170 171
c283 171 0 1.38532e-19 $X=12.2 $Y=2.035
c284 161 0 3.07445e-20 $X=10.375 $Y=1.92
c285 156 0 3.07333e-20 $X=9.475 $Y=1.92
c286 151 0 3.07333e-20 $X=8.575 $Y=1.92
c287 146 0 3.07333e-20 $X=7.675 $Y=1.92
c288 141 0 3.07333e-20 $X=6.775 $Y=1.92
c289 132 0 9.40629e-20 $X=12.18 $Y=1.15
c290 53 0 1.0086e-19 $X=5.825 $Y=2.085
c291 51 0 4.00291e-19 $X=5.8 $Y=0.515
r292 170 172 0.769762 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=12.225 $Y=2.035
+ $X2=12.225 $Y2=2.02
r293 170 171 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.2 $Y=2.035
+ $X2=12.2 $Y2=2.035
r294 168 171 0.590276 $w=2.3e-07 $l=9.2e-07 $layer=MET1_cond $X=11.28 $Y=2.035
+ $X2=12.2 $Y2=2.035
r295 165 168 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=2.035
+ $X2=11.28 $Y2=2.035
r296 165 166 4.36643 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=11.275 $Y=2.005
+ $X2=11.275 $Y2=1.92
r297 163 168 0.577444 $w=2.3e-07 $l=9e-07 $layer=MET1_cond $X=10.38 $Y=2.035
+ $X2=11.28 $Y2=2.035
r298 160 163 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.38 $Y=2.035
+ $X2=10.38 $Y2=2.035
r299 160 161 5.17556 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=10.375 $Y=2.005
+ $X2=10.375 $Y2=1.92
r300 158 163 0.571028 $w=2.3e-07 $l=8.9e-07 $layer=MET1_cond $X=9.49 $Y=2.035
+ $X2=10.38 $Y2=2.035
r301 155 158 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.49 $Y=2.035
+ $X2=9.49 $Y2=2.035
r302 155 156 5.66838 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=9.475 $Y=2.005
+ $X2=9.475 $Y2=1.92
r303 150 153 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.57 $Y=2.035
+ $X2=8.57 $Y2=2.035
r304 150 151 5.66838 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=8.575 $Y=2.005
+ $X2=8.575 $Y2=1.92
r305 148 153 0.571028 $w=2.3e-07 $l=8.9e-07 $layer=MET1_cond $X=7.68 $Y=2.035
+ $X2=8.57 $Y2=2.035
r306 145 148 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.68 $Y=2.035
+ $X2=7.68 $Y2=2.035
r307 145 146 5.66838 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=7.675 $Y=2.005
+ $X2=7.675 $Y2=1.92
r308 143 148 0.590276 $w=2.3e-07 $l=9.2e-07 $layer=MET1_cond $X=6.76 $Y=2.035
+ $X2=7.68 $Y2=2.035
r309 140 143 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.76 $Y=2.035
+ $X2=6.76 $Y2=2.035
r310 140 141 5.66838 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=6.775 $Y=2.005
+ $X2=6.775 $Y2=1.92
r311 138 143 0.587068 $w=2.3e-07 $l=9.15e-07 $layer=MET1_cond $X=5.845 $Y=2.035
+ $X2=6.76 $Y2=2.035
r312 136 138 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.845 $Y=2.035
+ $X2=5.845 $Y2=2.035
r313 133 158 0.288722 $w=2.3e-07 $l=4.5e-07 $layer=MET1_cond $X=9.04 $Y=2.035
+ $X2=9.49 $Y2=2.035
r314 133 153 0.301554 $w=2.3e-07 $l=4.7e-07 $layer=MET1_cond $X=9.04 $Y=2.035
+ $X2=8.57 $Y2=2.035
r315 131 161 16.1867 $w=1.83e-07 $l=2.7e-07 $layer=LI1_cond $X=10.302 $Y=1.65
+ $X2=10.302 $Y2=1.92
r316 130 156 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=9.395 $Y=1.65
+ $X2=9.395 $Y2=1.92
r317 129 151 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=8.495 $Y=1.65
+ $X2=8.495 $Y2=1.92
r318 128 146 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=7.595 $Y=1.65
+ $X2=7.595 $Y2=1.92
r319 127 141 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=6.695 $Y=1.65
+ $X2=6.695 $Y2=1.92
r320 123 170 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=12.225 $Y=2.185
+ $X2=12.225 $Y2=2.035
r321 123 125 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=12.225 $Y=2.185
+ $X2=12.225 $Y2=2.4
r322 122 172 1.41528 $w=2.83e-07 $l=3.5e-08 $layer=LI1_cond $X=12.202 $Y=1.985
+ $X2=12.202 $Y2=2.02
r323 122 132 33.7646 $w=2.83e-07 $l=8.35e-07 $layer=LI1_cond $X=12.202 $Y=1.985
+ $X2=12.202 $Y2=1.15
r324 115 132 6.00814 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=12.18 $Y=0.985
+ $X2=12.18 $Y2=1.15
r325 115 117 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=12.18 $Y=0.985
+ $X2=12.18 $Y2=0.515
r326 111 165 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=11.275 $Y=2.085
+ $X2=11.275 $Y2=2.005
r327 111 113 25.4934 $w=3.28e-07 $l=7.3e-07 $layer=LI1_cond $X=11.275 $Y=2.085
+ $X2=11.275 $Y2=2.815
r328 109 166 75.3108 $w=2.13e-07 $l=1.405e-06 $layer=LI1_cond $X=11.217 $Y=0.515
+ $X2=11.217 $Y2=1.92
r329 103 160 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=10.375 $Y=2.085
+ $X2=10.375 $Y2=2.005
r330 103 105 25.4934 $w=3.28e-07 $l=7.3e-07 $layer=LI1_cond $X=10.375 $Y=2.085
+ $X2=10.375 $Y2=2.815
r331 97 131 6.56491 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=10.27 $Y=1.525
+ $X2=10.27 $Y2=1.65
r332 97 99 46.5587 $w=2.48e-07 $l=1.01e-06 $layer=LI1_cond $X=10.27 $Y=1.525
+ $X2=10.27 $Y2=0.515
r333 93 155 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=9.475 $Y=2.085
+ $X2=9.475 $Y2=2.005
r334 93 95 25.4934 $w=3.28e-07 $l=7.3e-07 $layer=LI1_cond $X=9.475 $Y=2.085
+ $X2=9.475 $Y2=2.815
r335 87 130 7.21712 $w=2.63e-07 $l=1.32e-07 $layer=LI1_cond $X=9.347 $Y=1.518
+ $X2=9.347 $Y2=1.65
r336 87 89 43.6189 $w=2.63e-07 $l=1.003e-06 $layer=LI1_cond $X=9.347 $Y=1.518
+ $X2=9.347 $Y2=0.515
r337 83 150 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=8.575 $Y=2.085
+ $X2=8.575 $Y2=2.005
r338 83 85 25.4934 $w=3.28e-07 $l=7.3e-07 $layer=LI1_cond $X=8.575 $Y=2.085
+ $X2=8.575 $Y2=2.815
r339 77 129 7.79447 $w=2.93e-07 $l=1.47e-07 $layer=LI1_cond $X=8.432 $Y=1.503
+ $X2=8.432 $Y2=1.65
r340 77 79 38.5971 $w=2.93e-07 $l=9.88e-07 $layer=LI1_cond $X=8.432 $Y=1.503
+ $X2=8.432 $Y2=0.515
r341 73 145 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=7.675 $Y=2.085
+ $X2=7.675 $Y2=2.005
r342 73 75 25.4934 $w=3.28e-07 $l=7.3e-07 $layer=LI1_cond $X=7.675 $Y=2.085
+ $X2=7.675 $Y2=2.815
r343 67 128 7.79447 $w=2.93e-07 $l=1.47e-07 $layer=LI1_cond $X=7.532 $Y=1.503
+ $X2=7.532 $Y2=1.65
r344 67 69 38.5971 $w=2.93e-07 $l=9.88e-07 $layer=LI1_cond $X=7.532 $Y=1.503
+ $X2=7.532 $Y2=0.515
r345 63 140 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=6.775 $Y=2.085
+ $X2=6.775 $Y2=2.005
r346 63 65 25.4934 $w=3.28e-07 $l=7.3e-07 $layer=LI1_cond $X=6.775 $Y=2.085
+ $X2=6.775 $Y2=2.815
r347 57 127 6.82988 $w=2.43e-07 $l=1.22e-07 $layer=LI1_cond $X=6.657 $Y=1.528
+ $X2=6.657 $Y2=1.65
r348 57 59 47.65 $w=2.43e-07 $l=1.013e-06 $layer=LI1_cond $X=6.657 $Y=1.528
+ $X2=6.657 $Y2=0.515
r349 53 136 2.98307 $w=3.3e-07 $l=8.12404e-08 $layer=LI1_cond $X=5.825 $Y=2.085
+ $X2=5.812 $Y2=2.01
r350 53 55 25.4934 $w=3.28e-07 $l=7.3e-07 $layer=LI1_cond $X=5.825 $Y=2.085
+ $X2=5.825 $Y2=2.815
r351 49 136 10.152 $w=2.9e-07 $l=2.59702e-07 $layer=LI1_cond $X=5.76 $Y=1.775
+ $X2=5.812 $Y2=2.01
r352 49 51 58.0831 $w=2.48e-07 $l=1.26e-06 $layer=LI1_cond $X=5.76 $Y=1.775
+ $X2=5.76 $Y2=0.515
r353 16 125 300 $w=1.7e-07 $l=6.5238e-07 $layer=licon1_PDIFF $count=2 $X=12.025
+ $Y=1.84 $X2=12.225 $Y2=2.4
r354 16 122 600 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=1 $X=12.025
+ $Y=1.84 $X2=12.225 $Y2=1.985
r355 15 165 400 $w=1.7e-07 $l=2.2798e-07 $layer=licon1_PDIFF $count=1 $X=11.125
+ $Y=1.84 $X2=11.275 $Y2=2.005
r356 15 113 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=11.125
+ $Y=1.84 $X2=11.275 $Y2=2.815
r357 14 160 400 $w=1.7e-07 $l=2.2798e-07 $layer=licon1_PDIFF $count=1 $X=10.225
+ $Y=1.84 $X2=10.375 $Y2=2.005
r358 14 105 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=10.225
+ $Y=1.84 $X2=10.375 $Y2=2.815
r359 13 155 400 $w=1.7e-07 $l=2.2798e-07 $layer=licon1_PDIFF $count=1 $X=9.325
+ $Y=1.84 $X2=9.475 $Y2=2.005
r360 13 95 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=9.325
+ $Y=1.84 $X2=9.475 $Y2=2.815
r361 12 150 400 $w=1.7e-07 $l=2.2798e-07 $layer=licon1_PDIFF $count=1 $X=8.425
+ $Y=1.84 $X2=8.575 $Y2=2.005
r362 12 85 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=8.425
+ $Y=1.84 $X2=8.575 $Y2=2.815
r363 11 145 400 $w=1.7e-07 $l=2.2798e-07 $layer=licon1_PDIFF $count=1 $X=7.525
+ $Y=1.84 $X2=7.675 $Y2=2.005
r364 11 75 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=7.525
+ $Y=1.84 $X2=7.675 $Y2=2.815
r365 10 140 400 $w=1.7e-07 $l=2.2798e-07 $layer=licon1_PDIFF $count=1 $X=6.625
+ $Y=1.84 $X2=6.775 $Y2=2.005
r366 10 65 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=6.625
+ $Y=1.84 $X2=6.775 $Y2=2.815
r367 9 136 400 $w=1.7e-07 $l=2.33238e-07 $layer=licon1_PDIFF $count=1 $X=5.675
+ $Y=1.84 $X2=5.825 $Y2=2.01
r368 9 55 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=5.675
+ $Y=1.84 $X2=5.825 $Y2=2.815
r369 8 117 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=12.04
+ $Y=0.37 $X2=12.18 $Y2=0.515
r370 7 109 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=11.1
+ $Y=0.37 $X2=11.24 $Y2=0.515
r371 6 99 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.17
+ $Y=0.37 $X2=10.31 $Y2=0.515
r372 5 89 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.24
+ $Y=0.37 $X2=9.38 $Y2=0.515
r373 4 79 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.31
+ $Y=0.37 $X2=8.45 $Y2=0.515
r374 3 69 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.38
+ $Y=0.37 $X2=7.52 $Y2=0.515
r375 2 59 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.52
+ $Y=0.37 $X2=6.66 $Y2=0.515
r376 1 51 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.66
+ $Y=0.37 $X2=5.8 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__BUFBUF_16%VGND 1 2 3 4 5 6 7 8 9 10 11 12 13 14 45
+ 49 53 57 61 65 69 71 75 77 81 85 89 93 97 99 101 104 105 107 108 110 111 113
+ 114 115 116 118 119 120 122 131 148 153 158 167 172 175 178 181 184 187 190
+ 194
r222 193 194 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r223 190 191 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=0
+ $X2=10.8 $Y2=0
r224 187 188 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0
+ $X2=9.84 $Y2=0
r225 184 185 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r226 181 182 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r227 179 182 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=0
+ $X2=7.92 $Y2=0
r228 178 179 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r229 175 176 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r230 172 173 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0
+ $X2=0.72 $Y2=0
r231 170 194 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=12.72 $Y2=0
r232 169 170 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r233 167 193 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=12.515 $Y=0
+ $X2=12.737 $Y2=0
r234 167 169 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=12.515 $Y=0
+ $X2=12.24 $Y2=0
r235 166 170 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=12.24 $Y2=0
r236 166 191 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=10.8 $Y2=0
r237 165 166 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r238 163 190 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.905 $Y=0
+ $X2=10.74 $Y2=0
r239 163 165 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=10.905 $Y=0
+ $X2=11.28 $Y2=0
r240 162 191 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=10.8 $Y2=0
r241 162 188 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=9.84 $Y2=0
r242 161 162 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r243 159 187 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=9.975 $Y=0
+ $X2=9.82 $Y2=0
r244 159 161 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=9.975 $Y=0
+ $X2=10.32 $Y2=0
r245 158 190 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.575 $Y=0
+ $X2=10.74 $Y2=0
r246 158 161 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=10.575 $Y=0
+ $X2=10.32 $Y2=0
r247 157 188 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=9.84 $Y2=0
r248 157 185 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=8.88 $Y2=0
r249 156 157 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r250 154 184 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=9.045 $Y=0
+ $X2=8.897 $Y2=0
r251 154 156 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=9.045 $Y=0
+ $X2=9.36 $Y2=0
r252 153 187 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=9.665 $Y=0
+ $X2=9.82 $Y2=0
r253 153 156 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=9.665 $Y=0
+ $X2=9.36 $Y2=0
r254 152 185 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0
+ $X2=8.88 $Y2=0
r255 152 182 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0
+ $X2=7.92 $Y2=0
r256 151 152 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r257 149 181 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=8.115 $Y=0
+ $X2=7.982 $Y2=0
r258 149 151 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=8.115 $Y=0
+ $X2=8.4 $Y2=0
r259 148 184 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=8.75 $Y=0
+ $X2=8.897 $Y2=0
r260 148 151 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=8.75 $Y=0 $X2=8.4
+ $Y2=0
r261 146 147 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6
+ $Y2=0
r262 144 147 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=6
+ $Y2=0
r263 143 144 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r264 141 144 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0
+ $X2=5.04 $Y2=0
r265 140 141 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r266 138 141 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0
+ $X2=4.08 $Y2=0
r267 138 176 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0
+ $X2=2.64 $Y2=0
r268 137 138 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r269 135 175 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.745 $Y=0
+ $X2=2.58 $Y2=0
r270 135 137 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=2.745 $Y=0
+ $X2=3.12 $Y2=0
r271 134 176 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=2.64 $Y2=0
r272 133 134 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r273 131 175 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.415 $Y=0
+ $X2=2.58 $Y2=0
r274 131 133 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.415 $Y=0
+ $X2=2.16 $Y2=0
r275 130 134 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0
+ $X2=2.16 $Y2=0
r276 130 173 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0
+ $X2=0.72 $Y2=0
r277 129 130 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r278 127 172 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.89 $Y=0
+ $X2=0.725 $Y2=0
r279 127 129 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.89 $Y=0 $X2=1.2
+ $Y2=0
r280 125 173 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0
+ $X2=0.72 $Y2=0
r281 124 125 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r282 122 172 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.56 $Y=0
+ $X2=0.725 $Y2=0
r283 122 124 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.56 $Y=0 $X2=0.24
+ $Y2=0
r284 120 179 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0
+ $X2=6.96 $Y2=0
r285 120 147 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r286 118 165 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=11.505 $Y=0
+ $X2=11.28 $Y2=0
r287 118 119 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.505 $Y=0
+ $X2=11.67 $Y2=0
r288 117 169 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=11.835 $Y=0
+ $X2=12.24 $Y2=0
r289 117 119 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.835 $Y=0
+ $X2=11.67 $Y2=0
r290 115 146 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=6.065 $Y=0 $X2=6
+ $Y2=0
r291 115 116 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.065 $Y=0
+ $X2=6.19 $Y2=0
r292 113 143 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=5.275 $Y=0
+ $X2=5.04 $Y2=0
r293 113 114 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=5.275 $Y=0 $X2=5.365
+ $Y2=0
r294 112 146 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=5.455 $Y=0 $X2=6
+ $Y2=0
r295 112 114 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=5.455 $Y=0 $X2=5.365
+ $Y2=0
r296 110 140 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=4.275 $Y=0
+ $X2=4.08 $Y2=0
r297 110 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.275 $Y=0
+ $X2=4.44 $Y2=0
r298 109 143 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=4.605 $Y=0
+ $X2=5.04 $Y2=0
r299 109 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.605 $Y=0
+ $X2=4.44 $Y2=0
r300 107 137 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=3.345 $Y=0
+ $X2=3.12 $Y2=0
r301 107 108 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.345 $Y=0
+ $X2=3.51 $Y2=0
r302 106 140 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=3.675 $Y=0
+ $X2=4.08 $Y2=0
r303 106 108 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.675 $Y=0
+ $X2=3.51 $Y2=0
r304 104 129 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=1.42 $Y=0 $X2=1.2
+ $Y2=0
r305 104 105 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.42 $Y=0
+ $X2=1.545 $Y2=0
r306 103 133 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=1.67 $Y=0
+ $X2=2.16 $Y2=0
r307 103 105 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.67 $Y=0
+ $X2=1.545 $Y2=0
r308 99 193 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=12.68 $Y=0.085
+ $X2=12.737 $Y2=0
r309 99 101 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=12.68 $Y=0.085
+ $X2=12.68 $Y2=0.515
r310 95 119 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.67 $Y=0.085
+ $X2=11.67 $Y2=0
r311 95 97 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=11.67 $Y=0.085
+ $X2=11.67 $Y2=0.515
r312 91 190 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.74 $Y=0.085
+ $X2=10.74 $Y2=0
r313 91 93 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=10.74 $Y=0.085
+ $X2=10.74 $Y2=0.515
r314 87 187 0.701276 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=9.82 $Y=0.085
+ $X2=9.82 $Y2=0
r315 87 89 15.9855 $w=3.08e-07 $l=4.3e-07 $layer=LI1_cond $X=9.82 $Y=0.085
+ $X2=9.82 $Y2=0.515
r316 83 184 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=8.897 $Y=0.085
+ $X2=8.897 $Y2=0
r317 83 85 16.7983 $w=2.93e-07 $l=4.3e-07 $layer=LI1_cond $X=8.897 $Y=0.085
+ $X2=8.897 $Y2=0.515
r318 79 181 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=7.982 $Y=0.085
+ $X2=7.982 $Y2=0
r319 79 81 18.7 $w=2.63e-07 $l=4.3e-07 $layer=LI1_cond $X=7.982 $Y=0.085
+ $X2=7.982 $Y2=0.515
r320 78 178 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=7.175 $Y=0
+ $X2=7.067 $Y2=0
r321 77 181 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=7.85 $Y=0
+ $X2=7.982 $Y2=0
r322 77 78 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=7.85 $Y=0
+ $X2=7.175 $Y2=0
r323 73 178 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=7.067 $Y=0.085
+ $X2=7.067 $Y2=0
r324 73 75 23.0489 $w=2.13e-07 $l=4.3e-07 $layer=LI1_cond $X=7.067 $Y=0.085
+ $X2=7.067 $Y2=0.515
r325 72 116 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.315 $Y=0
+ $X2=6.19 $Y2=0
r326 71 178 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=6.96 $Y=0
+ $X2=7.067 $Y2=0
r327 71 72 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=6.96 $Y=0
+ $X2=6.315 $Y2=0
r328 67 116 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.19 $Y=0.085
+ $X2=6.19 $Y2=0
r329 67 69 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=6.19 $Y=0.085
+ $X2=6.19 $Y2=0.515
r330 63 114 1.13756 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=5.365 $Y=0.085
+ $X2=5.365 $Y2=0
r331 63 65 30.5 $w=1.78e-07 $l=4.95e-07 $layer=LI1_cond $X=5.365 $Y=0.085
+ $X2=5.365 $Y2=0.58
r332 59 111 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.44 $Y=0.085
+ $X2=4.44 $Y2=0
r333 59 61 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=4.44 $Y=0.085
+ $X2=4.44 $Y2=0.645
r334 55 108 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.51 $Y=0.085
+ $X2=3.51 $Y2=0
r335 55 57 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=3.51 $Y=0.085
+ $X2=3.51 $Y2=0.645
r336 51 175 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.58 $Y=0.085
+ $X2=2.58 $Y2=0
r337 51 53 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.58 $Y=0.085
+ $X2=2.58 $Y2=0.515
r338 47 105 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.545 $Y=0.085
+ $X2=1.545 $Y2=0
r339 47 49 24.8928 $w=2.48e-07 $l=5.4e-07 $layer=LI1_cond $X=1.545 $Y=0.085
+ $X2=1.545 $Y2=0.625
r340 43 172 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.725 $Y=0.085
+ $X2=0.725 $Y2=0
r341 43 45 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=0.725 $Y=0.085
+ $X2=0.725 $Y2=0.625
r342 14 101 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=12.47
+ $Y=0.37 $X2=12.68 $Y2=0.515
r343 13 97 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=11.53
+ $Y=0.37 $X2=11.67 $Y2=0.515
r344 12 93 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.6
+ $Y=0.37 $X2=10.74 $Y2=0.515
r345 11 89 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.67
+ $Y=0.37 $X2=9.81 $Y2=0.515
r346 10 85 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.74
+ $Y=0.37 $X2=8.88 $Y2=0.515
r347 9 81 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.81
+ $Y=0.37 $X2=7.95 $Y2=0.515
r348 8 75 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.95
+ $Y=0.37 $X2=7.09 $Y2=0.515
r349 7 69 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.09
+ $Y=0.37 $X2=6.23 $Y2=0.515
r350 6 65 91 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=2 $X=5.23
+ $Y=0.37 $X2=5.37 $Y2=0.58
r351 5 61 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=4.3
+ $Y=0.37 $X2=4.44 $Y2=0.645
r352 4 57 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=3.37
+ $Y=0.37 $X2=3.51 $Y2=0.645
r353 3 53 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=2.435
+ $Y=0.37 $X2=2.58 $Y2=0.515
r354 2 49 182 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=1 $X=1.445
+ $Y=0.37 $X2=1.585 $Y2=0.625
r355 1 45 182 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=1 $X=0.585
+ $Y=0.37 $X2=0.725 $Y2=0.625
.ends

