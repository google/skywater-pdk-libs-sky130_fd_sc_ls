* File: sky130_fd_sc_ls__decaphe_4.pxi.spice
* Created: Wed Sep  2 10:59:54 2020
* 
x_PM_SKY130_FD_SC_LS__DECAPHE_4%VGND N_VGND_M1000_s N_VGND_M1001_g VGND
+ N_VGND_c_12_n N_VGND_c_13_n N_VGND_c_14_n PM_SKY130_FD_SC_LS__DECAPHE_4%VGND
x_PM_SKY130_FD_SC_LS__DECAPHE_4%VPWR N_VPWR_M1001_s N_VPWR_M1000_g N_VPWR_c_26_n
+ VPWR N_VPWR_c_28_n N_VPWR_c_29_n VPWR PM_SKY130_FD_SC_LS__DECAPHE_4%VPWR
cc_1 VNB N_VGND_c_12_n 0.0323905f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=1.515
cc_2 VNB N_VGND_c_13_n 0.12642f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=0
cc_3 VNB N_VGND_c_14_n 0.146162f $X=-0.19 $Y=-0.245 $X2=0.26 $Y2=0.38
cc_4 VNB N_VPWR_c_26_n 0.0950012f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=1.71
cc_5 VNB VPWR 0.0840719f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_VPWR_c_28_n 0.0374636f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=1.515
cc_7 VNB N_VPWR_c_29_n 0.0257206f $X=-0.19 $Y=-0.245 $X2=1.66 $Y2=0.38
cc_8 VPB N_VGND_M1001_g 0.0950353f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=2.467
cc_9 VPB N_VGND_c_12_n 0.00562362f $X=-0.19 $Y=1.66 $X2=0.575 $Y2=1.515
cc_10 VPB VPWR 0.0423484f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_11 VPB N_VPWR_c_29_n 0.161239f $X=-0.19 $Y=1.66 $X2=1.66 $Y2=0.38
cc_12 N_VGND_M1001_g N_VPWR_c_26_n 0.00784274f $X=0.96 $Y=2.467 $X2=0 $Y2=0
cc_13 N_VGND_c_12_n N_VPWR_c_26_n 0.0225662f $X=0.575 $Y=1.515 $X2=0 $Y2=0
cc_14 N_VGND_c_14_n N_VPWR_c_26_n 0.157908f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_15 N_VGND_M1001_g N_VPWR_c_28_n 0.0219121f $X=0.96 $Y=2.467 $X2=0 $Y2=0
cc_16 N_VGND_c_12_n N_VPWR_c_28_n 0.00347831f $X=0.575 $Y=1.515 $X2=0 $Y2=0
cc_17 N_VGND_c_14_n N_VPWR_c_28_n 0.00531025f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_18 N_VGND_M1001_g N_VPWR_c_29_n 0.212228f $X=0.96 $Y=2.467 $X2=0 $Y2=0
cc_19 N_VGND_c_12_n N_VPWR_c_29_n 0.00518926f $X=0.575 $Y=1.515 $X2=0 $Y2=0
cc_20 N_VGND_c_14_n N_VPWR_c_29_n 0.173407f $X=0.26 $Y=0.38 $X2=0 $Y2=0
