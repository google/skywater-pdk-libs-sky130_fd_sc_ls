* File: sky130_fd_sc_ls__dlrbp_2.pxi.spice
* Created: Wed Sep  2 11:03:31 2020
* 
x_PM_SKY130_FD_SC_LS__DLRBP_2%D N_D_M1012_g N_D_c_173_n N_D_M1019_g D
+ PM_SKY130_FD_SC_LS__DLRBP_2%D
x_PM_SKY130_FD_SC_LS__DLRBP_2%GATE N_GATE_M1009_g N_GATE_c_208_n N_GATE_c_213_n
+ N_GATE_M1015_g GATE N_GATE_c_210_n N_GATE_c_211_n
+ PM_SKY130_FD_SC_LS__DLRBP_2%GATE
x_PM_SKY130_FD_SC_LS__DLRBP_2%A_230_74# N_A_230_74#_M1009_d N_A_230_74#_M1015_d
+ N_A_230_74#_c_248_n N_A_230_74#_c_249_n N_A_230_74#_c_250_n
+ N_A_230_74#_c_251_n N_A_230_74#_M1000_g N_A_230_74#_c_262_n
+ N_A_230_74#_M1025_g N_A_230_74#_c_263_n N_A_230_74#_M1010_g
+ N_A_230_74#_c_264_n N_A_230_74#_c_265_n N_A_230_74#_M1001_g
+ N_A_230_74#_c_267_n N_A_230_74#_c_253_n N_A_230_74#_c_254_n
+ N_A_230_74#_c_255_n N_A_230_74#_c_256_n N_A_230_74#_c_257_n
+ N_A_230_74#_c_268_n N_A_230_74#_c_258_n N_A_230_74#_c_259_n
+ N_A_230_74#_c_260_n PM_SKY130_FD_SC_LS__DLRBP_2%A_230_74#
x_PM_SKY130_FD_SC_LS__DLRBP_2%A_27_112# N_A_27_112#_M1012_s N_A_27_112#_M1019_s
+ N_A_27_112#_c_389_n N_A_27_112#_M1016_g N_A_27_112#_M1002_g
+ N_A_27_112#_c_391_n N_A_27_112#_c_396_n N_A_27_112#_c_397_n
+ N_A_27_112#_c_398_n N_A_27_112#_c_392_n N_A_27_112#_c_393_n
+ N_A_27_112#_c_400_n N_A_27_112#_c_394_n PM_SKY130_FD_SC_LS__DLRBP_2%A_27_112#
x_PM_SKY130_FD_SC_LS__DLRBP_2%A_363_82# N_A_363_82#_M1000_s N_A_363_82#_M1025_s
+ N_A_363_82#_M1022_g N_A_363_82#_c_478_n N_A_363_82#_M1020_g
+ N_A_363_82#_c_471_n N_A_363_82#_c_472_n N_A_363_82#_c_473_n
+ N_A_363_82#_c_474_n N_A_363_82#_c_481_n N_A_363_82#_c_482_n
+ N_A_363_82#_c_483_n N_A_363_82#_c_484_n N_A_363_82#_c_475_n
+ N_A_363_82#_c_476_n N_A_363_82#_c_477_n PM_SKY130_FD_SC_LS__DLRBP_2%A_363_82#
x_PM_SKY130_FD_SC_LS__DLRBP_2%A_821_98# N_A_821_98#_M1013_s N_A_821_98#_M1027_d
+ N_A_821_98#_c_587_n N_A_821_98#_M1017_g N_A_821_98#_c_588_n
+ N_A_821_98#_c_601_n N_A_821_98#_M1021_g N_A_821_98#_M1023_g
+ N_A_821_98#_c_602_n N_A_821_98#_M1003_g N_A_821_98#_M1024_g
+ N_A_821_98#_c_603_n N_A_821_98#_M1026_g N_A_821_98#_c_591_n
+ N_A_821_98#_c_592_n N_A_821_98#_c_605_n N_A_821_98#_M1008_g
+ N_A_821_98#_M1004_g N_A_821_98#_c_594_n N_A_821_98#_c_595_n
+ N_A_821_98#_c_607_n N_A_821_98#_c_596_n N_A_821_98#_c_608_n
+ N_A_821_98#_c_609_n N_A_821_98#_c_597_n N_A_821_98#_c_707_p
+ N_A_821_98#_c_598_n N_A_821_98#_c_611_n N_A_821_98#_c_599_n
+ PM_SKY130_FD_SC_LS__DLRBP_2%A_821_98#
x_PM_SKY130_FD_SC_LS__DLRBP_2%A_641_80# N_A_641_80#_M1022_d N_A_641_80#_M1010_d
+ N_A_641_80#_c_746_n N_A_641_80#_M1027_g N_A_641_80#_M1013_g
+ N_A_641_80#_c_748_n N_A_641_80#_c_760_n N_A_641_80#_c_755_n
+ N_A_641_80#_c_749_n N_A_641_80#_c_750_n N_A_641_80#_c_751_n
+ N_A_641_80#_c_752_n PM_SKY130_FD_SC_LS__DLRBP_2%A_641_80#
x_PM_SKY130_FD_SC_LS__DLRBP_2%RESET_B N_RESET_B_c_829_n N_RESET_B_M1006_g
+ N_RESET_B_c_830_n N_RESET_B_M1005_g RESET_B N_RESET_B_c_831_n
+ PM_SKY130_FD_SC_LS__DLRBP_2%RESET_B
x_PM_SKY130_FD_SC_LS__DLRBP_2%A_1449_368# N_A_1449_368#_M1004_s
+ N_A_1449_368#_M1008_s N_A_1449_368#_c_871_n N_A_1449_368#_M1011_g
+ N_A_1449_368#_M1007_g N_A_1449_368#_c_872_n N_A_1449_368#_M1018_g
+ N_A_1449_368#_M1014_g N_A_1449_368#_c_865_n N_A_1449_368#_c_866_n
+ N_A_1449_368#_c_867_n N_A_1449_368#_c_868_n N_A_1449_368#_c_869_n
+ N_A_1449_368#_c_885_n N_A_1449_368#_c_870_n
+ PM_SKY130_FD_SC_LS__DLRBP_2%A_1449_368#
x_PM_SKY130_FD_SC_LS__DLRBP_2%VPWR N_VPWR_M1019_d N_VPWR_M1025_d N_VPWR_M1021_d
+ N_VPWR_M1005_d N_VPWR_M1026_d N_VPWR_M1008_d N_VPWR_M1018_s N_VPWR_c_934_n
+ N_VPWR_c_935_n N_VPWR_c_936_n N_VPWR_c_937_n N_VPWR_c_938_n N_VPWR_c_939_n
+ N_VPWR_c_940_n N_VPWR_c_941_n N_VPWR_c_942_n N_VPWR_c_943_n N_VPWR_c_944_n
+ VPWR N_VPWR_c_945_n N_VPWR_c_946_n N_VPWR_c_947_n N_VPWR_c_948_n
+ N_VPWR_c_949_n N_VPWR_c_950_n N_VPWR_c_951_n N_VPWR_c_952_n N_VPWR_c_933_n
+ PM_SKY130_FD_SC_LS__DLRBP_2%VPWR
x_PM_SKY130_FD_SC_LS__DLRBP_2%Q N_Q_M1023_d N_Q_M1003_s N_Q_c_1047_n
+ N_Q_c_1051_n N_Q_c_1052_n N_Q_c_1053_n N_Q_c_1048_n N_Q_c_1049_n Q
+ PM_SKY130_FD_SC_LS__DLRBP_2%Q
x_PM_SKY130_FD_SC_LS__DLRBP_2%Q_N N_Q_N_M1007_d N_Q_N_M1011_d N_Q_N_c_1102_n
+ N_Q_N_c_1103_n Q_N Q_N N_Q_N_c_1104_n PM_SKY130_FD_SC_LS__DLRBP_2%Q_N
x_PM_SKY130_FD_SC_LS__DLRBP_2%VGND N_VGND_M1012_d N_VGND_M1000_d N_VGND_M1017_d
+ N_VGND_M1006_d N_VGND_M1024_s N_VGND_M1004_d N_VGND_M1014_s N_VGND_c_1132_n
+ N_VGND_c_1133_n N_VGND_c_1134_n N_VGND_c_1135_n N_VGND_c_1136_n
+ N_VGND_c_1137_n N_VGND_c_1138_n N_VGND_c_1139_n N_VGND_c_1140_n
+ N_VGND_c_1141_n N_VGND_c_1142_n N_VGND_c_1143_n N_VGND_c_1144_n
+ N_VGND_c_1145_n VGND N_VGND_c_1146_n N_VGND_c_1147_n N_VGND_c_1148_n
+ N_VGND_c_1149_n N_VGND_c_1150_n N_VGND_c_1151_n
+ PM_SKY130_FD_SC_LS__DLRBP_2%VGND
cc_1 VNB N_D_M1012_g 0.0375151f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.835
cc_2 VNB N_D_c_173_n 0.0219514f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.885
cc_3 VNB D 0.00242107f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_4 VNB N_GATE_c_208_n 0.00639429f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.885
cc_5 VNB GATE 0.0061593f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_GATE_c_210_n 0.0351696f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.615
cc_7 VNB N_GATE_c_211_n 0.0226366f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_230_74#_c_248_n 0.0153485f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.38
cc_9 VNB N_A_230_74#_c_249_n 0.0150746f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_230_74#_c_250_n 0.00785243f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.615
cc_11 VNB N_A_230_74#_c_251_n 0.0187611f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.615
cc_12 VNB N_A_230_74#_M1001_g 0.0417255f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_230_74#_c_253_n 0.00580127f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_230_74#_c_254_n 0.00163151f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_230_74#_c_255_n 0.00874055f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_230_74#_c_256_n 0.0446354f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_230_74#_c_257_n 0.0163502f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_230_74#_c_258_n 0.00543595f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_230_74#_c_259_n 0.00643839f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_230_74#_c_260_n 0.0272613f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_27_112#_c_389_n 0.020867f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.38
cc_22 VNB N_A_27_112#_M1002_g 0.0326722f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.615
cc_23 VNB N_A_27_112#_c_391_n 0.0201039f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_27_112#_c_392_n 0.00196261f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_27_112#_c_393_n 0.013652f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_27_112#_c_394_n 0.0253939f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_363_82#_c_471_n 0.00623344f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.615
cc_28 VNB N_A_363_82#_c_472_n 0.00153466f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_363_82#_c_473_n 0.0177304f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.615
cc_30 VNB N_A_363_82#_c_474_n 0.00287888f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_363_82#_c_475_n 0.00746834f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_363_82#_c_476_n 0.0308969f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_363_82#_c_477_n 0.0159056f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_821_98#_c_587_n 0.0171346f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.38
cc_35 VNB N_A_821_98#_c_588_n 0.0227549f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.615
cc_36 VNB N_A_821_98#_M1023_g 0.0223246f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_821_98#_M1024_g 0.0227941f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_821_98#_c_591_n 0.0808111f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_821_98#_c_592_n 0.0426054f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_821_98#_M1004_g 0.0259366f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_821_98#_c_594_n 0.0198739f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_821_98#_c_595_n 0.0119774f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_821_98#_c_596_n 0.00813778f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_821_98#_c_597_n 0.00536874f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_821_98#_c_598_n 0.00577602f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_821_98#_c_599_n 0.00387127f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_641_80#_c_746_n 0.012578f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.38
cc_48 VNB N_A_641_80#_M1013_g 0.0266521f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.615
cc_49 VNB N_A_641_80#_c_748_n 0.0311649f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.615
cc_50 VNB N_A_641_80#_c_749_n 0.00574196f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_641_80#_c_750_n 0.0140086f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_641_80#_c_751_n 0.007314f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_641_80#_c_752_n 0.00856244f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_RESET_B_c_829_n 0.0172008f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.45
cc_55 VNB N_RESET_B_c_830_n 0.0342434f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_RESET_B_c_831_n 0.00860315f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.615
cc_57 VNB N_A_1449_368#_M1007_g 0.0229007f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.615
cc_58 VNB N_A_1449_368#_M1014_g 0.0260184f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_1449_368#_c_865_n 0.00924021f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_1449_368#_c_866_n 0.00129392f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_1449_368#_c_867_n 2.15008e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_1449_368#_c_868_n 0.00569931f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_1449_368#_c_869_n 0.00140993f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_1449_368#_c_870_n 0.0742336f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VPWR_c_933_n 0.382608f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_Q_c_1047_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_Q_c_1048_n 0.00849508f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_Q_c_1049_n 0.00230427f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB Q 0.00348326f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_Q_N_c_1102_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_Q_N_c_1103_n 0.00429087f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.615
cc_72 VNB N_Q_N_c_1104_n 0.00141953f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1132_n 0.0168478f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1133_n 0.0219756f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1134_n 0.00650187f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1135_n 0.0171896f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1136_n 0.0166669f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1137_n 0.010678f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1138_n 0.0505285f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1139_n 0.0514319f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1140_n 0.0393212f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1141_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1142_n 0.0294964f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1143_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1144_n 0.0199677f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1145_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1146_n 0.020108f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1147_n 0.0221748f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1148_n 0.0189349f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1149_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_VGND_c_1150_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_VGND_c_1151_n 0.519539f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VPB N_D_c_173_n 0.0431196f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.885
cc_94 VPB D 0.00201744f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_95 VPB N_GATE_c_208_n 0.00832545f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.885
cc_96 VPB N_GATE_c_213_n 0.0275386f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.38
cc_97 VPB N_A_230_74#_c_250_n 0.00840691f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.615
cc_98 VPB N_A_230_74#_c_262_n 0.0277505f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB N_A_230_74#_c_263_n 0.0148583f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 VPB N_A_230_74#_c_264_n 0.0407751f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB N_A_230_74#_c_265_n 0.0107396f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_102 VPB N_A_230_74#_M1001_g 0.00178447f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 VPB N_A_230_74#_c_267_n 0.00639058f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB N_A_230_74#_c_268_n 0.0104636f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_105 VPB N_A_230_74#_c_258_n 0.007206f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_A_230_74#_c_260_n 0.0100279f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB N_A_27_112#_c_389_n 0.0382768f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.38
cc_108 VPB N_A_27_112#_c_396_n 0.00900146f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_109 VPB N_A_27_112#_c_397_n 0.0094938f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_110 VPB N_A_27_112#_c_398_n 0.0226171f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_A_27_112#_c_392_n 0.0011664f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_A_27_112#_c_400_n 0.0138013f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_A_27_112#_c_394_n 0.0138058f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_A_363_82#_c_478_n 0.0646292f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.615
cc_115 VPB N_A_363_82#_c_472_n 0.00382513f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_A_363_82#_c_474_n 0.00199723f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_A_363_82#_c_481_n 0.00595538f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_A_363_82#_c_482_n 0.00172818f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_A_363_82#_c_483_n 0.00463593f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_A_363_82#_c_484_n 0.00518455f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_A_821_98#_c_588_n 0.0240193f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.615
cc_122 VPB N_A_821_98#_c_601_n 0.061562f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.615
cc_123 VPB N_A_821_98#_c_602_n 0.0161151f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_A_821_98#_c_603_n 0.017277f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_A_821_98#_c_592_n 0.013608f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 VPB N_A_821_98#_c_605_n 0.0179607f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_127 VPB N_A_821_98#_c_595_n 0.00862332f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_A_821_98#_c_607_n 0.0085437f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_129 VPB N_A_821_98#_c_608_n 0.00289722f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_A_821_98#_c_609_n 0.00648491f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_A_821_98#_c_597_n 8.46891e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_A_821_98#_c_611_n 0.00760266f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_A_821_98#_c_599_n 6.12609e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_A_641_80#_c_746_n 0.0239864f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.38
cc_135 VPB N_A_641_80#_c_748_n 0.013129f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.615
cc_136 VPB N_A_641_80#_c_755_n 0.00481761f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_A_641_80#_c_750_n 0.0101815f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_A_641_80#_c_751_n 2.16397e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_A_641_80#_c_752_n 0.00406817f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_140 VPB N_RESET_B_c_830_n 0.0230301f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_141 VPB N_A_1449_368#_c_871_n 0.0163314f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.38
cc_142 VPB N_A_1449_368#_c_872_n 0.017357f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_143 VPB N_A_1449_368#_c_867_n 0.00476876f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_144 VPB N_A_1449_368#_c_870_n 0.016936f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_145 VPB N_VPWR_c_934_n 0.0212796f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_146 VPB N_VPWR_c_935_n 0.0130706f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_147 VPB N_VPWR_c_936_n 0.00823722f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_148 VPB N_VPWR_c_937_n 0.0174685f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_149 VPB N_VPWR_c_938_n 0.0176636f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_150 VPB N_VPWR_c_939_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_151 VPB N_VPWR_c_940_n 0.0644986f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_152 VPB N_VPWR_c_941_n 0.0185677f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_153 VPB N_VPWR_c_942_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_154 VPB N_VPWR_c_943_n 0.0175592f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_155 VPB N_VPWR_c_944_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_156 VPB N_VPWR_c_945_n 0.0428961f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_157 VPB N_VPWR_c_946_n 0.0443982f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_158 VPB N_VPWR_c_947_n 0.0212658f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_159 VPB N_VPWR_c_948_n 0.0194151f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_160 VPB N_VPWR_c_949_n 0.0270908f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_161 VPB N_VPWR_c_950_n 0.00681636f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_162 VPB N_VPWR_c_951_n 0.0180078f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_163 VPB N_VPWR_c_952_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_164 VPB N_VPWR_c_933_n 0.126582f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_165 VPB N_Q_c_1051_n 0.0018149f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.615
cc_166 VPB N_Q_c_1052_n 0.00722366f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_167 VPB N_Q_c_1053_n 0.00133363f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_168 VPB Q 0.00234812f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_169 VPB Q_N 0.00198321f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_170 VPB Q_N 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_171 VPB N_Q_N_c_1104_n 0.00104928f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_172 N_D_c_173_n N_GATE_c_208_n 0.013221f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_173 D N_GATE_c_208_n 0.00243125f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_174 N_D_c_173_n N_GATE_c_213_n 0.0237484f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_175 N_D_M1012_g GATE 0.00204708f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_176 D GATE 0.00792655f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_177 N_D_M1012_g N_GATE_c_210_n 0.00769876f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_178 N_D_c_173_n N_GATE_c_210_n 0.0062543f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_179 D N_GATE_c_210_n 5.77592e-19 $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_180 N_D_M1012_g N_GATE_c_211_n 0.0167806f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_181 N_D_c_173_n N_A_230_74#_c_268_n 0.00108229f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_182 D N_A_230_74#_c_258_n 0.00736576f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_183 N_D_M1012_g N_A_27_112#_c_391_n 0.00673958f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_184 N_D_c_173_n N_A_27_112#_c_396_n 0.0057145f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_185 N_D_c_173_n N_A_27_112#_c_397_n 0.0139311f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_186 D N_A_27_112#_c_397_n 0.00920867f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_187 N_D_c_173_n N_A_27_112#_c_398_n 0.00769688f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_188 N_D_M1012_g N_A_27_112#_c_393_n 0.00583243f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_189 D N_A_27_112#_c_393_n 9.01811e-19 $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_190 N_D_c_173_n N_A_27_112#_c_400_n 0.00477742f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_191 D N_A_27_112#_c_400_n 0.00153915f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_192 N_D_M1012_g N_A_27_112#_c_394_n 0.00927701f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_193 N_D_c_173_n N_A_27_112#_c_394_n 0.0117627f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_194 D N_A_27_112#_c_394_n 0.0250412f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_195 N_D_c_173_n N_VPWR_c_934_n 0.0043785f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_196 N_D_c_173_n N_VPWR_c_949_n 0.00457243f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_197 N_D_c_173_n N_VPWR_c_933_n 0.0049649f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_198 N_D_M1012_g N_VGND_c_1132_n 0.00610345f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_199 N_D_c_173_n N_VGND_c_1132_n 0.00252403f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_200 D N_VGND_c_1132_n 0.00727791f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_201 N_D_M1012_g N_VGND_c_1146_n 0.0043356f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_202 N_D_M1012_g N_VGND_c_1151_n 0.00487769f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_203 N_GATE_c_213_n N_A_230_74#_c_267_n 0.00528874f $X=1.125 $Y=1.885 $X2=0
+ $Y2=0
cc_204 GATE N_A_230_74#_c_257_n 0.0110796f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_205 N_GATE_c_210_n N_A_230_74#_c_257_n 0.00124558f $X=1.13 $Y=1.385 $X2=0
+ $Y2=0
cc_206 N_GATE_c_211_n N_A_230_74#_c_257_n 0.0080587f $X=1.13 $Y=1.22 $X2=0 $Y2=0
cc_207 N_GATE_c_213_n N_A_230_74#_c_268_n 0.00665365f $X=1.125 $Y=1.885 $X2=0
+ $Y2=0
cc_208 GATE N_A_230_74#_c_268_n 0.00411005f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_209 N_GATE_c_210_n N_A_230_74#_c_268_n 7.65906e-19 $X=1.13 $Y=1.385 $X2=0
+ $Y2=0
cc_210 N_GATE_c_208_n N_A_230_74#_c_258_n 0.00358524f $X=1.125 $Y=1.795 $X2=0
+ $Y2=0
cc_211 GATE N_A_230_74#_c_259_n 0.0289292f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_212 N_GATE_c_210_n N_A_230_74#_c_259_n 0.00404058f $X=1.13 $Y=1.385 $X2=0
+ $Y2=0
cc_213 N_GATE_c_211_n N_A_230_74#_c_259_n 0.00376199f $X=1.13 $Y=1.22 $X2=0
+ $Y2=0
cc_214 N_GATE_c_208_n N_A_230_74#_c_260_n 0.00418042f $X=1.125 $Y=1.795 $X2=0
+ $Y2=0
cc_215 GATE N_A_230_74#_c_260_n 2.22836e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_216 N_GATE_c_210_n N_A_230_74#_c_260_n 0.0110794f $X=1.13 $Y=1.385 $X2=0
+ $Y2=0
cc_217 N_GATE_c_211_n N_A_27_112#_c_391_n 6.40098e-19 $X=1.13 $Y=1.22 $X2=0
+ $Y2=0
cc_218 N_GATE_c_213_n N_A_27_112#_c_397_n 0.0186743f $X=1.125 $Y=1.885 $X2=0
+ $Y2=0
cc_219 N_GATE_c_213_n N_A_27_112#_c_398_n 7.68188e-19 $X=1.125 $Y=1.885 $X2=0
+ $Y2=0
cc_220 N_GATE_c_213_n N_A_27_112#_c_400_n 0.00178664f $X=1.125 $Y=1.885 $X2=0
+ $Y2=0
cc_221 N_GATE_c_213_n N_A_363_82#_c_484_n 3.43801e-19 $X=1.125 $Y=1.885 $X2=0
+ $Y2=0
cc_222 N_GATE_c_213_n N_VPWR_c_934_n 0.00663705f $X=1.125 $Y=1.885 $X2=0 $Y2=0
cc_223 N_GATE_c_213_n N_VPWR_c_945_n 0.00469064f $X=1.125 $Y=1.885 $X2=0 $Y2=0
cc_224 N_GATE_c_213_n N_VPWR_c_933_n 0.0049649f $X=1.125 $Y=1.885 $X2=0 $Y2=0
cc_225 N_GATE_c_211_n N_VGND_c_1132_n 0.00984417f $X=1.13 $Y=1.22 $X2=0 $Y2=0
cc_226 N_GATE_c_211_n N_VGND_c_1139_n 0.00434272f $X=1.13 $Y=1.22 $X2=0 $Y2=0
cc_227 N_GATE_c_211_n N_VGND_c_1151_n 0.00830058f $X=1.13 $Y=1.22 $X2=0 $Y2=0
cc_228 N_A_230_74#_c_249_n N_A_27_112#_c_389_n 0.0196982f $X=2.185 $Y=1.49 $X2=0
+ $Y2=0
cc_229 N_A_230_74#_c_262_n N_A_27_112#_c_389_n 0.0237573f $X=2.185 $Y=1.885
+ $X2=0 $Y2=0
cc_230 N_A_230_74#_c_263_n N_A_27_112#_c_389_n 0.0511533f $X=3.175 $Y=1.885
+ $X2=0 $Y2=0
cc_231 N_A_230_74#_c_265_n N_A_27_112#_c_389_n 0.0100872f $X=3.265 $Y=1.765
+ $X2=0 $Y2=0
cc_232 N_A_230_74#_c_249_n N_A_27_112#_M1002_g 0.00760431f $X=2.185 $Y=1.49
+ $X2=0 $Y2=0
cc_233 N_A_230_74#_c_251_n N_A_27_112#_M1002_g 0.0247978f $X=2.175 $Y=1.225
+ $X2=0 $Y2=0
cc_234 N_A_230_74#_c_253_n N_A_27_112#_M1002_g 0.00971882f $X=2.81 $Y=0.665
+ $X2=0 $Y2=0
cc_235 N_A_230_74#_c_254_n N_A_27_112#_M1002_g 0.00982733f $X=2.98 $Y=0.382
+ $X2=0 $Y2=0
cc_236 N_A_230_74#_c_255_n N_A_27_112#_M1002_g 2.18501e-19 $X=3.73 $Y=0.345
+ $X2=0 $Y2=0
cc_237 N_A_230_74#_M1015_d N_A_27_112#_c_397_n 0.0101873f $X=1.2 $Y=1.96 $X2=0
+ $Y2=0
cc_238 N_A_230_74#_c_262_n N_A_27_112#_c_397_n 0.0160246f $X=2.185 $Y=1.885
+ $X2=0 $Y2=0
cc_239 N_A_230_74#_c_268_n N_A_27_112#_c_397_n 0.0287578f $X=1.54 $Y=2.065 $X2=0
+ $Y2=0
cc_240 N_A_230_74#_c_260_n N_A_27_112#_c_397_n 0.00207455f $X=1.7 $Y=1.415 $X2=0
+ $Y2=0
cc_241 N_A_230_74#_c_249_n N_A_27_112#_c_392_n 0.00110392f $X=2.185 $Y=1.49
+ $X2=0 $Y2=0
cc_242 N_A_230_74#_c_262_n N_A_27_112#_c_392_n 0.00702891f $X=2.185 $Y=1.885
+ $X2=0 $Y2=0
cc_243 N_A_230_74#_c_263_n N_A_27_112#_c_392_n 4.70704e-19 $X=3.175 $Y=1.885
+ $X2=0 $Y2=0
cc_244 N_A_230_74#_c_253_n N_A_363_82#_M1000_s 0.00689956f $X=2.81 $Y=0.665
+ $X2=-0.19 $Y2=-0.245
cc_245 N_A_230_74#_c_263_n N_A_363_82#_c_478_n 0.0191917f $X=3.175 $Y=1.885
+ $X2=0 $Y2=0
cc_246 N_A_230_74#_c_264_n N_A_363_82#_c_478_n 0.0163016f $X=3.715 $Y=1.765
+ $X2=0 $Y2=0
cc_247 N_A_230_74#_c_249_n N_A_363_82#_c_471_n 0.00189668f $X=2.185 $Y=1.49
+ $X2=0 $Y2=0
cc_248 N_A_230_74#_c_251_n N_A_363_82#_c_471_n 0.00934554f $X=2.175 $Y=1.225
+ $X2=0 $Y2=0
cc_249 N_A_230_74#_c_253_n N_A_363_82#_c_471_n 0.0267031f $X=2.81 $Y=0.665 $X2=0
+ $Y2=0
cc_250 N_A_230_74#_c_257_n N_A_363_82#_c_471_n 0.0209634f $X=1.29 $Y=0.515 $X2=0
+ $Y2=0
cc_251 N_A_230_74#_c_258_n N_A_363_82#_c_471_n 0.00539606f $X=1.7 $Y=1.505 $X2=0
+ $Y2=0
cc_252 N_A_230_74#_c_259_n N_A_363_82#_c_471_n 0.00596096f $X=1.66 $Y=1.34 $X2=0
+ $Y2=0
cc_253 N_A_230_74#_c_260_n N_A_363_82#_c_471_n 0.00663024f $X=1.7 $Y=1.415 $X2=0
+ $Y2=0
cc_254 N_A_230_74#_c_248_n N_A_363_82#_c_472_n 0.00541098f $X=2.095 $Y=1.415
+ $X2=0 $Y2=0
cc_255 N_A_230_74#_c_249_n N_A_363_82#_c_472_n 0.00546978f $X=2.185 $Y=1.49
+ $X2=0 $Y2=0
cc_256 N_A_230_74#_c_250_n N_A_363_82#_c_472_n 0.00830621f $X=2.185 $Y=1.795
+ $X2=0 $Y2=0
cc_257 N_A_230_74#_c_262_n N_A_363_82#_c_472_n 0.00544217f $X=2.185 $Y=1.885
+ $X2=0 $Y2=0
cc_258 N_A_230_74#_c_267_n N_A_363_82#_c_472_n 0.0110444f $X=1.54 $Y=1.94 $X2=0
+ $Y2=0
cc_259 N_A_230_74#_c_258_n N_A_363_82#_c_472_n 0.0246582f $X=1.7 $Y=1.505 $X2=0
+ $Y2=0
cc_260 N_A_230_74#_c_259_n N_A_363_82#_c_472_n 0.00159827f $X=1.66 $Y=1.34 $X2=0
+ $Y2=0
cc_261 N_A_230_74#_c_260_n N_A_363_82#_c_472_n 9.9735e-19 $X=1.7 $Y=1.415 $X2=0
+ $Y2=0
cc_262 N_A_230_74#_c_249_n N_A_363_82#_c_473_n 0.00507959f $X=2.185 $Y=1.49
+ $X2=0 $Y2=0
cc_263 N_A_230_74#_c_251_n N_A_363_82#_c_473_n 0.00284581f $X=2.175 $Y=1.225
+ $X2=0 $Y2=0
cc_264 N_A_230_74#_c_253_n N_A_363_82#_c_473_n 0.0204051f $X=2.81 $Y=0.665 $X2=0
+ $Y2=0
cc_265 N_A_230_74#_c_254_n N_A_363_82#_c_473_n 0.005856f $X=2.98 $Y=0.382 $X2=0
+ $Y2=0
cc_266 N_A_230_74#_c_263_n N_A_363_82#_c_474_n 0.0200078f $X=3.175 $Y=1.885
+ $X2=0 $Y2=0
cc_267 N_A_230_74#_c_265_n N_A_363_82#_c_474_n 0.0054456f $X=3.265 $Y=1.765
+ $X2=0 $Y2=0
cc_268 N_A_230_74#_M1001_g N_A_363_82#_c_474_n 8.84971e-19 $X=3.79 $Y=0.83 $X2=0
+ $Y2=0
cc_269 N_A_230_74#_c_263_n N_A_363_82#_c_481_n 0.00926804f $X=3.175 $Y=1.885
+ $X2=0 $Y2=0
cc_270 N_A_230_74#_c_263_n N_A_363_82#_c_482_n 0.00205079f $X=3.175 $Y=1.885
+ $X2=0 $Y2=0
cc_271 N_A_230_74#_c_263_n N_A_363_82#_c_483_n 7.07247e-19 $X=3.175 $Y=1.885
+ $X2=0 $Y2=0
cc_272 N_A_230_74#_c_264_n N_A_363_82#_c_483_n 6.37973e-19 $X=3.715 $Y=1.765
+ $X2=0 $Y2=0
cc_273 N_A_230_74#_c_248_n N_A_363_82#_c_484_n 0.00469925f $X=2.095 $Y=1.415
+ $X2=0 $Y2=0
cc_274 N_A_230_74#_c_262_n N_A_363_82#_c_484_n 0.00645464f $X=2.185 $Y=1.885
+ $X2=0 $Y2=0
cc_275 N_A_230_74#_c_268_n N_A_363_82#_c_484_n 0.0216496f $X=1.54 $Y=2.065 $X2=0
+ $Y2=0
cc_276 N_A_230_74#_c_258_n N_A_363_82#_c_484_n 0.00379671f $X=1.7 $Y=1.505 $X2=0
+ $Y2=0
cc_277 N_A_230_74#_c_260_n N_A_363_82#_c_484_n 4.58946e-19 $X=1.7 $Y=1.415 $X2=0
+ $Y2=0
cc_278 N_A_230_74#_c_265_n N_A_363_82#_c_475_n 0.00124259f $X=3.265 $Y=1.765
+ $X2=0 $Y2=0
cc_279 N_A_230_74#_M1001_g N_A_363_82#_c_475_n 4.00544e-19 $X=3.79 $Y=0.83 $X2=0
+ $Y2=0
cc_280 N_A_230_74#_c_255_n N_A_363_82#_c_475_n 0.00497076f $X=3.73 $Y=0.345
+ $X2=0 $Y2=0
cc_281 N_A_230_74#_c_265_n N_A_363_82#_c_476_n 0.019332f $X=3.265 $Y=1.765 $X2=0
+ $Y2=0
cc_282 N_A_230_74#_M1001_g N_A_363_82#_c_476_n 0.0113395f $X=3.79 $Y=0.83 $X2=0
+ $Y2=0
cc_283 N_A_230_74#_M1001_g N_A_363_82#_c_477_n 0.0147384f $X=3.79 $Y=0.83 $X2=0
+ $Y2=0
cc_284 N_A_230_74#_c_254_n N_A_363_82#_c_477_n 0.00569577f $X=2.98 $Y=0.382
+ $X2=0 $Y2=0
cc_285 N_A_230_74#_c_255_n N_A_363_82#_c_477_n 0.0137397f $X=3.73 $Y=0.345 $X2=0
+ $Y2=0
cc_286 N_A_230_74#_c_256_n N_A_363_82#_c_477_n 0.00778027f $X=3.73 $Y=0.345
+ $X2=0 $Y2=0
cc_287 N_A_230_74#_M1001_g N_A_821_98#_c_587_n 0.0393303f $X=3.79 $Y=0.83 $X2=0
+ $Y2=0
cc_288 N_A_230_74#_c_256_n N_A_821_98#_c_587_n 0.00120024f $X=3.73 $Y=0.345
+ $X2=0 $Y2=0
cc_289 N_A_230_74#_M1001_g N_A_821_98#_c_588_n 0.0188158f $X=3.79 $Y=0.83 $X2=0
+ $Y2=0
cc_290 N_A_230_74#_c_255_n N_A_641_80#_M1022_d 0.0024671f $X=3.73 $Y=0.345
+ $X2=-0.19 $Y2=-0.245
cc_291 N_A_230_74#_M1001_g N_A_641_80#_c_760_n 0.00630606f $X=3.79 $Y=0.83 $X2=0
+ $Y2=0
cc_292 N_A_230_74#_c_255_n N_A_641_80#_c_760_n 0.0227491f $X=3.73 $Y=0.345 $X2=0
+ $Y2=0
cc_293 N_A_230_74#_c_256_n N_A_641_80#_c_760_n 0.00305359f $X=3.73 $Y=0.345
+ $X2=0 $Y2=0
cc_294 N_A_230_74#_c_263_n N_A_641_80#_c_755_n 0.00408166f $X=3.175 $Y=1.885
+ $X2=0 $Y2=0
cc_295 N_A_230_74#_c_264_n N_A_641_80#_c_755_n 0.00595711f $X=3.715 $Y=1.765
+ $X2=0 $Y2=0
cc_296 N_A_230_74#_c_265_n N_A_641_80#_c_755_n 0.00102991f $X=3.265 $Y=1.765
+ $X2=0 $Y2=0
cc_297 N_A_230_74#_c_264_n N_A_641_80#_c_749_n 0.00150476f $X=3.715 $Y=1.765
+ $X2=0 $Y2=0
cc_298 N_A_230_74#_M1001_g N_A_641_80#_c_749_n 0.0202191f $X=3.79 $Y=0.83 $X2=0
+ $Y2=0
cc_299 N_A_230_74#_c_264_n N_A_641_80#_c_750_n 0.00422622f $X=3.715 $Y=1.765
+ $X2=0 $Y2=0
cc_300 N_A_230_74#_M1001_g N_A_641_80#_c_750_n 0.00648948f $X=3.79 $Y=0.83 $X2=0
+ $Y2=0
cc_301 N_A_230_74#_c_264_n N_A_641_80#_c_751_n 0.0187322f $X=3.715 $Y=1.765
+ $X2=0 $Y2=0
cc_302 N_A_230_74#_M1001_g N_A_641_80#_c_751_n 9.81799e-19 $X=3.79 $Y=0.83 $X2=0
+ $Y2=0
cc_303 N_A_230_74#_c_262_n N_VPWR_c_935_n 0.00663011f $X=2.185 $Y=1.885 $X2=0
+ $Y2=0
cc_304 N_A_230_74#_c_263_n N_VPWR_c_935_n 4.20358e-19 $X=3.175 $Y=1.885 $X2=0
+ $Y2=0
cc_305 N_A_230_74#_c_262_n N_VPWR_c_945_n 0.00469064f $X=2.185 $Y=1.885 $X2=0
+ $Y2=0
cc_306 N_A_230_74#_c_263_n N_VPWR_c_946_n 0.00278227f $X=3.175 $Y=1.885 $X2=0
+ $Y2=0
cc_307 N_A_230_74#_c_262_n N_VPWR_c_933_n 0.0049649f $X=2.185 $Y=1.885 $X2=0
+ $Y2=0
cc_308 N_A_230_74#_c_263_n N_VPWR_c_933_n 0.00354419f $X=3.175 $Y=1.885 $X2=0
+ $Y2=0
cc_309 N_A_230_74#_c_253_n N_VGND_M1000_d 0.00930264f $X=2.81 $Y=0.665 $X2=0
+ $Y2=0
cc_310 N_A_230_74#_c_257_n N_VGND_c_1132_n 0.02718f $X=1.29 $Y=0.515 $X2=0 $Y2=0
cc_311 N_A_230_74#_M1001_g N_VGND_c_1133_n 0.00214993f $X=3.79 $Y=0.83 $X2=0
+ $Y2=0
cc_312 N_A_230_74#_c_255_n N_VGND_c_1133_n 0.01269f $X=3.73 $Y=0.345 $X2=0 $Y2=0
cc_313 N_A_230_74#_c_256_n N_VGND_c_1133_n 0.00337434f $X=3.73 $Y=0.345 $X2=0
+ $Y2=0
cc_314 N_A_230_74#_c_251_n N_VGND_c_1139_n 0.00794823f $X=2.175 $Y=1.225 $X2=0
+ $Y2=0
cc_315 N_A_230_74#_c_253_n N_VGND_c_1139_n 0.037305f $X=2.81 $Y=0.665 $X2=0
+ $Y2=0
cc_316 N_A_230_74#_c_254_n N_VGND_c_1139_n 0.0113147f $X=2.98 $Y=0.382 $X2=0
+ $Y2=0
cc_317 N_A_230_74#_c_257_n N_VGND_c_1139_n 0.0221178f $X=1.29 $Y=0.515 $X2=0
+ $Y2=0
cc_318 N_A_230_74#_c_253_n N_VGND_c_1140_n 0.00276577f $X=2.81 $Y=0.665 $X2=0
+ $Y2=0
cc_319 N_A_230_74#_c_254_n N_VGND_c_1140_n 0.0117598f $X=2.98 $Y=0.382 $X2=0
+ $Y2=0
cc_320 N_A_230_74#_c_255_n N_VGND_c_1140_n 0.0596213f $X=3.73 $Y=0.345 $X2=0
+ $Y2=0
cc_321 N_A_230_74#_c_256_n N_VGND_c_1140_n 0.00653686f $X=3.73 $Y=0.345 $X2=0
+ $Y2=0
cc_322 N_A_230_74#_c_251_n N_VGND_c_1151_n 0.00533081f $X=2.175 $Y=1.225 $X2=0
+ $Y2=0
cc_323 N_A_230_74#_c_253_n N_VGND_c_1151_n 0.0268131f $X=2.81 $Y=0.665 $X2=0
+ $Y2=0
cc_324 N_A_230_74#_c_254_n N_VGND_c_1151_n 0.00647831f $X=2.98 $Y=0.382 $X2=0
+ $Y2=0
cc_325 N_A_230_74#_c_255_n N_VGND_c_1151_n 0.0332028f $X=3.73 $Y=0.345 $X2=0
+ $Y2=0
cc_326 N_A_230_74#_c_256_n N_VGND_c_1151_n 0.0102677f $X=3.73 $Y=0.345 $X2=0
+ $Y2=0
cc_327 N_A_230_74#_c_257_n N_VGND_c_1151_n 0.0182647f $X=1.29 $Y=0.515 $X2=0
+ $Y2=0
cc_328 N_A_230_74#_c_254_n A_569_80# 0.00410008f $X=2.98 $Y=0.382 $X2=-0.19
+ $Y2=-0.245
cc_329 N_A_230_74#_c_255_n A_569_80# 6.30424e-19 $X=3.73 $Y=0.345 $X2=-0.19
+ $Y2=-0.245
cc_330 N_A_27_112#_c_397_n N_A_363_82#_M1025_s 0.00819116f $X=2.485 $Y=2.445
+ $X2=0 $Y2=0
cc_331 N_A_27_112#_M1002_g N_A_363_82#_c_471_n 0.00107979f $X=2.77 $Y=0.72 $X2=0
+ $Y2=0
cc_332 N_A_27_112#_c_389_n N_A_363_82#_c_472_n 0.00118244f $X=2.755 $Y=1.885
+ $X2=0 $Y2=0
cc_333 N_A_27_112#_M1002_g N_A_363_82#_c_472_n 8.52697e-19 $X=2.77 $Y=0.72 $X2=0
+ $Y2=0
cc_334 N_A_27_112#_c_392_n N_A_363_82#_c_472_n 0.0229906f $X=2.65 $Y=1.635 $X2=0
+ $Y2=0
cc_335 N_A_27_112#_c_389_n N_A_363_82#_c_473_n 0.00147151f $X=2.755 $Y=1.885
+ $X2=0 $Y2=0
cc_336 N_A_27_112#_M1002_g N_A_363_82#_c_473_n 0.0123903f $X=2.77 $Y=0.72 $X2=0
+ $Y2=0
cc_337 N_A_27_112#_c_392_n N_A_363_82#_c_473_n 0.0250055f $X=2.65 $Y=1.635 $X2=0
+ $Y2=0
cc_338 N_A_27_112#_c_389_n N_A_363_82#_c_474_n 0.0139713f $X=2.755 $Y=1.885
+ $X2=0 $Y2=0
cc_339 N_A_27_112#_c_397_n N_A_363_82#_c_474_n 0.0133618f $X=2.485 $Y=2.445
+ $X2=0 $Y2=0
cc_340 N_A_27_112#_c_389_n N_A_363_82#_c_482_n 0.00143578f $X=2.755 $Y=1.885
+ $X2=0 $Y2=0
cc_341 N_A_27_112#_c_389_n N_A_363_82#_c_484_n 2.27922e-19 $X=2.755 $Y=1.885
+ $X2=0 $Y2=0
cc_342 N_A_27_112#_c_397_n N_A_363_82#_c_484_n 0.0259159f $X=2.485 $Y=2.445
+ $X2=0 $Y2=0
cc_343 N_A_27_112#_c_392_n N_A_363_82#_c_484_n 0.0133854f $X=2.65 $Y=1.635 $X2=0
+ $Y2=0
cc_344 N_A_27_112#_M1002_g N_A_363_82#_c_475_n 0.0054138f $X=2.77 $Y=0.72 $X2=0
+ $Y2=0
cc_345 N_A_27_112#_c_392_n N_A_363_82#_c_475_n 0.0661442f $X=2.65 $Y=1.635 $X2=0
+ $Y2=0
cc_346 N_A_27_112#_c_389_n N_A_363_82#_c_476_n 0.0376213f $X=2.755 $Y=1.885
+ $X2=0 $Y2=0
cc_347 N_A_27_112#_M1002_g N_A_363_82#_c_477_n 0.0376213f $X=2.77 $Y=0.72 $X2=0
+ $Y2=0
cc_348 N_A_27_112#_M1002_g N_A_641_80#_c_760_n 8.37329e-19 $X=2.77 $Y=0.72 $X2=0
+ $Y2=0
cc_349 N_A_27_112#_c_397_n N_VPWR_M1019_d 0.0151265f $X=2.485 $Y=2.445 $X2=-0.19
+ $Y2=-0.245
cc_350 N_A_27_112#_c_397_n N_VPWR_M1025_d 0.0102836f $X=2.485 $Y=2.445 $X2=0
+ $Y2=0
cc_351 N_A_27_112#_c_392_n N_VPWR_M1025_d 0.00488198f $X=2.65 $Y=1.635 $X2=0
+ $Y2=0
cc_352 N_A_27_112#_c_397_n N_VPWR_c_934_n 0.0261153f $X=2.485 $Y=2.445 $X2=0
+ $Y2=0
cc_353 N_A_27_112#_c_398_n N_VPWR_c_934_n 0.00818236f $X=0.445 $Y=2.445 $X2=0
+ $Y2=0
cc_354 N_A_27_112#_c_389_n N_VPWR_c_935_n 0.00791234f $X=2.755 $Y=1.885 $X2=0
+ $Y2=0
cc_355 N_A_27_112#_c_397_n N_VPWR_c_935_n 0.0254379f $X=2.485 $Y=2.445 $X2=0
+ $Y2=0
cc_356 N_A_27_112#_c_389_n N_VPWR_c_946_n 0.00413917f $X=2.755 $Y=1.885 $X2=0
+ $Y2=0
cc_357 N_A_27_112#_c_398_n N_VPWR_c_949_n 0.00965232f $X=0.445 $Y=2.445 $X2=0
+ $Y2=0
cc_358 N_A_27_112#_c_389_n N_VPWR_c_933_n 0.00480856f $X=2.755 $Y=1.885 $X2=0
+ $Y2=0
cc_359 N_A_27_112#_c_397_n N_VPWR_c_933_n 0.0603658f $X=2.485 $Y=2.445 $X2=0
+ $Y2=0
cc_360 N_A_27_112#_c_398_n N_VPWR_c_933_n 0.0119361f $X=0.445 $Y=2.445 $X2=0
+ $Y2=0
cc_361 N_A_27_112#_c_391_n N_VGND_c_1132_n 0.0177942f $X=0.265 $Y=0.95 $X2=0
+ $Y2=0
cc_362 N_A_27_112#_M1002_g N_VGND_c_1139_n 0.00142194f $X=2.77 $Y=0.72 $X2=0
+ $Y2=0
cc_363 N_A_27_112#_M1002_g N_VGND_c_1140_n 0.00347067f $X=2.77 $Y=0.72 $X2=0
+ $Y2=0
cc_364 N_A_27_112#_c_391_n N_VGND_c_1146_n 0.00885135f $X=0.265 $Y=0.95 $X2=0
+ $Y2=0
cc_365 N_A_27_112#_M1002_g N_VGND_c_1151_n 0.00414706f $X=2.77 $Y=0.72 $X2=0
+ $Y2=0
cc_366 N_A_27_112#_c_391_n N_VGND_c_1151_n 0.0115776f $X=0.265 $Y=0.95 $X2=0
+ $Y2=0
cc_367 N_A_363_82#_c_478_n N_A_821_98#_c_601_n 0.0332545f $X=3.71 $Y=2.465 $X2=0
+ $Y2=0
cc_368 N_A_363_82#_c_481_n N_A_821_98#_c_601_n 0.00173515f $X=3.705 $Y=2.99
+ $X2=0 $Y2=0
cc_369 N_A_363_82#_c_483_n N_A_821_98#_c_601_n 0.00938739f $X=3.87 $Y=2.215
+ $X2=0 $Y2=0
cc_370 N_A_363_82#_c_478_n N_A_821_98#_c_607_n 9.76153e-19 $X=3.71 $Y=2.465
+ $X2=0 $Y2=0
cc_371 N_A_363_82#_c_483_n N_A_821_98#_c_607_n 0.0181165f $X=3.87 $Y=2.215 $X2=0
+ $Y2=0
cc_372 N_A_363_82#_c_481_n N_A_641_80#_M1010_d 0.00579062f $X=3.705 $Y=2.99
+ $X2=0 $Y2=0
cc_373 N_A_363_82#_c_475_n N_A_641_80#_c_760_n 0.0138103f $X=3.18 $Y=1.215 $X2=0
+ $Y2=0
cc_374 N_A_363_82#_c_476_n N_A_641_80#_c_760_n 0.00107163f $X=3.22 $Y=1.315
+ $X2=0 $Y2=0
cc_375 N_A_363_82#_c_477_n N_A_641_80#_c_760_n 0.00686671f $X=3.22 $Y=1.15 $X2=0
+ $Y2=0
cc_376 N_A_363_82#_c_478_n N_A_641_80#_c_755_n 0.00555548f $X=3.71 $Y=2.465
+ $X2=0 $Y2=0
cc_377 N_A_363_82#_c_474_n N_A_641_80#_c_755_n 0.0643116f $X=3.06 $Y=2.905 $X2=0
+ $Y2=0
cc_378 N_A_363_82#_c_481_n N_A_641_80#_c_755_n 0.012787f $X=3.705 $Y=2.99 $X2=0
+ $Y2=0
cc_379 N_A_363_82#_c_483_n N_A_641_80#_c_755_n 0.041442f $X=3.87 $Y=2.215 $X2=0
+ $Y2=0
cc_380 N_A_363_82#_c_474_n N_A_641_80#_c_749_n 0.00677684f $X=3.06 $Y=2.905
+ $X2=0 $Y2=0
cc_381 N_A_363_82#_c_475_n N_A_641_80#_c_749_n 0.0251828f $X=3.18 $Y=1.215 $X2=0
+ $Y2=0
cc_382 N_A_363_82#_c_476_n N_A_641_80#_c_749_n 0.00224196f $X=3.22 $Y=1.315
+ $X2=0 $Y2=0
cc_383 N_A_363_82#_c_477_n N_A_641_80#_c_749_n 0.00309916f $X=3.22 $Y=1.15 $X2=0
+ $Y2=0
cc_384 N_A_363_82#_c_478_n N_A_641_80#_c_750_n 0.00111766f $X=3.71 $Y=2.465
+ $X2=0 $Y2=0
cc_385 N_A_363_82#_c_478_n N_A_641_80#_c_751_n 8.23934e-19 $X=3.71 $Y=2.465
+ $X2=0 $Y2=0
cc_386 N_A_363_82#_c_474_n N_A_641_80#_c_751_n 0.0131205f $X=3.06 $Y=2.905 $X2=0
+ $Y2=0
cc_387 N_A_363_82#_c_483_n N_A_641_80#_c_751_n 0.0201952f $X=3.87 $Y=2.215 $X2=0
+ $Y2=0
cc_388 N_A_363_82#_c_475_n N_A_641_80#_c_751_n 0.00523479f $X=3.18 $Y=1.215
+ $X2=0 $Y2=0
cc_389 N_A_363_82#_c_476_n N_A_641_80#_c_751_n 2.01687e-19 $X=3.22 $Y=1.315
+ $X2=0 $Y2=0
cc_390 N_A_363_82#_c_474_n N_VPWR_c_935_n 0.010373f $X=3.06 $Y=2.905 $X2=0 $Y2=0
cc_391 N_A_363_82#_c_482_n N_VPWR_c_935_n 0.00984731f $X=3.145 $Y=2.99 $X2=0
+ $Y2=0
cc_392 N_A_363_82#_c_478_n N_VPWR_c_946_n 0.00278193f $X=3.71 $Y=2.465 $X2=0
+ $Y2=0
cc_393 N_A_363_82#_c_481_n N_VPWR_c_946_n 0.0588551f $X=3.705 $Y=2.99 $X2=0
+ $Y2=0
cc_394 N_A_363_82#_c_482_n N_VPWR_c_946_n 0.0119597f $X=3.145 $Y=2.99 $X2=0
+ $Y2=0
cc_395 N_A_363_82#_c_478_n N_VPWR_c_951_n 4.04476e-19 $X=3.71 $Y=2.465 $X2=0
+ $Y2=0
cc_396 N_A_363_82#_c_481_n N_VPWR_c_951_n 0.00796977f $X=3.705 $Y=2.99 $X2=0
+ $Y2=0
cc_397 N_A_363_82#_c_483_n N_VPWR_c_951_n 0.0109526f $X=3.87 $Y=2.215 $X2=0
+ $Y2=0
cc_398 N_A_363_82#_c_478_n N_VPWR_c_933_n 0.00356236f $X=3.71 $Y=2.465 $X2=0
+ $Y2=0
cc_399 N_A_363_82#_c_481_n N_VPWR_c_933_n 0.0327104f $X=3.705 $Y=2.99 $X2=0
+ $Y2=0
cc_400 N_A_363_82#_c_482_n N_VPWR_c_933_n 0.00639333f $X=3.145 $Y=2.99 $X2=0
+ $Y2=0
cc_401 N_A_363_82#_c_474_n A_566_392# 0.00874056f $X=3.06 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_402 N_A_363_82#_c_482_n A_566_392# 5.82339e-19 $X=3.145 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_403 N_A_363_82#_c_481_n A_757_508# 9.16612e-19 $X=3.705 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_404 N_A_363_82#_c_483_n A_757_508# 0.00589473f $X=3.87 $Y=2.215 $X2=-0.19
+ $Y2=-0.245
cc_405 N_A_363_82#_c_473_n N_VGND_M1000_d 0.00306155f $X=2.975 $Y=1.215 $X2=0
+ $Y2=0
cc_406 N_A_363_82#_c_477_n N_VGND_c_1140_n 9.29978e-19 $X=3.22 $Y=1.15 $X2=0
+ $Y2=0
cc_407 N_A_821_98#_c_588_n N_A_641_80#_c_746_n 0.00541465f $X=4.32 $Y=1.99 $X2=0
+ $Y2=0
cc_408 N_A_821_98#_c_601_n N_A_641_80#_c_746_n 0.0210627f $X=4.365 $Y=2.465
+ $X2=0 $Y2=0
cc_409 N_A_821_98#_c_607_n N_A_641_80#_c_746_n 0.0118128f $X=5.095 $Y=2.155
+ $X2=0 $Y2=0
cc_410 N_A_821_98#_c_608_n N_A_641_80#_c_746_n 0.00357621f $X=5.4 $Y=2.4 $X2=0
+ $Y2=0
cc_411 N_A_821_98#_c_611_n N_A_641_80#_c_746_n 0.028744f $X=5.33 $Y=1.805 $X2=0
+ $Y2=0
cc_412 N_A_821_98#_c_599_n N_A_641_80#_c_746_n 0.011448f $X=5.33 $Y=1.72 $X2=0
+ $Y2=0
cc_413 N_A_821_98#_c_594_n N_A_641_80#_M1013_g 0.00506044f $X=4.32 $Y=1.19 $X2=0
+ $Y2=0
cc_414 N_A_821_98#_c_596_n N_A_641_80#_M1013_g 0.0120602f $X=4.955 $Y=0.515
+ $X2=0 $Y2=0
cc_415 N_A_821_98#_c_598_n N_A_641_80#_M1013_g 0.00418289f $X=5.027 $Y=1.13
+ $X2=0 $Y2=0
cc_416 N_A_821_98#_c_599_n N_A_641_80#_M1013_g 0.0114535f $X=5.33 $Y=1.72 $X2=0
+ $Y2=0
cc_417 N_A_821_98#_c_588_n N_A_641_80#_c_748_n 0.0223372f $X=4.32 $Y=1.99 $X2=0
+ $Y2=0
cc_418 N_A_821_98#_c_607_n N_A_641_80#_c_748_n 0.00478787f $X=5.095 $Y=2.155
+ $X2=0 $Y2=0
cc_419 N_A_821_98#_c_598_n N_A_641_80#_c_748_n 0.00838546f $X=5.027 $Y=1.13
+ $X2=0 $Y2=0
cc_420 N_A_821_98#_c_587_n N_A_641_80#_c_760_n 4.80093e-19 $X=4.18 $Y=1.115
+ $X2=0 $Y2=0
cc_421 N_A_821_98#_c_587_n N_A_641_80#_c_749_n 0.00135697f $X=4.18 $Y=1.115
+ $X2=0 $Y2=0
cc_422 N_A_821_98#_c_588_n N_A_641_80#_c_749_n 0.00180539f $X=4.32 $Y=1.99 $X2=0
+ $Y2=0
cc_423 N_A_821_98#_c_588_n N_A_641_80#_c_750_n 0.0129508f $X=4.32 $Y=1.99 $X2=0
+ $Y2=0
cc_424 N_A_821_98#_c_601_n N_A_641_80#_c_750_n 0.00423928f $X=4.365 $Y=2.465
+ $X2=0 $Y2=0
cc_425 N_A_821_98#_c_594_n N_A_641_80#_c_750_n 0.00449484f $X=4.32 $Y=1.19 $X2=0
+ $Y2=0
cc_426 N_A_821_98#_c_607_n N_A_641_80#_c_750_n 0.0266186f $X=5.095 $Y=2.155
+ $X2=0 $Y2=0
cc_427 N_A_821_98#_c_588_n N_A_641_80#_c_752_n 0.00226349f $X=4.32 $Y=1.99 $X2=0
+ $Y2=0
cc_428 N_A_821_98#_c_607_n N_A_641_80#_c_752_n 0.027116f $X=5.095 $Y=2.155 $X2=0
+ $Y2=0
cc_429 N_A_821_98#_c_598_n N_A_641_80#_c_752_n 0.00950973f $X=5.027 $Y=1.13
+ $X2=0 $Y2=0
cc_430 N_A_821_98#_c_599_n N_A_641_80#_c_752_n 0.0345493f $X=5.33 $Y=1.72 $X2=0
+ $Y2=0
cc_431 N_A_821_98#_M1023_g N_RESET_B_c_829_n 0.0158216f $X=6.1 $Y=0.74 $X2=-0.19
+ $Y2=-0.245
cc_432 N_A_821_98#_c_596_n N_RESET_B_c_829_n 0.00349897f $X=4.955 $Y=0.515
+ $X2=-0.19 $Y2=-0.245
cc_433 N_A_821_98#_M1023_g N_RESET_B_c_830_n 0.0178261f $X=6.1 $Y=0.74 $X2=0
+ $Y2=0
cc_434 N_A_821_98#_c_602_n N_RESET_B_c_830_n 0.0199625f $X=6.155 $Y=1.765 $X2=0
+ $Y2=0
cc_435 N_A_821_98#_c_592_n N_RESET_B_c_830_n 0.00721062f $X=6.695 $Y=1.465 $X2=0
+ $Y2=0
cc_436 N_A_821_98#_c_608_n N_RESET_B_c_830_n 0.00698683f $X=5.4 $Y=2.4 $X2=0
+ $Y2=0
cc_437 N_A_821_98#_c_609_n N_RESET_B_c_830_n 0.0144567f $X=5.955 $Y=1.805 $X2=0
+ $Y2=0
cc_438 N_A_821_98#_c_597_n N_RESET_B_c_830_n 0.00425097f $X=6.125 $Y=1.465 $X2=0
+ $Y2=0
cc_439 N_A_821_98#_c_611_n N_RESET_B_c_830_n 0.0114554f $X=5.33 $Y=1.805 $X2=0
+ $Y2=0
cc_440 N_A_821_98#_c_599_n N_RESET_B_c_830_n 0.00410242f $X=5.33 $Y=1.72 $X2=0
+ $Y2=0
cc_441 N_A_821_98#_M1023_g N_RESET_B_c_831_n 0.00141176f $X=6.1 $Y=0.74 $X2=0
+ $Y2=0
cc_442 N_A_821_98#_c_592_n N_RESET_B_c_831_n 2.72691e-19 $X=6.695 $Y=1.465 $X2=0
+ $Y2=0
cc_443 N_A_821_98#_c_609_n N_RESET_B_c_831_n 0.0161187f $X=5.955 $Y=1.805 $X2=0
+ $Y2=0
cc_444 N_A_821_98#_c_597_n N_RESET_B_c_831_n 0.0188908f $X=6.125 $Y=1.465 $X2=0
+ $Y2=0
cc_445 N_A_821_98#_c_611_n N_RESET_B_c_831_n 0.010918f $X=5.33 $Y=1.805 $X2=0
+ $Y2=0
cc_446 N_A_821_98#_c_599_n N_RESET_B_c_831_n 0.0294391f $X=5.33 $Y=1.72 $X2=0
+ $Y2=0
cc_447 N_A_821_98#_c_605_n N_A_1449_368#_c_871_n 0.0252197f $X=7.615 $Y=1.765
+ $X2=0 $Y2=0
cc_448 N_A_821_98#_M1004_g N_A_1449_368#_M1007_g 0.0200925f $X=7.625 $Y=0.79
+ $X2=0 $Y2=0
cc_449 N_A_821_98#_M1024_g N_A_1449_368#_c_865_n 0.00494994f $X=6.53 $Y=0.74
+ $X2=0 $Y2=0
cc_450 N_A_821_98#_M1004_g N_A_1449_368#_c_865_n 0.005981f $X=7.625 $Y=0.79
+ $X2=0 $Y2=0
cc_451 N_A_821_98#_M1004_g N_A_1449_368#_c_866_n 0.00655853f $X=7.625 $Y=0.79
+ $X2=0 $Y2=0
cc_452 N_A_821_98#_c_603_n N_A_1449_368#_c_867_n 0.00594858f $X=6.605 $Y=1.765
+ $X2=0 $Y2=0
cc_453 N_A_821_98#_c_605_n N_A_1449_368#_c_867_n 0.013052f $X=7.615 $Y=1.765
+ $X2=0 $Y2=0
cc_454 N_A_821_98#_c_595_n N_A_1449_368#_c_867_n 0.00578318f $X=7.615 $Y=1.532
+ $X2=0 $Y2=0
cc_455 N_A_821_98#_c_595_n N_A_1449_368#_c_868_n 0.0210573f $X=7.615 $Y=1.532
+ $X2=0 $Y2=0
cc_456 N_A_821_98#_M1004_g N_A_1449_368#_c_869_n 0.00231106f $X=7.625 $Y=0.79
+ $X2=0 $Y2=0
cc_457 N_A_821_98#_c_591_n N_A_1449_368#_c_885_n 0.025616f $X=7.525 $Y=1.465
+ $X2=0 $Y2=0
cc_458 N_A_821_98#_c_595_n N_A_1449_368#_c_885_n 9.32228e-19 $X=7.615 $Y=1.532
+ $X2=0 $Y2=0
cc_459 N_A_821_98#_c_595_n N_A_1449_368#_c_870_n 0.0264068f $X=7.615 $Y=1.532
+ $X2=0 $Y2=0
cc_460 N_A_821_98#_c_607_n N_VPWR_M1021_d 0.00684417f $X=5.095 $Y=2.155 $X2=0
+ $Y2=0
cc_461 N_A_821_98#_c_609_n N_VPWR_M1005_d 0.00222173f $X=5.955 $Y=1.805 $X2=0
+ $Y2=0
cc_462 N_A_821_98#_c_597_n N_VPWR_M1005_d 8.60101e-19 $X=6.125 $Y=1.465 $X2=0
+ $Y2=0
cc_463 N_A_821_98#_c_602_n N_VPWR_c_936_n 0.00197331f $X=6.155 $Y=1.765 $X2=0
+ $Y2=0
cc_464 N_A_821_98#_c_609_n N_VPWR_c_936_n 0.016109f $X=5.955 $Y=1.805 $X2=0
+ $Y2=0
cc_465 N_A_821_98#_c_597_n N_VPWR_c_936_n 0.0059779f $X=6.125 $Y=1.465 $X2=0
+ $Y2=0
cc_466 N_A_821_98#_c_611_n N_VPWR_c_936_n 0.0358158f $X=5.33 $Y=1.805 $X2=0
+ $Y2=0
cc_467 N_A_821_98#_c_602_n N_VPWR_c_937_n 5.85463e-19 $X=6.155 $Y=1.765 $X2=0
+ $Y2=0
cc_468 N_A_821_98#_c_603_n N_VPWR_c_937_n 0.0160427f $X=6.605 $Y=1.765 $X2=0
+ $Y2=0
cc_469 N_A_821_98#_c_591_n N_VPWR_c_937_n 7.63246e-19 $X=7.525 $Y=1.465 $X2=0
+ $Y2=0
cc_470 N_A_821_98#_c_605_n N_VPWR_c_937_n 0.00412926f $X=7.615 $Y=1.765 $X2=0
+ $Y2=0
cc_471 N_A_821_98#_c_605_n N_VPWR_c_938_n 0.00954905f $X=7.615 $Y=1.765 $X2=0
+ $Y2=0
cc_472 N_A_821_98#_c_608_n N_VPWR_c_941_n 0.0145938f $X=5.4 $Y=2.4 $X2=0 $Y2=0
cc_473 N_A_821_98#_c_602_n N_VPWR_c_943_n 0.00461464f $X=6.155 $Y=1.765 $X2=0
+ $Y2=0
cc_474 N_A_821_98#_c_603_n N_VPWR_c_943_n 0.00413917f $X=6.605 $Y=1.765 $X2=0
+ $Y2=0
cc_475 N_A_821_98#_c_601_n N_VPWR_c_946_n 0.00415318f $X=4.365 $Y=2.465 $X2=0
+ $Y2=0
cc_476 N_A_821_98#_c_605_n N_VPWR_c_947_n 0.00481995f $X=7.615 $Y=1.765 $X2=0
+ $Y2=0
cc_477 N_A_821_98#_c_601_n N_VPWR_c_951_n 0.0182121f $X=4.365 $Y=2.465 $X2=0
+ $Y2=0
cc_478 N_A_821_98#_c_607_n N_VPWR_c_951_n 0.0286097f $X=5.095 $Y=2.155 $X2=0
+ $Y2=0
cc_479 N_A_821_98#_c_608_n N_VPWR_c_951_n 0.0144922f $X=5.4 $Y=2.4 $X2=0 $Y2=0
cc_480 N_A_821_98#_c_601_n N_VPWR_c_933_n 0.0085718f $X=4.365 $Y=2.465 $X2=0
+ $Y2=0
cc_481 N_A_821_98#_c_602_n N_VPWR_c_933_n 0.00908585f $X=6.155 $Y=1.765 $X2=0
+ $Y2=0
cc_482 N_A_821_98#_c_603_n N_VPWR_c_933_n 0.00817726f $X=6.605 $Y=1.765 $X2=0
+ $Y2=0
cc_483 N_A_821_98#_c_605_n N_VPWR_c_933_n 0.00508379f $X=7.615 $Y=1.765 $X2=0
+ $Y2=0
cc_484 N_A_821_98#_c_608_n N_VPWR_c_933_n 0.0120466f $X=5.4 $Y=2.4 $X2=0 $Y2=0
cc_485 N_A_821_98#_M1023_g N_Q_c_1047_n 0.00802514f $X=6.1 $Y=0.74 $X2=0 $Y2=0
cc_486 N_A_821_98#_M1024_g N_Q_c_1047_n 0.0131993f $X=6.53 $Y=0.74 $X2=0 $Y2=0
cc_487 N_A_821_98#_c_602_n N_Q_c_1051_n 0.0053278f $X=6.155 $Y=1.765 $X2=0 $Y2=0
cc_488 N_A_821_98#_c_603_n N_Q_c_1051_n 0.00624195f $X=6.605 $Y=1.765 $X2=0
+ $Y2=0
cc_489 N_A_821_98#_c_603_n N_Q_c_1052_n 0.0149886f $X=6.605 $Y=1.765 $X2=0 $Y2=0
cc_490 N_A_821_98#_c_591_n N_Q_c_1052_n 0.00407439f $X=7.525 $Y=1.465 $X2=0
+ $Y2=0
cc_491 N_A_821_98#_c_592_n N_Q_c_1052_n 0.00233698f $X=6.695 $Y=1.465 $X2=0
+ $Y2=0
cc_492 N_A_821_98#_c_605_n N_Q_c_1052_n 3.9824e-19 $X=7.615 $Y=1.765 $X2=0 $Y2=0
cc_493 N_A_821_98#_c_707_p N_Q_c_1052_n 0.0134169f $X=6.53 $Y=1.465 $X2=0 $Y2=0
cc_494 N_A_821_98#_c_602_n N_Q_c_1053_n 0.00268578f $X=6.155 $Y=1.765 $X2=0
+ $Y2=0
cc_495 N_A_821_98#_c_592_n N_Q_c_1053_n 0.00435468f $X=6.695 $Y=1.465 $X2=0
+ $Y2=0
cc_496 N_A_821_98#_c_597_n N_Q_c_1053_n 0.00717337f $X=6.125 $Y=1.465 $X2=0
+ $Y2=0
cc_497 N_A_821_98#_c_707_p N_Q_c_1053_n 0.0143367f $X=6.53 $Y=1.465 $X2=0 $Y2=0
cc_498 N_A_821_98#_M1024_g N_Q_c_1048_n 0.0128805f $X=6.53 $Y=0.74 $X2=0 $Y2=0
cc_499 N_A_821_98#_c_591_n N_Q_c_1048_n 0.00407439f $X=7.525 $Y=1.465 $X2=0
+ $Y2=0
cc_500 N_A_821_98#_M1004_g N_Q_c_1048_n 3.42629e-19 $X=7.625 $Y=0.79 $X2=0 $Y2=0
cc_501 N_A_821_98#_c_707_p N_Q_c_1048_n 0.0122755f $X=6.53 $Y=1.465 $X2=0 $Y2=0
cc_502 N_A_821_98#_M1023_g N_Q_c_1049_n 0.00374068f $X=6.1 $Y=0.74 $X2=0 $Y2=0
cc_503 N_A_821_98#_M1024_g N_Q_c_1049_n 9.7541e-19 $X=6.53 $Y=0.74 $X2=0 $Y2=0
cc_504 N_A_821_98#_c_592_n N_Q_c_1049_n 0.00232957f $X=6.695 $Y=1.465 $X2=0
+ $Y2=0
cc_505 N_A_821_98#_c_707_p N_Q_c_1049_n 0.0276081f $X=6.53 $Y=1.465 $X2=0 $Y2=0
cc_506 N_A_821_98#_M1024_g Q 0.00556303f $X=6.53 $Y=0.74 $X2=0 $Y2=0
cc_507 N_A_821_98#_c_603_n Q 0.00121312f $X=6.605 $Y=1.765 $X2=0 $Y2=0
cc_508 N_A_821_98#_c_591_n Q 0.0259674f $X=7.525 $Y=1.465 $X2=0 $Y2=0
cc_509 N_A_821_98#_c_592_n Q 0.00499466f $X=6.695 $Y=1.465 $X2=0 $Y2=0
cc_510 N_A_821_98#_M1004_g Q 6.46089e-19 $X=7.625 $Y=0.79 $X2=0 $Y2=0
cc_511 N_A_821_98#_c_595_n Q 5.40572e-19 $X=7.615 $Y=1.532 $X2=0 $Y2=0
cc_512 N_A_821_98#_c_707_p Q 0.0223699f $X=6.53 $Y=1.465 $X2=0 $Y2=0
cc_513 N_A_821_98#_c_587_n N_VGND_c_1133_n 0.0144666f $X=4.18 $Y=1.115 $X2=0
+ $Y2=0
cc_514 N_A_821_98#_c_594_n N_VGND_c_1133_n 0.00540622f $X=4.32 $Y=1.19 $X2=0
+ $Y2=0
cc_515 N_A_821_98#_c_596_n N_VGND_c_1133_n 0.0491859f $X=4.955 $Y=0.515 $X2=0
+ $Y2=0
cc_516 N_A_821_98#_M1023_g N_VGND_c_1134_n 0.00889628f $X=6.1 $Y=0.74 $X2=0
+ $Y2=0
cc_517 N_A_821_98#_c_596_n N_VGND_c_1134_n 0.0145513f $X=4.955 $Y=0.515 $X2=0
+ $Y2=0
cc_518 N_A_821_98#_M1024_g N_VGND_c_1135_n 0.013225f $X=6.53 $Y=0.74 $X2=0 $Y2=0
cc_519 N_A_821_98#_c_591_n N_VGND_c_1135_n 7.73684e-19 $X=7.525 $Y=1.465 $X2=0
+ $Y2=0
cc_520 N_A_821_98#_M1004_g N_VGND_c_1135_n 0.00336635f $X=7.625 $Y=0.79 $X2=0
+ $Y2=0
cc_521 N_A_821_98#_M1004_g N_VGND_c_1136_n 0.0074703f $X=7.625 $Y=0.79 $X2=0
+ $Y2=0
cc_522 N_A_821_98#_c_587_n N_VGND_c_1140_n 0.00347405f $X=4.18 $Y=1.115 $X2=0
+ $Y2=0
cc_523 N_A_821_98#_c_596_n N_VGND_c_1142_n 0.0206573f $X=4.955 $Y=0.515 $X2=0
+ $Y2=0
cc_524 N_A_821_98#_M1023_g N_VGND_c_1144_n 0.00434272f $X=6.1 $Y=0.74 $X2=0
+ $Y2=0
cc_525 N_A_821_98#_M1024_g N_VGND_c_1144_n 0.00434272f $X=6.53 $Y=0.74 $X2=0
+ $Y2=0
cc_526 N_A_821_98#_M1004_g N_VGND_c_1147_n 0.00485498f $X=7.625 $Y=0.79 $X2=0
+ $Y2=0
cc_527 N_A_821_98#_c_587_n N_VGND_c_1151_n 0.00395485f $X=4.18 $Y=1.115 $X2=0
+ $Y2=0
cc_528 N_A_821_98#_M1023_g N_VGND_c_1151_n 0.00821985f $X=6.1 $Y=0.74 $X2=0
+ $Y2=0
cc_529 N_A_821_98#_M1024_g N_VGND_c_1151_n 0.00825059f $X=6.53 $Y=0.74 $X2=0
+ $Y2=0
cc_530 N_A_821_98#_M1004_g N_VGND_c_1151_n 0.00514438f $X=7.625 $Y=0.79 $X2=0
+ $Y2=0
cc_531 N_A_821_98#_c_596_n N_VGND_c_1151_n 0.016746f $X=4.955 $Y=0.515 $X2=0
+ $Y2=0
cc_532 N_A_641_80#_M1013_g N_RESET_B_c_829_n 0.0496133f $X=5.17 $Y=0.74
+ $X2=-0.19 $Y2=-0.245
cc_533 N_A_641_80#_c_746_n N_RESET_B_c_830_n 0.0339789f $X=5.125 $Y=1.765 $X2=0
+ $Y2=0
cc_534 N_A_641_80#_M1013_g N_RESET_B_c_830_n 0.0181352f $X=5.17 $Y=0.74 $X2=0
+ $Y2=0
cc_535 N_A_641_80#_M1013_g N_RESET_B_c_831_n 0.00101423f $X=5.17 $Y=0.74 $X2=0
+ $Y2=0
cc_536 N_A_641_80#_c_746_n N_VPWR_c_941_n 0.00415318f $X=5.125 $Y=1.765 $X2=0
+ $Y2=0
cc_537 N_A_641_80#_c_746_n N_VPWR_c_951_n 0.0144285f $X=5.125 $Y=1.765 $X2=0
+ $Y2=0
cc_538 N_A_641_80#_c_746_n N_VPWR_c_933_n 0.00818241f $X=5.125 $Y=1.765 $X2=0
+ $Y2=0
cc_539 N_A_641_80#_M1013_g N_VGND_c_1133_n 0.00414178f $X=5.17 $Y=0.74 $X2=0
+ $Y2=0
cc_540 N_A_641_80#_c_760_n N_VGND_c_1133_n 0.00562511f $X=3.57 $Y=0.875 $X2=0
+ $Y2=0
cc_541 N_A_641_80#_c_749_n N_VGND_c_1133_n 0.00300042f $X=3.655 $Y=1.65 $X2=0
+ $Y2=0
cc_542 N_A_641_80#_c_750_n N_VGND_c_1133_n 0.0109219f $X=4.605 $Y=1.735 $X2=0
+ $Y2=0
cc_543 N_A_641_80#_M1013_g N_VGND_c_1134_n 0.00125099f $X=5.17 $Y=0.74 $X2=0
+ $Y2=0
cc_544 N_A_641_80#_M1013_g N_VGND_c_1142_n 0.00291513f $X=5.17 $Y=0.74 $X2=0
+ $Y2=0
cc_545 N_A_641_80#_M1013_g N_VGND_c_1151_n 0.00363725f $X=5.17 $Y=0.74 $X2=0
+ $Y2=0
cc_546 N_RESET_B_c_830_n N_VPWR_c_936_n 0.00709895f $X=5.625 $Y=1.765 $X2=0
+ $Y2=0
cc_547 N_RESET_B_c_830_n N_VPWR_c_941_n 0.00445602f $X=5.625 $Y=1.765 $X2=0
+ $Y2=0
cc_548 N_RESET_B_c_830_n N_VPWR_c_951_n 4.22856e-19 $X=5.625 $Y=1.765 $X2=0
+ $Y2=0
cc_549 N_RESET_B_c_830_n N_VPWR_c_933_n 0.00858186f $X=5.625 $Y=1.765 $X2=0
+ $Y2=0
cc_550 N_RESET_B_c_829_n N_Q_c_1049_n 3.46348e-19 $X=5.56 $Y=1.22 $X2=0 $Y2=0
cc_551 N_RESET_B_c_829_n N_VGND_c_1134_n 0.0136038f $X=5.56 $Y=1.22 $X2=0 $Y2=0
cc_552 N_RESET_B_c_830_n N_VGND_c_1134_n 9.00702e-19 $X=5.625 $Y=1.765 $X2=0
+ $Y2=0
cc_553 N_RESET_B_c_831_n N_VGND_c_1134_n 0.0124443f $X=5.62 $Y=1.385 $X2=0 $Y2=0
cc_554 N_RESET_B_c_829_n N_VGND_c_1142_n 0.00383152f $X=5.56 $Y=1.22 $X2=0 $Y2=0
cc_555 N_RESET_B_c_829_n N_VGND_c_1151_n 0.0075725f $X=5.56 $Y=1.22 $X2=0 $Y2=0
cc_556 N_A_1449_368#_c_867_n N_VPWR_c_937_n 0.0444757f $X=7.39 $Y=1.985 $X2=0
+ $Y2=0
cc_557 N_A_1449_368#_c_871_n N_VPWR_c_938_n 0.0118632f $X=8.165 $Y=1.765 $X2=0
+ $Y2=0
cc_558 N_A_1449_368#_c_867_n N_VPWR_c_938_n 0.0402324f $X=7.39 $Y=1.985 $X2=0
+ $Y2=0
cc_559 N_A_1449_368#_c_868_n N_VPWR_c_938_n 0.026236f $X=8.08 $Y=1.465 $X2=0
+ $Y2=0
cc_560 N_A_1449_368#_c_870_n N_VPWR_c_938_n 0.00320573f $X=8.615 $Y=1.532 $X2=0
+ $Y2=0
cc_561 N_A_1449_368#_c_872_n N_VPWR_c_940_n 0.00954146f $X=8.615 $Y=1.765 $X2=0
+ $Y2=0
cc_562 N_A_1449_368#_c_867_n N_VPWR_c_947_n 0.00919855f $X=7.39 $Y=1.985 $X2=0
+ $Y2=0
cc_563 N_A_1449_368#_c_871_n N_VPWR_c_948_n 0.00445602f $X=8.165 $Y=1.765 $X2=0
+ $Y2=0
cc_564 N_A_1449_368#_c_872_n N_VPWR_c_948_n 0.00411612f $X=8.615 $Y=1.765 $X2=0
+ $Y2=0
cc_565 N_A_1449_368#_c_871_n N_VPWR_c_933_n 0.00861719f $X=8.165 $Y=1.765 $X2=0
+ $Y2=0
cc_566 N_A_1449_368#_c_872_n N_VPWR_c_933_n 0.00751023f $X=8.615 $Y=1.765 $X2=0
+ $Y2=0
cc_567 N_A_1449_368#_c_867_n N_VPWR_c_933_n 0.0105074f $X=7.39 $Y=1.985 $X2=0
+ $Y2=0
cc_568 N_A_1449_368#_c_867_n N_Q_c_1052_n 0.0147754f $X=7.39 $Y=1.985 $X2=0
+ $Y2=0
cc_569 N_A_1449_368#_c_865_n N_Q_c_1048_n 0.0149965f $X=7.41 $Y=0.615 $X2=0
+ $Y2=0
cc_570 N_A_1449_368#_c_866_n Q 0.0135906f $X=7.4 $Y=1.3 $X2=0 $Y2=0
cc_571 N_A_1449_368#_c_867_n Q 0.0136317f $X=7.39 $Y=1.985 $X2=0 $Y2=0
cc_572 N_A_1449_368#_c_885_n Q 0.0256724f $X=7.4 $Y=1.465 $X2=0 $Y2=0
cc_573 N_A_1449_368#_M1007_g N_Q_N_c_1102_n 0.00746865f $X=8.195 $Y=0.74 $X2=0
+ $Y2=0
cc_574 N_A_1449_368#_M1014_g N_Q_N_c_1102_n 0.0081896f $X=8.625 $Y=0.74 $X2=0
+ $Y2=0
cc_575 N_A_1449_368#_M1007_g N_Q_N_c_1103_n 0.00316221f $X=8.195 $Y=0.74 $X2=0
+ $Y2=0
cc_576 N_A_1449_368#_M1014_g N_Q_N_c_1103_n 0.00215589f $X=8.625 $Y=0.74 $X2=0
+ $Y2=0
cc_577 N_A_1449_368#_c_870_n N_Q_N_c_1103_n 0.00244427f $X=8.615 $Y=1.532 $X2=0
+ $Y2=0
cc_578 N_A_1449_368#_c_871_n Q_N 0.00218574f $X=8.165 $Y=1.765 $X2=0 $Y2=0
cc_579 N_A_1449_368#_c_872_n Q_N 0.00240464f $X=8.615 $Y=1.765 $X2=0 $Y2=0
cc_580 N_A_1449_368#_c_868_n Q_N 0.00140951f $X=8.08 $Y=1.465 $X2=0 $Y2=0
cc_581 N_A_1449_368#_c_870_n Q_N 0.00807114f $X=8.615 $Y=1.532 $X2=0 $Y2=0
cc_582 N_A_1449_368#_c_871_n Q_N 0.0104214f $X=8.165 $Y=1.765 $X2=0 $Y2=0
cc_583 N_A_1449_368#_c_872_n Q_N 0.0130738f $X=8.615 $Y=1.765 $X2=0 $Y2=0
cc_584 N_A_1449_368#_M1007_g N_Q_N_c_1104_n 0.0025553f $X=8.195 $Y=0.74 $X2=0
+ $Y2=0
cc_585 N_A_1449_368#_c_872_n N_Q_N_c_1104_n 0.0030228f $X=8.615 $Y=1.765 $X2=0
+ $Y2=0
cc_586 N_A_1449_368#_M1014_g N_Q_N_c_1104_n 0.00866774f $X=8.625 $Y=0.74 $X2=0
+ $Y2=0
cc_587 N_A_1449_368#_c_868_n N_Q_N_c_1104_n 0.0249855f $X=8.08 $Y=1.465 $X2=0
+ $Y2=0
cc_588 N_A_1449_368#_c_870_n N_Q_N_c_1104_n 0.0359686f $X=8.615 $Y=1.532 $X2=0
+ $Y2=0
cc_589 N_A_1449_368#_c_865_n N_VGND_c_1135_n 0.0207909f $X=7.41 $Y=0.615 $X2=0
+ $Y2=0
cc_590 N_A_1449_368#_M1007_g N_VGND_c_1136_n 0.0093706f $X=8.195 $Y=0.74 $X2=0
+ $Y2=0
cc_591 N_A_1449_368#_c_865_n N_VGND_c_1136_n 0.0270587f $X=7.41 $Y=0.615 $X2=0
+ $Y2=0
cc_592 N_A_1449_368#_c_868_n N_VGND_c_1136_n 0.028359f $X=8.08 $Y=1.465 $X2=0
+ $Y2=0
cc_593 N_A_1449_368#_c_870_n N_VGND_c_1136_n 0.00370401f $X=8.615 $Y=1.532 $X2=0
+ $Y2=0
cc_594 N_A_1449_368#_M1014_g N_VGND_c_1138_n 0.00646793f $X=8.625 $Y=0.74 $X2=0
+ $Y2=0
cc_595 N_A_1449_368#_c_865_n N_VGND_c_1147_n 0.0103491f $X=7.41 $Y=0.615 $X2=0
+ $Y2=0
cc_596 N_A_1449_368#_M1007_g N_VGND_c_1148_n 0.00434272f $X=8.195 $Y=0.74 $X2=0
+ $Y2=0
cc_597 N_A_1449_368#_M1014_g N_VGND_c_1148_n 0.00422942f $X=8.625 $Y=0.74 $X2=0
+ $Y2=0
cc_598 N_A_1449_368#_M1007_g N_VGND_c_1151_n 0.00825059f $X=8.195 $Y=0.74 $X2=0
+ $Y2=0
cc_599 N_A_1449_368#_M1014_g N_VGND_c_1151_n 0.00787255f $X=8.625 $Y=0.74 $X2=0
+ $Y2=0
cc_600 N_A_1449_368#_c_865_n N_VGND_c_1151_n 0.0113354f $X=7.41 $Y=0.615 $X2=0
+ $Y2=0
cc_601 N_VPWR_c_936_n N_Q_c_1051_n 0.027389f $X=5.9 $Y=2.145 $X2=0 $Y2=0
cc_602 N_VPWR_c_937_n N_Q_c_1051_n 0.0547423f $X=6.83 $Y=2.305 $X2=0 $Y2=0
cc_603 N_VPWR_c_943_n N_Q_c_1051_n 0.00749631f $X=6.665 $Y=3.33 $X2=0 $Y2=0
cc_604 N_VPWR_c_933_n N_Q_c_1051_n 0.0062048f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_605 N_VPWR_M1026_d N_Q_c_1052_n 0.00340353f $X=6.68 $Y=1.84 $X2=0 $Y2=0
cc_606 N_VPWR_c_937_n N_Q_c_1052_n 0.0232758f $X=6.83 $Y=2.305 $X2=0 $Y2=0
cc_607 N_VPWR_c_938_n Q_N 0.0456525f $X=7.89 $Y=1.985 $X2=0 $Y2=0
cc_608 N_VPWR_c_940_n Q_N 0.0887573f $X=8.84 $Y=1.985 $X2=0 $Y2=0
cc_609 N_VPWR_c_948_n Q_N 0.0158009f $X=8.755 $Y=3.33 $X2=0 $Y2=0
cc_610 N_VPWR_c_933_n Q_N 0.0129424f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_611 N_Q_c_1048_n N_VGND_M1024_s 0.00464869f $X=6.845 $Y=1.045 $X2=0 $Y2=0
cc_612 N_Q_c_1047_n N_VGND_c_1134_n 0.0402483f $X=6.315 $Y=0.515 $X2=0 $Y2=0
cc_613 N_Q_c_1049_n N_VGND_c_1134_n 0.00349775f $X=6.48 $Y=1.045 $X2=0 $Y2=0
cc_614 N_Q_c_1047_n N_VGND_c_1135_n 0.0173003f $X=6.315 $Y=0.515 $X2=0 $Y2=0
cc_615 N_Q_c_1048_n N_VGND_c_1135_n 0.027001f $X=6.845 $Y=1.045 $X2=0 $Y2=0
cc_616 N_Q_c_1047_n N_VGND_c_1144_n 0.0144922f $X=6.315 $Y=0.515 $X2=0 $Y2=0
cc_617 N_Q_c_1047_n N_VGND_c_1151_n 0.0118826f $X=6.315 $Y=0.515 $X2=0 $Y2=0
cc_618 N_Q_N_c_1102_n N_VGND_c_1136_n 0.0309448f $X=8.41 $Y=0.515 $X2=0 $Y2=0
cc_619 N_Q_N_c_1102_n N_VGND_c_1138_n 0.0308798f $X=8.41 $Y=0.515 $X2=0 $Y2=0
cc_620 N_Q_N_c_1102_n N_VGND_c_1148_n 0.0149085f $X=8.41 $Y=0.515 $X2=0 $Y2=0
cc_621 N_Q_N_c_1102_n N_VGND_c_1151_n 0.0122037f $X=8.41 $Y=0.515 $X2=0 $Y2=0
