* File: sky130_fd_sc_ls__or3_1.pxi.spice
* Created: Fri Aug 28 13:58:13 2020
* 
x_PM_SKY130_FD_SC_LS__OR3_1%C N_C_M1006_g N_C_c_50_n N_C_M1004_g C N_C_c_51_n
+ PM_SKY130_FD_SC_LS__OR3_1%C
x_PM_SKY130_FD_SC_LS__OR3_1%B N_B_c_75_n N_B_M1000_g N_B_M1002_g B
+ PM_SKY130_FD_SC_LS__OR3_1%B
x_PM_SKY130_FD_SC_LS__OR3_1%A N_A_c_108_n N_A_M1007_g N_A_M1001_g A N_A_c_106_n
+ N_A_c_107_n PM_SKY130_FD_SC_LS__OR3_1%A
x_PM_SKY130_FD_SC_LS__OR3_1%A_27_74# N_A_27_74#_M1006_s N_A_27_74#_M1002_d
+ N_A_27_74#_M1004_s N_A_27_74#_c_140_n N_A_27_74#_M1005_g N_A_27_74#_M1003_g
+ N_A_27_74#_c_142_n N_A_27_74#_c_143_n N_A_27_74#_c_155_n N_A_27_74#_c_144_n
+ N_A_27_74#_c_145_n N_A_27_74#_c_146_n N_A_27_74#_c_151_n N_A_27_74#_c_147_n
+ N_A_27_74#_c_148_n PM_SKY130_FD_SC_LS__OR3_1%A_27_74#
x_PM_SKY130_FD_SC_LS__OR3_1%VPWR N_VPWR_M1007_d N_VPWR_c_226_n VPWR
+ N_VPWR_c_227_n N_VPWR_c_228_n N_VPWR_c_225_n N_VPWR_c_230_n
+ PM_SKY130_FD_SC_LS__OR3_1%VPWR
x_PM_SKY130_FD_SC_LS__OR3_1%X N_X_M1003_d N_X_M1005_d N_X_c_254_n N_X_c_255_n
+ N_X_c_251_n X X X PM_SKY130_FD_SC_LS__OR3_1%X
x_PM_SKY130_FD_SC_LS__OR3_1%VGND N_VGND_M1006_d N_VGND_M1001_d N_VGND_c_275_n
+ N_VGND_c_276_n VGND N_VGND_c_277_n N_VGND_c_278_n N_VGND_c_279_n
+ N_VGND_c_280_n N_VGND_c_281_n N_VGND_c_282_n PM_SKY130_FD_SC_LS__OR3_1%VGND
cc_1 VNB N_C_M1006_g 0.0444924f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.645
cc_2 VNB N_C_c_50_n 0.0279672f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_3 VNB N_C_c_51_n 0.0153111f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.515
cc_4 VNB N_B_c_75_n 0.022865f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.35
cc_5 VNB N_B_M1002_g 0.0402646f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.34
cc_6 VNB B 0.00552308f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_7 VNB N_A_M1001_g 0.0411168f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.34
cc_8 VNB N_A_c_106_n 0.0363017f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.515
cc_9 VNB N_A_c_107_n 0.00231998f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.565
cc_10 VNB N_A_27_74#_c_140_n 0.0355378f $X=-0.19 $Y=-0.245 $X2=0.41 $Y2=1.515
cc_11 VNB N_A_27_74#_M1003_g 0.0287882f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_74#_c_142_n 0.0277943f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_74#_c_143_n 0.00992268f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_74#_c_144_n 0.00979143f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_74#_c_145_n 0.00746217f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_27_74#_c_146_n 4.2489e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_27_74#_c_147_n 0.0161083f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_27_74#_c_148_n 0.0109349f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_VPWR_c_225_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_X_c_251_n 0.0247379f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB X 0.0267037f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.565
cc_22 VNB X 0.0139384f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_275_n 0.00651905f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_276_n 0.00981015f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.565
cc_25 VNB N_VGND_c_277_n 0.0173909f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_278_n 0.028973f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_279_n 0.0190372f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_280_n 0.186353f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_281_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_282_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VPB N_C_c_50_n 0.0330009f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_32 VPB N_C_c_51_n 0.00759236f $X=-0.19 $Y=1.66 $X2=0.405 $Y2=1.515
cc_33 VPB N_B_c_75_n 0.0264967f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.35
cc_34 VPB B 0.0046645f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_35 VPB N_A_c_108_n 0.0181457f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.35
cc_36 VPB N_A_c_106_n 0.0167473f $X=-0.19 $Y=1.66 $X2=0.405 $Y2=1.515
cc_37 VPB N_A_c_107_n 0.00311553f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.565
cc_38 VPB N_A_27_74#_c_140_n 0.0304506f $X=-0.19 $Y=1.66 $X2=0.41 $Y2=1.515
cc_39 VPB N_A_27_74#_c_146_n 0.00336149f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_40 VPB N_A_27_74#_c_151_n 0.0389799f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_41 VPB N_VPWR_c_226_n 0.0145621f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.34
cc_42 VPB N_VPWR_c_227_n 0.0496025f $X=-0.19 $Y=1.66 $X2=0.41 $Y2=1.515
cc_43 VPB N_VPWR_c_228_n 0.017793f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_44 VPB N_VPWR_c_225_n 0.0880907f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_45 VPB N_VPWR_c_230_n 0.0144122f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_X_c_254_n 0.0101094f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.34
cc_47 VPB N_X_c_255_n 0.0417436f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 VPB N_X_c_251_n 0.00756921f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 N_C_c_50_n N_B_c_75_n 0.0785041f $X=0.505 $Y=1.765 $X2=-0.19 $Y2=-0.245
cc_50 N_C_c_51_n N_B_c_75_n 5.45764e-19 $X=0.405 $Y=1.515 $X2=-0.19 $Y2=-0.245
cc_51 N_C_M1006_g N_B_M1002_g 0.0293272f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_52 N_C_c_50_n B 7.89422e-19 $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_53 N_C_c_51_n B 0.0239141f $X=0.405 $Y=1.515 $X2=0 $Y2=0
cc_54 N_C_M1006_g N_A_27_74#_c_142_n 0.00712316f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_55 N_C_c_50_n N_A_27_74#_c_143_n 0.00291196f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_56 N_C_c_51_n N_A_27_74#_c_143_n 0.0211058f $X=0.405 $Y=1.515 $X2=0 $Y2=0
cc_57 N_C_c_50_n N_A_27_74#_c_155_n 0.0120413f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_58 N_C_c_51_n N_A_27_74#_c_155_n 0.00908651f $X=0.405 $Y=1.515 $X2=0 $Y2=0
cc_59 N_C_c_50_n N_A_27_74#_c_151_n 0.018692f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_60 N_C_c_51_n N_A_27_74#_c_151_n 0.0255992f $X=0.405 $Y=1.515 $X2=0 $Y2=0
cc_61 N_C_M1006_g N_A_27_74#_c_147_n 0.0160891f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_62 N_C_c_50_n N_A_27_74#_c_147_n 0.00153002f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_63 N_C_c_51_n N_A_27_74#_c_147_n 0.0151257f $X=0.405 $Y=1.515 $X2=0 $Y2=0
cc_64 N_C_M1006_g N_A_27_74#_c_148_n 8.67149e-19 $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_65 N_C_c_50_n N_VPWR_c_227_n 0.00481995f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_66 N_C_c_50_n N_VPWR_c_225_n 0.00508379f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_67 N_C_M1006_g N_VGND_c_275_n 0.0130729f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_68 N_C_M1006_g N_VGND_c_277_n 0.00383152f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_69 N_C_M1006_g N_VGND_c_280_n 0.00761198f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_70 N_B_c_75_n N_A_c_108_n 0.0371947f $X=0.925 $Y=1.765 $X2=-0.19 $Y2=-0.245
cc_71 N_B_M1002_g N_A_M1001_g 0.0120173f $X=0.995 $Y=0.645 $X2=0 $Y2=0
cc_72 N_B_c_75_n N_A_c_106_n 0.0198431f $X=0.925 $Y=1.765 $X2=0 $Y2=0
cc_73 B N_A_c_106_n 0.00328391f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_74 N_B_c_75_n N_A_c_107_n 3.53813e-19 $X=0.925 $Y=1.765 $X2=0 $Y2=0
cc_75 B N_A_c_107_n 0.0350348f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_76 N_B_c_75_n N_A_27_74#_c_155_n 0.0163537f $X=0.925 $Y=1.765 $X2=0 $Y2=0
cc_77 B N_A_27_74#_c_155_n 0.0346145f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_78 N_B_c_75_n N_A_27_74#_c_151_n 0.00355341f $X=0.925 $Y=1.765 $X2=0 $Y2=0
cc_79 N_B_c_75_n N_A_27_74#_c_147_n 0.00219783f $X=0.925 $Y=1.765 $X2=0 $Y2=0
cc_80 N_B_M1002_g N_A_27_74#_c_147_n 0.0114826f $X=0.995 $Y=0.645 $X2=0 $Y2=0
cc_81 B N_A_27_74#_c_147_n 0.0392242f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_82 N_B_c_75_n N_A_27_74#_c_148_n 0.00221201f $X=0.925 $Y=1.765 $X2=0 $Y2=0
cc_83 N_B_M1002_g N_A_27_74#_c_148_n 0.0163295f $X=0.995 $Y=0.645 $X2=0 $Y2=0
cc_84 N_B_c_75_n N_VPWR_c_226_n 0.00302472f $X=0.925 $Y=1.765 $X2=0 $Y2=0
cc_85 N_B_c_75_n N_VPWR_c_227_n 0.0049405f $X=0.925 $Y=1.765 $X2=0 $Y2=0
cc_86 N_B_c_75_n N_VPWR_c_225_n 0.00508379f $X=0.925 $Y=1.765 $X2=0 $Y2=0
cc_87 N_B_M1002_g N_VGND_c_275_n 0.00593102f $X=0.995 $Y=0.645 $X2=0 $Y2=0
cc_88 N_B_M1002_g N_VGND_c_278_n 0.00435437f $X=0.995 $Y=0.645 $X2=0 $Y2=0
cc_89 N_B_M1002_g N_VGND_c_280_n 0.0082237f $X=0.995 $Y=0.645 $X2=0 $Y2=0
cc_90 N_A_M1001_g N_A_27_74#_c_140_n 0.0177468f $X=1.81 $Y=0.645 $X2=0 $Y2=0
cc_91 N_A_c_106_n N_A_27_74#_c_140_n 0.00193517f $X=1.65 $Y=1.515 $X2=0 $Y2=0
cc_92 N_A_c_107_n N_A_27_74#_c_140_n 3.03321e-19 $X=1.65 $Y=1.515 $X2=0 $Y2=0
cc_93 N_A_M1001_g N_A_27_74#_M1003_g 0.0220159f $X=1.81 $Y=0.645 $X2=0 $Y2=0
cc_94 N_A_c_108_n N_A_27_74#_c_155_n 0.0191733f $X=1.495 $Y=1.765 $X2=0 $Y2=0
cc_95 N_A_c_106_n N_A_27_74#_c_155_n 0.00381302f $X=1.65 $Y=1.515 $X2=0 $Y2=0
cc_96 N_A_c_107_n N_A_27_74#_c_155_n 0.0236066f $X=1.65 $Y=1.515 $X2=0 $Y2=0
cc_97 N_A_M1001_g N_A_27_74#_c_144_n 0.0135443f $X=1.81 $Y=0.645 $X2=0 $Y2=0
cc_98 N_A_M1001_g N_A_27_74#_c_145_n 0.00572869f $X=1.81 $Y=0.645 $X2=0 $Y2=0
cc_99 N_A_c_107_n N_A_27_74#_c_145_n 0.0156671f $X=1.65 $Y=1.515 $X2=0 $Y2=0
cc_100 N_A_c_108_n N_A_27_74#_c_146_n 0.00408171f $X=1.495 $Y=1.765 $X2=0 $Y2=0
cc_101 N_A_c_106_n N_A_27_74#_c_146_n 6.56864e-19 $X=1.65 $Y=1.515 $X2=0 $Y2=0
cc_102 N_A_c_107_n N_A_27_74#_c_146_n 0.00827245f $X=1.65 $Y=1.515 $X2=0 $Y2=0
cc_103 N_A_M1001_g N_A_27_74#_c_148_n 0.0162445f $X=1.81 $Y=0.645 $X2=0 $Y2=0
cc_104 N_A_c_106_n N_A_27_74#_c_148_n 0.00583308f $X=1.65 $Y=1.515 $X2=0 $Y2=0
cc_105 N_A_c_107_n N_A_27_74#_c_148_n 0.0273553f $X=1.65 $Y=1.515 $X2=0 $Y2=0
cc_106 N_A_c_108_n N_VPWR_c_226_n 0.01807f $X=1.495 $Y=1.765 $X2=0 $Y2=0
cc_107 N_A_c_108_n N_VPWR_c_227_n 0.00443511f $X=1.495 $Y=1.765 $X2=0 $Y2=0
cc_108 N_A_c_108_n N_VPWR_c_225_n 0.00460931f $X=1.495 $Y=1.765 $X2=0 $Y2=0
cc_109 N_A_M1001_g X 7.18714e-19 $X=1.81 $Y=0.645 $X2=0 $Y2=0
cc_110 N_A_M1001_g N_VGND_c_276_n 0.00642087f $X=1.81 $Y=0.645 $X2=0 $Y2=0
cc_111 N_A_M1001_g N_VGND_c_278_n 0.00435437f $X=1.81 $Y=0.645 $X2=0 $Y2=0
cc_112 N_A_M1001_g N_VGND_c_280_n 0.0082291f $X=1.81 $Y=0.645 $X2=0 $Y2=0
cc_113 N_A_27_74#_c_155_n A_116_368# 0.0119045f $X=2.09 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_114 N_A_27_74#_c_155_n A_200_368# 0.016602f $X=2.09 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_115 N_A_27_74#_c_155_n N_VPWR_M1007_d 0.0214124f $X=2.09 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_116 N_A_27_74#_c_146_n N_VPWR_M1007_d 0.00262568f $X=2.175 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_117 N_A_27_74#_c_140_n N_VPWR_c_226_n 0.0177874f $X=2.375 $Y=1.765 $X2=0
+ $Y2=0
cc_118 N_A_27_74#_c_155_n N_VPWR_c_226_n 0.0524065f $X=2.09 $Y=2.035 $X2=0 $Y2=0
cc_119 N_A_27_74#_c_145_n N_VPWR_c_226_n 8.31827e-19 $X=2.175 $Y=1.63 $X2=0
+ $Y2=0
cc_120 N_A_27_74#_c_151_n N_VPWR_c_227_n 0.0097982f $X=0.28 $Y=2.115 $X2=0 $Y2=0
cc_121 N_A_27_74#_c_140_n N_VPWR_c_228_n 0.00413917f $X=2.375 $Y=1.765 $X2=0
+ $Y2=0
cc_122 N_A_27_74#_c_140_n N_VPWR_c_225_n 0.00821221f $X=2.375 $Y=1.765 $X2=0
+ $Y2=0
cc_123 N_A_27_74#_c_151_n N_VPWR_c_225_n 0.0111907f $X=0.28 $Y=2.115 $X2=0 $Y2=0
cc_124 N_A_27_74#_c_140_n N_X_c_254_n 0.00916662f $X=2.375 $Y=1.765 $X2=0 $Y2=0
cc_125 N_A_27_74#_c_146_n N_X_c_254_n 0.00434166f $X=2.175 $Y=1.95 $X2=0 $Y2=0
cc_126 N_A_27_74#_c_140_n N_X_c_251_n 0.010619f $X=2.375 $Y=1.765 $X2=0 $Y2=0
cc_127 N_A_27_74#_M1003_g N_X_c_251_n 0.0025312f $X=2.38 $Y=0.74 $X2=0 $Y2=0
cc_128 N_A_27_74#_c_145_n N_X_c_251_n 0.0304389f $X=2.175 $Y=1.63 $X2=0 $Y2=0
cc_129 N_A_27_74#_c_146_n N_X_c_251_n 0.00616973f $X=2.175 $Y=1.95 $X2=0 $Y2=0
cc_130 N_A_27_74#_M1003_g X 0.00941145f $X=2.38 $Y=0.74 $X2=0 $Y2=0
cc_131 N_A_27_74#_c_148_n X 0.0050994f $X=1.76 $Y=0.817 $X2=0 $Y2=0
cc_132 N_A_27_74#_c_140_n X 4.6089e-19 $X=2.375 $Y=1.765 $X2=0 $Y2=0
cc_133 N_A_27_74#_M1003_g X 0.0032303f $X=2.38 $Y=0.74 $X2=0 $Y2=0
cc_134 N_A_27_74#_c_145_n X 0.00740597f $X=2.175 $Y=1.63 $X2=0 $Y2=0
cc_135 N_A_27_74#_c_144_n N_VGND_M1001_d 5.19034e-19 $X=2.09 $Y=1.095 $X2=0
+ $Y2=0
cc_136 N_A_27_74#_c_145_n N_VGND_M1001_d 0.00275048f $X=2.175 $Y=1.63 $X2=0
+ $Y2=0
cc_137 N_A_27_74#_c_142_n N_VGND_c_275_n 0.017215f $X=0.28 $Y=0.645 $X2=0 $Y2=0
cc_138 N_A_27_74#_c_147_n N_VGND_c_275_n 0.0211984f $X=1.045 $Y=0.817 $X2=0
+ $Y2=0
cc_139 N_A_27_74#_c_140_n N_VGND_c_276_n 5.51659e-19 $X=2.375 $Y=1.765 $X2=0
+ $Y2=0
cc_140 N_A_27_74#_M1003_g N_VGND_c_276_n 0.00604382f $X=2.38 $Y=0.74 $X2=0 $Y2=0
cc_141 N_A_27_74#_c_144_n N_VGND_c_276_n 0.0111634f $X=2.09 $Y=1.095 $X2=0 $Y2=0
cc_142 N_A_27_74#_c_145_n N_VGND_c_276_n 0.0126115f $X=2.175 $Y=1.63 $X2=0 $Y2=0
cc_143 N_A_27_74#_c_142_n N_VGND_c_277_n 0.011066f $X=0.28 $Y=0.645 $X2=0 $Y2=0
cc_144 N_A_27_74#_c_148_n N_VGND_c_278_n 0.0198465f $X=1.76 $Y=0.817 $X2=0 $Y2=0
cc_145 N_A_27_74#_M1003_g N_VGND_c_279_n 0.00434272f $X=2.38 $Y=0.74 $X2=0 $Y2=0
cc_146 N_A_27_74#_M1003_g N_VGND_c_280_n 0.00824987f $X=2.38 $Y=0.74 $X2=0 $Y2=0
cc_147 N_A_27_74#_c_142_n N_VGND_c_280_n 0.00915947f $X=0.28 $Y=0.645 $X2=0
+ $Y2=0
cc_148 N_A_27_74#_c_148_n N_VGND_c_280_n 0.0243841f $X=1.76 $Y=0.817 $X2=0 $Y2=0
cc_149 N_VPWR_c_226_n N_X_c_255_n 0.0493647f $X=2.15 $Y=2.375 $X2=0 $Y2=0
cc_150 N_VPWR_c_228_n N_X_c_255_n 0.0124046f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_151 N_VPWR_c_225_n N_X_c_255_n 0.0102675f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_152 X N_VGND_c_276_n 0.0183192f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_153 X N_VGND_c_279_n 0.0161257f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_154 X N_VGND_c_280_n 0.013291f $X=2.555 $Y=0.47 $X2=0 $Y2=0
