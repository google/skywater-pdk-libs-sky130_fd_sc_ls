* File: sky130_fd_sc_ls__and4_1.pxi.spice
* Created: Wed Sep  2 10:55:25 2020
* 
x_PM_SKY130_FD_SC_LS__AND4_1%A N_A_c_76_n N_A_c_77_n N_A_M1005_g N_A_M1007_g
+ N_A_c_71_n N_A_c_72_n N_A_c_73_n A A N_A_c_74_n N_A_c_75_n
+ PM_SKY130_FD_SC_LS__AND4_1%A
x_PM_SKY130_FD_SC_LS__AND4_1%B N_B_c_114_n N_B_c_115_n N_B_M1003_g N_B_M1008_g B
+ B B B N_B_c_113_n PM_SKY130_FD_SC_LS__AND4_1%B
x_PM_SKY130_FD_SC_LS__AND4_1%C N_C_M1006_g N_C_c_158_n N_C_c_159_n N_C_M1009_g
+ N_C_c_153_n N_C_c_154_n N_C_c_155_n C C C C N_C_c_157_n
+ PM_SKY130_FD_SC_LS__AND4_1%C
x_PM_SKY130_FD_SC_LS__AND4_1%D N_D_M1001_g N_D_c_200_n N_D_c_201_n N_D_M1000_g D
+ N_D_c_198_n N_D_c_199_n PM_SKY130_FD_SC_LS__AND4_1%D
x_PM_SKY130_FD_SC_LS__AND4_1%A_96_74# N_A_96_74#_M1007_s N_A_96_74#_M1005_d
+ N_A_96_74#_M1009_d N_A_96_74#_M1002_g N_A_96_74#_c_244_n N_A_96_74#_M1004_g
+ N_A_96_74#_c_245_n N_A_96_74#_c_251_n N_A_96_74#_c_252_n N_A_96_74#_c_253_n
+ N_A_96_74#_c_254_n N_A_96_74#_c_255_n N_A_96_74#_c_256_n N_A_96_74#_c_246_n
+ N_A_96_74#_c_247_n N_A_96_74#_c_258_n N_A_96_74#_c_259_n N_A_96_74#_c_248_n
+ PM_SKY130_FD_SC_LS__AND4_1%A_96_74#
x_PM_SKY130_FD_SC_LS__AND4_1%VPWR N_VPWR_M1005_s N_VPWR_M1003_d N_VPWR_M1000_d
+ N_VPWR_c_340_n N_VPWR_c_341_n N_VPWR_c_342_n N_VPWR_c_343_n VPWR
+ N_VPWR_c_344_n N_VPWR_c_345_n N_VPWR_c_346_n N_VPWR_c_339_n N_VPWR_c_348_n
+ N_VPWR_c_349_n PM_SKY130_FD_SC_LS__AND4_1%VPWR
x_PM_SKY130_FD_SC_LS__AND4_1%X N_X_M1002_d N_X_M1004_d N_X_c_389_n N_X_c_390_n
+ N_X_c_387_n X X N_X_c_388_n PM_SKY130_FD_SC_LS__AND4_1%X
x_PM_SKY130_FD_SC_LS__AND4_1%VGND N_VGND_M1001_d N_VGND_c_413_n N_VGND_c_414_n
+ N_VGND_c_415_n VGND N_VGND_c_416_n N_VGND_c_417_n
+ PM_SKY130_FD_SC_LS__AND4_1%VGND
cc_1 VNB N_A_c_71_n 0.0197349f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=1.085
cc_2 VNB N_A_c_72_n 0.0283042f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=1.235
cc_3 VNB N_A_c_73_n 0.00242775f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.79
cc_4 VNB N_A_c_74_n 0.0285305f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.285
cc_5 VNB N_A_c_75_n 0.00270112f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.285
cc_6 VNB N_B_M1008_g 0.0311068f $X=-0.19 $Y=-0.245 $X2=0.82 $Y2=0.69
cc_7 VNB B 0.00634804f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=1.085
cc_8 VNB N_B_c_113_n 0.0192404f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.285
cc_9 VNB N_C_c_153_n 0.018087f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=1.085
cc_10 VNB N_C_c_154_n 0.0233773f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=1.235
cc_11 VNB N_C_c_155_n 0.00238742f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.625
cc_12 VNB C 0.00115257f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.79
cc_13 VNB N_C_c_157_n 0.0167979f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_D_M1001_g 0.0315323f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=2.045
cc_15 VNB N_D_c_198_n 0.0243034f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.79
cc_16 VNB N_D_c_199_n 0.00563353f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_17 VNB N_A_96_74#_M1002_g 0.0299488f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.625
cc_18 VNB N_A_96_74#_c_244_n 0.0336591f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_19 VNB N_A_96_74#_c_245_n 0.0343689f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.285
cc_20 VNB N_A_96_74#_c_246_n 2.32711e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_96_74#_c_247_n 0.046163f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_96_74#_c_248_n 0.00358525f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VPWR_c_339_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_X_c_387_n 0.0252035f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_25 VNB N_X_c_388_n 0.0501995f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.285
cc_26 VNB N_VGND_c_413_n 0.007389f $X=-0.19 $Y=-0.245 $X2=0.82 $Y2=1.085
cc_27 VNB N_VGND_c_414_n 0.0630343f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.235
cc_28 VNB N_VGND_c_415_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=1.085
cc_29 VNB N_VGND_c_416_n 0.0236772f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.285
cc_30 VNB N_VGND_c_417_n 0.22352f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VPB N_A_c_76_n 0.0102912f $X=-0.19 $Y=1.66 $X2=0.555 $Y2=1.955
cc_32 VPB N_A_c_77_n 0.0235434f $X=-0.19 $Y=1.66 $X2=0.555 $Y2=2.045
cc_33 VPB N_A_c_73_n 0.0132698f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.79
cc_34 VPB N_A_c_75_n 0.00279274f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.285
cc_35 VPB N_B_c_114_n 0.00996873f $X=-0.19 $Y=1.66 $X2=0.555 $Y2=1.955
cc_36 VPB N_B_c_115_n 0.0225719f $X=-0.19 $Y=1.66 $X2=0.555 $Y2=2.045
cc_37 VPB B 0.00158699f $X=-0.19 $Y=1.66 $X2=0.66 $Y2=1.085
cc_38 VPB N_B_c_113_n 0.0151864f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.285
cc_39 VPB N_C_c_158_n 0.0109023f $X=-0.19 $Y=1.66 $X2=0.555 $Y2=2.54
cc_40 VPB N_C_c_159_n 0.0225453f $X=-0.19 $Y=1.66 $X2=0.82 $Y2=1.085
cc_41 VPB N_C_c_155_n 0.0135871f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.625
cc_42 VPB C 0.00144048f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.79
cc_43 VPB N_D_c_200_n 0.0161825f $X=-0.19 $Y=1.66 $X2=0.82 $Y2=1.085
cc_44 VPB N_D_c_201_n 0.0221675f $X=-0.19 $Y=1.66 $X2=0.82 $Y2=0.69
cc_45 VPB N_D_c_198_n 0.00560585f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.79
cc_46 VPB N_D_c_199_n 0.00303823f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_47 VPB N_A_96_74#_c_244_n 0.0295996f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_48 VPB N_A_96_74#_c_245_n 0.0152455f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.285
cc_49 VPB N_A_96_74#_c_251_n 0.00623619f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.285
cc_50 VPB N_A_96_74#_c_252_n 0.00928151f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.285
cc_51 VPB N_A_96_74#_c_253_n 0.00289722f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=1.295
cc_52 VPB N_A_96_74#_c_254_n 0.0113743f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=1.665
cc_53 VPB N_A_96_74#_c_255_n 0.00289722f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_A_96_74#_c_256_n 0.00423688f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_A_96_74#_c_246_n 0.00278511f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_A_96_74#_c_258_n 0.0066013f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_A_96_74#_c_259_n 0.00803253f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_340_n 0.0121909f $X=-0.19 $Y=1.66 $X2=0.66 $Y2=1.085
cc_59 VPB N_VPWR_c_341_n 0.0372498f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.625
cc_60 VPB N_VPWR_c_342_n 0.00552382f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_343_n 0.00978361f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.285
cc_62 VPB N_VPWR_c_344_n 0.0185368f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_345_n 0.0196506f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_346_n 0.0190372f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_339_n 0.0600116f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_348_n 0.010962f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_349_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_X_c_389_n 0.0418938f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.235
cc_69 VPB N_X_c_390_n 0.0141454f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_70 VPB N_X_c_387_n 0.00756817f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_71 N_A_c_77_n N_B_c_114_n 0.00553917f $X=0.555 $Y=2.045 $X2=0 $Y2=0
cc_72 N_A_c_77_n N_B_c_115_n 0.0196664f $X=0.555 $Y=2.045 $X2=0 $Y2=0
cc_73 N_A_c_71_n N_B_M1008_g 0.050914f $X=0.66 $Y=1.085 $X2=0 $Y2=0
cc_74 N_A_c_74_n N_B_M1008_g 0.00716063f $X=0.59 $Y=1.285 $X2=0 $Y2=0
cc_75 N_A_c_75_n N_B_M1008_g 7.58023e-19 $X=0.59 $Y=1.285 $X2=0 $Y2=0
cc_76 N_A_c_71_n B 0.0088638f $X=0.66 $Y=1.085 $X2=0 $Y2=0
cc_77 N_A_c_74_n B 0.00111998f $X=0.59 $Y=1.285 $X2=0 $Y2=0
cc_78 N_A_c_75_n B 0.0547116f $X=0.59 $Y=1.285 $X2=0 $Y2=0
cc_79 N_A_c_76_n N_B_c_113_n 0.00553917f $X=0.555 $Y=1.955 $X2=0 $Y2=0
cc_80 N_A_c_74_n N_B_c_113_n 0.0196867f $X=0.59 $Y=1.285 $X2=0 $Y2=0
cc_81 N_A_c_75_n N_B_c_113_n 0.00189366f $X=0.59 $Y=1.285 $X2=0 $Y2=0
cc_82 N_A_c_76_n N_A_96_74#_c_245_n 0.00614356f $X=0.555 $Y=1.955 $X2=0 $Y2=0
cc_83 N_A_c_71_n N_A_96_74#_c_245_n 0.00256672f $X=0.66 $Y=1.085 $X2=0 $Y2=0
cc_84 N_A_c_72_n N_A_96_74#_c_245_n 0.016551f $X=0.66 $Y=1.235 $X2=0 $Y2=0
cc_85 N_A_c_75_n N_A_96_74#_c_245_n 0.0509289f $X=0.59 $Y=1.285 $X2=0 $Y2=0
cc_86 N_A_c_77_n N_A_96_74#_c_251_n 0.0140657f $X=0.555 $Y=2.045 $X2=0 $Y2=0
cc_87 N_A_c_73_n N_A_96_74#_c_251_n 2.66536e-19 $X=0.59 $Y=1.79 $X2=0 $Y2=0
cc_88 N_A_c_75_n N_A_96_74#_c_251_n 0.0135474f $X=0.59 $Y=1.285 $X2=0 $Y2=0
cc_89 N_A_c_77_n N_A_96_74#_c_253_n 0.0159605f $X=0.555 $Y=2.045 $X2=0 $Y2=0
cc_90 N_A_c_71_n N_A_96_74#_c_247_n 0.00816713f $X=0.66 $Y=1.085 $X2=0 $Y2=0
cc_91 N_A_c_72_n N_A_96_74#_c_247_n 0.00885728f $X=0.66 $Y=1.235 $X2=0 $Y2=0
cc_92 N_A_c_75_n N_A_96_74#_c_247_n 0.0270622f $X=0.59 $Y=1.285 $X2=0 $Y2=0
cc_93 N_A_c_77_n N_A_96_74#_c_258_n 0.00309497f $X=0.555 $Y=2.045 $X2=0 $Y2=0
cc_94 N_A_c_73_n N_A_96_74#_c_258_n 8.51503e-19 $X=0.59 $Y=1.79 $X2=0 $Y2=0
cc_95 N_A_c_75_n N_A_96_74#_c_258_n 0.0167547f $X=0.59 $Y=1.285 $X2=0 $Y2=0
cc_96 N_A_c_77_n N_VPWR_c_341_n 0.0163913f $X=0.555 $Y=2.045 $X2=0 $Y2=0
cc_97 N_A_c_77_n N_VPWR_c_342_n 5.64706e-19 $X=0.555 $Y=2.045 $X2=0 $Y2=0
cc_98 N_A_c_77_n N_VPWR_c_344_n 0.00445602f $X=0.555 $Y=2.045 $X2=0 $Y2=0
cc_99 N_A_c_77_n N_VPWR_c_339_n 0.00861081f $X=0.555 $Y=2.045 $X2=0 $Y2=0
cc_100 N_A_c_71_n N_VGND_c_414_n 0.00433274f $X=0.66 $Y=1.085 $X2=0 $Y2=0
cc_101 N_A_c_71_n N_VGND_c_417_n 0.00822417f $X=0.66 $Y=1.085 $X2=0 $Y2=0
cc_102 N_B_c_114_n N_C_c_158_n 0.00306838f $X=1.055 $Y=1.955 $X2=0 $Y2=0
cc_103 N_B_c_113_n N_C_c_158_n 5.46201e-19 $X=1.15 $Y=1.64 $X2=0 $Y2=0
cc_104 N_B_c_115_n N_C_c_159_n 0.0212619f $X=1.055 $Y=2.045 $X2=0 $Y2=0
cc_105 N_B_M1008_g N_C_c_153_n 0.0643574f $X=1.21 $Y=0.69 $X2=0 $Y2=0
cc_106 B N_C_c_153_n 0.00429553f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_107 B N_C_c_154_n 0.00109427f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_108 N_B_c_113_n N_C_c_154_n 0.0192516f $X=1.15 $Y=1.64 $X2=0 $Y2=0
cc_109 N_B_M1008_g C 0.00126134f $X=1.21 $Y=0.69 $X2=0 $Y2=0
cc_110 B C 0.0693141f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_111 N_B_c_113_n C 0.0011086f $X=1.15 $Y=1.64 $X2=0 $Y2=0
cc_112 N_B_c_115_n N_A_96_74#_c_253_n 0.00450743f $X=1.055 $Y=2.045 $X2=0 $Y2=0
cc_113 N_B_c_115_n N_A_96_74#_c_254_n 0.0176436f $X=1.055 $Y=2.045 $X2=0 $Y2=0
cc_114 B N_A_96_74#_c_254_n 0.0256177f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_115 N_B_c_113_n N_A_96_74#_c_254_n 0.00117818f $X=1.15 $Y=1.64 $X2=0 $Y2=0
cc_116 N_B_M1008_g N_A_96_74#_c_247_n 8.33395e-19 $X=1.21 $Y=0.69 $X2=0 $Y2=0
cc_117 B N_A_96_74#_c_247_n 0.0349867f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_118 N_B_c_115_n N_VPWR_c_342_n 0.0234691f $X=1.055 $Y=2.045 $X2=0 $Y2=0
cc_119 N_B_c_115_n N_VPWR_c_344_n 0.00413917f $X=1.055 $Y=2.045 $X2=0 $Y2=0
cc_120 N_B_c_115_n N_VPWR_c_339_n 0.00818241f $X=1.055 $Y=2.045 $X2=0 $Y2=0
cc_121 B A_179_74# 0.00666137f $X=1.115 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_122 N_B_M1008_g N_VGND_c_414_n 0.00303293f $X=1.21 $Y=0.69 $X2=0 $Y2=0
cc_123 B N_VGND_c_414_n 0.00887369f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_124 N_B_M1008_g N_VGND_c_417_n 0.003711f $X=1.21 $Y=0.69 $X2=0 $Y2=0
cc_125 B N_VGND_c_417_n 0.0106888f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_126 N_C_c_153_n N_D_M1001_g 0.0217572f $X=1.69 $Y=1.12 $X2=0 $Y2=0
cc_127 C N_D_M1001_g 0.00862137f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_128 N_C_c_157_n N_D_M1001_g 0.0127959f $X=1.69 $Y=1.285 $X2=0 $Y2=0
cc_129 N_C_c_155_n N_D_c_200_n 0.00748003f $X=1.69 $Y=1.79 $X2=0 $Y2=0
cc_130 N_C_c_158_n N_D_c_201_n 0.00748003f $X=1.765 $Y=1.955 $X2=0 $Y2=0
cc_131 N_C_c_159_n N_D_c_201_n 0.0196951f $X=1.765 $Y=2.045 $X2=0 $Y2=0
cc_132 N_C_c_154_n N_D_c_198_n 0.0206633f $X=1.69 $Y=1.625 $X2=0 $Y2=0
cc_133 C N_D_c_198_n 3.98767e-19 $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_134 N_C_c_154_n N_D_c_199_n 0.00259302f $X=1.69 $Y=1.625 $X2=0 $Y2=0
cc_135 C N_D_c_199_n 0.0314204f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_136 N_C_c_159_n N_A_96_74#_c_254_n 0.0171489f $X=1.765 $Y=2.045 $X2=0 $Y2=0
cc_137 N_C_c_155_n N_A_96_74#_c_254_n 0.00101795f $X=1.69 $Y=1.79 $X2=0 $Y2=0
cc_138 C N_A_96_74#_c_254_n 0.023903f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_139 N_C_c_159_n N_A_96_74#_c_255_n 0.00450743f $X=1.765 $Y=2.045 $X2=0 $Y2=0
cc_140 N_C_c_159_n N_A_96_74#_c_259_n 5.07271e-19 $X=1.765 $Y=2.045 $X2=0 $Y2=0
cc_141 N_C_c_159_n N_VPWR_c_342_n 0.0235524f $X=1.765 $Y=2.045 $X2=0 $Y2=0
cc_142 N_C_c_159_n N_VPWR_c_345_n 0.00413917f $X=1.765 $Y=2.045 $X2=0 $Y2=0
cc_143 N_C_c_159_n N_VPWR_c_339_n 0.00818241f $X=1.765 $Y=2.045 $X2=0 $Y2=0
cc_144 C A_335_74# 0.00857283f $X=1.595 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_145 N_C_c_153_n N_VGND_c_413_n 0.00143141f $X=1.69 $Y=1.12 $X2=0 $Y2=0
cc_146 C N_VGND_c_413_n 0.025502f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_147 N_C_c_153_n N_VGND_c_414_n 0.00304348f $X=1.69 $Y=1.12 $X2=0 $Y2=0
cc_148 C N_VGND_c_414_n 0.00930091f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_149 N_C_c_153_n N_VGND_c_417_n 0.00371612f $X=1.69 $Y=1.12 $X2=0 $Y2=0
cc_150 C N_VGND_c_417_n 0.0106938f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_151 N_D_M1001_g N_A_96_74#_M1002_g 0.0240727f $X=2.17 $Y=0.69 $X2=0 $Y2=0
cc_152 N_D_c_200_n N_A_96_74#_c_244_n 0.00781309f $X=2.265 $Y=1.955 $X2=0 $Y2=0
cc_153 N_D_c_201_n N_A_96_74#_c_244_n 0.0201473f $X=2.265 $Y=2.045 $X2=0 $Y2=0
cc_154 N_D_c_198_n N_A_96_74#_c_244_n 0.0195574f $X=2.23 $Y=1.515 $X2=0 $Y2=0
cc_155 N_D_c_199_n N_A_96_74#_c_244_n 3.48015e-19 $X=2.23 $Y=1.515 $X2=0 $Y2=0
cc_156 N_D_c_201_n N_A_96_74#_c_255_n 0.0123377f $X=2.265 $Y=2.045 $X2=0 $Y2=0
cc_157 N_D_c_201_n N_A_96_74#_c_256_n 0.0129378f $X=2.265 $Y=2.045 $X2=0 $Y2=0
cc_158 N_D_c_198_n N_A_96_74#_c_256_n 2.11278e-19 $X=2.23 $Y=1.515 $X2=0 $Y2=0
cc_159 N_D_c_199_n N_A_96_74#_c_256_n 0.0135189f $X=2.23 $Y=1.515 $X2=0 $Y2=0
cc_160 N_D_c_200_n N_A_96_74#_c_246_n 0.00409025f $X=2.265 $Y=1.955 $X2=0 $Y2=0
cc_161 N_D_c_198_n N_A_96_74#_c_246_n 2.16901e-19 $X=2.23 $Y=1.515 $X2=0 $Y2=0
cc_162 N_D_c_199_n N_A_96_74#_c_246_n 0.0100188f $X=2.23 $Y=1.515 $X2=0 $Y2=0
cc_163 N_D_c_201_n N_A_96_74#_c_259_n 0.00360435f $X=2.265 $Y=2.045 $X2=0 $Y2=0
cc_164 N_D_c_198_n N_A_96_74#_c_259_n 6.70927e-19 $X=2.23 $Y=1.515 $X2=0 $Y2=0
cc_165 N_D_c_199_n N_A_96_74#_c_259_n 0.0135593f $X=2.23 $Y=1.515 $X2=0 $Y2=0
cc_166 N_D_M1001_g N_A_96_74#_c_248_n 5.96922e-19 $X=2.17 $Y=0.69 $X2=0 $Y2=0
cc_167 N_D_c_198_n N_A_96_74#_c_248_n 0.0017071f $X=2.23 $Y=1.515 $X2=0 $Y2=0
cc_168 N_D_c_199_n N_A_96_74#_c_248_n 0.0235504f $X=2.23 $Y=1.515 $X2=0 $Y2=0
cc_169 N_D_c_201_n N_VPWR_c_342_n 7.45467e-19 $X=2.265 $Y=2.045 $X2=0 $Y2=0
cc_170 N_D_c_201_n N_VPWR_c_343_n 0.0096747f $X=2.265 $Y=2.045 $X2=0 $Y2=0
cc_171 N_D_c_201_n N_VPWR_c_345_n 0.00445602f $X=2.265 $Y=2.045 $X2=0 $Y2=0
cc_172 N_D_c_201_n N_VPWR_c_339_n 0.00859378f $X=2.265 $Y=2.045 $X2=0 $Y2=0
cc_173 N_D_c_201_n N_X_c_389_n 9.39142e-19 $X=2.265 $Y=2.045 $X2=0 $Y2=0
cc_174 N_D_M1001_g N_X_c_388_n 6.48878e-19 $X=2.17 $Y=0.69 $X2=0 $Y2=0
cc_175 N_D_M1001_g N_VGND_c_413_n 0.015634f $X=2.17 $Y=0.69 $X2=0 $Y2=0
cc_176 N_D_c_198_n N_VGND_c_413_n 0.00108304f $X=2.23 $Y=1.515 $X2=0 $Y2=0
cc_177 N_D_c_199_n N_VGND_c_413_n 0.00911635f $X=2.23 $Y=1.515 $X2=0 $Y2=0
cc_178 N_D_M1001_g N_VGND_c_414_n 0.00383152f $X=2.17 $Y=0.69 $X2=0 $Y2=0
cc_179 N_D_M1001_g N_VGND_c_417_n 0.00758792f $X=2.17 $Y=0.69 $X2=0 $Y2=0
cc_180 N_A_96_74#_c_251_n N_VPWR_M1005_s 0.00181377f $X=0.615 $Y=2.06 $X2=-0.19
+ $Y2=-0.245
cc_181 N_A_96_74#_c_252_n N_VPWR_M1005_s 0.001494f $X=0.255 $Y=2.06 $X2=-0.19
+ $Y2=-0.245
cc_182 N_A_96_74#_c_254_n N_VPWR_M1003_d 0.0049669f $X=1.875 $Y=2.06 $X2=0 $Y2=0
cc_183 N_A_96_74#_c_256_n N_VPWR_M1000_d 0.00778325f $X=2.57 $Y=2.045 $X2=0
+ $Y2=0
cc_184 N_A_96_74#_c_246_n N_VPWR_M1000_d 0.00239047f $X=2.655 $Y=1.96 $X2=0
+ $Y2=0
cc_185 N_A_96_74#_c_251_n N_VPWR_c_341_n 0.0136318f $X=0.615 $Y=2.06 $X2=0 $Y2=0
cc_186 N_A_96_74#_c_252_n N_VPWR_c_341_n 0.0125997f $X=0.255 $Y=2.06 $X2=0 $Y2=0
cc_187 N_A_96_74#_c_253_n N_VPWR_c_341_n 0.0257429f $X=0.78 $Y=2.28 $X2=0 $Y2=0
cc_188 N_A_96_74#_c_253_n N_VPWR_c_342_n 0.0280607f $X=0.78 $Y=2.28 $X2=0 $Y2=0
cc_189 N_A_96_74#_c_254_n N_VPWR_c_342_n 0.0384188f $X=1.875 $Y=2.06 $X2=0 $Y2=0
cc_190 N_A_96_74#_c_255_n N_VPWR_c_342_n 0.0280607f $X=2.04 $Y=2.28 $X2=0 $Y2=0
cc_191 N_A_96_74#_c_244_n N_VPWR_c_343_n 0.00803019f $X=2.85 $Y=1.765 $X2=0
+ $Y2=0
cc_192 N_A_96_74#_c_255_n N_VPWR_c_343_n 0.0457344f $X=2.04 $Y=2.28 $X2=0 $Y2=0
cc_193 N_A_96_74#_c_256_n N_VPWR_c_343_n 0.0258647f $X=2.57 $Y=2.045 $X2=0 $Y2=0
cc_194 N_A_96_74#_c_253_n N_VPWR_c_344_n 0.0145938f $X=0.78 $Y=2.28 $X2=0 $Y2=0
cc_195 N_A_96_74#_c_255_n N_VPWR_c_345_n 0.0145938f $X=2.04 $Y=2.28 $X2=0 $Y2=0
cc_196 N_A_96_74#_c_244_n N_VPWR_c_346_n 0.00445602f $X=2.85 $Y=1.765 $X2=0
+ $Y2=0
cc_197 N_A_96_74#_c_244_n N_VPWR_c_339_n 0.0086159f $X=2.85 $Y=1.765 $X2=0 $Y2=0
cc_198 N_A_96_74#_c_253_n N_VPWR_c_339_n 0.0120466f $X=0.78 $Y=2.28 $X2=0 $Y2=0
cc_199 N_A_96_74#_c_255_n N_VPWR_c_339_n 0.0120466f $X=2.04 $Y=2.28 $X2=0 $Y2=0
cc_200 N_A_96_74#_c_244_n N_X_c_389_n 0.0127662f $X=2.85 $Y=1.765 $X2=0 $Y2=0
cc_201 N_A_96_74#_c_244_n N_X_c_390_n 0.00288786f $X=2.85 $Y=1.765 $X2=0 $Y2=0
cc_202 N_A_96_74#_c_246_n N_X_c_390_n 0.00604965f $X=2.655 $Y=1.96 $X2=0 $Y2=0
cc_203 N_A_96_74#_c_248_n N_X_c_390_n 0.00196075f $X=2.77 $Y=1.485 $X2=0 $Y2=0
cc_204 N_A_96_74#_M1002_g N_X_c_387_n 0.00394404f $X=2.68 $Y=0.74 $X2=0 $Y2=0
cc_205 N_A_96_74#_c_244_n N_X_c_387_n 0.0101214f $X=2.85 $Y=1.765 $X2=0 $Y2=0
cc_206 N_A_96_74#_c_246_n N_X_c_387_n 0.00530743f $X=2.655 $Y=1.96 $X2=0 $Y2=0
cc_207 N_A_96_74#_c_248_n N_X_c_387_n 0.0249641f $X=2.77 $Y=1.485 $X2=0 $Y2=0
cc_208 N_A_96_74#_M1002_g N_X_c_388_n 0.0120059f $X=2.68 $Y=0.74 $X2=0 $Y2=0
cc_209 N_A_96_74#_c_244_n N_X_c_388_n 0.00498973f $X=2.85 $Y=1.765 $X2=0 $Y2=0
cc_210 N_A_96_74#_c_248_n N_X_c_388_n 0.0157141f $X=2.77 $Y=1.485 $X2=0 $Y2=0
cc_211 N_A_96_74#_M1002_g N_VGND_c_413_n 0.00668894f $X=2.68 $Y=0.74 $X2=0 $Y2=0
cc_212 N_A_96_74#_c_247_n N_VGND_c_414_n 0.0294787f $X=0.605 $Y=0.515 $X2=0
+ $Y2=0
cc_213 N_A_96_74#_M1002_g N_VGND_c_416_n 0.00434272f $X=2.68 $Y=0.74 $X2=0 $Y2=0
cc_214 N_A_96_74#_M1002_g N_VGND_c_417_n 0.00825221f $X=2.68 $Y=0.74 $X2=0 $Y2=0
cc_215 N_A_96_74#_c_247_n N_VGND_c_417_n 0.0249691f $X=0.605 $Y=0.515 $X2=0
+ $Y2=0
cc_216 N_VPWR_c_343_n N_X_c_389_n 0.0267024f $X=2.575 $Y=2.465 $X2=0 $Y2=0
cc_217 N_VPWR_c_346_n N_X_c_389_n 0.0161555f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_218 N_VPWR_c_339_n N_X_c_389_n 0.0133393f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_219 N_X_c_388_n N_VGND_c_413_n 0.0270745f $X=2.895 $Y=0.515 $X2=0 $Y2=0
cc_220 N_X_c_388_n N_VGND_c_416_n 0.0241574f $X=2.895 $Y=0.515 $X2=0 $Y2=0
cc_221 N_X_c_388_n N_VGND_c_417_n 0.019939f $X=2.895 $Y=0.515 $X2=0 $Y2=0
