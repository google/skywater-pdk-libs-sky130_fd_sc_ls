* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
M1000 a_233_384# A1_N VPWR VPB phighvt w=840000u l=150000u
+  ad=2.982e+11p pd=2.39e+06u as=1.704e+12p ps=9.65e+06u
M1001 VPWR A2_N a_233_384# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 VGND a_83_260# X VNB nshort w=740000u l=150000u
+  ad=6.211e+11p pd=4.59e+06u as=2.109e+11p ps=2.05e+06u
M1003 a_253_94# A1_N VGND VNB nshort w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1004 a_233_384# A2_N a_253_94# VNB nshort w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=0p ps=0u
M1005 a_588_74# a_233_384# a_83_260# VNB nshort w=640000u l=150000u
+  ad=3.616e+11p pd=3.69e+06u as=1.824e+11p ps=1.85e+06u
M1006 VPWR B1 a_693_384# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1007 VPWR a_83_260# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.304e+11p ps=2.83e+06u
M1008 a_83_260# a_233_384# VPWR VPB phighvt w=840000u l=150000u
+  ad=3.448e+11p pd=2.72e+06u as=0p ps=0u
M1009 a_693_384# B2 a_83_260# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_588_74# B1 VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND B2 a_588_74# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
