* File: sky130_fd_sc_ls__maj3_1.spice
* Created: Wed Sep  2 11:09:48 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__maj3_1.pex.spice"
.subckt sky130_fd_sc_ls__maj3_1  VNB VPB B C A X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A	A
* C	C
* B	B
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_A_84_74#_M1003_g N_X_M1003_s VNB NSHORT L=0.15 W=0.74
+ AD=0.148965 AS=0.2081 PD=1.21725 PS=2.05 NRD=14.592 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75002.4 A=0.111 P=1.78 MULT=1
MM1012 A_223_120# N_A_M1012_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.64 AD=0.0768
+ AS=0.128835 PD=0.88 PS=1.05275 NRD=12.18 NRS=4.68 M=1 R=4.26667 SA=75000.8
+ SB=75002.2 A=0.096 P=1.58 MULT=1
MM1004 N_A_84_74#_M1004_d N_B_M1004_g A_223_120# VNB NSHORT L=0.15 W=0.64
+ AD=0.1222 AS=0.0768 PD=1.08 PS=0.88 NRD=0 NRS=12.18 M=1 R=4.26667 SA=75001.1
+ SB=75001.9 A=0.096 P=1.58 MULT=1
MM1013 A_403_136# N_B_M1013_g N_A_84_74#_M1004_d VNB NSHORT L=0.15 W=0.64
+ AD=0.0768 AS=0.1222 PD=0.88 PS=1.08 NRD=12.18 NRS=15.468 M=1 R=4.26667
+ SA=75001.5 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1007 N_VGND_M1007_d N_C_M1007_g A_403_136# VNB NSHORT L=0.15 W=0.64 AD=0.1344
+ AS=0.0768 PD=1.06 PS=0.88 NRD=13.116 NRS=12.18 M=1 R=4.26667 SA=75001.9
+ SB=75001.2 A=0.096 P=1.58 MULT=1
MM1005 A_595_136# N_A_M1005_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.64 AD=0.0864
+ AS=0.1344 PD=0.91 PS=1.06 NRD=15 NRS=13.116 M=1 R=4.26667 SA=75002.4
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1008 N_A_84_74#_M1008_d N_C_M1008_g A_595_136# VNB NSHORT L=0.15 W=0.64
+ AD=0.1733 AS=0.0864 PD=1.85 PS=0.91 NRD=0 NRS=15 M=1 R=4.26667 SA=75002.8
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1009 N_VPWR_M1009_d N_A_84_74#_M1009_g N_X_M1009_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.204347 AS=0.3304 PD=1.55849 PS=2.83 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75002.7 A=0.168 P=2.54 MULT=1
MM1002 A_226_384# N_A_M1002_g N_VPWR_M1009_d VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.182453 PD=1.27 PS=1.39151 NRD=15.7403 NRS=2.9353 M=1 R=6.66667 SA=75000.7
+ SB=75002.5 A=0.15 P=2.3 MULT=1
MM1001 N_A_84_74#_M1001_d N_B_M1001_g A_226_384# VPB PHIGHVT L=0.15 W=1 AD=0.165
+ AS=0.135 PD=1.33 PS=1.27 NRD=7.8603 NRS=15.7403 M=1 R=6.66667 SA=75001.1
+ SB=75002.1 A=0.15 P=2.3 MULT=1
MM1010 A_406_384# N_B_M1010_g N_A_84_74#_M1001_d VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.165 PD=1.27 PS=1.33 NRD=15.7403 NRS=1.9503 M=1 R=6.66667 SA=75001.6
+ SB=75001.6 A=0.15 P=2.3 MULT=1
MM1006 N_VPWR_M1006_d N_C_M1006_g A_406_384# VPB PHIGHVT L=0.15 W=1 AD=0.195
+ AS=0.135 PD=1.39 PS=1.27 NRD=9.8303 NRS=15.7403 M=1 R=6.66667 SA=75002
+ SB=75001.2 A=0.15 P=2.3 MULT=1
MM1000 A_598_384# N_A_M1000_g N_VPWR_M1006_d VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.195 PD=1.27 PS=1.39 NRD=15.7403 NRS=11.8003 M=1 R=6.66667 SA=75002.6
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1011 N_A_84_74#_M1011_d N_C_M1011_g A_598_384# VPB PHIGHVT L=0.15 W=1 AD=0.295
+ AS=0.135 PD=2.59 PS=1.27 NRD=1.9503 NRS=15.7403 M=1 R=6.66667 SA=75003
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX14_noxref VNB VPB NWDIODE A=7.8492 P=12.16
*
.include "sky130_fd_sc_ls__maj3_1.pxi.spice"
*
.ends
*
*
