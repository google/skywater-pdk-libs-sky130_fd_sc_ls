* File: sky130_fd_sc_ls__nand3b_2.pxi.spice
* Created: Wed Sep  2 11:12:34 2020
* 
x_PM_SKY130_FD_SC_LS__NAND3B_2%A_N N_A_N_M1003_g N_A_N_c_74_n N_A_N_M1002_g A_N
+ N_A_N_c_72_n N_A_N_c_73_n PM_SKY130_FD_SC_LS__NAND3B_2%A_N
x_PM_SKY130_FD_SC_LS__NAND3B_2%C N_C_c_104_n N_C_M1001_g N_C_c_108_n N_C_M1000_g
+ N_C_c_105_n N_C_M1007_g N_C_c_109_n N_C_M1006_g C C N_C_c_107_n
+ PM_SKY130_FD_SC_LS__NAND3B_2%C
x_PM_SKY130_FD_SC_LS__NAND3B_2%A_27_94# N_A_27_94#_M1003_s N_A_27_94#_M1002_s
+ N_A_27_94#_c_174_n N_A_27_94#_M1008_g N_A_27_94#_c_165_n N_A_27_94#_M1004_g
+ N_A_27_94#_c_175_n N_A_27_94#_M1012_g N_A_27_94#_M1005_g N_A_27_94#_c_167_n
+ N_A_27_94#_c_176_n N_A_27_94#_c_168_n N_A_27_94#_c_169_n N_A_27_94#_c_170_n
+ N_A_27_94#_c_171_n N_A_27_94#_c_178_n N_A_27_94#_c_207_n N_A_27_94#_c_172_n
+ N_A_27_94#_c_173_n PM_SKY130_FD_SC_LS__NAND3B_2%A_27_94#
x_PM_SKY130_FD_SC_LS__NAND3B_2%B N_B_c_281_n N_B_M1010_g N_B_c_277_n N_B_M1009_g
+ N_B_c_282_n N_B_M1013_g N_B_c_278_n N_B_M1011_g B B B N_B_c_280_n
+ PM_SKY130_FD_SC_LS__NAND3B_2%B
x_PM_SKY130_FD_SC_LS__NAND3B_2%VPWR N_VPWR_M1002_d N_VPWR_M1006_s N_VPWR_M1012_s
+ N_VPWR_M1013_s N_VPWR_c_321_n N_VPWR_c_322_n N_VPWR_c_323_n N_VPWR_c_324_n
+ N_VPWR_c_325_n N_VPWR_c_326_n N_VPWR_c_327_n N_VPWR_c_328_n N_VPWR_c_329_n
+ N_VPWR_c_330_n N_VPWR_c_331_n VPWR N_VPWR_c_332_n N_VPWR_c_320_n
+ PM_SKY130_FD_SC_LS__NAND3B_2%VPWR
x_PM_SKY130_FD_SC_LS__NAND3B_2%Y N_Y_M1004_d N_Y_M1000_d N_Y_M1008_d N_Y_M1010_d
+ N_Y_c_388_n N_Y_c_383_n N_Y_c_394_n N_Y_c_384_n N_Y_c_404_n N_Y_c_405_n
+ N_Y_c_420_n N_Y_c_385_n N_Y_c_408_n Y PM_SKY130_FD_SC_LS__NAND3B_2%Y
x_PM_SKY130_FD_SC_LS__NAND3B_2%VGND N_VGND_M1003_d N_VGND_M1007_s N_VGND_c_449_n
+ N_VGND_c_450_n VGND N_VGND_c_451_n N_VGND_c_452_n N_VGND_c_453_n
+ N_VGND_c_454_n N_VGND_c_455_n N_VGND_c_456_n PM_SKY130_FD_SC_LS__NAND3B_2%VGND
x_PM_SKY130_FD_SC_LS__NAND3B_2%A_206_74# N_A_206_74#_M1001_d N_A_206_74#_M1009_d
+ N_A_206_74#_c_498_n N_A_206_74#_c_495_n N_A_206_74#_c_496_n
+ N_A_206_74#_c_497_n N_A_206_74#_c_515_n N_A_206_74#_c_511_n
+ PM_SKY130_FD_SC_LS__NAND3B_2%A_206_74#
x_PM_SKY130_FD_SC_LS__NAND3B_2%A_403_54# N_A_403_54#_M1004_s N_A_403_54#_M1005_s
+ N_A_403_54#_M1011_s N_A_403_54#_c_537_n N_A_403_54#_c_538_n
+ PM_SKY130_FD_SC_LS__NAND3B_2%A_403_54#
cc_1 VNB N_A_N_M1003_g 0.0391626f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=0.79
cc_2 VNB N_A_N_c_72_n 0.00895418f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_3 VNB N_A_N_c_73_n 0.0306339f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=1.667
cc_4 VNB N_C_c_104_n 0.0152719f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=1.45
cc_5 VNB N_C_c_105_n 0.0171557f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=2.46
cc_6 VNB C 0.00358799f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=1.667
cc_7 VNB N_C_c_107_n 0.0794831f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_27_94#_c_165_n 0.0182994f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.667
cc_9 VNB N_A_27_94#_M1005_g 0.0185822f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_10 VNB N_A_27_94#_c_167_n 0.0266041f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_27_94#_c_168_n 0.0022042f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_94#_c_169_n 0.0104221f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_94#_c_170_n 0.00531239f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_94#_c_171_n 0.0110158f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_94#_c_172_n 0.00729475f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_27_94#_c_173_n 0.0492544f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_B_c_277_n 0.0165885f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_B_c_278_n 0.0205306f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.667
cc_19 VNB B 0.0224642f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.615
cc_20 VNB N_B_c_280_n 0.0402273f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_VPWR_c_320_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB Y 0.00108338f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_449_n 0.0093225f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_450_n 0.0108515f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=1.667
cc_25 VNB N_VGND_c_451_n 0.0174171f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_452_n 0.0166891f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_453_n 0.0644788f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_454_n 0.261576f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_455_n 0.00557808f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_456_n 0.00613127f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_206_74#_c_495_n 0.00214855f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_206_74#_c_496_n 0.00617097f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_206_74#_c_497_n 0.00550897f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_34 VNB N_A_403_54#_c_537_n 0.0324263f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.667
cc_35 VNB N_A_403_54#_c_538_n 0.0265018f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_36 VPB N_A_N_c_74_n 0.0211953f $X=-0.19 $Y=1.66 $X2=0.695 $Y2=1.885
cc_37 VPB N_A_N_c_72_n 0.00811757f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.615
cc_38 VPB N_A_N_c_73_n 0.0336147f $X=-0.19 $Y=1.66 $X2=0.48 $Y2=1.667
cc_39 VPB N_C_c_108_n 0.0164949f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_40 VPB N_C_c_109_n 0.0165188f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.667
cc_41 VPB C 0.00716393f $X=-0.19 $Y=1.66 $X2=0.695 $Y2=1.667
cc_42 VPB N_C_c_107_n 0.0209666f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_43 VPB N_A_27_94#_c_174_n 0.0155892f $X=-0.19 $Y=1.66 $X2=0.695 $Y2=2.46
cc_44 VPB N_A_27_94#_c_175_n 0.0164171f $X=-0.19 $Y=1.66 $X2=0.48 $Y2=1.667
cc_45 VPB N_A_27_94#_c_176_n 0.0354741f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_A_27_94#_c_170_n 0.00163525f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB N_A_27_94#_c_178_n 0.00927352f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 VPB N_A_27_94#_c_172_n 0.00180391f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 VPB N_A_27_94#_c_173_n 0.0286473f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_B_c_281_n 0.0175631f $X=-0.19 $Y=1.66 $X2=0.48 $Y2=1.45
cc_51 VPB N_B_c_282_n 0.0192901f $X=-0.19 $Y=1.66 $X2=0.695 $Y2=2.46
cc_52 VPB B 0.0158991f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.615
cc_53 VPB N_B_c_280_n 0.0235574f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_321_n 0.00886591f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.615
cc_55 VPB N_VPWR_c_322_n 0.00595027f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_323_n 0.00916228f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_324_n 0.0120106f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_325_n 0.0489067f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_326_n 0.0259932f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_327_n 0.00468662f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_328_n 0.0202526f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_329_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_330_n 0.0186844f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_331_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_332_n 0.0212417f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_320_n 0.0800232f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_Y_c_383_n 0.0029595f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.615
cc_68 VPB N_Y_c_384_n 0.00216998f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_Y_c_385_n 0.00290527f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB Y 0.00322709f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 N_A_N_M1003_g N_C_c_104_n 0.021804f $X=0.48 $Y=0.79 $X2=-0.19 $Y2=-0.245
cc_72 N_A_N_c_74_n N_C_c_108_n 0.014553f $X=0.695 $Y=1.885 $X2=0 $Y2=0
cc_73 N_A_N_c_73_n N_C_c_108_n 0.00382403f $X=0.48 $Y=1.667 $X2=0 $Y2=0
cc_74 N_A_N_c_73_n C 5.01996e-19 $X=0.48 $Y=1.667 $X2=0 $Y2=0
cc_75 N_A_N_M1003_g N_C_c_107_n 0.00438823f $X=0.48 $Y=0.79 $X2=0 $Y2=0
cc_76 N_A_N_c_73_n N_C_c_107_n 0.00506017f $X=0.48 $Y=1.667 $X2=0 $Y2=0
cc_77 N_A_N_M1003_g N_A_27_94#_c_167_n 4.43891e-19 $X=0.48 $Y=0.79 $X2=0 $Y2=0
cc_78 N_A_N_c_74_n N_A_27_94#_c_176_n 0.0107686f $X=0.695 $Y=1.885 $X2=0 $Y2=0
cc_79 N_A_N_M1003_g N_A_27_94#_c_168_n 0.0157512f $X=0.48 $Y=0.79 $X2=0 $Y2=0
cc_80 N_A_N_c_72_n N_A_27_94#_c_168_n 0.0132391f $X=0.385 $Y=1.615 $X2=0 $Y2=0
cc_81 N_A_N_c_73_n N_A_27_94#_c_168_n 0.00638349f $X=0.48 $Y=1.667 $X2=0 $Y2=0
cc_82 N_A_N_c_72_n N_A_27_94#_c_169_n 0.0178519f $X=0.385 $Y=1.615 $X2=0 $Y2=0
cc_83 N_A_N_c_73_n N_A_27_94#_c_169_n 0.00299816f $X=0.48 $Y=1.667 $X2=0 $Y2=0
cc_84 N_A_N_M1003_g N_A_27_94#_c_170_n 0.00598746f $X=0.48 $Y=0.79 $X2=0 $Y2=0
cc_85 N_A_N_c_74_n N_A_27_94#_c_170_n 0.00339612f $X=0.695 $Y=1.885 $X2=0 $Y2=0
cc_86 N_A_N_c_72_n N_A_27_94#_c_170_n 0.0247013f $X=0.385 $Y=1.615 $X2=0 $Y2=0
cc_87 N_A_N_c_73_n N_A_27_94#_c_170_n 0.0111218f $X=0.48 $Y=1.667 $X2=0 $Y2=0
cc_88 N_A_N_c_74_n N_A_27_94#_c_178_n 0.014186f $X=0.695 $Y=1.885 $X2=0 $Y2=0
cc_89 N_A_N_c_72_n N_A_27_94#_c_178_n 0.0184134f $X=0.385 $Y=1.615 $X2=0 $Y2=0
cc_90 N_A_N_c_73_n N_A_27_94#_c_178_n 0.00871839f $X=0.48 $Y=1.667 $X2=0 $Y2=0
cc_91 N_A_N_c_74_n N_VPWR_c_321_n 0.00531965f $X=0.695 $Y=1.885 $X2=0 $Y2=0
cc_92 N_A_N_c_74_n N_VPWR_c_326_n 0.00445602f $X=0.695 $Y=1.885 $X2=0 $Y2=0
cc_93 N_A_N_c_74_n N_VPWR_c_320_n 0.00862008f $X=0.695 $Y=1.885 $X2=0 $Y2=0
cc_94 N_A_N_c_74_n N_Y_c_383_n 6.154e-19 $X=0.695 $Y=1.885 $X2=0 $Y2=0
cc_95 N_A_N_M1003_g N_VGND_c_449_n 0.0125975f $X=0.48 $Y=0.79 $X2=0 $Y2=0
cc_96 N_A_N_M1003_g N_VGND_c_451_n 0.00421418f $X=0.48 $Y=0.79 $X2=0 $Y2=0
cc_97 N_A_N_M1003_g N_VGND_c_454_n 0.00432128f $X=0.48 $Y=0.79 $X2=0 $Y2=0
cc_98 N_C_c_109_n N_A_27_94#_c_174_n 0.0299722f $X=1.695 $Y=1.765 $X2=0 $Y2=0
cc_99 C N_A_27_94#_c_174_n 3.25855e-19 $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_100 N_C_c_107_n N_A_27_94#_c_165_n 0.00235466f $X=1.615 $Y=1.515 $X2=0 $Y2=0
cc_101 N_C_c_108_n N_A_27_94#_c_176_n 6.25613e-19 $X=1.2 $Y=1.765 $X2=0 $Y2=0
cc_102 N_C_c_108_n N_A_27_94#_c_170_n 0.00341516f $X=1.2 $Y=1.765 $X2=0 $Y2=0
cc_103 C N_A_27_94#_c_170_n 0.0267651f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_104 N_C_c_107_n N_A_27_94#_c_170_n 0.00764977f $X=1.615 $Y=1.515 $X2=0 $Y2=0
cc_105 N_C_c_104_n N_A_27_94#_c_171_n 0.00771139f $X=0.955 $Y=1.185 $X2=0 $Y2=0
cc_106 N_C_c_105_n N_A_27_94#_c_171_n 0.00671798f $X=1.385 $Y=1.185 $X2=0 $Y2=0
cc_107 C N_A_27_94#_c_171_n 0.051126f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_108 N_C_c_107_n N_A_27_94#_c_171_n 0.0310057f $X=1.615 $Y=1.515 $X2=0 $Y2=0
cc_109 N_C_c_108_n N_A_27_94#_c_178_n 0.00147835f $X=1.2 $Y=1.765 $X2=0 $Y2=0
cc_110 N_C_c_104_n N_A_27_94#_c_207_n 0.00184514f $X=0.955 $Y=1.185 $X2=0 $Y2=0
cc_111 N_C_c_107_n N_A_27_94#_c_207_n 0.00108279f $X=1.615 $Y=1.515 $X2=0 $Y2=0
cc_112 C N_A_27_94#_c_172_n 0.0168746f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_113 N_C_c_107_n N_A_27_94#_c_172_n 0.0030545f $X=1.615 $Y=1.515 $X2=0 $Y2=0
cc_114 C N_A_27_94#_c_173_n 0.00306885f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_115 N_C_c_107_n N_A_27_94#_c_173_n 0.0213904f $X=1.615 $Y=1.515 $X2=0 $Y2=0
cc_116 N_C_c_108_n N_VPWR_c_321_n 0.00308391f $X=1.2 $Y=1.765 $X2=0 $Y2=0
cc_117 N_C_c_109_n N_VPWR_c_322_n 0.0068696f $X=1.695 $Y=1.765 $X2=0 $Y2=0
cc_118 N_C_c_108_n N_VPWR_c_328_n 0.00445602f $X=1.2 $Y=1.765 $X2=0 $Y2=0
cc_119 N_C_c_109_n N_VPWR_c_328_n 0.00445602f $X=1.695 $Y=1.765 $X2=0 $Y2=0
cc_120 N_C_c_108_n N_VPWR_c_320_n 0.00858226f $X=1.2 $Y=1.765 $X2=0 $Y2=0
cc_121 N_C_c_109_n N_VPWR_c_320_n 0.00857848f $X=1.695 $Y=1.765 $X2=0 $Y2=0
cc_122 N_C_c_108_n N_Y_c_388_n 0.00257496f $X=1.2 $Y=1.765 $X2=0 $Y2=0
cc_123 N_C_c_109_n N_Y_c_388_n 4.27055e-19 $X=1.695 $Y=1.765 $X2=0 $Y2=0
cc_124 C N_Y_c_388_n 0.0272413f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_125 N_C_c_107_n N_Y_c_388_n 0.00171365f $X=1.615 $Y=1.515 $X2=0 $Y2=0
cc_126 N_C_c_108_n N_Y_c_383_n 0.0104597f $X=1.2 $Y=1.765 $X2=0 $Y2=0
cc_127 N_C_c_109_n N_Y_c_383_n 0.0102374f $X=1.695 $Y=1.765 $X2=0 $Y2=0
cc_128 N_C_c_109_n N_Y_c_394_n 0.01222f $X=1.695 $Y=1.765 $X2=0 $Y2=0
cc_129 C N_Y_c_394_n 0.0107028f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_130 N_C_c_104_n N_VGND_c_449_n 0.00556327f $X=0.955 $Y=1.185 $X2=0 $Y2=0
cc_131 N_C_c_104_n N_VGND_c_450_n 3.69172e-19 $X=0.955 $Y=1.185 $X2=0 $Y2=0
cc_132 N_C_c_105_n N_VGND_c_450_n 0.00769205f $X=1.385 $Y=1.185 $X2=0 $Y2=0
cc_133 N_C_c_104_n N_VGND_c_452_n 0.00433834f $X=0.955 $Y=1.185 $X2=0 $Y2=0
cc_134 N_C_c_105_n N_VGND_c_452_n 0.00281141f $X=1.385 $Y=1.185 $X2=0 $Y2=0
cc_135 N_C_c_104_n N_VGND_c_454_n 0.00825089f $X=0.955 $Y=1.185 $X2=0 $Y2=0
cc_136 N_C_c_105_n N_VGND_c_454_n 0.00365066f $X=1.385 $Y=1.185 $X2=0 $Y2=0
cc_137 N_C_c_104_n N_A_206_74#_c_498_n 0.00221999f $X=0.955 $Y=1.185 $X2=0 $Y2=0
cc_138 N_C_c_107_n N_A_206_74#_c_498_n 6.05124e-19 $X=1.615 $Y=1.515 $X2=0 $Y2=0
cc_139 N_C_c_104_n N_A_206_74#_c_495_n 0.00498672f $X=0.955 $Y=1.185 $X2=0 $Y2=0
cc_140 N_C_c_105_n N_A_206_74#_c_495_n 2.93125e-19 $X=1.385 $Y=1.185 $X2=0 $Y2=0
cc_141 N_C_c_105_n N_A_206_74#_c_496_n 0.0118272f $X=1.385 $Y=1.185 $X2=0 $Y2=0
cc_142 N_C_c_107_n N_A_206_74#_c_496_n 0.00167114f $X=1.615 $Y=1.515 $X2=0 $Y2=0
cc_143 N_C_c_105_n N_A_206_74#_c_497_n 0.00212344f $X=1.385 $Y=1.185 $X2=0 $Y2=0
cc_144 N_C_c_105_n N_A_403_54#_c_537_n 4.19228e-19 $X=1.385 $Y=1.185 $X2=0 $Y2=0
cc_145 N_A_27_94#_c_175_n N_B_c_281_n 0.0211788f $X=2.645 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_146 N_A_27_94#_M1005_g N_B_c_277_n 0.0272472f $X=2.85 $Y=0.87 $X2=0 $Y2=0
cc_147 N_A_27_94#_M1005_g B 0.00344966f $X=2.85 $Y=0.87 $X2=0 $Y2=0
cc_148 N_A_27_94#_c_173_n B 3.47983e-19 $X=2.645 $Y=1.557 $X2=0 $Y2=0
cc_149 N_A_27_94#_M1005_g N_B_c_280_n 0.0122044f $X=2.85 $Y=0.87 $X2=0 $Y2=0
cc_150 N_A_27_94#_c_173_n N_B_c_280_n 0.00166512f $X=2.645 $Y=1.557 $X2=0 $Y2=0
cc_151 N_A_27_94#_c_170_n N_VPWR_M1002_d 0.00142439f $X=0.805 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_152 N_A_27_94#_c_178_n N_VPWR_M1002_d 0.00276864f $X=0.805 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_153 N_A_27_94#_c_176_n N_VPWR_c_321_n 0.0471307f $X=0.47 $Y=2.815 $X2=0 $Y2=0
cc_154 N_A_27_94#_c_178_n N_VPWR_c_321_n 0.00476368f $X=0.805 $Y=2.035 $X2=0
+ $Y2=0
cc_155 N_A_27_94#_c_174_n N_VPWR_c_322_n 0.011285f $X=2.195 $Y=1.765 $X2=0 $Y2=0
cc_156 N_A_27_94#_c_175_n N_VPWR_c_322_n 5.55734e-19 $X=2.645 $Y=1.765 $X2=0
+ $Y2=0
cc_157 N_A_27_94#_c_175_n N_VPWR_c_323_n 0.00903992f $X=2.645 $Y=1.765 $X2=0
+ $Y2=0
cc_158 N_A_27_94#_c_176_n N_VPWR_c_326_n 0.0145938f $X=0.47 $Y=2.815 $X2=0 $Y2=0
cc_159 N_A_27_94#_c_174_n N_VPWR_c_330_n 0.00413917f $X=2.195 $Y=1.765 $X2=0
+ $Y2=0
cc_160 N_A_27_94#_c_175_n N_VPWR_c_330_n 0.00445602f $X=2.645 $Y=1.765 $X2=0
+ $Y2=0
cc_161 N_A_27_94#_c_174_n N_VPWR_c_320_n 0.00817726f $X=2.195 $Y=1.765 $X2=0
+ $Y2=0
cc_162 N_A_27_94#_c_175_n N_VPWR_c_320_n 0.00859358f $X=2.645 $Y=1.765 $X2=0
+ $Y2=0
cc_163 N_A_27_94#_c_176_n N_VPWR_c_320_n 0.0120466f $X=0.47 $Y=2.815 $X2=0 $Y2=0
cc_164 N_A_27_94#_c_178_n N_Y_c_388_n 0.00794558f $X=0.805 $Y=2.035 $X2=0 $Y2=0
cc_165 N_A_27_94#_c_174_n N_Y_c_383_n 7.87134e-19 $X=2.195 $Y=1.765 $X2=0 $Y2=0
cc_166 N_A_27_94#_c_176_n N_Y_c_383_n 0.00435639f $X=0.47 $Y=2.815 $X2=0 $Y2=0
cc_167 N_A_27_94#_c_174_n N_Y_c_394_n 0.0134681f $X=2.195 $Y=1.765 $X2=0 $Y2=0
cc_168 N_A_27_94#_c_172_n N_Y_c_394_n 0.0141818f $X=2.19 $Y=1.175 $X2=0 $Y2=0
cc_169 N_A_27_94#_c_173_n N_Y_c_394_n 7.25013e-19 $X=2.645 $Y=1.557 $X2=0 $Y2=0
cc_170 N_A_27_94#_c_174_n N_Y_c_384_n 0.00610043f $X=2.195 $Y=1.765 $X2=0 $Y2=0
cc_171 N_A_27_94#_c_175_n N_Y_c_384_n 0.0111767f $X=2.645 $Y=1.765 $X2=0 $Y2=0
cc_172 N_A_27_94#_c_173_n N_Y_c_404_n 0.00466734f $X=2.645 $Y=1.557 $X2=0 $Y2=0
cc_173 N_A_27_94#_c_175_n N_Y_c_405_n 0.0118676f $X=2.645 $Y=1.765 $X2=0 $Y2=0
cc_174 N_A_27_94#_c_173_n N_Y_c_405_n 0.00640314f $X=2.645 $Y=1.557 $X2=0 $Y2=0
cc_175 N_A_27_94#_c_175_n N_Y_c_385_n 8.78853e-19 $X=2.645 $Y=1.765 $X2=0 $Y2=0
cc_176 N_A_27_94#_c_165_n N_Y_c_408_n 0.00594556f $X=2.42 $Y=1.35 $X2=0 $Y2=0
cc_177 N_A_27_94#_M1005_g N_Y_c_408_n 0.00207245f $X=2.85 $Y=0.87 $X2=0 $Y2=0
cc_178 N_A_27_94#_c_172_n N_Y_c_408_n 0.0051356f $X=2.19 $Y=1.175 $X2=0 $Y2=0
cc_179 N_A_27_94#_c_174_n Y 0.00153193f $X=2.195 $Y=1.765 $X2=0 $Y2=0
cc_180 N_A_27_94#_c_165_n Y 0.00157436f $X=2.42 $Y=1.35 $X2=0 $Y2=0
cc_181 N_A_27_94#_c_175_n Y 0.00521289f $X=2.645 $Y=1.765 $X2=0 $Y2=0
cc_182 N_A_27_94#_M1005_g Y 0.00539959f $X=2.85 $Y=0.87 $X2=0 $Y2=0
cc_183 N_A_27_94#_c_172_n Y 0.0319153f $X=2.19 $Y=1.175 $X2=0 $Y2=0
cc_184 N_A_27_94#_c_173_n Y 0.0223711f $X=2.645 $Y=1.557 $X2=0 $Y2=0
cc_185 N_A_27_94#_c_168_n N_VGND_M1003_d 0.00116505f $X=0.72 $Y=1.175 $X2=-0.19
+ $Y2=-0.245
cc_186 N_A_27_94#_c_207_n N_VGND_M1003_d 0.00112241f $X=0.805 $Y=1.175 $X2=-0.19
+ $Y2=-0.245
cc_187 N_A_27_94#_c_171_n N_VGND_M1007_s 0.00205663f $X=2.025 $Y=1.175 $X2=0
+ $Y2=0
cc_188 N_A_27_94#_c_167_n N_VGND_c_449_n 0.0168919f $X=0.265 $Y=0.615 $X2=0
+ $Y2=0
cc_189 N_A_27_94#_c_168_n N_VGND_c_449_n 0.0100896f $X=0.72 $Y=1.175 $X2=0 $Y2=0
cc_190 N_A_27_94#_c_207_n N_VGND_c_449_n 0.00855018f $X=0.805 $Y=1.175 $X2=0
+ $Y2=0
cc_191 N_A_27_94#_c_165_n N_VGND_c_450_n 0.00241358f $X=2.42 $Y=1.35 $X2=0 $Y2=0
cc_192 N_A_27_94#_c_167_n N_VGND_c_451_n 0.00787252f $X=0.265 $Y=0.615 $X2=0
+ $Y2=0
cc_193 N_A_27_94#_c_165_n N_VGND_c_453_n 7.84925e-19 $X=2.42 $Y=1.35 $X2=0 $Y2=0
cc_194 N_A_27_94#_M1005_g N_VGND_c_453_n 7.84925e-19 $X=2.85 $Y=0.87 $X2=0 $Y2=0
cc_195 N_A_27_94#_c_167_n N_VGND_c_454_n 0.0085887f $X=0.265 $Y=0.615 $X2=0
+ $Y2=0
cc_196 N_A_27_94#_c_171_n N_A_206_74#_M1001_d 0.00176461f $X=2.025 $Y=1.175
+ $X2=-0.19 $Y2=-0.245
cc_197 N_A_27_94#_c_171_n N_A_206_74#_c_498_n 0.0151918f $X=2.025 $Y=1.175 $X2=0
+ $Y2=0
cc_198 N_A_27_94#_c_171_n N_A_206_74#_c_496_n 0.0479995f $X=2.025 $Y=1.175 $X2=0
+ $Y2=0
cc_199 N_A_27_94#_c_165_n N_A_206_74#_c_497_n 0.00301228f $X=2.42 $Y=1.35 $X2=0
+ $Y2=0
cc_200 N_A_27_94#_c_172_n N_A_206_74#_c_497_n 0.00682868f $X=2.19 $Y=1.175 $X2=0
+ $Y2=0
cc_201 N_A_27_94#_c_173_n N_A_206_74#_c_497_n 3.24197e-19 $X=2.645 $Y=1.557
+ $X2=0 $Y2=0
cc_202 N_A_27_94#_c_165_n N_A_206_74#_c_511_n 0.0159728f $X=2.42 $Y=1.35 $X2=0
+ $Y2=0
cc_203 N_A_27_94#_M1005_g N_A_206_74#_c_511_n 0.0149272f $X=2.85 $Y=0.87 $X2=0
+ $Y2=0
cc_204 N_A_27_94#_c_172_n N_A_206_74#_c_511_n 0.00950299f $X=2.19 $Y=1.175 $X2=0
+ $Y2=0
cc_205 N_A_27_94#_c_173_n N_A_206_74#_c_511_n 0.00128252f $X=2.645 $Y=1.557
+ $X2=0 $Y2=0
cc_206 N_A_27_94#_c_172_n N_A_403_54#_M1004_s 0.0033664f $X=2.19 $Y=1.175
+ $X2=-0.19 $Y2=-0.245
cc_207 N_A_27_94#_c_165_n N_A_403_54#_c_537_n 0.0103526f $X=2.42 $Y=1.35 $X2=0
+ $Y2=0
cc_208 N_A_27_94#_M1005_g N_A_403_54#_c_537_n 0.00963483f $X=2.85 $Y=0.87 $X2=0
+ $Y2=0
cc_209 N_B_c_281_n N_VPWR_c_323_n 0.0101198f $X=3.305 $Y=1.765 $X2=0 $Y2=0
cc_210 N_B_c_281_n N_VPWR_c_325_n 7.74286e-19 $X=3.305 $Y=1.765 $X2=0 $Y2=0
cc_211 N_B_c_282_n N_VPWR_c_325_n 0.0153451f $X=3.815 $Y=1.765 $X2=0 $Y2=0
cc_212 B N_VPWR_c_325_n 0.0255179f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_213 N_B_c_281_n N_VPWR_c_332_n 0.00445602f $X=3.305 $Y=1.765 $X2=0 $Y2=0
cc_214 N_B_c_282_n N_VPWR_c_332_n 0.00413917f $X=3.815 $Y=1.765 $X2=0 $Y2=0
cc_215 N_B_c_281_n N_VPWR_c_320_n 0.00860555f $X=3.305 $Y=1.765 $X2=0 $Y2=0
cc_216 N_B_c_282_n N_VPWR_c_320_n 0.00818274f $X=3.815 $Y=1.765 $X2=0 $Y2=0
cc_217 N_B_c_281_n N_Y_c_384_n 8.6014e-19 $X=3.305 $Y=1.765 $X2=0 $Y2=0
cc_218 N_B_c_281_n N_Y_c_404_n 0.0128654f $X=3.305 $Y=1.765 $X2=0 $Y2=0
cc_219 B N_Y_c_404_n 0.0256676f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_220 N_B_c_281_n N_Y_c_420_n 4.27055e-19 $X=3.305 $Y=1.765 $X2=0 $Y2=0
cc_221 B N_Y_c_420_n 0.0259268f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_222 N_B_c_280_n N_Y_c_420_n 0.00169967f $X=3.815 $Y=1.557 $X2=0 $Y2=0
cc_223 N_B_c_281_n N_Y_c_385_n 0.0119606f $X=3.305 $Y=1.765 $X2=0 $Y2=0
cc_224 N_B_c_282_n N_Y_c_385_n 0.00465795f $X=3.815 $Y=1.765 $X2=0 $Y2=0
cc_225 N_B_c_277_n N_Y_c_408_n 8.93946e-19 $X=3.41 $Y=1.35 $X2=0 $Y2=0
cc_226 N_B_c_281_n Y 0.00311836f $X=3.305 $Y=1.765 $X2=0 $Y2=0
cc_227 B Y 0.0313542f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_228 N_B_c_280_n Y 4.91491e-19 $X=3.815 $Y=1.557 $X2=0 $Y2=0
cc_229 N_B_c_277_n N_VGND_c_453_n 7.84925e-19 $X=3.41 $Y=1.35 $X2=0 $Y2=0
cc_230 N_B_c_278_n N_VGND_c_453_n 7.84925e-19 $X=3.84 $Y=1.35 $X2=0 $Y2=0
cc_231 N_B_c_277_n N_A_206_74#_c_515_n 0.0187719f $X=3.41 $Y=1.35 $X2=0 $Y2=0
cc_232 N_B_c_278_n N_A_206_74#_c_515_n 0.00611925f $X=3.84 $Y=1.35 $X2=0 $Y2=0
cc_233 B N_A_206_74#_c_515_n 0.0574195f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_234 N_B_c_280_n N_A_206_74#_c_515_n 0.00462978f $X=3.815 $Y=1.557 $X2=0 $Y2=0
cc_235 N_B_c_277_n N_A_403_54#_c_537_n 0.00963483f $X=3.41 $Y=1.35 $X2=0 $Y2=0
cc_236 N_B_c_278_n N_A_403_54#_c_537_n 0.0140521f $X=3.84 $Y=1.35 $X2=0 $Y2=0
cc_237 B N_A_403_54#_c_538_n 0.020209f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_238 N_VPWR_c_321_n N_Y_c_383_n 0.0253838f $X=0.95 $Y=2.455 $X2=0 $Y2=0
cc_239 N_VPWR_c_322_n N_Y_c_383_n 0.0271924f $X=1.97 $Y=2.41 $X2=0 $Y2=0
cc_240 N_VPWR_c_328_n N_Y_c_383_n 0.0165599f $X=1.805 $Y=3.33 $X2=0 $Y2=0
cc_241 N_VPWR_c_320_n N_Y_c_383_n 0.0136411f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_242 N_VPWR_M1006_s N_Y_c_394_n 0.0104614f $X=1.77 $Y=1.84 $X2=0 $Y2=0
cc_243 N_VPWR_c_322_n N_Y_c_394_n 0.0202249f $X=1.97 $Y=2.41 $X2=0 $Y2=0
cc_244 N_VPWR_c_322_n N_Y_c_384_n 0.0462948f $X=1.97 $Y=2.41 $X2=0 $Y2=0
cc_245 N_VPWR_c_323_n N_Y_c_384_n 0.0454782f $X=2.955 $Y=2.41 $X2=0 $Y2=0
cc_246 N_VPWR_c_330_n N_Y_c_384_n 0.0110241f $X=2.79 $Y=3.33 $X2=0 $Y2=0
cc_247 N_VPWR_c_320_n N_Y_c_384_n 0.00909194f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_248 N_VPWR_M1012_s N_Y_c_404_n 0.0132318f $X=2.72 $Y=1.84 $X2=0 $Y2=0
cc_249 N_VPWR_M1012_s N_Y_c_405_n 6.74228e-19 $X=2.72 $Y=1.84 $X2=0 $Y2=0
cc_250 N_VPWR_c_323_n N_Y_c_405_n 0.0266127f $X=2.955 $Y=2.41 $X2=0 $Y2=0
cc_251 N_VPWR_c_323_n N_Y_c_385_n 0.0404971f $X=2.955 $Y=2.41 $X2=0 $Y2=0
cc_252 N_VPWR_c_325_n N_Y_c_385_n 0.0315827f $X=4.04 $Y=2.035 $X2=0 $Y2=0
cc_253 N_VPWR_c_332_n N_Y_c_385_n 0.0145938f $X=3.875 $Y=3.33 $X2=0 $Y2=0
cc_254 N_VPWR_c_320_n N_Y_c_385_n 0.0120466f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_255 N_VPWR_M1012_s Y 0.001752f $X=2.72 $Y=1.84 $X2=0 $Y2=0
cc_256 N_Y_M1004_d N_A_206_74#_c_511_n 0.00337414f $X=2.495 $Y=0.5 $X2=0 $Y2=0
cc_257 N_Y_c_408_n N_A_206_74#_c_511_n 0.0168934f $X=2.635 $Y=1.095 $X2=0 $Y2=0
cc_258 N_VGND_c_449_n N_A_206_74#_c_498_n 0.01223f $X=0.695 $Y=0.725 $X2=0 $Y2=0
cc_259 N_VGND_c_449_n N_A_206_74#_c_495_n 0.0296545f $X=0.695 $Y=0.725 $X2=0
+ $Y2=0
cc_260 N_VGND_c_450_n N_A_206_74#_c_495_n 0.0104546f $X=1.6 $Y=0.495 $X2=0 $Y2=0
cc_261 N_VGND_c_452_n N_A_206_74#_c_495_n 0.0118323f $X=1.435 $Y=0 $X2=0 $Y2=0
cc_262 N_VGND_c_454_n N_A_206_74#_c_495_n 0.00911095f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_263 N_VGND_M1007_s N_A_206_74#_c_496_n 0.00433153f $X=1.46 $Y=0.37 $X2=0
+ $Y2=0
cc_264 N_VGND_c_450_n N_A_206_74#_c_496_n 0.0212697f $X=1.6 $Y=0.495 $X2=0 $Y2=0
cc_265 N_VGND_c_452_n N_A_206_74#_c_496_n 0.00197156f $X=1.435 $Y=0 $X2=0 $Y2=0
cc_266 N_VGND_c_453_n N_A_206_74#_c_496_n 0.0024506f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_267 N_VGND_c_454_n N_A_206_74#_c_496_n 0.00976958f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_268 N_VGND_c_453_n N_A_206_74#_c_497_n 6.97459e-19 $X=4.08 $Y=0 $X2=0 $Y2=0
cc_269 N_VGND_c_454_n N_A_206_74#_c_497_n 0.00468475f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_270 N_VGND_c_450_n N_A_403_54#_c_537_n 0.0128051f $X=1.6 $Y=0.495 $X2=0 $Y2=0
cc_271 N_VGND_c_453_n N_A_403_54#_c_537_n 0.0990761f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_272 N_VGND_c_454_n N_A_403_54#_c_537_n 0.0808667f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_273 N_A_206_74#_c_497_n N_A_403_54#_M1004_s 0.00147525f $X=2.105 $Y=0.795
+ $X2=-0.19 $Y2=-0.245
cc_274 N_A_206_74#_c_511_n N_A_403_54#_M1004_s 0.00484861f $X=2.97 $Y=0.925
+ $X2=-0.19 $Y2=-0.245
cc_275 N_A_206_74#_c_515_n N_A_403_54#_M1005_s 0.00952501f $X=3.625 $Y=0.755
+ $X2=0 $Y2=0
cc_276 N_A_206_74#_c_497_n N_A_403_54#_c_537_n 0.11551f $X=2.105 $Y=0.795 $X2=0
+ $Y2=0
