* File: sky130_fd_sc_ls__nand3b_2.spice
* Created: Fri Aug 28 13:34:15 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__nand3b_2.pex.spice"
.subckt sky130_fd_sc_ls__nand3b_2  VNB VPB A_N C B VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B	B
* C	C
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_A_N_M1003_g N_A_27_94#_M1003_s VNB NSHORT L=0.15 W=0.64
+ AD=0.108058 AS=0.1728 PD=0.987826 PS=1.82 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75001.1 A=0.096 P=1.58 MULT=1
MM1001 N_A_206_74#_M1001_d N_C_M1001_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.124942 PD=1.02 PS=1.14217 NRD=0 NRS=7.296 M=1 R=4.93333
+ SA=75000.6 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1007 N_A_206_74#_M1001_d N_C_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.19445 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75001
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1004 N_Y_M1004_d N_A_27_94#_M1004_g N_A_403_54#_M1004_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.24845 PD=1.02 PS=2.6 NRD=0 NRS=45.516 M=1 R=4.93333
+ SA=75000.2 SB=75001.6 A=0.111 P=1.78 MULT=1
MM1005 N_Y_M1004_d N_A_27_94#_M1005_g N_A_403_54#_M1005_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1816 PD=1.02 PS=1.38 NRD=0 NRS=30.876 M=1 R=4.93333
+ SA=75000.6 SB=75001.2 A=0.111 P=1.78 MULT=1
MM1009 N_A_206_74#_M1009_d N_B_M1009_g N_A_403_54#_M1005_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1816 PD=1.02 PS=1.38 NRD=0 NRS=30.876 M=1 R=4.93333
+ SA=75001.2 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1011 N_A_206_74#_M1009_d N_B_M1011_g N_A_403_54#_M1011_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1998 PD=1.02 PS=2.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1002 N_VPWR_M1002_d N_A_N_M1002_g N_A_27_94#_M1002_s VPB PHIGHVT L=0.15 W=1
+ AD=0.182453 AS=0.295 PD=1.39151 PS=2.59 NRD=7.8603 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75003.3 A=0.15 P=2.3 MULT=1
MM1000 N_Y_M1000_d N_C_M1000_g N_VPWR_M1002_d VPB PHIGHVT L=0.15 W=1.12
+ AD=0.1932 AS=0.204347 PD=1.465 PS=1.55849 NRD=5.2599 NRS=6.1464 M=1 R=7.46667
+ SA=75000.7 SB=75002.8 A=0.168 P=2.54 MULT=1
MM1006 N_Y_M1000_d N_C_M1006_g N_VPWR_M1006_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.1932 AS=0.196 PD=1.465 PS=1.47 NRD=6.1464 NRS=10.5395 M=1 R=7.46667
+ SA=75001.2 SB=75002.3 A=0.168 P=2.54 MULT=1
MM1008 N_Y_M1008_d N_A_27_94#_M1008_g N_VPWR_M1006_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.7 SB=75001.8 A=0.168 P=2.54 MULT=1
MM1012 N_Y_M1008_d N_A_27_94#_M1012_g N_VPWR_M1012_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.2856 PD=1.42 PS=1.63 NRD=1.7533 NRS=16.7056 M=1 R=7.46667
+ SA=75002.1 SB=75001.4 A=0.168 P=2.54 MULT=1
MM1010 N_Y_M1010_d N_B_M1010_g N_VPWR_M1012_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.2016 AS=0.2856 PD=1.48 PS=1.63 NRD=1.7533 NRS=23.7385 M=1 R=7.46667
+ SA=75002.8 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1013 N_Y_M1010_d N_B_M1013_g N_VPWR_M1013_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.2016 AS=0.3304 PD=1.48 PS=2.83 NRD=12.2928 NRS=1.7533 M=1 R=7.46667
+ SA=75003.3 SB=75000.2 A=0.168 P=2.54 MULT=1
DX14_noxref VNB VPB NWDIODE A=8.742 P=13.12
*
.include "sky130_fd_sc_ls__nand3b_2.pxi.spice"
*
.ends
*
*
