* NGSPICE file created from sky130_fd_sc_ls__dlxbn_2.ext - technology: sky130A

.subckt sky130_fd_sc_ls__dlxbn_2 D GATE_N VGND VNB VPB VPWR Q Q_N
M1000 VPWR D a_27_136# VPB phighvt w=840000u l=150000u
+  ad=2.5372e+12p pd=1.986e+07u as=3.192e+11p ps=2.44e+06u
M1001 a_232_98# GATE_N VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=2.0325e+12p ps=1.669e+07u
M1002 Q a_887_270# VGND VNB nshort w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1003 VPWR a_887_270# Q VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.36e+11p ps=2.84e+06u
M1004 a_814_392# a_232_98# a_647_79# VPB phighvt w=420000u l=150000u
+  ad=1.596e+11p pd=1.6e+06u as=4.372e+11p ps=3.35e+06u
M1005 VGND a_232_98# a_343_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.817e+11p ps=2.29e+06u
M1006 a_232_98# GATE_N VPWR VPB phighvt w=840000u l=150000u
+  ad=2.478e+11p pd=2.27e+06u as=0p ps=0u
M1007 Q_N a_1442_94# VGND VNB nshort w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1008 VPWR a_232_98# a_343_74# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=2.478e+11p ps=2.27e+06u
M1009 VGND a_887_270# Q VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_1442_94# a_887_270# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.95e+11p pd=2.59e+06u as=0p ps=0u
M1011 Q_N a_1442_94# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=0p ps=0u
M1012 a_569_79# a_27_136# VGND VNB nshort w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1013 a_647_79# a_232_98# a_569_79# VNB nshort w=640000u l=150000u
+  ad=3.952e+11p pd=2.9e+06u as=0p ps=0u
M1014 a_647_79# a_343_74# a_565_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1015 VGND a_1442_94# Q_N VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_887_270# a_647_79# VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1017 a_1442_94# a_887_270# VGND VNB nshort w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=0p ps=0u
M1018 VPWR a_887_270# a_814_392# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_887_270# a_647_79# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=0p ps=0u
M1020 VPWR a_1442_94# Q_N VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND D a_27_136# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1022 a_565_392# a_27_136# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VGND a_887_270# a_839_123# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1024 Q a_887_270# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_839_123# a_343_74# a_647_79# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

