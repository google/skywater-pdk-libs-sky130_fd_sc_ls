* File: sky130_fd_sc_ls__dfbbp_1.spice
* Created: Wed Sep  2 11:00:37 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__dfbbp_1.pex.spice"
.subckt sky130_fd_sc_ls__dfbbp_1  VNB VPB CLK D SET_B RESET_B VPWR Q_N Q VGND
* 
* VGND	VGND
* Q	Q
* Q_N	Q_N
* VPWR	VPWR
* RESET_B	RESET_B
* SET_B	SET_B
* D	D
* CLK	CLK
* VPB	VPB
* VNB	VNB
MM1029 N_VGND_M1029_d N_CLK_M1029_g N_A_27_74#_M1029_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1295 AS=0.2109 PD=1.09 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1013 N_A_214_74#_M1013_d N_A_27_74#_M1013_g N_VGND_M1029_d VNB NSHORT L=0.15
+ W=0.74 AD=0.2109 AS=0.1295 PD=2.05 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.7 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1031 N_A_422_125#_M1031_d N_D_M1031_g N_VGND_M1031_s VNB NSHORT L=0.15 W=0.42
+ AD=0.088025 AS=0.1197 PD=0.95 PS=1.41 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.1 A=0.063 P=1.14 MULT=1
MM1006 N_A_520_87#_M1006_d N_A_27_74#_M1006_g N_A_422_125#_M1031_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.0588 AS=0.088025 PD=0.7 PS=0.95 NRD=0 NRS=18.564 M=1 R=2.8
+ SA=75000.5 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1025 A_606_87# N_A_214_74#_M1025_g N_A_520_87#_M1006_d VNB NSHORT L=0.15
+ W=0.42 AD=0.08225 AS=0.0588 PD=0.905 PS=0.7 NRD=40.236 NRS=0 M=1 R=2.8
+ SA=75000.9 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1034 N_VGND_M1034_d N_A_671_93#_M1034_g A_606_87# VNB NSHORT L=0.15 W=0.42
+ AD=0.205962 AS=0.08225 PD=1.31629 PS=0.905 NRD=124.392 NRS=40.236 M=1 R=2.8
+ SA=75001 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1035 N_A_872_119#_M1035_d N_SET_B_M1035_g N_VGND_M1034_d VNB NSHORT L=0.15
+ W=0.55 AD=0.192025 AS=0.269713 PD=1.335 PS=1.72371 NRD=64.164 NRS=94.992 M=1
+ R=3.66667 SA=75001.5 SB=75001.4 A=0.0825 P=1.4 MULT=1
MM1019 N_A_671_93#_M1019_d N_A_520_87#_M1019_g N_A_872_119#_M1035_d VNB NSHORT
+ L=0.15 W=0.55 AD=0.077 AS=0.192025 PD=0.83 PS=1.335 NRD=0 NRS=64.164 M=1
+ R=3.66667 SA=75002.1 SB=75000.7 A=0.0825 P=1.4 MULT=1
MM1032 N_A_872_119#_M1032_d N_A_1062_93#_M1032_g N_A_671_93#_M1019_d VNB NSHORT
+ L=0.15 W=0.55 AD=0.26245 AS=0.077 PD=2.29 PS=0.83 NRD=92.112 NRS=0 M=1
+ R=3.66667 SA=75002.6 SB=75000.3 A=0.0825 P=1.4 MULT=1
MM1007 A_1318_119# N_A_671_93#_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.55
+ AD=0.05775 AS=0.26105 PD=0.76 PS=2.28 NRD=10.908 NRS=0 M=1 R=3.66667
+ SA=75000.3 SB=75001.5 A=0.0825 P=1.4 MULT=1
MM1011 N_A_1311_424#_M1011_d N_A_214_74#_M1011_g A_1318_119# VNB NSHORT L=0.15
+ W=0.55 AD=0.131376 AS=0.05775 PD=1.32113 PS=0.76 NRD=0 NRS=10.908 M=1
+ R=3.66667 SA=75000.6 SB=75001.1 A=0.0825 P=1.4 MULT=1
MM1012 A_1498_74# N_A_27_74#_M1012_g N_A_1311_424#_M1011_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0819 AS=0.100324 PD=0.81 PS=1.00887 NRD=39.996 NRS=32.856 M=1
+ R=2.8 SA=75000.6 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1016 N_VGND_M1016_d N_A_1474_446#_M1016_g A_1498_74# VNB NSHORT L=0.15 W=0.42
+ AD=0.0877655 AS=0.0819 PD=0.796552 PS=0.81 NRD=22.848 NRS=39.996 M=1 R=2.8
+ SA=75001.2 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1033 N_A_1708_74#_M1033_d N_SET_B_M1033_g N_VGND_M1016_d VNB NSHORT L=0.15
+ W=0.74 AD=0.1295 AS=0.154634 PD=1.09 PS=1.40345 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75001.1 SB=75001.2 A=0.111 P=1.78 MULT=1
MM1027 N_A_1474_446#_M1027_d N_A_1311_424#_M1027_g N_A_1708_74#_M1033_d VNB
+ NSHORT L=0.15 W=0.74 AD=0.10545 AS=0.1295 PD=1.025 PS=1.09 NRD=0.804 NRS=0 M=1
+ R=4.93333 SA=75001.6 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1030 N_A_1708_74#_M1030_d N_A_1062_93#_M1030_g N_A_1474_446#_M1027_d VNB
+ NSHORT L=0.15 W=0.74 AD=0.2294 AS=0.10545 PD=2.1 PS=1.025 NRD=4.044 NRS=0 M=1
+ R=4.93333 SA=75002 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1008 N_VGND_M1008_d N_RESET_B_M1008_g N_A_1062_93#_M1008_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0943552 AS=0.1197 PD=0.847241 PS=1.41 NRD=22.848 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1003 N_Q_N_M1003_d N_A_1474_446#_M1003_g N_VGND_M1008_d VNB NSHORT L=0.15
+ W=0.74 AD=0.2109 AS=0.166245 PD=2.05 PS=1.49276 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75000.5 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1015 N_VGND_M1015_d N_A_1474_446#_M1015_g N_A_2320_410#_M1015_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0783879 AS=0.1197 PD=0.771207 PS=1.41 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1036 N_Q_M1036_d N_A_2320_410#_M1036_g N_VGND_M1015_d VNB NSHORT L=0.15 W=0.74
+ AD=0.1998 AS=0.138112 PD=2.02 PS=1.35879 NRD=0 NRS=7.296 M=1 R=4.93333
+ SA=75000.5 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1037 N_VPWR_M1037_d N_CLK_M1037_g N_A_27_74#_M1037_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.2408 AS=0.3304 PD=1.55 PS=2.83 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.8 A=0.168 P=2.54 MULT=1
MM1014 N_A_214_74#_M1014_d N_A_27_74#_M1014_g N_VPWR_M1037_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.308 AS=0.2408 PD=2.79 PS=1.55 NRD=1.7533 NRS=15.8191 M=1 R=7.46667
+ SA=75000.8 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1024 N_A_422_125#_M1024_d N_D_M1024_g N_VPWR_M1024_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.063 AS=0.2604 PD=0.72 PS=2.08 NRD=4.6886 NRS=7.0329 M=1 R=2.8 SA=75000.5
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1038 N_A_520_87#_M1038_d N_A_214_74#_M1038_g N_A_422_125#_M1024_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.11445 AS=0.063 PD=1.21 PS=0.72 NRD=102.007 NRS=4.6886 M=1
+ R=2.8 SA=75001 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1028 A_713_379# N_A_27_74#_M1028_g N_A_520_87#_M1038_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0504 AS=0.11445 PD=0.66 PS=1.21 NRD=30.4759 NRS=4.6886 M=1 R=2.8
+ SA=75000.2 SB=75002.9 A=0.063 P=1.14 MULT=1
MM1010 N_VPWR_M1010_d N_A_671_93#_M1010_g A_713_379# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0987 AS=0.0504 PD=0.853333 PS=0.66 NRD=4.6886 NRS=30.4759 M=1 R=2.8
+ SA=75000.6 SB=75002.5 A=0.063 P=1.14 MULT=1
MM1022 N_A_671_93#_M1022_d N_SET_B_M1022_g N_VPWR_M1010_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.1638 AS=0.1974 PD=1.23 PS=1.70667 NRD=23.443 NRS=35.1645 M=1 R=5.6
+ SA=75000.7 SB=75002.8 A=0.126 P=1.98 MULT=1
MM1001 A_1017_379# N_A_520_87#_M1001_g N_A_671_93#_M1022_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.1134 AS=0.1638 PD=1.11 PS=1.23 NRD=18.7544 NRS=2.3443 M=1 R=5.6
+ SA=75001.2 SB=75002.2 A=0.126 P=1.98 MULT=1
MM1021 N_VPWR_M1021_d N_A_1062_93#_M1021_g A_1017_379# VPB PHIGHVT L=0.15 W=0.84
+ AD=0.1512 AS=0.1134 PD=1.2 PS=1.11 NRD=9.3772 NRS=18.7544 M=1 R=5.6 SA=75001.6
+ SB=75001.8 A=0.126 P=1.98 MULT=1
MM1023 A_1203_379# N_A_671_93#_M1023_g N_VPWR_M1021_d VPB PHIGHVT L=0.15 W=0.84
+ AD=0.17955 AS=0.1512 PD=1.455 PS=1.2 NRD=37.2133 NRS=9.3772 M=1 R=5.6
+ SA=75002.2 SB=75001.3 A=0.126 P=1.98 MULT=1
MM1005 N_A_1311_424#_M1005_d N_A_27_74#_M1005_g A_1203_379# VPB PHIGHVT L=0.15
+ W=0.84 AD=0.1904 AS=0.17955 PD=1.63333 PS=1.455 NRD=2.3443 NRS=37.2133 M=1
+ R=5.6 SA=75001.9 SB=75001.7 A=0.126 P=1.98 MULT=1
MM1020 A_1418_508# N_A_214_74#_M1020_g N_A_1311_424#_M1005_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.06195 AS=0.0952 PD=0.715 PS=0.816667 NRD=43.3794 NRS=44.5417 M=1
+ R=2.8 SA=75001.7 SB=75002.6 A=0.063 P=1.14 MULT=1
MM1039 N_VPWR_M1039_d N_A_1474_446#_M1039_g A_1418_508# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.153537 AS=0.06195 PD=1.1062 PS=0.715 NRD=23.443 NRS=43.3794 M=1
+ R=2.8 SA=75002.1 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1004 N_A_1474_446#_M1004_d N_SET_B_M1004_g N_VPWR_M1039_d VPB PHIGHVT L=0.15
+ W=1 AD=0.1825 AS=0.365563 PD=1.365 PS=2.6338 NRD=14.775 NRS=1.9503 M=1
+ R=6.66667 SA=75001.4 SB=75001.1 A=0.15 P=2.3 MULT=1
MM1002 A_1814_392# N_A_1311_424#_M1002_g N_A_1474_446#_M1004_d VPB PHIGHVT
+ L=0.15 W=1 AD=0.1325 AS=0.1825 PD=1.265 PS=1.365 NRD=15.2478 NRS=1.9503 M=1
+ R=6.66667 SA=75001.9 SB=75000.6 A=0.15 P=2.3 MULT=1
MM1000 N_VPWR_M1000_d N_A_1062_93#_M1000_g A_1814_392# VPB PHIGHVT L=0.15 W=1
+ AD=0.295 AS=0.1325 PD=2.59 PS=1.265 NRD=1.9503 NRS=15.2478 M=1 R=6.66667
+ SA=75002.4 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1026 N_VPWR_M1026_d N_RESET_B_M1026_g N_A_1062_93#_M1026_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.132945 AS=0.176 PD=1.08 PS=1.83 NRD=47.0042 NRS=3.0732 M=1
+ R=4.26667 SA=75000.2 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1017 N_Q_N_M1017_d N_A_1474_446#_M1017_g N_VPWR_M1026_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.308 AS=0.232655 PD=2.79 PS=1.89 NRD=1.7533 NRS=1.7533 M=1
+ R=7.46667 SA=75000.5 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1009 N_VPWR_M1009_d N_A_1474_446#_M1009_g N_A_2320_410#_M1009_s VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.1644 AS=0.231 PD=1.27286 PS=2.23 NRD=34.0022 NRS=0 M=1
+ R=5.6 SA=75000.2 SB=75000.7 A=0.126 P=1.98 MULT=1
MM1018 N_Q_M1018_d N_A_2320_410#_M1018_g N_VPWR_M1009_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.3192 AS=0.2192 PD=2.81 PS=1.69714 NRD=1.7533 NRS=1.7533 M=1
+ R=7.46667 SA=75000.6 SB=75000.2 A=0.168 P=2.54 MULT=1
DX40_noxref VNB VPB NWDIODE A=24.8124 P=30.4
c_150 VNB 0 1.25678e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_ls__dfbbp_1.pxi.spice"
*
.ends
*
*
