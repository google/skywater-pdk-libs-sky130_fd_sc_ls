* File: sky130_fd_sc_ls__sdfsbp_1.spice
* Created: Fri Aug 28 14:03:53 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__sdfsbp_1.pex.spice"
.subckt sky130_fd_sc_ls__sdfsbp_1  VNB VPB SCE D SCD CLK SET_B VPWR Q_N Q VGND
* 
* VGND	VGND
* Q	Q
* Q_N	Q_N
* VPWR	VPWR
* SET_B	SET_B
* CLK	CLK
* SCD	SCD
* D	D
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1033 N_VGND_M1033_d N_SCE_M1033_g N_A_27_74#_M1033_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0882 AS=0.1197 PD=0.84 PS=1.41 NRD=19.992 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1036 A_228_74# N_A_27_74#_M1036_g N_VGND_M1033_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0882 PD=0.66 PS=0.84 NRD=18.564 NRS=19.992 M=1 R=2.8 SA=75000.8
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1037 N_A_290_464#_M1037_d N_D_M1037_g A_228_74# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0504 PD=0.7 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.2
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1011 A_392_74# N_SCE_M1011_g N_A_290_464#_M1037_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0588 PD=0.66 PS=0.7 NRD=18.564 NRS=0 M=1 R=2.8 SA=75001.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1012 N_VGND_M1012_d N_SCD_M1012_g A_392_74# VNB NSHORT L=0.15 W=0.42 AD=0.1197
+ AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75002 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1022 N_VGND_M1022_d N_CLK_M1022_g N_A_594_74#_M1022_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1295 AS=0.2109 PD=1.09 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1020 N_A_781_74#_M1020_d N_A_594_74#_M1020_g N_VGND_M1022_d VNB NSHORT L=0.15
+ W=0.74 AD=0.2109 AS=0.1295 PD=2.05 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75000.7 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1034 N_A_995_74#_M1034_d N_A_594_74#_M1034_g N_A_290_464#_M1034_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0945 AS=0.18665 PD=0.87 PS=1.8 NRD=48.564 NRS=24.276 M=1
+ R=2.8 SA=75000.3 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1004 A_1115_74# N_A_781_74#_M1004_g N_A_995_74#_M1034_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.0945 PD=0.66 PS=0.87 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75000.9 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_A_1163_48#_M1002_g A_1115_74# VNB NSHORT L=0.15 W=0.42
+ AD=0.17255 AS=0.0504 PD=1.68 PS=0.66 NRD=25.704 NRS=18.564 M=1 R=2.8
+ SA=75001.3 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1041 A_1411_74# N_A_995_74#_M1041_g N_A_1163_48#_M1041_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75004.2 A=0.063 P=1.14 MULT=1
MM1010 N_VGND_M1010_d N_SET_B_M1010_g A_1411_74# VNB NSHORT L=0.15 W=0.42
+ AD=0.20267 AS=0.0504 PD=1.16094 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.6
+ SB=75003.9 A=0.063 P=1.14 MULT=1
MM1023 A_1684_74# N_A_995_74#_M1023_g N_VGND_M1010_d VNB NSHORT L=0.15 W=0.64
+ AD=0.0768 AS=0.30883 PD=0.88 PS=1.76906 NRD=12.18 NRS=0 M=1 R=4.26667
+ SA=75001.3 SB=75002.1 A=0.096 P=1.58 MULT=1
MM1024 N_A_1762_74#_M1024_d N_A_781_74#_M1024_g A_1684_74# VNB NSHORT L=0.15
+ W=0.64 AD=0.144362 AS=0.0768 PD=1.28 PS=0.88 NRD=13.116 NRS=12.18 M=1
+ R=4.26667 SA=75001.7 SB=75001.7 A=0.096 P=1.58 MULT=1
MM1000 A_1876_74# N_A_594_74#_M1000_g N_A_1762_74#_M1024_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.0947377 PD=0.66 PS=0.84 NRD=18.564 NRS=20.712 M=1 R=2.8
+ SA=75002.5 SB=75001.9 A=0.063 P=1.14 MULT=1
MM1001 A_1954_74# N_A_1924_48#_M1001_g A_1876_74# VNB NSHORT L=0.15 W=0.42
+ AD=0.0819 AS=0.0504 PD=0.81 PS=0.66 NRD=39.996 NRS=18.564 M=1 R=2.8 SA=75002.9
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1007 N_VGND_M1007_d N_SET_B_M1007_g A_1954_74# VNB NSHORT L=0.15 W=0.42
+ AD=0.1323 AS=0.0819 PD=1.05 PS=0.81 NRD=0 NRS=39.996 M=1 R=2.8 SA=75003.5
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1003 N_A_1924_48#_M1003_d N_A_1762_74#_M1003_g N_VGND_M1007_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.1197 AS=0.1323 PD=1.41 PS=1.05 NRD=0 NRS=0 M=1 R=2.8
+ SA=75004.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1005 N_Q_N_M1005_d N_A_1762_74#_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15
+ W=0.74 AD=0.2109 AS=0.2627 PD=2.05 PS=2.19 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75000.3 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1016 N_VGND_M1016_d N_A_1762_74#_M1016_g N_A_2556_112#_M1016_s VNB NSHORT
+ L=0.15 W=0.55 AD=0.172973 AS=0.15675 PD=1.15543 PS=1.67 NRD=58.356 NRS=0 M=1
+ R=3.66667 SA=75000.2 SB=75001 A=0.0825 P=1.4 MULT=1
MM1028 N_Q_M1028_d N_A_2556_112#_M1028_g N_VGND_M1016_d VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.232727 PD=2.05 PS=1.55457 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75000.8 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1026 N_VPWR_M1026_d N_SCE_M1026_g N_A_27_74#_M1026_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.096 AS=0.1888 PD=0.94 PS=1.87 NRD=3.0732 NRS=3.0732 M=1 R=4.26667
+ SA=75000.2 SB=75002.2 A=0.096 P=1.58 MULT=1
MM1027 A_206_464# N_SCE_M1027_g N_VPWR_M1026_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0864 AS=0.096 PD=0.91 PS=0.94 NRD=24.625 NRS=3.0732 M=1 R=4.26667
+ SA=75000.7 SB=75001.7 A=0.096 P=1.58 MULT=1
MM1014 N_A_290_464#_M1014_d N_D_M1014_g A_206_464# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1536 AS=0.0864 PD=1.12 PS=0.91 NRD=30.7714 NRS=24.625 M=1 R=4.26667
+ SA=75001.1 SB=75001.3 A=0.096 P=1.58 MULT=1
MM1039 A_416_464# N_A_27_74#_M1039_g N_A_290_464#_M1014_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0864 AS=0.1536 PD=0.91 PS=1.12 NRD=24.625 NRS=30.7714 M=1
+ R=4.26667 SA=75001.7 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1031 N_VPWR_M1031_d N_SCD_M1031_g A_416_464# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.208 AS=0.0864 PD=1.93 PS=0.91 NRD=4.6098 NRS=24.625 M=1 R=4.26667
+ SA=75002.1 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1019 N_VPWR_M1019_d N_CLK_M1019_g N_A_594_74#_M1019_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.3248 PD=1.42 PS=2.82 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1029 N_A_781_74#_M1029_d N_A_594_74#_M1029_g N_VPWR_M1019_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.3192 AS=0.168 PD=2.81 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1017 N_A_995_74#_M1017_d N_A_781_74#_M1017_g N_A_290_464#_M1017_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.105862 AS=0.1197 PD=0.95 PS=1.41 NRD=39.8531 NRS=4.6886 M=1
+ R=2.8 SA=75000.2 SB=75002.6 A=0.063 P=1.14 MULT=1
MM1018 A_1133_478# N_A_594_74#_M1018_g N_A_995_74#_M1017_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0837 AS=0.105862 PD=0.865 PS=0.95 NRD=67.6695 NRS=42.1974 M=1
+ R=2.8 SA=75000.7 SB=75002.1 A=0.063 P=1.14 MULT=1
MM1025 N_VPWR_M1025_d N_A_1163_48#_M1025_g A_1133_478# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.11235 AS=0.0837 PD=0.955 PS=0.865 NRD=7.0329 NRS=67.6695 M=1 R=2.8
+ SA=75001.1 SB=75002 A=0.063 P=1.14 MULT=1
MM1040 N_A_1163_48#_M1040_d N_A_995_74#_M1040_g N_VPWR_M1025_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0924 AS=0.11235 PD=0.86 PS=0.955 NRD=4.6886 NRS=112.566 M=1
+ R=2.8 SA=75001.8 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1013 N_VPWR_M1013_d N_SET_B_M1013_g N_A_1163_48#_M1040_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0939085 AS=0.0924 PD=0.822254 PS=0.86 NRD=46.886 NRS=70.3487 M=1
+ R=2.8 SA=75002.4 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1008 N_A_1600_347#_M1008_d N_A_995_74#_M1008_g N_VPWR_M1013_d VPB PHIGHVT
+ L=0.15 W=1 AD=0.29 AS=0.223592 PD=2.58 PS=1.95775 NRD=1.9503 NRS=1.9503 M=1
+ R=6.66667 SA=75001.3 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1035 N_A_1762_74#_M1035_d N_A_781_74#_M1035_g N_A_1712_374#_M1035_s VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.0939085 AS=0.2526 PD=0.822254 PS=3.03 NRD=44.5417
+ NRS=256.297 M=1 R=2.8 SA=75000.2 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1009 N_A_1600_347#_M1009_d N_A_594_74#_M1009_g N_A_1762_74#_M1035_d VPB
+ PHIGHVT L=0.15 W=1 AD=0.29 AS=0.223592 PD=2.58 PS=1.95775 NRD=1.9503
+ NRS=2.9353 M=1 R=6.66667 SA=75000.4 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1006 N_VPWR_M1006_d N_A_1924_48#_M1006_g N_A_1712_374#_M1006_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.063 AS=0.1218 PD=0.72 PS=1.42 NRD=4.6886 NRS=4.6886 M=1
+ R=2.8 SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1015 N_A_1762_74#_M1015_d N_SET_B_M1015_g N_VPWR_M1006_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1218 AS=0.063 PD=1.42 PS=0.72 NRD=4.6886 NRS=4.6886 M=1 R=2.8
+ SA=75000.7 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1032 N_VPWR_M1032_d N_A_1762_74#_M1032_g N_A_1924_48#_M1032_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0912545 AS=0.1218 PD=0.804545 PS=1.42 NRD=4.6886 NRS=4.6886
+ M=1 R=2.8 SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1038 N_Q_N_M1038_d N_A_1762_74#_M1038_g N_VPWR_M1032_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.3248 AS=0.243345 PD=2.82 PS=2.14545 NRD=1.7533 NRS=11.426 M=1
+ R=7.46667 SA=75000.4 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1030 N_VPWR_M1030_d N_A_1762_74#_M1030_g N_A_2556_112#_M1030_s VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.1596 AS=0.2436 PD=1.26429 PS=2.26 NRD=2.3443 NRS=2.3443 M=1
+ R=5.6 SA=75000.2 SB=75000.7 A=0.126 P=1.98 MULT=1
MM1021 N_Q_M1021_d N_A_2556_112#_M1021_g N_VPWR_M1030_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.3248 AS=0.2128 PD=2.82 PS=1.68571 NRD=1.7533 NRS=11.426 M=1
+ R=7.46667 SA=75000.6 SB=75000.2 A=0.168 P=2.54 MULT=1
DX42_noxref VNB VPB NWDIODE A=27.6026 P=33.49
*
.include "sky130_fd_sc_ls__sdfsbp_1.pxi.spice"
*
.ends
*
*
