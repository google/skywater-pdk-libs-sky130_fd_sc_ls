* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
M1000 X a_31_387# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=9.038e+11p ps=5.98e+06u
M1001 a_209_74# B1 a_131_74# VNB nshort w=640000u l=150000u
+  ad=8.448e+11p pd=5.2e+06u as=1.536e+11p ps=1.76e+06u
M1002 a_131_74# C1 a_31_387# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1003 a_209_74# A3 VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=6.202e+11p ps=4.62e+06u
M1004 X a_31_387# VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1005 VGND A2 a_209_74# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR C1 a_31_387# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=5.95e+11p ps=5.19e+06u
M1007 VPWR A1 a_536_387# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=4.2e+11p ps=2.84e+06u
M1008 a_320_387# A3 a_31_387# VPB phighvt w=1e+06u l=150000u
+  ad=9.3e+11p pd=3.86e+06u as=0p ps=0u
M1009 a_31_387# B1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_536_387# A2 a_320_387# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND A1 a_209_74# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
