* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__and3b_1 A_N B C VGND VNB VPB VPWR X
M1000 X a_266_94# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=1.0458e+12p ps=7.86e+06u
M1001 VPWR a_114_74# a_266_94# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=5.04e+11p ps=4.56e+06u
M1002 X a_266_94# VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=5.5385e+11p ps=4.28e+06u
M1003 a_353_94# a_114_74# a_266_94# VNB nshort w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=1.824e+11p ps=1.85e+06u
M1004 a_431_94# B a_353_94# VNB nshort w=640000u l=150000u
+  ad=2.496e+11p pd=2.06e+06u as=0p ps=0u
M1005 a_266_94# B VPWR VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_114_74# A_N VPWR VPB phighvt w=840000u l=150000u
+  ad=2.856e+11p pd=2.36e+06u as=0p ps=0u
M1007 VPWR C a_266_94# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_114_74# A_N VGND VNB nshort w=550000u l=150000u
+  ad=1.9525e+11p pd=1.81e+06u as=0p ps=0u
M1009 VGND C a_431_94# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
