* File: sky130_fd_sc_ls__o2111ai_1.pex.spice
* Created: Wed Sep  2 11:16:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__O2111AI_1%D1 1 3 4 6 7
c25 7 0 4.41642e-20 $X=0.72 $Y=1.295
r26 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.745
+ $Y=1.385 $X2=0.745 $Y2=1.385
r27 7 11 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.745 $Y=1.295
+ $X2=0.745 $Y2=1.385
r28 4 10 38.9026 $w=2.7e-07 $l=2.05122e-07 $layer=POLY_cond $X=0.835 $Y=1.22
+ $X2=0.745 $Y2=1.385
r29 4 6 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.835 $Y=1.22 $X2=0.835
+ $Y2=0.74
r30 1 10 77.2841 $w=2.7e-07 $l=4.15812e-07 $layer=POLY_cond $X=0.82 $Y=1.765
+ $X2=0.745 $Y2=1.385
r31 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.82 $Y=1.765
+ $X2=0.82 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__O2111AI_1%C1 1 3 4 6 7 8 9
c34 1 0 3.10838e-19 $X=1.225 $Y=1.22
r35 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.285
+ $Y=1.385 $X2=1.285 $Y2=1.385
r36 9 15 3.05058 $w=3.38e-07 $l=9e-08 $layer=LI1_cond $X=1.255 $Y=1.295
+ $X2=1.255 $Y2=1.385
r37 8 9 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=1.255 $Y=0.925
+ $X2=1.255 $Y2=1.295
r38 7 8 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=1.255 $Y=0.555
+ $X2=1.255 $Y2=0.925
r39 4 14 77.2841 $w=2.7e-07 $l=3.87427e-07 $layer=POLY_cond $X=1.27 $Y=1.765
+ $X2=1.285 $Y2=1.385
r40 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.27 $Y=1.765
+ $X2=1.27 $Y2=2.4
r41 1 14 38.9026 $w=2.7e-07 $l=1.92678e-07 $layer=POLY_cond $X=1.225 $Y=1.22
+ $X2=1.285 $Y2=1.385
r42 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.225 $Y=1.22 $X2=1.225
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__O2111AI_1%B1 1 3 4 6 7 11
c29 11 0 2.68987e-19 $X=1.825 $Y=1.385
c30 1 0 3.90916e-20 $X=1.765 $Y=1.22
r31 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.825
+ $Y=1.385 $X2=1.825 $Y2=1.385
r32 7 11 4.51633 $w=3.68e-07 $l=1.45e-07 $layer=LI1_cond $X=1.68 $Y=1.365
+ $X2=1.825 $Y2=1.365
r33 4 10 77.2841 $w=2.7e-07 $l=4.15812e-07 $layer=POLY_cond $X=1.9 $Y=1.765
+ $X2=1.825 $Y2=1.385
r34 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.9 $Y=1.765 $X2=1.9
+ $Y2=2.4
r35 1 10 38.9026 $w=2.7e-07 $l=1.92678e-07 $layer=POLY_cond $X=1.765 $Y=1.22
+ $X2=1.825 $Y2=1.385
r36 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.765 $Y=1.22 $X2=1.765
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__O2111AI_1%A2 1 3 4 6 7
c29 7 0 3.90916e-20 $X=2.64 $Y=1.295
c30 1 0 1.79793e-19 $X=2.275 $Y=1.22
r31 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.365
+ $Y=1.385 $X2=2.365 $Y2=1.385
r32 7 11 8.56545 $w=3.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.64 $Y=1.365
+ $X2=2.365 $Y2=1.365
r33 4 10 77.2841 $w=2.7e-07 $l=3.84968e-07 $layer=POLY_cond $X=2.375 $Y=1.765
+ $X2=2.365 $Y2=1.385
r34 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.375 $Y=1.765
+ $X2=2.375 $Y2=2.4
r35 1 10 38.9026 $w=2.7e-07 $l=2.05122e-07 $layer=POLY_cond $X=2.275 $Y=1.22
+ $X2=2.365 $Y2=1.385
r36 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.275 $Y=1.22 $X2=2.275
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__O2111AI_1%A1 1 3 4 6 7
c23 7 0 2.40942e-20 $X=3.12 $Y=1.295
r24 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.09
+ $Y=1.385 $X2=3.09 $Y2=1.385
r25 7 11 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=3.09 $Y=1.295 $X2=3.09
+ $Y2=1.385
r26 4 10 39.2524 $w=3.82e-07 $l=2.21371e-07 $layer=POLY_cond $X=2.865 $Y=1.22
+ $X2=2.997 $Y2=1.385
r27 4 6 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.865 $Y=1.22 $X2=2.865
+ $Y2=0.74
r28 1 10 66.3807 $w=3.82e-07 $l=4.55917e-07 $layer=POLY_cond $X=2.83 $Y=1.765
+ $X2=2.997 $Y2=1.385
r29 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.83 $Y=1.765
+ $X2=2.83 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__O2111AI_1%VPWR 1 2 3 12 18 22 24 29 30 31 37 41 47
+ 51
r40 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r41 45 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r42 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r43 42 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.815 $Y=3.33
+ $X2=1.65 $Y2=3.33
r44 42 44 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=1.815 $Y=3.33
+ $X2=2.64 $Y2=3.33
r45 41 50 4.67962 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=2.89 $Y=3.33
+ $X2=3.125 $Y2=3.33
r46 41 44 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.89 $Y=3.33
+ $X2=2.64 $Y2=3.33
r47 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r48 37 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.485 $Y=3.33
+ $X2=1.65 $Y2=3.33
r49 37 39 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.485 $Y=3.33
+ $X2=1.2 $Y2=3.33
r50 35 40 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r51 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r52 31 45 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r53 31 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r54 31 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r55 29 34 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=0.38 $Y=3.33
+ $X2=0.24 $Y2=3.33
r56 29 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.38 $Y=3.33
+ $X2=0.545 $Y2=3.33
r57 28 39 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=0.71 $Y=3.33 $X2=1.2
+ $Y2=3.33
r58 28 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.71 $Y=3.33
+ $X2=0.545 $Y2=3.33
r59 24 27 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=3.055 $Y=1.985
+ $X2=3.055 $Y2=2.815
r60 22 50 3.08656 $w=3.3e-07 $l=1.14782e-07 $layer=LI1_cond $X=3.055 $Y=3.245
+ $X2=3.125 $Y2=3.33
r61 22 27 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.055 $Y=3.245
+ $X2=3.055 $Y2=2.815
r62 18 21 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.65 $Y=2.145
+ $X2=1.65 $Y2=2.825
r63 16 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.65 $Y=3.245
+ $X2=1.65 $Y2=3.33
r64 16 21 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=1.65 $Y=3.245
+ $X2=1.65 $Y2=2.825
r65 12 15 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.545 $Y=2.145
+ $X2=0.545 $Y2=2.825
r66 10 30 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.545 $Y=3.245
+ $X2=0.545 $Y2=3.33
r67 10 15 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=0.545 $Y=3.245
+ $X2=0.545 $Y2=2.825
r68 3 27 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.905
+ $Y=1.84 $X2=3.055 $Y2=2.815
r69 3 24 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.905
+ $Y=1.84 $X2=3.055 $Y2=1.985
r70 2 21 400 $w=1.7e-07 $l=1.12723e-06 $layer=licon1_PDIFF $count=1 $X=1.345
+ $Y=1.84 $X2=1.65 $Y2=2.825
r71 2 18 400 $w=1.7e-07 $l=4.31335e-07 $layer=licon1_PDIFF $count=1 $X=1.345
+ $Y=1.84 $X2=1.65 $Y2=2.145
r72 1 15 400 $w=1.7e-07 $l=1.05501e-06 $layer=licon1_PDIFF $count=1 $X=0.4
+ $Y=1.84 $X2=0.545 $Y2=2.825
r73 1 12 400 $w=1.7e-07 $l=3.70473e-07 $layer=licon1_PDIFF $count=1 $X=0.4
+ $Y=1.84 $X2=0.545 $Y2=2.145
.ends

.subckt PM_SKY130_FD_SC_LS__O2111AI_1%Y 1 2 3 11 12 13 14 18 25 28 29 30 31 36
r51 31 44 1.05972 $w=4.33e-07 $l=4e-08 $layer=LI1_cond $X=1.097 $Y=2.775
+ $X2=1.097 $Y2=2.815
r52 30 31 9.80239 $w=4.33e-07 $l=3.7e-07 $layer=LI1_cond $X=1.097 $Y=2.405
+ $X2=1.097 $Y2=2.775
r53 29 30 9.80239 $w=4.33e-07 $l=3.7e-07 $layer=LI1_cond $X=1.097 $Y=2.035
+ $X2=1.097 $Y2=2.405
r54 29 36 1.32465 $w=4.33e-07 $l=5e-08 $layer=LI1_cond $X=1.097 $Y=2.035
+ $X2=1.097 $Y2=1.985
r55 27 36 2.51683 $w=4.33e-07 $l=9.5e-08 $layer=LI1_cond $X=1.097 $Y=1.89
+ $X2=1.097 $Y2=1.985
r56 27 28 1.70358 $w=4.35e-07 $l=8.5e-08 $layer=LI1_cond $X=1.097 $Y=1.89
+ $X2=1.097 $Y2=1.805
r57 22 25 7.61141 $w=6.58e-07 $l=4.2e-07 $layer=LI1_cond $X=0.2 $Y=0.68 $X2=0.62
+ $Y2=0.68
r58 18 20 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=2.15 $Y=1.985
+ $X2=2.15 $Y2=2.815
r59 16 18 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=2.15 $Y=1.89
+ $X2=2.15 $Y2=1.985
r60 15 28 10.3577 $w=1.7e-07 $l=2.18e-07 $layer=LI1_cond $X=1.315 $Y=1.805
+ $X2=1.097 $Y2=1.805
r61 14 16 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.985 $Y=1.805
+ $X2=2.15 $Y2=1.89
r62 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.985 $Y=1.805
+ $X2=1.315 $Y2=1.805
r63 12 28 10.3577 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=0.88 $Y=1.805
+ $X2=1.097 $Y2=1.805
r64 12 13 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=0.88 $Y=1.805
+ $X2=0.285 $Y2=1.805
r65 11 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.2 $Y=1.72
+ $X2=0.285 $Y2=1.805
r66 10 22 8.93547 $w=1.7e-07 $l=3.3e-07 $layer=LI1_cond $X=0.2 $Y=1.01 $X2=0.2
+ $Y2=0.68
r67 10 11 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=0.2 $Y=1.01 $X2=0.2
+ $Y2=1.72
r68 3 20 400 $w=1.7e-07 $l=1.05889e-06 $layer=licon1_PDIFF $count=1 $X=1.975
+ $Y=1.84 $X2=2.15 $Y2=2.815
r69 3 18 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=1.975
+ $Y=1.84 $X2=2.15 $Y2=1.985
r70 2 44 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=0.895
+ $Y=1.84 $X2=1.045 $Y2=2.815
r71 2 36 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=0.895
+ $Y=1.84 $X2=1.045 $Y2=1.985
r72 1 25 45.5 $w=1.7e-07 $l=5.52766e-07 $layer=licon1_NDIFF $count=4 $X=0.135
+ $Y=0.37 $X2=0.62 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__O2111AI_1%A_368_74# 1 2 7 9 11 15
c28 7 0 1.53386e-19 $X=1.99 $Y=0.84
r29 13 15 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=3.08 $Y=0.84
+ $X2=3.08 $Y2=0.515
r30 12 18 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.155 $Y=0.925
+ $X2=1.99 $Y2=0.925
r31 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.915 $Y=0.925
+ $X2=3.08 $Y2=0.84
r32 11 12 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=2.915 $Y=0.925
+ $X2=2.155 $Y2=0.925
r33 7 18 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.99 $Y=0.84 $X2=1.99
+ $Y2=0.925
r34 7 9 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=1.99 $Y=0.84 $X2=1.99
+ $Y2=0.515
r35 2 15 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.94
+ $Y=0.37 $X2=3.08 $Y2=0.515
r36 1 18 182 $w=1.7e-07 $l=6.2552e-07 $layer=licon1_NDIFF $count=1 $X=1.84
+ $Y=0.37 $X2=1.99 $Y2=0.925
r37 1 9 182 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_NDIFF $count=1 $X=1.84
+ $Y=0.37 $X2=1.99 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__O2111AI_1%VGND 1 6 8 10 20 21 24
r31 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r32 21 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r33 20 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r34 18 24 10.1275 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=2.745 $Y=0 $X2=2.535
+ $Y2=0
r35 18 20 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=2.745 $Y=0 $X2=3.12
+ $Y2=0
r36 17 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r37 16 17 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r38 12 16 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=2.16
+ $Y2=0
r39 12 13 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r40 10 24 10.1275 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=2.325 $Y=0 $X2=2.535
+ $Y2=0
r41 10 16 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.325 $Y=0 $X2=2.16
+ $Y2=0
r42 8 17 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r43 8 13 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.24
+ $Y2=0
r44 4 24 1.60615 $w=4.2e-07 $l=8.5e-08 $layer=LI1_cond $X=2.535 $Y=0.085
+ $X2=2.535 $Y2=0
r45 4 6 11.7988 $w=4.18e-07 $l=4.3e-07 $layer=LI1_cond $X=2.535 $Y=0.085
+ $X2=2.535 $Y2=0.515
r46 1 6 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=2.35
+ $Y=0.37 $X2=2.535 $Y2=0.515
.ends

