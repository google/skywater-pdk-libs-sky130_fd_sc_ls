* File: sky130_fd_sc_ls__sdfbbn_2.pxi.spice
* Created: Wed Sep  2 11:26:39 2020
* 
x_PM_SKY130_FD_SC_LS__SDFBBN_2%SCD N_SCD_c_377_n N_SCD_c_382_n N_SCD_M1028_g
+ N_SCD_M1004_g SCD SCD N_SCD_c_378_n N_SCD_c_379_n N_SCD_c_380_n
+ PM_SKY130_FD_SC_LS__SDFBBN_2%SCD
x_PM_SKY130_FD_SC_LS__SDFBBN_2%D N_D_c_409_n N_D_M1000_g N_D_c_410_n N_D_M1042_g
+ N_D_c_411_n D N_D_c_408_n PM_SKY130_FD_SC_LS__SDFBBN_2%D
x_PM_SKY130_FD_SC_LS__SDFBBN_2%A_341_410# N_A_341_410#_M1037_d
+ N_A_341_410#_M1024_d N_A_341_410#_c_470_n N_A_341_410#_M1015_g
+ N_A_341_410#_c_471_n N_A_341_410#_c_472_n N_A_341_410#_M1025_g
+ N_A_341_410#_c_473_n N_A_341_410#_c_466_n N_A_341_410#_c_475_n
+ N_A_341_410#_c_467_n N_A_341_410#_c_468_n N_A_341_410#_c_469_n
+ N_A_341_410#_c_477_n N_A_341_410#_c_501_p
+ PM_SKY130_FD_SC_LS__SDFBBN_2%A_341_410#
x_PM_SKY130_FD_SC_LS__SDFBBN_2%SCE N_SCE_M1032_g N_SCE_c_558_n N_SCE_c_559_n
+ N_SCE_M1029_g N_SCE_c_548_n N_SCE_c_549_n N_SCE_c_560_n N_SCE_M1024_g
+ N_SCE_M1037_g N_SCE_c_551_n N_SCE_c_552_n N_SCE_c_561_n N_SCE_c_562_n
+ N_SCE_c_553_n N_SCE_c_554_n N_SCE_c_555_n SCE SCE N_SCE_c_556_n N_SCE_c_557_n
+ PM_SKY130_FD_SC_LS__SDFBBN_2%SCE
x_PM_SKY130_FD_SC_LS__SDFBBN_2%CLK_N N_CLK_N_c_651_n N_CLK_N_M1035_g
+ N_CLK_N_c_652_n N_CLK_N_M1036_g CLK_N N_CLK_N_c_653_n
+ PM_SKY130_FD_SC_LS__SDFBBN_2%CLK_N
x_PM_SKY130_FD_SC_LS__SDFBBN_2%A_1007_366# N_A_1007_366#_M1017_d
+ N_A_1007_366#_M1034_s N_A_1007_366#_M1049_d N_A_1007_366#_c_700_n
+ N_A_1007_366#_M1045_g N_A_1007_366#_c_691_n N_A_1007_366#_c_692_n
+ N_A_1007_366#_c_693_n N_A_1007_366#_c_694_n N_A_1007_366#_M1027_g
+ N_A_1007_366#_M1046_g N_A_1007_366#_c_702_n N_A_1007_366#_M1009_g
+ N_A_1007_366#_c_703_n N_A_1007_366#_c_704_n N_A_1007_366#_c_705_n
+ N_A_1007_366#_c_706_n N_A_1007_366#_c_696_n N_A_1007_366#_c_756_p
+ N_A_1007_366#_c_697_n N_A_1007_366#_c_770_p N_A_1007_366#_c_708_n
+ N_A_1007_366#_c_698_n N_A_1007_366#_c_699_n N_A_1007_366#_c_711_n
+ N_A_1007_366#_c_712_n N_A_1007_366#_c_713_n N_A_1007_366#_c_739_p
+ N_A_1007_366#_c_758_p N_A_1007_366#_c_714_n N_A_1007_366#_c_715_n
+ PM_SKY130_FD_SC_LS__SDFBBN_2%A_1007_366#
x_PM_SKY130_FD_SC_LS__SDFBBN_2%A_868_368# N_A_868_368#_M1043_d
+ N_A_868_368#_M1048_d N_A_868_368#_c_905_n N_A_868_368#_c_906_n
+ N_A_868_368#_M1039_g N_A_868_368#_M1006_g N_A_868_368#_c_907_n
+ N_A_868_368#_c_908_n N_A_868_368#_M1010_g N_A_868_368#_M1012_g
+ N_A_868_368#_c_909_n N_A_868_368#_c_929_n N_A_868_368#_c_891_n
+ N_A_868_368#_c_892_n N_A_868_368#_c_893_n N_A_868_368#_c_910_n
+ N_A_868_368#_c_894_n N_A_868_368#_c_895_n N_A_868_368#_c_896_n
+ N_A_868_368#_c_897_n N_A_868_368#_c_898_n N_A_868_368#_c_899_n
+ N_A_868_368#_c_900_n N_A_868_368#_c_988_p N_A_868_368#_c_901_n
+ N_A_868_368#_c_902_n N_A_868_368#_c_903_n N_A_868_368#_c_904_n
+ PM_SKY130_FD_SC_LS__SDFBBN_2%A_868_368#
x_PM_SKY130_FD_SC_LS__SDFBBN_2%A_1154_464# N_A_1154_464#_M1016_d
+ N_A_1154_464#_M1039_d N_A_1154_464#_c_1099_n N_A_1154_464#_c_1100_n
+ N_A_1154_464#_c_1101_n N_A_1154_464#_c_1109_n N_A_1154_464#_M1034_g
+ N_A_1154_464#_c_1102_n N_A_1154_464#_M1017_g N_A_1154_464#_c_1103_n
+ N_A_1154_464#_c_1110_n N_A_1154_464#_c_1111_n N_A_1154_464#_c_1112_n
+ N_A_1154_464#_c_1104_n N_A_1154_464#_c_1105_n N_A_1154_464#_c_1106_n
+ N_A_1154_464#_c_1113_n N_A_1154_464#_c_1107_n
+ PM_SKY130_FD_SC_LS__SDFBBN_2%A_1154_464#
x_PM_SKY130_FD_SC_LS__SDFBBN_2%A_1643_257# N_A_1643_257#_M1005_s
+ N_A_1643_257#_M1026_s N_A_1643_257#_c_1217_n N_A_1643_257#_M1030_g
+ N_A_1643_257#_M1018_g N_A_1643_257#_c_1201_n N_A_1643_257#_M1038_g
+ N_A_1643_257#_c_1219_n N_A_1643_257#_M1014_g N_A_1643_257#_c_1202_n
+ N_A_1643_257#_c_1203_n N_A_1643_257#_c_1204_n N_A_1643_257#_c_1205_n
+ N_A_1643_257#_c_1206_n N_A_1643_257#_c_1207_n N_A_1643_257#_c_1251_n
+ N_A_1643_257#_c_1301_p N_A_1643_257#_c_1252_n N_A_1643_257#_c_1277_p
+ N_A_1643_257#_c_1208_n N_A_1643_257#_c_1209_n N_A_1643_257#_c_1210_n
+ N_A_1643_257#_c_1211_n N_A_1643_257#_c_1212_n N_A_1643_257#_c_1255_n
+ N_A_1643_257#_c_1213_n N_A_1643_257#_c_1291_p N_A_1643_257#_c_1214_n
+ N_A_1643_257#_c_1215_n N_A_1643_257#_c_1223_n N_A_1643_257#_c_1216_n
+ PM_SKY130_FD_SC_LS__SDFBBN_2%A_1643_257#
x_PM_SKY130_FD_SC_LS__SDFBBN_2%SET_B N_SET_B_c_1415_n N_SET_B_c_1416_n
+ N_SET_B_M1049_g N_SET_B_M1047_g N_SET_B_c_1407_n N_SET_B_M1002_g
+ N_SET_B_c_1418_n N_SET_B_M1011_g N_SET_B_c_1408_n N_SET_B_c_1420_n
+ N_SET_B_c_1409_n SET_B N_SET_B_c_1411_n N_SET_B_c_1412_n N_SET_B_c_1413_n
+ N_SET_B_c_1414_n PM_SKY130_FD_SC_LS__SDFBBN_2%SET_B
x_PM_SKY130_FD_SC_LS__SDFBBN_2%A_688_98# N_A_688_98#_M1035_s N_A_688_98#_M1036_s
+ N_A_688_98#_c_1560_n N_A_688_98#_M1048_g N_A_688_98#_M1043_g
+ N_A_688_98#_c_1547_n N_A_688_98#_c_1548_n N_A_688_98#_M1016_g
+ N_A_688_98#_M1013_g N_A_688_98#_c_1550_n N_A_688_98#_M1020_g
+ N_A_688_98#_c_1552_n N_A_688_98#_c_1553_n N_A_688_98#_c_1562_n
+ N_A_688_98#_c_1563_n N_A_688_98#_c_1564_n N_A_688_98#_M1031_g
+ N_A_688_98#_c_1554_n N_A_688_98#_c_1565_n N_A_688_98#_c_1555_n
+ N_A_688_98#_c_1556_n N_A_688_98#_c_1567_n N_A_688_98#_c_1568_n
+ N_A_688_98#_c_1586_n N_A_688_98#_c_1569_n N_A_688_98#_c_1557_n
+ N_A_688_98#_c_1558_n N_A_688_98#_c_1559_n
+ PM_SKY130_FD_SC_LS__SDFBBN_2%A_688_98#
x_PM_SKY130_FD_SC_LS__SDFBBN_2%A_2216_410# N_A_2216_410#_M1038_d
+ N_A_2216_410#_M1011_s N_A_2216_410#_M1051_d N_A_2216_410#_c_1742_n
+ N_A_2216_410#_M1008_g N_A_2216_410#_c_1743_n N_A_2216_410#_c_1727_n
+ N_A_2216_410#_M1044_g N_A_2216_410#_c_1728_n N_A_2216_410#_c_1729_n
+ N_A_2216_410#_M1003_g N_A_2216_410#_c_1745_n N_A_2216_410#_M1023_g
+ N_A_2216_410#_M1021_g N_A_2216_410#_c_1746_n N_A_2216_410#_M1033_g
+ N_A_2216_410#_c_1732_n N_A_2216_410#_c_1733_n N_A_2216_410#_M1019_g
+ N_A_2216_410#_c_1735_n N_A_2216_410#_M1050_g N_A_2216_410#_c_1736_n
+ N_A_2216_410#_c_1749_n N_A_2216_410#_c_1769_n N_A_2216_410#_c_1737_n
+ N_A_2216_410#_c_1750_n N_A_2216_410#_c_1751_n N_A_2216_410#_c_1738_n
+ N_A_2216_410#_c_1752_n N_A_2216_410#_c_1753_n N_A_2216_410#_c_1754_n
+ N_A_2216_410#_c_1777_n N_A_2216_410#_c_1778_n N_A_2216_410#_c_1739_n
+ N_A_2216_410#_c_1740_n N_A_2216_410#_c_1741_n
+ PM_SKY130_FD_SC_LS__SDFBBN_2%A_2216_410#
x_PM_SKY130_FD_SC_LS__SDFBBN_2%A_1997_82# N_A_1997_82#_M1020_d
+ N_A_1997_82#_M1010_d N_A_1997_82#_c_1935_n N_A_1997_82#_M1051_g
+ N_A_1997_82#_M1007_g N_A_1997_82#_c_1942_n N_A_1997_82#_c_1943_n
+ N_A_1997_82#_c_1944_n N_A_1997_82#_c_1945_n N_A_1997_82#_c_1937_n
+ N_A_1997_82#_c_1938_n N_A_1997_82#_c_1947_n N_A_1997_82#_c_1948_n
+ N_A_1997_82#_c_1949_n N_A_1997_82#_c_1939_n N_A_1997_82#_c_1950_n
+ N_A_1997_82#_c_1951_n N_A_1997_82#_c_1940_n
+ PM_SKY130_FD_SC_LS__SDFBBN_2%A_1997_82#
x_PM_SKY130_FD_SC_LS__SDFBBN_2%RESET_B N_RESET_B_c_2095_n N_RESET_B_M1026_g
+ N_RESET_B_M1005_g RESET_B PM_SKY130_FD_SC_LS__SDFBBN_2%RESET_B
x_PM_SKY130_FD_SC_LS__SDFBBN_2%A_3272_94# N_A_3272_94#_M1019_s
+ N_A_3272_94#_M1050_s N_A_3272_94#_c_2133_n N_A_3272_94#_M1001_g
+ N_A_3272_94#_c_2127_n N_A_3272_94#_M1022_g N_A_3272_94#_c_2134_n
+ N_A_3272_94#_M1040_g N_A_3272_94#_c_2128_n N_A_3272_94#_M1041_g
+ N_A_3272_94#_c_2129_n N_A_3272_94#_c_2135_n N_A_3272_94#_c_2130_n
+ N_A_3272_94#_c_2131_n N_A_3272_94#_c_2132_n
+ PM_SKY130_FD_SC_LS__SDFBBN_2%A_3272_94#
x_PM_SKY130_FD_SC_LS__SDFBBN_2%A_27_464# N_A_27_464#_M1028_s N_A_27_464#_M1015_d
+ N_A_27_464#_c_2193_n N_A_27_464#_c_2228_p N_A_27_464#_c_2194_n
+ N_A_27_464#_c_2195_n N_A_27_464#_c_2196_n N_A_27_464#_c_2197_n
+ PM_SKY130_FD_SC_LS__SDFBBN_2%A_27_464#
x_PM_SKY130_FD_SC_LS__SDFBBN_2%VPWR N_VPWR_M1028_d N_VPWR_M1024_s N_VPWR_M1036_d
+ N_VPWR_M1045_s N_VPWR_M1030_d N_VPWR_M1009_s N_VPWR_M1008_d N_VPWR_M1011_d
+ N_VPWR_M1026_d N_VPWR_M1033_s N_VPWR_M1050_d N_VPWR_M1040_d N_VPWR_c_2235_n
+ N_VPWR_c_2236_n N_VPWR_c_2237_n N_VPWR_c_2238_n N_VPWR_c_2239_n
+ N_VPWR_c_2240_n N_VPWR_c_2241_n N_VPWR_c_2242_n N_VPWR_c_2243_n
+ N_VPWR_c_2244_n N_VPWR_c_2245_n N_VPWR_c_2246_n N_VPWR_c_2247_n
+ N_VPWR_c_2248_n N_VPWR_c_2249_n N_VPWR_c_2250_n N_VPWR_c_2251_n
+ N_VPWR_c_2252_n N_VPWR_c_2253_n N_VPWR_c_2254_n VPWR N_VPWR_c_2255_n
+ N_VPWR_c_2256_n N_VPWR_c_2257_n N_VPWR_c_2258_n N_VPWR_c_2259_n
+ N_VPWR_c_2260_n N_VPWR_c_2261_n N_VPWR_c_2262_n N_VPWR_c_2263_n
+ N_VPWR_c_2264_n N_VPWR_c_2265_n N_VPWR_c_2266_n N_VPWR_c_2267_n
+ N_VPWR_c_2268_n N_VPWR_c_2269_n N_VPWR_c_2270_n N_VPWR_c_2234_n
+ PM_SKY130_FD_SC_LS__SDFBBN_2%VPWR
x_PM_SKY130_FD_SC_LS__SDFBBN_2%A_197_119# N_A_197_119#_M1032_d
+ N_A_197_119#_M1006_d N_A_197_119#_M1000_d N_A_197_119#_M1013_d
+ N_A_197_119#_c_2470_n N_A_197_119#_c_2481_n N_A_197_119#_c_2482_n
+ N_A_197_119#_c_2446_n N_A_197_119#_c_2471_n N_A_197_119#_c_2472_n
+ N_A_197_119#_c_2447_n N_A_197_119#_c_2448_n N_A_197_119#_c_2449_n
+ N_A_197_119#_c_2450_n N_A_197_119#_c_2451_n N_A_197_119#_c_2452_n
+ N_A_197_119#_c_2453_n N_A_197_119#_c_2454_n N_A_197_119#_c_2546_n
+ N_A_197_119#_c_2455_n N_A_197_119#_c_2456_n N_A_197_119#_c_2457_n
+ N_A_197_119#_c_2458_n N_A_197_119#_c_2459_n N_A_197_119#_c_2460_n
+ N_A_197_119#_c_2461_n N_A_197_119#_c_2462_n N_A_197_119#_c_2463_n
+ N_A_197_119#_c_2464_n N_A_197_119#_c_2474_n N_A_197_119#_c_2465_n
+ N_A_197_119#_c_2466_n N_A_197_119#_c_2467_n N_A_197_119#_c_2468_n
+ N_A_197_119#_c_2476_n N_A_197_119#_c_2478_n N_A_197_119#_c_2469_n
+ N_A_197_119#_c_2477_n PM_SKY130_FD_SC_LS__SDFBBN_2%A_197_119#
x_PM_SKY130_FD_SC_LS__SDFBBN_2%Q_N N_Q_N_M1003_s N_Q_N_M1023_d N_Q_N_c_2675_n
+ N_Q_N_c_2678_n N_Q_N_c_2676_n Q_N N_Q_N_c_2677_n
+ PM_SKY130_FD_SC_LS__SDFBBN_2%Q_N
x_PM_SKY130_FD_SC_LS__SDFBBN_2%Q N_Q_M1022_d N_Q_M1001_s N_Q_c_2705_n
+ N_Q_c_2712_n Q Q N_Q_c_2706_n PM_SKY130_FD_SC_LS__SDFBBN_2%Q
x_PM_SKY130_FD_SC_LS__SDFBBN_2%VGND N_VGND_M1004_s N_VGND_M1025_d N_VGND_M1035_d
+ N_VGND_M1027_s N_VGND_M1047_d N_VGND_M1044_d N_VGND_M1005_d N_VGND_M1021_d
+ N_VGND_M1019_d N_VGND_M1041_s N_VGND_c_2732_n N_VGND_c_2733_n N_VGND_c_2734_n
+ N_VGND_c_2735_n N_VGND_c_2736_n N_VGND_c_2737_n N_VGND_c_2738_n
+ N_VGND_c_2739_n N_VGND_c_2740_n N_VGND_c_2741_n N_VGND_c_2742_n
+ N_VGND_c_2743_n N_VGND_c_2744_n N_VGND_c_2745_n N_VGND_c_2746_n
+ N_VGND_c_2747_n N_VGND_c_2748_n N_VGND_c_2749_n VGND N_VGND_c_2750_n
+ N_VGND_c_2751_n N_VGND_c_2752_n N_VGND_c_2753_n N_VGND_c_2754_n
+ N_VGND_c_2755_n N_VGND_c_2756_n N_VGND_c_2757_n N_VGND_c_2758_n
+ N_VGND_c_2759_n PM_SKY130_FD_SC_LS__SDFBBN_2%VGND
x_PM_SKY130_FD_SC_LS__SDFBBN_2%A_1473_73# N_A_1473_73#_M1017_s
+ N_A_1473_73#_M1018_d N_A_1473_73#_c_2925_n N_A_1473_73#_c_2926_n
+ N_A_1473_73#_c_2927_n N_A_1473_73#_c_2928_n
+ PM_SKY130_FD_SC_LS__SDFBBN_2%A_1473_73#
x_PM_SKY130_FD_SC_LS__SDFBBN_2%A_2452_74# N_A_2452_74#_M1002_d
+ N_A_2452_74#_M1007_d N_A_2452_74#_c_2972_n N_A_2452_74#_c_2973_n
+ N_A_2452_74#_c_2974_n PM_SKY130_FD_SC_LS__SDFBBN_2%A_2452_74#
cc_1 VNB N_SCD_c_377_n 0.0295087f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.948
cc_2 VNB N_SCD_c_378_n 0.0223236f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.29
cc_3 VNB N_SCD_c_379_n 0.0240257f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.29
cc_4 VNB N_SCD_c_380_n 0.0213135f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.125
cc_5 VNB N_D_M1042_g 0.0352886f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.805
cc_6 VNB D 0.00165697f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_D_c_408_n 0.0266813f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.97
cc_8 VNB N_A_341_410#_M1025_g 0.0473704f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.29
cc_9 VNB N_A_341_410#_c_466_n 0.0101103f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.97
cc_10 VNB N_A_341_410#_c_467_n 0.00177782f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_341_410#_c_468_n 0.0182972f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.665
cc_12 VNB N_A_341_410#_c_469_n 0.0148708f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_SCE_M1032_g 0.0337655f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.64
cc_14 VNB N_SCE_c_548_n 0.145345f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_15 VNB N_SCE_c_549_n 0.0125534f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_SCE_M1037_g 0.0278614f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.97
cc_17 VNB N_SCE_c_551_n 0.0319917f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.97
cc_18 VNB N_SCE_c_552_n 0.00799454f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.29
cc_19 VNB N_SCE_c_553_n 0.0210745f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.665
cc_20 VNB N_SCE_c_554_n 0.022701f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_SCE_c_555_n 0.00185471f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_SCE_c_556_n 0.0170718f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_SCE_c_557_n 0.00847737f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_CLK_N_c_651_n 0.0210886f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.312
cc_25 VNB N_CLK_N_c_652_n 0.0251987f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.64
cc_26 VNB N_CLK_N_c_653_n 0.00469313f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_1007_366#_c_691_n 0.0243827f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.29
cc_28 VNB N_A_1007_366#_c_692_n 0.0306125f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.29
cc_29 VNB N_A_1007_366#_c_693_n 0.00958068f $X=-0.19 $Y=-0.245 $X2=0.407
+ $Y2=1.125
cc_30 VNB N_A_1007_366#_c_694_n 0.015556f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.97
cc_31 VNB N_A_1007_366#_M1046_g 0.0343259f $X=-0.19 $Y=-0.245 $X2=0.337
+ $Y2=1.295
cc_32 VNB N_A_1007_366#_c_696_n 0.00287006f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_1007_366#_c_697_n 0.00167086f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_1007_366#_c_698_n 0.00297418f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_1007_366#_c_699_n 0.0177963f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_868_368#_M1006_g 0.0390394f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.29
cc_37 VNB N_A_868_368#_M1012_g 0.0353628f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_868_368#_c_891_n 0.0148677f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_868_368#_c_892_n 0.00996027f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_868_368#_c_893_n 0.029767f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_868_368#_c_894_n 0.00368308f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_868_368#_c_895_n 0.00651249f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_868_368#_c_896_n 8.9717e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_868_368#_c_897_n 0.0118036f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_868_368#_c_898_n 0.00205349f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_868_368#_c_899_n 0.0425307f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_868_368#_c_900_n 0.00227713f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_868_368#_c_901_n 0.00417801f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_868_368#_c_902_n 0.0132802f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_868_368#_c_903_n 0.0203321f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_868_368#_c_904_n 0.00547296f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_1154_464#_c_1099_n 0.0290087f $X=-0.19 $Y=-0.245 $X2=0.52
+ $Y2=0.805
cc_53 VNB N_A_1154_464#_c_1100_n 0.0172355f $X=-0.19 $Y=-0.245 $X2=0.52
+ $Y2=0.805
cc_54 VNB N_A_1154_464#_c_1101_n 0.01189f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_55 VNB N_A_1154_464#_c_1102_n 0.0161432f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.29
cc_56 VNB N_A_1154_464#_c_1103_n 0.00562192f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.97
cc_57 VNB N_A_1154_464#_c_1104_n 0.0041336f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_1154_464#_c_1105_n 0.0103846f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_1154_464#_c_1106_n 0.00178644f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_1154_464#_c_1107_n 0.0169021f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_1643_257#_c_1201_n 0.00627308f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.29
cc_62 VNB N_A_1643_257#_c_1202_n 0.0161443f $X=-0.19 $Y=-0.245 $X2=0.337
+ $Y2=1.295
cc_63 VNB N_A_1643_257#_c_1203_n 0.0129324f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_1643_257#_c_1204_n 0.00628362f $X=-0.19 $Y=-0.245 $X2=0.337
+ $Y2=1.97
cc_65 VNB N_A_1643_257#_c_1205_n 0.001484f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_1643_257#_c_1206_n 0.0159308f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_1643_257#_c_1207_n 0.0028989f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_1643_257#_c_1208_n 0.0204306f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_1643_257#_c_1209_n 0.00759669f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_1643_257#_c_1210_n 0.00514335f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_1643_257#_c_1211_n 0.00582598f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_1643_257#_c_1212_n 0.0152277f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_1643_257#_c_1213_n 0.00405091f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_1643_257#_c_1214_n 0.0316147f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_1643_257#_c_1215_n 0.00578916f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_1643_257#_c_1216_n 0.0162265f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_SET_B_M1047_g 0.0248332f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.805
cc_78 VNB N_SET_B_c_1407_n 0.00552638f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_SET_B_c_1408_n 0.0139983f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.97
cc_80 VNB N_SET_B_c_1409_n 0.00175115f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.295
cc_81 VNB SET_B 0.00247325f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.665
cc_82 VNB N_SET_B_c_1411_n 0.019444f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_SET_B_c_1412_n 0.0297443f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_SET_B_c_1413_n 0.00686408f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_SET_B_c_1414_n 0.0186418f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_688_98#_M1043_g 0.0238035f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.29
cc_87 VNB N_A_688_98#_c_1547_n 0.100209f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.29
cc_88 VNB N_A_688_98#_c_1548_n 0.0125579f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.29
cc_89 VNB N_A_688_98#_M1016_g 0.0552224f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.97
cc_90 VNB N_A_688_98#_c_1550_n 0.263428f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_688_98#_M1020_g 0.0174579f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_688_98#_c_1552_n 0.0501571f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_688_98#_c_1553_n 0.00977566f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_688_98#_c_1554_n 0.00749069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_688_98#_c_1555_n 0.0235246f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_688_98#_c_1556_n 0.00223776f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_688_98#_c_1557_n 0.00508715f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_A_688_98#_c_1558_n 0.0440049f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_A_688_98#_c_1559_n 0.00200664f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_A_2216_410#_c_1727_n 0.0152288f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.29
cc_101 VNB N_A_2216_410#_c_1728_n 0.0292958f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.97
cc_102 VNB N_A_2216_410#_c_1729_n 0.0263378f $X=-0.19 $Y=-0.245 $X2=0.337
+ $Y2=1.29
cc_103 VNB N_A_2216_410#_M1003_g 0.0262134f $X=-0.19 $Y=-0.245 $X2=0.337
+ $Y2=1.665
cc_104 VNB N_A_2216_410#_M1021_g 0.0261462f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_A_2216_410#_c_1732_n 0.0745959f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_A_2216_410#_c_1733_n 0.0411399f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_A_2216_410#_M1019_g 0.0279425f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_A_2216_410#_c_1735_n 0.0130722f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_A_2216_410#_c_1736_n 0.0160979f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_A_2216_410#_c_1737_n 0.0169864f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_A_2216_410#_c_1738_n 0.00916846f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_A_2216_410#_c_1739_n 0.00593009f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_A_2216_410#_c_1740_n 0.00559626f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_A_2216_410#_c_1741_n 0.0215319f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_A_1997_82#_c_1935_n 0.0203002f $X=-0.19 $Y=-0.245 $X2=0.52
+ $Y2=0.805
cc_116 VNB N_A_1997_82#_M1007_g 0.0337407f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_A_1997_82#_c_1937_n 0.00577836f $X=-0.19 $Y=-0.245 $X2=0.337
+ $Y2=1.97
cc_118 VNB N_A_1997_82#_c_1938_n 0.00459897f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_A_1997_82#_c_1939_n 0.0147718f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_A_1997_82#_c_1940_n 0.00165779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_RESET_B_c_2095_n 0.0148491f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.312
cc_122 VNB N_RESET_B_M1005_g 0.0257887f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.125
cc_123 VNB RESET_B 0.00217311f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.805
cc_124 VNB N_A_3272_94#_c_2127_n 0.0185525f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.58
cc_125 VNB N_A_3272_94#_c_2128_n 0.0199293f $X=-0.19 $Y=-0.245 $X2=0.407
+ $Y2=1.125
cc_126 VNB N_A_3272_94#_c_2129_n 0.00721335f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_A_3272_94#_c_2130_n 0.00785255f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_A_3272_94#_c_2131_n 0.00216442f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_A_3272_94#_c_2132_n 0.0801406f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_VPWR_c_2234_n 0.760753f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_A_197_119#_c_2446_n 0.00136531f $X=-0.19 $Y=-0.245 $X2=0.337
+ $Y2=1.29
cc_132 VNB N_A_197_119#_c_2447_n 0.0083752f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_A_197_119#_c_2448_n 0.00228786f $X=-0.19 $Y=-0.245 $X2=0.337
+ $Y2=1.97
cc_134 VNB N_A_197_119#_c_2449_n 0.00287473f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_A_197_119#_c_2450_n 0.015027f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_A_197_119#_c_2451_n 0.00245103f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_A_197_119#_c_2452_n 0.0155526f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB N_A_197_119#_c_2453_n 0.00159638f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VNB N_A_197_119#_c_2454_n 0.00354964f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_A_197_119#_c_2455_n 0.00408608f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_141 VNB N_A_197_119#_c_2456_n 0.00104052f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_142 VNB N_A_197_119#_c_2457_n 0.0156551f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_143 VNB N_A_197_119#_c_2458_n 0.00291013f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_144 VNB N_A_197_119#_c_2459_n 0.00956105f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_145 VNB N_A_197_119#_c_2460_n 0.00204055f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_146 VNB N_A_197_119#_c_2461_n 0.00353255f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_147 VNB N_A_197_119#_c_2462_n 0.00309253f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_148 VNB N_A_197_119#_c_2463_n 0.0161189f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_149 VNB N_A_197_119#_c_2464_n 0.00281216f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_150 VNB N_A_197_119#_c_2465_n 0.0128672f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_151 VNB N_A_197_119#_c_2466_n 0.00459078f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_152 VNB N_A_197_119#_c_2467_n 2.32436e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_153 VNB N_A_197_119#_c_2468_n 0.00433075f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_154 VNB N_A_197_119#_c_2469_n 0.00285092f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_155 VNB N_Q_N_c_2675_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_156 VNB N_Q_N_c_2676_n 0.00285092f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.97
cc_157 VNB N_Q_N_c_2677_n 0.0012244f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_158 VNB N_Q_c_2705_n 0.00240255f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_159 VNB N_Q_c_2706_n 0.00208476f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.97
cc_160 VNB N_VGND_c_2732_n 0.0130142f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_161 VNB N_VGND_c_2733_n 0.0375162f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_162 VNB N_VGND_c_2734_n 0.0105181f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_163 VNB N_VGND_c_2735_n 0.00706582f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_164 VNB N_VGND_c_2736_n 0.00426387f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_165 VNB N_VGND_c_2737_n 0.00753696f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_166 VNB N_VGND_c_2738_n 0.0682466f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_167 VNB N_VGND_c_2739_n 0.0304662f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_168 VNB N_VGND_c_2740_n 0.0263825f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_169 VNB N_VGND_c_2741_n 0.0135219f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_170 VNB N_VGND_c_2742_n 0.0105185f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_171 VNB N_VGND_c_2743_n 0.050708f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_172 VNB N_VGND_c_2744_n 0.0499949f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_173 VNB N_VGND_c_2745_n 0.00332923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_174 VNB N_VGND_c_2746_n 0.0711334f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_175 VNB N_VGND_c_2747_n 0.00548191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_176 VNB N_VGND_c_2748_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_177 VNB N_VGND_c_2749_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_178 VNB N_VGND_c_2750_n 0.0360368f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_179 VNB N_VGND_c_2751_n 0.0296999f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_180 VNB N_VGND_c_2752_n 0.0801927f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_181 VNB N_VGND_c_2753_n 0.0223582f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_182 VNB N_VGND_c_2754_n 0.0189739f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_183 VNB N_VGND_c_2755_n 0.00477852f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_184 VNB N_VGND_c_2756_n 0.00359556f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_185 VNB N_VGND_c_2757_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_186 VNB N_VGND_c_2758_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_187 VNB N_VGND_c_2759_n 0.906318f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_188 VNB N_A_1473_73#_c_2925_n 0.0202421f $X=-0.19 $Y=-0.245 $X2=0.52
+ $Y2=0.805
cc_189 VNB N_A_1473_73#_c_2926_n 0.00620629f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.58
cc_190 VNB N_A_1473_73#_c_2927_n 0.0120137f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_191 VNB N_A_1473_73#_c_2928_n 0.00262521f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.97
cc_192 VNB N_A_2452_74#_c_2972_n 0.00270494f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.21
cc_193 VNB N_A_2452_74#_c_2973_n 0.0122425f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.29
cc_194 VNB N_A_2452_74#_c_2974_n 0.00237811f $X=-0.19 $Y=-0.245 $X2=0.407
+ $Y2=1.125
cc_195 VPB N_SCD_c_377_n 0.024805f $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.948
cc_196 VPB N_SCD_c_382_n 0.0523285f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.245
cc_197 VPB N_SCD_c_379_n 0.0209687f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.29
cc_198 VPB N_D_c_409_n 0.0144146f $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.312
cc_199 VPB N_D_c_410_n 0.0149255f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.64
cc_200 VPB N_D_c_411_n 0.0169099f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_201 VPB D 0.00263664f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_202 VPB N_D_c_408_n 0.01835f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.97
cc_203 VPB N_A_341_410#_c_470_n 0.0184825f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=0.805
cc_204 VPB N_A_341_410#_c_471_n 0.0220567f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_205 VPB N_A_341_410#_c_472_n 0.0128955f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_206 VPB N_A_341_410#_c_473_n 0.020091f $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.97
cc_207 VPB N_A_341_410#_c_466_n 0.0316015f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.97
cc_208 VPB N_A_341_410#_c_475_n 0.00432096f $X=-0.19 $Y=1.66 $X2=0.337 $Y2=1.29
cc_209 VPB N_A_341_410#_c_468_n 0.0142764f $X=-0.19 $Y=1.66 $X2=0.337 $Y2=1.665
cc_210 VPB N_A_341_410#_c_477_n 0.0188772f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_211 VPB N_SCE_c_558_n 0.0202904f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.125
cc_212 VPB N_SCE_c_559_n 0.0205091f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=0.805
cc_213 VPB N_SCE_c_560_n 0.022135f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_214 VPB N_SCE_c_561_n 0.0345514f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_215 VPB N_SCE_c_562_n 0.015354f $X=-0.19 $Y=1.66 $X2=0.337 $Y2=1.295
cc_216 VPB N_SCE_c_553_n 0.0213015f $X=-0.19 $Y=1.66 $X2=0.337 $Y2=1.665
cc_217 VPB N_SCE_c_555_n 0.0125991f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_218 VPB N_SCE_c_557_n 0.00608076f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_219 VPB N_CLK_N_c_652_n 0.0299485f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.64
cc_220 VPB N_CLK_N_c_653_n 0.00333099f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_221 VPB N_A_1007_366#_c_700_n 0.0561716f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_222 VPB N_A_1007_366#_c_691_n 0.010135f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.29
cc_223 VPB N_A_1007_366#_c_702_n 0.0171426f $X=-0.19 $Y=1.66 $X2=0.337 $Y2=1.665
cc_224 VPB N_A_1007_366#_c_703_n 0.00594041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_225 VPB N_A_1007_366#_c_704_n 0.00385457f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_226 VPB N_A_1007_366#_c_705_n 0.00652179f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_227 VPB N_A_1007_366#_c_706_n 0.00519677f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_228 VPB N_A_1007_366#_c_696_n 0.00336349f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_229 VPB N_A_1007_366#_c_708_n 0.0154267f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_230 VPB N_A_1007_366#_c_698_n 6.31765e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_231 VPB N_A_1007_366#_c_699_n 0.0432422f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_232 VPB N_A_1007_366#_c_711_n 0.0143316f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_233 VPB N_A_1007_366#_c_712_n 0.0216849f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_234 VPB N_A_1007_366#_c_713_n 0.00112972f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_235 VPB N_A_1007_366#_c_714_n 0.00579482f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_236 VPB N_A_1007_366#_c_715_n 0.00885653f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_237 VPB N_A_868_368#_c_905_n 0.0182291f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=0.805
cc_238 VPB N_A_868_368#_c_906_n 0.0216834f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_239 VPB N_A_868_368#_c_907_n 0.0113128f $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.97
cc_240 VPB N_A_868_368#_c_908_n 0.0225614f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.97
cc_241 VPB N_A_868_368#_c_909_n 0.0164697f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_242 VPB N_A_868_368#_c_910_n 0.00453418f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_243 VPB N_A_868_368#_c_894_n 0.00350364f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_244 VPB N_A_868_368#_c_896_n 0.001441f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_245 VPB N_A_868_368#_c_897_n 0.019116f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_246 VPB N_A_868_368#_c_898_n 0.0024891f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_247 VPB N_A_868_368#_c_901_n 0.00185142f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_248 VPB N_A_868_368#_c_902_n 0.0156189f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_249 VPB N_A_868_368#_c_903_n 0.00987632f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_250 VPB N_A_868_368#_c_904_n 0.00564828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_251 VPB N_A_1154_464#_c_1101_n 0.0156057f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_252 VPB N_A_1154_464#_c_1109_n 0.0229156f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_253 VPB N_A_1154_464#_c_1110_n 0.00121847f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_254 VPB N_A_1154_464#_c_1111_n 0.0202408f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_255 VPB N_A_1154_464#_c_1112_n 0.00454222f $X=-0.19 $Y=1.66 $X2=0.337
+ $Y2=1.665
cc_256 VPB N_A_1154_464#_c_1113_n 0.00371793f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_257 VPB N_A_1154_464#_c_1107_n 0.0346499f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_258 VPB N_A_1643_257#_c_1217_n 0.0159492f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=0.805
cc_259 VPB N_A_1643_257#_c_1201_n 0.0068631f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.29
cc_260 VPB N_A_1643_257#_c_1219_n 0.0202174f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.97
cc_261 VPB N_A_1643_257#_c_1203_n 0.0288397f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_262 VPB N_A_1643_257#_c_1209_n 0.00816623f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_263 VPB N_A_1643_257#_c_1211_n 0.00460414f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_264 VPB N_A_1643_257#_c_1223_n 0.00648869f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_265 VPB N_SET_B_c_1415_n 0.0105479f $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.948
cc_266 VPB N_SET_B_c_1416_n 0.0259019f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.245
cc_267 VPB N_SET_B_c_1407_n 0.0069629f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_268 VPB N_SET_B_c_1418_n 0.0239997f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.29
cc_269 VPB N_SET_B_c_1408_n 0.0160556f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.97
cc_270 VPB N_SET_B_c_1420_n 0.00103621f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.97
cc_271 VPB N_SET_B_c_1409_n 0.00137382f $X=-0.19 $Y=1.66 $X2=0.337 $Y2=1.295
cc_272 VPB SET_B 0.00242819f $X=-0.19 $Y=1.66 $X2=0.337 $Y2=1.665
cc_273 VPB N_SET_B_c_1411_n 0.0126394f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_274 VPB N_SET_B_c_1413_n 0.00277883f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_275 VPB N_A_688_98#_c_1560_n 0.0167386f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=0.805
cc_276 VPB N_A_688_98#_M1016_g 0.026271f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.97
cc_277 VPB N_A_688_98#_c_1562_n 0.0065161f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_278 VPB N_A_688_98#_c_1563_n 0.0144457f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_279 VPB N_A_688_98#_c_1564_n 0.0228896f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_280 VPB N_A_688_98#_c_1565_n 0.033276f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_281 VPB N_A_688_98#_c_1555_n 0.0219303f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_282 VPB N_A_688_98#_c_1567_n 0.00206029f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_283 VPB N_A_688_98#_c_1568_n 0.00988356f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_284 VPB N_A_688_98#_c_1569_n 0.00123041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_285 VPB N_A_688_98#_c_1557_n 0.00231451f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_286 VPB N_A_688_98#_c_1558_n 0.0187864f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_287 VPB N_A_2216_410#_c_1742_n 0.0585362f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_288 VPB N_A_2216_410#_c_1743_n 0.0203062f $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.29
cc_289 VPB N_A_2216_410#_c_1728_n 0.0238508f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.97
cc_290 VPB N_A_2216_410#_c_1745_n 0.0166637f $X=-0.19 $Y=1.66 $X2=0.337 $Y2=1.97
cc_291 VPB N_A_2216_410#_c_1746_n 0.0176401f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_292 VPB N_A_2216_410#_c_1733_n 0.0141335f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_293 VPB N_A_2216_410#_c_1735_n 0.0315352f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_294 VPB N_A_2216_410#_c_1749_n 0.0136515f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_295 VPB N_A_2216_410#_c_1750_n 0.00276769f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_296 VPB N_A_2216_410#_c_1751_n 0.0156132f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_297 VPB N_A_2216_410#_c_1752_n 0.00536784f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_298 VPB N_A_2216_410#_c_1753_n 0.00151987f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_299 VPB N_A_2216_410#_c_1754_n 0.00912948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_300 VPB N_A_2216_410#_c_1739_n 0.00593009f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_301 VPB N_A_2216_410#_c_1741_n 0.0167723f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_302 VPB N_A_1997_82#_c_1935_n 0.0405845f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=0.805
cc_303 VPB N_A_1997_82#_c_1942_n 0.00550006f $X=-0.19 $Y=1.66 $X2=0.337 $Y2=1.29
cc_304 VPB N_A_1997_82#_c_1943_n 0.00207661f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_305 VPB N_A_1997_82#_c_1944_n 0.0149965f $X=-0.19 $Y=1.66 $X2=0.337 $Y2=1.665
cc_306 VPB N_A_1997_82#_c_1945_n 4.60744e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_307 VPB N_A_1997_82#_c_1938_n 0.00144126f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_308 VPB N_A_1997_82#_c_1947_n 0.00873063f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_309 VPB N_A_1997_82#_c_1948_n 0.00616851f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_310 VPB N_A_1997_82#_c_1949_n 0.0082052f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_311 VPB N_A_1997_82#_c_1950_n 0.00428128f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_312 VPB N_A_1997_82#_c_1951_n 0.00243246f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_313 VPB N_A_1997_82#_c_1940_n 0.0024738f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_314 VPB N_RESET_B_c_2095_n 0.043597f $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.312
cc_315 VPB RESET_B 0.00276636f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=0.805
cc_316 VPB N_A_3272_94#_c_2133_n 0.0159939f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=0.805
cc_317 VPB N_A_3272_94#_c_2134_n 0.0173548f $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.29
cc_318 VPB N_A_3272_94#_c_2135_n 0.0169933f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_319 VPB N_A_3272_94#_c_2132_n 0.0168827f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_320 VPB N_A_27_464#_c_2193_n 0.0112389f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_321 VPB N_A_27_464#_c_2194_n 0.00669267f $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.29
cc_322 VPB N_A_27_464#_c_2195_n 0.00197776f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.29
cc_323 VPB N_A_27_464#_c_2196_n 0.00740921f $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.97
cc_324 VPB N_A_27_464#_c_2197_n 0.0301618f $X=-0.19 $Y=1.66 $X2=0.337 $Y2=1.29
cc_325 VPB N_VPWR_c_2235_n 0.00396467f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_326 VPB N_VPWR_c_2236_n 0.0166421f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_327 VPB N_VPWR_c_2237_n 0.00396467f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_328 VPB N_VPWR_c_2238_n 0.0210102f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_329 VPB N_VPWR_c_2239_n 0.012173f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_330 VPB N_VPWR_c_2240_n 0.00660284f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_331 VPB N_VPWR_c_2241_n 0.0131965f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_332 VPB N_VPWR_c_2242_n 0.0105447f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_333 VPB N_VPWR_c_2243_n 0.00662307f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_334 VPB N_VPWR_c_2244_n 0.00248226f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_335 VPB N_VPWR_c_2245_n 0.0166714f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_336 VPB N_VPWR_c_2246_n 0.0111387f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_337 VPB N_VPWR_c_2247_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_338 VPB N_VPWR_c_2248_n 0.0637998f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_339 VPB N_VPWR_c_2249_n 0.021877f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_340 VPB N_VPWR_c_2250_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_341 VPB N_VPWR_c_2251_n 0.0210814f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_342 VPB N_VPWR_c_2252_n 0.00615051f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_343 VPB N_VPWR_c_2253_n 0.0186844f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_344 VPB N_VPWR_c_2254_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_345 VPB N_VPWR_c_2255_n 0.0180274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_346 VPB N_VPWR_c_2256_n 0.0373247f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_347 VPB N_VPWR_c_2257_n 0.0317045f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_348 VPB N_VPWR_c_2258_n 0.0753346f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_349 VPB N_VPWR_c_2259_n 0.0427226f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_350 VPB N_VPWR_c_2260_n 0.020899f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_351 VPB N_VPWR_c_2261_n 0.0180566f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_352 VPB N_VPWR_c_2262_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_353 VPB N_VPWR_c_2263_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_354 VPB N_VPWR_c_2264_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_355 VPB N_VPWR_c_2265_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_356 VPB N_VPWR_c_2266_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_357 VPB N_VPWR_c_2267_n 0.00610243f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_358 VPB N_VPWR_c_2268_n 0.0465718f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_359 VPB N_VPWR_c_2269_n 0.0348815f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_360 VPB N_VPWR_c_2270_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_361 VPB N_VPWR_c_2234_n 0.232659f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_362 VPB N_A_197_119#_c_2470_n 7.96979e-19 $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.29
cc_363 VPB N_A_197_119#_c_2471_n 0.00521557f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_364 VPB N_A_197_119#_c_2472_n 9.80635e-19 $X=-0.19 $Y=1.66 $X2=0.337
+ $Y2=1.665
cc_365 VPB N_A_197_119#_c_2449_n 0.0029261f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_366 VPB N_A_197_119#_c_2474_n 0.00630366f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_367 VPB N_A_197_119#_c_2468_n 0.00855178f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_368 VPB N_A_197_119#_c_2476_n 0.00256186f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_369 VPB N_A_197_119#_c_2477_n 0.00743479f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_370 VPB N_Q_N_c_2678_n 0.00273338f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.29
cc_371 VPB Q_N 0.00232002f $X=-0.19 $Y=1.66 $X2=0.337 $Y2=1.29
cc_372 VPB Q 0.00382657f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.29
cc_373 VPB Q 0.0024312f $X=-0.19 $Y=1.66 $X2=0.337 $Y2=1.29
cc_374 VPB N_Q_c_2706_n 0.00104928f $X=-0.19 $Y=1.66 $X2=0.337 $Y2=1.97
cc_375 N_SCD_c_380_n N_SCE_M1032_g 0.0344188f $X=0.407 $Y=1.125 $X2=0 $Y2=0
cc_376 N_SCD_c_377_n N_SCE_c_558_n 0.0116048f $X=0.407 $Y=1.948 $X2=0 $Y2=0
cc_377 N_SCD_c_379_n N_SCE_c_558_n 0.00197263f $X=0.385 $Y=1.29 $X2=0 $Y2=0
cc_378 N_SCD_c_382_n N_SCE_c_559_n 0.0322044f $X=0.505 $Y=2.245 $X2=0 $Y2=0
cc_379 N_SCD_c_377_n N_SCE_c_554_n 0.0207335f $X=0.407 $Y=1.948 $X2=0 $Y2=0
cc_380 N_SCD_c_378_n N_SCE_c_556_n 0.0207335f $X=0.385 $Y=1.29 $X2=0 $Y2=0
cc_381 N_SCD_c_379_n N_SCE_c_556_n 0.00217323f $X=0.385 $Y=1.29 $X2=0 $Y2=0
cc_382 N_SCD_c_378_n N_SCE_c_557_n 0.00246198f $X=0.385 $Y=1.29 $X2=0 $Y2=0
cc_383 N_SCD_c_379_n N_SCE_c_557_n 0.0382498f $X=0.385 $Y=1.29 $X2=0 $Y2=0
cc_384 N_SCD_c_382_n N_A_27_464#_c_2193_n 0.0125458f $X=0.505 $Y=2.245 $X2=0
+ $Y2=0
cc_385 N_SCD_c_379_n N_A_27_464#_c_2193_n 0.0142215f $X=0.385 $Y=1.29 $X2=0
+ $Y2=0
cc_386 N_SCD_c_382_n N_A_27_464#_c_2197_n 0.00625229f $X=0.505 $Y=2.245 $X2=0
+ $Y2=0
cc_387 N_SCD_c_379_n N_A_27_464#_c_2197_n 0.0217226f $X=0.385 $Y=1.29 $X2=0
+ $Y2=0
cc_388 N_SCD_c_382_n N_VPWR_c_2235_n 0.010249f $X=0.505 $Y=2.245 $X2=0 $Y2=0
cc_389 N_SCD_c_382_n N_VPWR_c_2255_n 0.00413917f $X=0.505 $Y=2.245 $X2=0 $Y2=0
cc_390 N_SCD_c_382_n N_VPWR_c_2234_n 0.00421383f $X=0.505 $Y=2.245 $X2=0 $Y2=0
cc_391 N_SCD_c_380_n N_A_197_119#_c_2478_n 9.24658e-19 $X=0.407 $Y=1.125 $X2=0
+ $Y2=0
cc_392 N_SCD_c_378_n N_VGND_c_2733_n 0.00158682f $X=0.385 $Y=1.29 $X2=0 $Y2=0
cc_393 N_SCD_c_379_n N_VGND_c_2733_n 0.0263818f $X=0.385 $Y=1.29 $X2=0 $Y2=0
cc_394 N_SCD_c_380_n N_VGND_c_2733_n 0.0117834f $X=0.407 $Y=1.125 $X2=0 $Y2=0
cc_395 N_SCD_c_380_n N_VGND_c_2744_n 0.0035863f $X=0.407 $Y=1.125 $X2=0 $Y2=0
cc_396 N_SCD_c_380_n N_VGND_c_2759_n 0.00401353f $X=0.407 $Y=1.125 $X2=0 $Y2=0
cc_397 N_D_c_409_n N_A_341_410#_c_470_n 0.0175254f $X=1.345 $Y=2.245 $X2=0 $Y2=0
cc_398 N_D_c_411_n N_A_341_410#_c_472_n 0.0110128f $X=1.345 $Y=2.14 $X2=0 $Y2=0
cc_399 N_D_c_408_n N_A_341_410#_c_472_n 0.00552732f $X=1.74 $Y=1.625 $X2=0 $Y2=0
cc_400 N_D_M1042_g N_A_341_410#_M1025_g 0.0344383f $X=1.74 $Y=0.805 $X2=0 $Y2=0
cc_401 D N_A_341_410#_M1025_g 3.65577e-19 $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_402 N_D_c_411_n N_A_341_410#_c_473_n 0.00201894f $X=1.345 $Y=2.14 $X2=0 $Y2=0
cc_403 N_D_c_410_n N_A_341_410#_c_475_n 0.00201894f $X=1.42 $Y=2.035 $X2=0 $Y2=0
cc_404 N_D_c_408_n N_A_341_410#_c_475_n 0.0344383f $X=1.74 $Y=1.625 $X2=0 $Y2=0
cc_405 N_D_M1042_g N_SCE_M1032_g 0.00443391f $X=1.74 $Y=0.805 $X2=0 $Y2=0
cc_406 N_D_c_410_n N_SCE_c_558_n 0.011174f $X=1.42 $Y=2.035 $X2=0 $Y2=0
cc_407 N_D_c_411_n N_SCE_c_558_n 0.0136488f $X=1.345 $Y=2.14 $X2=0 $Y2=0
cc_408 N_D_c_409_n N_SCE_c_559_n 0.039278f $X=1.345 $Y=2.245 $X2=0 $Y2=0
cc_409 N_D_M1042_g N_SCE_c_548_n 0.0103083f $X=1.74 $Y=0.805 $X2=0 $Y2=0
cc_410 D N_SCE_c_554_n 2.39818e-19 $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_411 N_D_c_408_n N_SCE_c_554_n 0.010556f $X=1.74 $Y=1.625 $X2=0 $Y2=0
cc_412 N_D_c_410_n N_SCE_c_555_n 0.010556f $X=1.42 $Y=2.035 $X2=0 $Y2=0
cc_413 N_D_M1042_g N_SCE_c_556_n 0.00564298f $X=1.74 $Y=0.805 $X2=0 $Y2=0
cc_414 N_D_M1042_g N_SCE_c_557_n 0.00231918f $X=1.74 $Y=0.805 $X2=0 $Y2=0
cc_415 N_D_c_411_n N_SCE_c_557_n 0.0025439f $X=1.345 $Y=2.14 $X2=0 $Y2=0
cc_416 D N_SCE_c_557_n 0.0270453f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_417 N_D_c_408_n N_SCE_c_557_n 0.00278654f $X=1.74 $Y=1.625 $X2=0 $Y2=0
cc_418 N_D_c_409_n N_A_27_464#_c_2193_n 7.08327e-19 $X=1.345 $Y=2.245 $X2=0
+ $Y2=0
cc_419 N_D_c_409_n N_A_27_464#_c_2194_n 0.0126939f $X=1.345 $Y=2.245 $X2=0 $Y2=0
cc_420 N_D_c_409_n N_A_27_464#_c_2196_n 6.63009e-19 $X=1.345 $Y=2.245 $X2=0
+ $Y2=0
cc_421 N_D_c_409_n N_VPWR_c_2235_n 2.96128e-19 $X=1.345 $Y=2.245 $X2=0 $Y2=0
cc_422 N_D_c_409_n N_VPWR_c_2256_n 0.00278271f $X=1.345 $Y=2.245 $X2=0 $Y2=0
cc_423 N_D_c_409_n N_VPWR_c_2234_n 0.00353419f $X=1.345 $Y=2.245 $X2=0 $Y2=0
cc_424 N_D_c_409_n N_A_197_119#_c_2470_n 0.00206961f $X=1.345 $Y=2.245 $X2=0
+ $Y2=0
cc_425 N_D_c_411_n N_A_197_119#_c_2470_n 0.0032068f $X=1.345 $Y=2.14 $X2=0 $Y2=0
cc_426 N_D_c_409_n N_A_197_119#_c_2481_n 0.0033192f $X=1.345 $Y=2.245 $X2=0
+ $Y2=0
cc_427 N_D_M1042_g N_A_197_119#_c_2482_n 0.00586537f $X=1.74 $Y=0.805 $X2=0
+ $Y2=0
cc_428 N_D_M1042_g N_A_197_119#_c_2446_n 0.00470158f $X=1.74 $Y=0.805 $X2=0
+ $Y2=0
cc_429 D N_A_197_119#_c_2471_n 0.011971f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_430 N_D_c_408_n N_A_197_119#_c_2471_n 6.80579e-19 $X=1.74 $Y=1.625 $X2=0
+ $Y2=0
cc_431 N_D_c_410_n N_A_197_119#_c_2472_n 0.00292224f $X=1.42 $Y=2.035 $X2=0
+ $Y2=0
cc_432 N_D_c_411_n N_A_197_119#_c_2472_n 0.00285853f $X=1.345 $Y=2.14 $X2=0
+ $Y2=0
cc_433 D N_A_197_119#_c_2472_n 0.0142813f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_434 N_D_c_408_n N_A_197_119#_c_2472_n 0.00126636f $X=1.74 $Y=1.625 $X2=0
+ $Y2=0
cc_435 N_D_M1042_g N_A_197_119#_c_2447_n 0.0106578f $X=1.74 $Y=0.805 $X2=0 $Y2=0
cc_436 D N_A_197_119#_c_2447_n 0.00886748f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_437 N_D_M1042_g N_A_197_119#_c_2448_n 0.00292725f $X=1.74 $Y=0.805 $X2=0
+ $Y2=0
cc_438 D N_A_197_119#_c_2448_n 0.0171437f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_439 N_D_c_408_n N_A_197_119#_c_2448_n 0.00140614f $X=1.74 $Y=1.625 $X2=0
+ $Y2=0
cc_440 N_D_c_410_n N_A_197_119#_c_2449_n 0.00263471f $X=1.42 $Y=2.035 $X2=0
+ $Y2=0
cc_441 N_D_M1042_g N_A_197_119#_c_2449_n 0.00366275f $X=1.74 $Y=0.805 $X2=0
+ $Y2=0
cc_442 D N_A_197_119#_c_2449_n 0.0248017f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_443 N_D_c_409_n N_A_197_119#_c_2476_n 0.00128638f $X=1.345 $Y=2.245 $X2=0
+ $Y2=0
cc_444 N_D_c_411_n N_A_197_119#_c_2476_n 0.00286955f $X=1.345 $Y=2.14 $X2=0
+ $Y2=0
cc_445 N_D_c_408_n N_A_197_119#_c_2478_n 0.00435793f $X=1.74 $Y=1.625 $X2=0
+ $Y2=0
cc_446 N_D_M1042_g N_VGND_c_2734_n 0.00171774f $X=1.74 $Y=0.805 $X2=0 $Y2=0
cc_447 N_D_M1042_g N_VGND_c_2759_n 9.39239e-19 $X=1.74 $Y=0.805 $X2=0 $Y2=0
cc_448 N_A_341_410#_M1025_g N_SCE_c_548_n 0.0103107f $X=2.13 $Y=0.805 $X2=0
+ $Y2=0
cc_449 N_A_341_410#_c_477_n N_SCE_c_560_n 0.0052938f $X=3.03 $Y=2.465 $X2=0
+ $Y2=0
cc_450 N_A_341_410#_M1025_g N_SCE_M1037_g 0.0102025f $X=2.13 $Y=0.805 $X2=0
+ $Y2=0
cc_451 N_A_341_410#_c_469_n N_SCE_M1037_g 0.00221787f $X=3.025 $Y=0.815 $X2=0
+ $Y2=0
cc_452 N_A_341_410#_c_469_n N_SCE_c_551_n 0.0189146f $X=3.025 $Y=0.815 $X2=0
+ $Y2=0
cc_453 N_A_341_410#_c_467_n N_SCE_c_552_n 0.00123218f $X=2.94 $Y=1.645 $X2=0
+ $Y2=0
cc_454 N_A_341_410#_c_468_n N_SCE_c_552_n 0.0117621f $X=2.77 $Y=1.645 $X2=0
+ $Y2=0
cc_455 N_A_341_410#_c_477_n N_SCE_c_561_n 0.0225628f $X=3.03 $Y=2.465 $X2=0
+ $Y2=0
cc_456 N_A_341_410#_c_471_n N_SCE_c_562_n 0.00485861f $X=2.055 $Y=2.125 $X2=0
+ $Y2=0
cc_457 N_A_341_410#_c_467_n N_SCE_c_562_n 0.00151184f $X=2.94 $Y=1.645 $X2=0
+ $Y2=0
cc_458 N_A_341_410#_c_468_n N_SCE_c_562_n 0.0130968f $X=2.77 $Y=1.645 $X2=0
+ $Y2=0
cc_459 N_A_341_410#_c_477_n N_SCE_c_562_n 0.00187562f $X=3.03 $Y=2.465 $X2=0
+ $Y2=0
cc_460 N_A_341_410#_c_468_n N_SCE_c_553_n 0.0181259f $X=2.77 $Y=1.645 $X2=0
+ $Y2=0
cc_461 N_A_341_410#_c_469_n N_SCE_c_553_n 0.00654003f $X=3.025 $Y=0.815 $X2=0
+ $Y2=0
cc_462 N_A_341_410#_c_477_n N_SCE_c_553_n 0.00664705f $X=3.03 $Y=2.465 $X2=0
+ $Y2=0
cc_463 N_A_341_410#_c_501_p N_SCE_c_553_n 0.00776514f $X=3.067 $Y=1.645 $X2=0
+ $Y2=0
cc_464 N_A_341_410#_c_469_n N_CLK_N_c_651_n 0.00429407f $X=3.025 $Y=0.815
+ $X2=-0.19 $Y2=-0.245
cc_465 N_A_341_410#_c_477_n N_CLK_N_c_652_n 5.62636e-19 $X=3.03 $Y=2.465 $X2=0
+ $Y2=0
cc_466 N_A_341_410#_c_501_p N_CLK_N_c_652_n 3.99371e-19 $X=3.067 $Y=1.645 $X2=0
+ $Y2=0
cc_467 N_A_341_410#_c_469_n N_CLK_N_c_653_n 0.00689029f $X=3.025 $Y=0.815 $X2=0
+ $Y2=0
cc_468 N_A_341_410#_c_501_p N_CLK_N_c_653_n 0.0169701f $X=3.067 $Y=1.645 $X2=0
+ $Y2=0
cc_469 N_A_341_410#_c_469_n N_A_688_98#_c_1556_n 0.0116565f $X=3.025 $Y=0.815
+ $X2=0 $Y2=0
cc_470 N_A_341_410#_c_477_n N_A_688_98#_c_1567_n 0.0111955f $X=3.03 $Y=2.465
+ $X2=0 $Y2=0
cc_471 N_A_341_410#_c_477_n N_A_688_98#_c_1568_n 0.0552314f $X=3.03 $Y=2.465
+ $X2=0 $Y2=0
cc_472 N_A_341_410#_c_470_n N_A_27_464#_c_2194_n 0.0134197f $X=1.795 $Y=2.245
+ $X2=0 $Y2=0
cc_473 N_A_341_410#_c_470_n N_A_27_464#_c_2196_n 0.00809535f $X=1.795 $Y=2.245
+ $X2=0 $Y2=0
cc_474 N_A_341_410#_c_471_n N_A_27_464#_c_2196_n 0.00813623f $X=2.055 $Y=2.125
+ $X2=0 $Y2=0
cc_475 N_A_341_410#_c_472_n N_A_27_464#_c_2196_n 3.63282e-19 $X=1.885 $Y=2.125
+ $X2=0 $Y2=0
cc_476 N_A_341_410#_c_470_n N_VPWR_c_2236_n 0.00193603f $X=1.795 $Y=2.245 $X2=0
+ $Y2=0
cc_477 N_A_341_410#_c_466_n N_VPWR_c_2236_n 0.00764644f $X=2.605 $Y=1.735 $X2=0
+ $Y2=0
cc_478 N_A_341_410#_c_467_n N_VPWR_c_2236_n 0.00524534f $X=2.94 $Y=1.645 $X2=0
+ $Y2=0
cc_479 N_A_341_410#_c_477_n N_VPWR_c_2236_n 0.0456538f $X=3.03 $Y=2.465 $X2=0
+ $Y2=0
cc_480 N_A_341_410#_c_470_n N_VPWR_c_2256_n 0.00278257f $X=1.795 $Y=2.245 $X2=0
+ $Y2=0
cc_481 N_A_341_410#_c_477_n N_VPWR_c_2257_n 0.011066f $X=3.03 $Y=2.465 $X2=0
+ $Y2=0
cc_482 N_A_341_410#_c_470_n N_VPWR_c_2234_n 0.00358707f $X=1.795 $Y=2.245 $X2=0
+ $Y2=0
cc_483 N_A_341_410#_c_477_n N_VPWR_c_2234_n 0.00915947f $X=3.03 $Y=2.465 $X2=0
+ $Y2=0
cc_484 N_A_341_410#_M1025_g N_A_197_119#_c_2482_n 9.40746e-19 $X=2.13 $Y=0.805
+ $X2=0 $Y2=0
cc_485 N_A_341_410#_M1025_g N_A_197_119#_c_2446_n 8.17804e-19 $X=2.13 $Y=0.805
+ $X2=0 $Y2=0
cc_486 N_A_341_410#_c_471_n N_A_197_119#_c_2471_n 0.00864033f $X=2.055 $Y=2.125
+ $X2=0 $Y2=0
cc_487 N_A_341_410#_c_472_n N_A_197_119#_c_2471_n 0.0106564f $X=1.885 $Y=2.125
+ $X2=0 $Y2=0
cc_488 N_A_341_410#_c_473_n N_A_197_119#_c_2471_n 0.00638474f $X=2.13 $Y=2.05
+ $X2=0 $Y2=0
cc_489 N_A_341_410#_M1025_g N_A_197_119#_c_2449_n 0.0142097f $X=2.13 $Y=0.805
+ $X2=0 $Y2=0
cc_490 N_A_341_410#_c_473_n N_A_197_119#_c_2449_n 0.00838483f $X=2.13 $Y=2.05
+ $X2=0 $Y2=0
cc_491 N_A_341_410#_c_475_n N_A_197_119#_c_2449_n 0.0056277f $X=2.13 $Y=1.735
+ $X2=0 $Y2=0
cc_492 N_A_341_410#_c_467_n N_A_197_119#_c_2449_n 0.0111722f $X=2.94 $Y=1.645
+ $X2=0 $Y2=0
cc_493 N_A_341_410#_c_468_n N_A_197_119#_c_2449_n 2.07375e-19 $X=2.77 $Y=1.645
+ $X2=0 $Y2=0
cc_494 N_A_341_410#_M1025_g N_A_197_119#_c_2450_n 0.00762767f $X=2.13 $Y=0.805
+ $X2=0 $Y2=0
cc_495 N_A_341_410#_c_466_n N_A_197_119#_c_2450_n 0.0110613f $X=2.605 $Y=1.735
+ $X2=0 $Y2=0
cc_496 N_A_341_410#_c_467_n N_A_197_119#_c_2450_n 0.0127989f $X=2.94 $Y=1.645
+ $X2=0 $Y2=0
cc_497 N_A_341_410#_c_468_n N_A_197_119#_c_2450_n 0.00322911f $X=2.77 $Y=1.645
+ $X2=0 $Y2=0
cc_498 N_A_341_410#_c_469_n N_A_197_119#_c_2450_n 0.0137468f $X=3.025 $Y=0.815
+ $X2=0 $Y2=0
cc_499 N_A_341_410#_M1025_g N_A_197_119#_c_2451_n 0.00374668f $X=2.13 $Y=0.805
+ $X2=0 $Y2=0
cc_500 N_A_341_410#_c_469_n N_A_197_119#_c_2451_n 0.0217676f $X=3.025 $Y=0.815
+ $X2=0 $Y2=0
cc_501 N_A_341_410#_c_469_n N_A_197_119#_c_2452_n 0.0195912f $X=3.025 $Y=0.815
+ $X2=0 $Y2=0
cc_502 N_A_341_410#_c_469_n N_A_197_119#_c_2454_n 0.00501222f $X=3.025 $Y=0.815
+ $X2=0 $Y2=0
cc_503 N_A_341_410#_c_469_n N_A_197_119#_c_2455_n 0.0147661f $X=3.025 $Y=0.815
+ $X2=0 $Y2=0
cc_504 N_A_341_410#_c_470_n N_A_197_119#_c_2476_n 0.00297969f $X=1.795 $Y=2.245
+ $X2=0 $Y2=0
cc_505 N_A_341_410#_c_472_n N_A_197_119#_c_2476_n 0.00276562f $X=1.885 $Y=2.125
+ $X2=0 $Y2=0
cc_506 N_A_341_410#_M1025_g N_A_197_119#_c_2469_n 0.00832057f $X=2.13 $Y=0.805
+ $X2=0 $Y2=0
cc_507 N_A_341_410#_M1025_g N_VGND_c_2734_n 0.0104567f $X=2.13 $Y=0.805 $X2=0
+ $Y2=0
cc_508 N_A_341_410#_M1025_g N_VGND_c_2759_n 7.88961e-19 $X=2.13 $Y=0.805 $X2=0
+ $Y2=0
cc_509 N_SCE_c_551_n N_CLK_N_c_651_n 0.00663801f $X=3.175 $Y=1.165 $X2=-0.19
+ $Y2=-0.245
cc_510 N_SCE_c_553_n N_CLK_N_c_652_n 0.0266707f $X=3.25 $Y=2.05 $X2=0 $Y2=0
cc_511 N_SCE_c_553_n N_CLK_N_c_653_n 0.0033514f $X=3.25 $Y=2.05 $X2=0 $Y2=0
cc_512 N_SCE_c_551_n N_A_688_98#_c_1556_n 9.33152e-19 $X=3.175 $Y=1.165 $X2=0
+ $Y2=0
cc_513 N_SCE_c_553_n N_A_688_98#_c_1567_n 0.00204886f $X=3.25 $Y=2.05 $X2=0
+ $Y2=0
cc_514 N_SCE_c_561_n N_A_688_98#_c_1568_n 8.81041e-19 $X=3.175 $Y=2.125 $X2=0
+ $Y2=0
cc_515 N_SCE_c_559_n N_A_27_464#_c_2193_n 0.0138987f $X=0.955 $Y=2.245 $X2=0
+ $Y2=0
cc_516 N_SCE_c_555_n N_A_27_464#_c_2193_n 8.83169e-19 $X=0.97 $Y=1.795 $X2=0
+ $Y2=0
cc_517 N_SCE_c_557_n N_A_27_464#_c_2193_n 0.0154717f $X=0.97 $Y=1.29 $X2=0 $Y2=0
cc_518 N_SCE_c_560_n N_A_27_464#_c_2194_n 5.94256e-19 $X=2.805 $Y=2.245 $X2=0
+ $Y2=0
cc_519 N_SCE_c_559_n N_A_27_464#_c_2195_n 0.00111115f $X=0.955 $Y=2.245 $X2=0
+ $Y2=0
cc_520 N_SCE_c_560_n N_A_27_464#_c_2196_n 0.00107404f $X=2.805 $Y=2.245 $X2=0
+ $Y2=0
cc_521 N_SCE_c_559_n N_VPWR_c_2235_n 0.00635214f $X=0.955 $Y=2.245 $X2=0 $Y2=0
cc_522 N_SCE_c_560_n N_VPWR_c_2236_n 0.0154281f $X=2.805 $Y=2.245 $X2=0 $Y2=0
cc_523 N_SCE_c_562_n N_VPWR_c_2236_n 4.50637e-19 $X=2.895 $Y=2.125 $X2=0 $Y2=0
cc_524 N_SCE_c_559_n N_VPWR_c_2256_n 0.00413917f $X=0.955 $Y=2.245 $X2=0 $Y2=0
cc_525 N_SCE_c_560_n N_VPWR_c_2257_n 0.00413917f $X=2.805 $Y=2.245 $X2=0 $Y2=0
cc_526 N_SCE_c_559_n N_VPWR_c_2234_n 0.00417401f $X=0.955 $Y=2.245 $X2=0 $Y2=0
cc_527 N_SCE_c_560_n N_VPWR_c_2234_n 0.00822528f $X=2.805 $Y=2.245 $X2=0 $Y2=0
cc_528 N_SCE_c_548_n N_A_197_119#_c_2482_n 0.00323516f $X=2.735 $Y=0.18 $X2=0
+ $Y2=0
cc_529 N_SCE_M1032_g N_A_197_119#_c_2446_n 0.00262466f $X=0.91 $Y=0.805 $X2=0
+ $Y2=0
cc_530 N_SCE_c_562_n N_A_197_119#_c_2471_n 4.74987e-19 $X=2.895 $Y=2.125 $X2=0
+ $Y2=0
cc_531 N_SCE_c_558_n N_A_197_119#_c_2472_n 7.46448e-19 $X=0.955 $Y=2.155 $X2=0
+ $Y2=0
cc_532 N_SCE_c_556_n N_A_197_119#_c_2448_n 5.06463e-19 $X=0.97 $Y=1.29 $X2=0
+ $Y2=0
cc_533 N_SCE_c_557_n N_A_197_119#_c_2448_n 0.0150638f $X=0.97 $Y=1.29 $X2=0
+ $Y2=0
cc_534 N_SCE_c_557_n N_A_197_119#_c_2449_n 0.00543475f $X=0.97 $Y=1.29 $X2=0
+ $Y2=0
cc_535 N_SCE_c_552_n N_A_197_119#_c_2450_n 0.00448737f $X=2.885 $Y=1.165 $X2=0
+ $Y2=0
cc_536 N_SCE_M1037_g N_A_197_119#_c_2451_n 0.0172045f $X=2.81 $Y=0.805 $X2=0
+ $Y2=0
cc_537 N_SCE_c_552_n N_A_197_119#_c_2451_n 8.26088e-19 $X=2.885 $Y=1.165 $X2=0
+ $Y2=0
cc_538 N_SCE_M1037_g N_A_197_119#_c_2452_n 0.0117849f $X=2.81 $Y=0.805 $X2=0
+ $Y2=0
cc_539 N_SCE_c_551_n N_A_197_119#_c_2452_n 0.00507912f $X=3.175 $Y=1.165 $X2=0
+ $Y2=0
cc_540 N_SCE_c_548_n N_A_197_119#_c_2453_n 0.0025317f $X=2.735 $Y=0.18 $X2=0
+ $Y2=0
cc_541 N_SCE_M1037_g N_A_197_119#_c_2453_n 0.00343628f $X=2.81 $Y=0.805 $X2=0
+ $Y2=0
cc_542 N_SCE_M1037_g N_A_197_119#_c_2454_n 0.00279325f $X=2.81 $Y=0.805 $X2=0
+ $Y2=0
cc_543 N_SCE_c_558_n N_A_197_119#_c_2476_n 2.27132e-19 $X=0.955 $Y=2.155 $X2=0
+ $Y2=0
cc_544 N_SCE_M1032_g N_A_197_119#_c_2478_n 0.00633316f $X=0.91 $Y=0.805 $X2=0
+ $Y2=0
cc_545 N_SCE_c_548_n N_A_197_119#_c_2478_n 0.00760631f $X=2.735 $Y=0.18 $X2=0
+ $Y2=0
cc_546 N_SCE_c_556_n N_A_197_119#_c_2478_n 9.53161e-19 $X=0.97 $Y=1.29 $X2=0
+ $Y2=0
cc_547 N_SCE_c_557_n N_A_197_119#_c_2478_n 0.0275487f $X=0.97 $Y=1.29 $X2=0
+ $Y2=0
cc_548 N_SCE_M1032_g N_VGND_c_2733_n 0.00173097f $X=0.91 $Y=0.805 $X2=0 $Y2=0
cc_549 N_SCE_c_549_n N_VGND_c_2733_n 0.00977077f $X=0.985 $Y=0.18 $X2=0 $Y2=0
cc_550 N_SCE_c_548_n N_VGND_c_2734_n 0.0209847f $X=2.735 $Y=0.18 $X2=0 $Y2=0
cc_551 N_SCE_M1037_g N_VGND_c_2734_n 0.0025199f $X=2.81 $Y=0.805 $X2=0 $Y2=0
cc_552 N_SCE_c_549_n N_VGND_c_2744_n 0.0404572f $X=0.985 $Y=0.18 $X2=0 $Y2=0
cc_553 N_SCE_c_548_n N_VGND_c_2750_n 0.0125913f $X=2.735 $Y=0.18 $X2=0 $Y2=0
cc_554 N_SCE_c_548_n N_VGND_c_2759_n 0.0582401f $X=2.735 $Y=0.18 $X2=0 $Y2=0
cc_555 N_SCE_c_549_n N_VGND_c_2759_n 0.010774f $X=0.985 $Y=0.18 $X2=0 $Y2=0
cc_556 N_CLK_N_c_652_n N_A_688_98#_c_1560_n 0.0235133f $X=3.815 $Y=1.765 $X2=0
+ $Y2=0
cc_557 N_CLK_N_c_651_n N_A_688_98#_M1043_g 0.0113528f $X=3.8 $Y=1.35 $X2=0 $Y2=0
cc_558 N_CLK_N_c_651_n N_A_688_98#_c_1556_n 0.00945736f $X=3.8 $Y=1.35 $X2=0
+ $Y2=0
cc_559 N_CLK_N_c_652_n N_A_688_98#_c_1556_n 9.85402e-19 $X=3.815 $Y=1.765 $X2=0
+ $Y2=0
cc_560 N_CLK_N_c_653_n N_A_688_98#_c_1556_n 0.026852f $X=3.73 $Y=1.515 $X2=0
+ $Y2=0
cc_561 N_CLK_N_c_652_n N_A_688_98#_c_1567_n 6.76544e-19 $X=3.815 $Y=1.765 $X2=0
+ $Y2=0
cc_562 N_CLK_N_c_653_n N_A_688_98#_c_1567_n 0.016785f $X=3.73 $Y=1.515 $X2=0
+ $Y2=0
cc_563 N_CLK_N_c_652_n N_A_688_98#_c_1568_n 0.00634858f $X=3.815 $Y=1.765 $X2=0
+ $Y2=0
cc_564 N_CLK_N_c_652_n N_A_688_98#_c_1586_n 0.012823f $X=3.815 $Y=1.765 $X2=0
+ $Y2=0
cc_565 N_CLK_N_c_653_n N_A_688_98#_c_1586_n 0.0142266f $X=3.73 $Y=1.515 $X2=0
+ $Y2=0
cc_566 N_CLK_N_c_652_n N_A_688_98#_c_1569_n 0.00355938f $X=3.815 $Y=1.765 $X2=0
+ $Y2=0
cc_567 N_CLK_N_c_652_n N_A_688_98#_c_1557_n 0.002416f $X=3.815 $Y=1.765 $X2=0
+ $Y2=0
cc_568 N_CLK_N_c_653_n N_A_688_98#_c_1557_n 0.0344492f $X=3.73 $Y=1.515 $X2=0
+ $Y2=0
cc_569 N_CLK_N_c_651_n N_A_688_98#_c_1558_n 4.794e-19 $X=3.8 $Y=1.35 $X2=0 $Y2=0
cc_570 N_CLK_N_c_652_n N_A_688_98#_c_1558_n 0.0241918f $X=3.815 $Y=1.765 $X2=0
+ $Y2=0
cc_571 N_CLK_N_c_653_n N_A_688_98#_c_1558_n 4.52373e-19 $X=3.73 $Y=1.515 $X2=0
+ $Y2=0
cc_572 N_CLK_N_c_651_n N_A_688_98#_c_1559_n 0.00424047f $X=3.8 $Y=1.35 $X2=0
+ $Y2=0
cc_573 N_CLK_N_c_652_n N_VPWR_c_2237_n 0.0140627f $X=3.815 $Y=1.765 $X2=0 $Y2=0
cc_574 N_CLK_N_c_652_n N_VPWR_c_2257_n 0.00413917f $X=3.815 $Y=1.765 $X2=0 $Y2=0
cc_575 N_CLK_N_c_652_n N_VPWR_c_2234_n 0.00822528f $X=3.815 $Y=1.765 $X2=0 $Y2=0
cc_576 N_CLK_N_c_651_n N_A_197_119#_c_2452_n 0.00148145f $X=3.8 $Y=1.35 $X2=0
+ $Y2=0
cc_577 N_CLK_N_c_651_n N_A_197_119#_c_2454_n 0.00704041f $X=3.8 $Y=1.35 $X2=0
+ $Y2=0
cc_578 N_CLK_N_c_651_n N_A_197_119#_c_2546_n 0.0144737f $X=3.8 $Y=1.35 $X2=0
+ $Y2=0
cc_579 N_CLK_N_c_651_n N_A_197_119#_c_2456_n 0.00291863f $X=3.8 $Y=1.35 $X2=0
+ $Y2=0
cc_580 N_CLK_N_c_651_n N_VGND_c_2735_n 0.00196633f $X=3.8 $Y=1.35 $X2=0 $Y2=0
cc_581 N_CLK_N_c_651_n N_VGND_c_2750_n 0.0038134f $X=3.8 $Y=1.35 $X2=0 $Y2=0
cc_582 N_CLK_N_c_651_n N_VGND_c_2759_n 0.00508379f $X=3.8 $Y=1.35 $X2=0 $Y2=0
cc_583 N_A_1007_366#_c_700_n N_A_868_368#_c_905_n 0.0199979f $X=5.275 $Y=2.245
+ $X2=0 $Y2=0
cc_584 N_A_1007_366#_c_711_n N_A_868_368#_c_905_n 0.00334717f $X=5.2 $Y=1.995
+ $X2=0 $Y2=0
cc_585 N_A_1007_366#_c_700_n N_A_868_368#_c_906_n 0.0229609f $X=5.275 $Y=2.245
+ $X2=0 $Y2=0
cc_586 N_A_1007_366#_c_703_n N_A_868_368#_c_906_n 0.00777057f $X=5.47 $Y=2.905
+ $X2=0 $Y2=0
cc_587 N_A_1007_366#_c_712_n N_A_868_368#_c_906_n 0.00796635f $X=6.9 $Y=2.902
+ $X2=0 $Y2=0
cc_588 N_A_1007_366#_c_708_n N_A_868_368#_c_907_n 6.34296e-19 $X=9.615 $Y=2.035
+ $X2=0 $Y2=0
cc_589 N_A_1007_366#_c_702_n N_A_868_368#_c_908_n 0.0523069f $X=9.855 $Y=2.045
+ $X2=0 $Y2=0
cc_590 N_A_1007_366#_c_708_n N_A_868_368#_c_908_n 0.00156841f $X=9.615 $Y=2.035
+ $X2=0 $Y2=0
cc_591 N_A_1007_366#_c_700_n N_A_868_368#_c_909_n 0.00452937f $X=5.275 $Y=2.245
+ $X2=0 $Y2=0
cc_592 N_A_1007_366#_c_703_n N_A_868_368#_c_909_n 0.0051238f $X=5.47 $Y=2.905
+ $X2=0 $Y2=0
cc_593 N_A_1007_366#_c_693_n N_A_868_368#_c_929_n 0.00139903f $X=5.355 $Y=1.195
+ $X2=0 $Y2=0
cc_594 N_A_1007_366#_c_700_n N_A_868_368#_c_891_n 9.75528e-19 $X=5.275 $Y=2.245
+ $X2=0 $Y2=0
cc_595 N_A_1007_366#_c_691_n N_A_868_368#_c_891_n 0.00757693f $X=5.28 $Y=1.83
+ $X2=0 $Y2=0
cc_596 N_A_1007_366#_c_692_n N_A_868_368#_c_891_n 0.00758806f $X=5.775 $Y=1.195
+ $X2=0 $Y2=0
cc_597 N_A_1007_366#_c_693_n N_A_868_368#_c_891_n 0.00384428f $X=5.355 $Y=1.195
+ $X2=0 $Y2=0
cc_598 N_A_1007_366#_c_711_n N_A_868_368#_c_891_n 0.017023f $X=5.2 $Y=1.995
+ $X2=0 $Y2=0
cc_599 N_A_1007_366#_c_700_n N_A_868_368#_c_894_n 0.00154949f $X=5.275 $Y=2.245
+ $X2=0 $Y2=0
cc_600 N_A_1007_366#_c_691_n N_A_868_368#_c_894_n 0.00954614f $X=5.28 $Y=1.83
+ $X2=0 $Y2=0
cc_601 N_A_1007_366#_c_711_n N_A_868_368#_c_894_n 0.0214227f $X=5.2 $Y=1.995
+ $X2=0 $Y2=0
cc_602 N_A_1007_366#_M1046_g N_A_868_368#_c_899_n 0.00302354f $X=9.435 $Y=0.9
+ $X2=0 $Y2=0
cc_603 N_A_1007_366#_c_696_n N_A_868_368#_c_899_n 0.0233215f $X=7.96 $Y=2.125
+ $X2=0 $Y2=0
cc_604 N_A_1007_366#_c_698_n N_A_868_368#_c_899_n 0.0068339f $X=9.78 $Y=1.745
+ $X2=0 $Y2=0
cc_605 N_A_1007_366#_c_699_n N_A_868_368#_c_899_n 0.00158735f $X=9.78 $Y=1.745
+ $X2=0 $Y2=0
cc_606 N_A_1007_366#_c_739_p N_A_868_368#_c_899_n 0.010897f $X=8.077 $Y=1.115
+ $X2=0 $Y2=0
cc_607 N_A_1007_366#_c_692_n N_A_868_368#_c_900_n 6.55392e-19 $X=5.775 $Y=1.195
+ $X2=0 $Y2=0
cc_608 N_A_1007_366#_M1046_g N_A_868_368#_c_901_n 0.00350432f $X=9.435 $Y=0.9
+ $X2=0 $Y2=0
cc_609 N_A_1007_366#_c_698_n N_A_868_368#_c_901_n 0.00944344f $X=9.78 $Y=1.745
+ $X2=0 $Y2=0
cc_610 N_A_1007_366#_c_699_n N_A_868_368#_c_901_n 6.28561e-19 $X=9.78 $Y=1.745
+ $X2=0 $Y2=0
cc_611 N_A_1007_366#_c_700_n N_A_868_368#_c_902_n 5.62442e-19 $X=5.275 $Y=2.245
+ $X2=0 $Y2=0
cc_612 N_A_1007_366#_c_691_n N_A_868_368#_c_902_n 0.0178578f $X=5.28 $Y=1.83
+ $X2=0 $Y2=0
cc_613 N_A_1007_366#_c_692_n N_A_868_368#_c_902_n 0.0181644f $X=5.775 $Y=1.195
+ $X2=0 $Y2=0
cc_614 N_A_1007_366#_M1046_g N_A_868_368#_c_903_n 0.00313065f $X=9.435 $Y=0.9
+ $X2=0 $Y2=0
cc_615 N_A_1007_366#_c_698_n N_A_868_368#_c_903_n 0.00190689f $X=9.78 $Y=1.745
+ $X2=0 $Y2=0
cc_616 N_A_1007_366#_c_699_n N_A_868_368#_c_903_n 0.03095f $X=9.78 $Y=1.745
+ $X2=0 $Y2=0
cc_617 N_A_1007_366#_c_691_n N_A_868_368#_c_904_n 0.00824257f $X=5.28 $Y=1.83
+ $X2=0 $Y2=0
cc_618 N_A_1007_366#_c_692_n N_A_868_368#_c_904_n 0.00988844f $X=5.775 $Y=1.195
+ $X2=0 $Y2=0
cc_619 N_A_1007_366#_c_711_n N_A_868_368#_c_904_n 6.13001e-19 $X=5.2 $Y=1.995
+ $X2=0 $Y2=0
cc_620 N_A_1007_366#_c_712_n N_A_1154_464#_M1039_d 0.00287371f $X=6.9 $Y=2.902
+ $X2=0 $Y2=0
cc_621 N_A_1007_366#_c_696_n N_A_1154_464#_c_1101_n 0.0106061f $X=7.96 $Y=2.125
+ $X2=0 $Y2=0
cc_622 N_A_1007_366#_c_696_n N_A_1154_464#_c_1109_n 0.00382104f $X=7.96 $Y=2.125
+ $X2=0 $Y2=0
cc_623 N_A_1007_366#_c_756_p N_A_1154_464#_c_1109_n 0.0141783f $X=7.96 $Y=2.73
+ $X2=0 $Y2=0
cc_624 N_A_1007_366#_c_713_n N_A_1154_464#_c_1109_n 0.0138077f $X=7.66 $Y=2.815
+ $X2=0 $Y2=0
cc_625 N_A_1007_366#_c_758_p N_A_1154_464#_c_1109_n 0.00443638f $X=7.96 $Y=2.21
+ $X2=0 $Y2=0
cc_626 N_A_1007_366#_c_696_n N_A_1154_464#_c_1102_n 0.00326187f $X=7.96 $Y=2.125
+ $X2=0 $Y2=0
cc_627 N_A_1007_366#_c_697_n N_A_1154_464#_c_1102_n 0.0102469f $X=8.115 $Y=0.86
+ $X2=0 $Y2=0
cc_628 N_A_1007_366#_c_739_p N_A_1154_464#_c_1102_n 0.00492568f $X=8.077
+ $Y=1.115 $X2=0 $Y2=0
cc_629 N_A_1007_366#_c_696_n N_A_1154_464#_c_1103_n 0.00359245f $X=7.96 $Y=2.125
+ $X2=0 $Y2=0
cc_630 N_A_1007_366#_c_703_n N_A_1154_464#_c_1110_n 0.0277246f $X=5.47 $Y=2.905
+ $X2=0 $Y2=0
cc_631 N_A_1007_366#_c_712_n N_A_1154_464#_c_1110_n 0.0206186f $X=6.9 $Y=2.902
+ $X2=0 $Y2=0
cc_632 N_A_1007_366#_M1034_s N_A_1154_464#_c_1111_n 0.00758356f $X=6.92 $Y=2.12
+ $X2=0 $Y2=0
cc_633 N_A_1007_366#_c_703_n N_A_1154_464#_c_1112_n 0.0017365f $X=5.47 $Y=2.905
+ $X2=0 $Y2=0
cc_634 N_A_1007_366#_c_711_n N_A_1154_464#_c_1112_n 0.00893001f $X=5.2 $Y=1.995
+ $X2=0 $Y2=0
cc_635 N_A_1007_366#_c_696_n N_A_1643_257#_c_1217_n 0.00159585f $X=7.96 $Y=2.125
+ $X2=0 $Y2=0
cc_636 N_A_1007_366#_c_756_p N_A_1643_257#_c_1217_n 0.00524388f $X=7.96 $Y=2.73
+ $X2=0 $Y2=0
cc_637 N_A_1007_366#_c_770_p N_A_1643_257#_c_1217_n 0.0150529f $X=8.905 $Y=2.21
+ $X2=0 $Y2=0
cc_638 N_A_1007_366#_c_713_n N_A_1643_257#_c_1217_n 0.00192993f $X=7.66 $Y=2.815
+ $X2=0 $Y2=0
cc_639 N_A_1007_366#_c_714_n N_A_1643_257#_c_1217_n 0.00114671f $X=9.07 $Y=2.035
+ $X2=0 $Y2=0
cc_640 N_A_1007_366#_c_715_n N_A_1643_257#_c_1217_n 2.0116e-19 $X=9.07 $Y=2.265
+ $X2=0 $Y2=0
cc_641 N_A_1007_366#_c_696_n N_A_1643_257#_c_1202_n 0.00116211f $X=7.96 $Y=2.125
+ $X2=0 $Y2=0
cc_642 N_A_1007_366#_c_697_n N_A_1643_257#_c_1202_n 0.00448089f $X=8.115 $Y=0.86
+ $X2=0 $Y2=0
cc_643 N_A_1007_366#_c_739_p N_A_1643_257#_c_1202_n 0.00456437f $X=8.077
+ $Y=1.115 $X2=0 $Y2=0
cc_644 N_A_1007_366#_c_696_n N_A_1643_257#_c_1203_n 0.00448477f $X=7.96 $Y=2.125
+ $X2=0 $Y2=0
cc_645 N_A_1007_366#_c_770_p N_A_1643_257#_c_1203_n 9.52862e-19 $X=8.905 $Y=2.21
+ $X2=0 $Y2=0
cc_646 N_A_1007_366#_c_714_n N_A_1643_257#_c_1203_n 4.18161e-19 $X=9.07 $Y=2.035
+ $X2=0 $Y2=0
cc_647 N_A_1007_366#_M1046_g N_A_1643_257#_c_1204_n 0.0148208f $X=9.435 $Y=0.9
+ $X2=0 $Y2=0
cc_648 N_A_1007_366#_c_708_n N_A_1643_257#_c_1204_n 0.00189168f $X=9.615
+ $Y=2.035 $X2=0 $Y2=0
cc_649 N_A_1007_366#_c_698_n N_A_1643_257#_c_1204_n 0.00410116f $X=9.78 $Y=1.745
+ $X2=0 $Y2=0
cc_650 N_A_1007_366#_c_699_n N_A_1643_257#_c_1204_n 0.00298923f $X=9.78 $Y=1.745
+ $X2=0 $Y2=0
cc_651 N_A_1007_366#_M1046_g N_A_1643_257#_c_1205_n 0.00337498f $X=9.435 $Y=0.9
+ $X2=0 $Y2=0
cc_652 N_A_1007_366#_c_696_n N_A_1643_257#_c_1211_n 0.0556415f $X=7.96 $Y=2.125
+ $X2=0 $Y2=0
cc_653 N_A_1007_366#_c_770_p N_A_1643_257#_c_1211_n 0.0290352f $X=8.905 $Y=2.21
+ $X2=0 $Y2=0
cc_654 N_A_1007_366#_c_739_p N_A_1643_257#_c_1211_n 0.00290063f $X=8.077
+ $Y=1.115 $X2=0 $Y2=0
cc_655 N_A_1007_366#_c_714_n N_A_1643_257#_c_1211_n 2.49034e-19 $X=9.07 $Y=2.035
+ $X2=0 $Y2=0
cc_656 N_A_1007_366#_c_696_n N_A_1643_257#_c_1212_n 5.71848e-19 $X=7.96 $Y=2.125
+ $X2=0 $Y2=0
cc_657 N_A_1007_366#_c_708_n N_SET_B_c_1415_n 3.22493e-19 $X=9.615 $Y=2.035
+ $X2=0 $Y2=0
cc_658 N_A_1007_366#_c_698_n N_SET_B_c_1415_n 0.00137285f $X=9.78 $Y=1.745 $X2=0
+ $Y2=0
cc_659 N_A_1007_366#_c_699_n N_SET_B_c_1415_n 0.0045314f $X=9.78 $Y=1.745 $X2=0
+ $Y2=0
cc_660 N_A_1007_366#_c_714_n N_SET_B_c_1415_n 4.1911e-19 $X=9.07 $Y=2.035 $X2=0
+ $Y2=0
cc_661 N_A_1007_366#_c_770_p N_SET_B_c_1416_n 0.0143374f $X=8.905 $Y=2.21 $X2=0
+ $Y2=0
cc_662 N_A_1007_366#_c_708_n N_SET_B_c_1416_n 2.45687e-19 $X=9.615 $Y=2.035
+ $X2=0 $Y2=0
cc_663 N_A_1007_366#_c_714_n N_SET_B_c_1416_n 0.0077824f $X=9.07 $Y=2.035 $X2=0
+ $Y2=0
cc_664 N_A_1007_366#_c_715_n N_SET_B_c_1416_n 0.0124644f $X=9.07 $Y=2.265 $X2=0
+ $Y2=0
cc_665 N_A_1007_366#_M1046_g N_SET_B_M1047_g 0.0260735f $X=9.435 $Y=0.9 $X2=0
+ $Y2=0
cc_666 N_A_1007_366#_c_697_n N_SET_B_M1047_g 7.78613e-19 $X=8.115 $Y=0.86 $X2=0
+ $Y2=0
cc_667 N_A_1007_366#_c_708_n N_SET_B_c_1408_n 0.00288187f $X=9.615 $Y=2.035
+ $X2=0 $Y2=0
cc_668 N_A_1007_366#_c_698_n N_SET_B_c_1408_n 0.0209753f $X=9.78 $Y=1.745 $X2=0
+ $Y2=0
cc_669 N_A_1007_366#_c_699_n N_SET_B_c_1408_n 0.0019492f $X=9.78 $Y=1.745 $X2=0
+ $Y2=0
cc_670 N_A_1007_366#_M1046_g N_SET_B_c_1420_n 0.00146728f $X=9.435 $Y=0.9 $X2=0
+ $Y2=0
cc_671 N_A_1007_366#_c_708_n N_SET_B_c_1420_n 0.00726112f $X=9.615 $Y=2.035
+ $X2=0 $Y2=0
cc_672 N_A_1007_366#_c_698_n N_SET_B_c_1420_n 0.0016174f $X=9.78 $Y=1.745 $X2=0
+ $Y2=0
cc_673 N_A_1007_366#_c_699_n N_SET_B_c_1420_n 0.00166115f $X=9.78 $Y=1.745 $X2=0
+ $Y2=0
cc_674 N_A_1007_366#_c_714_n N_SET_B_c_1420_n 5.39857e-19 $X=9.07 $Y=2.035 $X2=0
+ $Y2=0
cc_675 N_A_1007_366#_M1046_g N_SET_B_c_1409_n 0.00832335f $X=9.435 $Y=0.9 $X2=0
+ $Y2=0
cc_676 N_A_1007_366#_c_770_p N_SET_B_c_1409_n 0.00465613f $X=8.905 $Y=2.21 $X2=0
+ $Y2=0
cc_677 N_A_1007_366#_c_708_n N_SET_B_c_1409_n 0.0136834f $X=9.615 $Y=2.035 $X2=0
+ $Y2=0
cc_678 N_A_1007_366#_c_698_n N_SET_B_c_1409_n 0.0129338f $X=9.78 $Y=1.745 $X2=0
+ $Y2=0
cc_679 N_A_1007_366#_c_699_n N_SET_B_c_1409_n 0.00556251f $X=9.78 $Y=1.745 $X2=0
+ $Y2=0
cc_680 N_A_1007_366#_c_714_n N_SET_B_c_1409_n 0.0270009f $X=9.07 $Y=2.035 $X2=0
+ $Y2=0
cc_681 N_A_1007_366#_M1046_g N_SET_B_c_1411_n 0.0181567f $X=9.435 $Y=0.9 $X2=0
+ $Y2=0
cc_682 N_A_1007_366#_c_714_n N_SET_B_c_1411_n 0.00460551f $X=9.07 $Y=2.035 $X2=0
+ $Y2=0
cc_683 N_A_1007_366#_c_700_n N_A_688_98#_c_1560_n 0.00167644f $X=5.275 $Y=2.245
+ $X2=0 $Y2=0
cc_684 N_A_1007_366#_c_693_n N_A_688_98#_M1043_g 0.00485477f $X=5.355 $Y=1.195
+ $X2=0 $Y2=0
cc_685 N_A_1007_366#_c_694_n N_A_688_98#_c_1547_n 0.00862445f $X=5.85 $Y=1.12
+ $X2=0 $Y2=0
cc_686 N_A_1007_366#_c_694_n N_A_688_98#_M1016_g 0.0447055f $X=5.85 $Y=1.12
+ $X2=0 $Y2=0
cc_687 N_A_1007_366#_M1046_g N_A_688_98#_c_1550_n 0.00894529f $X=9.435 $Y=0.9
+ $X2=0 $Y2=0
cc_688 N_A_1007_366#_M1046_g N_A_688_98#_M1020_g 0.0204245f $X=9.435 $Y=0.9
+ $X2=0 $Y2=0
cc_689 N_A_1007_366#_c_698_n N_A_688_98#_c_1553_n 7.66191e-19 $X=9.78 $Y=1.745
+ $X2=0 $Y2=0
cc_690 N_A_1007_366#_c_699_n N_A_688_98#_c_1553_n 0.00332218f $X=9.78 $Y=1.745
+ $X2=0 $Y2=0
cc_691 N_A_1007_366#_c_703_n N_A_688_98#_c_1565_n 0.00103605f $X=5.47 $Y=2.905
+ $X2=0 $Y2=0
cc_692 N_A_1007_366#_c_706_n N_A_688_98#_c_1565_n 0.00456723f $X=7.072 $Y=2.902
+ $X2=0 $Y2=0
cc_693 N_A_1007_366#_c_712_n N_A_688_98#_c_1565_n 0.0174215f $X=6.9 $Y=2.902
+ $X2=0 $Y2=0
cc_694 N_A_1007_366#_c_691_n N_A_688_98#_c_1558_n 0.00485477f $X=5.28 $Y=1.83
+ $X2=0 $Y2=0
cc_695 N_A_1007_366#_c_702_n N_A_1997_82#_c_1942_n 0.00202904f $X=9.855 $Y=2.045
+ $X2=0 $Y2=0
cc_696 N_A_1007_366#_c_702_n N_A_1997_82#_c_1949_n 7.38698e-19 $X=9.855 $Y=2.045
+ $X2=0 $Y2=0
cc_697 N_A_1007_366#_c_708_n N_A_1997_82#_c_1949_n 9.59981e-19 $X=9.615 $Y=2.035
+ $X2=0 $Y2=0
cc_698 N_A_1007_366#_c_770_p N_VPWR_M1030_d 0.00899607f $X=8.905 $Y=2.21 $X2=0
+ $Y2=0
cc_699 N_A_1007_366#_c_708_n N_VPWR_M1009_s 0.00180215f $X=9.615 $Y=2.035 $X2=0
+ $Y2=0
cc_700 N_A_1007_366#_c_700_n N_VPWR_c_2239_n 0.00906771f $X=5.275 $Y=2.245 $X2=0
+ $Y2=0
cc_701 N_A_1007_366#_c_703_n N_VPWR_c_2239_n 0.0262296f $X=5.47 $Y=2.905 $X2=0
+ $Y2=0
cc_702 N_A_1007_366#_c_704_n N_VPWR_c_2239_n 0.0147459f $X=5.555 $Y=2.99 $X2=0
+ $Y2=0
cc_703 N_A_1007_366#_c_711_n N_VPWR_c_2239_n 0.01293f $X=5.2 $Y=1.995 $X2=0
+ $Y2=0
cc_704 N_A_1007_366#_c_756_p N_VPWR_c_2240_n 0.0120128f $X=7.96 $Y=2.73 $X2=0
+ $Y2=0
cc_705 N_A_1007_366#_c_770_p N_VPWR_c_2240_n 0.0219335f $X=8.905 $Y=2.21 $X2=0
+ $Y2=0
cc_706 N_A_1007_366#_c_713_n N_VPWR_c_2240_n 0.0140315f $X=7.66 $Y=2.815 $X2=0
+ $Y2=0
cc_707 N_A_1007_366#_c_715_n N_VPWR_c_2240_n 0.0340117f $X=9.07 $Y=2.265 $X2=0
+ $Y2=0
cc_708 N_A_1007_366#_c_702_n N_VPWR_c_2241_n 0.016195f $X=9.855 $Y=2.045 $X2=0
+ $Y2=0
cc_709 N_A_1007_366#_c_708_n N_VPWR_c_2241_n 0.0247912f $X=9.615 $Y=2.035 $X2=0
+ $Y2=0
cc_710 N_A_1007_366#_c_699_n N_VPWR_c_2241_n 9.66821e-19 $X=9.78 $Y=1.745 $X2=0
+ $Y2=0
cc_711 N_A_1007_366#_c_714_n N_VPWR_c_2241_n 0.0464852f $X=9.07 $Y=2.035 $X2=0
+ $Y2=0
cc_712 N_A_1007_366#_c_715_n N_VPWR_c_2249_n 0.0145938f $X=9.07 $Y=2.265 $X2=0
+ $Y2=0
cc_713 N_A_1007_366#_c_700_n N_VPWR_c_2258_n 0.00389876f $X=5.275 $Y=2.245 $X2=0
+ $Y2=0
cc_714 N_A_1007_366#_c_704_n N_VPWR_c_2258_n 0.0121867f $X=5.555 $Y=2.99 $X2=0
+ $Y2=0
cc_715 N_A_1007_366#_c_712_n N_VPWR_c_2258_n 0.137047f $X=6.9 $Y=2.902 $X2=0
+ $Y2=0
cc_716 N_A_1007_366#_c_713_n N_VPWR_c_2258_n 0.0176329f $X=7.66 $Y=2.815 $X2=0
+ $Y2=0
cc_717 N_A_1007_366#_c_702_n N_VPWR_c_2259_n 0.00413917f $X=9.855 $Y=2.045 $X2=0
+ $Y2=0
cc_718 N_A_1007_366#_c_700_n N_VPWR_c_2234_n 0.00434485f $X=5.275 $Y=2.245 $X2=0
+ $Y2=0
cc_719 N_A_1007_366#_c_702_n N_VPWR_c_2234_n 0.00817239f $X=9.855 $Y=2.045 $X2=0
+ $Y2=0
cc_720 N_A_1007_366#_c_704_n N_VPWR_c_2234_n 0.00660921f $X=5.555 $Y=2.99 $X2=0
+ $Y2=0
cc_721 N_A_1007_366#_c_712_n N_VPWR_c_2234_n 0.078629f $X=6.9 $Y=2.902 $X2=0
+ $Y2=0
cc_722 N_A_1007_366#_c_713_n N_VPWR_c_2234_n 0.0134714f $X=7.66 $Y=2.815 $X2=0
+ $Y2=0
cc_723 N_A_1007_366#_c_715_n N_VPWR_c_2234_n 0.0120466f $X=9.07 $Y=2.265 $X2=0
+ $Y2=0
cc_724 N_A_1007_366#_c_712_n N_A_197_119#_M1013_d 0.00356213f $X=6.9 $Y=2.902
+ $X2=0 $Y2=0
cc_725 N_A_1007_366#_c_694_n N_A_197_119#_c_2459_n 0.00293755f $X=5.85 $Y=1.12
+ $X2=0 $Y2=0
cc_726 N_A_1007_366#_c_693_n N_A_197_119#_c_2460_n 0.0105699f $X=5.355 $Y=1.195
+ $X2=0 $Y2=0
cc_727 N_A_1007_366#_c_694_n N_A_197_119#_c_2460_n 0.0108717f $X=5.85 $Y=1.12
+ $X2=0 $Y2=0
cc_728 N_A_1007_366#_c_693_n N_A_197_119#_c_2461_n 0.0021947f $X=5.355 $Y=1.195
+ $X2=0 $Y2=0
cc_729 N_A_1007_366#_c_694_n N_A_197_119#_c_2462_n 0.00170607f $X=5.85 $Y=1.12
+ $X2=0 $Y2=0
cc_730 N_A_1007_366#_M1034_s N_A_197_119#_c_2474_n 0.02781f $X=6.92 $Y=2.12
+ $X2=0 $Y2=0
cc_731 N_A_1007_366#_c_705_n N_A_197_119#_c_2474_n 0.0092162f $X=7.653 $Y=2.902
+ $X2=0 $Y2=0
cc_732 N_A_1007_366#_c_706_n N_A_197_119#_c_2474_n 0.0450538f $X=7.072 $Y=2.902
+ $X2=0 $Y2=0
cc_733 N_A_1007_366#_c_756_p N_A_197_119#_c_2474_n 0.0134181f $X=7.96 $Y=2.73
+ $X2=0 $Y2=0
cc_734 N_A_1007_366#_c_712_n N_A_197_119#_c_2474_n 0.00900428f $X=6.9 $Y=2.902
+ $X2=0 $Y2=0
cc_735 N_A_1007_366#_c_713_n N_A_197_119#_c_2474_n 0.00407712f $X=7.66 $Y=2.815
+ $X2=0 $Y2=0
cc_736 N_A_1007_366#_c_697_n N_A_197_119#_c_2466_n 0.00620554f $X=8.115 $Y=0.86
+ $X2=0 $Y2=0
cc_737 N_A_1007_366#_c_739_p N_A_197_119#_c_2466_n 0.00586459f $X=8.077 $Y=1.115
+ $X2=0 $Y2=0
cc_738 N_A_1007_366#_M1034_s N_A_197_119#_c_2468_n 0.0117748f $X=6.92 $Y=2.12
+ $X2=0 $Y2=0
cc_739 N_A_1007_366#_c_756_p N_A_197_119#_c_2468_n 0.00589718f $X=7.96 $Y=2.73
+ $X2=0 $Y2=0
cc_740 N_A_1007_366#_c_739_p N_A_197_119#_c_2468_n 0.0784277f $X=8.077 $Y=1.115
+ $X2=0 $Y2=0
cc_741 N_A_1007_366#_c_758_p N_A_197_119#_c_2468_n 0.0133617f $X=7.96 $Y=2.21
+ $X2=0 $Y2=0
cc_742 N_A_1007_366#_c_712_n N_A_197_119#_c_2477_n 0.0222541f $X=6.9 $Y=2.902
+ $X2=0 $Y2=0
cc_743 N_A_1007_366#_c_703_n A_1070_464# 0.00732705f $X=5.47 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_744 N_A_1007_366#_c_756_p A_1592_424# 0.00485784f $X=7.96 $Y=2.73 $X2=-0.19
+ $Y2=-0.245
cc_745 N_A_1007_366#_c_770_p A_1592_424# 0.00969151f $X=8.905 $Y=2.21 $X2=-0.19
+ $Y2=-0.245
cc_746 N_A_1007_366#_c_713_n A_1592_424# 0.00230347f $X=7.66 $Y=2.815 $X2=-0.19
+ $Y2=-0.245
cc_747 N_A_1007_366#_c_708_n A_1986_424# 6.1435e-19 $X=9.615 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_748 N_A_1007_366#_c_694_n N_VGND_c_2736_n 0.00386607f $X=5.85 $Y=1.12 $X2=0
+ $Y2=0
cc_749 N_A_1007_366#_M1046_g N_VGND_c_2737_n 0.00666708f $X=9.435 $Y=0.9 $X2=0
+ $Y2=0
cc_750 N_A_1007_366#_c_694_n N_VGND_c_2759_n 9.49986e-19 $X=5.85 $Y=1.12 $X2=0
+ $Y2=0
cc_751 N_A_1007_366#_M1046_g N_VGND_c_2759_n 7.97988e-19 $X=9.435 $Y=0.9 $X2=0
+ $Y2=0
cc_752 N_A_1007_366#_c_697_n N_A_1473_73#_c_2925_n 0.0253693f $X=8.115 $Y=0.86
+ $X2=0 $Y2=0
cc_753 N_A_1007_366#_c_739_p N_A_1473_73#_c_2925_n 0.00255767f $X=8.077 $Y=1.115
+ $X2=0 $Y2=0
cc_754 N_A_1007_366#_c_697_n N_A_1473_73#_c_2927_n 0.00329772f $X=8.115 $Y=0.86
+ $X2=0 $Y2=0
cc_755 N_A_1007_366#_c_697_n N_A_1473_73#_c_2928_n 0.0131504f $X=8.115 $Y=0.86
+ $X2=0 $Y2=0
cc_756 N_A_868_368#_c_899_n N_A_1154_464#_c_1099_n 0.0125145f $X=10.175 $Y=1.295
+ $X2=0 $Y2=0
cc_757 N_A_868_368#_M1006_g N_A_1154_464#_c_1100_n 0.0108764f $X=6.665 $Y=0.835
+ $X2=0 $Y2=0
cc_758 N_A_868_368#_c_899_n N_A_1154_464#_c_1102_n 0.0030464f $X=10.175 $Y=1.295
+ $X2=0 $Y2=0
cc_759 N_A_868_368#_c_899_n N_A_1154_464#_c_1103_n 0.00359786f $X=10.175
+ $Y=1.295 $X2=0 $Y2=0
cc_760 N_A_868_368#_c_906_n N_A_1154_464#_c_1110_n 0.00543049f $X=5.695 $Y=2.245
+ $X2=0 $Y2=0
cc_761 N_A_868_368#_c_896_n N_A_1154_464#_c_1111_n 0.023272f $X=6.66 $Y=1.69
+ $X2=0 $Y2=0
cc_762 N_A_868_368#_c_897_n N_A_1154_464#_c_1111_n 0.00790882f $X=6.66 $Y=1.69
+ $X2=0 $Y2=0
cc_763 N_A_868_368#_c_898_n N_A_1154_464#_c_1111_n 0.0219168f $X=6.495 $Y=1.69
+ $X2=0 $Y2=0
cc_764 N_A_868_368#_c_905_n N_A_1154_464#_c_1112_n 0.00194373f $X=5.695 $Y=2.155
+ $X2=0 $Y2=0
cc_765 N_A_868_368#_c_898_n N_A_1154_464#_c_1112_n 0.00402216f $X=6.495 $Y=1.69
+ $X2=0 $Y2=0
cc_766 N_A_868_368#_c_902_n N_A_1154_464#_c_1112_n 6.56837e-19 $X=5.76 $Y=1.675
+ $X2=0 $Y2=0
cc_767 N_A_868_368#_c_904_n N_A_1154_464#_c_1112_n 0.0224664f $X=5.855 $Y=1.265
+ $X2=0 $Y2=0
cc_768 N_A_868_368#_M1006_g N_A_1154_464#_c_1104_n 0.0139237f $X=6.665 $Y=0.835
+ $X2=0 $Y2=0
cc_769 N_A_868_368#_c_904_n N_A_1154_464#_c_1104_n 3.15813e-19 $X=5.855 $Y=1.265
+ $X2=0 $Y2=0
cc_770 N_A_868_368#_M1006_g N_A_1154_464#_c_1105_n 0.0115425f $X=6.665 $Y=0.835
+ $X2=0 $Y2=0
cc_771 N_A_868_368#_c_896_n N_A_1154_464#_c_1105_n 0.0133808f $X=6.66 $Y=1.69
+ $X2=0 $Y2=0
cc_772 N_A_868_368#_c_897_n N_A_1154_464#_c_1105_n 0.00186601f $X=6.66 $Y=1.69
+ $X2=0 $Y2=0
cc_773 N_A_868_368#_c_899_n N_A_1154_464#_c_1105_n 0.0298532f $X=10.175 $Y=1.295
+ $X2=0 $Y2=0
cc_774 N_A_868_368#_M1006_g N_A_1154_464#_c_1106_n 0.00271534f $X=6.665 $Y=0.835
+ $X2=0 $Y2=0
cc_775 N_A_868_368#_c_897_n N_A_1154_464#_c_1106_n 0.0021192f $X=6.66 $Y=1.69
+ $X2=0 $Y2=0
cc_776 N_A_868_368#_c_898_n N_A_1154_464#_c_1106_n 0.0228086f $X=6.495 $Y=1.69
+ $X2=0 $Y2=0
cc_777 N_A_868_368#_c_899_n N_A_1154_464#_c_1106_n 0.0241047f $X=10.175 $Y=1.295
+ $X2=0 $Y2=0
cc_778 N_A_868_368#_c_900_n N_A_1154_464#_c_1106_n 0.00104584f $X=6.145 $Y=1.295
+ $X2=0 $Y2=0
cc_779 N_A_868_368#_c_904_n N_A_1154_464#_c_1106_n 0.0118934f $X=5.855 $Y=1.265
+ $X2=0 $Y2=0
cc_780 N_A_868_368#_M1006_g N_A_1154_464#_c_1113_n 0.00107406f $X=6.665 $Y=0.835
+ $X2=0 $Y2=0
cc_781 N_A_868_368#_c_896_n N_A_1154_464#_c_1113_n 0.0221115f $X=6.66 $Y=1.69
+ $X2=0 $Y2=0
cc_782 N_A_868_368#_c_897_n N_A_1154_464#_c_1113_n 4.14293e-19 $X=6.66 $Y=1.69
+ $X2=0 $Y2=0
cc_783 N_A_868_368#_c_899_n N_A_1154_464#_c_1113_n 0.0181829f $X=10.175 $Y=1.295
+ $X2=0 $Y2=0
cc_784 N_A_868_368#_c_896_n N_A_1154_464#_c_1107_n 0.00114027f $X=6.66 $Y=1.69
+ $X2=0 $Y2=0
cc_785 N_A_868_368#_c_897_n N_A_1154_464#_c_1107_n 0.0207808f $X=6.66 $Y=1.69
+ $X2=0 $Y2=0
cc_786 N_A_868_368#_c_899_n N_A_1643_257#_c_1202_n 0.00629037f $X=10.175
+ $Y=1.295 $X2=0 $Y2=0
cc_787 N_A_868_368#_c_899_n N_A_1643_257#_c_1204_n 0.0494221f $X=10.175 $Y=1.295
+ $X2=0 $Y2=0
cc_788 N_A_868_368#_c_988_p N_A_1643_257#_c_1204_n 3.49597e-19 $X=10.32 $Y=1.295
+ $X2=0 $Y2=0
cc_789 N_A_868_368#_c_901_n N_A_1643_257#_c_1204_n 0.00320167f $X=10.32 $Y=1.295
+ $X2=0 $Y2=0
cc_790 N_A_868_368#_M1012_g N_A_1643_257#_c_1206_n 0.0128014f $X=11.16 $Y=0.62
+ $X2=0 $Y2=0
cc_791 N_A_868_368#_M1012_g N_A_1643_257#_c_1251_n 0.0036889f $X=11.16 $Y=0.62
+ $X2=0 $Y2=0
cc_792 N_A_868_368#_M1012_g N_A_1643_257#_c_1252_n 0.00129854f $X=11.16 $Y=0.62
+ $X2=0 $Y2=0
cc_793 N_A_868_368#_c_899_n N_A_1643_257#_c_1211_n 0.0360902f $X=10.175 $Y=1.295
+ $X2=0 $Y2=0
cc_794 N_A_868_368#_c_899_n N_A_1643_257#_c_1212_n 0.00121118f $X=10.175
+ $Y=1.295 $X2=0 $Y2=0
cc_795 N_A_868_368#_M1012_g N_A_1643_257#_c_1255_n 2.18093e-19 $X=11.16 $Y=0.62
+ $X2=0 $Y2=0
cc_796 N_A_868_368#_c_899_n N_SET_B_M1047_g 0.00243523f $X=10.175 $Y=1.295 $X2=0
+ $Y2=0
cc_797 N_A_868_368#_c_892_n N_SET_B_c_1408_n 0.0272571f $X=11.22 $Y=1.43 $X2=0
+ $Y2=0
cc_798 N_A_868_368#_c_893_n N_SET_B_c_1408_n 0.00602718f $X=11.22 $Y=1.43 $X2=0
+ $Y2=0
cc_799 N_A_868_368#_c_899_n N_SET_B_c_1408_n 0.0503643f $X=10.175 $Y=1.295 $X2=0
+ $Y2=0
cc_800 N_A_868_368#_c_988_p N_SET_B_c_1408_n 0.0229319f $X=10.32 $Y=1.295 $X2=0
+ $Y2=0
cc_801 N_A_868_368#_c_901_n N_SET_B_c_1408_n 0.0243046f $X=10.32 $Y=1.295 $X2=0
+ $Y2=0
cc_802 N_A_868_368#_c_903_n N_SET_B_c_1408_n 0.0013891f $X=10.32 $Y=1.59 $X2=0
+ $Y2=0
cc_803 N_A_868_368#_c_899_n N_SET_B_c_1420_n 0.0243346f $X=10.175 $Y=1.295 $X2=0
+ $Y2=0
cc_804 N_A_868_368#_c_899_n N_SET_B_c_1409_n 0.0129054f $X=10.175 $Y=1.295 $X2=0
+ $Y2=0
cc_805 N_A_868_368#_c_899_n N_SET_B_c_1411_n 0.00585216f $X=10.175 $Y=1.295
+ $X2=0 $Y2=0
cc_806 N_A_868_368#_c_910_n N_A_688_98#_c_1560_n 0.00845306f $X=4.49 $Y=2.005
+ $X2=0 $Y2=0
cc_807 N_A_868_368#_c_894_n N_A_688_98#_c_1560_n 0.00129893f $X=4.595 $Y=1.84
+ $X2=0 $Y2=0
cc_808 N_A_868_368#_c_929_n N_A_688_98#_M1043_g 0.0131546f $X=4.855 $Y=0.76
+ $X2=0 $Y2=0
cc_809 N_A_868_368#_c_895_n N_A_688_98#_M1043_g 0.00913092f $X=4.777 $Y=1.265
+ $X2=0 $Y2=0
cc_810 N_A_868_368#_c_905_n N_A_688_98#_M1016_g 0.00716615f $X=5.695 $Y=2.155
+ $X2=0 $Y2=0
cc_811 N_A_868_368#_M1006_g N_A_688_98#_M1016_g 0.024932f $X=6.665 $Y=0.835
+ $X2=0 $Y2=0
cc_812 N_A_868_368#_c_897_n N_A_688_98#_M1016_g 0.0212658f $X=6.66 $Y=1.69 $X2=0
+ $Y2=0
cc_813 N_A_868_368#_c_898_n N_A_688_98#_M1016_g 0.0125674f $X=6.495 $Y=1.69
+ $X2=0 $Y2=0
cc_814 N_A_868_368#_c_899_n N_A_688_98#_M1016_g 0.00700914f $X=10.175 $Y=1.295
+ $X2=0 $Y2=0
cc_815 N_A_868_368#_c_900_n N_A_688_98#_M1016_g 0.00383053f $X=6.145 $Y=1.295
+ $X2=0 $Y2=0
cc_816 N_A_868_368#_c_902_n N_A_688_98#_M1016_g 0.0212267f $X=5.76 $Y=1.675
+ $X2=0 $Y2=0
cc_817 N_A_868_368#_c_904_n N_A_688_98#_M1016_g 0.010272f $X=5.855 $Y=1.265
+ $X2=0 $Y2=0
cc_818 N_A_868_368#_M1006_g N_A_688_98#_c_1550_n 0.00737233f $X=6.665 $Y=0.835
+ $X2=0 $Y2=0
cc_819 N_A_868_368#_M1012_g N_A_688_98#_c_1552_n 0.0134642f $X=11.16 $Y=0.62
+ $X2=0 $Y2=0
cc_820 N_A_868_368#_c_892_n N_A_688_98#_c_1552_n 0.00521347f $X=11.22 $Y=1.43
+ $X2=0 $Y2=0
cc_821 N_A_868_368#_c_988_p N_A_688_98#_c_1552_n 0.00285289f $X=10.32 $Y=1.295
+ $X2=0 $Y2=0
cc_822 N_A_868_368#_c_901_n N_A_688_98#_c_1552_n 0.00649983f $X=10.32 $Y=1.295
+ $X2=0 $Y2=0
cc_823 N_A_868_368#_c_903_n N_A_688_98#_c_1552_n 0.0181286f $X=10.32 $Y=1.59
+ $X2=0 $Y2=0
cc_824 N_A_868_368#_c_899_n N_A_688_98#_c_1553_n 0.00695899f $X=10.175 $Y=1.295
+ $X2=0 $Y2=0
cc_825 N_A_868_368#_c_908_n N_A_688_98#_c_1562_n 0.00900277f $X=10.245 $Y=2.045
+ $X2=0 $Y2=0
cc_826 N_A_868_368#_c_892_n N_A_688_98#_c_1562_n 2.11037e-19 $X=11.22 $Y=1.43
+ $X2=0 $Y2=0
cc_827 N_A_868_368#_c_908_n N_A_688_98#_c_1564_n 0.0123454f $X=10.245 $Y=2.045
+ $X2=0 $Y2=0
cc_828 N_A_868_368#_c_906_n N_A_688_98#_c_1565_n 0.0184867f $X=5.695 $Y=2.245
+ $X2=0 $Y2=0
cc_829 N_A_868_368#_c_898_n N_A_688_98#_c_1565_n 2.19364e-19 $X=6.495 $Y=1.69
+ $X2=0 $Y2=0
cc_830 N_A_868_368#_c_907_n N_A_688_98#_c_1555_n 0.00834769f $X=10.245 $Y=1.955
+ $X2=0 $Y2=0
cc_831 N_A_868_368#_c_892_n N_A_688_98#_c_1555_n 0.0159935f $X=11.22 $Y=1.43
+ $X2=0 $Y2=0
cc_832 N_A_868_368#_c_893_n N_A_688_98#_c_1555_n 0.0214104f $X=11.22 $Y=1.43
+ $X2=0 $Y2=0
cc_833 N_A_868_368#_c_901_n N_A_688_98#_c_1555_n 0.00587313f $X=10.32 $Y=1.295
+ $X2=0 $Y2=0
cc_834 N_A_868_368#_c_903_n N_A_688_98#_c_1555_n 0.0220416f $X=10.32 $Y=1.59
+ $X2=0 $Y2=0
cc_835 N_A_868_368#_c_929_n N_A_688_98#_c_1556_n 0.00643303f $X=4.855 $Y=0.76
+ $X2=0 $Y2=0
cc_836 N_A_868_368#_c_910_n N_A_688_98#_c_1586_n 0.014113f $X=4.49 $Y=2.005
+ $X2=0 $Y2=0
cc_837 N_A_868_368#_c_910_n N_A_688_98#_c_1569_n 0.00819907f $X=4.49 $Y=2.005
+ $X2=0 $Y2=0
cc_838 N_A_868_368#_c_894_n N_A_688_98#_c_1569_n 0.00662407f $X=4.595 $Y=1.84
+ $X2=0 $Y2=0
cc_839 N_A_868_368#_c_910_n N_A_688_98#_c_1557_n 0.0031538f $X=4.49 $Y=2.005
+ $X2=0 $Y2=0
cc_840 N_A_868_368#_c_894_n N_A_688_98#_c_1557_n 0.0230802f $X=4.595 $Y=1.84
+ $X2=0 $Y2=0
cc_841 N_A_868_368#_c_895_n N_A_688_98#_c_1557_n 8.06475e-19 $X=4.777 $Y=1.265
+ $X2=0 $Y2=0
cc_842 N_A_868_368#_c_910_n N_A_688_98#_c_1558_n 0.00809743f $X=4.49 $Y=2.005
+ $X2=0 $Y2=0
cc_843 N_A_868_368#_c_894_n N_A_688_98#_c_1558_n 0.0146401f $X=4.595 $Y=1.84
+ $X2=0 $Y2=0
cc_844 N_A_868_368#_c_895_n N_A_688_98#_c_1558_n 4.16759e-19 $X=4.777 $Y=1.265
+ $X2=0 $Y2=0
cc_845 N_A_868_368#_c_929_n N_A_688_98#_c_1559_n 3.03589e-19 $X=4.855 $Y=0.76
+ $X2=0 $Y2=0
cc_846 N_A_868_368#_c_895_n N_A_688_98#_c_1559_n 0.00686048f $X=4.777 $Y=1.265
+ $X2=0 $Y2=0
cc_847 N_A_868_368#_c_893_n N_A_2216_410#_c_1742_n 0.00764195f $X=11.22 $Y=1.43
+ $X2=0 $Y2=0
cc_848 N_A_868_368#_M1012_g N_A_2216_410#_c_1727_n 0.0399286f $X=11.16 $Y=0.62
+ $X2=0 $Y2=0
cc_849 N_A_868_368#_M1012_g N_A_2216_410#_c_1728_n 0.00636512f $X=11.16 $Y=0.62
+ $X2=0 $Y2=0
cc_850 N_A_868_368#_c_892_n N_A_2216_410#_c_1728_n 3.44953e-19 $X=11.22 $Y=1.43
+ $X2=0 $Y2=0
cc_851 N_A_868_368#_c_893_n N_A_2216_410#_c_1728_n 0.0212501f $X=11.22 $Y=1.43
+ $X2=0 $Y2=0
cc_852 N_A_868_368#_c_908_n N_A_1997_82#_c_1942_n 0.0140341f $X=10.245 $Y=2.045
+ $X2=0 $Y2=0
cc_853 N_A_868_368#_c_907_n N_A_1997_82#_c_1943_n 6.88245e-19 $X=10.245 $Y=1.955
+ $X2=0 $Y2=0
cc_854 N_A_868_368#_c_908_n N_A_1997_82#_c_1943_n 2.90959e-19 $X=10.245 $Y=2.045
+ $X2=0 $Y2=0
cc_855 N_A_868_368#_c_892_n N_A_1997_82#_c_1944_n 0.0278715f $X=11.22 $Y=1.43
+ $X2=0 $Y2=0
cc_856 N_A_868_368#_c_893_n N_A_1997_82#_c_1944_n 0.00261045f $X=11.22 $Y=1.43
+ $X2=0 $Y2=0
cc_857 N_A_868_368#_c_907_n N_A_1997_82#_c_1945_n 9.0435e-19 $X=10.245 $Y=1.955
+ $X2=0 $Y2=0
cc_858 N_A_868_368#_c_892_n N_A_1997_82#_c_1945_n 0.010348f $X=11.22 $Y=1.43
+ $X2=0 $Y2=0
cc_859 N_A_868_368#_c_901_n N_A_1997_82#_c_1945_n 2.88219e-19 $X=10.32 $Y=1.295
+ $X2=0 $Y2=0
cc_860 N_A_868_368#_M1012_g N_A_1997_82#_c_1937_n 0.00924867f $X=11.16 $Y=0.62
+ $X2=0 $Y2=0
cc_861 N_A_868_368#_c_892_n N_A_1997_82#_c_1937_n 0.0193121f $X=11.22 $Y=1.43
+ $X2=0 $Y2=0
cc_862 N_A_868_368#_c_893_n N_A_1997_82#_c_1937_n 0.00342275f $X=11.22 $Y=1.43
+ $X2=0 $Y2=0
cc_863 N_A_868_368#_M1012_g N_A_1997_82#_c_1938_n 0.00276073f $X=11.16 $Y=0.62
+ $X2=0 $Y2=0
cc_864 N_A_868_368#_c_892_n N_A_1997_82#_c_1938_n 0.0238149f $X=11.22 $Y=1.43
+ $X2=0 $Y2=0
cc_865 N_A_868_368#_c_893_n N_A_1997_82#_c_1938_n 0.00152446f $X=11.22 $Y=1.43
+ $X2=0 $Y2=0
cc_866 N_A_868_368#_c_908_n N_A_1997_82#_c_1949_n 0.00403823f $X=10.245 $Y=2.045
+ $X2=0 $Y2=0
cc_867 N_A_868_368#_c_892_n N_A_1997_82#_c_1949_n 0.00399039f $X=11.22 $Y=1.43
+ $X2=0 $Y2=0
cc_868 N_A_868_368#_c_901_n N_A_1997_82#_c_1949_n 0.00685826f $X=10.32 $Y=1.295
+ $X2=0 $Y2=0
cc_869 N_A_868_368#_c_903_n N_A_1997_82#_c_1949_n 9.01994e-19 $X=10.32 $Y=1.59
+ $X2=0 $Y2=0
cc_870 N_A_868_368#_M1012_g N_A_1997_82#_c_1939_n 0.0103143f $X=11.16 $Y=0.62
+ $X2=0 $Y2=0
cc_871 N_A_868_368#_c_892_n N_A_1997_82#_c_1939_n 0.0322743f $X=11.22 $Y=1.43
+ $X2=0 $Y2=0
cc_872 N_A_868_368#_c_893_n N_A_1997_82#_c_1939_n 7.0447e-19 $X=11.22 $Y=1.43
+ $X2=0 $Y2=0
cc_873 N_A_868_368#_c_899_n N_A_1997_82#_c_1939_n 0.00757497f $X=10.175 $Y=1.295
+ $X2=0 $Y2=0
cc_874 N_A_868_368#_c_988_p N_A_1997_82#_c_1939_n 0.00211868f $X=10.32 $Y=1.295
+ $X2=0 $Y2=0
cc_875 N_A_868_368#_c_901_n N_A_1997_82#_c_1939_n 0.0108475f $X=10.32 $Y=1.295
+ $X2=0 $Y2=0
cc_876 N_A_868_368#_c_909_n N_VPWR_c_2237_n 0.0478153f $X=4.49 $Y=2.815 $X2=0
+ $Y2=0
cc_877 N_A_868_368#_c_909_n N_VPWR_c_2238_n 0.0168667f $X=4.49 $Y=2.815 $X2=0
+ $Y2=0
cc_878 N_A_868_368#_c_909_n N_VPWR_c_2239_n 0.0493206f $X=4.49 $Y=2.815 $X2=0
+ $Y2=0
cc_879 N_A_868_368#_c_908_n N_VPWR_c_2241_n 0.00248208f $X=10.245 $Y=2.045 $X2=0
+ $Y2=0
cc_880 N_A_868_368#_c_908_n N_VPWR_c_2259_n 0.00445602f $X=10.245 $Y=2.045 $X2=0
+ $Y2=0
cc_881 N_A_868_368#_c_908_n N_VPWR_c_2234_n 0.00858657f $X=10.245 $Y=2.045 $X2=0
+ $Y2=0
cc_882 N_A_868_368#_c_909_n N_VPWR_c_2234_n 0.0139608f $X=4.49 $Y=2.815 $X2=0
+ $Y2=0
cc_883 N_A_868_368#_c_929_n N_A_197_119#_c_2457_n 0.016761f $X=4.855 $Y=0.76
+ $X2=0 $Y2=0
cc_884 N_A_868_368#_c_929_n N_A_197_119#_c_2459_n 0.0186129f $X=4.855 $Y=0.76
+ $X2=0 $Y2=0
cc_885 N_A_868_368#_c_891_n N_A_197_119#_c_2460_n 0.0221874f $X=5.595 $Y=1.265
+ $X2=0 $Y2=0
cc_886 N_A_868_368#_c_900_n N_A_197_119#_c_2460_n 0.00209831f $X=6.145 $Y=1.295
+ $X2=0 $Y2=0
cc_887 N_A_868_368#_c_904_n N_A_197_119#_c_2460_n 0.0328006f $X=5.855 $Y=1.265
+ $X2=0 $Y2=0
cc_888 N_A_868_368#_c_929_n N_A_197_119#_c_2461_n 0.0145003f $X=4.855 $Y=0.76
+ $X2=0 $Y2=0
cc_889 N_A_868_368#_c_891_n N_A_197_119#_c_2461_n 0.0140745f $X=5.595 $Y=1.265
+ $X2=0 $Y2=0
cc_890 N_A_868_368#_M1006_g N_A_197_119#_c_2463_n 0.00330783f $X=6.665 $Y=0.835
+ $X2=0 $Y2=0
cc_891 N_A_868_368#_M1006_g N_A_197_119#_c_2465_n 0.00799322f $X=6.665 $Y=0.835
+ $X2=0 $Y2=0
cc_892 N_A_868_368#_c_899_n N_A_197_119#_c_2466_n 0.00913521f $X=10.175 $Y=1.295
+ $X2=0 $Y2=0
cc_893 N_A_868_368#_c_899_n N_A_197_119#_c_2467_n 0.00257612f $X=10.175 $Y=1.295
+ $X2=0 $Y2=0
cc_894 N_A_868_368#_c_899_n N_A_197_119#_c_2468_n 0.017403f $X=10.175 $Y=1.295
+ $X2=0 $Y2=0
cc_895 N_A_868_368#_c_899_n N_VGND_c_2737_n 0.00213546f $X=10.175 $Y=1.295 $X2=0
+ $Y2=0
cc_896 N_A_868_368#_M1012_g N_VGND_c_2738_n 9.08817e-19 $X=11.16 $Y=0.62 $X2=0
+ $Y2=0
cc_897 N_A_868_368#_c_899_n N_A_1473_73#_c_2927_n 0.00319761f $X=10.175 $Y=1.295
+ $X2=0 $Y2=0
cc_898 N_A_868_368#_c_899_n N_A_1473_73#_c_2928_n 0.00265792f $X=10.175 $Y=1.295
+ $X2=0 $Y2=0
cc_899 N_A_1154_464#_c_1109_n N_A_1643_257#_c_1217_n 0.0453692f $X=7.885
+ $Y=2.045 $X2=0 $Y2=0
cc_900 N_A_1154_464#_c_1102_n N_A_1643_257#_c_1202_n 0.0173121f $X=7.9 $Y=1.285
+ $X2=0 $Y2=0
cc_901 N_A_1154_464#_c_1101_n N_A_1643_257#_c_1203_n 0.0200671f $X=7.885
+ $Y=1.955 $X2=0 $Y2=0
cc_902 N_A_1154_464#_c_1101_n N_A_1643_257#_c_1211_n 5.19903e-19 $X=7.885
+ $Y=1.955 $X2=0 $Y2=0
cc_903 N_A_1154_464#_c_1103_n N_A_1643_257#_c_1211_n 2.66045e-19 $X=7.885
+ $Y=1.36 $X2=0 $Y2=0
cc_904 N_A_1154_464#_c_1103_n N_A_1643_257#_c_1212_n 0.0200671f $X=7.885 $Y=1.36
+ $X2=0 $Y2=0
cc_905 N_A_1154_464#_c_1111_n N_A_688_98#_M1016_g 0.00354424f $X=7.035 $Y=2.125
+ $X2=0 $Y2=0
cc_906 N_A_1154_464#_c_1112_n N_A_688_98#_M1016_g 0.00135573f $X=6.17 $Y=2.125
+ $X2=0 $Y2=0
cc_907 N_A_1154_464#_c_1104_n N_A_688_98#_M1016_g 0.00431122f $X=6.45 $Y=0.835
+ $X2=0 $Y2=0
cc_908 N_A_1154_464#_c_1106_n N_A_688_98#_M1016_g 0.00146824f $X=6.615 $Y=1.27
+ $X2=0 $Y2=0
cc_909 N_A_1154_464#_c_1102_n N_A_688_98#_c_1550_n 0.00737233f $X=7.9 $Y=1.285
+ $X2=0 $Y2=0
cc_910 N_A_1154_464#_c_1110_n N_A_688_98#_c_1565_n 0.0130895f $X=6.005 $Y=2.515
+ $X2=0 $Y2=0
cc_911 N_A_1154_464#_c_1111_n N_A_688_98#_c_1565_n 0.0113715f $X=7.035 $Y=2.125
+ $X2=0 $Y2=0
cc_912 N_A_1154_464#_c_1112_n N_A_688_98#_c_1565_n 0.0017429f $X=6.17 $Y=2.125
+ $X2=0 $Y2=0
cc_913 N_A_1154_464#_c_1109_n N_VPWR_c_2240_n 0.00100347f $X=7.885 $Y=2.045
+ $X2=0 $Y2=0
cc_914 N_A_1154_464#_c_1109_n N_VPWR_c_2258_n 0.00299636f $X=7.885 $Y=2.045
+ $X2=0 $Y2=0
cc_915 N_A_1154_464#_c_1109_n N_VPWR_c_2234_n 0.00373332f $X=7.885 $Y=2.045
+ $X2=0 $Y2=0
cc_916 N_A_1154_464#_c_1104_n N_A_197_119#_c_2462_n 0.0098261f $X=6.45 $Y=0.835
+ $X2=0 $Y2=0
cc_917 N_A_1154_464#_c_1104_n N_A_197_119#_c_2463_n 0.0258727f $X=6.45 $Y=0.835
+ $X2=0 $Y2=0
cc_918 N_A_1154_464#_c_1109_n N_A_197_119#_c_2474_n 0.00367705f $X=7.885
+ $Y=2.045 $X2=0 $Y2=0
cc_919 N_A_1154_464#_c_1111_n N_A_197_119#_c_2474_n 0.0268483f $X=7.035 $Y=2.125
+ $X2=0 $Y2=0
cc_920 N_A_1154_464#_c_1107_n N_A_197_119#_c_2474_n 0.00128531f $X=7.2 $Y=1.45
+ $X2=0 $Y2=0
cc_921 N_A_1154_464#_c_1104_n N_A_197_119#_c_2465_n 0.00979587f $X=6.45 $Y=0.835
+ $X2=0 $Y2=0
cc_922 N_A_1154_464#_c_1099_n N_A_197_119#_c_2466_n 0.0047529f $X=7.795 $Y=1.36
+ $X2=0 $Y2=0
cc_923 N_A_1154_464#_c_1100_n N_A_197_119#_c_2466_n 0.00134296f $X=7.365 $Y=1.36
+ $X2=0 $Y2=0
cc_924 N_A_1154_464#_c_1102_n N_A_197_119#_c_2466_n 0.00374247f $X=7.9 $Y=1.285
+ $X2=0 $Y2=0
cc_925 N_A_1154_464#_c_1105_n N_A_197_119#_c_2466_n 0.0194567f $X=7.035 $Y=1.27
+ $X2=0 $Y2=0
cc_926 N_A_1154_464#_c_1100_n N_A_197_119#_c_2467_n 4.86892e-19 $X=7.365 $Y=1.36
+ $X2=0 $Y2=0
cc_927 N_A_1154_464#_c_1105_n N_A_197_119#_c_2467_n 0.0250229f $X=7.035 $Y=1.27
+ $X2=0 $Y2=0
cc_928 N_A_1154_464#_c_1099_n N_A_197_119#_c_2468_n 0.0131848f $X=7.795 $Y=1.36
+ $X2=0 $Y2=0
cc_929 N_A_1154_464#_c_1101_n N_A_197_119#_c_2468_n 0.00636113f $X=7.885
+ $Y=1.955 $X2=0 $Y2=0
cc_930 N_A_1154_464#_c_1109_n N_A_197_119#_c_2468_n 0.00689017f $X=7.885
+ $Y=2.045 $X2=0 $Y2=0
cc_931 N_A_1154_464#_c_1102_n N_A_197_119#_c_2468_n 0.00523896f $X=7.9 $Y=1.285
+ $X2=0 $Y2=0
cc_932 N_A_1154_464#_c_1111_n N_A_197_119#_c_2468_n 0.014079f $X=7.035 $Y=2.125
+ $X2=0 $Y2=0
cc_933 N_A_1154_464#_c_1105_n N_A_197_119#_c_2468_n 0.0123301f $X=7.035 $Y=1.27
+ $X2=0 $Y2=0
cc_934 N_A_1154_464#_c_1113_n N_A_197_119#_c_2468_n 0.0513584f $X=7.2 $Y=1.45
+ $X2=0 $Y2=0
cc_935 N_A_1154_464#_c_1107_n N_A_197_119#_c_2468_n 0.00415297f $X=7.2 $Y=1.45
+ $X2=0 $Y2=0
cc_936 N_A_1154_464#_c_1111_n N_A_197_119#_c_2477_n 0.0520475f $X=7.035 $Y=2.125
+ $X2=0 $Y2=0
cc_937 N_A_1154_464#_c_1102_n N_A_1473_73#_c_2925_n 0.0023857f $X=7.9 $Y=1.285
+ $X2=0 $Y2=0
cc_938 N_A_1154_464#_c_1099_n N_A_1473_73#_c_2927_n 0.00207968f $X=7.795 $Y=1.36
+ $X2=0 $Y2=0
cc_939 N_A_1154_464#_c_1102_n N_A_1473_73#_c_2927_n 0.0061858f $X=7.9 $Y=1.285
+ $X2=0 $Y2=0
cc_940 N_A_1643_257#_c_1217_n N_SET_B_c_1416_n 0.0231197f $X=8.305 $Y=2.045
+ $X2=0 $Y2=0
cc_941 N_A_1643_257#_c_1203_n N_SET_B_c_1416_n 0.00328086f $X=8.38 $Y=1.79 $X2=0
+ $Y2=0
cc_942 N_A_1643_257#_c_1202_n N_SET_B_M1047_g 0.0131958f $X=8.38 $Y=1.285 $X2=0
+ $Y2=0
cc_943 N_A_1643_257#_c_1204_n N_SET_B_M1047_g 0.0140929f $X=9.555 $Y=1.195 $X2=0
+ $Y2=0
cc_944 N_A_1643_257#_c_1211_n N_SET_B_M1047_g 0.00329771f $X=8.38 $Y=1.45 $X2=0
+ $Y2=0
cc_945 N_A_1643_257#_c_1212_n N_SET_B_M1047_g 0.00630924f $X=8.38 $Y=1.45 $X2=0
+ $Y2=0
cc_946 N_A_1643_257#_c_1201_n N_SET_B_c_1407_n 0.00571788f $X=12.705 $Y=1.795
+ $X2=0 $Y2=0
cc_947 N_A_1643_257#_c_1219_n N_SET_B_c_1418_n 0.0385192f $X=12.705 $Y=1.885
+ $X2=0 $Y2=0
cc_948 N_A_1643_257#_c_1204_n N_SET_B_c_1408_n 5.02172e-19 $X=9.555 $Y=1.195
+ $X2=0 $Y2=0
cc_949 N_A_1643_257#_c_1204_n N_SET_B_c_1420_n 6.37746e-19 $X=9.555 $Y=1.195
+ $X2=0 $Y2=0
cc_950 N_A_1643_257#_c_1211_n N_SET_B_c_1420_n 7.94041e-19 $X=8.38 $Y=1.45 $X2=0
+ $Y2=0
cc_951 N_A_1643_257#_c_1203_n N_SET_B_c_1409_n 3.32748e-19 $X=8.38 $Y=1.79 $X2=0
+ $Y2=0
cc_952 N_A_1643_257#_c_1204_n N_SET_B_c_1409_n 0.0424892f $X=9.555 $Y=1.195
+ $X2=0 $Y2=0
cc_953 N_A_1643_257#_c_1211_n N_SET_B_c_1409_n 0.0273649f $X=8.38 $Y=1.45 $X2=0
+ $Y2=0
cc_954 N_A_1643_257#_c_1201_n SET_B 0.00306859f $X=12.705 $Y=1.795 $X2=0 $Y2=0
cc_955 N_A_1643_257#_c_1277_p SET_B 0.00272157f $X=12.495 $Y=0.855 $X2=0 $Y2=0
cc_956 N_A_1643_257#_c_1203_n N_SET_B_c_1411_n 0.030989f $X=8.38 $Y=1.79 $X2=0
+ $Y2=0
cc_957 N_A_1643_257#_c_1204_n N_SET_B_c_1411_n 0.00553531f $X=9.555 $Y=1.195
+ $X2=0 $Y2=0
cc_958 N_A_1643_257#_c_1211_n N_SET_B_c_1411_n 0.00635226f $X=8.38 $Y=1.45 $X2=0
+ $Y2=0
cc_959 N_A_1643_257#_c_1255_n N_SET_B_c_1412_n 6.60906e-19 $X=11.98 $Y=0.685
+ $X2=0 $Y2=0
cc_960 N_A_1643_257#_c_1213_n N_SET_B_c_1412_n 3.80681e-19 $X=12.66 $Y=1.215
+ $X2=0 $Y2=0
cc_961 N_A_1643_257#_c_1214_n N_SET_B_c_1412_n 0.0206294f $X=12.66 $Y=1.385
+ $X2=0 $Y2=0
cc_962 N_A_1643_257#_c_1201_n N_SET_B_c_1413_n 0.00267378f $X=12.705 $Y=1.795
+ $X2=0 $Y2=0
cc_963 N_A_1643_257#_c_1277_p N_SET_B_c_1413_n 0.0121625f $X=12.495 $Y=0.855
+ $X2=0 $Y2=0
cc_964 N_A_1643_257#_c_1255_n N_SET_B_c_1413_n 0.00691486f $X=11.98 $Y=0.685
+ $X2=0 $Y2=0
cc_965 N_A_1643_257#_c_1213_n N_SET_B_c_1413_n 0.0297148f $X=12.66 $Y=1.215
+ $X2=0 $Y2=0
cc_966 N_A_1643_257#_c_1214_n N_SET_B_c_1413_n 0.00188197f $X=12.66 $Y=1.385
+ $X2=0 $Y2=0
cc_967 N_A_1643_257#_c_1251_n N_SET_B_c_1414_n 7.62389e-19 $X=11.425 $Y=0.6
+ $X2=0 $Y2=0
cc_968 N_A_1643_257#_c_1277_p N_SET_B_c_1414_n 0.0116228f $X=12.495 $Y=0.855
+ $X2=0 $Y2=0
cc_969 N_A_1643_257#_c_1291_p N_SET_B_c_1414_n 0.00488698f $X=12.66 $Y=1.13
+ $X2=0 $Y2=0
cc_970 N_A_1643_257#_c_1216_n N_SET_B_c_1414_n 0.0191139f $X=12.66 $Y=1.22 $X2=0
+ $Y2=0
cc_971 N_A_1643_257#_c_1202_n N_A_688_98#_c_1550_n 0.00737233f $X=8.38 $Y=1.285
+ $X2=0 $Y2=0
cc_972 N_A_1643_257#_c_1206_n N_A_688_98#_c_1550_n 4.65214e-19 $X=11.34 $Y=0.345
+ $X2=0 $Y2=0
cc_973 N_A_1643_257#_c_1207_n N_A_688_98#_c_1550_n 0.0041955f $X=9.725 $Y=0.345
+ $X2=0 $Y2=0
cc_974 N_A_1643_257#_c_1205_n N_A_688_98#_M1020_g 0.012723f $X=9.64 $Y=1.11
+ $X2=0 $Y2=0
cc_975 N_A_1643_257#_c_1206_n N_A_688_98#_M1020_g 0.0169448f $X=11.34 $Y=0.345
+ $X2=0 $Y2=0
cc_976 N_A_1643_257#_c_1204_n N_A_688_98#_c_1553_n 0.00230751f $X=9.555 $Y=1.195
+ $X2=0 $Y2=0
cc_977 N_A_1643_257#_c_1206_n N_A_2216_410#_c_1727_n 0.00370663f $X=11.34
+ $Y=0.345 $X2=0 $Y2=0
cc_978 N_A_1643_257#_c_1251_n N_A_2216_410#_c_1727_n 0.00450139f $X=11.425
+ $Y=0.6 $X2=0 $Y2=0
cc_979 N_A_1643_257#_c_1301_p N_A_2216_410#_c_1727_n 0.00793623f $X=11.895
+ $Y=0.685 $X2=0 $Y2=0
cc_980 N_A_1643_257#_c_1252_n N_A_2216_410#_c_1727_n 0.00208735f $X=11.51
+ $Y=0.685 $X2=0 $Y2=0
cc_981 N_A_1643_257#_c_1255_n N_A_2216_410#_c_1727_n 0.00290549f $X=11.98
+ $Y=0.685 $X2=0 $Y2=0
cc_982 N_A_1643_257#_c_1301_p N_A_2216_410#_c_1736_n 0.00347296f $X=11.895
+ $Y=0.685 $X2=0 $Y2=0
cc_983 N_A_1643_257#_c_1255_n N_A_2216_410#_c_1736_n 7.95569e-19 $X=11.98
+ $Y=0.685 $X2=0 $Y2=0
cc_984 N_A_1643_257#_c_1219_n N_A_2216_410#_c_1769_n 0.0157446f $X=12.705
+ $Y=1.885 $X2=0 $Y2=0
cc_985 N_A_1643_257#_c_1208_n N_A_2216_410#_c_1737_n 0.0216222f $X=13.605
+ $Y=1.215 $X2=0 $Y2=0
cc_986 N_A_1643_257#_c_1210_n N_A_2216_410#_c_1737_n 0.0267417f $X=13.985
+ $Y=1.17 $X2=0 $Y2=0
cc_987 N_A_1643_257#_c_1215_n N_A_2216_410#_c_1737_n 0.0143583f $X=13.69 $Y=1.17
+ $X2=0 $Y2=0
cc_988 N_A_1643_257#_M1026_s N_A_2216_410#_c_1751_n 0.00331364f $X=13.765
+ $Y=1.995 $X2=0 $Y2=0
cc_989 N_A_1643_257#_c_1223_n N_A_2216_410#_c_1751_n 0.0318661f $X=13.91 $Y=2.17
+ $X2=0 $Y2=0
cc_990 N_A_1643_257#_c_1223_n N_A_2216_410#_c_1752_n 0.0126401f $X=13.91 $Y=2.17
+ $X2=0 $Y2=0
cc_991 N_A_1643_257#_c_1219_n N_A_2216_410#_c_1754_n 8.66265e-19 $X=12.705
+ $Y=1.885 $X2=0 $Y2=0
cc_992 N_A_1643_257#_c_1208_n N_A_2216_410#_c_1777_n 0.0169915f $X=13.605
+ $Y=1.215 $X2=0 $Y2=0
cc_993 N_A_1643_257#_c_1219_n N_A_2216_410#_c_1778_n 0.00291257f $X=12.705
+ $Y=1.885 $X2=0 $Y2=0
cc_994 N_A_1643_257#_c_1223_n N_A_2216_410#_c_1778_n 0.0226806f $X=13.91 $Y=2.17
+ $X2=0 $Y2=0
cc_995 N_A_1643_257#_c_1210_n N_A_2216_410#_c_1740_n 0.0151454f $X=13.985
+ $Y=1.17 $X2=0 $Y2=0
cc_996 N_A_1643_257#_c_1206_n N_A_1997_82#_M1020_d 0.0105494f $X=11.34 $Y=0.345
+ $X2=-0.19 $Y2=-0.245
cc_997 N_A_1643_257#_c_1201_n N_A_1997_82#_c_1935_n 0.018592f $X=12.705 $Y=1.795
+ $X2=0 $Y2=0
cc_998 N_A_1643_257#_c_1219_n N_A_1997_82#_c_1935_n 0.0550342f $X=12.705
+ $Y=1.885 $X2=0 $Y2=0
cc_999 N_A_1643_257#_c_1208_n N_A_1997_82#_c_1935_n 0.00125334f $X=13.605
+ $Y=1.215 $X2=0 $Y2=0
cc_1000 N_A_1643_257#_c_1209_n N_A_1997_82#_c_1935_n 0.00694786f $X=13.69
+ $Y=2.005 $X2=0 $Y2=0
cc_1001 N_A_1643_257#_c_1213_n N_A_1997_82#_c_1935_n 2.78633e-19 $X=12.66
+ $Y=1.215 $X2=0 $Y2=0
cc_1002 N_A_1643_257#_c_1214_n N_A_1997_82#_c_1935_n 0.00487525f $X=12.66
+ $Y=1.385 $X2=0 $Y2=0
cc_1003 N_A_1643_257#_c_1223_n N_A_1997_82#_c_1935_n 0.00124086f $X=13.91
+ $Y=2.17 $X2=0 $Y2=0
cc_1004 N_A_1643_257#_c_1208_n N_A_1997_82#_M1007_g 0.0140174f $X=13.605
+ $Y=1.215 $X2=0 $Y2=0
cc_1005 N_A_1643_257#_c_1209_n N_A_1997_82#_M1007_g 0.00361491f $X=13.69
+ $Y=2.005 $X2=0 $Y2=0
cc_1006 N_A_1643_257#_c_1213_n N_A_1997_82#_M1007_g 0.00123112f $X=12.66
+ $Y=1.215 $X2=0 $Y2=0
cc_1007 N_A_1643_257#_c_1291_p N_A_1997_82#_M1007_g 8.30634e-19 $X=12.66 $Y=1.13
+ $X2=0 $Y2=0
cc_1008 N_A_1643_257#_c_1214_n N_A_1997_82#_M1007_g 0.0141845f $X=12.66 $Y=1.385
+ $X2=0 $Y2=0
cc_1009 N_A_1643_257#_c_1215_n N_A_1997_82#_M1007_g 0.00499702f $X=13.69 $Y=1.17
+ $X2=0 $Y2=0
cc_1010 N_A_1643_257#_c_1216_n N_A_1997_82#_M1007_g 0.0264974f $X=12.66 $Y=1.22
+ $X2=0 $Y2=0
cc_1011 N_A_1643_257#_c_1206_n N_A_1997_82#_c_1937_n 0.00605937f $X=11.34
+ $Y=0.345 $X2=0 $Y2=0
cc_1012 N_A_1643_257#_c_1301_p N_A_1997_82#_c_1937_n 0.0140954f $X=11.895
+ $Y=0.685 $X2=0 $Y2=0
cc_1013 N_A_1643_257#_c_1252_n N_A_1997_82#_c_1937_n 0.0110616f $X=11.51
+ $Y=0.685 $X2=0 $Y2=0
cc_1014 N_A_1643_257#_c_1219_n N_A_1997_82#_c_1947_n 2.46149e-19 $X=12.705
+ $Y=1.885 $X2=0 $Y2=0
cc_1015 N_A_1643_257#_c_1201_n N_A_1997_82#_c_1948_n 0.00363067f $X=12.705
+ $Y=1.795 $X2=0 $Y2=0
cc_1016 N_A_1643_257#_c_1219_n N_A_1997_82#_c_1948_n 0.00494015f $X=12.705
+ $Y=1.885 $X2=0 $Y2=0
cc_1017 N_A_1643_257#_c_1208_n N_A_1997_82#_c_1948_n 0.00846624f $X=13.605
+ $Y=1.215 $X2=0 $Y2=0
cc_1018 N_A_1643_257#_c_1213_n N_A_1997_82#_c_1948_n 0.0117468f $X=12.66
+ $Y=1.215 $X2=0 $Y2=0
cc_1019 N_A_1643_257#_c_1214_n N_A_1997_82#_c_1948_n 2.04435e-19 $X=12.66
+ $Y=1.385 $X2=0 $Y2=0
cc_1020 N_A_1643_257#_c_1205_n N_A_1997_82#_c_1939_n 0.0151673f $X=9.64 $Y=1.11
+ $X2=0 $Y2=0
cc_1021 N_A_1643_257#_c_1206_n N_A_1997_82#_c_1939_n 0.0728842f $X=11.34
+ $Y=0.345 $X2=0 $Y2=0
cc_1022 N_A_1643_257#_c_1252_n N_A_1997_82#_c_1939_n 0.010457f $X=11.51 $Y=0.685
+ $X2=0 $Y2=0
cc_1023 N_A_1643_257#_c_1201_n N_A_1997_82#_c_1951_n 0.00182266f $X=12.705
+ $Y=1.795 $X2=0 $Y2=0
cc_1024 N_A_1643_257#_c_1219_n N_A_1997_82#_c_1951_n 0.00743416f $X=12.705
+ $Y=1.885 $X2=0 $Y2=0
cc_1025 N_A_1643_257#_c_1213_n N_A_1997_82#_c_1951_n 0.0140865f $X=12.66
+ $Y=1.215 $X2=0 $Y2=0
cc_1026 N_A_1643_257#_c_1214_n N_A_1997_82#_c_1951_n 8.91042e-19 $X=12.66
+ $Y=1.385 $X2=0 $Y2=0
cc_1027 N_A_1643_257#_c_1201_n N_A_1997_82#_c_1940_n 0.0012269f $X=12.705
+ $Y=1.795 $X2=0 $Y2=0
cc_1028 N_A_1643_257#_c_1208_n N_A_1997_82#_c_1940_n 0.0246745f $X=13.605
+ $Y=1.215 $X2=0 $Y2=0
cc_1029 N_A_1643_257#_c_1209_n N_A_1997_82#_c_1940_n 0.024772f $X=13.69 $Y=2.005
+ $X2=0 $Y2=0
cc_1030 N_A_1643_257#_c_1213_n N_A_1997_82#_c_1940_n 0.00506988f $X=12.66
+ $Y=1.215 $X2=0 $Y2=0
cc_1031 N_A_1643_257#_c_1214_n N_A_1997_82#_c_1940_n 2.78633e-19 $X=12.66
+ $Y=1.385 $X2=0 $Y2=0
cc_1032 N_A_1643_257#_c_1209_n N_RESET_B_c_2095_n 0.00648351f $X=13.69 $Y=2.005
+ $X2=-0.19 $Y2=-0.245
cc_1033 N_A_1643_257#_c_1210_n N_RESET_B_c_2095_n 0.00437319f $X=13.985 $Y=1.17
+ $X2=-0.19 $Y2=-0.245
cc_1034 N_A_1643_257#_c_1223_n N_RESET_B_c_2095_n 0.00784604f $X=13.91 $Y=2.17
+ $X2=-0.19 $Y2=-0.245
cc_1035 N_A_1643_257#_c_1209_n N_RESET_B_M1005_g 0.00477786f $X=13.69 $Y=2.005
+ $X2=0 $Y2=0
cc_1036 N_A_1643_257#_c_1210_n N_RESET_B_M1005_g 0.00589306f $X=13.985 $Y=1.17
+ $X2=0 $Y2=0
cc_1037 N_A_1643_257#_c_1209_n RESET_B 0.0247729f $X=13.69 $Y=2.005 $X2=0 $Y2=0
cc_1038 N_A_1643_257#_c_1210_n RESET_B 0.0161212f $X=13.985 $Y=1.17 $X2=0 $Y2=0
cc_1039 N_A_1643_257#_c_1223_n RESET_B 0.00772923f $X=13.91 $Y=2.17 $X2=0 $Y2=0
cc_1040 N_A_1643_257#_c_1217_n N_VPWR_c_2240_n 0.0127047f $X=8.305 $Y=2.045
+ $X2=0 $Y2=0
cc_1041 N_A_1643_257#_c_1219_n N_VPWR_c_2243_n 0.00968828f $X=12.705 $Y=1.885
+ $X2=0 $Y2=0
cc_1042 N_A_1643_257#_c_1217_n N_VPWR_c_2258_n 0.00413917f $X=8.305 $Y=2.045
+ $X2=0 $Y2=0
cc_1043 N_A_1643_257#_c_1219_n N_VPWR_c_2268_n 0.00444681f $X=12.705 $Y=1.885
+ $X2=0 $Y2=0
cc_1044 N_A_1643_257#_c_1217_n N_VPWR_c_2234_n 0.00817532f $X=8.305 $Y=2.045
+ $X2=0 $Y2=0
cc_1045 N_A_1643_257#_c_1219_n N_VPWR_c_2234_n 0.00877522f $X=12.705 $Y=1.885
+ $X2=0 $Y2=0
cc_1046 N_A_1643_257#_c_1204_n N_VGND_M1047_d 0.00250873f $X=9.555 $Y=1.195
+ $X2=0 $Y2=0
cc_1047 N_A_1643_257#_c_1301_p N_VGND_M1044_d 0.00967028f $X=11.895 $Y=0.685
+ $X2=0 $Y2=0
cc_1048 N_A_1643_257#_c_1255_n N_VGND_M1044_d 0.00817844f $X=11.98 $Y=0.685
+ $X2=0 $Y2=0
cc_1049 N_A_1643_257#_c_1204_n N_VGND_c_2737_n 0.0193447f $X=9.555 $Y=1.195
+ $X2=0 $Y2=0
cc_1050 N_A_1643_257#_c_1205_n N_VGND_c_2737_n 0.0266667f $X=9.64 $Y=1.11 $X2=0
+ $Y2=0
cc_1051 N_A_1643_257#_c_1207_n N_VGND_c_2737_n 0.0150383f $X=9.725 $Y=0.345
+ $X2=0 $Y2=0
cc_1052 N_A_1643_257#_c_1206_n N_VGND_c_2738_n 0.125559f $X=11.34 $Y=0.345 $X2=0
+ $Y2=0
cc_1053 N_A_1643_257#_c_1207_n N_VGND_c_2738_n 0.011809f $X=9.725 $Y=0.345 $X2=0
+ $Y2=0
cc_1054 N_A_1643_257#_c_1301_p N_VGND_c_2738_n 0.0186762f $X=11.895 $Y=0.685
+ $X2=0 $Y2=0
cc_1055 N_A_1643_257#_c_1255_n N_VGND_c_2738_n 0.0124527f $X=11.98 $Y=0.685
+ $X2=0 $Y2=0
cc_1056 N_A_1643_257#_c_1216_n N_VGND_c_2746_n 0.00279469f $X=12.66 $Y=1.22
+ $X2=0 $Y2=0
cc_1057 N_A_1643_257#_c_1206_n N_VGND_c_2759_n 0.0659229f $X=11.34 $Y=0.345
+ $X2=0 $Y2=0
cc_1058 N_A_1643_257#_c_1207_n N_VGND_c_2759_n 0.00591594f $X=9.725 $Y=0.345
+ $X2=0 $Y2=0
cc_1059 N_A_1643_257#_c_1301_p N_VGND_c_2759_n 0.00593218f $X=11.895 $Y=0.685
+ $X2=0 $Y2=0
cc_1060 N_A_1643_257#_c_1277_p N_VGND_c_2759_n 0.0061479f $X=12.495 $Y=0.855
+ $X2=0 $Y2=0
cc_1061 N_A_1643_257#_c_1255_n N_VGND_c_2759_n 0.001121f $X=11.98 $Y=0.685 $X2=0
+ $Y2=0
cc_1062 N_A_1643_257#_c_1216_n N_VGND_c_2759_n 0.00353488f $X=12.66 $Y=1.22
+ $X2=0 $Y2=0
cc_1063 N_A_1643_257#_c_1204_n N_A_1473_73#_M1018_d 0.00196293f $X=9.555
+ $Y=1.195 $X2=0 $Y2=0
cc_1064 N_A_1643_257#_c_1211_n N_A_1473_73#_M1018_d 0.001763f $X=8.38 $Y=1.45
+ $X2=0 $Y2=0
cc_1065 N_A_1643_257#_c_1202_n N_A_1473_73#_c_2925_n 0.00330783f $X=8.38
+ $Y=1.285 $X2=0 $Y2=0
cc_1066 N_A_1643_257#_c_1202_n N_A_1473_73#_c_2926_n 0.0028994f $X=8.38 $Y=1.285
+ $X2=0 $Y2=0
cc_1067 N_A_1643_257#_c_1202_n N_A_1473_73#_c_2928_n 0.00219422f $X=8.38
+ $Y=1.285 $X2=0 $Y2=0
cc_1068 N_A_1643_257#_c_1204_n N_A_1473_73#_c_2928_n 0.0141554f $X=9.555
+ $Y=1.195 $X2=0 $Y2=0
cc_1069 N_A_1643_257#_c_1211_n N_A_1473_73#_c_2928_n 0.0122474f $X=8.38 $Y=1.45
+ $X2=0 $Y2=0
cc_1070 N_A_1643_257#_c_1212_n N_A_1473_73#_c_2928_n 4.37138e-19 $X=8.38 $Y=1.45
+ $X2=0 $Y2=0
cc_1071 N_A_1643_257#_c_1204_n A_1902_125# 9.86779e-19 $X=9.555 $Y=1.195
+ $X2=-0.19 $Y2=-0.245
cc_1072 N_A_1643_257#_c_1205_n A_1902_125# 0.0109374f $X=9.64 $Y=1.11 $X2=-0.19
+ $Y2=-0.245
cc_1073 N_A_1643_257#_c_1206_n A_1902_125# 0.00198409f $X=11.34 $Y=0.345
+ $X2=-0.19 $Y2=-0.245
cc_1074 N_A_1643_257#_c_1206_n A_2247_82# 8.57957e-19 $X=11.34 $Y=0.345
+ $X2=-0.19 $Y2=-0.245
cc_1075 N_A_1643_257#_c_1251_n A_2247_82# 0.00187849f $X=11.425 $Y=0.6 $X2=-0.19
+ $Y2=-0.245
cc_1076 N_A_1643_257#_c_1252_n A_2247_82# 0.00241035f $X=11.51 $Y=0.685
+ $X2=-0.19 $Y2=-0.245
cc_1077 N_A_1643_257#_c_1277_p N_A_2452_74#_M1002_d 0.00826983f $X=12.495
+ $Y=0.855 $X2=-0.19 $Y2=-0.245
cc_1078 N_A_1643_257#_c_1291_p N_A_2452_74#_M1002_d 0.00205664f $X=12.66 $Y=1.13
+ $X2=-0.19 $Y2=-0.245
cc_1079 N_A_1643_257#_c_1277_p N_A_2452_74#_c_2972_n 0.0232142f $X=12.495
+ $Y=0.855 $X2=0 $Y2=0
cc_1080 N_A_1643_257#_c_1214_n N_A_2452_74#_c_2972_n 3.37831e-19 $X=12.66
+ $Y=1.385 $X2=0 $Y2=0
cc_1081 N_A_1643_257#_c_1216_n N_A_2452_74#_c_2972_n 0.00618812f $X=12.66
+ $Y=1.22 $X2=0 $Y2=0
cc_1082 N_A_1643_257#_c_1277_p N_A_2452_74#_c_2974_n 3.69705e-19 $X=12.495
+ $Y=0.855 $X2=0 $Y2=0
cc_1083 N_A_1643_257#_c_1216_n N_A_2452_74#_c_2974_n 0.0103546f $X=12.66 $Y=1.22
+ $X2=0 $Y2=0
cc_1084 N_SET_B_M1047_g N_A_688_98#_c_1550_n 0.00894519f $X=8.935 $Y=0.9 $X2=0
+ $Y2=0
cc_1085 N_SET_B_c_1408_n N_A_688_98#_c_1555_n 0.00646001f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_1086 N_SET_B_c_1418_n N_A_2216_410#_c_1742_n 0.00161456f $X=12.195 $Y=1.885
+ $X2=0 $Y2=0
cc_1087 N_SET_B_c_1414_n N_A_2216_410#_c_1727_n 0.0113438f $X=12.12 $Y=1.22
+ $X2=0 $Y2=0
cc_1088 N_SET_B_c_1407_n N_A_2216_410#_c_1728_n 0.0108751f $X=12.195 $Y=1.795
+ $X2=0 $Y2=0
cc_1089 N_SET_B_c_1418_n N_A_2216_410#_c_1728_n 0.0109889f $X=12.195 $Y=1.885
+ $X2=0 $Y2=0
cc_1090 N_SET_B_c_1408_n N_A_2216_410#_c_1728_n 0.00208814f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_1091 N_SET_B_c_1412_n N_A_2216_410#_c_1728_n 0.0190514f $X=12.12 $Y=1.385
+ $X2=0 $Y2=0
cc_1092 N_SET_B_c_1413_n N_A_2216_410#_c_1728_n 0.00245434f $X=12.12 $Y=1.385
+ $X2=0 $Y2=0
cc_1093 N_SET_B_c_1414_n N_A_2216_410#_c_1736_n 0.0104689f $X=12.12 $Y=1.22
+ $X2=0 $Y2=0
cc_1094 N_SET_B_c_1408_n N_A_2216_410#_c_1749_n 0.00125344f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_1095 N_SET_B_c_1418_n N_A_2216_410#_c_1769_n 0.0120695f $X=12.195 $Y=1.885
+ $X2=0 $Y2=0
cc_1096 N_SET_B_c_1418_n N_A_2216_410#_c_1754_n 0.0077283f $X=12.195 $Y=1.885
+ $X2=0 $Y2=0
cc_1097 N_SET_B_c_1408_n N_A_1997_82#_c_1944_n 0.0208248f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_1098 N_SET_B_c_1408_n N_A_1997_82#_c_1945_n 0.00477725f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_1099 N_SET_B_c_1408_n N_A_1997_82#_c_1937_n 0.00414645f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_1100 N_SET_B_c_1414_n N_A_1997_82#_c_1937_n 9.54794e-19 $X=12.12 $Y=1.22
+ $X2=0 $Y2=0
cc_1101 N_SET_B_c_1407_n N_A_1997_82#_c_1938_n 2.65996e-19 $X=12.195 $Y=1.795
+ $X2=0 $Y2=0
cc_1102 N_SET_B_c_1408_n N_A_1997_82#_c_1938_n 0.02011f $X=12.095 $Y=1.665 $X2=0
+ $Y2=0
cc_1103 SET_B N_A_1997_82#_c_1938_n 2.92235e-19 $X=12.155 $Y=1.58 $X2=0 $Y2=0
cc_1104 N_SET_B_c_1412_n N_A_1997_82#_c_1938_n 0.00111915f $X=12.12 $Y=1.385
+ $X2=0 $Y2=0
cc_1105 N_SET_B_c_1413_n N_A_1997_82#_c_1938_n 0.0314411f $X=12.12 $Y=1.385
+ $X2=0 $Y2=0
cc_1106 N_SET_B_c_1414_n N_A_1997_82#_c_1938_n 4.36939e-19 $X=12.12 $Y=1.22
+ $X2=0 $Y2=0
cc_1107 N_SET_B_c_1418_n N_A_1997_82#_c_1947_n 0.0115755f $X=12.195 $Y=1.885
+ $X2=0 $Y2=0
cc_1108 N_SET_B_c_1408_n N_A_1997_82#_c_1947_n 0.0102273f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_1109 SET_B N_A_1997_82#_c_1947_n 0.00873829f $X=12.155 $Y=1.58 $X2=0 $Y2=0
cc_1110 N_SET_B_c_1412_n N_A_1997_82#_c_1947_n 6.5626e-19 $X=12.12 $Y=1.385
+ $X2=0 $Y2=0
cc_1111 N_SET_B_c_1413_n N_A_1997_82#_c_1947_n 0.0248499f $X=12.12 $Y=1.385
+ $X2=0 $Y2=0
cc_1112 N_SET_B_c_1408_n N_A_1997_82#_c_1949_n 0.00714641f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_1113 N_SET_B_c_1407_n N_A_1997_82#_c_1950_n 0.0030679f $X=12.195 $Y=1.795
+ $X2=0 $Y2=0
cc_1114 N_SET_B_c_1418_n N_A_1997_82#_c_1950_n 7.86492e-19 $X=12.195 $Y=1.885
+ $X2=0 $Y2=0
cc_1115 N_SET_B_c_1408_n N_A_1997_82#_c_1950_n 0.00127856f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_1116 SET_B N_A_1997_82#_c_1950_n 0.00141707f $X=12.155 $Y=1.58 $X2=0 $Y2=0
cc_1117 N_SET_B_c_1407_n N_A_1997_82#_c_1951_n 0.0028047f $X=12.195 $Y=1.795
+ $X2=0 $Y2=0
cc_1118 N_SET_B_c_1418_n N_A_1997_82#_c_1951_n 8.87563e-19 $X=12.195 $Y=1.885
+ $X2=0 $Y2=0
cc_1119 SET_B N_A_1997_82#_c_1951_n 0.00254814f $X=12.155 $Y=1.58 $X2=0 $Y2=0
cc_1120 N_SET_B_c_1413_n N_A_1997_82#_c_1951_n 0.00197725f $X=12.12 $Y=1.385
+ $X2=0 $Y2=0
cc_1121 N_SET_B_c_1416_n N_VPWR_c_2240_n 0.00773228f $X=8.845 $Y=2.045 $X2=0
+ $Y2=0
cc_1122 N_SET_B_c_1416_n N_VPWR_c_2241_n 0.00427151f $X=8.845 $Y=2.045 $X2=0
+ $Y2=0
cc_1123 N_SET_B_c_1408_n N_VPWR_c_2241_n 9.40915e-19 $X=12.095 $Y=1.665 $X2=0
+ $Y2=0
cc_1124 N_SET_B_c_1418_n N_VPWR_c_2242_n 0.00337783f $X=12.195 $Y=1.885 $X2=0
+ $Y2=0
cc_1125 N_SET_B_c_1418_n N_VPWR_c_2243_n 0.00528294f $X=12.195 $Y=1.885 $X2=0
+ $Y2=0
cc_1126 N_SET_B_c_1416_n N_VPWR_c_2249_n 0.00445602f $X=8.845 $Y=2.045 $X2=0
+ $Y2=0
cc_1127 N_SET_B_c_1418_n N_VPWR_c_2251_n 0.00445602f $X=12.195 $Y=1.885 $X2=0
+ $Y2=0
cc_1128 N_SET_B_c_1416_n N_VPWR_c_2234_n 0.00863447f $X=8.845 $Y=2.045 $X2=0
+ $Y2=0
cc_1129 N_SET_B_c_1418_n N_VPWR_c_2234_n 0.00862315f $X=12.195 $Y=1.885 $X2=0
+ $Y2=0
cc_1130 N_SET_B_M1047_g N_VGND_c_2737_n 0.00322717f $X=8.935 $Y=0.9 $X2=0 $Y2=0
cc_1131 N_SET_B_c_1414_n N_VGND_c_2738_n 0.00248478f $X=12.12 $Y=1.22 $X2=0
+ $Y2=0
cc_1132 N_SET_B_c_1414_n N_VGND_c_2746_n 0.0043213f $X=12.12 $Y=1.22 $X2=0 $Y2=0
cc_1133 N_SET_B_M1047_g N_VGND_c_2759_n 9.49986e-19 $X=8.935 $Y=0.9 $X2=0 $Y2=0
cc_1134 N_SET_B_c_1414_n N_VGND_c_2759_n 0.0043699f $X=12.12 $Y=1.22 $X2=0 $Y2=0
cc_1135 N_SET_B_M1047_g N_A_1473_73#_c_2926_n 9.77356e-19 $X=8.935 $Y=0.9 $X2=0
+ $Y2=0
cc_1136 N_SET_B_M1047_g N_A_1473_73#_c_2928_n 0.00432596f $X=8.935 $Y=0.9 $X2=0
+ $Y2=0
cc_1137 N_SET_B_c_1414_n N_A_2452_74#_c_2972_n 0.00767947f $X=12.12 $Y=1.22
+ $X2=0 $Y2=0
cc_1138 N_A_688_98#_c_1562_n N_A_2216_410#_c_1742_n 0.0260087f $X=10.78 $Y=2.085
+ $X2=0 $Y2=0
cc_1139 N_A_688_98#_c_1564_n N_A_2216_410#_c_1742_n 0.0320085f $X=10.78 $Y=2.465
+ $X2=0 $Y2=0
cc_1140 N_A_688_98#_c_1563_n N_A_2216_410#_c_1753_n 8.04528e-19 $X=10.78
+ $Y=2.375 $X2=0 $Y2=0
cc_1141 N_A_688_98#_c_1563_n N_A_1997_82#_c_1942_n 0.00308241f $X=10.78 $Y=2.375
+ $X2=0 $Y2=0
cc_1142 N_A_688_98#_c_1564_n N_A_1997_82#_c_1942_n 0.00927397f $X=10.78 $Y=2.465
+ $X2=0 $Y2=0
cc_1143 N_A_688_98#_c_1562_n N_A_1997_82#_c_1943_n 0.00378556f $X=10.78 $Y=2.085
+ $X2=0 $Y2=0
cc_1144 N_A_688_98#_c_1563_n N_A_1997_82#_c_1943_n 8.5016e-19 $X=10.78 $Y=2.375
+ $X2=0 $Y2=0
cc_1145 N_A_688_98#_c_1555_n N_A_1997_82#_c_1943_n 0.00289557f $X=10.78 $Y=1.995
+ $X2=0 $Y2=0
cc_1146 N_A_688_98#_c_1555_n N_A_1997_82#_c_1945_n 0.0100134f $X=10.78 $Y=1.995
+ $X2=0 $Y2=0
cc_1147 N_A_688_98#_c_1563_n N_A_1997_82#_c_1949_n 0.0151046f $X=10.78 $Y=2.375
+ $X2=0 $Y2=0
cc_1148 N_A_688_98#_M1020_g N_A_1997_82#_c_1939_n 0.00368644f $X=9.91 $Y=0.685
+ $X2=0 $Y2=0
cc_1149 N_A_688_98#_c_1552_n N_A_1997_82#_c_1939_n 0.0225496f $X=10.695 $Y=1.11
+ $X2=0 $Y2=0
cc_1150 N_A_688_98#_c_1586_n N_VPWR_M1036_d 0.00644937f $X=4.065 $Y=2.035 $X2=0
+ $Y2=0
cc_1151 N_A_688_98#_c_1569_n N_VPWR_M1036_d 0.00126846f $X=4.15 $Y=1.95 $X2=0
+ $Y2=0
cc_1152 N_A_688_98#_c_1560_n N_VPWR_c_2237_n 0.0140621f $X=4.265 $Y=1.765 $X2=0
+ $Y2=0
cc_1153 N_A_688_98#_c_1568_n N_VPWR_c_2237_n 0.0462948f $X=3.59 $Y=2.815 $X2=0
+ $Y2=0
cc_1154 N_A_688_98#_c_1586_n N_VPWR_c_2237_n 0.0178169f $X=4.065 $Y=2.035 $X2=0
+ $Y2=0
cc_1155 N_A_688_98#_c_1560_n N_VPWR_c_2238_n 0.00413917f $X=4.265 $Y=1.765 $X2=0
+ $Y2=0
cc_1156 N_A_688_98#_c_1560_n N_VPWR_c_2239_n 0.00311538f $X=4.265 $Y=1.765 $X2=0
+ $Y2=0
cc_1157 N_A_688_98#_c_1564_n N_VPWR_c_2242_n 0.0016566f $X=10.78 $Y=2.465 $X2=0
+ $Y2=0
cc_1158 N_A_688_98#_c_1568_n N_VPWR_c_2257_n 0.011066f $X=3.59 $Y=2.815 $X2=0
+ $Y2=0
cc_1159 N_A_688_98#_c_1565_n N_VPWR_c_2258_n 0.00278271f $X=6.227 $Y=2.245 $X2=0
+ $Y2=0
cc_1160 N_A_688_98#_c_1564_n N_VPWR_c_2259_n 0.00461464f $X=10.78 $Y=2.465 $X2=0
+ $Y2=0
cc_1161 N_A_688_98#_c_1560_n N_VPWR_c_2234_n 0.00822528f $X=4.265 $Y=1.765 $X2=0
+ $Y2=0
cc_1162 N_A_688_98#_c_1564_n N_VPWR_c_2234_n 0.00982378f $X=10.78 $Y=2.465 $X2=0
+ $Y2=0
cc_1163 N_A_688_98#_c_1565_n N_VPWR_c_2234_n 0.00363426f $X=6.227 $Y=2.245 $X2=0
+ $Y2=0
cc_1164 N_A_688_98#_c_1568_n N_VPWR_c_2234_n 0.00915947f $X=3.59 $Y=2.815 $X2=0
+ $Y2=0
cc_1165 N_A_688_98#_M1035_s N_A_197_119#_c_2454_n 0.00286661f $X=3.44 $Y=0.49
+ $X2=0 $Y2=0
cc_1166 N_A_688_98#_M1035_s N_A_197_119#_c_2546_n 0.00373877f $X=3.44 $Y=0.49
+ $X2=0 $Y2=0
cc_1167 N_A_688_98#_c_1556_n N_A_197_119#_c_2546_n 0.0432119f $X=4.065 $Y=1.085
+ $X2=0 $Y2=0
cc_1168 N_A_688_98#_c_1557_n N_A_197_119#_c_2546_n 0.00684564f $X=4.28 $Y=1.505
+ $X2=0 $Y2=0
cc_1169 N_A_688_98#_c_1558_n N_A_197_119#_c_2546_n 0.00372791f $X=4.28 $Y=1.505
+ $X2=0 $Y2=0
cc_1170 N_A_688_98#_M1035_s N_A_197_119#_c_2455_n 0.00193137f $X=3.44 $Y=0.49
+ $X2=0 $Y2=0
cc_1171 N_A_688_98#_c_1556_n N_A_197_119#_c_2455_n 0.0092465f $X=4.065 $Y=1.085
+ $X2=0 $Y2=0
cc_1172 N_A_688_98#_M1043_g N_A_197_119#_c_2456_n 0.00261388f $X=4.64 $Y=0.86
+ $X2=0 $Y2=0
cc_1173 N_A_688_98#_M1043_g N_A_197_119#_c_2457_n 0.0163579f $X=4.64 $Y=0.86
+ $X2=0 $Y2=0
cc_1174 N_A_688_98#_c_1547_n N_A_197_119#_c_2457_n 0.0113624f $X=6.135 $Y=0.18
+ $X2=0 $Y2=0
cc_1175 N_A_688_98#_M1043_g N_A_197_119#_c_2459_n 0.00259659f $X=4.64 $Y=0.86
+ $X2=0 $Y2=0
cc_1176 N_A_688_98#_c_1547_n N_A_197_119#_c_2460_n 0.00511412f $X=6.135 $Y=0.18
+ $X2=0 $Y2=0
cc_1177 N_A_688_98#_M1016_g N_A_197_119#_c_2462_n 0.0040541f $X=6.21 $Y=0.835
+ $X2=0 $Y2=0
cc_1178 N_A_688_98#_M1016_g N_A_197_119#_c_2463_n 0.0174699f $X=6.21 $Y=0.835
+ $X2=0 $Y2=0
cc_1179 N_A_688_98#_c_1550_n N_A_197_119#_c_2463_n 0.015287f $X=9.835 $Y=0.18
+ $X2=0 $Y2=0
cc_1180 N_A_688_98#_c_1547_n N_A_197_119#_c_2464_n 0.00246334f $X=6.135 $Y=0.18
+ $X2=0 $Y2=0
cc_1181 N_A_688_98#_M1016_g N_A_197_119#_c_2465_n 0.00121318f $X=6.21 $Y=0.835
+ $X2=0 $Y2=0
cc_1182 N_A_688_98#_c_1550_n N_A_197_119#_c_2466_n 0.00529214f $X=9.835 $Y=0.18
+ $X2=0 $Y2=0
cc_1183 N_A_688_98#_c_1556_n N_VGND_M1035_d 0.0123255f $X=4.065 $Y=1.085 $X2=0
+ $Y2=0
cc_1184 N_A_688_98#_c_1559_n N_VGND_M1035_d 0.00144075f $X=4.255 $Y=1.34 $X2=0
+ $Y2=0
cc_1185 N_A_688_98#_M1043_g N_VGND_c_2735_n 7.43091e-19 $X=4.64 $Y=0.86 $X2=0
+ $Y2=0
cc_1186 N_A_688_98#_c_1548_n N_VGND_c_2735_n 0.00328096f $X=4.715 $Y=0.18 $X2=0
+ $Y2=0
cc_1187 N_A_688_98#_c_1547_n N_VGND_c_2736_n 0.0221124f $X=6.135 $Y=0.18 $X2=0
+ $Y2=0
cc_1188 N_A_688_98#_M1016_g N_VGND_c_2736_n 0.0012066f $X=6.21 $Y=0.835 $X2=0
+ $Y2=0
cc_1189 N_A_688_98#_c_1550_n N_VGND_c_2737_n 0.0256092f $X=9.835 $Y=0.18 $X2=0
+ $Y2=0
cc_1190 N_A_688_98#_M1020_g N_VGND_c_2737_n 9.32533e-19 $X=9.91 $Y=0.685 $X2=0
+ $Y2=0
cc_1191 N_A_688_98#_c_1550_n N_VGND_c_2738_n 0.0155404f $X=9.835 $Y=0.18 $X2=0
+ $Y2=0
cc_1192 N_A_688_98#_c_1548_n N_VGND_c_2751_n 0.0212479f $X=4.715 $Y=0.18 $X2=0
+ $Y2=0
cc_1193 N_A_688_98#_c_1547_n N_VGND_c_2752_n 0.0792334f $X=6.135 $Y=0.18 $X2=0
+ $Y2=0
cc_1194 N_A_688_98#_c_1547_n N_VGND_c_2759_n 0.0289617f $X=6.135 $Y=0.18 $X2=0
+ $Y2=0
cc_1195 N_A_688_98#_c_1548_n N_VGND_c_2759_n 0.00604517f $X=4.715 $Y=0.18 $X2=0
+ $Y2=0
cc_1196 N_A_688_98#_c_1550_n N_VGND_c_2759_n 0.0882651f $X=9.835 $Y=0.18 $X2=0
+ $Y2=0
cc_1197 N_A_688_98#_c_1554_n N_VGND_c_2759_n 0.00371014f $X=6.21 $Y=0.18 $X2=0
+ $Y2=0
cc_1198 N_A_688_98#_c_1550_n N_A_1473_73#_c_2925_n 0.0151187f $X=9.835 $Y=0.18
+ $X2=0 $Y2=0
cc_1199 N_A_688_98#_c_1550_n N_A_1473_73#_c_2927_n 0.0101915f $X=9.835 $Y=0.18
+ $X2=0 $Y2=0
cc_1200 N_A_688_98#_c_1550_n N_A_1473_73#_c_2928_n 0.00461421f $X=9.835 $Y=0.18
+ $X2=0 $Y2=0
cc_1201 N_A_2216_410#_c_1769_n N_A_1997_82#_c_1935_n 0.0131714f $X=13.185
+ $Y=2.345 $X2=0 $Y2=0
cc_1202 N_A_2216_410#_c_1750_n N_A_1997_82#_c_1935_n 0.00568183f $X=13.35
+ $Y=2.815 $X2=0 $Y2=0
cc_1203 N_A_2216_410#_c_1751_n N_A_1997_82#_c_1935_n 4.68534e-19 $X=14.485
+ $Y=2.59 $X2=0 $Y2=0
cc_1204 N_A_2216_410#_c_1778_n N_A_1997_82#_c_1935_n 0.013096f $X=13.35 $Y=2.225
+ $X2=0 $Y2=0
cc_1205 N_A_2216_410#_c_1737_n N_A_1997_82#_M1007_g 0.00945324f $X=14.32 $Y=0.75
+ $X2=0 $Y2=0
cc_1206 N_A_2216_410#_c_1777_n N_A_1997_82#_M1007_g 0.00919204f $X=13.085
+ $Y=0.777 $X2=0 $Y2=0
cc_1207 N_A_2216_410#_c_1753_n N_A_1997_82#_c_1942_n 0.00615248f $X=11.245
+ $Y=2.215 $X2=0 $Y2=0
cc_1208 N_A_2216_410#_c_1742_n N_A_1997_82#_c_1943_n 4.87001e-19 $X=11.17
+ $Y=2.465 $X2=0 $Y2=0
cc_1209 N_A_2216_410#_c_1728_n N_A_1997_82#_c_1943_n 6.12047e-19 $X=11.67
+ $Y=2.05 $X2=0 $Y2=0
cc_1210 N_A_2216_410#_c_1753_n N_A_1997_82#_c_1943_n 7.51566e-19 $X=11.245
+ $Y=2.215 $X2=0 $Y2=0
cc_1211 N_A_2216_410#_c_1742_n N_A_1997_82#_c_1944_n 0.00672329f $X=11.17
+ $Y=2.465 $X2=0 $Y2=0
cc_1212 N_A_2216_410#_c_1736_n N_A_1997_82#_c_1944_n 3.69566e-19 $X=11.67
+ $Y=0.98 $X2=0 $Y2=0
cc_1213 N_A_2216_410#_c_1749_n N_A_1997_82#_c_1944_n 0.00586426f $X=11.805
+ $Y=2.345 $X2=0 $Y2=0
cc_1214 N_A_2216_410#_c_1753_n N_A_1997_82#_c_1944_n 0.0233976f $X=11.245
+ $Y=2.215 $X2=0 $Y2=0
cc_1215 N_A_2216_410#_c_1728_n N_A_1997_82#_c_1937_n 0.00229815f $X=11.67
+ $Y=2.05 $X2=0 $Y2=0
cc_1216 N_A_2216_410#_c_1736_n N_A_1997_82#_c_1937_n 0.0106122f $X=11.67 $Y=0.98
+ $X2=0 $Y2=0
cc_1217 N_A_2216_410#_c_1728_n N_A_1997_82#_c_1938_n 0.0156997f $X=11.67 $Y=2.05
+ $X2=0 $Y2=0
cc_1218 N_A_2216_410#_M1011_s N_A_1997_82#_c_1947_n 0.00263709f $X=11.825
+ $Y=1.96 $X2=0 $Y2=0
cc_1219 N_A_2216_410#_c_1749_n N_A_1997_82#_c_1947_n 0.00393489f $X=11.805
+ $Y=2.345 $X2=0 $Y2=0
cc_1220 N_A_2216_410#_c_1769_n N_A_1997_82#_c_1947_n 0.0208133f $X=13.185
+ $Y=2.345 $X2=0 $Y2=0
cc_1221 N_A_2216_410#_c_1754_n N_A_1997_82#_c_1947_n 0.0214641f $X=11.97
+ $Y=2.425 $X2=0 $Y2=0
cc_1222 N_A_2216_410#_c_1769_n N_A_1997_82#_c_1948_n 0.0129802f $X=13.185
+ $Y=2.345 $X2=0 $Y2=0
cc_1223 N_A_2216_410#_c_1742_n N_A_1997_82#_c_1949_n 0.00106329f $X=11.17
+ $Y=2.465 $X2=0 $Y2=0
cc_1224 N_A_2216_410#_c_1753_n N_A_1997_82#_c_1949_n 0.0140315f $X=11.245
+ $Y=2.215 $X2=0 $Y2=0
cc_1225 N_A_2216_410#_c_1727_n N_A_1997_82#_c_1939_n 0.00101133f $X=11.55
+ $Y=0.905 $X2=0 $Y2=0
cc_1226 N_A_2216_410#_c_1743_n N_A_1997_82#_c_1950_n 0.00449844f $X=11.595
+ $Y=2.125 $X2=0 $Y2=0
cc_1227 N_A_2216_410#_c_1728_n N_A_1997_82#_c_1950_n 0.01315f $X=11.67 $Y=2.05
+ $X2=0 $Y2=0
cc_1228 N_A_2216_410#_c_1749_n N_A_1997_82#_c_1950_n 0.014174f $X=11.805
+ $Y=2.345 $X2=0 $Y2=0
cc_1229 N_A_2216_410#_c_1769_n N_A_1997_82#_c_1951_n 0.00842961f $X=13.185
+ $Y=2.345 $X2=0 $Y2=0
cc_1230 N_A_2216_410#_c_1778_n N_A_1997_82#_c_1951_n 8.39722e-19 $X=13.35
+ $Y=2.225 $X2=0 $Y2=0
cc_1231 N_A_2216_410#_c_1769_n N_A_1997_82#_c_1940_n 0.00563106f $X=13.185
+ $Y=2.345 $X2=0 $Y2=0
cc_1232 N_A_2216_410#_c_1778_n N_A_1997_82#_c_1940_n 0.0130707f $X=13.35
+ $Y=2.225 $X2=0 $Y2=0
cc_1233 N_A_2216_410#_c_1751_n N_RESET_B_c_2095_n 0.017337f $X=14.485 $Y=2.59
+ $X2=-0.19 $Y2=-0.245
cc_1234 N_A_2216_410#_c_1752_n N_RESET_B_c_2095_n 0.0172709f $X=14.57 $Y=2.505
+ $X2=-0.19 $Y2=-0.245
cc_1235 N_A_2216_410#_c_1778_n N_RESET_B_c_2095_n 0.00586581f $X=13.35 $Y=2.225
+ $X2=-0.19 $Y2=-0.245
cc_1236 N_A_2216_410#_c_1739_n N_RESET_B_c_2095_n 3.20825e-19 $X=14.65 $Y=1.595
+ $X2=-0.19 $Y2=-0.245
cc_1237 N_A_2216_410#_c_1737_n N_RESET_B_M1005_g 0.0098987f $X=14.32 $Y=0.75
+ $X2=0 $Y2=0
cc_1238 N_A_2216_410#_c_1738_n N_RESET_B_M1005_g 0.00478654f $X=14.57 $Y=1.005
+ $X2=0 $Y2=0
cc_1239 N_A_2216_410#_c_1739_n N_RESET_B_M1005_g 5.04769e-19 $X=14.65 $Y=1.595
+ $X2=0 $Y2=0
cc_1240 N_A_2216_410#_c_1740_n N_RESET_B_M1005_g 0.00967958f $X=14.65 $Y=1.43
+ $X2=0 $Y2=0
cc_1241 N_A_2216_410#_c_1741_n N_RESET_B_M1005_g 0.0217165f $X=14.65 $Y=1.537
+ $X2=0 $Y2=0
cc_1242 N_A_2216_410#_c_1737_n RESET_B 0.00272307f $X=14.32 $Y=0.75 $X2=0 $Y2=0
cc_1243 N_A_2216_410#_c_1751_n RESET_B 0.00394184f $X=14.485 $Y=2.59 $X2=0 $Y2=0
cc_1244 N_A_2216_410#_c_1739_n RESET_B 0.0208985f $X=14.65 $Y=1.595 $X2=0 $Y2=0
cc_1245 N_A_2216_410#_c_1741_n RESET_B 9.6319e-19 $X=14.65 $Y=1.537 $X2=0 $Y2=0
cc_1246 N_A_2216_410#_c_1735_n N_A_3272_94#_c_2133_n 0.0177582f $X=16.76
+ $Y=1.845 $X2=0 $Y2=0
cc_1247 N_A_2216_410#_M1019_g N_A_3272_94#_c_2127_n 0.0168621f $X=16.72 $Y=0.79
+ $X2=0 $Y2=0
cc_1248 N_A_2216_410#_M1021_g N_A_3272_94#_c_2129_n 0.00302515f $X=15.66 $Y=0.74
+ $X2=0 $Y2=0
cc_1249 N_A_2216_410#_M1019_g N_A_3272_94#_c_2129_n 0.0117319f $X=16.72 $Y=0.79
+ $X2=0 $Y2=0
cc_1250 N_A_2216_410#_c_1746_n N_A_3272_94#_c_2135_n 0.00438746f $X=15.765
+ $Y=1.765 $X2=0 $Y2=0
cc_1251 N_A_2216_410#_c_1732_n N_A_3272_94#_c_2135_n 0.0128835f $X=16.645
+ $Y=1.497 $X2=0 $Y2=0
cc_1252 N_A_2216_410#_c_1733_n N_A_3272_94#_c_2135_n 0.00207643f $X=15.855
+ $Y=1.497 $X2=0 $Y2=0
cc_1253 N_A_2216_410#_c_1735_n N_A_3272_94#_c_2135_n 0.0243353f $X=16.76
+ $Y=1.845 $X2=0 $Y2=0
cc_1254 N_A_2216_410#_M1019_g N_A_3272_94#_c_2130_n 0.00692483f $X=16.72 $Y=0.79
+ $X2=0 $Y2=0
cc_1255 N_A_2216_410#_c_1735_n N_A_3272_94#_c_2130_n 0.0116748f $X=16.76
+ $Y=1.845 $X2=0 $Y2=0
cc_1256 N_A_2216_410#_M1021_g N_A_3272_94#_c_2131_n 0.00339198f $X=15.66 $Y=0.74
+ $X2=0 $Y2=0
cc_1257 N_A_2216_410#_c_1732_n N_A_3272_94#_c_2131_n 0.0213836f $X=16.645
+ $Y=1.497 $X2=0 $Y2=0
cc_1258 N_A_2216_410#_M1019_g N_A_3272_94#_c_2131_n 0.0048318f $X=16.72 $Y=0.79
+ $X2=0 $Y2=0
cc_1259 N_A_2216_410#_c_1735_n N_A_3272_94#_c_2131_n 0.00103581f $X=16.76
+ $Y=1.845 $X2=0 $Y2=0
cc_1260 N_A_2216_410#_M1019_g N_A_3272_94#_c_2132_n 0.00713437f $X=16.72 $Y=0.79
+ $X2=0 $Y2=0
cc_1261 N_A_2216_410#_c_1735_n N_A_3272_94#_c_2132_n 0.0210248f $X=16.76
+ $Y=1.845 $X2=0 $Y2=0
cc_1262 N_A_2216_410#_c_1769_n N_VPWR_M1011_d 0.0051977f $X=13.185 $Y=2.345
+ $X2=0 $Y2=0
cc_1263 N_A_2216_410#_c_1751_n N_VPWR_M1026_d 0.0160022f $X=14.485 $Y=2.59 $X2=0
+ $Y2=0
cc_1264 N_A_2216_410#_c_1752_n N_VPWR_M1026_d 0.0160868f $X=14.57 $Y=2.505 $X2=0
+ $Y2=0
cc_1265 N_A_2216_410#_c_1742_n N_VPWR_c_2242_n 0.0125837f $X=11.17 $Y=2.465
+ $X2=0 $Y2=0
cc_1266 N_A_2216_410#_c_1749_n N_VPWR_c_2242_n 0.0123543f $X=11.805 $Y=2.345
+ $X2=0 $Y2=0
cc_1267 N_A_2216_410#_c_1753_n N_VPWR_c_2242_n 0.0127679f $X=11.245 $Y=2.215
+ $X2=0 $Y2=0
cc_1268 N_A_2216_410#_c_1754_n N_VPWR_c_2242_n 0.0245258f $X=11.97 $Y=2.425
+ $X2=0 $Y2=0
cc_1269 N_A_2216_410#_c_1769_n N_VPWR_c_2243_n 0.0201954f $X=13.185 $Y=2.345
+ $X2=0 $Y2=0
cc_1270 N_A_2216_410#_c_1754_n N_VPWR_c_2243_n 0.015049f $X=11.97 $Y=2.425 $X2=0
+ $Y2=0
cc_1271 N_A_2216_410#_c_1778_n N_VPWR_c_2243_n 0.0106303f $X=13.35 $Y=2.225
+ $X2=0 $Y2=0
cc_1272 N_A_2216_410#_c_1729_n N_VPWR_c_2244_n 0.0126913f $X=15.155 $Y=1.537
+ $X2=0 $Y2=0
cc_1273 N_A_2216_410#_c_1745_n N_VPWR_c_2244_n 0.0202255f $X=15.315 $Y=1.765
+ $X2=0 $Y2=0
cc_1274 N_A_2216_410#_c_1751_n N_VPWR_c_2244_n 0.0145234f $X=14.485 $Y=2.59
+ $X2=0 $Y2=0
cc_1275 N_A_2216_410#_c_1752_n N_VPWR_c_2244_n 0.0426554f $X=14.57 $Y=2.505
+ $X2=0 $Y2=0
cc_1276 N_A_2216_410#_c_1745_n N_VPWR_c_2245_n 6.81303e-19 $X=15.315 $Y=1.765
+ $X2=0 $Y2=0
cc_1277 N_A_2216_410#_c_1746_n N_VPWR_c_2245_n 0.0160518f $X=15.765 $Y=1.765
+ $X2=0 $Y2=0
cc_1278 N_A_2216_410#_c_1732_n N_VPWR_c_2245_n 0.0104745f $X=16.645 $Y=1.497
+ $X2=0 $Y2=0
cc_1279 N_A_2216_410#_c_1735_n N_VPWR_c_2245_n 0.0042597f $X=16.76 $Y=1.845
+ $X2=0 $Y2=0
cc_1280 N_A_2216_410#_c_1735_n N_VPWR_c_2246_n 0.0131658f $X=16.76 $Y=1.845
+ $X2=0 $Y2=0
cc_1281 N_A_2216_410#_c_1754_n N_VPWR_c_2251_n 0.0146549f $X=11.97 $Y=2.425
+ $X2=0 $Y2=0
cc_1282 N_A_2216_410#_c_1745_n N_VPWR_c_2253_n 0.00445602f $X=15.315 $Y=1.765
+ $X2=0 $Y2=0
cc_1283 N_A_2216_410#_c_1746_n N_VPWR_c_2253_n 0.00413917f $X=15.765 $Y=1.765
+ $X2=0 $Y2=0
cc_1284 N_A_2216_410#_c_1742_n N_VPWR_c_2259_n 0.00413917f $X=11.17 $Y=2.465
+ $X2=0 $Y2=0
cc_1285 N_A_2216_410#_c_1735_n N_VPWR_c_2260_n 0.00534256f $X=16.76 $Y=1.845
+ $X2=0 $Y2=0
cc_1286 N_A_2216_410#_c_1750_n N_VPWR_c_2268_n 0.0110241f $X=13.35 $Y=2.815
+ $X2=0 $Y2=0
cc_1287 N_A_2216_410#_c_1751_n N_VPWR_c_2268_n 0.0144354f $X=14.485 $Y=2.59
+ $X2=0 $Y2=0
cc_1288 N_A_2216_410#_c_1745_n N_VPWR_c_2269_n 0.00646036f $X=15.315 $Y=1.765
+ $X2=0 $Y2=0
cc_1289 N_A_2216_410#_c_1751_n N_VPWR_c_2269_n 0.0299125f $X=14.485 $Y=2.59
+ $X2=0 $Y2=0
cc_1290 N_A_2216_410#_c_1742_n N_VPWR_c_2234_n 0.00851932f $X=11.17 $Y=2.465
+ $X2=0 $Y2=0
cc_1291 N_A_2216_410#_c_1745_n N_VPWR_c_2234_n 0.00862481f $X=15.315 $Y=1.765
+ $X2=0 $Y2=0
cc_1292 N_A_2216_410#_c_1746_n N_VPWR_c_2234_n 0.00817726f $X=15.765 $Y=1.765
+ $X2=0 $Y2=0
cc_1293 N_A_2216_410#_c_1735_n N_VPWR_c_2234_n 0.00533081f $X=16.76 $Y=1.845
+ $X2=0 $Y2=0
cc_1294 N_A_2216_410#_c_1750_n N_VPWR_c_2234_n 0.00909194f $X=13.35 $Y=2.815
+ $X2=0 $Y2=0
cc_1295 N_A_2216_410#_c_1751_n N_VPWR_c_2234_n 0.0253264f $X=14.485 $Y=2.59
+ $X2=0 $Y2=0
cc_1296 N_A_2216_410#_c_1754_n N_VPWR_c_2234_n 0.0120704f $X=11.97 $Y=2.425
+ $X2=0 $Y2=0
cc_1297 N_A_2216_410#_c_1769_n A_2556_392# 0.00835497f $X=13.185 $Y=2.345
+ $X2=-0.19 $Y2=-0.245
cc_1298 N_A_2216_410#_M1003_g N_Q_N_c_2675_n 0.00868707f $X=15.23 $Y=0.74 $X2=0
+ $Y2=0
cc_1299 N_A_2216_410#_M1021_g N_Q_N_c_2675_n 0.00868707f $X=15.66 $Y=0.74 $X2=0
+ $Y2=0
cc_1300 N_A_2216_410#_c_1745_n N_Q_N_c_2678_n 0.0195341f $X=15.315 $Y=1.765
+ $X2=0 $Y2=0
cc_1301 N_A_2216_410#_c_1746_n N_Q_N_c_2678_n 0.00771123f $X=15.765 $Y=1.765
+ $X2=0 $Y2=0
cc_1302 N_A_2216_410#_M1003_g N_Q_N_c_2676_n 0.00528879f $X=15.23 $Y=0.74 $X2=0
+ $Y2=0
cc_1303 N_A_2216_410#_M1021_g N_Q_N_c_2676_n 0.00601183f $X=15.66 $Y=0.74 $X2=0
+ $Y2=0
cc_1304 N_A_2216_410#_c_1740_n N_Q_N_c_2676_n 0.00251143f $X=14.65 $Y=1.43 $X2=0
+ $Y2=0
cc_1305 N_A_2216_410#_c_1745_n Q_N 7.57488e-19 $X=15.315 $Y=1.765 $X2=0 $Y2=0
cc_1306 N_A_2216_410#_c_1746_n Q_N 0.00157942f $X=15.765 $Y=1.765 $X2=0 $Y2=0
cc_1307 N_A_2216_410#_c_1733_n Q_N 0.0281842f $X=15.855 $Y=1.497 $X2=0 $Y2=0
cc_1308 N_A_2216_410#_c_1741_n Q_N 3.87333e-19 $X=14.65 $Y=1.537 $X2=0 $Y2=0
cc_1309 N_A_2216_410#_M1003_g N_Q_N_c_2677_n 0.00321384f $X=15.23 $Y=0.74 $X2=0
+ $Y2=0
cc_1310 N_A_2216_410#_M1021_g N_Q_N_c_2677_n 0.0064747f $X=15.66 $Y=0.74 $X2=0
+ $Y2=0
cc_1311 N_A_2216_410#_c_1733_n N_Q_N_c_2677_n 0.0223956f $X=15.855 $Y=1.497
+ $X2=0 $Y2=0
cc_1312 N_A_2216_410#_c_1739_n N_Q_N_c_2677_n 0.00920625f $X=14.65 $Y=1.595
+ $X2=0 $Y2=0
cc_1313 N_A_2216_410#_c_1738_n N_VGND_M1005_d 0.00852738f $X=14.57 $Y=1.005
+ $X2=0 $Y2=0
cc_1314 N_A_2216_410#_c_1740_n N_VGND_M1005_d 0.0057756f $X=14.65 $Y=1.43 $X2=0
+ $Y2=0
cc_1315 N_A_2216_410#_c_1727_n N_VGND_c_2738_n 0.00484024f $X=11.55 $Y=0.905
+ $X2=0 $Y2=0
cc_1316 N_A_2216_410#_c_1729_n N_VGND_c_2739_n 0.0104813f $X=15.155 $Y=1.537
+ $X2=0 $Y2=0
cc_1317 N_A_2216_410#_M1003_g N_VGND_c_2739_n 0.00527975f $X=15.23 $Y=0.74 $X2=0
+ $Y2=0
cc_1318 N_A_2216_410#_c_1738_n N_VGND_c_2739_n 0.0230527f $X=14.57 $Y=1.005
+ $X2=0 $Y2=0
cc_1319 N_A_2216_410#_c_1740_n N_VGND_c_2739_n 0.00946423f $X=14.65 $Y=1.43
+ $X2=0 $Y2=0
cc_1320 N_A_2216_410#_M1021_g N_VGND_c_2740_n 0.00532106f $X=15.66 $Y=0.74 $X2=0
+ $Y2=0
cc_1321 N_A_2216_410#_c_1733_n N_VGND_c_2740_n 0.0118899f $X=15.855 $Y=1.497
+ $X2=0 $Y2=0
cc_1322 N_A_2216_410#_M1019_g N_VGND_c_2740_n 0.00532677f $X=16.72 $Y=0.79 $X2=0
+ $Y2=0
cc_1323 N_A_2216_410#_M1019_g N_VGND_c_2741_n 0.0106131f $X=16.72 $Y=0.79 $X2=0
+ $Y2=0
cc_1324 N_A_2216_410#_c_1737_n N_VGND_c_2746_n 0.0125015f $X=14.32 $Y=0.75 $X2=0
+ $Y2=0
cc_1325 N_A_2216_410#_c_1738_n N_VGND_c_2746_n 0.00307629f $X=14.57 $Y=1.005
+ $X2=0 $Y2=0
cc_1326 N_A_2216_410#_M1003_g N_VGND_c_2748_n 0.00434272f $X=15.23 $Y=0.74 $X2=0
+ $Y2=0
cc_1327 N_A_2216_410#_M1021_g N_VGND_c_2748_n 0.00434272f $X=15.66 $Y=0.74 $X2=0
+ $Y2=0
cc_1328 N_A_2216_410#_M1019_g N_VGND_c_2753_n 0.00486866f $X=16.72 $Y=0.79 $X2=0
+ $Y2=0
cc_1329 N_A_2216_410#_c_1727_n N_VGND_c_2759_n 0.00408695f $X=11.55 $Y=0.905
+ $X2=0 $Y2=0
cc_1330 N_A_2216_410#_M1003_g N_VGND_c_2759_n 0.00825059f $X=15.23 $Y=0.74 $X2=0
+ $Y2=0
cc_1331 N_A_2216_410#_M1021_g N_VGND_c_2759_n 0.00825059f $X=15.66 $Y=0.74 $X2=0
+ $Y2=0
cc_1332 N_A_2216_410#_M1019_g N_VGND_c_2759_n 0.00514438f $X=16.72 $Y=0.79 $X2=0
+ $Y2=0
cc_1333 N_A_2216_410#_c_1737_n N_VGND_c_2759_n 0.0213693f $X=14.32 $Y=0.75 $X2=0
+ $Y2=0
cc_1334 N_A_2216_410#_c_1738_n N_VGND_c_2759_n 0.0114279f $X=14.57 $Y=1.005
+ $X2=0 $Y2=0
cc_1335 N_A_2216_410#_c_1737_n N_A_2452_74#_M1007_d 0.00899529f $X=14.32 $Y=0.75
+ $X2=0 $Y2=0
cc_1336 N_A_2216_410#_c_1727_n N_A_2452_74#_c_2972_n 7.73746e-19 $X=11.55
+ $Y=0.905 $X2=0 $Y2=0
cc_1337 N_A_2216_410#_c_1737_n N_A_2452_74#_c_2973_n 0.023391f $X=14.32 $Y=0.75
+ $X2=0 $Y2=0
cc_1338 N_A_2216_410#_M1038_d N_A_2452_74#_c_2974_n 0.00176891f $X=12.78 $Y=0.37
+ $X2=0 $Y2=0
cc_1339 N_A_2216_410#_c_1737_n N_A_2452_74#_c_2974_n 0.00605639f $X=14.32
+ $Y=0.75 $X2=0 $Y2=0
cc_1340 N_A_2216_410#_c_1777_n N_A_2452_74#_c_2974_n 0.0136435f $X=13.085
+ $Y=0.777 $X2=0 $Y2=0
cc_1341 N_A_1997_82#_c_1935_n N_RESET_B_c_2095_n 0.00421082f $X=13.125 $Y=1.885
+ $X2=-0.19 $Y2=-0.245
cc_1342 N_A_1997_82#_c_1947_n N_VPWR_M1011_d 0.00209889f $X=12.495 $Y=2.005
+ $X2=0 $Y2=0
cc_1343 N_A_1997_82#_c_1951_n N_VPWR_M1011_d 0.00115596f $X=12.58 $Y=1.805 $X2=0
+ $Y2=0
cc_1344 N_A_1997_82#_c_1942_n N_VPWR_c_2241_n 0.0211074f $X=10.47 $Y=2.815 $X2=0
+ $Y2=0
cc_1345 N_A_1997_82#_c_1942_n N_VPWR_c_2242_n 0.0110165f $X=10.47 $Y=2.815 $X2=0
+ $Y2=0
cc_1346 N_A_1997_82#_c_1935_n N_VPWR_c_2243_n 0.00161227f $X=13.125 $Y=1.885
+ $X2=0 $Y2=0
cc_1347 N_A_1997_82#_c_1942_n N_VPWR_c_2259_n 0.0146399f $X=10.47 $Y=2.815 $X2=0
+ $Y2=0
cc_1348 N_A_1997_82#_c_1935_n N_VPWR_c_2268_n 0.00445602f $X=13.125 $Y=1.885
+ $X2=0 $Y2=0
cc_1349 N_A_1997_82#_c_1935_n N_VPWR_c_2234_n 0.00862959f $X=13.125 $Y=1.885
+ $X2=0 $Y2=0
cc_1350 N_A_1997_82#_c_1942_n N_VPWR_c_2234_n 0.0120646f $X=10.47 $Y=2.815 $X2=0
+ $Y2=0
cc_1351 N_A_1997_82#_M1007_g N_VGND_c_2746_n 0.00278271f $X=13.135 $Y=0.74 $X2=0
+ $Y2=0
cc_1352 N_A_1997_82#_M1007_g N_VGND_c_2759_n 0.00358525f $X=13.135 $Y=0.74 $X2=0
+ $Y2=0
cc_1353 N_A_1997_82#_M1007_g N_A_2452_74#_c_2972_n 7.51897e-19 $X=13.135 $Y=0.74
+ $X2=0 $Y2=0
cc_1354 N_A_1997_82#_M1007_g N_A_2452_74#_c_2974_n 0.0110587f $X=13.135 $Y=0.74
+ $X2=0 $Y2=0
cc_1355 N_RESET_B_c_2095_n N_VPWR_c_2244_n 0.0032988f $X=14.135 $Y=1.92 $X2=0
+ $Y2=0
cc_1356 N_RESET_B_c_2095_n N_VPWR_c_2268_n 0.00296344f $X=14.135 $Y=1.92 $X2=0
+ $Y2=0
cc_1357 N_RESET_B_c_2095_n N_VPWR_c_2234_n 0.0045051f $X=14.135 $Y=1.92 $X2=0
+ $Y2=0
cc_1358 N_RESET_B_M1005_g N_VGND_c_2739_n 6.60505e-19 $X=14.2 $Y=1.11 $X2=0
+ $Y2=0
cc_1359 N_RESET_B_M1005_g N_VGND_c_2746_n 4.65242e-19 $X=14.2 $Y=1.11 $X2=0
+ $Y2=0
cc_1360 N_A_3272_94#_c_2135_n N_VPWR_c_2245_n 0.0781858f $X=16.535 $Y=2.065
+ $X2=0 $Y2=0
cc_1361 N_A_3272_94#_c_2133_n N_VPWR_c_2246_n 0.0158737f $X=17.285 $Y=1.765
+ $X2=0 $Y2=0
cc_1362 N_A_3272_94#_c_2134_n N_VPWR_c_2246_n 6.79664e-19 $X=17.735 $Y=1.765
+ $X2=0 $Y2=0
cc_1363 N_A_3272_94#_c_2135_n N_VPWR_c_2246_n 0.0788767f $X=16.535 $Y=2.065
+ $X2=0 $Y2=0
cc_1364 N_A_3272_94#_c_2130_n N_VPWR_c_2246_n 0.0201266f $X=17.2 $Y=1.385 $X2=0
+ $Y2=0
cc_1365 N_A_3272_94#_c_2132_n N_VPWR_c_2246_n 0.00399876f $X=17.735 $Y=1.492
+ $X2=0 $Y2=0
cc_1366 N_A_3272_94#_c_2134_n N_VPWR_c_2248_n 0.0082329f $X=17.735 $Y=1.765
+ $X2=0 $Y2=0
cc_1367 N_A_3272_94#_c_2135_n N_VPWR_c_2260_n 0.0137187f $X=16.535 $Y=2.065
+ $X2=0 $Y2=0
cc_1368 N_A_3272_94#_c_2133_n N_VPWR_c_2261_n 0.00413917f $X=17.285 $Y=1.765
+ $X2=0 $Y2=0
cc_1369 N_A_3272_94#_c_2134_n N_VPWR_c_2261_n 0.00411612f $X=17.735 $Y=1.765
+ $X2=0 $Y2=0
cc_1370 N_A_3272_94#_c_2133_n N_VPWR_c_2234_n 0.00817726f $X=17.285 $Y=1.765
+ $X2=0 $Y2=0
cc_1371 N_A_3272_94#_c_2134_n N_VPWR_c_2234_n 0.00751023f $X=17.735 $Y=1.765
+ $X2=0 $Y2=0
cc_1372 N_A_3272_94#_c_2135_n N_VPWR_c_2234_n 0.0128859f $X=16.535 $Y=2.065
+ $X2=0 $Y2=0
cc_1373 N_A_3272_94#_c_2135_n Q_N 0.00643638f $X=16.535 $Y=2.065 $X2=0 $Y2=0
cc_1374 N_A_3272_94#_c_2127_n N_Q_c_2705_n 0.00597104f $X=17.32 $Y=1.22 $X2=0
+ $Y2=0
cc_1375 N_A_3272_94#_c_2128_n N_Q_c_2705_n 0.00643254f $X=17.75 $Y=1.22 $X2=0
+ $Y2=0
cc_1376 N_A_3272_94#_c_2127_n N_Q_c_2712_n 0.00292633f $X=17.32 $Y=1.22 $X2=0
+ $Y2=0
cc_1377 N_A_3272_94#_c_2128_n N_Q_c_2712_n 0.00185771f $X=17.75 $Y=1.22 $X2=0
+ $Y2=0
cc_1378 N_A_3272_94#_c_2132_n N_Q_c_2712_n 0.00221432f $X=17.735 $Y=1.492 $X2=0
+ $Y2=0
cc_1379 N_A_3272_94#_c_2133_n Q 5.45961e-19 $X=17.285 $Y=1.765 $X2=0 $Y2=0
cc_1380 N_A_3272_94#_c_2134_n Q 0.00205881f $X=17.735 $Y=1.765 $X2=0 $Y2=0
cc_1381 N_A_3272_94#_c_2132_n Q 0.00286568f $X=17.735 $Y=1.492 $X2=0 $Y2=0
cc_1382 N_A_3272_94#_c_2134_n Q 0.0132088f $X=17.735 $Y=1.765 $X2=0 $Y2=0
cc_1383 N_A_3272_94#_c_2127_n N_Q_c_2706_n 0.00257108f $X=17.32 $Y=1.22 $X2=0
+ $Y2=0
cc_1384 N_A_3272_94#_c_2134_n N_Q_c_2706_n 0.0030228f $X=17.735 $Y=1.765 $X2=0
+ $Y2=0
cc_1385 N_A_3272_94#_c_2128_n N_Q_c_2706_n 0.0056016f $X=17.75 $Y=1.22 $X2=0
+ $Y2=0
cc_1386 N_A_3272_94#_c_2130_n N_Q_c_2706_n 0.0249855f $X=17.2 $Y=1.385 $X2=0
+ $Y2=0
cc_1387 N_A_3272_94#_c_2132_n N_Q_c_2706_n 0.0395125f $X=17.735 $Y=1.492 $X2=0
+ $Y2=0
cc_1388 N_A_3272_94#_c_2129_n N_VGND_c_2740_n 0.0397772f $X=16.505 $Y=0.645
+ $X2=0 $Y2=0
cc_1389 N_A_3272_94#_c_2127_n N_VGND_c_2741_n 0.00907221f $X=17.32 $Y=1.22 $X2=0
+ $Y2=0
cc_1390 N_A_3272_94#_c_2129_n N_VGND_c_2741_n 0.0349326f $X=16.505 $Y=0.645
+ $X2=0 $Y2=0
cc_1391 N_A_3272_94#_c_2130_n N_VGND_c_2741_n 0.0272668f $X=17.2 $Y=1.385 $X2=0
+ $Y2=0
cc_1392 N_A_3272_94#_c_2132_n N_VGND_c_2741_n 0.00379679f $X=17.735 $Y=1.492
+ $X2=0 $Y2=0
cc_1393 N_A_3272_94#_c_2128_n N_VGND_c_2743_n 0.00647103f $X=17.75 $Y=1.22 $X2=0
+ $Y2=0
cc_1394 N_A_3272_94#_c_2129_n N_VGND_c_2753_n 0.00720482f $X=16.505 $Y=0.645
+ $X2=0 $Y2=0
cc_1395 N_A_3272_94#_c_2127_n N_VGND_c_2754_n 0.00434272f $X=17.32 $Y=1.22 $X2=0
+ $Y2=0
cc_1396 N_A_3272_94#_c_2128_n N_VGND_c_2754_n 0.00428607f $X=17.75 $Y=1.22 $X2=0
+ $Y2=0
cc_1397 N_A_3272_94#_c_2127_n N_VGND_c_2759_n 0.00825059f $X=17.32 $Y=1.22 $X2=0
+ $Y2=0
cc_1398 N_A_3272_94#_c_2128_n N_VGND_c_2759_n 0.00805581f $X=17.75 $Y=1.22 $X2=0
+ $Y2=0
cc_1399 N_A_3272_94#_c_2129_n N_VGND_c_2759_n 0.010626f $X=16.505 $Y=0.645 $X2=0
+ $Y2=0
cc_1400 N_A_27_464#_c_2193_n N_VPWR_M1028_d 0.00195252f $X=1.065 $Y=2.39
+ $X2=-0.19 $Y2=1.66
cc_1401 N_A_27_464#_c_2193_n N_VPWR_c_2235_n 0.0168243f $X=1.065 $Y=2.39 $X2=0
+ $Y2=0
cc_1402 N_A_27_464#_c_2195_n N_VPWR_c_2235_n 0.0117237f $X=1.235 $Y=2.99 $X2=0
+ $Y2=0
cc_1403 N_A_27_464#_c_2197_n N_VPWR_c_2235_n 0.0224916f $X=0.28 $Y=2.47 $X2=0
+ $Y2=0
cc_1404 N_A_27_464#_c_2194_n N_VPWR_c_2236_n 0.0121617f $X=1.855 $Y=2.99 $X2=0
+ $Y2=0
cc_1405 N_A_27_464#_c_2196_n N_VPWR_c_2236_n 0.0407546f $X=2.02 $Y=2.465 $X2=0
+ $Y2=0
cc_1406 N_A_27_464#_c_2197_n N_VPWR_c_2255_n 0.01106f $X=0.28 $Y=2.47 $X2=0
+ $Y2=0
cc_1407 N_A_27_464#_c_2194_n N_VPWR_c_2256_n 0.0626582f $X=1.855 $Y=2.99 $X2=0
+ $Y2=0
cc_1408 N_A_27_464#_c_2195_n N_VPWR_c_2256_n 0.0121867f $X=1.235 $Y=2.99 $X2=0
+ $Y2=0
cc_1409 N_A_27_464#_c_2193_n N_VPWR_c_2234_n 0.0117086f $X=1.065 $Y=2.39 $X2=0
+ $Y2=0
cc_1410 N_A_27_464#_c_2194_n N_VPWR_c_2234_n 0.0347672f $X=1.855 $Y=2.99 $X2=0
+ $Y2=0
cc_1411 N_A_27_464#_c_2195_n N_VPWR_c_2234_n 0.00660921f $X=1.235 $Y=2.99 $X2=0
+ $Y2=0
cc_1412 N_A_27_464#_c_2197_n N_VPWR_c_2234_n 0.00915715f $X=0.28 $Y=2.47 $X2=0
+ $Y2=0
cc_1413 N_A_27_464#_c_2228_p A_206_464# 5.61252e-19 $X=1.15 $Y=2.905 $X2=-0.19
+ $Y2=1.66
cc_1414 N_A_27_464#_c_2194_n N_A_197_119#_M1000_d 0.00222494f $X=1.855 $Y=2.99
+ $X2=0 $Y2=0
cc_1415 N_A_27_464#_c_2193_n N_A_197_119#_c_2470_n 0.00675867f $X=1.065 $Y=2.39
+ $X2=0 $Y2=0
cc_1416 N_A_27_464#_c_2196_n N_A_197_119#_c_2470_n 0.0291626f $X=2.02 $Y=2.465
+ $X2=0 $Y2=0
cc_1417 N_A_27_464#_c_2194_n N_A_197_119#_c_2481_n 0.014415f $X=1.855 $Y=2.99
+ $X2=0 $Y2=0
cc_1418 N_A_27_464#_c_2196_n N_A_197_119#_c_2471_n 0.0253885f $X=2.02 $Y=2.465
+ $X2=0 $Y2=0
cc_1419 N_VPWR_c_2244_n N_Q_N_c_2678_n 0.059157f $X=15.005 $Y=2.15 $X2=0 $Y2=0
cc_1420 N_VPWR_c_2245_n N_Q_N_c_2678_n 0.0690922f $X=15.99 $Y=2.115 $X2=0 $Y2=0
cc_1421 N_VPWR_c_2253_n N_Q_N_c_2678_n 0.0110241f $X=15.825 $Y=3.33 $X2=0 $Y2=0
cc_1422 N_VPWR_c_2269_n N_Q_N_c_2678_n 0.00943121f $X=15.17 $Y=3.13 $X2=0 $Y2=0
cc_1423 N_VPWR_c_2234_n N_Q_N_c_2678_n 0.00909194f $X=18 $Y=3.33 $X2=0 $Y2=0
cc_1424 N_VPWR_c_2246_n Q 0.045092f $X=17.06 $Y=2.045 $X2=0 $Y2=0
cc_1425 N_VPWR_c_2248_n Q 0.0877598f $X=17.96 $Y=1.985 $X2=0 $Y2=0
cc_1426 N_VPWR_c_2261_n Q 0.0136117f $X=17.875 $Y=3.33 $X2=0 $Y2=0
cc_1427 N_VPWR_c_2234_n Q 0.0111632f $X=18 $Y=3.33 $X2=0 $Y2=0
cc_1428 N_A_197_119#_c_2451_n N_VGND_M1025_d 0.00415254f $X=2.685 $Y=1.12 $X2=0
+ $Y2=0
cc_1429 N_A_197_119#_c_2546_n N_VGND_M1035_d 0.017252f $X=4.35 $Y=0.745 $X2=0
+ $Y2=0
cc_1430 N_A_197_119#_c_2456_n N_VGND_M1035_d 0.00323892f $X=4.435 $Y=0.66 $X2=0
+ $Y2=0
cc_1431 N_A_197_119#_c_2460_n N_VGND_M1027_s 0.00757503f $X=5.945 $Y=0.925 $X2=0
+ $Y2=0
cc_1432 N_A_197_119#_c_2478_n N_VGND_c_2733_n 0.0110205f $X=1.525 $Y=0.79 $X2=0
+ $Y2=0
cc_1433 N_A_197_119#_c_2482_n N_VGND_c_2734_n 0.0107049f $X=1.587 $Y=0.955 $X2=0
+ $Y2=0
cc_1434 N_A_197_119#_c_2450_n N_VGND_c_2734_n 0.0177503f $X=2.6 $Y=1.205 $X2=0
+ $Y2=0
cc_1435 N_A_197_119#_c_2451_n N_VGND_c_2734_n 0.0396995f $X=2.685 $Y=1.12 $X2=0
+ $Y2=0
cc_1436 N_A_197_119#_c_2453_n N_VGND_c_2734_n 0.0147449f $X=2.77 $Y=0.34 $X2=0
+ $Y2=0
cc_1437 N_A_197_119#_c_2452_n N_VGND_c_2735_n 0.00820222f $X=3.365 $Y=0.34 $X2=0
+ $Y2=0
cc_1438 N_A_197_119#_c_2454_n N_VGND_c_2735_n 0.00278228f $X=3.45 $Y=0.66 $X2=0
+ $Y2=0
cc_1439 N_A_197_119#_c_2546_n N_VGND_c_2735_n 0.0190193f $X=4.35 $Y=0.745 $X2=0
+ $Y2=0
cc_1440 N_A_197_119#_c_2456_n N_VGND_c_2735_n 0.00491052f $X=4.435 $Y=0.66 $X2=0
+ $Y2=0
cc_1441 N_A_197_119#_c_2458_n N_VGND_c_2735_n 0.0145006f $X=4.52 $Y=0.34 $X2=0
+ $Y2=0
cc_1442 N_A_197_119#_c_2457_n N_VGND_c_2736_n 0.0147306f $X=5.11 $Y=0.34 $X2=0
+ $Y2=0
cc_1443 N_A_197_119#_c_2459_n N_VGND_c_2736_n 0.0187223f $X=5.195 $Y=0.84 $X2=0
+ $Y2=0
cc_1444 N_A_197_119#_c_2460_n N_VGND_c_2736_n 0.0212468f $X=5.945 $Y=0.925 $X2=0
+ $Y2=0
cc_1445 N_A_197_119#_c_2462_n N_VGND_c_2736_n 0.0120826f $X=6.03 $Y=0.84 $X2=0
+ $Y2=0
cc_1446 N_A_197_119#_c_2464_n N_VGND_c_2736_n 0.012174f $X=6.115 $Y=0.35 $X2=0
+ $Y2=0
cc_1447 N_A_197_119#_c_2482_n N_VGND_c_2744_n 0.00344134f $X=1.587 $Y=0.955
+ $X2=0 $Y2=0
cc_1448 N_A_197_119#_c_2478_n N_VGND_c_2744_n 0.00925972f $X=1.525 $Y=0.79 $X2=0
+ $Y2=0
cc_1449 N_A_197_119#_c_2452_n N_VGND_c_2750_n 0.0499722f $X=3.365 $Y=0.34 $X2=0
+ $Y2=0
cc_1450 N_A_197_119#_c_2453_n N_VGND_c_2750_n 0.0115566f $X=2.77 $Y=0.34 $X2=0
+ $Y2=0
cc_1451 N_A_197_119#_c_2546_n N_VGND_c_2750_n 0.00552268f $X=4.35 $Y=0.745 $X2=0
+ $Y2=0
cc_1452 N_A_197_119#_c_2546_n N_VGND_c_2751_n 0.00279509f $X=4.35 $Y=0.745 $X2=0
+ $Y2=0
cc_1453 N_A_197_119#_c_2457_n N_VGND_c_2751_n 0.0490946f $X=5.11 $Y=0.34 $X2=0
+ $Y2=0
cc_1454 N_A_197_119#_c_2458_n N_VGND_c_2751_n 0.0120335f $X=4.52 $Y=0.34 $X2=0
+ $Y2=0
cc_1455 N_A_197_119#_c_2463_n N_VGND_c_2752_n 0.0623722f $X=6.785 $Y=0.35 $X2=0
+ $Y2=0
cc_1456 N_A_197_119#_c_2464_n N_VGND_c_2752_n 0.0114593f $X=6.115 $Y=0.35 $X2=0
+ $Y2=0
cc_1457 N_A_197_119#_c_2482_n N_VGND_c_2759_n 0.00540954f $X=1.587 $Y=0.955
+ $X2=0 $Y2=0
cc_1458 N_A_197_119#_c_2452_n N_VGND_c_2759_n 0.0284203f $X=3.365 $Y=0.34 $X2=0
+ $Y2=0
cc_1459 N_A_197_119#_c_2453_n N_VGND_c_2759_n 0.00579705f $X=2.77 $Y=0.34 $X2=0
+ $Y2=0
cc_1460 N_A_197_119#_c_2546_n N_VGND_c_2759_n 0.0168022f $X=4.35 $Y=0.745 $X2=0
+ $Y2=0
cc_1461 N_A_197_119#_c_2457_n N_VGND_c_2759_n 0.0257198f $X=5.11 $Y=0.34 $X2=0
+ $Y2=0
cc_1462 N_A_197_119#_c_2458_n N_VGND_c_2759_n 0.00658039f $X=4.52 $Y=0.34 $X2=0
+ $Y2=0
cc_1463 N_A_197_119#_c_2460_n N_VGND_c_2759_n 0.0125365f $X=5.945 $Y=0.925 $X2=0
+ $Y2=0
cc_1464 N_A_197_119#_c_2463_n N_VGND_c_2759_n 0.0336647f $X=6.785 $Y=0.35 $X2=0
+ $Y2=0
cc_1465 N_A_197_119#_c_2464_n N_VGND_c_2759_n 0.00589978f $X=6.115 $Y=0.35 $X2=0
+ $Y2=0
cc_1466 N_A_197_119#_c_2466_n N_VGND_c_2759_n 0.00732007f $X=7.535 $Y=0.93 $X2=0
+ $Y2=0
cc_1467 N_A_197_119#_c_2478_n N_VGND_c_2759_n 0.0133937f $X=1.525 $Y=0.79 $X2=0
+ $Y2=0
cc_1468 N_A_197_119#_c_2460_n A_1185_125# 9.645e-19 $X=5.945 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_1469 N_A_197_119#_c_2466_n N_A_1473_73#_M1017_s 0.00873925f $X=7.535 $Y=0.93
+ $X2=-0.19 $Y2=-0.245
cc_1470 N_A_197_119#_c_2468_n N_A_1473_73#_M1017_s 0.00816566f $X=7.62 $Y=2.38
+ $X2=-0.19 $Y2=-0.245
cc_1471 N_A_197_119#_c_2463_n N_A_1473_73#_c_2927_n 0.0123861f $X=6.785 $Y=0.35
+ $X2=0 $Y2=0
cc_1472 N_A_197_119#_c_2465_n N_A_1473_73#_c_2927_n 0.0164625f $X=6.95 $Y=0.81
+ $X2=0 $Y2=0
cc_1473 N_A_197_119#_c_2466_n N_A_1473_73#_c_2927_n 0.0279978f $X=7.535 $Y=0.93
+ $X2=0 $Y2=0
cc_1474 N_Q_N_c_2675_n N_VGND_c_2739_n 0.0307762f $X=15.445 $Y=0.515 $X2=0 $Y2=0
cc_1475 N_Q_N_c_2675_n N_VGND_c_2740_n 0.0308109f $X=15.445 $Y=0.515 $X2=0 $Y2=0
cc_1476 N_Q_N_c_2675_n N_VGND_c_2748_n 0.0144922f $X=15.445 $Y=0.515 $X2=0 $Y2=0
cc_1477 N_Q_N_c_2675_n N_VGND_c_2759_n 0.0118826f $X=15.445 $Y=0.515 $X2=0 $Y2=0
cc_1478 N_Q_c_2705_n N_VGND_c_2741_n 0.0270791f $X=17.535 $Y=0.515 $X2=0 $Y2=0
cc_1479 N_Q_c_2705_n N_VGND_c_2743_n 0.0301698f $X=17.535 $Y=0.515 $X2=0 $Y2=0
cc_1480 N_Q_c_2705_n N_VGND_c_2754_n 0.0147156f $X=17.535 $Y=0.515 $X2=0 $Y2=0
cc_1481 N_Q_c_2705_n N_VGND_c_2759_n 0.0120492f $X=17.535 $Y=0.515 $X2=0 $Y2=0
cc_1482 N_VGND_c_2737_n N_A_1473_73#_c_2925_n 0.00783795f $X=9.22 $Y=0.77 $X2=0
+ $Y2=0
cc_1483 N_VGND_c_2752_n N_A_1473_73#_c_2925_n 0.0520824f $X=9.055 $Y=0 $X2=0
+ $Y2=0
cc_1484 N_VGND_c_2759_n N_A_1473_73#_c_2925_n 0.0284814f $X=18 $Y=0 $X2=0 $Y2=0
cc_1485 N_VGND_c_2737_n N_A_1473_73#_c_2926_n 0.00699789f $X=9.22 $Y=0.77 $X2=0
+ $Y2=0
cc_1486 N_VGND_c_2752_n N_A_1473_73#_c_2927_n 0.0274584f $X=9.055 $Y=0 $X2=0
+ $Y2=0
cc_1487 N_VGND_c_2759_n N_A_1473_73#_c_2927_n 0.014464f $X=18 $Y=0 $X2=0 $Y2=0
cc_1488 N_VGND_c_2737_n N_A_1473_73#_c_2928_n 0.0136607f $X=9.22 $Y=0.77 $X2=0
+ $Y2=0
cc_1489 N_VGND_c_2752_n N_A_1473_73#_c_2928_n 0.00536382f $X=9.055 $Y=0 $X2=0
+ $Y2=0
cc_1490 N_VGND_c_2759_n N_A_1473_73#_c_2928_n 0.00689759f $X=18 $Y=0 $X2=0 $Y2=0
cc_1491 N_VGND_c_2738_n N_A_2452_74#_c_2972_n 0.0111522f $X=11.68 $Y=0 $X2=0
+ $Y2=0
cc_1492 N_VGND_c_2746_n N_A_2452_74#_c_2972_n 0.0283431f $X=14.825 $Y=0 $X2=0
+ $Y2=0
cc_1493 N_VGND_c_2759_n N_A_2452_74#_c_2972_n 0.0157587f $X=18 $Y=0 $X2=0 $Y2=0
cc_1494 N_VGND_c_2746_n N_A_2452_74#_c_2974_n 0.0602407f $X=14.825 $Y=0 $X2=0
+ $Y2=0
cc_1495 N_VGND_c_2759_n N_A_2452_74#_c_2974_n 0.0341799f $X=18 $Y=0 $X2=0 $Y2=0
