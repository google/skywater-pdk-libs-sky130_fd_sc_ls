* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__dfrbp_2 CLK D RESET_B VGND VNB VPB VPWR Q Q_N
X0 a_156_74# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_70_74# a_728_331# a_298_294# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_818_418# a_728_331# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X3 a_1800_291# a_1586_149# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 a_298_294# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 a_818_418# a_728_331# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X6 VPWR a_2363_352# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X7 VGND a_2363_352# Q VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X8 a_1586_149# a_818_418# a_331_392# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X9 VGND a_1586_149# a_2363_352# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X10 Q a_2363_352# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X11 a_1499_149# a_1800_291# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 VGND CLK a_728_331# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X13 VPWR a_1586_149# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X14 VGND RESET_B a_1974_74# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 a_1755_389# a_1800_291# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X16 VGND a_1586_149# Q_N VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X17 a_70_74# D a_156_74# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 Q_N a_1586_149# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X19 VPWR a_331_392# a_683_485# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X20 a_1586_149# a_818_418# a_1755_389# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X21 a_1974_74# a_1586_149# a_1800_291# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X22 a_298_294# a_818_418# a_70_74# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X23 VPWR CLK a_728_331# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X24 VPWR a_1586_149# a_2363_352# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X25 Q a_2363_352# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X26 VGND a_298_294# a_331_392# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X27 a_70_74# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X28 VPWR D a_70_74# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X29 a_298_294# a_818_418# a_614_81# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X30 VGND RESET_B a_536_81# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X31 Q_N a_1586_149# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X32 VPWR a_298_294# a_331_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X33 a_331_392# a_728_331# a_1586_149# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X34 a_536_81# a_331_392# a_614_81# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X35 VPWR RESET_B a_1800_291# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X36 a_1499_149# a_728_331# a_1586_149# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X37 a_683_485# a_728_331# a_298_294# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
.ends
