* File: sky130_fd_sc_ls__nor4bb_2.pxi.spice
* Created: Wed Sep  2 11:16:12 2020
* 
x_PM_SKY130_FD_SC_LS__NOR4BB_2%C_N N_C_N_c_110_n N_C_N_M1014_g N_C_N_M1016_g C_N
+ C_N N_C_N_c_109_n PM_SKY130_FD_SC_LS__NOR4BB_2%C_N
x_PM_SKY130_FD_SC_LS__NOR4BB_2%D_N N_D_N_c_140_n N_D_N_M1004_g N_D_N_c_143_n
+ N_D_N_M1012_g D_N N_D_N_c_142_n PM_SKY130_FD_SC_LS__NOR4BB_2%D_N
x_PM_SKY130_FD_SC_LS__NOR4BB_2%A_311_124# N_A_311_124#_M1004_d
+ N_A_311_124#_M1012_d N_A_311_124#_c_181_n N_A_311_124#_M1001_g
+ N_A_311_124#_M1000_g N_A_311_124#_M1010_g N_A_311_124#_c_182_n
+ N_A_311_124#_M1015_g N_A_311_124#_c_178_n N_A_311_124#_c_183_n
+ N_A_311_124#_c_202_p N_A_311_124#_c_184_n N_A_311_124#_c_185_n
+ N_A_311_124#_c_179_n N_A_311_124#_c_180_n
+ PM_SKY130_FD_SC_LS__NOR4BB_2%A_311_124#
x_PM_SKY130_FD_SC_LS__NOR4BB_2%A_27_392# N_A_27_392#_M1016_s N_A_27_392#_M1014_s
+ N_A_27_392#_c_265_n N_A_27_392#_M1005_g N_A_27_392#_M1002_g
+ N_A_27_392#_c_266_n N_A_27_392#_M1008_g N_A_27_392#_M1011_g
+ N_A_27_392#_c_267_n N_A_27_392#_c_268_n N_A_27_392#_c_253_n
+ N_A_27_392#_c_254_n N_A_27_392#_c_255_n N_A_27_392#_c_256_n
+ N_A_27_392#_c_257_n N_A_27_392#_c_258_n N_A_27_392#_c_259_n
+ N_A_27_392#_c_260_n N_A_27_392#_c_261_n N_A_27_392#_c_262_n
+ N_A_27_392#_c_263_n N_A_27_392#_c_264_n PM_SKY130_FD_SC_LS__NOR4BB_2%A_27_392#
x_PM_SKY130_FD_SC_LS__NOR4BB_2%B N_B_M1007_g N_B_M1019_g N_B_c_392_n N_B_M1009_g
+ N_B_c_393_n N_B_M1013_g B B N_B_c_391_n N_B_c_398_n
+ PM_SKY130_FD_SC_LS__NOR4BB_2%B
x_PM_SKY130_FD_SC_LS__NOR4BB_2%A N_A_M1006_g N_A_c_451_n N_A_M1003_g N_A_c_452_n
+ N_A_M1018_g N_A_M1017_g A A N_A_c_450_n PM_SKY130_FD_SC_LS__NOR4BB_2%A
x_PM_SKY130_FD_SC_LS__NOR4BB_2%VPWR N_VPWR_M1014_d N_VPWR_M1003_s N_VPWR_c_495_n
+ N_VPWR_c_496_n N_VPWR_c_497_n N_VPWR_c_498_n VPWR N_VPWR_c_499_n
+ N_VPWR_c_500_n N_VPWR_c_494_n N_VPWR_c_502_n PM_SKY130_FD_SC_LS__NOR4BB_2%VPWR
x_PM_SKY130_FD_SC_LS__NOR4BB_2%A_493_368# N_A_493_368#_M1001_d
+ N_A_493_368#_M1015_d N_A_493_368#_M1008_s N_A_493_368#_c_557_n
+ N_A_493_368#_c_553_n N_A_493_368#_c_554_n N_A_493_368#_c_568_n
+ N_A_493_368#_c_569_n N_A_493_368#_c_571_n N_A_493_368#_c_555_n
+ PM_SKY130_FD_SC_LS__NOR4BB_2%A_493_368#
x_PM_SKY130_FD_SC_LS__NOR4BB_2%Y N_Y_M1000_d N_Y_M1002_s N_Y_M1007_s N_Y_M1006_d
+ N_Y_M1001_s N_Y_c_608_n N_Y_c_609_n N_Y_c_627_n N_Y_c_596_n N_Y_c_597_n
+ N_Y_c_598_n N_Y_c_599_n N_Y_c_600_n N_Y_c_601_n N_Y_c_612_n N_Y_c_602_n
+ N_Y_c_603_n N_Y_c_606_n N_Y_c_604_n Y PM_SKY130_FD_SC_LS__NOR4BB_2%Y
x_PM_SKY130_FD_SC_LS__NOR4BB_2%A_772_368# N_A_772_368#_M1005_d
+ N_A_772_368#_M1009_d N_A_772_368#_c_726_n N_A_772_368#_c_712_n
+ N_A_772_368#_c_713_n N_A_772_368#_c_718_n
+ PM_SKY130_FD_SC_LS__NOR4BB_2%A_772_368#
x_PM_SKY130_FD_SC_LS__NOR4BB_2%A_985_368# N_A_985_368#_M1009_s
+ N_A_985_368#_M1013_s N_A_985_368#_M1018_d N_A_985_368#_c_739_n
+ N_A_985_368#_c_740_n N_A_985_368#_c_749_n N_A_985_368#_c_741_n
+ N_A_985_368#_c_758_n N_A_985_368#_c_742_n N_A_985_368#_c_743_n
+ N_A_985_368#_c_755_n PM_SKY130_FD_SC_LS__NOR4BB_2%A_985_368#
x_PM_SKY130_FD_SC_LS__NOR4BB_2%VGND N_VGND_M1016_d N_VGND_M1000_s N_VGND_M1010_s
+ N_VGND_M1011_d N_VGND_M1019_d N_VGND_M1017_s N_VGND_c_784_n N_VGND_c_785_n
+ N_VGND_c_786_n N_VGND_c_787_n N_VGND_c_788_n VGND N_VGND_c_789_n
+ N_VGND_c_790_n N_VGND_c_791_n N_VGND_c_792_n N_VGND_c_793_n N_VGND_c_794_n
+ N_VGND_c_795_n N_VGND_c_796_n N_VGND_c_797_n PM_SKY130_FD_SC_LS__NOR4BB_2%VGND
cc_1 VNB N_C_N_M1016_g 0.0481849f $X=-0.19 $Y=-0.245 $X2=0.865 $Y2=0.69
cc_2 VNB C_N 0.00306502f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_3 VNB N_C_N_c_109_n 0.0401836f $X=-0.19 $Y=-0.245 $X2=0.865 $Y2=1.677
cc_4 VNB N_D_N_c_140_n 0.045888f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.885
cc_5 VNB D_N 0.00293047f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_D_N_c_142_n 0.0269274f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_311_124#_M1000_g 0.0263535f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.677
cc_8 VNB N_A_311_124#_M1010_g 0.0258625f $X=-0.19 $Y=-0.245 $X2=1.03 $Y2=1.635
cc_9 VNB N_A_311_124#_c_178_n 0.0150347f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.635
cc_10 VNB N_A_311_124#_c_179_n 0.0424258f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_311_124#_c_180_n 0.0298372f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_392#_M1002_g 0.0261479f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.677
cc_13 VNB N_A_27_392#_M1011_g 0.0237682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_392#_c_253_n 0.0134205f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_392#_c_254_n 0.0149407f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_27_392#_c_255_n 0.0159433f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_27_392#_c_256_n 0.00987904f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_27_392#_c_257_n 0.00769251f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_27_392#_c_258_n 0.00857814f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_27_392#_c_259_n 0.0179867f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_27_392#_c_260_n 0.00704942f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_27_392#_c_261_n 0.00199894f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_27_392#_c_262_n 6.67662e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_27_392#_c_263_n 0.00295901f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_27_392#_c_264_n 0.0474555f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_B_M1007_g 0.023712f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.46
cc_27 VNB N_B_M1019_g 0.0297486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB B 0.00615235f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.635
cc_29 VNB N_B_c_391_n 0.0604396f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_M1006_g 0.0304733f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.46
cc_31 VNB N_A_M1017_g 0.032403f $X=-0.19 $Y=-0.245 $X2=0.865 $Y2=1.677
cc_32 VNB A 0.0135557f $X=-0.19 $Y=-0.245 $X2=1.03 $Y2=1.635
cc_33 VNB N_A_c_450_n 0.0513016f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VPWR_c_494_n 0.302998f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_Y_c_596_n 0.00125292f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_Y_c_597_n 0.00616913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_Y_c_598_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_Y_c_599_n 0.0110441f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_Y_c_600_n 0.00253236f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_Y_c_601_n 0.00238751f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_Y_c_602_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_Y_c_603_n 0.00176983f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_Y_c_604_n 0.00178779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB Y 0.00422131f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_784_n 0.00811375f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.635
cc_46 VNB N_VGND_c_785_n 0.00578139f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_786_n 0.0120272f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_787_n 0.0410035f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_788_n 0.0422414f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_789_n 0.0484972f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_790_n 0.0186085f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_791_n 0.0182584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_792_n 0.016966f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_793_n 0.016966f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_794_n 0.00718138f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_795_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_796_n 0.0275348f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_797_n 0.395051f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VPB N_C_N_c_110_n 0.0219367f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.885
cc_60 VPB C_N 0.00195622f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_61 VPB N_C_N_c_109_n 0.0406789f $X=-0.19 $Y=1.66 $X2=0.865 $Y2=1.677
cc_62 VPB N_D_N_c_143_n 0.0204358f $X=-0.19 $Y=1.66 $X2=0.865 $Y2=1.47
cc_63 VPB D_N 0.00280121f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_D_N_c_142_n 0.0314886f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_A_311_124#_c_181_n 0.0174519f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_A_311_124#_c_182_n 0.0152894f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_A_311_124#_c_183_n 0.0107464f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_A_311_124#_c_184_n 0.00644823f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_A_311_124#_c_185_n 0.00607539f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_A_311_124#_c_179_n 0.0211875f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_A_311_124#_c_180_n 0.0221435f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_A_27_392#_c_265_n 0.0161065f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_A_27_392#_c_266_n 0.0184063f $X=-0.19 $Y=1.66 $X2=1.03 $Y2=1.677
cc_74 VPB N_A_27_392#_c_267_n 0.00626527f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_A_27_392#_c_268_n 0.0348264f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_A_27_392#_c_259_n 0.0147077f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_A_27_392#_c_262_n 0.00138164f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_A_27_392#_c_264_n 0.025076f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 VPB N_B_c_392_n 0.018203f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_80 VPB N_B_c_393_n 0.0158237f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.677
cc_81 VPB B 0.00748815f $X=-0.19 $Y=1.66 $X2=1.2 $Y2=1.635
cc_82 VPB N_B_c_391_n 0.0373831f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 VPB N_A_c_451_n 0.0162195f $X=-0.19 $Y=1.66 $X2=0.865 $Y2=0.69
cc_84 VPB N_A_c_452_n 0.0208611f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_85 VPB A 0.0104885f $X=-0.19 $Y=1.66 $X2=1.03 $Y2=1.635
cc_86 VPB N_A_c_450_n 0.0273696f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_495_n 0.0180076f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_88 VPB N_VPWR_c_496_n 0.00799266f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_497_n 0.114199f $X=-0.19 $Y=1.66 $X2=1.2 $Y2=1.635
cc_90 VPB N_VPWR_c_498_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_499_n 0.0191515f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_500_n 0.0201062f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_494_n 0.0961603f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_502_n 0.0211323f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_95 VPB N_A_493_368#_c_553_n 0.00467121f $X=-0.19 $Y=1.66 $X2=1.03 $Y2=1.635
cc_96 VPB N_A_493_368#_c_554_n 0.00404126f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.635
cc_97 VPB N_A_493_368#_c_555_n 0.00526828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_Y_c_606_n 0.00162905f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB Y 0.00634508f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 VPB N_A_772_368#_c_712_n 0.0194809f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB N_A_772_368#_c_713_n 0.00321292f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.677
cc_102 VPB N_A_985_368#_c_739_n 0.00607444f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 VPB N_A_985_368#_c_740_n 0.00599038f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.677
cc_104 VPB N_A_985_368#_c_741_n 0.00289633f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_105 VPB N_A_985_368#_c_742_n 0.0075506f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_A_985_368#_c_743_n 0.035396f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 N_C_N_M1016_g N_D_N_c_140_n 0.0297753f $X=0.865 $Y=0.69 $X2=-0.19
+ $Y2=-0.245
cc_108 C_N D_N 0.0264922f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_109 N_C_N_c_109_n D_N 2.80835e-19 $X=0.865 $Y=1.677 $X2=0 $Y2=0
cc_110 C_N N_D_N_c_142_n 0.00255377f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_111 N_C_N_c_109_n N_D_N_c_142_n 0.0212069f $X=0.865 $Y=1.677 $X2=0 $Y2=0
cc_112 N_C_N_c_110_n N_A_27_392#_c_267_n 0.00198043f $X=0.505 $Y=1.885 $X2=0
+ $Y2=0
cc_113 N_C_N_c_110_n N_A_27_392#_c_268_n 0.00893538f $X=0.505 $Y=1.885 $X2=0
+ $Y2=0
cc_114 N_C_N_M1016_g N_A_27_392#_c_253_n 0.00828957f $X=0.865 $Y=0.69 $X2=0
+ $Y2=0
cc_115 C_N N_A_27_392#_c_253_n 0.0243439f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_116 N_C_N_c_109_n N_A_27_392#_c_253_n 0.0108906f $X=0.865 $Y=1.677 $X2=0
+ $Y2=0
cc_117 N_C_N_M1016_g N_A_27_392#_c_255_n 0.00587382f $X=0.865 $Y=0.69 $X2=0
+ $Y2=0
cc_118 N_C_N_M1016_g N_A_27_392#_c_256_n 0.00761094f $X=0.865 $Y=0.69 $X2=0
+ $Y2=0
cc_119 N_C_N_M1016_g N_A_27_392#_c_257_n 0.0111064f $X=0.865 $Y=0.69 $X2=0 $Y2=0
cc_120 C_N N_A_27_392#_c_257_n 0.0132706f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_121 N_C_N_c_109_n N_A_27_392#_c_257_n 0.00395761f $X=0.865 $Y=1.677 $X2=0
+ $Y2=0
cc_122 N_C_N_c_110_n N_A_27_392#_c_259_n 0.00278118f $X=0.505 $Y=1.885 $X2=0
+ $Y2=0
cc_123 N_C_N_M1016_g N_A_27_392#_c_259_n 0.00407288f $X=0.865 $Y=0.69 $X2=0
+ $Y2=0
cc_124 C_N N_A_27_392#_c_259_n 0.0201997f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_125 N_C_N_c_109_n N_A_27_392#_c_259_n 0.0125307f $X=0.865 $Y=1.677 $X2=0
+ $Y2=0
cc_126 N_C_N_M1016_g N_A_27_392#_c_260_n 3.84191e-19 $X=0.865 $Y=0.69 $X2=0
+ $Y2=0
cc_127 N_C_N_c_110_n N_VPWR_c_495_n 0.00565407f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_128 C_N N_VPWR_c_495_n 0.0572746f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_129 N_C_N_c_109_n N_VPWR_c_495_n 0.0140158f $X=0.865 $Y=1.677 $X2=0 $Y2=0
cc_130 N_C_N_c_110_n N_VPWR_c_499_n 0.00445602f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_131 N_C_N_c_110_n N_VPWR_c_494_n 0.00865213f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_132 N_C_N_M1016_g N_VGND_c_789_n 0.00831433f $X=0.865 $Y=0.69 $X2=0 $Y2=0
cc_133 N_C_N_M1016_g N_VGND_c_797_n 0.00424622f $X=0.865 $Y=0.69 $X2=0 $Y2=0
cc_134 N_D_N_c_140_n N_A_311_124#_c_178_n 0.0127302f $X=1.48 $Y=1.47 $X2=0 $Y2=0
cc_135 D_N N_A_311_124#_c_178_n 0.0301611f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_136 N_D_N_c_142_n N_A_311_124#_c_178_n 0.00591586f $X=1.66 $Y=1.635 $X2=0
+ $Y2=0
cc_137 N_D_N_c_143_n N_A_311_124#_c_183_n 0.00888556f $X=1.825 $Y=1.885 $X2=0
+ $Y2=0
cc_138 N_D_N_c_143_n N_A_311_124#_c_184_n 0.00203024f $X=1.825 $Y=1.885 $X2=0
+ $Y2=0
cc_139 N_D_N_c_143_n N_A_311_124#_c_185_n 0.00247102f $X=1.825 $Y=1.885 $X2=0
+ $Y2=0
cc_140 N_D_N_c_142_n N_A_311_124#_c_185_n 0.00565736f $X=1.66 $Y=1.635 $X2=0
+ $Y2=0
cc_141 N_D_N_c_140_n N_A_311_124#_c_179_n 0.00282376f $X=1.48 $Y=1.47 $X2=0
+ $Y2=0
cc_142 D_N N_A_311_124#_c_179_n 7.79116e-19 $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_143 N_D_N_c_142_n N_A_311_124#_c_179_n 0.0121608f $X=1.66 $Y=1.635 $X2=0
+ $Y2=0
cc_144 N_D_N_c_140_n N_A_27_392#_c_253_n 7.52115e-19 $X=1.48 $Y=1.47 $X2=0 $Y2=0
cc_145 N_D_N_c_140_n N_A_27_392#_c_255_n 8.70511e-19 $X=1.48 $Y=1.47 $X2=0 $Y2=0
cc_146 N_D_N_c_140_n N_A_27_392#_c_256_n 0.00110957f $X=1.48 $Y=1.47 $X2=0 $Y2=0
cc_147 N_D_N_c_140_n N_A_27_392#_c_257_n 0.0173011f $X=1.48 $Y=1.47 $X2=0 $Y2=0
cc_148 D_N N_A_27_392#_c_257_n 0.00250074f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_149 N_D_N_c_142_n N_A_27_392#_c_257_n 3.6161e-19 $X=1.66 $Y=1.635 $X2=0 $Y2=0
cc_150 N_D_N_c_143_n N_VPWR_c_495_n 0.00565407f $X=1.825 $Y=1.885 $X2=0 $Y2=0
cc_151 D_N N_VPWR_c_495_n 0.0171462f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_152 N_D_N_c_142_n N_VPWR_c_495_n 0.00605928f $X=1.66 $Y=1.635 $X2=0 $Y2=0
cc_153 N_D_N_c_143_n N_VPWR_c_497_n 0.00445602f $X=1.825 $Y=1.885 $X2=0 $Y2=0
cc_154 N_D_N_c_143_n N_VPWR_c_494_n 0.00866521f $X=1.825 $Y=1.885 $X2=0 $Y2=0
cc_155 N_D_N_c_143_n N_A_493_368#_c_554_n 0.00271992f $X=1.825 $Y=1.885 $X2=0
+ $Y2=0
cc_156 N_D_N_c_140_n N_VGND_c_788_n 0.00808015f $X=1.48 $Y=1.47 $X2=0 $Y2=0
cc_157 N_D_N_c_140_n N_VGND_c_789_n 0.0241121f $X=1.48 $Y=1.47 $X2=0 $Y2=0
cc_158 N_D_N_c_140_n N_VGND_c_797_n 0.00122193f $X=1.48 $Y=1.47 $X2=0 $Y2=0
cc_159 N_A_311_124#_c_182_n N_A_27_392#_c_265_n 0.0304639f $X=3.285 $Y=1.765
+ $X2=0 $Y2=0
cc_160 N_A_311_124#_M1010_g N_A_27_392#_M1002_g 0.021145f $X=3.27 $Y=0.74 $X2=0
+ $Y2=0
cc_161 N_A_311_124#_M1004_d N_A_27_392#_c_257_n 0.0115648f $X=1.555 $Y=0.62
+ $X2=0 $Y2=0
cc_162 N_A_311_124#_c_178_n N_A_27_392#_c_257_n 0.0544489f $X=2.155 $Y=1.175
+ $X2=0 $Y2=0
cc_163 N_A_311_124#_c_202_p N_A_27_392#_c_257_n 0.00570404f $X=3 $Y=1.515 $X2=0
+ $Y2=0
cc_164 N_A_311_124#_c_179_n N_A_27_392#_c_257_n 0.00368582f $X=2.745 $Y=1.515
+ $X2=0 $Y2=0
cc_165 N_A_311_124#_M1000_g N_A_27_392#_c_258_n 0.0150458f $X=2.84 $Y=0.74 $X2=0
+ $Y2=0
cc_166 N_A_311_124#_M1010_g N_A_27_392#_c_258_n 0.0133835f $X=3.27 $Y=0.74 $X2=0
+ $Y2=0
cc_167 N_A_311_124#_c_202_p N_A_27_392#_c_258_n 0.0369816f $X=3 $Y=1.515 $X2=0
+ $Y2=0
cc_168 N_A_311_124#_c_179_n N_A_27_392#_c_258_n 0.00225781f $X=2.745 $Y=1.515
+ $X2=0 $Y2=0
cc_169 N_A_311_124#_c_180_n N_A_27_392#_c_258_n 0.0029606f $X=3.27 $Y=1.557
+ $X2=0 $Y2=0
cc_170 N_A_311_124#_M1000_g N_A_27_392#_c_261_n 0.0102303f $X=2.84 $Y=0.74 $X2=0
+ $Y2=0
cc_171 N_A_311_124#_c_178_n N_A_27_392#_c_261_n 0.00962897f $X=2.155 $Y=1.175
+ $X2=0 $Y2=0
cc_172 N_A_311_124#_c_202_p N_A_27_392#_c_261_n 0.0137448f $X=3 $Y=1.515 $X2=0
+ $Y2=0
cc_173 N_A_311_124#_c_179_n N_A_27_392#_c_261_n 0.00386621f $X=2.745 $Y=1.515
+ $X2=0 $Y2=0
cc_174 N_A_311_124#_c_202_p N_A_27_392#_c_262_n 0.0118608f $X=3 $Y=1.515 $X2=0
+ $Y2=0
cc_175 N_A_311_124#_c_180_n N_A_27_392#_c_262_n 0.0015832f $X=3.27 $Y=1.557
+ $X2=0 $Y2=0
cc_176 N_A_311_124#_M1010_g N_A_27_392#_c_263_n 0.00337019f $X=3.27 $Y=0.74
+ $X2=0 $Y2=0
cc_177 N_A_311_124#_c_202_p N_A_27_392#_c_264_n 0.00105222f $X=3 $Y=1.515 $X2=0
+ $Y2=0
cc_178 N_A_311_124#_c_180_n N_A_27_392#_c_264_n 0.0227948f $X=3.27 $Y=1.557
+ $X2=0 $Y2=0
cc_179 N_A_311_124#_c_184_n N_VPWR_c_495_n 0.0390291f $X=2.05 $Y=2.135 $X2=0
+ $Y2=0
cc_180 N_A_311_124#_c_181_n N_VPWR_c_497_n 0.00278257f $X=2.835 $Y=1.765 $X2=0
+ $Y2=0
cc_181 N_A_311_124#_c_182_n N_VPWR_c_497_n 0.00278271f $X=3.285 $Y=1.765 $X2=0
+ $Y2=0
cc_182 N_A_311_124#_c_183_n N_VPWR_c_497_n 0.0145938f $X=2.05 $Y=2.815 $X2=0
+ $Y2=0
cc_183 N_A_311_124#_c_181_n N_VPWR_c_494_n 0.00358623f $X=2.835 $Y=1.765 $X2=0
+ $Y2=0
cc_184 N_A_311_124#_c_182_n N_VPWR_c_494_n 0.00354337f $X=3.285 $Y=1.765 $X2=0
+ $Y2=0
cc_185 N_A_311_124#_c_183_n N_VPWR_c_494_n 0.0120466f $X=2.05 $Y=2.815 $X2=0
+ $Y2=0
cc_186 N_A_311_124#_c_181_n N_A_493_368#_c_557_n 0.0127774f $X=2.835 $Y=1.765
+ $X2=0 $Y2=0
cc_187 N_A_311_124#_c_182_n N_A_493_368#_c_557_n 7.89375e-19 $X=3.285 $Y=1.765
+ $X2=0 $Y2=0
cc_188 N_A_311_124#_c_183_n N_A_493_368#_c_557_n 0.0432034f $X=2.05 $Y=2.815
+ $X2=0 $Y2=0
cc_189 N_A_311_124#_c_202_p N_A_493_368#_c_557_n 0.0202808f $X=3 $Y=1.515 $X2=0
+ $Y2=0
cc_190 N_A_311_124#_c_185_n N_A_493_368#_c_557_n 0.0232212f $X=2.105 $Y=1.97
+ $X2=0 $Y2=0
cc_191 N_A_311_124#_c_179_n N_A_493_368#_c_557_n 0.00565239f $X=2.745 $Y=1.515
+ $X2=0 $Y2=0
cc_192 N_A_311_124#_c_181_n N_A_493_368#_c_553_n 0.0108414f $X=2.835 $Y=1.765
+ $X2=0 $Y2=0
cc_193 N_A_311_124#_c_182_n N_A_493_368#_c_553_n 0.013742f $X=3.285 $Y=1.765
+ $X2=0 $Y2=0
cc_194 N_A_311_124#_c_181_n N_A_493_368#_c_554_n 0.00253887f $X=2.835 $Y=1.765
+ $X2=0 $Y2=0
cc_195 N_A_311_124#_c_183_n N_A_493_368#_c_554_n 0.00457905f $X=2.05 $Y=2.815
+ $X2=0 $Y2=0
cc_196 N_A_311_124#_M1010_g N_Y_c_608_n 0.010397f $X=3.27 $Y=0.74 $X2=0 $Y2=0
cc_197 N_A_311_124#_c_182_n N_Y_c_609_n 0.0141859f $X=3.285 $Y=1.765 $X2=0 $Y2=0
cc_198 N_A_311_124#_M1000_g N_Y_c_601_n 0.0131323f $X=2.84 $Y=0.74 $X2=0 $Y2=0
cc_199 N_A_311_124#_M1010_g N_Y_c_601_n 0.00825973f $X=3.27 $Y=0.74 $X2=0 $Y2=0
cc_200 N_A_311_124#_c_181_n N_Y_c_612_n 0.00318422f $X=2.835 $Y=1.765 $X2=0
+ $Y2=0
cc_201 N_A_311_124#_c_182_n N_Y_c_612_n 0.0106928f $X=3.285 $Y=1.765 $X2=0 $Y2=0
cc_202 N_A_311_124#_c_202_p N_Y_c_612_n 0.0151518f $X=3 $Y=1.515 $X2=0 $Y2=0
cc_203 N_A_311_124#_c_180_n N_Y_c_612_n 0.00547037f $X=3.27 $Y=1.557 $X2=0 $Y2=0
cc_204 N_A_311_124#_M1010_g N_Y_c_602_n 0.00160592f $X=3.27 $Y=0.74 $X2=0 $Y2=0
cc_205 N_A_311_124#_c_178_n N_VGND_M1000_s 0.00212811f $X=2.155 $Y=1.175 $X2=0
+ $Y2=0
cc_206 N_A_311_124#_M1010_g N_VGND_c_784_n 0.00436974f $X=3.27 $Y=0.74 $X2=0
+ $Y2=0
cc_207 N_A_311_124#_M1000_g N_VGND_c_788_n 0.00856324f $X=2.84 $Y=0.74 $X2=0
+ $Y2=0
cc_208 N_A_311_124#_M1000_g N_VGND_c_790_n 0.00434272f $X=2.84 $Y=0.74 $X2=0
+ $Y2=0
cc_209 N_A_311_124#_M1010_g N_VGND_c_790_n 0.00324657f $X=3.27 $Y=0.74 $X2=0
+ $Y2=0
cc_210 N_A_311_124#_M1000_g N_VGND_c_797_n 0.00825283f $X=2.84 $Y=0.74 $X2=0
+ $Y2=0
cc_211 N_A_311_124#_M1010_g N_VGND_c_797_n 0.00411452f $X=3.27 $Y=0.74 $X2=0
+ $Y2=0
cc_212 N_A_27_392#_M1011_g N_B_M1007_g 0.0171226f $X=4.335 $Y=0.74 $X2=0 $Y2=0
cc_213 N_A_27_392#_c_264_n N_B_c_391_n 0.0225964f $X=4.285 $Y=1.557 $X2=0 $Y2=0
cc_214 N_A_27_392#_c_264_n N_B_c_398_n 9.08473e-19 $X=4.285 $Y=1.557 $X2=0 $Y2=0
cc_215 N_A_27_392#_c_267_n N_VPWR_c_495_n 0.0387421f $X=0.28 $Y=2.135 $X2=0
+ $Y2=0
cc_216 N_A_27_392#_c_265_n N_VPWR_c_497_n 0.0044313f $X=3.785 $Y=1.765 $X2=0
+ $Y2=0
cc_217 N_A_27_392#_c_266_n N_VPWR_c_497_n 0.00278271f $X=4.285 $Y=1.765 $X2=0
+ $Y2=0
cc_218 N_A_27_392#_c_268_n N_VPWR_c_499_n 0.0145938f $X=0.28 $Y=2.815 $X2=0
+ $Y2=0
cc_219 N_A_27_392#_c_265_n N_VPWR_c_494_n 0.00855098f $X=3.785 $Y=1.765 $X2=0
+ $Y2=0
cc_220 N_A_27_392#_c_266_n N_VPWR_c_494_n 0.00359085f $X=4.285 $Y=1.765 $X2=0
+ $Y2=0
cc_221 N_A_27_392#_c_268_n N_VPWR_c_494_n 0.0120466f $X=0.28 $Y=2.815 $X2=0
+ $Y2=0
cc_222 N_A_27_392#_c_265_n N_A_493_368#_c_553_n 0.00327969f $X=3.785 $Y=1.765
+ $X2=0 $Y2=0
cc_223 N_A_27_392#_c_265_n N_A_493_368#_c_568_n 4.27055e-19 $X=3.785 $Y=1.765
+ $X2=0 $Y2=0
cc_224 N_A_27_392#_c_265_n N_A_493_368#_c_569_n 0.00755948f $X=3.785 $Y=1.765
+ $X2=0 $Y2=0
cc_225 N_A_27_392#_c_266_n N_A_493_368#_c_569_n 5.31972e-19 $X=4.285 $Y=1.765
+ $X2=0 $Y2=0
cc_226 N_A_27_392#_c_265_n N_A_493_368#_c_571_n 0.0122806f $X=3.785 $Y=1.765
+ $X2=0 $Y2=0
cc_227 N_A_27_392#_c_266_n N_A_493_368#_c_571_n 0.0102892f $X=4.285 $Y=1.765
+ $X2=0 $Y2=0
cc_228 N_A_27_392#_c_264_n N_A_493_368#_c_571_n 4.45802e-19 $X=4.285 $Y=1.557
+ $X2=0 $Y2=0
cc_229 N_A_27_392#_c_265_n N_A_493_368#_c_555_n 5.62223e-19 $X=3.785 $Y=1.765
+ $X2=0 $Y2=0
cc_230 N_A_27_392#_c_266_n N_A_493_368#_c_555_n 0.00580253f $X=4.285 $Y=1.765
+ $X2=0 $Y2=0
cc_231 N_A_27_392#_c_258_n N_Y_M1000_d 0.00176461f $X=3.615 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_232 N_A_27_392#_M1002_g N_Y_c_608_n 0.012023f $X=3.905 $Y=0.74 $X2=0 $Y2=0
cc_233 N_A_27_392#_c_258_n N_Y_c_608_n 0.0367463f $X=3.615 $Y=1.095 $X2=0 $Y2=0
cc_234 N_A_27_392#_c_262_n N_Y_c_608_n 0.00401767f $X=3.78 $Y=1.515 $X2=0 $Y2=0
cc_235 N_A_27_392#_c_264_n N_Y_c_608_n 5.55922e-19 $X=4.285 $Y=1.557 $X2=0 $Y2=0
cc_236 N_A_27_392#_c_265_n N_Y_c_609_n 0.0106888f $X=3.785 $Y=1.765 $X2=0 $Y2=0
cc_237 N_A_27_392#_c_266_n N_Y_c_609_n 3.00121e-19 $X=4.285 $Y=1.765 $X2=0 $Y2=0
cc_238 N_A_27_392#_c_258_n N_Y_c_609_n 0.00917652f $X=3.615 $Y=1.095 $X2=0 $Y2=0
cc_239 N_A_27_392#_c_262_n N_Y_c_609_n 0.020545f $X=3.78 $Y=1.515 $X2=0 $Y2=0
cc_240 N_A_27_392#_c_264_n N_Y_c_609_n 0.0061371f $X=4.285 $Y=1.557 $X2=0 $Y2=0
cc_241 N_A_27_392#_M1002_g N_Y_c_627_n 0.00358524f $X=3.905 $Y=0.74 $X2=0 $Y2=0
cc_242 N_A_27_392#_M1011_g N_Y_c_627_n 0.00324256f $X=4.335 $Y=0.74 $X2=0 $Y2=0
cc_243 N_A_27_392#_M1002_g N_Y_c_596_n 0.00132575f $X=3.905 $Y=0.74 $X2=0 $Y2=0
cc_244 N_A_27_392#_M1011_g N_Y_c_596_n 0.00426553f $X=4.335 $Y=0.74 $X2=0 $Y2=0
cc_245 N_A_27_392#_c_262_n N_Y_c_596_n 0.0235323f $X=3.78 $Y=1.515 $X2=0 $Y2=0
cc_246 N_A_27_392#_c_263_n N_Y_c_596_n 0.007992f $X=3.78 $Y=1.35 $X2=0 $Y2=0
cc_247 N_A_27_392#_c_264_n N_Y_c_596_n 0.0104007f $X=4.285 $Y=1.557 $X2=0 $Y2=0
cc_248 N_A_27_392#_M1011_g N_Y_c_597_n 0.0121595f $X=4.335 $Y=0.74 $X2=0 $Y2=0
cc_249 N_A_27_392#_M1002_g N_Y_c_601_n 8.5656e-19 $X=3.905 $Y=0.74 $X2=0 $Y2=0
cc_250 N_A_27_392#_c_258_n N_Y_c_601_n 0.01663f $X=3.615 $Y=1.095 $X2=0 $Y2=0
cc_251 N_A_27_392#_c_261_n N_Y_c_601_n 0.00773618f $X=2.58 $Y=0.795 $X2=0 $Y2=0
cc_252 N_A_27_392#_c_265_n N_Y_c_612_n 8.78539e-19 $X=3.785 $Y=1.765 $X2=0 $Y2=0
cc_253 N_A_27_392#_c_258_n N_Y_c_612_n 9.44131e-19 $X=3.615 $Y=1.095 $X2=0 $Y2=0
cc_254 N_A_27_392#_M1002_g N_Y_c_602_n 0.00731716f $X=3.905 $Y=0.74 $X2=0 $Y2=0
cc_255 N_A_27_392#_M1011_g N_Y_c_602_n 0.00619455f $X=4.335 $Y=0.74 $X2=0 $Y2=0
cc_256 N_A_27_392#_M1002_g N_Y_c_603_n 0.00323058f $X=3.905 $Y=0.74 $X2=0 $Y2=0
cc_257 N_A_27_392#_M1011_g N_Y_c_603_n 0.00121492f $X=4.335 $Y=0.74 $X2=0 $Y2=0
cc_258 N_A_27_392#_c_258_n N_Y_c_603_n 0.0104256f $X=3.615 $Y=1.095 $X2=0 $Y2=0
cc_259 N_A_27_392#_c_264_n N_Y_c_603_n 0.00135793f $X=4.285 $Y=1.557 $X2=0 $Y2=0
cc_260 N_A_27_392#_c_265_n N_Y_c_606_n 0.00180311f $X=3.785 $Y=1.765 $X2=0 $Y2=0
cc_261 N_A_27_392#_c_266_n N_Y_c_606_n 0.00988825f $X=4.285 $Y=1.765 $X2=0 $Y2=0
cc_262 N_A_27_392#_c_264_n N_Y_c_606_n 0.00933825f $X=4.285 $Y=1.557 $X2=0 $Y2=0
cc_263 N_A_27_392#_c_266_n Y 0.00211858f $X=4.285 $Y=1.765 $X2=0 $Y2=0
cc_264 N_A_27_392#_c_264_n Y 0.00958836f $X=4.285 $Y=1.557 $X2=0 $Y2=0
cc_265 N_A_27_392#_c_266_n N_A_772_368#_c_712_n 0.0128758f $X=4.285 $Y=1.765
+ $X2=0 $Y2=0
cc_266 N_A_27_392#_c_265_n N_A_772_368#_c_713_n 0.00136321f $X=3.785 $Y=1.765
+ $X2=0 $Y2=0
cc_267 N_A_27_392#_c_266_n N_A_985_368#_c_739_n 0.00545516f $X=4.285 $Y=1.765
+ $X2=0 $Y2=0
cc_268 N_A_27_392#_c_257_n N_VGND_M1016_d 0.0115959f $X=2.495 $Y=0.795 $X2=-0.19
+ $Y2=-0.245
cc_269 N_A_27_392#_c_257_n N_VGND_M1000_s 0.00942815f $X=2.495 $Y=0.795 $X2=0
+ $Y2=0
cc_270 N_A_27_392#_c_258_n N_VGND_M1000_s 0.00104037f $X=3.615 $Y=1.095 $X2=0
+ $Y2=0
cc_271 N_A_27_392#_c_261_n N_VGND_M1000_s 0.0152615f $X=2.58 $Y=0.795 $X2=0
+ $Y2=0
cc_272 N_A_27_392#_c_258_n N_VGND_M1010_s 0.00530094f $X=3.615 $Y=1.095 $X2=0
+ $Y2=0
cc_273 N_A_27_392#_M1002_g N_VGND_c_784_n 0.00436974f $X=3.905 $Y=0.74 $X2=0
+ $Y2=0
cc_274 N_A_27_392#_M1011_g N_VGND_c_785_n 0.00571035f $X=4.335 $Y=0.74 $X2=0
+ $Y2=0
cc_275 N_A_27_392#_c_257_n N_VGND_c_788_n 0.033238f $X=2.495 $Y=0.795 $X2=0
+ $Y2=0
cc_276 N_A_27_392#_c_258_n N_VGND_c_788_n 0.0016343f $X=3.615 $Y=1.095 $X2=0
+ $Y2=0
cc_277 N_A_27_392#_c_261_n N_VGND_c_788_n 0.0140889f $X=2.58 $Y=0.795 $X2=0
+ $Y2=0
cc_278 N_A_27_392#_c_255_n N_VGND_c_789_n 0.0209923f $X=0.65 $Y=0.525 $X2=0
+ $Y2=0
cc_279 N_A_27_392#_c_257_n N_VGND_c_789_n 0.040123f $X=2.495 $Y=0.795 $X2=0
+ $Y2=0
cc_280 N_A_27_392#_M1002_g N_VGND_c_791_n 0.00324657f $X=3.905 $Y=0.74 $X2=0
+ $Y2=0
cc_281 N_A_27_392#_M1011_g N_VGND_c_791_n 0.00434272f $X=4.335 $Y=0.74 $X2=0
+ $Y2=0
cc_282 N_A_27_392#_M1002_g N_VGND_c_797_n 0.00411452f $X=3.905 $Y=0.74 $X2=0
+ $Y2=0
cc_283 N_A_27_392#_M1011_g N_VGND_c_797_n 0.00820772f $X=4.335 $Y=0.74 $X2=0
+ $Y2=0
cc_284 N_A_27_392#_c_255_n N_VGND_c_797_n 0.0119247f $X=0.65 $Y=0.525 $X2=0
+ $Y2=0
cc_285 N_A_27_392#_c_257_n N_VGND_c_797_n 0.0255197f $X=2.495 $Y=0.795 $X2=0
+ $Y2=0
cc_286 N_A_27_392#_c_261_n N_VGND_c_797_n 7.23349e-19 $X=2.58 $Y=0.795 $X2=0
+ $Y2=0
cc_287 N_B_c_393_n N_A_c_451_n 0.0228597f $X=5.745 $Y=1.765 $X2=0 $Y2=0
cc_288 B A 0.034382f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_289 N_B_c_391_n A 2.83596e-19 $X=5.64 $Y=1.515 $X2=0 $Y2=0
cc_290 B N_A_c_450_n 0.00479375f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_291 N_B_c_391_n N_A_c_450_n 0.0135817f $X=5.64 $Y=1.515 $X2=0 $Y2=0
cc_292 N_B_c_392_n N_VPWR_c_497_n 0.00278257f $X=5.295 $Y=1.765 $X2=0 $Y2=0
cc_293 N_B_c_393_n N_VPWR_c_497_n 0.0044313f $X=5.745 $Y=1.765 $X2=0 $Y2=0
cc_294 N_B_c_392_n N_VPWR_c_494_n 0.00358623f $X=5.295 $Y=1.765 $X2=0 $Y2=0
cc_295 N_B_c_393_n N_VPWR_c_494_n 0.00854637f $X=5.745 $Y=1.765 $X2=0 $Y2=0
cc_296 N_B_M1007_g N_Y_c_627_n 7.28304e-19 $X=4.835 $Y=0.74 $X2=0 $Y2=0
cc_297 N_B_M1007_g N_Y_c_596_n 8.18227e-19 $X=4.835 $Y=0.74 $X2=0 $Y2=0
cc_298 N_B_c_398_n N_Y_c_596_n 0.00554962f $X=5.405 $Y=1.565 $X2=0 $Y2=0
cc_299 N_B_M1007_g N_Y_c_597_n 0.0162328f $X=4.835 $Y=0.74 $X2=0 $Y2=0
cc_300 N_B_c_398_n N_Y_c_597_n 0.00758f $X=5.405 $Y=1.565 $X2=0 $Y2=0
cc_301 N_B_M1007_g N_Y_c_598_n 3.97481e-19 $X=4.835 $Y=0.74 $X2=0 $Y2=0
cc_302 N_B_M1019_g N_Y_c_598_n 0.0132814f $X=5.265 $Y=0.74 $X2=0 $Y2=0
cc_303 N_B_M1019_g N_Y_c_599_n 0.0131358f $X=5.265 $Y=0.74 $X2=0 $Y2=0
cc_304 N_B_c_391_n N_Y_c_599_n 0.0111596f $X=5.64 $Y=1.515 $X2=0 $Y2=0
cc_305 N_B_c_398_n N_Y_c_599_n 0.0693712f $X=5.405 $Y=1.565 $X2=0 $Y2=0
cc_306 N_B_c_391_n N_Y_c_606_n 8.18227e-19 $X=5.64 $Y=1.515 $X2=0 $Y2=0
cc_307 N_B_M1019_g N_Y_c_604_n 0.00157732f $X=5.265 $Y=0.74 $X2=0 $Y2=0
cc_308 N_B_c_391_n N_Y_c_604_n 0.00232957f $X=5.64 $Y=1.515 $X2=0 $Y2=0
cc_309 N_B_c_398_n N_Y_c_604_n 0.0207638f $X=5.405 $Y=1.565 $X2=0 $Y2=0
cc_310 N_B_c_392_n Y 3.47741e-19 $X=5.295 $Y=1.765 $X2=0 $Y2=0
cc_311 N_B_c_391_n Y 0.00456209f $X=5.64 $Y=1.515 $X2=0 $Y2=0
cc_312 N_B_c_398_n Y 0.00664505f $X=5.405 $Y=1.565 $X2=0 $Y2=0
cc_313 N_B_c_392_n N_A_772_368#_c_712_n 0.0145139f $X=5.295 $Y=1.765 $X2=0 $Y2=0
cc_314 N_B_c_393_n N_A_772_368#_c_712_n 0.00416253f $X=5.745 $Y=1.765 $X2=0
+ $Y2=0
cc_315 N_B_c_392_n N_A_772_368#_c_718_n 0.0121561f $X=5.295 $Y=1.765 $X2=0 $Y2=0
cc_316 N_B_c_393_n N_A_772_368#_c_718_n 0.00604065f $X=5.745 $Y=1.765 $X2=0
+ $Y2=0
cc_317 N_B_c_392_n N_A_985_368#_c_739_n 0.00314968f $X=5.295 $Y=1.765 $X2=0
+ $Y2=0
cc_318 N_B_c_391_n N_A_985_368#_c_739_n 0.00671543f $X=5.64 $Y=1.515 $X2=0 $Y2=0
cc_319 N_B_c_398_n N_A_985_368#_c_739_n 0.0195868f $X=5.405 $Y=1.565 $X2=0 $Y2=0
cc_320 N_B_c_392_n N_A_985_368#_c_740_n 0.00881943f $X=5.295 $Y=1.765 $X2=0
+ $Y2=0
cc_321 N_B_c_392_n N_A_985_368#_c_749_n 0.0134968f $X=5.295 $Y=1.765 $X2=0 $Y2=0
cc_322 N_B_c_393_n N_A_985_368#_c_749_n 0.0150982f $X=5.745 $Y=1.765 $X2=0 $Y2=0
cc_323 B N_A_985_368#_c_749_n 0.0306997f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_324 N_B_c_391_n N_A_985_368#_c_749_n 0.00235538f $X=5.64 $Y=1.515 $X2=0 $Y2=0
cc_325 N_B_c_398_n N_A_985_368#_c_749_n 0.00882073f $X=5.405 $Y=1.565 $X2=0
+ $Y2=0
cc_326 N_B_c_393_n N_A_985_368#_c_741_n 0.00464012f $X=5.745 $Y=1.765 $X2=0
+ $Y2=0
cc_327 B N_A_985_368#_c_755_n 0.0219062f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_328 N_B_M1007_g N_VGND_c_785_n 0.0108107f $X=4.835 $Y=0.74 $X2=0 $Y2=0
cc_329 N_B_M1019_g N_VGND_c_785_n 5.17822e-19 $X=5.265 $Y=0.74 $X2=0 $Y2=0
cc_330 N_B_M1007_g N_VGND_c_792_n 0.00383152f $X=4.835 $Y=0.74 $X2=0 $Y2=0
cc_331 N_B_M1019_g N_VGND_c_792_n 0.00434272f $X=5.265 $Y=0.74 $X2=0 $Y2=0
cc_332 N_B_M1019_g N_VGND_c_796_n 0.00596513f $X=5.265 $Y=0.74 $X2=0 $Y2=0
cc_333 N_B_M1007_g N_VGND_c_797_n 0.0075754f $X=4.835 $Y=0.74 $X2=0 $Y2=0
cc_334 N_B_M1019_g N_VGND_c_797_n 0.00825059f $X=5.265 $Y=0.74 $X2=0 $Y2=0
cc_335 N_A_c_451_n N_VPWR_c_496_n 0.00486623f $X=6.245 $Y=1.765 $X2=0 $Y2=0
cc_336 N_A_c_452_n N_VPWR_c_496_n 0.00486623f $X=6.695 $Y=1.765 $X2=0 $Y2=0
cc_337 N_A_c_451_n N_VPWR_c_497_n 0.00445602f $X=6.245 $Y=1.765 $X2=0 $Y2=0
cc_338 N_A_c_452_n N_VPWR_c_500_n 0.00445602f $X=6.695 $Y=1.765 $X2=0 $Y2=0
cc_339 N_A_c_451_n N_VPWR_c_494_n 0.00858104f $X=6.245 $Y=1.765 $X2=0 $Y2=0
cc_340 N_A_c_452_n N_VPWR_c_494_n 0.00861084f $X=6.695 $Y=1.765 $X2=0 $Y2=0
cc_341 N_A_M1006_g N_Y_c_599_n 0.0203499f $X=6.23 $Y=0.74 $X2=0 $Y2=0
cc_342 N_A_M1017_g N_Y_c_599_n 0.00178479f $X=6.705 $Y=0.74 $X2=0 $Y2=0
cc_343 A N_Y_c_599_n 0.0225881f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_344 N_A_c_450_n N_Y_c_599_n 0.00337787f $X=6.705 $Y=1.557 $X2=0 $Y2=0
cc_345 N_A_M1006_g N_Y_c_600_n 4.74419e-19 $X=6.23 $Y=0.74 $X2=0 $Y2=0
cc_346 N_A_M1017_g N_Y_c_600_n 4.44219e-19 $X=6.705 $Y=0.74 $X2=0 $Y2=0
cc_347 N_A_c_451_n N_A_772_368#_c_712_n 4.63564e-19 $X=6.245 $Y=1.765 $X2=0
+ $Y2=0
cc_348 N_A_c_451_n N_A_985_368#_c_741_n 0.0103949f $X=6.245 $Y=1.765 $X2=0 $Y2=0
cc_349 N_A_c_452_n N_A_985_368#_c_741_n 6.45594e-19 $X=6.695 $Y=1.765 $X2=0
+ $Y2=0
cc_350 N_A_c_451_n N_A_985_368#_c_758_n 0.0157945f $X=6.245 $Y=1.765 $X2=0 $Y2=0
cc_351 N_A_c_452_n N_A_985_368#_c_758_n 0.0120074f $X=6.695 $Y=1.765 $X2=0 $Y2=0
cc_352 A N_A_985_368#_c_758_n 0.0303009f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_353 N_A_c_450_n N_A_985_368#_c_758_n 0.00131177f $X=6.705 $Y=1.557 $X2=0
+ $Y2=0
cc_354 N_A_c_452_n N_A_985_368#_c_742_n 4.27055e-19 $X=6.695 $Y=1.765 $X2=0
+ $Y2=0
cc_355 A N_A_985_368#_c_742_n 0.0255992f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_356 N_A_c_450_n N_A_985_368#_c_742_n 0.00109667f $X=6.705 $Y=1.557 $X2=0
+ $Y2=0
cc_357 N_A_c_451_n N_A_985_368#_c_743_n 6.45594e-19 $X=6.245 $Y=1.765 $X2=0
+ $Y2=0
cc_358 N_A_c_452_n N_A_985_368#_c_743_n 0.0105912f $X=6.695 $Y=1.765 $X2=0 $Y2=0
cc_359 N_A_c_451_n N_A_985_368#_c_755_n 9.50925e-19 $X=6.245 $Y=1.765 $X2=0
+ $Y2=0
cc_360 N_A_M1006_g N_VGND_c_787_n 5.53719e-19 $X=6.23 $Y=0.74 $X2=0 $Y2=0
cc_361 N_A_M1017_g N_VGND_c_787_n 0.0152652f $X=6.705 $Y=0.74 $X2=0 $Y2=0
cc_362 A N_VGND_c_787_n 0.022893f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_363 N_A_c_450_n N_VGND_c_787_n 0.00454352f $X=6.705 $Y=1.557 $X2=0 $Y2=0
cc_364 N_A_M1006_g N_VGND_c_793_n 0.00461464f $X=6.23 $Y=0.74 $X2=0 $Y2=0
cc_365 N_A_M1017_g N_VGND_c_793_n 0.00383152f $X=6.705 $Y=0.74 $X2=0 $Y2=0
cc_366 N_A_M1006_g N_VGND_c_796_n 0.0063291f $X=6.23 $Y=0.74 $X2=0 $Y2=0
cc_367 N_A_M1006_g N_VGND_c_797_n 0.00912532f $X=6.23 $Y=0.74 $X2=0 $Y2=0
cc_368 N_A_M1017_g N_VGND_c_797_n 0.00757973f $X=6.705 $Y=0.74 $X2=0 $Y2=0
cc_369 N_VPWR_c_497_n N_A_493_368#_c_553_n 0.0626582f $X=6.385 $Y=3.33 $X2=0
+ $Y2=0
cc_370 N_VPWR_c_494_n N_A_493_368#_c_553_n 0.0347672f $X=6.96 $Y=3.33 $X2=0
+ $Y2=0
cc_371 N_VPWR_c_497_n N_A_493_368#_c_554_n 0.0200196f $X=6.385 $Y=3.33 $X2=0
+ $Y2=0
cc_372 N_VPWR_c_494_n N_A_493_368#_c_554_n 0.0108171f $X=6.96 $Y=3.33 $X2=0
+ $Y2=0
cc_373 N_VPWR_c_497_n N_A_772_368#_c_712_n 0.0986536f $X=6.385 $Y=3.33 $X2=0
+ $Y2=0
cc_374 N_VPWR_c_494_n N_A_772_368#_c_712_n 0.0557499f $X=6.96 $Y=3.33 $X2=0
+ $Y2=0
cc_375 N_VPWR_c_497_n N_A_772_368#_c_713_n 0.0197429f $X=6.385 $Y=3.33 $X2=0
+ $Y2=0
cc_376 N_VPWR_c_494_n N_A_772_368#_c_713_n 0.0108239f $X=6.96 $Y=3.33 $X2=0
+ $Y2=0
cc_377 N_VPWR_c_496_n N_A_985_368#_c_741_n 0.0449718f $X=6.47 $Y=2.455 $X2=0
+ $Y2=0
cc_378 N_VPWR_c_497_n N_A_985_368#_c_741_n 0.0145938f $X=6.385 $Y=3.33 $X2=0
+ $Y2=0
cc_379 N_VPWR_c_494_n N_A_985_368#_c_741_n 0.0120466f $X=6.96 $Y=3.33 $X2=0
+ $Y2=0
cc_380 N_VPWR_M1003_s N_A_985_368#_c_758_n 0.00408911f $X=6.32 $Y=1.84 $X2=0
+ $Y2=0
cc_381 N_VPWR_c_496_n N_A_985_368#_c_758_n 0.0136682f $X=6.47 $Y=2.455 $X2=0
+ $Y2=0
cc_382 N_VPWR_c_496_n N_A_985_368#_c_743_n 0.0449718f $X=6.47 $Y=2.455 $X2=0
+ $Y2=0
cc_383 N_VPWR_c_500_n N_A_985_368#_c_743_n 0.0145938f $X=6.96 $Y=3.33 $X2=0
+ $Y2=0
cc_384 N_VPWR_c_494_n N_A_985_368#_c_743_n 0.0120466f $X=6.96 $Y=3.33 $X2=0
+ $Y2=0
cc_385 N_A_493_368#_c_553_n N_Y_M1001_s 0.00222494f $X=3.395 $Y=2.99 $X2=0 $Y2=0
cc_386 N_A_493_368#_M1015_d N_Y_c_609_n 0.00699639f $X=3.36 $Y=1.84 $X2=0 $Y2=0
cc_387 N_A_493_368#_c_568_n N_Y_c_609_n 0.0203011f $X=3.56 $Y=2.36 $X2=0 $Y2=0
cc_388 N_A_493_368#_c_571_n N_Y_c_609_n 0.0234979f $X=4.345 $Y=2.275 $X2=0 $Y2=0
cc_389 N_A_493_368#_c_557_n N_Y_c_612_n 0.0595639f $X=2.61 $Y=2.015 $X2=0 $Y2=0
cc_390 N_A_493_368#_c_553_n N_Y_c_612_n 0.0144323f $X=3.395 $Y=2.99 $X2=0 $Y2=0
cc_391 N_A_493_368#_c_571_n N_Y_c_606_n 0.00864724f $X=4.345 $Y=2.275 $X2=0
+ $Y2=0
cc_392 N_A_493_368#_c_571_n Y 0.00203023f $X=4.345 $Y=2.275 $X2=0 $Y2=0
cc_393 N_A_493_368#_c_555_n Y 0.0131966f $X=4.51 $Y=2.275 $X2=0 $Y2=0
cc_394 N_A_493_368#_c_571_n N_A_772_368#_M1005_d 0.00474045f $X=4.345 $Y=2.275
+ $X2=-0.19 $Y2=1.66
cc_395 N_A_493_368#_c_571_n N_A_772_368#_c_726_n 0.0188586f $X=4.345 $Y=2.275
+ $X2=0 $Y2=0
cc_396 N_A_493_368#_M1008_s N_A_772_368#_c_712_n 0.00287371f $X=4.36 $Y=1.84
+ $X2=0 $Y2=0
cc_397 N_A_493_368#_c_571_n N_A_772_368#_c_712_n 0.00347925f $X=4.345 $Y=2.275
+ $X2=0 $Y2=0
cc_398 N_A_493_368#_c_555_n N_A_772_368#_c_712_n 0.0202301f $X=4.51 $Y=2.275
+ $X2=0 $Y2=0
cc_399 N_A_493_368#_c_553_n N_A_772_368#_c_713_n 0.0125323f $X=3.395 $Y=2.99
+ $X2=0 $Y2=0
cc_400 N_A_493_368#_c_555_n N_A_985_368#_c_740_n 0.036653f $X=4.51 $Y=2.275
+ $X2=0 $Y2=0
cc_401 N_Y_c_609_n N_A_772_368#_M1005_d 0.00510366f $X=4.115 $Y=1.935 $X2=-0.19
+ $Y2=-0.245
cc_402 N_Y_c_606_n N_A_772_368#_M1005_d 9.64364e-19 $X=4.285 $Y=1.665 $X2=-0.19
+ $Y2=-0.245
cc_403 N_Y_c_606_n N_A_985_368#_c_739_n 0.00575161f $X=4.285 $Y=1.665 $X2=0
+ $Y2=0
cc_404 N_Y_c_608_n N_VGND_M1010_s 0.00873456f $X=3.955 $Y=0.755 $X2=0 $Y2=0
cc_405 N_Y_c_597_n N_VGND_M1011_d 0.00250873f $X=4.965 $Y=1.095 $X2=0 $Y2=0
cc_406 N_Y_c_599_n N_VGND_M1019_d 0.00994502f $X=6.325 $Y=1.095 $X2=0 $Y2=0
cc_407 N_Y_c_608_n N_VGND_c_784_n 0.0285862f $X=3.955 $Y=0.755 $X2=0 $Y2=0
cc_408 N_Y_c_601_n N_VGND_c_784_n 0.00615024f $X=3.055 $Y=0.675 $X2=0 $Y2=0
cc_409 N_Y_c_602_n N_VGND_c_784_n 0.00615024f $X=4.12 $Y=0.515 $X2=0 $Y2=0
cc_410 N_Y_c_597_n N_VGND_c_785_n 0.0209867f $X=4.965 $Y=1.095 $X2=0 $Y2=0
cc_411 N_Y_c_598_n N_VGND_c_785_n 0.0182902f $X=5.05 $Y=0.515 $X2=0 $Y2=0
cc_412 N_Y_c_602_n N_VGND_c_785_n 0.0191765f $X=4.12 $Y=0.515 $X2=0 $Y2=0
cc_413 N_Y_c_599_n N_VGND_c_787_n 0.00517071f $X=6.325 $Y=1.095 $X2=0 $Y2=0
cc_414 N_Y_c_600_n N_VGND_c_787_n 0.0243832f $X=6.49 $Y=0.515 $X2=0 $Y2=0
cc_415 N_Y_c_601_n N_VGND_c_788_n 0.00762189f $X=3.055 $Y=0.675 $X2=0 $Y2=0
cc_416 N_Y_c_608_n N_VGND_c_790_n 0.0023667f $X=3.955 $Y=0.755 $X2=0 $Y2=0
cc_417 N_Y_c_601_n N_VGND_c_790_n 0.0141563f $X=3.055 $Y=0.675 $X2=0 $Y2=0
cc_418 N_Y_c_608_n N_VGND_c_791_n 0.0023667f $X=3.955 $Y=0.755 $X2=0 $Y2=0
cc_419 N_Y_c_602_n N_VGND_c_791_n 0.0144922f $X=4.12 $Y=0.515 $X2=0 $Y2=0
cc_420 N_Y_c_598_n N_VGND_c_792_n 0.0109942f $X=5.05 $Y=0.515 $X2=0 $Y2=0
cc_421 N_Y_c_600_n N_VGND_c_793_n 0.011066f $X=6.49 $Y=0.515 $X2=0 $Y2=0
cc_422 N_Y_c_598_n N_VGND_c_796_n 0.0185022f $X=5.05 $Y=0.515 $X2=0 $Y2=0
cc_423 N_Y_c_599_n N_VGND_c_796_n 0.0570323f $X=6.325 $Y=1.095 $X2=0 $Y2=0
cc_424 N_Y_c_600_n N_VGND_c_796_n 0.0183526f $X=6.49 $Y=0.515 $X2=0 $Y2=0
cc_425 N_Y_c_608_n N_VGND_c_797_n 0.0104088f $X=3.955 $Y=0.755 $X2=0 $Y2=0
cc_426 N_Y_c_598_n N_VGND_c_797_n 0.00904371f $X=5.05 $Y=0.515 $X2=0 $Y2=0
cc_427 N_Y_c_600_n N_VGND_c_797_n 0.00915947f $X=6.49 $Y=0.515 $X2=0 $Y2=0
cc_428 N_Y_c_601_n N_VGND_c_797_n 0.0117515f $X=3.055 $Y=0.675 $X2=0 $Y2=0
cc_429 N_Y_c_602_n N_VGND_c_797_n 0.0118826f $X=4.12 $Y=0.515 $X2=0 $Y2=0
cc_430 N_A_772_368#_c_712_n N_A_985_368#_M1009_s 0.00308328f $X=5.355 $Y=2.99
+ $X2=-0.19 $Y2=1.66
cc_431 N_A_772_368#_c_712_n N_A_985_368#_c_740_n 0.018931f $X=5.355 $Y=2.99
+ $X2=0 $Y2=0
cc_432 N_A_772_368#_c_718_n N_A_985_368#_c_740_n 0.0298377f $X=5.52 $Y=2.455
+ $X2=0 $Y2=0
cc_433 N_A_772_368#_M1009_d N_A_985_368#_c_749_n 0.00359365f $X=5.37 $Y=1.84
+ $X2=0 $Y2=0
cc_434 N_A_772_368#_c_718_n N_A_985_368#_c_749_n 0.0171813f $X=5.52 $Y=2.455
+ $X2=0 $Y2=0
cc_435 N_A_772_368#_c_712_n N_A_985_368#_c_741_n 0.00395311f $X=5.355 $Y=2.99
+ $X2=0 $Y2=0
