* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
X0 VPWR a_310_392# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X1 a_310_392# B2 a_41_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 VGND B2 a_27_74# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X3 VPWR B1 a_41_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 a_476_48# A2_N a_835_94# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X5 a_41_392# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 a_835_94# A1_N VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X7 VGND a_310_392# X VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X8 X a_310_392# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X9 a_310_392# a_476_48# a_27_74# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X10 VGND B1 a_27_74# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X11 a_27_74# a_476_48# a_310_392# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X12 a_27_74# B2 VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X13 VPWR a_476_48# a_310_392# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X14 X a_310_392# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X15 a_41_392# B2 a_310_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 a_476_48# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X17 VGND a_310_392# X VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X18 X a_310_392# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X19 VPWR A2_N a_476_48# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X20 VPWR a_310_392# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X21 X a_310_392# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X22 a_27_74# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X23 a_310_392# a_476_48# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
.ends
