* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__ha_1 A B VGND VNB VPB VPWR COUT SUM
M1000 a_695_119# B a_239_294# VNB nshort w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=1.824e+11p ps=1.85e+06u
M1001 VPWR A a_239_294# VPB phighvt w=840000u l=150000u
+  ad=1.732e+12p pd=1.002e+07u as=2.52e+11p ps=2.28e+06u
M1002 a_83_260# a_239_294# VPWR VPB phighvt w=840000u l=150000u
+  ad=3.406e+11p pd=2.71e+06u as=0p ps=0u
M1003 a_386_392# B a_83_260# VPB phighvt w=1e+06u l=150000u
+  ad=4.2e+11p pd=2.84e+06u as=0p ps=0u
M1004 COUT a_239_294# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=0p ps=0u
M1005 COUT a_239_294# VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=6.95225e+11p ps=6.36e+06u
M1006 VPWR a_83_260# SUM VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.304e+11p ps=2.83e+06u
M1007 a_305_130# a_239_294# a_83_260# VNB nshort w=640000u l=150000u
+  ad=3.616e+11p pd=3.69e+06u as=1.726e+11p ps=1.85e+06u
M1008 VGND B a_305_130# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND A a_695_119# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_239_294# B VPWR VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND a_83_260# SUM VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1012 VPWR A a_386_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_305_130# A VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
