* File: sky130_fd_sc_ls__sdlclkp_2.pex.spice
* Created: Wed Sep  2 11:28:56 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__SDLCLKP_2%SCE 2 5 7 9 10 13 14
r32 13 15 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=0.402 $Y=1.455
+ $X2=0.402 $Y2=1.29
r33 13 14 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.385
+ $Y=1.455 $X2=0.385 $Y2=1.455
r34 10 14 2.58853 $w=6.68e-07 $l=1.45e-07 $layer=LI1_cond $X=0.24 $Y=1.625
+ $X2=0.385 $Y2=1.625
r35 7 9 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.495 $Y=2.045
+ $X2=0.495 $Y2=2.54
r36 5 15 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=0.495 $Y=0.835
+ $X2=0.495 $Y2=1.29
r37 2 7 42.0569 $w=3.06e-07 $l=3.10032e-07 $layer=POLY_cond $X=0.402 $Y=1.778
+ $X2=0.495 $Y2=2.045
r38 1 13 2.68759 $w=3.65e-07 $l=1.7e-08 $layer=POLY_cond $X=0.402 $Y=1.472
+ $X2=0.402 $Y2=1.455
r39 1 2 48.3767 $w=3.65e-07 $l=3.06e-07 $layer=POLY_cond $X=0.402 $Y=1.472
+ $X2=0.402 $Y2=1.778
.ends

.subckt PM_SKY130_FD_SC_LS__SDLCLKP_2%GATE 1 3 6 8 12
r38 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.96
+ $Y=1.795 $X2=0.96 $Y2=1.795
r39 8 12 5.68433 $w=5.03e-07 $l=2.4e-07 $layer=LI1_cond $X=1.047 $Y=2.035
+ $X2=1.047 $Y2=1.795
r40 4 11 38.5562 $w=2.99e-07 $l=1.81659e-07 $layer=POLY_cond $X=0.925 $Y=1.63
+ $X2=0.96 $Y2=1.795
r41 4 6 407.649 $w=1.5e-07 $l=7.95e-07 $layer=POLY_cond $X=0.925 $Y=1.63
+ $X2=0.925 $Y2=0.835
r42 1 11 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=0.885 $Y=2.045
+ $X2=0.96 $Y2=1.795
r43 1 3 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.885 $Y=2.045
+ $X2=0.885 $Y2=2.54
.ends

.subckt PM_SKY130_FD_SC_LS__SDLCLKP_2%A_318_74# 1 2 7 9 12 15 16 21 27 29 35
c84 35 0 1.42669e-19 $X=2.94 $Y=1.507
c85 29 0 4.32489e-20 $X=2.855 $Y=1.55
c86 12 0 3.10502e-20 $X=3.35 $Y=0.615
r87 30 35 11.349 $w=3.61e-07 $l=8.5e-08 $layer=POLY_cond $X=2.855 $Y=1.507
+ $X2=2.94 $Y2=1.507
r88 29 32 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=2.855 $Y=1.55 $X2=2.855
+ $Y2=1.63
r89 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.855
+ $Y=1.55 $X2=2.855 $Y2=1.55
r90 26 27 10.1887 $w=6.03e-07 $l=1.65e-07 $layer=LI1_cond $X=2.175 $Y=1.847
+ $X2=2.34 $Y2=1.847
r91 19 21 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.73 $Y=0.965
+ $X2=1.895 $Y2=0.965
r92 16 32 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.69 $Y=1.63
+ $X2=2.855 $Y2=1.63
r93 16 27 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=2.69 $Y=1.63
+ $X2=2.34 $Y2=1.63
r94 15 26 5.53557 $w=6.03e-07 $l=2.8e-07 $layer=LI1_cond $X=1.895 $Y=1.847
+ $X2=2.175 $Y2=1.847
r95 14 21 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.895 $Y=1.05
+ $X2=1.895 $Y2=0.965
r96 14 15 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=1.895 $Y=1.05
+ $X2=1.895 $Y2=1.545
r97 10 35 54.7424 $w=3.61e-07 $l=5.44077e-07 $layer=POLY_cond $X=3.35 $Y=1.195
+ $X2=2.94 $Y2=1.507
r98 10 12 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.35 $Y=1.195
+ $X2=3.35 $Y2=0.615
r99 7 35 23.3725 $w=1.5e-07 $l=3.13e-07 $layer=POLY_cond $X=2.94 $Y=1.82
+ $X2=2.94 $Y2=1.507
r100 7 9 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.94 $Y=1.82 $X2=2.94
+ $Y2=2.315
r101 2 26 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.025
+ $Y=1.84 $X2=2.175 $Y2=1.985
r102 1 19 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=1.59
+ $Y=0.37 $X2=1.73 $Y2=0.965
.ends

.subckt PM_SKY130_FD_SC_LS__SDLCLKP_2%A_288_48# 1 2 7 9 10 11 13 14 15 16 19 20
+ 21 22 23 24 26 27 28 29 31 33 34 35 37 38 39 41 42 43 47 51 54 56 57
c168 57 0 1.08887e-19 $X=5.152 $Y=1.72
c169 47 0 1.44698e-19 $X=5.195 $Y=0.515
c170 43 0 1.9008e-19 $X=4.38 $Y=0.34
c171 42 0 9.22391e-20 $X=4.995 $Y=0.34
c172 33 0 3.10502e-20 $X=2.63 $Y=1.03
r173 56 57 8.46257 $w=3.13e-07 $l=1.65e-07 $layer=LI1_cond $X=5.152 $Y=1.885
+ $X2=5.152 $Y2=1.72
r174 54 57 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=5.08 $Y=1.01
+ $X2=5.08 $Y2=1.72
r175 51 53 14.6122 $w=2.63e-07 $l=3.15e-07 $layer=LI1_cond $X=2.315 $Y=1.195
+ $X2=2.63 $Y2=1.195
r176 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.315
+ $Y=1.195 $X2=2.315 $Y2=1.195
r177 45 54 9.06106 $w=3.63e-07 $l=1.82e-07 $layer=LI1_cond $X=5.177 $Y=0.828
+ $X2=5.177 $Y2=1.01
r178 45 47 9.88259 $w=3.63e-07 $l=3.13e-07 $layer=LI1_cond $X=5.177 $Y=0.828
+ $X2=5.177 $Y2=0.515
r179 44 47 2.84164 $w=3.63e-07 $l=9e-08 $layer=LI1_cond $X=5.177 $Y=0.425
+ $X2=5.177 $Y2=0.515
r180 42 44 8.06639 $w=1.7e-07 $l=2.2044e-07 $layer=LI1_cond $X=4.995 $Y=0.34
+ $X2=5.177 $Y2=0.425
r181 42 43 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=4.995 $Y=0.34
+ $X2=4.38 $Y2=0.34
r182 40 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.295 $Y=0.425
+ $X2=4.38 $Y2=0.34
r183 40 41 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=4.295 $Y=0.425
+ $X2=4.295 $Y2=0.905
r184 38 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.21 $Y=0.99
+ $X2=4.295 $Y2=0.905
r185 38 39 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=4.21 $Y=0.99
+ $X2=3.7 $Y2=0.99
r186 37 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.615 $Y=0.905
+ $X2=3.7 $Y2=0.99
r187 36 37 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=3.615 $Y=0.425
+ $X2=3.615 $Y2=0.905
r188 34 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.53 $Y=0.34
+ $X2=3.615 $Y2=0.425
r189 34 35 53.1711 $w=1.68e-07 $l=8.15e-07 $layer=LI1_cond $X=3.53 $Y=0.34
+ $X2=2.715 $Y2=0.34
r190 33 53 3.29066 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.63 $Y=1.03
+ $X2=2.63 $Y2=1.195
r191 32 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.63 $Y=0.425
+ $X2=2.715 $Y2=0.34
r192 32 33 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=2.63 $Y=0.425
+ $X2=2.63 $Y2=1.03
r193 29 31 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.465 $Y=2.75
+ $X2=3.465 $Y2=2.465
r194 27 29 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.465 $Y=2.84
+ $X2=3.465 $Y2=2.75
r195 27 28 91.3468 $w=1.8e-07 $l=2.35e-07 $layer=POLY_cond $X=3.465 $Y=2.84
+ $X2=3.465 $Y2=3.075
r196 24 26 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=2.825 $Y=0.995
+ $X2=2.825 $Y2=0.645
r197 23 52 39.0383 $w=2.64e-07 $l=2.11849e-07 $layer=POLY_cond $X=2.48 $Y=1.07
+ $X2=2.315 $Y2=1.177
r198 22 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.75 $Y=1.07
+ $X2=2.825 $Y2=0.995
r199 22 23 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.75 $Y=1.07
+ $X2=2.48 $Y2=1.07
r200 20 28 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=3.375 $Y=3.15
+ $X2=3.465 $Y2=3.075
r201 20 21 684.543 $w=1.5e-07 $l=1.335e-06 $layer=POLY_cond $X=3.375 $Y=3.15
+ $X2=2.04 $Y2=3.15
r202 17 19 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.95 $Y=2.755
+ $X2=1.95 $Y2=2.26
r203 16 19 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.95 $Y=1.765
+ $X2=1.95 $Y2=2.26
r204 15 21 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=1.95 $Y=3.075
+ $X2=2.04 $Y2=3.15
r205 14 17 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.95 $Y=2.845
+ $X2=1.95 $Y2=2.755
r206 14 15 89.4032 $w=1.8e-07 $l=2.3e-07 $layer=POLY_cond $X=1.95 $Y=2.845
+ $X2=1.95 $Y2=3.075
r207 13 16 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.95 $Y=1.675
+ $X2=1.95 $Y2=1.765
r208 12 52 66.6402 $w=2.64e-07 $l=4.47236e-07 $layer=POLY_cond $X=1.95 $Y=1.36
+ $X2=2.315 $Y2=1.177
r209 12 13 122.444 $w=1.8e-07 $l=3.15e-07 $layer=POLY_cond $X=1.95 $Y=1.36
+ $X2=1.95 $Y2=1.675
r210 10 12 25.3451 $w=2.64e-07 $l=1.21861e-07 $layer=POLY_cond $X=1.86 $Y=1.285
+ $X2=1.95 $Y2=1.36
r211 10 11 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=1.86 $Y=1.285
+ $X2=1.59 $Y2=1.285
r212 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.515 $Y=1.21
+ $X2=1.59 $Y2=1.285
r213 7 9 151.027 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=1.515 $Y=1.21
+ $X2=1.515 $Y2=0.74
r214 2 56 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=5.01
+ $Y=1.74 $X2=5.145 $Y2=1.885
r215 1 47 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=5.05
+ $Y=0.37 $X2=5.195 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__SDLCLKP_2%A_706_317# 1 2 9 12 13 15 18 20 22 23 26
+ 31 35 38 39 42 43 45 49 54 55 56 60
c135 49 0 1.42669e-19 $X=3.695 $Y=1.75
c136 42 0 1.37146e-19 $X=5.92 $Y=2.22
c137 20 0 1.93704e-19 $X=6.565 $Y=1.795
c138 9 0 4.32489e-20 $X=3.74 $Y=0.615
r139 59 60 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=3.74 $Y=1.75
+ $X2=3.855 $Y2=1.75
r140 50 59 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=3.695 $Y=1.75
+ $X2=3.74 $Y2=1.75
r141 49 52 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=3.695 $Y=1.75
+ $X2=3.695 $Y2=1.84
r142 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.695
+ $Y=1.75 $X2=3.695 $Y2=1.75
r143 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.365
+ $Y=1.465 $X2=6.365 $Y2=1.465
r144 43 45 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=6.005 $Y=1.465
+ $X2=6.365 $Y2=1.465
r145 41 43 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.92 $Y=1.63
+ $X2=6.005 $Y2=1.465
r146 41 42 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=5.92 $Y=1.63
+ $X2=5.92 $Y2=2.22
r147 40 55 4.39717 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=4.825 $Y=2.305
+ $X2=4.632 $Y2=2.305
r148 39 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.835 $Y=2.305
+ $X2=5.92 $Y2=2.22
r149 39 40 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=5.835 $Y=2.305
+ $X2=4.825 $Y2=2.305
r150 38 54 3.37808 $w=2.77e-07 $l=1.44375e-07 $layer=LI1_cond $X=4.74 $Y=1.755
+ $X2=4.632 $Y2=1.84
r151 38 56 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.74 $Y=1.755
+ $X2=4.74 $Y2=1.075
r152 33 56 7.41084 $w=2.73e-07 $l=1.37e-07 $layer=LI1_cond $X=4.687 $Y=0.938
+ $X2=4.687 $Y2=1.075
r153 33 35 4.31642 $w=2.73e-07 $l=1.03e-07 $layer=LI1_cond $X=4.687 $Y=0.938
+ $X2=4.687 $Y2=0.835
r154 29 55 2.50573 $w=3.85e-07 $l=8.5e-08 $layer=LI1_cond $X=4.632 $Y=2.39
+ $X2=4.632 $Y2=2.305
r155 29 31 10.9258 $w=3.83e-07 $l=3.65e-07 $layer=LI1_cond $X=4.632 $Y=2.39
+ $X2=4.632 $Y2=2.755
r156 28 54 3.37808 $w=2.77e-07 $l=8.5e-08 $layer=LI1_cond $X=4.632 $Y=1.925
+ $X2=4.632 $Y2=1.84
r157 26 55 2.50573 $w=3.85e-07 $l=8.5e-08 $layer=LI1_cond $X=4.632 $Y=2.22
+ $X2=4.632 $Y2=2.305
r158 26 28 8.83041 $w=3.83e-07 $l=2.95e-07 $layer=LI1_cond $X=4.632 $Y=2.22
+ $X2=4.632 $Y2=1.925
r159 24 52 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.86 $Y=1.84
+ $X2=3.695 $Y2=1.84
r160 23 54 3.15366 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=4.44 $Y=1.84
+ $X2=4.632 $Y2=1.84
r161 23 24 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=4.44 $Y=1.84
+ $X2=3.86 $Y2=1.84
r162 20 46 60.8611 $w=3.63e-07 $l=3.92989e-07 $layer=POLY_cond $X=6.565 $Y=1.795
+ $X2=6.427 $Y2=1.465
r163 20 22 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.565 $Y=1.795
+ $X2=6.565 $Y2=2.37
r164 16 46 38.952 $w=3.63e-07 $l=2.28703e-07 $layer=POLY_cond $X=6.275 $Y=1.3
+ $X2=6.427 $Y2=1.465
r165 16 18 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=6.275 $Y=1.3
+ $X2=6.275 $Y2=0.74
r166 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.855 $Y=2.18
+ $X2=3.855 $Y2=2.465
r167 12 13 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.855 $Y=2.09
+ $X2=3.855 $Y2=2.18
r168 11 60 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.855 $Y=1.915
+ $X2=3.855 $Y2=1.75
r169 11 12 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=3.855 $Y=1.915
+ $X2=3.855 $Y2=2.09
r170 7 59 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.74 $Y=1.585
+ $X2=3.74 $Y2=1.75
r171 7 9 497.383 $w=1.5e-07 $l=9.7e-07 $layer=POLY_cond $X=3.74 $Y=1.585
+ $X2=3.74 $Y2=0.615
r172 2 31 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=4.455
+ $Y=1.78 $X2=4.605 $Y2=2.755
r173 2 28 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=4.455
+ $Y=1.78 $X2=4.605 $Y2=1.925
r174 1 35 182 $w=1.7e-07 $l=4.95076e-07 $layer=licon1_NDIFF $count=1 $X=4.495
+ $Y=0.405 $X2=4.635 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_LS__SDLCLKP_2%A_580_74# 1 2 7 9 10 12 13 18 21 24 25 27
+ 28
r84 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.32
+ $Y=1.42 $X2=4.32 $Y2=1.42
r85 28 31 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=4.32 $Y=1.33 $X2=4.32
+ $Y2=1.42
r86 24 25 10.5918 $w=3.58e-07 $l=2.3e-07 $layer=LI1_cond $X=3.18 $Y=2.465
+ $X2=3.18 $Y2=2.235
r87 22 27 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.36 $Y=1.33
+ $X2=3.275 $Y2=1.33
r88 21 28 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.155 $Y=1.33
+ $X2=4.32 $Y2=1.33
r89 21 22 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=4.155 $Y=1.33
+ $X2=3.36 $Y2=1.33
r90 19 27 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.275 $Y=1.415
+ $X2=3.275 $Y2=1.33
r91 19 25 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=3.275 $Y=1.415
+ $X2=3.275 $Y2=2.235
r92 18 27 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.275 $Y=1.245
+ $X2=3.275 $Y2=1.33
r93 17 18 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=3.275 $Y=0.845
+ $X2=3.275 $Y2=1.245
r94 13 17 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.19 $Y=0.72
+ $X2=3.275 $Y2=0.845
r95 13 15 6.45368 $w=2.48e-07 $l=1.4e-07 $layer=LI1_cond $X=3.19 $Y=0.72
+ $X2=3.05 $Y2=0.72
r96 10 32 38.5662 $w=2.97e-07 $l=2.07123e-07 $layer=POLY_cond $X=4.42 $Y=1.255
+ $X2=4.325 $Y2=1.42
r97 10 12 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.42 $Y=1.255
+ $X2=4.42 $Y2=0.775
r98 7 32 58.0409 $w=2.97e-07 $l=3.11288e-07 $layer=POLY_cond $X=4.38 $Y=1.705
+ $X2=4.325 $Y2=1.42
r99 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.38 $Y=1.705
+ $X2=4.38 $Y2=2.34
r100 2 24 600 $w=1.7e-07 $l=6.40625e-07 $layer=licon1_PDIFF $count=1 $X=3.015
+ $Y=1.895 $X2=3.165 $Y2=2.465
r101 1 15 182 $w=1.7e-07 $l=3.77624e-07 $layer=licon1_NDIFF $count=1 $X=2.9
+ $Y=0.37 $X2=3.05 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_LS__SDLCLKP_2%CLK 1 3 4 6 7 8 9 11 12 14 15
c56 15 0 1.1118e-19 $X=5.52 $Y=1.295
c57 12 0 2.36937e-19 $X=5.915 $Y=1.22
c58 7 0 1.37146e-19 $X=5.9 $Y=1.55
c59 1 0 1.08887e-19 $X=5.37 $Y=1.665
r60 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.5
+ $Y=1.385 $X2=5.5 $Y2=1.385
r61 18 20 12.0836 $w=3.59e-07 $l=9e-08 $layer=POLY_cond $X=5.41 $Y=1.442 $X2=5.5
+ $Y2=1.442
r62 17 18 5.37047 $w=3.59e-07 $l=4e-08 $layer=POLY_cond $X=5.37 $Y=1.442
+ $X2=5.41 $Y2=1.442
r63 15 21 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=5.5 $Y=1.295 $X2=5.5
+ $Y2=1.385
r64 12 23 23.2387 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=5.915 $Y=1.22
+ $X2=5.915 $Y2=1.442
r65 12 14 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.915 $Y=1.22
+ $X2=5.915 $Y2=0.74
r66 9 11 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.9 $Y=1.795 $X2=5.9
+ $Y2=2.37
r67 8 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.9 $Y=1.705 $X2=5.9
+ $Y2=1.795
r68 7 23 2.01393 $w=3.59e-07 $l=1.5e-08 $layer=POLY_cond $X=5.9 $Y=1.442
+ $X2=5.915 $Y2=1.442
r69 7 20 53.7047 $w=3.59e-07 $l=4e-07 $layer=POLY_cond $X=5.9 $Y=1.442 $X2=5.5
+ $Y2=1.442
r70 7 8 60.25 $w=1.8e-07 $l=1.55e-07 $layer=POLY_cond $X=5.9 $Y=1.55 $X2=5.9
+ $Y2=1.705
r71 4 18 23.2387 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=5.41 $Y=1.22
+ $X2=5.41 $Y2=1.442
r72 4 6 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.41 $Y=1.22 $X2=5.41
+ $Y2=0.74
r73 1 17 23.2387 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=5.37 $Y=1.665
+ $X2=5.37 $Y2=1.442
r74 1 3 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=5.37 $Y=1.665 $X2=5.37
+ $Y2=2.16
.ends

.subckt PM_SKY130_FD_SC_LS__SDLCLKP_2%A_1195_374# 1 2 7 9 12 14 16 19 23 29 31
+ 32 33 34 38 40 42 47
c87 38 0 8.25245e-20 $X=6.955 $Y=1.8
r88 47 48 9.66578 $w=3.74e-07 $l=7.5e-08 $layer=POLY_cond $X=7.6 $Y=1.532
+ $X2=7.675 $Y2=1.532
r89 46 47 45.7513 $w=3.74e-07 $l=3.55e-07 $layer=POLY_cond $X=7.245 $Y=1.532
+ $X2=7.6 $Y2=1.532
r90 45 46 12.2433 $w=3.74e-07 $l=9.5e-08 $layer=POLY_cond $X=7.15 $Y=1.532
+ $X2=7.245 $Y2=1.532
r91 41 45 11.5989 $w=3.74e-07 $l=9e-08 $layer=POLY_cond $X=7.06 $Y=1.532
+ $X2=7.15 $Y2=1.532
r92 40 43 8.49906 $w=3.53e-07 $l=1.65e-07 $layer=LI1_cond $X=7.047 $Y=1.465
+ $X2=7.047 $Y2=1.63
r93 40 42 8.49906 $w=3.53e-07 $l=1.65e-07 $layer=LI1_cond $X=7.047 $Y=1.465
+ $X2=7.047 $Y2=1.3
r94 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.06
+ $Y=1.465 $X2=7.06 $Y2=1.465
r95 38 43 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=6.955 $Y=1.8
+ $X2=6.955 $Y2=1.63
r96 35 42 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=6.955 $Y=1.13
+ $X2=6.955 $Y2=1.3
r97 33 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.87 $Y=1.045
+ $X2=6.955 $Y2=1.13
r98 33 34 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=6.87 $Y=1.045
+ $X2=6.655 $Y2=1.045
r99 31 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.87 $Y=1.885
+ $X2=6.955 $Y2=1.8
r100 31 32 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=6.87 $Y=1.885
+ $X2=6.505 $Y2=1.885
r101 27 34 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.49 $Y=0.96
+ $X2=6.655 $Y2=1.045
r102 27 29 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=6.49 $Y=0.96
+ $X2=6.49 $Y2=0.515
r103 23 25 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=6.34 $Y=2.015
+ $X2=6.34 $Y2=2.725
r104 21 32 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.34 $Y=1.97
+ $X2=6.505 $Y2=1.885
r105 21 23 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=6.34 $Y=1.97
+ $X2=6.34 $Y2=2.015
r106 17 48 24.2268 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=7.675 $Y=1.3
+ $X2=7.675 $Y2=1.532
r107 17 19 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=7.675 $Y=1.3
+ $X2=7.675 $Y2=0.74
r108 14 47 24.2268 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=7.6 $Y=1.765
+ $X2=7.6 $Y2=1.532
r109 14 16 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.6 $Y=1.765
+ $X2=7.6 $Y2=2.4
r110 10 46 24.2268 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=7.245 $Y=1.3
+ $X2=7.245 $Y2=1.532
r111 10 12 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=7.245 $Y=1.3
+ $X2=7.245 $Y2=0.74
r112 7 45 24.2268 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=7.15 $Y=1.765
+ $X2=7.15 $Y2=1.532
r113 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.15 $Y=1.765
+ $X2=7.15 $Y2=2.4
r114 2 25 400 $w=1.7e-07 $l=1.02132e-06 $layer=licon1_PDIFF $count=1 $X=5.975
+ $Y=1.87 $X2=6.34 $Y2=2.725
r115 2 23 400 $w=1.7e-07 $l=4.31451e-07 $layer=licon1_PDIFF $count=1 $X=5.975
+ $Y=1.87 $X2=6.34 $Y2=2.015
r116 1 29 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.35
+ $Y=0.37 $X2=6.49 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__SDLCLKP_2%VPWR 1 2 3 4 5 6 19 21 25 29 35 39 43 45
+ 50 51 52 54 59 67 76 84 87 90 94
r95 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r96 90 91 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r97 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r98 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r99 79 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r100 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r101 76 93 3.94754 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=7.74 $Y=3.33
+ $X2=7.95 $Y2=3.33
r102 76 78 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=7.74 $Y=3.33 $X2=7.44
+ $Y2=3.33
r103 75 79 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=7.44 $Y2=3.33
r104 75 91 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=5.52 $Y2=3.33
r105 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r106 72 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.84 $Y=3.33
+ $X2=5.675 $Y2=3.33
r107 72 74 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=5.84 $Y=3.33
+ $X2=6.48 $Y2=3.33
r108 71 91 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r109 70 71 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r110 68 87 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.24 $Y=3.33
+ $X2=4.115 $Y2=3.33
r111 68 70 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=4.24 $Y=3.33
+ $X2=4.56 $Y2=3.33
r112 67 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.51 $Y=3.33
+ $X2=5.675 $Y2=3.33
r113 67 70 61.9786 $w=1.68e-07 $l=9.5e-07 $layer=LI1_cond $X=5.51 $Y=3.33
+ $X2=4.56 $Y2=3.33
r114 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r115 63 66 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.6 $Y2=3.33
r116 63 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r117 62 65 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=3.6 $Y2=3.33
r118 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r119 60 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.815 $Y=3.33
+ $X2=1.65 $Y2=3.33
r120 60 62 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.815 $Y=3.33
+ $X2=2.16 $Y2=3.33
r121 59 87 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.99 $Y=3.33
+ $X2=4.115 $Y2=3.33
r122 59 65 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=3.99 $Y=3.33
+ $X2=3.6 $Y2=3.33
r123 58 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r124 58 82 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.24 $Y2=3.33
r125 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r126 55 81 4.75569 $w=1.7e-07 $l=2.18e-07 $layer=LI1_cond $X=0.435 $Y=3.33
+ $X2=0.217 $Y2=3.33
r127 55 57 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=0.435 $Y=3.33
+ $X2=1.2 $Y2=3.33
r128 54 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.485 $Y=3.33
+ $X2=1.65 $Y2=3.33
r129 54 57 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.485 $Y=3.33
+ $X2=1.2 $Y2=3.33
r130 52 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r131 52 66 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r132 52 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r133 50 74 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=6.71 $Y=3.33
+ $X2=6.48 $Y2=3.33
r134 50 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.71 $Y=3.33
+ $X2=6.875 $Y2=3.33
r135 49 78 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=7.04 $Y=3.33 $X2=7.44
+ $Y2=3.33
r136 49 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.04 $Y=3.33
+ $X2=6.875 $Y2=3.33
r137 45 48 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=7.865 $Y=1.985
+ $X2=7.865 $Y2=2.815
r138 43 93 3.19563 $w=2.5e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.865 $Y=3.245
+ $X2=7.95 $Y2=3.33
r139 43 48 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=7.865 $Y=3.245
+ $X2=7.865 $Y2=2.815
r140 39 42 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=6.875 $Y=2.305
+ $X2=6.875 $Y2=2.815
r141 37 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.875 $Y=3.245
+ $X2=6.875 $Y2=3.33
r142 37 42 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=6.875 $Y=3.245
+ $X2=6.875 $Y2=2.815
r143 33 90 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.675 $Y=3.245
+ $X2=5.675 $Y2=3.33
r144 33 35 18.1597 $w=3.28e-07 $l=5.2e-07 $layer=LI1_cond $X=5.675 $Y=3.245
+ $X2=5.675 $Y2=2.725
r145 29 32 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=4.115 $Y=2.26
+ $X2=4.115 $Y2=2.755
r146 27 87 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.115 $Y=3.245
+ $X2=4.115 $Y2=3.33
r147 27 32 22.5879 $w=2.48e-07 $l=4.9e-07 $layer=LI1_cond $X=4.115 $Y=3.245
+ $X2=4.115 $Y2=2.755
r148 23 84 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.65 $Y=3.245
+ $X2=1.65 $Y2=3.33
r149 23 25 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=1.65 $Y=3.245
+ $X2=1.65 $Y2=2.825
r150 19 81 3.01048 $w=3.3e-07 $l=1.08305e-07 $layer=LI1_cond $X=0.27 $Y=3.245
+ $X2=0.217 $Y2=3.33
r151 19 21 33.1764 $w=3.28e-07 $l=9.5e-07 $layer=LI1_cond $X=0.27 $Y=3.245
+ $X2=0.27 $Y2=2.295
r152 6 48 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=7.675
+ $Y=1.84 $X2=7.825 $Y2=2.815
r153 6 45 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=7.675
+ $Y=1.84 $X2=7.825 $Y2=1.985
r154 5 42 600 $w=1.7e-07 $l=1.05598e-06 $layer=licon1_PDIFF $count=1 $X=6.64
+ $Y=1.87 $X2=6.875 $Y2=2.815
r155 5 39 600 $w=1.7e-07 $l=5.39861e-07 $layer=licon1_PDIFF $count=1 $X=6.64
+ $Y=1.87 $X2=6.875 $Y2=2.305
r156 4 35 600 $w=1.7e-07 $l=1.09397e-06 $layer=licon1_PDIFF $count=1 $X=5.445
+ $Y=1.74 $X2=5.675 $Y2=2.725
r157 3 32 600 $w=1.7e-07 $l=6.0208e-07 $layer=licon1_PDIFF $count=1 $X=3.93
+ $Y=2.255 $X2=4.155 $Y2=2.755
r158 3 29 600 $w=1.7e-07 $l=2.27486e-07 $layer=licon1_PDIFF $count=1 $X=3.93
+ $Y=2.255 $X2=4.155 $Y2=2.26
r159 2 25 600 $w=1.7e-07 $l=1.05033e-06 $layer=licon1_PDIFF $count=1 $X=1.515
+ $Y=1.84 $X2=1.65 $Y2=2.825
r160 1 21 300 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.12 $X2=0.27 $Y2=2.295
.ends

.subckt PM_SKY130_FD_SC_LS__SDLCLKP_2%A_114_112# 1 2 3 4 14 16 17 18 19 23 26 27
+ 31 35 36 38
r99 38 40 4.37928 $w=2.48e-07 $l=9.5e-08 $layer=LI1_cond $X=2.25 $Y=0.53
+ $X2=2.25 $Y2=0.625
r100 29 31 12.4464 $w=2.48e-07 $l=2.7e-07 $layer=LI1_cond $X=2.675 $Y=2.32
+ $X2=2.675 $Y2=2.05
r101 28 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.64 $Y=2.405
+ $X2=1.555 $Y2=2.405
r102 27 29 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.55 $Y=2.405
+ $X2=2.675 $Y2=2.32
r103 27 28 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=2.55 $Y=2.405
+ $X2=1.64 $Y2=2.405
r104 26 36 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.555 $Y=2.32
+ $X2=1.555 $Y2=2.405
r105 25 26 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=1.555 $Y=1.39
+ $X2=1.555 $Y2=2.32
r106 24 35 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.275 $Y=2.405
+ $X2=1.11 $Y2=2.405
r107 23 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.47 $Y=2.405
+ $X2=1.555 $Y2=2.405
r108 23 24 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=1.47 $Y=2.405
+ $X2=1.275 $Y2=2.405
r109 20 33 2.70854 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=0.89 $Y=1.305
+ $X2=0.72 $Y2=1.305
r110 19 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.47 $Y=1.305
+ $X2=1.555 $Y2=1.39
r111 19 20 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=1.47 $Y=1.305
+ $X2=0.89 $Y2=1.305
r112 17 40 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.125 $Y=0.625
+ $X2=2.25 $Y2=0.625
r113 17 18 80.5722 $w=1.68e-07 $l=1.235e-06 $layer=LI1_cond $X=2.125 $Y=0.625
+ $X2=0.89 $Y2=0.625
r114 14 33 13.8085 $w=3.45e-07 $l=3.58497e-07 $layer=LI1_cond $X=0.717 $Y=0.948
+ $X2=0.72 $Y2=1.305
r115 14 16 3.94169 $w=3.43e-07 $l=1.18e-07 $layer=LI1_cond $X=0.717 $Y=0.948
+ $X2=0.717 $Y2=0.83
r116 13 18 7.89393 $w=1.7e-07 $l=2.11268e-07 $layer=LI1_cond $X=0.717 $Y=0.71
+ $X2=0.89 $Y2=0.625
r117 13 16 4.0085 $w=3.43e-07 $l=1.2e-07 $layer=LI1_cond $X=0.717 $Y=0.71
+ $X2=0.717 $Y2=0.83
r118 4 31 300 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=2 $X=2.58
+ $Y=1.895 $X2=2.715 $Y2=2.05
r119 3 35 300 $w=1.7e-07 $l=3.52101e-07 $layer=licon1_PDIFF $count=2 $X=0.96
+ $Y=2.12 $X2=1.11 $Y2=2.405
r120 2 38 182 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=1 $X=2.145
+ $Y=0.37 $X2=2.29 $Y2=0.53
r121 1 16 182 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.56 $X2=0.71 $Y2=0.83
.ends

.subckt PM_SKY130_FD_SC_LS__SDLCLKP_2%GCLK 1 2 9 13 14 15 16 23 32
r37 21 23 1.2336 $w=3.53e-07 $l=3.8e-08 $layer=LI1_cond $X=7.387 $Y=1.997
+ $X2=7.387 $Y2=2.035
r38 15 16 12.0114 $w=3.53e-07 $l=3.7e-07 $layer=LI1_cond $X=7.387 $Y=2.405
+ $X2=7.387 $Y2=2.775
r39 14 21 0.779116 $w=3.53e-07 $l=2.4e-08 $layer=LI1_cond $X=7.387 $Y=1.973
+ $X2=7.387 $Y2=1.997
r40 14 32 8.1095 $w=3.53e-07 $l=1.53e-07 $layer=LI1_cond $X=7.387 $Y=1.973
+ $X2=7.387 $Y2=1.82
r41 14 15 11.2647 $w=3.53e-07 $l=3.47e-07 $layer=LI1_cond $X=7.387 $Y=2.058
+ $X2=7.387 $Y2=2.405
r42 14 23 0.746653 $w=3.53e-07 $l=2.3e-08 $layer=LI1_cond $X=7.387 $Y=2.058
+ $X2=7.387 $Y2=2.035
r43 13 32 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=7.48 $Y=1.13 $X2=7.48
+ $Y2=1.82
r44 7 13 7.30505 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.46 $Y=0.965
+ $X2=7.46 $Y2=1.13
r45 7 9 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=7.46 $Y=0.965 $X2=7.46
+ $Y2=0.515
r46 2 14 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=7.225
+ $Y=1.84 $X2=7.375 $Y2=1.985
r47 2 16 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=7.225
+ $Y=1.84 $X2=7.375 $Y2=2.815
r48 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.32
+ $Y=0.37 $X2=7.46 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__SDLCLKP_2%VGND 1 2 3 4 5 6 19 21 25 29 33 35 37 40
+ 41 43 44 45 47 65 69 79 85 89
c93 3 0 1.9008e-19 $X=3.815 $Y=0.405
r94 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r95 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r96 79 82 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=1.22 $Y=0 $X2=1.22
+ $Y2=0.285
r97 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r98 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r99 73 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=7.92
+ $Y2=0
r100 73 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=6.96
+ $Y2=0
r101 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r102 70 85 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.115 $Y=0 $X2=6.99
+ $Y2=0
r103 70 72 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=7.115 $Y=0
+ $X2=7.44 $Y2=0
r104 69 88 4.02656 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=7.805 $Y=0
+ $X2=7.982 $Y2=0
r105 69 72 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=7.805 $Y=0
+ $X2=7.44 $Y2=0
r106 68 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6.96
+ $Y2=0
r107 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r108 65 85 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.865 $Y=0 $X2=6.99
+ $Y2=0
r109 65 67 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=6.865 $Y=0
+ $X2=6.48 $Y2=0
r110 64 68 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6.48
+ $Y2=0
r111 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r112 60 63 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=4.08 $Y=0 $X2=5.52
+ $Y2=0
r113 57 58 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r114 55 58 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=1.68 $Y=0 $X2=3.6
+ $Y2=0
r115 55 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r116 54 57 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.68 $Y=0 $X2=3.6
+ $Y2=0
r117 54 55 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.68 $Y=0
+ $X2=1.68 $Y2=0
r118 52 79 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.385 $Y=0 $X2=1.22
+ $Y2=0
r119 52 54 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.385 $Y=0 $X2=1.68
+ $Y2=0
r120 51 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r121 51 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r122 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r123 48 75 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=0
+ $X2=0.182 $Y2=0
r124 48 50 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=0
+ $X2=0.72 $Y2=0
r125 47 79 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.055 $Y=0 $X2=1.22
+ $Y2=0
r126 47 50 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.055 $Y=0
+ $X2=0.72 $Y2=0
r127 45 64 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.08 $Y=0
+ $X2=5.52 $Y2=0
r128 45 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r129 45 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r130 43 63 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=5.53 $Y=0 $X2=5.52
+ $Y2=0
r131 43 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.53 $Y=0 $X2=5.695
+ $Y2=0
r132 42 67 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=5.86 $Y=0 $X2=6.48
+ $Y2=0
r133 42 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.86 $Y=0 $X2=5.695
+ $Y2=0
r134 40 57 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=3.87 $Y=0 $X2=3.6
+ $Y2=0
r135 40 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.87 $Y=0 $X2=3.955
+ $Y2=0
r136 39 60 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=4.04 $Y=0 $X2=4.08
+ $Y2=0
r137 39 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.04 $Y=0 $X2=3.955
+ $Y2=0
r138 35 88 3.1166 $w=2.5e-07 $l=1.07912e-07 $layer=LI1_cond $X=7.93 $Y=0.085
+ $X2=7.982 $Y2=0
r139 35 37 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=7.93 $Y=0.085
+ $X2=7.93 $Y2=0.515
r140 31 85 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.99 $Y=0.085
+ $X2=6.99 $Y2=0
r141 31 33 22.3574 $w=2.48e-07 $l=4.85e-07 $layer=LI1_cond $X=6.99 $Y=0.085
+ $X2=6.99 $Y2=0.57
r142 27 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.695 $Y=0.085
+ $X2=5.695 $Y2=0
r143 27 29 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=5.695 $Y=0.085
+ $X2=5.695 $Y2=0.515
r144 23 41 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.955 $Y=0.085
+ $X2=3.955 $Y2=0
r145 23 25 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=3.955 $Y=0.085
+ $X2=3.955 $Y2=0.56
r146 19 75 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.182 $Y2=0
r147 19 21 34.3428 $w=2.48e-07 $l=7.45e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.24 $Y2=0.83
r148 6 37 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.75
+ $Y=0.37 $X2=7.89 $Y2=0.515
r149 5 33 182 $w=1.7e-07 $l=2.58844e-07 $layer=licon1_NDIFF $count=1 $X=6.895
+ $Y=0.37 $X2=7.03 $Y2=0.57
r150 4 29 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=5.485
+ $Y=0.37 $X2=5.695 $Y2=0.515
r151 3 25 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=3.815
+ $Y=0.405 $X2=3.955 $Y2=0.56
r152 2 82 182 $w=1.7e-07 $l=3.68951e-07 $layer=licon1_NDIFF $count=1 $X=1
+ $Y=0.56 $X2=1.22 $Y2=0.285
r153 1 21 182 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.56 $X2=0.28 $Y2=0.83
.ends

