* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__nand3_4 A B C VGND VNB VPB VPWR Y
X0 a_27_82# B a_456_82# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X1 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X2 a_27_82# A Y VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X3 a_456_82# B a_27_82# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X4 a_456_82# C VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X5 VGND C a_456_82# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X6 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X7 a_456_82# C VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X8 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X9 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X10 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X11 Y A a_27_82# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X12 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X13 a_27_82# A Y VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X14 Y A a_27_82# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X15 a_27_82# B a_456_82# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X16 a_456_82# B a_27_82# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X17 VGND C a_456_82# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
.ends
