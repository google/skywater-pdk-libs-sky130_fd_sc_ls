* NGSPICE file created from sky130_fd_sc_ls__o22ai_1.ext - technology: sky130A

.subckt sky130_fd_sc_ls__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
M1000 a_142_368# B1 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.024e+11p pd=2.78e+06u as=7.952e+11p ps=5.9e+06u
M1001 VGND A2 a_27_74# VNB nshort w=740000u l=150000u
+  ad=3.108e+11p pd=2.32e+06u as=6.808e+11p ps=6.28e+06u
M1002 a_27_74# B2 Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=4.255e+11p ps=2.63e+06u
M1003 a_27_74# A1 VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR A1 a_340_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=4.704e+11p ps=3.08e+06u
M1005 Y B2 a_142_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=4.704e+11p pd=3.08e+06u as=0p ps=0u
M1006 a_340_368# A2 Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y B1 a_27_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

