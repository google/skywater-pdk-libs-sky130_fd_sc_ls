* File: sky130_fd_sc_ls__nor2_4.spice
* Created: Fri Aug 28 13:37:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__nor2_4.pex.spice"
.subckt sky130_fd_sc_ls__nor2_4  VNB VPB A B VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1001 N_VGND_M1001_d N_A_M1001_g N_Y_M1001_s VNB NSHORT L=0.15 W=0.74 AD=0.2294
+ AS=0.4218 PD=2.1 PS=1.88 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2 SB=75003.5
+ A=0.111 P=1.78 MULT=1
MM1003 N_VGND_M1003_d N_A_M1003_g N_Y_M1001_s VNB NSHORT L=0.15 W=0.74 AD=0.1221
+ AS=0.4218 PD=1.07 PS=1.88 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5 SB=75002.2
+ A=0.111 P=1.78 MULT=1
MM1004 N_Y_M1004_d N_B_M1004_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.74 AD=0.111
+ AS=0.1221 PD=1.04 PS=1.07 NRD=3.24 NRS=8.1 M=1 R=4.93333 SA=75002 SB=75001.7
+ A=0.111 P=1.78 MULT=1
MM1006 N_Y_M1004_d N_B_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.74 AD=0.111
+ AS=1.0138 PD=1.04 PS=4.22 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.5 SB=75001.3
+ A=0.111 P=1.78 MULT=1
MM1000 N_A_27_368#_M1000_d N_A_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75003.5 A=0.168 P=2.54 MULT=1
MM1007 N_A_27_368#_M1007_d N_A_M1007_g N_VPWR_M1000_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75003.1 A=0.168 P=2.54 MULT=1
MM1008 N_A_27_368#_M1007_d N_A_M1008_g N_VPWR_M1008_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75002.6 A=0.168 P=2.54 MULT=1
MM1010 N_A_27_368#_M1010_d N_A_M1010_g N_VPWR_M1008_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.6 SB=75002.2 A=0.168 P=2.54 MULT=1
MM1002 N_Y_M1002_d N_B_M1002_g N_A_27_368#_M1010_d VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75002
+ SB=75001.7 A=0.168 P=2.54 MULT=1
MM1005 N_Y_M1002_d N_B_M1005_g N_A_27_368#_M1005_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75002.5 SB=75001.3 A=0.168 P=2.54 MULT=1
MM1009 N_Y_M1009_d N_B_M1009_g N_A_27_368#_M1005_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.196 AS=0.196 PD=1.47 PS=1.47 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75003 SB=75000.8 A=0.168 P=2.54 MULT=1
MM1011 N_Y_M1009_d N_B_M1011_g N_A_27_368#_M1011_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.196 AS=0.3976 PD=1.47 PS=2.95 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75003.5 SB=75000.3 A=0.168 P=2.54 MULT=1
DX12_noxref VNB VPB NWDIODE A=8.742 P=13.12
*
.include "sky130_fd_sc_ls__nor2_4.pxi.spice"
*
.ends
*
*
