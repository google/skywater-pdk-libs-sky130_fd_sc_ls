* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
X0 Y D1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X1 VPWR D1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X2 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X3 a_472_74# B1 a_841_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X4 Y D1 a_27_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X5 a_27_74# C1 a_472_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X6 a_841_74# B1 a_472_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X7 a_472_74# B1 a_841_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X8 a_954_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X9 a_954_368# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X10 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X11 Y A2 a_954_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X12 a_472_74# C1 a_27_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X13 VGND A1 a_841_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X14 a_841_74# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X15 VGND A2 a_841_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X16 a_27_74# C1 a_472_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X17 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X18 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X19 a_472_74# C1 a_27_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X20 a_841_74# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X21 VGND A2 a_841_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X22 a_954_368# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X23 VPWR A1 a_954_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X24 a_841_74# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X25 VGND A1 a_841_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X26 a_841_74# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X27 a_27_74# D1 Y VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X28 Y D1 a_27_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X29 a_841_74# B1 a_472_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X30 VPWR A1 a_954_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X31 a_27_74# D1 Y VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X32 Y A2 a_954_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X33 a_954_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
.ends
