* File: sky130_fd_sc_ls__bufinv_16.spice
* Created: Fri Aug 28 13:08:04 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__bufinv_16.pex.spice"
.subckt sky130_fd_sc_ls__bufinv_16  VNB VPB A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1025 N_VGND_M1025_d N_A_M1025_g N_A_27_74#_M1025_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1258 AS=0.2109 PD=1.08 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75011.2 A=0.111 P=1.78 MULT=1
MM1041 N_VGND_M1025_d N_A_M1041_g N_A_27_74#_M1041_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1258 AS=0.1036 PD=1.08 PS=1.02 NRD=9.72 NRS=0 M=1 R=4.93333 SA=75000.7
+ SB=75010.7 A=0.111 P=1.78 MULT=1
MM1049 N_VGND_M1049_d N_A_M1049_g N_A_27_74#_M1041_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75010.3 A=0.111 P=1.78 MULT=1
MM1003 N_A_384_74#_M1003_d N_A_27_74#_M1003_g N_VGND_M1049_d VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.6 SB=75009.9 A=0.111 P=1.78 MULT=1
MM1007 N_A_384_74#_M1003_d N_A_27_74#_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002
+ SB=75009.4 A=0.111 P=1.78 MULT=1
MM1008 N_A_384_74#_M1008_d N_A_27_74#_M1008_g N_VGND_M1007_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75002.4 SB=75009 A=0.111 P=1.78 MULT=1
MM1016 N_A_384_74#_M1008_d N_A_27_74#_M1016_g N_VGND_M1016_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75002.9 SB=75008.6 A=0.111 P=1.78 MULT=1
MM1044 N_A_384_74#_M1044_d N_A_27_74#_M1044_g N_VGND_M1016_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75003.3 SB=75008.1 A=0.111 P=1.78 MULT=1
MM1045 N_A_384_74#_M1044_d N_A_27_74#_M1045_g N_VGND_M1045_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75003.8 SB=75007.6 A=0.111 P=1.78 MULT=1
MM1000 N_VGND_M1045_s N_A_384_74#_M1000_g N_Y_M1000_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75004.3
+ SB=75007.2 A=0.111 P=1.78 MULT=1
MM1002 N_VGND_M1002_d N_A_384_74#_M1002_g N_Y_M1000_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75004.7
+ SB=75006.7 A=0.111 P=1.78 MULT=1
MM1005 N_VGND_M1002_d N_A_384_74#_M1005_g N_Y_M1005_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75005.1
+ SB=75006.3 A=0.111 P=1.78 MULT=1
MM1009 N_VGND_M1009_d N_A_384_74#_M1009_g N_Y_M1005_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75005.6
+ SB=75005.9 A=0.111 P=1.78 MULT=1
MM1011 N_VGND_M1009_d N_A_384_74#_M1011_g N_Y_M1011_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75006.1
+ SB=75005.4 A=0.111 P=1.78 MULT=1
MM1012 N_VGND_M1012_d N_A_384_74#_M1012_g N_Y_M1011_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75006.5
+ SB=75004.9 A=0.111 P=1.78 MULT=1
MM1018 N_VGND_M1012_d N_A_384_74#_M1018_g N_Y_M1018_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75007
+ SB=75004.4 A=0.111 P=1.78 MULT=1
MM1019 N_VGND_M1019_d N_A_384_74#_M1019_g N_Y_M1018_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75007.4
+ SB=75004 A=0.111 P=1.78 MULT=1
MM1020 N_VGND_M1019_d N_A_384_74#_M1020_g N_Y_M1020_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75007.9
+ SB=75003.5 A=0.111 P=1.78 MULT=1
MM1026 N_VGND_M1026_d N_A_384_74#_M1026_g N_Y_M1020_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75008.4
+ SB=75003.1 A=0.111 P=1.78 MULT=1
MM1030 N_VGND_M1026_d N_A_384_74#_M1030_g N_Y_M1030_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75008.9
+ SB=75002.6 A=0.111 P=1.78 MULT=1
MM1031 N_VGND_M1031_d N_A_384_74#_M1031_g N_Y_M1030_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75009.3
+ SB=75002.1 A=0.111 P=1.78 MULT=1
MM1032 N_VGND_M1031_d N_A_384_74#_M1032_g N_Y_M1032_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75009.8
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1033 N_VGND_M1033_d N_A_384_74#_M1033_g N_Y_M1032_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75010.2
+ SB=75001.2 A=0.111 P=1.78 MULT=1
MM1038 N_VGND_M1033_d N_A_384_74#_M1038_g N_Y_M1038_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75010.7
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1040 N_VGND_M1040_d N_A_384_74#_M1040_g N_Y_M1038_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2627 AS=0.1036 PD=2.19 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75011.1
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1021 N_VPWR_M1021_d N_A_M1021_g N_A_27_74#_M1021_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75011.2 A=0.168 P=2.54 MULT=1
MM1022 N_VPWR_M1021_d N_A_M1022_g N_A_27_74#_M1022_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75010.7 A=0.168 P=2.54 MULT=1
MM1034 N_VPWR_M1034_d N_A_M1034_g N_A_27_74#_M1022_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75010.3 A=0.168 P=2.54 MULT=1
MM1004 N_VPWR_M1034_d N_A_27_74#_M1004_g N_A_384_74#_M1004_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.1792 PD=1.42 PS=1.44 NRD=1.7533 NRS=5.2599 M=1 R=7.46667
+ SA=75001.6 SB=75009.8 A=0.168 P=2.54 MULT=1
MM1014 N_VPWR_M1014_d N_A_27_74#_M1014_g N_A_384_74#_M1004_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.1792 PD=1.42 PS=1.44 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002 SB=75009.4 A=0.168 P=2.54 MULT=1
MM1027 N_VPWR_M1014_d N_A_27_74#_M1027_g N_A_384_74#_M1027_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.5 SB=75008.9 A=0.168 P=2.54 MULT=1
MM1035 N_VPWR_M1035_d N_A_27_74#_M1035_g N_A_384_74#_M1027_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.9 SB=75008.5 A=0.168 P=2.54 MULT=1
MM1046 N_VPWR_M1035_d N_A_27_74#_M1046_g N_A_384_74#_M1046_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75003.4 SB=75008 A=0.168 P=2.54 MULT=1
MM1048 N_VPWR_M1048_d N_A_27_74#_M1048_g N_A_384_74#_M1046_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75003.8 SB=75007.6 A=0.168 P=2.54 MULT=1
MM1001 N_Y_M1001_d N_A_384_74#_M1001_g N_VPWR_M1048_d VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75004.3 SB=75007.1 A=0.168 P=2.54 MULT=1
MM1006 N_Y_M1001_d N_A_384_74#_M1006_g N_VPWR_M1006_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75004.7 SB=75006.7 A=0.168 P=2.54 MULT=1
MM1010 N_Y_M1010_d N_A_384_74#_M1010_g N_VPWR_M1006_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75005.2 SB=75006.2 A=0.168 P=2.54 MULT=1
MM1013 N_Y_M1010_d N_A_384_74#_M1013_g N_VPWR_M1013_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75005.6 SB=75005.8 A=0.168 P=2.54 MULT=1
MM1015 N_Y_M1015_d N_A_384_74#_M1015_g N_VPWR_M1013_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75006.1 SB=75005.3 A=0.168 P=2.54 MULT=1
MM1017 N_Y_M1015_d N_A_384_74#_M1017_g N_VPWR_M1017_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75006.5 SB=75004.9 A=0.168 P=2.54 MULT=1
MM1023 N_Y_M1023_d N_A_384_74#_M1023_g N_VPWR_M1017_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75007
+ SB=75004.4 A=0.168 P=2.54 MULT=1
MM1024 N_Y_M1023_d N_A_384_74#_M1024_g N_VPWR_M1024_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75007.4 SB=75004 A=0.168 P=2.54 MULT=1
MM1028 N_Y_M1028_d N_A_384_74#_M1028_g N_VPWR_M1024_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75007.9 SB=75003.5 A=0.168 P=2.54 MULT=1
MM1029 N_Y_M1028_d N_A_384_74#_M1029_g N_VPWR_M1029_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75008.3 SB=75003.1 A=0.168 P=2.54 MULT=1
MM1036 N_Y_M1036_d N_A_384_74#_M1036_g N_VPWR_M1029_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75008.8 SB=75002.6 A=0.168 P=2.54 MULT=1
MM1037 N_Y_M1036_d N_A_384_74#_M1037_g N_VPWR_M1037_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75009.3 SB=75002.1 A=0.168 P=2.54 MULT=1
MM1039 N_Y_M1039_d N_A_384_74#_M1039_g N_VPWR_M1037_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75009.8 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1042 N_Y_M1039_d N_A_384_74#_M1042_g N_VPWR_M1042_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.1736 PD=1.42 PS=1.43 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75010.2 SB=75001.2 A=0.168 P=2.54 MULT=1
MM1043 N_Y_M1043_d N_A_384_74#_M1043_g N_VPWR_M1042_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.1904 AS=0.1736 PD=1.46 PS=1.43 NRD=8.7862 NRS=3.5066 M=1 R=7.46667
+ SA=75010.7 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1047 N_Y_M1043_d N_A_384_74#_M1047_g N_VPWR_M1047_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.1904 AS=0.3304 PD=1.46 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75011.2 SB=75000.2 A=0.168 P=2.54 MULT=1
DX50_noxref VNB VPB NWDIODE A=23.0268 P=28.48
*
.include "sky130_fd_sc_ls__bufinv_16.pxi.spice"
*
.ends
*
*
