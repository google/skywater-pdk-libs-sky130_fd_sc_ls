* File: sky130_fd_sc_ls__fa_4.pex.spice
* Created: Wed Sep  2 11:07:44 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__FA_4%B 1 3 6 10 12 14 17 19 21 22 24 27 29 32 35 36
+ 37 40 43 47 50 52 54 55
c226 55 0 1.6719e-19 $X=6.48 $Y=1.665
c227 52 0 1.25803e-19 $X=4.62 $Y=1.805
c228 47 0 6.12639e-20 $X=4.115 $Y=1.41
c229 40 0 1.17721e-19 $X=2.645 $Y=1.41
c230 29 0 1.19152e-19 $X=1.665 $Y=1.417
r231 65 66 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.175
+ $Y=1.41 $X2=6.175 $Y2=1.41
r232 55 66 8.49543 $w=4.38e-07 $l=3.05e-07 $layer=LI1_cond $X=6.48 $Y=1.575
+ $X2=6.175 $Y2=1.575
r233 54 66 4.87443 $w=4.38e-07 $l=1.75e-07 $layer=LI1_cond $X=6 $Y=1.575
+ $X2=6.175 $Y2=1.575
r234 52 54 72.095 $w=1.98e-07 $l=1.295e-06 $layer=LI1_cond $X=4.62 $Y=1.805
+ $X2=5.915 $Y2=1.805
r235 50 51 10.3347 $w=2.42e-07 $l=2.05e-07 $layer=LI1_cond $X=2.645 $Y=1.83
+ $X2=2.645 $Y2=2.035
r236 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.115
+ $Y=1.41 $X2=4.115 $Y2=1.41
r237 45 52 35.0057 $w=1.76e-07 $l=5.10965e-07 $layer=LI1_cond $X=4.115 $Y=1.817
+ $X2=4.62 $Y2=1.805
r238 45 47 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.115 $Y=1.745
+ $X2=4.115 $Y2=1.41
r239 44 50 2.80567 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.81 $Y=1.83
+ $X2=2.645 $Y2=1.83
r240 43 45 11.4375 $w=1.76e-07 $l=1.71377e-07 $layer=LI1_cond $X=3.95 $Y=1.83
+ $X2=4.115 $Y2=1.817
r241 43 44 74.3743 $w=1.68e-07 $l=1.14e-06 $layer=LI1_cond $X=3.95 $Y=1.83
+ $X2=2.81 $Y2=1.83
r242 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.645
+ $Y=1.41 $X2=2.645 $Y2=1.41
r243 38 50 4.03333 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.645 $Y=1.745
+ $X2=2.645 $Y2=1.83
r244 38 40 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.645 $Y=1.745
+ $X2=2.645 $Y2=1.41
r245 36 51 2.80567 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.48 $Y=2.035
+ $X2=2.645 $Y2=2.035
r246 36 37 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=2.48 $Y=2.035
+ $X2=1.835 $Y2=2.035
r247 35 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.75 $Y=1.95
+ $X2=1.835 $Y2=2.035
r248 34 35 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.75 $Y=1.575
+ $X2=1.75 $Y2=1.95
r249 32 61 10.1831 $w=3.55e-07 $l=7.5e-08 $layer=POLY_cond $X=1.51 $Y=1.452
+ $X2=1.585 $Y2=1.452
r250 32 59 48.2 $w=3.55e-07 $l=3.55e-07 $layer=POLY_cond $X=1.51 $Y=1.452
+ $X2=1.155 $Y2=1.452
r251 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.51
+ $Y=1.41 $X2=1.51 $Y2=1.41
r252 29 34 7.64049 $w=3.15e-07 $l=1.95944e-07 $layer=LI1_cond $X=1.665 $Y=1.417
+ $X2=1.75 $Y2=1.575
r253 29 31 5.67075 $w=3.13e-07 $l=1.55e-07 $layer=LI1_cond $X=1.665 $Y=1.417
+ $X2=1.51 $Y2=1.417
r254 25 65 38.5562 $w=2.99e-07 $l=1.92678e-07 $layer=POLY_cond $X=6.115 $Y=1.245
+ $X2=6.175 $Y2=1.41
r255 25 27 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=6.115 $Y=1.245
+ $X2=6.115 $Y2=0.74
r256 22 65 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=6.1 $Y=1.66
+ $X2=6.175 $Y2=1.41
r257 22 24 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.1 $Y=1.66
+ $X2=6.1 $Y2=2.235
r258 19 48 52.2586 $w=2.99e-07 $l=2.76134e-07 $layer=POLY_cond $X=4.06 $Y=1.66
+ $X2=4.115 $Y2=1.41
r259 19 21 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=4.06 $Y=1.66
+ $X2=4.06 $Y2=2.235
r260 15 48 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=4.025 $Y=1.245
+ $X2=4.115 $Y2=1.41
r261 15 17 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=4.025 $Y=1.245
+ $X2=4.025 $Y2=0.74
r262 12 41 52.2586 $w=2.99e-07 $l=2.7157e-07 $layer=POLY_cond $X=2.6 $Y=1.66
+ $X2=2.645 $Y2=1.41
r263 12 14 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.6 $Y=1.66
+ $X2=2.6 $Y2=2.235
r264 8 41 38.5562 $w=2.99e-07 $l=1.92678e-07 $layer=POLY_cond $X=2.585 $Y=1.245
+ $X2=2.645 $Y2=1.41
r265 8 10 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=2.585 $Y=1.245
+ $X2=2.585 $Y2=0.74
r266 4 61 22.9692 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.585 $Y=1.245
+ $X2=1.585 $Y2=1.452
r267 4 6 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=1.585 $Y=1.245
+ $X2=1.585 $Y2=0.74
r268 1 59 22.9692 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.155 $Y=1.66
+ $X2=1.155 $Y2=1.452
r269 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.155 $Y=1.66
+ $X2=1.155 $Y2=2.235
.ends

.subckt PM_SKY130_FD_SC_LS__FA_4%CIN 1 3 4 6 9 11 13 14 16 17 19 22 25 26 27 28
+ 33 34 36 46 55
c151 34 0 9.09194e-20 $X=5.52 $Y=1.295
c152 14 0 1.48729e-19 $X=5.63 $Y=1.66
c153 9 0 1.78103e-19 $X=3.595 $Y=0.74
r154 39 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.105
+ $Y=1.385 $X2=2.105 $Y2=1.385
r155 36 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=1.295
+ $X2=2.16 $Y2=1.295
r156 34 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.635
+ $Y=1.385 $X2=5.635 $Y2=1.385
r157 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=1.295
+ $X2=5.52 $Y2=1.295
r158 31 55 3.27739 $w=3.93e-07 $l=9.5e-08 $layer=LI1_cond $X=3.12 $Y=1.377
+ $X2=3.215 $Y2=1.377
r159 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=1.295
+ $X2=3.12 $Y2=1.295
r160 28 30 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.265 $Y=1.295
+ $X2=3.12 $Y2=1.295
r161 27 33 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.375 $Y=1.295
+ $X2=5.52 $Y2=1.295
r162 27 28 2.61138 $w=1.4e-07 $l=2.11e-06 $layer=MET1_cond $X=5.375 $Y=1.295
+ $X2=3.265 $Y2=1.295
r163 26 36 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.305 $Y=1.295
+ $X2=2.16 $Y2=1.295
r164 25 30 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.975 $Y=1.295
+ $X2=3.12 $Y2=1.295
r165 25 26 0.829206 $w=1.4e-07 $l=6.7e-07 $layer=MET1_cond $X=2.975 $Y=1.295
+ $X2=2.305 $Y2=1.295
r166 22 55 13.1708 $w=3.13e-07 $l=3.6e-07 $layer=LI1_cond $X=3.575 $Y=1.417
+ $X2=3.215 $Y2=1.417
r167 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.575
+ $Y=1.41 $X2=3.575 $Y2=1.41
r168 17 43 38.5991 $w=2.92e-07 $l=2.05122e-07 $layer=POLY_cond $X=5.725 $Y=1.22
+ $X2=5.635 $Y2=1.385
r169 17 19 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.725 $Y=1.22
+ $X2=5.725 $Y2=0.74
r170 14 43 56.7567 $w=2.92e-07 $l=2.77489e-07 $layer=POLY_cond $X=5.63 $Y=1.66
+ $X2=5.635 $Y2=1.385
r171 14 16 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.63 $Y=1.66
+ $X2=5.63 $Y2=2.235
r172 11 23 52.2586 $w=2.99e-07 $l=2.66927e-07 $layer=POLY_cond $X=3.61 $Y=1.66
+ $X2=3.575 $Y2=1.41
r173 11 13 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.61 $Y=1.66
+ $X2=3.61 $Y2=2.235
r174 7 23 38.5562 $w=2.99e-07 $l=1.74714e-07 $layer=POLY_cond $X=3.595 $Y=1.245
+ $X2=3.575 $Y2=1.41
r175 7 9 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=3.595 $Y=1.245
+ $X2=3.595 $Y2=0.74
r176 4 39 56.7567 $w=2.92e-07 $l=2.96648e-07 $layer=POLY_cond $X=2.15 $Y=1.66
+ $X2=2.105 $Y2=1.385
r177 4 6 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.15 $Y=1.66
+ $X2=2.15 $Y2=2.235
r178 1 39 38.5991 $w=2.92e-07 $l=2.05122e-07 $layer=POLY_cond $X=2.015 $Y=1.22
+ $X2=2.105 $Y2=1.385
r179 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.015 $Y=1.22
+ $X2=2.015 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__FA_4%A_418_74# 1 2 7 9 10 12 13 15 18 20 22 25 27 29
+ 32 34 36 39 42 44 46 47 48 49 53 57 60 61 62 64 65 66 68 69 74 79 81 82 84 85
+ 90 91 92 105
c293 92 0 2.88491e-20 $X=5.095 $Y=1.005
c294 42 0 1.41883e-19 $X=1.09 $Y=1.745
c295 10 0 1.25803e-19 $X=5.13 $Y=1.66
c296 7 0 2.53523e-19 $X=5.045 $Y=1.22
r297 105 106 7.712 $w=3.75e-07 $l=6e-08 $layer=POLY_cond $X=10.485 $Y=1.542
+ $X2=10.545 $Y2=1.542
r298 104 105 47.5573 $w=3.75e-07 $l=3.7e-07 $layer=POLY_cond $X=10.115 $Y=1.542
+ $X2=10.485 $Y2=1.542
r299 103 104 10.2827 $w=3.75e-07 $l=8e-08 $layer=POLY_cond $X=10.035 $Y=1.542
+ $X2=10.115 $Y2=1.542
r300 100 101 19.28 $w=3.75e-07 $l=1.5e-07 $layer=POLY_cond $X=9.535 $Y=1.542
+ $X2=9.685 $Y2=1.542
r301 99 100 35.9893 $w=3.75e-07 $l=2.8e-07 $layer=POLY_cond $X=9.255 $Y=1.542
+ $X2=9.535 $Y2=1.542
r302 94 95 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.095
+ $Y=1.385 $X2=5.095 $Y2=1.385
r303 92 94 14.1774 $w=3.27e-07 $l=3.8e-07 $layer=LI1_cond $X=5.095 $Y=1.005
+ $X2=5.095 $Y2=1.385
r304 90 91 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=3.385 $Y=0.965
+ $X2=3.555 $Y2=0.965
r305 85 88 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=2.375 $Y=2.375
+ $X2=2.375 $Y2=2.455
r306 81 82 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=1.665 $Y=0.965
+ $X2=1.835 $Y2=0.965
r307 77 79 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.09 $Y=1.83
+ $X2=1.41 $Y2=1.83
r308 75 103 25.064 $w=3.75e-07 $l=1.95e-07 $layer=POLY_cond $X=9.84 $Y=1.542
+ $X2=10.035 $Y2=1.542
r309 75 101 19.9227 $w=3.75e-07 $l=1.55e-07 $layer=POLY_cond $X=9.84 $Y=1.542
+ $X2=9.685 $Y2=1.542
r310 74 75 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=9.84
+ $Y=1.485 $X2=9.84 $Y2=1.485
r311 72 99 12.2107 $w=3.75e-07 $l=9.5e-08 $layer=POLY_cond $X=9.16 $Y=1.542
+ $X2=9.255 $Y2=1.542
r312 72 97 9.64 $w=3.75e-07 $l=7.5e-08 $layer=POLY_cond $X=9.16 $Y=1.542
+ $X2=9.085 $Y2=1.542
r313 71 74 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=9.16 $Y=1.485
+ $X2=9.84 $Y2=1.485
r314 71 72 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=9.16
+ $Y=1.485 $X2=9.16 $Y2=1.485
r315 69 71 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=9.135 $Y=1.485
+ $X2=9.16 $Y2=1.485
r316 68 69 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.05 $Y=1.32
+ $X2=9.135 $Y2=1.485
r317 67 68 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=9.05 $Y=0.75
+ $X2=9.05 $Y2=1.32
r318 65 67 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.965 $Y=0.665
+ $X2=9.05 $Y2=0.75
r319 65 66 165.711 $w=1.68e-07 $l=2.54e-06 $layer=LI1_cond $X=8.965 $Y=0.665
+ $X2=6.425 $Y2=0.665
r320 64 66 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.34 $Y=0.58
+ $X2=6.425 $Y2=0.665
r321 63 64 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=6.34 $Y=0.425
+ $X2=6.34 $Y2=0.58
r322 61 63 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.255 $Y=0.34
+ $X2=6.34 $Y2=0.425
r323 61 62 65.2406 $w=1.68e-07 $l=1e-06 $layer=LI1_cond $X=6.255 $Y=0.34
+ $X2=5.255 $Y2=0.34
r324 60 92 5.97199 $w=3.27e-07 $l=1.16619e-07 $layer=LI1_cond $X=5.17 $Y=0.92
+ $X2=5.095 $Y2=1.005
r325 59 62 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.17 $Y=0.425
+ $X2=5.255 $Y2=0.34
r326 59 60 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=5.17 $Y=0.425
+ $X2=5.17 $Y2=0.92
r327 57 92 4.5696 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.93 $Y=1.005
+ $X2=5.095 $Y2=1.005
r328 57 91 89.7059 $w=1.68e-07 $l=1.375e-06 $layer=LI1_cond $X=4.93 $Y=1.005
+ $X2=3.555 $Y2=1.005
r329 56 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.465 $Y=0.925
+ $X2=2.3 $Y2=0.925
r330 56 90 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.465 $Y=0.925
+ $X2=3.385 $Y2=0.925
r331 51 84 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.3 $Y=0.84 $X2=2.3
+ $Y2=0.925
r332 51 53 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=2.3 $Y=0.84
+ $X2=2.3 $Y2=0.515
r333 49 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.135 $Y=0.925
+ $X2=2.3 $Y2=0.925
r334 49 82 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=2.135 $Y=0.925
+ $X2=1.835 $Y2=0.925
r335 47 85 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.21 $Y=2.375
+ $X2=2.375 $Y2=2.375
r336 47 48 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=2.21 $Y=2.375
+ $X2=1.495 $Y2=2.375
r337 46 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.41 $Y=2.29
+ $X2=1.495 $Y2=2.375
r338 45 79 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.41 $Y=1.915
+ $X2=1.41 $Y2=1.83
r339 45 46 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.41 $Y=1.915
+ $X2=1.41 $Y2=2.29
r340 44 81 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=1.175 $Y=1.005
+ $X2=1.665 $Y2=1.005
r341 42 77 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.09 $Y=1.745
+ $X2=1.09 $Y2=1.83
r342 41 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.09 $Y=1.09
+ $X2=1.175 $Y2=1.005
r343 41 42 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=1.09 $Y=1.09
+ $X2=1.09 $Y2=1.745
r344 37 106 24.2915 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=10.545 $Y=1.32
+ $X2=10.545 $Y2=1.542
r345 37 39 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=10.545 $Y=1.32
+ $X2=10.545 $Y2=0.78
r346 34 105 24.2915 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=10.485 $Y=1.765
+ $X2=10.485 $Y2=1.542
r347 34 36 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=10.485 $Y=1.765
+ $X2=10.485 $Y2=2.4
r348 30 104 24.2915 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=10.115 $Y=1.32
+ $X2=10.115 $Y2=1.542
r349 30 32 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=10.115 $Y=1.32
+ $X2=10.115 $Y2=0.78
r350 27 103 24.2915 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=10.035 $Y=1.765
+ $X2=10.035 $Y2=1.542
r351 27 29 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=10.035 $Y=1.765
+ $X2=10.035 $Y2=2.4
r352 23 101 24.2915 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=9.685 $Y=1.32
+ $X2=9.685 $Y2=1.542
r353 23 25 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=9.685 $Y=1.32
+ $X2=9.685 $Y2=0.78
r354 20 100 24.2915 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=9.535 $Y=1.765
+ $X2=9.535 $Y2=1.542
r355 20 22 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=9.535 $Y=1.765
+ $X2=9.535 $Y2=2.4
r356 16 99 24.2915 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=9.255 $Y=1.32
+ $X2=9.255 $Y2=1.542
r357 16 18 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=9.255 $Y=1.32
+ $X2=9.255 $Y2=0.78
r358 13 97 24.2915 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=9.085 $Y=1.765
+ $X2=9.085 $Y2=1.542
r359 13 15 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=9.085 $Y=1.765
+ $X2=9.085 $Y2=2.4
r360 10 95 56.7567 $w=2.92e-07 $l=2.91976e-07 $layer=POLY_cond $X=5.13 $Y=1.66
+ $X2=5.095 $Y2=1.385
r361 10 12 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.13 $Y=1.66
+ $X2=5.13 $Y2=2.235
r362 7 95 38.5991 $w=2.92e-07 $l=1.88348e-07 $layer=POLY_cond $X=5.045 $Y=1.22
+ $X2=5.095 $Y2=1.385
r363 7 9 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.045 $Y=1.22
+ $X2=5.045 $Y2=0.74
r364 2 88 600 $w=1.7e-07 $l=7.91454e-07 $layer=licon1_PDIFF $count=1 $X=2.225
+ $Y=1.735 $X2=2.375 $Y2=2.455
r365 1 84 182 $w=1.7e-07 $l=6.51594e-07 $layer=licon1_NDIFF $count=1 $X=2.09
+ $Y=0.37 $X2=2.3 $Y2=0.925
r366 1 53 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=2.09
+ $Y=0.37 $X2=2.3 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__FA_4%A 2 5 7 10 11 12 13 14 15 16 17 20 23 24 28 29
+ 30 31 32 33 36 37 41 43 46 47 48 49 50 52 54 55 62
c201 46 0 6.3363e-20 $X=6.64 $Y=2.34
c202 41 0 1.30844e-19 $X=6.625 $Y=0.74
c203 20 0 1.37405e-19 $X=3.11 $Y=2.235
r204 62 63 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.63
+ $Y=1.41 $X2=0.63 $Y2=1.41
r205 60 62 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=0.505 $Y=1.41
+ $X2=0.63 $Y2=1.41
r206 58 60 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.505 $Y2=1.41
r207 55 63 2.01209 $w=5.33e-07 $l=9e-08 $layer=LI1_cond $X=0.72 $Y=1.512
+ $X2=0.63 $Y2=1.512
r208 54 63 8.71908 $w=5.33e-07 $l=3.9e-07 $layer=LI1_cond $X=0.24 $Y=1.512
+ $X2=0.63 $Y2=1.512
r209 44 52 93.4966 $w=1.8e-07 $l=2.35e-07 $layer=POLY_cond $X=6.64 $Y=2.915
+ $X2=6.64 $Y2=3.15
r210 44 46 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.64 $Y=2.915
+ $X2=6.64 $Y2=2.34
r211 43 51 58.3064 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=6.64 $Y=1.765
+ $X2=6.64 $Y2=1.615
r212 43 46 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.64 $Y=1.765
+ $X2=6.64 $Y2=2.34
r213 41 51 448.67 $w=1.5e-07 $l=8.75e-07 $layer=POLY_cond $X=6.625 $Y=0.74
+ $X2=6.625 $Y2=1.615
r214 38 50 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.72 $Y=3.15 $X2=4.63
+ $Y2=3.15
r215 37 52 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=6.55 $Y=3.15 $X2=6.64
+ $Y2=3.15
r216 37 38 938.362 $w=1.5e-07 $l=1.83e-06 $layer=POLY_cond $X=6.55 $Y=3.15
+ $X2=4.72 $Y2=3.15
r217 34 36 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=4.63 $Y=2.81
+ $X2=4.63 $Y2=2.235
r218 33 36 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=4.63 $Y=1.66
+ $X2=4.63 $Y2=2.235
r219 32 50 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=4.63 $Y=3.075
+ $X2=4.63 $Y2=3.15
r220 31 34 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=4.63 $Y=2.9 $X2=4.63
+ $Y2=2.81
r221 31 32 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=4.63 $Y=2.9
+ $X2=4.63 $Y2=3.075
r222 30 33 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=4.63 $Y=1.57 $X2=4.63
+ $Y2=1.66
r223 29 49 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=4.63 $Y=1.275
+ $X2=4.63 $Y2=1.185
r224 29 30 114.669 $w=1.8e-07 $l=2.95e-07 $layer=POLY_cond $X=4.63 $Y=1.275
+ $X2=4.63 $Y2=1.57
r225 28 49 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=4.615 $Y=0.74
+ $X2=4.615 $Y2=1.185
r226 25 48 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.2 $Y=3.15 $X2=3.11
+ $Y2=3.15
r227 24 50 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.54 $Y=3.15 $X2=4.63
+ $Y2=3.15
r228 24 25 687.106 $w=1.5e-07 $l=1.34e-06 $layer=POLY_cond $X=4.54 $Y=3.15
+ $X2=3.2 $Y2=3.15
r229 23 47 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=3.125 $Y=0.74
+ $X2=3.125 $Y2=1.185
r230 18 20 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.11 $Y=2.81
+ $X2=3.11 $Y2=2.235
r231 17 20 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.11 $Y=1.66
+ $X2=3.11 $Y2=2.235
r232 16 48 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=3.11 $Y=3.075
+ $X2=3.11 $Y2=3.15
r233 15 18 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.11 $Y=2.9 $X2=3.11
+ $Y2=2.81
r234 15 16 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=3.11 $Y=2.9
+ $X2=3.11 $Y2=3.075
r235 14 17 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.11 $Y=1.57 $X2=3.11
+ $Y2=1.66
r236 13 47 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.11 $Y=1.275
+ $X2=3.11 $Y2=1.185
r237 13 14 114.669 $w=1.8e-07 $l=2.95e-07 $layer=POLY_cond $X=3.11 $Y=1.275
+ $X2=3.11 $Y2=1.57
r238 11 48 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.02 $Y=3.15 $X2=3.11
+ $Y2=3.15
r239 11 12 1243.46 $w=1.5e-07 $l=2.425e-06 $layer=POLY_cond $X=3.02 $Y=3.15
+ $X2=0.595 $Y2=3.15
r240 8 12 26.9307 $w=1.5e-07 $l=1.53542e-07 $layer=POLY_cond $X=0.505 $Y=3.035
+ $X2=0.595 $Y2=3.15
r241 8 10 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.505 $Y=3.035
+ $X2=0.505 $Y2=2.46
r242 7 10 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.505 $Y=1.885
+ $X2=0.505 $Y2=2.46
r243 3 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.245
+ $X2=0.495 $Y2=1.41
r244 3 5 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=0.495 $Y=1.245
+ $X2=0.495 $Y2=0.74
r245 2 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.505 $Y=1.795
+ $X2=0.505 $Y2=1.885
r246 1 60 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.575
+ $X2=0.505 $Y2=1.41
r247 1 2 85.5161 $w=1.8e-07 $l=2.2e-07 $layer=POLY_cond $X=0.505 $Y=1.575
+ $X2=0.505 $Y2=1.795
.ends

.subckt PM_SKY130_FD_SC_LS__FA_4%A_1024_74# 1 2 7 9 12 14 16 19 21 23 26 28 30
+ 33 37 41 43 46 48 54 58 60 64 65 66 70 79
c159 79 0 1.38341e-19 $X=8.585 $Y=1.552
c160 70 0 7.54566e-20 $X=6.99 $Y=1.505
r161 79 80 10.5934 $w=3.64e-07 $l=8e-08 $layer=POLY_cond $X=8.585 $Y=1.552
+ $X2=8.665 $Y2=1.552
r162 78 79 46.3462 $w=3.64e-07 $l=3.5e-07 $layer=POLY_cond $X=8.235 $Y=1.552
+ $X2=8.585 $Y2=1.552
r163 77 78 13.2418 $w=3.64e-07 $l=1e-07 $layer=POLY_cond $X=8.135 $Y=1.552
+ $X2=8.235 $Y2=1.552
r164 74 75 1.32418 $w=3.64e-07 $l=1e-08 $layer=POLY_cond $X=7.635 $Y=1.552
+ $X2=7.645 $Y2=1.552
r165 71 72 3.97253 $w=3.64e-07 $l=3e-08 $layer=POLY_cond $X=7.185 $Y=1.552
+ $X2=7.215 $Y2=1.552
r166 66 68 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=6.34 $Y=2.035
+ $X2=6.34 $Y2=2.145
r167 64 65 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=5.915 $Y=0.965
+ $X2=6.085 $Y2=0.965
r168 60 62 5.76222 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=5.55 $Y=0.8
+ $X2=5.55 $Y2=0.925
r169 55 77 25.8214 $w=3.64e-07 $l=1.95e-07 $layer=POLY_cond $X=7.94 $Y=1.552
+ $X2=8.135 $Y2=1.552
r170 55 75 39.0632 $w=3.64e-07 $l=2.95e-07 $layer=POLY_cond $X=7.94 $Y=1.552
+ $X2=7.645 $Y2=1.552
r171 54 55 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=7.94
+ $Y=1.505 $X2=7.94 $Y2=1.505
r172 52 74 49.6566 $w=3.64e-07 $l=3.75e-07 $layer=POLY_cond $X=7.26 $Y=1.552
+ $X2=7.635 $Y2=1.552
r173 52 72 5.95879 $w=3.64e-07 $l=4.5e-08 $layer=POLY_cond $X=7.26 $Y=1.552
+ $X2=7.215 $Y2=1.552
r174 51 54 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=7.26 $Y=1.505
+ $X2=7.94 $Y2=1.505
r175 51 52 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=7.26
+ $Y=1.505 $X2=7.26 $Y2=1.505
r176 49 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.075 $Y=1.505
+ $X2=6.99 $Y2=1.505
r177 49 51 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=7.075 $Y=1.505
+ $X2=7.26 $Y2=1.505
r178 47 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.99 $Y=1.67
+ $X2=6.99 $Y2=1.505
r179 47 48 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=6.99 $Y=1.67
+ $X2=6.99 $Y2=1.95
r180 46 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.99 $Y=1.34
+ $X2=6.99 $Y2=1.505
r181 45 46 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=6.99 $Y=1.09
+ $X2=6.99 $Y2=1.34
r182 44 66 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.425 $Y=2.035
+ $X2=6.34 $Y2=2.035
r183 43 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.905 $Y=2.035
+ $X2=6.99 $Y2=1.95
r184 43 44 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=6.905 $Y=2.035
+ $X2=6.425 $Y2=2.035
r185 41 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.905 $Y=1.005
+ $X2=6.99 $Y2=1.09
r186 41 65 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=6.905 $Y=1.005
+ $X2=6.085 $Y2=1.005
r187 40 62 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.675 $Y=0.925
+ $X2=5.55 $Y2=0.925
r188 40 64 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=5.675 $Y=0.925
+ $X2=5.915 $Y2=0.925
r189 38 58 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.57 $Y=2.145
+ $X2=5.405 $Y2=2.145
r190 37 68 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.255 $Y=2.145
+ $X2=6.34 $Y2=2.145
r191 37 38 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=6.255 $Y=2.145
+ $X2=5.57 $Y2=2.145
r192 31 80 23.572 $w=1.5e-07 $l=2.12e-07 $layer=POLY_cond $X=8.665 $Y=1.34
+ $X2=8.665 $Y2=1.552
r193 31 33 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=8.665 $Y=1.34
+ $X2=8.665 $Y2=0.78
r194 28 79 23.572 $w=1.5e-07 $l=2.13e-07 $layer=POLY_cond $X=8.585 $Y=1.765
+ $X2=8.585 $Y2=1.552
r195 28 30 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.585 $Y=1.765
+ $X2=8.585 $Y2=2.4
r196 24 78 23.572 $w=1.5e-07 $l=2.12e-07 $layer=POLY_cond $X=8.235 $Y=1.34
+ $X2=8.235 $Y2=1.552
r197 24 26 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=8.235 $Y=1.34
+ $X2=8.235 $Y2=0.78
r198 21 77 23.572 $w=1.5e-07 $l=2.13e-07 $layer=POLY_cond $X=8.135 $Y=1.765
+ $X2=8.135 $Y2=1.552
r199 21 23 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.135 $Y=1.765
+ $X2=8.135 $Y2=2.4
r200 17 75 23.572 $w=1.5e-07 $l=2.12e-07 $layer=POLY_cond $X=7.645 $Y=1.34
+ $X2=7.645 $Y2=1.552
r201 17 19 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=7.645 $Y=1.34
+ $X2=7.645 $Y2=0.78
r202 14 74 23.572 $w=1.5e-07 $l=2.13e-07 $layer=POLY_cond $X=7.635 $Y=1.765
+ $X2=7.635 $Y2=1.552
r203 14 16 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.635 $Y=1.765
+ $X2=7.635 $Y2=2.4
r204 10 72 23.572 $w=1.5e-07 $l=2.12e-07 $layer=POLY_cond $X=7.215 $Y=1.34
+ $X2=7.215 $Y2=1.552
r205 10 12 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=7.215 $Y=1.34
+ $X2=7.215 $Y2=0.78
r206 7 71 23.572 $w=1.5e-07 $l=2.13e-07 $layer=POLY_cond $X=7.185 $Y=1.765
+ $X2=7.185 $Y2=1.552
r207 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.185 $Y=1.765
+ $X2=7.185 $Y2=2.4
r208 2 58 300 $w=1.7e-07 $l=5.001e-07 $layer=licon1_PDIFF $count=2 $X=5.205
+ $Y=1.735 $X2=5.405 $Y2=2.145
r209 1 60 182 $w=1.7e-07 $l=5.93801e-07 $layer=licon1_NDIFF $count=1 $X=5.12
+ $Y=0.37 $X2=5.51 $Y2=0.8
.ends

.subckt PM_SKY130_FD_SC_LS__FA_4%A_27_392# 1 2 7 9 11 14 15 19
r51 17 19 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=1.465 $Y=2.795
+ $X2=1.84 $Y2=2.795
r52 15 17 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=1.155 $Y=2.795
+ $X2=1.465 $Y2=2.795
r53 14 15 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.07 $Y=2.63
+ $X2=1.155 $Y2=2.795
r54 13 14 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.07 $Y=2.255
+ $X2=1.07 $Y2=2.63
r55 12 22 4.68787 $w=1.7e-07 $l=1.96074e-07 $layer=LI1_cond $X=0.445 $Y=2.17
+ $X2=0.28 $Y2=2.102
r56 11 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.985 $Y=2.17
+ $X2=1.07 $Y2=2.255
r57 11 12 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=0.985 $Y=2.17
+ $X2=0.445 $Y2=2.17
r58 7 22 3.0783 $w=3.3e-07 $l=1.53e-07 $layer=LI1_cond $X=0.28 $Y=2.255 $X2=0.28
+ $Y2=2.102
r59 7 9 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=0.28 $Y=2.255 $X2=0.28
+ $Y2=2.815
r60 2 19 600 $w=1.7e-07 $l=1.33049e-06 $layer=licon1_PDIFF $count=1 $X=1.23
+ $Y=1.735 $X2=1.84 $Y2=2.795
r61 2 17 600 $w=1.7e-07 $l=1.17162e-06 $layer=licon1_PDIFF $count=1 $X=1.23
+ $Y=1.735 $X2=1.465 $Y2=2.795
r62 1 22 400 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.28 $Y2=2.115
r63 1 9 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.28 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_LS__FA_4%VPWR 1 2 3 4 5 6 7 8 29 33 37 41 47 51 57 59 61
+ 66 67 68 77 81 86 91 96 101 107 110 113 116 119 122 126
c150 3 0 6.12639e-20 $X=4.135 $Y=1.735
c151 1 0 1.41883e-19 $X=0.58 $Y=1.96
r152 125 126 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r153 122 123 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r154 119 120 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r155 116 117 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r156 113 114 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r157 110 111 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r158 107 108 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r159 105 126 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=10.8 $Y2=3.33
r160 105 123 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=9.84 $Y2=3.33
r161 104 105 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r162 102 122 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.925 $Y=3.33
+ $X2=9.8 $Y2=3.33
r163 102 104 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=9.925 $Y=3.33
+ $X2=10.32 $Y2=3.33
r164 101 125 3.95357 $w=1.7e-07 $l=2.07e-07 $layer=LI1_cond $X=10.625 $Y=3.33
+ $X2=10.832 $Y2=3.33
r165 101 104 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=10.625 $Y=3.33
+ $X2=10.32 $Y2=3.33
r166 100 123 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=9.84 $Y2=3.33
r167 100 120 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=8.88 $Y2=3.33
r168 99 100 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r169 97 119 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.975 $Y=3.33
+ $X2=8.85 $Y2=3.33
r170 97 99 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=8.975 $Y=3.33
+ $X2=9.36 $Y2=3.33
r171 96 122 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.675 $Y=3.33
+ $X2=9.8 $Y2=3.33
r172 96 99 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=9.675 $Y=3.33
+ $X2=9.36 $Y2=3.33
r173 95 120 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=8.88 $Y2=3.33
r174 95 117 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=7.92 $Y2=3.33
r175 94 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33 $X2=8.4
+ $Y2=3.33
r176 92 116 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.025 $Y=3.33
+ $X2=7.9 $Y2=3.33
r177 92 94 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=8.025 $Y=3.33
+ $X2=8.4 $Y2=3.33
r178 91 119 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.725 $Y=3.33
+ $X2=8.85 $Y2=3.33
r179 91 94 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=8.725 $Y=3.33
+ $X2=8.4 $Y2=3.33
r180 90 117 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r181 90 114 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6.96 $Y2=3.33
r182 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r183 87 113 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.045 $Y=3.33
+ $X2=6.92 $Y2=3.33
r184 87 89 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=7.045 $Y=3.33
+ $X2=7.44 $Y2=3.33
r185 86 116 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.775 $Y=3.33
+ $X2=7.9 $Y2=3.33
r186 86 89 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=7.775 $Y=3.33
+ $X2=7.44 $Y2=3.33
r187 85 114 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6.96 $Y2=3.33
r188 84 85 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r189 82 110 9.81116 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=4.57 $Y=3.33 $X2=4.37
+ $Y2=3.33
r190 82 84 124.61 $w=1.68e-07 $l=1.91e-06 $layer=LI1_cond $X=4.57 $Y=3.33
+ $X2=6.48 $Y2=3.33
r191 81 113 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.795 $Y=3.33
+ $X2=6.92 $Y2=3.33
r192 81 84 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=6.795 $Y=3.33
+ $X2=6.48 $Y2=3.33
r193 80 111 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r194 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r195 77 110 9.81116 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=4.17 $Y=3.33 $X2=4.37
+ $Y2=3.33
r196 77 79 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=4.17 $Y=3.33 $X2=4.08
+ $Y2=3.33
r197 76 80 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r198 75 76 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r199 73 76 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=3.12 $Y2=3.33
r200 73 108 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r201 72 75 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=3.12 $Y2=3.33
r202 72 73 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r203 70 107 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=3.33
+ $X2=0.73 $Y2=3.33
r204 70 72 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.815 $Y=3.33
+ $X2=1.2 $Y2=3.33
r205 68 85 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6.48 $Y2=3.33
r206 68 111 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=4.56 $Y2=3.33
r207 66 75 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=3.17 $Y=3.33 $X2=3.12
+ $Y2=3.33
r208 66 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.17 $Y=3.33
+ $X2=3.335 $Y2=3.33
r209 65 79 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=3.5 $Y=3.33
+ $X2=4.08 $Y2=3.33
r210 65 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.5 $Y=3.33
+ $X2=3.335 $Y2=3.33
r211 61 64 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=10.75 $Y=1.985
+ $X2=10.75 $Y2=2.815
r212 59 125 3.18959 $w=2.5e-07 $l=1.19143e-07 $layer=LI1_cond $X=10.75 $Y=3.245
+ $X2=10.832 $Y2=3.33
r213 59 64 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=10.75 $Y=3.245
+ $X2=10.75 $Y2=2.815
r214 55 122 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.8 $Y=3.245
+ $X2=9.8 $Y2=3.33
r215 55 57 42.4099 $w=2.48e-07 $l=9.2e-07 $layer=LI1_cond $X=9.8 $Y=3.245
+ $X2=9.8 $Y2=2.325
r216 51 54 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=8.85 $Y=1.985
+ $X2=8.85 $Y2=2.815
r217 49 119 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.85 $Y=3.245
+ $X2=8.85 $Y2=3.33
r218 49 54 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=8.85 $Y=3.245
+ $X2=8.85 $Y2=2.815
r219 45 116 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.9 $Y=3.245
+ $X2=7.9 $Y2=3.33
r220 45 47 41.4879 $w=2.48e-07 $l=9e-07 $layer=LI1_cond $X=7.9 $Y=3.245 $X2=7.9
+ $Y2=2.345
r221 41 44 16.5952 $w=2.48e-07 $l=3.6e-07 $layer=LI1_cond $X=6.92 $Y=2.455
+ $X2=6.92 $Y2=2.815
r222 39 113 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.92 $Y=3.245
+ $X2=6.92 $Y2=3.33
r223 39 44 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=6.92 $Y=3.245
+ $X2=6.92 $Y2=2.815
r224 35 110 1.46811 $w=4e-07 $l=8.5e-08 $layer=LI1_cond $X=4.37 $Y=3.245
+ $X2=4.37 $Y2=3.33
r225 35 37 18.8713 $w=3.98e-07 $l=6.55e-07 $layer=LI1_cond $X=4.37 $Y=3.245
+ $X2=4.37 $Y2=2.59
r226 31 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.335 $Y=3.245
+ $X2=3.335 $Y2=3.33
r227 31 33 37.5417 $w=3.28e-07 $l=1.075e-06 $layer=LI1_cond $X=3.335 $Y=3.245
+ $X2=3.335 $Y2=2.17
r228 27 107 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=3.33
r229 27 29 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=2.59
r230 8 64 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=10.56
+ $Y=1.84 $X2=10.71 $Y2=2.815
r231 8 61 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=10.56
+ $Y=1.84 $X2=10.71 $Y2=1.985
r232 7 57 300 $w=1.7e-07 $l=5.54955e-07 $layer=licon1_PDIFF $count=2 $X=9.61
+ $Y=1.84 $X2=9.76 $Y2=2.325
r233 6 54 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=8.66
+ $Y=1.84 $X2=8.81 $Y2=2.815
r234 6 51 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=8.66
+ $Y=1.84 $X2=8.81 $Y2=1.985
r235 5 47 300 $w=1.7e-07 $l=5.7513e-07 $layer=licon1_PDIFF $count=2 $X=7.71
+ $Y=1.84 $X2=7.86 $Y2=2.345
r236 4 44 600 $w=1.7e-07 $l=1.09064e-06 $layer=licon1_PDIFF $count=1 $X=6.715
+ $Y=1.84 $X2=6.96 $Y2=2.815
r237 4 41 600 $w=1.7e-07 $l=7.27255e-07 $layer=licon1_PDIFF $count=1 $X=6.715
+ $Y=1.84 $X2=6.96 $Y2=2.455
r238 3 37 600 $w=1.7e-07 $l=9.65376e-07 $layer=licon1_PDIFF $count=1 $X=4.135
+ $Y=1.735 $X2=4.37 $Y2=2.59
r239 2 33 300 $w=1.7e-07 $l=5.04455e-07 $layer=licon1_PDIFF $count=2 $X=3.185
+ $Y=1.735 $X2=3.335 $Y2=2.17
r240 1 29 600 $w=1.7e-07 $l=7.00999e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.96 $X2=0.73 $Y2=2.59
.ends

.subckt PM_SKY130_FD_SC_LS__FA_4%A_737_347# 1 2 9 11 13 16
c29 16 0 1.37405e-19 $X=3.835 $Y=2.17
c30 13 0 1.48729e-19 $X=4.905 $Y=2.59
r31 11 18 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.905 $Y=2.255
+ $X2=4.905 $Y2=2.17
r32 11 13 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.905 $Y=2.255
+ $X2=4.905 $Y2=2.59
r33 10 16 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4 $Y=2.17 $X2=3.835
+ $Y2=2.17
r34 9 18 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.74 $Y=2.17
+ $X2=4.905 $Y2=2.17
r35 9 10 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=4.74 $Y=2.17 $X2=4
+ $Y2=2.17
r36 2 18 600 $w=1.7e-07 $l=5.25571e-07 $layer=licon1_PDIFF $count=1 $X=4.705
+ $Y=1.735 $X2=4.905 $Y2=2.17
r37 2 13 600 $w=1.7e-07 $l=9.4975e-07 $layer=licon1_PDIFF $count=1 $X=4.705
+ $Y=1.735 $X2=4.905 $Y2=2.59
r38 1 16 300 $w=1.7e-07 $l=5.04455e-07 $layer=licon1_PDIFF $count=2 $X=3.685
+ $Y=1.735 $X2=3.835 $Y2=2.17
.ends

.subckt PM_SKY130_FD_SC_LS__FA_4%SUM 1 2 3 4 13 15 17 21 23 24 29 30 31 38
c63 29 0 1.61113e-19 $X=8.315 $Y=1.95
c64 17 0 1.30844e-19 $X=8.285 $Y=1.045
c65 13 0 6.3363e-20 $X=7.41 $Y=2.01
r66 36 38 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=8.36 $Y=2.01
+ $X2=8.36 $Y2=2.035
r67 30 31 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=8.36 $Y=2.405
+ $X2=8.36 $Y2=2.775
r68 29 36 3.29812 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=8.36 $Y=1.925
+ $X2=8.36 $Y2=2.01
r69 29 30 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=8.36 $Y=2.065
+ $X2=8.36 $Y2=2.405
r70 29 38 1.04768 $w=3.28e-07 $l=3e-08 $layer=LI1_cond $X=8.36 $Y=2.065 $X2=8.36
+ $Y2=2.035
r71 24 29 3.29812 $w=2.85e-07 $l=1.05119e-07 $layer=LI1_cond $X=8.405 $Y=1.84
+ $X2=8.36 $Y2=1.925
r72 23 28 3.46099 $w=2.4e-07 $l=1.45774e-07 $layer=LI1_cond $X=8.405 $Y=1.17
+ $X2=8.45 $Y2=1.045
r73 23 24 32.1724 $w=2.38e-07 $l=6.7e-07 $layer=LI1_cond $X=8.405 $Y=1.17
+ $X2=8.405 $Y2=1.84
r74 22 26 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.575 $Y=1.925
+ $X2=7.41 $Y2=1.925
r75 21 29 3.25423 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.195 $Y=1.925
+ $X2=8.36 $Y2=1.925
r76 21 22 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=8.195 $Y=1.925
+ $X2=7.575 $Y2=1.925
r77 17 28 3.3592 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=8.285 $Y=1.045
+ $X2=8.45 $Y2=1.045
r78 17 19 39.4136 $w=2.48e-07 $l=8.55e-07 $layer=LI1_cond $X=8.285 $Y=1.045
+ $X2=7.43 $Y2=1.045
r79 13 26 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.41 $Y=2.01 $X2=7.41
+ $Y2=1.925
r80 13 15 28.1126 $w=3.28e-07 $l=8.05e-07 $layer=LI1_cond $X=7.41 $Y=2.01
+ $X2=7.41 $Y2=2.815
r81 4 29 400 $w=1.7e-07 $l=2.2798e-07 $layer=licon1_PDIFF $count=1 $X=8.21
+ $Y=1.84 $X2=8.36 $Y2=2.005
r82 4 31 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=8.21
+ $Y=1.84 $X2=8.36 $Y2=2.815
r83 3 26 400 $w=1.7e-07 $l=2.2798e-07 $layer=licon1_PDIFF $count=1 $X=7.26
+ $Y=1.84 $X2=7.41 $Y2=2.005
r84 3 15 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=7.26
+ $Y=1.84 $X2=7.41 $Y2=2.815
r85 2 28 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=8.31
+ $Y=0.41 $X2=8.45 $Y2=1.005
r86 1 19 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=7.29
+ $Y=0.41 $X2=7.43 $Y2=1.005
.ends

.subckt PM_SKY130_FD_SC_LS__FA_4%COUT 1 2 3 4 13 15 19 21 23 24 27 30 33 34 35
+ 36 37 43 45
c69 43 0 9.5881e-20 $X=10.265 $Y=1.99
r70 43 45 1.52529 $w=3.38e-07 $l=4.5e-08 $layer=LI1_cond $X=10.265 $Y=1.99
+ $X2=10.265 $Y2=2.035
r71 36 37 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=10.265 $Y=2.405
+ $X2=10.265 $Y2=2.775
r72 35 43 0.944793 $w=3.4e-07 $l=2e-08 $layer=LI1_cond $X=10.265 $Y=1.97
+ $X2=10.265 $Y2=1.99
r73 35 55 2.67003 $w=2.97e-07 $l=6.5e-08 $layer=LI1_cond $X=10.265 $Y=1.97
+ $X2=10.265 $Y2=1.905
r74 35 36 11.8634 $w=3.38e-07 $l=3.5e-07 $layer=LI1_cond $X=10.265 $Y=2.055
+ $X2=10.265 $Y2=2.405
r75 35 45 0.677908 $w=3.38e-07 $l=2e-08 $layer=LI1_cond $X=10.265 $Y=2.055
+ $X2=10.265 $Y2=2.035
r76 34 55 9.85859 $w=2.97e-07 $l=2.4e-07 $layer=LI1_cond $X=10.265 $Y=1.665
+ $X2=10.265 $Y2=1.905
r77 30 34 4.94494 $w=2.97e-07 $l=1.29132e-07 $layer=LI1_cond $X=10.295 $Y=1.55
+ $X2=10.265 $Y2=1.665
r78 29 33 3.58051 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=10.295 $Y=1.15
+ $X2=10.295 $Y2=1.065
r79 29 30 17.7299 $w=2.58e-07 $l=4e-07 $layer=LI1_cond $X=10.295 $Y=1.15
+ $X2=10.295 $Y2=1.55
r80 25 33 3.58051 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=10.295 $Y=0.98
+ $X2=10.295 $Y2=1.065
r81 25 27 18.838 $w=2.58e-07 $l=4.25e-07 $layer=LI1_cond $X=10.295 $Y=0.98
+ $X2=10.295 $Y2=0.555
r82 23 33 2.90867 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=10.165 $Y=1.065
+ $X2=10.295 $Y2=1.065
r83 23 24 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=10.165 $Y=1.065
+ $X2=9.555 $Y2=1.065
r84 22 32 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.475 $Y=1.905
+ $X2=9.31 $Y2=1.905
r85 21 55 4.00195 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=10.095 $Y=1.905
+ $X2=10.265 $Y2=1.905
r86 21 22 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=10.095 $Y=1.905
+ $X2=9.475 $Y2=1.905
r87 17 24 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=9.43 $Y=0.98
+ $X2=9.555 $Y2=1.065
r88 17 19 19.5915 $w=2.48e-07 $l=4.25e-07 $layer=LI1_cond $X=9.43 $Y=0.98
+ $X2=9.43 $Y2=0.555
r89 13 32 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.31 $Y=1.99 $X2=9.31
+ $Y2=1.905
r90 13 15 28.8111 $w=3.28e-07 $l=8.25e-07 $layer=LI1_cond $X=9.31 $Y=1.99
+ $X2=9.31 $Y2=2.815
r91 4 35 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=10.11
+ $Y=1.84 $X2=10.26 $Y2=1.985
r92 4 37 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=10.11
+ $Y=1.84 $X2=10.26 $Y2=2.815
r93 3 32 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=9.16
+ $Y=1.84 $X2=9.31 $Y2=1.985
r94 3 15 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=9.16
+ $Y=1.84 $X2=9.31 $Y2=2.815
r95 2 27 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.19
+ $Y=0.41 $X2=10.33 $Y2=0.555
r96 1 19 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.33
+ $Y=0.41 $X2=9.47 $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_LS__FA_4%A_27_74# 1 2 11 14 18 19
r32 18 19 8.64032 $w=3.18e-07 $l=1.7e-07 $layer=LI1_cond $X=1.325 $Y=0.55
+ $X2=1.495 $Y2=0.55
r33 14 16 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=0.28 $Y=0.515
+ $X2=0.28 $Y2=0.665
r34 11 19 10.9842 $w=3.18e-07 $l=3.05e-07 $layer=LI1_cond $X=1.8 $Y=0.51
+ $X2=1.495 $Y2=0.51
r35 8 16 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.445 $Y=0.665
+ $X2=0.28 $Y2=0.665
r36 8 18 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=0.445 $Y=0.665
+ $X2=1.325 $Y2=0.665
r37 2 11 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=1.66 $Y=0.37
+ $X2=1.8 $Y2=0.55
r38 1 14 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__FA_4%VGND 1 2 3 4 5 6 7 8 27 31 33 35 38 39 40 41 47
+ 64 71 76 81 86 94 97 100 107 114 120 124
r146 123 124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=0
+ $X2=10.8 $Y2=0
r147 120 121 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0
+ $X2=9.84 $Y2=0
r148 114 117 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=8.96 $Y=0
+ $X2=8.96 $Y2=0.325
r149 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r150 107 110 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=7.94 $Y=0
+ $X2=7.94 $Y2=0.325
r151 107 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r152 100 103 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=6.92 $Y=0
+ $X2=6.92 $Y2=0.325
r153 100 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r154 96 97 11.9029 $w=4.93e-07 $l=2.65e-07 $layer=LI1_cond $X=0.89 $Y=0.162
+ $X2=1.155 $Y2=0.162
r155 92 96 4.10774 $w=4.93e-07 $l=1.7e-07 $layer=LI1_cond $X=0.72 $Y=0.162
+ $X2=0.89 $Y2=0.162
r156 92 94 7.79514 $w=4.93e-07 $l=9.5e-08 $layer=LI1_cond $X=0.72 $Y=0.162
+ $X2=0.625 $Y2=0.162
r157 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r158 90 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=10.8 $Y2=0
r159 90 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=9.84 $Y2=0
r160 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r161 87 120 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.985 $Y=0
+ $X2=9.86 $Y2=0
r162 87 89 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=9.985 $Y=0
+ $X2=10.32 $Y2=0
r163 86 123 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=10.595 $Y=0
+ $X2=10.817 $Y2=0
r164 86 89 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=10.595 $Y=0
+ $X2=10.32 $Y2=0
r165 85 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=9.84 $Y2=0
r166 85 115 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=8.88 $Y2=0
r167 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r168 82 114 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.125 $Y=0
+ $X2=8.96 $Y2=0
r169 82 84 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=9.125 $Y=0
+ $X2=9.36 $Y2=0
r170 81 120 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.735 $Y=0
+ $X2=9.86 $Y2=0
r171 81 84 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=9.735 $Y=0
+ $X2=9.36 $Y2=0
r172 80 115 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=8.88
+ $Y2=0
r173 80 108 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=7.92
+ $Y2=0
r174 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r175 77 107 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.105 $Y=0
+ $X2=7.94 $Y2=0
r176 77 79 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=8.105 $Y=0 $X2=8.4
+ $Y2=0
r177 76 114 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.795 $Y=0
+ $X2=8.96 $Y2=0
r178 76 79 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=8.795 $Y=0 $X2=8.4
+ $Y2=0
r179 75 108 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=7.92 $Y2=0
r180 75 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=6.96 $Y2=0
r181 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r182 72 100 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.085 $Y=0
+ $X2=6.92 $Y2=0
r183 72 74 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=7.085 $Y=0
+ $X2=7.44 $Y2=0
r184 71 107 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.775 $Y=0
+ $X2=7.94 $Y2=0
r185 71 74 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=7.775 $Y=0
+ $X2=7.44 $Y2=0
r186 70 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0
+ $X2=6.96 $Y2=0
r187 69 70 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r188 66 69 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.56 $Y=0 $X2=6.48
+ $Y2=0
r189 66 67 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r190 64 100 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.755 $Y=0
+ $X2=6.92 $Y2=0
r191 64 69 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.755 $Y=0
+ $X2=6.48 $Y2=0
r192 63 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r193 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r194 60 63 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r195 59 60 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r196 57 60 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r197 57 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r198 56 59 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r199 56 97 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=1.2 $Y=0 $X2=1.155
+ $Y2=0
r200 56 57 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r201 52 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r202 51 94 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.24 $Y=0
+ $X2=0.625 $Y2=0
r203 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r204 47 70 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6.48
+ $Y2=0
r205 47 67 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=4.56
+ $Y2=0
r206 43 66 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=4.485 $Y=0 $X2=4.56
+ $Y2=0
r207 41 62 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=4.155 $Y=0 $X2=4.08
+ $Y2=0
r208 40 45 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=4.32 $Y=0 $X2=4.32
+ $Y2=0.325
r209 40 43 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.32 $Y=0 $X2=4.485
+ $Y2=0
r210 40 41 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.32 $Y=0 $X2=4.155
+ $Y2=0
r211 38 59 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=3.175 $Y=0 $X2=3.12
+ $Y2=0
r212 38 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.175 $Y=0 $X2=3.34
+ $Y2=0
r213 37 62 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=3.505 $Y=0
+ $X2=4.08 $Y2=0
r214 37 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.505 $Y=0 $X2=3.34
+ $Y2=0
r215 33 123 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=10.76 $Y=0.085
+ $X2=10.817 $Y2=0
r216 33 35 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=10.76 $Y=0.085
+ $X2=10.76 $Y2=0.555
r217 29 120 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.86 $Y=0.085
+ $X2=9.86 $Y2=0
r218 29 31 25.8147 $w=2.48e-07 $l=5.6e-07 $layer=LI1_cond $X=9.86 $Y=0.085
+ $X2=9.86 $Y2=0.645
r219 25 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.34 $Y=0.085
+ $X2=3.34 $Y2=0
r220 25 27 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=3.34 $Y=0.085
+ $X2=3.34 $Y2=0.55
r221 8 35 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.62
+ $Y=0.41 $X2=10.76 $Y2=0.555
r222 7 31 182 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=1 $X=9.76
+ $Y=0.41 $X2=9.9 $Y2=0.645
r223 6 117 182 $w=1.7e-07 $l=2.59037e-07 $layer=licon1_NDIFF $count=1 $X=8.74
+ $Y=0.41 $X2=8.96 $Y2=0.325
r224 5 110 182 $w=1.7e-07 $l=2.59037e-07 $layer=licon1_NDIFF $count=1 $X=7.72
+ $Y=0.41 $X2=7.94 $Y2=0.325
r225 4 103 182 $w=1.7e-07 $l=2.41454e-07 $layer=licon1_NDIFF $count=1 $X=6.7
+ $Y=0.37 $X2=6.92 $Y2=0.325
r226 3 45 182 $w=1.7e-07 $l=2.41454e-07 $layer=licon1_NDIFF $count=1 $X=4.1
+ $Y=0.37 $X2=4.32 $Y2=0.325
r227 2 27 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=3.2 $Y=0.37
+ $X2=3.34 $Y2=0.55
r228 1 96 182 $w=1.7e-07 $l=3.4176e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.89 $Y2=0.325
.ends

.subckt PM_SKY130_FD_SC_LS__FA_4%A_734_74# 1 2 7 10 15
c26 15 0 1.62604e-19 $X=4.83 $Y=0.55
c27 10 0 1.78103e-19 $X=3.81 $Y=0.55
r28 15 17 5.30124 $w=2.48e-07 $l=1.15e-07 $layer=LI1_cond $X=4.79 $Y=0.55
+ $X2=4.79 $Y2=0.665
r29 10 12 5.30124 $w=2.48e-07 $l=1.15e-07 $layer=LI1_cond $X=3.85 $Y=0.55
+ $X2=3.85 $Y2=0.665
r30 8 12 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.975 $Y=0.665
+ $X2=3.85 $Y2=0.665
r31 7 17 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.665 $Y=0.665
+ $X2=4.79 $Y2=0.665
r32 7 8 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.665 $Y=0.665
+ $X2=3.975 $Y2=0.665
r33 2 15 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=4.69 $Y=0.37
+ $X2=4.83 $Y2=0.55
r34 1 10 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=3.67 $Y=0.37
+ $X2=3.81 $Y2=0.55
.ends

