* File: sky130_fd_sc_ls__a211o_4.pxi.spice
* Created: Fri Aug 28 12:49:13 2020
* 
x_PM_SKY130_FD_SC_LS__A211O_4%A_105_280# N_A_105_280#_M1005_d
+ N_A_105_280#_M1021_s N_A_105_280#_M1002_d N_A_105_280#_M1004_d
+ N_A_105_280#_c_140_n N_A_105_280#_M1008_g N_A_105_280#_c_124_n
+ N_A_105_280#_c_141_n N_A_105_280#_M1013_g N_A_105_280#_M1001_g
+ N_A_105_280#_c_142_n N_A_105_280#_M1016_g N_A_105_280#_c_126_n
+ N_A_105_280#_M1010_g N_A_105_280#_c_143_n N_A_105_280#_M1019_g
+ N_A_105_280#_c_127_n N_A_105_280#_M1011_g N_A_105_280#_c_128_n
+ N_A_105_280#_M1018_g N_A_105_280#_c_129_n N_A_105_280#_c_130_n
+ N_A_105_280#_c_131_n N_A_105_280#_c_132_n N_A_105_280#_c_133_n
+ N_A_105_280#_c_147_n N_A_105_280#_c_151_p N_A_105_280#_c_134_n
+ N_A_105_280#_c_174_p N_A_105_280#_c_135_n N_A_105_280#_c_136_n
+ N_A_105_280#_c_137_n N_A_105_280#_c_138_n N_A_105_280#_c_139_n
+ PM_SKY130_FD_SC_LS__A211O_4%A_105_280#
x_PM_SKY130_FD_SC_LS__A211O_4%B1 N_B1_c_294_n N_B1_M1003_g N_B1_M1005_g
+ N_B1_c_296_n N_B1_M1023_g N_B1_M1015_g N_B1_c_302_n N_B1_c_298_n B1 B1
+ PM_SKY130_FD_SC_LS__A211O_4%B1
x_PM_SKY130_FD_SC_LS__A211O_4%C1 N_C1_M1020_g N_C1_c_391_n N_C1_c_397_n
+ N_C1_M1004_g N_C1_c_392_n N_C1_c_399_n N_C1_M1009_g N_C1_c_393_n N_C1_M1021_g
+ C1 N_C1_c_395_n PM_SKY130_FD_SC_LS__A211O_4%C1
x_PM_SKY130_FD_SC_LS__A211O_4%A1 N_A1_c_457_n N_A1_M1007_g N_A1_M1002_g
+ N_A1_c_458_n N_A1_M1012_g N_A1_M1017_g A1 A1 A1 N_A1_c_456_n
+ PM_SKY130_FD_SC_LS__A211O_4%A1
x_PM_SKY130_FD_SC_LS__A211O_4%A2 N_A2_c_505_n N_A2_c_516_n N_A2_M1006_g
+ N_A2_c_506_n N_A2_c_507_n N_A2_M1000_g N_A2_c_509_n N_A2_c_510_n N_A2_c_511_n
+ N_A2_c_518_n N_A2_M1014_g N_A2_M1022_g A2 N_A2_c_514_n
+ PM_SKY130_FD_SC_LS__A211O_4%A2
x_PM_SKY130_FD_SC_LS__A211O_4%VPWR N_VPWR_M1008_d N_VPWR_M1013_d N_VPWR_M1019_d
+ N_VPWR_M1006_d N_VPWR_M1012_d N_VPWR_c_573_n N_VPWR_c_574_n N_VPWR_c_575_n
+ N_VPWR_c_576_n N_VPWR_c_577_n N_VPWR_c_578_n N_VPWR_c_579_n N_VPWR_c_580_n
+ N_VPWR_c_581_n N_VPWR_c_582_n VPWR N_VPWR_c_583_n N_VPWR_c_584_n
+ N_VPWR_c_572_n N_VPWR_c_586_n N_VPWR_c_587_n N_VPWR_c_588_n
+ PM_SKY130_FD_SC_LS__A211O_4%VPWR
x_PM_SKY130_FD_SC_LS__A211O_4%X N_X_M1001_d N_X_M1011_d N_X_M1008_s N_X_M1016_s
+ N_X_c_665_n N_X_c_671_n N_X_c_666_n N_X_c_667_n N_X_c_672_n N_X_c_668_n
+ N_X_c_673_n N_X_c_694_n N_X_c_697_n N_X_c_699_n X X N_X_c_702_n N_X_c_669_n
+ PM_SKY130_FD_SC_LS__A211O_4%X
x_PM_SKY130_FD_SC_LS__A211O_4%A_517_392# N_A_517_392#_M1003_d
+ N_A_517_392#_M1023_d N_A_517_392#_M1007_s N_A_517_392#_M1014_s
+ N_A_517_392#_c_746_n N_A_517_392#_c_748_n N_A_517_392#_c_757_n
+ N_A_517_392#_c_736_n N_A_517_392#_c_766_n N_A_517_392#_c_737_n
+ N_A_517_392#_c_738_n N_A_517_392#_c_739_n N_A_517_392#_c_740_n
+ N_A_517_392#_c_741_n N_A_517_392#_c_760_n N_A_517_392#_c_742_n
+ PM_SKY130_FD_SC_LS__A211O_4%A_517_392#
x_PM_SKY130_FD_SC_LS__A211O_4%A_602_392# N_A_602_392#_M1003_s
+ N_A_602_392#_M1009_s N_A_602_392#_c_807_n
+ PM_SKY130_FD_SC_LS__A211O_4%A_602_392#
x_PM_SKY130_FD_SC_LS__A211O_4%VGND N_VGND_M1001_s N_VGND_M1010_s N_VGND_M1018_s
+ N_VGND_M1020_d N_VGND_M1015_s N_VGND_M1022_s N_VGND_c_821_n N_VGND_c_822_n
+ N_VGND_c_823_n N_VGND_c_824_n N_VGND_c_825_n N_VGND_c_826_n N_VGND_c_827_n
+ N_VGND_c_828_n N_VGND_c_829_n N_VGND_c_830_n N_VGND_c_831_n N_VGND_c_832_n
+ VGND N_VGND_c_833_n N_VGND_c_834_n N_VGND_c_835_n N_VGND_c_836_n
+ N_VGND_c_837_n N_VGND_c_838_n N_VGND_c_839_n N_VGND_c_840_n
+ PM_SKY130_FD_SC_LS__A211O_4%VGND
x_PM_SKY130_FD_SC_LS__A211O_4%A_1064_123# N_A_1064_123#_M1000_d
+ N_A_1064_123#_M1017_s N_A_1064_123#_c_925_n N_A_1064_123#_c_922_n
+ N_A_1064_123#_c_923_n PM_SKY130_FD_SC_LS__A211O_4%A_1064_123#
cc_1 VNB N_A_105_280#_c_124_n 0.0144728f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.475
cc_2 VNB N_A_105_280#_M1001_g 0.0325584f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=0.74
cc_3 VNB N_A_105_280#_c_126_n 0.0155441f $X=-0.19 $Y=-0.245 $X2=1.63 $Y2=1.22
cc_4 VNB N_A_105_280#_c_127_n 0.0157624f $X=-0.19 $Y=-0.245 $X2=2.06 $Y2=1.22
cc_5 VNB N_A_105_280#_c_128_n 0.0176521f $X=-0.19 $Y=-0.245 $X2=2.49 $Y2=1.22
cc_6 VNB N_A_105_280#_c_129_n 0.0290413f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.475
cc_7 VNB N_A_105_280#_c_130_n 0.0104143f $X=-0.19 $Y=-0.245 $X2=2.445 $Y2=1.34
cc_8 VNB N_A_105_280#_c_131_n 0.10066f $X=-0.19 $Y=-0.245 $X2=2.13 $Y2=1.385
cc_9 VNB N_A_105_280#_c_132_n 0.00244339f $X=-0.19 $Y=-0.245 $X2=2.53 $Y2=2.06
cc_10 VNB N_A_105_280#_c_133_n 0.00983787f $X=-0.19 $Y=-0.245 $X2=3.04 $Y2=1.215
cc_11 VNB N_A_105_280#_c_134_n 0.00241387f $X=-0.19 $Y=-0.245 $X2=3.195
+ $Y2=0.615
cc_12 VNB N_A_105_280#_c_135_n 0.0138404f $X=-0.19 $Y=-0.245 $X2=5.725 $Y2=1.195
cc_13 VNB N_A_105_280#_c_136_n 0.00306752f $X=-0.19 $Y=-0.245 $X2=2.53 $Y2=1.34
cc_14 VNB N_A_105_280#_c_137_n 0.0042379f $X=-0.19 $Y=-0.245 $X2=3.195 $Y2=0.965
cc_15 VNB N_A_105_280#_c_138_n 0.00283233f $X=-0.19 $Y=-0.245 $X2=4.14 $Y2=0.895
cc_16 VNB N_A_105_280#_c_139_n 0.00225819f $X=-0.19 $Y=-0.245 $X2=5.89 $Y2=1.105
cc_17 VNB N_B1_c_294_n 0.020508f $X=-0.19 $Y=-0.245 $X2=3.055 $Y2=0.47
cc_18 VNB N_B1_M1005_g 0.0301204f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_B1_c_296_n 0.0156372f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_B1_M1015_g 0.0248495f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.765
cc_21 VNB N_B1_c_298_n 0.00156376f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=1.765
cc_22 VNB B1 0.00539681f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_C1_M1020_g 0.0210426f $X=-0.19 $Y=-0.245 $X2=5.75 $Y2=0.615
cc_24 VNB N_C1_c_391_n 0.00209214f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_C1_c_392_n 0.00180727f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_C1_c_393_n 0.0176663f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=2.4
cc_27 VNB C1 0.00323687f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=1.765
cc_28 VNB N_C1_c_395_n 0.0410167f $X=-0.19 $Y=-0.245 $X2=1.515 $Y2=2.4
cc_29 VNB N_A1_M1002_g 0.019291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A1_M1017_g 0.0193558f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.765
cc_31 VNB A1 0.00339878f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=1.475
cc_32 VNB N_A1_c_456_n 0.0270195f $X=-0.19 $Y=-0.245 $X2=1.515 $Y2=2.4
cc_33 VNB N_A2_c_505_n 0.0113836f $X=-0.19 $Y=-0.245 $X2=3.975 $Y2=0.54
cc_34 VNB N_A2_c_506_n 0.0266867f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A2_c_507_n 0.0102689f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A2_M1000_g 0.0116349f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A2_c_509_n 0.0902248f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A2_c_510_n 0.00927219f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=2.4
cc_39 VNB N_A2_c_511_n 0.0156508f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=2.4
cc_40 VNB N_A2_M1022_g 0.0375929f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=0.74
cc_41 VNB A2 0.0135013f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A2_c_514_n 0.047283f $X=-0.19 $Y=-0.245 $X2=1.515 $Y2=2.4
cc_43 VNB N_VPWR_c_572_n 0.302998f $X=-0.19 $Y=-0.245 $X2=2.53 $Y2=1.34
cc_44 VNB N_X_c_665_n 0.00104623f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=2.4
cc_45 VNB N_X_c_666_n 0.00375064f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.4
cc_46 VNB N_X_c_667_n 0.0134757f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=0.74
cc_47 VNB N_X_c_668_n 0.00178908f $X=-0.19 $Y=-0.245 $X2=1.515 $Y2=2.4
cc_48 VNB N_X_c_669_n 0.00209458f $X=-0.19 $Y=-0.245 $X2=3.66 $Y2=2.145
cc_49 VNB N_VGND_c_821_n 0.0358565f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.4
cc_50 VNB N_VGND_c_822_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=0.74
cc_51 VNB N_VGND_c_823_n 0.00250542f $X=-0.19 $Y=-0.245 $X2=1.515 $Y2=2.4
cc_52 VNB N_VGND_c_824_n 0.00634533f $X=-0.19 $Y=-0.245 $X2=1.965 $Y2=1.765
cc_53 VNB N_VGND_c_825_n 0.0100309f $X=-0.19 $Y=-0.245 $X2=2.49 $Y2=1.22
cc_54 VNB N_VGND_c_826_n 0.0131973f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_827_n 0.0495565f $X=-0.19 $Y=-0.245 $X2=2.13 $Y2=1.385
cc_56 VNB N_VGND_c_828_n 0.0282373f $X=-0.19 $Y=-0.245 $X2=2.53 $Y2=1.55
cc_57 VNB N_VGND_c_829_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=2.53 $Y2=2.06
cc_58 VNB N_VGND_c_830_n 0.0112126f $X=-0.19 $Y=-0.245 $X2=3.04 $Y2=1.215
cc_59 VNB N_VGND_c_831_n 0.0487363f $X=-0.19 $Y=-0.245 $X2=2.615 $Y2=1.215
cc_60 VNB N_VGND_c_832_n 0.00528596f $X=-0.19 $Y=-0.245 $X2=2.615 $Y2=2.145
cc_61 VNB N_VGND_c_833_n 0.0154855f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_834_n 0.0171837f $X=-0.19 $Y=-0.245 $X2=2.53 $Y2=1.34
cc_63 VNB N_VGND_c_835_n 0.0187793f $X=-0.19 $Y=-0.245 $X2=4.102 $Y2=0.895
cc_64 VNB N_VGND_c_836_n 0.422175f $X=-0.19 $Y=-0.245 $X2=1.63 $Y2=1.492
cc_65 VNB N_VGND_c_837_n 0.00601765f $X=-0.19 $Y=-0.245 $X2=2.06 $Y2=1.492
cc_66 VNB N_VGND_c_838_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_839_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_840_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_1064_123#_c_922_n 0.00186167f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_1064_123#_c_923_n 0.00326506f $X=-0.19 $Y=-0.245 $X2=0.615
+ $Y2=1.765
cc_71 VPB N_A_105_280#_c_140_n 0.0174317f $X=-0.19 $Y=1.66 $X2=0.615 $Y2=1.765
cc_72 VPB N_A_105_280#_c_141_n 0.0144458f $X=-0.19 $Y=1.66 $X2=1.065 $Y2=1.765
cc_73 VPB N_A_105_280#_c_142_n 0.0149585f $X=-0.19 $Y=1.66 $X2=1.515 $Y2=1.765
cc_74 VPB N_A_105_280#_c_143_n 0.0163149f $X=-0.19 $Y=1.66 $X2=1.965 $Y2=1.765
cc_75 VPB N_A_105_280#_c_129_n 0.00958277f $X=-0.19 $Y=1.66 $X2=0.615 $Y2=1.475
cc_76 VPB N_A_105_280#_c_131_n 0.0202335f $X=-0.19 $Y=1.66 $X2=2.13 $Y2=1.385
cc_77 VPB N_A_105_280#_c_132_n 0.00765216f $X=-0.19 $Y=1.66 $X2=2.53 $Y2=2.06
cc_78 VPB N_A_105_280#_c_147_n 0.00650326f $X=-0.19 $Y=1.66 $X2=2.615 $Y2=2.145
cc_79 VPB N_B1_c_294_n 0.0395926f $X=-0.19 $Y=1.66 $X2=3.055 $Y2=0.47
cc_80 VPB N_B1_c_296_n 0.0330788f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_B1_c_302_n 0.0121673f $X=-0.19 $Y=1.66 $X2=0.615 $Y2=2.4
cc_82 VPB N_B1_c_298_n 0.00257084f $X=-0.19 $Y=1.66 $X2=1.065 $Y2=1.765
cc_83 VPB B1 0.0061444f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_84 VPB N_C1_c_391_n 0.006437f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_C1_c_397_n 0.0210495f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_C1_c_392_n 0.00590434f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_C1_c_399_n 0.0206091f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_A1_c_457_n 0.0171333f $X=-0.19 $Y=1.66 $X2=3.055 $Y2=0.47
cc_89 VPB N_A1_c_458_n 0.0150798f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB A1 0.00962019f $X=-0.19 $Y=1.66 $X2=0.705 $Y2=1.475
cc_91 VPB N_A1_c_456_n 0.0348023f $X=-0.19 $Y=1.66 $X2=1.515 $Y2=2.4
cc_92 VPB N_A2_c_505_n 0.00854871f $X=-0.19 $Y=1.66 $X2=3.975 $Y2=0.54
cc_93 VPB N_A2_c_516_n 0.0243379f $X=-0.19 $Y=1.66 $X2=5.75 $Y2=0.615
cc_94 VPB N_A2_c_511_n 0.0113925f $X=-0.19 $Y=1.66 $X2=0.615 $Y2=2.4
cc_95 VPB N_A2_c_518_n 0.0285533f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.475
cc_96 VPB N_VPWR_c_573_n 0.0141609f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.475
cc_97 VPB N_VPWR_c_574_n 0.0647052f $X=-0.19 $Y=1.66 $X2=1.065 $Y2=1.765
cc_98 VPB N_VPWR_c_575_n 0.0185253f $X=-0.19 $Y=1.66 $X2=1.2 $Y2=0.74
cc_99 VPB N_VPWR_c_576_n 0.00514362f $X=-0.19 $Y=1.66 $X2=1.515 $Y2=2.4
cc_100 VPB N_VPWR_c_577_n 0.0206041f $X=-0.19 $Y=1.66 $X2=1.63 $Y2=1.22
cc_101 VPB N_VPWR_c_578_n 0.0103038f $X=-0.19 $Y=1.66 $X2=1.965 $Y2=2.4
cc_102 VPB N_VPWR_c_579_n 0.00640809f $X=-0.19 $Y=1.66 $X2=2.49 $Y2=0.74
cc_103 VPB N_VPWR_c_580_n 0.00329801f $X=-0.19 $Y=1.66 $X2=2.445 $Y2=1.34
cc_104 VPB N_VPWR_c_581_n 0.0160978f $X=-0.19 $Y=1.66 $X2=2.13 $Y2=1.385
cc_105 VPB N_VPWR_c_582_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_VPWR_c_583_n 0.0680039f $X=-0.19 $Y=1.66 $X2=3.04 $Y2=1.215
cc_107 VPB N_VPWR_c_584_n 0.0233618f $X=-0.19 $Y=1.66 $X2=4.245 $Y2=1.195
cc_108 VPB N_VPWR_c_572_n 0.105181f $X=-0.19 $Y=1.66 $X2=2.53 $Y2=1.34
cc_109 VPB N_VPWR_c_586_n 0.00460249f $X=-0.19 $Y=1.66 $X2=4.14 $Y2=0.895
cc_110 VPB N_VPWR_c_587_n 0.00324402f $X=-0.19 $Y=1.66 $X2=4.102 $Y2=1.195
cc_111 VPB N_VPWR_c_588_n 0.0126062f $X=-0.19 $Y=1.66 $X2=5.89 $Y2=1.105
cc_112 VPB N_X_c_665_n 5.61158e-19 $X=-0.19 $Y=1.66 $X2=0.615 $Y2=2.4
cc_113 VPB N_X_c_671_n 0.00216998f $X=-0.19 $Y=1.66 $X2=0.705 $Y2=1.475
cc_114 VPB N_X_c_672_n 0.00737223f $X=-0.19 $Y=1.66 $X2=1.2 $Y2=0.74
cc_115 VPB N_X_c_673_n 0.00257348f $X=-0.19 $Y=1.66 $X2=1.965 $Y2=1.765
cc_116 VPB N_A_517_392#_c_736_n 0.00232042f $X=-0.19 $Y=1.66 $X2=1.065 $Y2=2.4
cc_117 VPB N_A_517_392#_c_737_n 0.0023786f $X=-0.19 $Y=1.66 $X2=1.515 $Y2=1.765
cc_118 VPB N_A_517_392#_c_738_n 0.00633583f $X=-0.19 $Y=1.66 $X2=1.515 $Y2=2.4
cc_119 VPB N_A_517_392#_c_739_n 0.0129448f $X=-0.19 $Y=1.66 $X2=1.63 $Y2=0.74
cc_120 VPB N_A_517_392#_c_740_n 0.0352805f $X=-0.19 $Y=1.66 $X2=1.965 $Y2=1.765
cc_121 VPB N_A_517_392#_c_741_n 0.00459713f $X=-0.19 $Y=1.66 $X2=1.965 $Y2=2.4
cc_122 VPB N_A_517_392#_c_742_n 0.00162378f $X=-0.19 $Y=1.66 $X2=2.445 $Y2=1.34
cc_123 VPB N_A_602_392#_c_807_n 0.00824035f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 N_A_105_280#_c_131_n N_B1_c_294_n 0.00360108f $X=2.13 $Y=1.385 $X2=-0.19
+ $Y2=-0.245
cc_125 N_A_105_280#_c_132_n N_B1_c_294_n 0.00908203f $X=2.53 $Y=2.06 $X2=-0.19
+ $Y2=-0.245
cc_126 N_A_105_280#_c_133_n N_B1_c_294_n 0.00124746f $X=3.04 $Y=1.215 $X2=-0.19
+ $Y2=-0.245
cc_127 N_A_105_280#_c_151_p N_B1_c_294_n 0.013426f $X=3.66 $Y=2.145 $X2=-0.19
+ $Y2=-0.245
cc_128 N_A_105_280#_c_136_n N_B1_c_294_n 7.62508e-19 $X=2.53 $Y=1.34 $X2=-0.19
+ $Y2=-0.245
cc_129 N_A_105_280#_c_137_n N_B1_c_294_n 3.87822e-19 $X=3.195 $Y=0.965 $X2=-0.19
+ $Y2=-0.245
cc_130 N_A_105_280#_c_128_n N_B1_M1005_g 0.0217726f $X=2.49 $Y=1.22 $X2=0 $Y2=0
cc_131 N_A_105_280#_c_131_n N_B1_M1005_g 0.00124571f $X=2.13 $Y=1.385 $X2=0
+ $Y2=0
cc_132 N_A_105_280#_c_133_n N_B1_M1005_g 0.0127351f $X=3.04 $Y=1.215 $X2=0 $Y2=0
cc_133 N_A_105_280#_c_134_n N_B1_M1005_g 0.00433283f $X=3.195 $Y=0.615 $X2=0
+ $Y2=0
cc_134 N_A_105_280#_c_136_n N_B1_M1005_g 0.00427034f $X=2.53 $Y=1.34 $X2=0 $Y2=0
cc_135 N_A_105_280#_c_137_n N_B1_M1005_g 0.006532f $X=3.195 $Y=0.965 $X2=0 $Y2=0
cc_136 N_A_105_280#_c_151_p N_B1_c_296_n 2.57215e-19 $X=3.66 $Y=2.145 $X2=0
+ $Y2=0
cc_137 N_A_105_280#_c_135_n N_B1_c_296_n 8.24154e-19 $X=5.725 $Y=1.195 $X2=0
+ $Y2=0
cc_138 N_A_105_280#_c_138_n N_B1_c_296_n 4.58199e-19 $X=4.14 $Y=0.895 $X2=0
+ $Y2=0
cc_139 N_A_105_280#_c_135_n N_B1_M1015_g 0.0147131f $X=5.725 $Y=1.195 $X2=0
+ $Y2=0
cc_140 N_A_105_280#_c_138_n N_B1_M1015_g 0.00104272f $X=4.14 $Y=0.895 $X2=0
+ $Y2=0
cc_141 N_A_105_280#_c_151_p N_B1_c_302_n 0.0459576f $X=3.66 $Y=2.145 $X2=0 $Y2=0
cc_142 N_A_105_280#_c_137_n N_B1_c_302_n 0.00784836f $X=3.195 $Y=0.965 $X2=0
+ $Y2=0
cc_143 N_A_105_280#_c_132_n N_B1_c_298_n 0.0258245f $X=2.53 $Y=2.06 $X2=0 $Y2=0
cc_144 N_A_105_280#_c_133_n N_B1_c_298_n 0.0190372f $X=3.04 $Y=1.215 $X2=0 $Y2=0
cc_145 N_A_105_280#_c_151_p N_B1_c_298_n 0.0202392f $X=3.66 $Y=2.145 $X2=0 $Y2=0
cc_146 N_A_105_280#_c_136_n N_B1_c_298_n 0.00670748f $X=2.53 $Y=1.34 $X2=0 $Y2=0
cc_147 N_A_105_280#_c_137_n N_B1_c_298_n 0.00536516f $X=3.195 $Y=0.965 $X2=0
+ $Y2=0
cc_148 N_A_105_280#_c_135_n B1 0.0185247f $X=5.725 $Y=1.195 $X2=0 $Y2=0
cc_149 N_A_105_280#_c_138_n B1 0.023578f $X=4.14 $Y=0.895 $X2=0 $Y2=0
cc_150 N_A_105_280#_c_174_p N_C1_M1020_g 0.0158149f $X=3.96 $Y=0.955 $X2=0 $Y2=0
cc_151 N_A_105_280#_c_137_n N_C1_M1020_g 0.00318964f $X=3.195 $Y=0.965 $X2=0
+ $Y2=0
cc_152 N_A_105_280#_c_138_n N_C1_M1020_g 0.00147283f $X=4.14 $Y=0.895 $X2=0
+ $Y2=0
cc_153 N_A_105_280#_c_151_p N_C1_c_397_n 0.00877535f $X=3.66 $Y=2.145 $X2=0
+ $Y2=0
cc_154 N_A_105_280#_c_151_p N_C1_c_399_n 0.0026585f $X=3.66 $Y=2.145 $X2=0 $Y2=0
cc_155 N_A_105_280#_c_174_p N_C1_c_393_n 0.0164949f $X=3.96 $Y=0.955 $X2=0 $Y2=0
cc_156 N_A_105_280#_c_138_n N_C1_c_393_n 0.0122258f $X=4.14 $Y=0.895 $X2=0 $Y2=0
cc_157 N_A_105_280#_c_174_p C1 0.0230486f $X=3.96 $Y=0.955 $X2=0 $Y2=0
cc_158 N_A_105_280#_c_137_n C1 0.00690772f $X=3.195 $Y=0.965 $X2=0 $Y2=0
cc_159 N_A_105_280#_c_138_n C1 0.00525028f $X=4.14 $Y=0.895 $X2=0 $Y2=0
cc_160 N_A_105_280#_c_174_p N_C1_c_395_n 9.07417e-19 $X=3.96 $Y=0.955 $X2=0
+ $Y2=0
cc_161 N_A_105_280#_c_135_n N_A1_M1002_g 0.00877195f $X=5.725 $Y=1.195 $X2=0
+ $Y2=0
cc_162 N_A_105_280#_c_139_n N_A1_M1002_g 0.00357018f $X=5.89 $Y=1.105 $X2=0
+ $Y2=0
cc_163 N_A_105_280#_c_139_n N_A1_M1017_g 0.00370955f $X=5.89 $Y=1.105 $X2=0
+ $Y2=0
cc_164 N_A_105_280#_c_135_n A1 0.0599227f $X=5.725 $Y=1.195 $X2=0 $Y2=0
cc_165 N_A_105_280#_c_139_n A1 0.0254529f $X=5.89 $Y=1.105 $X2=0 $Y2=0
cc_166 N_A_105_280#_c_135_n N_A1_c_456_n 0.00180587f $X=5.725 $Y=1.195 $X2=0
+ $Y2=0
cc_167 N_A_105_280#_c_139_n N_A1_c_456_n 0.00226744f $X=5.89 $Y=1.105 $X2=0
+ $Y2=0
cc_168 N_A_105_280#_c_135_n N_A2_c_507_n 0.0146175f $X=5.725 $Y=1.195 $X2=0
+ $Y2=0
cc_169 N_A_105_280#_c_135_n N_A2_M1000_g 0.013753f $X=5.725 $Y=1.195 $X2=0 $Y2=0
cc_170 N_A_105_280#_c_139_n N_A2_M1000_g 5.447e-19 $X=5.89 $Y=1.105 $X2=0 $Y2=0
cc_171 N_A_105_280#_c_135_n A2 0.0108974f $X=5.725 $Y=1.195 $X2=0 $Y2=0
cc_172 N_A_105_280#_c_135_n N_A2_c_514_n 5.5067e-19 $X=5.725 $Y=1.195 $X2=0
+ $Y2=0
cc_173 N_A_105_280#_c_140_n N_VPWR_c_574_n 0.0087819f $X=0.615 $Y=1.765 $X2=0
+ $Y2=0
cc_174 N_A_105_280#_c_140_n N_VPWR_c_575_n 0.00445602f $X=0.615 $Y=1.765 $X2=0
+ $Y2=0
cc_175 N_A_105_280#_c_141_n N_VPWR_c_575_n 0.00413917f $X=1.065 $Y=1.765 $X2=0
+ $Y2=0
cc_176 N_A_105_280#_c_140_n N_VPWR_c_576_n 6.4972e-19 $X=0.615 $Y=1.765 $X2=0
+ $Y2=0
cc_177 N_A_105_280#_c_141_n N_VPWR_c_576_n 0.0150725f $X=1.065 $Y=1.765 $X2=0
+ $Y2=0
cc_178 N_A_105_280#_c_142_n N_VPWR_c_576_n 0.0069311f $X=1.515 $Y=1.765 $X2=0
+ $Y2=0
cc_179 N_A_105_280#_c_142_n N_VPWR_c_577_n 0.00445602f $X=1.515 $Y=1.765 $X2=0
+ $Y2=0
cc_180 N_A_105_280#_c_143_n N_VPWR_c_577_n 0.00445602f $X=1.965 $Y=1.765 $X2=0
+ $Y2=0
cc_181 N_A_105_280#_c_143_n N_VPWR_c_578_n 0.0095569f $X=1.965 $Y=1.765 $X2=0
+ $Y2=0
cc_182 N_A_105_280#_c_130_n N_VPWR_c_578_n 0.010202f $X=2.445 $Y=1.34 $X2=0
+ $Y2=0
cc_183 N_A_105_280#_c_131_n N_VPWR_c_578_n 0.00412269f $X=2.13 $Y=1.385 $X2=0
+ $Y2=0
cc_184 N_A_105_280#_c_132_n N_VPWR_c_578_n 0.0177407f $X=2.53 $Y=2.06 $X2=0
+ $Y2=0
cc_185 N_A_105_280#_c_147_n N_VPWR_c_578_n 0.0141316f $X=2.615 $Y=2.145 $X2=0
+ $Y2=0
cc_186 N_A_105_280#_c_140_n N_VPWR_c_572_n 0.00861395f $X=0.615 $Y=1.765 $X2=0
+ $Y2=0
cc_187 N_A_105_280#_c_141_n N_VPWR_c_572_n 0.00817726f $X=1.065 $Y=1.765 $X2=0
+ $Y2=0
cc_188 N_A_105_280#_c_142_n N_VPWR_c_572_n 0.00857589f $X=1.515 $Y=1.765 $X2=0
+ $Y2=0
cc_189 N_A_105_280#_c_143_n N_VPWR_c_572_n 0.00862391f $X=1.965 $Y=1.765 $X2=0
+ $Y2=0
cc_190 N_A_105_280#_c_124_n N_X_c_665_n 0.01145f $X=0.975 $Y=1.475 $X2=0 $Y2=0
cc_191 N_A_105_280#_c_129_n N_X_c_665_n 0.0146874f $X=0.615 $Y=1.475 $X2=0 $Y2=0
cc_192 N_A_105_280#_c_131_n N_X_c_665_n 0.00438049f $X=2.13 $Y=1.385 $X2=0 $Y2=0
cc_193 N_A_105_280#_c_140_n N_X_c_671_n 0.0125133f $X=0.615 $Y=1.765 $X2=0 $Y2=0
cc_194 N_A_105_280#_c_141_n N_X_c_671_n 0.00504132f $X=1.065 $Y=1.765 $X2=0
+ $Y2=0
cc_195 N_A_105_280#_c_124_n N_X_c_666_n 0.00172879f $X=0.975 $Y=1.475 $X2=0
+ $Y2=0
cc_196 N_A_105_280#_M1001_g N_X_c_666_n 0.0135219f $X=1.2 $Y=0.74 $X2=0 $Y2=0
cc_197 N_A_105_280#_c_131_n N_X_c_666_n 0.00873843f $X=2.13 $Y=1.385 $X2=0 $Y2=0
cc_198 N_A_105_280#_c_124_n N_X_c_667_n 0.00405513f $X=0.975 $Y=1.475 $X2=0
+ $Y2=0
cc_199 N_A_105_280#_c_129_n N_X_c_667_n 0.00100704f $X=0.615 $Y=1.475 $X2=0
+ $Y2=0
cc_200 N_A_105_280#_c_141_n N_X_c_672_n 0.0103758f $X=1.065 $Y=1.765 $X2=0 $Y2=0
cc_201 N_A_105_280#_c_142_n N_X_c_672_n 0.0101302f $X=1.515 $Y=1.765 $X2=0 $Y2=0
cc_202 N_A_105_280#_c_143_n N_X_c_672_n 0.0027144f $X=1.965 $Y=1.765 $X2=0 $Y2=0
cc_203 N_A_105_280#_c_131_n N_X_c_672_n 0.0194814f $X=2.13 $Y=1.385 $X2=0 $Y2=0
cc_204 N_A_105_280#_c_132_n N_X_c_672_n 0.00329969f $X=2.53 $Y=2.06 $X2=0 $Y2=0
cc_205 N_A_105_280#_M1001_g N_X_c_668_n 3.92313e-19 $X=1.2 $Y=0.74 $X2=0 $Y2=0
cc_206 N_A_105_280#_c_126_n N_X_c_668_n 3.92313e-19 $X=1.63 $Y=1.22 $X2=0 $Y2=0
cc_207 N_A_105_280#_c_141_n N_X_c_673_n 8.28592e-19 $X=1.065 $Y=1.765 $X2=0
+ $Y2=0
cc_208 N_A_105_280#_c_142_n N_X_c_673_n 0.0135168f $X=1.515 $Y=1.765 $X2=0 $Y2=0
cc_209 N_A_105_280#_c_143_n N_X_c_673_n 0.0127167f $X=1.965 $Y=1.765 $X2=0 $Y2=0
cc_210 N_A_105_280#_c_127_n N_X_c_694_n 0.00952589f $X=2.06 $Y=1.22 $X2=0 $Y2=0
cc_211 N_A_105_280#_c_130_n N_X_c_694_n 0.0137302f $X=2.445 $Y=1.34 $X2=0 $Y2=0
cc_212 N_A_105_280#_c_131_n N_X_c_694_n 0.0037328f $X=2.13 $Y=1.385 $X2=0 $Y2=0
cc_213 N_A_105_280#_c_140_n N_X_c_697_n 0.00418463f $X=0.615 $Y=1.765 $X2=0
+ $Y2=0
cc_214 N_A_105_280#_c_129_n N_X_c_697_n 0.00304999f $X=0.615 $Y=1.475 $X2=0
+ $Y2=0
cc_215 N_A_105_280#_c_130_n N_X_c_699_n 0.0150761f $X=2.445 $Y=1.34 $X2=0 $Y2=0
cc_216 N_A_105_280#_c_131_n N_X_c_699_n 6.02637e-19 $X=2.13 $Y=1.385 $X2=0 $Y2=0
cc_217 N_A_105_280#_c_126_n X 0.00785688f $X=1.63 $Y=1.22 $X2=0 $Y2=0
cc_218 N_A_105_280#_c_130_n N_X_c_702_n 0.0143588f $X=2.445 $Y=1.34 $X2=0 $Y2=0
cc_219 N_A_105_280#_c_131_n N_X_c_702_n 0.0185894f $X=2.13 $Y=1.385 $X2=0 $Y2=0
cc_220 N_A_105_280#_M1001_g N_X_c_669_n 0.00371782f $X=1.2 $Y=0.74 $X2=0 $Y2=0
cc_221 N_A_105_280#_c_126_n N_X_c_669_n 0.00610015f $X=1.63 $Y=1.22 $X2=0 $Y2=0
cc_222 N_A_105_280#_c_127_n N_X_c_669_n 0.00449938f $X=2.06 $Y=1.22 $X2=0 $Y2=0
cc_223 N_A_105_280#_c_130_n N_X_c_669_n 0.00966603f $X=2.445 $Y=1.34 $X2=0 $Y2=0
cc_224 N_A_105_280#_c_131_n N_X_c_669_n 8.70522e-19 $X=2.13 $Y=1.385 $X2=0 $Y2=0
cc_225 N_A_105_280#_c_132_n N_A_517_392#_M1003_d 0.00136467f $X=2.53 $Y=2.06
+ $X2=-0.19 $Y2=-0.245
cc_226 N_A_105_280#_c_147_n N_A_517_392#_M1003_d 6.03208e-19 $X=2.615 $Y=2.145
+ $X2=-0.19 $Y2=-0.245
cc_227 N_A_105_280#_c_151_p N_A_517_392#_M1003_d 0.00892986f $X=3.66 $Y=2.145
+ $X2=-0.19 $Y2=-0.245
cc_228 N_A_105_280#_M1004_d N_A_517_392#_c_746_n 0.00392274f $X=3.51 $Y=1.96
+ $X2=0 $Y2=0
cc_229 N_A_105_280#_c_151_p N_A_517_392#_c_746_n 0.0509176f $X=3.66 $Y=2.145
+ $X2=0 $Y2=0
cc_230 N_A_105_280#_c_151_p N_A_517_392#_c_748_n 0.00235846f $X=3.66 $Y=2.145
+ $X2=0 $Y2=0
cc_231 N_A_105_280#_c_147_n N_A_517_392#_c_741_n 0.00604908f $X=2.615 $Y=2.145
+ $X2=0 $Y2=0
cc_232 N_A_105_280#_c_151_p N_A_517_392#_c_741_n 0.0155391f $X=3.66 $Y=2.145
+ $X2=0 $Y2=0
cc_233 N_A_105_280#_c_151_p N_A_602_392#_M1003_s 0.00494431f $X=3.66 $Y=2.145
+ $X2=-0.19 $Y2=-0.245
cc_234 N_A_105_280#_M1004_d N_A_602_392#_c_807_n 0.00200574f $X=3.51 $Y=1.96
+ $X2=0 $Y2=0
cc_235 N_A_105_280#_c_174_p N_VGND_M1020_d 0.0044804f $X=3.96 $Y=0.955 $X2=0
+ $Y2=0
cc_236 N_A_105_280#_c_135_n N_VGND_M1015_s 0.0149463f $X=5.725 $Y=1.195 $X2=0
+ $Y2=0
cc_237 N_A_105_280#_c_124_n N_VGND_c_821_n 0.00152058f $X=0.975 $Y=1.475 $X2=0
+ $Y2=0
cc_238 N_A_105_280#_M1001_g N_VGND_c_821_n 0.0138061f $X=1.2 $Y=0.74 $X2=0 $Y2=0
cc_239 N_A_105_280#_c_126_n N_VGND_c_821_n 4.56715e-19 $X=1.63 $Y=1.22 $X2=0
+ $Y2=0
cc_240 N_A_105_280#_M1001_g N_VGND_c_822_n 0.00383152f $X=1.2 $Y=0.74 $X2=0
+ $Y2=0
cc_241 N_A_105_280#_c_126_n N_VGND_c_822_n 0.00383152f $X=1.63 $Y=1.22 $X2=0
+ $Y2=0
cc_242 N_A_105_280#_M1001_g N_VGND_c_823_n 4.05984e-19 $X=1.2 $Y=0.74 $X2=0
+ $Y2=0
cc_243 N_A_105_280#_c_126_n N_VGND_c_823_n 0.00706531f $X=1.63 $Y=1.22 $X2=0
+ $Y2=0
cc_244 N_A_105_280#_c_127_n N_VGND_c_823_n 0.00843621f $X=2.06 $Y=1.22 $X2=0
+ $Y2=0
cc_245 N_A_105_280#_c_128_n N_VGND_c_823_n 9.20677e-19 $X=2.49 $Y=1.22 $X2=0
+ $Y2=0
cc_246 N_A_105_280#_c_127_n N_VGND_c_824_n 9.69054e-19 $X=2.06 $Y=1.22 $X2=0
+ $Y2=0
cc_247 N_A_105_280#_c_128_n N_VGND_c_824_n 0.0126826f $X=2.49 $Y=1.22 $X2=0
+ $Y2=0
cc_248 N_A_105_280#_c_133_n N_VGND_c_824_n 0.0197087f $X=3.04 $Y=1.215 $X2=0
+ $Y2=0
cc_249 N_A_105_280#_c_134_n N_VGND_c_824_n 0.0189796f $X=3.195 $Y=0.615 $X2=0
+ $Y2=0
cc_250 N_A_105_280#_c_136_n N_VGND_c_824_n 0.00433174f $X=2.53 $Y=1.34 $X2=0
+ $Y2=0
cc_251 N_A_105_280#_c_134_n N_VGND_c_825_n 0.00968381f $X=3.195 $Y=0.615 $X2=0
+ $Y2=0
cc_252 N_A_105_280#_c_174_p N_VGND_c_825_n 0.0201731f $X=3.96 $Y=0.955 $X2=0
+ $Y2=0
cc_253 N_A_105_280#_c_135_n N_VGND_c_826_n 0.0218816f $X=5.725 $Y=1.195 $X2=0
+ $Y2=0
cc_254 N_A_105_280#_c_138_n N_VGND_c_826_n 0.0131078f $X=4.14 $Y=0.895 $X2=0
+ $Y2=0
cc_255 N_A_105_280#_c_127_n N_VGND_c_833_n 0.00383152f $X=2.06 $Y=1.22 $X2=0
+ $Y2=0
cc_256 N_A_105_280#_c_128_n N_VGND_c_833_n 0.00383152f $X=2.49 $Y=1.22 $X2=0
+ $Y2=0
cc_257 N_A_105_280#_c_134_n N_VGND_c_834_n 0.00751838f $X=3.195 $Y=0.615 $X2=0
+ $Y2=0
cc_258 N_A_105_280#_c_138_n N_VGND_c_835_n 0.0053849f $X=4.14 $Y=0.895 $X2=0
+ $Y2=0
cc_259 N_A_105_280#_M1001_g N_VGND_c_836_n 0.0075754f $X=1.2 $Y=0.74 $X2=0 $Y2=0
cc_260 N_A_105_280#_c_126_n N_VGND_c_836_n 0.00373265f $X=1.63 $Y=1.22 $X2=0
+ $Y2=0
cc_261 N_A_105_280#_c_127_n N_VGND_c_836_n 0.00373475f $X=2.06 $Y=1.22 $X2=0
+ $Y2=0
cc_262 N_A_105_280#_c_128_n N_VGND_c_836_n 0.0075754f $X=2.49 $Y=1.22 $X2=0
+ $Y2=0
cc_263 N_A_105_280#_c_134_n N_VGND_c_836_n 0.00822849f $X=3.195 $Y=0.615 $X2=0
+ $Y2=0
cc_264 N_A_105_280#_c_138_n N_VGND_c_836_n 0.00883028f $X=4.14 $Y=0.895 $X2=0
+ $Y2=0
cc_265 N_A_105_280#_c_135_n N_A_1064_123#_M1000_d 0.00216063f $X=5.725 $Y=1.195
+ $X2=-0.19 $Y2=-0.245
cc_266 N_A_105_280#_M1002_d N_A_1064_123#_c_925_n 0.00407798f $X=5.75 $Y=0.615
+ $X2=0 $Y2=0
cc_267 N_A_105_280#_c_135_n N_A_1064_123#_c_925_n 0.0157791f $X=5.725 $Y=1.195
+ $X2=0 $Y2=0
cc_268 N_A_105_280#_c_139_n N_A_1064_123#_c_925_n 0.015847f $X=5.89 $Y=1.105
+ $X2=0 $Y2=0
cc_269 N_A_105_280#_c_139_n N_A_1064_123#_c_923_n 0.0100053f $X=5.89 $Y=1.105
+ $X2=0 $Y2=0
cc_270 N_B1_M1005_g N_C1_M1020_g 0.0217088f $X=2.98 $Y=0.79 $X2=0 $Y2=0
cc_271 N_B1_c_294_n N_C1_c_391_n 0.00998934f $X=2.935 $Y=1.885 $X2=0 $Y2=0
cc_272 N_B1_c_302_n N_C1_c_391_n 0.00852551f $X=3.965 $Y=1.805 $X2=0 $Y2=0
cc_273 N_B1_c_298_n N_C1_c_391_n 7.13761e-19 $X=2.94 $Y=1.635 $X2=0 $Y2=0
cc_274 B1 N_C1_c_391_n 4.51928e-19 $X=3.995 $Y=1.95 $X2=0 $Y2=0
cc_275 N_B1_c_294_n N_C1_c_397_n 0.0411776f $X=2.935 $Y=1.885 $X2=0 $Y2=0
cc_276 N_B1_c_302_n N_C1_c_397_n 0.00600113f $X=3.965 $Y=1.805 $X2=0 $Y2=0
cc_277 N_B1_c_302_n N_C1_c_392_n 0.00946445f $X=3.965 $Y=1.805 $X2=0 $Y2=0
cc_278 B1 N_C1_c_392_n 0.00348543f $X=3.995 $Y=1.95 $X2=0 $Y2=0
cc_279 N_B1_c_296_n N_C1_c_399_n 0.0347373f $X=4.36 $Y=1.885 $X2=0 $Y2=0
cc_280 N_B1_c_302_n N_C1_c_399_n 0.00628739f $X=3.965 $Y=1.805 $X2=0 $Y2=0
cc_281 B1 N_C1_c_399_n 0.00405267f $X=3.995 $Y=1.95 $X2=0 $Y2=0
cc_282 N_B1_M1015_g N_C1_c_393_n 0.0226577f $X=4.375 $Y=0.935 $X2=0 $Y2=0
cc_283 N_B1_c_294_n C1 2.43307e-19 $X=2.935 $Y=1.885 $X2=0 $Y2=0
cc_284 N_B1_M1005_g C1 9.1033e-19 $X=2.98 $Y=0.79 $X2=0 $Y2=0
cc_285 N_B1_M1015_g C1 7.59958e-19 $X=4.375 $Y=0.935 $X2=0 $Y2=0
cc_286 N_B1_c_302_n C1 0.0245545f $X=3.965 $Y=1.805 $X2=0 $Y2=0
cc_287 N_B1_c_298_n C1 0.00339543f $X=2.94 $Y=1.635 $X2=0 $Y2=0
cc_288 B1 C1 0.00586513f $X=3.995 $Y=1.95 $X2=0 $Y2=0
cc_289 N_B1_c_294_n N_C1_c_395_n 0.00920115f $X=2.935 $Y=1.885 $X2=0 $Y2=0
cc_290 N_B1_c_296_n N_C1_c_395_n 0.021345f $X=4.36 $Y=1.885 $X2=0 $Y2=0
cc_291 N_B1_c_302_n N_C1_c_395_n 0.00263852f $X=3.965 $Y=1.805 $X2=0 $Y2=0
cc_292 N_B1_c_298_n N_C1_c_395_n 8.77101e-19 $X=2.94 $Y=1.635 $X2=0 $Y2=0
cc_293 B1 N_C1_c_395_n 0.00626662f $X=3.995 $Y=1.95 $X2=0 $Y2=0
cc_294 B1 A1 0.0139741f $X=3.995 $Y=1.95 $X2=0 $Y2=0
cc_295 N_B1_c_296_n N_A2_c_516_n 0.0118858f $X=4.36 $Y=1.885 $X2=0 $Y2=0
cc_296 B1 N_A2_c_516_n 0.00236668f $X=3.995 $Y=1.95 $X2=0 $Y2=0
cc_297 N_B1_c_296_n N_A2_c_507_n 0.0198771f $X=4.36 $Y=1.885 $X2=0 $Y2=0
cc_298 N_B1_M1015_g N_A2_c_507_n 0.00796009f $X=4.375 $Y=0.935 $X2=0 $Y2=0
cc_299 B1 N_A2_c_507_n 0.00126105f $X=3.995 $Y=1.95 $X2=0 $Y2=0
cc_300 N_B1_M1015_g N_A2_M1000_g 0.00842148f $X=4.375 $Y=0.935 $X2=0 $Y2=0
cc_301 N_B1_M1015_g A2 3.51473e-19 $X=4.375 $Y=0.935 $X2=0 $Y2=0
cc_302 N_B1_M1015_g N_A2_c_514_n 3.35183e-19 $X=4.375 $Y=0.935 $X2=0 $Y2=0
cc_303 N_B1_c_294_n N_VPWR_c_578_n 0.0116548f $X=2.935 $Y=1.885 $X2=0 $Y2=0
cc_304 N_B1_c_296_n N_VPWR_c_579_n 5.84978e-19 $X=4.36 $Y=1.885 $X2=0 $Y2=0
cc_305 N_B1_c_294_n N_VPWR_c_583_n 0.00337764f $X=2.935 $Y=1.885 $X2=0 $Y2=0
cc_306 N_B1_c_296_n N_VPWR_c_583_n 0.00334159f $X=4.36 $Y=1.885 $X2=0 $Y2=0
cc_307 N_B1_c_294_n N_VPWR_c_572_n 0.00444032f $X=2.935 $Y=1.885 $X2=0 $Y2=0
cc_308 N_B1_c_296_n N_VPWR_c_572_n 0.00436743f $X=4.36 $Y=1.885 $X2=0 $Y2=0
cc_309 N_B1_c_294_n N_A_517_392#_c_746_n 0.0102662f $X=2.935 $Y=1.885 $X2=0
+ $Y2=0
cc_310 N_B1_c_296_n N_A_517_392#_c_746_n 0.0111642f $X=4.36 $Y=1.885 $X2=0 $Y2=0
cc_311 N_B1_c_302_n N_A_517_392#_c_746_n 0.00380194f $X=3.965 $Y=1.805 $X2=0
+ $Y2=0
cc_312 B1 N_A_517_392#_c_746_n 0.0172389f $X=3.995 $Y=1.95 $X2=0 $Y2=0
cc_313 N_B1_c_296_n N_A_517_392#_c_748_n 0.00289278f $X=4.36 $Y=1.885 $X2=0
+ $Y2=0
cc_314 B1 N_A_517_392#_c_748_n 0.0114465f $X=3.995 $Y=1.95 $X2=0 $Y2=0
cc_315 N_B1_c_296_n N_A_517_392#_c_757_n 0.00301296f $X=4.36 $Y=1.885 $X2=0
+ $Y2=0
cc_316 N_B1_c_296_n N_A_517_392#_c_736_n 0.00444146f $X=4.36 $Y=1.885 $X2=0
+ $Y2=0
cc_317 N_B1_c_294_n N_A_517_392#_c_741_n 0.00513486f $X=2.935 $Y=1.885 $X2=0
+ $Y2=0
cc_318 N_B1_c_296_n N_A_517_392#_c_760_n 5.77764e-19 $X=4.36 $Y=1.885 $X2=0
+ $Y2=0
cc_319 B1 N_A_602_392#_M1009_s 0.0050902f $X=3.995 $Y=1.95 $X2=0 $Y2=0
cc_320 N_B1_c_294_n N_A_602_392#_c_807_n 0.00210745f $X=2.935 $Y=1.885 $X2=0
+ $Y2=0
cc_321 N_B1_c_296_n N_A_602_392#_c_807_n 0.00323776f $X=4.36 $Y=1.885 $X2=0
+ $Y2=0
cc_322 N_B1_M1005_g N_VGND_c_824_n 0.00435179f $X=2.98 $Y=0.79 $X2=0 $Y2=0
cc_323 N_B1_M1005_g N_VGND_c_825_n 4.1551e-19 $X=2.98 $Y=0.79 $X2=0 $Y2=0
cc_324 N_B1_M1015_g N_VGND_c_826_n 0.00879011f $X=4.375 $Y=0.935 $X2=0 $Y2=0
cc_325 N_B1_M1005_g N_VGND_c_834_n 0.00494504f $X=2.98 $Y=0.79 $X2=0 $Y2=0
cc_326 N_B1_M1015_g N_VGND_c_835_n 0.00349617f $X=4.375 $Y=0.935 $X2=0 $Y2=0
cc_327 N_B1_M1005_g N_VGND_c_836_n 0.00514438f $X=2.98 $Y=0.79 $X2=0 $Y2=0
cc_328 N_B1_M1015_g N_VGND_c_836_n 0.00396651f $X=4.375 $Y=0.935 $X2=0 $Y2=0
cc_329 N_C1_c_397_n N_VPWR_c_583_n 0.00290288f $X=3.435 $Y=1.885 $X2=0 $Y2=0
cc_330 N_C1_c_399_n N_VPWR_c_583_n 0.00290288f $X=3.885 $Y=1.885 $X2=0 $Y2=0
cc_331 N_C1_c_397_n N_VPWR_c_572_n 0.00359019f $X=3.435 $Y=1.885 $X2=0 $Y2=0
cc_332 N_C1_c_399_n N_VPWR_c_572_n 0.00358808f $X=3.885 $Y=1.885 $X2=0 $Y2=0
cc_333 N_C1_c_397_n N_A_517_392#_c_746_n 0.0109348f $X=3.435 $Y=1.885 $X2=0
+ $Y2=0
cc_334 N_C1_c_399_n N_A_517_392#_c_746_n 0.0123386f $X=3.885 $Y=1.885 $X2=0
+ $Y2=0
cc_335 N_C1_c_399_n N_A_517_392#_c_748_n 2.68578e-19 $X=3.885 $Y=1.885 $X2=0
+ $Y2=0
cc_336 N_C1_c_399_n N_A_517_392#_c_757_n 7.94878e-19 $X=3.885 $Y=1.885 $X2=0
+ $Y2=0
cc_337 N_C1_c_397_n N_A_517_392#_c_741_n 6.19408e-19 $X=3.435 $Y=1.885 $X2=0
+ $Y2=0
cc_338 N_C1_c_397_n N_A_602_392#_c_807_n 0.0104484f $X=3.435 $Y=1.885 $X2=0
+ $Y2=0
cc_339 N_C1_c_399_n N_A_602_392#_c_807_n 0.0104761f $X=3.885 $Y=1.885 $X2=0
+ $Y2=0
cc_340 N_C1_M1020_g N_VGND_c_825_n 0.00758501f $X=3.41 $Y=0.79 $X2=0 $Y2=0
cc_341 N_C1_c_393_n N_VGND_c_825_n 0.00282961f $X=3.9 $Y=1.29 $X2=0 $Y2=0
cc_342 N_C1_c_393_n N_VGND_c_826_n 0.00179111f $X=3.9 $Y=1.29 $X2=0 $Y2=0
cc_343 N_C1_M1020_g N_VGND_c_834_n 0.00421418f $X=3.41 $Y=0.79 $X2=0 $Y2=0
cc_344 N_C1_c_393_n N_VGND_c_835_n 0.00452791f $X=3.9 $Y=1.29 $X2=0 $Y2=0
cc_345 N_C1_M1020_g N_VGND_c_836_n 0.00432128f $X=3.41 $Y=0.79 $X2=0 $Y2=0
cc_346 N_C1_c_393_n N_VGND_c_836_n 0.00493565f $X=3.9 $Y=1.29 $X2=0 $Y2=0
cc_347 A1 N_A2_c_505_n 0.00539784f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_348 N_A1_c_456_n N_A2_c_505_n 0.00602007f $X=6.07 $Y=1.667 $X2=0 $Y2=0
cc_349 N_A1_c_457_n N_A2_c_516_n 0.00881086f $X=5.62 $Y=1.885 $X2=0 $Y2=0
cc_350 A1 N_A2_c_506_n 0.013926f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_351 N_A1_c_456_n N_A2_c_506_n 0.00197579f $X=6.07 $Y=1.667 $X2=0 $Y2=0
cc_352 N_A1_M1002_g N_A2_c_509_n 0.00985192f $X=5.675 $Y=0.935 $X2=0 $Y2=0
cc_353 N_A1_M1017_g N_A2_c_509_n 0.00985192f $X=6.105 $Y=0.935 $X2=0 $Y2=0
cc_354 N_A1_M1017_g N_A2_c_510_n 0.011445f $X=6.105 $Y=0.935 $X2=0 $Y2=0
cc_355 A1 N_A2_c_510_n 0.00183891f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_356 N_A1_c_456_n N_A2_c_511_n 0.0170847f $X=6.07 $Y=1.667 $X2=0 $Y2=0
cc_357 N_A1_c_458_n N_A2_c_518_n 0.0197382f $X=6.07 $Y=1.885 $X2=0 $Y2=0
cc_358 N_A1_M1017_g N_A2_M1022_g 0.0119526f $X=6.105 $Y=0.935 $X2=0 $Y2=0
cc_359 N_A1_M1002_g N_A2_c_514_n 0.0302298f $X=5.675 $Y=0.935 $X2=0 $Y2=0
cc_360 N_A1_c_457_n N_VPWR_c_579_n 0.0100617f $X=5.62 $Y=1.885 $X2=0 $Y2=0
cc_361 N_A1_c_458_n N_VPWR_c_579_n 4.69752e-19 $X=6.07 $Y=1.885 $X2=0 $Y2=0
cc_362 N_A1_c_457_n N_VPWR_c_580_n 5.07136e-19 $X=5.62 $Y=1.885 $X2=0 $Y2=0
cc_363 N_A1_c_458_n N_VPWR_c_580_n 0.011138f $X=6.07 $Y=1.885 $X2=0 $Y2=0
cc_364 N_A1_c_457_n N_VPWR_c_581_n 0.00429299f $X=5.62 $Y=1.885 $X2=0 $Y2=0
cc_365 N_A1_c_458_n N_VPWR_c_581_n 0.00413917f $X=6.07 $Y=1.885 $X2=0 $Y2=0
cc_366 N_A1_c_457_n N_VPWR_c_572_n 0.00847721f $X=5.62 $Y=1.885 $X2=0 $Y2=0
cc_367 N_A1_c_458_n N_VPWR_c_572_n 0.00817726f $X=6.07 $Y=1.885 $X2=0 $Y2=0
cc_368 N_A1_c_457_n N_A_517_392#_c_766_n 0.014438f $X=5.62 $Y=1.885 $X2=0 $Y2=0
cc_369 A1 N_A_517_392#_c_766_n 0.0382707f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_370 N_A1_c_458_n N_A_517_392#_c_738_n 0.0136012f $X=6.07 $Y=1.885 $X2=0 $Y2=0
cc_371 A1 N_A_517_392#_c_738_n 0.0111998f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_372 N_A1_c_456_n N_A_517_392#_c_738_n 0.00250266f $X=6.07 $Y=1.667 $X2=0
+ $Y2=0
cc_373 N_A1_c_457_n N_A_517_392#_c_742_n 0.00625797f $X=5.62 $Y=1.885 $X2=0
+ $Y2=0
cc_374 A1 N_A_517_392#_c_742_n 0.0231322f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_375 N_A1_c_456_n N_A_517_392#_c_742_n 0.00683203f $X=6.07 $Y=1.667 $X2=0
+ $Y2=0
cc_376 N_A1_M1017_g N_VGND_c_827_n 5.60436e-19 $X=6.105 $Y=0.935 $X2=0 $Y2=0
cc_377 N_A1_M1002_g N_VGND_c_836_n 9.15321e-19 $X=5.675 $Y=0.935 $X2=0 $Y2=0
cc_378 N_A1_M1017_g N_VGND_c_836_n 9.15321e-19 $X=6.105 $Y=0.935 $X2=0 $Y2=0
cc_379 N_A1_M1002_g N_A_1064_123#_c_925_n 0.00929401f $X=5.675 $Y=0.935 $X2=0
+ $Y2=0
cc_380 N_A1_M1017_g N_A_1064_123#_c_925_n 0.0116895f $X=6.105 $Y=0.935 $X2=0
+ $Y2=0
cc_381 A1 N_A_1064_123#_c_925_n 0.00154834f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_382 N_A1_M1017_g N_A_1064_123#_c_922_n 4.59247e-19 $X=6.105 $Y=0.935 $X2=0
+ $Y2=0
cc_383 N_A2_c_516_n N_VPWR_c_579_n 0.0101755f $X=4.815 $Y=1.885 $X2=0 $Y2=0
cc_384 N_A2_c_518_n N_VPWR_c_580_n 0.0141474f $X=6.52 $Y=1.885 $X2=0 $Y2=0
cc_385 N_A2_c_516_n N_VPWR_c_583_n 0.00429299f $X=4.815 $Y=1.885 $X2=0 $Y2=0
cc_386 N_A2_c_518_n N_VPWR_c_584_n 0.00413917f $X=6.52 $Y=1.885 $X2=0 $Y2=0
cc_387 N_A2_c_516_n N_VPWR_c_572_n 0.0084785f $X=4.815 $Y=1.885 $X2=0 $Y2=0
cc_388 N_A2_c_518_n N_VPWR_c_572_n 0.00821673f $X=6.52 $Y=1.885 $X2=0 $Y2=0
cc_389 N_A2_c_516_n N_A_517_392#_c_736_n 2.32562e-19 $X=4.815 $Y=1.885 $X2=0
+ $Y2=0
cc_390 N_A2_c_516_n N_A_517_392#_c_766_n 0.0186387f $X=4.815 $Y=1.885 $X2=0
+ $Y2=0
cc_391 N_A2_c_506_n N_A_517_392#_c_766_n 0.00140678f $X=5.17 $Y=1.405 $X2=0
+ $Y2=0
cc_392 N_A2_c_518_n N_A_517_392#_c_738_n 0.0162564f $X=6.52 $Y=1.885 $X2=0 $Y2=0
cc_393 N_A2_c_518_n N_A_517_392#_c_739_n 0.00248775f $X=6.52 $Y=1.885 $X2=0
+ $Y2=0
cc_394 N_A2_c_518_n N_A_517_392#_c_740_n 4.53441e-19 $X=6.52 $Y=1.885 $X2=0
+ $Y2=0
cc_395 A2 N_VGND_M1015_s 0.00344879f $X=4.955 $Y=0.47 $X2=0 $Y2=0
cc_396 N_A2_M1000_g N_VGND_c_826_n 0.00390703f $X=5.245 $Y=0.935 $X2=0 $Y2=0
cc_397 A2 N_VGND_c_826_n 0.0343402f $X=4.955 $Y=0.47 $X2=0 $Y2=0
cc_398 N_A2_c_514_n N_VGND_c_826_n 0.0052481f $X=5.155 $Y=0.2 $X2=0 $Y2=0
cc_399 N_A2_c_509_n N_VGND_c_827_n 0.00811888f $X=6.46 $Y=0.2 $X2=0 $Y2=0
cc_400 N_A2_M1022_g N_VGND_c_827_n 0.0259975f $X=6.535 $Y=0.935 $X2=0 $Y2=0
cc_401 A2 N_VGND_c_831_n 0.0257682f $X=4.955 $Y=0.47 $X2=0 $Y2=0
cc_402 N_A2_c_514_n N_VGND_c_831_n 0.0403962f $X=5.155 $Y=0.2 $X2=0 $Y2=0
cc_403 N_A2_c_509_n N_VGND_c_836_n 0.0406735f $X=6.46 $Y=0.2 $X2=0 $Y2=0
cc_404 A2 N_VGND_c_836_n 0.0135719f $X=4.955 $Y=0.47 $X2=0 $Y2=0
cc_405 N_A2_c_514_n N_VGND_c_836_n 0.0100036f $X=5.155 $Y=0.2 $X2=0 $Y2=0
cc_406 N_A2_M1000_g N_A_1064_123#_c_925_n 0.00405878f $X=5.245 $Y=0.935 $X2=0
+ $Y2=0
cc_407 N_A2_c_509_n N_A_1064_123#_c_925_n 0.00827463f $X=6.46 $Y=0.2 $X2=0 $Y2=0
cc_408 A2 N_A_1064_123#_c_925_n 0.00164856f $X=4.955 $Y=0.47 $X2=0 $Y2=0
cc_409 N_A2_c_509_n N_A_1064_123#_c_922_n 0.00275881f $X=6.46 $Y=0.2 $X2=0 $Y2=0
cc_410 N_VPWR_c_574_n N_X_c_671_n 0.0715879f $X=0.39 $Y=1.985 $X2=0 $Y2=0
cc_411 N_VPWR_c_575_n N_X_c_671_n 0.0110241f $X=1.125 $Y=3.33 $X2=0 $Y2=0
cc_412 N_VPWR_c_576_n N_X_c_671_n 0.060454f $X=1.29 $Y=2.225 $X2=0 $Y2=0
cc_413 N_VPWR_c_572_n N_X_c_671_n 0.00909194f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_414 N_VPWR_M1013_d N_X_c_672_n 0.00222494f $X=1.14 $Y=1.84 $X2=0 $Y2=0
cc_415 N_VPWR_c_576_n N_X_c_672_n 0.0154248f $X=1.29 $Y=2.225 $X2=0 $Y2=0
cc_416 N_VPWR_c_578_n N_X_c_672_n 0.00487617f $X=2.19 $Y=1.985 $X2=0 $Y2=0
cc_417 N_VPWR_c_576_n N_X_c_673_n 0.0617165f $X=1.29 $Y=2.225 $X2=0 $Y2=0
cc_418 N_VPWR_c_577_n N_X_c_673_n 0.014552f $X=2.105 $Y=3.33 $X2=0 $Y2=0
cc_419 N_VPWR_c_578_n N_X_c_673_n 0.0709936f $X=2.19 $Y=1.985 $X2=0 $Y2=0
cc_420 N_VPWR_c_572_n N_X_c_673_n 0.0119791f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_421 N_VPWR_c_574_n N_X_c_697_n 0.00501285f $X=0.39 $Y=1.985 $X2=0 $Y2=0
cc_422 N_VPWR_c_583_n N_A_517_392#_c_746_n 0.00340729f $X=4.88 $Y=3.33 $X2=0
+ $Y2=0
cc_423 N_VPWR_c_572_n N_A_517_392#_c_746_n 0.00814829f $X=6.96 $Y=3.33 $X2=0
+ $Y2=0
cc_424 N_VPWR_c_579_n N_A_517_392#_c_736_n 0.0187075f $X=5.39 $Y=2.485 $X2=0
+ $Y2=0
cc_425 N_VPWR_c_583_n N_A_517_392#_c_736_n 0.00966867f $X=4.88 $Y=3.33 $X2=0
+ $Y2=0
cc_426 N_VPWR_c_572_n N_A_517_392#_c_736_n 0.007728f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_427 N_VPWR_M1006_d N_A_517_392#_c_766_n 0.0152098f $X=4.89 $Y=1.96 $X2=0
+ $Y2=0
cc_428 N_VPWR_c_579_n N_A_517_392#_c_766_n 0.0453019f $X=5.39 $Y=2.485 $X2=0
+ $Y2=0
cc_429 N_VPWR_c_579_n N_A_517_392#_c_737_n 0.0250292f $X=5.39 $Y=2.485 $X2=0
+ $Y2=0
cc_430 N_VPWR_c_580_n N_A_517_392#_c_737_n 0.0266413f $X=6.295 $Y=2.375 $X2=0
+ $Y2=0
cc_431 N_VPWR_c_581_n N_A_517_392#_c_737_n 0.0103967f $X=6.13 $Y=3.33 $X2=0
+ $Y2=0
cc_432 N_VPWR_c_572_n N_A_517_392#_c_737_n 0.00860547f $X=6.96 $Y=3.33 $X2=0
+ $Y2=0
cc_433 N_VPWR_M1012_d N_A_517_392#_c_738_n 0.00197722f $X=6.145 $Y=1.96 $X2=0
+ $Y2=0
cc_434 N_VPWR_c_580_n N_A_517_392#_c_738_n 0.0171814f $X=6.295 $Y=2.375 $X2=0
+ $Y2=0
cc_435 N_VPWR_c_580_n N_A_517_392#_c_740_n 0.0266615f $X=6.295 $Y=2.375 $X2=0
+ $Y2=0
cc_436 N_VPWR_c_584_n N_A_517_392#_c_740_n 0.0124046f $X=6.96 $Y=3.33 $X2=0
+ $Y2=0
cc_437 N_VPWR_c_572_n N_A_517_392#_c_740_n 0.0102675f $X=6.96 $Y=3.33 $X2=0
+ $Y2=0
cc_438 N_VPWR_c_578_n N_A_517_392#_c_741_n 0.0212872f $X=2.19 $Y=1.985 $X2=0
+ $Y2=0
cc_439 N_VPWR_c_583_n N_A_517_392#_c_741_n 0.00681978f $X=4.88 $Y=3.33 $X2=0
+ $Y2=0
cc_440 N_VPWR_c_572_n N_A_517_392#_c_741_n 0.0102611f $X=6.96 $Y=3.33 $X2=0
+ $Y2=0
cc_441 N_VPWR_c_583_n N_A_517_392#_c_760_n 7.17652e-19 $X=4.88 $Y=3.33 $X2=0
+ $Y2=0
cc_442 N_VPWR_c_572_n N_A_517_392#_c_760_n 0.00209261f $X=6.96 $Y=3.33 $X2=0
+ $Y2=0
cc_443 N_VPWR_c_583_n N_A_602_392#_c_807_n 0.053277f $X=4.88 $Y=3.33 $X2=0 $Y2=0
cc_444 N_VPWR_c_572_n N_A_602_392#_c_807_n 0.0436645f $X=6.96 $Y=3.33 $X2=0
+ $Y2=0
cc_445 N_X_c_694_n N_VGND_M1010_s 0.00386728f $X=2.18 $Y=0.875 $X2=0 $Y2=0
cc_446 X N_VGND_M1010_s 3.57684e-19 $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_447 N_X_c_669_n N_VGND_M1010_s 0.00197831f $X=1.415 $Y=0.965 $X2=0 $Y2=0
cc_448 N_X_c_666_n N_VGND_c_821_n 0.0144939f $X=1.33 $Y=1.325 $X2=0 $Y2=0
cc_449 N_X_c_667_n N_VGND_c_821_n 0.00888458f $X=0.925 $Y=1.325 $X2=0 $Y2=0
cc_450 N_X_c_668_n N_VGND_c_821_n 0.0164567f $X=1.415 $Y=0.515 $X2=0 $Y2=0
cc_451 N_X_c_668_n N_VGND_c_822_n 0.00749631f $X=1.415 $Y=0.515 $X2=0 $Y2=0
cc_452 N_X_c_668_n N_VGND_c_823_n 0.0103637f $X=1.415 $Y=0.515 $X2=0 $Y2=0
cc_453 N_X_c_694_n N_VGND_c_823_n 0.0122752f $X=2.18 $Y=0.875 $X2=0 $Y2=0
cc_454 X N_VGND_c_823_n 0.00479967f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_455 N_X_c_699_n N_VGND_c_833_n 0.00408057f $X=2.275 $Y=0.745 $X2=0 $Y2=0
cc_456 N_X_c_668_n N_VGND_c_836_n 0.0062048f $X=1.415 $Y=0.515 $X2=0 $Y2=0
cc_457 N_X_c_694_n N_VGND_c_836_n 0.00594702f $X=2.18 $Y=0.875 $X2=0 $Y2=0
cc_458 N_X_c_699_n N_VGND_c_836_n 0.00596517f $X=2.275 $Y=0.745 $X2=0 $Y2=0
cc_459 X N_VGND_c_836_n 0.00681138f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_460 N_A_517_392#_c_746_n N_A_602_392#_M1003_s 0.00493283f $X=4.42 $Y=2.485
+ $X2=-0.19 $Y2=1.66
cc_461 N_A_517_392#_c_746_n N_A_602_392#_M1009_s 0.00496373f $X=4.42 $Y=2.485
+ $X2=0 $Y2=0
cc_462 N_A_517_392#_c_746_n N_A_602_392#_c_807_n 0.0669824f $X=4.42 $Y=2.485
+ $X2=0 $Y2=0
cc_463 N_A_517_392#_c_736_n N_A_602_392#_c_807_n 0.017478f $X=4.585 $Y=2.825
+ $X2=0 $Y2=0
cc_464 N_A_517_392#_c_739_n N_VGND_c_827_n 0.0113511f $X=6.77 $Y=2.12 $X2=0
+ $Y2=0
cc_465 N_A_517_392#_c_738_n N_A_1064_123#_c_923_n 0.00539705f $X=6.58 $Y=2.035
+ $X2=0 $Y2=0
cc_466 N_VGND_c_826_n N_A_1064_123#_c_925_n 0.00559098f $X=4.59 $Y=0.765 $X2=0
+ $Y2=0
cc_467 N_VGND_c_831_n N_A_1064_123#_c_925_n 0.0122684f $X=6.585 $Y=0 $X2=0 $Y2=0
cc_468 N_VGND_c_836_n N_A_1064_123#_c_925_n 0.0214259f $X=6.96 $Y=0 $X2=0 $Y2=0
cc_469 N_VGND_c_827_n N_A_1064_123#_c_922_n 0.0096909f $X=6.75 $Y=0.76 $X2=0
+ $Y2=0
cc_470 N_VGND_c_831_n N_A_1064_123#_c_922_n 0.00374365f $X=6.585 $Y=0 $X2=0
+ $Y2=0
cc_471 N_VGND_c_836_n N_A_1064_123#_c_922_n 0.00464028f $X=6.96 $Y=0 $X2=0 $Y2=0
cc_472 N_VGND_c_827_n N_A_1064_123#_c_923_n 0.0160983f $X=6.75 $Y=0.76 $X2=0
+ $Y2=0
