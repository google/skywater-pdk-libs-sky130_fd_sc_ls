* File: sky130_fd_sc_ls__dlclkp_1.pxi.spice
* Created: Wed Sep  2 11:02:47 2020
* 
x_PM_SKY130_FD_SC_LS__DLCLKP_1%A_83_260# N_A_83_260#_M1019_d N_A_83_260#_M1013_d
+ N_A_83_260#_M1015_g N_A_83_260#_c_122_n N_A_83_260#_M1010_g
+ N_A_83_260#_c_123_n N_A_83_260#_c_124_n N_A_83_260#_c_125_n
+ N_A_83_260#_c_133_p N_A_83_260#_c_184_p N_A_83_260#_c_126_n
+ N_A_83_260#_c_134_p N_A_83_260#_c_180_p N_A_83_260#_c_147_p
+ N_A_83_260#_c_135_p N_A_83_260#_c_148_p PM_SKY130_FD_SC_LS__DLCLKP_1%A_83_260#
x_PM_SKY130_FD_SC_LS__DLCLKP_1%GATE N_GATE_c_205_n N_GATE_M1017_g N_GATE_M1018_g
+ GATE PM_SKY130_FD_SC_LS__DLCLKP_1%GATE
x_PM_SKY130_FD_SC_LS__DLCLKP_1%A_315_54# N_A_315_54#_M1002_s N_A_315_54#_M1004_s
+ N_A_315_54#_c_244_n N_A_315_54#_M1019_g N_A_315_54#_c_251_n
+ N_A_315_54#_M1006_g N_A_315_54#_c_245_n N_A_315_54#_M1016_g
+ N_A_315_54#_M1003_g N_A_315_54#_c_247_n N_A_315_54#_c_248_n
+ N_A_315_54#_c_254_n N_A_315_54#_c_270_n N_A_315_54#_c_255_n
+ N_A_315_54#_c_256_n N_A_315_54#_c_249_n N_A_315_54#_c_258_n
+ N_A_315_54#_c_259_n N_A_315_54#_c_250_n N_A_315_54#_c_327_p
+ PM_SKY130_FD_SC_LS__DLCLKP_1%A_315_54#
x_PM_SKY130_FD_SC_LS__DLCLKP_1%A_309_338# N_A_309_338#_M1003_d
+ N_A_309_338#_M1016_d N_A_309_338#_c_367_n N_A_309_338#_M1013_g
+ N_A_309_338#_c_368_n N_A_309_338#_c_369_n N_A_309_338#_M1001_g
+ N_A_309_338#_c_360_n N_A_309_338#_c_361_n N_A_309_338#_c_362_n
+ N_A_309_338#_c_363_n N_A_309_338#_c_364_n N_A_309_338#_c_365_n
+ N_A_309_338#_c_373_n N_A_309_338#_c_366_n
+ PM_SKY130_FD_SC_LS__DLCLKP_1%A_309_338#
x_PM_SKY130_FD_SC_LS__DLCLKP_1%CLK N_CLK_c_440_n N_CLK_M1004_g N_CLK_c_436_n
+ N_CLK_M1002_g N_CLK_M1011_g N_CLK_c_441_n N_CLK_M1009_g CLK CLK N_CLK_c_439_n
+ PM_SKY130_FD_SC_LS__DLCLKP_1%CLK
x_PM_SKY130_FD_SC_LS__DLCLKP_1%A_27_74# N_A_27_74#_M1015_s N_A_27_74#_M1010_s
+ N_A_27_74#_M1014_g N_A_27_74#_c_497_n N_A_27_74#_c_498_n N_A_27_74#_M1005_g
+ N_A_27_74#_c_484_n N_A_27_74#_M1008_g N_A_27_74#_c_486_n N_A_27_74#_c_500_n
+ N_A_27_74#_M1007_g N_A_27_74#_c_487_n N_A_27_74#_c_488_n N_A_27_74#_c_502_n
+ N_A_27_74#_c_489_n N_A_27_74#_c_490_n N_A_27_74#_c_503_n N_A_27_74#_c_510_n
+ N_A_27_74#_c_514_n N_A_27_74#_c_491_n N_A_27_74#_c_492_n N_A_27_74#_c_504_n
+ N_A_27_74#_c_493_n N_A_27_74#_c_494_n N_A_27_74#_c_495_n N_A_27_74#_c_496_n
+ PM_SKY130_FD_SC_LS__DLCLKP_1%A_27_74#
x_PM_SKY130_FD_SC_LS__DLCLKP_1%A_987_393# N_A_987_393#_M1008_d
+ N_A_987_393#_M1009_d N_A_987_393#_c_623_n N_A_987_393#_M1000_g
+ N_A_987_393#_M1012_g N_A_987_393#_c_625_n N_A_987_393#_c_626_n
+ N_A_987_393#_c_627_n N_A_987_393#_c_628_n N_A_987_393#_c_632_n
+ N_A_987_393#_c_638_n N_A_987_393#_c_629_n
+ PM_SKY130_FD_SC_LS__DLCLKP_1%A_987_393#
x_PM_SKY130_FD_SC_LS__DLCLKP_1%VPWR N_VPWR_M1010_d N_VPWR_M1005_d N_VPWR_M1004_d
+ N_VPWR_M1007_d N_VPWR_c_688_n N_VPWR_c_689_n N_VPWR_c_690_n N_VPWR_c_691_n
+ N_VPWR_c_692_n N_VPWR_c_693_n VPWR N_VPWR_c_694_n N_VPWR_c_695_n
+ N_VPWR_c_696_n N_VPWR_c_697_n N_VPWR_c_687_n N_VPWR_c_699_n N_VPWR_c_700_n
+ N_VPWR_c_701_n PM_SKY130_FD_SC_LS__DLCLKP_1%VPWR
x_PM_SKY130_FD_SC_LS__DLCLKP_1%GCLK N_GCLK_M1012_d N_GCLK_M1000_d N_GCLK_c_773_n
+ GCLK GCLK GCLK GCLK N_GCLK_c_776_n PM_SKY130_FD_SC_LS__DLCLKP_1%GCLK
x_PM_SKY130_FD_SC_LS__DLCLKP_1%VGND N_VGND_M1015_d N_VGND_M1014_d N_VGND_M1002_d
+ N_VGND_M1012_s N_VGND_c_791_n N_VGND_c_806_n N_VGND_c_792_n N_VGND_c_793_n
+ N_VGND_c_794_n N_VGND_c_795_n N_VGND_c_796_n VGND N_VGND_c_797_n
+ N_VGND_c_798_n N_VGND_c_799_n N_VGND_c_800_n N_VGND_c_801_n N_VGND_c_802_n
+ N_VGND_c_803_n N_VGND_c_804_n PM_SKY130_FD_SC_LS__DLCLKP_1%VGND
cc_1 VNB N_A_83_260#_M1015_g 0.030146f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_A_83_260#_c_122_n 0.0376037f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_3 VNB N_A_83_260#_c_123_n 0.00759181f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.63
cc_4 VNB N_A_83_260#_c_124_n 4.07393e-19 $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.97
cc_5 VNB N_A_83_260#_c_125_n 0.0146521f $X=-0.19 $Y=-0.245 $X2=1.385 $Y2=1.215
cc_6 VNB N_A_83_260#_c_126_n 0.00159251f $X=-0.19 $Y=-0.245 $X2=1.47 $Y2=1.13
cc_7 VNB N_GATE_c_205_n 0.0205983f $X=-0.19 $Y=-0.245 $X2=1.725 $Y2=0.4
cc_8 VNB N_GATE_M1018_g 0.0345308f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB GATE 0.00166024f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_10 VNB N_A_315_54#_c_244_n 0.0180708f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.3
cc_11 VNB N_A_315_54#_c_245_n 0.025399f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_12 VNB N_A_315_54#_M1003_g 0.0207868f $X=-0.19 $Y=-0.245 $X2=1.385 $Y2=2.055
cc_13 VNB N_A_315_54#_c_247_n 0.00535921f $X=-0.19 $Y=-0.245 $X2=1.47 $Y2=2.14
cc_14 VNB N_A_315_54#_c_248_n 0.0395251f $X=-0.19 $Y=-0.245 $X2=1.47 $Y2=2.55
cc_15 VNB N_A_315_54#_c_249_n 0.0132503f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.465
cc_16 VNB N_A_315_54#_c_250_n 0.00584675f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_309_338#_M1001_g 0.0339887f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.63
cc_18 VNB N_A_309_338#_c_360_n 0.00319078f $X=-0.19 $Y=-0.245 $X2=1.385
+ $Y2=2.055
cc_19 VNB N_A_309_338#_c_361_n 0.0165635f $X=-0.19 $Y=-0.245 $X2=0.785 $Y2=2.055
cc_20 VNB N_A_309_338#_c_362_n 0.0152503f $X=-0.19 $Y=-0.245 $X2=1.47 $Y2=1.13
cc_21 VNB N_A_309_338#_c_363_n 0.00748342f $X=-0.19 $Y=-0.245 $X2=1.47 $Y2=2.14
cc_22 VNB N_A_309_338#_c_364_n 0.0105451f $X=-0.19 $Y=-0.245 $X2=1.98 $Y2=0.815
cc_23 VNB N_A_309_338#_c_365_n 0.00878008f $X=-0.19 $Y=-0.245 $X2=1.555
+ $Y2=2.715
cc_24 VNB N_A_309_338#_c_366_n 0.00173862f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.465
cc_25 VNB N_CLK_c_436_n 0.0187791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_CLK_M1011_g 0.0209903f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_27 VNB CLK 0.0101706f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.97
cc_28 VNB N_CLK_c_439_n 0.0418332f $X=-0.19 $Y=-0.245 $X2=1.47 $Y2=2.55
cc_29 VNB N_A_27_74#_M1014_g 0.0108504f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_27_74#_c_484_n 0.184715f $X=-0.19 $Y=-0.245 $X2=1.385 $Y2=2.055
cc_31 VNB N_A_27_74#_M1008_g 0.0294989f $X=-0.19 $Y=-0.245 $X2=1.47 $Y2=2.55
cc_32 VNB N_A_27_74#_c_486_n 0.0092132f $X=-0.19 $Y=-0.245 $X2=1.98 $Y2=0.815
cc_33 VNB N_A_27_74#_c_487_n 0.015735f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_27_74#_c_488_n 0.0271016f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.465
cc_35 VNB N_A_27_74#_c_489_n 0.0136994f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.465
cc_36 VNB N_A_27_74#_c_490_n 0.0199695f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_27_74#_c_491_n 0.0022869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_27_74#_c_492_n 0.019497f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_27_74#_c_493_n 0.0246006f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_27_74#_c_494_n 0.00496022f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_27_74#_c_495_n 0.025466f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_27_74#_c_496_n 0.0493903f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_987_393#_c_623_n 0.0244484f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.3
cc_44 VNB N_A_987_393#_M1012_g 0.0293558f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_45 VNB N_A_987_393#_c_625_n 0.038908f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.97
cc_46 VNB N_A_987_393#_c_626_n 0.00849579f $X=-0.19 $Y=-0.245 $X2=1.47 $Y2=0.98
cc_47 VNB N_A_987_393#_c_627_n 3.54303e-19 $X=-0.19 $Y=-0.245 $X2=1.47 $Y2=2.55
cc_48 VNB N_A_987_393#_c_628_n 0.00663381f $X=-0.19 $Y=-0.245 $X2=1.98 $Y2=0.815
cc_49 VNB N_A_987_393#_c_629_n 0.00656085f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.465
cc_50 VNB N_VPWR_c_687_n 0.283096f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_GCLK_c_773_n 0.0505628f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_52 VNB GCLK 0.00521116f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_53 VNB N_VGND_c_791_n 0.00805223f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.97
cc_54 VNB N_VGND_c_792_n 0.0115327f $X=-0.19 $Y=-0.245 $X2=1.47 $Y2=2.14
cc_55 VNB N_VGND_c_793_n 0.0153007f $X=-0.19 $Y=-0.245 $X2=1.98 $Y2=0.815
cc_56 VNB N_VGND_c_794_n 0.0196172f $X=-0.19 $Y=-0.245 $X2=1.99 $Y2=2.715
cc_57 VNB N_VGND_c_795_n 0.0517199f $X=-0.19 $Y=-0.245 $X2=0.785 $Y2=1.215
cc_58 VNB N_VGND_c_796_n 0.00226387f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.465
cc_59 VNB N_VGND_c_797_n 0.0193135f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.465
cc_60 VNB N_VGND_c_798_n 0.0310734f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_799_n 0.0332986f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_800_n 0.0194697f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_801_n 0.364249f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_802_n 0.00478372f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_803_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_804_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VPB N_A_83_260#_c_122_n 0.0301608f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_68 VPB N_A_83_260#_c_124_n 0.00292699f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.97
cc_69 VPB N_GATE_c_205_n 0.039028f $X=-0.19 $Y=1.66 $X2=1.725 $Y2=0.4
cc_70 VPB GATE 0.00137271f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_71 VPB N_A_315_54#_c_251_n 0.0552606f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_A_315_54#_c_245_n 0.0334719f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_73 VPB N_A_315_54#_c_247_n 0.00920932f $X=-0.19 $Y=1.66 $X2=1.47 $Y2=2.14
cc_74 VPB N_A_315_54#_c_254_n 0.0231456f $X=-0.19 $Y=1.66 $X2=1.98 $Y2=0.815
cc_75 VPB N_A_315_54#_c_255_n 0.0029468f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_A_315_54#_c_256_n 0.0199098f $X=-0.19 $Y=1.66 $X2=0.785 $Y2=1.215
cc_77 VPB N_A_315_54#_c_249_n 0.00331749f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.465
cc_78 VPB N_A_315_54#_c_258_n 0.00244941f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 VPB N_A_315_54#_c_259_n 0.00338564f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 VPB N_A_315_54#_c_250_n 0.00100914f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_A_309_338#_c_367_n 0.0173488f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.3
cc_82 VPB N_A_309_338#_c_368_n 0.0321781f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 VPB N_A_309_338#_c_369_n 0.0128531f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_84 VPB N_A_309_338#_c_360_n 0.00243131f $X=-0.19 $Y=1.66 $X2=1.385 $Y2=2.055
cc_85 VPB N_A_309_338#_c_361_n 0.0146979f $X=-0.19 $Y=1.66 $X2=0.785 $Y2=2.055
cc_86 VPB N_A_309_338#_c_365_n 0.00514213f $X=-0.19 $Y=1.66 $X2=1.555 $Y2=2.715
cc_87 VPB N_A_309_338#_c_373_n 0.00292336f $X=-0.19 $Y=1.66 $X2=0.785 $Y2=1.215
cc_88 VPB N_CLK_c_440_n 0.01932f $X=-0.19 $Y=1.66 $X2=1.725 $Y2=0.4
cc_89 VPB N_CLK_c_441_n 0.015908f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_90 VPB CLK 0.00294547f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.97
cc_91 VPB N_CLK_c_439_n 0.0247209f $X=-0.19 $Y=1.66 $X2=1.47 $Y2=2.55
cc_92 VPB N_A_27_74#_c_497_n 0.00661569f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_93 VPB N_A_27_74#_c_498_n 0.0235063f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_94 VPB N_A_27_74#_c_486_n 0.00856377f $X=-0.19 $Y=1.66 $X2=1.98 $Y2=0.815
cc_95 VPB N_A_27_74#_c_500_n 0.0234309f $X=-0.19 $Y=1.66 $X2=1.98 $Y2=0.815
cc_96 VPB N_A_27_74#_c_488_n 0.0215507f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.465
cc_97 VPB N_A_27_74#_c_502_n 0.0105142f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.465
cc_98 VPB N_A_27_74#_c_503_n 0.0413071f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB N_A_27_74#_c_504_n 0.0131772f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 VPB N_A_27_74#_c_493_n 0.00751948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB N_A_987_393#_c_623_n 0.0305113f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.3
cc_102 VPB N_A_987_393#_c_627_n 0.00364593f $X=-0.19 $Y=1.66 $X2=1.47 $Y2=2.55
cc_103 VPB N_A_987_393#_c_632_n 0.00342231f $X=-0.19 $Y=1.66 $X2=1.99 $Y2=2.715
cc_104 VPB N_VPWR_c_688_n 0.00994497f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.97
cc_105 VPB N_VPWR_c_689_n 0.0115779f $X=-0.19 $Y=1.66 $X2=0.785 $Y2=2.055
cc_106 VPB N_VPWR_c_690_n 0.0228511f $X=-0.19 $Y=1.66 $X2=1.47 $Y2=2.55
cc_107 VPB N_VPWR_c_691_n 0.0160896f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_VPWR_c_692_n 0.0280909f $X=-0.19 $Y=1.66 $X2=0.785 $Y2=1.215
cc_109 VPB N_VPWR_c_693_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.465
cc_110 VPB N_VPWR_c_694_n 0.0189953f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.465
cc_111 VPB N_VPWR_c_695_n 0.0541543f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_696_n 0.03837f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_VPWR_c_697_n 0.0208322f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_VPWR_c_687_n 0.120975f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_VPWR_c_699_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_VPWR_c_700_n 0.00615076f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_701_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB GCLK 0.00406323f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_119 VPB N_GCLK_c_776_n 0.0546484f $X=-0.19 $Y=1.66 $X2=1.47 $Y2=2.14
cc_120 N_A_83_260#_c_122_n N_GATE_c_205_n 0.0302036f $X=0.505 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_121 N_A_83_260#_c_123_n N_GATE_c_205_n 9.81638e-19 $X=0.7 $Y=1.63 $X2=-0.19
+ $Y2=-0.245
cc_122 N_A_83_260#_c_124_n N_GATE_c_205_n 0.00446738f $X=0.7 $Y=1.97 $X2=-0.19
+ $Y2=-0.245
cc_123 N_A_83_260#_c_125_n N_GATE_c_205_n 0.0012572f $X=1.385 $Y=1.215 $X2=-0.19
+ $Y2=-0.245
cc_124 N_A_83_260#_c_133_p N_GATE_c_205_n 0.0164359f $X=1.385 $Y=2.055 $X2=-0.19
+ $Y2=-0.245
cc_125 N_A_83_260#_c_134_p N_GATE_c_205_n 0.00612497f $X=1.47 $Y=2.55 $X2=-0.19
+ $Y2=-0.245
cc_126 N_A_83_260#_c_135_p N_GATE_c_205_n 0.0039481f $X=1.555 $Y=2.715 $X2=-0.19
+ $Y2=-0.245
cc_127 N_A_83_260#_M1015_g N_GATE_M1018_g 0.0146085f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_128 N_A_83_260#_c_122_n N_GATE_M1018_g 0.00413511f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_129 N_A_83_260#_c_123_n N_GATE_M1018_g 0.00326474f $X=0.7 $Y=1.63 $X2=0 $Y2=0
cc_130 N_A_83_260#_c_125_n N_GATE_M1018_g 0.0146591f $X=1.385 $Y=1.215 $X2=0
+ $Y2=0
cc_131 N_A_83_260#_c_126_n N_GATE_M1018_g 0.00229553f $X=1.47 $Y=1.13 $X2=0
+ $Y2=0
cc_132 N_A_83_260#_c_123_n GATE 0.0105342f $X=0.7 $Y=1.63 $X2=0 $Y2=0
cc_133 N_A_83_260#_c_124_n GATE 0.0105003f $X=0.7 $Y=1.97 $X2=0 $Y2=0
cc_134 N_A_83_260#_c_125_n GATE 0.0242156f $X=1.385 $Y=1.215 $X2=0 $Y2=0
cc_135 N_A_83_260#_c_133_p GATE 0.0202935f $X=1.385 $Y=2.055 $X2=0 $Y2=0
cc_136 N_A_83_260#_c_125_n N_A_315_54#_c_244_n 0.00202048f $X=1.385 $Y=1.215
+ $X2=0 $Y2=0
cc_137 N_A_83_260#_c_126_n N_A_315_54#_c_244_n 0.00239048f $X=1.47 $Y=1.13 $X2=0
+ $Y2=0
cc_138 N_A_83_260#_c_147_p N_A_315_54#_c_244_n 0.0220414f $X=1.98 $Y=0.815 $X2=0
+ $Y2=0
cc_139 N_A_83_260#_c_148_p N_A_315_54#_c_251_n 0.0151374f $X=1.99 $Y=2.715 $X2=0
+ $Y2=0
cc_140 N_A_83_260#_M1013_d N_A_315_54#_c_247_n 3.0177e-19 $X=1.71 $Y=1.96 $X2=0
+ $Y2=0
cc_141 N_A_83_260#_c_125_n N_A_315_54#_c_247_n 0.0124767f $X=1.385 $Y=1.215
+ $X2=0 $Y2=0
cc_142 N_A_83_260#_c_147_p N_A_315_54#_c_247_n 0.0198287f $X=1.98 $Y=0.815 $X2=0
+ $Y2=0
cc_143 N_A_83_260#_c_147_p N_A_315_54#_c_248_n 0.00184334f $X=1.98 $Y=0.815
+ $X2=0 $Y2=0
cc_144 N_A_83_260#_c_148_p N_A_315_54#_c_254_n 0.0207213f $X=1.99 $Y=2.715 $X2=0
+ $Y2=0
cc_145 N_A_83_260#_M1013_d N_A_315_54#_c_270_n 0.0056801f $X=1.71 $Y=1.96 $X2=0
+ $Y2=0
cc_146 N_A_83_260#_c_148_p N_A_315_54#_c_270_n 0.0194061f $X=1.99 $Y=2.715 $X2=0
+ $Y2=0
cc_147 N_A_83_260#_c_148_p N_A_309_338#_c_367_n 0.0226435f $X=1.99 $Y=2.715
+ $X2=0 $Y2=0
cc_148 N_A_83_260#_c_125_n N_A_309_338#_c_369_n 2.0815e-19 $X=1.385 $Y=1.215
+ $X2=0 $Y2=0
cc_149 N_A_83_260#_c_147_p N_A_309_338#_M1001_g 0.0121375f $X=1.98 $Y=0.815
+ $X2=0 $Y2=0
cc_150 N_A_83_260#_c_147_p N_A_309_338#_c_363_n 0.00324967f $X=1.98 $Y=0.815
+ $X2=0 $Y2=0
cc_151 N_A_83_260#_c_147_p N_A_27_74#_M1014_g 0.00109152f $X=1.98 $Y=0.815 $X2=0
+ $Y2=0
cc_152 N_A_83_260#_c_148_p N_A_27_74#_c_498_n 0.00128241f $X=1.99 $Y=2.715 $X2=0
+ $Y2=0
cc_153 N_A_83_260#_M1015_g N_A_27_74#_c_490_n 0.00835019f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_154 N_A_83_260#_c_122_n N_A_27_74#_c_503_n 0.0132247f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_155 N_A_83_260#_M1015_g N_A_27_74#_c_510_n 0.0110265f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_156 N_A_83_260#_c_122_n N_A_27_74#_c_510_n 6.82831e-19 $X=0.505 $Y=1.765
+ $X2=0 $Y2=0
cc_157 N_A_83_260#_c_123_n N_A_27_74#_c_510_n 0.0198027f $X=0.7 $Y=1.63 $X2=0
+ $Y2=0
cc_158 N_A_83_260#_c_125_n N_A_27_74#_c_510_n 0.030488f $X=1.385 $Y=1.215 $X2=0
+ $Y2=0
cc_159 N_A_83_260#_M1015_g N_A_27_74#_c_514_n 0.00154004f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_160 N_A_83_260#_M1015_g N_A_27_74#_c_492_n 0.00963393f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_161 N_A_83_260#_c_122_n N_A_27_74#_c_492_n 2.30445e-19 $X=0.505 $Y=1.765
+ $X2=0 $Y2=0
cc_162 N_A_83_260#_c_123_n N_A_27_74#_c_492_n 7.22171e-19 $X=0.7 $Y=1.63 $X2=0
+ $Y2=0
cc_163 N_A_83_260#_c_122_n N_A_27_74#_c_504_n 0.00330026f $X=0.505 $Y=1.765
+ $X2=0 $Y2=0
cc_164 N_A_83_260#_c_123_n N_A_27_74#_c_504_n 6.59918e-19 $X=0.7 $Y=1.63 $X2=0
+ $Y2=0
cc_165 N_A_83_260#_c_124_n N_A_27_74#_c_504_n 0.00639412f $X=0.7 $Y=1.97 $X2=0
+ $Y2=0
cc_166 N_A_83_260#_M1015_g N_A_27_74#_c_493_n 0.00256037f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_167 N_A_83_260#_c_122_n N_A_27_74#_c_493_n 0.0107701f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_168 N_A_83_260#_c_123_n N_A_27_74#_c_493_n 0.0311509f $X=0.7 $Y=1.63 $X2=0
+ $Y2=0
cc_169 N_A_83_260#_c_124_n N_A_27_74#_c_493_n 0.00635208f $X=0.7 $Y=1.97 $X2=0
+ $Y2=0
cc_170 N_A_83_260#_M1019_d N_A_27_74#_c_495_n 0.00241797f $X=1.725 $Y=0.4 $X2=0
+ $Y2=0
cc_171 N_A_83_260#_c_180_p N_A_27_74#_c_495_n 0.00750924f $X=1.555 $Y=0.815
+ $X2=0 $Y2=0
cc_172 N_A_83_260#_c_147_p N_A_27_74#_c_495_n 0.0336011f $X=1.98 $Y=0.815 $X2=0
+ $Y2=0
cc_173 N_A_83_260#_c_124_n N_VPWR_M1010_d 0.00278448f $X=0.7 $Y=1.97 $X2=-0.19
+ $Y2=-0.245
cc_174 N_A_83_260#_c_133_p N_VPWR_M1010_d 0.0135858f $X=1.385 $Y=2.055 $X2=-0.19
+ $Y2=-0.245
cc_175 N_A_83_260#_c_184_p N_VPWR_M1010_d 0.00301935f $X=0.785 $Y=2.055
+ $X2=-0.19 $Y2=-0.245
cc_176 N_A_83_260#_c_122_n N_VPWR_c_688_n 0.00909918f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_177 N_A_83_260#_c_133_p N_VPWR_c_688_n 0.0128995f $X=1.385 $Y=2.055 $X2=0
+ $Y2=0
cc_178 N_A_83_260#_c_184_p N_VPWR_c_688_n 0.0132989f $X=0.785 $Y=2.055 $X2=0
+ $Y2=0
cc_179 N_A_83_260#_c_134_p N_VPWR_c_688_n 0.00905739f $X=1.47 $Y=2.55 $X2=0
+ $Y2=0
cc_180 N_A_83_260#_c_135_p N_VPWR_c_688_n 0.0138684f $X=1.555 $Y=2.715 $X2=0
+ $Y2=0
cc_181 N_A_83_260#_c_148_p N_VPWR_c_689_n 0.00451977f $X=1.99 $Y=2.715 $X2=0
+ $Y2=0
cc_182 N_A_83_260#_c_122_n N_VPWR_c_694_n 0.00445602f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_183 N_A_83_260#_c_135_p N_VPWR_c_695_n 0.00447406f $X=1.555 $Y=2.715 $X2=0
+ $Y2=0
cc_184 N_A_83_260#_c_148_p N_VPWR_c_695_n 0.0195114f $X=1.99 $Y=2.715 $X2=0
+ $Y2=0
cc_185 N_A_83_260#_c_122_n N_VPWR_c_687_n 0.00862362f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_186 N_A_83_260#_c_135_p N_VPWR_c_687_n 0.00588029f $X=1.555 $Y=2.715 $X2=0
+ $Y2=0
cc_187 N_A_83_260#_c_148_p N_VPWR_c_687_n 0.023752f $X=1.99 $Y=2.715 $X2=0 $Y2=0
cc_188 N_A_83_260#_c_133_p A_258_392# 0.00480556f $X=1.385 $Y=2.055 $X2=-0.19
+ $Y2=-0.245
cc_189 N_A_83_260#_c_134_p A_258_392# 0.00544755f $X=1.47 $Y=2.55 $X2=-0.19
+ $Y2=-0.245
cc_190 N_A_83_260#_c_135_p A_258_392# 0.00586186f $X=1.555 $Y=2.715 $X2=-0.19
+ $Y2=-0.245
cc_191 N_A_83_260#_M1015_g N_VGND_c_791_n 0.00578197f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_192 N_A_83_260#_c_147_p N_VGND_c_806_n 0.00866412f $X=1.98 $Y=0.815 $X2=0
+ $Y2=0
cc_193 N_A_83_260#_M1015_g N_VGND_c_797_n 0.00434272f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_194 N_A_83_260#_M1015_g N_VGND_c_801_n 0.00443309f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_195 N_A_83_260#_c_180_p A_267_80# 0.00151363f $X=1.555 $Y=0.815 $X2=-0.19
+ $Y2=-0.245
cc_196 N_GATE_M1018_g N_A_315_54#_c_244_n 0.0312233f $X=1.26 $Y=0.72 $X2=0 $Y2=0
cc_197 N_GATE_c_205_n N_A_315_54#_c_247_n 0.00455885f $X=1.215 $Y=1.885 $X2=0
+ $Y2=0
cc_198 N_GATE_M1018_g N_A_315_54#_c_247_n 9.40021e-19 $X=1.26 $Y=0.72 $X2=0
+ $Y2=0
cc_199 GATE N_A_315_54#_c_247_n 0.0133585f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_200 N_GATE_c_205_n N_A_315_54#_c_248_n 0.0312233f $X=1.215 $Y=1.885 $X2=0
+ $Y2=0
cc_201 N_GATE_c_205_n N_A_309_338#_c_367_n 0.0505077f $X=1.215 $Y=1.885 $X2=0
+ $Y2=0
cc_202 N_GATE_c_205_n N_A_309_338#_c_369_n 0.0123452f $X=1.215 $Y=1.885 $X2=0
+ $Y2=0
cc_203 GATE N_A_309_338#_c_369_n 4.953e-19 $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_204 N_GATE_c_205_n N_A_27_74#_c_503_n 8.03191e-19 $X=1.215 $Y=1.885 $X2=0
+ $Y2=0
cc_205 N_GATE_M1018_g N_A_27_74#_c_510_n 0.00554112f $X=1.26 $Y=0.72 $X2=0 $Y2=0
cc_206 N_GATE_M1018_g N_A_27_74#_c_514_n 0.00991337f $X=1.26 $Y=0.72 $X2=0 $Y2=0
cc_207 N_GATE_M1018_g N_A_27_74#_c_491_n 0.00285373f $X=1.26 $Y=0.72 $X2=0 $Y2=0
cc_208 N_GATE_M1018_g N_A_27_74#_c_495_n 0.010234f $X=1.26 $Y=0.72 $X2=0 $Y2=0
cc_209 N_GATE_c_205_n N_VPWR_c_688_n 0.0117996f $X=1.215 $Y=1.885 $X2=0 $Y2=0
cc_210 N_GATE_c_205_n N_VPWR_c_695_n 0.00461464f $X=1.215 $Y=1.885 $X2=0 $Y2=0
cc_211 N_GATE_c_205_n N_VPWR_c_687_n 0.00911469f $X=1.215 $Y=1.885 $X2=0 $Y2=0
cc_212 N_GATE_M1018_g N_VGND_c_791_n 0.0010533f $X=1.26 $Y=0.72 $X2=0 $Y2=0
cc_213 N_GATE_M1018_g N_VGND_c_795_n 9.48944e-19 $X=1.26 $Y=0.72 $X2=0 $Y2=0
cc_214 N_A_315_54#_c_256_n N_A_309_338#_M1016_d 0.0081007f $X=3.945 $Y=2.475
+ $X2=0 $Y2=0
cc_215 N_A_315_54#_c_251_n N_A_309_338#_c_367_n 0.0227084f $X=2.345 $Y=2.465
+ $X2=0 $Y2=0
cc_216 N_A_315_54#_c_247_n N_A_309_338#_c_367_n 0.00497441f $X=1.83 $Y=1.315
+ $X2=0 $Y2=0
cc_217 N_A_315_54#_c_251_n N_A_309_338#_c_368_n 0.0214699f $X=2.345 $Y=2.465
+ $X2=0 $Y2=0
cc_218 N_A_315_54#_c_247_n N_A_309_338#_c_368_n 0.0168228f $X=1.83 $Y=1.315
+ $X2=0 $Y2=0
cc_219 N_A_315_54#_c_254_n N_A_309_338#_c_368_n 0.00542654f $X=3.03 $Y=2.215
+ $X2=0 $Y2=0
cc_220 N_A_315_54#_c_247_n N_A_309_338#_c_369_n 0.00200055f $X=1.83 $Y=1.315
+ $X2=0 $Y2=0
cc_221 N_A_315_54#_c_248_n N_A_309_338#_c_369_n 0.0298557f $X=1.83 $Y=1.315
+ $X2=0 $Y2=0
cc_222 N_A_315_54#_c_244_n N_A_309_338#_M1001_g 0.0150689f $X=1.65 $Y=1.15 $X2=0
+ $Y2=0
cc_223 N_A_315_54#_c_247_n N_A_309_338#_M1001_g 6.52036e-19 $X=1.83 $Y=1.315
+ $X2=0 $Y2=0
cc_224 N_A_315_54#_c_248_n N_A_309_338#_M1001_g 0.0177805f $X=1.83 $Y=1.315
+ $X2=0 $Y2=0
cc_225 N_A_315_54#_c_251_n N_A_309_338#_c_360_n 9.88384e-19 $X=2.345 $Y=2.465
+ $X2=0 $Y2=0
cc_226 N_A_315_54#_c_247_n N_A_309_338#_c_360_n 0.0334095f $X=1.83 $Y=1.315
+ $X2=0 $Y2=0
cc_227 N_A_315_54#_c_248_n N_A_309_338#_c_360_n 9.37391e-19 $X=1.83 $Y=1.315
+ $X2=0 $Y2=0
cc_228 N_A_315_54#_c_254_n N_A_309_338#_c_360_n 0.0223796f $X=3.03 $Y=2.215
+ $X2=0 $Y2=0
cc_229 N_A_315_54#_c_255_n N_A_309_338#_c_360_n 3.35121e-19 $X=3.115 $Y=2.05
+ $X2=0 $Y2=0
cc_230 N_A_315_54#_c_250_n N_A_309_338#_c_360_n 0.0118744f $X=3.27 $Y=1.665
+ $X2=0 $Y2=0
cc_231 N_A_315_54#_c_247_n N_A_309_338#_c_361_n 0.00398033f $X=1.83 $Y=1.315
+ $X2=0 $Y2=0
cc_232 N_A_315_54#_c_254_n N_A_309_338#_c_361_n 8.18206e-19 $X=3.03 $Y=2.215
+ $X2=0 $Y2=0
cc_233 N_A_315_54#_c_245_n N_A_309_338#_c_362_n 0.00346492f $X=3.31 $Y=1.915
+ $X2=0 $Y2=0
cc_234 N_A_315_54#_M1003_g N_A_309_338#_c_362_n 0.0122329f $X=3.335 $Y=0.995
+ $X2=0 $Y2=0
cc_235 N_A_315_54#_c_250_n N_A_309_338#_c_362_n 0.0268373f $X=3.27 $Y=1.665
+ $X2=0 $Y2=0
cc_236 N_A_315_54#_c_247_n N_A_309_338#_c_363_n 0.0120735f $X=1.83 $Y=1.315
+ $X2=0 $Y2=0
cc_237 N_A_315_54#_c_248_n N_A_309_338#_c_363_n 0.00116112f $X=1.83 $Y=1.315
+ $X2=0 $Y2=0
cc_238 N_A_315_54#_M1003_g N_A_309_338#_c_364_n 5.39498e-19 $X=3.335 $Y=0.995
+ $X2=0 $Y2=0
cc_239 N_A_315_54#_c_249_n N_A_309_338#_c_364_n 0.00850585f $X=4.115 $Y=1.22
+ $X2=0 $Y2=0
cc_240 N_A_315_54#_c_245_n N_A_309_338#_c_365_n 0.00590021f $X=3.31 $Y=1.915
+ $X2=0 $Y2=0
cc_241 N_A_315_54#_M1003_g N_A_309_338#_c_365_n 0.00513868f $X=3.335 $Y=0.995
+ $X2=0 $Y2=0
cc_242 N_A_315_54#_c_255_n N_A_309_338#_c_365_n 0.00771087f $X=3.115 $Y=2.05
+ $X2=0 $Y2=0
cc_243 N_A_315_54#_c_249_n N_A_309_338#_c_365_n 0.0560684f $X=4.115 $Y=1.22
+ $X2=0 $Y2=0
cc_244 N_A_315_54#_c_250_n N_A_309_338#_c_365_n 0.0251647f $X=3.27 $Y=1.665
+ $X2=0 $Y2=0
cc_245 N_A_315_54#_c_245_n N_A_309_338#_c_373_n 0.00201359f $X=3.31 $Y=1.915
+ $X2=0 $Y2=0
cc_246 N_A_315_54#_c_256_n N_A_309_338#_c_373_n 0.0253855f $X=3.945 $Y=2.475
+ $X2=0 $Y2=0
cc_247 N_A_315_54#_c_258_n N_A_309_338#_c_373_n 0.0141831f $X=4.102 $Y=2.102
+ $X2=0 $Y2=0
cc_248 N_A_315_54#_c_250_n N_A_309_338#_c_373_n 0.00237071f $X=3.27 $Y=1.665
+ $X2=0 $Y2=0
cc_249 N_A_315_54#_c_249_n N_A_309_338#_c_366_n 0.0147863f $X=4.115 $Y=1.22
+ $X2=0 $Y2=0
cc_250 N_A_315_54#_c_256_n N_CLK_c_440_n 0.00659227f $X=3.945 $Y=2.475 $X2=-0.19
+ $Y2=-0.245
cc_251 N_A_315_54#_c_249_n N_CLK_c_440_n 0.00224171f $X=4.115 $Y=1.22 $X2=-0.19
+ $Y2=-0.245
cc_252 N_A_315_54#_c_258_n N_CLK_c_440_n 0.0028454f $X=4.102 $Y=2.102 $X2=-0.19
+ $Y2=-0.245
cc_253 N_A_315_54#_c_259_n N_CLK_c_440_n 0.00443109f $X=4.095 $Y=2.11 $X2=-0.19
+ $Y2=-0.245
cc_254 N_A_315_54#_c_249_n N_CLK_c_436_n 0.00445076f $X=4.115 $Y=1.22 $X2=0
+ $Y2=0
cc_255 N_A_315_54#_c_249_n CLK 0.0209126f $X=4.115 $Y=1.22 $X2=0 $Y2=0
cc_256 N_A_315_54#_c_249_n N_CLK_c_439_n 0.015011f $X=4.115 $Y=1.22 $X2=0 $Y2=0
cc_257 N_A_315_54#_c_258_n N_CLK_c_439_n 7.74196e-19 $X=4.102 $Y=2.102 $X2=0
+ $Y2=0
cc_258 N_A_315_54#_M1003_g N_A_27_74#_M1014_g 0.0131462f $X=3.335 $Y=0.995 $X2=0
+ $Y2=0
cc_259 N_A_315_54#_c_245_n N_A_27_74#_c_497_n 0.00612277f $X=3.31 $Y=1.915 $X2=0
+ $Y2=0
cc_260 N_A_315_54#_c_254_n N_A_27_74#_c_497_n 0.00559679f $X=3.03 $Y=2.215 $X2=0
+ $Y2=0
cc_261 N_A_315_54#_c_251_n N_A_27_74#_c_498_n 0.0338785f $X=2.345 $Y=2.465 $X2=0
+ $Y2=0
cc_262 N_A_315_54#_c_245_n N_A_27_74#_c_498_n 0.00906853f $X=3.31 $Y=1.915 $X2=0
+ $Y2=0
cc_263 N_A_315_54#_c_254_n N_A_27_74#_c_498_n 0.00783014f $X=3.03 $Y=2.215 $X2=0
+ $Y2=0
cc_264 N_A_315_54#_c_327_p N_A_27_74#_c_498_n 0.00501994f $X=3.115 $Y=2.305
+ $X2=0 $Y2=0
cc_265 N_A_315_54#_M1003_g N_A_27_74#_c_484_n 0.00889043f $X=3.335 $Y=0.995
+ $X2=0 $Y2=0
cc_266 N_A_315_54#_M1003_g N_A_27_74#_c_487_n 0.0138204f $X=3.335 $Y=0.995 $X2=0
+ $Y2=0
cc_267 N_A_315_54#_c_251_n N_A_27_74#_c_488_n 0.00134234f $X=2.345 $Y=2.465
+ $X2=0 $Y2=0
cc_268 N_A_315_54#_c_245_n N_A_27_74#_c_488_n 0.0309611f $X=3.31 $Y=1.915 $X2=0
+ $Y2=0
cc_269 N_A_315_54#_c_254_n N_A_27_74#_c_488_n 0.00821606f $X=3.03 $Y=2.215 $X2=0
+ $Y2=0
cc_270 N_A_315_54#_c_255_n N_A_27_74#_c_488_n 0.0047439f $X=3.115 $Y=2.05 $X2=0
+ $Y2=0
cc_271 N_A_315_54#_c_250_n N_A_27_74#_c_488_n 0.00331054f $X=3.27 $Y=1.665 $X2=0
+ $Y2=0
cc_272 N_A_315_54#_c_251_n N_A_27_74#_c_502_n 0.0193573f $X=2.345 $Y=2.465 $X2=0
+ $Y2=0
cc_273 N_A_315_54#_c_254_n N_A_27_74#_c_502_n 0.00793908f $X=3.03 $Y=2.215 $X2=0
+ $Y2=0
cc_274 N_A_315_54#_c_244_n N_A_27_74#_c_514_n 0.00124375f $X=1.65 $Y=1.15 $X2=0
+ $Y2=0
cc_275 N_A_315_54#_c_244_n N_A_27_74#_c_495_n 0.0119481f $X=1.65 $Y=1.15 $X2=0
+ $Y2=0
cc_276 N_A_315_54#_M1003_g N_A_27_74#_c_496_n 6.13725e-19 $X=3.335 $Y=0.995
+ $X2=0 $Y2=0
cc_277 N_A_315_54#_c_254_n N_VPWR_M1005_d 0.0033399f $X=3.03 $Y=2.215 $X2=0
+ $Y2=0
cc_278 N_A_315_54#_c_255_n N_VPWR_M1005_d 8.97844e-19 $X=3.115 $Y=2.05 $X2=0
+ $Y2=0
cc_279 N_A_315_54#_c_327_p N_VPWR_M1005_d 0.00530672f $X=3.115 $Y=2.305 $X2=0
+ $Y2=0
cc_280 N_A_315_54#_c_251_n N_VPWR_c_689_n 0.00143234f $X=2.345 $Y=2.465 $X2=0
+ $Y2=0
cc_281 N_A_315_54#_c_245_n N_VPWR_c_689_n 0.00644269f $X=3.31 $Y=1.915 $X2=0
+ $Y2=0
cc_282 N_A_315_54#_c_254_n N_VPWR_c_689_n 0.00828406f $X=3.03 $Y=2.215 $X2=0
+ $Y2=0
cc_283 N_A_315_54#_c_327_p N_VPWR_c_689_n 0.0116666f $X=3.115 $Y=2.305 $X2=0
+ $Y2=0
cc_284 N_A_315_54#_c_256_n N_VPWR_c_690_n 0.0178843f $X=3.945 $Y=2.475 $X2=0
+ $Y2=0
cc_285 N_A_315_54#_c_251_n N_VPWR_c_695_n 0.00445785f $X=2.345 $Y=2.465 $X2=0
+ $Y2=0
cc_286 N_A_315_54#_c_245_n N_VPWR_c_696_n 0.00487664f $X=3.31 $Y=1.915 $X2=0
+ $Y2=0
cc_287 N_A_315_54#_c_256_n N_VPWR_c_696_n 0.00854871f $X=3.945 $Y=2.475 $X2=0
+ $Y2=0
cc_288 N_A_315_54#_c_251_n N_VPWR_c_687_n 0.00892591f $X=2.345 $Y=2.465 $X2=0
+ $Y2=0
cc_289 N_A_315_54#_c_245_n N_VPWR_c_687_n 0.00505379f $X=3.31 $Y=1.915 $X2=0
+ $Y2=0
cc_290 N_A_315_54#_c_256_n N_VPWR_c_687_n 0.0373199f $X=3.945 $Y=2.475 $X2=0
+ $Y2=0
cc_291 N_A_315_54#_c_327_p N_VPWR_c_687_n 0.00202923f $X=3.115 $Y=2.305 $X2=0
+ $Y2=0
cc_292 N_A_315_54#_M1003_g N_VGND_c_806_n 0.00774033f $X=3.335 $Y=0.995 $X2=0
+ $Y2=0
cc_293 N_A_315_54#_M1003_g N_VGND_c_792_n 0.00779576f $X=3.335 $Y=0.995 $X2=0
+ $Y2=0
cc_294 N_A_315_54#_c_244_n N_VGND_c_795_n 9.29978e-19 $X=1.65 $Y=1.15 $X2=0
+ $Y2=0
cc_295 N_A_315_54#_M1003_g N_VGND_c_801_n 7.34656e-19 $X=3.335 $Y=0.995 $X2=0
+ $Y2=0
cc_296 N_A_309_338#_c_364_n N_CLK_c_436_n 0.00722606f $X=3.55 $Y=0.77 $X2=0
+ $Y2=0
cc_297 N_A_309_338#_c_364_n N_A_27_74#_c_484_n 0.0061136f $X=3.55 $Y=0.77 $X2=0
+ $Y2=0
cc_298 N_A_309_338#_c_362_n N_A_27_74#_c_487_n 0.0119084f $X=3.465 $Y=1.245
+ $X2=0 $Y2=0
cc_299 N_A_309_338#_M1001_g N_A_27_74#_c_488_n 0.0072772f $X=2.31 $Y=0.83 $X2=0
+ $Y2=0
cc_300 N_A_309_338#_c_360_n N_A_27_74#_c_488_n 0.00526915f $X=2.37 $Y=1.675
+ $X2=0 $Y2=0
cc_301 N_A_309_338#_c_361_n N_A_27_74#_c_488_n 0.02065f $X=2.37 $Y=1.675 $X2=0
+ $Y2=0
cc_302 N_A_309_338#_c_362_n N_A_27_74#_c_488_n 0.00932416f $X=3.465 $Y=1.245
+ $X2=0 $Y2=0
cc_303 N_A_309_338#_c_362_n N_A_27_74#_c_494_n 0.00285995f $X=3.465 $Y=1.245
+ $X2=0 $Y2=0
cc_304 N_A_309_338#_M1001_g N_A_27_74#_c_495_n 0.00658236f $X=2.31 $Y=0.83 $X2=0
+ $Y2=0
cc_305 N_A_309_338#_M1001_g N_A_27_74#_c_496_n 0.0418981f $X=2.31 $Y=0.83 $X2=0
+ $Y2=0
cc_306 N_A_309_338#_c_367_n N_VPWR_c_695_n 0.00304676f $X=1.635 $Y=1.885 $X2=0
+ $Y2=0
cc_307 N_A_309_338#_c_367_n N_VPWR_c_687_n 0.00375764f $X=1.635 $Y=1.885 $X2=0
+ $Y2=0
cc_308 N_A_309_338#_c_362_n N_VGND_M1014_d 0.00469367f $X=3.465 $Y=1.245 $X2=0
+ $Y2=0
cc_309 N_A_309_338#_M1001_g N_VGND_c_806_n 7.00177e-19 $X=2.31 $Y=0.83 $X2=0
+ $Y2=0
cc_310 N_A_309_338#_c_362_n N_VGND_c_806_n 0.0279461f $X=3.465 $Y=1.245 $X2=0
+ $Y2=0
cc_311 N_A_309_338#_c_364_n N_VGND_c_792_n 0.00346039f $X=3.55 $Y=0.77 $X2=0
+ $Y2=0
cc_312 N_A_309_338#_c_364_n N_VGND_c_793_n 0.0134733f $X=3.55 $Y=0.77 $X2=0
+ $Y2=0
cc_313 N_A_309_338#_c_364_n N_VGND_c_798_n 0.00663535f $X=3.55 $Y=0.77 $X2=0
+ $Y2=0
cc_314 N_A_309_338#_c_364_n N_VGND_c_801_n 0.00833855f $X=3.55 $Y=0.77 $X2=0
+ $Y2=0
cc_315 N_CLK_c_436_n N_A_27_74#_c_484_n 0.00894529f $X=4.335 $Y=1.475 $X2=0
+ $Y2=0
cc_316 N_CLK_M1011_g N_A_27_74#_c_484_n 0.00907339f $X=4.845 $Y=0.945 $X2=0
+ $Y2=0
cc_317 N_CLK_M1011_g N_A_27_74#_M1008_g 0.0253528f $X=4.845 $Y=0.945 $X2=0 $Y2=0
cc_318 CLK N_A_27_74#_c_486_n 0.00281307f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_319 N_CLK_c_439_n N_A_27_74#_c_486_n 0.0159521f $X=4.845 $Y=1.682 $X2=0 $Y2=0
cc_320 N_CLK_c_441_n N_A_27_74#_c_500_n 0.0135311f $X=4.86 $Y=1.89 $X2=0 $Y2=0
cc_321 N_CLK_c_439_n N_A_27_74#_c_489_n 0.0253528f $X=4.845 $Y=1.682 $X2=0 $Y2=0
cc_322 N_CLK_M1011_g N_A_987_393#_c_626_n 0.00151317f $X=4.845 $Y=0.945 $X2=0
+ $Y2=0
cc_323 N_CLK_c_441_n N_A_987_393#_c_627_n 3.88984e-19 $X=4.86 $Y=1.89 $X2=0
+ $Y2=0
cc_324 CLK N_A_987_393#_c_627_n 0.0119738f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_325 N_CLK_c_439_n N_A_987_393#_c_627_n 6.16305e-19 $X=4.845 $Y=1.682 $X2=0
+ $Y2=0
cc_326 N_CLK_c_441_n N_A_987_393#_c_632_n 0.00795337f $X=4.86 $Y=1.89 $X2=0
+ $Y2=0
cc_327 N_CLK_c_441_n N_A_987_393#_c_638_n 0.00150219f $X=4.86 $Y=1.89 $X2=0
+ $Y2=0
cc_328 CLK N_A_987_393#_c_638_n 0.0153408f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_329 N_CLK_M1011_g N_A_987_393#_c_629_n 0.0010598f $X=4.845 $Y=0.945 $X2=0
+ $Y2=0
cc_330 CLK N_A_987_393#_c_629_n 0.0116912f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_331 N_CLK_c_440_n N_VPWR_c_690_n 0.0082344f $X=4.32 $Y=1.89 $X2=0 $Y2=0
cc_332 N_CLK_c_441_n N_VPWR_c_690_n 0.00421592f $X=4.86 $Y=1.89 $X2=0 $Y2=0
cc_333 CLK N_VPWR_c_690_n 0.0242246f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_334 N_CLK_c_439_n N_VPWR_c_690_n 0.00900791f $X=4.845 $Y=1.682 $X2=0 $Y2=0
cc_335 N_CLK_c_441_n N_VPWR_c_692_n 0.0046892f $X=4.86 $Y=1.89 $X2=0 $Y2=0
cc_336 N_CLK_c_440_n N_VPWR_c_696_n 0.00460155f $X=4.32 $Y=1.89 $X2=0 $Y2=0
cc_337 N_CLK_c_440_n N_VPWR_c_687_n 0.0049796f $X=4.32 $Y=1.89 $X2=0 $Y2=0
cc_338 N_CLK_c_441_n N_VPWR_c_687_n 0.0049796f $X=4.86 $Y=1.89 $X2=0 $Y2=0
cc_339 N_CLK_c_436_n N_VGND_c_793_n 0.0200137f $X=4.335 $Y=1.475 $X2=0 $Y2=0
cc_340 N_CLK_M1011_g N_VGND_c_793_n 0.00730266f $X=4.845 $Y=0.945 $X2=0 $Y2=0
cc_341 CLK N_VGND_c_793_n 0.0212606f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_342 N_CLK_c_439_n N_VGND_c_793_n 0.00436753f $X=4.845 $Y=1.682 $X2=0 $Y2=0
cc_343 N_CLK_c_436_n N_VGND_c_801_n 7.97988e-19 $X=4.335 $Y=1.475 $X2=0 $Y2=0
cc_344 N_CLK_M1011_g N_VGND_c_801_n 9.49986e-19 $X=4.845 $Y=0.945 $X2=0 $Y2=0
cc_345 N_A_27_74#_c_486_n N_A_987_393#_c_623_n 0.00314054f $X=5.32 $Y=1.8 $X2=0
+ $Y2=0
cc_346 N_A_27_74#_c_500_n N_A_987_393#_c_623_n 0.00988243f $X=5.32 $Y=1.89 $X2=0
+ $Y2=0
cc_347 N_A_27_74#_M1008_g N_A_987_393#_c_625_n 9.88035e-19 $X=5.235 $Y=0.945
+ $X2=0 $Y2=0
cc_348 N_A_27_74#_c_489_n N_A_987_393#_c_625_n 0.012306f $X=5.285 $Y=1.49 $X2=0
+ $Y2=0
cc_349 N_A_27_74#_M1008_g N_A_987_393#_c_626_n 0.0100958f $X=5.235 $Y=0.945
+ $X2=0 $Y2=0
cc_350 N_A_27_74#_c_486_n N_A_987_393#_c_627_n 0.00438577f $X=5.32 $Y=1.8 $X2=0
+ $Y2=0
cc_351 N_A_27_74#_c_500_n N_A_987_393#_c_627_n 0.00580919f $X=5.32 $Y=1.89 $X2=0
+ $Y2=0
cc_352 N_A_27_74#_c_500_n N_A_987_393#_c_632_n 0.0136103f $X=5.32 $Y=1.89 $X2=0
+ $Y2=0
cc_353 N_A_27_74#_c_500_n N_A_987_393#_c_638_n 0.0159564f $X=5.32 $Y=1.89 $X2=0
+ $Y2=0
cc_354 N_A_27_74#_c_489_n N_A_987_393#_c_638_n 0.001564f $X=5.285 $Y=1.49 $X2=0
+ $Y2=0
cc_355 N_A_27_74#_M1008_g N_A_987_393#_c_629_n 0.00624269f $X=5.235 $Y=0.945
+ $X2=0 $Y2=0
cc_356 N_A_27_74#_c_486_n N_A_987_393#_c_629_n 0.003544f $X=5.32 $Y=1.8 $X2=0
+ $Y2=0
cc_357 N_A_27_74#_c_489_n N_A_987_393#_c_629_n 0.00927392f $X=5.285 $Y=1.49
+ $X2=0 $Y2=0
cc_358 N_A_27_74#_c_503_n N_VPWR_c_688_n 0.0261579f $X=0.28 $Y=2.815 $X2=0 $Y2=0
cc_359 N_A_27_74#_c_498_n N_VPWR_c_689_n 0.00861583f $X=2.765 $Y=2.465 $X2=0
+ $Y2=0
cc_360 N_A_27_74#_c_500_n N_VPWR_c_691_n 0.0100062f $X=5.32 $Y=1.89 $X2=0 $Y2=0
cc_361 N_A_27_74#_c_500_n N_VPWR_c_692_n 0.00460952f $X=5.32 $Y=1.89 $X2=0 $Y2=0
cc_362 N_A_27_74#_c_503_n N_VPWR_c_694_n 0.0154862f $X=0.28 $Y=2.815 $X2=0 $Y2=0
cc_363 N_A_27_74#_c_498_n N_VPWR_c_695_n 0.00444681f $X=2.765 $Y=2.465 $X2=0
+ $Y2=0
cc_364 N_A_27_74#_c_498_n N_VPWR_c_687_n 0.00911827f $X=2.765 $Y=2.465 $X2=0
+ $Y2=0
cc_365 N_A_27_74#_c_500_n N_VPWR_c_687_n 0.0049796f $X=5.32 $Y=1.89 $X2=0 $Y2=0
cc_366 N_A_27_74#_c_503_n N_VPWR_c_687_n 0.0127853f $X=0.28 $Y=2.815 $X2=0 $Y2=0
cc_367 N_A_27_74#_c_510_n N_VGND_M1015_d 0.0132019f $X=1.045 $Y=0.875 $X2=-0.19
+ $Y2=-0.245
cc_368 N_A_27_74#_c_514_n N_VGND_M1015_d 0.00441864f $X=1.13 $Y=0.79 $X2=-0.19
+ $Y2=-0.245
cc_369 N_A_27_74#_c_491_n N_VGND_M1015_d 2.44449e-19 $X=1.215 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_370 N_A_27_74#_c_490_n N_VGND_c_791_n 0.0104927f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_371 N_A_27_74#_c_510_n N_VGND_c_791_n 0.0196232f $X=1.045 $Y=0.875 $X2=0
+ $Y2=0
cc_372 N_A_27_74#_c_514_n N_VGND_c_791_n 0.0145482f $X=1.13 $Y=0.79 $X2=0 $Y2=0
cc_373 N_A_27_74#_c_491_n N_VGND_c_791_n 0.0145354f $X=1.215 $Y=0.34 $X2=0 $Y2=0
cc_374 N_A_27_74#_M1014_g N_VGND_c_806_n 0.00917897f $X=2.7 $Y=0.83 $X2=0 $Y2=0
cc_375 N_A_27_74#_c_484_n N_VGND_c_806_n 0.00138507f $X=5.16 $Y=0.18 $X2=0 $Y2=0
cc_376 N_A_27_74#_c_487_n N_VGND_c_806_n 0.00126939f $X=2.82 $Y=1.19 $X2=0 $Y2=0
cc_377 N_A_27_74#_c_494_n N_VGND_c_806_n 0.0122171f $X=2.79 $Y=0.345 $X2=0 $Y2=0
cc_378 N_A_27_74#_c_496_n N_VGND_c_806_n 0.00251883f $X=2.79 $Y=0.18 $X2=0 $Y2=0
cc_379 N_A_27_74#_M1014_g N_VGND_c_792_n 0.00316397f $X=2.7 $Y=0.83 $X2=0 $Y2=0
cc_380 N_A_27_74#_c_484_n N_VGND_c_792_n 0.0163869f $X=5.16 $Y=0.18 $X2=0 $Y2=0
cc_381 N_A_27_74#_c_494_n N_VGND_c_792_n 0.0198501f $X=2.79 $Y=0.345 $X2=0 $Y2=0
cc_382 N_A_27_74#_c_496_n N_VGND_c_792_n 0.00172991f $X=2.79 $Y=0.18 $X2=0 $Y2=0
cc_383 N_A_27_74#_c_484_n N_VGND_c_793_n 0.0257165f $X=5.16 $Y=0.18 $X2=0 $Y2=0
cc_384 N_A_27_74#_M1008_g N_VGND_c_793_n 0.00806567f $X=5.235 $Y=0.945 $X2=0
+ $Y2=0
cc_385 N_A_27_74#_c_484_n N_VGND_c_794_n 0.0111053f $X=5.16 $Y=0.18 $X2=0 $Y2=0
cc_386 N_A_27_74#_M1008_g N_VGND_c_794_n 8.98699e-19 $X=5.235 $Y=0.945 $X2=0
+ $Y2=0
cc_387 N_A_27_74#_c_491_n N_VGND_c_795_n 0.0122203f $X=1.215 $Y=0.34 $X2=0 $Y2=0
cc_388 N_A_27_74#_c_495_n N_VGND_c_795_n 0.111626f $X=2.625 $Y=0.382 $X2=0 $Y2=0
cc_389 N_A_27_74#_c_496_n N_VGND_c_795_n 0.0121847f $X=2.79 $Y=0.18 $X2=0 $Y2=0
cc_390 N_A_27_74#_c_490_n N_VGND_c_797_n 0.0154563f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_391 N_A_27_74#_c_484_n N_VGND_c_798_n 0.0350534f $X=5.16 $Y=0.18 $X2=0 $Y2=0
cc_392 N_A_27_74#_c_484_n N_VGND_c_799_n 0.0215943f $X=5.16 $Y=0.18 $X2=0 $Y2=0
cc_393 N_A_27_74#_c_484_n N_VGND_c_801_n 0.0817763f $X=5.16 $Y=0.18 $X2=0 $Y2=0
cc_394 N_A_27_74#_c_490_n N_VGND_c_801_n 0.012737f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_395 N_A_27_74#_c_510_n N_VGND_c_801_n 0.0126469f $X=1.045 $Y=0.875 $X2=0
+ $Y2=0
cc_396 N_A_27_74#_c_491_n N_VGND_c_801_n 0.00661553f $X=1.215 $Y=0.34 $X2=0
+ $Y2=0
cc_397 N_A_27_74#_c_495_n N_VGND_c_801_n 0.0640172f $X=2.625 $Y=0.382 $X2=0
+ $Y2=0
cc_398 N_A_27_74#_c_496_n N_VGND_c_801_n 0.0102842f $X=2.79 $Y=0.18 $X2=0 $Y2=0
cc_399 N_A_27_74#_c_495_n A_267_80# 0.00151475f $X=2.625 $Y=0.382 $X2=-0.19
+ $Y2=-0.245
cc_400 N_A_987_393#_c_627_n N_VPWR_M1007_d 3.38187e-19 $X=5.45 $Y=1.975 $X2=0
+ $Y2=0
cc_401 N_A_987_393#_c_638_n N_VPWR_M1007_d 0.00503912f $X=5.45 $Y=2.06 $X2=0
+ $Y2=0
cc_402 N_A_987_393#_c_632_n N_VPWR_c_690_n 0.0263057f $X=5.095 $Y=2.14 $X2=0
+ $Y2=0
cc_403 N_A_987_393#_c_623_n N_VPWR_c_691_n 0.0145077f $X=6.145 $Y=1.765 $X2=0
+ $Y2=0
cc_404 N_A_987_393#_c_625_n N_VPWR_c_691_n 0.00693494f $X=6.055 $Y=1.465 $X2=0
+ $Y2=0
cc_405 N_A_987_393#_c_627_n N_VPWR_c_691_n 0.0023498f $X=5.45 $Y=1.975 $X2=0
+ $Y2=0
cc_406 N_A_987_393#_c_628_n N_VPWR_c_691_n 0.0163051f $X=5.87 $Y=1.465 $X2=0
+ $Y2=0
cc_407 N_A_987_393#_c_632_n N_VPWR_c_691_n 0.0251369f $X=5.095 $Y=2.14 $X2=0
+ $Y2=0
cc_408 N_A_987_393#_c_638_n N_VPWR_c_691_n 0.0141779f $X=5.45 $Y=2.06 $X2=0
+ $Y2=0
cc_409 N_A_987_393#_c_632_n N_VPWR_c_692_n 0.00890943f $X=5.095 $Y=2.14 $X2=0
+ $Y2=0
cc_410 N_A_987_393#_c_623_n N_VPWR_c_697_n 0.00445602f $X=6.145 $Y=1.765 $X2=0
+ $Y2=0
cc_411 N_A_987_393#_c_623_n N_VPWR_c_687_n 0.00865423f $X=6.145 $Y=1.765 $X2=0
+ $Y2=0
cc_412 N_A_987_393#_c_632_n N_VPWR_c_687_n 0.0109157f $X=5.095 $Y=2.14 $X2=0
+ $Y2=0
cc_413 N_A_987_393#_c_623_n N_GCLK_c_773_n 0.00953446f $X=6.145 $Y=1.765 $X2=0
+ $Y2=0
cc_414 N_A_987_393#_M1012_g N_GCLK_c_773_n 0.0179032f $X=6.225 $Y=0.74 $X2=0
+ $Y2=0
cc_415 N_A_987_393#_c_628_n N_GCLK_c_773_n 0.0154371f $X=5.87 $Y=1.465 $X2=0
+ $Y2=0
cc_416 N_A_987_393#_c_629_n N_GCLK_c_773_n 0.00478285f $X=5.285 $Y=1.12 $X2=0
+ $Y2=0
cc_417 N_A_987_393#_c_623_n GCLK 0.0119702f $X=6.145 $Y=1.765 $X2=0 $Y2=0
cc_418 N_A_987_393#_c_627_n GCLK 0.00836825f $X=5.45 $Y=1.975 $X2=0 $Y2=0
cc_419 N_A_987_393#_c_628_n GCLK 0.00638763f $X=5.87 $Y=1.465 $X2=0 $Y2=0
cc_420 N_A_987_393#_c_623_n N_GCLK_c_776_n 0.018353f $X=6.145 $Y=1.765 $X2=0
+ $Y2=0
cc_421 N_A_987_393#_c_626_n N_VGND_c_793_n 0.0074529f $X=5.45 $Y=0.77 $X2=0
+ $Y2=0
cc_422 N_A_987_393#_c_629_n N_VGND_c_793_n 0.00326799f $X=5.285 $Y=1.12 $X2=0
+ $Y2=0
cc_423 N_A_987_393#_M1012_g N_VGND_c_794_n 0.00647412f $X=6.225 $Y=0.74 $X2=0
+ $Y2=0
cc_424 N_A_987_393#_c_625_n N_VGND_c_794_n 0.00712404f $X=6.055 $Y=1.465 $X2=0
+ $Y2=0
cc_425 N_A_987_393#_c_626_n N_VGND_c_794_n 0.0339721f $X=5.45 $Y=0.77 $X2=0
+ $Y2=0
cc_426 N_A_987_393#_c_628_n N_VGND_c_794_n 0.015939f $X=5.87 $Y=1.465 $X2=0
+ $Y2=0
cc_427 N_A_987_393#_c_629_n N_VGND_c_794_n 6.6261e-19 $X=5.285 $Y=1.12 $X2=0
+ $Y2=0
cc_428 N_A_987_393#_c_626_n N_VGND_c_799_n 0.00702137f $X=5.45 $Y=0.77 $X2=0
+ $Y2=0
cc_429 N_A_987_393#_M1012_g N_VGND_c_800_n 0.00434272f $X=6.225 $Y=0.74 $X2=0
+ $Y2=0
cc_430 N_A_987_393#_M1012_g N_VGND_c_801_n 0.00828941f $X=6.225 $Y=0.74 $X2=0
+ $Y2=0
cc_431 N_A_987_393#_c_626_n N_VGND_c_801_n 0.0100521f $X=5.45 $Y=0.77 $X2=0
+ $Y2=0
cc_432 N_VPWR_c_691_n N_GCLK_c_776_n 0.0407863f $X=5.87 $Y=2.11 $X2=0 $Y2=0
cc_433 N_VPWR_c_697_n N_GCLK_c_776_n 0.0177173f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_434 N_VPWR_c_687_n N_GCLK_c_776_n 0.0146319f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_435 N_GCLK_c_773_n N_VGND_c_794_n 0.0294122f $X=6.44 $Y=0.515 $X2=0 $Y2=0
cc_436 N_GCLK_c_773_n N_VGND_c_800_n 0.0145639f $X=6.44 $Y=0.515 $X2=0 $Y2=0
cc_437 N_GCLK_c_773_n N_VGND_c_801_n 0.0119984f $X=6.44 $Y=0.515 $X2=0 $Y2=0
