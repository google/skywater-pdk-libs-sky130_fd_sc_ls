* File: sky130_fd_sc_ls__mux2_4.pex.spice
* Created: Fri Aug 28 13:30:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__MUX2_4%S 1 3 6 10 12 14 17 19 21 23 24 25 26 29 30
+ 32 35 39 43 47
c138 47 0 1.32825e-20 $X=3.97 $Y=1.657
c139 32 0 1.42621e-19 $X=3.58 $Y=1.6
r140 47 48 1.85385 $w=3.9e-07 $l=1.5e-08 $layer=POLY_cond $X=3.97 $Y=1.657
+ $X2=3.985 $Y2=1.657
r141 44 45 8.03333 $w=3.9e-07 $l=6.5e-08 $layer=POLY_cond $X=3.47 $Y=1.657
+ $X2=3.535 $Y2=1.657
r142 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.59
+ $Y=1.515 $X2=0.59 $Y2=1.515
r143 39 53 7.28531 $w=4.08e-07 $l=1.15e-07 $layer=LI1_cond $X=0.63 $Y=1.665
+ $X2=0.63 $Y2=1.78
r144 39 43 4.21625 $w=4.08e-07 $l=1.5e-07 $layer=LI1_cond $X=0.63 $Y=1.665
+ $X2=0.63 $Y2=1.515
r145 35 37 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=1.59 $Y=2.135
+ $X2=1.59 $Y2=2.24
r146 33 47 48.2 $w=3.9e-07 $l=3.9e-07 $layer=POLY_cond $X=3.58 $Y=1.657 $X2=3.97
+ $Y2=1.657
r147 33 45 5.56154 $w=3.9e-07 $l=4.5e-08 $layer=POLY_cond $X=3.58 $Y=1.657
+ $X2=3.535 $Y2=1.657
r148 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.58
+ $Y=1.6 $X2=3.58 $Y2=1.6
r149 30 32 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=3.165 $Y=1.6
+ $X2=3.58 $Y2=1.6
r150 28 30 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.08 $Y=1.765
+ $X2=3.165 $Y2=1.6
r151 28 29 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=3.08 $Y=1.765
+ $X2=3.08 $Y2=2.155
r152 27 37 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.675 $Y=2.24
+ $X2=1.59 $Y2=2.24
r153 26 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.995 $Y=2.24
+ $X2=3.08 $Y2=2.155
r154 26 27 86.1176 $w=1.68e-07 $l=1.32e-06 $layer=LI1_cond $X=2.995 $Y=2.24
+ $X2=1.675 $Y2=2.24
r155 24 35 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.505 $Y=2.135
+ $X2=1.59 $Y2=2.135
r156 24 25 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.505 $Y=2.135
+ $X2=0.835 $Y2=2.135
r157 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.75 $Y=2.05
+ $X2=0.835 $Y2=2.135
r158 23 53 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.75 $Y=2.05
+ $X2=0.75 $Y2=1.78
r159 19 48 25.2441 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=3.985 $Y=1.88
+ $X2=3.985 $Y2=1.657
r160 19 21 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.985 $Y=1.88
+ $X2=3.985 $Y2=2.455
r161 15 47 25.2441 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=3.97 $Y=1.435
+ $X2=3.97 $Y2=1.657
r162 15 17 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=3.97 $Y=1.435
+ $X2=3.97 $Y2=0.915
r163 12 45 25.2441 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=3.535 $Y=1.88
+ $X2=3.535 $Y2=1.657
r164 12 14 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.535 $Y=1.88
+ $X2=3.535 $Y2=2.455
r165 8 44 25.2441 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=3.47 $Y=1.435
+ $X2=3.47 $Y2=1.657
r166 8 10 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=3.47 $Y=1.435
+ $X2=3.47 $Y2=0.915
r167 4 42 38.5336 $w=3.07e-07 $l=1.94808e-07 $layer=POLY_cond $X=0.65 $Y=1.35
+ $X2=0.585 $Y2=1.515
r168 4 6 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=0.65 $Y=1.35 $X2=0.65
+ $Y2=0.81
r169 1 42 51.8789 $w=3.07e-07 $l=2.87228e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.585 $Y2=1.515
r170 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_LS__MUX2_4%A_27_368# 1 2 7 9 12 16 18 20 24 25 26 27 30
+ 31 32 34 35 37 41 45 46 47 54
c137 54 0 1.42621e-19 $X=5.04 $Y=1.657
c138 45 0 1.47598e-19 $X=0.28 $Y=2.115
c139 27 0 5.64602e-20 $X=3.335 $Y=2.58
r140 54 55 1.90765 $w=3.79e-07 $l=1.5e-08 $layer=POLY_cond $X=5.04 $Y=1.657
+ $X2=5.055 $Y2=1.657
r141 51 52 0.635884 $w=3.79e-07 $l=5e-09 $layer=POLY_cond $X=4.605 $Y=1.657
+ $X2=4.61 $Y2=1.657
r142 47 49 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=1.25 $Y=2.475
+ $X2=1.25 $Y2=2.58
r143 45 46 8.51103 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=0.265 $Y=2.115
+ $X2=0.265 $Y2=1.95
r144 43 46 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=0.17 $Y=1.15 $X2=0.17
+ $Y2=1.95
r145 41 43 17.7387 $w=5.13e-07 $l=5.15e-07 $layer=LI1_cond $X=0.342 $Y=0.635
+ $X2=0.342 $Y2=1.15
r146 38 54 27.9789 $w=3.79e-07 $l=2.2e-07 $layer=POLY_cond $X=4.82 $Y=1.657
+ $X2=5.04 $Y2=1.657
r147 38 52 26.7071 $w=3.79e-07 $l=2.1e-07 $layer=POLY_cond $X=4.82 $Y=1.657
+ $X2=4.61 $Y2=1.657
r148 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.82
+ $Y=1.6 $X2=4.82 $Y2=1.6
r149 35 37 25.668 $w=3.28e-07 $l=7.35e-07 $layer=LI1_cond $X=4.085 $Y=1.6
+ $X2=4.82 $Y2=1.6
r150 33 35 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=4 $Y=1.765
+ $X2=4.085 $Y2=1.6
r151 33 34 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4 $Y=1.765 $X2=4
+ $Y2=1.935
r152 31 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.915 $Y=2.02
+ $X2=4 $Y2=1.935
r153 31 32 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=3.915 $Y=2.02
+ $X2=3.505 $Y2=2.02
r154 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.42 $Y=2.105
+ $X2=3.505 $Y2=2.02
r155 29 30 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=3.42 $Y=2.105
+ $X2=3.42 $Y2=2.495
r156 28 49 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.335 $Y=2.58
+ $X2=1.25 $Y2=2.58
r157 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.335 $Y=2.58
+ $X2=3.42 $Y2=2.495
r158 27 28 130.481 $w=1.68e-07 $l=2e-06 $layer=LI1_cond $X=3.335 $Y=2.58
+ $X2=1.335 $Y2=2.58
r159 25 47 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.165 $Y=2.475
+ $X2=1.25 $Y2=2.475
r160 25 26 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=1.165 $Y=2.475
+ $X2=0.445 $Y2=2.475
r161 24 26 8.02311 $w=1.7e-07 $l=2.18403e-07 $layer=LI1_cond $X=0.265 $Y=2.39
+ $X2=0.445 $Y2=2.475
r162 23 45 0.480185 $w=3.58e-07 $l=1.5e-08 $layer=LI1_cond $X=0.265 $Y=2.13
+ $X2=0.265 $Y2=2.115
r163 23 24 8.3232 $w=3.58e-07 $l=2.6e-07 $layer=LI1_cond $X=0.265 $Y=2.13
+ $X2=0.265 $Y2=2.39
r164 18 55 24.5487 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=5.055 $Y=1.88
+ $X2=5.055 $Y2=1.657
r165 18 20 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.055 $Y=1.88
+ $X2=5.055 $Y2=2.455
r166 14 54 24.5487 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=5.04 $Y=1.435
+ $X2=5.04 $Y2=1.657
r167 14 16 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=5.04 $Y=1.435
+ $X2=5.04 $Y2=0.915
r168 10 52 24.5487 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=4.61 $Y=1.435
+ $X2=4.61 $Y2=1.657
r169 10 12 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=4.61 $Y=1.435
+ $X2=4.61 $Y2=0.915
r170 7 51 24.5487 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=4.605 $Y=1.88
+ $X2=4.605 $Y2=1.657
r171 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=4.605 $Y=1.88
+ $X2=4.605 $Y2=2.455
r172 2 45 300 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.115
r173 1 41 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.29
+ $Y=0.49 $X2=0.435 $Y2=0.635
.ends

.subckt PM_SKY130_FD_SC_LS__MUX2_4%A_193_241# 1 2 3 4 5 6 20 21 23 27 28 29 30
+ 31 32 34 38 39 44 45 46 47 49 50 55 56 58 59 60 62 64 67 70 71 73 78 85 89 90
+ 91 96 100 102 107 110 113 115 116 117 118 120 121
c231 45 0 5.9954e-20 $X=2.295 $Y=1.295
c232 21 0 1.47598e-19 $X=1.055 $Y=1.765
c233 20 0 1.62123e-19 $X=1.055 $Y=1.675
r234 121 126 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=5.78 $Y=1.615
+ $X2=5.705 $Y2=1.615
r235 115 116 8.4794 $w=3.43e-07 $l=1.65e-07 $layer=LI1_cond $X=6.425 $Y=0.427
+ $X2=6.59 $Y2=0.427
r236 113 120 5.16603 $w=2.5e-07 $l=1.60078e-07 $layer=LI1_cond $X=8.44 $Y=1.95
+ $X2=8.36 $Y2=2.075
r237 113 118 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=8.44 $Y=1.95
+ $X2=8.44 $Y2=1.03
r238 108 120 5.16603 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=8.36 $Y=2.2
+ $X2=8.36 $Y2=2.075
r239 108 110 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=8.36 $Y=2.2
+ $X2=8.36 $Y2=2.465
r240 105 118 8.53494 $w=3.33e-07 $l=1.67e-07 $layer=LI1_cond $X=8.357 $Y=0.863
+ $X2=8.357 $Y2=1.03
r241 105 107 11.9716 $w=3.33e-07 $l=3.48e-07 $layer=LI1_cond $X=8.357 $Y=0.863
+ $X2=8.357 $Y2=0.515
r242 104 107 3.09612 $w=3.33e-07 $l=9e-08 $layer=LI1_cond $X=8.357 $Y=0.425
+ $X2=8.357 $Y2=0.515
r243 103 117 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.59 $Y=0.34
+ $X2=7.425 $Y2=0.34
r244 102 104 7.80856 $w=1.7e-07 $l=2.05144e-07 $layer=LI1_cond $X=8.19 $Y=0.34
+ $X2=8.357 $Y2=0.425
r245 102 103 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=8.19 $Y=0.34
+ $X2=7.59 $Y2=0.34
r246 98 117 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.425 $Y=0.425
+ $X2=7.425 $Y2=0.34
r247 98 100 2.44458 $w=3.28e-07 $l=7e-08 $layer=LI1_cond $X=7.425 $Y=0.425
+ $X2=7.425 $Y2=0.495
r248 96 117 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.26 $Y=0.34
+ $X2=7.425 $Y2=0.34
r249 96 116 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.26 $Y=0.34
+ $X2=6.59 $Y2=0.34
r250 93 95 42.6404 $w=2.48e-07 $l=9.25e-07 $layer=LI1_cond $X=6.48 $Y=2.075
+ $X2=7.405 $Y2=2.075
r251 91 93 0.460977 $w=2.48e-07 $l=1e-08 $layer=LI1_cond $X=6.47 $Y=2.075
+ $X2=6.48 $Y2=2.075
r252 90 120 1.34256 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=8.195 $Y=2.075
+ $X2=8.36 $Y2=2.075
r253 90 95 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=8.195 $Y=2.075
+ $X2=7.405 $Y2=2.075
r254 89 91 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.385 $Y=1.95
+ $X2=6.47 $Y2=2.075
r255 88 89 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=6.385 $Y=1.78
+ $X2=6.385 $Y2=1.95
r256 85 121 78.6876 $w=3.3e-07 $l=4.5e-07 $layer=POLY_cond $X=6.23 $Y=1.615
+ $X2=5.78 $Y2=1.615
r257 84 85 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=6.23
+ $Y=1.615 $X2=6.23 $Y2=1.615
r258 81 126 27.1035 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=5.55 $Y=1.615
+ $X2=5.705 $Y2=1.615
r259 80 84 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=5.55 $Y=1.615
+ $X2=6.23 $Y2=1.615
r260 80 81 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=5.55
+ $Y=1.615 $X2=5.55 $Y2=1.615
r261 78 88 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.3 $Y=1.615
+ $X2=6.385 $Y2=1.78
r262 78 84 2.44458 $w=3.28e-07 $l=7e-08 $layer=LI1_cond $X=6.3 $Y=1.615 $X2=6.23
+ $Y2=1.615
r263 64 126 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.705 $Y=1.45
+ $X2=5.705 $Y2=1.615
r264 63 64 612.755 $w=1.5e-07 $l=1.195e-06 $layer=POLY_cond $X=5.705 $Y=0.255
+ $X2=5.705 $Y2=1.45
r265 60 62 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.915 $Y=1.765
+ $X2=2.915 $Y2=2.4
r266 59 60 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.915 $Y=1.675
+ $X2=2.915 $Y2=1.765
r267 58 74 105.117 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=2.915 $Y=1.385
+ $X2=2.71 $Y2=1.385
r268 58 59 83.5726 $w=1.8e-07 $l=2.15e-07 $layer=POLY_cond $X=2.915 $Y=1.46
+ $X2=2.915 $Y2=1.675
r269 57 73 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.785 $Y=0.18
+ $X2=2.71 $Y2=0.18
r270 56 63 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.63 $Y=0.18
+ $X2=5.705 $Y2=0.255
r271 56 57 1458.82 $w=1.5e-07 $l=2.845e-06 $layer=POLY_cond $X=5.63 $Y=0.18
+ $X2=2.785 $Y2=0.18
r272 53 74 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.71 $Y=1.31
+ $X2=2.71 $Y2=1.385
r273 53 55 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.71 $Y=1.31
+ $X2=2.71 $Y2=0.76
r274 52 73 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.71 $Y=0.255
+ $X2=2.71 $Y2=0.18
r275 52 55 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=2.71 $Y=0.255
+ $X2=2.71 $Y2=0.76
r276 51 71 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.355 $Y=0.18
+ $X2=2.28 $Y2=0.18
r277 50 73 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.635 $Y=0.18
+ $X2=2.71 $Y2=0.18
r278 50 51 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.635 $Y=0.18
+ $X2=2.355 $Y2=0.18
r279 47 49 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.295 $Y=1.765
+ $X2=2.295 $Y2=2.4
r280 46 47 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.295 $Y=1.675
+ $X2=2.295 $Y2=1.765
r281 45 72 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.295 $Y=1.295
+ $X2=2.295 $Y2=1.205
r282 45 46 147.71 $w=1.8e-07 $l=3.8e-07 $layer=POLY_cond $X=2.295 $Y=1.295
+ $X2=2.295 $Y2=1.675
r283 44 72 228.181 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.28 $Y=0.76
+ $X2=2.28 $Y2=1.205
r284 41 71 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.28 $Y=0.255
+ $X2=2.28 $Y2=0.18
r285 41 44 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=2.28 $Y=0.255
+ $X2=2.28 $Y2=0.76
r286 40 70 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.765 $Y=0.18
+ $X2=1.69 $Y2=0.18
r287 39 71 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.205 $Y=0.18
+ $X2=2.28 $Y2=0.18
r288 39 40 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=2.205 $Y=0.18
+ $X2=1.765 $Y2=0.18
r289 38 69 228.181 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.69 $Y=0.76
+ $X2=1.69 $Y2=1.205
r290 35 70 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.69 $Y=0.255
+ $X2=1.69 $Y2=0.18
r291 35 38 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=1.69 $Y=0.255
+ $X2=1.69 $Y2=0.76
r292 32 34 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.675 $Y=1.765
+ $X2=1.675 $Y2=2.4
r293 31 32 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.675 $Y=1.675
+ $X2=1.675 $Y2=1.765
r294 30 69 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.675 $Y=1.295
+ $X2=1.675 $Y2=1.205
r295 30 31 147.71 $w=1.8e-07 $l=3.8e-07 $layer=POLY_cond $X=1.675 $Y=1.295
+ $X2=1.675 $Y2=1.675
r296 28 70 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.615 $Y=0.18
+ $X2=1.69 $Y2=0.18
r297 28 29 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.615 $Y=0.18
+ $X2=1.295 $Y2=0.18
r298 25 67 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.22 $Y=1.205
+ $X2=1.22 $Y2=1.28
r299 25 27 228.181 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.22 $Y=1.205
+ $X2=1.22 $Y2=0.76
r300 24 29 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.22 $Y=0.255
+ $X2=1.295 $Y2=0.18
r301 24 27 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=1.22 $Y=0.255
+ $X2=1.22 $Y2=0.76
r302 21 23 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.055 $Y=1.765
+ $X2=1.055 $Y2=2.4
r303 20 21 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.055 $Y=1.675
+ $X2=1.055 $Y2=1.765
r304 19 67 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.055 $Y=1.28
+ $X2=1.22 $Y2=1.28
r305 19 20 124.387 $w=1.8e-07 $l=3.2e-07 $layer=POLY_cond $X=1.055 $Y=1.355
+ $X2=1.055 $Y2=1.675
r306 6 120 600 $w=1.7e-07 $l=2.66458e-07 $layer=licon1_PDIFF $count=1 $X=8.16
+ $Y=1.96 $X2=8.36 $Y2=2.115
r307 6 110 300 $w=1.7e-07 $l=5.96678e-07 $layer=licon1_PDIFF $count=2 $X=8.16
+ $Y=1.96 $X2=8.36 $Y2=2.465
r308 5 95 600 $w=1.7e-07 $l=2.19203e-07 $layer=licon1_PDIFF $count=1 $X=7.25
+ $Y=1.96 $X2=7.405 $Y2=2.115
r309 4 93 600 $w=1.7e-07 $l=2.24499e-07 $layer=licon1_PDIFF $count=1 $X=6.32
+ $Y=1.96 $X2=6.48 $Y2=2.115
r310 3 107 91 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_NDIFF $count=2 $X=8.175
+ $Y=0.37 $X2=8.355 $Y2=0.515
r311 2 100 91 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_NDIFF $count=2 $X=7.235
+ $Y=0.37 $X2=7.425 $Y2=0.495
r312 1 115 91 $w=1.7e-07 $l=6.38396e-07 $layer=licon1_NDIFF $count=2 $X=5.855
+ $Y=0.37 $X2=6.425 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__MUX2_4%A0 3 5 7 10 12 14 15 22
r45 22 23 1.89267 $w=3.82e-07 $l=1.5e-08 $layer=POLY_cond $X=7.16 $Y=1.667
+ $X2=7.175 $Y2=1.667
r46 20 22 44.7932 $w=3.82e-07 $l=3.55e-07 $layer=POLY_cond $X=6.805 $Y=1.667
+ $X2=7.16 $Y2=1.667
r47 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.805
+ $Y=1.615 $X2=6.805 $Y2=1.615
r48 18 20 10.0942 $w=3.82e-07 $l=8e-08 $layer=POLY_cond $X=6.725 $Y=1.667
+ $X2=6.805 $Y2=1.667
r49 17 18 1.89267 $w=3.82e-07 $l=1.5e-08 $layer=POLY_cond $X=6.71 $Y=1.667
+ $X2=6.725 $Y2=1.667
r50 15 21 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=6.96 $Y=1.615
+ $X2=6.805 $Y2=1.615
r51 12 23 24.74 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=7.175 $Y=1.885
+ $X2=7.175 $Y2=1.667
r52 12 14 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=7.175 $Y=1.885
+ $X2=7.175 $Y2=2.46
r53 8 22 24.74 $w=1.5e-07 $l=2.17e-07 $layer=POLY_cond $X=7.16 $Y=1.45 $X2=7.16
+ $Y2=1.667
r54 8 10 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=7.16 $Y=1.45 $X2=7.16
+ $Y2=0.69
r55 5 18 24.74 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=6.725 $Y=1.885
+ $X2=6.725 $Y2=1.667
r56 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.725 $Y=1.885
+ $X2=6.725 $Y2=2.46
r57 1 17 24.74 $w=1.5e-07 $l=2.17e-07 $layer=POLY_cond $X=6.71 $Y=1.45 $X2=6.71
+ $Y2=1.667
r58 1 3 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=6.71 $Y=1.45 $X2=6.71
+ $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_LS__MUX2_4%A1 1 3 6 8 10 13 15 16 23 24
r47 24 25 1.87306 $w=3.86e-07 $l=1.5e-08 $layer=POLY_cond $X=8.085 $Y=1.667
+ $X2=8.1 $Y2=1.667
r48 22 24 9.36528 $w=3.86e-07 $l=7.5e-08 $layer=POLY_cond $X=8.01 $Y=1.667
+ $X2=8.085 $Y2=1.667
r49 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.01
+ $Y=1.615 $X2=8.01 $Y2=1.615
r50 20 22 46.2021 $w=3.86e-07 $l=3.7e-07 $layer=POLY_cond $X=7.64 $Y=1.667
+ $X2=8.01 $Y2=1.667
r51 19 20 0.624352 $w=3.86e-07 $l=5e-09 $layer=POLY_cond $X=7.635 $Y=1.667
+ $X2=7.64 $Y2=1.667
r52 16 23 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=7.92 $Y=1.615 $X2=8.01
+ $Y2=1.615
r53 15 16 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=7.44 $Y=1.615
+ $X2=7.92 $Y2=1.615
r54 11 25 24.9932 $w=1.5e-07 $l=2.17e-07 $layer=POLY_cond $X=8.1 $Y=1.45 $X2=8.1
+ $Y2=1.667
r55 11 13 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=8.1 $Y=1.45 $X2=8.1
+ $Y2=0.69
r56 8 24 24.9932 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=8.085 $Y=1.885
+ $X2=8.085 $Y2=1.667
r57 8 10 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=8.085 $Y=1.885
+ $X2=8.085 $Y2=2.46
r58 4 20 24.9932 $w=1.5e-07 $l=2.17e-07 $layer=POLY_cond $X=7.64 $Y=1.45
+ $X2=7.64 $Y2=1.667
r59 4 6 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=7.64 $Y=1.45 $X2=7.64
+ $Y2=0.69
r60 1 19 24.9932 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=7.635 $Y=1.885
+ $X2=7.635 $Y2=1.667
r61 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=7.635 $Y=1.885
+ $X2=7.635 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_LS__MUX2_4%VPWR 1 2 3 4 5 20 24 28 32 36 39 40 42 43 45
+ 46 47 53 68 69 72 75
r101 75 76 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r102 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r103 68 69 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r104 66 69 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=8.4 $Y2=3.33
r105 65 68 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=5.52 $Y=3.33
+ $X2=8.4 $Y2=3.33
r106 65 66 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r107 63 66 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r108 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r109 60 76 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.12 $Y2=3.33
r110 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r111 57 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.39 $Y=3.33
+ $X2=3.225 $Y2=3.33
r112 57 59 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.39 $Y=3.33
+ $X2=4.08 $Y2=3.33
r113 56 76 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r114 55 56 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r115 53 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.06 $Y=3.33
+ $X2=3.225 $Y2=3.33
r116 53 55 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=3.06 $Y=3.33 $X2=2.16
+ $Y2=3.33
r117 52 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r118 52 73 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r119 51 52 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r120 49 72 8.88104 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.995 $Y=3.33
+ $X2=0.822 $Y2=3.33
r121 49 51 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=0.995 $Y=3.33
+ $X2=1.68 $Y2=3.33
r122 47 63 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=4.32 $Y=3.33
+ $X2=5.04 $Y2=3.33
r123 47 60 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=3.33
+ $X2=4.08 $Y2=3.33
r124 45 62 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=5.2 $Y=3.33
+ $X2=5.04 $Y2=3.33
r125 45 46 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.2 $Y=3.33
+ $X2=5.325 $Y2=3.33
r126 44 65 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=5.45 $Y=3.33 $X2=5.52
+ $Y2=3.33
r127 44 46 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.45 $Y=3.33
+ $X2=5.325 $Y2=3.33
r128 42 59 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=4.13 $Y=3.33 $X2=4.08
+ $Y2=3.33
r129 42 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.13 $Y=3.33
+ $X2=4.295 $Y2=3.33
r130 41 62 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=4.46 $Y=3.33
+ $X2=5.04 $Y2=3.33
r131 41 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.46 $Y=3.33
+ $X2=4.295 $Y2=3.33
r132 39 51 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=1.82 $Y=3.33
+ $X2=1.68 $Y2=3.33
r133 39 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.82 $Y=3.33
+ $X2=1.985 $Y2=3.33
r134 38 55 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=2.15 $Y=3.33
+ $X2=2.16 $Y2=3.33
r135 38 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.15 $Y=3.33
+ $X2=1.985 $Y2=3.33
r136 34 46 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.325 $Y=3.245
+ $X2=5.325 $Y2=3.33
r137 34 36 14.0598 $w=2.48e-07 $l=3.05e-07 $layer=LI1_cond $X=5.325 $Y=3.245
+ $X2=5.325 $Y2=2.94
r138 30 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.295 $Y=3.245
+ $X2=4.295 $Y2=3.33
r139 30 32 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=4.295 $Y=3.245
+ $X2=4.295 $Y2=2.94
r140 26 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.225 $Y=3.245
+ $X2=3.225 $Y2=3.33
r141 26 28 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=3.225 $Y=3.245
+ $X2=3.225 $Y2=3
r142 22 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.985 $Y=3.245
+ $X2=1.985 $Y2=3.33
r143 22 24 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=1.985 $Y=3.245
+ $X2=1.985 $Y2=3
r144 18 72 1.03204 $w=3.45e-07 $l=8.5e-08 $layer=LI1_cond $X=0.822 $Y=3.245
+ $X2=0.822 $Y2=3.33
r145 18 20 14.3638 $w=3.43e-07 $l=4.3e-07 $layer=LI1_cond $X=0.822 $Y=3.245
+ $X2=0.822 $Y2=2.815
r146 5 36 600 $w=1.7e-07 $l=1.09622e-06 $layer=licon1_PDIFF $count=1 $X=5.13
+ $Y=1.955 $X2=5.365 $Y2=2.94
r147 4 32 600 $w=1.7e-07 $l=1.09622e-06 $layer=licon1_PDIFF $count=1 $X=4.06
+ $Y=1.955 $X2=4.295 $Y2=2.94
r148 3 28 600 $w=1.7e-07 $l=1.27208e-06 $layer=licon1_PDIFF $count=1 $X=2.99
+ $Y=1.84 $X2=3.225 $Y2=3
r149 2 24 600 $w=1.7e-07 $l=1.27208e-06 $layer=licon1_PDIFF $count=1 $X=1.75
+ $Y=1.84 $X2=1.985 $Y2=3
r150 1 20 600 $w=1.7e-07 $l=1.0884e-06 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.84 $X2=0.82 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_LS__MUX2_4%X 1 2 3 4 13 15 17 19 21 23 24 30 33
c64 30 0 2.54869e-20 $X=2.33 $Y=1.625
c65 17 0 1.32825e-20 $X=2.542 $Y=1.37
c66 15 0 1.62123e-19 $X=1.475 $Y=0.535
c67 13 0 3.09733e-20 $X=1.475 $Y=1.37
r68 31 33 0.938101 $w=5.08e-07 $l=4e-08 $layer=LI1_cond $X=1.64 $Y=1.625
+ $X2=1.68 $Y2=1.625
r69 24 30 3.19265 $w=5.1e-07 $l=2.44622e-07 $layer=LI1_cond $X=2.55 $Y=1.677
+ $X2=2.33 $Y2=1.625
r70 23 30 3.98693 $w=5.08e-07 $l=1.7e-07 $layer=LI1_cond $X=2.16 $Y=1.625
+ $X2=2.33 $Y2=1.625
r71 21 31 3.11208 $w=5.1e-07 $l=2.78e-07 $layer=LI1_cond $X=1.362 $Y=1.625
+ $X2=1.64 $Y2=1.625
r72 21 23 10.7413 $w=5.08e-07 $l=4.58e-07 $layer=LI1_cond $X=1.702 $Y=1.625
+ $X2=2.16 $Y2=1.625
r73 21 33 0.515955 $w=5.08e-07 $l=2.2e-08 $layer=LI1_cond $X=1.702 $Y=1.625
+ $X2=1.68 $Y2=1.625
r74 17 24 3.69737 $w=4.25e-07 $l=3.10974e-07 $layer=LI1_cond $X=2.542 $Y=1.37
+ $X2=2.55 $Y2=1.677
r75 17 19 22.6421 $w=4.23e-07 $l=8.35e-07 $layer=LI1_cond $X=2.542 $Y=1.37
+ $X2=2.542 $Y2=0.535
r76 13 21 4.11959 $w=3.3e-07 $l=3.06333e-07 $layer=LI1_cond $X=1.475 $Y=1.37
+ $X2=1.362 $Y2=1.625
r77 13 15 29.1603 $w=3.28e-07 $l=8.35e-07 $layer=LI1_cond $X=1.475 $Y=1.37
+ $X2=1.475 $Y2=0.535
r78 4 24 600 $w=1.7e-07 $l=2.63296e-07 $layer=licon1_PDIFF $count=1 $X=2.37
+ $Y=1.84 $X2=2.605 $Y2=1.9
r79 3 21 600 $w=1.7e-07 $l=2.56515e-07 $layer=licon1_PDIFF $count=1 $X=1.13
+ $Y=1.84 $X2=1.365 $Y2=1.795
r80 2 19 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.355
+ $Y=0.39 $X2=2.495 $Y2=0.535
r81 1 15 91 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_NDIFF $count=2 $X=1.295
+ $Y=0.39 $X2=1.475 $Y2=0.535
.ends

.subckt PM_SKY130_FD_SC_LS__MUX2_4%A_722_391# 1 2 9 13 16 17
r49 11 17 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=5.705 $Y=2.845
+ $X2=5.705 $Y2=2.52
r50 11 13 49.5124 $w=2.68e-07 $l=1.16e-06 $layer=LI1_cond $X=5.79 $Y=2.845
+ $X2=6.95 $Y2=2.845
r51 10 16 3.9577 $w=1.7e-07 $l=1.60078e-07 $layer=LI1_cond $X=3.925 $Y=2.52
+ $X2=3.8 $Y2=2.44
r52 9 17 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.62 $Y=2.52
+ $X2=5.705 $Y2=2.52
r53 9 10 110.583 $w=1.68e-07 $l=1.695e-06 $layer=LI1_cond $X=5.62 $Y=2.52
+ $X2=3.925 $Y2=2.52
r54 2 13 600 $w=1.7e-07 $l=9.16938e-07 $layer=licon1_PDIFF $count=1 $X=6.8
+ $Y=1.96 $X2=6.95 $Y2=2.805
r55 1 16 300 $w=1.7e-07 $l=5.54955e-07 $layer=licon1_PDIFF $count=2 $X=3.61
+ $Y=1.955 $X2=3.76 $Y2=2.44
.ends

.subckt PM_SKY130_FD_SC_LS__MUX2_4%A_936_391# 1 2 7 9 16 17 22
r46 17 19 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.045 $Y=2.18
+ $X2=6.045 $Y2=2.455
r47 14 16 13.5259 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=4.83 $Y=2.1 $X2=5.14
+ $Y2=2.1
r48 10 19 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.13 $Y=2.455
+ $X2=6.045 $Y2=2.455
r49 9 22 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.695 $Y=2.455
+ $X2=7.86 $Y2=2.455
r50 9 10 102.102 $w=1.68e-07 $l=1.565e-06 $layer=LI1_cond $X=7.695 $Y=2.455
+ $X2=6.13 $Y2=2.455
r51 7 17 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.96 $Y=2.18
+ $X2=6.045 $Y2=2.18
r52 7 16 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=5.96 $Y=2.18 $X2=5.14
+ $Y2=2.18
r53 2 22 300 $w=1.7e-07 $l=5.65044e-07 $layer=licon1_PDIFF $count=2 $X=7.71
+ $Y=1.96 $X2=7.86 $Y2=2.455
r54 1 14 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=4.68
+ $Y=1.955 $X2=4.83 $Y2=2.1
.ends

.subckt PM_SKY130_FD_SC_LS__MUX2_4%VGND 1 2 3 4 5 18 22 26 30 34 38 41 42 44 45
+ 46 55 59 66 67 70 73 76
c106 26 0 5.9954e-20 $X=3.09 $Y=0.535
r107 76 77 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r108 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r109 71 74 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r110 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r111 67 77 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=8.4 $Y=0 $X2=5.52
+ $Y2=0
r112 66 67 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=8.4 $Y=0
+ $X2=8.4 $Y2=0
r113 64 76 9.89127 $w=1.7e-07 $l=2.03e-07 $layer=LI1_cond $X=5.575 $Y=0
+ $X2=5.372 $Y2=0
r114 64 66 184.305 $w=1.68e-07 $l=2.825e-06 $layer=LI1_cond $X=5.575 $Y=0
+ $X2=8.4 $Y2=0
r115 63 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r116 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r117 60 73 10.873 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=4.49 $Y=0 $X2=4.255
+ $Y2=0
r118 60 62 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=4.49 $Y=0 $X2=5.04
+ $Y2=0
r119 59 76 9.89127 $w=1.7e-07 $l=2.02e-07 $layer=LI1_cond $X=5.17 $Y=0 $X2=5.372
+ $Y2=0
r120 59 62 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=5.17 $Y=0 $X2=5.04
+ $Y2=0
r121 58 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r122 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r123 55 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.925 $Y=0 $X2=3.09
+ $Y2=0
r124 55 57 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.925 $Y=0
+ $X2=2.64 $Y2=0
r125 54 58 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r126 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r127 50 54 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r128 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r129 46 63 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=4.32 $Y=0 $X2=5.04
+ $Y2=0
r130 46 74 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=0
+ $X2=4.08 $Y2=0
r131 44 53 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=1.81 $Y=0 $X2=1.68
+ $Y2=0
r132 44 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.81 $Y=0 $X2=1.975
+ $Y2=0
r133 43 57 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=2.14 $Y=0 $X2=2.64
+ $Y2=0
r134 43 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.14 $Y=0 $X2=1.975
+ $Y2=0
r135 41 49 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=0.77 $Y=0 $X2=0.72
+ $Y2=0
r136 41 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.77 $Y=0 $X2=0.935
+ $Y2=0
r137 40 53 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=1.1 $Y=0 $X2=1.68
+ $Y2=0
r138 40 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.1 $Y=0 $X2=0.935
+ $Y2=0
r139 36 76 1.50354 $w=4.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.372 $Y=0.085
+ $X2=5.372 $Y2=0
r140 36 38 11.809 $w=4.03e-07 $l=4.15e-07 $layer=LI1_cond $X=5.372 $Y=0.085
+ $X2=5.372 $Y2=0.5
r141 32 73 1.91284 $w=4.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.255 $Y=0.085
+ $X2=4.255 $Y2=0
r142 32 34 16.6688 $w=4.68e-07 $l=6.55e-07 $layer=LI1_cond $X=4.255 $Y=0.085
+ $X2=4.255 $Y2=0.74
r143 31 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.255 $Y=0 $X2=3.09
+ $Y2=0
r144 30 73 10.873 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=4.02 $Y=0 $X2=4.255
+ $Y2=0
r145 30 31 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=4.02 $Y=0
+ $X2=3.255 $Y2=0
r146 26 28 19.382 $w=3.28e-07 $l=5.55e-07 $layer=LI1_cond $X=3.09 $Y=0.535
+ $X2=3.09 $Y2=1.09
r147 24 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.09 $Y=0.085
+ $X2=3.09 $Y2=0
r148 24 26 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=3.09 $Y=0.085
+ $X2=3.09 $Y2=0.535
r149 20 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.975 $Y=0.085
+ $X2=1.975 $Y2=0
r150 20 22 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=1.975 $Y=0.085
+ $X2=1.975 $Y2=0.535
r151 16 42 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.935 $Y=0.085
+ $X2=0.935 $Y2=0
r152 16 18 19.2074 $w=3.28e-07 $l=5.5e-07 $layer=LI1_cond $X=0.935 $Y=0.085
+ $X2=0.935 $Y2=0.635
r153 5 38 182 $w=1.7e-07 $l=2.98747e-07 $layer=licon1_NDIFF $count=1 $X=5.115
+ $Y=0.595 $X2=5.37 $Y2=0.5
r154 4 34 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=4.045
+ $Y=0.595 $X2=4.255 $Y2=0.74
r155 3 28 182 $w=1.7e-07 $l=8.38749e-07 $layer=licon1_NDIFF $count=1 $X=2.785
+ $Y=0.39 $X2=3.09 $Y2=1.09
r156 3 26 182 $w=1.7e-07 $l=3.70473e-07 $layer=licon1_NDIFF $count=1 $X=2.785
+ $Y=0.39 $X2=3.09 $Y2=0.535
r157 2 22 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=1.765
+ $Y=0.39 $X2=1.975 $Y2=0.535
r158 1 18 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=0.725
+ $Y=0.49 $X2=0.935 $Y2=0.635
.ends

.subckt PM_SKY130_FD_SC_LS__MUX2_4%A_709_119# 1 2 9 12 13 17 19 20
r60 19 20 10.1916 $w=1.83e-07 $l=1.7e-07 $layer=LI1_cond $X=5.155 $Y=1.187
+ $X2=5.325 $Y2=1.187
r61 15 17 13.8293 $w=2.48e-07 $l=3e-07 $layer=LI1_cond $X=7.895 $Y=1.11
+ $X2=7.895 $Y2=0.81
r62 13 15 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=7.77 $Y=1.195
+ $X2=7.895 $Y2=1.11
r63 13 20 159.513 $w=1.68e-07 $l=2.445e-06 $layer=LI1_cond $X=7.77 $Y=1.195
+ $X2=5.325 $Y2=1.195
r64 12 19 85.139 $w=1.68e-07 $l=1.305e-06 $layer=LI1_cond $X=3.85 $Y=1.18
+ $X2=5.155 $Y2=1.18
r65 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.685 $Y=1.095
+ $X2=3.85 $Y2=1.18
r66 7 9 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=3.685 $Y=1.095
+ $X2=3.685 $Y2=0.74
r67 2 17 182 $w=1.7e-07 $l=5.05173e-07 $layer=licon1_NDIFF $count=1 $X=7.715
+ $Y=0.37 $X2=7.855 $Y2=0.81
r68 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.545
+ $Y=0.595 $X2=3.685 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__MUX2_4%A_937_119# 1 2 9 12 16 17 19
r39 19 21 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=6.925 $Y=0.765
+ $X2=6.925 $Y2=0.855
r40 16 17 10.1916 $w=1.83e-07 $l=1.7e-07 $layer=LI1_cond $X=5.495 $Y=0.847
+ $X2=5.665 $Y2=0.847
r41 12 14 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=4.825 $Y=0.75
+ $X2=4.825 $Y2=0.84
r42 9 21 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.76 $Y=0.855
+ $X2=6.925 $Y2=0.855
r43 9 17 71.4385 $w=1.68e-07 $l=1.095e-06 $layer=LI1_cond $X=6.76 $Y=0.855
+ $X2=5.665 $Y2=0.855
r44 8 14 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.99 $Y=0.84
+ $X2=4.825 $Y2=0.84
r45 8 16 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=4.99 $Y=0.84
+ $X2=5.495 $Y2=0.84
r46 2 19 182 $w=1.7e-07 $l=4.59701e-07 $layer=licon1_NDIFF $count=1 $X=6.785
+ $Y=0.37 $X2=6.925 $Y2=0.765
r47 1 12 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=4.685
+ $Y=0.595 $X2=4.825 $Y2=0.75
.ends

