* File: sky130_fd_sc_ls__mux4_1.spice
* Created: Fri Aug 28 13:31:02 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__mux4_1.pex.spice"
.subckt sky130_fd_sc_ls__mux4_1  VNB VPB A0 A1 A2 S0 A3 S1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* S1	S1
* A3	A3
* S0	S0
* A2	A2
* A1	A1
* A0	A0
* VPB	VPB
* VNB	VNB
MM1020 N_VGND_M1020_d N_S0_M1020_g N_A_27_74#_M1020_s VNB NSHORT L=0.15 W=0.64
+ AD=0.192 AS=0.1824 PD=1.24 PS=1.85 NRD=34.68 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75004.9 A=0.096 P=1.58 MULT=1
MM1007 A_264_74# N_A0_M1007_g N_VGND_M1020_d VNB NSHORT L=0.15 W=0.64 AD=0.0768
+ AS=0.192 PD=0.88 PS=1.24 NRD=12.18 NRS=25.308 M=1 R=4.26667 SA=75001
+ SB=75004.2 A=0.096 P=1.58 MULT=1
MM1008 N_A_342_74#_M1008_d N_A_27_74#_M1008_g A_264_74# VNB NSHORT L=0.15 W=0.64
+ AD=0.1248 AS=0.0768 PD=1.03 PS=0.88 NRD=20.616 NRS=12.18 M=1 R=4.26667
+ SA=75001.3 SB=75003.8 A=0.096 P=1.58 MULT=1
MM1018 A_450_74# N_S0_M1018_g N_A_342_74#_M1008_d VNB NSHORT L=0.15 W=0.64
+ AD=0.24 AS=0.1248 PD=1.39 PS=1.03 NRD=60 NRS=0 M=1 R=4.26667 SA=75001.9
+ SB=75003.2 A=0.096 P=1.58 MULT=1
MM1000 N_VGND_M1000_d N_A1_M1000_g A_450_74# VNB NSHORT L=0.15 W=0.64 AD=0.1728
+ AS=0.24 PD=1.18 PS=1.39 NRD=24.372 NRS=60 M=1 R=4.26667 SA=75002.8 SB=75002.3
+ A=0.096 P=1.58 MULT=1
MM1023 A_768_74# N_A2_M1023_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.64 AD=0.0768
+ AS=0.1728 PD=0.88 PS=1.18 NRD=12.18 NRS=24.372 M=1 R=4.26667 SA=75003.5
+ SB=75001.7 A=0.096 P=1.58 MULT=1
MM1021 N_A_846_74#_M1021_d N_A_27_74#_M1021_g A_768_74# VNB NSHORT L=0.15 W=0.64
+ AD=0.1648 AS=0.0768 PD=1.155 PS=0.88 NRD=21.552 NRS=12.18 M=1 R=4.26667
+ SA=75003.9 SB=75001.3 A=0.096 P=1.58 MULT=1
MM1001 A_979_74# N_S0_M1001_g N_A_846_74#_M1021_d VNB NSHORT L=0.15 W=0.64
+ AD=0.0768 AS=0.1648 PD=0.88 PS=1.155 NRD=12.18 NRS=22.488 M=1 R=4.26667
+ SA=75004.5 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1025 N_VGND_M1025_d N_A3_M1025_g A_979_74# VNB NSHORT L=0.15 W=0.64 AD=0.1824
+ AS=0.0768 PD=1.85 PS=0.88 NRD=0 NRS=12.18 M=1 R=4.26667 SA=75004.9 SB=75000.2
+ A=0.096 P=1.58 MULT=1
MM1003 N_A_1338_125#_M1003_d N_S1_M1003_g N_A_846_74#_M1003_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0928 AS=0.454475 PD=0.93 PS=3.19 NRD=0.936 NRS=46.872 M=1
+ R=4.26667 SA=75000.3 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1024 N_A_342_74#_M1024_d N_A_1396_99#_M1024_g N_A_1338_125#_M1003_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.1824 AS=0.0928 PD=1.85 PS=0.93 NRD=0 NRS=0.936 M=1
+ R=4.26667 SA=75000.8 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1005 N_VGND_M1005_d N_S1_M1005_g N_A_1396_99#_M1005_s VNB NSHORT L=0.15 W=0.64
+ AD=0.136255 AS=0.1824 PD=1.07594 PS=1.85 NRD=13.116 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1012 N_X_M1012_d N_A_1338_125#_M1012_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.157545 PD=2.05 PS=1.24406 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75000.7 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1011 N_VPWR_M1011_d N_S0_M1011_g N_A_27_74#_M1011_s VPB PHIGHVT L=0.15 W=1
+ AD=0.229312 AS=0.295 PD=1.57 PS=2.59 NRD=11.8003 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75004.4 A=0.15 P=2.3 MULT=1
MM1004 A_255_341# N_A0_M1004_g N_VPWR_M1011_d VPB PHIGHVT L=0.15 W=1 AD=0.405
+ AS=0.229312 PD=1.81 PS=1.57 NRD=68.9303 NRS=19.0302 M=1 R=6.66667 SA=75000.7
+ SB=75004.2 A=0.15 P=2.3 MULT=1
MM1009 N_A_342_74#_M1009_d N_S0_M1009_g A_255_341# VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.405 PD=1.3 PS=1.81 NRD=1.9503 NRS=68.9303 M=1 R=6.66667
+ SA=75001.7 SB=75003.3 A=0.15 P=2.3 MULT=1
MM1016 A_537_341# N_A_27_74#_M1016_g N_A_342_74#_M1009_d VPB PHIGHVT L=0.15 W=1
+ AD=0.18 AS=0.15 PD=1.36 PS=1.3 NRD=24.6053 NRS=1.9503 M=1 R=6.66667 SA=75002.1
+ SB=75002.8 A=0.15 P=2.3 MULT=1
MM1017 N_VPWR_M1017_d N_A1_M1017_g A_537_341# VPB PHIGHVT L=0.15 W=1 AD=0.2756
+ AS=0.18 PD=1.75 PS=1.36 NRD=43.4385 NRS=24.6053 M=1 R=6.66667 SA=75002.6
+ SB=75002.3 A=0.15 P=2.3 MULT=1
MM1006 A_763_341# N_A2_M1006_g N_VPWR_M1017_d VPB PHIGHVT L=0.15 W=1 AD=0.197625
+ AS=0.2756 PD=1.585 PS=1.75 NRD=28.0922 NRS=43.4385 M=1 R=6.66667 SA=75003.3
+ SB=75001.7 A=0.15 P=2.3 MULT=1
MM1013 N_A_846_74#_M1013_d N_S0_M1013_g A_763_341# VPB PHIGHVT L=0.15 W=1
+ AD=0.4275 AS=0.197625 PD=1.855 PS=1.585 NRD=1.9503 NRS=28.0922 M=1 R=6.66667
+ SA=75003 SB=75001.6 A=0.15 P=2.3 MULT=1
MM1019 A_1065_387# N_A_27_74#_M1019_g N_A_846_74#_M1013_d VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.4275 PD=1.27 PS=1.855 NRD=15.7403 NRS=1.9503 M=1 R=6.66667
+ SA=75004 SB=75000.6 A=0.15 P=2.3 MULT=1
MM1015 N_VPWR_M1015_d N_A3_M1015_g A_1065_387# VPB PHIGHVT L=0.15 W=1 AD=0.295
+ AS=0.135 PD=2.59 PS=1.27 NRD=1.9503 NRS=15.7403 M=1 R=6.66667 SA=75004.4
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1014 N_A_1338_125#_M1014_d N_S1_M1014_g N_A_342_74#_M1014_s VPB PHIGHVT L=0.15
+ W=1 AD=0.175 AS=0.295 PD=1.35 PS=2.59 NRD=11.8003 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75000.8 A=0.15 P=2.3 MULT=1
MM1022 N_A_846_74#_M1022_d N_A_1396_99#_M1022_g N_A_1338_125#_M1014_d VPB
+ PHIGHVT L=0.15 W=1 AD=0.345 AS=0.175 PD=2.69 PS=1.35 NRD=11.8003 NRS=1.9503
+ M=1 R=6.66667 SA=75000.7 SB=75000.3 A=0.15 P=2.3 MULT=1
MM1002 N_VPWR_M1002_d N_S1_M1002_g N_A_1396_99#_M1002_s VPB PHIGHVT L=0.15 W=1
+ AD=0.317241 AS=0.345 PD=1.66038 PS=2.69 NRD=68.95 NRS=11.8003 M=1 R=6.66667
+ SA=75000.3 SB=75001 A=0.15 P=2.3 MULT=1
MM1010 N_X_M1010_d N_A_1338_125#_M1010_g N_VPWR_M1002_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.3472 AS=0.355309 PD=2.86 PS=1.85962 NRD=2.6201 NRS=1.7533 M=1
+ R=7.46667 SA=75001 SB=75000.2 A=0.168 P=2.54 MULT=1
DX26_noxref VNB VPB NWDIODE A=19.0461 P=23.95
c_180 VPB 0 1.25754e-19 $X=0 $Y=3.085
c_1219 A_1065_387# 0 5.47968e-20 $X=5.325 $Y=1.935
*
.include "sky130_fd_sc_ls__mux4_1.pxi.spice"
*
.ends
*
*
