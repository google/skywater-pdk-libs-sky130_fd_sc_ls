# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ls__a311o_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_ls__a311o_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 0.440000 2.335000 0.670000 ;
        RECT 2.005000 0.255000 2.335000 0.440000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 1.450000 1.905000 1.780000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.115000 1.450000 1.365000 1.780000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525000 0.255000 2.875000 0.505000 ;
        RECT 2.525000 0.505000 2.725000 0.670000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.385000 0.255000 3.715000 0.670000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.504100 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.010000 0.605000 1.180000 ;
        RECT 0.125000 1.180000 0.295000 1.850000 ;
        RECT 0.125000 1.850000 0.475000 2.980000 ;
        RECT 0.355000 0.480000 0.605000 1.010000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.480000  1.350000 0.945000 1.680000 ;
      RECT 0.645000  1.950000 1.105000 3.245000 ;
      RECT 0.775000  1.110000 2.570000 1.280000 ;
      RECT 0.775000  1.280000 0.945000 1.350000 ;
      RECT 0.785000  0.085000 1.115000 0.940000 ;
      RECT 1.275000  1.950000 2.595000 2.120000 ;
      RECT 1.275000  2.120000 1.605000 2.980000 ;
      RECT 1.805000  2.290000 2.095000 3.245000 ;
      RECT 2.240000  0.840000 2.570000 1.110000 ;
      RECT 2.240000  1.280000 2.570000 1.445000 ;
      RECT 2.240000  1.445000 3.575000 1.615000 ;
      RECT 2.265000  1.940000 2.595000 1.950000 ;
      RECT 2.265000  2.120000 2.595000 2.980000 ;
      RECT 2.750000  0.855000 3.075000 1.185000 ;
      RECT 2.895000  0.675000 3.215000 0.845000 ;
      RECT 2.895000  0.845000 3.075000 0.855000 ;
      RECT 3.045000  0.085000 3.215000 0.675000 ;
      RECT 3.105000  1.940000 3.575000 2.980000 ;
      RECT 3.245000  1.015000 3.575000 1.445000 ;
      RECT 3.245000  1.615000 3.575000 1.940000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_ls__a311o_1
END LIBRARY
