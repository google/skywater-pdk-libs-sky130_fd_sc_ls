# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ls__o41ai_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ls__o41ai_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.08000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.285000 1.180000 9.955000 1.550000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.365000 1.180000 8.035000 1.550000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.395000 1.180000 6.115000 1.550000 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.180000 3.160000 1.550000 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.780000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.180000 1.145000 1.550000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.586200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.615000 1.720000 3.330000 1.890000 ;
        RECT 0.615000 1.890000 0.945000 2.980000 ;
        RECT 0.625000 0.595000 0.795000 0.840000 ;
        RECT 0.625000 0.840000 1.805000 1.010000 ;
        RECT 1.475000 0.595000 1.805000 0.840000 ;
        RECT 1.475000 1.010000 1.805000 1.720000 ;
        RECT 2.150000 1.890000 3.330000 2.150000 ;
        RECT 2.150000 2.150000 2.430000 2.735000 ;
        RECT 3.050000 2.150000 3.330000 2.735000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 10.080000 0.085000 ;
        RECT 2.475000  0.085000  2.990000 0.600000 ;
        RECT 3.670000  0.085000  3.840000 1.130000 ;
        RECT 4.520000  0.085000  4.850000 0.670000 ;
        RECT 5.450000  0.085000  5.780000 0.670000 ;
        RECT 6.380000  0.085000  6.710000 0.670000 ;
        RECT 7.240000  0.085000  7.570000 0.670000 ;
        RECT 8.205000  0.085000  8.535000 0.670000 ;
        RECT 9.205000  0.085000  9.535000 0.670000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
        RECT 6.395000 -0.085000 6.565000 0.085000 ;
        RECT 6.875000 -0.085000 7.045000 0.085000 ;
        RECT 7.355000 -0.085000 7.525000 0.085000 ;
        RECT 7.835000 -0.085000 8.005000 0.085000 ;
        RECT 8.315000 -0.085000 8.485000 0.085000 ;
        RECT 8.795000 -0.085000 8.965000 0.085000 ;
        RECT 9.275000 -0.085000 9.445000 0.085000 ;
        RECT 9.755000 -0.085000 9.925000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.080000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 10.080000 3.415000 ;
        RECT 0.115000 1.820000  0.445000 3.245000 ;
        RECT 1.115000 2.060000  1.445000 3.245000 ;
        RECT 8.185000 2.060000  8.515000 3.245000 ;
        RECT 9.185000 2.060000  9.515000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
        RECT 6.395000 3.245000 6.565000 3.415000 ;
        RECT 6.875000 3.245000 7.045000 3.415000 ;
        RECT 7.355000 3.245000 7.525000 3.415000 ;
        RECT 7.835000 3.245000 8.005000 3.415000 ;
        RECT 8.315000 3.245000 8.485000 3.415000 ;
        RECT 8.795000 3.245000 8.965000 3.415000 ;
        RECT 9.275000 3.245000 9.445000 3.415000 ;
        RECT 9.755000 3.245000 9.925000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 10.080000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.115000 0.255000 2.305000 0.425000 ;
      RECT 0.115000 0.425000 0.445000 1.010000 ;
      RECT 0.975000 0.425000 1.305000 0.670000 ;
      RECT 1.675000 2.060000 1.980000 2.905000 ;
      RECT 1.675000 2.905000 5.705000 3.075000 ;
      RECT 1.975000 0.425000 2.305000 0.840000 ;
      RECT 1.975000 0.840000 3.500000 1.010000 ;
      RECT 2.600000 2.320000 2.880000 2.905000 ;
      RECT 3.160000 0.350000 3.500000 0.840000 ;
      RECT 3.330000 1.010000 3.500000 1.300000 ;
      RECT 3.330000 1.300000 4.190000 1.470000 ;
      RECT 3.500000 1.800000 3.805000 2.905000 ;
      RECT 3.975000 1.720000 7.565000 1.890000 ;
      RECT 3.975000 1.890000 4.305000 2.735000 ;
      RECT 4.020000 0.350000 4.350000 0.840000 ;
      RECT 4.020000 0.840000 9.965000 1.010000 ;
      RECT 4.020000 1.010000 4.190000 1.300000 ;
      RECT 4.475000 2.060000 4.805000 2.905000 ;
      RECT 4.975000 1.890000 5.205000 2.735000 ;
      RECT 5.030000 0.350000 5.280000 0.840000 ;
      RECT 5.375000 2.060000 5.705000 2.905000 ;
      RECT 5.935000 2.060000 6.265000 2.890000 ;
      RECT 5.935000 2.890000 7.165000 2.905000 ;
      RECT 5.935000 2.905000 8.015000 3.075000 ;
      RECT 5.960000 0.350000 6.210000 0.840000 ;
      RECT 6.435000 1.890000 6.665000 2.720000 ;
      RECT 6.835000 2.060000 7.165000 2.890000 ;
      RECT 6.890000 0.350000 7.060000 0.840000 ;
      RECT 7.335000 1.890000 7.565000 2.735000 ;
      RECT 7.735000 1.720000 9.965000 1.890000 ;
      RECT 7.735000 1.890000 8.015000 2.905000 ;
      RECT 7.785000 0.350000 8.035000 0.840000 ;
      RECT 8.685000 1.890000 9.015000 3.000000 ;
      RECT 8.705000 0.350000 9.035000 0.840000 ;
      RECT 9.685000 1.890000 9.965000 3.000000 ;
      RECT 9.715000 0.350000 9.965000 0.840000 ;
  END
END sky130_fd_sc_ls__o41ai_4
