* File: sky130_fd_sc_ls__and4_2.pxi.spice
* Created: Fri Aug 28 13:05:09 2020
* 
x_PM_SKY130_FD_SC_LS__AND4_2%A N_A_c_69_n N_A_c_75_n N_A_M1002_g N_A_M1007_g
+ N_A_c_71_n N_A_c_72_n A N_A_c_73_n PM_SKY130_FD_SC_LS__AND4_2%A
x_PM_SKY130_FD_SC_LS__AND4_2%B N_B_M1000_g N_B_c_101_n N_B_c_106_n N_B_M1011_g B
+ B B N_B_c_103_n N_B_c_104_n PM_SKY130_FD_SC_LS__AND4_2%B
x_PM_SKY130_FD_SC_LS__AND4_2%C N_C_M1010_g N_C_c_143_n N_C_c_148_n N_C_M1005_g C
+ C C N_C_c_145_n N_C_c_146_n PM_SKY130_FD_SC_LS__AND4_2%C
x_PM_SKY130_FD_SC_LS__AND4_2%D N_D_M1008_g N_D_M1006_g N_D_c_182_n N_D_c_187_n D
+ N_D_c_183_n N_D_c_184_n N_D_c_185_n PM_SKY130_FD_SC_LS__AND4_2%D
x_PM_SKY130_FD_SC_LS__AND4_2%A_56_74# N_A_56_74#_M1007_s N_A_56_74#_M1002_d
+ N_A_56_74#_M1005_d N_A_56_74#_M1003_g N_A_56_74#_c_231_n N_A_56_74#_M1001_g
+ N_A_56_74#_M1009_g N_A_56_74#_c_232_n N_A_56_74#_M1004_g N_A_56_74#_c_225_n
+ N_A_56_74#_c_226_n N_A_56_74#_c_227_n N_A_56_74#_c_235_n N_A_56_74#_c_236_n
+ N_A_56_74#_c_262_n N_A_56_74#_c_237_n N_A_56_74#_c_238_n N_A_56_74#_c_228_n
+ N_A_56_74#_c_229_n N_A_56_74#_c_230_n N_A_56_74#_c_240_n N_A_56_74#_c_275_n
+ PM_SKY130_FD_SC_LS__AND4_2%A_56_74#
x_PM_SKY130_FD_SC_LS__AND4_2%VPWR N_VPWR_M1002_s N_VPWR_M1011_d N_VPWR_M1008_d
+ N_VPWR_M1004_s N_VPWR_c_338_n N_VPWR_c_339_n N_VPWR_c_340_n N_VPWR_c_341_n
+ N_VPWR_c_342_n N_VPWR_c_343_n N_VPWR_c_344_n N_VPWR_c_345_n N_VPWR_c_346_n
+ N_VPWR_c_347_n VPWR N_VPWR_c_348_n N_VPWR_c_337_n
+ PM_SKY130_FD_SC_LS__AND4_2%VPWR
x_PM_SKY130_FD_SC_LS__AND4_2%X N_X_M1003_s N_X_M1001_d X X X X N_X_c_388_n
+ PM_SKY130_FD_SC_LS__AND4_2%X
x_PM_SKY130_FD_SC_LS__AND4_2%VGND N_VGND_M1006_d N_VGND_M1009_d N_VGND_c_411_n
+ N_VGND_c_412_n N_VGND_c_413_n N_VGND_c_414_n N_VGND_c_415_n N_VGND_c_416_n
+ N_VGND_c_417_n VGND N_VGND_c_418_n N_VGND_c_419_n
+ PM_SKY130_FD_SC_LS__AND4_2%VGND
cc_1 VNB N_A_c_69_n 0.00155843f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.795
cc_2 VNB N_A_M1007_g 0.0287743f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=0.74
cc_3 VNB N_A_c_71_n 0.0547136f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.465
cc_4 VNB N_A_c_72_n 0.0132577f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.3
cc_5 VNB N_A_c_73_n 0.0086234f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.465
cc_6 VNB N_B_c_101_n 0.00695258f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=2.46
cc_7 VNB B 0.00459753f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_B_c_103_n 0.0308072f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.465
cc_9 VNB N_B_c_104_n 0.0180773f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.465
cc_10 VNB N_C_c_143_n 0.00710459f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=2.46
cc_11 VNB C 0.00242177f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_C_c_145_n 0.0326377f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.465
cc_13 VNB N_C_c_146_n 0.0195889f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.465
cc_14 VNB N_D_c_182_n 0.00655899f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_D_c_183_n 0.033522f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.465
cc_16 VNB N_D_c_184_n 0.0101128f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.465
cc_17 VNB N_D_c_185_n 0.0197696f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.465
cc_18 VNB N_A_56_74#_M1003_g 0.0225826f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_19 VNB N_A_56_74#_M1009_g 0.0273222f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_56_74#_c_225_n 0.0467635f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_56_74#_c_226_n 0.0258829f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_56_74#_c_227_n 0.00377606f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_56_74#_c_228_n 0.00710428f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_56_74#_c_229_n 0.0577987f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_56_74#_c_230_n 0.0094188f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VPWR_c_337_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB X 0.00144878f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=0.74
cc_28 VNB N_X_c_388_n 7.53866e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_411_n 0.0091706f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_412_n 0.016267f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.3
cc_31 VNB N_VGND_c_413_n 0.0111347f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_32 VNB N_VGND_c_414_n 0.0182112f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.465
cc_33 VNB N_VGND_c_415_n 0.0671414f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.465
cc_34 VNB N_VGND_c_416_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_417_n 0.00867839f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_418_n 0.0196671f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_419_n 0.258397f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VPB N_A_c_69_n 0.0075559f $X=-0.19 $Y=1.66 $X2=0.595 $Y2=1.795
cc_39 VPB N_A_c_75_n 0.0262416f $X=-0.19 $Y=1.66 $X2=0.595 $Y2=1.885
cc_40 VPB N_A_c_73_n 0.00823058f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=1.465
cc_41 VPB N_B_c_101_n 0.00766537f $X=-0.19 $Y=1.66 $X2=0.595 $Y2=2.46
cc_42 VPB N_B_c_106_n 0.0224387f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.3
cc_43 VPB N_C_c_143_n 0.00778252f $X=-0.19 $Y=1.66 $X2=0.595 $Y2=2.46
cc_44 VPB N_C_c_148_n 0.0224923f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.3
cc_45 VPB N_D_c_182_n 0.00741153f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_D_c_187_n 0.0230513f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.465
cc_47 VPB N_A_56_74#_c_231_n 0.0167666f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=1.465
cc_48 VPB N_A_56_74#_c_232_n 0.0161592f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 VPB N_A_56_74#_c_225_n 0.0134803f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_A_56_74#_c_227_n 5.66269e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_51 VPB N_A_56_74#_c_235_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_A_56_74#_c_236_n 0.0275577f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_A_56_74#_c_237_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_A_56_74#_c_238_n 0.00748573f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_A_56_74#_c_228_n 0.026493f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_A_56_74#_c_240_n 0.00692367f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_338_n 0.0121909f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_339_n 0.0539929f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=1.465
cc_59 VPB N_VPWR_c_340_n 0.00988978f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_341_n 0.00993905f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_342_n 0.0126718f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_343_n 0.025422f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_344_n 0.0215645f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_345_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_346_n 0.0213997f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_347_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_348_n 0.0234846f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_337_n 0.0661765f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 N_A_c_69_n N_B_c_101_n 0.00653161f $X=0.595 $Y=1.795 $X2=0 $Y2=0
cc_70 N_A_c_75_n N_B_c_106_n 0.0147625f $X=0.595 $Y=1.885 $X2=0 $Y2=0
cc_71 N_A_M1007_g B 0.00235149f $X=0.64 $Y=0.74 $X2=0 $Y2=0
cc_72 N_A_c_72_n N_B_c_103_n 0.0369205f $X=0.505 $Y=1.3 $X2=0 $Y2=0
cc_73 N_A_M1007_g N_B_c_104_n 0.0303889f $X=0.64 $Y=0.74 $X2=0 $Y2=0
cc_74 N_A_M1007_g N_A_56_74#_c_226_n 0.0109243f $X=0.64 $Y=0.74 $X2=0 $Y2=0
cc_75 N_A_c_69_n N_A_56_74#_c_227_n 0.00179792f $X=0.595 $Y=1.795 $X2=0 $Y2=0
cc_76 N_A_M1007_g N_A_56_74#_c_227_n 0.00887397f $X=0.64 $Y=0.74 $X2=0 $Y2=0
cc_77 N_A_c_72_n N_A_56_74#_c_227_n 0.00952112f $X=0.505 $Y=1.3 $X2=0 $Y2=0
cc_78 N_A_c_73_n N_A_56_74#_c_227_n 0.030293f $X=0.28 $Y=1.465 $X2=0 $Y2=0
cc_79 N_A_c_75_n N_A_56_74#_c_235_n 0.0174114f $X=0.595 $Y=1.885 $X2=0 $Y2=0
cc_80 N_A_M1007_g N_A_56_74#_c_230_n 0.0116482f $X=0.64 $Y=0.74 $X2=0 $Y2=0
cc_81 N_A_c_71_n N_A_56_74#_c_230_n 0.00604202f $X=0.505 $Y=1.465 $X2=0 $Y2=0
cc_82 N_A_c_73_n N_A_56_74#_c_230_n 0.0143044f $X=0.28 $Y=1.465 $X2=0 $Y2=0
cc_83 N_A_c_69_n N_A_56_74#_c_240_n 0.00243422f $X=0.595 $Y=1.795 $X2=0 $Y2=0
cc_84 N_A_c_75_n N_A_56_74#_c_240_n 0.00600565f $X=0.595 $Y=1.885 $X2=0 $Y2=0
cc_85 N_A_c_73_n N_A_56_74#_c_240_n 0.00503427f $X=0.28 $Y=1.465 $X2=0 $Y2=0
cc_86 N_A_c_75_n N_VPWR_c_339_n 0.0269837f $X=0.595 $Y=1.885 $X2=0 $Y2=0
cc_87 N_A_c_71_n N_VPWR_c_339_n 0.00181048f $X=0.505 $Y=1.465 $X2=0 $Y2=0
cc_88 N_A_c_73_n N_VPWR_c_339_n 0.0299469f $X=0.28 $Y=1.465 $X2=0 $Y2=0
cc_89 N_A_c_75_n N_VPWR_c_344_n 0.00400282f $X=0.595 $Y=1.885 $X2=0 $Y2=0
cc_90 N_A_c_75_n N_VPWR_c_337_n 0.00714906f $X=0.595 $Y=1.885 $X2=0 $Y2=0
cc_91 N_A_M1007_g N_VGND_c_415_n 0.00434272f $X=0.64 $Y=0.74 $X2=0 $Y2=0
cc_92 N_A_M1007_g N_VGND_c_419_n 0.0082504f $X=0.64 $Y=0.74 $X2=0 $Y2=0
cc_93 N_B_c_101_n N_C_c_143_n 0.00440326f $X=1.045 $Y=1.795 $X2=0 $Y2=0
cc_94 N_B_c_106_n N_C_c_148_n 0.0223942f $X=1.045 $Y=1.885 $X2=0 $Y2=0
cc_95 B C 0.0744187f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_96 N_B_c_103_n C 3.9854e-19 $X=1.12 $Y=1.385 $X2=0 $Y2=0
cc_97 N_B_c_104_n C 7.46328e-19 $X=1.12 $Y=1.22 $X2=0 $Y2=0
cc_98 N_B_c_103_n N_C_c_145_n 0.0175135f $X=1.12 $Y=1.385 $X2=0 $Y2=0
cc_99 B N_C_c_146_n 0.00774327f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_100 N_B_c_104_n N_C_c_146_n 0.024906f $X=1.12 $Y=1.22 $X2=0 $Y2=0
cc_101 B N_A_56_74#_c_226_n 0.0212655f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_102 N_B_c_104_n N_A_56_74#_c_226_n 0.00182282f $X=1.12 $Y=1.22 $X2=0 $Y2=0
cc_103 B N_A_56_74#_c_227_n 0.031739f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_104 N_B_c_104_n N_A_56_74#_c_227_n 0.00586721f $X=1.12 $Y=1.22 $X2=0 $Y2=0
cc_105 N_B_c_106_n N_A_56_74#_c_235_n 0.0151124f $X=1.045 $Y=1.885 $X2=0 $Y2=0
cc_106 N_B_c_101_n N_A_56_74#_c_236_n 0.00431415f $X=1.045 $Y=1.795 $X2=0 $Y2=0
cc_107 N_B_c_106_n N_A_56_74#_c_236_n 0.00898393f $X=1.045 $Y=1.885 $X2=0 $Y2=0
cc_108 B N_A_56_74#_c_236_n 0.025829f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_109 N_B_c_103_n N_A_56_74#_c_236_n 0.00105742f $X=1.12 $Y=1.385 $X2=0 $Y2=0
cc_110 N_B_c_106_n N_A_56_74#_c_262_n 7.77169e-19 $X=1.045 $Y=1.885 $X2=0 $Y2=0
cc_111 B N_A_56_74#_c_230_n 0.0137062f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_112 N_B_c_104_n N_A_56_74#_c_230_n 9.65577e-19 $X=1.12 $Y=1.22 $X2=0 $Y2=0
cc_113 N_B_c_101_n N_A_56_74#_c_240_n 0.00146745f $X=1.045 $Y=1.795 $X2=0 $Y2=0
cc_114 N_B_c_106_n N_A_56_74#_c_240_n 0.00165207f $X=1.045 $Y=1.885 $X2=0 $Y2=0
cc_115 B N_A_56_74#_c_240_n 0.00245488f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_116 N_B_c_106_n N_VPWR_c_340_n 0.0126176f $X=1.045 $Y=1.885 $X2=0 $Y2=0
cc_117 N_B_c_106_n N_VPWR_c_344_n 0.00445602f $X=1.045 $Y=1.885 $X2=0 $Y2=0
cc_118 N_B_c_106_n N_VPWR_c_337_n 0.00860001f $X=1.045 $Y=1.885 $X2=0 $Y2=0
cc_119 B A_221_74# 0.00939544f $X=1.115 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_120 B N_VGND_c_415_n 0.0102495f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_121 N_B_c_104_n N_VGND_c_415_n 0.00304348f $X=1.12 $Y=1.22 $X2=0 $Y2=0
cc_122 B N_VGND_c_419_n 0.0117398f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_123 N_B_c_104_n N_VGND_c_419_n 0.00371612f $X=1.12 $Y=1.22 $X2=0 $Y2=0
cc_124 N_C_c_143_n N_D_c_182_n 0.0110466f $X=1.705 $Y=1.795 $X2=0 $Y2=0
cc_125 N_C_c_143_n N_D_c_187_n 0.00416562f $X=1.705 $Y=1.795 $X2=0 $Y2=0
cc_126 N_C_c_148_n N_D_c_187_n 0.00821772f $X=1.705 $Y=1.885 $X2=0 $Y2=0
cc_127 C N_D_c_183_n 3.80049e-19 $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_128 N_C_c_145_n N_D_c_183_n 0.0174582f $X=1.69 $Y=1.385 $X2=0 $Y2=0
cc_129 C N_D_c_184_n 0.0273797f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_130 N_C_c_145_n N_D_c_184_n 0.00202602f $X=1.69 $Y=1.385 $X2=0 $Y2=0
cc_131 C N_D_c_185_n 0.00922273f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_132 N_C_c_146_n N_D_c_185_n 0.0242189f $X=1.69 $Y=1.22 $X2=0 $Y2=0
cc_133 N_C_c_148_n N_A_56_74#_c_235_n 9.17041e-19 $X=1.705 $Y=1.885 $X2=0 $Y2=0
cc_134 N_C_c_143_n N_A_56_74#_c_236_n 0.00582404f $X=1.705 $Y=1.795 $X2=0 $Y2=0
cc_135 N_C_c_148_n N_A_56_74#_c_236_n 0.0106833f $X=1.705 $Y=1.885 $X2=0 $Y2=0
cc_136 C N_A_56_74#_c_236_n 0.0263044f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_137 N_C_c_145_n N_A_56_74#_c_236_n 0.00108599f $X=1.69 $Y=1.385 $X2=0 $Y2=0
cc_138 N_C_c_148_n N_A_56_74#_c_262_n 0.00722962f $X=1.705 $Y=1.885 $X2=0 $Y2=0
cc_139 N_C_c_148_n N_A_56_74#_c_237_n 0.00572924f $X=1.705 $Y=1.885 $X2=0 $Y2=0
cc_140 N_C_c_148_n N_A_56_74#_c_275_n 0.00186907f $X=1.705 $Y=1.885 $X2=0 $Y2=0
cc_141 N_C_c_148_n N_VPWR_c_340_n 0.0127027f $X=1.705 $Y=1.885 $X2=0 $Y2=0
cc_142 N_C_c_148_n N_VPWR_c_346_n 0.00445602f $X=1.705 $Y=1.885 $X2=0 $Y2=0
cc_143 N_C_c_148_n N_VPWR_c_337_n 0.00859777f $X=1.705 $Y=1.885 $X2=0 $Y2=0
cc_144 C A_335_74# 0.0102591f $X=1.595 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_145 C N_VGND_c_415_n 0.00930091f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_146 N_C_c_146_n N_VGND_c_415_n 0.00304348f $X=1.69 $Y=1.22 $X2=0 $Y2=0
cc_147 C N_VGND_c_419_n 0.0106938f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_148 N_C_c_146_n N_VGND_c_419_n 0.00373154f $X=1.69 $Y=1.22 $X2=0 $Y2=0
cc_149 N_D_c_183_n N_A_56_74#_M1003_g 0.0181812f $X=2.26 $Y=1.385 $X2=0 $Y2=0
cc_150 N_D_c_184_n N_A_56_74#_M1003_g 0.00180549f $X=2.26 $Y=1.385 $X2=0 $Y2=0
cc_151 N_D_c_185_n N_A_56_74#_M1003_g 0.0138101f $X=2.26 $Y=1.22 $X2=0 $Y2=0
cc_152 N_D_c_182_n N_A_56_74#_c_231_n 0.00275438f $X=2.162 $Y=1.79 $X2=0 $Y2=0
cc_153 N_D_c_187_n N_A_56_74#_c_231_n 0.0255426f $X=2.162 $Y=1.885 $X2=0 $Y2=0
cc_154 N_D_c_182_n N_A_56_74#_c_225_n 0.00636274f $X=2.162 $Y=1.79 $X2=0 $Y2=0
cc_155 N_D_c_182_n N_A_56_74#_c_236_n 0.00235788f $X=2.162 $Y=1.79 $X2=0 $Y2=0
cc_156 N_D_c_187_n N_A_56_74#_c_236_n 0.00348199f $X=2.162 $Y=1.885 $X2=0 $Y2=0
cc_157 N_D_c_184_n N_A_56_74#_c_236_n 0.0044594f $X=2.26 $Y=1.385 $X2=0 $Y2=0
cc_158 N_D_c_187_n N_A_56_74#_c_262_n 0.00957073f $X=2.162 $Y=1.885 $X2=0 $Y2=0
cc_159 N_D_c_187_n N_A_56_74#_c_237_n 0.00719071f $X=2.162 $Y=1.885 $X2=0 $Y2=0
cc_160 N_D_c_187_n N_A_56_74#_c_238_n 0.0139895f $X=2.162 $Y=1.885 $X2=0 $Y2=0
cc_161 N_D_c_187_n N_A_56_74#_c_275_n 2.24111e-19 $X=2.162 $Y=1.885 $X2=0 $Y2=0
cc_162 N_D_c_187_n N_VPWR_c_341_n 0.00636186f $X=2.162 $Y=1.885 $X2=0 $Y2=0
cc_163 N_D_c_187_n N_VPWR_c_346_n 0.00445602f $X=2.162 $Y=1.885 $X2=0 $Y2=0
cc_164 N_D_c_187_n N_VPWR_c_337_n 0.00454315f $X=2.162 $Y=1.885 $X2=0 $Y2=0
cc_165 N_D_c_182_n X 0.00145145f $X=2.162 $Y=1.79 $X2=0 $Y2=0
cc_166 N_D_c_187_n X 0.00115345f $X=2.162 $Y=1.885 $X2=0 $Y2=0
cc_167 N_D_c_183_n X 2.48447e-19 $X=2.26 $Y=1.385 $X2=0 $Y2=0
cc_168 N_D_c_184_n X 0.0146227f $X=2.26 $Y=1.385 $X2=0 $Y2=0
cc_169 N_D_c_185_n N_X_c_388_n 3.54267e-19 $X=2.26 $Y=1.22 $X2=0 $Y2=0
cc_170 N_D_c_183_n N_VGND_c_411_n 0.00103009f $X=2.26 $Y=1.385 $X2=0 $Y2=0
cc_171 N_D_c_184_n N_VGND_c_411_n 0.0122839f $X=2.26 $Y=1.385 $X2=0 $Y2=0
cc_172 N_D_c_185_n N_VGND_c_411_n 0.00413006f $X=2.26 $Y=1.22 $X2=0 $Y2=0
cc_173 N_D_c_185_n N_VGND_c_415_n 0.00461464f $X=2.26 $Y=1.22 $X2=0 $Y2=0
cc_174 N_D_c_185_n N_VGND_c_419_n 0.00910053f $X=2.26 $Y=1.22 $X2=0 $Y2=0
cc_175 N_A_56_74#_c_238_n N_VPWR_M1008_d 0.0186086f $X=3.405 $Y=2.405 $X2=0
+ $Y2=0
cc_176 N_A_56_74#_c_238_n N_VPWR_M1004_s 0.00685378f $X=3.405 $Y=2.405 $X2=0
+ $Y2=0
cc_177 N_A_56_74#_c_228_n N_VPWR_M1004_s 0.0117108f $X=3.57 $Y=1.465 $X2=0 $Y2=0
cc_178 N_A_56_74#_c_235_n N_VPWR_c_339_n 0.0806812f $X=0.82 $Y=2.105 $X2=0 $Y2=0
cc_179 N_A_56_74#_c_235_n N_VPWR_c_340_n 0.0571325f $X=0.82 $Y=2.105 $X2=0 $Y2=0
cc_180 N_A_56_74#_c_236_n N_VPWR_c_340_n 0.0271222f $X=1.765 $Y=1.805 $X2=0
+ $Y2=0
cc_181 N_A_56_74#_c_262_n N_VPWR_c_340_n 0.0165245f $X=1.93 $Y=2.105 $X2=0 $Y2=0
cc_182 N_A_56_74#_c_237_n N_VPWR_c_340_n 0.0312009f $X=1.93 $Y=2.815 $X2=0 $Y2=0
cc_183 N_A_56_74#_c_275_n N_VPWR_c_340_n 0.0114735f $X=1.93 $Y=2.405 $X2=0 $Y2=0
cc_184 N_A_56_74#_c_231_n N_VPWR_c_341_n 0.0123794f $X=2.775 $Y=1.765 $X2=0
+ $Y2=0
cc_185 N_A_56_74#_c_237_n N_VPWR_c_341_n 0.0215387f $X=1.93 $Y=2.815 $X2=0 $Y2=0
cc_186 N_A_56_74#_c_238_n N_VPWR_c_341_n 0.0261009f $X=3.405 $Y=2.405 $X2=0
+ $Y2=0
cc_187 N_A_56_74#_c_232_n N_VPWR_c_343_n 0.0179113f $X=3.225 $Y=1.765 $X2=0
+ $Y2=0
cc_188 N_A_56_74#_c_238_n N_VPWR_c_343_n 0.0307621f $X=3.405 $Y=2.405 $X2=0
+ $Y2=0
cc_189 N_A_56_74#_c_235_n N_VPWR_c_344_n 0.0162172f $X=0.82 $Y=2.105 $X2=0 $Y2=0
cc_190 N_A_56_74#_c_237_n N_VPWR_c_346_n 0.014552f $X=1.93 $Y=2.815 $X2=0 $Y2=0
cc_191 N_A_56_74#_c_231_n N_VPWR_c_348_n 0.00461464f $X=2.775 $Y=1.765 $X2=0
+ $Y2=0
cc_192 N_A_56_74#_c_232_n N_VPWR_c_348_n 0.00461464f $X=3.225 $Y=1.765 $X2=0
+ $Y2=0
cc_193 N_A_56_74#_c_231_n N_VPWR_c_337_n 0.00465735f $X=2.775 $Y=1.765 $X2=0
+ $Y2=0
cc_194 N_A_56_74#_c_232_n N_VPWR_c_337_n 0.00468139f $X=3.225 $Y=1.765 $X2=0
+ $Y2=0
cc_195 N_A_56_74#_c_235_n N_VPWR_c_337_n 0.0132635f $X=0.82 $Y=2.105 $X2=0 $Y2=0
cc_196 N_A_56_74#_c_237_n N_VPWR_c_337_n 0.0119791f $X=1.93 $Y=2.815 $X2=0 $Y2=0
cc_197 N_A_56_74#_c_238_n N_VPWR_c_337_n 0.0323619f $X=3.405 $Y=2.405 $X2=0
+ $Y2=0
cc_198 N_A_56_74#_c_238_n N_X_M1001_d 0.00571673f $X=3.405 $Y=2.405 $X2=0 $Y2=0
cc_199 N_A_56_74#_M1003_g X 0.00294214f $X=2.74 $Y=0.74 $X2=0 $Y2=0
cc_200 N_A_56_74#_c_231_n X 0.00908633f $X=2.775 $Y=1.765 $X2=0 $Y2=0
cc_201 N_A_56_74#_M1009_g X 0.0106301f $X=3.17 $Y=0.74 $X2=0 $Y2=0
cc_202 N_A_56_74#_c_232_n X 0.00776126f $X=3.225 $Y=1.765 $X2=0 $Y2=0
cc_203 N_A_56_74#_c_225_n X 0.0395251f $X=3.315 $Y=1.465 $X2=0 $Y2=0
cc_204 N_A_56_74#_c_238_n X 0.0225136f $X=3.405 $Y=2.405 $X2=0 $Y2=0
cc_205 N_A_56_74#_c_228_n X 0.0663603f $X=3.57 $Y=1.465 $X2=0 $Y2=0
cc_206 N_A_56_74#_M1003_g N_X_c_388_n 0.00713606f $X=2.74 $Y=0.74 $X2=0 $Y2=0
cc_207 N_A_56_74#_M1009_g N_X_c_388_n 0.0119323f $X=3.17 $Y=0.74 $X2=0 $Y2=0
cc_208 N_A_56_74#_c_230_n A_143_74# 0.00178387f $X=0.7 $Y=1.045 $X2=-0.19
+ $Y2=-0.245
cc_209 N_A_56_74#_M1003_g N_VGND_c_411_n 0.0125291f $X=2.74 $Y=0.74 $X2=0 $Y2=0
cc_210 N_A_56_74#_M1003_g N_VGND_c_413_n 0.00110029f $X=2.74 $Y=0.74 $X2=0 $Y2=0
cc_211 N_A_56_74#_M1009_g N_VGND_c_413_n 0.00595376f $X=3.17 $Y=0.74 $X2=0 $Y2=0
cc_212 N_A_56_74#_M1009_g N_VGND_c_414_n 0.0103157f $X=3.17 $Y=0.74 $X2=0 $Y2=0
cc_213 N_A_56_74#_c_228_n N_VGND_c_414_n 0.0178142f $X=3.57 $Y=1.465 $X2=0 $Y2=0
cc_214 N_A_56_74#_c_229_n N_VGND_c_414_n 0.00190129f $X=3.57 $Y=1.465 $X2=0
+ $Y2=0
cc_215 N_A_56_74#_c_226_n N_VGND_c_415_n 0.0144497f $X=0.425 $Y=0.515 $X2=0
+ $Y2=0
cc_216 N_A_56_74#_M1009_g N_VGND_c_417_n 0.00481221f $X=3.17 $Y=0.74 $X2=0 $Y2=0
cc_217 N_A_56_74#_c_225_n N_VGND_c_417_n 0.00343719f $X=3.315 $Y=1.465 $X2=0
+ $Y2=0
cc_218 N_A_56_74#_M1003_g N_VGND_c_418_n 0.00461464f $X=2.74 $Y=0.74 $X2=0 $Y2=0
cc_219 N_A_56_74#_M1009_g N_VGND_c_418_n 0.00383152f $X=3.17 $Y=0.74 $X2=0 $Y2=0
cc_220 N_A_56_74#_M1003_g N_VGND_c_419_n 0.00835925f $X=2.74 $Y=0.74 $X2=0 $Y2=0
cc_221 N_A_56_74#_M1009_g N_VGND_c_419_n 0.0036906f $X=3.17 $Y=0.74 $X2=0 $Y2=0
cc_222 N_A_56_74#_c_226_n N_VGND_c_419_n 0.0119539f $X=0.425 $Y=0.515 $X2=0
+ $Y2=0
cc_223 N_X_c_388_n N_VGND_c_411_n 0.017139f $X=2.955 $Y=0.91 $X2=0 $Y2=0
cc_224 N_X_c_388_n N_VGND_c_414_n 0.0241034f $X=2.955 $Y=0.91 $X2=0 $Y2=0
cc_225 N_X_c_388_n N_VGND_c_417_n 0.00106652f $X=2.955 $Y=0.91 $X2=0 $Y2=0
cc_226 N_X_c_388_n N_VGND_c_419_n 0.0167375f $X=2.955 $Y=0.91 $X2=0 $Y2=0
