* NGSPICE file created from sky130_fd_sc_ls__einvp_2.ext - technology: sky130A

.subckt sky130_fd_sc_ls__einvp_2 A TE VGND VNB VPB VPWR Z
M1000 a_27_368# a_263_323# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=9.912e+11p pd=8.49e+06u as=5.248e+11p ps=4.71e+06u
M1001 a_36_74# A Z VNB nshort w=740000u l=150000u
+  ad=6.29e+11p pd=6.14e+06u as=2.072e+11p ps=2.04e+06u
M1002 VPWR TE a_263_323# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.856e+11p ps=1.86e+06u
M1003 VGND TE a_36_74# VNB nshort w=740000u l=150000u
+  ad=3.332e+11p pd=3.48e+06u as=0p ps=0u
M1004 Z A a_27_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=0p ps=0u
M1005 a_27_368# A Z VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR a_263_323# a_27_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_36_74# TE VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Z A a_36_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND TE a_263_323# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
.ends

