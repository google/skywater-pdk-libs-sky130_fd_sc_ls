* NGSPICE file created from sky130_fd_sc_ls__nand2b_4.ext - technology: sky130A

.subckt sky130_fd_sc_ls__nand2b_4 A_N B VGND VNB VPB VPWR Y
M1000 VGND B a_243_74# VNB nshort w=740000u l=150000u
+  ad=1.0286e+12p pd=7.22e+06u as=1.0434e+12p ps=1.022e+07u
M1001 Y a_31_74# a_243_74# VNB nshort w=740000u l=150000u
+  ad=5.143e+11p pd=4.35e+06u as=0p ps=0u
M1002 Y a_31_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=1.12e+12p pd=6.48e+06u as=3.0716e+12p ps=1.425e+07u
M1003 a_243_74# B VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR B Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND B a_243_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_243_74# a_31_74# Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND A_N a_31_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1008 a_31_74# A_N VPWR VPB phighvt w=840000u l=150000u
+  ad=2.52e+11p pd=2.28e+06u as=0p ps=0u
M1009 Y B VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_243_74# a_31_74# Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR a_31_74# Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR A_N a_31_74# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 Y a_31_74# a_243_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_243_74# B VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

