* File: sky130_fd_sc_ls__dfrtp_2.spice
* Created: Wed Sep  2 11:01:13 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__dfrtp_2.pex.spice"
.subckt sky130_fd_sc_ls__dfrtp_2  VNB VPB D CLK RESET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* RESET_B	RESET_B
* CLK	CLK
* D	D
* VPB	VPB
* VNB	VNB
MM1025 A_117_78# N_D_M1025_g N_A_30_78#_M1025_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1009 N_VGND_M1009_d N_RESET_B_M1009_g A_117_78# VNB NSHORT L=0.15 W=0.42
+ AD=0.1344 AS=0.0504 PD=1.48 PS=0.66 NRD=9.996 NRS=18.564 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1015 N_VGND_M1015_d N_CLK_M1015_g N_A_309_390#_M1015_s VNB NSHORT L=0.15
+ W=0.74 AD=0.162375 AS=0.2646 PD=1.255 PS=2.4 NRD=9.72 NRS=5.268 M=1 R=4.93333
+ SA=75000.2 SB=75000.8 A=0.111 P=1.78 MULT=1
MM1012 N_A_495_390#_M1012_d N_A_309_390#_M1012_g N_VGND_M1015_d VNB NSHORT
+ L=0.15 W=0.74 AD=0.20885 AS=0.162375 PD=2.07 PS=1.255 NRD=1.62 NRS=9.72 M=1
+ R=4.93333 SA=75000.8 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1016 N_A_697_463#_M1016_d N_A_309_390#_M1016_g N_A_30_78#_M1016_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0735 AS=0.1197 PD=0.77 PS=1.41 NRD=19.992 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75003.7 A=0.063 P=1.14 MULT=1
MM1014 A_823_138# N_A_495_390#_M1014_g N_A_697_463#_M1016_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.0735 PD=0.66 PS=0.77 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75000.7 SB=75003.2 A=0.063 P=1.14 MULT=1
MM1006 A_901_138# N_A_839_359#_M1006_g A_823_138# VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0504 PD=0.63 PS=0.66 NRD=14.28 NRS=18.564 M=1 R=2.8 SA=75001.1
+ SB=75002.8 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_RESET_B_M1001_g A_901_138# VNB NSHORT L=0.15 W=0.42
+ AD=0.255829 AS=0.0441 PD=1.33241 PS=0.63 NRD=158.316 NRS=14.28 M=1 R=2.8
+ SA=75001.5 SB=75002.4 A=0.063 P=1.14 MULT=1
MM1020 N_A_839_359#_M1020_d N_A_697_463#_M1020_g N_VGND_M1001_d VNB NSHORT
+ L=0.15 W=0.74 AD=0.12025 AS=0.450746 PD=1.065 PS=2.34759 NRD=0 NRS=89.856 M=1
+ R=4.93333 SA=75001.7 SB=75002 A=0.111 P=1.78 MULT=1
MM1003 N_A_1271_74#_M1003_d N_A_495_390#_M1003_g N_A_839_359#_M1020_d VNB NSHORT
+ L=0.15 W=0.74 AD=0.292172 AS=0.12025 PD=2.09241 PS=1.065 NRD=4.044 NRS=7.296
+ M=1 R=4.93333 SA=75002.2 SB=75001.5 A=0.111 P=1.78 MULT=1
MM1031 A_1481_81# N_A_309_390#_M1031_g N_A_1271_74#_M1003_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.165828 PD=0.66 PS=1.18759 NRD=18.564 NRS=47.136 M=1
+ R=2.8 SA=75002.8 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1005_d N_A_1525_212#_M1005_g A_1481_81# VNB NSHORT L=0.15 W=0.42
+ AD=0.0777 AS=0.0504 PD=0.79 PS=0.66 NRD=12.852 NRS=18.564 M=1 R=2.8 SA=75003.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1017 A_1663_81# N_RESET_B_M1017_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0777 PD=0.66 PS=0.79 NRD=18.564 NRS=12.852 M=1 R=2.8 SA=75003.7
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1018 N_A_1525_212#_M1018_d N_A_1271_74#_M1018_g A_1663_81# VNB NSHORT L=0.15
+ W=0.42 AD=0.1176 AS=0.0504 PD=1.4 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8
+ SA=75004.1 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1019 N_A_1921_409#_M1019_d N_A_1271_74#_M1019_g N_VGND_M1019_s VNB NSHORT
+ L=0.15 W=0.74 AD=0.2109 AS=0.2072 PD=2.05 PS=2.04 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1029 N_Q_M1029_d N_A_1921_409#_M1029_g N_VGND_M1029_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1032 N_Q_M1029_d N_A_1921_409#_M1032_g N_VGND_M1032_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.2072 PD=1.02 PS=2.04 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1022 N_A_30_78#_M1022_d N_D_M1022_g N_VPWR_M1022_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.063 AS=0.1197 PD=0.72 PS=1.41 NRD=4.6886 NRS=4.6886 M=1 R=2.8 SA=75000.2
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1023 N_VPWR_M1023_d N_RESET_B_M1023_g N_A_30_78#_M1022_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1197 AS=0.063 PD=1.41 PS=0.72 NRD=9.3772 NRS=4.6886 M=1 R=2.8
+ SA=75000.7 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1027 N_VPWR_M1027_d N_CLK_M1027_g N_A_309_390#_M1027_s VPB PHIGHVT L=0.15 W=1
+ AD=0.1725 AS=0.2688 PD=1.345 PS=2.57 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75000.7 A=0.15 P=2.3 MULT=1
MM1004 N_A_495_390#_M1004_d N_A_309_390#_M1004_g N_VPWR_M1027_d VPB PHIGHVT
+ L=0.15 W=1 AD=0.265 AS=0.1725 PD=2.53 PS=1.345 NRD=0 NRS=12.7853 M=1 R=6.66667
+ SA=75000.7 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1008 N_A_697_463#_M1008_d N_A_495_390#_M1008_g N_A_30_78#_M1008_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.07455 AS=0.1113 PD=0.775 PS=1.37 NRD=16.4101 NRS=0 M=1
+ R=2.8 SA=75000.2 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1011 A_798_463# N_A_309_390#_M1011_g N_A_697_463#_M1008_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.07455 PD=0.63 PS=0.775 NRD=23.443 NRS=18.7544 M=1 R=2.8
+ SA=75000.7 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1010 N_VPWR_M1010_d N_A_839_359#_M1010_g A_798_463# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.13495 AS=0.0441 PD=1.14 PS=0.63 NRD=124.898 NRS=23.443 M=1 R=2.8
+ SA=75001.1 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1007 N_A_697_463#_M1007_d N_RESET_B_M1007_g N_VPWR_M1010_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1239 AS=0.13495 PD=1.43 PS=1.14 NRD=4.6886 NRS=124.898 M=1 R=2.8
+ SA=75001.7 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1028 N_A_839_359#_M1028_d N_A_697_463#_M1028_g N_VPWR_M1028_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.184062 AS=0.295 PD=1.43 PS=2.59 NRD=11.8003 NRS=1.9503 M=1
+ R=6.66667 SA=75000.2 SB=75001.5 A=0.15 P=2.3 MULT=1
MM1013 N_A_1271_74#_M1013_d N_A_309_390#_M1013_g N_A_839_359#_M1028_d VPB
+ PHIGHVT L=0.15 W=1 AD=0.319665 AS=0.184062 PD=2.57746 PS=1.43 NRD=10.8153
+ NRS=2.9353 M=1 R=6.66667 SA=75000.7 SB=75001.3 A=0.15 P=2.3 MULT=1
MM1002 A_1478_493# N_A_495_390#_M1002_g N_A_1271_74#_M1013_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0567 AS=0.13426 PD=0.69 PS=1.08254 NRD=37.5088 NRS=4.6886 M=1
+ R=2.8 SA=75001.3 SB=75002.4 A=0.063 P=1.14 MULT=1
MM1026 N_VPWR_M1026_d N_A_1525_212#_M1026_g A_1478_493# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0735 AS=0.0567 PD=0.77 PS=0.69 NRD=4.6886 NRS=37.5088 M=1 R=2.8
+ SA=75001.7 SB=75002 A=0.063 P=1.14 MULT=1
MM1000 N_A_1525_212#_M1000_d N_RESET_B_M1000_g N_VPWR_M1026_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1176 AS=0.0735 PD=0.98 PS=0.77 NRD=65.6601 NRS=28.1316 M=1 R=2.8
+ SA=75002.2 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1033 N_VPWR_M1033_d N_A_1271_74#_M1033_g N_A_1525_212#_M1000_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.1092 AS=0.1176 PD=0.85 PS=0.98 NRD=44.5417 NRS=65.6601 M=1
+ R=2.8 SA=75002.9 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1024 N_A_1921_409#_M1024_d N_A_1271_74#_M1024_g N_VPWR_M1033_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.2478 AS=0.2184 PD=2.27 PS=1.7 NRD=2.3443 NRS=14.0658 M=1
+ R=5.6 SA=75001.9 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1021 N_Q_M1021_d N_A_1921_409#_M1021_g N_VPWR_M1021_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.3584 PD=1.42 PS=2.88 NRD=1.7533 NRS=6.1464 M=1 R=7.46667
+ SA=75000.2 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1030 N_Q_M1021_d N_A_1921_409#_M1030_g N_VPWR_M1030_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75000.2 A=0.168 P=2.54 MULT=1
DX34_noxref VNB VPB NWDIODE A=22.4853 P=27.76
c_118 VNB 0 9.16943e-20 $X=0 $Y=0
c_242 VPB 0 1.1997e-19 $X=0 $Y=3.085
c_1745 A_1478_493# 0 1.15577e-19 $X=7.39 $Y=2.465
*
.include "sky130_fd_sc_ls__dfrtp_2.pxi.spice"
*
.ends
*
*
