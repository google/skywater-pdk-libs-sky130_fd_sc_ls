* File: sky130_fd_sc_ls__a21o_1.spice
* Created: Wed Sep  2 10:48:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__a21o_1.pex.spice"
.subckt sky130_fd_sc_ls__a21o_1  VNB VPB B1 A1 A2 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A2	A2
* A1	A1
* B1	B1
* VPB	VPB
* VNB	VNB
MM1001 N_VGND_M1001_d N_A_81_264#_M1001_g N_X_M1001_s VNB NSHORT L=0.15 W=0.74
+ AD=0.152558 AS=0.1961 PD=1.22261 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.5 A=0.111 P=1.78 MULT=1
MM1004 N_A_81_264#_M1004_d N_B1_M1004_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.131942 PD=0.92 PS=1.05739 NRD=0 NRS=22.488 M=1 R=4.26667
+ SA=75000.7 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1005 A_452_136# N_A1_M1005_g N_A_81_264#_M1004_d VNB NSHORT L=0.15 W=0.64
+ AD=0.104 AS=0.0896 PD=0.965 PS=0.92 NRD=20.148 NRS=0 M=1 R=4.26667 SA=75001.2
+ SB=75000.7 A=0.096 P=1.58 MULT=1
MM1003 N_VGND_M1003_d N_A2_M1003_g A_452_136# VNB NSHORT L=0.15 W=0.64 AD=0.1696
+ AS=0.104 PD=1.81 PS=0.965 NRD=0 NRS=20.148 M=1 R=4.26667 SA=75001.6 SB=75000.2
+ A=0.096 P=1.58 MULT=1
MM1007 N_VPWR_M1007_d N_A_81_264#_M1007_g N_X_M1007_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.308 AS=0.308 PD=2.79 PS=2.79 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1002 N_A_364_392#_M1002_d N_B1_M1002_g N_A_81_264#_M1002_s VPB PHIGHVT L=0.15
+ W=1 AD=0.15 AS=0.275 PD=1.3 PS=2.55 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75001.1 A=0.15 P=2.3 MULT=1
MM1006 N_VPWR_M1006_d N_A1_M1006_g N_A_364_392#_M1002_d VPB PHIGHVT L=0.15 W=1
+ AD=0.165 AS=0.15 PD=1.33 PS=1.3 NRD=4.9053 NRS=1.9503 M=1 R=6.66667 SA=75000.6
+ SB=75000.7 A=0.15 P=2.3 MULT=1
MM1000 N_A_364_392#_M1000_d N_A2_M1000_g N_VPWR_M1006_d VPB PHIGHVT L=0.15 W=1
+ AD=0.275 AS=0.165 PD=2.55 PS=1.33 NRD=1.9503 NRS=4.9053 M=1 R=6.66667
+ SA=75001.1 SB=75000.2 A=0.15 P=2.3 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.9564 P=11.2
c_33 VNB 0 1.84796e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_ls__a21o_1.pxi.spice"
*
.ends
*
*
