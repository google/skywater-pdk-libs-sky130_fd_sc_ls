* File: sky130_fd_sc_ls__and4bb_1.pxi.spice
* Created: Wed Sep  2 10:56:04 2020
* 
x_PM_SKY130_FD_SC_LS__AND4BB_1%A_N N_A_N_M1012_g N_A_N_c_98_n N_A_N_M1008_g A_N
+ N_A_N_c_99_n PM_SKY130_FD_SC_LS__AND4BB_1%A_N
x_PM_SKY130_FD_SC_LS__AND4BB_1%A_179_48# N_A_179_48#_M1004_s N_A_179_48#_M1009_d
+ N_A_179_48#_M1001_d N_A_179_48#_M1002_g N_A_179_48#_c_124_n
+ N_A_179_48#_M1011_g N_A_179_48#_c_125_n N_A_179_48#_c_126_n
+ N_A_179_48#_c_127_n N_A_179_48#_c_128_n N_A_179_48#_c_134_n
+ N_A_179_48#_c_135_n N_A_179_48#_c_136_n N_A_179_48#_c_129_n
+ N_A_179_48#_c_130_n N_A_179_48#_c_131_n N_A_179_48#_c_137_n
+ PM_SKY130_FD_SC_LS__AND4BB_1%A_179_48#
x_PM_SKY130_FD_SC_LS__AND4BB_1%A_27_74# N_A_27_74#_M1012_s N_A_27_74#_M1008_s
+ N_A_27_74#_c_228_n N_A_27_74#_M1009_g N_A_27_74#_M1004_g N_A_27_74#_c_230_n
+ N_A_27_74#_c_231_n N_A_27_74#_c_232_n N_A_27_74#_c_233_n N_A_27_74#_c_237_n
+ N_A_27_74#_c_234_n N_A_27_74#_c_239_n PM_SKY130_FD_SC_LS__AND4BB_1%A_27_74#
x_PM_SKY130_FD_SC_LS__AND4BB_1%A_503_48# N_A_503_48#_M1007_d N_A_503_48#_M1003_d
+ N_A_503_48#_M1005_g N_A_503_48#_c_318_n N_A_503_48#_c_319_n
+ N_A_503_48#_M1013_g N_A_503_48#_c_310_n N_A_503_48#_c_311_n
+ N_A_503_48#_c_312_n N_A_503_48#_c_313_n N_A_503_48#_c_314_n
+ N_A_503_48#_c_337_n N_A_503_48#_c_315_n N_A_503_48#_c_323_n
+ N_A_503_48#_c_324_n N_A_503_48#_c_316_n N_A_503_48#_c_317_n
+ PM_SKY130_FD_SC_LS__AND4BB_1%A_503_48#
x_PM_SKY130_FD_SC_LS__AND4BB_1%C N_C_M1010_g N_C_c_406_n N_C_M1001_g N_C_c_403_n
+ C N_C_c_404_n N_C_c_405_n PM_SKY130_FD_SC_LS__AND4BB_1%C
x_PM_SKY130_FD_SC_LS__AND4BB_1%D N_D_M1000_g N_D_c_446_n N_D_M1006_g N_D_c_443_n
+ D N_D_c_444_n N_D_c_445_n PM_SKY130_FD_SC_LS__AND4BB_1%D
x_PM_SKY130_FD_SC_LS__AND4BB_1%B_N N_B_N_c_485_n N_B_N_c_490_n N_B_N_M1003_g
+ N_B_N_M1007_g B_N N_B_N_c_487_n N_B_N_c_488_n PM_SKY130_FD_SC_LS__AND4BB_1%B_N
x_PM_SKY130_FD_SC_LS__AND4BB_1%VPWR N_VPWR_M1008_d N_VPWR_M1009_s N_VPWR_M1013_d
+ N_VPWR_M1006_d N_VPWR_c_519_n N_VPWR_c_520_n N_VPWR_c_521_n N_VPWR_c_522_n
+ N_VPWR_c_523_n N_VPWR_c_524_n N_VPWR_c_525_n N_VPWR_c_526_n N_VPWR_c_527_n
+ N_VPWR_c_528_n VPWR N_VPWR_c_529_n N_VPWR_c_518_n N_VPWR_c_531_n
+ PM_SKY130_FD_SC_LS__AND4BB_1%VPWR
x_PM_SKY130_FD_SC_LS__AND4BB_1%X N_X_M1002_d N_X_M1011_d N_X_c_582_n N_X_c_583_n
+ N_X_c_584_n N_X_c_588_n X N_X_c_586_n PM_SKY130_FD_SC_LS__AND4BB_1%X
x_PM_SKY130_FD_SC_LS__AND4BB_1%VGND N_VGND_M1012_d N_VGND_M1000_d N_VGND_c_617_n
+ N_VGND_c_618_n N_VGND_c_619_n N_VGND_c_620_n VGND N_VGND_c_621_n
+ N_VGND_c_622_n N_VGND_c_623_n N_VGND_c_624_n PM_SKY130_FD_SC_LS__AND4BB_1%VGND
cc_1 VNB N_A_N_M1012_g 0.0410018f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.645
cc_2 VNB N_A_N_c_98_n 0.0597667f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_3 VNB N_A_N_c_99_n 0.00427511f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_4 VNB N_A_179_48#_M1002_g 0.027508f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_5 VNB N_A_179_48#_c_124_n 0.0193298f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_A_179_48#_c_125_n 0.00566753f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_179_48#_c_126_n 0.0108078f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_179_48#_c_127_n 0.00552356f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_179_48#_c_128_n 0.00371726f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_179_48#_c_129_n 0.0429901f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_179_48#_c_130_n 0.00402396f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_179_48#_c_131_n 0.0156032f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_74#_c_228_n 0.0418726f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.26
cc_14 VNB N_A_27_74#_M1004_g 0.0304942f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_15 VNB N_A_27_74#_c_230_n 0.0252878f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_27_74#_c_231_n 0.00307298f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_27_74#_c_232_n 0.00912492f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_27_74#_c_233_n 0.00471389f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_27_74#_c_234_n 0.00288195f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_503_48#_c_310_n 0.0180921f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_503_48#_c_311_n 0.0233755f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_503_48#_c_312_n 0.0024279f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_503_48#_c_313_n 0.00106996f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_503_48#_c_314_n 0.0166374f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_503_48#_c_315_n 0.00741585f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_503_48#_c_316_n 0.0290446f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_503_48#_c_317_n 0.0184362f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_C_M1010_g 0.0235303f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.645
cc_29 VNB N_C_c_403_n 0.0187725f $X=-0.19 $Y=-0.245 $X2=0.35 $Y2=1.465
cc_30 VNB N_C_c_404_n 0.0152048f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_C_c_405_n 0.00452729f $X=-0.19 $Y=-0.245 $X2=0.252 $Y2=1.665
cc_32 VNB N_D_M1000_g 0.0243691f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.645
cc_33 VNB N_D_c_443_n 0.0191427f $X=-0.19 $Y=-0.245 $X2=0.35 $Y2=1.465
cc_34 VNB N_D_c_444_n 0.0153308f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_D_c_445_n 0.0035566f $X=-0.19 $Y=-0.245 $X2=0.252 $Y2=1.665
cc_36 VNB N_B_N_c_485_n 0.00151951f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.645
cc_37 VNB N_B_N_M1007_g 0.0394675f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_38 VNB N_B_N_c_487_n 0.0607038f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_B_N_c_488_n 0.00477584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VPWR_c_518_n 0.203486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_X_c_582_n 0.00354223f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_42 VNB N_X_c_583_n 0.00216891f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_43 VNB N_X_c_584_n 0.00202082f $X=-0.19 $Y=-0.245 $X2=0.252 $Y2=1.665
cc_44 VNB N_VGND_c_617_n 0.00647573f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_618_n 0.00961301f $X=-0.19 $Y=-0.245 $X2=0.252 $Y2=1.465
cc_46 VNB N_VGND_c_619_n 0.0844452f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_620_n 0.007312f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_621_n 0.0173909f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_622_n 0.0219533f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_623_n 0.295025f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_624_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VPB N_A_N_c_98_n 0.0277647f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_53 VPB N_A_N_c_99_n 0.00810654f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_54 VPB N_A_179_48#_c_124_n 0.0269547f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_A_179_48#_c_128_n 0.00312957f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_A_179_48#_c_134_n 0.00289722f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_A_179_48#_c_135_n 0.0139431f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_A_179_48#_c_136_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_A_179_48#_c_137_n 0.00606315f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_A_27_74#_c_228_n 0.0629782f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.26
cc_61 VPB N_A_27_74#_c_233_n 0.00110566f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_A_27_74#_c_237_n 0.0131844f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_A_27_74#_c_234_n 0.00538803f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_A_27_74#_c_239_n 0.0345873f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_A_503_48#_c_318_n 0.0098842f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_66 VPB N_A_503_48#_c_319_n 0.0226511f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_67 VPB N_A_503_48#_c_312_n 0.0132216f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_A_503_48#_c_313_n 0.00115078f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_A_503_48#_c_315_n 0.00242007f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_A_503_48#_c_323_n 0.0144694f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_A_503_48#_c_324_n 0.0360197f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_C_c_406_n 0.016008f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_73 VPB N_C_c_403_n 0.0285498f $X=-0.19 $Y=1.66 $X2=0.35 $Y2=1.465
cc_74 VPB N_C_c_405_n 0.00289358f $X=-0.19 $Y=1.66 $X2=0.252 $Y2=1.665
cc_75 VPB N_D_c_446_n 0.0165427f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_76 VPB N_D_c_443_n 0.0305808f $X=-0.19 $Y=1.66 $X2=0.35 $Y2=1.465
cc_77 VPB N_D_c_445_n 0.00194081f $X=-0.19 $Y=1.66 $X2=0.252 $Y2=1.665
cc_78 VPB N_B_N_c_485_n 0.0202878f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.645
cc_79 VPB N_B_N_c_490_n 0.0271315f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.645
cc_80 VPB N_B_N_c_488_n 0.00929358f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_519_n 0.0170949f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_520_n 0.0121322f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_521_n 0.00900305f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_522_n 0.00976973f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_523_n 0.0257133f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_524_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_525_n 0.0185368f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_526_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_527_n 0.0193312f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_528_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_529_n 0.0204244f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_518_n 0.0782942f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_531_n 0.0274851f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB N_X_c_582_n 0.00103408f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_95 VPB N_X_c_586_n 0.00653284f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 N_A_N_M1012_g N_A_179_48#_M1002_g 0.0215682f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_97 N_A_N_c_98_n N_A_179_48#_c_124_n 0.0435145f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_98 N_A_N_M1012_g N_A_27_74#_c_230_n 0.00509125f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_99 N_A_N_M1012_g N_A_27_74#_c_231_n 0.0197086f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_100 N_A_N_c_98_n N_A_27_74#_c_231_n 0.00103462f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_101 N_A_N_c_99_n N_A_27_74#_c_231_n 0.00260541f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_102 N_A_N_c_98_n N_A_27_74#_c_232_n 0.00197868f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_103 N_A_N_c_99_n N_A_27_74#_c_232_n 0.0217424f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_104 N_A_N_M1012_g N_A_27_74#_c_233_n 0.00443834f $X=0.495 $Y=0.645 $X2=0
+ $Y2=0
cc_105 N_A_N_c_98_n N_A_27_74#_c_233_n 0.0201799f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_106 N_A_N_c_99_n N_A_27_74#_c_233_n 0.0345406f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_107 N_A_N_c_98_n N_A_27_74#_c_239_n 0.0305969f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_108 N_A_N_c_99_n N_A_27_74#_c_239_n 0.0242922f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_109 N_A_N_c_98_n N_VPWR_c_519_n 0.00343137f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_110 N_A_N_c_98_n N_VPWR_c_518_n 0.00462577f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_111 N_A_N_c_98_n N_VPWR_c_531_n 0.00393265f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_112 N_A_N_c_98_n N_X_c_582_n 0.00102122f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_113 N_A_N_c_98_n N_X_c_588_n 2.90832e-19 $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_114 N_A_N_M1012_g N_VGND_c_617_n 0.0124836f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_115 N_A_N_M1012_g N_VGND_c_621_n 0.00383152f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_116 N_A_N_M1012_g N_VGND_c_623_n 0.00761198f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_117 N_A_179_48#_c_124_n N_A_27_74#_c_228_n 0.0047992f $X=1.04 $Y=1.765 $X2=0
+ $Y2=0
cc_118 N_A_179_48#_c_126_n N_A_27_74#_c_228_n 0.00121947f $X=1.82 $Y=0.945 $X2=0
+ $Y2=0
cc_119 N_A_179_48#_c_128_n N_A_27_74#_c_228_n 0.0181507f $X=2.3 $Y=2.03 $X2=0
+ $Y2=0
cc_120 N_A_179_48#_c_134_n N_A_27_74#_c_228_n 0.00421477f $X=2.46 $Y=2.265 $X2=0
+ $Y2=0
cc_121 N_A_179_48#_c_129_n N_A_27_74#_c_228_n 0.0213513f $X=1.38 $Y=1.465 $X2=0
+ $Y2=0
cc_122 N_A_179_48#_c_130_n N_A_27_74#_c_228_n 0.00207719f $X=1.525 $Y=1.465
+ $X2=0 $Y2=0
cc_123 N_A_179_48#_c_131_n N_A_27_74#_c_228_n 0.00516793f $X=1.985 $Y=0.515
+ $X2=0 $Y2=0
cc_124 N_A_179_48#_c_137_n N_A_27_74#_c_228_n 0.00701831f $X=2.42 $Y=2.115 $X2=0
+ $Y2=0
cc_125 N_A_179_48#_c_125_n N_A_27_74#_M1004_g 0.00398916f $X=1.525 $Y=1.3 $X2=0
+ $Y2=0
cc_126 N_A_179_48#_c_128_n N_A_27_74#_M1004_g 0.0074719f $X=2.3 $Y=2.03 $X2=0
+ $Y2=0
cc_127 N_A_179_48#_c_131_n N_A_27_74#_M1004_g 0.0201006f $X=1.985 $Y=0.515 $X2=0
+ $Y2=0
cc_128 N_A_179_48#_M1002_g N_A_27_74#_c_231_n 0.00122398f $X=0.97 $Y=0.74 $X2=0
+ $Y2=0
cc_129 N_A_179_48#_M1002_g N_A_27_74#_c_233_n 0.00215077f $X=0.97 $Y=0.74 $X2=0
+ $Y2=0
cc_130 N_A_179_48#_c_124_n N_A_27_74#_c_233_n 0.00151261f $X=1.04 $Y=1.765 $X2=0
+ $Y2=0
cc_131 N_A_179_48#_c_124_n N_A_27_74#_c_237_n 0.0142912f $X=1.04 $Y=1.765 $X2=0
+ $Y2=0
cc_132 N_A_179_48#_c_124_n N_A_27_74#_c_234_n 0.00527556f $X=1.04 $Y=1.765 $X2=0
+ $Y2=0
cc_133 N_A_179_48#_c_125_n N_A_27_74#_c_234_n 7.3914e-19 $X=1.525 $Y=1.3 $X2=0
+ $Y2=0
cc_134 N_A_179_48#_c_126_n N_A_27_74#_c_234_n 0.00226272f $X=1.82 $Y=0.945 $X2=0
+ $Y2=0
cc_135 N_A_179_48#_c_128_n N_A_27_74#_c_234_n 0.0521712f $X=2.3 $Y=2.03 $X2=0
+ $Y2=0
cc_136 N_A_179_48#_c_129_n N_A_27_74#_c_234_n 3.42035e-19 $X=1.38 $Y=1.465 $X2=0
+ $Y2=0
cc_137 N_A_179_48#_c_130_n N_A_27_74#_c_234_n 0.0258568f $X=1.525 $Y=1.465 $X2=0
+ $Y2=0
cc_138 N_A_179_48#_c_131_n N_A_27_74#_c_234_n 0.0144437f $X=1.985 $Y=0.515 $X2=0
+ $Y2=0
cc_139 N_A_179_48#_c_137_n N_A_27_74#_c_234_n 0.0138749f $X=2.42 $Y=2.115 $X2=0
+ $Y2=0
cc_140 N_A_179_48#_c_124_n N_A_27_74#_c_239_n 0.00576749f $X=1.04 $Y=1.765 $X2=0
+ $Y2=0
cc_141 N_A_179_48#_c_128_n N_A_503_48#_c_318_n 0.00411263f $X=2.3 $Y=2.03 $X2=0
+ $Y2=0
cc_142 N_A_179_48#_c_134_n N_A_503_48#_c_319_n 0.0114968f $X=2.46 $Y=2.265 $X2=0
+ $Y2=0
cc_143 N_A_179_48#_c_135_n N_A_503_48#_c_319_n 0.0133045f $X=3.295 $Y=2.115
+ $X2=0 $Y2=0
cc_144 N_A_179_48#_c_136_n N_A_503_48#_c_319_n 6.47235e-19 $X=3.46 $Y=2.265
+ $X2=0 $Y2=0
cc_145 N_A_179_48#_c_137_n N_A_503_48#_c_319_n 0.00236345f $X=2.42 $Y=2.115
+ $X2=0 $Y2=0
cc_146 N_A_179_48#_c_131_n N_A_503_48#_c_310_n 0.00961636f $X=1.985 $Y=0.515
+ $X2=0 $Y2=0
cc_147 N_A_179_48#_c_128_n N_A_503_48#_c_311_n 0.00961636f $X=2.3 $Y=2.03 $X2=0
+ $Y2=0
cc_148 N_A_179_48#_c_135_n N_A_503_48#_c_312_n 4.47545e-19 $X=3.295 $Y=2.115
+ $X2=0 $Y2=0
cc_149 N_A_179_48#_c_137_n N_A_503_48#_c_312_n 0.00213307f $X=2.42 $Y=2.115
+ $X2=0 $Y2=0
cc_150 N_A_179_48#_c_135_n N_A_503_48#_c_313_n 0.012887f $X=3.295 $Y=2.115 $X2=0
+ $Y2=0
cc_151 N_A_179_48#_c_131_n N_A_503_48#_c_313_n 0.0571916f $X=1.985 $Y=0.515
+ $X2=0 $Y2=0
cc_152 N_A_179_48#_c_137_n N_A_503_48#_c_313_n 0.00460395f $X=2.42 $Y=2.115
+ $X2=0 $Y2=0
cc_153 N_A_179_48#_c_131_n N_A_503_48#_c_337_n 0.0145967f $X=1.985 $Y=0.515
+ $X2=0 $Y2=0
cc_154 N_A_179_48#_c_135_n N_A_503_48#_c_323_n 0.00384588f $X=3.295 $Y=2.115
+ $X2=0 $Y2=0
cc_155 N_A_179_48#_c_134_n N_C_c_406_n 6.47235e-19 $X=2.46 $Y=2.265 $X2=0 $Y2=0
cc_156 N_A_179_48#_c_135_n N_C_c_406_n 0.0113102f $X=3.295 $Y=2.115 $X2=0 $Y2=0
cc_157 N_A_179_48#_c_136_n N_C_c_406_n 0.0115316f $X=3.46 $Y=2.265 $X2=0 $Y2=0
cc_158 N_A_179_48#_c_135_n N_C_c_403_n 0.00646084f $X=3.295 $Y=2.115 $X2=0 $Y2=0
cc_159 N_A_179_48#_c_128_n N_C_c_405_n 0.0022031f $X=2.3 $Y=2.03 $X2=0 $Y2=0
cc_160 N_A_179_48#_c_135_n N_C_c_405_n 0.0260806f $X=3.295 $Y=2.115 $X2=0 $Y2=0
cc_161 N_A_179_48#_c_135_n N_D_c_446_n 0.00377778f $X=3.295 $Y=2.115 $X2=0 $Y2=0
cc_162 N_A_179_48#_c_136_n N_D_c_446_n 0.0110868f $X=3.46 $Y=2.265 $X2=0 $Y2=0
cc_163 N_A_179_48#_c_135_n N_D_c_443_n 0.00124348f $X=3.295 $Y=2.115 $X2=0 $Y2=0
cc_164 N_A_179_48#_c_135_n N_D_c_445_n 0.00997848f $X=3.295 $Y=2.115 $X2=0 $Y2=0
cc_165 N_A_179_48#_c_135_n N_B_N_c_490_n 4.40222e-19 $X=3.295 $Y=2.115 $X2=0
+ $Y2=0
cc_166 N_A_179_48#_c_136_n N_B_N_c_490_n 5.50696e-19 $X=3.46 $Y=2.265 $X2=0
+ $Y2=0
cc_167 N_A_179_48#_c_135_n N_VPWR_M1013_d 0.00308396f $X=3.295 $Y=2.115 $X2=0
+ $Y2=0
cc_168 N_A_179_48#_c_124_n N_VPWR_c_519_n 0.0212893f $X=1.04 $Y=1.765 $X2=0
+ $Y2=0
cc_169 N_A_179_48#_c_124_n N_VPWR_c_520_n 0.0093841f $X=1.04 $Y=1.765 $X2=0
+ $Y2=0
cc_170 N_A_179_48#_c_134_n N_VPWR_c_520_n 0.0127976f $X=2.46 $Y=2.265 $X2=0
+ $Y2=0
cc_171 N_A_179_48#_c_134_n N_VPWR_c_521_n 0.0236791f $X=2.46 $Y=2.265 $X2=0
+ $Y2=0
cc_172 N_A_179_48#_c_135_n N_VPWR_c_521_n 0.0232685f $X=3.295 $Y=2.115 $X2=0
+ $Y2=0
cc_173 N_A_179_48#_c_136_n N_VPWR_c_521_n 0.0236791f $X=3.46 $Y=2.265 $X2=0
+ $Y2=0
cc_174 N_A_179_48#_c_136_n N_VPWR_c_522_n 0.0244142f $X=3.46 $Y=2.265 $X2=0
+ $Y2=0
cc_175 N_A_179_48#_c_124_n N_VPWR_c_523_n 0.00413917f $X=1.04 $Y=1.765 $X2=0
+ $Y2=0
cc_176 N_A_179_48#_c_134_n N_VPWR_c_525_n 0.0145938f $X=2.46 $Y=2.265 $X2=0
+ $Y2=0
cc_177 N_A_179_48#_c_136_n N_VPWR_c_527_n 0.014552f $X=3.46 $Y=2.265 $X2=0 $Y2=0
cc_178 N_A_179_48#_c_124_n N_VPWR_c_518_n 0.00419307f $X=1.04 $Y=1.765 $X2=0
+ $Y2=0
cc_179 N_A_179_48#_c_134_n N_VPWR_c_518_n 0.0120466f $X=2.46 $Y=2.265 $X2=0
+ $Y2=0
cc_180 N_A_179_48#_c_136_n N_VPWR_c_518_n 0.0119791f $X=3.46 $Y=2.265 $X2=0
+ $Y2=0
cc_181 N_A_179_48#_M1002_g N_X_c_582_n 0.00581287f $X=0.97 $Y=0.74 $X2=0 $Y2=0
cc_182 N_A_179_48#_c_124_n N_X_c_582_n 0.0193255f $X=1.04 $Y=1.765 $X2=0 $Y2=0
cc_183 N_A_179_48#_c_125_n N_X_c_582_n 0.00761824f $X=1.525 $Y=1.3 $X2=0 $Y2=0
cc_184 N_A_179_48#_c_130_n N_X_c_582_n 0.023711f $X=1.525 $Y=1.465 $X2=0 $Y2=0
cc_185 N_A_179_48#_M1002_g N_X_c_583_n 0.00163355f $X=0.97 $Y=0.74 $X2=0 $Y2=0
cc_186 N_A_179_48#_c_127_n N_X_c_583_n 0.00798712f $X=1.61 $Y=0.945 $X2=0 $Y2=0
cc_187 N_A_179_48#_c_131_n N_X_c_583_n 0.0181191f $X=1.985 $Y=0.515 $X2=0 $Y2=0
cc_188 N_A_179_48#_M1002_g N_X_c_584_n 0.0096135f $X=0.97 $Y=0.74 $X2=0 $Y2=0
cc_189 N_A_179_48#_c_124_n N_X_c_584_n 0.0071813f $X=1.04 $Y=1.765 $X2=0 $Y2=0
cc_190 N_A_179_48#_c_125_n N_X_c_584_n 0.00777787f $X=1.525 $Y=1.3 $X2=0 $Y2=0
cc_191 N_A_179_48#_c_127_n N_X_c_584_n 0.0057961f $X=1.61 $Y=0.945 $X2=0 $Y2=0
cc_192 N_A_179_48#_c_130_n N_X_c_584_n 0.00150313f $X=1.525 $Y=1.465 $X2=0 $Y2=0
cc_193 N_A_179_48#_c_124_n N_X_c_588_n 0.00751788f $X=1.04 $Y=1.765 $X2=0 $Y2=0
cc_194 N_A_179_48#_c_124_n N_X_c_586_n 0.0104764f $X=1.04 $Y=1.765 $X2=0 $Y2=0
cc_195 N_A_179_48#_c_129_n N_X_c_586_n 0.01137f $X=1.38 $Y=1.465 $X2=0 $Y2=0
cc_196 N_A_179_48#_c_130_n N_X_c_586_n 0.0230181f $X=1.525 $Y=1.465 $X2=0 $Y2=0
cc_197 N_A_179_48#_M1002_g N_VGND_c_617_n 0.00364992f $X=0.97 $Y=0.74 $X2=0
+ $Y2=0
cc_198 N_A_179_48#_M1002_g N_VGND_c_619_n 0.00461464f $X=0.97 $Y=0.74 $X2=0
+ $Y2=0
cc_199 N_A_179_48#_c_131_n N_VGND_c_619_n 0.0246732f $X=1.985 $Y=0.515 $X2=0
+ $Y2=0
cc_200 N_A_179_48#_M1002_g N_VGND_c_623_n 0.00913048f $X=0.97 $Y=0.74 $X2=0
+ $Y2=0
cc_201 N_A_179_48#_c_126_n N_VGND_c_623_n 0.00711624f $X=1.82 $Y=0.945 $X2=0
+ $Y2=0
cc_202 N_A_179_48#_c_127_n N_VGND_c_623_n 0.00631461f $X=1.61 $Y=0.945 $X2=0
+ $Y2=0
cc_203 N_A_179_48#_c_131_n N_VGND_c_623_n 0.02007f $X=1.985 $Y=0.515 $X2=0 $Y2=0
cc_204 N_A_179_48#_c_131_n A_455_74# 0.00765047f $X=1.985 $Y=0.515 $X2=-0.19
+ $Y2=-0.245
cc_205 N_A_27_74#_c_228_n N_A_503_48#_c_318_n 0.00888341f $X=2.185 $Y=2.045
+ $X2=0 $Y2=0
cc_206 N_A_27_74#_c_228_n N_A_503_48#_c_319_n 0.0201462f $X=2.185 $Y=2.045 $X2=0
+ $Y2=0
cc_207 N_A_27_74#_M1004_g N_A_503_48#_c_310_n 0.0397166f $X=2.2 $Y=0.69 $X2=0
+ $Y2=0
cc_208 N_A_27_74#_c_228_n N_A_503_48#_c_311_n 0.0397166f $X=2.185 $Y=2.045 $X2=0
+ $Y2=0
cc_209 N_A_27_74#_M1004_g N_A_503_48#_c_313_n 7.44855e-19 $X=2.2 $Y=0.69 $X2=0
+ $Y2=0
cc_210 N_A_27_74#_c_233_n N_VPWR_M1008_d 9.28557e-19 $X=0.655 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_211 N_A_27_74#_c_237_n N_VPWR_M1008_d 0.00835563f $X=1.78 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_212 N_A_27_74#_c_239_n N_VPWR_M1008_d 0.00546216f $X=0.28 $Y=2.115 $X2=-0.19
+ $Y2=-0.245
cc_213 N_A_27_74#_c_237_n N_VPWR_M1009_s 0.00624981f $X=1.78 $Y=2.405 $X2=0
+ $Y2=0
cc_214 N_A_27_74#_c_234_n N_VPWR_M1009_s 0.00398414f $X=1.92 $Y=1.455 $X2=0
+ $Y2=0
cc_215 N_A_27_74#_c_237_n N_VPWR_c_519_n 0.0143351f $X=1.78 $Y=2.405 $X2=0 $Y2=0
cc_216 N_A_27_74#_c_239_n N_VPWR_c_519_n 0.0105191f $X=0.28 $Y=2.115 $X2=0 $Y2=0
cc_217 N_A_27_74#_c_228_n N_VPWR_c_520_n 0.0102595f $X=2.185 $Y=2.045 $X2=0
+ $Y2=0
cc_218 N_A_27_74#_c_237_n N_VPWR_c_520_n 0.021932f $X=1.78 $Y=2.405 $X2=0 $Y2=0
cc_219 N_A_27_74#_c_228_n N_VPWR_c_525_n 0.00413917f $X=2.185 $Y=2.045 $X2=0
+ $Y2=0
cc_220 N_A_27_74#_c_228_n N_VPWR_c_518_n 0.00818241f $X=2.185 $Y=2.045 $X2=0
+ $Y2=0
cc_221 N_A_27_74#_c_237_n N_VPWR_c_518_n 0.0289854f $X=1.78 $Y=2.405 $X2=0 $Y2=0
cc_222 N_A_27_74#_c_239_n N_VPWR_c_518_n 0.0178324f $X=0.28 $Y=2.115 $X2=0 $Y2=0
cc_223 N_A_27_74#_c_239_n N_VPWR_c_531_n 0.00671799f $X=0.28 $Y=2.115 $X2=0
+ $Y2=0
cc_224 N_A_27_74#_c_237_n N_X_M1011_d 0.0135333f $X=1.78 $Y=2.405 $X2=0 $Y2=0
cc_225 N_A_27_74#_c_228_n N_X_c_582_n 0.00109827f $X=2.185 $Y=2.045 $X2=0 $Y2=0
cc_226 N_A_27_74#_c_233_n N_X_c_582_n 0.0506332f $X=0.655 $Y=1.95 $X2=0 $Y2=0
cc_227 N_A_27_74#_c_231_n N_X_c_584_n 0.0139665f $X=0.57 $Y=1.045 $X2=0 $Y2=0
cc_228 N_A_27_74#_c_233_n N_X_c_588_n 0.00561338f $X=0.655 $Y=1.95 $X2=0 $Y2=0
cc_229 N_A_27_74#_c_237_n N_X_c_588_n 0.00871803f $X=1.78 $Y=2.405 $X2=0 $Y2=0
cc_230 N_A_27_74#_c_228_n N_X_c_586_n 0.00168619f $X=2.185 $Y=2.045 $X2=0 $Y2=0
cc_231 N_A_27_74#_c_237_n N_X_c_586_n 0.032553f $X=1.78 $Y=2.405 $X2=0 $Y2=0
cc_232 N_A_27_74#_c_234_n N_X_c_586_n 0.0235675f $X=1.92 $Y=1.455 $X2=0 $Y2=0
cc_233 N_A_27_74#_c_231_n N_VGND_M1012_d 0.00233685f $X=0.57 $Y=1.045 $X2=-0.19
+ $Y2=-0.245
cc_234 N_A_27_74#_c_230_n N_VGND_c_617_n 0.0164982f $X=0.28 $Y=0.645 $X2=0 $Y2=0
cc_235 N_A_27_74#_c_231_n N_VGND_c_617_n 0.0146425f $X=0.57 $Y=1.045 $X2=0 $Y2=0
cc_236 N_A_27_74#_M1004_g N_VGND_c_619_n 0.00291513f $X=2.2 $Y=0.69 $X2=0 $Y2=0
cc_237 N_A_27_74#_c_230_n N_VGND_c_621_n 0.011066f $X=0.28 $Y=0.645 $X2=0 $Y2=0
cc_238 N_A_27_74#_M1004_g N_VGND_c_623_n 0.00363725f $X=2.2 $Y=0.69 $X2=0 $Y2=0
cc_239 N_A_27_74#_c_230_n N_VGND_c_623_n 0.00915947f $X=0.28 $Y=0.645 $X2=0
+ $Y2=0
cc_240 N_A_503_48#_c_310_n N_C_M1010_g 0.0281202f $X=2.68 $Y=1.12 $X2=0 $Y2=0
cc_241 N_A_503_48#_c_313_n N_C_M1010_g 0.00266937f $X=2.68 $Y=1.285 $X2=0 $Y2=0
cc_242 N_A_503_48#_c_314_n N_C_M1010_g 0.00388845f $X=2.68 $Y=1.285 $X2=0 $Y2=0
cc_243 N_A_503_48#_c_317_n N_C_M1010_g 0.0129618f $X=4.06 $Y=0.94 $X2=0 $Y2=0
cc_244 N_A_503_48#_c_319_n N_C_c_406_n 0.023586f $X=2.685 $Y=2.045 $X2=0 $Y2=0
cc_245 N_A_503_48#_c_318_n N_C_c_403_n 0.0102658f $X=2.685 $Y=1.955 $X2=0 $Y2=0
cc_246 N_A_503_48#_c_311_n N_C_c_403_n 0.0186915f $X=2.68 $Y=1.625 $X2=0 $Y2=0
cc_247 N_A_503_48#_c_313_n N_C_c_404_n 6.90861e-19 $X=2.68 $Y=1.285 $X2=0 $Y2=0
cc_248 N_A_503_48#_c_314_n N_C_c_404_n 0.0186915f $X=2.68 $Y=1.285 $X2=0 $Y2=0
cc_249 N_A_503_48#_c_317_n N_C_c_404_n 0.00265283f $X=4.06 $Y=0.94 $X2=0 $Y2=0
cc_250 N_A_503_48#_c_318_n N_C_c_405_n 6.97875e-19 $X=2.685 $Y=1.955 $X2=0 $Y2=0
cc_251 N_A_503_48#_c_313_n N_C_c_405_n 0.0469689f $X=2.68 $Y=1.285 $X2=0 $Y2=0
cc_252 N_A_503_48#_c_314_n N_C_c_405_n 0.00337482f $X=2.68 $Y=1.285 $X2=0 $Y2=0
cc_253 N_A_503_48#_c_317_n N_C_c_405_n 0.0257971f $X=4.06 $Y=0.94 $X2=0 $Y2=0
cc_254 N_A_503_48#_c_315_n N_D_M1000_g 0.00303034f $X=4.145 $Y=1.95 $X2=0 $Y2=0
cc_255 N_A_503_48#_c_316_n N_D_M1000_g 0.001133f $X=4.52 $Y=0.85 $X2=0 $Y2=0
cc_256 N_A_503_48#_c_317_n N_D_M1000_g 0.0129805f $X=4.06 $Y=0.94 $X2=0 $Y2=0
cc_257 N_A_503_48#_c_323_n N_D_c_446_n 6.62548e-19 $X=4.48 $Y=2.12 $X2=0 $Y2=0
cc_258 N_A_503_48#_c_324_n N_D_c_446_n 8.97107e-19 $X=4.48 $Y=2.265 $X2=0 $Y2=0
cc_259 N_A_503_48#_c_315_n N_D_c_443_n 0.00171772f $X=4.145 $Y=1.95 $X2=0 $Y2=0
cc_260 N_A_503_48#_c_323_n N_D_c_443_n 0.00204631f $X=4.48 $Y=2.12 $X2=0 $Y2=0
cc_261 N_A_503_48#_c_315_n N_D_c_444_n 0.00418923f $X=4.145 $Y=1.95 $X2=0 $Y2=0
cc_262 N_A_503_48#_c_317_n N_D_c_444_n 0.00521595f $X=4.06 $Y=0.94 $X2=0 $Y2=0
cc_263 N_A_503_48#_c_315_n N_D_c_445_n 0.050868f $X=4.145 $Y=1.95 $X2=0 $Y2=0
cc_264 N_A_503_48#_c_317_n N_D_c_445_n 0.0295937f $X=4.06 $Y=0.94 $X2=0 $Y2=0
cc_265 N_A_503_48#_c_315_n N_B_N_c_485_n 0.0117678f $X=4.145 $Y=1.95 $X2=0 $Y2=0
cc_266 N_A_503_48#_c_323_n N_B_N_c_485_n 0.00538323f $X=4.48 $Y=2.12 $X2=0 $Y2=0
cc_267 N_A_503_48#_c_323_n N_B_N_c_490_n 0.0138437f $X=4.48 $Y=2.12 $X2=0 $Y2=0
cc_268 N_A_503_48#_c_324_n N_B_N_c_490_n 0.0138153f $X=4.48 $Y=2.265 $X2=0 $Y2=0
cc_269 N_A_503_48#_c_315_n N_B_N_M1007_g 0.00739013f $X=4.145 $Y=1.95 $X2=0
+ $Y2=0
cc_270 N_A_503_48#_c_316_n N_B_N_M1007_g 0.0261445f $X=4.52 $Y=0.85 $X2=0 $Y2=0
cc_271 N_A_503_48#_c_315_n N_B_N_c_487_n 0.00949279f $X=4.145 $Y=1.95 $X2=0
+ $Y2=0
cc_272 N_A_503_48#_c_323_n N_B_N_c_487_n 0.0031002f $X=4.48 $Y=2.12 $X2=0 $Y2=0
cc_273 N_A_503_48#_c_316_n N_B_N_c_487_n 0.00276952f $X=4.52 $Y=0.85 $X2=0 $Y2=0
cc_274 N_A_503_48#_c_315_n N_B_N_c_488_n 0.0345409f $X=4.145 $Y=1.95 $X2=0 $Y2=0
cc_275 N_A_503_48#_c_323_n N_B_N_c_488_n 0.0200264f $X=4.48 $Y=2.12 $X2=0 $Y2=0
cc_276 N_A_503_48#_c_316_n N_B_N_c_488_n 0.0156602f $X=4.52 $Y=0.85 $X2=0 $Y2=0
cc_277 N_A_503_48#_c_319_n N_VPWR_c_520_n 4.22589e-19 $X=2.685 $Y=2.045 $X2=0
+ $Y2=0
cc_278 N_A_503_48#_c_319_n N_VPWR_c_521_n 0.00551009f $X=2.685 $Y=2.045 $X2=0
+ $Y2=0
cc_279 N_A_503_48#_c_323_n N_VPWR_c_522_n 0.00596561f $X=4.48 $Y=2.12 $X2=0
+ $Y2=0
cc_280 N_A_503_48#_c_324_n N_VPWR_c_522_n 0.0266809f $X=4.48 $Y=2.265 $X2=0
+ $Y2=0
cc_281 N_A_503_48#_c_319_n N_VPWR_c_525_n 0.00445602f $X=2.685 $Y=2.045 $X2=0
+ $Y2=0
cc_282 N_A_503_48#_c_324_n N_VPWR_c_529_n 0.0145938f $X=4.48 $Y=2.265 $X2=0
+ $Y2=0
cc_283 N_A_503_48#_c_319_n N_VPWR_c_518_n 0.00858339f $X=2.685 $Y=2.045 $X2=0
+ $Y2=0
cc_284 N_A_503_48#_c_324_n N_VPWR_c_518_n 0.0120466f $X=4.48 $Y=2.265 $X2=0
+ $Y2=0
cc_285 N_A_503_48#_c_316_n N_VGND_M1000_d 0.00182175f $X=4.52 $Y=0.85 $X2=0
+ $Y2=0
cc_286 N_A_503_48#_c_317_n N_VGND_M1000_d 0.00379698f $X=4.06 $Y=0.94 $X2=0
+ $Y2=0
cc_287 N_A_503_48#_c_316_n N_VGND_c_618_n 0.0142603f $X=4.52 $Y=0.85 $X2=0 $Y2=0
cc_288 N_A_503_48#_c_317_n N_VGND_c_618_n 0.0262201f $X=4.06 $Y=0.94 $X2=0 $Y2=0
cc_289 N_A_503_48#_c_310_n N_VGND_c_619_n 0.00461464f $X=2.68 $Y=1.12 $X2=0
+ $Y2=0
cc_290 N_A_503_48#_c_316_n N_VGND_c_622_n 0.0102877f $X=4.52 $Y=0.85 $X2=0 $Y2=0
cc_291 N_A_503_48#_c_310_n N_VGND_c_623_n 0.00585788f $X=2.68 $Y=1.12 $X2=0
+ $Y2=0
cc_292 N_A_503_48#_c_337_n N_VGND_c_623_n 0.0104896f $X=2.845 $Y=0.935 $X2=0
+ $Y2=0
cc_293 N_A_503_48#_c_316_n N_VGND_c_623_n 0.0193098f $X=4.52 $Y=0.85 $X2=0 $Y2=0
cc_294 N_A_503_48#_c_317_n N_VGND_c_623_n 0.029238f $X=4.06 $Y=0.94 $X2=0 $Y2=0
cc_295 N_A_503_48#_c_337_n A_533_74# 0.00294599f $X=2.845 $Y=0.935 $X2=-0.19
+ $Y2=-0.245
cc_296 N_A_503_48#_c_317_n A_533_74# 0.00398078f $X=4.06 $Y=0.94 $X2=-0.19
+ $Y2=-0.245
cc_297 N_A_503_48#_c_317_n A_647_74# 0.00498776f $X=4.06 $Y=0.94 $X2=-0.19
+ $Y2=-0.245
cc_298 N_C_M1010_g N_D_M1000_g 0.034747f $X=3.16 $Y=0.69 $X2=0 $Y2=0
cc_299 N_C_c_406_n N_D_c_446_n 0.0147471f $X=3.235 $Y=2.045 $X2=0 $Y2=0
cc_300 N_C_c_403_n N_D_c_443_n 0.0306548f $X=3.22 $Y=1.695 $X2=0 $Y2=0
cc_301 N_C_c_404_n N_D_c_444_n 0.020772f $X=3.22 $Y=1.355 $X2=0 $Y2=0
cc_302 N_C_c_405_n N_D_c_444_n 6.62791e-19 $X=3.22 $Y=1.355 $X2=0 $Y2=0
cc_303 N_C_c_404_n N_D_c_445_n 0.00412737f $X=3.22 $Y=1.355 $X2=0 $Y2=0
cc_304 N_C_c_405_n N_D_c_445_n 0.0535897f $X=3.22 $Y=1.355 $X2=0 $Y2=0
cc_305 N_C_c_406_n N_VPWR_c_521_n 0.00689824f $X=3.235 $Y=2.045 $X2=0 $Y2=0
cc_306 N_C_c_406_n N_VPWR_c_527_n 0.00445602f $X=3.235 $Y=2.045 $X2=0 $Y2=0
cc_307 N_C_c_406_n N_VPWR_c_518_n 0.00857909f $X=3.235 $Y=2.045 $X2=0 $Y2=0
cc_308 N_C_M1010_g N_VGND_c_618_n 0.00207664f $X=3.16 $Y=0.69 $X2=0 $Y2=0
cc_309 N_C_M1010_g N_VGND_c_619_n 0.00461464f $X=3.16 $Y=0.69 $X2=0 $Y2=0
cc_310 N_C_M1010_g N_VGND_c_623_n 0.00469123f $X=3.16 $Y=0.69 $X2=0 $Y2=0
cc_311 N_D_c_443_n N_B_N_c_485_n 0.0195515f $X=3.76 $Y=1.695 $X2=0 $Y2=0
cc_312 N_D_c_446_n N_B_N_c_490_n 0.0212652f $X=3.685 $Y=2.045 $X2=0 $Y2=0
cc_313 N_D_M1000_g N_B_N_M1007_g 0.0168987f $X=3.67 $Y=0.69 $X2=0 $Y2=0
cc_314 N_D_c_444_n N_B_N_M1007_g 0.00363085f $X=3.76 $Y=1.355 $X2=0 $Y2=0
cc_315 N_D_c_444_n N_B_N_c_487_n 0.0146356f $X=3.76 $Y=1.355 $X2=0 $Y2=0
cc_316 N_D_c_445_n N_B_N_c_487_n 5.47444e-19 $X=3.76 $Y=1.355 $X2=0 $Y2=0
cc_317 N_D_c_446_n N_VPWR_c_522_n 0.00732073f $X=3.685 $Y=2.045 $X2=0 $Y2=0
cc_318 N_D_c_443_n N_VPWR_c_522_n 0.00293286f $X=3.76 $Y=1.695 $X2=0 $Y2=0
cc_319 N_D_c_445_n N_VPWR_c_522_n 0.00311272f $X=3.76 $Y=1.355 $X2=0 $Y2=0
cc_320 N_D_c_446_n N_VPWR_c_527_n 0.00445602f $X=3.685 $Y=2.045 $X2=0 $Y2=0
cc_321 N_D_c_446_n N_VPWR_c_518_n 0.00858504f $X=3.685 $Y=2.045 $X2=0 $Y2=0
cc_322 N_D_M1000_g N_VGND_c_618_n 0.0168272f $X=3.67 $Y=0.69 $X2=0 $Y2=0
cc_323 N_D_M1000_g N_VGND_c_619_n 0.00383152f $X=3.67 $Y=0.69 $X2=0 $Y2=0
cc_324 N_D_M1000_g N_VGND_c_623_n 0.00386851f $X=3.67 $Y=0.69 $X2=0 $Y2=0
cc_325 N_B_N_c_490_n N_VPWR_c_522_n 0.0075701f $X=4.255 $Y=2.045 $X2=0 $Y2=0
cc_326 N_B_N_c_490_n N_VPWR_c_529_n 0.00445602f $X=4.255 $Y=2.045 $X2=0 $Y2=0
cc_327 N_B_N_c_490_n N_VPWR_c_518_n 0.00861592f $X=4.255 $Y=2.045 $X2=0 $Y2=0
cc_328 N_B_N_M1007_g N_VGND_c_618_n 0.00548248f $X=4.305 $Y=0.735 $X2=0 $Y2=0
cc_329 N_B_N_M1007_g N_VGND_c_622_n 0.00491683f $X=4.305 $Y=0.735 $X2=0 $Y2=0
cc_330 N_B_N_M1007_g N_VGND_c_623_n 0.00517496f $X=4.305 $Y=0.735 $X2=0 $Y2=0
cc_331 N_X_c_583_n N_VGND_c_617_n 0.00133028f $X=1.185 $Y=0.515 $X2=0 $Y2=0
cc_332 N_X_c_583_n N_VGND_c_619_n 0.00832263f $X=1.185 $Y=0.515 $X2=0 $Y2=0
cc_333 N_X_c_583_n N_VGND_c_623_n 0.00691792f $X=1.185 $Y=0.515 $X2=0 $Y2=0
