# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ls__dlrtn_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ls__dlrtn_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.600000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.208500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 1.450000 0.805000 1.780000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  1.198400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.545000 1.960000 9.475000 1.970000 ;
        RECT 7.545000 1.970000 8.875000 2.130000 ;
        RECT 7.545000 2.130000 7.875000 2.980000 ;
        RECT 7.935000 0.360000 8.125000 0.960000 ;
        RECT 7.935000 0.960000 9.475000 1.130000 ;
        RECT 8.545000 1.800000 9.475000 1.960000 ;
        RECT 8.545000 2.130000 8.875000 2.980000 ;
        RECT 8.795000 0.360000 8.985000 0.800000 ;
        RECT 8.795000 0.800000 9.475000 0.960000 ;
        RECT 9.245000 1.130000 9.475000 1.800000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.444000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.320000 1.120000 7.555000 1.450000 ;
    END
  END RESET_B
  PIN GATE_N
    ANTENNAGATEAREA  0.237000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.975000 1.450000 1.290000 1.780000 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 9.600000 0.085000 ;
        RECT 0.625000  0.085000 0.955000 0.490000 ;
        RECT 2.310000  0.085000 3.125000 0.490000 ;
        RECT 4.595000  0.085000 4.925000 0.680000 ;
        RECT 6.445000  0.085000 6.775000 0.600000 ;
        RECT 7.435000  0.085000 7.765000 0.950000 ;
        RECT 8.295000  0.085000 8.625000 0.790000 ;
        RECT 9.155000  0.085000 9.485000 0.630000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
        RECT 6.395000 -0.085000 6.565000 0.085000 ;
        RECT 6.875000 -0.085000 7.045000 0.085000 ;
        RECT 7.355000 -0.085000 7.525000 0.085000 ;
        RECT 7.835000 -0.085000 8.005000 0.085000 ;
        RECT 8.315000 -0.085000 8.485000 0.085000 ;
        RECT 8.795000 -0.085000 8.965000 0.085000 ;
        RECT 9.275000 -0.085000 9.445000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 9.600000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 9.600000 3.415000 ;
        RECT 0.645000 1.950000 0.975000 3.245000 ;
        RECT 2.255000 2.940000 2.585000 3.245000 ;
        RECT 4.590000 2.630000 5.320000 3.245000 ;
        RECT 5.990000 2.080000 6.320000 3.245000 ;
        RECT 7.045000 2.080000 7.375000 3.245000 ;
        RECT 8.045000 2.300000 8.375000 3.245000 ;
        RECT 9.045000 2.140000 9.375000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
        RECT 6.395000 3.245000 6.565000 3.415000 ;
        RECT 6.875000 3.245000 7.045000 3.415000 ;
        RECT 7.355000 3.245000 7.525000 3.415000 ;
        RECT 7.835000 3.245000 8.005000 3.415000 ;
        RECT 8.315000 3.245000 8.485000 3.415000 ;
        RECT 8.795000 3.245000 8.965000 3.415000 ;
        RECT 9.275000 3.245000 9.445000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 9.600000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085000 0.660000 2.820000 0.830000 ;
      RECT 0.085000 0.830000 0.445000 1.250000 ;
      RECT 0.085000 1.250000 0.255000 1.950000 ;
      RECT 0.085000 1.950000 0.475000 2.830000 ;
      RECT 1.135000 1.000000 1.630000 1.250000 ;
      RECT 1.145000 1.950000 1.630000 2.600000 ;
      RECT 1.145000 2.600000 4.200000 2.770000 ;
      RECT 1.145000 2.770000 1.630000 2.830000 ;
      RECT 1.460000 1.250000 1.630000 1.420000 ;
      RECT 1.460000 1.420000 1.865000 1.750000 ;
      RECT 1.460000 1.750000 1.630000 1.950000 ;
      RECT 1.800000 1.000000 2.205000 1.250000 ;
      RECT 1.800000 1.920000 3.360000 2.090000 ;
      RECT 1.800000 2.090000 2.205000 2.430000 ;
      RECT 2.035000 1.250000 2.205000 1.920000 ;
      RECT 2.490000 0.830000 2.820000 1.670000 ;
      RECT 3.030000 1.190000 4.260000 1.520000 ;
      RECT 3.030000 1.520000 3.360000 1.920000 ;
      RECT 3.180000 2.260000 3.700000 2.430000 ;
      RECT 3.530000 1.690000 5.220000 1.860000 ;
      RECT 3.530000 1.860000 3.700000 2.260000 ;
      RECT 3.740000 0.400000 4.070000 0.850000 ;
      RECT 3.740000 0.850000 4.985000 1.020000 ;
      RECT 3.870000 2.030000 4.200000 2.600000 ;
      RECT 4.440000 2.030000 5.820000 2.360000 ;
      RECT 4.815000 1.020000 4.985000 1.120000 ;
      RECT 4.815000 1.120000 5.220000 1.690000 ;
      RECT 5.155000 0.255000 6.265000 0.425000 ;
      RECT 5.155000 0.425000 5.485000 0.950000 ;
      RECT 5.490000 1.620000 9.075000 1.630000 ;
      RECT 5.490000 1.630000 7.895000 1.790000 ;
      RECT 5.490000 1.790000 5.820000 2.030000 ;
      RECT 5.490000 2.360000 5.820000 2.960000 ;
      RECT 5.665000 0.595000 5.835000 1.620000 ;
      RECT 6.015000 0.425000 6.265000 0.770000 ;
      RECT 6.015000 0.770000 7.205000 0.950000 ;
      RECT 6.490000 1.790000 6.820000 2.960000 ;
      RECT 6.945000 0.355000 7.205000 0.770000 ;
      RECT 7.725000 1.300000 9.075000 1.620000 ;
  END
END sky130_fd_sc_ls__dlrtn_4
