* File: sky130_fd_sc_ls__o31a_2.pxi.spice
* Created: Fri Aug 28 13:52:50 2020
* 
x_PM_SKY130_FD_SC_LS__O31A_2%A_55_264# N_A_55_264#_M1002_d N_A_55_264#_M1011_d
+ N_A_55_264#_c_69_n N_A_55_264#_M1007_g N_A_55_264#_M1005_g N_A_55_264#_c_71_n
+ N_A_55_264#_M1006_g N_A_55_264#_c_73_n N_A_55_264#_c_82_n N_A_55_264#_M1008_g
+ N_A_55_264#_c_74_n N_A_55_264#_c_75_n N_A_55_264#_c_91_p N_A_55_264#_c_121_p
+ N_A_55_264#_c_76_n N_A_55_264#_c_77_n N_A_55_264#_c_78_n N_A_55_264#_c_84_n
+ N_A_55_264#_c_79_n N_A_55_264#_c_86_n PM_SKY130_FD_SC_LS__O31A_2%A_55_264#
x_PM_SKY130_FD_SC_LS__O31A_2%A1 N_A1_M1010_g N_A1_c_175_n N_A1_M1004_g A1 A1
+ N_A1_c_176_n PM_SKY130_FD_SC_LS__O31A_2%A1
x_PM_SKY130_FD_SC_LS__O31A_2%A2 N_A2_M1000_g N_A2_c_215_n N_A2_M1001_g A2 A2
+ PM_SKY130_FD_SC_LS__O31A_2%A2
x_PM_SKY130_FD_SC_LS__O31A_2%A3 N_A3_M1009_g N_A3_c_250_n N_A3_c_255_n
+ N_A3_M1011_g A3 N_A3_c_252_n N_A3_c_253_n PM_SKY130_FD_SC_LS__O31A_2%A3
x_PM_SKY130_FD_SC_LS__O31A_2%B1 N_B1_M1003_g N_B1_M1002_g N_B1_c_293_n
+ N_B1_c_297_n B1 N_B1_c_294_n N_B1_c_295_n PM_SKY130_FD_SC_LS__O31A_2%B1
x_PM_SKY130_FD_SC_LS__O31A_2%VPWR N_VPWR_M1007_d N_VPWR_M1008_d N_VPWR_M1003_d
+ N_VPWR_c_326_n N_VPWR_c_327_n N_VPWR_c_328_n N_VPWR_c_329_n N_VPWR_c_330_n
+ VPWR N_VPWR_c_331_n N_VPWR_c_332_n N_VPWR_c_333_n N_VPWR_c_325_n
+ PM_SKY130_FD_SC_LS__O31A_2%VPWR
x_PM_SKY130_FD_SC_LS__O31A_2%X N_X_M1005_d N_X_M1007_s N_X_c_368_n N_X_c_369_n
+ N_X_c_370_n X N_X_c_372_n PM_SKY130_FD_SC_LS__O31A_2%X
x_PM_SKY130_FD_SC_LS__O31A_2%VGND N_VGND_M1005_s N_VGND_M1006_s N_VGND_M1000_d
+ N_VGND_c_407_n N_VGND_c_408_n N_VGND_c_409_n N_VGND_c_410_n N_VGND_c_411_n
+ VGND N_VGND_c_412_n N_VGND_c_413_n N_VGND_c_414_n N_VGND_c_415_n
+ N_VGND_c_416_n PM_SKY130_FD_SC_LS__O31A_2%VGND
x_PM_SKY130_FD_SC_LS__O31A_2%A_328_74# N_A_328_74#_M1010_d N_A_328_74#_M1009_d
+ N_A_328_74#_c_455_n N_A_328_74#_c_456_n N_A_328_74#_c_465_n
+ N_A_328_74#_c_458_n PM_SKY130_FD_SC_LS__O31A_2%A_328_74#
cc_1 VNB N_A_55_264#_c_69_n 0.0378189f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_2 VNB N_A_55_264#_M1005_g 0.028293f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.74
cc_3 VNB N_A_55_264#_c_71_n 0.0148764f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=1.395
cc_4 VNB N_A_55_264#_M1006_g 0.0234109f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_5 VNB N_A_55_264#_c_73_n 0.00998306f $X=-0.19 $Y=-0.245 $X2=1.01 $Y2=1.675
cc_6 VNB N_A_55_264#_c_74_n 0.00775857f $X=-0.19 $Y=-0.245 $X2=1.01 $Y2=1.395
cc_7 VNB N_A_55_264#_c_75_n 5.59499e-19 $X=-0.19 $Y=-0.245 $X2=0.31 $Y2=2.32
cc_8 VNB N_A_55_264#_c_76_n 0.0100621f $X=-0.19 $Y=-0.245 $X2=3.56 $Y2=0.96
cc_9 VNB N_A_55_264#_c_77_n 0.0264193f $X=-0.19 $Y=-0.245 $X2=3.56 $Y2=0.515
cc_10 VNB N_A_55_264#_c_78_n 0.0130668f $X=-0.19 $Y=-0.245 $X2=0.44 $Y2=1.485
cc_11 VNB N_A_55_264#_c_79_n 0.00441108f $X=-0.19 $Y=-0.245 $X2=2.995 $Y2=1.94
cc_12 VNB N_A1_M1010_g 0.0273181f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A1_c_175_n 0.0260373f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A1_c_176_n 0.00624344f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=1.395
cc_15 VNB N_A2_M1000_g 0.0336545f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A2_c_215_n 0.0185605f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB A2 0.00275083f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_18 VNB N_A3_c_250_n 0.00649324f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB A3 0.0105601f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_20 VNB N_A3_c_252_n 0.0324936f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.74
cc_21 VNB N_A3_c_253_n 0.0202699f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=1.395
cc_22 VNB N_B1_M1002_g 0.0309473f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_23 VNB N_B1_c_293_n 0.00159338f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.32
cc_24 VNB N_B1_c_294_n 0.0716888f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_25 VNB N_B1_c_295_n 0.00435854f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VPWR_c_325_n 0.163682f $X=-0.19 $Y=-0.245 $X2=2.995 $Y2=2.405
cc_27 VNB N_X_c_368_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_28 VNB N_X_c_369_n 0.00291266f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.74
cc_29 VNB N_X_c_370_n 0.00418437f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_407_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.32
cc_31 VNB N_VGND_c_408_n 0.0477751f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.74
cc_32 VNB N_VGND_c_409_n 0.021169f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.32
cc_33 VNB N_VGND_c_410_n 0.0185368f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_34 VNB N_VGND_c_411_n 0.00673484f $X=-0.19 $Y=-0.245 $X2=1.01 $Y2=1.765
cc_35 VNB N_VGND_c_412_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0.31 $Y2=1.65
cc_36 VNB N_VGND_c_413_n 0.0384742f $X=-0.19 $Y=-0.245 $X2=3.56 $Y2=0.515
cc_37 VNB N_VGND_c_414_n 0.228611f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_415_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_416_n 0.0073872f $X=-0.19 $Y=-0.245 $X2=2.995 $Y2=1.94
cc_40 VNB N_A_328_74#_c_455_n 0.00760749f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_41 VNB N_A_328_74#_c_456_n 0.00280429f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_42 VPB N_A_55_264#_c_69_n 0.0246228f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_43 VPB N_A_55_264#_c_73_n 7.64023e-19 $X=-0.19 $Y=1.66 $X2=1.01 $Y2=1.675
cc_44 VPB N_A_55_264#_c_82_n 0.0227335f $X=-0.19 $Y=1.66 $X2=1.01 $Y2=1.765
cc_45 VPB N_A_55_264#_c_75_n 0.00756917f $X=-0.19 $Y=1.66 $X2=0.31 $Y2=2.32
cc_46 VPB N_A_55_264#_c_84_n 0.00834388f $X=-0.19 $Y=1.66 $X2=2.93 $Y2=2.105
cc_47 VPB N_A_55_264#_c_79_n 0.00303792f $X=-0.19 $Y=1.66 $X2=2.995 $Y2=1.94
cc_48 VPB N_A_55_264#_c_86_n 0.00326634f $X=-0.19 $Y=1.66 $X2=2.93 $Y2=2.46
cc_49 VPB N_A1_c_175_n 0.0324004f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_A1_c_176_n 0.00458039f $X=-0.19 $Y=1.66 $X2=0.92 $Y2=1.395
cc_51 VPB N_A2_c_215_n 0.035697f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB A2 0.00221071f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_53 VPB N_A3_c_250_n 0.00789082f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_A3_c_255_n 0.0245478f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_B1_c_293_n 0.00731593f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=1.32
cc_56 VPB N_B1_c_297_n 0.0275843f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=0.74
cc_57 VPB N_B1_c_295_n 0.00824274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_326_n 0.0120106f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=1.32
cc_59 VPB N_VPWR_c_327_n 0.0216574f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=0.74
cc_60 VPB N_VPWR_c_328_n 0.00478709f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=1.32
cc_61 VPB N_VPWR_c_329_n 0.0121909f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=0.74
cc_62 VPB N_VPWR_c_330_n 0.0540256f $X=-0.19 $Y=1.66 $X2=1.01 $Y2=1.47
cc_63 VPB N_VPWR_c_331_n 0.0195091f $X=-0.19 $Y=1.66 $X2=0.31 $Y2=1.65
cc_64 VPB N_VPWR_c_332_n 0.0534801f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_333_n 0.00971174f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_325_n 0.0672969f $X=-0.19 $Y=1.66 $X2=2.995 $Y2=2.405
cc_67 VPB N_X_c_369_n 0.00173426f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=0.74
cc_68 VPB N_X_c_372_n 0.0024942f $X=-0.19 $Y=1.66 $X2=1.01 $Y2=1.47
cc_69 N_A_55_264#_M1006_g N_A1_M1010_g 0.0226424f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_70 N_A_55_264#_c_74_n N_A1_M1010_g 0.00111862f $X=1.01 $Y=1.395 $X2=0 $Y2=0
cc_71 N_A_55_264#_c_82_n N_A1_c_175_n 0.0309064f $X=1.01 $Y=1.765 $X2=0 $Y2=0
cc_72 N_A_55_264#_c_74_n N_A1_c_175_n 0.0126587f $X=1.01 $Y=1.395 $X2=0 $Y2=0
cc_73 N_A_55_264#_c_91_p N_A1_c_175_n 0.0129544f $X=2.765 $Y=2.405 $X2=0 $Y2=0
cc_74 N_A_55_264#_c_82_n N_A1_c_176_n 0.00419315f $X=1.01 $Y=1.765 $X2=0 $Y2=0
cc_75 N_A_55_264#_c_74_n N_A1_c_176_n 0.00139611f $X=1.01 $Y=1.395 $X2=0 $Y2=0
cc_76 N_A_55_264#_c_91_p N_A1_c_176_n 0.0207012f $X=2.765 $Y=2.405 $X2=0 $Y2=0
cc_77 N_A_55_264#_c_91_p N_A2_c_215_n 0.0128905f $X=2.765 $Y=2.405 $X2=0 $Y2=0
cc_78 N_A_55_264#_c_91_p A2 0.0201317f $X=2.765 $Y=2.405 $X2=0 $Y2=0
cc_79 N_A_55_264#_c_84_n A2 0.00455465f $X=2.93 $Y=2.105 $X2=0 $Y2=0
cc_80 N_A_55_264#_c_79_n N_A3_c_250_n 0.00611211f $X=2.995 $Y=1.94 $X2=0 $Y2=0
cc_81 N_A_55_264#_c_91_p N_A3_c_255_n 0.0162548f $X=2.765 $Y=2.405 $X2=0 $Y2=0
cc_82 N_A_55_264#_c_84_n N_A3_c_255_n 0.00233406f $X=2.93 $Y=2.105 $X2=0 $Y2=0
cc_83 N_A_55_264#_c_79_n N_A3_c_255_n 9.6311e-19 $X=2.995 $Y=1.94 $X2=0 $Y2=0
cc_84 N_A_55_264#_c_86_n N_A3_c_255_n 0.00327892f $X=2.93 $Y=2.46 $X2=0 $Y2=0
cc_85 N_A_55_264#_c_84_n A3 0.00541843f $X=2.93 $Y=2.105 $X2=0 $Y2=0
cc_86 N_A_55_264#_c_79_n A3 0.0281608f $X=2.995 $Y=1.94 $X2=0 $Y2=0
cc_87 N_A_55_264#_c_84_n N_A3_c_252_n 8.3549e-19 $X=2.93 $Y=2.105 $X2=0 $Y2=0
cc_88 N_A_55_264#_c_79_n N_A3_c_252_n 0.00194886f $X=2.995 $Y=1.94 $X2=0 $Y2=0
cc_89 N_A_55_264#_c_76_n N_A3_c_253_n 0.00396327f $X=3.56 $Y=0.96 $X2=0 $Y2=0
cc_90 N_A_55_264#_c_79_n N_A3_c_253_n 0.00100883f $X=2.995 $Y=1.94 $X2=0 $Y2=0
cc_91 N_A_55_264#_c_76_n N_B1_M1002_g 0.0191744f $X=3.56 $Y=0.96 $X2=0 $Y2=0
cc_92 N_A_55_264#_c_77_n N_B1_M1002_g 0.0122539f $X=3.56 $Y=0.515 $X2=0 $Y2=0
cc_93 N_A_55_264#_c_79_n N_B1_M1002_g 0.00855406f $X=2.995 $Y=1.94 $X2=0 $Y2=0
cc_94 N_A_55_264#_c_79_n N_B1_c_293_n 0.00394106f $X=2.995 $Y=1.94 $X2=0 $Y2=0
cc_95 N_A_55_264#_c_84_n N_B1_c_297_n 0.00972136f $X=2.93 $Y=2.105 $X2=0 $Y2=0
cc_96 N_A_55_264#_c_79_n N_B1_c_297_n 0.00843713f $X=2.995 $Y=1.94 $X2=0 $Y2=0
cc_97 N_A_55_264#_c_86_n N_B1_c_297_n 0.0094783f $X=2.93 $Y=2.46 $X2=0 $Y2=0
cc_98 N_A_55_264#_c_76_n N_B1_c_294_n 0.0043993f $X=3.56 $Y=0.96 $X2=0 $Y2=0
cc_99 N_A_55_264#_c_79_n N_B1_c_294_n 0.0105781f $X=2.995 $Y=1.94 $X2=0 $Y2=0
cc_100 N_A_55_264#_c_76_n N_B1_c_295_n 0.0254991f $X=3.56 $Y=0.96 $X2=0 $Y2=0
cc_101 N_A_55_264#_c_79_n N_B1_c_295_n 0.0348575f $X=2.995 $Y=1.94 $X2=0 $Y2=0
cc_102 N_A_55_264#_c_75_n N_VPWR_M1007_d 0.0209621f $X=0.31 $Y=2.32 $X2=-0.19
+ $Y2=-0.245
cc_103 N_A_55_264#_c_121_p N_VPWR_M1007_d 0.00950867f $X=0.395 $Y=2.405
+ $X2=-0.19 $Y2=-0.245
cc_104 N_A_55_264#_c_91_p N_VPWR_M1008_d 0.0167554f $X=2.765 $Y=2.405 $X2=0
+ $Y2=0
cc_105 N_A_55_264#_c_69_n N_VPWR_c_327_n 0.0111125f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_106 N_A_55_264#_c_82_n N_VPWR_c_327_n 0.00130785f $X=1.01 $Y=1.765 $X2=0
+ $Y2=0
cc_107 N_A_55_264#_c_91_p N_VPWR_c_327_n 0.00100103f $X=2.765 $Y=2.405 $X2=0
+ $Y2=0
cc_108 N_A_55_264#_c_121_p N_VPWR_c_327_n 0.0129795f $X=0.395 $Y=2.405 $X2=0
+ $Y2=0
cc_109 N_A_55_264#_c_69_n N_VPWR_c_328_n 0.00130463f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_110 N_A_55_264#_c_82_n N_VPWR_c_328_n 0.0160434f $X=1.01 $Y=1.765 $X2=0 $Y2=0
cc_111 N_A_55_264#_c_91_p N_VPWR_c_328_n 0.0324048f $X=2.765 $Y=2.405 $X2=0
+ $Y2=0
cc_112 N_A_55_264#_c_84_n N_VPWR_c_330_n 0.0819742f $X=2.93 $Y=2.105 $X2=0 $Y2=0
cc_113 N_A_55_264#_c_69_n N_VPWR_c_331_n 0.00413917f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_114 N_A_55_264#_c_82_n N_VPWR_c_331_n 0.00413917f $X=1.01 $Y=1.765 $X2=0
+ $Y2=0
cc_115 N_A_55_264#_c_86_n N_VPWR_c_332_n 0.0200956f $X=2.93 $Y=2.46 $X2=0 $Y2=0
cc_116 N_A_55_264#_c_69_n N_VPWR_c_325_n 0.0041501f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_117 N_A_55_264#_c_82_n N_VPWR_c_325_n 0.0041501f $X=1.01 $Y=1.765 $X2=0 $Y2=0
cc_118 N_A_55_264#_c_91_p N_VPWR_c_325_n 0.0588629f $X=2.765 $Y=2.405 $X2=0
+ $Y2=0
cc_119 N_A_55_264#_c_121_p N_VPWR_c_325_n 6.15054e-19 $X=0.395 $Y=2.405 $X2=0
+ $Y2=0
cc_120 N_A_55_264#_c_86_n N_VPWR_c_325_n 0.0163656f $X=2.93 $Y=2.46 $X2=0 $Y2=0
cc_121 N_A_55_264#_c_91_p N_X_M1007_s 0.00738143f $X=2.765 $Y=2.405 $X2=0 $Y2=0
cc_122 N_A_55_264#_M1005_g N_X_c_368_n 0.00772833f $X=0.565 $Y=0.74 $X2=0 $Y2=0
cc_123 N_A_55_264#_M1006_g N_X_c_368_n 0.00752022f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_124 N_A_55_264#_c_69_n N_X_c_369_n 0.00262965f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_125 N_A_55_264#_M1005_g N_X_c_369_n 0.00408016f $X=0.565 $Y=0.74 $X2=0 $Y2=0
cc_126 N_A_55_264#_c_71_n N_X_c_369_n 0.00833621f $X=0.92 $Y=1.395 $X2=0 $Y2=0
cc_127 N_A_55_264#_M1006_g N_X_c_369_n 0.00495702f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_128 N_A_55_264#_c_73_n N_X_c_369_n 0.00503245f $X=1.01 $Y=1.675 $X2=0 $Y2=0
cc_129 N_A_55_264#_c_82_n N_X_c_369_n 0.00399275f $X=1.01 $Y=1.765 $X2=0 $Y2=0
cc_130 N_A_55_264#_c_74_n N_X_c_369_n 0.00266977f $X=1.01 $Y=1.395 $X2=0 $Y2=0
cc_131 N_A_55_264#_c_75_n N_X_c_369_n 0.00731165f $X=0.31 $Y=2.32 $X2=0 $Y2=0
cc_132 N_A_55_264#_c_78_n N_X_c_369_n 0.0244835f $X=0.44 $Y=1.485 $X2=0 $Y2=0
cc_133 N_A_55_264#_M1005_g N_X_c_370_n 0.00316168f $X=0.565 $Y=0.74 $X2=0 $Y2=0
cc_134 N_A_55_264#_c_71_n N_X_c_370_n 0.00181038f $X=0.92 $Y=1.395 $X2=0 $Y2=0
cc_135 N_A_55_264#_M1006_g N_X_c_370_n 0.00193058f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_136 N_A_55_264#_c_69_n N_X_c_372_n 0.00623195f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_137 N_A_55_264#_c_71_n N_X_c_372_n 0.00512017f $X=0.92 $Y=1.395 $X2=0 $Y2=0
cc_138 N_A_55_264#_c_82_n N_X_c_372_n 0.00630519f $X=1.01 $Y=1.765 $X2=0 $Y2=0
cc_139 N_A_55_264#_c_75_n N_X_c_372_n 0.013351f $X=0.31 $Y=2.32 $X2=0 $Y2=0
cc_140 N_A_55_264#_c_91_p N_X_c_372_n 0.020485f $X=2.765 $Y=2.405 $X2=0 $Y2=0
cc_141 N_A_55_264#_c_78_n N_X_c_372_n 0.00310399f $X=0.44 $Y=1.485 $X2=0 $Y2=0
cc_142 N_A_55_264#_c_91_p A_346_392# 0.00889595f $X=2.765 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_143 N_A_55_264#_c_91_p A_430_392# 0.0153203f $X=2.765 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_144 N_A_55_264#_c_69_n N_VGND_c_408_n 0.00397263f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_145 N_A_55_264#_M1005_g N_VGND_c_408_n 0.0184907f $X=0.565 $Y=0.74 $X2=0
+ $Y2=0
cc_146 N_A_55_264#_c_78_n N_VGND_c_408_n 0.0171976f $X=0.44 $Y=1.485 $X2=0 $Y2=0
cc_147 N_A_55_264#_M1006_g N_VGND_c_409_n 0.00666821f $X=0.995 $Y=0.74 $X2=0
+ $Y2=0
cc_148 N_A_55_264#_M1005_g N_VGND_c_412_n 0.00434272f $X=0.565 $Y=0.74 $X2=0
+ $Y2=0
cc_149 N_A_55_264#_M1006_g N_VGND_c_412_n 0.00434272f $X=0.995 $Y=0.74 $X2=0
+ $Y2=0
cc_150 N_A_55_264#_c_77_n N_VGND_c_413_n 0.0145203f $X=3.56 $Y=0.515 $X2=0 $Y2=0
cc_151 N_A_55_264#_M1005_g N_VGND_c_414_n 0.00823934f $X=0.565 $Y=0.74 $X2=0
+ $Y2=0
cc_152 N_A_55_264#_M1006_g N_VGND_c_414_n 0.00821312f $X=0.995 $Y=0.74 $X2=0
+ $Y2=0
cc_153 N_A_55_264#_c_77_n N_VGND_c_414_n 0.0120696f $X=3.56 $Y=0.515 $X2=0 $Y2=0
cc_154 N_A_55_264#_c_76_n N_A_328_74#_M1009_d 0.00329864f $X=3.56 $Y=0.96 $X2=0
+ $Y2=0
cc_155 N_A_55_264#_c_76_n N_A_328_74#_c_458_n 0.00855261f $X=3.56 $Y=0.96 $X2=0
+ $Y2=0
cc_156 N_A1_M1010_g N_A2_M1000_g 0.0252626f $X=1.565 $Y=0.74 $X2=0 $Y2=0
cc_157 N_A1_c_175_n N_A2_M1000_g 0.027699f $X=1.655 $Y=1.885 $X2=0 $Y2=0
cc_158 N_A1_c_176_n N_A2_M1000_g 0.00530086f $X=1.58 $Y=1.515 $X2=0 $Y2=0
cc_159 N_A1_c_175_n N_A2_c_215_n 0.0587416f $X=1.655 $Y=1.885 $X2=0 $Y2=0
cc_160 N_A1_c_176_n N_A2_c_215_n 9.40794e-19 $X=1.58 $Y=1.515 $X2=0 $Y2=0
cc_161 N_A1_c_175_n A2 8.4161e-19 $X=1.655 $Y=1.885 $X2=0 $Y2=0
cc_162 N_A1_c_176_n A2 0.0435211f $X=1.58 $Y=1.515 $X2=0 $Y2=0
cc_163 N_A1_c_176_n N_VPWR_M1008_d 0.00384295f $X=1.58 $Y=1.515 $X2=0 $Y2=0
cc_164 N_A1_c_175_n N_VPWR_c_328_n 0.0159146f $X=1.655 $Y=1.885 $X2=0 $Y2=0
cc_165 N_A1_c_175_n N_VPWR_c_332_n 0.00413917f $X=1.655 $Y=1.885 $X2=0 $Y2=0
cc_166 N_A1_c_175_n N_VPWR_c_325_n 0.00414311f $X=1.655 $Y=1.885 $X2=0 $Y2=0
cc_167 N_A1_M1010_g N_X_c_368_n 0.00115542f $X=1.565 $Y=0.74 $X2=0 $Y2=0
cc_168 N_A1_c_175_n N_X_c_369_n 0.00116914f $X=1.655 $Y=1.885 $X2=0 $Y2=0
cc_169 N_A1_c_176_n N_X_c_369_n 0.0154056f $X=1.58 $Y=1.515 $X2=0 $Y2=0
cc_170 N_A1_c_175_n N_X_c_372_n 2.80093e-19 $X=1.655 $Y=1.885 $X2=0 $Y2=0
cc_171 N_A1_c_176_n N_X_c_372_n 0.0122126f $X=1.58 $Y=1.515 $X2=0 $Y2=0
cc_172 N_A1_c_176_n A_346_392# 0.00179993f $X=1.58 $Y=1.515 $X2=-0.19 $Y2=-0.245
cc_173 N_A1_M1010_g N_VGND_c_409_n 0.00666787f $X=1.565 $Y=0.74 $X2=0 $Y2=0
cc_174 N_A1_c_175_n N_VGND_c_409_n 2.14662e-19 $X=1.655 $Y=1.885 $X2=0 $Y2=0
cc_175 N_A1_c_176_n N_VGND_c_409_n 0.00205464f $X=1.58 $Y=1.515 $X2=0 $Y2=0
cc_176 N_A1_M1010_g N_VGND_c_410_n 0.00434272f $X=1.565 $Y=0.74 $X2=0 $Y2=0
cc_177 N_A1_M1010_g N_VGND_c_411_n 4.1081e-19 $X=1.565 $Y=0.74 $X2=0 $Y2=0
cc_178 N_A1_M1010_g N_VGND_c_414_n 0.00821983f $X=1.565 $Y=0.74 $X2=0 $Y2=0
cc_179 N_A1_M1010_g N_A_328_74#_c_455_n 0.00437183f $X=1.565 $Y=0.74 $X2=0 $Y2=0
cc_180 N_A1_c_175_n N_A_328_74#_c_455_n 7.96959e-19 $X=1.655 $Y=1.885 $X2=0
+ $Y2=0
cc_181 N_A1_c_176_n N_A_328_74#_c_455_n 0.0132489f $X=1.58 $Y=1.515 $X2=0 $Y2=0
cc_182 N_A1_M1010_g N_A_328_74#_c_456_n 0.00549371f $X=1.565 $Y=0.74 $X2=0 $Y2=0
cc_183 A2 N_A3_c_250_n 0.00164156f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_184 N_A2_c_215_n N_A3_c_255_n 0.0367877f $X=2.075 $Y=1.885 $X2=0 $Y2=0
cc_185 A2 N_A3_c_255_n 0.00510705f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_186 N_A2_M1000_g A3 0.00565381f $X=2.06 $Y=0.74 $X2=0 $Y2=0
cc_187 N_A2_c_215_n A3 4.91538e-19 $X=2.075 $Y=1.885 $X2=0 $Y2=0
cc_188 A2 A3 0.00544377f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_189 N_A2_c_215_n N_A3_c_252_n 0.0183284f $X=2.075 $Y=1.885 $X2=0 $Y2=0
cc_190 N_A2_M1000_g N_A3_c_253_n 0.0270404f $X=2.06 $Y=0.74 $X2=0 $Y2=0
cc_191 N_A2_c_215_n N_VPWR_c_328_n 0.00206865f $X=2.075 $Y=1.885 $X2=0 $Y2=0
cc_192 N_A2_c_215_n N_VPWR_c_332_n 0.00461464f $X=2.075 $Y=1.885 $X2=0 $Y2=0
cc_193 N_A2_c_215_n N_VPWR_c_325_n 0.00465844f $X=2.075 $Y=1.885 $X2=0 $Y2=0
cc_194 A2 A_430_392# 0.00371845f $X=2.075 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_195 N_A2_M1000_g N_VGND_c_410_n 0.00398535f $X=2.06 $Y=0.74 $X2=0 $Y2=0
cc_196 N_A2_M1000_g N_VGND_c_411_n 0.00710985f $X=2.06 $Y=0.74 $X2=0 $Y2=0
cc_197 N_A2_M1000_g N_VGND_c_414_n 0.00384527f $X=2.06 $Y=0.74 $X2=0 $Y2=0
cc_198 N_A2_M1000_g N_A_328_74#_c_455_n 0.00143395f $X=2.06 $Y=0.74 $X2=0 $Y2=0
cc_199 N_A2_M1000_g N_A_328_74#_c_456_n 0.00224861f $X=2.06 $Y=0.74 $X2=0 $Y2=0
cc_200 N_A2_M1000_g N_A_328_74#_c_465_n 0.0142189f $X=2.06 $Y=0.74 $X2=0 $Y2=0
cc_201 N_A2_c_215_n N_A_328_74#_c_465_n 7.72429e-19 $X=2.075 $Y=1.885 $X2=0
+ $Y2=0
cc_202 A2 N_A_328_74#_c_465_n 0.00933039f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_203 N_A2_M1000_g N_A_328_74#_c_458_n 5.02222e-19 $X=2.06 $Y=0.74 $X2=0 $Y2=0
cc_204 N_A3_c_252_n N_B1_M1002_g 0.002904f $X=2.72 $Y=1.385 $X2=0 $Y2=0
cc_205 N_A3_c_253_n N_B1_M1002_g 0.0197735f $X=2.72 $Y=1.22 $X2=0 $Y2=0
cc_206 N_A3_c_250_n N_B1_c_297_n 0.0026884f $X=2.645 $Y=1.795 $X2=0 $Y2=0
cc_207 N_A3_c_255_n N_B1_c_297_n 0.0174149f $X=2.645 $Y=1.885 $X2=0 $Y2=0
cc_208 N_A3_c_250_n N_B1_c_294_n 0.00641549f $X=2.645 $Y=1.795 $X2=0 $Y2=0
cc_209 A3 N_B1_c_294_n 2.74107e-19 $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_210 N_A3_c_252_n N_B1_c_294_n 0.0132146f $X=2.72 $Y=1.385 $X2=0 $Y2=0
cc_211 N_A3_c_255_n N_VPWR_c_332_n 0.00461464f $X=2.645 $Y=1.885 $X2=0 $Y2=0
cc_212 N_A3_c_255_n N_VPWR_c_325_n 0.0046687f $X=2.645 $Y=1.885 $X2=0 $Y2=0
cc_213 N_A3_c_253_n N_VGND_c_411_n 0.0052684f $X=2.72 $Y=1.22 $X2=0 $Y2=0
cc_214 N_A3_c_253_n N_VGND_c_413_n 0.0043552f $X=2.72 $Y=1.22 $X2=0 $Y2=0
cc_215 N_A3_c_253_n N_VGND_c_414_n 0.00436921f $X=2.72 $Y=1.22 $X2=0 $Y2=0
cc_216 A3 N_A_328_74#_c_465_n 0.0078091f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_217 N_A3_c_253_n N_A_328_74#_c_465_n 0.00931502f $X=2.72 $Y=1.22 $X2=0 $Y2=0
cc_218 A3 N_A_328_74#_c_458_n 0.010823f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_219 N_A3_c_252_n N_A_328_74#_c_458_n 9.87553e-19 $X=2.72 $Y=1.385 $X2=0 $Y2=0
cc_220 N_A3_c_253_n N_A_328_74#_c_458_n 0.01381f $X=2.72 $Y=1.22 $X2=0 $Y2=0
cc_221 N_B1_c_297_n N_VPWR_c_330_n 0.025097f $X=3.192 $Y=1.885 $X2=0 $Y2=0
cc_222 N_B1_c_294_n N_VPWR_c_330_n 0.00181048f $X=3.56 $Y=1.465 $X2=0 $Y2=0
cc_223 N_B1_c_295_n N_VPWR_c_330_n 0.0299469f $X=3.56 $Y=1.465 $X2=0 $Y2=0
cc_224 N_B1_c_297_n N_VPWR_c_332_n 0.00332301f $X=3.192 $Y=1.885 $X2=0 $Y2=0
cc_225 N_B1_c_297_n N_VPWR_c_325_n 0.0049621f $X=3.192 $Y=1.885 $X2=0 $Y2=0
cc_226 N_B1_M1002_g N_VGND_c_413_n 0.0043552f $X=3.275 $Y=0.74 $X2=0 $Y2=0
cc_227 N_B1_M1002_g N_VGND_c_414_n 0.00825941f $X=3.275 $Y=0.74 $X2=0 $Y2=0
cc_228 N_B1_M1002_g N_A_328_74#_c_458_n 0.0115428f $X=3.275 $Y=0.74 $X2=0 $Y2=0
cc_229 N_X_c_368_n N_VGND_c_408_n 0.0308109f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_230 N_X_c_368_n N_VGND_c_409_n 0.0308109f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_231 N_X_c_368_n N_VGND_c_412_n 0.0144922f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_232 N_X_c_368_n N_VGND_c_414_n 0.0118826f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_233 N_VGND_c_409_n N_A_328_74#_c_455_n 0.0151247f $X=1.28 $Y=0.515 $X2=0
+ $Y2=0
cc_234 N_VGND_c_409_n N_A_328_74#_c_456_n 0.0165124f $X=1.28 $Y=0.515 $X2=0
+ $Y2=0
cc_235 N_VGND_c_410_n N_A_328_74#_c_456_n 0.0145639f $X=2.115 $Y=0 $X2=0 $Y2=0
cc_236 N_VGND_c_411_n N_A_328_74#_c_456_n 0.0104328f $X=2.31 $Y=0.515 $X2=0
+ $Y2=0
cc_237 N_VGND_c_414_n N_A_328_74#_c_456_n 0.0119984f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_238 N_VGND_M1000_d N_A_328_74#_c_465_n 0.0126964f $X=2.135 $Y=0.37 $X2=0
+ $Y2=0
cc_239 N_VGND_c_411_n N_A_328_74#_c_465_n 0.0255658f $X=2.31 $Y=0.515 $X2=0
+ $Y2=0
cc_240 N_VGND_c_414_n N_A_328_74#_c_465_n 0.0120739f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_241 N_VGND_c_413_n N_A_328_74#_c_458_n 0.0140542f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_242 N_VGND_c_414_n N_A_328_74#_c_458_n 0.0180651f $X=3.6 $Y=0 $X2=0 $Y2=0
