* File: sky130_fd_sc_ls__o211ai_1.pex.spice
* Created: Fri Aug 28 13:43:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__O211AI_1%A1 1 3 6 8 12
c24 1 0 1.96061e-19 $X=0.505 $Y=1.765
r25 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.465 $X2=0.27 $Y2=1.465
r26 8 12 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=0.27 $Y=1.665 $X2=0.27
+ $Y2=1.465
r27 4 11 39.5853 $w=4e-07 $l=2.33345e-07 $layer=POLY_cond $X=0.515 $Y=1.3
+ $X2=0.35 $Y2=1.465
r28 4 6 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.515 $Y=1.3 $X2=0.515
+ $Y2=0.74
r29 1 11 55.8528 $w=4e-07 $l=3.69459e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.35 $Y2=1.465
r30 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__O211AI_1%A2 1 3 6 8 9 10 11 22
r35 20 22 1.75372 $w=2.28e-07 $l=3.5e-08 $layer=LI1_cond $X=0.72 $Y=1.63
+ $X2=0.72 $Y2=1.665
r36 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1 $Y=1.465
+ $X2=1 $Y2=1.465
r37 10 11 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.72 $Y=2.405
+ $X2=0.72 $Y2=2.775
r38 9 10 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.72 $Y=2.035
+ $X2=0.72 $Y2=2.405
r39 8 19 11.2739 $w=3.03e-07 $l=2.8e-07 $layer=LI1_cond $X=0.72 $Y=1.465 $X2=1
+ $Y2=1.465
r40 8 20 2.35376 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=0.72 $Y=1.465
+ $X2=0.72 $Y2=1.63
r41 8 9 17.2866 $w=2.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.72 $Y=1.69 $X2=0.72
+ $Y2=2.035
r42 8 22 1.25266 $w=2.28e-07 $l=2.5e-08 $layer=LI1_cond $X=0.72 $Y=1.69 $X2=0.72
+ $Y2=1.665
r43 4 18 38.6549 $w=2.86e-07 $l=1.72337e-07 $layer=POLY_cond $X=1.015 $Y=1.3
+ $X2=1 $Y2=1.465
r44 4 6 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.015 $Y=1.3 $X2=1.015
+ $Y2=0.74
r45 1 18 61.4066 $w=2.86e-07 $l=3.3541e-07 $layer=POLY_cond $X=0.925 $Y=1.765
+ $X2=1 $Y2=1.465
r46 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.925 $Y=1.765
+ $X2=0.925 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__O211AI_1%B1 3 5 7 8 9 10 26
c35 3 0 1.83455e-19 $X=1.48 $Y=0.74
r36 18 26 0.250531 $w=2.28e-07 $l=5e-09 $layer=LI1_cond $X=1.68 $Y=1.3 $X2=1.68
+ $Y2=1.295
r37 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.57
+ $Y=1.465 $X2=1.57 $Y2=1.465
r38 10 17 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=1.68 $Y=1.465
+ $X2=1.57 $Y2=1.465
r39 10 18 2.85155 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=1.68 $Y=1.465
+ $X2=1.68 $Y2=1.3
r40 10 26 2.00425 $w=2.28e-07 $l=4e-08 $layer=LI1_cond $X=1.68 $Y=1.255 $X2=1.68
+ $Y2=1.295
r41 9 10 16.5351 $w=2.28e-07 $l=3.3e-07 $layer=LI1_cond $X=1.68 $Y=0.925
+ $X2=1.68 $Y2=1.255
r42 8 9 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.68 $Y=0.555 $X2=1.68
+ $Y2=0.925
r43 5 16 61.4066 $w=2.86e-07 $l=3.3541e-07 $layer=POLY_cond $X=1.645 $Y=1.765
+ $X2=1.57 $Y2=1.465
r44 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.645 $Y=1.765
+ $X2=1.645 $Y2=2.4
r45 1 16 38.6549 $w=2.86e-07 $l=2.05122e-07 $layer=POLY_cond $X=1.48 $Y=1.3
+ $X2=1.57 $Y2=1.465
r46 1 3 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.48 $Y=1.3 $X2=1.48
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__O211AI_1%C1 1 3 4 6 7
r27 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.14
+ $Y=1.385 $X2=2.14 $Y2=1.385
r28 7 11 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=2.14 $Y=1.295 $X2=2.14
+ $Y2=1.385
r29 4 10 77.2841 $w=2.7e-07 $l=3.82492e-07 $layer=POLY_cond $X=2.145 $Y=1.765
+ $X2=2.14 $Y2=1.385
r30 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.145 $Y=1.765
+ $X2=2.145 $Y2=2.4
r31 1 10 38.9026 $w=2.7e-07 $l=2.05122e-07 $layer=POLY_cond $X=2.05 $Y=1.22
+ $X2=2.14 $Y2=1.385
r32 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.05 $Y=1.22 $X2=2.05
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__O211AI_1%VPWR 1 2 7 9 15 18 19 20 30 31
r30 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r31 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r32 28 31 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r33 27 28 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r34 25 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r35 24 27 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=3.33 $X2=1.68
+ $Y2=3.33
r36 24 25 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r37 22 34 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.182 $Y2=3.33
r38 22 24 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.72 $Y2=3.33
r39 20 28 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.68 $Y2=3.33
r40 20 25 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=0.72 $Y2=3.33
r41 18 27 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=1.705 $Y=3.33
+ $X2=1.68 $Y2=3.33
r42 18 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.705 $Y=3.33
+ $X2=1.87 $Y2=3.33
r43 17 30 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=2.035 $Y=3.33
+ $X2=2.64 $Y2=3.33
r44 17 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.035 $Y=3.33
+ $X2=1.87 $Y2=3.33
r45 13 19 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.87 $Y=3.245
+ $X2=1.87 $Y2=3.33
r46 13 15 32.8272 $w=3.28e-07 $l=9.4e-07 $layer=LI1_cond $X=1.87 $Y=3.245
+ $X2=1.87 $Y2=2.305
r47 9 12 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=0.24 $Y=2.115 $X2=0.24
+ $Y2=2.815
r48 7 34 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.182 $Y2=3.33
r49 7 12 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.24 $Y=3.245 $X2=0.24
+ $Y2=2.815
r50 2 15 300 $w=1.7e-07 $l=5.34766e-07 $layer=licon1_PDIFF $count=2 $X=1.72
+ $Y=1.84 $X2=1.87 $Y2=2.305
r51 1 12 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r52 1 9 400 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_LS__O211AI_1%Y 1 2 3 12 16 17 20 25 26 27 28 37
r41 28 37 1.61576 $w=5.68e-07 $l=7.7e-08 $layer=LI1_cond $X=2.605 $Y=0.725
+ $X2=2.682 $Y2=0.725
r42 27 28 9.3378 $w=5.68e-07 $l=4.45e-07 $layer=LI1_cond $X=2.16 $Y=0.725
+ $X2=2.605 $Y2=0.725
r43 25 26 2.59952 $w=3.7e-07 $l=2.33666e-07 $layer=LI1_cond $X=2.682 $Y=1.8
+ $X2=2.487 $Y2=1.885
r44 24 37 7.81285 $w=1.75e-07 $l=2.85e-07 $layer=LI1_cond $X=2.682 $Y=1.01
+ $X2=2.682 $Y2=0.725
r45 24 25 50.0675 $w=1.73e-07 $l=7.9e-07 $layer=LI1_cond $X=2.682 $Y=1.01
+ $X2=2.682 $Y2=1.8
r46 20 22 17.5707 $w=5.63e-07 $l=8.3e-07 $layer=LI1_cond $X=2.487 $Y=1.985
+ $X2=2.487 $Y2=2.815
r47 18 26 2.59952 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.487 $Y=1.97
+ $X2=2.487 $Y2=1.885
r48 18 20 0.317543 $w=5.63e-07 $l=1.5e-08 $layer=LI1_cond $X=2.487 $Y=1.97
+ $X2=2.487 $Y2=1.985
r49 16 26 4.24538 $w=1.7e-07 $l=2.82e-07 $layer=LI1_cond $X=2.205 $Y=1.885
+ $X2=2.487 $Y2=1.885
r50 16 17 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=2.205 $Y=1.885
+ $X2=1.455 $Y2=1.885
r51 12 14 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=1.29 $Y=1.985
+ $X2=1.29 $Y2=2.815
r52 10 17 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.29 $Y=1.97
+ $X2=1.455 $Y2=1.885
r53 10 12 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=1.29 $Y=1.97
+ $X2=1.29 $Y2=1.985
r54 3 22 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.22
+ $Y=1.84 $X2=2.37 $Y2=2.815
r55 3 20 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.22
+ $Y=1.84 $X2=2.37 $Y2=1.985
r56 2 14 400 $w=1.7e-07 $l=1.11057e-06 $layer=licon1_PDIFF $count=1 $X=1 $Y=1.84
+ $X2=1.29 $Y2=2.815
r57 2 12 400 $w=1.7e-07 $l=3.55176e-07 $layer=licon1_PDIFF $count=1 $X=1 $Y=1.84
+ $X2=1.29 $Y2=1.985
r58 1 28 45.5 $w=1.7e-07 $l=5.67098e-07 $layer=licon1_NDIFF $count=4 $X=2.125
+ $Y=0.37 $X2=2.605 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_LS__O211AI_1%A_31_74# 1 2 9 11 12 15
c25 11 0 3.79516e-19 $X=1.145 $Y=1.045
r26 13 15 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=1.27 $Y=0.96
+ $X2=1.27 $Y2=0.515
r27 11 13 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.145 $Y=1.045
+ $X2=1.27 $Y2=0.96
r28 11 12 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.145 $Y=1.045
+ $X2=0.465 $Y2=1.045
r29 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.3 $Y=0.96
+ $X2=0.465 $Y2=1.045
r30 7 9 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=0.3 $Y=0.96 $X2=0.3
+ $Y2=0.515
r31 2 15 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.09
+ $Y=0.37 $X2=1.23 $Y2=0.515
r32 1 9 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.155
+ $Y=0.37 $X2=0.3 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__O211AI_1%VGND 1 6 8 10 20 21 24
r28 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r29 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r30 18 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r31 17 20 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r32 17 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r33 15 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.965 $Y=0 $X2=0.8
+ $Y2=0
r34 15 17 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=0.965 $Y=0 $X2=1.2
+ $Y2=0
r35 13 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r36 12 13 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r37 10 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.635 $Y=0 $X2=0.8
+ $Y2=0
r38 10 12 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=0.635 $Y=0 $X2=0.24
+ $Y2=0
r39 8 21 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.44 $Y=0 $X2=2.64
+ $Y2=0
r40 8 18 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.2
+ $Y2=0
r41 4 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.8 $Y=0.085 $X2=0.8
+ $Y2=0
r42 4 6 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=0.8 $Y=0.085 $X2=0.8
+ $Y2=0.615
r43 1 6 182 $w=1.7e-07 $l=3.33879e-07 $layer=licon1_NDIFF $count=1 $X=0.59
+ $Y=0.37 $X2=0.8 $Y2=0.615
.ends

