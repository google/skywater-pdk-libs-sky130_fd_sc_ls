* File: sky130_fd_sc_ls__and4b_2.pxi.spice
* Created: Fri Aug 28 13:05:50 2020
* 
x_PM_SKY130_FD_SC_LS__AND4B_2%A_N N_A_N_M1005_g N_A_N_c_73_n N_A_N_M1008_g A_N
+ N_A_N_c_74_n PM_SKY130_FD_SC_LS__AND4B_2%A_N
x_PM_SKY130_FD_SC_LS__AND4B_2%A_186_48# N_A_186_48#_M1007_d N_A_186_48#_M1002_d
+ N_A_186_48#_M1006_d N_A_186_48#_M1003_g N_A_186_48#_c_108_n
+ N_A_186_48#_M1009_g N_A_186_48#_M1011_g N_A_186_48#_c_109_n
+ N_A_186_48#_M1012_g N_A_186_48#_c_102_n N_A_186_48#_c_103_n
+ N_A_186_48#_c_171_p N_A_186_48#_c_153_p N_A_186_48#_c_118_p
+ N_A_186_48#_c_104_n N_A_186_48#_c_105_n N_A_186_48#_c_106_n
+ N_A_186_48#_c_107_n PM_SKY130_FD_SC_LS__AND4B_2%A_186_48#
x_PM_SKY130_FD_SC_LS__AND4B_2%D N_D_c_205_n N_D_M1002_g N_D_M1001_g D
+ N_D_c_207_n PM_SKY130_FD_SC_LS__AND4B_2%D
x_PM_SKY130_FD_SC_LS__AND4B_2%C N_C_c_236_n N_C_M1010_g N_C_M1000_g C
+ N_C_c_238_n PM_SKY130_FD_SC_LS__AND4B_2%C
x_PM_SKY130_FD_SC_LS__AND4B_2%B N_B_M1004_g N_B_c_264_n N_B_M1006_g B
+ N_B_c_265_n PM_SKY130_FD_SC_LS__AND4B_2%B
x_PM_SKY130_FD_SC_LS__AND4B_2%A_27_112# N_A_27_112#_M1005_s N_A_27_112#_M1008_s
+ N_A_27_112#_M1007_g N_A_27_112#_c_292_n N_A_27_112#_M1013_g
+ N_A_27_112#_c_293_n N_A_27_112#_c_294_n N_A_27_112#_c_295_n
+ N_A_27_112#_c_296_n N_A_27_112#_c_324_n N_A_27_112#_c_300_n
+ N_A_27_112#_c_301_n N_A_27_112#_c_297_n PM_SKY130_FD_SC_LS__AND4B_2%A_27_112#
x_PM_SKY130_FD_SC_LS__AND4B_2%VPWR N_VPWR_M1008_d N_VPWR_M1012_s N_VPWR_M1010_d
+ N_VPWR_M1013_d N_VPWR_c_375_n N_VPWR_c_376_n N_VPWR_c_377_n N_VPWR_c_378_n
+ N_VPWR_c_379_n N_VPWR_c_380_n N_VPWR_c_381_n N_VPWR_c_382_n VPWR
+ N_VPWR_c_383_n N_VPWR_c_384_n N_VPWR_c_385_n N_VPWR_c_374_n
+ PM_SKY130_FD_SC_LS__AND4B_2%VPWR
x_PM_SKY130_FD_SC_LS__AND4B_2%X N_X_M1003_s N_X_M1009_d N_X_c_428_n N_X_c_429_n
+ N_X_c_430_n X PM_SKY130_FD_SC_LS__AND4B_2%X
x_PM_SKY130_FD_SC_LS__AND4B_2%VGND N_VGND_M1005_d N_VGND_M1011_d N_VGND_c_465_n
+ N_VGND_c_466_n VGND N_VGND_c_467_n N_VGND_c_468_n N_VGND_c_469_n
+ N_VGND_c_470_n N_VGND_c_471_n N_VGND_c_472_n PM_SKY130_FD_SC_LS__AND4B_2%VGND
cc_1 VNB N_A_N_M1005_g 0.0304431f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.835
cc_2 VNB N_A_N_c_73_n 0.0605514f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_3 VNB N_A_N_c_74_n 0.00385705f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_4 VNB N_A_186_48#_M1003_g 0.021717f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_5 VNB N_A_186_48#_M1011_g 0.0244852f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_A_186_48#_c_102_n 4.01658e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_186_48#_c_103_n 0.0433786f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_186_48#_c_104_n 0.02581f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_186_48#_c_105_n 0.00578534f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_186_48#_c_106_n 0.00320654f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_186_48#_c_107_n 0.0636355f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_D_c_205_n 0.0267808f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.3
cc_13 VNB N_D_M1001_g 0.0266603f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.26
cc_14 VNB N_D_c_207_n 0.00182951f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_15 VNB N_C_c_236_n 0.0266079f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.3
cc_16 VNB N_C_M1000_g 0.0256596f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.26
cc_17 VNB N_C_c_238_n 0.00181929f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_18 VNB N_B_M1004_g 0.0276909f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.835
cc_19 VNB N_B_c_264_n 0.0246959f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_20 VNB N_B_c_265_n 0.00442487f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_21 VNB N_A_27_112#_M1007_g 0.0358374f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_27_112#_c_292_n 0.0273588f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_23 VNB N_A_27_112#_c_293_n 0.0195128f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_27_112#_c_294_n 0.00140869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_27_112#_c_295_n 0.00927871f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_27_112#_c_296_n 0.00959177f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_27_112#_c_297_n 0.0141382f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VPWR_c_374_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_X_c_428_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_X_c_429_n 0.00156999f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_31 VNB N_X_c_430_n 0.00417716f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_32 VNB N_VGND_c_465_n 0.0157594f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_466_n 0.00951062f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_34 VNB N_VGND_c_467_n 0.0202692f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_468_n 0.019013f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_469_n 0.0679994f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_470_n 0.292092f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_471_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_472_n 0.0115483f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VPB N_A_N_c_73_n 0.0296463f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_41 VPB N_A_N_c_74_n 0.00730438f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.465
cc_42 VPB N_A_186_48#_c_108_n 0.0169158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_43 VPB N_A_186_48#_c_109_n 0.0166172f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_44 VPB N_A_186_48#_c_102_n 0.00289025f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_45 VPB N_A_186_48#_c_107_n 0.0137528f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_D_c_205_n 0.0275707f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.3
cc_47 VPB N_D_c_207_n 0.00301842f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.465
cc_48 VPB N_C_c_236_n 0.0279903f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.3
cc_49 VPB N_C_c_238_n 0.00241094f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.465
cc_50 VPB N_B_c_264_n 0.0275524f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_51 VPB N_B_c_265_n 0.00394399f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.465
cc_52 VPB N_A_27_112#_c_292_n 0.0280322f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.465
cc_53 VPB N_A_27_112#_c_296_n 0.00320132f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_A_27_112#_c_300_n 0.00692485f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_A_27_112#_c_301_n 0.0352878f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_A_27_112#_c_297_n 9.55674e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_375_n 0.0165704f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_376_n 0.02094f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_377_n 0.0136955f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_378_n 0.0191737f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_379_n 0.0126731f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_380_n 0.0289141f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_381_n 0.0242802f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_382_n 0.00632279f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_383_n 0.0247575f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_384_n 0.0274955f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_385_n 0.00632279f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_374_n 0.0771067f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_X_c_429_n 0.00157267f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.465
cc_70 VPB X 0.00222f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 N_A_N_M1005_g N_A_186_48#_M1003_g 0.0179601f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_72 N_A_N_c_73_n N_A_186_48#_c_108_n 0.0244097f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_73 N_A_N_c_73_n N_A_186_48#_c_107_n 0.0136501f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_74 N_A_N_M1005_g N_A_27_112#_c_293_n 0.00822581f $X=0.495 $Y=0.835 $X2=0
+ $Y2=0
cc_75 N_A_N_M1005_g N_A_27_112#_c_294_n 0.0142232f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_76 N_A_N_c_73_n N_A_27_112#_c_294_n 0.00100324f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_77 N_A_N_c_74_n N_A_27_112#_c_294_n 6.31955e-19 $X=0.29 $Y=1.465 $X2=0 $Y2=0
cc_78 N_A_N_M1005_g N_A_27_112#_c_295_n 0.00275868f $X=0.495 $Y=0.835 $X2=0
+ $Y2=0
cc_79 N_A_N_c_73_n N_A_27_112#_c_295_n 0.00228716f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_80 N_A_N_c_74_n N_A_27_112#_c_295_n 0.0273182f $X=0.29 $Y=1.465 $X2=0 $Y2=0
cc_81 N_A_N_M1005_g N_A_27_112#_c_296_n 0.00420609f $X=0.495 $Y=0.835 $X2=0
+ $Y2=0
cc_82 N_A_N_c_73_n N_A_27_112#_c_296_n 0.00673346f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_83 N_A_N_c_74_n N_A_27_112#_c_296_n 0.0360322f $X=0.29 $Y=1.465 $X2=0 $Y2=0
cc_84 N_A_N_c_73_n N_A_27_112#_c_301_n 0.0314022f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_85 N_A_N_c_74_n N_A_27_112#_c_301_n 0.0265948f $X=0.29 $Y=1.465 $X2=0 $Y2=0
cc_86 N_A_N_c_73_n N_VPWR_c_375_n 0.00280117f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_87 N_A_N_c_73_n N_VPWR_c_384_n 0.00393265f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_88 N_A_N_c_73_n N_VPWR_c_374_n 0.00462577f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_89 N_A_N_M1005_g N_X_c_428_n 7.4905e-19 $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_90 N_A_N_c_73_n X 2.15414e-19 $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_91 N_A_N_M1005_g N_VGND_c_465_n 0.00430723f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_92 N_A_N_M1005_g N_VGND_c_467_n 0.0043356f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_93 N_A_N_M1005_g N_VGND_c_470_n 0.00487769f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_94 N_A_186_48#_c_109_n N_D_c_205_n 0.0263411f $X=1.5 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_95 N_A_186_48#_c_102_n N_D_c_205_n 0.00369938f $X=1.695 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_96 N_A_186_48#_c_103_n N_D_c_205_n 0.00118632f $X=3.74 $Y=1.045 $X2=-0.19
+ $Y2=-0.245
cc_97 N_A_186_48#_c_118_p N_D_c_205_n 0.0122189f $X=3.46 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_98 N_A_186_48#_c_105_n N_D_c_205_n 0.00208763f $X=1.56 $Y=1.465 $X2=-0.19
+ $Y2=-0.245
cc_99 N_A_186_48#_c_107_n N_D_c_205_n 0.017885f $X=1.5 $Y=1.532 $X2=-0.19
+ $Y2=-0.245
cc_100 N_A_186_48#_M1011_g N_D_M1001_g 0.00908327f $X=1.435 $Y=0.74 $X2=0 $Y2=0
cc_101 N_A_186_48#_c_103_n N_D_M1001_g 0.0156497f $X=3.74 $Y=1.045 $X2=0 $Y2=0
cc_102 N_A_186_48#_c_106_n N_D_M1001_g 0.00418176f $X=1.587 $Y=1.3 $X2=0 $Y2=0
cc_103 N_A_186_48#_c_107_n N_D_M1001_g 0.00120051f $X=1.5 $Y=1.532 $X2=0 $Y2=0
cc_104 N_A_186_48#_c_103_n N_D_c_207_n 0.0202397f $X=3.74 $Y=1.045 $X2=0 $Y2=0
cc_105 N_A_186_48#_c_118_p N_D_c_207_n 0.0215009f $X=3.46 $Y=2.035 $X2=0 $Y2=0
cc_106 N_A_186_48#_c_105_n N_D_c_207_n 0.032015f $X=1.56 $Y=1.465 $X2=0 $Y2=0
cc_107 N_A_186_48#_c_107_n N_D_c_207_n 3.17162e-19 $X=1.5 $Y=1.532 $X2=0 $Y2=0
cc_108 N_A_186_48#_c_103_n N_C_c_236_n 0.00118651f $X=3.74 $Y=1.045 $X2=-0.19
+ $Y2=-0.245
cc_109 N_A_186_48#_c_118_p N_C_c_236_n 0.0125786f $X=3.46 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_110 N_A_186_48#_c_103_n N_C_M1000_g 0.0155906f $X=3.74 $Y=1.045 $X2=0 $Y2=0
cc_111 N_A_186_48#_c_103_n N_C_c_238_n 0.0202359f $X=3.74 $Y=1.045 $X2=0 $Y2=0
cc_112 N_A_186_48#_c_118_p N_C_c_238_n 0.0231626f $X=3.46 $Y=2.035 $X2=0 $Y2=0
cc_113 N_A_186_48#_c_103_n N_B_M1004_g 0.0164071f $X=3.74 $Y=1.045 $X2=0 $Y2=0
cc_114 N_A_186_48#_c_104_n N_B_M1004_g 0.00282462f $X=3.905 $Y=0.515 $X2=0 $Y2=0
cc_115 N_A_186_48#_c_103_n N_B_c_264_n 0.00118914f $X=3.74 $Y=1.045 $X2=0 $Y2=0
cc_116 N_A_186_48#_c_118_p N_B_c_264_n 0.0124926f $X=3.46 $Y=2.035 $X2=0 $Y2=0
cc_117 N_A_186_48#_c_103_n N_B_c_265_n 0.0249816f $X=3.74 $Y=1.045 $X2=0 $Y2=0
cc_118 N_A_186_48#_c_118_p N_B_c_265_n 0.0272543f $X=3.46 $Y=2.035 $X2=0 $Y2=0
cc_119 N_A_186_48#_c_103_n N_A_27_112#_M1007_g 0.0131028f $X=3.74 $Y=1.045 $X2=0
+ $Y2=0
cc_120 N_A_186_48#_c_104_n N_A_27_112#_M1007_g 0.0139597f $X=3.905 $Y=0.515
+ $X2=0 $Y2=0
cc_121 N_A_186_48#_c_103_n N_A_27_112#_c_292_n 0.00415604f $X=3.74 $Y=1.045
+ $X2=0 $Y2=0
cc_122 N_A_186_48#_c_118_p N_A_27_112#_c_292_n 0.00292652f $X=3.46 $Y=2.035
+ $X2=0 $Y2=0
cc_123 N_A_186_48#_M1003_g N_A_27_112#_c_293_n 5.13233e-19 $X=1.005 $Y=0.74
+ $X2=0 $Y2=0
cc_124 N_A_186_48#_M1003_g N_A_27_112#_c_294_n 0.00156766f $X=1.005 $Y=0.74
+ $X2=0 $Y2=0
cc_125 N_A_186_48#_M1003_g N_A_27_112#_c_296_n 0.00275641f $X=1.005 $Y=0.74
+ $X2=0 $Y2=0
cc_126 N_A_186_48#_c_108_n N_A_27_112#_c_296_n 0.00140973f $X=1.05 $Y=1.765
+ $X2=0 $Y2=0
cc_127 N_A_186_48#_c_107_n N_A_27_112#_c_296_n 0.00272225f $X=1.5 $Y=1.532 $X2=0
+ $Y2=0
cc_128 N_A_186_48#_M1002_d N_A_27_112#_c_324_n 0.006278f $X=2.195 $Y=1.84 $X2=0
+ $Y2=0
cc_129 N_A_186_48#_M1006_d N_A_27_112#_c_324_n 0.00671576f $X=3.29 $Y=1.84 $X2=0
+ $Y2=0
cc_130 N_A_186_48#_c_108_n N_A_27_112#_c_324_n 0.0147359f $X=1.05 $Y=1.765 $X2=0
+ $Y2=0
cc_131 N_A_186_48#_c_109_n N_A_27_112#_c_324_n 0.016816f $X=1.5 $Y=1.765 $X2=0
+ $Y2=0
cc_132 N_A_186_48#_c_153_p N_A_27_112#_c_324_n 0.0119962f $X=1.78 $Y=2.075 $X2=0
+ $Y2=0
cc_133 N_A_186_48#_c_118_p N_A_27_112#_c_324_n 0.107165f $X=3.46 $Y=2.035 $X2=0
+ $Y2=0
cc_134 N_A_186_48#_c_108_n N_A_27_112#_c_301_n 0.00749533f $X=1.05 $Y=1.765
+ $X2=0 $Y2=0
cc_135 N_A_186_48#_c_103_n N_A_27_112#_c_297_n 0.0243261f $X=3.74 $Y=1.045 $X2=0
+ $Y2=0
cc_136 N_A_186_48#_c_118_p N_A_27_112#_c_297_n 0.00112569f $X=3.46 $Y=2.035
+ $X2=0 $Y2=0
cc_137 N_A_186_48#_c_102_n N_VPWR_M1012_s 0.0022467f $X=1.695 $Y=1.95 $X2=0
+ $Y2=0
cc_138 N_A_186_48#_c_153_p N_VPWR_M1012_s 0.00361743f $X=1.78 $Y=2.075 $X2=0
+ $Y2=0
cc_139 N_A_186_48#_c_118_p N_VPWR_M1012_s 0.0109741f $X=3.46 $Y=2.035 $X2=0
+ $Y2=0
cc_140 N_A_186_48#_c_118_p N_VPWR_M1010_d 0.0139764f $X=3.46 $Y=2.035 $X2=0
+ $Y2=0
cc_141 N_A_186_48#_c_108_n N_VPWR_c_375_n 0.00956311f $X=1.05 $Y=1.765 $X2=0
+ $Y2=0
cc_142 N_A_186_48#_c_109_n N_VPWR_c_375_n 0.00114115f $X=1.5 $Y=1.765 $X2=0
+ $Y2=0
cc_143 N_A_186_48#_c_108_n N_VPWR_c_376_n 0.00444681f $X=1.05 $Y=1.765 $X2=0
+ $Y2=0
cc_144 N_A_186_48#_c_109_n N_VPWR_c_376_n 0.00461464f $X=1.5 $Y=1.765 $X2=0
+ $Y2=0
cc_145 N_A_186_48#_c_109_n N_VPWR_c_377_n 0.00765649f $X=1.5 $Y=1.765 $X2=0
+ $Y2=0
cc_146 N_A_186_48#_c_108_n N_VPWR_c_374_n 0.00432688f $X=1.05 $Y=1.765 $X2=0
+ $Y2=0
cc_147 N_A_186_48#_c_109_n N_VPWR_c_374_n 0.00456645f $X=1.5 $Y=1.765 $X2=0
+ $Y2=0
cc_148 N_A_186_48#_M1003_g N_X_c_428_n 0.00909182f $X=1.005 $Y=0.74 $X2=0 $Y2=0
cc_149 N_A_186_48#_M1011_g N_X_c_428_n 0.0132513f $X=1.435 $Y=0.74 $X2=0 $Y2=0
cc_150 N_A_186_48#_c_171_p N_X_c_428_n 0.0113177f $X=1.78 $Y=1.045 $X2=0 $Y2=0
cc_151 N_A_186_48#_M1003_g N_X_c_429_n 0.00331189f $X=1.005 $Y=0.74 $X2=0 $Y2=0
cc_152 N_A_186_48#_c_108_n N_X_c_429_n 0.00140832f $X=1.05 $Y=1.765 $X2=0 $Y2=0
cc_153 N_A_186_48#_M1011_g N_X_c_429_n 0.00142748f $X=1.435 $Y=0.74 $X2=0 $Y2=0
cc_154 N_A_186_48#_c_109_n N_X_c_429_n 4.17329e-19 $X=1.5 $Y=1.765 $X2=0 $Y2=0
cc_155 N_A_186_48#_c_102_n N_X_c_429_n 0.00807649f $X=1.695 $Y=1.95 $X2=0 $Y2=0
cc_156 N_A_186_48#_c_105_n N_X_c_429_n 0.0238617f $X=1.56 $Y=1.465 $X2=0 $Y2=0
cc_157 N_A_186_48#_c_106_n N_X_c_429_n 0.00718069f $X=1.587 $Y=1.3 $X2=0 $Y2=0
cc_158 N_A_186_48#_c_107_n N_X_c_429_n 0.0201326f $X=1.5 $Y=1.532 $X2=0 $Y2=0
cc_159 N_A_186_48#_M1003_g N_X_c_430_n 0.00225198f $X=1.005 $Y=0.74 $X2=0 $Y2=0
cc_160 N_A_186_48#_M1011_g N_X_c_430_n 0.00339002f $X=1.435 $Y=0.74 $X2=0 $Y2=0
cc_161 N_A_186_48#_c_107_n N_X_c_430_n 0.00199986f $X=1.5 $Y=1.532 $X2=0 $Y2=0
cc_162 N_A_186_48#_c_108_n X 0.00725312f $X=1.05 $Y=1.765 $X2=0 $Y2=0
cc_163 N_A_186_48#_c_109_n X 0.00431584f $X=1.5 $Y=1.765 $X2=0 $Y2=0
cc_164 N_A_186_48#_c_102_n X 0.00566346f $X=1.695 $Y=1.95 $X2=0 $Y2=0
cc_165 N_A_186_48#_c_105_n X 0.00319041f $X=1.56 $Y=1.465 $X2=0 $Y2=0
cc_166 N_A_186_48#_c_107_n X 0.00848106f $X=1.5 $Y=1.532 $X2=0 $Y2=0
cc_167 N_A_186_48#_c_103_n N_VGND_M1011_d 0.00478095f $X=3.74 $Y=1.045 $X2=0
+ $Y2=0
cc_168 N_A_186_48#_c_171_p N_VGND_M1011_d 0.00472321f $X=1.78 $Y=1.045 $X2=0
+ $Y2=0
cc_169 N_A_186_48#_M1003_g N_VGND_c_465_n 0.00603022f $X=1.005 $Y=0.74 $X2=0
+ $Y2=0
cc_170 N_A_186_48#_M1011_g N_VGND_c_466_n 0.00456117f $X=1.435 $Y=0.74 $X2=0
+ $Y2=0
cc_171 N_A_186_48#_c_103_n N_VGND_c_466_n 0.0264272f $X=3.74 $Y=1.045 $X2=0
+ $Y2=0
cc_172 N_A_186_48#_c_171_p N_VGND_c_466_n 0.0153275f $X=1.78 $Y=1.045 $X2=0
+ $Y2=0
cc_173 N_A_186_48#_c_105_n N_VGND_c_466_n 0.00168337f $X=1.56 $Y=1.465 $X2=0
+ $Y2=0
cc_174 N_A_186_48#_c_107_n N_VGND_c_466_n 7.53724e-19 $X=1.5 $Y=1.532 $X2=0
+ $Y2=0
cc_175 N_A_186_48#_M1003_g N_VGND_c_468_n 0.00434272f $X=1.005 $Y=0.74 $X2=0
+ $Y2=0
cc_176 N_A_186_48#_M1011_g N_VGND_c_468_n 0.00434272f $X=1.435 $Y=0.74 $X2=0
+ $Y2=0
cc_177 N_A_186_48#_c_104_n N_VGND_c_469_n 0.0145639f $X=3.905 $Y=0.515 $X2=0
+ $Y2=0
cc_178 N_A_186_48#_M1003_g N_VGND_c_470_n 0.00825283f $X=1.005 $Y=0.74 $X2=0
+ $Y2=0
cc_179 N_A_186_48#_M1011_g N_VGND_c_470_n 0.00822601f $X=1.435 $Y=0.74 $X2=0
+ $Y2=0
cc_180 N_A_186_48#_c_104_n N_VGND_c_470_n 0.0119984f $X=3.905 $Y=0.515 $X2=0
+ $Y2=0
cc_181 N_A_186_48#_c_103_n A_459_74# 0.0048076f $X=3.74 $Y=1.045 $X2=-0.19
+ $Y2=-0.245
cc_182 N_A_186_48#_c_103_n A_537_74# 0.0107783f $X=3.74 $Y=1.045 $X2=-0.19
+ $Y2=-0.245
cc_183 N_A_186_48#_c_103_n A_645_74# 0.0107783f $X=3.74 $Y=1.045 $X2=-0.19
+ $Y2=-0.245
cc_184 N_D_c_205_n N_C_c_236_n 0.0558997f $X=2.12 $Y=1.765 $X2=-0.19 $Y2=-0.245
cc_185 N_D_c_207_n N_C_c_236_n 0.00173456f $X=2.13 $Y=1.515 $X2=-0.19 $Y2=-0.245
cc_186 N_D_M1001_g N_C_M1000_g 0.0614519f $X=2.22 $Y=0.74 $X2=0 $Y2=0
cc_187 N_D_c_205_n N_C_c_238_n 0.00129012f $X=2.12 $Y=1.765 $X2=0 $Y2=0
cc_188 N_D_c_207_n N_C_c_238_n 0.0277336f $X=2.13 $Y=1.515 $X2=0 $Y2=0
cc_189 N_D_c_205_n N_A_27_112#_c_324_n 0.012707f $X=2.12 $Y=1.765 $X2=0 $Y2=0
cc_190 N_D_c_205_n N_VPWR_c_377_n 0.00750276f $X=2.12 $Y=1.765 $X2=0 $Y2=0
cc_191 N_D_c_205_n N_VPWR_c_381_n 0.0049405f $X=2.12 $Y=1.765 $X2=0 $Y2=0
cc_192 N_D_c_205_n N_VPWR_c_374_n 0.00508379f $X=2.12 $Y=1.765 $X2=0 $Y2=0
cc_193 N_D_M1001_g N_VGND_c_466_n 0.0145292f $X=2.22 $Y=0.74 $X2=0 $Y2=0
cc_194 N_D_M1001_g N_VGND_c_469_n 0.00398535f $X=2.22 $Y=0.74 $X2=0 $Y2=0
cc_195 N_D_M1001_g N_VGND_c_470_n 0.00787244f $X=2.22 $Y=0.74 $X2=0 $Y2=0
cc_196 N_C_M1000_g N_B_M1004_g 0.0402276f $X=2.61 $Y=0.74 $X2=0 $Y2=0
cc_197 N_C_c_236_n N_B_c_264_n 0.0490624f $X=2.595 $Y=1.765 $X2=0 $Y2=0
cc_198 N_C_c_238_n N_B_c_264_n 6.60228e-19 $X=2.67 $Y=1.515 $X2=0 $Y2=0
cc_199 N_C_c_236_n N_B_c_265_n 0.00231399f $X=2.595 $Y=1.765 $X2=0 $Y2=0
cc_200 N_C_c_238_n N_B_c_265_n 0.03497f $X=2.67 $Y=1.515 $X2=0 $Y2=0
cc_201 N_C_c_236_n N_A_27_112#_c_324_n 0.012707f $X=2.595 $Y=1.765 $X2=0 $Y2=0
cc_202 N_C_c_236_n N_VPWR_c_378_n 0.00750276f $X=2.595 $Y=1.765 $X2=0 $Y2=0
cc_203 N_C_c_236_n N_VPWR_c_381_n 0.0049405f $X=2.595 $Y=1.765 $X2=0 $Y2=0
cc_204 N_C_c_236_n N_VPWR_c_374_n 0.00508379f $X=2.595 $Y=1.765 $X2=0 $Y2=0
cc_205 N_C_M1000_g N_VGND_c_466_n 0.00269307f $X=2.61 $Y=0.74 $X2=0 $Y2=0
cc_206 N_C_M1000_g N_VGND_c_469_n 0.00461464f $X=2.61 $Y=0.74 $X2=0 $Y2=0
cc_207 N_C_M1000_g N_VGND_c_470_n 0.00910057f $X=2.61 $Y=0.74 $X2=0 $Y2=0
cc_208 N_B_M1004_g N_A_27_112#_M1007_g 0.0370849f $X=3.15 $Y=0.74 $X2=0 $Y2=0
cc_209 N_B_c_264_n N_A_27_112#_c_292_n 0.0538299f $X=3.215 $Y=1.765 $X2=0 $Y2=0
cc_210 N_B_c_265_n N_A_27_112#_c_292_n 0.00130265f $X=3.24 $Y=1.515 $X2=0 $Y2=0
cc_211 N_B_c_264_n N_A_27_112#_c_324_n 0.0127845f $X=3.215 $Y=1.765 $X2=0 $Y2=0
cc_212 N_B_c_265_n N_A_27_112#_c_300_n 0.00436153f $X=3.24 $Y=1.515 $X2=0 $Y2=0
cc_213 N_B_c_264_n N_A_27_112#_c_297_n 0.00114347f $X=3.215 $Y=1.765 $X2=0 $Y2=0
cc_214 N_B_c_265_n N_A_27_112#_c_297_n 0.0213706f $X=3.24 $Y=1.515 $X2=0 $Y2=0
cc_215 N_B_c_264_n N_VPWR_c_378_n 0.00750276f $X=3.215 $Y=1.765 $X2=0 $Y2=0
cc_216 N_B_c_264_n N_VPWR_c_383_n 0.0049405f $X=3.215 $Y=1.765 $X2=0 $Y2=0
cc_217 N_B_c_264_n N_VPWR_c_374_n 0.00508379f $X=3.215 $Y=1.765 $X2=0 $Y2=0
cc_218 N_B_M1004_g N_VGND_c_469_n 0.00461464f $X=3.15 $Y=0.74 $X2=0 $Y2=0
cc_219 N_B_M1004_g N_VGND_c_470_n 0.00911376f $X=3.15 $Y=0.74 $X2=0 $Y2=0
cc_220 N_A_27_112#_c_296_n N_VPWR_M1008_d 0.00128827f $X=0.71 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_221 N_A_27_112#_c_324_n N_VPWR_M1008_d 0.00592885f $X=3.815 $Y=2.455
+ $X2=-0.19 $Y2=-0.245
cc_222 N_A_27_112#_c_301_n N_VPWR_M1008_d 0.00795497f $X=0.28 $Y=2.115 $X2=-0.19
+ $Y2=-0.245
cc_223 N_A_27_112#_c_324_n N_VPWR_M1012_s 0.00874987f $X=3.815 $Y=2.455 $X2=0
+ $Y2=0
cc_224 N_A_27_112#_c_324_n N_VPWR_M1010_d 0.00869819f $X=3.815 $Y=2.455 $X2=0
+ $Y2=0
cc_225 N_A_27_112#_c_324_n N_VPWR_M1013_d 0.00966782f $X=3.815 $Y=2.455 $X2=0
+ $Y2=0
cc_226 N_A_27_112#_c_300_n N_VPWR_M1013_d 0.0231221f $X=3.9 $Y=2.37 $X2=0 $Y2=0
cc_227 N_A_27_112#_c_324_n N_VPWR_c_375_n 0.00999279f $X=3.815 $Y=2.455 $X2=0
+ $Y2=0
cc_228 N_A_27_112#_c_301_n N_VPWR_c_375_n 0.0126312f $X=0.28 $Y=2.115 $X2=0
+ $Y2=0
cc_229 N_A_27_112#_c_324_n N_VPWR_c_377_n 0.0260584f $X=3.815 $Y=2.455 $X2=0
+ $Y2=0
cc_230 N_A_27_112#_c_324_n N_VPWR_c_378_n 0.0260584f $X=3.815 $Y=2.455 $X2=0
+ $Y2=0
cc_231 N_A_27_112#_c_292_n N_VPWR_c_380_n 0.0108539f $X=3.705 $Y=1.765 $X2=0
+ $Y2=0
cc_232 N_A_27_112#_c_324_n N_VPWR_c_380_n 0.0117196f $X=3.815 $Y=2.455 $X2=0
+ $Y2=0
cc_233 N_A_27_112#_c_292_n N_VPWR_c_383_n 0.0049405f $X=3.705 $Y=1.765 $X2=0
+ $Y2=0
cc_234 N_A_27_112#_c_301_n N_VPWR_c_384_n 0.00671799f $X=0.28 $Y=2.115 $X2=0
+ $Y2=0
cc_235 N_A_27_112#_c_292_n N_VPWR_c_374_n 0.00508379f $X=3.705 $Y=1.765 $X2=0
+ $Y2=0
cc_236 N_A_27_112#_c_324_n N_VPWR_c_374_n 0.0793995f $X=3.815 $Y=2.455 $X2=0
+ $Y2=0
cc_237 N_A_27_112#_c_301_n N_VPWR_c_374_n 0.0184551f $X=0.28 $Y=2.115 $X2=0
+ $Y2=0
cc_238 N_A_27_112#_c_324_n N_X_M1009_d 0.00556049f $X=3.815 $Y=2.455 $X2=0 $Y2=0
cc_239 N_A_27_112#_c_293_n N_X_c_428_n 0.00441257f $X=0.28 $Y=0.835 $X2=0 $Y2=0
cc_240 N_A_27_112#_c_294_n N_X_c_428_n 0.0101363f $X=0.625 $Y=1.045 $X2=0 $Y2=0
cc_241 N_A_27_112#_c_296_n N_X_c_429_n 0.035856f $X=0.71 $Y=1.95 $X2=0 $Y2=0
cc_242 N_A_27_112#_c_296_n X 0.00697858f $X=0.71 $Y=1.95 $X2=0 $Y2=0
cc_243 N_A_27_112#_c_324_n X 0.0203978f $X=3.815 $Y=2.455 $X2=0 $Y2=0
cc_244 N_A_27_112#_c_301_n X 0.0150414f $X=0.28 $Y=2.115 $X2=0 $Y2=0
cc_245 N_A_27_112#_c_294_n N_VGND_M1005_d 0.00376661f $X=0.625 $Y=1.045
+ $X2=-0.19 $Y2=-0.245
cc_246 N_A_27_112#_c_293_n N_VGND_c_465_n 0.0096883f $X=0.28 $Y=0.835 $X2=0
+ $Y2=0
cc_247 N_A_27_112#_c_294_n N_VGND_c_465_n 0.0151472f $X=0.625 $Y=1.045 $X2=0
+ $Y2=0
cc_248 N_A_27_112#_c_293_n N_VGND_c_467_n 0.00806442f $X=0.28 $Y=0.835 $X2=0
+ $Y2=0
cc_249 N_A_27_112#_M1007_g N_VGND_c_469_n 0.00434272f $X=3.69 $Y=0.74 $X2=0
+ $Y2=0
cc_250 N_A_27_112#_M1007_g N_VGND_c_470_n 0.00826337f $X=3.69 $Y=0.74 $X2=0
+ $Y2=0
cc_251 N_A_27_112#_c_293_n N_VGND_c_470_n 0.0105742f $X=0.28 $Y=0.835 $X2=0
+ $Y2=0
cc_252 N_X_c_428_n N_VGND_c_465_n 0.0164982f $X=1.22 $Y=0.515 $X2=0 $Y2=0
cc_253 N_X_c_428_n N_VGND_c_466_n 0.0173772f $X=1.22 $Y=0.515 $X2=0 $Y2=0
cc_254 N_X_c_428_n N_VGND_c_468_n 0.0144922f $X=1.22 $Y=0.515 $X2=0 $Y2=0
cc_255 N_X_c_428_n N_VGND_c_470_n 0.0118826f $X=1.22 $Y=0.515 $X2=0 $Y2=0
