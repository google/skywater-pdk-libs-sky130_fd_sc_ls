* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
M1000 a_27_368# A3 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=1.7808e+12p pd=1.438e+07u as=1.0752e+12p ps=8.64e+06u
M1001 Y B1 a_27_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=0p ps=0u
M1002 Y B1 VGND VNB nshort w=740000u l=150000u
+  ad=7.548e+11p pd=5e+06u as=5.217e+11p ps=4.37e+06u
M1003 a_27_368# B1 Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_27_368# A2 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y A1 a_200_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=4.773e+11p ps=4.25e+06u
M1006 VPWR A1 a_27_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR A3 a_27_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND A3 a_114_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=4.662e+11p ps=4.22e+06u
M1009 a_27_368# A1 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_114_74# A2 a_200_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR A2 a_27_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_114_74# A3 VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_200_74# A2 a_114_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_200_74# A1 Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
