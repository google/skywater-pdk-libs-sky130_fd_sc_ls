* File: sky130_fd_sc_ls__a311o_2.pxi.spice
* Created: Fri Aug 28 12:57:32 2020
* 
x_PM_SKY130_FD_SC_LS__A311O_2%A_21_270# N_A_21_270#_M1012_d N_A_21_270#_M1008_d
+ N_A_21_270#_M1002_d N_A_21_270#_c_93_n N_A_21_270#_M1007_g N_A_21_270#_M1003_g
+ N_A_21_270#_c_82_n N_A_21_270#_c_83_n N_A_21_270#_c_84_n N_A_21_270#_c_96_n
+ N_A_21_270#_M1010_g N_A_21_270#_M1009_g N_A_21_270#_c_86_n N_A_21_270#_c_87_n
+ N_A_21_270#_c_88_n N_A_21_270#_c_159_p N_A_21_270#_c_99_n N_A_21_270#_c_89_n
+ N_A_21_270#_c_113_p N_A_21_270#_c_209_p N_A_21_270#_c_101_n N_A_21_270#_c_90_n
+ N_A_21_270#_c_91_n N_A_21_270#_c_102_n N_A_21_270#_c_103_n N_A_21_270#_c_92_n
+ N_A_21_270#_c_110_p N_A_21_270#_c_131_p PM_SKY130_FD_SC_LS__A311O_2%A_21_270#
x_PM_SKY130_FD_SC_LS__A311O_2%A3 N_A3_c_230_n N_A3_c_235_n N_A3_M1013_g
+ N_A3_M1006_g A3 N_A3_c_232_n N_A3_c_233_n PM_SKY130_FD_SC_LS__A311O_2%A3
x_PM_SKY130_FD_SC_LS__A311O_2%A2 N_A2_M1001_g N_A2_c_271_n N_A2_M1000_g A2
+ PM_SKY130_FD_SC_LS__A311O_2%A2
x_PM_SKY130_FD_SC_LS__A311O_2%A1 N_A1_M1012_g N_A1_c_301_n N_A1_M1011_g A1
+ PM_SKY130_FD_SC_LS__A311O_2%A1
x_PM_SKY130_FD_SC_LS__A311O_2%B1 N_B1_M1004_g N_B1_c_334_n N_B1_c_338_n
+ N_B1_M1005_g B1 B1 N_B1_c_336_n PM_SKY130_FD_SC_LS__A311O_2%B1
x_PM_SKY130_FD_SC_LS__A311O_2%C1 N_C1_c_375_n N_C1_M1002_g N_C1_M1008_g
+ N_C1_c_372_n C1 N_C1_c_374_n PM_SKY130_FD_SC_LS__A311O_2%C1
x_PM_SKY130_FD_SC_LS__A311O_2%VPWR N_VPWR_M1007_d N_VPWR_M1010_d N_VPWR_M1000_d
+ N_VPWR_c_405_n N_VPWR_c_406_n N_VPWR_c_407_n N_VPWR_c_408_n VPWR
+ N_VPWR_c_409_n N_VPWR_c_410_n N_VPWR_c_404_n N_VPWR_c_412_n N_VPWR_c_413_n
+ PM_SKY130_FD_SC_LS__A311O_2%VPWR
x_PM_SKY130_FD_SC_LS__A311O_2%X N_X_M1003_s N_X_M1007_s N_X_c_461_n N_X_c_462_n
+ X PM_SKY130_FD_SC_LS__A311O_2%X
x_PM_SKY130_FD_SC_LS__A311O_2%A_330_392# N_A_330_392#_M1013_d
+ N_A_330_392#_M1011_d N_A_330_392#_c_488_n N_A_330_392#_c_484_n
+ N_A_330_392#_c_491_n N_A_330_392#_c_492_n N_A_330_392#_c_485_n
+ PM_SKY130_FD_SC_LS__A311O_2%A_330_392#
x_PM_SKY130_FD_SC_LS__A311O_2%VGND N_VGND_M1003_d N_VGND_M1009_d N_VGND_M1004_d
+ N_VGND_c_518_n N_VGND_c_519_n N_VGND_c_520_n N_VGND_c_521_n N_VGND_c_522_n
+ N_VGND_c_523_n N_VGND_c_524_n N_VGND_c_525_n N_VGND_c_526_n VGND
+ N_VGND_c_527_n N_VGND_c_528_n PM_SKY130_FD_SC_LS__A311O_2%VGND
cc_1 VNB N_A_21_270#_M1003_g 0.0298485f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=0.74
cc_2 VNB N_A_21_270#_c_82_n 0.0121213f $X=-0.19 $Y=-0.245 $X2=0.965 $Y2=1.425
cc_3 VNB N_A_21_270#_c_83_n 0.0134848f $X=-0.19 $Y=-0.245 $X2=0.755 $Y2=1.425
cc_4 VNB N_A_21_270#_c_84_n 0.00777664f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=1.675
cc_5 VNB N_A_21_270#_M1009_g 0.0239659f $X=-0.19 $Y=-0.245 $X2=1.11 $Y2=0.74
cc_6 VNB N_A_21_270#_c_86_n 0.0418684f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.515
cc_7 VNB N_A_21_270#_c_87_n 0.00694108f $X=-0.19 $Y=-0.245 $X2=1.075 $Y2=1.425
cc_8 VNB N_A_21_270#_c_88_n 0.00930993f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.515
cc_9 VNB N_A_21_270#_c_89_n 0.00482179f $X=-0.19 $Y=-0.245 $X2=1.25 $Y2=1.95
cc_10 VNB N_A_21_270#_c_90_n 0.00317749f $X=-0.19 $Y=-0.245 $X2=2.815 $Y2=0.515
cc_11 VNB N_A_21_270#_c_91_n 0.00752401f $X=-0.19 $Y=-0.245 $X2=3.71 $Y2=1.005
cc_12 VNB N_A_21_270#_c_92_n 0.0246973f $X=-0.19 $Y=-0.245 $X2=3.875 $Y2=0.515
cc_13 VNB N_A3_c_230_n 0.00374859f $X=-0.19 $Y=-0.245 $X2=3.735 $Y2=0.37
cc_14 VNB N_A3_M1006_g 0.0197804f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A3_c_232_n 0.0299527f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=1.35
cc_16 VNB N_A3_c_233_n 0.00451054f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=0.74
cc_17 VNB N_A2_M1001_g 0.030979f $X=-0.19 $Y=-0.245 $X2=3.72 $Y2=1.96
cc_18 VNB N_A2_c_271_n 0.019683f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB A2 0.00224383f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A1_M1012_g 0.0339807f $X=-0.19 $Y=-0.245 $X2=3.72 $Y2=1.96
cc_21 VNB N_A1_c_301_n 0.0196759f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB A1 0.00224095f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_B1_M1004_g 0.0214481f $X=-0.19 $Y=-0.245 $X2=3.72 $Y2=1.96
cc_24 VNB N_B1_c_334_n 0.00318739f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB B1 0.00614412f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=2.4
cc_26 VNB N_B1_c_336_n 0.0284591f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=0.74
cc_27 VNB N_C1_M1008_g 0.0417252f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_C1_c_372_n 0.00592792f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB C1 0.00841732f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.765
cc_30 VNB N_C1_c_374_n 0.0366622f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=1.35
cc_31 VNB N_VPWR_c_404_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=1.557
cc_32 VNB N_X_c_461_n 0.00150157f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.765
cc_33 VNB N_X_c_462_n 0.00239859f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=2.4
cc_34 VNB N_VGND_c_518_n 0.043308f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=2.4
cc_35 VNB N_VGND_c_519_n 0.00718188f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_520_n 0.00685406f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=1.675
cc_37 VNB N_VGND_c_521_n 0.0116899f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=2.4
cc_38 VNB N_VGND_c_522_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=1.11 $Y2=1.35
cc_39 VNB N_VGND_c_523_n 0.019013f $X=-0.19 $Y=-0.245 $X2=1.11 $Y2=0.74
cc_40 VNB N_VGND_c_524_n 0.00750435f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_525_n 0.0457514f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.557
cc_42 VNB N_VGND_c_526_n 0.0069273f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=1.557
cc_43 VNB N_VGND_c_527_n 0.0244021f $X=-0.19 $Y=-0.245 $X2=2.815 $Y2=0.515
cc_44 VNB N_VGND_c_528_n 0.282418f $X=-0.19 $Y=-0.245 $X2=2.815 $Y2=0.515
cc_45 VPB N_A_21_270#_c_93_n 0.0168943f $X=-0.19 $Y=1.66 $X2=0.605 $Y2=1.765
cc_46 VPB N_A_21_270#_c_83_n 0.00788081f $X=-0.19 $Y=1.66 $X2=0.755 $Y2=1.425
cc_47 VPB N_A_21_270#_c_84_n 7.0174e-19 $X=-0.19 $Y=1.66 $X2=1.055 $Y2=1.675
cc_48 VPB N_A_21_270#_c_96_n 0.0210041f $X=-0.19 $Y=1.66 $X2=1.055 $Y2=1.765
cc_49 VPB N_A_21_270#_c_86_n 0.0138413f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=1.515
cc_50 VPB N_A_21_270#_c_88_n 0.0234375f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.515
cc_51 VPB N_A_21_270#_c_99_n 0.0127531f $X=-0.19 $Y=1.66 $X2=0.435 $Y2=2.315
cc_52 VPB N_A_21_270#_c_89_n 0.00319924f $X=-0.19 $Y=1.66 $X2=1.25 $Y2=1.95
cc_53 VPB N_A_21_270#_c_101_n 0.0269422f $X=-0.19 $Y=1.66 $X2=3.705 $Y2=2.035
cc_54 VPB N_A_21_270#_c_102_n 0.0100184f $X=-0.19 $Y=1.66 $X2=3.87 $Y2=2.12
cc_55 VPB N_A_21_270#_c_103_n 0.0360166f $X=-0.19 $Y=1.66 $X2=3.87 $Y2=2.815
cc_56 VPB N_A3_c_230_n 0.00737631f $X=-0.19 $Y=1.66 $X2=3.735 $Y2=0.37
cc_57 VPB N_A3_c_235_n 0.0229699f $X=-0.19 $Y=1.66 $X2=3.72 $Y2=1.96
cc_58 VPB N_A3_c_233_n 0.00193345f $X=-0.19 $Y=1.66 $X2=0.68 $Y2=0.74
cc_59 VPB N_A2_c_271_n 0.038398f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB A2 0.00138199f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_A1_c_301_n 0.0383607f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB A1 0.00138199f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_B1_c_334_n 0.00625192f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_B1_c_338_n 0.0219876f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB B1 0.00419635f $X=-0.19 $Y=1.66 $X2=0.605 $Y2=2.4
cc_66 VPB N_C1_c_375_n 0.0209993f $X=-0.19 $Y=1.66 $X2=2.655 $Y2=0.37
cc_67 VPB N_C1_c_372_n 0.0142876f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB C1 0.00850711f $X=-0.19 $Y=1.66 $X2=0.605 $Y2=1.765
cc_69 VPB N_C1_c_374_n 0.0246274f $X=-0.19 $Y=1.66 $X2=0.68 $Y2=1.35
cc_70 VPB N_VPWR_c_405_n 0.0152004f $X=-0.19 $Y=1.66 $X2=0.605 $Y2=1.765
cc_71 VPB N_VPWR_c_406_n 0.0248846f $X=-0.19 $Y=1.66 $X2=0.605 $Y2=2.4
cc_72 VPB N_VPWR_c_407_n 0.00591275f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_408_n 0.0187618f $X=-0.19 $Y=1.66 $X2=0.755 $Y2=1.425
cc_74 VPB N_VPWR_c_409_n 0.0177589f $X=-0.19 $Y=1.66 $X2=1.055 $Y2=2.4
cc_75 VPB N_VPWR_c_410_n 0.0491146f $X=-0.19 $Y=1.66 $X2=0.605 $Y2=1.557
cc_76 VPB N_VPWR_c_404_n 0.0892858f $X=-0.19 $Y=1.66 $X2=0.68 $Y2=1.557
cc_77 VPB N_VPWR_c_412_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_413_n 0.0222783f $X=-0.19 $Y=1.66 $X2=1.25 $Y2=1.09
cc_79 VPB N_A_330_392#_c_484_n 0.00290264f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 VPB N_A_330_392#_c_485_n 0.00290264f $X=-0.19 $Y=1.66 $X2=0.68 $Y2=0.74
cc_81 N_A_21_270#_c_84_n N_A3_c_230_n 0.00476241f $X=1.055 $Y=1.675 $X2=0 $Y2=0
cc_82 N_A_21_270#_c_96_n N_A3_c_230_n 0.00301393f $X=1.055 $Y=1.765 $X2=0 $Y2=0
cc_83 N_A_21_270#_c_89_n N_A3_c_230_n 0.00357281f $X=1.25 $Y=1.95 $X2=0 $Y2=0
cc_84 N_A_21_270#_c_96_n N_A3_c_235_n 0.0272987f $X=1.055 $Y=1.765 $X2=0 $Y2=0
cc_85 N_A_21_270#_c_89_n N_A3_c_235_n 0.00141317f $X=1.25 $Y=1.95 $X2=0 $Y2=0
cc_86 N_A_21_270#_c_101_n N_A3_c_235_n 0.0157789f $X=3.705 $Y=2.035 $X2=0 $Y2=0
cc_87 N_A_21_270#_c_110_p N_A3_c_235_n 0.00481502f $X=1.25 $Y=2.035 $X2=0 $Y2=0
cc_88 N_A_21_270#_M1009_g N_A3_M1006_g 0.0199253f $X=1.11 $Y=0.74 $X2=0 $Y2=0
cc_89 N_A_21_270#_c_89_n N_A3_M1006_g 0.00329937f $X=1.25 $Y=1.95 $X2=0 $Y2=0
cc_90 N_A_21_270#_c_113_p N_A3_M1006_g 0.0144802f $X=2.63 $Y=1.005 $X2=0 $Y2=0
cc_91 N_A_21_270#_c_84_n N_A3_c_232_n 0.0033774f $X=1.055 $Y=1.675 $X2=0 $Y2=0
cc_92 N_A_21_270#_M1009_g N_A3_c_232_n 0.0124913f $X=1.11 $Y=0.74 $X2=0 $Y2=0
cc_93 N_A_21_270#_c_89_n N_A3_c_232_n 0.00225453f $X=1.25 $Y=1.95 $X2=0 $Y2=0
cc_94 N_A_21_270#_c_113_p N_A3_c_232_n 0.0036783f $X=2.63 $Y=1.005 $X2=0 $Y2=0
cc_95 N_A_21_270#_c_101_n N_A3_c_232_n 0.00224107f $X=3.705 $Y=2.035 $X2=0 $Y2=0
cc_96 N_A_21_270#_M1009_g N_A3_c_233_n 2.03914e-19 $X=1.11 $Y=0.74 $X2=0 $Y2=0
cc_97 N_A_21_270#_c_89_n N_A3_c_233_n 0.0386594f $X=1.25 $Y=1.95 $X2=0 $Y2=0
cc_98 N_A_21_270#_c_113_p N_A3_c_233_n 0.0184565f $X=2.63 $Y=1.005 $X2=0 $Y2=0
cc_99 N_A_21_270#_c_101_n N_A3_c_233_n 0.0225571f $X=3.705 $Y=2.035 $X2=0 $Y2=0
cc_100 N_A_21_270#_c_113_p N_A2_M1001_g 0.0161078f $X=2.63 $Y=1.005 $X2=0 $Y2=0
cc_101 N_A_21_270#_c_90_n N_A2_M1001_g 0.00263562f $X=2.815 $Y=0.515 $X2=0 $Y2=0
cc_102 N_A_21_270#_c_113_p N_A2_c_271_n 8.99171e-19 $X=2.63 $Y=1.005 $X2=0 $Y2=0
cc_103 N_A_21_270#_c_101_n N_A2_c_271_n 0.0137064f $X=3.705 $Y=2.035 $X2=0 $Y2=0
cc_104 N_A_21_270#_c_113_p A2 0.0120888f $X=2.63 $Y=1.005 $X2=0 $Y2=0
cc_105 N_A_21_270#_c_101_n A2 0.0242115f $X=3.705 $Y=2.035 $X2=0 $Y2=0
cc_106 N_A_21_270#_c_113_p N_A1_M1012_g 0.0125062f $X=2.63 $Y=1.005 $X2=0 $Y2=0
cc_107 N_A_21_270#_c_90_n N_A1_M1012_g 0.0122227f $X=2.815 $Y=0.515 $X2=0 $Y2=0
cc_108 N_A_21_270#_c_131_p N_A1_M1012_g 9.09362e-19 $X=2.815 $Y=1.005 $X2=0
+ $Y2=0
cc_109 N_A_21_270#_c_101_n N_A1_c_301_n 0.0136482f $X=3.705 $Y=2.035 $X2=0 $Y2=0
cc_110 N_A_21_270#_c_131_p N_A1_c_301_n 0.0010368f $X=2.815 $Y=1.005 $X2=0 $Y2=0
cc_111 N_A_21_270#_c_113_p A1 0.00484352f $X=2.63 $Y=1.005 $X2=0 $Y2=0
cc_112 N_A_21_270#_c_101_n A1 0.0242115f $X=3.705 $Y=2.035 $X2=0 $Y2=0
cc_113 N_A_21_270#_c_131_p A1 0.00792052f $X=2.815 $Y=1.005 $X2=0 $Y2=0
cc_114 N_A_21_270#_c_90_n N_B1_M1004_g 0.00331992f $X=2.815 $Y=0.515 $X2=0 $Y2=0
cc_115 N_A_21_270#_c_91_n N_B1_M1004_g 0.0153799f $X=3.71 $Y=1.005 $X2=0 $Y2=0
cc_116 N_A_21_270#_c_92_n N_B1_M1004_g 8.17215e-19 $X=3.875 $Y=0.515 $X2=0 $Y2=0
cc_117 N_A_21_270#_c_101_n N_B1_c_338_n 0.0156212f $X=3.705 $Y=2.035 $X2=0 $Y2=0
cc_118 N_A_21_270#_c_103_n N_B1_c_338_n 0.00280486f $X=3.87 $Y=2.815 $X2=0 $Y2=0
cc_119 N_A_21_270#_c_101_n B1 0.0550228f $X=3.705 $Y=2.035 $X2=0 $Y2=0
cc_120 N_A_21_270#_c_91_n B1 0.049173f $X=3.71 $Y=1.005 $X2=0 $Y2=0
cc_121 N_A_21_270#_c_102_n B1 8.25396e-19 $X=3.87 $Y=2.12 $X2=0 $Y2=0
cc_122 N_A_21_270#_c_101_n N_B1_c_336_n 6.69993e-19 $X=3.705 $Y=2.035 $X2=0
+ $Y2=0
cc_123 N_A_21_270#_c_91_n N_B1_c_336_n 0.00437192f $X=3.71 $Y=1.005 $X2=0 $Y2=0
cc_124 N_A_21_270#_c_101_n N_C1_c_375_n 0.0117808f $X=3.705 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_125 N_A_21_270#_c_102_n N_C1_c_375_n 8.1278e-19 $X=3.87 $Y=2.12 $X2=-0.19
+ $Y2=-0.245
cc_126 N_A_21_270#_c_103_n N_C1_c_375_n 0.0151063f $X=3.87 $Y=2.815 $X2=-0.19
+ $Y2=-0.245
cc_127 N_A_21_270#_c_91_n N_C1_M1008_g 0.0131131f $X=3.71 $Y=1.005 $X2=0 $Y2=0
cc_128 N_A_21_270#_c_92_n N_C1_M1008_g 0.00850118f $X=3.875 $Y=0.515 $X2=0 $Y2=0
cc_129 N_A_21_270#_c_101_n N_C1_c_372_n 3.37059e-19 $X=3.705 $Y=2.035 $X2=0
+ $Y2=0
cc_130 N_A_21_270#_c_102_n N_C1_c_372_n 8.13785e-19 $X=3.87 $Y=2.12 $X2=0 $Y2=0
cc_131 N_A_21_270#_c_91_n C1 0.00741042f $X=3.71 $Y=1.005 $X2=0 $Y2=0
cc_132 N_A_21_270#_c_102_n C1 0.0132673f $X=3.87 $Y=2.12 $X2=0 $Y2=0
cc_133 N_A_21_270#_c_91_n N_C1_c_374_n 0.00549698f $X=3.71 $Y=1.005 $X2=0 $Y2=0
cc_134 N_A_21_270#_c_102_n N_C1_c_374_n 0.0077648f $X=3.87 $Y=2.12 $X2=0 $Y2=0
cc_135 N_A_21_270#_c_88_n N_VPWR_M1007_d 0.00662212f $X=0.27 $Y=1.515 $X2=-0.19
+ $Y2=-0.245
cc_136 N_A_21_270#_c_159_p N_VPWR_M1007_d 9.88419e-19 $X=1.165 $Y=2.315
+ $X2=-0.19 $Y2=-0.245
cc_137 N_A_21_270#_c_99_n N_VPWR_M1007_d 0.00287476f $X=0.435 $Y=2.315 $X2=-0.19
+ $Y2=-0.245
cc_138 N_A_21_270#_c_89_n N_VPWR_M1010_d 0.00205762f $X=1.25 $Y=1.95 $X2=0 $Y2=0
cc_139 N_A_21_270#_c_101_n N_VPWR_M1010_d 0.00492339f $X=3.705 $Y=2.035 $X2=0
+ $Y2=0
cc_140 N_A_21_270#_c_110_p N_VPWR_M1010_d 0.00616934f $X=1.25 $Y=2.035 $X2=0
+ $Y2=0
cc_141 N_A_21_270#_c_101_n N_VPWR_M1000_d 0.00612363f $X=3.705 $Y=2.035 $X2=0
+ $Y2=0
cc_142 N_A_21_270#_c_93_n N_VPWR_c_406_n 0.0128316f $X=0.605 $Y=1.765 $X2=0
+ $Y2=0
cc_143 N_A_21_270#_c_96_n N_VPWR_c_406_n 0.00153724f $X=1.055 $Y=1.765 $X2=0
+ $Y2=0
cc_144 N_A_21_270#_c_159_p N_VPWR_c_406_n 0.00407948f $X=1.165 $Y=2.315 $X2=0
+ $Y2=0
cc_145 N_A_21_270#_c_99_n N_VPWR_c_406_n 0.0198382f $X=0.435 $Y=2.315 $X2=0
+ $Y2=0
cc_146 N_A_21_270#_c_93_n N_VPWR_c_407_n 0.00153724f $X=0.605 $Y=1.765 $X2=0
+ $Y2=0
cc_147 N_A_21_270#_c_96_n N_VPWR_c_407_n 0.0115864f $X=1.055 $Y=1.765 $X2=0
+ $Y2=0
cc_148 N_A_21_270#_c_159_p N_VPWR_c_407_n 0.00102433f $X=1.165 $Y=2.315 $X2=0
+ $Y2=0
cc_149 N_A_21_270#_c_101_n N_VPWR_c_407_n 0.00427241f $X=3.705 $Y=2.035 $X2=0
+ $Y2=0
cc_150 N_A_21_270#_c_110_p N_VPWR_c_407_n 0.0132538f $X=1.25 $Y=2.035 $X2=0
+ $Y2=0
cc_151 N_A_21_270#_c_93_n N_VPWR_c_409_n 0.00413917f $X=0.605 $Y=1.765 $X2=0
+ $Y2=0
cc_152 N_A_21_270#_c_96_n N_VPWR_c_409_n 0.00413917f $X=1.055 $Y=1.765 $X2=0
+ $Y2=0
cc_153 N_A_21_270#_c_103_n N_VPWR_c_410_n 0.0145938f $X=3.87 $Y=2.815 $X2=0
+ $Y2=0
cc_154 N_A_21_270#_c_93_n N_VPWR_c_404_n 0.00817726f $X=0.605 $Y=1.765 $X2=0
+ $Y2=0
cc_155 N_A_21_270#_c_96_n N_VPWR_c_404_n 0.00817726f $X=1.055 $Y=1.765 $X2=0
+ $Y2=0
cc_156 N_A_21_270#_c_103_n N_VPWR_c_404_n 0.0120466f $X=3.87 $Y=2.815 $X2=0
+ $Y2=0
cc_157 N_A_21_270#_c_159_p N_X_M1007_s 0.00905546f $X=1.165 $Y=2.315 $X2=0 $Y2=0
cc_158 N_A_21_270#_M1003_g N_X_c_461_n 0.016013f $X=0.68 $Y=0.74 $X2=0 $Y2=0
cc_159 N_A_21_270#_c_82_n N_X_c_461_n 0.010131f $X=0.965 $Y=1.425 $X2=0 $Y2=0
cc_160 N_A_21_270#_c_83_n N_X_c_461_n 0.00463964f $X=0.755 $Y=1.425 $X2=0 $Y2=0
cc_161 N_A_21_270#_c_84_n N_X_c_461_n 9.79881e-19 $X=1.055 $Y=1.675 $X2=0 $Y2=0
cc_162 N_A_21_270#_M1009_g N_X_c_461_n 0.00197084f $X=1.11 $Y=0.74 $X2=0 $Y2=0
cc_163 N_A_21_270#_c_87_n N_X_c_461_n 0.00237831f $X=1.075 $Y=1.425 $X2=0 $Y2=0
cc_164 N_A_21_270#_c_88_n N_X_c_461_n 0.00947676f $X=0.27 $Y=1.515 $X2=0 $Y2=0
cc_165 N_A_21_270#_c_89_n N_X_c_461_n 0.0629389f $X=1.25 $Y=1.95 $X2=0 $Y2=0
cc_166 N_A_21_270#_M1003_g N_X_c_462_n 0.00555206f $X=0.68 $Y=0.74 $X2=0 $Y2=0
cc_167 N_A_21_270#_M1009_g N_X_c_462_n 0.00648554f $X=1.11 $Y=0.74 $X2=0 $Y2=0
cc_168 N_A_21_270#_c_93_n X 0.00609323f $X=0.605 $Y=1.765 $X2=0 $Y2=0
cc_169 N_A_21_270#_c_83_n X 0.0149968f $X=0.755 $Y=1.425 $X2=0 $Y2=0
cc_170 N_A_21_270#_c_84_n X 0.00253974f $X=1.055 $Y=1.675 $X2=0 $Y2=0
cc_171 N_A_21_270#_c_96_n X 0.00628315f $X=1.055 $Y=1.765 $X2=0 $Y2=0
cc_172 N_A_21_270#_c_88_n X 0.0399512f $X=0.27 $Y=1.515 $X2=0 $Y2=0
cc_173 N_A_21_270#_c_159_p X 0.0216202f $X=1.165 $Y=2.315 $X2=0 $Y2=0
cc_174 N_A_21_270#_c_101_n N_A_330_392#_M1013_d 0.00229612f $X=3.705 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_175 N_A_21_270#_c_101_n N_A_330_392#_M1011_d 0.00229612f $X=3.705 $Y=2.035
+ $X2=0 $Y2=0
cc_176 N_A_21_270#_c_96_n N_A_330_392#_c_488_n 7.08343e-19 $X=1.055 $Y=1.765
+ $X2=0 $Y2=0
cc_177 N_A_21_270#_c_101_n N_A_330_392#_c_488_n 0.0186962f $X=3.705 $Y=2.035
+ $X2=0 $Y2=0
cc_178 N_A_21_270#_c_110_p N_A_330_392#_c_488_n 0.00557251f $X=1.25 $Y=2.035
+ $X2=0 $Y2=0
cc_179 N_A_21_270#_c_101_n N_A_330_392#_c_491_n 0.0532125f $X=3.705 $Y=2.035
+ $X2=0 $Y2=0
cc_180 N_A_21_270#_c_101_n N_A_330_392#_c_492_n 0.0186962f $X=3.705 $Y=2.035
+ $X2=0 $Y2=0
cc_181 N_A_21_270#_c_103_n N_A_330_392#_c_492_n 0.00863451f $X=3.87 $Y=2.815
+ $X2=0 $Y2=0
cc_182 N_A_21_270#_c_103_n N_A_330_392#_c_485_n 0.0119084f $X=3.87 $Y=2.815
+ $X2=0 $Y2=0
cc_183 N_A_21_270#_c_101_n A_660_392# 0.00595227f $X=3.705 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_184 N_A_21_270#_c_89_n N_VGND_M1009_d 2.38044e-19 $X=1.25 $Y=1.95 $X2=0 $Y2=0
cc_185 N_A_21_270#_c_113_p N_VGND_M1009_d 0.00746768f $X=2.63 $Y=1.005 $X2=0
+ $Y2=0
cc_186 N_A_21_270#_c_209_p N_VGND_M1009_d 0.00102916f $X=1.335 $Y=1.005 $X2=0
+ $Y2=0
cc_187 N_A_21_270#_c_91_n N_VGND_M1004_d 0.0058594f $X=3.71 $Y=1.005 $X2=0 $Y2=0
cc_188 N_A_21_270#_M1003_g N_VGND_c_518_n 0.00647412f $X=0.68 $Y=0.74 $X2=0
+ $Y2=0
cc_189 N_A_21_270#_c_86_n N_VGND_c_518_n 0.00592994f $X=0.515 $Y=1.515 $X2=0
+ $Y2=0
cc_190 N_A_21_270#_c_88_n N_VGND_c_518_n 0.00975954f $X=0.27 $Y=1.515 $X2=0
+ $Y2=0
cc_191 N_A_21_270#_M1009_g N_VGND_c_519_n 0.00579414f $X=1.11 $Y=0.74 $X2=0
+ $Y2=0
cc_192 N_A_21_270#_c_113_p N_VGND_c_519_n 0.019079f $X=2.63 $Y=1.005 $X2=0 $Y2=0
cc_193 N_A_21_270#_c_209_p N_VGND_c_519_n 0.00838504f $X=1.335 $Y=1.005 $X2=0
+ $Y2=0
cc_194 N_A_21_270#_c_90_n N_VGND_c_520_n 0.0160784f $X=2.815 $Y=0.515 $X2=0
+ $Y2=0
cc_195 N_A_21_270#_c_91_n N_VGND_c_520_n 0.024241f $X=3.71 $Y=1.005 $X2=0 $Y2=0
cc_196 N_A_21_270#_c_92_n N_VGND_c_520_n 0.0158132f $X=3.875 $Y=0.515 $X2=0
+ $Y2=0
cc_197 N_A_21_270#_M1003_g N_VGND_c_523_n 0.00434272f $X=0.68 $Y=0.74 $X2=0
+ $Y2=0
cc_198 N_A_21_270#_M1009_g N_VGND_c_523_n 0.00434272f $X=1.11 $Y=0.74 $X2=0
+ $Y2=0
cc_199 N_A_21_270#_c_90_n N_VGND_c_525_n 0.0163488f $X=2.815 $Y=0.515 $X2=0
+ $Y2=0
cc_200 N_A_21_270#_c_92_n N_VGND_c_527_n 0.0145639f $X=3.875 $Y=0.515 $X2=0
+ $Y2=0
cc_201 N_A_21_270#_M1003_g N_VGND_c_528_n 0.00824428f $X=0.68 $Y=0.74 $X2=0
+ $Y2=0
cc_202 N_A_21_270#_M1009_g N_VGND_c_528_n 0.00821312f $X=1.11 $Y=0.74 $X2=0
+ $Y2=0
cc_203 N_A_21_270#_c_90_n N_VGND_c_528_n 0.0134757f $X=2.815 $Y=0.515 $X2=0
+ $Y2=0
cc_204 N_A_21_270#_c_92_n N_VGND_c_528_n 0.0119984f $X=3.875 $Y=0.515 $X2=0
+ $Y2=0
cc_205 N_A_21_270#_c_113_p A_351_74# 0.00732587f $X=2.63 $Y=1.005 $X2=-0.19
+ $Y2=-0.245
cc_206 N_A_21_270#_c_113_p A_423_74# 0.0181941f $X=2.63 $Y=1.005 $X2=-0.19
+ $Y2=-0.245
cc_207 N_A3_M1006_g N_A2_M1001_g 0.042114f $X=1.68 $Y=0.74 $X2=0 $Y2=0
cc_208 N_A3_c_233_n N_A2_M1001_g 0.00626927f $X=1.59 $Y=1.425 $X2=0 $Y2=0
cc_209 N_A3_c_230_n N_A2_c_271_n 0.0121574f $X=1.575 $Y=1.795 $X2=0 $Y2=0
cc_210 N_A3_c_235_n N_A2_c_271_n 0.0180709f $X=1.575 $Y=1.885 $X2=0 $Y2=0
cc_211 N_A3_c_232_n N_A2_c_271_n 0.042114f $X=1.59 $Y=1.425 $X2=0 $Y2=0
cc_212 N_A3_c_233_n A2 0.0258501f $X=1.59 $Y=1.425 $X2=0 $Y2=0
cc_213 N_A3_c_235_n N_VPWR_c_407_n 0.00534351f $X=1.575 $Y=1.885 $X2=0 $Y2=0
cc_214 N_A3_c_235_n N_VPWR_c_408_n 0.00445602f $X=1.575 $Y=1.885 $X2=0 $Y2=0
cc_215 N_A3_c_235_n N_VPWR_c_404_n 0.00858388f $X=1.575 $Y=1.885 $X2=0 $Y2=0
cc_216 N_A3_c_235_n N_A_330_392#_c_488_n 0.00505325f $X=1.575 $Y=1.885 $X2=0
+ $Y2=0
cc_217 N_A3_c_235_n N_A_330_392#_c_484_n 0.00494057f $X=1.575 $Y=1.885 $X2=0
+ $Y2=0
cc_218 N_A3_M1006_g N_VGND_c_519_n 0.012001f $X=1.68 $Y=0.74 $X2=0 $Y2=0
cc_219 N_A3_M1006_g N_VGND_c_525_n 0.00383152f $X=1.68 $Y=0.74 $X2=0 $Y2=0
cc_220 N_A3_M1006_g N_VGND_c_528_n 0.0075694f $X=1.68 $Y=0.74 $X2=0 $Y2=0
cc_221 N_A2_M1001_g N_A1_M1012_g 0.0410548f $X=2.04 $Y=0.74 $X2=0 $Y2=0
cc_222 N_A2_c_271_n N_A1_c_301_n 0.0465434f $X=2.055 $Y=1.885 $X2=0 $Y2=0
cc_223 A2 N_A1_c_301_n 0.00114936f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_224 N_A2_c_271_n A1 0.00114936f $X=2.055 $Y=1.885 $X2=0 $Y2=0
cc_225 A2 A1 0.0209133f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_226 N_A2_c_271_n N_VPWR_c_408_n 0.00339044f $X=2.055 $Y=1.885 $X2=0 $Y2=0
cc_227 N_A2_c_271_n N_VPWR_c_404_n 0.0044506f $X=2.055 $Y=1.885 $X2=0 $Y2=0
cc_228 N_A2_c_271_n N_VPWR_c_413_n 0.00582408f $X=2.055 $Y=1.885 $X2=0 $Y2=0
cc_229 N_A2_c_271_n N_A_330_392#_c_484_n 3.83538e-19 $X=2.055 $Y=1.885 $X2=0
+ $Y2=0
cc_230 N_A2_c_271_n N_A_330_392#_c_491_n 0.0148466f $X=2.055 $Y=1.885 $X2=0
+ $Y2=0
cc_231 N_A2_M1001_g N_VGND_c_519_n 0.00256807f $X=2.04 $Y=0.74 $X2=0 $Y2=0
cc_232 N_A2_M1001_g N_VGND_c_525_n 0.00461464f $X=2.04 $Y=0.74 $X2=0 $Y2=0
cc_233 N_A2_M1001_g N_VGND_c_528_n 0.00909747f $X=2.04 $Y=0.74 $X2=0 $Y2=0
cc_234 N_A1_M1012_g N_B1_M1004_g 0.0237799f $X=2.58 $Y=0.74 $X2=0 $Y2=0
cc_235 N_A1_c_301_n N_B1_c_334_n 0.0125479f $X=2.745 $Y=1.885 $X2=0 $Y2=0
cc_236 N_A1_c_301_n N_B1_c_338_n 0.0191334f $X=2.745 $Y=1.885 $X2=0 $Y2=0
cc_237 N_A1_M1012_g B1 0.00436692f $X=2.58 $Y=0.74 $X2=0 $Y2=0
cc_238 N_A1_c_301_n B1 0.0022363f $X=2.745 $Y=1.885 $X2=0 $Y2=0
cc_239 A1 B1 0.0278455f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_240 N_A1_c_301_n N_B1_c_336_n 0.00875058f $X=2.745 $Y=1.885 $X2=0 $Y2=0
cc_241 N_A1_c_301_n N_VPWR_c_410_n 0.00339044f $X=2.745 $Y=1.885 $X2=0 $Y2=0
cc_242 N_A1_c_301_n N_VPWR_c_404_n 0.0044506f $X=2.745 $Y=1.885 $X2=0 $Y2=0
cc_243 N_A1_c_301_n N_VPWR_c_413_n 0.00582408f $X=2.745 $Y=1.885 $X2=0 $Y2=0
cc_244 N_A1_c_301_n N_A_330_392#_c_491_n 0.0148466f $X=2.745 $Y=1.885 $X2=0
+ $Y2=0
cc_245 N_A1_c_301_n N_A_330_392#_c_485_n 3.83538e-19 $X=2.745 $Y=1.885 $X2=0
+ $Y2=0
cc_246 N_A1_M1012_g N_VGND_c_520_n 6.23202e-19 $X=2.58 $Y=0.74 $X2=0 $Y2=0
cc_247 N_A1_M1012_g N_VGND_c_525_n 0.00434272f $X=2.58 $Y=0.74 $X2=0 $Y2=0
cc_248 N_A1_M1012_g N_VGND_c_528_n 0.00823328f $X=2.58 $Y=0.74 $X2=0 $Y2=0
cc_249 N_B1_c_338_n N_C1_c_375_n 0.0544714f $X=3.225 $Y=1.885 $X2=-0.19
+ $Y2=-0.245
cc_250 N_B1_M1004_g N_C1_M1008_g 0.0232223f $X=3.12 $Y=0.74 $X2=0 $Y2=0
cc_251 B1 N_C1_M1008_g 0.0133809f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_252 N_B1_c_336_n N_C1_M1008_g 0.0213711f $X=3.21 $Y=1.425 $X2=0 $Y2=0
cc_253 N_B1_c_334_n N_C1_c_372_n 0.015845f $X=3.225 $Y=1.795 $X2=0 $Y2=0
cc_254 B1 N_C1_c_372_n 0.0155352f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_255 B1 C1 0.0271915f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_256 N_B1_c_338_n N_VPWR_c_410_n 0.00445602f $X=3.225 $Y=1.885 $X2=0 $Y2=0
cc_257 N_B1_c_338_n N_VPWR_c_404_n 0.00858504f $X=3.225 $Y=1.885 $X2=0 $Y2=0
cc_258 N_B1_c_338_n N_A_330_392#_c_492_n 0.0049297f $X=3.225 $Y=1.885 $X2=0
+ $Y2=0
cc_259 N_B1_c_338_n N_A_330_392#_c_485_n 0.00774064f $X=3.225 $Y=1.885 $X2=0
+ $Y2=0
cc_260 N_B1_M1004_g N_VGND_c_520_n 0.00917877f $X=3.12 $Y=0.74 $X2=0 $Y2=0
cc_261 N_B1_M1004_g N_VGND_c_525_n 0.00383152f $X=3.12 $Y=0.74 $X2=0 $Y2=0
cc_262 N_B1_M1004_g N_VGND_c_528_n 0.00758569f $X=3.12 $Y=0.74 $X2=0 $Y2=0
cc_263 N_C1_c_375_n N_VPWR_c_410_n 0.00445602f $X=3.645 $Y=1.885 $X2=0 $Y2=0
cc_264 N_C1_c_375_n N_VPWR_c_404_n 0.00862094f $X=3.645 $Y=1.885 $X2=0 $Y2=0
cc_265 N_C1_c_375_n N_A_330_392#_c_492_n 8.04855e-19 $X=3.645 $Y=1.885 $X2=0
+ $Y2=0
cc_266 N_C1_c_375_n N_A_330_392#_c_485_n 0.00118224f $X=3.645 $Y=1.885 $X2=0
+ $Y2=0
cc_267 N_C1_M1008_g N_VGND_c_520_n 0.0055626f $X=3.66 $Y=0.74 $X2=0 $Y2=0
cc_268 N_C1_M1008_g N_VGND_c_527_n 0.00434272f $X=3.66 $Y=0.74 $X2=0 $Y2=0
cc_269 N_C1_M1008_g N_VGND_c_528_n 0.00825192f $X=3.66 $Y=0.74 $X2=0 $Y2=0
cc_270 N_VPWR_c_407_n N_A_330_392#_c_484_n 0.0147692f $X=1.28 $Y=2.735 $X2=0
+ $Y2=0
cc_271 N_VPWR_c_408_n N_A_330_392#_c_484_n 0.0146094f $X=2.135 $Y=3.33 $X2=0
+ $Y2=0
cc_272 N_VPWR_c_404_n N_A_330_392#_c_484_n 0.0120527f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_273 N_VPWR_c_413_n N_A_330_392#_c_484_n 0.00163961f $X=2.4 $Y=2.825 $X2=0
+ $Y2=0
cc_274 N_VPWR_M1000_d N_A_330_392#_c_491_n 0.0116313f $X=2.13 $Y=1.96 $X2=0
+ $Y2=0
cc_275 N_VPWR_c_408_n N_A_330_392#_c_491_n 0.00206097f $X=2.135 $Y=3.33 $X2=0
+ $Y2=0
cc_276 N_VPWR_c_410_n N_A_330_392#_c_491_n 0.00206097f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_277 N_VPWR_c_404_n N_A_330_392#_c_491_n 0.00953739f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_278 N_VPWR_c_413_n N_A_330_392#_c_491_n 0.0347384f $X=2.4 $Y=2.825 $X2=0
+ $Y2=0
cc_279 N_VPWR_c_410_n N_A_330_392#_c_485_n 0.0146094f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_280 N_VPWR_c_404_n N_A_330_392#_c_485_n 0.0120527f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_281 N_VPWR_c_413_n N_A_330_392#_c_485_n 0.00163961f $X=2.4 $Y=2.825 $X2=0
+ $Y2=0
cc_282 N_X_c_462_n N_VGND_c_518_n 0.0289274f $X=0.895 $Y=0.495 $X2=0 $Y2=0
cc_283 N_X_c_462_n N_VGND_c_519_n 0.0158228f $X=0.895 $Y=0.495 $X2=0 $Y2=0
cc_284 N_X_c_462_n N_VGND_c_523_n 0.0143908f $X=0.895 $Y=0.495 $X2=0 $Y2=0
cc_285 N_X_c_462_n N_VGND_c_528_n 0.0118422f $X=0.895 $Y=0.495 $X2=0 $Y2=0
