* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__xnor2_2 A B VGND VNB VPB VPWR Y
M1000 a_133_368# A VPWR VPB phighvt w=1e+06u l=150000u
+  ad=3.45e+11p pd=2.69e+06u as=2.25905e+12p ps=1.319e+07u
M1001 Y a_133_368# a_340_107# VNB nshort w=740000u l=150000u
+  ad=4.008e+11p pd=2.67e+06u as=8.30525e+11p ps=8.22e+06u
M1002 Y B a_638_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=6.72e+11p pd=5.68e+06u as=9.566e+11p ps=6.32e+06u
M1003 VGND B a_340_107# VNB nshort w=740000u l=150000u
+  ad=1.024e+12p pd=7.92e+06u as=0p ps=0u
M1004 Y a_133_368# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_340_107# A VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND A a_340_107# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR B a_133_368# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_638_368# B Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR a_133_368# Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR A a_638_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_638_368# A VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_133_368# B a_151_74# VNB nshort w=740000u l=150000u
+  ad=2.06875e+11p pd=2.05e+06u as=1.776e+11p ps=1.96e+06u
M1013 a_151_74# A VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_340_107# a_133_368# Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_340_107# B VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
