* File: sky130_fd_sc_ls__o22ai_4.spice
* Created: Wed Sep  2 11:20:26 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__o22ai_4.pex.spice"
.subckt sky130_fd_sc_ls__o22ai_4  VNB VPB A1 A2 B1 B2 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B2	B2
* B1	B1
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1008 N_A_27_74#_M1008_d N_A1_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.1295 PD=2.05 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75000.2
+ SB=75007.4 A=0.111 P=1.78 MULT=1
MM1021 N_A_27_74#_M1021_d N_A1_M1021_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.7
+ SB=75006.9 A=0.111 P=1.78 MULT=1
MM1026 N_A_27_74#_M1021_d N_A1_M1026_g N_VGND_M1026_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.1
+ SB=75006.4 A=0.111 P=1.78 MULT=1
MM1002 N_A_27_74#_M1002_d N_A2_M1002_g N_VGND_M1026_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.6
+ SB=75005.9 A=0.111 P=1.78 MULT=1
MM1005 N_A_27_74#_M1002_d N_A2_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75002.1
+ SB=75005.5 A=0.111 P=1.78 MULT=1
MM1017 N_A_27_74#_M1017_d N_A2_M1017_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1184 AS=0.1295 PD=1.06 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.6
+ SB=75005 A=0.111 P=1.78 MULT=1
MM1027 N_A_27_74#_M1017_d N_A2_M1027_g N_VGND_M1027_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1184 AS=0.1406 PD=1.06 PS=1.12 NRD=6.48 NRS=4.86 M=1 R=4.93333 SA=75003
+ SB=75004.5 A=0.111 P=1.78 MULT=1
MM1029 N_A_27_74#_M1029_d N_A1_M1029_g N_VGND_M1027_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1073 AS=0.1406 PD=1.03 PS=1.12 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75003.6
+ SB=75004 A=0.111 P=1.78 MULT=1
MM1003 N_A_27_74#_M1029_d N_B1_M1003_g N_Y_M1003_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1073 AS=0.1258 PD=1.03 PS=1.08 NRD=1.62 NRS=9.72 M=1 R=4.93333 SA=75004
+ SB=75003.6 A=0.111 P=1.78 MULT=1
MM1010 N_A_27_74#_M1010_d N_B1_M1010_g N_Y_M1003_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1073 AS=0.1258 PD=1.03 PS=1.08 NRD=0.804 NRS=0 M=1 R=4.93333 SA=75004.5
+ SB=75003.1 A=0.111 P=1.78 MULT=1
MM1019 N_A_27_74#_M1010_d N_B1_M1019_g N_Y_M1019_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1073 AS=0.1036 PD=1.03 PS=1.02 NRD=0.804 NRS=0 M=1 R=4.93333 SA=75004.9
+ SB=75002.6 A=0.111 P=1.78 MULT=1
MM1009 N_A_27_74#_M1009_d N_B2_M1009_g N_Y_M1019_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75005.4
+ SB=75002.2 A=0.111 P=1.78 MULT=1
MM1014 N_A_27_74#_M1009_d N_B2_M1014_g N_Y_M1014_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75005.8
+ SB=75001.8 A=0.111 P=1.78 MULT=1
MM1018 N_A_27_74#_M1018_d N_B2_M1018_g N_Y_M1014_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1295 AS=0.1295 PD=1.09 PS=1.09 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75006.3
+ SB=75001.3 A=0.111 P=1.78 MULT=1
MM1022 N_A_27_74#_M1018_d N_B2_M1022_g N_Y_M1022_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1295 AS=0.1295 PD=1.09 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75006.8
+ SB=75000.8 A=0.111 P=1.78 MULT=1
MM1024 N_A_27_74#_M1024_d N_B1_M1024_g N_Y_M1022_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2991 AS=0.1295 PD=2.41 PS=1.09 NRD=13.776 NRS=0 M=1 R=4.93333 SA=75007.3
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1011 N_A_117_368#_M1011_d N_A1_M1011_g N_VPWR_M1011_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75007.3 A=0.168 P=2.54 MULT=1
MM1012 N_A_117_368#_M1011_d N_A1_M1012_g N_VPWR_M1012_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75006.9 A=0.168 P=2.54 MULT=1
MM1020 N_A_117_368#_M1020_d N_A1_M1020_g N_VPWR_M1012_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75001.2 SB=75006.4 A=0.168 P=2.54 MULT=1
MM1001 N_A_117_368#_M1020_d N_A2_M1001_g N_Y_M1001_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75001.6 SB=75005.9 A=0.168 P=2.54 MULT=1
MM1007 N_A_117_368#_M1007_d N_A2_M1007_g N_Y_M1001_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.1 SB=75005.4 A=0.168 P=2.54 MULT=1
MM1015 N_A_117_368#_M1007_d N_A2_M1015_g N_Y_M1015_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.6 SB=75005 A=0.168 P=2.54 MULT=1
MM1028 N_A_117_368#_M1028_d N_A2_M1028_g N_Y_M1015_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75003
+ SB=75004.5 A=0.168 P=2.54 MULT=1
MM1025 N_A_117_368#_M1028_d N_A1_M1025_g N_VPWR_M1025_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.224 PD=1.42 PS=1.52 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75003.5 SB=75004.1 A=0.168 P=2.54 MULT=1
MM1000 N_A_877_368#_M1000_d N_B1_M1000_g N_VPWR_M1025_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.224 PD=1.42 PS=1.52 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75004 SB=75003.5 A=0.168 P=2.54 MULT=1
MM1004 N_A_877_368#_M1000_d N_B1_M1004_g N_VPWR_M1004_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75004.5 SB=75003.1 A=0.168 P=2.54 MULT=1
MM1006 N_A_877_368#_M1006_d N_B1_M1006_g N_VPWR_M1004_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.196 AS=0.168 PD=1.47 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75004.9 SB=75002.6 A=0.168 P=2.54 MULT=1
MM1013 N_Y_M1013_d N_B2_M1013_g N_A_877_368#_M1006_d VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75005.4 SB=75002.1 A=0.168 P=2.54 MULT=1
MM1016 N_Y_M1013_d N_B2_M1016_g N_A_877_368#_M1016_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75005.9 SB=75001.7 A=0.168 P=2.54 MULT=1
MM1023 N_Y_M1023_d N_B2_M1023_g N_A_877_368#_M1016_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.1736 AS=0.168 PD=1.43 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75006.3 SB=75001.2 A=0.168 P=2.54 MULT=1
MM1030 N_Y_M1023_d N_B2_M1030_g N_A_877_368#_M1030_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.1736 AS=0.1904 PD=1.43 PS=1.46 NRD=3.5066 NRS=8.7862 M=1 R=7.46667
+ SA=75006.8 SB=75000.8 A=0.168 P=2.54 MULT=1
MM1031 N_A_877_368#_M1030_s N_B1_M1031_g N_VPWR_M1031_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.1904 AS=0.3864 PD=1.46 PS=2.93 NRD=1.7533 NRS=10.5395 M=1
+ R=7.46667 SA=75007.3 SB=75000.3 A=0.168 P=2.54 MULT=1
DX32_noxref VNB VPB NWDIODE A=15.8844 P=20.8
*
.include "sky130_fd_sc_ls__o22ai_4.pxi.spice"
*
.ends
*
*
