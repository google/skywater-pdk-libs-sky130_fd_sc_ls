* File: sky130_fd_sc_ls__nand2_8.spice
* Created: Wed Sep  2 11:11:36 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__nand2_8.pex.spice"
.subckt sky130_fd_sc_ls__nand2_8  VNB VPB B A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* B	B
* VPB	VPB
* VNB	VNB
MM1000 N_VGND_M1000_d N_B_M1000_g N_A_27_74#_M1000_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.2035 PD=1.02 PS=2.03 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75007.4 A=0.111 P=1.78 MULT=1
MM1010 N_VGND_M1000_d N_B_M1010_g N_A_27_74#_M1010_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75006.9 A=0.111 P=1.78 MULT=1
MM1011 N_VGND_M1011_d N_B_M1011_g N_A_27_74#_M1010_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75006.5 A=0.111 P=1.78 MULT=1
MM1012 N_VGND_M1011_d N_B_M1012_g N_A_27_74#_M1012_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75006.1 A=0.111 P=1.78 MULT=1
MM1015 N_VGND_M1015_d N_B_M1015_g N_A_27_74#_M1012_s VNB NSHORT L=0.15 W=0.74
+ AD=0.222 AS=0.1036 PD=1.34 PS=1.02 NRD=25.944 NRS=0 M=1 R=4.93333 SA=75001.9
+ SB=75005.6 A=0.111 P=1.78 MULT=1
MM1016 N_VGND_M1015_d N_B_M1016_g N_A_27_74#_M1016_s VNB NSHORT L=0.15 W=0.74
+ AD=0.222 AS=0.1184 PD=1.34 PS=1.06 NRD=25.944 NRS=3.24 M=1 R=4.93333
+ SA=75002.7 SB=75004.9 A=0.111 P=1.78 MULT=1
MM1021 N_VGND_M1021_d N_B_M1021_g N_A_27_74#_M1016_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1184 PD=1.02 PS=1.06 NRD=0 NRS=3.24 M=1 R=4.93333 SA=75003.1
+ SB=75004.4 A=0.111 P=1.78 MULT=1
MM1022 N_VGND_M1021_d N_B_M1022_g N_A_27_74#_M1022_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75003.6
+ SB=75004 A=0.111 P=1.78 MULT=1
MM1001 N_A_27_74#_M1022_s N_A_M1001_g N_Y_M1001_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75004
+ SB=75003.6 A=0.111 P=1.78 MULT=1
MM1002 N_A_27_74#_M1002_d N_A_M1002_g N_Y_M1001_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75004.4
+ SB=75003.1 A=0.111 P=1.78 MULT=1
MM1005 N_A_27_74#_M1002_d N_A_M1005_g N_Y_M1005_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75004.9
+ SB=75002.7 A=0.111 P=1.78 MULT=1
MM1008 N_A_27_74#_M1008_d N_A_M1008_g N_Y_M1005_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75005.3
+ SB=75002.3 A=0.111 P=1.78 MULT=1
MM1013 N_A_27_74#_M1008_d N_A_M1013_g N_Y_M1013_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75005.7
+ SB=75001.8 A=0.111 P=1.78 MULT=1
MM1014 N_A_27_74#_M1014_d N_A_M1014_g N_Y_M1013_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2368 AS=0.1036 PD=1.38 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75006.1
+ SB=75001.4 A=0.111 P=1.78 MULT=1
MM1017 N_A_27_74#_M1014_d N_A_M1017_g N_Y_M1017_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2368 AS=0.1036 PD=1.38 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75006.9
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1020 N_A_27_74#_M1020_d N_A_M1020_g N_Y_M1017_s VNB NSHORT L=0.15 W=0.74
+ AD=0.19805 AS=0.1036 PD=2.07 PS=1.02 NRD=0.804 NRS=0 M=1 R=4.93333 SA=75007.4
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1003 N_VPWR_M1003_d N_B_M1003_g N_Y_M1003_s VPB PHIGHVT L=0.15 W=1.12
+ AD=1.4952 AS=0.196 PD=4.91 PS=1.47 NRD=2.6201 NRS=1.7533 M=1 R=7.46667
+ SA=75001.3 SB=75003 A=0.168 P=2.54 MULT=1
MM1004 N_VPWR_M1004_d N_B_M1004_g N_Y_M1003_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.8904 AS=0.196 PD=2.71 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75001.8 SB=75002.5 A=0.168 P=2.54 MULT=1
MM1018 N_VPWR_M1004_d N_B_M1018_g N_Y_M1018_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.8904 AS=0.168 PD=2.71 PS=1.42 NRD=2.6201 NRS=1.7533 M=1 R=7.46667
+ SA=75003.5 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1019 N_VPWR_M1019_d N_B_M1019_g N_Y_M1018_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3864 AS=0.168 PD=2.93 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75003.9 SB=75000.3 A=0.168 P=2.54 MULT=1
MM1006 N_Y_M1006_d N_A_M1006_g N_VPWR_M1006_s VPB PHIGHVT L=0.15 W=1.12 AD=0.196
+ AS=0.3864 PD=1.47 PS=2.93 NRD=1.7533 NRS=10.5395 M=1 R=7.46667 SA=75000.3
+ SB=75002 A=0.168 P=2.54 MULT=1
MM1007 N_Y_M1006_d N_A_M1007_g N_VPWR_M1007_s VPB PHIGHVT L=0.15 W=1.12 AD=0.196
+ AS=0.3808 PD=1.47 PS=1.8 NRD=10.5395 NRS=1.7533 M=1 R=7.46667 SA=75000.8
+ SB=75001.5 A=0.168 P=2.54 MULT=1
MM1009 N_Y_M1009_d N_A_M1009_g N_VPWR_M1007_s VPB PHIGHVT L=0.15 W=1.12 AD=0.168
+ AS=0.3808 PD=1.42 PS=1.8 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75001.6
+ SB=75000.7 A=0.168 P=2.54 MULT=1
MM1023 N_Y_M1009_d N_A_M1023_g N_VPWR_M1023_s VPB PHIGHVT L=0.15 W=1.12 AD=0.168
+ AS=0.3248 PD=1.42 PS=2.82 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75002
+ SB=75000.2 A=0.168 P=2.54 MULT=1
DX24_noxref VNB VPB NWDIODE A=15.8844 P=20.8
*
.include "sky130_fd_sc_ls__nand2_8.pxi.spice"
*
.ends
*
*
