# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_ls__sdfxtp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_ls__sdfxtp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.04000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.455000 1.655000 1.785000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.528300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.600000 0.370000 10.935000 2.980000 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.405000 1.470000 2.740000 2.140000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 0.955000 2.250000 1.285000 ;
        RECT 1.085000 0.810000 1.315000 0.900000 ;
        RECT 1.085000 0.900000 2.250000 0.955000 ;
    END
  END SCE
  PIN VNB
    PORT
      LAYER pwell ;
        RECT 0.000000 0.000000 11.040000 0.245000 ;
    END
  END VNB
  PIN VPB
    PORT
      LAYER nwell ;
        RECT -0.190000 1.660000 11.230000 3.520000 ;
    END
  END VPB
  PIN CLK
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.250000 1.180000 3.685000 1.550000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 11.040000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 11.040000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.040000 0.085000 ;
      RECT  0.000000  3.245000 11.040000 3.415000 ;
      RECT  0.085000  0.350000  0.405000 0.785000 ;
      RECT  0.085000  0.785000  0.255000 1.525000 ;
      RECT  0.085000  1.525000  0.825000 1.955000 ;
      RECT  0.085000  1.955000  2.195000 2.125000 ;
      RECT  0.085000  2.125000  0.555000 2.980000 ;
      RECT  0.585000  0.085000  0.915000 0.785000 ;
      RECT  0.725000  2.300000  1.055000 3.245000 ;
      RECT  1.485000  0.400000  2.590000 0.730000 ;
      RECT  1.595000  2.310000  4.395000 2.390000 ;
      RECT  1.595000  2.390000  4.705000 2.480000 ;
      RECT  1.595000  2.480000  1.925000 2.980000 ;
      RECT  1.865000  1.470000  2.195000 1.955000 ;
      RECT  1.865000  2.125000  2.195000 2.140000 ;
      RECT  2.420000  0.730000  2.590000 1.130000 ;
      RECT  2.420000  1.130000  3.080000 1.300000 ;
      RECT  2.670000  2.650000  3.175000 3.245000 ;
      RECT  2.775000  0.085000  2.945000 0.790000 ;
      RECT  2.910000  1.300000  3.080000 2.310000 ;
      RECT  3.125000  0.350000  3.455000 0.790000 ;
      RECT  3.125000  0.790000  4.025000 0.960000 ;
      RECT  3.295000  1.820000  4.055000 2.140000 ;
      RECT  3.345000  2.480000  4.705000 2.560000 ;
      RECT  3.685000  0.085000  4.015000 0.620000 ;
      RECT  3.855000  0.960000  4.025000 1.300000 ;
      RECT  3.855000  1.300000  4.055000 1.820000 ;
      RECT  3.855000  2.730000  4.365000 3.245000 ;
      RECT  4.195000  0.255000  5.905000 0.425000 ;
      RECT  4.195000  0.425000  4.445000 1.130000 ;
      RECT  4.225000  1.480000  4.785000 1.650000 ;
      RECT  4.225000  1.650000  4.395000 2.310000 ;
      RECT  4.535000  2.560000  4.705000 2.710000 ;
      RECT  4.535000  2.710000  5.375000 2.980000 ;
      RECT  4.565000  1.820000  4.815000 2.050000 ;
      RECT  4.565000  2.050000  5.225000 2.220000 ;
      RECT  4.615000  0.595000  4.885000 0.940000 ;
      RECT  4.615000  0.940000  4.785000 1.480000 ;
      RECT  4.955000  2.220000  5.225000 2.380000 ;
      RECT  5.055000  0.425000  5.225000 2.050000 ;
      RECT  5.395000  0.595000  5.565000 1.530000 ;
      RECT  5.395000  1.530000  6.975000 1.700000 ;
      RECT  5.395000  1.700000  5.565000 2.370000 ;
      RECT  5.395000  2.370000  5.875000 2.540000 ;
      RECT  5.545000  2.540000  5.875000 2.980000 ;
      RECT  5.735000  0.425000  5.905000 0.690000 ;
      RECT  5.735000  0.690000  6.975000 0.860000 ;
      RECT  5.735000  0.860000  5.985000 1.360000 ;
      RECT  5.735000  1.870000  6.215000 2.200000 ;
      RECT  6.045000  2.200000  6.215000 2.520000 ;
      RECT  6.045000  2.520000  7.715000 2.690000 ;
      RECT  6.195000  1.030000  7.315000 1.360000 ;
      RECT  6.385000  0.085000  6.635000 0.520000 ;
      RECT  6.480000  2.860000  6.810000 3.245000 ;
      RECT  6.645000  1.700000  6.975000 1.930000 ;
      RECT  6.805000  0.255000  7.815000 0.425000 ;
      RECT  6.805000  0.425000  6.975000 0.690000 ;
      RECT  7.015000  2.100000  7.375000 2.350000 ;
      RECT  7.145000  0.595000  7.475000 0.860000 ;
      RECT  7.145000  0.860000  7.315000 1.030000 ;
      RECT  7.145000  1.360000  7.315000 2.100000 ;
      RECT  7.485000  1.030000  7.815000 1.190000 ;
      RECT  7.485000  1.190000  8.240000 1.320000 ;
      RECT  7.485000  1.320000  8.555000 1.360000 ;
      RECT  7.545000  1.600000  7.900000 1.930000 ;
      RECT  7.545000  1.930000  7.715000 2.520000 ;
      RECT  7.645000  0.425000  7.815000 1.030000 ;
      RECT  7.885000  2.100000  8.135000 2.245000 ;
      RECT  7.885000  2.245000  8.895000 2.415000 ;
      RECT  7.885000  2.415000  8.135000 2.980000 ;
      RECT  7.985000  0.480000  8.315000 0.770000 ;
      RECT  7.985000  0.770000  8.580000 0.940000 ;
      RECT  8.070000  1.360000  8.555000 1.490000 ;
      RECT  8.305000  1.490000  8.555000 2.075000 ;
      RECT  8.410000  0.940000  8.580000 0.980000 ;
      RECT  8.410000  0.980000  8.895000 1.150000 ;
      RECT  8.725000  1.150000  8.895000 1.600000 ;
      RECT  8.725000  1.600000  9.595000 1.930000 ;
      RECT  8.725000  1.930000  8.895000 2.245000 ;
      RECT  8.805000  0.085000  9.480000 0.810000 ;
      RECT  8.845000  2.650000  9.420000 3.245000 ;
      RECT  9.065000  1.030000  9.980000 1.320000 ;
      RECT  9.065000  1.320000 10.245000 1.360000 ;
      RECT  9.590000  2.100000  9.935000 2.980000 ;
      RECT  9.650000  0.350000  9.980000 1.030000 ;
      RECT  9.765000  1.360000 10.245000 1.650000 ;
      RECT  9.765000  1.650000  9.935000 2.100000 ;
      RECT 10.150000  1.820000 10.400000 3.245000 ;
      RECT 10.175000  0.085000 10.425000 1.150000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
  END
END sky130_fd_sc_ls__sdfxtp_1
END LIBRARY
