* File: sky130_fd_sc_ls__einvp_4.pex.spice
* Created: Wed Sep  2 11:07:18 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__EINVP_4%A 3 5 7 10 12 14 15 17 20 22 23 25 26 28 31
+ 33 34 35 36 49
r93 50 51 1.95935 $w=3.69e-07 $l=1.5e-08 $layer=POLY_cond $X=1.505 $Y=1.557
+ $X2=1.52 $Y2=1.557
r94 48 50 31.3496 $w=3.69e-07 $l=2.4e-07 $layer=POLY_cond $X=1.265 $Y=1.557
+ $X2=1.505 $Y2=1.557
r95 48 49 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.265
+ $Y=1.515 $X2=1.265 $Y2=1.515
r96 46 48 33.9621 $w=3.69e-07 $l=2.6e-07 $layer=POLY_cond $X=1.005 $Y=1.557
+ $X2=1.265 $Y2=1.557
r97 45 46 1.30623 $w=3.69e-07 $l=1e-08 $layer=POLY_cond $X=0.995 $Y=1.557
+ $X2=1.005 $Y2=1.557
r98 43 45 53.5556 $w=3.69e-07 $l=4.1e-07 $layer=POLY_cond $X=0.585 $Y=1.557
+ $X2=0.995 $Y2=1.557
r99 43 44 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.585
+ $Y=1.515 $X2=0.585 $Y2=1.515
r100 41 43 9.79675 $w=3.69e-07 $l=7.5e-08 $layer=POLY_cond $X=0.51 $Y=1.557
+ $X2=0.585 $Y2=1.557
r101 40 41 1.95935 $w=3.69e-07 $l=1.5e-08 $layer=POLY_cond $X=0.495 $Y=1.557
+ $X2=0.51 $Y2=1.557
r102 36 49 1.74206 $w=4.28e-07 $l=6.5e-08 $layer=LI1_cond $X=1.2 $Y=1.565
+ $X2=1.265 $Y2=1.565
r103 35 36 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=1.2 $Y2=1.565
r104 35 44 3.61813 $w=4.28e-07 $l=1.35e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=0.585 $Y2=1.565
r105 34 44 9.24634 $w=4.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.24 $Y=1.565
+ $X2=0.585 $Y2=1.565
r106 29 33 18.8402 $w=1.65e-07 $l=8.7892e-08 $layer=POLY_cond $X=1.995 $Y=1.35
+ $X2=1.967 $Y2=1.425
r107 29 31 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.995 $Y=1.35
+ $X2=1.995 $Y2=0.74
r108 26 28 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.955 $Y=1.765
+ $X2=1.955 $Y2=2.4
r109 25 26 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.955 $Y=1.675
+ $X2=1.955 $Y2=1.765
r110 24 33 18.8402 $w=1.65e-07 $l=8.07775e-08 $layer=POLY_cond $X=1.955 $Y=1.5
+ $X2=1.967 $Y2=1.425
r111 24 25 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=1.955 $Y=1.5
+ $X2=1.955 $Y2=1.675
r112 23 51 27.2843 $w=3.69e-07 $l=1.653e-07 $layer=POLY_cond $X=1.595 $Y=1.425
+ $X2=1.52 $Y2=1.557
r113 22 33 6.66866 $w=1.5e-07 $l=1.02e-07 $layer=POLY_cond $X=1.865 $Y=1.425
+ $X2=1.967 $Y2=1.425
r114 22 23 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=1.865 $Y=1.425
+ $X2=1.595 $Y2=1.425
r115 18 51 23.9013 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.52 $Y=1.35
+ $X2=1.52 $Y2=1.557
r116 18 20 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.52 $Y=1.35
+ $X2=1.52 $Y2=0.74
r117 15 50 23.9013 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.505 $Y=1.765
+ $X2=1.505 $Y2=1.557
r118 15 17 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.505 $Y=1.765
+ $X2=1.505 $Y2=2.4
r119 12 46 23.9013 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.005 $Y=1.765
+ $X2=1.005 $Y2=1.557
r120 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.005 $Y=1.765
+ $X2=1.005 $Y2=2.4
r121 8 45 23.9013 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.995 $Y=1.35
+ $X2=0.995 $Y2=1.557
r122 8 10 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.995 $Y=1.35
+ $X2=0.995 $Y2=0.74
r123 5 41 23.9013 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.51 $Y=1.765
+ $X2=0.51 $Y2=1.557
r124 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.51 $Y=1.765
+ $X2=0.51 $Y2=2.4
r125 1 40 23.9013 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=1.557
r126 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__EINVP_4%A_473_323# 1 2 7 9 10 11 12 14 15 17 19 20
+ 22 24 25 27 28 29 33 36 39 43 47
c113 25 0 1.57571e-20 $X=4.395 $Y=1.69
c114 7 0 2.41426e-19 $X=2.455 $Y=1.765
r115 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.56
+ $Y=2.825 $X2=4.56 $Y2=2.825
r116 43 45 0.16442 $w=7.42e-07 $l=1e-08 $layer=LI1_cond $X=4.795 $Y=2.815
+ $X2=4.795 $Y2=2.825
r117 41 43 13.6469 $w=7.42e-07 $l=8.3e-07 $layer=LI1_cond $X=4.795 $Y=1.985
+ $X2=4.795 $Y2=2.815
r118 39 46 178.359 $w=3.3e-07 $l=1.02e-06 $layer=POLY_cond $X=4.56 $Y=1.805
+ $X2=4.56 $Y2=2.825
r119 38 41 2.95957 $w=7.42e-07 $l=3.1229e-07 $layer=LI1_cond $X=4.56 $Y=1.805
+ $X2=4.795 $Y2=1.985
r120 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.56
+ $Y=1.805 $X2=4.56 $Y2=1.805
r121 36 38 11.294 $w=7.42e-07 $l=2.24332e-07 $layer=LI1_cond $X=4.7 $Y=1.64
+ $X2=4.56 $Y2=1.805
r122 36 47 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=4.7 $Y=1.64 $X2=4.7
+ $Y2=1.13
r123 31 47 9.49412 $w=3.88e-07 $l=1.95e-07 $layer=LI1_cond $X=4.81 $Y=0.935
+ $X2=4.81 $Y2=1.13
r124 31 33 12.4109 $w=3.88e-07 $l=4.2e-07 $layer=LI1_cond $X=4.81 $Y=0.935
+ $X2=4.81 $Y2=0.515
r125 30 39 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=4.56 $Y=1.765
+ $X2=4.56 $Y2=1.805
r126 26 29 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.94 $Y=1.69
+ $X2=3.865 $Y2=1.69
r127 25 30 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=4.395 $Y=1.69
+ $X2=4.56 $Y2=1.765
r128 25 26 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=4.395 $Y=1.69
+ $X2=3.94 $Y2=1.69
r129 22 29 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.865 $Y=1.765
+ $X2=3.865 $Y2=1.69
r130 22 24 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.865 $Y=1.765
+ $X2=3.865 $Y2=2.4
r131 21 28 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.48 $Y=1.69
+ $X2=3.405 $Y2=1.69
r132 20 29 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.79 $Y=1.69
+ $X2=3.865 $Y2=1.69
r133 20 21 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=3.79 $Y=1.69
+ $X2=3.48 $Y2=1.69
r134 17 28 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.405 $Y=1.765
+ $X2=3.405 $Y2=1.69
r135 17 19 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.405 $Y=1.765
+ $X2=3.405 $Y2=2.4
r136 16 27 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.03 $Y=1.69
+ $X2=2.955 $Y2=1.69
r137 15 28 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.33 $Y=1.69
+ $X2=3.405 $Y2=1.69
r138 15 16 153.83 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=3.33 $Y=1.69 $X2=3.03
+ $Y2=1.69
r139 12 27 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.955 $Y=1.765
+ $X2=2.955 $Y2=1.69
r140 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.955 $Y=1.765
+ $X2=2.955 $Y2=2.4
r141 10 27 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.88 $Y=1.69
+ $X2=2.955 $Y2=1.69
r142 10 11 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=2.88 $Y=1.69
+ $X2=2.53 $Y2=1.69
r143 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.455 $Y=1.765
+ $X2=2.53 $Y2=1.69
r144 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.455 $Y=1.765
+ $X2=2.455 $Y2=2.4
r145 2 43 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=4.885
+ $Y=1.84 $X2=5.03 $Y2=2.815
r146 2 41 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=4.885
+ $Y=1.84 $X2=5.03 $Y2=1.985
r147 1 33 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=4.695
+ $Y=0.37 $X2=4.84 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__EINVP_4%TE 1 3 4 5 6 8 9 11 13 14 16 18 19 21 23 24
+ 26 27 28 29 32 35 38
c100 38 0 1.57571e-20 $X=5.485 $Y=1.465
c101 5 0 1.65243e-20 $X=2.57 $Y=1.3
c102 1 0 1.81908e-19 $X=2.495 $Y=1.225
r103 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.485
+ $Y=1.465 $X2=5.485 $Y2=1.465
r104 35 37 25.1383 $w=4.41e-07 $l=2.3e-07 $layer=POLY_cond $X=5.255 $Y=1.495
+ $X2=5.485 $Y2=1.495
r105 34 35 21.8594 $w=4.41e-07 $l=2e-07 $layer=POLY_cond $X=5.055 $Y=1.495
+ $X2=5.255 $Y2=1.495
r106 32 38 0.930283 $w=4.48e-07 $l=3.5e-08 $layer=LI1_cond $X=5.52 $Y=1.405
+ $X2=5.485 $Y2=1.405
r107 24 35 28.2648 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=5.255 $Y=1.765
+ $X2=5.255 $Y2=1.495
r108 24 26 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.255 $Y=1.765
+ $X2=5.255 $Y2=2.4
r109 21 34 28.2648 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=5.055 $Y=1.225
+ $X2=5.055 $Y2=1.495
r110 21 23 155.847 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=5.055 $Y=1.225
+ $X2=5.055 $Y2=0.74
r111 20 29 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.14 $Y=1.3
+ $X2=4.065 $Y2=1.3
r112 19 34 30.6324 $w=4.41e-07 $l=2.29456e-07 $layer=POLY_cond $X=4.98 $Y=1.3
+ $X2=5.055 $Y2=1.495
r113 19 20 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=4.98 $Y=1.3
+ $X2=4.14 $Y2=1.3
r114 16 29 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.065 $Y=1.225
+ $X2=4.065 $Y2=1.3
r115 16 18 155.847 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=4.065 $Y=1.225
+ $X2=4.065 $Y2=0.74
r116 15 28 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.57 $Y=1.3
+ $X2=3.495 $Y2=1.3
r117 14 29 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.99 $Y=1.3
+ $X2=4.065 $Y2=1.3
r118 14 15 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=3.99 $Y=1.3
+ $X2=3.57 $Y2=1.3
r119 11 28 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.495 $Y=1.225
+ $X2=3.495 $Y2=1.3
r120 11 13 155.847 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=3.495 $Y=1.225
+ $X2=3.495 $Y2=0.74
r121 10 27 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.14 $Y=1.3
+ $X2=3.065 $Y2=1.3
r122 9 28 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.42 $Y=1.3
+ $X2=3.495 $Y2=1.3
r123 9 10 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.42 $Y=1.3 $X2=3.14
+ $Y2=1.3
r124 6 27 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.065 $Y=1.225
+ $X2=3.065 $Y2=1.3
r125 6 8 155.847 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=3.065 $Y=1.225
+ $X2=3.065 $Y2=0.74
r126 4 27 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.99 $Y=1.3
+ $X2=3.065 $Y2=1.3
r127 4 5 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=2.99 $Y=1.3 $X2=2.57
+ $Y2=1.3
r128 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.495 $Y=1.225
+ $X2=2.57 $Y2=1.3
r129 1 3 155.847 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=2.495 $Y=1.225
+ $X2=2.495 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__EINVP_4%A_27_368# 1 2 3 4 5 18 22 23 26 28 33 36 37
+ 40 44 48 52 53
r91 48 50 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=4.05 $Y=1.985
+ $X2=4.05 $Y2=2.815
r92 46 48 8.0671 $w=2.48e-07 $l=1.75e-07 $layer=LI1_cond $X=4.05 $Y=1.81
+ $X2=4.05 $Y2=1.985
r93 45 53 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.265 $Y=1.725
+ $X2=3.14 $Y2=1.725
r94 44 46 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.925 $Y=1.725
+ $X2=4.05 $Y2=1.81
r95 44 45 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=3.925 $Y=1.725
+ $X2=3.265 $Y2=1.725
r96 40 42 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=3.14 $Y=1.985
+ $X2=3.14 $Y2=2.815
r97 38 53 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.14 $Y=1.81
+ $X2=3.14 $Y2=1.725
r98 38 40 8.0671 $w=2.48e-07 $l=1.75e-07 $layer=LI1_cond $X=3.14 $Y=1.81
+ $X2=3.14 $Y2=1.985
r99 36 53 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.015 $Y=1.725
+ $X2=3.14 $Y2=1.725
r100 36 37 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=3.015 $Y=1.725
+ $X2=2.395 $Y2=1.725
r101 33 35 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=2.23 $Y=1.985
+ $X2=2.23 $Y2=2.815
r102 31 35 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=2.23 $Y=2.905
+ $X2=2.23 $Y2=2.815
r103 30 37 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.23 $Y=1.81
+ $X2=2.395 $Y2=1.725
r104 30 33 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=2.23 $Y=1.81
+ $X2=2.23 $Y2=1.985
r105 29 52 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.365 $Y=2.99
+ $X2=1.24 $Y2=2.99
r106 28 31 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.065 $Y=2.99
+ $X2=2.23 $Y2=2.905
r107 28 29 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=2.065 $Y=2.99
+ $X2=1.365 $Y2=2.99
r108 24 52 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.24 $Y=2.905
+ $X2=1.24 $Y2=2.99
r109 24 26 20.744 $w=2.48e-07 $l=4.5e-07 $layer=LI1_cond $X=1.24 $Y=2.905
+ $X2=1.24 $Y2=2.455
r110 22 52 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.115 $Y=2.99
+ $X2=1.24 $Y2=2.99
r111 22 23 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.115 $Y=2.99
+ $X2=0.445 $Y2=2.99
r112 18 21 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=0.28 $Y=2.035
+ $X2=0.28 $Y2=2.815
r113 16 23 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=2.905
+ $X2=0.445 $Y2=2.99
r114 16 21 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.28 $Y=2.905
+ $X2=0.28 $Y2=2.815
r115 5 50 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=3.94
+ $Y=1.84 $X2=4.09 $Y2=2.815
r116 5 48 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=3.94
+ $Y=1.84 $X2=4.09 $Y2=1.985
r117 4 42 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=3.03
+ $Y=1.84 $X2=3.18 $Y2=2.815
r118 4 40 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=3.03
+ $Y=1.84 $X2=3.18 $Y2=1.985
r119 3 35 400 $w=1.7e-07 $l=1.07034e-06 $layer=licon1_PDIFF $count=1 $X=2.03
+ $Y=1.84 $X2=2.23 $Y2=2.815
r120 3 33 400 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=1 $X=2.03
+ $Y=1.84 $X2=2.23 $Y2=1.985
r121 2 26 300 $w=1.7e-07 $l=7.07972e-07 $layer=licon1_PDIFF $count=2 $X=1.08
+ $Y=1.84 $X2=1.28 $Y2=2.455
r122 1 21 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r123 1 18 400 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.035
.ends

.subckt PM_SKY130_FD_SC_LS__EINVP_4%Z 1 2 3 4 15 19 20 21 25 28 30 33 34 35
c61 35 0 1.63851e-19 $X=1.68 $Y=2.405
c62 34 0 7.17626e-20 $X=1.78 $Y=1.095
c63 28 0 9.40992e-20 $X=1.755 $Y=1.95
c64 25 0 1.10145e-19 $X=1.78 $Y=0.825
r65 31 35 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=1.73 $Y=2.12
+ $X2=1.73 $Y2=2.405
r66 31 33 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.73 $Y=2.12
+ $X2=1.73 $Y2=2.035
r67 28 33 3.10218 $w=3.05e-07 $l=9.66954e-08 $layer=LI1_cond $X=1.755 $Y=1.95
+ $X2=1.73 $Y2=2.035
r68 27 34 3.10218 $w=3.05e-07 $l=9.66954e-08 $layer=LI1_cond $X=1.755 $Y=1.18
+ $X2=1.78 $Y2=1.095
r69 27 28 31.6922 $w=2.78e-07 $l=7.7e-07 $layer=LI1_cond $X=1.755 $Y=1.18
+ $X2=1.755 $Y2=1.95
r70 23 34 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.78 $Y=1.01
+ $X2=1.78 $Y2=1.095
r71 23 25 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=1.78 $Y=1.01
+ $X2=1.78 $Y2=0.825
r72 22 30 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=2.035
+ $X2=0.78 $Y2=2.035
r73 21 33 3.51065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.565 $Y=2.035
+ $X2=1.73 $Y2=2.035
r74 21 22 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=1.565 $Y=2.035
+ $X2=0.945 $Y2=2.035
r75 19 34 3.51065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.615 $Y=1.095
+ $X2=1.78 $Y2=1.095
r76 19 20 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.615 $Y=1.095
+ $X2=0.945 $Y2=1.095
r77 13 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.78 $Y=1.01
+ $X2=0.945 $Y2=1.095
r78 13 15 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=0.78 $Y=1.01
+ $X2=0.78 $Y2=0.825
r79 4 33 300 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=2 $X=1.58
+ $Y=1.84 $X2=1.73 $Y2=2.035
r80 3 30 300 $w=1.7e-07 $l=2.75772e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.84 $X2=0.78 $Y2=2.035
r81 2 25 182 $w=1.7e-07 $l=5.3963e-07 $layer=licon1_NDIFF $count=1 $X=1.595
+ $Y=0.37 $X2=1.78 $Y2=0.825
r82 1 15 182 $w=1.7e-07 $l=5.50068e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.78 $Y2=0.825
.ends

.subckt PM_SKY130_FD_SC_LS__EINVP_4%VPWR 1 2 3 12 18 22 24 28 30 35 40 49 52 56
r62 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r63 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r64 49 50 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r65 47 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r66 46 47 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r67 44 47 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r68 44 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r69 43 46 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.08 $Y=3.33 $X2=5.04
+ $Y2=3.33
r70 43 44 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r71 41 52 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.725 $Y=3.33
+ $X2=3.595 $Y2=3.33
r72 41 43 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=3.725 $Y=3.33
+ $X2=4.08 $Y2=3.33
r73 40 55 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=5.395 $Y=3.33
+ $X2=5.577 $Y2=3.33
r74 40 46 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=5.395 $Y=3.33
+ $X2=5.04 $Y2=3.33
r75 39 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r76 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r77 36 49 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.815 $Y=3.33
+ $X2=2.69 $Y2=3.33
r78 36 38 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.815 $Y=3.33
+ $X2=3.12 $Y2=3.33
r79 35 52 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.465 $Y=3.33
+ $X2=3.595 $Y2=3.33
r80 35 38 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=3.465 $Y=3.33
+ $X2=3.12 $Y2=3.33
r81 33 50 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=2.64 $Y2=3.33
r82 32 33 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r83 30 49 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.565 $Y=3.33
+ $X2=2.69 $Y2=3.33
r84 30 32 151.684 $w=1.68e-07 $l=2.325e-06 $layer=LI1_cond $X=2.565 $Y=3.33
+ $X2=0.24 $Y2=3.33
r85 28 39 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=3.12 $Y2=3.33
r86 28 50 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=2.64 $Y2=3.33
r87 24 27 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=5.52 $Y=1.985
+ $X2=5.52 $Y2=2.815
r88 22 55 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=5.52 $Y=3.245
+ $X2=5.577 $Y2=3.33
r89 22 27 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=5.52 $Y=3.245
+ $X2=5.52 $Y2=2.815
r90 18 21 30.1408 $w=2.58e-07 $l=6.8e-07 $layer=LI1_cond $X=3.595 $Y=2.145
+ $X2=3.595 $Y2=2.825
r91 16 52 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.595 $Y=3.245
+ $X2=3.595 $Y2=3.33
r92 16 21 18.6164 $w=2.58e-07 $l=4.2e-07 $layer=LI1_cond $X=3.595 $Y=3.245
+ $X2=3.595 $Y2=2.825
r93 12 15 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=2.69 $Y=2.145
+ $X2=2.69 $Y2=2.825
r94 10 49 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.69 $Y=3.245
+ $X2=2.69 $Y2=3.33
r95 10 15 19.361 $w=2.48e-07 $l=4.2e-07 $layer=LI1_cond $X=2.69 $Y=3.245
+ $X2=2.69 $Y2=2.825
r96 3 27 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=5.33
+ $Y=1.84 $X2=5.48 $Y2=2.815
r97 3 24 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=5.33
+ $Y=1.84 $X2=5.48 $Y2=1.985
r98 2 21 400 $w=1.7e-07 $l=1.05967e-06 $layer=licon1_PDIFF $count=1 $X=3.48
+ $Y=1.84 $X2=3.635 $Y2=2.825
r99 2 18 400 $w=1.7e-07 $l=3.74566e-07 $layer=licon1_PDIFF $count=1 $X=3.48
+ $Y=1.84 $X2=3.635 $Y2=2.145
r100 1 15 400 $w=1.7e-07 $l=1.08038e-06 $layer=licon1_PDIFF $count=1 $X=2.53
+ $Y=1.84 $X2=2.73 $Y2=2.825
r101 1 12 400 $w=1.7e-07 $l=3.9246e-07 $layer=licon1_PDIFF $count=1 $X=2.53
+ $Y=1.84 $X2=2.73 $Y2=2.145
.ends

.subckt PM_SKY130_FD_SC_LS__EINVP_4%A_27_74# 1 2 3 4 5 18 20 21 24 26 31 32 33
+ 36 38 42 44 45
r96 40 42 27.4142 $w=3.28e-07 $l=7.85e-07 $layer=LI1_cond $X=4.28 $Y=1.3
+ $X2=4.28 $Y2=0.515
r97 39 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.445 $Y=1.385
+ $X2=3.28 $Y2=1.385
r98 38 40 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.115 $Y=1.385
+ $X2=4.28 $Y2=1.3
r99 38 39 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.115 $Y=1.385
+ $X2=3.445 $Y2=1.385
r100 34 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.28 $Y=1.3 $X2=3.28
+ $Y2=1.385
r101 34 36 27.4142 $w=3.28e-07 $l=7.85e-07 $layer=LI1_cond $X=3.28 $Y=1.3
+ $X2=3.28 $Y2=0.515
r102 32 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.115 $Y=1.385
+ $X2=3.28 $Y2=1.385
r103 32 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.115 $Y=1.385
+ $X2=2.445 $Y2=1.385
r104 29 33 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.28 $Y=1.3
+ $X2=2.445 $Y2=1.385
r105 29 31 27.4142 $w=3.28e-07 $l=7.85e-07 $layer=LI1_cond $X=2.28 $Y=1.3
+ $X2=2.28 $Y2=0.515
r106 28 31 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=2.28 $Y=0.425
+ $X2=2.28 $Y2=0.515
r107 27 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.445 $Y=0.34
+ $X2=1.28 $Y2=0.34
r108 26 28 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.115 $Y=0.34
+ $X2=2.28 $Y2=0.425
r109 26 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.115 $Y=0.34
+ $X2=1.445 $Y2=0.34
r110 22 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.28 $Y=0.425
+ $X2=1.28 $Y2=0.34
r111 22 24 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=1.28 $Y=0.425
+ $X2=1.28 $Y2=0.635
r112 20 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.115 $Y=0.34
+ $X2=1.28 $Y2=0.34
r113 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.115 $Y=0.34
+ $X2=0.445 $Y2=0.34
r114 16 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=0.425
+ $X2=0.445 $Y2=0.34
r115 16 18 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.28 $Y=0.425
+ $X2=0.28 $Y2=0.515
r116 5 42 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.14
+ $Y=0.37 $X2=4.28 $Y2=0.515
r117 4 36 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.14
+ $Y=0.37 $X2=3.28 $Y2=0.515
r118 3 31 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=2.07
+ $Y=0.37 $X2=2.28 $Y2=0.515
r119 2 24 182 $w=1.7e-07 $l=3.54789e-07 $layer=licon1_NDIFF $count=1 $X=1.07
+ $Y=0.37 $X2=1.28 $Y2=0.635
r120 1 18 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__EINVP_4%VGND 1 2 3 12 16 18 20 23 24 25 27 36 44 48
r60 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r61 44 45 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r62 42 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r63 41 42 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r64 39 42 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=5.04
+ $Y2=0
r65 38 41 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.08 $Y=0 $X2=5.04
+ $Y2=0
r66 38 39 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r67 36 47 4.49945 $w=1.7e-07 $l=2.92e-07 $layer=LI1_cond $X=5.175 $Y=0 $X2=5.467
+ $Y2=0
r68 36 41 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=5.175 $Y=0 $X2=5.04
+ $Y2=0
r69 35 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r70 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r71 32 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.945 $Y=0 $X2=2.78
+ $Y2=0
r72 32 34 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=2.945 $Y=0 $X2=3.6
+ $Y2=0
r73 30 45 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=0.24 $Y=0 $X2=2.64
+ $Y2=0
r74 29 30 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r75 27 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.615 $Y=0 $X2=2.78
+ $Y2=0
r76 27 29 154.947 $w=1.68e-07 $l=2.375e-06 $layer=LI1_cond $X=2.615 $Y=0
+ $X2=0.24 $Y2=0
r77 25 35 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.88 $Y=0 $X2=3.6
+ $Y2=0
r78 25 45 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=0 $X2=2.64
+ $Y2=0
r79 23 34 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=3.615 $Y=0 $X2=3.6
+ $Y2=0
r80 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.615 $Y=0 $X2=3.78
+ $Y2=0
r81 22 38 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=3.945 $Y=0 $X2=4.08
+ $Y2=0
r82 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.945 $Y=0 $X2=3.78
+ $Y2=0
r83 18 47 3.26672 $w=3.3e-07 $l=1.64085e-07 $layer=LI1_cond $X=5.34 $Y=0.085
+ $X2=5.467 $Y2=0
r84 18 20 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=5.34 $Y=0.085
+ $X2=5.34 $Y2=0.515
r85 14 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.78 $Y=0.085
+ $X2=3.78 $Y2=0
r86 14 16 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.78 $Y=0.085
+ $X2=3.78 $Y2=0.515
r87 10 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.78 $Y=0.085
+ $X2=2.78 $Y2=0
r88 10 12 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.78 $Y=0.085
+ $X2=2.78 $Y2=0.515
r89 3 20 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=5.13
+ $Y=0.37 $X2=5.34 $Y2=0.515
r90 2 16 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=3.57
+ $Y=0.37 $X2=3.78 $Y2=0.515
r91 1 12 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=2.57
+ $Y=0.37 $X2=2.78 $Y2=0.515
.ends

