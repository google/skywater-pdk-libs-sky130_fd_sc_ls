* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
X0 VPWR D1 a_82_48# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X1 a_82_48# A2 a_600_381# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_82_48# D1 a_321_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X3 a_82_48# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X4 VPWR B1 a_82_48# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X5 X a_82_48# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X6 X a_82_48# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X7 a_393_74# B1 a_471_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X8 a_471_74# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X9 VGND A1 a_471_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X10 a_321_74# C1 a_393_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X11 a_600_381# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends
