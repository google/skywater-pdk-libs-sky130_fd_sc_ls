* File: sky130_fd_sc_ls__sdfrtp_1.pex.spice
* Created: Fri Aug 28 14:03:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__SDFRTP_1%SCE 2 5 7 9 11 12 14 19 20 21 22 25 26 30
+ 31 32 40 44 46 55 57
c96 40 0 9.7872e-20 $X=0.96 $Y=1.67
c97 26 0 1.56864e-19 $X=2.51 $Y=1.425
c98 25 0 2.15287e-19 $X=2.51 $Y=1.425
r99 46 55 1.90404 $w=3.43e-07 $l=5.7e-08 $layer=LI1_cond $X=1.623 $Y=1.662
+ $X2=1.68 $Y2=1.662
r100 40 42 6.6128 $w=3.28e-07 $l=4.5e-08 $layer=POLY_cond $X=0.96 $Y=1.67
+ $X2=1.005 $Y2=1.67
r101 40 41 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.96
+ $Y=1.67 $X2=0.96 $Y2=1.67
r102 38 40 66.8628 $w=3.28e-07 $l=4.55e-07 $layer=POLY_cond $X=0.505 $Y=1.67
+ $X2=0.96 $Y2=1.67
r103 37 38 1.46951 $w=3.28e-07 $l=1e-08 $layer=POLY_cond $X=0.495 $Y=1.67
+ $X2=0.505 $Y2=1.67
r104 32 57 6.34154 $w=3.43e-07 $l=1.01e-07 $layer=LI1_cond $X=1.694 $Y=1.662
+ $X2=1.795 $Y2=1.662
r105 32 55 0.467658 $w=3.43e-07 $l=1.4e-08 $layer=LI1_cond $X=1.694 $Y=1.662
+ $X2=1.68 $Y2=1.662
r106 32 46 0.467658 $w=3.43e-07 $l=1.4e-08 $layer=LI1_cond $X=1.609 $Y=1.662
+ $X2=1.623 $Y2=1.662
r107 31 32 13.6623 $w=3.43e-07 $l=4.09e-07 $layer=LI1_cond $X=1.2 $Y=1.662
+ $X2=1.609 $Y2=1.662
r108 31 41 8.01699 $w=3.43e-07 $l=2.4e-07 $layer=LI1_cond $X=1.2 $Y=1.662
+ $X2=0.96 $Y2=1.662
r109 30 41 8.01699 $w=3.43e-07 $l=2.4e-07 $layer=LI1_cond $X=0.72 $Y=1.662
+ $X2=0.96 $Y2=1.662
r110 26 44 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.51 $Y=1.425
+ $X2=2.51 $Y2=1.26
r111 25 28 4.54912 $w=3.78e-07 $l=1.5e-07 $layer=LI1_cond $X=2.535 $Y=1.425
+ $X2=2.535 $Y2=1.575
r112 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.51
+ $Y=1.425 $X2=2.51 $Y2=1.425
r113 22 28 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.345 $Y=1.575
+ $X2=2.535 $Y2=1.575
r114 22 57 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=2.345 $Y=1.575
+ $X2=1.795 $Y2=1.575
r115 21 44 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=2.6 $Y=1.05 $X2=2.6
+ $Y2=1.26
r116 20 21 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=2.625 $Y=0.9
+ $X2=2.625 $Y2=1.05
r117 19 20 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.65 $Y=0.615
+ $X2=2.65 $Y2=0.9
r118 12 14 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.005 $Y=2.245
+ $X2=1.005 $Y2=2.64
r119 11 12 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.005 $Y=2.155
+ $X2=1.005 $Y2=2.245
r120 10 42 16.7902 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.005 $Y=1.835
+ $X2=1.005 $Y2=1.67
r121 10 11 124.387 $w=1.8e-07 $l=3.2e-07 $layer=POLY_cond $X=1.005 $Y=1.835
+ $X2=1.005 $Y2=2.155
r122 7 9 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.505 $Y=2.245
+ $X2=0.505 $Y2=2.64
r123 3 37 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.505
+ $X2=0.495 $Y2=1.67
r124 3 5 438.415 $w=1.5e-07 $l=8.55e-07 $layer=POLY_cond $X=0.495 $Y=1.505
+ $X2=0.495 $Y2=0.65
r125 2 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.505 $Y=2.155
+ $X2=0.505 $Y2=2.245
r126 1 38 16.7902 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.835
+ $X2=0.505 $Y2=1.67
r127 1 2 124.387 $w=1.8e-07 $l=3.2e-07 $layer=POLY_cond $X=0.505 $Y=1.835
+ $X2=0.505 $Y2=2.155
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTP_1%A_27_88# 1 2 7 9 12 14 17 20 23 25 29 31 34
+ 35 37 38 42
c84 37 0 9.7872e-20 $X=1.21 $Y=1.1
c85 7 0 3.56444e-20 $X=1.485 $Y=0.935
r86 37 40 1.99058 $w=3.28e-07 $l=5.7e-08 $layer=LI1_cond $X=1.21 $Y=1.1 $X2=1.21
+ $Y2=1.157
r87 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.21
+ $Y=1.1 $X2=1.21 $Y2=1.1
r88 31 32 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.51
+ $Y=1.995 $X2=2.51 $Y2=1.995
r89 29 42 8.71323 $w=3.43e-07 $l=1.72e-07 $layer=LI1_cond $X=2.207 $Y=2.002
+ $X2=2.035 $Y2=2.002
r90 29 31 10.1215 $w=3.43e-07 $l=3.03e-07 $layer=LI1_cond $X=2.207 $Y=2.002
+ $X2=2.51 $Y2=2.002
r91 28 35 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.445 $Y=2.09
+ $X2=0.28 $Y2=2.09
r92 28 42 103.733 $w=1.68e-07 $l=1.59e-06 $layer=LI1_cond $X=0.445 $Y=2.09
+ $X2=2.035 $Y2=2.09
r93 26 34 1.25797 $w=2.15e-07 $l=1.25e-07 $layer=LI1_cond $X=0.365 $Y=1.157
+ $X2=0.24 $Y2=1.157
r94 25 40 3.26307 $w=2.15e-07 $l=1.65e-07 $layer=LI1_cond $X=1.045 $Y=1.157
+ $X2=1.21 $Y2=1.157
r95 25 26 36.4494 $w=2.13e-07 $l=6.8e-07 $layer=LI1_cond $X=1.045 $Y=1.157
+ $X2=0.365 $Y2=1.157
r96 21 35 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.28 $Y=2.175
+ $X2=0.28 $Y2=2.09
r97 21 23 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=0.28 $Y=2.175
+ $X2=0.28 $Y2=2.465
r98 20 35 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=0.2 $Y=2.005
+ $X2=0.28 $Y2=2.09
r99 19 34 5.26796 $w=2.1e-07 $l=1.26428e-07 $layer=LI1_cond $X=0.2 $Y=1.265
+ $X2=0.24 $Y2=1.157
r100 19 20 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=0.2 $Y=1.265
+ $X2=0.2 $Y2=2.005
r101 15 34 5.26796 $w=2.1e-07 $l=1.07e-07 $layer=LI1_cond $X=0.24 $Y=1.05
+ $X2=0.24 $Y2=1.157
r102 15 17 18.4391 $w=2.48e-07 $l=4e-07 $layer=LI1_cond $X=0.24 $Y=1.05 $X2=0.24
+ $Y2=0.65
r103 14 32 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=2.525 $Y=1.995
+ $X2=2.51 $Y2=1.995
r104 10 14 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=2.6 $Y=2.16
+ $X2=2.525 $Y2=1.995
r105 10 12 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.6 $Y=2.16 $X2=2.6
+ $Y2=2.64
r106 7 38 50.0189 $w=2.65e-07 $l=3.47851e-07 $layer=POLY_cond $X=1.485 $Y=0.935
+ $X2=1.21 $Y2=1.1
r107 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.485 $Y=0.935
+ $X2=1.485 $Y2=0.615
r108 2 23 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.32 $X2=0.28 $Y2=2.465
r109 1 17 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.44 $X2=0.28 $Y2=0.65
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTP_1%D 1 3 5 7 10 11 15 17 20 21 22
c57 15 0 6.10037e-20 $X=1.845 $Y=1.515
c58 5 0 1.54283e-19 $X=1.69 $Y=2.075
r59 20 23 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.935 $Y=1.1
+ $X2=1.935 $Y2=1.265
r60 20 22 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.935 $Y=1.1
+ $X2=1.935 $Y2=0.935
r61 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.935
+ $Y=1.1 $X2=1.935 $Y2=1.1
r62 17 21 6.7033 $w=4.53e-07 $l=2.55e-07 $layer=LI1_cond $X=1.68 $Y=1.037
+ $X2=1.935 $Y2=1.037
r63 13 15 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=1.69 $Y=1.515
+ $X2=1.845 $Y2=1.515
r64 11 12 80.8418 $w=1.58e-07 $l=2.65e-07 $layer=POLY_cond $X=1.425 $Y=2.16
+ $X2=1.69 $Y2=2.16
r65 10 22 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.875 $Y=0.615
+ $X2=1.875 $Y2=0.935
r66 7 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.845 $Y=1.44
+ $X2=1.845 $Y2=1.515
r67 7 23 89.734 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=1.845 $Y=1.44
+ $X2=1.845 $Y2=1.265
r68 5 12 4.07462 $w=1.5e-07 $l=8.5e-08 $layer=POLY_cond $X=1.69 $Y=2.075
+ $X2=1.69 $Y2=2.16
r69 4 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.69 $Y=1.59 $X2=1.69
+ $Y2=1.515
r70 4 5 248.691 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=1.69 $Y=1.59 $X2=1.69
+ $Y2=2.075
r71 1 11 4.07462 $w=1.5e-07 $l=8.5e-08 $layer=POLY_cond $X=1.425 $Y=2.245
+ $X2=1.425 $Y2=2.16
r72 1 3 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.425 $Y=2.245
+ $X2=1.425 $Y2=2.64
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTP_1%SCD 3 6 10 11 12 13 17
c41 12 0 1.56864e-19 $X=3.12 $Y=1.665
c42 11 0 8.81023e-20 $X=3.05 $Y=2.245
c43 6 0 1.93733e-19 $X=3.04 $Y=0.615
r44 12 13 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.11 $Y=1.605
+ $X2=3.11 $Y2=2.035
r45 12 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.05
+ $Y=1.605 $X2=3.05 $Y2=1.605
r46 10 17 83.0591 $w=3.3e-07 $l=4.75e-07 $layer=POLY_cond $X=3.05 $Y=2.08
+ $X2=3.05 $Y2=1.605
r47 10 11 38.3209 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.05 $Y=2.08
+ $X2=3.05 $Y2=2.245
r48 9 17 38.0424 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.05 $Y=1.44
+ $X2=3.05 $Y2=1.605
r49 6 9 423.032 $w=1.5e-07 $l=8.25e-07 $layer=POLY_cond $X=3.04 $Y=0.615
+ $X2=3.04 $Y2=1.44
r50 3 11 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.035 $Y=2.64
+ $X2=3.035 $Y2=2.245
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTP_1%CLK 1 2 3 5 7 10 12 13 16 19 20
c67 20 0 3.52919e-20 $X=3.95 $Y=1.115
c68 13 0 1.4151e-19 $X=4.62 $Y=1.885
c69 3 0 4.1107e-20 $X=4.595 $Y=1.41
c70 1 0 2.74116e-20 $X=4.52 $Y=1.515
r71 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.95
+ $Y=1.115 $X2=3.95 $Y2=1.115
r72 16 20 5.05951 $w=4.08e-07 $l=1.8e-07 $layer=LI1_cond $X=3.99 $Y=1.295
+ $X2=3.99 $Y2=1.115
r73 11 19 51.5841 $w=3.3e-07 $l=2.95e-07 $layer=POLY_cond $X=3.95 $Y=1.41
+ $X2=3.95 $Y2=1.115
r74 10 13 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=4.645 $Y=2.46
+ $X2=4.645 $Y2=1.885
r75 7 13 37.4512 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=4.62 $Y=1.785 $X2=4.62
+ $Y2=1.885
r76 6 12 23.6879 $w=1.75e-07 $l=1.05e-07 $layer=POLY_cond $X=4.62 $Y=1.62
+ $X2=4.62 $Y2=1.515
r77 6 7 54.7102 $w=2e-07 $l=1.65e-07 $layer=POLY_cond $X=4.62 $Y=1.62 $X2=4.62
+ $Y2=1.785
r78 3 12 23.6879 $w=1.75e-07 $l=1.16833e-07 $layer=POLY_cond $X=4.595 $Y=1.41
+ $X2=4.62 $Y2=1.515
r79 3 5 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=4.595 $Y=1.41
+ $X2=4.595 $Y2=0.965
r80 2 11 28.6974 $w=2.1e-07 $l=2.11069e-07 $layer=POLY_cond $X=4.115 $Y=1.515
+ $X2=3.95 $Y2=1.41
r81 1 12 2.7459 $w=2.1e-07 $l=1e-07 $layer=POLY_cond $X=4.52 $Y=1.515 $X2=4.62
+ $Y2=1.515
r82 1 2 127.894 $w=2.1e-07 $l=4.05e-07 $layer=POLY_cond $X=4.52 $Y=1.515
+ $X2=4.115 $Y2=1.515
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTP_1%A_1034_392# 1 2 8 9 11 12 16 18 20 22 23 25
+ 26 33 35 36 37 38 40 44 45 46 48 49 50 52 54 55 57 61 69 70 72 77
c220 70 0 1.39473e-19 $X=9.33 $Y=1.105
c221 61 0 4.1107e-20 $X=5.422 $Y=1.285
c222 46 0 1.61901e-19 $X=7.22 $Y=0.665
c223 9 0 1.93993e-19 $X=6.135 $Y=2.21
r224 69 77 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.25 $Y=1.105
+ $X2=9.085 $Y2=1.105
r225 68 70 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=9.25 $Y=1.105 $X2=9.33
+ $Y2=1.105
r226 68 69 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.25
+ $Y=1.105 $X2=9.25 $Y2=1.105
r227 65 68 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=9.15 $Y=1.105
+ $X2=9.25 $Y2=1.105
r228 60 61 9.72653 $w=4.03e-07 $l=2.15e-07 $layer=LI1_cond $X=5.422 $Y=1.07
+ $X2=5.422 $Y2=1.285
r229 57 58 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.81
+ $Y=2.215 $X2=9.81 $Y2=2.215
r230 55 57 17.8516 $w=2.53e-07 $l=3.95e-07 $layer=LI1_cond $X=9.415 $Y=2.252
+ $X2=9.81 $Y2=2.252
r231 54 55 7.17723 $w=2.55e-07 $l=1.64085e-07 $layer=LI1_cond $X=9.33 $Y=2.125
+ $X2=9.415 $Y2=2.252
r232 53 70 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.33 $Y=1.27
+ $X2=9.33 $Y2=1.105
r233 53 54 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=9.33 $Y=1.27
+ $X2=9.33 $Y2=2.125
r234 52 65 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.15 $Y=0.94
+ $X2=9.15 $Y2=1.105
r235 51 52 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=9.15 $Y=0.425
+ $X2=9.15 $Y2=0.94
r236 49 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.065 $Y=0.34
+ $X2=9.15 $Y2=0.425
r237 49 50 62.9572 $w=1.68e-07 $l=9.65e-07 $layer=LI1_cond $X=9.065 $Y=0.34
+ $X2=8.1 $Y2=0.34
r238 47 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.015 $Y=0.425
+ $X2=8.1 $Y2=0.34
r239 47 48 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=8.015 $Y=0.425
+ $X2=8.015 $Y2=0.58
r240 45 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.93 $Y=0.665
+ $X2=8.015 $Y2=0.58
r241 45 46 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=7.93 $Y=0.665
+ $X2=7.22 $Y2=0.665
r242 44 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.135 $Y=0.58
+ $X2=7.22 $Y2=0.665
r243 43 44 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=7.135 $Y=0.425
+ $X2=7.135 $Y2=0.58
r244 41 75 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.085 $Y=1.71
+ $X2=6.085 $Y2=1.875
r245 41 72 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=6.085 $Y=1.71
+ $X2=6.085 $Y2=1.635
r246 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.085
+ $Y=1.71 $X2=6.085 $Y2=1.71
r247 38 40 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=5.63 $Y=1.71
+ $X2=6.085 $Y2=1.71
r248 36 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.05 $Y=0.34
+ $X2=7.135 $Y2=0.425
r249 36 37 93.2941 $w=1.68e-07 $l=1.43e-06 $layer=LI1_cond $X=7.05 $Y=0.34
+ $X2=5.62 $Y2=0.34
r250 35 38 10.1667 $w=1.78e-07 $l=1.65e-07 $layer=LI1_cond $X=5.54 $Y=1.545
+ $X2=5.54 $Y2=1.71
r251 35 61 16.0202 $w=1.78e-07 $l=2.6e-07 $layer=LI1_cond $X=5.54 $Y=1.545
+ $X2=5.54 $Y2=1.285
r252 33 60 8.25206 $w=4.03e-07 $l=2.9e-07 $layer=LI1_cond $X=5.417 $Y=0.78
+ $X2=5.417 $Y2=1.07
r253 30 37 8.41448 $w=1.7e-07 $l=2.41793e-07 $layer=LI1_cond $X=5.417 $Y=0.425
+ $X2=5.62 $Y2=0.34
r254 30 33 10.1017 $w=4.03e-07 $l=3.55e-07 $layer=LI1_cond $X=5.417 $Y=0.425
+ $X2=5.417 $Y2=0.78
r255 26 38 23.1061 $w=1.78e-07 $l=3.75e-07 $layer=LI1_cond $X=5.54 $Y=2.085
+ $X2=5.54 $Y2=1.71
r256 26 28 5.76222 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=5.45 $Y=2.085
+ $X2=5.32 $Y2=2.085
r257 23 58 52.063 $w=3.03e-07 $l=2.86356e-07 $layer=POLY_cond $X=9.89 $Y=2.465
+ $X2=9.812 $Y2=2.215
r258 23 25 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=9.89 $Y=2.465
+ $X2=9.89 $Y2=2.75
r259 22 77 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=8.725 $Y=1.16
+ $X2=9.085 $Y2=1.16
r260 18 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.65 $Y=1.085
+ $X2=8.725 $Y2=1.16
r261 18 20 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=8.65 $Y=1.085
+ $X2=8.65 $Y2=0.69
r262 14 16 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=6.525 $Y=1.545
+ $X2=6.525 $Y2=0.805
r263 13 72 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.25 $Y=1.635
+ $X2=6.085 $Y2=1.635
r264 12 14 27.2212 $w=1.8e-07 $l=1.21861e-07 $layer=POLY_cond $X=6.45 $Y=1.635
+ $X2=6.525 $Y2=1.545
r265 12 13 77.7419 $w=1.8e-07 $l=2e-07 $layer=POLY_cond $X=6.45 $Y=1.635
+ $X2=6.25 $Y2=1.635
r266 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.135 $Y=2.21
+ $X2=6.135 $Y2=2.495
r267 8 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.135 $Y=2.12 $X2=6.135
+ $Y2=2.21
r268 8 75 95.2339 $w=1.8e-07 $l=2.45e-07 $layer=POLY_cond $X=6.135 $Y=2.12
+ $X2=6.135 $Y2=1.875
r269 2 28 600 $w=1.7e-07 $l=2.33238e-07 $layer=licon1_PDIFF $count=1 $X=5.17
+ $Y=1.96 $X2=5.32 $Y2=2.13
r270 1 33 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=5.22
+ $Y=0.595 $X2=5.36 $Y2=0.78
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTP_1%A_1367_93# 1 2 9 12 13 15 18 19 21 22 25 27
+ 32 34
c112 18 0 4.99889e-20 $X=7.185 $Y=1.64
c113 9 0 1.55517e-19 $X=6.91 $Y=0.805
r114 35 37 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=6.91 $Y=1.64
+ $X2=7.06 $Y2=1.64
r115 27 29 29.2227 $w=2.78e-07 $l=7.1e-07 $layer=LI1_cond $X=8.865 $Y=1.88
+ $X2=8.865 $Y2=2.59
r116 25 34 7.52792 $w=2.78e-07 $l=1.4e-07 $layer=LI1_cond $X=8.865 $Y=1.855
+ $X2=8.865 $Y2=1.715
r117 25 27 1.02897 $w=2.78e-07 $l=2.5e-08 $layer=LI1_cond $X=8.865 $Y=1.855
+ $X2=8.865 $Y2=1.88
r118 23 32 12.3649 $w=3.7e-07 $l=4.83348e-07 $layer=LI1_cond $X=8.81 $Y=1.09
+ $X2=8.435 $Y2=0.842
r119 23 34 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=8.81 $Y=1.09
+ $X2=8.81 $Y2=1.715
r120 21 32 9.03936 $w=3.7e-07 $l=2.32637e-07 $layer=LI1_cond $X=8.27 $Y=1.005
+ $X2=8.435 $Y2=0.842
r121 21 22 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=8.27 $Y=1.005
+ $X2=7.325 $Y2=1.005
r122 19 37 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=7.185 $Y=1.64
+ $X2=7.06 $Y2=1.64
r123 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.185
+ $Y=1.64 $X2=7.185 $Y2=1.64
r124 16 22 7.32204 $w=1.7e-07 $l=1.75425e-07 $layer=LI1_cond $X=7.187 $Y=1.09
+ $X2=7.325 $Y2=1.005
r125 16 18 23.0489 $w=2.73e-07 $l=5.5e-07 $layer=LI1_cond $X=7.187 $Y=1.09
+ $X2=7.187 $Y2=1.64
r126 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.06 $Y=2.23
+ $X2=7.06 $Y2=2.515
r127 12 13 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=7.06 $Y=2.14 $X2=7.06
+ $Y2=2.23
r128 11 37 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.06 $Y=1.805
+ $X2=7.06 $Y2=1.64
r129 11 12 130.218 $w=1.8e-07 $l=3.35e-07 $layer=POLY_cond $X=7.06 $Y=1.805
+ $X2=7.06 $Y2=2.14
r130 7 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.91 $Y=1.475
+ $X2=6.91 $Y2=1.64
r131 7 9 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=6.91 $Y=1.475
+ $X2=6.91 $Y2=0.805
r132 2 29 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=8.77
+ $Y=1.735 $X2=8.92 $Y2=2.59
r133 2 27 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=8.77
+ $Y=1.735 $X2=8.92 $Y2=1.88
r134 1 32 182 $w=1.7e-07 $l=5.05173e-07 $layer=licon1_NDIFF $count=1 $X=8.295
+ $Y=0.37 $X2=8.435 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTP_1%RESET_B 4 7 8 9 10 11 15 16 17 19 20 22 25
+ 28 30 31 33 36 39 41 42 43 44 51 52 56 58 66 67
c230 56 0 1.4151e-19 $X=3.95 $Y=1.995
c231 43 0 1.37312e-19 $X=10.655 $Y=2.035
c232 42 0 2.74116e-20 $X=4.225 $Y=2.035
c233 39 0 6.31244e-20 $X=10.715 $Y=1.375
c234 36 0 9.37604e-20 $X=3.56 $Y=2.245
c235 25 0 5.21422e-20 $X=10.6 $Y=0.58
c236 15 0 1.88097e-19 $X=7.3 $Y=0.805
r237 65 67 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=10.805 $Y=1.985
+ $X2=10.885 $Y2=1.985
r238 65 66 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.805
+ $Y=1.985 $X2=10.805 $Y2=1.985
r239 62 65 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=10.715 $Y=1.985
+ $X2=10.805 $Y2=1.985
r240 58 60 42.6489 $w=3.56e-07 $l=3.15e-07 $layer=POLY_cond $X=7.685 $Y=2.022
+ $X2=8 $Y2=2.022
r241 57 58 2.0309 $w=3.56e-07 $l=1.5e-08 $layer=POLY_cond $X=7.67 $Y=2.022
+ $X2=7.685 $Y2=2.022
r242 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.95
+ $Y=1.995 $X2=3.95 $Y2=1.995
r243 52 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=2.035
+ $X2=10.8 $Y2=2.035
r244 51 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8 $Y=1.98
+ $X2=8 $Y2=1.98
r245 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=2.035
+ $X2=7.92 $Y2=2.035
r246 46 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=2.035
+ $X2=4.08 $Y2=2.035
r247 44 50 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.065 $Y=2.035
+ $X2=7.92 $Y2=2.035
r248 43 52 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=10.655 $Y=2.035
+ $X2=10.8 $Y2=2.035
r249 43 44 3.20544 $w=1.4e-07 $l=2.59e-06 $layer=MET1_cond $X=10.655 $Y=2.035
+ $X2=8.065 $Y2=2.035
r250 42 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.225 $Y=2.035
+ $X2=4.08 $Y2=2.035
r251 41 50 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.775 $Y=2.035
+ $X2=7.92 $Y2=2.035
r252 41 42 4.39356 $w=1.4e-07 $l=3.55e-06 $layer=MET1_cond $X=7.775 $Y=2.035
+ $X2=4.225 $Y2=2.035
r253 37 39 58.9681 $w=1.5e-07 $l=1.15e-07 $layer=POLY_cond $X=10.6 $Y=1.375
+ $X2=10.715 $Y2=1.375
r254 31 33 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=10.885 $Y=2.465
+ $X2=10.885 $Y2=2.75
r255 30 31 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=10.885 $Y=2.375
+ $X2=10.885 $Y2=2.465
r256 29 67 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=10.885 $Y=2.15
+ $X2=10.885 $Y2=1.985
r257 29 30 87.4597 $w=1.8e-07 $l=2.25e-07 $layer=POLY_cond $X=10.885 $Y=2.15
+ $X2=10.885 $Y2=2.375
r258 28 62 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.715 $Y=1.82
+ $X2=10.715 $Y2=1.985
r259 27 39 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.715 $Y=1.45
+ $X2=10.715 $Y2=1.375
r260 27 28 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=10.715 $Y=1.45
+ $X2=10.715 $Y2=1.82
r261 23 37 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.6 $Y=1.3
+ $X2=10.6 $Y2=1.375
r262 23 25 369.191 $w=1.5e-07 $l=7.2e-07 $layer=POLY_cond $X=10.6 $Y=1.3
+ $X2=10.6 $Y2=0.58
r263 20 58 23.0368 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=7.685 $Y=2.23
+ $X2=7.685 $Y2=2.022
r264 20 22 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.685 $Y=2.23
+ $X2=7.685 $Y2=2.515
r265 19 57 23.0368 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.67 $Y=1.815
+ $X2=7.67 $Y2=2.022
r266 18 19 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=7.67 $Y=1.265
+ $X2=7.67 $Y2=1.815
r267 16 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.595 $Y=1.19
+ $X2=7.67 $Y2=1.265
r268 16 17 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=7.595 $Y=1.19
+ $X2=7.375 $Y2=1.19
r269 13 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.3 $Y=1.115
+ $X2=7.375 $Y2=1.19
r270 13 15 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=7.3 $Y=1.115
+ $X2=7.3 $Y2=0.805
r271 12 15 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=7.3 $Y=0.255
+ $X2=7.3 $Y2=0.805
r272 11 36 67.3007 $w=2.7e-07 $l=2.5e-07 $layer=POLY_cond $X=3.56 $Y=1.995
+ $X2=3.56 $Y2=2.245
r273 11 35 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.56 $Y=1.995
+ $X2=3.56 $Y2=1.83
r274 10 55 2.92121 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=3.93 $Y=1.995
+ $X2=3.95 $Y2=1.995
r275 10 11 41.0924 $w=3.3e-07 $l=2.35e-07 $layer=POLY_cond $X=3.93 $Y=1.995
+ $X2=3.695 $Y2=1.995
r276 8 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.225 $Y=0.18
+ $X2=7.3 $Y2=0.255
r277 8 9 1871.6 $w=1.5e-07 $l=3.65e-06 $layer=POLY_cond $X=7.225 $Y=0.18
+ $X2=3.575 $Y2=0.18
r278 7 36 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.605 $Y=2.64
+ $X2=3.605 $Y2=2.245
r279 4 35 623.011 $w=1.5e-07 $l=1.215e-06 $layer=POLY_cond $X=3.5 $Y=0.615
+ $X2=3.5 $Y2=1.83
r280 1 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.5 $Y=0.255
+ $X2=3.575 $Y2=0.18
r281 1 4 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=3.5 $Y=0.255 $X2=3.5
+ $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTP_1%A_1234_119# 1 2 3 12 14 16 18 19 23 26 27
+ 30 31 33 34 37 41
c136 41 0 1.93993e-19 $X=6.795 $Y=2.522
c137 34 0 4.99889e-20 $X=8.15 $Y=1.41
c138 30 0 7.00504e-20 $X=7.58 $Y=2.32
c139 26 0 3.72382e-19 $X=6.795 $Y=2.32
c140 23 0 1.51838e-20 $X=6.71 $Y=0.945
r141 37 39 4.78707 $w=3.23e-07 $l=1.35e-07 $layer=LI1_cond $X=6.307 $Y=0.81
+ $X2=6.307 $Y2=0.945
r142 34 46 16.6207 $w=3.19e-07 $l=1.1e-07 $layer=POLY_cond $X=8.15 $Y=1.41
+ $X2=8.15 $Y2=1.52
r143 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.15
+ $Y=1.41 $X2=8.15 $Y2=1.41
r144 31 33 17.744 $w=3.13e-07 $l=4.85e-07 $layer=LI1_cond $X=7.665 $Y=1.417
+ $X2=8.15 $Y2=1.417
r145 30 44 12.781 $w=3.15e-07 $l=4.22918e-07 $layer=LI1_cond $X=7.58 $Y=2.32
+ $X2=7.91 $Y2=2.532
r146 29 31 7.64049 $w=3.15e-07 $l=1.95944e-07 $layer=LI1_cond $X=7.58 $Y=1.575
+ $X2=7.665 $Y2=1.417
r147 29 30 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=7.58 $Y=1.575
+ $X2=7.58 $Y2=2.32
r148 28 41 3.64284 $w=2.55e-07 $l=1.53734e-07 $layer=LI1_cond $X=6.88 $Y=2.405
+ $X2=6.795 $Y2=2.522
r149 27 30 5.86024 $w=3.15e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.495 $Y=2.405
+ $X2=7.58 $Y2=2.32
r150 27 28 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=7.495 $Y=2.405
+ $X2=6.88 $Y2=2.405
r151 26 41 2.83584 $w=1.7e-07 $l=2.02e-07 $layer=LI1_cond $X=6.795 $Y=2.32
+ $X2=6.795 $Y2=2.522
r152 25 26 84.1604 $w=1.68e-07 $l=1.29e-06 $layer=LI1_cond $X=6.795 $Y=1.03
+ $X2=6.795 $Y2=2.32
r153 24 39 4.53325 $w=1.7e-07 $l=1.63e-07 $layer=LI1_cond $X=6.47 $Y=0.945
+ $X2=6.307 $Y2=0.945
r154 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.71 $Y=0.945
+ $X2=6.795 $Y2=1.03
r155 23 24 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=6.71 $Y=0.945
+ $X2=6.47 $Y2=0.945
r156 19 41 3.64284 $w=2.55e-07 $l=1.0015e-07 $layer=LI1_cond $X=6.71 $Y=2.555
+ $X2=6.795 $Y2=2.522
r157 19 21 9.99914 $w=3.38e-07 $l=2.95e-07 $layer=LI1_cond $X=6.71 $Y=2.555
+ $X2=6.415 $Y2=2.555
r158 16 18 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=8.695 $Y=1.66
+ $X2=8.695 $Y2=2.235
r159 15 46 20.418 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.315 $Y=1.52
+ $X2=8.15 $Y2=1.52
r160 14 16 26.9307 $w=1.5e-07 $l=1.79444e-07 $layer=POLY_cond $X=8.605 $Y=1.52
+ $X2=8.695 $Y2=1.66
r161 14 15 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=8.605 $Y=1.52
+ $X2=8.315 $Y2=1.52
r162 10 34 38.5462 $w=3.19e-07 $l=1.96914e-07 $layer=POLY_cond $X=8.22 $Y=1.245
+ $X2=8.15 $Y2=1.41
r163 10 12 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=8.22 $Y=1.245
+ $X2=8.22 $Y2=0.69
r164 3 44 600 $w=1.7e-07 $l=2.90474e-07 $layer=licon1_PDIFF $count=1 $X=7.76
+ $Y=2.305 $X2=7.91 $Y2=2.53
r165 2 21 600 $w=1.7e-07 $l=3.5812e-07 $layer=licon1_PDIFF $count=1 $X=6.21
+ $Y=2.285 $X2=6.415 $Y2=2.555
r166 1 37 182 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=1 $X=6.17
+ $Y=0.595 $X2=6.31 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTP_1%A_835_98# 1 2 7 9 10 12 14 15 16 17 19 21
+ 22 23 24 26 27 29 30 34 35 36 38 41 43 46 49 50 51 53 57 61 64
c201 61 0 1.29052e-19 $X=4.927 $Y=1.852
c202 41 0 2.96321e-20 $X=9.785 $Y=0.58
c203 35 0 1.09841e-19 $X=9.625 $Y=1.585
c204 19 0 1.51838e-20 $X=6.095 $Y=1.115
c205 7 0 1.94423e-19 $X=5.095 $Y=1.875
r206 63 64 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.115
+ $Y=1.635 $X2=5.115 $Y2=1.635
r207 61 63 5.297 $w=4.33e-07 $l=2.96454e-07 $layer=LI1_cond $X=4.927 $Y=1.852
+ $X2=5.115 $Y2=1.635
r208 60 61 14.285 $w=4.33e-07 $l=5.07e-07 $layer=LI1_cond $X=4.42 $Y=1.852
+ $X2=4.927 $Y2=1.852
r209 55 57 5.9927 $w=2.48e-07 $l=1.3e-07 $layer=LI1_cond $X=4.32 $Y=0.625
+ $X2=4.45 $Y2=0.625
r210 53 61 4.32933 $w=2.35e-07 $l=3.97e-07 $layer=LI1_cond $X=4.927 $Y=1.455
+ $X2=4.927 $Y2=1.852
r211 52 53 17.8996 $w=2.33e-07 $l=3.65e-07 $layer=LI1_cond $X=4.927 $Y=1.09
+ $X2=4.927 $Y2=1.455
r212 50 52 7.04737 $w=1.7e-07 $l=1.53734e-07 $layer=LI1_cond $X=4.81 $Y=1.005
+ $X2=4.927 $Y2=1.09
r213 50 51 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.81 $Y=1.005
+ $X2=4.535 $Y2=1.005
r214 49 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.45 $Y=0.92
+ $X2=4.535 $Y2=1.005
r215 48 57 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.45 $Y=0.75
+ $X2=4.45 $Y2=0.625
r216 48 49 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.45 $Y=0.75
+ $X2=4.45 $Y2=0.92
r217 44 46 43.5851 $w=1.5e-07 $l=8.5e-08 $layer=POLY_cond $X=9.7 $Y=1.045
+ $X2=9.785 $Y2=1.045
r218 39 46 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.785 $Y=0.97
+ $X2=9.785 $Y2=1.045
r219 39 41 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=9.785 $Y=0.97
+ $X2=9.785 $Y2=0.58
r220 37 44 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.7 $Y=1.12 $X2=9.7
+ $Y2=1.045
r221 37 38 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=9.7 $Y=1.12 $X2=9.7
+ $Y2=1.51
r222 35 38 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.625 $Y=1.585
+ $X2=9.7 $Y2=1.51
r223 35 36 207.67 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=9.625 $Y=1.585
+ $X2=9.22 $Y2=1.585
r224 32 34 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=9.145 $Y=2.81
+ $X2=9.145 $Y2=2.235
r225 31 36 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.145 $Y=1.66
+ $X2=9.22 $Y2=1.585
r226 31 34 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=9.145 $Y=1.66
+ $X2=9.145 $Y2=2.235
r227 29 32 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=9.145 $Y=2.9
+ $X2=9.145 $Y2=2.81
r228 29 30 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=9.145 $Y=2.9
+ $X2=9.145 $Y2=3.075
r229 28 43 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=6.73 $Y=3.15 $X2=6.64
+ $Y2=3.15
r230 27 30 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=9.055 $Y=3.15
+ $X2=9.145 $Y2=3.075
r231 27 28 1192.18 $w=1.5e-07 $l=2.325e-06 $layer=POLY_cond $X=9.055 $Y=3.15
+ $X2=6.73 $Y2=3.15
r232 24 26 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.64 $Y=2.8 $X2=6.64
+ $Y2=2.515
r233 23 43 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=6.64 $Y=3.075
+ $X2=6.64 $Y2=3.15
r234 22 24 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.64 $Y=2.89 $X2=6.64
+ $Y2=2.8
r235 22 23 71.9113 $w=1.8e-07 $l=1.85e-07 $layer=POLY_cond $X=6.64 $Y=2.89
+ $X2=6.64 $Y2=3.075
r236 19 21 99.6133 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=6.095 $Y=1.115
+ $X2=6.095 $Y2=0.805
r237 18 64 37.7859 $w=5.23e-07 $l=5.69122e-07 $layer=POLY_cond $X=5.71 $Y=1.225
+ $X2=5.33 $Y2=1.635
r238 17 19 28.2037 $w=2.2e-07 $l=1.42653e-07 $layer=POLY_cond $X=6.02 $Y=1.225
+ $X2=6.095 $Y2=1.115
r239 17 18 90.4236 $w=2.2e-07 $l=3.1e-07 $layer=POLY_cond $X=6.02 $Y=1.225
+ $X2=5.71 $Y2=1.225
r240 15 43 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=6.55 $Y=3.15 $X2=6.64
+ $Y2=3.15
r241 15 16 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=6.55 $Y=3.15
+ $X2=5.69 $Y2=3.15
r242 14 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.615 $Y=3.075
+ $X2=5.69 $Y2=3.15
r243 13 64 46.2206 $w=2.61e-07 $l=3.86814e-07 $layer=POLY_cond $X=5.615 $Y=1.875
+ $X2=5.33 $Y2=1.635
r244 13 14 615.319 $w=1.5e-07 $l=1.2e-06 $layer=POLY_cond $X=5.615 $Y=1.875
+ $X2=5.615 $Y2=3.075
r245 10 18 44.3687 $w=5.23e-07 $l=6.50961e-07 $layer=POLY_cond $X=5.145 $Y=1.41
+ $X2=5.71 $Y2=1.225
r246 10 12 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=5.145 $Y=1.41
+ $X2=5.145 $Y2=0.965
r247 7 64 46.2206 $w=2.61e-07 $l=3.37639e-07 $layer=POLY_cond $X=5.095 $Y=1.875
+ $X2=5.33 $Y2=1.635
r248 7 9 187.98 $w=1.5e-07 $l=5.85e-07 $layer=POLY_cond $X=5.095 $Y=1.875
+ $X2=5.095 $Y2=2.46
r249 2 60 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=4.275
+ $Y=1.96 $X2=4.42 $Y2=2.085
r250 1 55 182 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_NDIFF $count=1 $X=4.175
+ $Y=0.49 $X2=4.32 $Y2=0.665
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTP_1%A_1997_272# 1 2 9 11 12 13 15 16 20 24 26
+ 27 29 34 36 37 39
c117 34 0 6.31244e-20 $X=10.315 $Y=1.525
c118 29 0 1.53844e-19 $X=11.65 $Y=1.445
c119 16 0 6.72618e-20 $X=11.14 $Y=1.53
r120 36 37 10.5766 $w=3.63e-07 $l=2.3e-07 $layer=LI1_cond $X=11.127 $Y=2.75
+ $X2=11.127 $Y2=2.52
r121 31 34 10.2135 $w=1.78e-07 $l=1.65e-07 $layer=LI1_cond $X=10.15 $Y=1.525
+ $X2=10.315 $Y2=1.525
r122 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.15
+ $Y=1.525 $X2=10.15 $Y2=1.525
r123 28 29 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=11.65 $Y=0.925
+ $X2=11.65 $Y2=1.445
r124 26 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.565 $Y=0.84
+ $X2=11.65 $Y2=0.925
r125 26 27 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=11.565 $Y=0.84
+ $X2=11.34 $Y2=0.84
r126 25 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.31 $Y=1.53
+ $X2=11.225 $Y2=1.53
r127 24 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.565 $Y=1.53
+ $X2=11.65 $Y2=1.445
r128 24 25 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=11.565 $Y=1.53
+ $X2=11.31 $Y2=1.53
r129 22 39 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.225 $Y=1.615
+ $X2=11.225 $Y2=1.53
r130 22 37 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=11.225 $Y=1.615
+ $X2=11.225 $Y2=2.52
r131 18 27 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=11.175 $Y=0.755
+ $X2=11.34 $Y2=0.84
r132 18 20 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=11.175 $Y=0.755
+ $X2=11.175 $Y2=0.58
r133 16 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.14 $Y=1.53
+ $X2=11.225 $Y2=1.53
r134 16 34 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=11.14 $Y=1.53
+ $X2=10.315 $Y2=1.53
r135 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=10.31 $Y=2.465
+ $X2=10.31 $Y2=2.75
r136 12 13 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=10.31 $Y=2.375
+ $X2=10.31 $Y2=2.465
r137 11 32 58.2622 $w=3e-07 $l=3.69317e-07 $layer=POLY_cond $X=10.31 $Y=1.84
+ $X2=10.192 $Y2=1.525
r138 11 12 207.96 $w=1.8e-07 $l=5.35e-07 $layer=POLY_cond $X=10.31 $Y=1.84
+ $X2=10.31 $Y2=2.375
r139 7 32 38.5519 $w=3e-07 $l=1.87029e-07 $layer=POLY_cond $X=10.145 $Y=1.36
+ $X2=10.192 $Y2=1.525
r140 7 9 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=10.145 $Y=1.36
+ $X2=10.145 $Y2=0.58
r141 2 36 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=10.96
+ $Y=2.54 $X2=11.11 $Y2=2.75
r142 1 20 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=11.035
+ $Y=0.37 $X2=11.175 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTP_1%A_1745_74# 1 2 9 12 14 15 17 18 19 20 22 24
+ 27 29 30 35 37 40 41 43 45 48 50 52
c167 50 0 5.21422e-20 $X=11.23 $Y=1.185
c168 43 0 1.05093e-19 $X=10.23 $Y=2.55
c169 12 0 1.53844e-19 $X=11.32 $Y=1.84
r170 51 56 13.6415 $w=3.18e-07 $l=9e-08 $layer=POLY_cond $X=11.23 $Y=1.145
+ $X2=11.32 $Y2=1.145
r171 50 52 10.2135 $w=1.78e-07 $l=1.65e-07 $layer=LI1_cond $X=11.23 $Y=1.185
+ $X2=11.065 $Y2=1.185
r172 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.23
+ $Y=1.185 $X2=11.23 $Y2=1.185
r173 45 47 9.9702 $w=3.48e-07 $l=2.1e-07 $layer=LI1_cond $X=9.58 $Y=0.56
+ $X2=9.58 $Y2=0.77
r174 42 43 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=10.23 $Y=1.955
+ $X2=10.23 $Y2=2.55
r175 40 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.145 $Y=1.87
+ $X2=10.23 $Y2=1.955
r176 40 41 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=10.145 $Y=1.87
+ $X2=9.755 $Y2=1.87
r177 39 48 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.755 $Y=1.18
+ $X2=9.67 $Y2=1.18
r178 39 52 85.4652 $w=1.68e-07 $l=1.31e-06 $layer=LI1_cond $X=9.755 $Y=1.18
+ $X2=11.065 $Y2=1.18
r179 37 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.67 $Y=1.785
+ $X2=9.755 $Y2=1.87
r180 36 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.67 $Y=1.265
+ $X2=9.67 $Y2=1.18
r181 36 37 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=9.67 $Y=1.265
+ $X2=9.67 $Y2=1.785
r182 35 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.67 $Y=1.095
+ $X2=9.67 $Y2=1.18
r183 35 47 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=9.67 $Y=1.095
+ $X2=9.67 $Y2=0.77
r184 30 43 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=10.145 $Y=2.715
+ $X2=10.23 $Y2=2.55
r185 30 32 20.4297 $w=3.28e-07 $l=5.85e-07 $layer=LI1_cond $X=10.145 $Y=2.715
+ $X2=9.56 $Y2=2.715
r186 25 27 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=11.955 $Y=1.2
+ $X2=11.955 $Y2=0.645
r187 22 24 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=11.92 $Y=2.045
+ $X2=11.92 $Y2=2.54
r188 21 29 6.66866 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=11.425 $Y=1.915
+ $X2=11.335 $Y2=1.915
r189 20 22 26.9307 $w=1.5e-07 $l=1.69115e-07 $layer=POLY_cond $X=11.83 $Y=1.915
+ $X2=11.92 $Y2=2.045
r190 20 21 207.67 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=11.83 $Y=1.915
+ $X2=11.425 $Y2=1.915
r191 19 56 24.9017 $w=3.18e-07 $l=1.63248e-07 $layer=POLY_cond $X=11.395
+ $Y=1.275 $X2=11.32 $Y2=1.145
r192 18 25 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=11.88 $Y=1.275
+ $X2=11.955 $Y2=1.2
r193 18 19 248.691 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=11.88 $Y=1.275
+ $X2=11.395 $Y2=1.275
r194 15 17 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=11.335 $Y=2.465
+ $X2=11.335 $Y2=2.75
r195 14 15 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=11.335 $Y=2.375
+ $X2=11.335 $Y2=2.465
r196 13 29 18.8402 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=11.335 $Y=1.99
+ $X2=11.335 $Y2=1.915
r197 13 14 149.653 $w=1.8e-07 $l=3.85e-07 $layer=POLY_cond $X=11.335 $Y=1.99
+ $X2=11.335 $Y2=2.375
r198 12 29 18.8402 $w=1.65e-07 $l=8.21584e-08 $layer=POLY_cond $X=11.32 $Y=1.84
+ $X2=11.335 $Y2=1.915
r199 11 56 20.3436 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=11.32 $Y=1.35
+ $X2=11.32 $Y2=1.145
r200 11 12 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=11.32 $Y=1.35
+ $X2=11.32 $Y2=1.84
r201 7 51 40.9245 $w=3.18e-07 $l=3.5812e-07 $layer=POLY_cond $X=10.96 $Y=0.94
+ $X2=11.23 $Y2=1.145
r202 7 9 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=10.96 $Y=0.94
+ $X2=10.96 $Y2=0.58
r203 2 32 600 $w=1.7e-07 $l=1.13737e-06 $layer=licon1_PDIFF $count=1 $X=9.22
+ $Y=1.735 $X2=9.56 $Y2=2.715
r204 1 45 182 $w=1.7e-07 $l=9.35187e-07 $layer=licon1_NDIFF $count=1 $X=8.725
+ $Y=0.37 $X2=9.57 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTP_1%A_2399_424# 1 2 7 9 12 15 19 23 29 32 33
r47 29 30 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=12.745
+ $Y=1.465 $X2=12.745 $Y2=1.465
r48 27 33 0.189605 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=12.335 $Y=1.465
+ $X2=12.21 $Y2=1.465
r49 27 29 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=12.335 $Y=1.465
+ $X2=12.745 $Y2=1.465
r50 25 33 6.72893 $w=2.37e-07 $l=1.71377e-07 $layer=LI1_cond $X=12.197 $Y=1.63
+ $X2=12.21 $Y2=1.465
r51 25 32 24.0733 $w=2.23e-07 $l=4.7e-07 $layer=LI1_cond $X=12.197 $Y=1.63
+ $X2=12.197 $Y2=2.1
r52 21 33 6.72893 $w=2.37e-07 $l=1.65e-07 $layer=LI1_cond $X=12.21 $Y=1.3
+ $X2=12.21 $Y2=1.465
r53 21 23 30.194 $w=2.48e-07 $l=6.55e-07 $layer=LI1_cond $X=12.21 $Y=1.3
+ $X2=12.21 $Y2=0.645
r54 19 32 6.93655 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=12.145 $Y=2.265
+ $X2=12.145 $Y2=2.1
r55 15 30 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=12.84 $Y=1.465
+ $X2=12.745 $Y2=1.465
r56 15 16 66.2869 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=12.93 $Y=1.465
+ $X2=12.93 $Y2=1.3
r57 12 16 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=12.945 $Y=0.74
+ $X2=12.945 $Y2=1.3
r58 7 15 118.763 $w=1.8e-07 $l=3e-07 $layer=POLY_cond $X=12.93 $Y=1.765
+ $X2=12.93 $Y2=1.465
r59 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=12.93 $Y=1.765
+ $X2=12.93 $Y2=2.4
r60 2 19 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=11.995
+ $Y=2.12 $X2=12.145 $Y2=2.265
r61 1 23 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=12.03
+ $Y=0.37 $X2=12.17 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTP_1%VPWR 1 2 3 4 5 6 7 8 27 31 35 39 41 45 51
+ 55 61 66 67 69 70 72 73 74 76 81 93 110 116 117 120 123 126 129 132
c167 2 0 1.19423e-19 $X=3.11 $Y=2.32
r168 132 133 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r169 129 130 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r170 127 130 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=8.4 $Y2=3.33
r171 126 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r172 123 124 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r173 120 121 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r174 117 133 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=3.33
+ $X2=12.72 $Y2=3.33
r175 116 117 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=3.33
+ $X2=13.2 $Y2=3.33
r176 114 132 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.87 $Y=3.33
+ $X2=12.705 $Y2=3.33
r177 114 116 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=12.87 $Y=3.33
+ $X2=13.2 $Y2=3.33
r178 113 133 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=12.72 $Y2=3.33
r179 112 113 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r180 110 132 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.54 $Y=3.33
+ $X2=12.705 $Y2=3.33
r181 110 112 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=12.54 $Y=3.33
+ $X2=12.24 $Y2=3.33
r182 109 113 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=12.24 $Y2=3.33
r183 108 109 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r184 106 109 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=11.28 $Y2=3.33
r185 105 106 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r186 103 106 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=10.32 $Y2=3.33
r187 103 130 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=8.4 $Y2=3.33
r188 102 105 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=8.88 $Y=3.33
+ $X2=10.32 $Y2=3.33
r189 102 103 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r190 100 129 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.555 $Y=3.33
+ $X2=8.47 $Y2=3.33
r191 100 102 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=8.555 $Y=3.33
+ $X2=8.88 $Y2=3.33
r192 99 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.44 $Y2=3.33
r193 98 99 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r194 95 98 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=5.04 $Y=3.33
+ $X2=6.96 $Y2=3.33
r195 95 96 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r196 93 126 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=7.205 $Y=3.33
+ $X2=7.372 $Y2=3.33
r197 93 98 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=7.205 $Y=3.33
+ $X2=6.96 $Y2=3.33
r198 92 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r199 91 92 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r200 89 92 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r201 89 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r202 88 91 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.6 $Y=3.33 $X2=4.56
+ $Y2=3.33
r203 88 89 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r204 86 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.425 $Y=3.33
+ $X2=3.26 $Y2=3.33
r205 86 88 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.425 $Y=3.33
+ $X2=3.6 $Y2=3.33
r206 85 124 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=3.12 $Y2=3.33
r207 85 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r208 84 85 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r209 82 120 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=0.78 $Y2=3.33
r210 82 84 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=1.2 $Y2=3.33
r211 81 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.095 $Y=3.33
+ $X2=3.26 $Y2=3.33
r212 81 84 123.631 $w=1.68e-07 $l=1.895e-06 $layer=LI1_cond $X=3.095 $Y=3.33
+ $X2=1.2 $Y2=3.33
r213 79 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r214 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r215 76 120 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.78 $Y2=3.33
r216 76 78 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.24 $Y2=3.33
r217 74 99 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=6.72 $Y=3.33
+ $X2=6.96 $Y2=3.33
r218 74 96 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=6.72 $Y=3.33
+ $X2=5.04 $Y2=3.33
r219 72 108 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=11.48 $Y=3.33
+ $X2=11.28 $Y2=3.33
r220 72 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.48 $Y=3.33
+ $X2=11.645 $Y2=3.33
r221 71 112 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=11.81 $Y=3.33
+ $X2=12.24 $Y2=3.33
r222 71 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.81 $Y=3.33
+ $X2=11.645 $Y2=3.33
r223 69 105 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=10.485 $Y=3.33
+ $X2=10.32 $Y2=3.33
r224 69 70 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.485 $Y=3.33
+ $X2=10.61 $Y2=3.33
r225 68 108 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=10.735 $Y=3.33
+ $X2=11.28 $Y2=3.33
r226 68 70 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.735 $Y=3.33
+ $X2=10.61 $Y2=3.33
r227 66 91 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=4.705 $Y=3.33
+ $X2=4.56 $Y2=3.33
r228 66 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.705 $Y=3.33
+ $X2=4.87 $Y2=3.33
r229 65 95 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=5.035 $Y=3.33
+ $X2=5.04 $Y2=3.33
r230 65 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.035 $Y=3.33
+ $X2=4.87 $Y2=3.33
r231 61 64 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=12.705 $Y=1.985
+ $X2=12.705 $Y2=2.815
r232 59 132 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.705 $Y=3.245
+ $X2=12.705 $Y2=3.33
r233 59 64 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=12.705 $Y=3.245
+ $X2=12.705 $Y2=2.815
r234 55 58 19.2074 $w=3.28e-07 $l=5.5e-07 $layer=LI1_cond $X=11.645 $Y=2.265
+ $X2=11.645 $Y2=2.815
r235 53 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.645 $Y=3.245
+ $X2=11.645 $Y2=3.33
r236 53 58 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=11.645 $Y=3.245
+ $X2=11.645 $Y2=2.815
r237 49 70 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=10.61 $Y=3.245
+ $X2=10.61 $Y2=3.33
r238 49 51 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=10.61 $Y=3.245
+ $X2=10.61 $Y2=2.75
r239 45 48 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=8.47 $Y=1.91
+ $X2=8.47 $Y2=2.59
r240 43 129 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.47 $Y=3.245
+ $X2=8.47 $Y2=3.33
r241 43 48 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=8.47 $Y=3.245
+ $X2=8.47 $Y2=2.59
r242 42 126 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=7.54 $Y=3.33
+ $X2=7.372 $Y2=3.33
r243 41 129 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.385 $Y=3.33
+ $X2=8.47 $Y2=3.33
r244 41 42 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=8.385 $Y=3.33
+ $X2=7.54 $Y2=3.33
r245 37 126 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=7.372 $Y=3.245
+ $X2=7.372 $Y2=3.33
r246 37 39 14.4485 $w=3.33e-07 $l=4.2e-07 $layer=LI1_cond $X=7.372 $Y=3.245
+ $X2=7.372 $Y2=2.825
r247 33 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.87 $Y=3.245
+ $X2=4.87 $Y2=3.33
r248 33 35 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=4.87 $Y=3.245
+ $X2=4.87 $Y2=2.835
r249 29 123 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.26 $Y=3.245
+ $X2=3.26 $Y2=3.33
r250 29 31 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=3.26 $Y=3.245
+ $X2=3.26 $Y2=2.79
r251 25 120 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=3.245
+ $X2=0.78 $Y2=3.33
r252 25 27 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=0.78 $Y=3.245
+ $X2=0.78 $Y2=2.465
r253 8 64 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=12.56
+ $Y=1.84 $X2=12.705 $Y2=2.815
r254 8 61 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=12.56
+ $Y=1.84 $X2=12.705 $Y2=1.985
r255 7 58 600 $w=1.7e-07 $l=3.745e-07 $layer=licon1_PDIFF $count=1 $X=11.41
+ $Y=2.54 $X2=11.645 $Y2=2.815
r256 7 55 600 $w=1.7e-07 $l=3.745e-07 $layer=licon1_PDIFF $count=1 $X=11.41
+ $Y=2.54 $X2=11.645 $Y2=2.265
r257 6 51 600 $w=1.7e-07 $l=2.8801e-07 $layer=licon1_PDIFF $count=1 $X=10.385
+ $Y=2.54 $X2=10.57 $Y2=2.75
r258 5 48 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=8.325
+ $Y=1.735 $X2=8.47 $Y2=2.59
r259 5 45 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=8.325
+ $Y=1.735 $X2=8.47 $Y2=1.91
r260 4 39 600 $w=1.7e-07 $l=6.26578e-07 $layer=licon1_PDIFF $count=1 $X=7.135
+ $Y=2.305 $X2=7.37 $Y2=2.825
r261 3 35 600 $w=1.7e-07 $l=9.47035e-07 $layer=licon1_PDIFF $count=1 $X=4.72
+ $Y=1.96 $X2=4.87 $Y2=2.835
r262 2 31 600 $w=1.7e-07 $l=5.39815e-07 $layer=licon1_PDIFF $count=1 $X=3.11
+ $Y=2.32 $X2=3.26 $Y2=2.79
r263 1 27 300 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=2 $X=0.58
+ $Y=2.32 $X2=0.78 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTP_1%A_300_464# 1 2 3 4 5 16 20 22 25 28 29 30
+ 34 37 39 40 41 42 43 45 48 50 56
c169 56 0 8.81023e-20 $X=3.83 $Y=2.475
c170 40 0 1.55517e-19 $X=6.37 $Y=1.285
c171 28 0 1.94423e-19 $X=4.555 $Y=2.52
c172 25 0 1.19423e-19 $X=3.53 $Y=2.33
r173 54 56 15.9825 $w=2.29e-07 $l=3e-07 $layer=LI1_cond $X=3.53 $Y=2.475
+ $X2=3.83 $Y2=2.475
r174 50 52 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=2.435 $Y=0.68
+ $X2=2.435 $Y2=1.005
r175 47 48 10.4785 $w=6.33e-07 $l=1.7e-07 $layer=LI1_cond $X=2.385 $Y=2.662
+ $X2=2.555 $Y2=2.662
r176 44 45 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=6.455 $Y=1.37
+ $X2=6.455 $Y2=2.045
r177 42 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.37 $Y=2.13
+ $X2=6.455 $Y2=2.045
r178 42 43 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=6.37 $Y=2.13
+ $X2=6.075 $Y2=2.13
r179 40 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.37 $Y=1.285
+ $X2=6.455 $Y2=1.37
r180 40 41 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=6.37 $Y=1.285
+ $X2=5.975 $Y2=1.285
r181 39 59 3.21189 $w=2.5e-07 $l=1.7e-07 $layer=LI1_cond $X=5.95 $Y=2.385
+ $X2=5.95 $Y2=2.555
r182 38 43 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.95 $Y=2.215
+ $X2=6.075 $Y2=2.13
r183 38 39 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=5.95 $Y=2.215
+ $X2=5.95 $Y2=2.385
r184 37 41 6.81835 $w=1.7e-07 $l=1.23386e-07 $layer=LI1_cond $X=5.887 $Y=1.2
+ $X2=5.975 $Y2=1.285
r185 37 57 12.9922 $w=1.73e-07 $l=2.05e-07 $layer=LI1_cond $X=5.887 $Y=1.2
+ $X2=5.887 $Y2=0.995
r186 32 57 5.54545 $w=1.78e-07 $l=9e-08 $layer=LI1_cond $X=5.885 $Y=0.905
+ $X2=5.885 $Y2=0.995
r187 32 34 5.85354 $w=1.78e-07 $l=9.5e-08 $layer=LI1_cond $X=5.885 $Y=0.905
+ $X2=5.885 $Y2=0.81
r188 30 59 3.74091 $w=1.95e-07 $l=1.57321e-07 $layer=LI1_cond $X=5.825 $Y=2.482
+ $X2=5.95 $Y2=2.555
r189 30 31 67.1142 $w=1.93e-07 $l=1.18e-06 $layer=LI1_cond $X=5.825 $Y=2.482
+ $X2=4.645 $Y2=2.482
r190 29 56 22.6032 $w=2.29e-07 $l=4.41928e-07 $layer=LI1_cond $X=4.25 $Y=2.52
+ $X2=3.83 $Y2=2.475
r191 28 31 5.46269 $w=2.01e-07 $l=1.07331e-07 $layer=LI1_cond $X=4.555 $Y=2.52
+ $X2=4.645 $Y2=2.482
r192 28 29 16.9136 $w=1.98e-07 $l=3.05e-07 $layer=LI1_cond $X=4.555 $Y=2.52
+ $X2=4.25 $Y2=2.52
r193 25 54 2.48377 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=3.53 $Y=2.33
+ $X2=3.53 $Y2=2.475
r194 24 25 80.8984 $w=1.68e-07 $l=1.24e-06 $layer=LI1_cond $X=3.53 $Y=1.09
+ $X2=3.53 $Y2=2.33
r195 23 52 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.6 $Y=1.005
+ $X2=2.435 $Y2=1.005
r196 22 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.445 $Y=1.005
+ $X2=3.53 $Y2=1.09
r197 22 23 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=3.445 $Y=1.005
+ $X2=2.6 $Y2=1.005
r198 20 54 5.36381 $w=2.29e-07 $l=1.05119e-07 $layer=LI1_cond $X=3.445 $Y=2.43
+ $X2=3.53 $Y2=2.475
r199 20 48 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=3.445 $Y=2.43
+ $X2=2.555 $Y2=2.43
r200 16 47 2.76887 $w=6.33e-07 $l=1.47e-07 $layer=LI1_cond $X=2.238 $Y=2.662
+ $X2=2.385 $Y2=2.662
r201 16 18 11.0755 $w=6.33e-07 $l=5.88e-07 $layer=LI1_cond $X=2.238 $Y=2.662
+ $X2=1.65 $Y2=2.662
r202 5 59 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=5.765
+ $Y=2.285 $X2=5.91 $Y2=2.495
r203 4 56 300 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=2 $X=3.68
+ $Y=2.32 $X2=3.83 $Y2=2.475
r204 3 47 200 $w=1.7e-07 $l=9.54751e-07 $layer=licon1_PDIFF $count=3 $X=1.5
+ $Y=2.32 $X2=2.385 $Y2=2.465
r205 3 18 200 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=3 $X=1.5
+ $Y=2.32 $X2=1.65 $Y2=2.465
r206 2 34 182 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_NDIFF $count=1 $X=5.755
+ $Y=0.595 $X2=5.88 $Y2=0.81
r207 1 50 182 $w=1.7e-07 $l=6.07124e-07 $layer=licon1_NDIFF $count=1 $X=1.95
+ $Y=0.405 $X2=2.435 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTP_1%Q 1 2 7 8 9 10 11 12 13 29
r15 22 29 1.3969 $w=3.28e-07 $l=4e-08 $layer=LI1_cond $X=13.16 $Y=0.965
+ $X2=13.16 $Y2=0.925
r16 12 13 16.7217 $w=2.53e-07 $l=3.7e-07 $layer=LI1_cond $X=13.197 $Y=2.405
+ $X2=13.197 $Y2=2.775
r17 11 12 18.9814 $w=2.53e-07 $l=4.2e-07 $layer=LI1_cond $X=13.197 $Y=1.985
+ $X2=13.197 $Y2=2.405
r18 10 11 14.462 $w=2.53e-07 $l=3.2e-07 $layer=LI1_cond $X=13.197 $Y=1.665
+ $X2=13.197 $Y2=1.985
r19 9 10 16.7217 $w=2.53e-07 $l=3.7e-07 $layer=LI1_cond $X=13.197 $Y=1.295
+ $X2=13.197 $Y2=1.665
r20 9 45 7.45698 $w=2.53e-07 $l=1.65e-07 $layer=LI1_cond $X=13.197 $Y=1.295
+ $X2=13.197 $Y2=1.13
r21 8 45 5.6192 $w=3.28e-07 $l=1.43e-07 $layer=LI1_cond $X=13.16 $Y=0.987
+ $X2=13.16 $Y2=1.13
r22 8 22 0.768295 $w=3.28e-07 $l=2.2e-08 $layer=LI1_cond $X=13.16 $Y=0.987
+ $X2=13.16 $Y2=0.965
r23 8 29 0.803218 $w=3.28e-07 $l=2.3e-08 $layer=LI1_cond $X=13.16 $Y=0.902
+ $X2=13.16 $Y2=0.925
r24 7 8 13.515 $w=3.28e-07 $l=3.87e-07 $layer=LI1_cond $X=13.16 $Y=0.515
+ $X2=13.16 $Y2=0.902
r25 2 13 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=13.005
+ $Y=1.84 $X2=13.155 $Y2=2.815
r26 2 11 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=13.005
+ $Y=1.84 $X2=13.155 $Y2=1.985
r27 1 7 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=13.02
+ $Y=0.37 $X2=13.16 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTP_1%VGND 1 2 3 4 5 6 7 24 28 32 36 40 44 47 48
+ 49 51 56 65 69 77 82 89 90 93 96 100 106 109 112
c133 90 0 7.12888e-20 $X=13.2 $Y=0
c134 28 0 1.58089e-19 $X=3.715 $Y=0.565
r135 112 113 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r136 109 110 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r137 106 107 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r138 100 103 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=7.595 $Y=0
+ $X2=7.595 $Y2=0.325
r139 100 101 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r140 96 97 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r141 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r142 90 113 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=0
+ $X2=12.72 $Y2=0
r143 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=0 $X2=13.2
+ $Y2=0
r144 87 112 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.815 $Y=0
+ $X2=12.69 $Y2=0
r145 87 89 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=12.815 $Y=0
+ $X2=13.2 $Y2=0
r146 86 113 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=12.72 $Y2=0
r147 86 110 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=11.76 $Y2=0
r148 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r149 83 109 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=11.905 $Y=0
+ $X2=11.737 $Y2=0
r150 83 85 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=11.905 $Y=0
+ $X2=12.24 $Y2=0
r151 82 112 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.565 $Y=0
+ $X2=12.69 $Y2=0
r152 82 85 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=12.565 $Y=0
+ $X2=12.24 $Y2=0
r153 81 110 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=11.76 $Y2=0
r154 81 107 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=10.32 $Y2=0
r155 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r156 78 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.525 $Y=0
+ $X2=10.36 $Y2=0
r157 78 80 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=10.525 $Y=0
+ $X2=11.28 $Y2=0
r158 77 109 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=11.57 $Y=0
+ $X2=11.737 $Y2=0
r159 77 80 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=11.57 $Y=0
+ $X2=11.28 $Y2=0
r160 76 107 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=10.32 $Y2=0
r161 75 76 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=9.84 $Y=0
+ $X2=9.84 $Y2=0
r162 73 76 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=7.92 $Y=0
+ $X2=9.84 $Y2=0
r163 73 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0
+ $X2=7.44 $Y2=0
r164 72 75 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=7.92 $Y=0 $X2=9.84
+ $Y2=0
r165 72 73 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r166 70 100 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.76 $Y=0
+ $X2=7.595 $Y2=0
r167 70 72 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=7.76 $Y=0 $X2=7.92
+ $Y2=0
r168 69 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.195 $Y=0
+ $X2=10.36 $Y2=0
r169 69 75 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=10.195 $Y=0
+ $X2=9.84 $Y2=0
r170 67 68 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r171 65 100 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.43 $Y=0
+ $X2=7.595 $Y2=0
r172 65 67 155.925 $w=1.68e-07 $l=2.39e-06 $layer=LI1_cond $X=7.43 $Y=0 $X2=5.04
+ $Y2=0
r173 64 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r174 64 97 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=3.6
+ $Y2=0
r175 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r176 61 96 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=3.88 $Y=0 $X2=3.735
+ $Y2=0
r177 61 63 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.88 $Y=0 $X2=4.56
+ $Y2=0
r178 60 97 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=3.6
+ $Y2=0
r179 60 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r180 59 60 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r181 57 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=0.71
+ $Y2=0
r182 57 59 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=1.2
+ $Y2=0
r183 56 96 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=3.59 $Y=0 $X2=3.735
+ $Y2=0
r184 56 59 155.925 $w=1.68e-07 $l=2.39e-06 $layer=LI1_cond $X=3.59 $Y=0 $X2=1.2
+ $Y2=0
r185 54 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r186 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r187 51 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.71
+ $Y2=0
r188 51 53 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0
+ $X2=0.24 $Y2=0
r189 49 101 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=6.72 $Y=0
+ $X2=7.44 $Y2=0
r190 49 68 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=6.72 $Y=0
+ $X2=5.04 $Y2=0
r191 47 63 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=4.705 $Y=0
+ $X2=4.56 $Y2=0
r192 47 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.705 $Y=0 $X2=4.87
+ $Y2=0
r193 46 67 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=5.035 $Y=0 $X2=5.04
+ $Y2=0
r194 46 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.035 $Y=0 $X2=4.87
+ $Y2=0
r195 42 112 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=12.69 $Y=0.085
+ $X2=12.69 $Y2=0
r196 42 44 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=12.69 $Y=0.085
+ $X2=12.69 $Y2=0.515
r197 38 109 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=11.737 $Y=0.085
+ $X2=11.737 $Y2=0
r198 38 40 14.2765 $w=3.33e-07 $l=4.15e-07 $layer=LI1_cond $X=11.737 $Y=0.085
+ $X2=11.737 $Y2=0.5
r199 34 106 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.36 $Y=0.085
+ $X2=10.36 $Y2=0
r200 34 36 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=10.36 $Y=0.085
+ $X2=10.36 $Y2=0.58
r201 30 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.87 $Y=0.085
+ $X2=4.87 $Y2=0
r202 30 32 20.2551 $w=3.28e-07 $l=5.8e-07 $layer=LI1_cond $X=4.87 $Y=0.085
+ $X2=4.87 $Y2=0.665
r203 26 96 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.735 $Y=0.085
+ $X2=3.735 $Y2=0
r204 26 28 19.0749 $w=2.88e-07 $l=4.8e-07 $layer=LI1_cond $X=3.735 $Y=0.085
+ $X2=3.735 $Y2=0.565
r205 22 93 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0
r206 22 24 19.7312 $w=3.28e-07 $l=5.65e-07 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0.65
r207 7 44 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=12.585
+ $Y=0.37 $X2=12.73 $Y2=0.515
r208 6 40 182 $w=1.7e-07 $l=1.99687e-07 $layer=licon1_NDIFF $count=1 $X=11.59
+ $Y=0.37 $X2=11.735 $Y2=0.5
r209 5 36 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=10.22
+ $Y=0.37 $X2=10.36 $Y2=0.58
r210 4 103 182 $w=1.7e-07 $l=3.63731e-07 $layer=licon1_NDIFF $count=1 $X=7.375
+ $Y=0.595 $X2=7.595 $Y2=0.325
r211 3 32 182 $w=1.7e-07 $l=2.32379e-07 $layer=licon1_NDIFF $count=1 $X=4.67
+ $Y=0.595 $X2=4.87 $Y2=0.665
r212 2 28 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=3.575
+ $Y=0.405 $X2=3.715 $Y2=0.565
r213 1 24 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.44 $X2=0.71 $Y2=0.65
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTP_1%noxref_24 1 2 7 9 14
r32 14 17 7.40856 $w=3.48e-07 $l=2.25e-07 $layer=LI1_cond $X=3.235 $Y=0.34
+ $X2=3.235 $Y2=0.565
r33 9 12 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=1.27 $Y=0.34 $X2=1.27
+ $Y2=0.55
r34 8 9 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.435 $Y=0.34 $X2=1.27
+ $Y2=0.34
r35 7 14 4.974 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=3.06 $Y=0.34 $X2=3.235
+ $Y2=0.34
r36 7 8 106.016 $w=1.68e-07 $l=1.625e-06 $layer=LI1_cond $X=3.06 $Y=0.34
+ $X2=1.435 $Y2=0.34
r37 2 17 182 $w=1.7e-07 $l=2.22711e-07 $layer=licon1_NDIFF $count=1 $X=3.115
+ $Y=0.405 $X2=3.265 $Y2=0.565
r38 1 12 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=1.125
+ $Y=0.405 $X2=1.27 $Y2=0.55
.ends

