* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
X0 VGND A3 a_355_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X1 a_45_264# B1 a_661_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X2 a_346_368# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 a_661_74# B2 VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X4 VPWR a_45_264# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X5 VPWR A1 a_346_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 X a_45_264# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X7 VPWR A3 a_346_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 a_355_74# A2 a_433_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X9 VGND a_45_264# X VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X10 X a_45_264# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X11 a_346_368# B1 a_45_264# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 a_45_264# B2 a_346_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 a_433_74# A1 a_45_264# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
.ends
