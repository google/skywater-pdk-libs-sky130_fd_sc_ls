* File: sky130_fd_sc_ls__a2111o_2.pex.spice
* Created: Fri Aug 28 12:47:31 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__A2111O_2%A_91_244# 1 2 3 4 13 15 16 18 19 21 22 24
+ 25 26 27 29 30 31 33 37 39 43 45 49 57 58 62
c111 58 0 1.10806e-19 $X=2.885 $Y=1.095
c112 31 0 1.74446e-19 $X=1.92 $Y=2.12
c113 25 0 1.60145e-19 $X=1.275 $Y=1.55
r114 61 62 0.580723 $w=4.15e-07 $l=5e-09 $layer=POLY_cond $X=0.99 $Y=1.492
+ $X2=0.995 $Y2=1.492
r115 60 61 49.9422 $w=4.15e-07 $l=4.3e-07 $layer=POLY_cond $X=0.56 $Y=1.492
+ $X2=0.99 $Y2=1.492
r116 59 60 1.74217 $w=4.15e-07 $l=1.5e-08 $layer=POLY_cond $X=0.545 $Y=1.492
+ $X2=0.56 $Y2=1.492
r117 54 62 23.2289 $w=4.15e-07 $l=2e-07 $layer=POLY_cond $X=1.195 $Y=1.492
+ $X2=0.995 $Y2=1.492
r118 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.195
+ $Y=1.385 $X2=1.195 $Y2=1.385
r119 51 53 13.2509 $w=2.67e-07 $l=2.9e-07 $layer=LI1_cond $X=1.195 $Y=1.095
+ $X2=1.195 $Y2=1.385
r120 47 49 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=4.355 $Y=1.01
+ $X2=4.355 $Y2=0.515
r121 46 58 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.01 $Y=1.095
+ $X2=2.885 $Y2=1.095
r122 45 47 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.19 $Y=1.095
+ $X2=4.355 $Y2=1.01
r123 45 46 76.984 $w=1.68e-07 $l=1.18e-06 $layer=LI1_cond $X=4.19 $Y=1.095
+ $X2=3.01 $Y2=1.095
r124 41 58 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.885 $Y=1.01
+ $X2=2.885 $Y2=1.095
r125 41 43 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=2.885 $Y=1.01
+ $X2=2.885 $Y2=0.515
r126 40 57 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.03 $Y=1.095
+ $X2=1.905 $Y2=1.095
r127 39 58 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.76 $Y=1.095
+ $X2=2.885 $Y2=1.095
r128 39 40 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=2.76 $Y=1.095
+ $X2=2.03 $Y2=1.095
r129 35 57 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.905 $Y=1.01
+ $X2=1.905 $Y2=1.095
r130 35 37 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=1.905 $Y=1.01
+ $X2=1.905 $Y2=0.515
r131 31 56 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.92 $Y=2.12 $X2=1.92
+ $Y2=2.035
r132 31 33 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=1.92 $Y=2.12
+ $X2=1.92 $Y2=2.815
r133 29 56 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.755 $Y=2.035
+ $X2=1.92 $Y2=2.035
r134 29 30 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.755 $Y=2.035
+ $X2=1.36 $Y2=2.035
r135 28 51 3.37873 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.36 $Y=1.095
+ $X2=1.195 $Y2=1.095
r136 27 57 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.78 $Y=1.095
+ $X2=1.905 $Y2=1.095
r137 27 28 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=1.78 $Y=1.095
+ $X2=1.36 $Y2=1.095
r138 26 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.275 $Y=1.95
+ $X2=1.36 $Y2=2.035
r139 25 53 9.14344 $w=2.67e-07 $l=2.0106e-07 $layer=LI1_cond $X=1.275 $Y=1.55
+ $X2=1.195 $Y2=1.385
r140 25 26 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=1.275 $Y=1.55
+ $X2=1.275 $Y2=1.95
r141 22 62 26.7644 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=0.995 $Y=1.765
+ $X2=0.995 $Y2=1.492
r142 22 24 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.995 $Y=1.765
+ $X2=0.995 $Y2=2.4
r143 19 61 26.7644 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=0.99 $Y=1.22
+ $X2=0.99 $Y2=1.492
r144 19 21 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.99 $Y=1.22
+ $X2=0.99 $Y2=0.74
r145 16 60 26.7644 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=0.56 $Y=1.22
+ $X2=0.56 $Y2=1.492
r146 16 18 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.56 $Y=1.22
+ $X2=0.56 $Y2=0.74
r147 13 59 26.7644 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=0.545 $Y=1.765
+ $X2=0.545 $Y2=1.492
r148 13 15 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.545 $Y=1.765
+ $X2=0.545 $Y2=2.4
r149 4 56 400 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=1.795
+ $Y=1.84 $X2=1.92 $Y2=2.115
r150 4 33 400 $w=1.7e-07 $l=1.03562e-06 $layer=licon1_PDIFF $count=1 $X=1.795
+ $Y=1.84 $X2=1.92 $Y2=2.815
r151 3 49 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.215
+ $Y=0.37 $X2=4.355 $Y2=0.515
r152 2 43 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.705
+ $Y=0.37 $X2=2.845 $Y2=0.515
r153 1 37 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=1.82
+ $Y=0.37 $X2=1.945 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__A2111O_2%D1 1 3 6 8 9
c32 1 0 1.60145e-19 $X=2.145 $Y=1.765
r33 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.07
+ $Y=1.515 $X2=2.07 $Y2=1.515
r34 9 14 2.41209 $w=4.28e-07 $l=9e-08 $layer=LI1_cond $X=2.16 $Y=1.565 $X2=2.07
+ $Y2=1.565
r35 8 14 10.4524 $w=4.28e-07 $l=3.9e-07 $layer=LI1_cond $X=1.68 $Y=1.565
+ $X2=2.07 $Y2=1.565
r36 4 13 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=2.16 $Y=1.35
+ $X2=2.07 $Y2=1.515
r37 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.16 $Y=1.35 $X2=2.16
+ $Y2=0.74
r38 1 13 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=2.145 $Y=1.765
+ $X2=2.07 $Y2=1.515
r39 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.145 $Y=1.765
+ $X2=2.145 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__A2111O_2%C1 1 3 6 8 9 10 11 18
c32 1 0 4.31819e-19 $X=2.535 $Y=1.765
r33 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.61
+ $Y=1.515 $X2=2.61 $Y2=1.515
r34 10 11 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.61 $Y=2.405
+ $X2=2.61 $Y2=2.775
r35 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.61 $Y=2.035
+ $X2=2.61 $Y2=2.405
r36 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.61 $Y=1.665 $X2=2.61
+ $Y2=2.035
r37 8 18 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=2.61 $Y=1.665
+ $X2=2.61 $Y2=1.515
r38 4 17 38.5562 $w=2.99e-07 $l=1.74714e-07 $layer=POLY_cond $X=2.63 $Y=1.35
+ $X2=2.61 $Y2=1.515
r39 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.63 $Y=1.35 $X2=2.63
+ $Y2=0.74
r40 1 17 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=2.535 $Y=1.765
+ $X2=2.61 $Y2=1.515
r41 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.535 $Y=1.765
+ $X2=2.535 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__A2111O_2%B1 3 5 7 8 12
r31 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.15
+ $Y=1.515 $X2=3.15 $Y2=1.515
r32 8 12 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=3.15 $Y=1.665
+ $X2=3.15 $Y2=1.515
r33 5 11 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=3.075 $Y=1.765
+ $X2=3.15 $Y2=1.515
r34 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.075 $Y=1.765
+ $X2=3.075 $Y2=2.4
r35 1 11 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=3.06 $Y=1.35
+ $X2=3.15 $Y2=1.515
r36 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.06 $Y=1.35 $X2=3.06
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__A2111O_2%A2 1 3 6 8 9
c31 1 0 1.56668e-19 $X=3.615 $Y=1.765
r32 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.69
+ $Y=1.515 $X2=3.69 $Y2=1.515
r33 9 14 10.4524 $w=4.28e-07 $l=3.9e-07 $layer=LI1_cond $X=4.08 $Y=1.565
+ $X2=3.69 $Y2=1.565
r34 8 14 2.41209 $w=4.28e-07 $l=9e-08 $layer=LI1_cond $X=3.6 $Y=1.565 $X2=3.69
+ $Y2=1.565
r35 4 13 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=3.78 $Y=1.35
+ $X2=3.69 $Y2=1.515
r36 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.78 $Y=1.35 $X2=3.78
+ $Y2=0.74
r37 1 13 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=3.615 $Y=1.765
+ $X2=3.69 $Y2=1.515
r38 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.615 $Y=1.765
+ $X2=3.615 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__A2111O_2%A1 3 5 7 9 10 13 14
c30 14 0 1.56668e-19 $X=4.53 $Y=1.515
r31 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.53
+ $Y=1.515 $X2=4.53 $Y2=1.515
r32 10 14 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=4.53 $Y=1.665
+ $X2=4.53 $Y2=1.515
r33 8 13 49.8355 $w=3.3e-07 $l=2.85e-07 $layer=POLY_cond $X=4.245 $Y=1.515
+ $X2=4.53 $Y2=1.515
r34 8 9 5.03009 $w=3.3e-07 $l=1.08995e-07 $layer=POLY_cond $X=4.245 $Y=1.515
+ $X2=4.155 $Y2=1.557
r35 5 9 37.0704 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=4.155 $Y=1.765
+ $X2=4.155 $Y2=1.557
r36 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.155 $Y=1.765
+ $X2=4.155 $Y2=2.4
r37 1 9 37.0704 $w=1.5e-07 $l=2.14369e-07 $layer=POLY_cond $X=4.14 $Y=1.35
+ $X2=4.155 $Y2=1.557
r38 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.14 $Y=1.35 $X2=4.14
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__A2111O_2%VPWR 1 2 3 10 12 18 22 25 26 27 29 42 43 49
r53 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r54 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r55 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r56 40 43 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r57 39 40 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r58 37 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r59 36 39 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.68 $Y=3.33
+ $X2=3.6 $Y2=3.33
r60 36 37 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r61 34 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.385 $Y=3.33
+ $X2=1.22 $Y2=3.33
r62 34 36 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.385 $Y=3.33
+ $X2=1.68 $Y2=3.33
r63 33 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r64 33 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r65 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r66 30 46 3.96192 $w=1.7e-07 $l=2.03e-07 $layer=LI1_cond $X=0.405 $Y=3.33
+ $X2=0.202 $Y2=3.33
r67 30 32 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.405 $Y=3.33
+ $X2=0.72 $Y2=3.33
r68 29 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.055 $Y=3.33
+ $X2=1.22 $Y2=3.33
r69 29 32 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.055 $Y=3.33
+ $X2=0.72 $Y2=3.33
r70 27 40 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=2.4 $Y=3.33 $X2=3.6
+ $Y2=3.33
r71 27 37 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=1.68 $Y2=3.33
r72 25 39 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=3.675 $Y=3.33
+ $X2=3.6 $Y2=3.33
r73 25 26 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=3.675 $Y=3.33
+ $X2=3.86 $Y2=3.33
r74 24 42 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=4.045 $Y=3.33
+ $X2=4.56 $Y2=3.33
r75 24 26 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=4.045 $Y=3.33
+ $X2=3.86 $Y2=3.33
r76 20 26 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.86 $Y=3.245
+ $X2=3.86 $Y2=3.33
r77 20 22 24.6062 $w=3.68e-07 $l=7.9e-07 $layer=LI1_cond $X=3.86 $Y=3.245
+ $X2=3.86 $Y2=2.455
r78 16 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=3.245
+ $X2=1.22 $Y2=3.33
r79 16 18 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=1.22 $Y=3.245
+ $X2=1.22 $Y2=2.455
r80 12 15 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=0.28 $Y=1.985
+ $X2=0.28 $Y2=2.815
r81 10 46 3.18124 $w=2.5e-07 $l=1.17707e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.202 $Y2=3.33
r82 10 15 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.28 $Y2=2.815
r83 3 22 300 $w=1.7e-07 $l=6.9482e-07 $layer=licon1_PDIFF $count=2 $X=3.69
+ $Y=1.84 $X2=3.86 $Y2=2.455
r84 2 18 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=1.07
+ $Y=1.84 $X2=1.22 $Y2=2.455
r85 1 15 400 $w=1.7e-07 $l=1.03562e-06 $layer=licon1_PDIFF $count=1 $X=0.195
+ $Y=1.84 $X2=0.32 $Y2=2.815
r86 1 12 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.195
+ $Y=1.84 $X2=0.32 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_LS__A2111O_2%X 1 2 9 11 12 13 14 34
c20 11 0 1.2388e-19 $X=0.635 $Y=1.58
r21 20 34 0.542326 $w=2.53e-07 $l=1.2e-08 $layer=LI1_cond $X=0.732 $Y=1.677
+ $X2=0.732 $Y2=1.665
r22 13 14 16.7217 $w=2.53e-07 $l=3.7e-07 $layer=LI1_cond $X=0.732 $Y=2.405
+ $X2=0.732 $Y2=2.775
r23 12 13 18.9814 $w=2.53e-07 $l=4.2e-07 $layer=LI1_cond $X=0.732 $Y=1.985
+ $X2=0.732 $Y2=2.405
r24 11 34 1.67217 $w=2.53e-07 $l=3.7e-08 $layer=LI1_cond $X=0.732 $Y=1.628
+ $X2=0.732 $Y2=1.665
r25 11 32 4.80861 $w=2.53e-07 $l=7.8e-08 $layer=LI1_cond $X=0.732 $Y=1.628
+ $X2=0.732 $Y2=1.55
r26 11 12 12.2927 $w=2.53e-07 $l=2.72e-07 $layer=LI1_cond $X=0.732 $Y=1.713
+ $X2=0.732 $Y2=1.985
r27 11 20 1.62698 $w=2.53e-07 $l=3.6e-08 $layer=LI1_cond $X=0.732 $Y=1.713
+ $X2=0.732 $Y2=1.677
r28 9 32 67.5241 $w=1.68e-07 $l=1.035e-06 $layer=LI1_cond $X=0.775 $Y=0.515
+ $X2=0.775 $Y2=1.55
r29 2 14 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=0.62
+ $Y=1.84 $X2=0.77 $Y2=2.815
r30 2 12 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=0.62
+ $Y=1.84 $X2=0.77 $Y2=1.985
r31 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.635
+ $Y=0.37 $X2=0.775 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__A2111O_2%A_630_368# 1 2 7 9 11 13 15
c26 7 0 1.46567e-19 $X=3.32 $Y=2.12
r27 13 20 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.38 $Y=2.12 $X2=4.38
+ $Y2=2.035
r28 13 15 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=4.38 $Y=2.12
+ $X2=4.38 $Y2=2.815
r29 12 18 5.55669 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=3.505 $Y=2.035
+ $X2=3.32 $Y2=2.035
r30 11 20 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.215 $Y=2.035
+ $X2=4.38 $Y2=2.035
r31 11 12 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=4.215 $Y=2.035
+ $X2=3.505 $Y2=2.035
r32 7 18 2.55307 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.32 $Y=2.12 $X2=3.32
+ $Y2=2.035
r33 7 9 21.6472 $w=3.68e-07 $l=6.95e-07 $layer=LI1_cond $X=3.32 $Y=2.12 $X2=3.32
+ $Y2=2.815
r34 2 20 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=4.23
+ $Y=1.84 $X2=4.38 $Y2=2.115
r35 2 15 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=4.23
+ $Y=1.84 $X2=4.38 $Y2=2.815
r36 1 18 400 $w=1.7e-07 $l=3.49821e-07 $layer=licon1_PDIFF $count=1 $X=3.15
+ $Y=1.84 $X2=3.32 $Y2=2.115
r37 1 9 400 $w=1.7e-07 $l=1.05659e-06 $layer=licon1_PDIFF $count=1 $X=3.15
+ $Y=1.84 $X2=3.32 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_LS__A2111O_2%VGND 1 2 3 4 13 15 19 23 27 30 31 32 34 43
+ 49 50 56 59
r61 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r62 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r63 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r64 50 60 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=3.6
+ $Y2=0
r65 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r66 47 59 11.9488 $w=1.7e-07 $l=2.75e-07 $layer=LI1_cond $X=3.73 $Y=0 $X2=3.455
+ $Y2=0
r67 47 49 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=3.73 $Y=0 $X2=4.56
+ $Y2=0
r68 46 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r69 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r70 43 59 11.9488 $w=1.7e-07 $l=2.75e-07 $layer=LI1_cond $X=3.18 $Y=0 $X2=3.455
+ $Y2=0
r71 43 45 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=3.18 $Y=0 $X2=3.12
+ $Y2=0
r72 42 57 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.2
+ $Y2=0
r73 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r74 39 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.37 $Y=0 $X2=1.205
+ $Y2=0
r75 39 41 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=1.37 $Y=0 $X2=2.16
+ $Y2=0
r76 38 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r77 38 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r78 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r79 35 53 4.60552 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=0.51 $Y=0 $X2=0.255
+ $Y2=0
r80 35 37 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=0.51 $Y=0 $X2=0.72
+ $Y2=0
r81 34 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.04 $Y=0 $X2=1.205
+ $Y2=0
r82 34 37 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.04 $Y=0 $X2=0.72
+ $Y2=0
r83 32 46 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=3.12
+ $Y2=0
r84 32 42 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=2.16
+ $Y2=0
r85 30 41 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=2.21 $Y=0 $X2=2.16
+ $Y2=0
r86 30 31 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=2.21 $Y=0 $X2=2.395
+ $Y2=0
r87 29 45 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=2.58 $Y=0 $X2=3.12
+ $Y2=0
r88 29 31 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=2.58 $Y=0 $X2=2.395
+ $Y2=0
r89 25 59 2.31338 $w=5.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.455 $Y=0.085
+ $X2=3.455 $Y2=0
r90 25 27 12.8307 $w=5.48e-07 $l=5.9e-07 $layer=LI1_cond $X=3.455 $Y=0.085
+ $X2=3.455 $Y2=0.675
r91 21 31 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.395 $Y=0.085
+ $X2=2.395 $Y2=0
r92 21 23 18.3768 $w=3.68e-07 $l=5.9e-07 $layer=LI1_cond $X=2.395 $Y=0.085
+ $X2=2.395 $Y2=0.675
r93 17 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=0.085
+ $X2=1.205 $Y2=0
r94 17 19 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=1.205 $Y=0.085
+ $X2=1.205 $Y2=0.675
r95 13 53 3.16065 $w=3.3e-07 $l=1.25499e-07 $layer=LI1_cond $X=0.345 $Y=0.085
+ $X2=0.255 $Y2=0
r96 13 15 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.345 $Y=0.085
+ $X2=0.345 $Y2=0.515
r97 4 27 182 $w=1.7e-07 $l=4.36635e-07 $layer=licon1_NDIFF $count=1 $X=3.135
+ $Y=0.37 $X2=3.445 $Y2=0.675
r98 3 23 182 $w=1.7e-07 $l=3.76597e-07 $layer=licon1_NDIFF $count=1 $X=2.235
+ $Y=0.37 $X2=2.395 $Y2=0.675
r99 2 19 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=1.065
+ $Y=0.37 $X2=1.205 $Y2=0.675
r100 1 15 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.22
+ $Y=0.37 $X2=0.345 $Y2=0.515
.ends

