* File: sky130_fd_sc_ls__a31o_2.pex.spice
* Created: Fri Aug 28 12:58:46 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__A31O_2%A_97_296# 1 2 9 11 13 16 18 20 22 23 24 25 27
+ 29 33 38 46
c102 18 0 3.54614e-20 $X=1.025 $Y=1.765
r103 45 46 3.71722 $w=3.89e-07 $l=3e-08 $layer=POLY_cond $X=0.995 $Y=1.532
+ $X2=1.025 $Y2=1.532
r104 44 45 52.0411 $w=3.89e-07 $l=4.2e-07 $layer=POLY_cond $X=0.575 $Y=1.532
+ $X2=0.995 $Y2=1.532
r105 43 44 1.23907 $w=3.89e-07 $l=1e-08 $layer=POLY_cond $X=0.565 $Y=1.532
+ $X2=0.575 $Y2=1.532
r106 39 46 11.7712 $w=3.89e-07 $l=9.5e-08 $layer=POLY_cond $X=1.12 $Y=1.532
+ $X2=1.025 $Y2=1.532
r107 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.12
+ $Y=1.465 $X2=1.12 $Y2=1.465
r108 33 35 24.0657 $w=3.38e-07 $l=7.1e-07 $layer=LI1_cond $X=3.555 $Y=1.985
+ $X2=3.555 $Y2=2.695
r109 31 33 3.22006 $w=3.38e-07 $l=9.5e-08 $layer=LI1_cond $X=3.555 $Y=1.89
+ $X2=3.555 $Y2=1.985
r110 27 42 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.015 $Y=0.84
+ $X2=3.015 $Y2=0.925
r111 27 29 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=3.015 $Y=0.84
+ $X2=3.015 $Y2=0.495
r112 26 38 15.363 $w=2.7e-07 $l=4.1845e-07 $layer=LI1_cond $X=1.305 $Y=1.805
+ $X2=1.13 $Y2=1.465
r113 25 31 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=3.385 $Y=1.805
+ $X2=3.555 $Y2=1.89
r114 25 26 135.701 $w=1.68e-07 $l=2.08e-06 $layer=LI1_cond $X=3.385 $Y=1.805
+ $X2=1.305 $Y2=1.805
r115 23 42 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.85 $Y=0.925
+ $X2=3.015 $Y2=0.925
r116 23 24 100.797 $w=1.68e-07 $l=1.545e-06 $layer=LI1_cond $X=2.85 $Y=0.925
+ $X2=1.305 $Y2=0.925
r117 22 38 9.12098 $w=2.7e-07 $l=2.05122e-07 $layer=LI1_cond $X=1.22 $Y=1.3
+ $X2=1.13 $Y2=1.465
r118 21 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.22 $Y=1.01
+ $X2=1.305 $Y2=0.925
r119 21 22 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.22 $Y=1.01
+ $X2=1.22 $Y2=1.3
r120 18 46 25.1816 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=1.025 $Y=1.765
+ $X2=1.025 $Y2=1.532
r121 18 20 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.025 $Y=1.765
+ $X2=1.025 $Y2=2.4
r122 14 45 25.1816 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=0.995 $Y=1.3
+ $X2=0.995 $Y2=1.532
r123 14 16 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.995 $Y=1.3
+ $X2=0.995 $Y2=0.74
r124 11 44 25.1816 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=0.575 $Y=1.765
+ $X2=0.575 $Y2=1.532
r125 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.575 $Y=1.765
+ $X2=0.575 $Y2=2.4
r126 7 43 25.1816 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=0.565 $Y=1.3
+ $X2=0.565 $Y2=1.532
r127 7 9 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.565 $Y=1.3
+ $X2=0.565 $Y2=0.74
r128 2 35 400 $w=1.7e-07 $l=9.29274e-07 $layer=licon1_PDIFF $count=1 $X=3.4
+ $Y=1.84 $X2=3.555 $Y2=2.695
r129 2 33 400 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=1 $X=3.4
+ $Y=1.84 $X2=3.555 $Y2=1.985
r130 1 42 182 $w=1.7e-07 $l=6.47321e-07 $layer=licon1_NDIFF $count=1 $X=2.815
+ $Y=0.37 $X2=3.015 $Y2=0.925
r131 1 29 182 $w=1.7e-07 $l=2.54951e-07 $layer=licon1_NDIFF $count=1 $X=2.815
+ $Y=0.37 $X2=3.015 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LS__A31O_2%A3 1 3 4 6 7
r31 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.69
+ $Y=1.385 $X2=1.69 $Y2=1.385
r32 7 11 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=1.69 $Y=1.295 $X2=1.69
+ $Y2=1.385
r33 4 10 38.9026 $w=2.7e-07 $l=2.05122e-07 $layer=POLY_cond $X=1.78 $Y=1.22
+ $X2=1.69 $Y2=1.385
r34 4 6 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.78 $Y=1.22 $X2=1.78
+ $Y2=0.74
r35 1 10 77.2841 $w=2.7e-07 $l=4.01871e-07 $layer=POLY_cond $X=1.735 $Y=1.765
+ $X2=1.69 $Y2=1.385
r36 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.735 $Y=1.765
+ $X2=1.735 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_LS__A31O_2%A2 1 3 4 6 7 11
c28 11 0 1.63365e-19 $X=2.26 $Y=1.385
c29 1 0 3.78493e-20 $X=2.17 $Y=1.22
r30 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.26
+ $Y=1.385 $X2=2.26 $Y2=1.385
r31 7 11 3.11471 $w=3.68e-07 $l=1e-07 $layer=LI1_cond $X=2.16 $Y=1.365 $X2=2.26
+ $Y2=1.365
r32 4 10 77.2841 $w=2.7e-07 $l=4.15812e-07 $layer=POLY_cond $X=2.185 $Y=1.765
+ $X2=2.26 $Y2=1.385
r33 4 6 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.185 $Y=1.765
+ $X2=2.185 $Y2=2.34
r34 1 10 38.9026 $w=2.7e-07 $l=2.05122e-07 $layer=POLY_cond $X=2.17 $Y=1.22
+ $X2=2.26 $Y2=1.385
r35 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.17 $Y=1.22 $X2=2.17
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__A31O_2%A1 1 3 4 6 7
c31 7 0 3.78493e-20 $X=3.12 $Y=1.295
c32 1 0 1.63365e-19 $X=2.74 $Y=1.22
r33 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.83
+ $Y=1.385 $X2=2.83 $Y2=1.385
r34 7 11 9.03266 $w=3.68e-07 $l=2.9e-07 $layer=LI1_cond $X=3.12 $Y=1.365
+ $X2=2.83 $Y2=1.365
r35 4 10 77.2841 $w=2.7e-07 $l=3.82492e-07 $layer=POLY_cond $X=2.825 $Y=1.765
+ $X2=2.83 $Y2=1.385
r36 4 6 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.825 $Y=1.765
+ $X2=2.825 $Y2=2.34
r37 1 10 38.9026 $w=2.7e-07 $l=2.05122e-07 $layer=POLY_cond $X=2.74 $Y=1.22
+ $X2=2.83 $Y2=1.385
r38 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.74 $Y=1.22 $X2=2.74
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__A31O_2%B1 1 3 4 6 7
r21 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.57
+ $Y=1.385 $X2=3.57 $Y2=1.385
r22 7 11 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=3.57 $Y=1.295 $X2=3.57
+ $Y2=1.385
r23 4 10 66.8857 $w=3.73e-07 $l=4.5299e-07 $layer=POLY_cond $X=3.325 $Y=1.765
+ $X2=3.485 $Y2=1.385
r24 4 6 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.325 $Y=1.765
+ $X2=3.325 $Y2=2.34
r25 1 10 39.1028 $w=3.73e-07 $l=2.43926e-07 $layer=POLY_cond $X=3.31 $Y=1.22
+ $X2=3.485 $Y2=1.385
r26 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.31 $Y=1.22 $X2=3.31
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__A31O_2%VPWR 1 2 3 10 12 18 24 26 28 33 40 41 47 50
r50 50 51 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r51 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r52 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r53 41 51 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=2.64 $Y2=3.33
r54 40 41 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r55 38 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.68 $Y=3.33
+ $X2=2.515 $Y2=3.33
r56 38 40 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.68 $Y=3.33 $X2=3.6
+ $Y2=3.33
r57 37 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r58 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r59 34 47 11.757 $w=1.7e-07 $l=2.68e-07 $layer=LI1_cond $X=1.625 $Y=3.33
+ $X2=1.357 $Y2=3.33
r60 34 36 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=1.625 $Y=3.33
+ $X2=2.16 $Y2=3.33
r61 33 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.35 $Y=3.33
+ $X2=2.515 $Y2=3.33
r62 33 36 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=2.35 $Y=3.33
+ $X2=2.16 $Y2=3.33
r63 32 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r64 32 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r65 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r66 29 44 3.93235 $w=1.7e-07 $l=2.18e-07 $layer=LI1_cond $X=0.435 $Y=3.33
+ $X2=0.217 $Y2=3.33
r67 29 31 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.435 $Y=3.33
+ $X2=0.72 $Y2=3.33
r68 28 47 11.757 $w=1.7e-07 $l=2.67e-07 $layer=LI1_cond $X=1.09 $Y=3.33
+ $X2=1.357 $Y2=3.33
r69 28 31 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.09 $Y=3.33 $X2=0.72
+ $Y2=3.33
r70 26 37 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.16 $Y2=3.33
r71 26 48 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.2 $Y2=3.33
r72 22 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.515 $Y=3.245
+ $X2=2.515 $Y2=3.33
r73 22 24 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=2.515 $Y=3.245
+ $X2=2.515 $Y2=2.565
r74 18 21 15.4261 $w=5.33e-07 $l=6.9e-07 $layer=LI1_cond $X=1.357 $Y=2.145
+ $X2=1.357 $Y2=2.835
r75 16 47 2.24534 $w=5.35e-07 $l=8.5e-08 $layer=LI1_cond $X=1.357 $Y=3.245
+ $X2=1.357 $Y2=3.33
r76 16 21 9.16621 $w=5.33e-07 $l=4.1e-07 $layer=LI1_cond $X=1.357 $Y=3.245
+ $X2=1.357 $Y2=2.835
r77 12 15 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=0.31 $Y=1.985
+ $X2=0.31 $Y2=2.815
r78 10 44 3.21082 $w=2.5e-07 $l=1.28662e-07 $layer=LI1_cond $X=0.31 $Y=3.245
+ $X2=0.217 $Y2=3.33
r79 10 15 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.31 $Y=3.245
+ $X2=0.31 $Y2=2.815
r80 3 24 600 $w=1.7e-07 $l=8.42912e-07 $layer=licon1_PDIFF $count=1 $X=2.26
+ $Y=1.84 $X2=2.515 $Y2=2.565
r81 2 21 400 $w=1.7e-07 $l=1.0697e-06 $layer=licon1_PDIFF $count=1 $X=1.1
+ $Y=1.84 $X2=1.255 $Y2=2.835
r82 2 18 400 $w=1.7e-07 $l=3.74566e-07 $layer=licon1_PDIFF $count=1 $X=1.1
+ $Y=1.84 $X2=1.255 $Y2=2.145
r83 1 15 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.205
+ $Y=1.84 $X2=0.35 $Y2=2.815
r84 1 12 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.205
+ $Y=1.84 $X2=0.35 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_LS__A31O_2%X 1 2 9 13 14 15 16 24 33
c30 33 0 3.54614e-20 $X=0.762 $Y=1.82
r31 21 24 0.292684 $w=3.13e-07 $l=8e-09 $layer=LI1_cond $X=0.762 $Y=1.977
+ $X2=0.762 $Y2=1.985
r32 15 16 13.5366 $w=3.13e-07 $l=3.7e-07 $layer=LI1_cond $X=0.762 $Y=2.405
+ $X2=0.762 $Y2=2.775
r33 14 21 0.512197 $w=3.13e-07 $l=1.4e-08 $layer=LI1_cond $X=0.762 $Y=1.963
+ $X2=0.762 $Y2=1.977
r34 14 33 7.65769 $w=3.13e-07 $l=1.43e-07 $layer=LI1_cond $X=0.762 $Y=1.963
+ $X2=0.762 $Y2=1.82
r35 14 15 13.061 $w=3.13e-07 $l=3.57e-07 $layer=LI1_cond $X=0.762 $Y=2.048
+ $X2=0.762 $Y2=2.405
r36 14 24 2.30489 $w=3.13e-07 $l=6.3e-08 $layer=LI1_cond $X=0.762 $Y=2.048
+ $X2=0.762 $Y2=1.985
r37 13 33 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=0.7 $Y=1.13 $X2=0.7
+ $Y2=1.82
r38 7 13 7.41084 $w=2.73e-07 $l=1.37e-07 $layer=LI1_cond $X=0.752 $Y=0.993
+ $X2=0.752 $Y2=1.13
r39 7 9 20.0316 $w=2.73e-07 $l=4.78e-07 $layer=LI1_cond $X=0.752 $Y=0.993
+ $X2=0.752 $Y2=0.515
r40 2 16 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=0.65
+ $Y=1.84 $X2=0.8 $Y2=2.815
r41 2 24 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=0.65
+ $Y=1.84 $X2=0.8 $Y2=1.985
r42 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.64
+ $Y=0.37 $X2=0.78 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__A31O_2%A_362_368# 1 2 9 14 16
r26 10 14 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.125 $Y=2.145
+ $X2=1.96 $Y2=2.145
r27 9 16 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.885 $Y=2.145
+ $X2=3.05 $Y2=2.145
r28 9 10 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=2.885 $Y=2.145
+ $X2=2.125 $Y2=2.145
r29 2 16 300 $w=1.7e-07 $l=3.97995e-07 $layer=licon1_PDIFF $count=2 $X=2.9
+ $Y=1.84 $X2=3.05 $Y2=2.17
r30 1 14 300 $w=1.7e-07 $l=3.87814e-07 $layer=licon1_PDIFF $count=2 $X=1.81
+ $Y=1.84 $X2=1.96 $Y2=2.16
.ends

.subckt PM_SKY130_FD_SC_LS__A31O_2%VGND 1 2 3 10 12 14 16 18 20 25 35 44
r44 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r45 36 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r46 35 40 9.19374 $w=6.68e-07 $l=5.15e-07 $layer=LI1_cond $X=1.395 $Y=0
+ $X2=1.395 $Y2=0.515
r47 35 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r48 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r49 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r50 29 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r51 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r52 26 35 9.03384 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=1.73 $Y=0 $X2=1.395
+ $Y2=0
r53 26 28 90.6845 $w=1.68e-07 $l=1.39e-06 $layer=LI1_cond $X=1.73 $Y=0 $X2=3.12
+ $Y2=0
r54 25 43 4.65971 $w=1.7e-07 $l=2.4e-07 $layer=LI1_cond $X=3.36 $Y=0 $X2=3.6
+ $Y2=0
r55 25 28 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=3.36 $Y=0 $X2=3.12
+ $Y2=0
r56 24 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r57 24 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r58 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r59 21 31 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.222
+ $Y2=0
r60 21 23 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.72
+ $Y2=0
r61 20 35 9.03384 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=1.06 $Y=0 $X2=1.395
+ $Y2=0
r62 20 23 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.06 $Y=0 $X2=0.72
+ $Y2=0
r63 18 29 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.92 $Y=0 $X2=3.12
+ $Y2=0
r64 18 38 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r65 14 43 3.10647 $w=3.3e-07 $l=1.16619e-07 $layer=LI1_cond $X=3.525 $Y=0.085
+ $X2=3.6 $Y2=0
r66 14 16 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.525 $Y=0.085
+ $X2=3.525 $Y2=0.515
r67 10 31 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.222 $Y2=0
r68 10 12 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.28 $Y2=0.515
r69 3 16 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.385
+ $Y=0.37 $X2=3.525 $Y2=0.515
r70 2 40 91 $w=1.7e-07 $l=5.6285e-07 $layer=licon1_NDIFF $count=2 $X=1.07
+ $Y=0.37 $X2=1.565 $Y2=0.515
r71 1 12 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

