* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__and4b_2 A_N B C D VGND VNB VPB VPWR X
X0 a_459_74# C a_537_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X1 VPWR B a_186_48# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_537_74# B a_645_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X3 VPWR D a_186_48# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 a_186_48# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 VGND a_186_48# X VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X6 X a_186_48# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X7 a_645_74# a_27_112# a_186_48# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X8 VPWR a_186_48# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X9 a_186_48# a_27_112# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_27_112# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X11 VGND D a_459_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X12 X a_186_48# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X13 a_27_112# A_N VGND VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
.ends
