* NGSPICE file created from sky130_fd_sc_ls__sdfxbp_2.ext - technology: sky130A

.subckt sky130_fd_sc_ls__sdfxbp_2 CLK D SCD SCE VGND VNB VPB VPWR Q Q_N
M1000 a_630_74# CLK VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=2.2043e+12p ps=1.954e+07u
M1001 a_630_74# CLK VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=5.656e+11p pd=3.25e+06u as=3.1895e+12p ps=2.586e+07u
M1002 VPWR a_2322_368# Q_N VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.36e+11p ps=2.84e+06u
M1003 a_301_74# D a_238_453# VPB phighvt w=640000u l=150000u
+  ad=3.511e+11p pd=3.42e+06u as=1.728e+11p ps=1.82e+06u
M1004 VPWR a_1243_48# a_1217_499# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1005 VPWR a_1711_48# a_2322_368# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.85e+11p ps=2.57e+06u
M1006 a_423_453# a_36_74# a_301_74# VPB phighvt w=640000u l=150000u
+  ad=2.144e+11p pd=1.95e+06u as=0p ps=0u
M1007 a_1711_48# a_1511_74# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.85e+11p pd=2.57e+06u as=0p ps=0u
M1008 a_1663_74# a_630_74# a_1511_74# VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=2.887e+11p ps=2.32e+06u
M1009 VGND a_1711_48# a_1663_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 Q a_1711_48# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=0p ps=0u
M1011 a_828_74# a_630_74# VGND VNB nshort w=740000u l=150000u
+  ad=1.998e+11p pd=2.02e+06u as=0p ps=0u
M1012 a_223_74# a_36_74# VGND VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1013 a_301_74# D a_223_74# VNB nshort w=420000u l=150000u
+  ad=3.654e+11p pd=3.42e+06u as=0p ps=0u
M1014 VGND a_1243_48# a_1173_97# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.6425e+11p ps=1.77e+06u
M1015 a_1217_499# a_630_74# a_1021_97# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.617e+11p ps=1.61e+06u
M1016 a_1511_74# a_630_74# a_1243_48# VPB phighvt w=840000u l=150000u
+  ad=2.856e+11p pd=2.45e+06u as=5.418e+11p ps=2.97e+06u
M1017 a_1021_97# a_630_74# a_301_74# VNB nshort w=420000u l=150000u
+  ad=2.562e+11p pd=2.06e+06u as=0p ps=0u
M1018 a_1243_48# a_1021_97# VGND VNB nshort w=550000u l=150000u
+  ad=1.54e+11p pd=1.66e+06u as=0p ps=0u
M1019 Q_N a_2322_368# VGND VNB nshort w=740000u l=150000u
+  ad=2.183e+11p pd=2.07e+06u as=0p ps=0u
M1020 VPWR a_1711_48# Q VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND a_1711_48# a_2322_368# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1022 Q a_1711_48# VGND VNB nshort w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1023 VPWR SCE a_36_74# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=2.432e+11p ps=2.04e+06u
M1024 VGND SCD a_450_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1025 a_1711_48# a_1511_74# VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1026 a_450_74# SCE a_301_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VPWR SCD a_423_453# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_1173_97# a_828_74# a_1021_97# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPWR a_1711_48# a_1691_508# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1030 a_238_453# SCE VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_828_74# a_630_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=0p ps=0u
M1032 VGND SCE a_36_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1033 a_1511_74# a_828_74# a_1243_48# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 Q_N a_2322_368# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_1021_97# a_828_74# a_301_74# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_1691_508# a_828_74# a_1511_74# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 VGND a_1711_48# Q VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 a_1243_48# a_1021_97# VPWR VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 VGND a_2322_368# Q_N VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

