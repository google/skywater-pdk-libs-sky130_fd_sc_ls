* File: sky130_fd_sc_ls__o32ai_1.pex.spice
* Created: Wed Sep  2 11:23:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__O32AI_1%B1 1 3 4 6 7
r23 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.28
+ $Y=1.385 $X2=0.28 $Y2=1.385
r24 7 11 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.28 $Y=1.295 $X2=0.28
+ $Y2=1.385
r25 4 10 67.1244 $w=3.69e-07 $l=4.61302e-07 $layer=POLY_cond $X=0.565 $Y=1.765
+ $X2=0.385 $Y2=1.385
r26 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.565 $Y=1.765
+ $X2=0.565 $Y2=2.4
r27 1 10 39.0404 $w=3.69e-07 $l=2.13014e-07 $layer=POLY_cond $X=0.495 $Y=1.22
+ $X2=0.385 $Y2=1.385
r28 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.495 $Y=1.22 $X2=0.495
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__O32AI_1%B2 1 3 6 8 12
r27 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.14
+ $Y=1.515 $X2=1.14 $Y2=1.515
r28 8 12 5.08431 $w=3.38e-07 $l=1.5e-07 $layer=LI1_cond $X=1.145 $Y=1.665
+ $X2=1.145 $Y2=1.515
r29 4 11 38.9379 $w=3.62e-07 $l=2.20624e-07 $layer=POLY_cond $X=1.23 $Y=1.35
+ $X2=1.1 $Y2=1.515
r30 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.23 $Y=1.35 $X2=1.23
+ $Y2=0.74
r31 1 11 50.2556 $w=3.62e-07 $l=3.02076e-07 $layer=POLY_cond $X=0.985 $Y=1.765
+ $X2=1.1 $Y2=1.515
r32 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.985 $Y=1.765
+ $X2=0.985 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__O32AI_1%A3 1 3 6 8 9 10 16
r32 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.71
+ $Y=1.515 $X2=1.71 $Y2=1.515
r33 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.71 $Y=2.035
+ $X2=1.71 $Y2=2.405
r34 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.71 $Y=1.665 $X2=1.71
+ $Y2=2.035
r35 8 16 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.71 $Y=1.665
+ $X2=1.71 $Y2=1.515
r36 4 15 38.5562 $w=2.99e-07 $l=1.74714e-07 $layer=POLY_cond $X=1.73 $Y=1.35
+ $X2=1.71 $Y2=1.515
r37 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.73 $Y=1.35 $X2=1.73
+ $Y2=0.74
r38 1 15 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=1.635 $Y=1.765
+ $X2=1.71 $Y2=1.515
r39 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.635 $Y=1.765
+ $X2=1.635 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__O32AI_1%A2 1 3 6 8 9 10 11 18
r33 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.28
+ $Y=1.515 $X2=2.28 $Y2=1.515
r34 10 11 10.6601 $w=3.98e-07 $l=3.7e-07 $layer=LI1_cond $X=2.245 $Y=2.405
+ $X2=2.245 $Y2=2.775
r35 9 10 10.6601 $w=3.98e-07 $l=3.7e-07 $layer=LI1_cond $X=2.245 $Y=2.035
+ $X2=2.245 $Y2=2.405
r36 8 9 10.6601 $w=3.98e-07 $l=3.7e-07 $layer=LI1_cond $X=2.245 $Y=1.665
+ $X2=2.245 $Y2=2.035
r37 8 18 4.32166 $w=3.98e-07 $l=1.5e-07 $layer=LI1_cond $X=2.245 $Y=1.665
+ $X2=2.245 $Y2=1.515
r38 4 17 38.5562 $w=2.99e-07 $l=1.88348e-07 $layer=POLY_cond $X=2.33 $Y=1.35
+ $X2=2.28 $Y2=1.515
r39 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.33 $Y=1.35 $X2=2.33
+ $Y2=0.74
r40 1 17 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=2.205 $Y=1.765
+ $X2=2.28 $Y2=1.515
r41 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.205 $Y=1.765
+ $X2=2.205 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__O32AI_1%A1 1 3 4 6 7
r21 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.045
+ $Y=1.385 $X2=3.045 $Y2=1.385
r22 7 11 2.92169 $w=3.53e-07 $l=9e-08 $layer=LI1_cond $X=3.057 $Y=1.295
+ $X2=3.057 $Y2=1.385
r23 4 10 66.0675 $w=3.88e-07 $l=4.57996e-07 $layer=POLY_cond $X=2.775 $Y=1.765
+ $X2=2.947 $Y2=1.385
r24 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.775 $Y=1.765
+ $X2=2.775 $Y2=2.4
r25 1 10 39.3587 $w=3.88e-07 $l=2.56562e-07 $layer=POLY_cond $X=2.76 $Y=1.22
+ $X2=2.947 $Y2=1.385
r26 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.76 $Y=1.22 $X2=2.76
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__O32AI_1%VPWR 1 2 7 9 13 15 19 21 34
r29 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r30 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r31 28 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r32 27 28 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r33 25 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r34 24 27 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.72 $Y=3.33
+ $X2=2.64 $Y2=3.33
r35 24 25 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r36 22 30 4.68787 $w=1.7e-07 $l=2.33e-07 $layer=LI1_cond $X=0.465 $Y=3.33
+ $X2=0.232 $Y2=3.33
r37 22 24 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.465 $Y=3.33
+ $X2=0.72 $Y2=3.33
r38 21 33 4.58274 $w=1.7e-07 $l=2.62e-07 $layer=LI1_cond $X=2.835 $Y=3.33
+ $X2=3.097 $Y2=3.33
r39 21 27 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=2.835 $Y=3.33
+ $X2=2.64 $Y2=3.33
r40 19 28 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r41 19 25 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r42 15 18 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=3 $Y=1.985 $X2=3
+ $Y2=2.815
r43 13 33 3.18343 $w=3.3e-07 $l=1.32868e-07 $layer=LI1_cond $X=3 $Y=3.245
+ $X2=3.097 $Y2=3.33
r44 13 18 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3 $Y=3.245 $X2=3
+ $Y2=2.815
r45 9 12 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=0.3 $Y=1.985 $X2=0.3
+ $Y2=2.815
r46 7 30 3.0783 $w=3.3e-07 $l=1.14039e-07 $layer=LI1_cond $X=0.3 $Y=3.245
+ $X2=0.232 $Y2=3.33
r47 7 12 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.3 $Y=3.245 $X2=0.3
+ $Y2=2.815
r48 2 18 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.85
+ $Y=1.84 $X2=3 $Y2=2.815
r49 2 15 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.85
+ $Y=1.84 $X2=3 $Y2=1.985
r50 1 12 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.155
+ $Y=1.84 $X2=0.3 $Y2=2.815
r51 1 9 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.155
+ $Y=1.84 $X2=0.3 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_LS__O32AI_1%Y 1 2 12 14 17 18
r29 17 18 11.0599 $w=7.38e-07 $l=1.65e-07 $layer=LI1_cond $X=1.005 $Y=2.115
+ $X2=1.005 $Y2=1.95
r30 14 17 10.6677 $w=7.38e-07 $l=6.6e-07 $layer=LI1_cond $X=1.005 $Y=2.775
+ $X2=1.005 $Y2=2.115
r31 9 12 4.91896 $w=4.08e-07 $l=1.75e-07 $layer=LI1_cond $X=0.72 $Y=0.925
+ $X2=0.895 $Y2=0.925
r32 7 9 5.92876 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=0.72 $Y=1.13 $X2=0.72
+ $Y2=0.925
r33 7 18 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=0.72 $Y=1.13 $X2=0.72
+ $Y2=1.95
r34 2 14 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.06
+ $Y=1.84 $X2=1.21 $Y2=2.815
r35 2 17 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=1.06
+ $Y=1.84 $X2=1.21 $Y2=2.115
r36 1 12 182 $w=1.7e-07 $l=6.83447e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.895 $Y2=0.91
.ends

.subckt PM_SKY130_FD_SC_LS__O32AI_1%A_27_74# 1 2 3 12 14 15 16 17 20 23
r45 18 20 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=2.545 $Y=1.01
+ $X2=2.545 $Y2=0.515
r46 16 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.38 $Y=1.095
+ $X2=2.545 $Y2=1.01
r47 16 17 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=2.38 $Y=1.095 $X2=1.68
+ $Y2=1.095
r48 15 17 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.515 $Y=1.01
+ $X2=1.68 $Y2=1.095
r49 14 25 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.515 $Y=0.52
+ $X2=1.515 $Y2=0.435
r50 14 15 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=1.515 $Y=0.52
+ $X2=1.515 $Y2=1.01
r51 13 23 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.445 $Y=0.435
+ $X2=0.28 $Y2=0.435
r52 12 25 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.35 $Y=0.435
+ $X2=1.515 $Y2=0.435
r53 12 13 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=1.35 $Y=0.435
+ $X2=0.445 $Y2=0.435
r54 3 20 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.405
+ $Y=0.37 $X2=2.545 $Y2=0.515
r55 2 25 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=1.305
+ $Y=0.37 $X2=1.515 $Y2=0.515
r56 1 23 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__O32AI_1%VGND 1 2 9 11 13 16 17 18 27 33
r35 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r36 30 33 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r37 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r38 27 32 3.97916 $w=1.7e-07 $l=2.4e-07 $layer=LI1_cond $X=2.88 $Y=0 $X2=3.12
+ $Y2=0
r39 27 29 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=2.88 $Y=0 $X2=2.64
+ $Y2=0
r40 21 25 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=1.68
+ $Y2=0
r41 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r42 18 30 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r43 18 22 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.24
+ $Y2=0
r44 18 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r45 16 25 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.85 $Y=0 $X2=1.68
+ $Y2=0
r46 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.85 $Y=0 $X2=2.015
+ $Y2=0
r47 15 29 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=2.18 $Y=0 $X2=2.64
+ $Y2=0
r48 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.18 $Y=0 $X2=2.015
+ $Y2=0
r49 11 32 3.23306 $w=2.6e-07 $l=1.46458e-07 $layer=LI1_cond $X=3.01 $Y=0.085
+ $X2=3.12 $Y2=0
r50 11 13 18.6164 $w=2.58e-07 $l=4.2e-07 $layer=LI1_cond $X=3.01 $Y=0.085
+ $X2=3.01 $Y2=0.505
r51 7 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.015 $Y=0.085
+ $X2=2.015 $Y2=0
r52 7 9 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=2.015 $Y=0.085
+ $X2=2.015 $Y2=0.645
r53 2 13 91 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=2 $X=2.835
+ $Y=0.37 $X2=2.975 $Y2=0.505
r54 1 9 182 $w=1.7e-07 $l=3.65205e-07 $layer=licon1_NDIFF $count=1 $X=1.805
+ $Y=0.37 $X2=2.015 $Y2=0.645
.ends

