* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__o41ai_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
M1000 a_132_74# A4 VGND VNB nshort w=740000u l=150000u
+  ad=1.4245e+12p pd=1.273e+07u as=1.0397e+12p ps=8.73e+06u
M1001 VGND A4 a_132_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_607_368# A2 a_807_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=6.72e+11p pd=5.68e+06u as=9.744e+11p ps=8.46e+06u
M1003 a_132_74# B1 Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.072e+11p ps=2.04e+06u
M1004 VGND A3 a_132_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_132_74# A3 VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_607_368# A3 a_314_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=1.1144e+12p ps=8.71e+06u
M1007 a_132_74# A2 VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_132_74# A1 VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_807_368# A2 a_607_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR A1 a_807_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=9.688e+11p pd=8.45e+06u as=0p ps=0u
M1011 Y A4 a_314_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=6.72e+11p pd=5.68e+06u as=0p ps=0u
M1012 a_314_368# A3 a_607_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND A1 a_132_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_807_368# A1 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y B1 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR B1 Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_314_368# A4 Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND A2 a_132_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 Y B1 a_132_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
