* File: sky130_fd_sc_ls__a311oi_2.pxi.spice
* Created: Wed Sep  2 10:51:55 2020
* 
x_PM_SKY130_FD_SC_LS__A311OI_2%A3 N_A3_c_93_n N_A3_M1007_g N_A3_c_89_n
+ N_A3_M1004_g N_A3_c_90_n N_A3_M1005_g N_A3_c_94_n N_A3_M1008_g A3 N_A3_c_92_n
+ PM_SKY130_FD_SC_LS__A311OI_2%A3
x_PM_SKY130_FD_SC_LS__A311OI_2%A2 N_A2_c_130_n N_A2_M1002_g N_A2_c_135_n
+ N_A2_M1010_g N_A2_c_131_n N_A2_M1012_g N_A2_c_136_n N_A2_M1016_g N_A2_c_132_n
+ A2 N_A2_c_133_n N_A2_c_134_n PM_SKY130_FD_SC_LS__A311OI_2%A2
x_PM_SKY130_FD_SC_LS__A311OI_2%A1 N_A1_c_190_n N_A1_M1009_g N_A1_c_191_n
+ N_A1_M1011_g N_A1_M1006_g N_A1_M1015_g N_A1_c_188_n A1 N_A1_c_189_n
+ PM_SKY130_FD_SC_LS__A311OI_2%A1
x_PM_SKY130_FD_SC_LS__A311OI_2%B1 N_B1_M1014_g N_B1_c_240_n N_B1_M1000_g
+ N_B1_c_241_n N_B1_M1013_g B1 B1 B1 N_B1_c_239_n
+ PM_SKY130_FD_SC_LS__A311OI_2%B1
x_PM_SKY130_FD_SC_LS__A311OI_2%C1 N_C1_M1017_g N_C1_c_288_n N_C1_M1001_g
+ N_C1_c_289_n N_C1_M1003_g C1 N_C1_c_286_n N_C1_c_287_n
+ PM_SKY130_FD_SC_LS__A311OI_2%C1
x_PM_SKY130_FD_SC_LS__A311OI_2%VPWR N_VPWR_M1007_s N_VPWR_M1008_s N_VPWR_M1016_s
+ N_VPWR_M1011_s N_VPWR_c_328_n N_VPWR_c_329_n N_VPWR_c_330_n N_VPWR_c_331_n
+ N_VPWR_c_332_n N_VPWR_c_333_n VPWR N_VPWR_c_334_n N_VPWR_c_335_n
+ N_VPWR_c_336_n N_VPWR_c_327_n N_VPWR_c_338_n N_VPWR_c_339_n N_VPWR_c_340_n
+ PM_SKY130_FD_SC_LS__A311OI_2%VPWR
x_PM_SKY130_FD_SC_LS__A311OI_2%A_127_368# N_A_127_368#_M1007_d
+ N_A_127_368#_M1010_d N_A_127_368#_M1009_d N_A_127_368#_M1000_s
+ N_A_127_368#_c_399_n N_A_127_368#_c_400_n N_A_127_368#_c_401_n
+ N_A_127_368#_c_402_n N_A_127_368#_c_403_n N_A_127_368#_c_404_n
+ N_A_127_368#_c_405_n N_A_127_368#_c_406_n N_A_127_368#_c_407_n
+ N_A_127_368#_c_443_n PM_SKY130_FD_SC_LS__A311OI_2%A_127_368#
x_PM_SKY130_FD_SC_LS__A311OI_2%A_692_368# N_A_692_368#_M1000_d
+ N_A_692_368#_M1013_d N_A_692_368#_M1003_s N_A_692_368#_c_471_n
+ N_A_692_368#_c_472_n N_A_692_368#_c_473_n N_A_692_368#_c_484_n
+ N_A_692_368#_c_474_n N_A_692_368#_c_475_n N_A_692_368#_c_476_n
+ PM_SKY130_FD_SC_LS__A311OI_2%A_692_368#
x_PM_SKY130_FD_SC_LS__A311OI_2%Y N_Y_M1006_d N_Y_M1015_d N_Y_M1017_d N_Y_M1001_d
+ N_Y_c_518_n N_Y_c_519_n N_Y_c_524_n N_Y_c_520_n N_Y_c_542_n Y Y Y N_Y_c_523_n
+ PM_SKY130_FD_SC_LS__A311OI_2%Y
x_PM_SKY130_FD_SC_LS__A311OI_2%A_45_74# N_A_45_74#_M1004_s N_A_45_74#_M1005_s
+ N_A_45_74#_M1012_d N_A_45_74#_c_576_n N_A_45_74#_c_581_n N_A_45_74#_c_577_n
+ N_A_45_74#_c_578_n N_A_45_74#_c_587_n N_A_45_74#_c_579_n N_A_45_74#_c_591_n
+ PM_SKY130_FD_SC_LS__A311OI_2%A_45_74#
x_PM_SKY130_FD_SC_LS__A311OI_2%VGND N_VGND_M1004_d N_VGND_M1014_d N_VGND_c_611_n
+ N_VGND_c_612_n VGND N_VGND_c_613_n N_VGND_c_614_n N_VGND_c_615_n
+ N_VGND_c_616_n N_VGND_c_617_n N_VGND_c_618_n PM_SKY130_FD_SC_LS__A311OI_2%VGND
x_PM_SKY130_FD_SC_LS__A311OI_2%A_300_74# N_A_300_74#_M1002_s N_A_300_74#_M1006_s
+ N_A_300_74#_c_661_n N_A_300_74#_c_662_n PM_SKY130_FD_SC_LS__A311OI_2%A_300_74#
cc_1 VNB N_A3_c_89_n 0.022852f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.22
cc_2 VNB N_A3_c_90_n 0.0168728f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.22
cc_3 VNB A3 0.0155644f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_4 VNB N_A3_c_92_n 0.059158f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.492
cc_5 VNB N_A2_c_130_n 0.0174681f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=1.765
cc_6 VNB N_A2_c_131_n 0.022624f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.22
cc_7 VNB N_A2_c_132_n 0.00595132f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.385
cc_8 VNB N_A2_c_133_n 0.0586322f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A2_c_134_n 0.00814841f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A1_M1006_g 0.0285804f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_11 VNB N_A1_M1015_g 0.0236097f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_12 VNB N_A1_c_188_n 0.003533f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=1.492
cc_13 VNB N_A1_c_189_n 0.0806997f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_B1_M1014_g 0.0281458f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=2.4
cc_15 VNB B1 0.00612637f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_16 VNB N_B1_c_239_n 0.0429774f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.492
cc_17 VNB N_C1_M1017_g 0.0346834f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=2.4
cc_18 VNB N_C1_c_286_n 0.0486353f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.492
cc_19 VNB N_C1_c_287_n 0.00305603f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.492
cc_20 VNB N_VPWR_c_327_n 0.243291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_Y_c_518_n 0.0126151f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_22 VNB N_Y_c_519_n 0.00206055f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.385
cc_23 VNB N_Y_c_520_n 0.00198283f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB Y 0.0734368f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB Y 0.0265258f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_Y_c_523_n 0.00555748f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_45_74#_c_576_n 0.0207156f $X=-0.19 $Y=-0.245 $X2=1.01 $Y2=2.4
cc_28 VNB N_A_45_74#_c_577_n 0.0102706f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=1.492
cc_29 VNB N_A_45_74#_c_578_n 0.00216743f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.385
cc_30 VNB N_A_45_74#_c_579_n 0.00469816f $X=-0.19 $Y=-0.245 $X2=0.652 $Y2=1.385
cc_31 VNB N_VGND_c_611_n 0.00396467f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_32 VNB N_VGND_c_612_n 0.0127126f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_33 VNB N_VGND_c_613_n 0.0196185f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.492
cc_34 VNB N_VGND_c_614_n 0.0766417f $X=-0.19 $Y=-0.245 $X2=0.652 $Y2=1.295
cc_35 VNB N_VGND_c_615_n 0.0343549f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_616_n 0.323383f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_617_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_618_n 0.0115409f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_300_74#_c_661_n 0.002374f $X=-0.19 $Y=-0.245 $X2=1.01 $Y2=2.4
cc_40 VNB N_A_300_74#_c_662_n 0.0263182f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_41 VPB N_A3_c_93_n 0.0174349f $X=-0.19 $Y=1.66 $X2=0.56 $Y2=1.765
cc_42 VPB N_A3_c_94_n 0.0151654f $X=-0.19 $Y=1.66 $X2=1.01 $Y2=1.765
cc_43 VPB N_A3_c_92_n 0.0160648f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=1.492
cc_44 VPB N_A2_c_135_n 0.0151654f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=1.22
cc_45 VPB N_A2_c_136_n 0.0153802f $X=-0.19 $Y=1.66 $X2=1.01 $Y2=1.765
cc_46 VPB N_A2_c_133_n 0.0124937f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB N_A1_c_190_n 0.0146815f $X=-0.19 $Y=1.66 $X2=0.56 $Y2=1.765
cc_48 VPB N_A1_c_191_n 0.0187985f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=1.22
cc_49 VPB N_A1_c_188_n 0.00394407f $X=-0.19 $Y=1.66 $X2=0.56 $Y2=1.492
cc_50 VPB N_A1_c_189_n 0.0282956f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_51 VPB N_B1_c_240_n 0.018461f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=0.74
cc_52 VPB N_B1_c_241_n 0.0147854f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=0.74
cc_53 VPB B1 0.010884f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_54 VPB N_B1_c_239_n 0.0215624f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=1.492
cc_55 VPB N_C1_c_288_n 0.0148335f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=0.74
cc_56 VPB N_C1_c_289_n 0.0170355f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=0.74
cc_57 VPB N_C1_c_286_n 0.0233284f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=1.492
cc_58 VPB N_C1_c_287_n 0.00276432f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.492
cc_59 VPB N_VPWR_c_328_n 0.0124065f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_60 VPB N_VPWR_c_329_n 0.0654039f $X=-0.19 $Y=1.66 $X2=0.56 $Y2=1.492
cc_61 VPB N_VPWR_c_330_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.385
cc_62 VPB N_VPWR_c_331_n 0.00799266f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_332_n 0.00537498f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_333_n 0.0121236f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_334_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_335_n 0.0164465f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_336_n 0.0619548f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_327_n 0.0922127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_338_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_339_n 0.00517953f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_340_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_A_127_368#_c_399_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0.56 $Y2=1.492
cc_73 VPB N_A_127_368#_c_400_n 0.00242893f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.385
cc_74 VPB N_A_127_368#_c_401_n 0.00490377f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=1.492
cc_75 VPB N_A_127_368#_c_402_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_A_127_368#_c_403_n 0.00573492f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_A_127_368#_c_404_n 0.00180921f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_A_127_368#_c_405_n 0.0125008f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 VPB N_A_127_368#_c_406_n 0.00224287f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 VPB N_A_127_368#_c_407_n 0.00215641f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_A_692_368#_c_471_n 0.00587339f $X=-0.19 $Y=1.66 $X2=1.01 $Y2=2.4
cc_82 VPB N_A_692_368#_c_472_n 0.00213603f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 VPB N_A_692_368#_c_473_n 0.00424137f $X=-0.19 $Y=1.66 $X2=0.56 $Y2=1.492
cc_84 VPB N_A_692_368#_c_474_n 0.0120084f $X=-0.19 $Y=1.66 $X2=0.652 $Y2=1.295
cc_85 VPB N_A_692_368#_c_475_n 0.0241341f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_A_692_368#_c_476_n 0.0021839f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_Y_c_524_n 0.011537f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB Y 0.01369f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 N_A3_c_90_n N_A2_c_130_n 0.0103348f $X=0.995 $Y=1.22 $X2=-0.19 $Y2=-0.245
cc_90 N_A3_c_94_n N_A2_c_135_n 0.0208942f $X=1.01 $Y=1.765 $X2=0 $Y2=0
cc_91 A3 N_A2_c_133_n 2.0669e-19 $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_92 N_A3_c_92_n N_A2_c_133_n 0.0289262f $X=0.995 $Y=1.492 $X2=0 $Y2=0
cc_93 N_A3_c_90_n N_A2_c_134_n 0.00444493f $X=0.995 $Y=1.22 $X2=0 $Y2=0
cc_94 A3 N_A2_c_134_n 0.0233695f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_95 N_A3_c_92_n N_A2_c_134_n 3.87575e-19 $X=0.995 $Y=1.492 $X2=0 $Y2=0
cc_96 N_A3_c_93_n N_VPWR_c_329_n 0.0100905f $X=0.56 $Y=1.765 $X2=0 $Y2=0
cc_97 N_A3_c_93_n N_VPWR_c_330_n 0.00445602f $X=0.56 $Y=1.765 $X2=0 $Y2=0
cc_98 N_A3_c_94_n N_VPWR_c_330_n 0.00445602f $X=1.01 $Y=1.765 $X2=0 $Y2=0
cc_99 N_A3_c_94_n N_VPWR_c_331_n 0.00646778f $X=1.01 $Y=1.765 $X2=0 $Y2=0
cc_100 N_A3_c_93_n N_VPWR_c_327_n 0.00861252f $X=0.56 $Y=1.765 $X2=0 $Y2=0
cc_101 N_A3_c_94_n N_VPWR_c_327_n 0.00857673f $X=1.01 $Y=1.765 $X2=0 $Y2=0
cc_102 N_A3_c_93_n N_A_127_368#_c_399_n 0.0127167f $X=0.56 $Y=1.765 $X2=0 $Y2=0
cc_103 N_A3_c_94_n N_A_127_368#_c_399_n 0.0133148f $X=1.01 $Y=1.765 $X2=0 $Y2=0
cc_104 N_A3_c_94_n N_A_127_368#_c_400_n 0.00899835f $X=1.01 $Y=1.765 $X2=0 $Y2=0
cc_105 N_A3_c_92_n N_A_127_368#_c_400_n 0.00735489f $X=0.995 $Y=1.492 $X2=0
+ $Y2=0
cc_106 N_A3_c_93_n N_A_127_368#_c_401_n 0.00418463f $X=0.56 $Y=1.765 $X2=0 $Y2=0
cc_107 N_A3_c_94_n N_A_127_368#_c_401_n 0.00109449f $X=1.01 $Y=1.765 $X2=0 $Y2=0
cc_108 A3 N_A_127_368#_c_401_n 0.0182301f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_109 N_A3_c_92_n N_A_127_368#_c_401_n 0.00678516f $X=0.995 $Y=1.492 $X2=0
+ $Y2=0
cc_110 N_A3_c_94_n N_A_127_368#_c_402_n 7.15508e-19 $X=1.01 $Y=1.765 $X2=0 $Y2=0
cc_111 N_A3_c_89_n N_A_45_74#_c_576_n 4.43891e-19 $X=0.565 $Y=1.22 $X2=0 $Y2=0
cc_112 N_A3_c_89_n N_A_45_74#_c_581_n 0.00979433f $X=0.565 $Y=1.22 $X2=0 $Y2=0
cc_113 N_A3_c_90_n N_A_45_74#_c_581_n 0.014168f $X=0.995 $Y=1.22 $X2=0 $Y2=0
cc_114 A3 N_A_45_74#_c_581_n 0.0234443f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_115 N_A3_c_92_n N_A_45_74#_c_581_n 6.29572e-19 $X=0.995 $Y=1.492 $X2=0 $Y2=0
cc_116 N_A3_c_90_n N_A_45_74#_c_578_n 2.82517e-19 $X=0.995 $Y=1.22 $X2=0 $Y2=0
cc_117 N_A3_c_89_n N_VGND_c_611_n 0.010528f $X=0.565 $Y=1.22 $X2=0 $Y2=0
cc_118 N_A3_c_90_n N_VGND_c_611_n 0.00755236f $X=0.995 $Y=1.22 $X2=0 $Y2=0
cc_119 N_A3_c_89_n N_VGND_c_613_n 0.00383152f $X=0.565 $Y=1.22 $X2=0 $Y2=0
cc_120 N_A3_c_90_n N_VGND_c_614_n 0.00383152f $X=0.995 $Y=1.22 $X2=0 $Y2=0
cc_121 N_A3_c_89_n N_VGND_c_616_n 0.00387841f $X=0.565 $Y=1.22 $X2=0 $Y2=0
cc_122 N_A3_c_90_n N_VGND_c_616_n 0.00384065f $X=0.995 $Y=1.22 $X2=0 $Y2=0
cc_123 N_A2_c_136_n N_A1_c_190_n 0.0198677f $X=1.91 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_124 N_A2_c_132_n N_A1_c_188_n 0.0139406f $X=1.925 $Y=1.385 $X2=0 $Y2=0
cc_125 N_A2_c_133_n N_A1_c_188_n 2.46355e-19 $X=1.91 $Y=1.492 $X2=0 $Y2=0
cc_126 N_A2_c_132_n N_A1_c_189_n 6.33995e-19 $X=1.925 $Y=1.385 $X2=0 $Y2=0
cc_127 N_A2_c_133_n N_A1_c_189_n 0.0273979f $X=1.91 $Y=1.492 $X2=0 $Y2=0
cc_128 N_A2_c_135_n N_VPWR_c_331_n 0.00646778f $X=1.46 $Y=1.765 $X2=0 $Y2=0
cc_129 N_A2_c_136_n N_VPWR_c_332_n 0.00719936f $X=1.91 $Y=1.765 $X2=0 $Y2=0
cc_130 N_A2_c_135_n N_VPWR_c_334_n 0.00445602f $X=1.46 $Y=1.765 $X2=0 $Y2=0
cc_131 N_A2_c_136_n N_VPWR_c_334_n 0.00445602f $X=1.91 $Y=1.765 $X2=0 $Y2=0
cc_132 N_A2_c_135_n N_VPWR_c_327_n 0.00857673f $X=1.46 $Y=1.765 $X2=0 $Y2=0
cc_133 N_A2_c_136_n N_VPWR_c_327_n 0.00857936f $X=1.91 $Y=1.765 $X2=0 $Y2=0
cc_134 N_A2_c_135_n N_A_127_368#_c_399_n 7.15508e-19 $X=1.46 $Y=1.765 $X2=0
+ $Y2=0
cc_135 N_A2_c_135_n N_A_127_368#_c_400_n 0.00899835f $X=1.46 $Y=1.765 $X2=0
+ $Y2=0
cc_136 N_A2_c_133_n N_A_127_368#_c_400_n 0.00349848f $X=1.91 $Y=1.492 $X2=0
+ $Y2=0
cc_137 N_A2_c_134_n N_A_127_368#_c_400_n 0.0333429f $X=1.315 $Y=1.365 $X2=0
+ $Y2=0
cc_138 N_A2_c_135_n N_A_127_368#_c_402_n 0.0133148f $X=1.46 $Y=1.765 $X2=0 $Y2=0
cc_139 N_A2_c_136_n N_A_127_368#_c_402_n 0.0134918f $X=1.91 $Y=1.765 $X2=0 $Y2=0
cc_140 N_A2_c_136_n N_A_127_368#_c_403_n 0.00911718f $X=1.91 $Y=1.765 $X2=0
+ $Y2=0
cc_141 N_A2_c_132_n N_A_127_368#_c_403_n 0.0174421f $X=1.925 $Y=1.385 $X2=0
+ $Y2=0
cc_142 N_A2_c_133_n N_A_127_368#_c_403_n 0.00547177f $X=1.91 $Y=1.492 $X2=0
+ $Y2=0
cc_143 N_A2_c_135_n N_A_127_368#_c_406_n 0.00109449f $X=1.46 $Y=1.765 $X2=0
+ $Y2=0
cc_144 N_A2_c_136_n N_A_127_368#_c_406_n 0.00109449f $X=1.91 $Y=1.765 $X2=0
+ $Y2=0
cc_145 N_A2_c_132_n N_A_127_368#_c_406_n 0.0275631f $X=1.925 $Y=1.385 $X2=0
+ $Y2=0
cc_146 N_A2_c_133_n N_A_127_368#_c_406_n 0.00517401f $X=1.91 $Y=1.492 $X2=0
+ $Y2=0
cc_147 N_A2_c_131_n N_Y_c_518_n 0.00316716f $X=1.855 $Y=1.22 $X2=0 $Y2=0
cc_148 N_A2_c_130_n N_A_45_74#_c_578_n 6.33564e-19 $X=1.425 $Y=1.22 $X2=0 $Y2=0
cc_149 N_A2_c_134_n N_A_45_74#_c_587_n 0.014682f $X=1.315 $Y=1.365 $X2=0 $Y2=0
cc_150 N_A2_c_131_n N_A_45_74#_c_579_n 0.00192588f $X=1.855 $Y=1.22 $X2=0 $Y2=0
cc_151 N_A2_c_132_n N_A_45_74#_c_579_n 0.0118504f $X=1.925 $Y=1.385 $X2=0 $Y2=0
cc_152 N_A2_c_133_n N_A_45_74#_c_579_n 0.00374323f $X=1.91 $Y=1.492 $X2=0 $Y2=0
cc_153 N_A2_c_130_n N_A_45_74#_c_591_n 0.0116093f $X=1.425 $Y=1.22 $X2=0 $Y2=0
cc_154 N_A2_c_131_n N_A_45_74#_c_591_n 0.00924272f $X=1.855 $Y=1.22 $X2=0 $Y2=0
cc_155 N_A2_c_132_n N_A_45_74#_c_591_n 0.0324746f $X=1.925 $Y=1.385 $X2=0 $Y2=0
cc_156 N_A2_c_133_n N_A_45_74#_c_591_n 0.00239267f $X=1.91 $Y=1.492 $X2=0 $Y2=0
cc_157 N_A2_c_130_n N_VGND_c_611_n 5.54504e-19 $X=1.425 $Y=1.22 $X2=0 $Y2=0
cc_158 N_A2_c_130_n N_VGND_c_614_n 0.00433162f $X=1.425 $Y=1.22 $X2=0 $Y2=0
cc_159 N_A2_c_131_n N_VGND_c_614_n 0.00291649f $X=1.855 $Y=1.22 $X2=0 $Y2=0
cc_160 N_A2_c_130_n N_VGND_c_616_n 0.00432528f $X=1.425 $Y=1.22 $X2=0 $Y2=0
cc_161 N_A2_c_131_n N_VGND_c_616_n 0.0036412f $X=1.855 $Y=1.22 $X2=0 $Y2=0
cc_162 N_A2_c_130_n N_A_300_74#_c_662_n 0.00337267f $X=1.425 $Y=1.22 $X2=0 $Y2=0
cc_163 N_A2_c_131_n N_A_300_74#_c_662_n 0.0132302f $X=1.855 $Y=1.22 $X2=0 $Y2=0
cc_164 N_A1_M1015_g N_B1_M1014_g 0.0200484f $X=3.365 $Y=0.74 $X2=0 $Y2=0
cc_165 N_A1_c_188_n B1 0.0284542f $X=2.87 $Y=1.45 $X2=0 $Y2=0
cc_166 N_A1_c_189_n B1 0.00280225f $X=3.035 $Y=1.515 $X2=0 $Y2=0
cc_167 N_A1_c_188_n N_B1_c_239_n 9.99318e-19 $X=2.87 $Y=1.45 $X2=0 $Y2=0
cc_168 N_A1_c_189_n N_B1_c_239_n 0.0120684f $X=3.035 $Y=1.515 $X2=0 $Y2=0
cc_169 N_A1_c_190_n N_VPWR_c_332_n 0.0153393f $X=2.39 $Y=1.765 $X2=0 $Y2=0
cc_170 N_A1_c_191_n N_VPWR_c_332_n 5.89254e-19 $X=2.84 $Y=1.765 $X2=0 $Y2=0
cc_171 N_A1_c_190_n N_VPWR_c_333_n 5.35985e-19 $X=2.39 $Y=1.765 $X2=0 $Y2=0
cc_172 N_A1_c_191_n N_VPWR_c_333_n 0.0124262f $X=2.84 $Y=1.765 $X2=0 $Y2=0
cc_173 N_A1_c_190_n N_VPWR_c_335_n 0.00413917f $X=2.39 $Y=1.765 $X2=0 $Y2=0
cc_174 N_A1_c_191_n N_VPWR_c_335_n 0.00413917f $X=2.84 $Y=1.765 $X2=0 $Y2=0
cc_175 N_A1_c_190_n N_VPWR_c_327_n 0.00817726f $X=2.39 $Y=1.765 $X2=0 $Y2=0
cc_176 N_A1_c_191_n N_VPWR_c_327_n 0.00817726f $X=2.84 $Y=1.765 $X2=0 $Y2=0
cc_177 N_A1_c_190_n N_A_127_368#_c_402_n 0.00108467f $X=2.39 $Y=1.765 $X2=0
+ $Y2=0
cc_178 N_A1_c_190_n N_A_127_368#_c_403_n 0.0099355f $X=2.39 $Y=1.765 $X2=0 $Y2=0
cc_179 N_A1_c_188_n N_A_127_368#_c_403_n 0.0159735f $X=2.87 $Y=1.45 $X2=0 $Y2=0
cc_180 N_A1_c_189_n N_A_127_368#_c_403_n 0.00579656f $X=3.035 $Y=1.515 $X2=0
+ $Y2=0
cc_181 N_A1_c_191_n N_A_127_368#_c_405_n 0.015443f $X=2.84 $Y=1.765 $X2=0 $Y2=0
cc_182 N_A1_c_188_n N_A_127_368#_c_405_n 0.0316215f $X=2.87 $Y=1.45 $X2=0 $Y2=0
cc_183 N_A1_c_189_n N_A_127_368#_c_405_n 0.0088446f $X=3.035 $Y=1.515 $X2=0
+ $Y2=0
cc_184 N_A1_c_190_n N_A_127_368#_c_407_n 0.00667324f $X=2.39 $Y=1.765 $X2=0
+ $Y2=0
cc_185 N_A1_c_191_n N_A_127_368#_c_407_n 0.00947771f $X=2.84 $Y=1.765 $X2=0
+ $Y2=0
cc_186 N_A1_c_188_n N_A_127_368#_c_407_n 0.0182032f $X=2.87 $Y=1.45 $X2=0 $Y2=0
cc_187 N_A1_c_189_n N_A_127_368#_c_407_n 0.00512635f $X=3.035 $Y=1.515 $X2=0
+ $Y2=0
cc_188 N_A1_c_191_n N_A_692_368#_c_471_n 9.88057e-19 $X=2.84 $Y=1.765 $X2=0
+ $Y2=0
cc_189 N_A1_c_191_n N_A_692_368#_c_473_n 5.75404e-19 $X=2.84 $Y=1.765 $X2=0
+ $Y2=0
cc_190 N_A1_M1006_g N_Y_c_518_n 0.0144828f $X=2.935 $Y=0.74 $X2=0 $Y2=0
cc_191 N_A1_M1015_g N_Y_c_518_n 0.0192938f $X=3.365 $Y=0.74 $X2=0 $Y2=0
cc_192 N_A1_c_188_n N_Y_c_518_n 0.0528772f $X=2.87 $Y=1.45 $X2=0 $Y2=0
cc_193 N_A1_c_189_n N_Y_c_518_n 0.00867365f $X=3.035 $Y=1.515 $X2=0 $Y2=0
cc_194 N_A1_M1015_g N_Y_c_519_n 4.15473e-19 $X=3.365 $Y=0.74 $X2=0 $Y2=0
cc_195 N_A1_M1006_g N_VGND_c_614_n 0.00291649f $X=2.935 $Y=0.74 $X2=0 $Y2=0
cc_196 N_A1_M1015_g N_VGND_c_614_n 0.00433162f $X=3.365 $Y=0.74 $X2=0 $Y2=0
cc_197 N_A1_M1006_g N_VGND_c_616_n 0.0036412f $X=2.935 $Y=0.74 $X2=0 $Y2=0
cc_198 N_A1_M1015_g N_VGND_c_616_n 0.00449183f $X=3.365 $Y=0.74 $X2=0 $Y2=0
cc_199 N_A1_M1006_g N_A_300_74#_c_661_n 0.00479781f $X=2.935 $Y=0.74 $X2=0 $Y2=0
cc_200 N_A1_M1015_g N_A_300_74#_c_661_n 0.00420713f $X=3.365 $Y=0.74 $X2=0 $Y2=0
cc_201 N_A1_M1006_g N_A_300_74#_c_662_n 0.0122192f $X=2.935 $Y=0.74 $X2=0 $Y2=0
cc_202 N_B1_M1014_g N_C1_M1017_g 0.0105379f $X=3.795 $Y=0.74 $X2=0 $Y2=0
cc_203 N_B1_c_241_n N_C1_c_288_n 0.0105683f $X=4.26 $Y=1.765 $X2=0 $Y2=0
cc_204 B1 N_C1_c_288_n 0.00178648f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_205 B1 N_C1_c_286_n 0.0163092f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_206 N_B1_c_239_n N_C1_c_286_n 0.0256033f $X=4.185 $Y=1.515 $X2=0 $Y2=0
cc_207 B1 N_C1_c_287_n 0.0345267f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_208 N_B1_c_240_n N_VPWR_c_333_n 0.00181484f $X=3.81 $Y=1.765 $X2=0 $Y2=0
cc_209 N_B1_c_240_n N_VPWR_c_336_n 0.00278252f $X=3.81 $Y=1.765 $X2=0 $Y2=0
cc_210 N_B1_c_241_n N_VPWR_c_336_n 0.00278257f $X=4.26 $Y=1.765 $X2=0 $Y2=0
cc_211 N_B1_c_240_n N_VPWR_c_327_n 0.00358623f $X=3.81 $Y=1.765 $X2=0 $Y2=0
cc_212 N_B1_c_241_n N_VPWR_c_327_n 0.00353905f $X=4.26 $Y=1.765 $X2=0 $Y2=0
cc_213 N_B1_c_240_n N_A_127_368#_c_405_n 0.0144529f $X=3.81 $Y=1.765 $X2=0 $Y2=0
cc_214 B1 N_A_127_368#_c_405_n 0.0304867f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_215 N_B1_c_241_n N_A_127_368#_c_443_n 0.00228378f $X=4.26 $Y=1.765 $X2=0
+ $Y2=0
cc_216 B1 N_A_127_368#_c_443_n 0.0164744f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_217 N_B1_c_239_n N_A_127_368#_c_443_n 0.00115938f $X=4.185 $Y=1.515 $X2=0
+ $Y2=0
cc_218 N_B1_c_240_n N_A_692_368#_c_471_n 0.00772703f $X=3.81 $Y=1.765 $X2=0
+ $Y2=0
cc_219 N_B1_c_241_n N_A_692_368#_c_471_n 5.56897e-19 $X=4.26 $Y=1.765 $X2=0
+ $Y2=0
cc_220 N_B1_c_240_n N_A_692_368#_c_472_n 0.0105163f $X=3.81 $Y=1.765 $X2=0 $Y2=0
cc_221 N_B1_c_241_n N_A_692_368#_c_472_n 0.0108414f $X=4.26 $Y=1.765 $X2=0 $Y2=0
cc_222 N_B1_c_240_n N_A_692_368#_c_473_n 0.00273404f $X=3.81 $Y=1.765 $X2=0
+ $Y2=0
cc_223 N_B1_c_240_n N_A_692_368#_c_484_n 6.2215e-19 $X=3.81 $Y=1.765 $X2=0 $Y2=0
cc_224 N_B1_c_241_n N_A_692_368#_c_484_n 0.0110801f $X=4.26 $Y=1.765 $X2=0 $Y2=0
cc_225 B1 N_A_692_368#_c_484_n 0.0235972f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_226 N_B1_c_241_n N_A_692_368#_c_476_n 0.00171731f $X=4.26 $Y=1.765 $X2=0
+ $Y2=0
cc_227 B1 N_Y_c_518_n 8.08061e-19 $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_228 N_B1_M1014_g N_Y_c_519_n 0.00654828f $X=3.795 $Y=0.74 $X2=0 $Y2=0
cc_229 N_B1_M1014_g N_Y_c_520_n 0.00909025f $X=3.795 $Y=0.74 $X2=0 $Y2=0
cc_230 B1 N_Y_c_520_n 0.0221514f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_231 N_B1_c_239_n N_Y_c_520_n 9.31826e-19 $X=4.185 $Y=1.515 $X2=0 $Y2=0
cc_232 N_B1_M1014_g N_Y_c_523_n 0.0104686f $X=3.795 $Y=0.74 $X2=0 $Y2=0
cc_233 B1 N_Y_c_523_n 0.0720188f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_234 N_B1_c_239_n N_Y_c_523_n 0.0114608f $X=4.185 $Y=1.515 $X2=0 $Y2=0
cc_235 N_B1_M1014_g N_VGND_c_612_n 0.00509642f $X=3.795 $Y=0.74 $X2=0 $Y2=0
cc_236 N_B1_M1014_g N_VGND_c_614_n 0.00434272f $X=3.795 $Y=0.74 $X2=0 $Y2=0
cc_237 N_B1_M1014_g N_VGND_c_616_n 0.00822954f $X=3.795 $Y=0.74 $X2=0 $Y2=0
cc_238 N_C1_c_288_n N_VPWR_c_336_n 0.00278257f $X=4.71 $Y=1.765 $X2=0 $Y2=0
cc_239 N_C1_c_289_n N_VPWR_c_336_n 0.00278257f $X=5.16 $Y=1.765 $X2=0 $Y2=0
cc_240 N_C1_c_288_n N_VPWR_c_327_n 0.00353905f $X=4.71 $Y=1.765 $X2=0 $Y2=0
cc_241 N_C1_c_289_n N_VPWR_c_327_n 0.00357591f $X=5.16 $Y=1.765 $X2=0 $Y2=0
cc_242 N_C1_c_288_n N_A_692_368#_c_484_n 0.0110935f $X=4.71 $Y=1.765 $X2=0 $Y2=0
cc_243 N_C1_c_289_n N_A_692_368#_c_484_n 6.23098e-19 $X=5.16 $Y=1.765 $X2=0
+ $Y2=0
cc_244 N_C1_c_286_n N_A_692_368#_c_484_n 2.60261e-19 $X=5.01 $Y=1.515 $X2=0
+ $Y2=0
cc_245 N_C1_c_288_n N_A_692_368#_c_474_n 0.0108414f $X=4.71 $Y=1.765 $X2=0 $Y2=0
cc_246 N_C1_c_289_n N_A_692_368#_c_474_n 0.0134708f $X=5.16 $Y=1.765 $X2=0 $Y2=0
cc_247 N_C1_c_288_n N_A_692_368#_c_475_n 5.7112e-19 $X=4.71 $Y=1.765 $X2=0 $Y2=0
cc_248 N_C1_c_289_n N_A_692_368#_c_475_n 0.00766499f $X=5.16 $Y=1.765 $X2=0
+ $Y2=0
cc_249 N_C1_c_288_n N_A_692_368#_c_476_n 0.00171731f $X=4.71 $Y=1.765 $X2=0
+ $Y2=0
cc_250 N_C1_c_289_n N_Y_c_524_n 0.015921f $X=5.16 $Y=1.765 $X2=0 $Y2=0
cc_251 N_C1_c_287_n N_Y_c_524_n 0.00957882f $X=5.01 $Y=1.515 $X2=0 $Y2=0
cc_252 N_C1_c_288_n N_Y_c_542_n 0.00222151f $X=4.71 $Y=1.765 $X2=0 $Y2=0
cc_253 N_C1_c_289_n N_Y_c_542_n 0.00497407f $X=5.16 $Y=1.765 $X2=0 $Y2=0
cc_254 N_C1_c_286_n N_Y_c_542_n 0.00104557f $X=5.01 $Y=1.515 $X2=0 $Y2=0
cc_255 N_C1_c_287_n N_Y_c_542_n 0.0150976f $X=5.01 $Y=1.515 $X2=0 $Y2=0
cc_256 N_C1_M1017_g Y 0.0186914f $X=4.635 $Y=0.74 $X2=0 $Y2=0
cc_257 N_C1_c_286_n Y 0.012565f $X=5.01 $Y=1.515 $X2=0 $Y2=0
cc_258 N_C1_c_287_n Y 0.0281815f $X=5.01 $Y=1.515 $X2=0 $Y2=0
cc_259 N_C1_M1017_g Y 0.00350742f $X=4.635 $Y=0.74 $X2=0 $Y2=0
cc_260 N_C1_c_289_n Y 0.00629738f $X=5.16 $Y=1.765 $X2=0 $Y2=0
cc_261 N_C1_c_286_n Y 0.0108744f $X=5.01 $Y=1.515 $X2=0 $Y2=0
cc_262 N_C1_c_287_n Y 0.026353f $X=5.01 $Y=1.515 $X2=0 $Y2=0
cc_263 N_C1_M1017_g N_Y_c_523_n 0.010805f $X=4.635 $Y=0.74 $X2=0 $Y2=0
cc_264 N_C1_M1017_g N_VGND_c_612_n 0.00511882f $X=4.635 $Y=0.74 $X2=0 $Y2=0
cc_265 N_C1_M1017_g N_VGND_c_615_n 0.00433162f $X=4.635 $Y=0.74 $X2=0 $Y2=0
cc_266 N_C1_M1017_g N_VGND_c_616_n 0.00824204f $X=4.635 $Y=0.74 $X2=0 $Y2=0
cc_267 N_VPWR_c_329_n N_A_127_368#_c_399_n 0.0730823f $X=0.335 $Y=1.985 $X2=0
+ $Y2=0
cc_268 N_VPWR_c_330_n N_A_127_368#_c_399_n 0.014552f $X=1.15 $Y=3.33 $X2=0 $Y2=0
cc_269 N_VPWR_c_331_n N_A_127_368#_c_399_n 0.0599532f $X=1.235 $Y=2.225 $X2=0
+ $Y2=0
cc_270 N_VPWR_c_327_n N_A_127_368#_c_399_n 0.0119791f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_271 N_VPWR_M1008_s N_A_127_368#_c_400_n 0.00247267f $X=1.085 $Y=1.84 $X2=0
+ $Y2=0
cc_272 N_VPWR_c_331_n N_A_127_368#_c_400_n 0.0136682f $X=1.235 $Y=2.225 $X2=0
+ $Y2=0
cc_273 N_VPWR_c_329_n N_A_127_368#_c_401_n 0.00501285f $X=0.335 $Y=1.985 $X2=0
+ $Y2=0
cc_274 N_VPWR_c_331_n N_A_127_368#_c_402_n 0.0599532f $X=1.235 $Y=2.225 $X2=0
+ $Y2=0
cc_275 N_VPWR_c_332_n N_A_127_368#_c_402_n 0.0622532f $X=2.15 $Y=2.225 $X2=0
+ $Y2=0
cc_276 N_VPWR_c_334_n N_A_127_368#_c_402_n 0.014552f $X=2.05 $Y=3.33 $X2=0 $Y2=0
cc_277 N_VPWR_c_327_n N_A_127_368#_c_402_n 0.0119791f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_278 N_VPWR_M1016_s N_A_127_368#_c_403_n 0.00254385f $X=1.985 $Y=1.84 $X2=0
+ $Y2=0
cc_279 N_VPWR_c_332_n N_A_127_368#_c_403_n 0.0178655f $X=2.15 $Y=2.225 $X2=0
+ $Y2=0
cc_280 N_VPWR_c_333_n N_A_127_368#_c_404_n 0.0449718f $X=3.065 $Y=2.405 $X2=0
+ $Y2=0
cc_281 N_VPWR_c_335_n N_A_127_368#_c_404_n 0.00749631f $X=2.9 $Y=3.33 $X2=0
+ $Y2=0
cc_282 N_VPWR_c_327_n N_A_127_368#_c_404_n 0.0062048f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_283 N_VPWR_M1011_s N_A_127_368#_c_405_n 0.0050911f $X=2.915 $Y=1.84 $X2=0
+ $Y2=0
cc_284 N_VPWR_c_333_n N_A_127_368#_c_405_n 0.0220544f $X=3.065 $Y=2.405 $X2=0
+ $Y2=0
cc_285 N_VPWR_c_332_n N_A_127_368#_c_407_n 0.0591677f $X=2.15 $Y=2.225 $X2=0
+ $Y2=0
cc_286 N_VPWR_c_333_n N_A_692_368#_c_471_n 0.0473719f $X=3.065 $Y=2.405 $X2=0
+ $Y2=0
cc_287 N_VPWR_c_336_n N_A_692_368#_c_472_n 0.0355725f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_288 N_VPWR_c_327_n N_A_692_368#_c_472_n 0.0200299f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_289 N_VPWR_c_333_n N_A_692_368#_c_473_n 0.0139f $X=3.065 $Y=2.405 $X2=0 $Y2=0
cc_290 N_VPWR_c_336_n N_A_692_368#_c_473_n 0.0239448f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_291 N_VPWR_c_327_n N_A_692_368#_c_473_n 0.0129325f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_292 N_VPWR_c_336_n N_A_692_368#_c_474_n 0.0594839f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_293 N_VPWR_c_327_n N_A_692_368#_c_474_n 0.0329562f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_294 N_VPWR_c_336_n N_A_692_368#_c_476_n 0.0235512f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_295 N_VPWR_c_327_n N_A_692_368#_c_476_n 0.0126924f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_296 N_A_127_368#_c_405_n N_A_692_368#_M1000_d 0.00621129f $X=3.925 $Y=2.035
+ $X2=-0.19 $Y2=1.66
cc_297 N_A_127_368#_c_405_n N_A_692_368#_c_471_n 0.0224353f $X=3.925 $Y=2.035
+ $X2=0 $Y2=0
cc_298 N_A_127_368#_M1000_s N_A_692_368#_c_472_n 0.00222494f $X=3.885 $Y=1.84
+ $X2=0 $Y2=0
cc_299 N_A_127_368#_c_443_n N_A_692_368#_c_472_n 0.013472f $X=4.035 $Y=2.115
+ $X2=0 $Y2=0
cc_300 N_A_127_368#_c_443_n N_A_692_368#_c_484_n 0.0528196f $X=4.035 $Y=2.115
+ $X2=0 $Y2=0
cc_301 N_A_127_368#_c_403_n N_A_45_74#_c_579_n 0.00418019f $X=2.53 $Y=1.805
+ $X2=0 $Y2=0
cc_302 N_A_692_368#_c_474_n N_Y_M1001_d 0.00247267f $X=5.22 $Y=2.99 $X2=0 $Y2=0
cc_303 N_A_692_368#_M1003_s N_Y_c_524_n 0.0075088f $X=5.235 $Y=1.84 $X2=0 $Y2=0
cc_304 N_A_692_368#_c_475_n N_Y_c_524_n 0.0232575f $X=5.385 $Y=2.425 $X2=0 $Y2=0
cc_305 N_A_692_368#_c_484_n N_Y_c_542_n 0.0524087f $X=4.485 $Y=2.07 $X2=0 $Y2=0
cc_306 N_A_692_368#_c_474_n N_Y_c_542_n 0.012787f $X=5.22 $Y=2.99 $X2=0 $Y2=0
cc_307 N_A_692_368#_c_475_n N_Y_c_542_n 0.0289859f $X=5.385 $Y=2.425 $X2=0 $Y2=0
cc_308 N_A_692_368#_M1003_s Y 0.00188446f $X=5.235 $Y=1.84 $X2=0 $Y2=0
cc_309 N_Y_c_518_n N_A_45_74#_c_579_n 0.0118023f $X=3.495 $Y=1.015 $X2=0 $Y2=0
cc_310 N_Y_c_523_n N_VGND_M1014_d 0.00793129f $X=4.685 $Y=0.765 $X2=0 $Y2=0
cc_311 N_Y_c_519_n N_VGND_c_612_n 0.0184853f $X=3.58 $Y=0.515 $X2=0 $Y2=0
cc_312 Y N_VGND_c_612_n 0.0214218f $X=5.435 $Y=0.47 $X2=0 $Y2=0
cc_313 N_Y_c_523_n N_VGND_c_612_n 0.0468625f $X=4.685 $Y=0.765 $X2=0 $Y2=0
cc_314 N_Y_c_519_n N_VGND_c_614_n 0.0109942f $X=3.58 $Y=0.515 $X2=0 $Y2=0
cc_315 Y N_VGND_c_615_n 0.0421459f $X=5.435 $Y=0.47 $X2=0 $Y2=0
cc_316 N_Y_c_518_n N_VGND_c_616_n 0.00699508f $X=3.495 $Y=1.015 $X2=0 $Y2=0
cc_317 N_Y_c_519_n N_VGND_c_616_n 0.00904371f $X=3.58 $Y=0.515 $X2=0 $Y2=0
cc_318 Y N_VGND_c_616_n 0.0349449f $X=5.435 $Y=0.47 $X2=0 $Y2=0
cc_319 N_Y_c_518_n N_A_300_74#_M1006_s 0.00178215f $X=3.495 $Y=1.015 $X2=0 $Y2=0
cc_320 N_Y_c_518_n N_A_300_74#_c_661_n 0.0165836f $X=3.495 $Y=1.015 $X2=0 $Y2=0
cc_321 N_Y_c_519_n N_A_300_74#_c_661_n 0.0135554f $X=3.58 $Y=0.515 $X2=0 $Y2=0
cc_322 N_Y_M1006_d N_A_300_74#_c_662_n 0.00374227f $X=2.595 $Y=0.37 $X2=0 $Y2=0
cc_323 N_Y_c_518_n N_A_300_74#_c_662_n 0.0201119f $X=3.495 $Y=1.015 $X2=0 $Y2=0
cc_324 N_A_45_74#_c_581_n N_VGND_M1004_d 0.00406005f $X=1.125 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_325 N_A_45_74#_c_576_n N_VGND_c_611_n 0.0121972f $X=0.35 $Y=0.515 $X2=0 $Y2=0
cc_326 N_A_45_74#_c_581_n N_VGND_c_611_n 0.0167019f $X=1.125 $Y=0.925 $X2=0
+ $Y2=0
cc_327 N_A_45_74#_c_578_n N_VGND_c_611_n 0.0135953f $X=1.21 $Y=0.495 $X2=0 $Y2=0
cc_328 N_A_45_74#_c_576_n N_VGND_c_613_n 0.0110895f $X=0.35 $Y=0.515 $X2=0 $Y2=0
cc_329 N_A_45_74#_c_578_n N_VGND_c_614_n 0.00814895f $X=1.21 $Y=0.495 $X2=0
+ $Y2=0
cc_330 N_A_45_74#_c_576_n N_VGND_c_616_n 0.00916858f $X=0.35 $Y=0.515 $X2=0
+ $Y2=0
cc_331 N_A_45_74#_c_581_n N_VGND_c_616_n 0.0116543f $X=1.125 $Y=0.925 $X2=0
+ $Y2=0
cc_332 N_A_45_74#_c_578_n N_VGND_c_616_n 0.00627841f $X=1.21 $Y=0.495 $X2=0
+ $Y2=0
cc_333 N_A_45_74#_c_591_n N_VGND_c_616_n 0.0070825f $X=1.905 $Y=0.91 $X2=0 $Y2=0
cc_334 N_A_45_74#_c_591_n N_A_300_74#_M1002_s 0.0034629f $X=1.905 $Y=0.91
+ $X2=-0.19 $Y2=-0.245
cc_335 N_A_45_74#_M1012_d N_A_300_74#_c_662_n 0.0032303f $X=1.93 $Y=0.37 $X2=0
+ $Y2=0
cc_336 N_A_45_74#_c_578_n N_A_300_74#_c_662_n 0.010629f $X=1.21 $Y=0.495 $X2=0
+ $Y2=0
cc_337 N_A_45_74#_c_591_n N_A_300_74#_c_662_n 0.0430812f $X=1.905 $Y=0.91 $X2=0
+ $Y2=0
cc_338 N_VGND_c_614_n N_A_300_74#_c_662_n 0.0755134f $X=3.915 $Y=0 $X2=0 $Y2=0
cc_339 N_VGND_c_616_n N_A_300_74#_c_662_n 0.064201f $X=5.52 $Y=0 $X2=0 $Y2=0
