* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
M1000 a_1525_212# RESET_B VPWR VPB phighvt w=420000u l=150000u
+  ad=2.352e+11p pd=1.96e+06u as=2.3127e+12p ps=2.018e+07u
M1001 VGND RESET_B a_901_138# VNB nshort w=420000u l=150000u
+  ad=1.94642e+12p pd=1.538e+07u as=8.82e+10p ps=1.26e+06u
M1002 a_1478_493# a_495_390# a_1271_74# VPB phighvt w=420000u l=150000u
+  ad=1.134e+11p pd=1.38e+06u as=4.53925e+11p ps=3.66e+06u
M1003 a_1271_74# a_495_390# a_839_359# VNB nshort w=740000u l=150000u
+  ad=4.58e+11p pd=3.28e+06u as=2.405e+11p ps=2.13e+06u
M1004 a_495_390# a_309_390# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.65e+11p pd=2.53e+06u as=0p ps=0u
M1005 VGND a_1525_212# a_1481_81# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1006 a_901_138# a_839_359# a_823_138# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1007 a_697_463# RESET_B VPWR VPB phighvt w=420000u l=150000u
+  ad=2.73e+11p pd=2.98e+06u as=0p ps=0u
M1008 a_697_463# a_495_390# a_30_78# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=2.373e+11p ps=2.81e+06u
M1009 VGND RESET_B a_117_78# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1010 VPWR a_839_359# a_798_463# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1011 a_798_463# a_309_390# a_697_463# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_495_390# a_309_390# VGND VNB nshort w=740000u l=150000u
+  ad=2.0885e+11p pd=2.07e+06u as=0p ps=0u
M1013 a_1271_74# a_309_390# a_839_359# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=3.68125e+11p ps=2.86e+06u
M1014 a_823_138# a_495_390# a_697_463# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.47e+11p ps=1.54e+06u
M1015 VGND CLK a_309_390# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.646e+11p ps=2.4e+06u
M1016 a_697_463# a_309_390# a_30_78# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=2.394e+11p ps=2.82e+06u
M1017 a_1663_81# RESET_B VGND VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1018 a_1525_212# a_1271_74# a_1663_81# VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1019 a_1921_409# a_1271_74# VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1020 a_839_359# a_697_463# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 Q a_1921_409# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=0p ps=0u
M1022 a_30_78# D VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VPWR RESET_B a_30_78# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_1921_409# a_1271_74# VPWR VPB phighvt w=840000u l=150000u
+  ad=2.478e+11p pd=2.27e+06u as=0p ps=0u
M1025 a_117_78# D a_30_78# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VPWR a_1525_212# a_1478_493# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VPWR CLK a_309_390# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.688e+11p ps=2.57e+06u
M1028 a_839_359# a_697_463# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 Q a_1921_409# VGND VNB nshort w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1030 VPWR a_1921_409# Q VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_1481_81# a_309_390# a_1271_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 VGND a_1921_409# Q VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VPWR a_1271_74# a_1525_212# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
