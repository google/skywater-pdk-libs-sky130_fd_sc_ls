* NGSPICE file created from sky130_fd_sc_ls__and4bb_2.ext - technology: sky130A

.subckt sky130_fd_sc_ls__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
M1000 VPWR A_N a_27_74# VPB phighvt w=840000u l=150000u
+  ad=1.9728e+12p pd=1.236e+07u as=2.478e+11p ps=2.27e+06u
M1001 X a_225_82# VGND VNB nshort w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=1.0454e+12p ps=7.35e+06u
M1002 a_312_82# a_27_74# a_225_82# VNB nshort w=740000u l=150000u
+  ad=1.776e+11p pd=1.96e+06u as=2.109e+11p ps=2.05e+06u
M1003 a_390_82# a_354_252# a_312_82# VNB nshort w=740000u l=150000u
+  ad=2.886e+11p pd=2.26e+06u as=0p ps=0u
M1004 a_354_252# B_N VPWR VPB phighvt w=840000u l=150000u
+  ad=2.604e+11p pd=2.3e+06u as=0p ps=0u
M1005 a_354_252# B_N VGND VNB nshort w=550000u l=150000u
+  ad=1.5675e+11p pd=1.67e+06u as=0p ps=0u
M1006 a_225_82# C VPWR VPB phighvt w=1e+06u l=150000u
+  ad=8.7e+11p pd=5.74e+06u as=0p ps=0u
M1007 X a_225_82# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=0p ps=0u
M1008 VGND a_225_82# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR a_354_252# a_225_82# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_498_82# C a_390_82# VNB nshort w=740000u l=150000u
+  ad=2.664e+11p pd=2.2e+06u as=0p ps=0u
M1011 VPWR D a_225_82# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR a_225_82# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND D a_498_82# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_225_82# a_27_74# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND A_N a_27_74# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
.ends

