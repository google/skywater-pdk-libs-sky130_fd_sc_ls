* File: sky130_fd_sc_ls__a22o_4.pxi.spice
* Created: Fri Aug 28 12:55:16 2020
* 
x_PM_SKY130_FD_SC_LS__A22O_4%A_95_306# N_A_95_306#_M1000_d N_A_95_306#_M1003_d
+ N_A_95_306#_M1009_d N_A_95_306#_M1014_d N_A_95_306#_c_147_n
+ N_A_95_306#_M1007_g N_A_95_306#_c_131_n N_A_95_306#_c_149_n
+ N_A_95_306#_M1008_g N_A_95_306#_c_132_n N_A_95_306#_M1002_g
+ N_A_95_306#_c_151_n N_A_95_306#_M1013_g N_A_95_306#_c_134_n
+ N_A_95_306#_c_135_n N_A_95_306#_c_136_n N_A_95_306#_M1004_g
+ N_A_95_306#_c_154_n N_A_95_306#_M1019_g N_A_95_306#_c_137_n
+ N_A_95_306#_M1017_g N_A_95_306#_c_138_n N_A_95_306#_M1020_g
+ N_A_95_306#_c_139_n N_A_95_306#_c_140_n N_A_95_306#_c_221_p
+ N_A_95_306#_c_141_n N_A_95_306#_c_158_n N_A_95_306#_c_159_n
+ N_A_95_306#_c_160_n N_A_95_306#_c_142_n N_A_95_306#_c_162_n
+ N_A_95_306#_c_163_n N_A_95_306#_c_143_n N_A_95_306#_c_144_n
+ N_A_95_306#_c_145_n N_A_95_306#_c_146_n PM_SKY130_FD_SC_LS__A22O_4%A_95_306#
x_PM_SKY130_FD_SC_LS__A22O_4%B2 N_B2_c_323_n N_B2_M1009_g N_B2_M1021_g
+ N_B2_c_325_n N_B2_M1015_g N_B2_M1023_g N_B2_c_332_n N_B2_c_333_n N_B2_c_327_n
+ N_B2_c_328_n N_B2_c_329_n N_B2_c_359_n B2 B2 N_B2_c_336_n
+ PM_SKY130_FD_SC_LS__A22O_4%B2
x_PM_SKY130_FD_SC_LS__A22O_4%B1 N_B1_c_423_n N_B1_M1010_g N_B1_M1000_g
+ N_B1_M1018_g N_B1_c_424_n N_B1_M1014_g B1 N_B1_c_422_n
+ PM_SKY130_FD_SC_LS__A22O_4%B1
x_PM_SKY130_FD_SC_LS__A22O_4%A1 N_A1_c_477_n N_A1_M1005_g N_A1_M1003_g
+ N_A1_c_478_n N_A1_M1011_g N_A1_M1016_g A1 A1 N_A1_c_476_n
+ PM_SKY130_FD_SC_LS__A22O_4%A1
x_PM_SKY130_FD_SC_LS__A22O_4%A2 N_A2_c_526_n N_A2_c_536_n N_A2_M1006_g
+ N_A2_M1001_g N_A2_c_528_n N_A2_c_529_n N_A2_c_530_n N_A2_c_538_n N_A2_M1012_g
+ N_A2_M1022_g N_A2_c_532_n A2 N_A2_c_534_n PM_SKY130_FD_SC_LS__A22O_4%A2
x_PM_SKY130_FD_SC_LS__A22O_4%VPWR N_VPWR_M1007_s N_VPWR_M1008_s N_VPWR_M1019_s
+ N_VPWR_M1006_d N_VPWR_M1011_d N_VPWR_c_594_n N_VPWR_c_595_n N_VPWR_c_596_n
+ N_VPWR_c_597_n N_VPWR_c_598_n N_VPWR_c_599_n N_VPWR_c_600_n N_VPWR_c_601_n
+ VPWR N_VPWR_c_602_n N_VPWR_c_603_n N_VPWR_c_604_n N_VPWR_c_605_n
+ N_VPWR_c_593_n N_VPWR_c_607_n N_VPWR_c_608_n N_VPWR_c_609_n
+ PM_SKY130_FD_SC_LS__A22O_4%VPWR
x_PM_SKY130_FD_SC_LS__A22O_4%X N_X_M1002_d N_X_M1017_d N_X_M1007_d N_X_M1013_d
+ N_X_c_687_n N_X_c_682_n N_X_c_688_n N_X_c_706_n N_X_c_683_n N_X_c_684_n
+ N_X_c_718_n X X N_X_c_686_n PM_SKY130_FD_SC_LS__A22O_4%X
x_PM_SKY130_FD_SC_LS__A22O_4%A_555_392# N_A_555_392#_M1009_s
+ N_A_555_392#_M1010_s N_A_555_392#_M1015_s N_A_555_392#_M1005_s
+ N_A_555_392#_M1012_s N_A_555_392#_c_749_n N_A_555_392#_c_763_n
+ N_A_555_392#_c_750_n N_A_555_392#_c_784_n N_A_555_392#_c_751_n
+ N_A_555_392#_c_752_n N_A_555_392#_c_753_n N_A_555_392#_c_754_n
+ N_A_555_392#_c_755_n N_A_555_392#_c_768_n N_A_555_392#_c_756_n
+ N_A_555_392#_c_757_n PM_SKY130_FD_SC_LS__A22O_4%A_555_392#
x_PM_SKY130_FD_SC_LS__A22O_4%VGND N_VGND_M1002_s N_VGND_M1004_s N_VGND_M1020_s
+ N_VGND_M1023_d N_VGND_M1022_s N_VGND_c_825_n N_VGND_c_826_n N_VGND_c_827_n
+ N_VGND_c_828_n N_VGND_c_829_n N_VGND_c_830_n N_VGND_c_831_n N_VGND_c_832_n
+ N_VGND_c_833_n N_VGND_c_834_n N_VGND_c_835_n N_VGND_c_836_n N_VGND_c_837_n
+ N_VGND_c_838_n VGND N_VGND_c_839_n N_VGND_c_840_n N_VGND_c_841_n
+ PM_SKY130_FD_SC_LS__A22O_4%VGND
x_PM_SKY130_FD_SC_LS__A22O_4%A_645_120# N_A_645_120#_M1021_s
+ N_A_645_120#_M1018_s N_A_645_120#_c_913_n N_A_645_120#_c_914_n
+ PM_SKY130_FD_SC_LS__A22O_4%A_645_120#
x_PM_SKY130_FD_SC_LS__A22O_4%A_1064_123# N_A_1064_123#_M1001_d
+ N_A_1064_123#_M1016_s N_A_1064_123#_c_933_n N_A_1064_123#_c_930_n
+ N_A_1064_123#_c_931_n PM_SKY130_FD_SC_LS__A22O_4%A_1064_123#
cc_1 VNB N_A_95_306#_c_131_n 0.0110061f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.605
cc_2 VNB N_A_95_306#_c_132_n 0.00734144f $X=-0.19 $Y=-0.245 $X2=1.28 $Y2=1.605
cc_3 VNB N_A_95_306#_M1002_g 0.0278837f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=0.87
cc_4 VNB N_A_95_306#_c_134_n 0.00394382f $X=-0.19 $Y=-0.245 $X2=1.71 $Y2=1.605
cc_5 VNB N_A_95_306#_c_135_n 0.00479405f $X=-0.19 $Y=-0.245 $X2=1.555 $Y2=1.605
cc_6 VNB N_A_95_306#_c_136_n 0.0153169f $X=-0.19 $Y=-0.245 $X2=1.785 $Y2=1.35
cc_7 VNB N_A_95_306#_c_137_n 0.0162201f $X=-0.19 $Y=-0.245 $X2=2.215 $Y2=1.35
cc_8 VNB N_A_95_306#_c_138_n 0.0172571f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=1.35
cc_9 VNB N_A_95_306#_c_139_n 0.014179f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.605
cc_10 VNB N_A_95_306#_c_140_n 0.00762258f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=1.605
cc_11 VNB N_A_95_306#_c_141_n 0.00322996f $X=-0.19 $Y=-0.245 $X2=2.56 $Y2=1.68
cc_12 VNB N_A_95_306#_c_142_n 0.0443678f $X=-0.19 $Y=-0.245 $X2=2.555 $Y2=1.515
cc_13 VNB N_A_95_306#_c_143_n 0.00618103f $X=-0.19 $Y=-0.245 $X2=3.63 $Y2=1.132
cc_14 VNB N_A_95_306#_c_144_n 0.00304687f $X=-0.19 $Y=-0.245 $X2=3.96 $Y2=1.132
cc_15 VNB N_A_95_306#_c_145_n 0.00229391f $X=-0.19 $Y=-0.245 $X2=5.89 $Y2=1.105
cc_16 VNB N_A_95_306#_c_146_n 0.0141457f $X=-0.19 $Y=-0.245 $X2=5.725 $Y2=1.145
cc_17 VNB N_B2_c_323_n 0.0184292f $X=-0.19 $Y=-0.245 $X2=3.655 $Y2=0.6
cc_18 VNB N_B2_M1021_g 0.02243f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_B2_c_325_n 0.0165592f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_B2_M1023_g 0.0230208f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.765
cc_21 VNB N_B2_c_327_n 7.59216e-19 $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=2.4
cc_22 VNB N_B2_c_328_n 0.0037501f $X=-0.19 $Y=-0.245 $X2=1.28 $Y2=1.605
cc_23 VNB N_B2_c_329_n 0.00181489f $X=-0.19 $Y=-0.245 $X2=1.465 $Y2=2.4
cc_24 VNB N_B1_M1000_g 0.0210564f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_B1_M1018_g 0.0217123f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB B1 8.16208e-19 $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=2.4
cc_27 VNB N_B1_c_422_n 0.0251107f $X=-0.19 $Y=-0.245 $X2=1.105 $Y2=1.605
cc_28 VNB N_A1_M1003_g 0.0194032f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A1_M1016_g 0.0193298f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.765
cc_30 VNB A1 0.00392757f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.605
cc_31 VNB N_A1_c_476_n 0.0265391f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=0.87
cc_32 VNB N_A2_c_526_n 0.0109566f $X=-0.19 $Y=-0.245 $X2=5.75 $Y2=0.615
cc_33 VNB N_A2_M1001_g 0.0114364f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A2_c_528_n 0.0902248f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A2_c_529_n 0.00930145f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A2_c_530_n 0.0203142f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.765
cc_37 VNB N_A2_M1022_g 0.0330549f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=2.4
cc_38 VNB N_A2_c_532_n 0.0285121f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=1.53
cc_39 VNB A2 0.0131334f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A2_c_534_n 0.0472248f $X=-0.19 $Y=-0.245 $X2=1.465 $Y2=2.4
cc_41 VNB N_VPWR_c_593_n 0.302998f $X=-0.19 $Y=-0.245 $X2=3.35 $Y2=2.867
cc_42 VNB N_X_c_682_n 0.00251264f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=1.53
cc_43 VNB N_X_c_683_n 0.00252589f $X=-0.19 $Y=-0.245 $X2=1.915 $Y2=1.765
cc_44 VNB N_X_c_684_n 0.00571544f $X=-0.19 $Y=-0.245 $X2=2.215 $Y2=1.35
cc_45 VNB X 0.0131314f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=0.87
cc_46 VNB N_X_c_686_n 0.0457248f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_825_n 0.0371369f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=1.765
cc_48 VNB N_VGND_c_826_n 0.00886349f $X=-0.19 $Y=-0.245 $X2=1.105 $Y2=1.605
cc_49 VNB N_VGND_c_827_n 0.0176237f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_828_n 0.0172788f $X=-0.19 $Y=-0.245 $X2=1.71 $Y2=1.605
cc_51 VNB N_VGND_c_829_n 0.049564f $X=-0.19 $Y=-0.245 $X2=1.785 $Y2=0.87
cc_52 VNB N_VGND_c_830_n 0.0331697f $X=-0.19 $Y=-0.245 $X2=1.915 $Y2=2.4
cc_53 VNB N_VGND_c_831_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=2.215 $Y2=1.35
cc_54 VNB N_VGND_c_832_n 0.0178473f $X=-0.19 $Y=-0.245 $X2=2.215 $Y2=0.87
cc_55 VNB N_VGND_c_833_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=1.35
cc_56 VNB N_VGND_c_834_n 0.0178473f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=0.87
cc_57 VNB N_VGND_c_835_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.605
cc_58 VNB N_VGND_c_836_n 0.0112126f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_837_n 0.0480638f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=1.605
cc_60 VNB N_VGND_c_838_n 0.00528596f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_839_n 0.042264f $X=-0.19 $Y=-0.245 $X2=4.25 $Y2=2.78
cc_62 VNB N_VGND_c_840_n 0.442195f $X=-0.19 $Y=-0.245 $X2=3.795 $Y2=1.09
cc_63 VNB N_VGND_c_841_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=3.96 $Y2=1.132
cc_64 VNB N_A_645_120#_c_913_n 0.00288446f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_645_120#_c_914_n 0.00740647f $X=-0.19 $Y=-0.245 $X2=0.565
+ $Y2=1.765
cc_66 VNB N_A_1064_123#_c_930_n 0.00186167f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_1064_123#_c_931_n 0.00325899f $X=-0.19 $Y=-0.245 $X2=0.565
+ $Y2=1.765
cc_68 VPB N_A_95_306#_c_147_n 0.0190854f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=1.765
cc_69 VPB N_A_95_306#_c_131_n 0.0100889f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.605
cc_70 VPB N_A_95_306#_c_149_n 0.0149757f $X=-0.19 $Y=1.66 $X2=1.015 $Y2=1.765
cc_71 VPB N_A_95_306#_c_132_n 0.00416132f $X=-0.19 $Y=1.66 $X2=1.28 $Y2=1.605
cc_72 VPB N_A_95_306#_c_151_n 0.0152868f $X=-0.19 $Y=1.66 $X2=1.465 $Y2=1.765
cc_73 VPB N_A_95_306#_c_134_n 0.00469763f $X=-0.19 $Y=1.66 $X2=1.71 $Y2=1.605
cc_74 VPB N_A_95_306#_c_135_n 0.00995703f $X=-0.19 $Y=1.66 $X2=1.555 $Y2=1.605
cc_75 VPB N_A_95_306#_c_154_n 0.016533f $X=-0.19 $Y=1.66 $X2=1.915 $Y2=1.765
cc_76 VPB N_A_95_306#_c_139_n 0.00969622f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=1.605
cc_77 VPB N_A_95_306#_c_140_n 0.00594789f $X=-0.19 $Y=1.66 $X2=1.015 $Y2=1.605
cc_78 VPB N_A_95_306#_c_141_n 0.00727707f $X=-0.19 $Y=1.66 $X2=2.56 $Y2=1.68
cc_79 VPB N_A_95_306#_c_158_n 0.0253988f $X=-0.19 $Y=1.66 $X2=2.56 $Y2=2.905
cc_80 VPB N_A_95_306#_c_159_n 0.00354206f $X=-0.19 $Y=1.66 $X2=2.645 $Y2=2.99
cc_81 VPB N_A_95_306#_c_160_n 0.00508424f $X=-0.19 $Y=1.66 $X2=4.25 $Y2=2.78
cc_82 VPB N_A_95_306#_c_142_n 0.0371223f $X=-0.19 $Y=1.66 $X2=2.555 $Y2=1.515
cc_83 VPB N_A_95_306#_c_162_n 0.00851027f $X=-0.19 $Y=1.66 $X2=3.185 $Y2=2.867
cc_84 VPB N_A_95_306#_c_163_n 0.00216917f $X=-0.19 $Y=1.66 $X2=3.515 $Y2=2.867
cc_85 VPB N_B2_c_323_n 0.0364935f $X=-0.19 $Y=1.66 $X2=3.655 $Y2=0.6
cc_86 VPB N_B2_c_325_n 0.0345218f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_B2_c_332_n 0.00175595f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.605
cc_88 VPB N_B2_c_333_n 0.00182275f $X=-0.19 $Y=1.66 $X2=1.015 $Y2=1.765
cc_89 VPB N_B2_c_328_n 0.0032539f $X=-0.19 $Y=1.66 $X2=1.28 $Y2=1.605
cc_90 VPB N_B2_c_329_n 7.66814e-19 $X=-0.19 $Y=1.66 $X2=1.465 $Y2=2.4
cc_91 VPB N_B2_c_336_n 0.00508342f $X=-0.19 $Y=1.66 $X2=2.215 $Y2=1.35
cc_92 VPB N_B1_c_423_n 0.0149201f $X=-0.19 $Y=1.66 $X2=3.655 $Y2=0.6
cc_93 VPB N_B1_c_424_n 0.0152356f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB B1 0.00147474f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=2.4
cc_95 VPB N_B1_c_422_n 0.0312056f $X=-0.19 $Y=1.66 $X2=1.105 $Y2=1.605
cc_96 VPB N_A1_c_477_n 0.0170887f $X=-0.19 $Y=1.66 $X2=3.655 $Y2=0.6
cc_97 VPB N_A1_c_478_n 0.0150823f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB A1 0.00275828f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.605
cc_99 VPB N_A1_c_476_n 0.0340818f $X=-0.19 $Y=1.66 $X2=1.355 $Y2=0.87
cc_100 VPB N_A2_c_526_n 0.00828065f $X=-0.19 $Y=1.66 $X2=5.75 $Y2=0.615
cc_101 VPB N_A2_c_536_n 0.0243148f $X=-0.19 $Y=1.66 $X2=3.2 $Y2=1.96
cc_102 VPB N_A2_c_530_n 0.0113925f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=1.765
cc_103 VPB N_A2_c_538_n 0.0284588f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=2.4
cc_104 VPB N_VPWR_c_594_n 0.0139245f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.605
cc_105 VPB N_VPWR_c_595_n 0.0510315f $X=-0.19 $Y=1.66 $X2=1.015 $Y2=1.765
cc_106 VPB N_VPWR_c_596_n 0.00660498f $X=-0.19 $Y=1.66 $X2=1.355 $Y2=0.87
cc_107 VPB N_VPWR_c_597_n 0.021328f $X=-0.19 $Y=1.66 $X2=1.71 $Y2=1.605
cc_108 VPB N_VPWR_c_598_n 0.0105344f $X=-0.19 $Y=1.66 $X2=1.915 $Y2=2.4
cc_109 VPB N_VPWR_c_599_n 0.00335558f $X=-0.19 $Y=1.66 $X2=2.215 $Y2=0.87
cc_110 VPB N_VPWR_c_600_n 0.0175706f $X=-0.19 $Y=1.66 $X2=2.645 $Y2=0.87
cc_111 VPB N_VPWR_c_601_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=1.605
cc_112 VPB N_VPWR_c_602_n 0.0164465f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_VPWR_c_603_n 0.0206041f $X=-0.19 $Y=1.66 $X2=2.56 $Y2=1.68
cc_114 VPB N_VPWR_c_604_n 0.0677928f $X=-0.19 $Y=1.66 $X2=2.855 $Y2=1.18
cc_115 VPB N_VPWR_c_605_n 0.0235962f $X=-0.19 $Y=1.66 $X2=2.555 $Y2=1.515
cc_116 VPB N_VPWR_c_593_n 0.101648f $X=-0.19 $Y=1.66 $X2=3.35 $Y2=2.867
cc_117 VPB N_VPWR_c_607_n 0.00460249f $X=-0.19 $Y=1.66 $X2=3.63 $Y2=1.132
cc_118 VPB N_VPWR_c_608_n 0.0047828f $X=-0.19 $Y=1.66 $X2=5.89 $Y2=1.105
cc_119 VPB N_VPWR_c_609_n 0.00911062f $X=-0.19 $Y=1.66 $X2=1.785 $Y2=1.557
cc_120 VPB N_X_c_687_n 0.0045716f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=2.4
cc_121 VPB N_X_c_688_n 0.00257348f $X=-0.19 $Y=1.66 $X2=1.465 $Y2=1.765
cc_122 VPB N_A_555_392#_c_749_n 0.00279505f $X=-0.19 $Y=1.66 $X2=1.015 $Y2=1.765
cc_123 VPB N_A_555_392#_c_750_n 0.00419391f $X=-0.19 $Y=1.66 $X2=1.355 $Y2=0.87
cc_124 VPB N_A_555_392#_c_751_n 0.00789967f $X=-0.19 $Y=1.66 $X2=1.465 $Y2=2.4
cc_125 VPB N_A_555_392#_c_752_n 0.00216998f $X=-0.19 $Y=1.66 $X2=1.785 $Y2=1.35
cc_126 VPB N_A_555_392#_c_753_n 0.00746248f $X=-0.19 $Y=1.66 $X2=1.785 $Y2=0.87
cc_127 VPB N_A_555_392#_c_754_n 0.0120331f $X=-0.19 $Y=1.66 $X2=1.915 $Y2=2.4
cc_128 VPB N_A_555_392#_c_755_n 0.0345863f $X=-0.19 $Y=1.66 $X2=2.215 $Y2=1.35
cc_129 VPB N_A_555_392#_c_756_n 0.00253596f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_A_555_392#_c_757_n 0.00143967f $X=-0.19 $Y=1.66 $X2=1.465 $Y2=1.647
cc_131 N_A_95_306#_c_141_n N_B2_c_323_n 0.00182761f $X=2.56 $Y=1.68 $X2=-0.19
+ $Y2=-0.245
cc_132 N_A_95_306#_c_158_n N_B2_c_323_n 0.0082586f $X=2.56 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_133 N_A_95_306#_c_142_n N_B2_c_323_n 0.0139355f $X=2.555 $Y=1.515 $X2=-0.19
+ $Y2=-0.245
cc_134 N_A_95_306#_c_162_n N_B2_c_323_n 0.00966378f $X=3.185 $Y=2.867 $X2=-0.19
+ $Y2=-0.245
cc_135 N_A_95_306#_c_163_n N_B2_c_323_n 0.0059392f $X=3.515 $Y=2.867 $X2=-0.19
+ $Y2=-0.245
cc_136 N_A_95_306#_c_143_n N_B2_c_323_n 0.00497072f $X=3.63 $Y=1.132 $X2=-0.19
+ $Y2=-0.245
cc_137 N_A_95_306#_c_138_n N_B2_M1021_g 0.0233895f $X=2.645 $Y=1.35 $X2=0 $Y2=0
cc_138 N_A_95_306#_c_141_n N_B2_M1021_g 0.00398423f $X=2.56 $Y=1.68 $X2=0 $Y2=0
cc_139 N_A_95_306#_c_143_n N_B2_M1021_g 0.0145118f $X=3.63 $Y=1.132 $X2=0 $Y2=0
cc_140 N_A_95_306#_c_144_n N_B2_M1021_g 4.59187e-19 $X=3.96 $Y=1.132 $X2=0 $Y2=0
cc_141 N_A_95_306#_c_160_n N_B2_c_325_n 0.00382887f $X=4.25 $Y=2.78 $X2=0 $Y2=0
cc_142 N_A_95_306#_c_146_n N_B2_c_325_n 0.00409036f $X=5.725 $Y=1.145 $X2=0
+ $Y2=0
cc_143 N_A_95_306#_c_144_n N_B2_M1023_g 4.50172e-19 $X=3.96 $Y=1.132 $X2=0 $Y2=0
cc_144 N_A_95_306#_c_146_n N_B2_M1023_g 0.015625f $X=5.725 $Y=1.145 $X2=0 $Y2=0
cc_145 N_A_95_306#_c_158_n N_B2_c_332_n 0.00530737f $X=2.56 $Y=2.905 $X2=0 $Y2=0
cc_146 N_A_95_306#_M1014_d N_B2_c_333_n 0.00286492f $X=4.1 $Y=1.96 $X2=0 $Y2=0
cc_147 N_A_95_306#_c_146_n N_B2_c_327_n 0.0134773f $X=5.725 $Y=1.145 $X2=0 $Y2=0
cc_148 N_A_95_306#_c_146_n N_B2_c_328_n 0.0337589f $X=5.725 $Y=1.145 $X2=0 $Y2=0
cc_149 N_A_95_306#_c_141_n N_B2_c_329_n 0.0205422f $X=2.56 $Y=1.68 $X2=0 $Y2=0
cc_150 N_A_95_306#_c_158_n N_B2_c_329_n 0.00342481f $X=2.56 $Y=2.905 $X2=0 $Y2=0
cc_151 N_A_95_306#_c_142_n N_B2_c_329_n 2.0818e-19 $X=2.555 $Y=1.515 $X2=0 $Y2=0
cc_152 N_A_95_306#_c_143_n N_B2_c_329_n 0.0221918f $X=3.63 $Y=1.132 $X2=0 $Y2=0
cc_153 N_A_95_306#_M1009_d N_B2_c_359_n 7.30474e-19 $X=3.2 $Y=1.96 $X2=0 $Y2=0
cc_154 N_A_95_306#_M1009_d N_B2_c_336_n 0.00125583f $X=3.2 $Y=1.96 $X2=0 $Y2=0
cc_155 N_A_95_306#_c_143_n N_B2_c_336_n 0.0103756f $X=3.63 $Y=1.132 $X2=0 $Y2=0
cc_156 N_A_95_306#_c_160_n N_B1_c_423_n 0.0112503f $X=4.25 $Y=2.78 $X2=-0.19
+ $Y2=-0.245
cc_157 N_A_95_306#_c_163_n N_B1_c_423_n 0.00392126f $X=3.515 $Y=2.867 $X2=-0.19
+ $Y2=-0.245
cc_158 N_A_95_306#_c_143_n N_B1_M1000_g 0.0077677f $X=3.63 $Y=1.132 $X2=0 $Y2=0
cc_159 N_A_95_306#_c_144_n N_B1_M1000_g 0.00306707f $X=3.96 $Y=1.132 $X2=0 $Y2=0
cc_160 N_A_95_306#_c_144_n N_B1_M1018_g 0.00347829f $X=3.96 $Y=1.132 $X2=0 $Y2=0
cc_161 N_A_95_306#_c_146_n N_B1_M1018_g 0.00900647f $X=5.725 $Y=1.145 $X2=0
+ $Y2=0
cc_162 N_A_95_306#_c_160_n N_B1_c_424_n 0.012279f $X=4.25 $Y=2.78 $X2=0 $Y2=0
cc_163 N_A_95_306#_c_163_n N_B1_c_424_n 4.4235e-19 $X=3.515 $Y=2.867 $X2=0 $Y2=0
cc_164 N_A_95_306#_c_143_n B1 0.0246846f $X=3.63 $Y=1.132 $X2=0 $Y2=0
cc_165 N_A_95_306#_c_143_n N_B1_c_422_n 3.7993e-19 $X=3.63 $Y=1.132 $X2=0 $Y2=0
cc_166 N_A_95_306#_c_144_n N_B1_c_422_n 0.0011658f $X=3.96 $Y=1.132 $X2=0 $Y2=0
cc_167 N_A_95_306#_c_146_n N_B1_c_422_n 7.55386e-19 $X=5.725 $Y=1.145 $X2=0
+ $Y2=0
cc_168 N_A_95_306#_c_145_n N_A1_M1003_g 0.00290472f $X=5.89 $Y=1.105 $X2=0 $Y2=0
cc_169 N_A_95_306#_c_146_n N_A1_M1003_g 0.00778018f $X=5.725 $Y=1.145 $X2=0
+ $Y2=0
cc_170 N_A_95_306#_c_145_n N_A1_M1016_g 0.00358331f $X=5.89 $Y=1.105 $X2=0 $Y2=0
cc_171 N_A_95_306#_c_145_n A1 0.0248801f $X=5.89 $Y=1.105 $X2=0 $Y2=0
cc_172 N_A_95_306#_c_146_n A1 0.0225843f $X=5.725 $Y=1.145 $X2=0 $Y2=0
cc_173 N_A_95_306#_c_145_n N_A1_c_476_n 0.00225781f $X=5.89 $Y=1.105 $X2=0 $Y2=0
cc_174 N_A_95_306#_c_146_n N_A1_c_476_n 0.00178691f $X=5.725 $Y=1.145 $X2=0
+ $Y2=0
cc_175 N_A_95_306#_c_145_n N_A2_M1001_g 4.29877e-19 $X=5.89 $Y=1.105 $X2=0 $Y2=0
cc_176 N_A_95_306#_c_146_n N_A2_M1001_g 0.0172761f $X=5.725 $Y=1.145 $X2=0 $Y2=0
cc_177 N_A_95_306#_c_146_n N_A2_c_532_n 0.0131284f $X=5.725 $Y=1.145 $X2=0 $Y2=0
cc_178 N_A_95_306#_c_146_n A2 0.0099843f $X=5.725 $Y=1.145 $X2=0 $Y2=0
cc_179 N_A_95_306#_c_146_n N_A2_c_534_n 5.55026e-19 $X=5.725 $Y=1.145 $X2=0
+ $Y2=0
cc_180 N_A_95_306#_c_147_n N_VPWR_c_595_n 0.0170804f $X=0.565 $Y=1.765 $X2=0
+ $Y2=0
cc_181 N_A_95_306#_c_149_n N_VPWR_c_595_n 6.54535e-19 $X=1.015 $Y=1.765 $X2=0
+ $Y2=0
cc_182 N_A_95_306#_c_147_n N_VPWR_c_596_n 6.81676e-19 $X=0.565 $Y=1.765 $X2=0
+ $Y2=0
cc_183 N_A_95_306#_c_149_n N_VPWR_c_596_n 0.016107f $X=1.015 $Y=1.765 $X2=0
+ $Y2=0
cc_184 N_A_95_306#_c_132_n N_VPWR_c_596_n 0.00483147f $X=1.28 $Y=1.605 $X2=0
+ $Y2=0
cc_185 N_A_95_306#_c_151_n N_VPWR_c_596_n 0.00718907f $X=1.465 $Y=1.765 $X2=0
+ $Y2=0
cc_186 N_A_95_306#_c_140_n N_VPWR_c_596_n 3.76561e-19 $X=1.015 $Y=1.605 $X2=0
+ $Y2=0
cc_187 N_A_95_306#_c_154_n N_VPWR_c_597_n 0.00904085f $X=1.915 $Y=1.765 $X2=0
+ $Y2=0
cc_188 N_A_95_306#_c_221_p N_VPWR_c_597_n 0.0205483f $X=2.475 $Y=1.515 $X2=0
+ $Y2=0
cc_189 N_A_95_306#_c_158_n N_VPWR_c_597_n 0.0817995f $X=2.56 $Y=2.905 $X2=0
+ $Y2=0
cc_190 N_A_95_306#_c_159_n N_VPWR_c_597_n 0.0147457f $X=2.645 $Y=2.99 $X2=0
+ $Y2=0
cc_191 N_A_95_306#_c_142_n N_VPWR_c_597_n 0.00675548f $X=2.555 $Y=1.515 $X2=0
+ $Y2=0
cc_192 N_A_95_306#_c_147_n N_VPWR_c_602_n 0.00413917f $X=0.565 $Y=1.765 $X2=0
+ $Y2=0
cc_193 N_A_95_306#_c_149_n N_VPWR_c_602_n 0.00413917f $X=1.015 $Y=1.765 $X2=0
+ $Y2=0
cc_194 N_A_95_306#_c_151_n N_VPWR_c_603_n 0.00445602f $X=1.465 $Y=1.765 $X2=0
+ $Y2=0
cc_195 N_A_95_306#_c_154_n N_VPWR_c_603_n 0.00445602f $X=1.915 $Y=1.765 $X2=0
+ $Y2=0
cc_196 N_A_95_306#_c_159_n N_VPWR_c_604_n 0.0121867f $X=2.645 $Y=2.99 $X2=0
+ $Y2=0
cc_197 N_A_95_306#_c_160_n N_VPWR_c_604_n 0.037076f $X=4.25 $Y=2.78 $X2=0 $Y2=0
cc_198 N_A_95_306#_c_162_n N_VPWR_c_604_n 0.0568899f $X=3.185 $Y=2.867 $X2=0
+ $Y2=0
cc_199 N_A_95_306#_c_147_n N_VPWR_c_593_n 0.00817726f $X=0.565 $Y=1.765 $X2=0
+ $Y2=0
cc_200 N_A_95_306#_c_149_n N_VPWR_c_593_n 0.00817726f $X=1.015 $Y=1.765 $X2=0
+ $Y2=0
cc_201 N_A_95_306#_c_151_n N_VPWR_c_593_n 0.00857589f $X=1.465 $Y=1.765 $X2=0
+ $Y2=0
cc_202 N_A_95_306#_c_154_n N_VPWR_c_593_n 0.00862391f $X=1.915 $Y=1.765 $X2=0
+ $Y2=0
cc_203 N_A_95_306#_c_159_n N_VPWR_c_593_n 0.00660921f $X=2.645 $Y=2.99 $X2=0
+ $Y2=0
cc_204 N_A_95_306#_c_160_n N_VPWR_c_593_n 0.0309707f $X=4.25 $Y=2.78 $X2=0 $Y2=0
cc_205 N_A_95_306#_c_162_n N_VPWR_c_593_n 0.0322058f $X=3.185 $Y=2.867 $X2=0
+ $Y2=0
cc_206 N_A_95_306#_c_147_n N_X_c_687_n 0.00666212f $X=0.565 $Y=1.765 $X2=0 $Y2=0
cc_207 N_A_95_306#_c_131_n N_X_c_687_n 0.00645686f $X=0.925 $Y=1.605 $X2=0 $Y2=0
cc_208 N_A_95_306#_c_149_n N_X_c_687_n 0.00475527f $X=1.015 $Y=1.765 $X2=0 $Y2=0
cc_209 N_A_95_306#_c_139_n N_X_c_687_n 0.00204495f $X=0.565 $Y=1.605 $X2=0 $Y2=0
cc_210 N_A_95_306#_c_140_n N_X_c_687_n 0.00110515f $X=1.015 $Y=1.605 $X2=0 $Y2=0
cc_211 N_A_95_306#_M1002_g N_X_c_682_n 0.00813435f $X=1.355 $Y=0.87 $X2=0 $Y2=0
cc_212 N_A_95_306#_c_135_n N_X_c_682_n 2.21462e-19 $X=1.555 $Y=1.605 $X2=0 $Y2=0
cc_213 N_A_95_306#_c_136_n N_X_c_682_n 3.97481e-19 $X=1.785 $Y=1.35 $X2=0 $Y2=0
cc_214 N_A_95_306#_c_149_n N_X_c_688_n 5.57044e-19 $X=1.015 $Y=1.765 $X2=0 $Y2=0
cc_215 N_A_95_306#_c_151_n N_X_c_688_n 0.0147312f $X=1.465 $Y=1.765 $X2=0 $Y2=0
cc_216 N_A_95_306#_c_134_n N_X_c_688_n 0.00469357f $X=1.71 $Y=1.605 $X2=0 $Y2=0
cc_217 N_A_95_306#_c_135_n N_X_c_688_n 0.00409733f $X=1.555 $Y=1.605 $X2=0 $Y2=0
cc_218 N_A_95_306#_c_154_n N_X_c_688_n 0.0158231f $X=1.915 $Y=1.765 $X2=0 $Y2=0
cc_219 N_A_95_306#_c_140_n N_X_c_688_n 2.56101e-19 $X=1.015 $Y=1.605 $X2=0 $Y2=0
cc_220 N_A_95_306#_c_221_p N_X_c_688_n 0.00231492f $X=2.475 $Y=1.515 $X2=0 $Y2=0
cc_221 N_A_95_306#_c_158_n N_X_c_688_n 0.00474642f $X=2.56 $Y=2.905 $X2=0 $Y2=0
cc_222 N_A_95_306#_c_142_n N_X_c_688_n 0.00743235f $X=2.555 $Y=1.515 $X2=0 $Y2=0
cc_223 N_A_95_306#_c_136_n N_X_c_706_n 0.00202331f $X=1.785 $Y=1.35 $X2=0 $Y2=0
cc_224 N_A_95_306#_c_137_n N_X_c_706_n 0.01168f $X=2.215 $Y=1.35 $X2=0 $Y2=0
cc_225 N_A_95_306#_c_221_p N_X_c_706_n 0.0299782f $X=2.475 $Y=1.515 $X2=0 $Y2=0
cc_226 N_A_95_306#_c_141_n N_X_c_706_n 0.00341346f $X=2.56 $Y=1.68 $X2=0 $Y2=0
cc_227 N_A_95_306#_c_142_n N_X_c_706_n 0.00580258f $X=2.555 $Y=1.515 $X2=0 $Y2=0
cc_228 N_A_95_306#_c_136_n N_X_c_683_n 6.0186e-19 $X=1.785 $Y=1.35 $X2=0 $Y2=0
cc_229 N_A_95_306#_c_137_n N_X_c_683_n 0.00736569f $X=2.215 $Y=1.35 $X2=0 $Y2=0
cc_230 N_A_95_306#_c_131_n N_X_c_684_n 0.00357743f $X=0.925 $Y=1.605 $X2=0 $Y2=0
cc_231 N_A_95_306#_c_132_n N_X_c_684_n 0.00662608f $X=1.28 $Y=1.605 $X2=0 $Y2=0
cc_232 N_A_95_306#_M1002_g N_X_c_684_n 0.0199862f $X=1.355 $Y=0.87 $X2=0 $Y2=0
cc_233 N_A_95_306#_c_135_n N_X_c_684_n 0.00513294f $X=1.555 $Y=1.605 $X2=0 $Y2=0
cc_234 N_A_95_306#_c_140_n N_X_c_684_n 0.0136613f $X=1.015 $Y=1.605 $X2=0 $Y2=0
cc_235 N_A_95_306#_M1002_g N_X_c_718_n 0.0105486f $X=1.355 $Y=0.87 $X2=0 $Y2=0
cc_236 N_A_95_306#_c_134_n N_X_c_718_n 0.00364852f $X=1.71 $Y=1.605 $X2=0 $Y2=0
cc_237 N_A_95_306#_c_135_n N_X_c_718_n 0.00880219f $X=1.555 $Y=1.605 $X2=0 $Y2=0
cc_238 N_A_95_306#_c_136_n N_X_c_718_n 0.0148936f $X=1.785 $Y=1.35 $X2=0 $Y2=0
cc_239 N_A_95_306#_c_137_n N_X_c_718_n 0.00103837f $X=2.215 $Y=1.35 $X2=0 $Y2=0
cc_240 N_A_95_306#_c_221_p N_X_c_718_n 0.025226f $X=2.475 $Y=1.515 $X2=0 $Y2=0
cc_241 N_A_95_306#_c_142_n N_X_c_718_n 0.0109931f $X=2.555 $Y=1.515 $X2=0 $Y2=0
cc_242 N_A_95_306#_c_131_n X 0.0110935f $X=0.925 $Y=1.605 $X2=0 $Y2=0
cc_243 N_A_95_306#_c_139_n N_X_c_686_n 0.00956398f $X=0.565 $Y=1.605 $X2=0 $Y2=0
cc_244 N_A_95_306#_c_162_n N_A_555_392#_M1009_s 0.00376506f $X=3.185 $Y=2.867
+ $X2=-0.19 $Y2=-0.245
cc_245 N_A_95_306#_c_160_n N_A_555_392#_M1010_s 0.00202102f $X=4.25 $Y=2.78
+ $X2=0 $Y2=0
cc_246 N_A_95_306#_c_141_n N_A_555_392#_c_749_n 0.0026803f $X=2.56 $Y=1.68 $X2=0
+ $Y2=0
cc_247 N_A_95_306#_c_158_n N_A_555_392#_c_749_n 0.0587927f $X=2.56 $Y=2.905
+ $X2=0 $Y2=0
cc_248 N_A_95_306#_c_143_n N_A_555_392#_c_749_n 0.00410878f $X=3.63 $Y=1.132
+ $X2=0 $Y2=0
cc_249 N_A_95_306#_M1009_d N_A_555_392#_c_763_n 0.0039169f $X=3.2 $Y=1.96 $X2=0
+ $Y2=0
cc_250 N_A_95_306#_M1014_d N_A_555_392#_c_763_n 0.00512165f $X=4.1 $Y=1.96 $X2=0
+ $Y2=0
cc_251 N_A_95_306#_c_162_n N_A_555_392#_c_763_n 0.0040366f $X=3.185 $Y=2.867
+ $X2=0 $Y2=0
cc_252 N_A_95_306#_c_163_n N_A_555_392#_c_763_n 0.0645696f $X=3.515 $Y=2.867
+ $X2=0 $Y2=0
cc_253 N_A_95_306#_c_146_n N_A_555_392#_c_750_n 0.00674632f $X=5.725 $Y=1.145
+ $X2=0 $Y2=0
cc_254 N_A_95_306#_c_162_n N_A_555_392#_c_768_n 0.012787f $X=3.185 $Y=2.867
+ $X2=0 $Y2=0
cc_255 N_A_95_306#_c_163_n N_A_555_392#_c_768_n 0.00512594f $X=3.515 $Y=2.867
+ $X2=0 $Y2=0
cc_256 N_A_95_306#_c_160_n N_A_555_392#_c_756_n 0.0226667f $X=4.25 $Y=2.78 $X2=0
+ $Y2=0
cc_257 N_A_95_306#_c_141_n N_VGND_M1020_s 8.59214e-19 $X=2.56 $Y=1.68 $X2=0
+ $Y2=0
cc_258 N_A_95_306#_c_143_n N_VGND_M1020_s 0.00172209f $X=3.63 $Y=1.132 $X2=0
+ $Y2=0
cc_259 N_A_95_306#_c_146_n N_VGND_M1023_d 0.0128721f $X=5.725 $Y=1.145 $X2=0
+ $Y2=0
cc_260 N_A_95_306#_M1002_g N_VGND_c_825_n 0.00564714f $X=1.355 $Y=0.87 $X2=0
+ $Y2=0
cc_261 N_A_95_306#_c_140_n N_VGND_c_825_n 8.79152e-19 $X=1.015 $Y=1.605 $X2=0
+ $Y2=0
cc_262 N_A_95_306#_M1002_g N_VGND_c_826_n 4.52371e-19 $X=1.355 $Y=0.87 $X2=0
+ $Y2=0
cc_263 N_A_95_306#_c_136_n N_VGND_c_826_n 0.00782105f $X=1.785 $Y=1.35 $X2=0
+ $Y2=0
cc_264 N_A_95_306#_c_137_n N_VGND_c_826_n 0.00159705f $X=2.215 $Y=1.35 $X2=0
+ $Y2=0
cc_265 N_A_95_306#_c_137_n N_VGND_c_827_n 4.76302e-19 $X=2.215 $Y=1.35 $X2=0
+ $Y2=0
cc_266 N_A_95_306#_c_138_n N_VGND_c_827_n 0.0105834f $X=2.645 $Y=1.35 $X2=0
+ $Y2=0
cc_267 N_A_95_306#_c_141_n N_VGND_c_827_n 0.00892131f $X=2.56 $Y=1.68 $X2=0
+ $Y2=0
cc_268 N_A_95_306#_c_143_n N_VGND_c_827_n 0.013225f $X=3.63 $Y=1.132 $X2=0 $Y2=0
cc_269 N_A_95_306#_c_146_n N_VGND_c_828_n 0.015373f $X=5.725 $Y=1.145 $X2=0
+ $Y2=0
cc_270 N_A_95_306#_M1002_g N_VGND_c_832_n 0.00467453f $X=1.355 $Y=0.87 $X2=0
+ $Y2=0
cc_271 N_A_95_306#_c_136_n N_VGND_c_832_n 0.00405273f $X=1.785 $Y=1.35 $X2=0
+ $Y2=0
cc_272 N_A_95_306#_c_137_n N_VGND_c_834_n 0.00467453f $X=2.215 $Y=1.35 $X2=0
+ $Y2=0
cc_273 N_A_95_306#_c_138_n N_VGND_c_834_n 0.00405273f $X=2.645 $Y=1.35 $X2=0
+ $Y2=0
cc_274 N_A_95_306#_M1002_g N_VGND_c_840_n 0.00505379f $X=1.355 $Y=0.87 $X2=0
+ $Y2=0
cc_275 N_A_95_306#_c_136_n N_VGND_c_840_n 0.00424518f $X=1.785 $Y=1.35 $X2=0
+ $Y2=0
cc_276 N_A_95_306#_c_137_n N_VGND_c_840_n 0.00505379f $X=2.215 $Y=1.35 $X2=0
+ $Y2=0
cc_277 N_A_95_306#_c_138_n N_VGND_c_840_n 0.00424518f $X=2.645 $Y=1.35 $X2=0
+ $Y2=0
cc_278 N_A_95_306#_c_143_n N_A_645_120#_M1021_s 0.00216063f $X=3.63 $Y=1.132
+ $X2=-0.19 $Y2=-0.245
cc_279 N_A_95_306#_c_146_n N_A_645_120#_M1018_s 0.00224844f $X=5.725 $Y=1.145
+ $X2=0 $Y2=0
cc_280 N_A_95_306#_c_146_n N_A_645_120#_c_913_n 0.0161813f $X=5.725 $Y=1.145
+ $X2=0 $Y2=0
cc_281 N_A_95_306#_M1000_d N_A_645_120#_c_914_n 0.00169898f $X=3.655 $Y=0.6
+ $X2=0 $Y2=0
cc_282 N_A_95_306#_c_143_n N_A_645_120#_c_914_n 0.0162287f $X=3.63 $Y=1.132
+ $X2=0 $Y2=0
cc_283 N_A_95_306#_c_144_n N_A_645_120#_c_914_n 0.0163695f $X=3.96 $Y=1.132
+ $X2=0 $Y2=0
cc_284 N_A_95_306#_c_146_n N_A_645_120#_c_914_n 0.00607509f $X=5.725 $Y=1.145
+ $X2=0 $Y2=0
cc_285 N_A_95_306#_c_146_n N_A_1064_123#_M1001_d 0.00210096f $X=5.725 $Y=1.145
+ $X2=-0.19 $Y2=-0.245
cc_286 N_A_95_306#_M1003_d N_A_1064_123#_c_933_n 0.00408194f $X=5.75 $Y=0.615
+ $X2=0 $Y2=0
cc_287 N_A_95_306#_c_145_n N_A_1064_123#_c_933_n 0.0158841f $X=5.89 $Y=1.105
+ $X2=0 $Y2=0
cc_288 N_A_95_306#_c_146_n N_A_1064_123#_c_933_n 0.0164704f $X=5.725 $Y=1.145
+ $X2=0 $Y2=0
cc_289 N_A_95_306#_c_145_n N_A_1064_123#_c_931_n 0.0106625f $X=5.89 $Y=1.105
+ $X2=0 $Y2=0
cc_290 N_B2_c_323_n N_B1_c_423_n 0.0346236f $X=3.125 $Y=1.885 $X2=-0.19
+ $Y2=-0.245
cc_291 N_B2_c_332_n N_B1_c_423_n 0.0010174f $X=3.24 $Y=1.935 $X2=-0.19
+ $Y2=-0.245
cc_292 N_B2_c_333_n N_B1_c_423_n 2.59595e-19 $X=4.11 $Y=1.935 $X2=-0.19
+ $Y2=-0.245
cc_293 N_B2_c_336_n N_B1_c_423_n 0.0123645f $X=4.025 $Y=2.042 $X2=-0.19
+ $Y2=-0.245
cc_294 N_B2_M1021_g N_B1_M1000_g 0.0291033f $X=3.15 $Y=0.92 $X2=0 $Y2=0
cc_295 N_B2_M1023_g N_B1_M1018_g 0.0246028f $X=4.485 $Y=0.935 $X2=0 $Y2=0
cc_296 N_B2_c_325_n N_B1_c_424_n 0.0344067f $X=4.475 $Y=1.885 $X2=0 $Y2=0
cc_297 N_B2_c_333_n N_B1_c_424_n 0.00529793f $X=4.11 $Y=1.935 $X2=0 $Y2=0
cc_298 N_B2_c_336_n N_B1_c_424_n 0.0073645f $X=4.025 $Y=2.042 $X2=0 $Y2=0
cc_299 N_B2_c_323_n B1 3.6348e-19 $X=3.125 $Y=1.885 $X2=0 $Y2=0
cc_300 N_B2_c_327_n B1 0.0226234f $X=4.195 $Y=1.605 $X2=0 $Y2=0
cc_301 N_B2_c_329_n B1 0.0258902f $X=3.24 $Y=1.6 $X2=0 $Y2=0
cc_302 N_B2_c_336_n B1 0.0246438f $X=4.025 $Y=2.042 $X2=0 $Y2=0
cc_303 N_B2_c_323_n N_B1_c_422_n 0.0268045f $X=3.125 $Y=1.885 $X2=0 $Y2=0
cc_304 N_B2_c_325_n N_B1_c_422_n 0.0264761f $X=4.475 $Y=1.885 $X2=0 $Y2=0
cc_305 N_B2_M1023_g N_B1_c_422_n 2.32253e-19 $X=4.485 $Y=0.935 $X2=0 $Y2=0
cc_306 N_B2_c_332_n N_B1_c_422_n 0.00251579f $X=3.24 $Y=1.935 $X2=0 $Y2=0
cc_307 N_B2_c_333_n N_B1_c_422_n 0.00407615f $X=4.11 $Y=1.935 $X2=0 $Y2=0
cc_308 N_B2_c_327_n N_B1_c_422_n 0.0119783f $X=4.195 $Y=1.605 $X2=0 $Y2=0
cc_309 N_B2_c_329_n N_B1_c_422_n 0.00203145f $X=3.24 $Y=1.6 $X2=0 $Y2=0
cc_310 N_B2_c_336_n N_B1_c_422_n 0.00606449f $X=4.025 $Y=2.042 $X2=0 $Y2=0
cc_311 N_B2_c_325_n N_A2_c_526_n 0.00523896f $X=4.475 $Y=1.885 $X2=0 $Y2=0
cc_312 N_B2_c_325_n N_A2_c_536_n 0.00760542f $X=4.475 $Y=1.885 $X2=0 $Y2=0
cc_313 N_B2_M1023_g N_A2_M1001_g 0.0108695f $X=4.485 $Y=0.935 $X2=0 $Y2=0
cc_314 N_B2_c_325_n N_A2_c_532_n 0.0200398f $X=4.475 $Y=1.885 $X2=0 $Y2=0
cc_315 N_B2_M1023_g N_A2_c_532_n 0.00562171f $X=4.485 $Y=0.935 $X2=0 $Y2=0
cc_316 N_B2_c_328_n N_A2_c_532_n 0.00222306f $X=4.49 $Y=1.605 $X2=0 $Y2=0
cc_317 N_B2_M1023_g A2 3.85498e-19 $X=4.485 $Y=0.935 $X2=0 $Y2=0
cc_318 N_B2_M1023_g N_A2_c_534_n 4.96786e-19 $X=4.485 $Y=0.935 $X2=0 $Y2=0
cc_319 N_B2_c_323_n N_VPWR_c_604_n 0.00278271f $X=3.125 $Y=1.885 $X2=0 $Y2=0
cc_320 N_B2_c_325_n N_VPWR_c_604_n 0.00444483f $X=4.475 $Y=1.885 $X2=0 $Y2=0
cc_321 N_B2_c_323_n N_VPWR_c_593_n 0.00358708f $X=3.125 $Y=1.885 $X2=0 $Y2=0
cc_322 N_B2_c_325_n N_VPWR_c_593_n 0.00454867f $X=4.475 $Y=1.885 $X2=0 $Y2=0
cc_323 N_B2_c_336_n N_A_555_392#_M1010_s 0.00199645f $X=4.025 $Y=2.042 $X2=0
+ $Y2=0
cc_324 N_B2_c_323_n N_A_555_392#_c_749_n 0.00582136f $X=3.125 $Y=1.885 $X2=0
+ $Y2=0
cc_325 N_B2_c_359_n N_A_555_392#_c_749_n 0.0165318f $X=3.325 $Y=2.042 $X2=0
+ $Y2=0
cc_326 N_B2_c_323_n N_A_555_392#_c_763_n 0.0127027f $X=3.125 $Y=1.885 $X2=0
+ $Y2=0
cc_327 N_B2_c_325_n N_A_555_392#_c_763_n 0.0131928f $X=4.475 $Y=1.885 $X2=0
+ $Y2=0
cc_328 N_B2_c_333_n N_A_555_392#_c_763_n 0.00879415f $X=4.11 $Y=1.935 $X2=0
+ $Y2=0
cc_329 N_B2_c_328_n N_A_555_392#_c_763_n 0.0108057f $X=4.49 $Y=1.605 $X2=0 $Y2=0
cc_330 N_B2_c_329_n N_A_555_392#_c_763_n 0.00322388f $X=3.24 $Y=1.6 $X2=0 $Y2=0
cc_331 N_B2_c_359_n N_A_555_392#_c_763_n 0.00852115f $X=3.325 $Y=2.042 $X2=0
+ $Y2=0
cc_332 N_B2_c_336_n N_A_555_392#_c_763_n 0.0378665f $X=4.025 $Y=2.042 $X2=0
+ $Y2=0
cc_333 N_B2_c_325_n N_A_555_392#_c_750_n 0.00251422f $X=4.475 $Y=1.885 $X2=0
+ $Y2=0
cc_334 N_B2_c_333_n N_A_555_392#_c_750_n 0.00831476f $X=4.11 $Y=1.935 $X2=0
+ $Y2=0
cc_335 N_B2_c_328_n N_A_555_392#_c_750_n 0.00337333f $X=4.49 $Y=1.605 $X2=0
+ $Y2=0
cc_336 N_B2_c_333_n N_A_555_392#_c_784_n 0.00126147f $X=4.11 $Y=1.935 $X2=0
+ $Y2=0
cc_337 N_B2_c_323_n N_A_555_392#_c_768_n 4.48201e-19 $X=3.125 $Y=1.885 $X2=0
+ $Y2=0
cc_338 N_B2_c_325_n N_A_555_392#_c_756_n 0.00481991f $X=4.475 $Y=1.885 $X2=0
+ $Y2=0
cc_339 N_B2_M1021_g N_VGND_c_827_n 0.00499212f $X=3.15 $Y=0.92 $X2=0 $Y2=0
cc_340 N_B2_M1023_g N_VGND_c_828_n 0.008067f $X=4.485 $Y=0.935 $X2=0 $Y2=0
cc_341 N_B2_M1021_g N_VGND_c_839_n 0.00411835f $X=3.15 $Y=0.92 $X2=0 $Y2=0
cc_342 N_B2_M1023_g N_VGND_c_839_n 0.00349617f $X=4.485 $Y=0.935 $X2=0 $Y2=0
cc_343 N_B2_M1021_g N_VGND_c_840_n 0.00476395f $X=3.15 $Y=0.92 $X2=0 $Y2=0
cc_344 N_B2_M1023_g N_VGND_c_840_n 0.00396651f $X=4.485 $Y=0.935 $X2=0 $Y2=0
cc_345 N_B2_M1023_g N_A_645_120#_c_913_n 2.97537e-19 $X=4.485 $Y=0.935 $X2=0
+ $Y2=0
cc_346 N_B2_M1021_g N_A_645_120#_c_914_n 0.00359638f $X=3.15 $Y=0.92 $X2=0 $Y2=0
cc_347 N_B1_c_423_n N_VPWR_c_604_n 0.00290311f $X=3.575 $Y=1.885 $X2=0 $Y2=0
cc_348 N_B1_c_424_n N_VPWR_c_604_n 0.00291649f $X=4.025 $Y=1.885 $X2=0 $Y2=0
cc_349 N_B1_c_423_n N_VPWR_c_593_n 0.0035903f $X=3.575 $Y=1.885 $X2=0 $Y2=0
cc_350 N_B1_c_424_n N_VPWR_c_593_n 0.00359599f $X=4.025 $Y=1.885 $X2=0 $Y2=0
cc_351 N_B1_c_423_n N_A_555_392#_c_763_n 0.00850597f $X=3.575 $Y=1.885 $X2=0
+ $Y2=0
cc_352 N_B1_c_424_n N_A_555_392#_c_763_n 0.00848923f $X=4.025 $Y=1.885 $X2=0
+ $Y2=0
cc_353 N_B1_M1018_g N_VGND_c_828_n 9.3562e-19 $X=4.01 $Y=0.92 $X2=0 $Y2=0
cc_354 N_B1_M1000_g N_VGND_c_839_n 0.00327294f $X=3.58 $Y=0.92 $X2=0 $Y2=0
cc_355 N_B1_M1018_g N_VGND_c_839_n 0.00327294f $X=4.01 $Y=0.92 $X2=0 $Y2=0
cc_356 N_B1_M1000_g N_VGND_c_840_n 0.00476395f $X=3.58 $Y=0.92 $X2=0 $Y2=0
cc_357 N_B1_M1018_g N_VGND_c_840_n 0.00476395f $X=4.01 $Y=0.92 $X2=0 $Y2=0
cc_358 N_B1_M1000_g N_A_645_120#_c_914_n 0.0114295f $X=3.58 $Y=0.92 $X2=0 $Y2=0
cc_359 N_B1_M1018_g N_A_645_120#_c_914_n 0.0114847f $X=4.01 $Y=0.92 $X2=0 $Y2=0
cc_360 A1 N_A2_c_526_n 0.00707418f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_361 N_A1_c_476_n N_A2_c_526_n 0.00916309f $X=6.07 $Y=1.667 $X2=0 $Y2=0
cc_362 N_A1_c_477_n N_A2_c_536_n 0.0192726f $X=5.62 $Y=1.885 $X2=0 $Y2=0
cc_363 N_A1_M1003_g N_A2_c_528_n 0.00985192f $X=5.675 $Y=0.935 $X2=0 $Y2=0
cc_364 N_A1_M1016_g N_A2_c_528_n 0.00985192f $X=6.105 $Y=0.935 $X2=0 $Y2=0
cc_365 N_A1_M1016_g N_A2_c_529_n 0.0130116f $X=6.105 $Y=0.935 $X2=0 $Y2=0
cc_366 A1 N_A2_c_530_n 0.00184168f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_367 N_A1_c_476_n N_A2_c_530_n 0.0186513f $X=6.07 $Y=1.667 $X2=0 $Y2=0
cc_368 N_A1_c_478_n N_A2_c_538_n 0.0197812f $X=6.07 $Y=1.885 $X2=0 $Y2=0
cc_369 N_A1_M1016_g N_A2_M1022_g 0.00918444f $X=6.105 $Y=0.935 $X2=0 $Y2=0
cc_370 A1 N_A2_c_532_n 8.81484e-19 $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_371 N_A1_c_476_n N_A2_c_532_n 0.00192331f $X=6.07 $Y=1.667 $X2=0 $Y2=0
cc_372 N_A1_M1003_g N_A2_c_534_n 0.0301212f $X=5.675 $Y=0.935 $X2=0 $Y2=0
cc_373 N_A1_c_477_n N_VPWR_c_598_n 0.00709964f $X=5.62 $Y=1.885 $X2=0 $Y2=0
cc_374 N_A1_c_477_n N_VPWR_c_599_n 5.51351e-19 $X=5.62 $Y=1.885 $X2=0 $Y2=0
cc_375 N_A1_c_478_n N_VPWR_c_599_n 0.0116936f $X=6.07 $Y=1.885 $X2=0 $Y2=0
cc_376 N_A1_c_477_n N_VPWR_c_600_n 0.00445602f $X=5.62 $Y=1.885 $X2=0 $Y2=0
cc_377 N_A1_c_478_n N_VPWR_c_600_n 0.00413917f $X=6.07 $Y=1.885 $X2=0 $Y2=0
cc_378 N_A1_c_477_n N_VPWR_c_593_n 0.00858604f $X=5.62 $Y=1.885 $X2=0 $Y2=0
cc_379 N_A1_c_478_n N_VPWR_c_593_n 0.00817726f $X=6.07 $Y=1.885 $X2=0 $Y2=0
cc_380 N_A1_c_477_n N_A_555_392#_c_751_n 0.0128815f $X=5.62 $Y=1.885 $X2=0 $Y2=0
cc_381 A1 N_A_555_392#_c_751_n 0.0206447f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_382 N_A1_c_476_n N_A_555_392#_c_751_n 4.03117e-19 $X=6.07 $Y=1.667 $X2=0
+ $Y2=0
cc_383 N_A1_c_477_n N_A_555_392#_c_752_n 0.0104895f $X=5.62 $Y=1.885 $X2=0 $Y2=0
cc_384 N_A1_c_478_n N_A_555_392#_c_752_n 0.00605728f $X=6.07 $Y=1.885 $X2=0
+ $Y2=0
cc_385 N_A1_c_478_n N_A_555_392#_c_753_n 0.0136663f $X=6.07 $Y=1.885 $X2=0 $Y2=0
cc_386 A1 N_A_555_392#_c_753_n 0.0134169f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_387 N_A1_c_476_n N_A_555_392#_c_753_n 0.00325188f $X=6.07 $Y=1.667 $X2=0
+ $Y2=0
cc_388 N_A1_c_477_n N_A_555_392#_c_757_n 5.56417e-19 $X=5.62 $Y=1.885 $X2=0
+ $Y2=0
cc_389 A1 N_A_555_392#_c_757_n 0.0210155f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_390 N_A1_c_476_n N_A_555_392#_c_757_n 0.00610137f $X=6.07 $Y=1.667 $X2=0
+ $Y2=0
cc_391 N_A1_M1016_g N_VGND_c_829_n 5.60436e-19 $X=6.105 $Y=0.935 $X2=0 $Y2=0
cc_392 N_A1_M1003_g N_VGND_c_840_n 9.15321e-19 $X=5.675 $Y=0.935 $X2=0 $Y2=0
cc_393 N_A1_M1016_g N_VGND_c_840_n 9.15321e-19 $X=6.105 $Y=0.935 $X2=0 $Y2=0
cc_394 N_A1_M1003_g N_A_1064_123#_c_933_n 0.00924024f $X=5.675 $Y=0.935 $X2=0
+ $Y2=0
cc_395 N_A1_M1016_g N_A_1064_123#_c_933_n 0.0116768f $X=6.105 $Y=0.935 $X2=0
+ $Y2=0
cc_396 A1 N_A_1064_123#_c_933_n 0.00149839f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_397 N_A1_M1016_g N_A_1064_123#_c_930_n 4.59247e-19 $X=6.105 $Y=0.935 $X2=0
+ $Y2=0
cc_398 N_A2_c_536_n N_VPWR_c_598_n 0.0091384f $X=4.955 $Y=1.885 $X2=0 $Y2=0
cc_399 N_A2_c_538_n N_VPWR_c_599_n 0.0146851f $X=6.52 $Y=1.885 $X2=0 $Y2=0
cc_400 N_A2_c_536_n N_VPWR_c_604_n 0.00461464f $X=4.955 $Y=1.885 $X2=0 $Y2=0
cc_401 N_A2_c_538_n N_VPWR_c_605_n 0.00413917f $X=6.52 $Y=1.885 $X2=0 $Y2=0
cc_402 N_A2_c_536_n N_VPWR_c_593_n 0.0090964f $X=4.955 $Y=1.885 $X2=0 $Y2=0
cc_403 N_A2_c_538_n N_VPWR_c_593_n 0.00821673f $X=6.52 $Y=1.885 $X2=0 $Y2=0
cc_404 N_A2_c_536_n N_A_555_392#_c_750_n 2.78055e-19 $X=4.955 $Y=1.885 $X2=0
+ $Y2=0
cc_405 N_A2_c_536_n N_A_555_392#_c_751_n 0.0197548f $X=4.955 $Y=1.885 $X2=0
+ $Y2=0
cc_406 N_A2_c_532_n N_A_555_392#_c_751_n 0.00766307f $X=5.245 $Y=1.405 $X2=0
+ $Y2=0
cc_407 N_A2_c_536_n N_A_555_392#_c_752_n 8.33866e-19 $X=4.955 $Y=1.885 $X2=0
+ $Y2=0
cc_408 N_A2_c_538_n N_A_555_392#_c_753_n 0.0184423f $X=6.52 $Y=1.885 $X2=0 $Y2=0
cc_409 N_A2_c_538_n N_A_555_392#_c_754_n 4.02768e-19 $X=6.52 $Y=1.885 $X2=0
+ $Y2=0
cc_410 N_A2_c_538_n N_A_555_392#_c_755_n 0.00634858f $X=6.52 $Y=1.885 $X2=0
+ $Y2=0
cc_411 A2 N_VGND_M1023_d 0.00292336f $X=4.955 $Y=0.47 $X2=0 $Y2=0
cc_412 N_A2_M1001_g N_VGND_c_828_n 0.00341364f $X=5.245 $Y=0.935 $X2=0 $Y2=0
cc_413 A2 N_VGND_c_828_n 0.0333508f $X=4.955 $Y=0.47 $X2=0 $Y2=0
cc_414 N_A2_c_534_n N_VGND_c_828_n 0.00545095f $X=5.155 $Y=0.2 $X2=0 $Y2=0
cc_415 N_A2_c_528_n N_VGND_c_829_n 0.00811888f $X=6.46 $Y=0.2 $X2=0 $Y2=0
cc_416 N_A2_M1022_g N_VGND_c_829_n 0.0259946f $X=6.535 $Y=0.935 $X2=0 $Y2=0
cc_417 A2 N_VGND_c_837_n 0.0236953f $X=4.955 $Y=0.47 $X2=0 $Y2=0
cc_418 N_A2_c_534_n N_VGND_c_837_n 0.0403962f $X=5.155 $Y=0.2 $X2=0 $Y2=0
cc_419 N_A2_c_528_n N_VGND_c_840_n 0.0406735f $X=6.46 $Y=0.2 $X2=0 $Y2=0
cc_420 A2 N_VGND_c_840_n 0.0124201f $X=4.955 $Y=0.47 $X2=0 $Y2=0
cc_421 N_A2_c_534_n N_VGND_c_840_n 0.0100036f $X=5.155 $Y=0.2 $X2=0 $Y2=0
cc_422 N_A2_M1001_g N_A_1064_123#_c_933_n 0.00393563f $X=5.245 $Y=0.935 $X2=0
+ $Y2=0
cc_423 N_A2_c_528_n N_A_1064_123#_c_933_n 0.00827463f $X=6.46 $Y=0.2 $X2=0 $Y2=0
cc_424 A2 N_A_1064_123#_c_933_n 0.00164856f $X=4.955 $Y=0.47 $X2=0 $Y2=0
cc_425 N_A2_c_528_n N_A_1064_123#_c_930_n 0.00275881f $X=6.46 $Y=0.2 $X2=0 $Y2=0
cc_426 N_VPWR_c_595_n N_X_c_687_n 0.0703751f $X=0.34 $Y=1.985 $X2=0 $Y2=0
cc_427 N_VPWR_c_596_n N_X_c_687_n 0.0740216f $X=1.24 $Y=1.985 $X2=0 $Y2=0
cc_428 N_VPWR_c_602_n N_X_c_687_n 0.00749631f $X=1.075 $Y=3.33 $X2=0 $Y2=0
cc_429 N_VPWR_c_593_n N_X_c_687_n 0.0062048f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_430 N_VPWR_c_596_n N_X_c_688_n 0.0778383f $X=1.24 $Y=1.985 $X2=0 $Y2=0
cc_431 N_VPWR_c_597_n N_X_c_688_n 0.0757973f $X=2.14 $Y=2.015 $X2=0 $Y2=0
cc_432 N_VPWR_c_603_n N_X_c_688_n 0.014552f $X=2.055 $Y=3.33 $X2=0 $Y2=0
cc_433 N_VPWR_c_593_n N_X_c_688_n 0.0119791f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_434 N_VPWR_c_596_n N_X_c_684_n 0.0214136f $X=1.24 $Y=1.985 $X2=0 $Y2=0
cc_435 N_VPWR_c_595_n N_X_c_686_n 0.0119353f $X=0.34 $Y=1.985 $X2=0 $Y2=0
cc_436 N_VPWR_c_593_n N_A_555_392#_c_763_n 0.00807103f $X=6.96 $Y=3.33 $X2=0
+ $Y2=0
cc_437 N_VPWR_M1006_d N_A_555_392#_c_751_n 0.00562682f $X=5.03 $Y=1.96 $X2=0
+ $Y2=0
cc_438 N_VPWR_c_598_n N_A_555_392#_c_751_n 0.0326248f $X=5.27 $Y=2.375 $X2=0
+ $Y2=0
cc_439 N_VPWR_c_598_n N_A_555_392#_c_752_n 0.0256472f $X=5.27 $Y=2.375 $X2=0
+ $Y2=0
cc_440 N_VPWR_c_599_n N_A_555_392#_c_752_n 0.0462948f $X=6.295 $Y=2.375 $X2=0
+ $Y2=0
cc_441 N_VPWR_c_600_n N_A_555_392#_c_752_n 0.0110241f $X=6.13 $Y=3.33 $X2=0
+ $Y2=0
cc_442 N_VPWR_c_593_n N_A_555_392#_c_752_n 0.00909194f $X=6.96 $Y=3.33 $X2=0
+ $Y2=0
cc_443 N_VPWR_M1011_d N_A_555_392#_c_753_n 0.00197722f $X=6.145 $Y=1.96 $X2=0
+ $Y2=0
cc_444 N_VPWR_c_599_n N_A_555_392#_c_753_n 0.0171814f $X=6.295 $Y=2.375 $X2=0
+ $Y2=0
cc_445 N_VPWR_c_599_n N_A_555_392#_c_755_n 0.0462948f $X=6.295 $Y=2.375 $X2=0
+ $Y2=0
cc_446 N_VPWR_c_605_n N_A_555_392#_c_755_n 0.011066f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_447 N_VPWR_c_593_n N_A_555_392#_c_755_n 0.00915947f $X=6.96 $Y=3.33 $X2=0
+ $Y2=0
cc_448 N_VPWR_c_598_n N_A_555_392#_c_756_n 0.00159314f $X=5.27 $Y=2.375 $X2=0
+ $Y2=0
cc_449 N_VPWR_c_604_n N_A_555_392#_c_756_n 0.011066f $X=5.035 $Y=3.33 $X2=0
+ $Y2=0
cc_450 N_VPWR_c_593_n N_A_555_392#_c_756_n 0.00915947f $X=6.96 $Y=3.33 $X2=0
+ $Y2=0
cc_451 N_X_c_684_n N_VGND_M1002_s 0.00275278f $X=1.405 $Y=1.33 $X2=-0.19
+ $Y2=-0.245
cc_452 N_X_c_706_n N_VGND_M1004_s 0.0044545f $X=2.265 $Y=1.095 $X2=0 $Y2=0
cc_453 N_X_c_682_n N_VGND_c_825_n 0.0175587f $X=1.57 $Y=0.645 $X2=0 $Y2=0
cc_454 N_X_c_684_n N_VGND_c_825_n 0.0218366f $X=1.405 $Y=1.33 $X2=0 $Y2=0
cc_455 N_X_c_682_n N_VGND_c_826_n 0.0130934f $X=1.57 $Y=0.645 $X2=0 $Y2=0
cc_456 N_X_c_683_n N_VGND_c_826_n 0.0130934f $X=2.43 $Y=0.645 $X2=0 $Y2=0
cc_457 N_X_c_718_n N_VGND_c_826_n 0.0154032f $X=1.855 $Y=1.33 $X2=0 $Y2=0
cc_458 N_X_c_683_n N_VGND_c_827_n 0.0166774f $X=2.43 $Y=0.645 $X2=0 $Y2=0
cc_459 N_X_c_682_n N_VGND_c_832_n 0.00704565f $X=1.57 $Y=0.645 $X2=0 $Y2=0
cc_460 N_X_c_683_n N_VGND_c_834_n 0.00718756f $X=2.43 $Y=0.645 $X2=0 $Y2=0
cc_461 N_X_c_682_n N_VGND_c_840_n 0.00830435f $X=1.57 $Y=0.645 $X2=0 $Y2=0
cc_462 N_X_c_683_n N_VGND_c_840_n 0.0083989f $X=2.43 $Y=0.645 $X2=0 $Y2=0
cc_463 N_A_555_392#_c_753_n N_VGND_c_829_n 0.00221723f $X=6.66 $Y=2.035 $X2=0
+ $Y2=0
cc_464 N_A_555_392#_c_754_n N_VGND_c_829_n 0.00898193f $X=6.785 $Y=2.12 $X2=0
+ $Y2=0
cc_465 N_A_555_392#_c_753_n N_A_1064_123#_c_931_n 0.00539705f $X=6.66 $Y=2.035
+ $X2=0 $Y2=0
cc_466 N_VGND_c_828_n N_A_645_120#_c_913_n 0.0133114f $X=4.7 $Y=0.76 $X2=0 $Y2=0
cc_467 N_VGND_c_827_n N_A_645_120#_c_914_n 0.0109419f $X=2.86 $Y=0.75 $X2=0
+ $Y2=0
cc_468 N_VGND_c_839_n N_A_645_120#_c_914_n 0.0238447f $X=4.535 $Y=0 $X2=0 $Y2=0
cc_469 N_VGND_c_840_n N_A_645_120#_c_914_n 0.0346781f $X=6.96 $Y=0 $X2=0 $Y2=0
cc_470 N_VGND_c_828_n N_A_1064_123#_c_933_n 0.00574236f $X=4.7 $Y=0.76 $X2=0
+ $Y2=0
cc_471 N_VGND_c_837_n N_A_1064_123#_c_933_n 0.0122684f $X=6.585 $Y=0 $X2=0 $Y2=0
cc_472 N_VGND_c_840_n N_A_1064_123#_c_933_n 0.0214259f $X=6.96 $Y=0 $X2=0 $Y2=0
cc_473 N_VGND_c_829_n N_A_1064_123#_c_930_n 0.0096909f $X=6.75 $Y=0.76 $X2=0
+ $Y2=0
cc_474 N_VGND_c_837_n N_A_1064_123#_c_930_n 0.00374365f $X=6.585 $Y=0 $X2=0
+ $Y2=0
cc_475 N_VGND_c_840_n N_A_1064_123#_c_930_n 0.00464028f $X=6.96 $Y=0 $X2=0 $Y2=0
cc_476 N_VGND_c_829_n N_A_1064_123#_c_931_n 0.0160983f $X=6.75 $Y=0.76 $X2=0
+ $Y2=0
