* File: sky130_fd_sc_ls__decap_4.pxi.spice
* Created: Fri Aug 28 13:11:35 2020
* 
x_PM_SKY130_FD_SC_LS__DECAP_4%VGND N_VGND_M1001_s N_VGND_M1000_g N_VGND_c_22_n
+ N_VGND_c_23_n N_VGND_c_24_n N_VGND_c_25_n N_VGND_c_26_n N_VGND_c_27_n
+ N_VGND_c_28_n VGND N_VGND_c_29_n N_VGND_c_30_n
+ PM_SKY130_FD_SC_LS__DECAP_4%VGND
x_PM_SKY130_FD_SC_LS__DECAP_4%VPWR N_VPWR_M1000_s N_VPWR_M1001_g N_VPWR_c_50_n
+ N_VPWR_c_54_n N_VPWR_c_55_n N_VPWR_c_51_n N_VPWR_c_52_n VPWR N_VPWR_c_57_n
+ N_VPWR_c_58_n N_VPWR_c_53_n PM_SKY130_FD_SC_LS__DECAP_4%VPWR
cc_1 VNB N_VGND_c_22_n 0.021048f $X=-0.19 $Y=-0.245 $X2=0.547 $Y2=0.085
cc_2 VNB N_VGND_c_23_n 0.0103014f $X=-0.19 $Y=-0.245 $X2=0.547 $Y2=0.408
cc_3 VNB N_VGND_c_24_n 0.00972132f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.42
cc_4 VNB N_VGND_c_25_n 0.0504669f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.42
cc_5 VNB N_VGND_c_26_n 0.0145229f $X=-0.19 $Y=-0.245 $X2=1.552 $Y2=0.085
cc_6 VNB N_VGND_c_27_n 0.0102976f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=0.55
cc_7 VNB N_VGND_c_28_n 7.08202e-19 $X=-0.19 $Y=-0.245 $X2=0.325 $Y2=0.55
cc_8 VNB N_VGND_c_29_n 0.0176931f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=0
cc_9 VNB N_VGND_c_30_n 0.13936f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=0
cc_10 VNB N_VPWR_c_50_n 0.122413f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=1.83
cc_11 VNB N_VPWR_c_51_n 0.00369168f $X=-0.19 $Y=-0.245 $X2=1.552 $Y2=0.085
cc_12 VNB N_VPWR_c_52_n 0.0665683f $X=-0.19 $Y=-0.245 $X2=1.552 $Y2=0.55
cc_13 VNB N_VPWR_c_53_n 0.0840719f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=0
cc_14 VPB N_VGND_M1000_g 0.0982527f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=2.46
cc_15 VPB N_VGND_c_25_n 0.0201326f $X=-0.19 $Y=1.66 $X2=0.69 $Y2=1.42
cc_16 VPB N_VPWR_c_54_n 0.0144452f $X=-0.19 $Y=1.66 $X2=0.547 $Y2=0.408
cc_17 VPB N_VPWR_c_55_n 0.00826885f $X=-0.19 $Y=1.66 $X2=0.73 $Y2=1.42
cc_18 VPB N_VPWR_c_51_n 0.00788492f $X=-0.19 $Y=1.66 $X2=1.552 $Y2=0.085
cc_19 VPB N_VPWR_c_57_n 0.0179171f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_20 VPB N_VPWR_c_58_n 0.0299848f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=0
cc_21 VPB N_VPWR_c_53_n 0.0552469f $X=-0.19 $Y=1.66 $X2=1.68 $Y2=0
cc_22 N_VGND_c_23_n N_VPWR_c_50_n 0.0220411f $X=0.547 $Y=0.408 $X2=0 $Y2=0
cc_23 N_VGND_c_24_n N_VPWR_c_50_n 0.0377444f $X=0.69 $Y=1.42 $X2=0 $Y2=0
cc_24 N_VGND_c_25_n N_VPWR_c_50_n 0.0280007f $X=0.69 $Y=1.42 $X2=0 $Y2=0
cc_25 N_VGND_c_27_n N_VPWR_c_50_n 0.0198293f $X=1.595 $Y=0.55 $X2=0 $Y2=0
cc_26 N_VGND_c_28_n N_VPWR_c_50_n 0.0226114f $X=0.325 $Y=0.55 $X2=0 $Y2=0
cc_27 N_VGND_c_29_n N_VPWR_c_50_n 0.0176625f $X=1.425 $Y=0 $X2=0 $Y2=0
cc_28 N_VGND_c_30_n N_VPWR_c_50_n 0.0344366f $X=1.68 $Y=0 $X2=0 $Y2=0
cc_29 N_VGND_M1000_g N_VPWR_c_55_n 0.0164803f $X=0.96 $Y=2.46 $X2=0 $Y2=0
cc_30 N_VGND_M1000_g N_VPWR_c_51_n 0.0931345f $X=0.96 $Y=2.46 $X2=0 $Y2=0
cc_31 N_VGND_c_24_n N_VPWR_c_51_n 0.0203862f $X=0.69 $Y=1.42 $X2=0 $Y2=0
cc_32 N_VGND_c_25_n N_VPWR_c_51_n 0.0106588f $X=0.69 $Y=1.42 $X2=0 $Y2=0
cc_33 N_VGND_M1000_g N_VPWR_c_52_n 0.0235629f $X=0.96 $Y=2.46 $X2=0 $Y2=0
cc_34 N_VGND_c_24_n N_VPWR_c_52_n 0.00912536f $X=0.69 $Y=1.42 $X2=0 $Y2=0
cc_35 N_VGND_c_25_n N_VPWR_c_52_n 0.0203515f $X=0.69 $Y=1.42 $X2=0 $Y2=0
cc_36 N_VGND_M1000_g N_VPWR_c_57_n 0.0176614f $X=0.96 $Y=2.46 $X2=0 $Y2=0
cc_37 N_VGND_M1000_g N_VPWR_c_58_n 0.0444836f $X=0.96 $Y=2.46 $X2=0 $Y2=0
cc_38 N_VGND_M1000_g N_VPWR_c_53_n 0.0346242f $X=0.96 $Y=2.46 $X2=0 $Y2=0
