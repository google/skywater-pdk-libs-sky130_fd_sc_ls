* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
X0 X a_187_338# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X1 a_187_338# a_29_392# VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X2 X a_187_338# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X3 a_864_123# A1 a_187_338# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X4 a_596_392# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 X a_187_338# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X6 VPWR A2 a_596_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 a_596_392# a_29_392# a_187_338# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 VGND a_29_392# a_187_338# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X9 a_187_338# A1 a_864_123# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X10 a_29_392# B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 VPWR a_187_338# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X12 VGND A2 a_864_123# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X13 VPWR a_187_338# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X14 VPWR A1 a_596_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 a_864_123# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X16 a_187_338# a_29_392# a_596_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X17 X a_187_338# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X18 a_596_392# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 a_29_392# B1_N VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X20 VGND a_187_338# X VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X21 VGND a_187_338# X VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
.ends
