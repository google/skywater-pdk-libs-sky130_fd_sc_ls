* NGSPICE file created from sky130_fd_sc_ls__o22a_2.ext - technology: sky130A

.subckt sky130_fd_sc_ls__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
M1000 VPWR a_82_48# X VPB phighvt w=1.12e+06u l=150000u
+  ad=1.3764e+12p pd=9.08e+06u as=3.36e+11p ps=2.84e+06u
M1001 a_383_384# B1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=3e+11p pd=2.6e+06u as=0p ps=0u
M1002 a_82_48# B1 a_307_74# VNB nshort w=740000u l=150000u
+  ad=2.294e+11p pd=2.1e+06u as=6.649e+11p ps=6.26e+06u
M1003 X a_82_48# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_82_48# B2 a_383_384# VPB phighvt w=1e+06u l=150000u
+  ad=3.6e+11p pd=2.72e+06u as=0p ps=0u
M1005 a_575_384# A2 a_82_48# VPB phighvt w=1e+06u l=150000u
+  ad=3.9e+11p pd=2.78e+06u as=0p ps=0u
M1006 X a_82_48# VGND VNB nshort w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=6.5575e+11p ps=6.24e+06u
M1007 a_307_74# A1 VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND a_82_48# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR A1 a_575_384# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND A2 a_307_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_307_74# B2 a_82_48# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

