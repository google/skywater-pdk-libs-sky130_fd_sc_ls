* NGSPICE file created from sky130_fd_sc_ls__o21bai_4.ext - technology: sky130A

.subckt sky130_fd_sc_ls__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
M1000 VPWR a_828_48# Y VPB phighvt w=1.12e+06u l=150000u
+  ad=1.5204e+12p pd=1.309e+07u as=1.3888e+12p ps=1.144e+07u
M1001 a_27_74# A2 VGND VNB nshort w=740000u l=150000u
+  ad=1.6132e+12p pd=1.472e+07u as=1.2473e+12p ps=1.099e+07u
M1002 Y a_828_48# a_27_74# VNB nshort w=740000u l=150000u
+  ad=4.662e+11p pd=4.22e+06u as=0p ps=0u
M1003 VGND A2 a_27_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND A1 a_27_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND B1_N a_828_48# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1006 Y A2 a_28_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=1.7248e+12p ps=1.428e+07u
M1007 VPWR B1_N a_828_48# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=2.52e+11p ps=2.28e+06u
M1008 a_27_74# a_828_48# Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_28_368# A2 Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_27_74# A2 VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR A1 a_28_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_28_368# A1 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_27_74# A1 VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_27_74# A1 VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y A2 a_28_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR A1 a_28_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 Y a_828_48# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND A1 a_27_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND A2 a_27_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_28_368# A2 Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_28_368# A1 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_828_48# B1_N VPWR VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 Y a_828_48# a_27_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_27_74# a_828_48# Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

