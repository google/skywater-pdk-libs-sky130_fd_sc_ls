* File: sky130_fd_sc_ls__nor4bb_2.pex.spice
* Created: Wed Sep  2 11:16:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__NOR4BB_2%C_N 1 3 6 8 9 13
r33 15 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.03
+ $Y=1.635 $X2=1.03 $Y2=1.635
r34 13 15 22.788 $w=3.49e-07 $l=1.65e-07 $layer=POLY_cond $X=0.865 $Y=1.677
+ $X2=1.03 $Y2=1.677
r35 12 13 49.7192 $w=3.49e-07 $l=3.6e-07 $layer=POLY_cond $X=0.505 $Y=1.677
+ $X2=0.865 $Y2=1.677
r36 9 16 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=1.2 $Y=1.635 $X2=1.03
+ $Y2=1.635
r37 8 16 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=0.72 $Y=1.635 $X2=1.03
+ $Y2=1.635
r38 4 13 22.56 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.865 $Y=1.47
+ $X2=0.865 $Y2=1.677
r39 4 6 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=0.865 $Y=1.47
+ $X2=0.865 $Y2=0.69
r40 1 12 22.56 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.505 $Y=1.885
+ $X2=0.505 $Y2=1.677
r41 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.505 $Y=1.885
+ $X2=0.505 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_LS__NOR4BB_2%D_N 1 3 4 6 7 11
r36 11 13 22.0917 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=1.66 $Y=1.677
+ $X2=1.825 $Y2=1.677
r37 9 11 24.1 $w=3.6e-07 $l=1.8e-07 $layer=POLY_cond $X=1.48 $Y=1.677 $X2=1.66
+ $Y2=1.677
r38 7 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.66
+ $Y=1.635 $X2=1.66 $Y2=1.635
r39 4 13 23.3057 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.825 $Y=1.885
+ $X2=1.825 $Y2=1.677
r40 4 6 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.825 $Y=1.885
+ $X2=1.825 $Y2=2.46
r41 1 9 23.3057 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.48 $Y=1.47 $X2=1.48
+ $Y2=1.677
r42 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.48 $Y=1.47 $X2=1.48
+ $Y2=0.94
.ends

.subckt PM_SKY130_FD_SC_LS__NOR4BB_2%A_311_124# 1 2 7 9 12 16 18 20 21 27 33 37
+ 38 45 51
c75 16 0 1.04248e-19 $X=3.27 $Y=0.74
r76 51 52 1.94879 $w=3.71e-07 $l=1.5e-08 $layer=POLY_cond $X=3.27 $Y=1.557
+ $X2=3.285 $Y2=1.557
r77 48 49 0.649596 $w=3.71e-07 $l=5e-09 $layer=POLY_cond $X=2.835 $Y=1.557
+ $X2=2.84 $Y2=1.557
r78 45 48 12.3959 $w=3.71e-07 $l=1.08995e-07 $layer=POLY_cond $X=2.745 $Y=1.515
+ $X2=2.835 $Y2=1.557
r79 44 45 74.316 $w=3.3e-07 $l=4.25e-07 $layer=POLY_cond $X=2.32 $Y=1.515
+ $X2=2.745 $Y2=1.515
r80 43 44 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.32
+ $Y=1.515 $X2=2.32 $Y2=1.515
r81 37 39 0.877092 $w=4.38e-07 $l=5e-09 $layer=LI1_cond $X=2.105 $Y=2.135
+ $X2=2.105 $Y2=2.14
r82 37 38 8.83531 $w=4.38e-07 $l=1.65e-07 $layer=LI1_cond $X=2.105 $Y=2.135
+ $X2=2.105 $Y2=1.97
r83 34 51 35.0782 $w=3.71e-07 $l=2.7e-07 $layer=POLY_cond $X=3 $Y=1.557 $X2=3.27
+ $Y2=1.557
r84 34 49 20.7871 $w=3.71e-07 $l=1.6e-07 $layer=POLY_cond $X=3 $Y=1.557 $X2=2.84
+ $Y2=1.557
r85 33 43 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=3 $Y=1.515
+ $X2=2.325 $Y2=1.515
r86 33 34 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3
+ $Y=1.515 $X2=3 $Y2=1.515
r87 29 43 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.24 $Y=1.68
+ $X2=2.24 $Y2=1.515
r88 29 38 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=2.24 $Y=1.68
+ $X2=2.24 $Y2=1.97
r89 27 39 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.05 $Y=2.815
+ $X2=2.05 $Y2=2.14
r90 21 43 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.24 $Y=1.175
+ $X2=2.24 $Y2=1.515
r91 21 23 16.8257 $w=2.48e-07 $l=3.65e-07 $layer=LI1_cond $X=2.155 $Y=1.175
+ $X2=1.79 $Y2=1.175
r92 18 52 24.032 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.285 $Y=1.765
+ $X2=3.285 $Y2=1.557
r93 18 20 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.285 $Y=1.765
+ $X2=3.285 $Y2=2.4
r94 14 51 24.032 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.27 $Y=1.35
+ $X2=3.27 $Y2=1.557
r95 14 16 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.27 $Y=1.35
+ $X2=3.27 $Y2=0.74
r96 10 49 24.032 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.84 $Y=1.35
+ $X2=2.84 $Y2=1.557
r97 10 12 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.84 $Y=1.35
+ $X2=2.84 $Y2=0.74
r98 7 48 24.032 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.835 $Y=1.765
+ $X2=2.835 $Y2=1.557
r99 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.835 $Y=1.765
+ $X2=2.835 $Y2=2.4
r100 2 37 400 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=1 $X=1.9
+ $Y=1.96 $X2=2.05 $Y2=2.135
r101 2 27 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=1.9
+ $Y=1.96 $X2=2.05 $Y2=2.815
r102 1 23 182 $w=1.7e-07 $l=6.2149e-07 $layer=licon1_NDIFF $count=1 $X=1.555
+ $Y=0.62 $X2=1.79 $Y2=1.135
.ends

.subckt PM_SKY130_FD_SC_LS__NOR4BB_2%A_27_392# 1 2 7 9 12 14 16 19 25 27 29 30
+ 33 36 37 39 43 44 45 50 52 57
c137 19 0 3.67831e-20 $X=4.335 $Y=0.74
c138 14 0 1.13845e-19 $X=4.285 $Y=1.765
r139 57 58 6.69444 $w=3.6e-07 $l=5e-08 $layer=POLY_cond $X=4.285 $Y=1.557
+ $X2=4.335 $Y2=1.557
r140 56 57 50.8778 $w=3.6e-07 $l=3.8e-07 $layer=POLY_cond $X=3.905 $Y=1.557
+ $X2=4.285 $Y2=1.557
r141 55 56 16.0667 $w=3.6e-07 $l=1.2e-07 $layer=POLY_cond $X=3.785 $Y=1.557
+ $X2=3.905 $Y2=1.557
r142 51 55 0.669444 $w=3.6e-07 $l=5e-09 $layer=POLY_cond $X=3.78 $Y=1.557
+ $X2=3.785 $Y2=1.557
r143 50 52 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.78 $Y=1.515
+ $X2=3.78 $Y2=1.35
r144 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.78
+ $Y=1.515 $X2=3.78 $Y2=1.515
r145 45 47 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=2.58 $Y=0.795
+ $X2=2.58 $Y2=1.095
r146 41 52 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.7 $Y=1.18 $X2=3.7
+ $Y2=1.35
r147 40 47 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.665 $Y=1.095
+ $X2=2.58 $Y2=1.095
r148 39 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.615 $Y=1.095
+ $X2=3.7 $Y2=1.18
r149 39 40 61.9786 $w=1.68e-07 $l=9.5e-07 $layer=LI1_cond $X=3.615 $Y=1.095
+ $X2=2.665 $Y2=1.095
r150 38 44 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.815 $Y=0.795
+ $X2=0.65 $Y2=0.795
r151 37 45 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.495 $Y=0.795
+ $X2=2.58 $Y2=0.795
r152 37 38 109.604 $w=1.68e-07 $l=1.68e-06 $layer=LI1_cond $X=2.495 $Y=0.795
+ $X2=0.815 $Y2=0.795
r153 35 44 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.65 $Y=0.88
+ $X2=0.65 $Y2=0.795
r154 35 36 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=0.65 $Y=0.88
+ $X2=0.65 $Y2=1.13
r155 31 44 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.65 $Y=0.71
+ $X2=0.65 $Y2=0.795
r156 31 33 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=0.65 $Y=0.71
+ $X2=0.65 $Y2=0.525
r157 29 36 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.485 $Y=1.215
+ $X2=0.65 $Y2=1.13
r158 29 30 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=0.485 $Y=1.215
+ $X2=0.285 $Y2=1.215
r159 25 43 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.28 $Y=2.135
+ $X2=0.28 $Y2=1.97
r160 25 27 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.28 $Y=2.135
+ $X2=0.28 $Y2=2.815
r161 21 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.2 $Y=1.3
+ $X2=0.285 $Y2=1.215
r162 21 43 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.2 $Y=1.3 $X2=0.2
+ $Y2=1.97
r163 17 58 23.3057 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.335 $Y=1.35
+ $X2=4.335 $Y2=1.557
r164 17 19 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.335 $Y=1.35
+ $X2=4.335 $Y2=0.74
r165 14 57 23.3057 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=4.285 $Y=1.765
+ $X2=4.285 $Y2=1.557
r166 14 16 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.285 $Y=1.765
+ $X2=4.285 $Y2=2.4
r167 10 56 23.3057 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.905 $Y=1.35
+ $X2=3.905 $Y2=1.557
r168 10 12 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.905 $Y=1.35
+ $X2=3.905 $Y2=0.74
r169 7 55 23.3057 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.785 $Y=1.765
+ $X2=3.785 $Y2=1.557
r170 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.785 $Y=1.765
+ $X2=3.785 $Y2=2.4
r171 2 27 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.28 $Y2=2.815
r172 2 25 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.28 $Y2=2.135
r173 1 33 91 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=2 $X=0.505
+ $Y=0.37 $X2=0.65 $Y2=0.525
.ends

.subckt PM_SKY130_FD_SC_LS__NOR4BB_2%B 3 7 9 11 12 14 20 21 29 33
c59 21 0 1.27327e-19 $X=6 $Y=1.665
c60 3 0 1.75889e-19 $X=4.835 $Y=0.74
r61 29 31 14.3778 $w=3.52e-07 $l=1.05e-07 $layer=POLY_cond $X=5.64 $Y=1.557
+ $X2=5.745 $Y2=1.557
r62 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.64
+ $Y=1.515 $X2=5.64 $Y2=1.515
r63 27 29 47.2415 $w=3.52e-07 $l=3.45e-07 $layer=POLY_cond $X=5.295 $Y=1.557
+ $X2=5.64 $Y2=1.557
r64 26 27 4.10795 $w=3.52e-07 $l=3e-08 $layer=POLY_cond $X=5.265 $Y=1.557
+ $X2=5.295 $Y2=1.557
r65 21 30 9.64836 $w=4.28e-07 $l=3.6e-07 $layer=LI1_cond $X=6 $Y=1.565 $X2=5.64
+ $Y2=1.565
r66 20 30 3.21612 $w=4.28e-07 $l=1.2e-07 $layer=LI1_cond $X=5.52 $Y=1.565
+ $X2=5.64 $Y2=1.565
r67 20 33 4.39439 $w=4.28e-07 $l=1.15e-07 $layer=LI1_cond $X=5.52 $Y=1.565
+ $X2=5.405 $Y2=1.565
r68 18 26 32.8636 $w=3.52e-07 $l=2.4e-07 $layer=POLY_cond $X=5.025 $Y=1.557
+ $X2=5.265 $Y2=1.557
r69 18 24 26.017 $w=3.52e-07 $l=1.9e-07 $layer=POLY_cond $X=5.025 $Y=1.557
+ $X2=4.835 $Y2=1.557
r70 17 33 15.3659 $w=2.83e-07 $l=3.8e-07 $layer=LI1_cond $X=5.025 $Y=1.492
+ $X2=5.405 $Y2=1.492
r71 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.025
+ $Y=1.515 $X2=5.025 $Y2=1.515
r72 12 31 22.7654 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=5.745 $Y=1.765
+ $X2=5.745 $Y2=1.557
r73 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.745 $Y=1.765
+ $X2=5.745 $Y2=2.4
r74 9 27 22.7654 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=5.295 $Y=1.765
+ $X2=5.295 $Y2=1.557
r75 9 11 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.295 $Y=1.765
+ $X2=5.295 $Y2=2.4
r76 5 26 22.7654 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.265 $Y=1.35
+ $X2=5.265 $Y2=1.557
r77 5 7 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.265 $Y=1.35
+ $X2=5.265 $Y2=0.74
r78 1 24 22.7654 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.835 $Y=1.35
+ $X2=4.835 $Y2=1.557
r79 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.835 $Y=1.35
+ $X2=4.835 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__NOR4BB_2%A 3 5 7 8 10 13 15 16 22
c47 5 0 1.27327e-19 $X=6.245 $Y=1.765
r48 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.815
+ $Y=1.515 $X2=6.815 $Y2=1.515
r49 22 24 14.4469 $w=3.67e-07 $l=1.1e-07 $layer=POLY_cond $X=6.705 $Y=1.557
+ $X2=6.815 $Y2=1.557
r50 21 22 1.31335 $w=3.67e-07 $l=1e-08 $layer=POLY_cond $X=6.695 $Y=1.557
+ $X2=6.705 $Y2=1.557
r51 20 21 59.1008 $w=3.67e-07 $l=4.5e-07 $layer=POLY_cond $X=6.245 $Y=1.557
+ $X2=6.695 $Y2=1.557
r52 19 20 1.97003 $w=3.67e-07 $l=1.5e-08 $layer=POLY_cond $X=6.23 $Y=1.557
+ $X2=6.245 $Y2=1.557
r53 16 25 3.88615 $w=4.28e-07 $l=1.45e-07 $layer=LI1_cond $X=6.96 $Y=1.565
+ $X2=6.815 $Y2=1.565
r54 15 25 8.97834 $w=4.28e-07 $l=3.35e-07 $layer=LI1_cond $X=6.48 $Y=1.565
+ $X2=6.815 $Y2=1.565
r55 11 22 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.705 $Y=1.35
+ $X2=6.705 $Y2=1.557
r56 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.705 $Y=1.35
+ $X2=6.705 $Y2=0.74
r57 8 21 23.77 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=6.695 $Y=1.765
+ $X2=6.695 $Y2=1.557
r58 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.695 $Y=1.765
+ $X2=6.695 $Y2=2.4
r59 5 20 23.77 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=6.245 $Y=1.765
+ $X2=6.245 $Y2=1.557
r60 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.245 $Y=1.765
+ $X2=6.245 $Y2=2.4
r61 1 19 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.23 $Y=1.35 $X2=6.23
+ $Y2=1.557
r62 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.23 $Y=1.35 $X2=6.23
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__NOR4BB_2%VPWR 1 2 9 18 21 22 23 25 35 36 39
r59 40 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r60 39 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r61 39 40 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r62 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r63 33 36 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.96
+ $Y2=3.33
r64 32 33 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r65 30 39 17.0061 $w=1.7e-07 $l=5.5e-07 $layer=LI1_cond $X=1.715 $Y=3.33
+ $X2=1.165 $Y2=3.33
r66 30 32 279.556 $w=1.68e-07 $l=4.285e-06 $layer=LI1_cond $X=1.715 $Y=3.33
+ $X2=6 $Y2=3.33
r67 28 42 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r68 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r69 25 39 17.0061 $w=1.7e-07 $l=5.5e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=1.165 $Y2=3.33
r70 25 27 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.24 $Y2=3.33
r71 23 33 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=3.6 $Y=3.33 $X2=6
+ $Y2=3.33
r72 23 40 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=1.68 $Y2=3.33
r73 21 32 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=6.385 $Y=3.33 $X2=6
+ $Y2=3.33
r74 21 22 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.385 $Y=3.33
+ $X2=6.47 $Y2=3.33
r75 20 35 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=6.555 $Y=3.33
+ $X2=6.96 $Y2=3.33
r76 20 22 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.555 $Y=3.33
+ $X2=6.47 $Y2=3.33
r77 16 22 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.47 $Y=3.245
+ $X2=6.47 $Y2=3.33
r78 16 18 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=6.47 $Y=3.245
+ $X2=6.47 $Y2=2.455
r79 12 15 3.77091 $w=1.098e-06 $l=3.4e-07 $layer=LI1_cond $X=1.165 $Y=2.475
+ $X2=1.165 $Y2=2.815
r80 9 12 3.77091 $w=1.098e-06 $l=3.4e-07 $layer=LI1_cond $X=1.165 $Y=2.135
+ $X2=1.165 $Y2=2.475
r81 7 39 3.68071 $w=1.1e-06 $l=8.5e-08 $layer=LI1_cond $X=1.165 $Y=3.245
+ $X2=1.165 $Y2=3.33
r82 7 15 4.76909 $w=1.098e-06 $l=4.3e-07 $layer=LI1_cond $X=1.165 $Y=3.245
+ $X2=1.165 $Y2=2.815
r83 2 18 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=6.32
+ $Y=1.84 $X2=6.47 $Y2=2.455
r84 1 15 266.667 $w=1.7e-07 $l=1.10959e-06 $layer=licon1_PDIFF $count=2 $X=0.58
+ $Y=1.96 $X2=1.165 $Y2=2.815
r85 1 12 266.667 $w=1.7e-07 $l=1.25128e-06 $layer=licon1_PDIFF $count=2 $X=0.58
+ $Y=1.96 $X2=1.6 $Y2=2.475
r86 1 12 266.667 $w=1.7e-07 $l=5.85214e-07 $layer=licon1_PDIFF $count=2 $X=0.58
+ $Y=1.96 $X2=0.73 $Y2=2.475
r87 1 9 266.667 $w=1.7e-07 $l=6.66783e-07 $layer=licon1_PDIFF $count=2 $X=0.58
+ $Y=1.96 $X2=1.165 $Y2=2.135
.ends

.subckt PM_SKY130_FD_SC_LS__NOR4BB_2%A_493_368# 1 2 3 12 16 17 18 19 20 27
c43 16 0 1.13845e-19 $X=3.395 $Y=2.99
r44 21 25 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.725 $Y=2.275
+ $X2=3.56 $Y2=2.275
r45 20 27 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.345 $Y=2.275
+ $X2=4.51 $Y2=2.275
r46 20 21 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=4.345 $Y=2.275
+ $X2=3.725 $Y2=2.275
r47 18 25 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.56 $Y=2.36 $X2=3.56
+ $Y2=2.275
r48 18 19 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=3.56 $Y=2.36
+ $X2=3.56 $Y2=2.905
r49 16 19 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.395 $Y=2.99
+ $X2=3.56 $Y2=2.905
r50 16 17 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=3.395 $Y=2.99
+ $X2=2.775 $Y2=2.99
r51 12 15 32.9269 $w=2.78e-07 $l=8e-07 $layer=LI1_cond $X=2.635 $Y=2.015
+ $X2=2.635 $Y2=2.815
r52 10 17 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=2.635 $Y=2.905
+ $X2=2.775 $Y2=2.99
r53 10 15 3.70428 $w=2.78e-07 $l=9e-08 $layer=LI1_cond $X=2.635 $Y=2.905
+ $X2=2.635 $Y2=2.815
r54 3 27 300 $w=1.7e-07 $l=5.04455e-07 $layer=licon1_PDIFF $count=2 $X=4.36
+ $Y=1.84 $X2=4.51 $Y2=2.275
r55 2 25 300 $w=1.7e-07 $l=6.06815e-07 $layer=licon1_PDIFF $count=2 $X=3.36
+ $Y=1.84 $X2=3.56 $Y2=2.355
r56 1 15 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=2.465
+ $Y=1.84 $X2=2.61 $Y2=2.815
r57 1 12 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=2.465
+ $Y=1.84 $X2=2.61 $Y2=2.015
.ends

.subckt PM_SKY130_FD_SC_LS__NOR4BB_2%Y 1 2 3 4 5 18 20 23 25 26 30 32 36 39 44
+ 46 49 51 54 55
c116 49 0 1.04248e-19 $X=4.12 $Y=1.095
c117 46 0 1.75889e-19 $X=4.12 $Y=0.515
c118 18 0 3.67831e-20 $X=3.955 $Y=0.755
r119 51 55 13.7792 $w=2.28e-07 $l=2.75e-07 $layer=LI1_cond $X=4.285 $Y=1.665
+ $X2=4.56 $Y2=1.665
r120 51 52 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=4.2 $Y=1.665 $X2=4.2
+ $Y2=1.935
r121 46 48 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=4.12 $Y=0.515
+ $X2=4.12 $Y2=0.755
r122 39 41 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=3.055 $Y=0.675
+ $X2=3.055 $Y2=0.755
r123 34 36 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=6.45 $Y=1.01
+ $X2=6.45 $Y2=0.515
r124 33 54 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.215 $Y=1.095
+ $X2=5.09 $Y2=1.095
r125 32 34 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.325 $Y=1.095
+ $X2=6.45 $Y2=1.01
r126 32 33 72.4171 $w=1.68e-07 $l=1.11e-06 $layer=LI1_cond $X=6.325 $Y=1.095
+ $X2=5.215 $Y2=1.095
r127 28 54 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.09 $Y=1.01
+ $X2=5.09 $Y2=1.095
r128 28 30 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=5.09 $Y=1.01
+ $X2=5.09 $Y2=0.515
r129 27 49 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.285 $Y=1.095
+ $X2=4.12 $Y2=1.095
r130 26 54 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.965 $Y=1.095
+ $X2=5.09 $Y2=1.095
r131 26 27 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.965 $Y=1.095
+ $X2=4.285 $Y2=1.095
r132 25 51 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=4.2 $Y=1.55
+ $X2=4.2 $Y2=1.665
r133 24 49 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=4.2 $Y=1.18
+ $X2=4.12 $Y2=1.095
r134 24 25 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=4.2 $Y=1.18 $X2=4.2
+ $Y2=1.55
r135 23 49 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.12 $Y=1.01
+ $X2=4.12 $Y2=1.095
r136 22 48 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=4.12 $Y=0.84
+ $X2=4.12 $Y2=0.755
r137 22 23 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=4.12 $Y=0.84
+ $X2=4.12 $Y2=1.01
r138 21 44 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.225 $Y=1.935
+ $X2=3.1 $Y2=1.935
r139 20 52 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.115 $Y=1.935
+ $X2=4.2 $Y2=1.935
r140 20 21 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=4.115 $Y=1.935
+ $X2=3.225 $Y2=1.935
r141 19 41 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.22 $Y=0.755
+ $X2=3.055 $Y2=0.755
r142 18 48 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.955 $Y=0.755
+ $X2=4.12 $Y2=0.755
r143 18 19 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=3.955 $Y=0.755
+ $X2=3.22 $Y2=0.755
r144 5 44 300 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=2 $X=2.91
+ $Y=1.84 $X2=3.06 $Y2=2.015
r145 4 36 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=6.305
+ $Y=0.37 $X2=6.49 $Y2=0.515
r146 3 30 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.91
+ $Y=0.37 $X2=5.05 $Y2=0.515
r147 2 46 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.98
+ $Y=0.37 $X2=4.12 $Y2=0.515
r148 1 39 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=2.915
+ $Y=0.37 $X2=3.055 $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_LS__NOR4BB_2%A_772_368# 1 2 9 11 12 15
r27 13 15 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=5.52 $Y=2.905
+ $X2=5.52 $Y2=2.455
r28 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.355 $Y=2.99
+ $X2=5.52 $Y2=2.905
r29 11 12 76.984 $w=1.68e-07 $l=1.18e-06 $layer=LI1_cond $X=5.355 $Y=2.99
+ $X2=4.175 $Y2=2.99
r30 7 12 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=4.035 $Y=2.905
+ $X2=4.175 $Y2=2.99
r31 7 9 8.64332 $w=2.78e-07 $l=2.1e-07 $layer=LI1_cond $X=4.035 $Y=2.905
+ $X2=4.035 $Y2=2.695
r32 2 15 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=5.37
+ $Y=1.84 $X2=5.52 $Y2=2.455
r33 1 9 600 $w=1.7e-07 $l=9.4975e-07 $layer=licon1_PDIFF $count=1 $X=3.86
+ $Y=1.84 $X2=4.06 $Y2=2.695
.ends

.subckt PM_SKY130_FD_SC_LS__NOR4BB_2%A_985_368# 1 2 3 10 12 14 18 20 22 24 29
r45 22 31 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.92 $Y=2.12 $X2=6.92
+ $Y2=2.035
r46 22 24 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=6.92 $Y=2.12
+ $X2=6.92 $Y2=2.815
r47 21 29 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.185 $Y=2.035
+ $X2=6.02 $Y2=2.035
r48 20 31 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.755 $Y=2.035
+ $X2=6.92 $Y2=2.035
r49 20 21 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=6.755 $Y=2.035
+ $X2=6.185 $Y2=2.035
r50 16 29 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.02 $Y=2.12 $X2=6.02
+ $Y2=2.035
r51 16 18 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=6.02 $Y=2.12 $X2=6.02
+ $Y2=2.43
r52 15 27 3.99177 $w=1.7e-07 $l=1.5411e-07 $layer=LI1_cond $X=5.155 $Y=2.035
+ $X2=5.03 $Y2=1.97
r53 14 29 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.855 $Y=2.035
+ $X2=6.02 $Y2=2.035
r54 14 15 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=5.855 $Y=2.035
+ $X2=5.155 $Y2=2.035
r55 10 27 3.1514 $w=2.5e-07 $l=1.5e-07 $layer=LI1_cond $X=5.03 $Y=2.12 $X2=5.03
+ $Y2=1.97
r56 10 12 20.744 $w=2.48e-07 $l=4.5e-07 $layer=LI1_cond $X=5.03 $Y=2.12 $X2=5.03
+ $Y2=2.57
r57 3 31 400 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=6.77
+ $Y=1.84 $X2=6.92 $Y2=2.035
r58 3 24 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=6.77
+ $Y=1.84 $X2=6.92 $Y2=2.815
r59 2 29 600 $w=1.7e-07 $l=2.81069e-07 $layer=licon1_PDIFF $count=1 $X=5.82
+ $Y=1.84 $X2=6.02 $Y2=2.035
r60 2 18 300 $w=1.7e-07 $l=6.82715e-07 $layer=licon1_PDIFF $count=2 $X=5.82
+ $Y=1.84 $X2=6.02 $Y2=2.43
r61 1 27 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=4.925
+ $Y=1.84 $X2=5.07 $Y2=1.985
r62 1 12 600 $w=1.7e-07 $l=7.99218e-07 $layer=licon1_PDIFF $count=1 $X=4.925
+ $Y=1.84 $X2=5.07 $Y2=2.57
.ends

.subckt PM_SKY130_FD_SC_LS__NOR4BB_2%VGND 1 2 3 4 5 6 21 25 27 29 32 38 40 49 53
+ 58 63 76 79 83 92
r87 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r88 84 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r89 83 88 10.4851 $w=7.68e-07 $l=6.75e-07 $layer=LI1_cond $X=5.77 $Y=0 $X2=5.77
+ $Y2=0.675
r90 83 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r91 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r92 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r93 67 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6.96
+ $Y2=0
r94 67 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r95 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r96 64 83 9.95332 $w=1.7e-07 $l=3.85e-07 $layer=LI1_cond $X=6.155 $Y=0 $X2=5.77
+ $Y2=0
r97 64 66 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=6.155 $Y=0 $X2=6.48
+ $Y2=0
r98 63 91 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=6.755 $Y=0 $X2=6.977
+ $Y2=0
r99 63 66 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.755 $Y=0 $X2=6.48
+ $Y2=0
r100 62 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r101 62 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.56
+ $Y2=0
r102 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r103 59 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.785 $Y=0 $X2=4.62
+ $Y2=0
r104 59 61 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=4.785 $Y=0
+ $X2=5.04 $Y2=0
r105 58 83 9.95332 $w=1.7e-07 $l=3.85e-07 $layer=LI1_cond $X=5.385 $Y=0 $X2=5.77
+ $Y2=0
r106 58 61 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=5.385 $Y=0 $X2=5.04
+ $Y2=0
r107 57 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r108 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r109 54 76 9.39981 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=3.775 $Y=0
+ $X2=3.587 $Y2=0
r110 54 56 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.775 $Y=0
+ $X2=4.08 $Y2=0
r111 53 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.455 $Y=0 $X2=4.62
+ $Y2=0
r112 53 56 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=4.455 $Y=0
+ $X2=4.08 $Y2=0
r113 51 52 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r114 49 76 9.39981 $w=1.7e-07 $l=1.87e-07 $layer=LI1_cond $X=3.4 $Y=0 $X2=3.587
+ $Y2=0
r115 49 51 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=3.4 $Y=0 $X2=3.12
+ $Y2=0
r116 48 52 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r117 48 71 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.2
+ $Y2=0
r118 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r119 45 47 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=1.515 $Y=0
+ $X2=2.16 $Y2=0
r120 43 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r121 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r122 40 73 10.2521 $w=5.23e-07 $l=4.5e-07 $layer=LI1_cond $X=1.252 $Y=0
+ $X2=1.252 $Y2=0.45
r123 40 45 7.46409 $w=1.7e-07 $l=2.63e-07 $layer=LI1_cond $X=1.252 $Y=0
+ $X2=1.515 $Y2=0
r124 40 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r125 40 42 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.99 $Y=0 $X2=0.72
+ $Y2=0
r126 38 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r127 38 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r128 38 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r129 34 51 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=2.71 $Y=0 $X2=3.12
+ $Y2=0
r130 32 47 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=2.195 $Y=0 $X2=2.16
+ $Y2=0
r131 32 36 8.70931 $w=5.13e-07 $l=3.75e-07 $layer=LI1_cond $X=2.452 $Y=0
+ $X2=2.452 $Y2=0.375
r132 32 34 7.34265 $w=1.7e-07 $l=2.58e-07 $layer=LI1_cond $X=2.452 $Y=0 $X2=2.71
+ $Y2=0
r133 27 91 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=6.92 $Y=0.085
+ $X2=6.977 $Y2=0
r134 27 29 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=6.92 $Y=0.085
+ $X2=6.92 $Y2=0.515
r135 23 79 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.62 $Y=0.085
+ $X2=4.62 $Y2=0
r136 23 25 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=4.62 $Y=0.085
+ $X2=4.62 $Y2=0.675
r137 19 76 1.28102 $w=3.75e-07 $l=8.5e-08 $layer=LI1_cond $X=3.587 $Y=0.085
+ $X2=3.587 $Y2=0
r138 19 21 7.68295 $w=3.73e-07 $l=2.5e-07 $layer=LI1_cond $X=3.587 $Y=0.085
+ $X2=3.587 $Y2=0.335
r139 6 29 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.78
+ $Y=0.37 $X2=6.92 $Y2=0.515
r140 5 88 91 $w=1.7e-07 $l=8.13326e-07 $layer=licon1_NDIFF $count=2 $X=5.34
+ $Y=0.37 $X2=6.015 $Y2=0.675
r141 4 25 182 $w=1.7e-07 $l=3.96327e-07 $layer=licon1_NDIFF $count=1 $X=4.41
+ $Y=0.37 $X2=4.62 $Y2=0.675
r142 3 21 182 $w=1.7e-07 $l=2.56905e-07 $layer=licon1_NDIFF $count=1 $X=3.345
+ $Y=0.37 $X2=3.585 $Y2=0.335
r143 2 36 182 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_NDIFF $count=1 $X=2.215
+ $Y=0.23 $X2=2.45 $Y2=0.375
r144 1 73 182 $w=1.7e-07 $l=2.56905e-07 $layer=licon1_NDIFF $count=1 $X=0.94
+ $Y=0.37 $X2=1.16 $Y2=0.45
.ends

