* File: sky130_fd_sc_ls__or4_4.spice
* Created: Fri Aug 28 13:59:54 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__or4_4.pex.spice"
.subckt sky130_fd_sc_ls__or4_4  VNB VPB B A C D VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* D	D
* C	C
* A	A
* B	B
* VPB	VPB
* VNB	VNB
MM1000 N_VGND_M1000_d N_A_83_264#_M1000_g N_X_M1000_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2627 AS=0.1036 PD=2.19 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.3
+ SB=75005 A=0.111 P=1.78 MULT=1
MM1004 N_VGND_M1004_d N_A_83_264#_M1004_g N_X_M1000_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.7
+ SB=75004.6 A=0.111 P=1.78 MULT=1
MM1007 N_VGND_M1004_d N_A_83_264#_M1007_g N_X_M1007_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1295 AS=0.22385 PD=1.09 PS=1.345 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.2
+ SB=75004.1 A=0.111 P=1.78 MULT=1
MM1008 N_VGND_M1008_d N_A_83_264#_M1008_g N_X_M1007_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1835 AS=0.22385 PD=1.27 PS=1.345 NRD=16.212 NRS=41.34 M=1 R=4.93333
+ SA=75002 SB=75003.4 A=0.111 P=1.78 MULT=1
MM1003 N_A_83_264#_M1003_d N_B_M1003_g N_VGND_M1008_d VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1835 PD=1.02 PS=1.27 NRD=0 NRS=16.212 M=1 R=4.93333 SA=75002.6
+ SB=75002.7 A=0.111 P=1.78 MULT=1
MM1010 N_VGND_M1010_d N_A_M1010_g N_A_83_264#_M1003_d VNB NSHORT L=0.15 W=0.74
+ AD=0.5035 AS=0.1036 PD=2.07 PS=1.02 NRD=13.776 NRS=0 M=1 R=4.93333 SA=75003
+ SB=75002.3 A=0.111 P=1.78 MULT=1
MM1013 N_A_83_264#_M1013_d N_C_M1013_g N_VGND_M1010_d VNB NSHORT L=0.15 W=0.74
+ AD=0.1295 AS=0.5035 PD=1.09 PS=2.07 NRD=0 NRS=13.776 M=1 R=4.93333 SA=75004.4
+ SB=75000.9 A=0.111 P=1.78 MULT=1
MM1005 N_VGND_M1005_d N_D_M1005_g N_A_83_264#_M1013_d VNB NSHORT L=0.15 W=0.74
+ AD=0.3445 AS=0.1295 PD=3.08 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75004.9
+ SB=75000.4 A=0.111 P=1.78 MULT=1
MM1001 N_VPWR_M1001_d N_A_83_264#_M1001_g N_X_M1001_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1011 N_VPWR_M1011_d N_A_83_264#_M1011_g N_X_M1001_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1012 N_VPWR_M1011_d N_A_83_264#_M1012_g N_X_M1012_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1016 N_VPWR_M1016_d N_A_83_264#_M1016_g N_X_M1012_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.6 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1009 N_A_588_392#_M1009_d N_B_M1009_g N_A_499_392#_M1009_s VPB PHIGHVT L=0.15
+ W=1 AD=0.15 AS=0.295 PD=1.3 PS=2.59 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75003.5 A=0.15 P=2.3 MULT=1
MM1015 N_VPWR_M1015_d N_A_M1015_g N_A_588_392#_M1009_d VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75000.7
+ SB=75003.1 A=0.15 P=2.3 MULT=1
MM1018 N_VPWR_M1015_d N_A_M1018_g N_A_588_392#_M1018_s VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.16 PD=1.3 PS=1.32 NRD=1.9503 NRS=3.9203 M=1 R=6.66667 SA=75001.1
+ SB=75002.6 A=0.15 P=2.3 MULT=1
MM1014 N_A_588_392#_M1018_s N_B_M1014_g N_A_499_392#_M1014_s VPB PHIGHVT L=0.15
+ W=1 AD=0.16 AS=0.175 PD=1.32 PS=1.35 NRD=3.9203 NRS=11.8003 M=1 R=6.66667
+ SA=75001.6 SB=75002.2 A=0.15 P=2.3 MULT=1
MM1006 N_A_499_392#_M1014_s N_C_M1006_g N_A_962_392#_M1006_s VPB PHIGHVT L=0.15
+ W=1 AD=0.175 AS=0.175 PD=1.35 PS=1.35 NRD=1.9503 NRS=11.8003 M=1 R=6.66667
+ SA=75002.1 SB=75001.7 A=0.15 P=2.3 MULT=1
MM1002 N_A_962_392#_M1006_s N_D_M1002_g N_A_83_264#_M1002_s VPB PHIGHVT L=0.15
+ W=1 AD=0.175 AS=0.15 PD=1.35 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75002.6 SB=75001.2 A=0.15 P=2.3 MULT=1
MM1019 N_A_962_392#_M1019_d N_D_M1019_g N_A_83_264#_M1002_s VPB PHIGHVT L=0.15
+ W=1 AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75003
+ SB=75000.7 A=0.15 P=2.3 MULT=1
MM1017 N_A_499_392#_M1017_d N_C_M1017_g N_A_962_392#_M1019_d VPB PHIGHVT L=0.15
+ W=1 AD=0.345 AS=0.15 PD=2.69 PS=1.3 NRD=11.8003 NRS=1.9503 M=1 R=6.66667
+ SA=75003.5 SB=75000.3 A=0.15 P=2.3 MULT=1
DX20_noxref VNB VPB NWDIODE A=13.206 P=17.92
*
.include "sky130_fd_sc_ls__or4_4.pxi.spice"
*
.ends
*
*
