* File: sky130_fd_sc_ls__o21a_4.pex.spice
* Created: Wed Sep  2 11:18:06 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__O21A_4%A2 3 5 7 10 12 14 15 21 22
c52 21 0 1.27326e-19 $X=1.34 $Y=1.61
c53 3 0 1.92186e-19 $X=1 $Y=0.945
r54 22 23 3.23056 $w=3.73e-07 $l=2.5e-08 $layer=POLY_cond $X=1.43 $Y=1.652
+ $X2=1.455 $Y2=1.652
r55 20 22 11.63 $w=3.73e-07 $l=9e-08 $layer=POLY_cond $X=1.34 $Y=1.652 $X2=1.43
+ $Y2=1.652
r56 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.34
+ $Y=1.61 $X2=1.34 $Y2=1.61
r57 18 20 43.2895 $w=3.73e-07 $l=3.35e-07 $layer=POLY_cond $X=1.005 $Y=1.652
+ $X2=1.34 $Y2=1.652
r58 17 18 0.646113 $w=3.73e-07 $l=5e-09 $layer=POLY_cond $X=1 $Y=1.652 $X2=1.005
+ $Y2=1.652
r59 15 21 0.981855 $w=6.68e-07 $l=5.5e-08 $layer=LI1_cond $X=1.17 $Y=1.665
+ $X2=1.17 $Y2=1.61
r60 12 23 24.162 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.455 $Y=1.86
+ $X2=1.455 $Y2=1.652
r61 12 14 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.455 $Y=1.86
+ $X2=1.455 $Y2=2.435
r62 8 22 24.162 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.43 $Y=1.445
+ $X2=1.43 $Y2=1.652
r63 8 10 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=1.43 $Y=1.445 $X2=1.43
+ $Y2=0.945
r64 5 18 24.162 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.005 $Y=1.86
+ $X2=1.005 $Y2=1.652
r65 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.005 $Y=1.86
+ $X2=1.005 $Y2=2.435
r66 1 17 24.162 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1 $Y=1.445 $X2=1
+ $Y2=1.652
r67 1 3 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=1 $Y=1.445 $X2=1
+ $Y2=0.945
.ends

.subckt PM_SKY130_FD_SC_LS__O21A_4%A1 1 2 6 7 9 10 11 12 14 18 20
c65 7 0 1.27326e-19 $X=0.505 $Y=1.86
c66 1 0 1.85268e-19 $X=0.505 $Y=1.43
r67 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.96
+ $Y=1.61 $X2=1.96 $Y2=1.61
r68 20 24 6.88026 $w=3.33e-07 $l=2e-07 $layer=LI1_cond $X=2.16 $Y=1.612 $X2=1.96
+ $Y2=1.612
r69 16 23 38.5562 $w=2.99e-07 $l=1.88348e-07 $layer=POLY_cond $X=2.01 $Y=1.445
+ $X2=1.96 $Y2=1.61
r70 16 18 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=2.01 $Y=1.445 $X2=2.01
+ $Y2=0.945
r71 15 18 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.01 $Y=0.255
+ $X2=2.01 $Y2=0.945
r72 12 23 52.2586 $w=2.99e-07 $l=2.52488e-07 $layer=POLY_cond $X=1.955 $Y=1.86
+ $X2=1.96 $Y2=1.61
r73 12 14 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.955 $Y=1.86
+ $X2=1.955 $Y2=2.435
r74 10 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.935 $Y=0.18
+ $X2=2.01 $Y2=0.255
r75 10 11 699.926 $w=1.5e-07 $l=1.365e-06 $layer=POLY_cond $X=1.935 $Y=0.18
+ $X2=0.57 $Y2=0.18
r76 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.505 $Y=1.86
+ $X2=0.505 $Y2=2.435
r77 6 19 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.495 $Y=0.945
+ $X2=0.495 $Y2=1.34
r78 3 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.495 $Y=0.255
+ $X2=0.57 $Y2=0.18
r79 3 6 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.495 $Y=0.255
+ $X2=0.495 $Y2=0.945
r80 2 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.505 $Y=1.77 $X2=0.505
+ $Y2=1.86
r81 1 19 36.5962 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.505 $Y=1.43 $X2=0.505
+ $Y2=1.34
r82 1 2 132.161 $w=1.8e-07 $l=3.4e-07 $layer=POLY_cond $X=0.505 $Y=1.43
+ $X2=0.505 $Y2=1.77
.ends

.subckt PM_SKY130_FD_SC_LS__O21A_4%B1 3 5 7 10 12 14 15 16 23
c53 16 0 1.26926e-19 $X=3.12 $Y=1.665
c54 10 0 5.40193e-20 $X=2.87 $Y=0.945
c55 5 0 6.40318e-20 $X=2.495 $Y=1.86
c56 3 0 1.44963e-19 $X=2.44 $Y=0.945
r57 23 25 9.77027 $w=3.7e-07 $l=7.5e-08 $layer=POLY_cond $X=2.95 $Y=1.652
+ $X2=3.025 $Y2=1.652
r58 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.95
+ $Y=1.61 $X2=2.95 $Y2=1.61
r59 21 23 10.4216 $w=3.7e-07 $l=8e-08 $layer=POLY_cond $X=2.87 $Y=1.652 $X2=2.95
+ $Y2=1.652
r60 20 21 48.8514 $w=3.7e-07 $l=3.75e-07 $layer=POLY_cond $X=2.495 $Y=1.652
+ $X2=2.87 $Y2=1.652
r61 19 20 7.16487 $w=3.7e-07 $l=5.5e-08 $layer=POLY_cond $X=2.44 $Y=1.652
+ $X2=2.495 $Y2=1.652
r62 16 24 7.39303 $w=2.63e-07 $l=1.7e-07 $layer=LI1_cond $X=3.12 $Y=1.647
+ $X2=2.95 $Y2=1.647
r63 15 24 13.4814 $w=2.63e-07 $l=3.1e-07 $layer=LI1_cond $X=2.64 $Y=1.647
+ $X2=2.95 $Y2=1.647
r64 12 25 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.025 $Y=1.86
+ $X2=3.025 $Y2=1.652
r65 12 14 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=3.025 $Y=1.86
+ $X2=3.025 $Y2=2.355
r66 8 21 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.87 $Y=1.445
+ $X2=2.87 $Y2=1.652
r67 8 10 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=2.87 $Y=1.445 $X2=2.87
+ $Y2=0.945
r68 5 20 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.495 $Y=1.86
+ $X2=2.495 $Y2=1.652
r69 5 7 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.495 $Y=1.86
+ $X2=2.495 $Y2=2.355
r70 1 19 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.44 $Y=1.445
+ $X2=2.44 $Y2=1.652
r71 1 3 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=2.44 $Y=1.445 $X2=2.44
+ $Y2=0.945
.ends

.subckt PM_SKY130_FD_SC_LS__O21A_4%A_216_387# 1 2 3 10 12 13 15 16 18 19 21 22
+ 24 25 27 28 30 31 33 36 42 44 45 46 49 58 62 64 65 75
c142 75 0 1.26926e-19 $X=5.205 $Y=1.492
c143 64 0 6.40318e-20 $X=2.73 $Y=2.115
c144 42 0 1.44963e-19 $X=2.655 $Y=0.77
r145 75 76 6.61785 $w=4.37e-07 $l=6e-08 $layer=POLY_cond $X=5.205 $Y=1.492
+ $X2=5.265 $Y2=1.492
r146 74 75 40.8101 $w=4.37e-07 $l=3.7e-07 $layer=POLY_cond $X=4.835 $Y=1.492
+ $X2=5.205 $Y2=1.492
r147 73 74 8.8238 $w=4.37e-07 $l=8e-08 $layer=POLY_cond $X=4.755 $Y=1.492
+ $X2=4.835 $Y2=1.492
r148 70 71 18.1991 $w=4.37e-07 $l=1.65e-07 $layer=POLY_cond $X=4.205 $Y=1.492
+ $X2=4.37 $Y2=1.492
r149 67 68 20.405 $w=4.37e-07 $l=1.85e-07 $layer=POLY_cond $X=3.755 $Y=1.492
+ $X2=3.94 $Y2=1.492
r150 59 73 13.7872 $w=4.37e-07 $l=1.25e-07 $layer=POLY_cond $X=4.63 $Y=1.492
+ $X2=4.755 $Y2=1.492
r151 59 71 28.6773 $w=4.37e-07 $l=2.6e-07 $layer=POLY_cond $X=4.63 $Y=1.492
+ $X2=4.37 $Y2=1.492
r152 58 59 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=4.63
+ $Y=1.385 $X2=4.63 $Y2=1.385
r153 56 70 28.1259 $w=4.37e-07 $l=2.55e-07 $layer=POLY_cond $X=3.95 $Y=1.492
+ $X2=4.205 $Y2=1.492
r154 56 68 1.10297 $w=4.37e-07 $l=1e-08 $layer=POLY_cond $X=3.95 $Y=1.492
+ $X2=3.94 $Y2=1.492
r155 55 58 20.8976 $w=3.73e-07 $l=6.8e-07 $layer=LI1_cond $X=3.95 $Y=1.362
+ $X2=4.63 $Y2=1.362
r156 55 56 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.95
+ $Y=1.385 $X2=3.95 $Y2=1.385
r157 53 67 15.9931 $w=4.37e-07 $l=1.45e-07 $layer=POLY_cond $X=3.61 $Y=1.492
+ $X2=3.755 $Y2=1.492
r158 52 55 10.4488 $w=3.73e-07 $l=3.4e-07 $layer=LI1_cond $X=3.61 $Y=1.362
+ $X2=3.95 $Y2=1.362
r159 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.61
+ $Y=1.385 $X2=3.61 $Y2=1.385
r160 50 65 3.43356 $w=2.72e-07 $l=8.5e-08 $layer=LI1_cond $X=3.575 $Y=1.362
+ $X2=3.49 $Y2=1.362
r161 50 52 1.07561 $w=3.73e-07 $l=3.5e-08 $layer=LI1_cond $X=3.575 $Y=1.362
+ $X2=3.61 $Y2=1.362
r162 48 65 3.08518 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=3.49 $Y=1.55
+ $X2=3.49 $Y2=1.362
r163 48 49 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=3.49 $Y=1.55 $X2=3.49
+ $Y2=1.95
r164 47 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.895 $Y=2.035
+ $X2=2.73 $Y2=2.035
r165 46 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.405 $Y=2.035
+ $X2=3.49 $Y2=1.95
r166 46 47 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=3.405 $Y=2.035
+ $X2=2.895 $Y2=2.035
r167 44 65 3.43356 $w=2.72e-07 $l=1.38109e-07 $layer=LI1_cond $X=3.405 $Y=1.26
+ $X2=3.49 $Y2=1.362
r168 44 45 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=3.405 $Y=1.26
+ $X2=2.82 $Y2=1.26
r169 40 45 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.695 $Y=1.175
+ $X2=2.82 $Y2=1.26
r170 40 42 18.6696 $w=2.48e-07 $l=4.05e-07 $layer=LI1_cond $X=2.695 $Y=1.175
+ $X2=2.695 $Y2=0.77
r171 37 62 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.395 $Y=2.035
+ $X2=1.23 $Y2=2.035
r172 36 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.565 $Y=2.035
+ $X2=2.73 $Y2=2.035
r173 36 37 76.3316 $w=1.68e-07 $l=1.17e-06 $layer=LI1_cond $X=2.565 $Y=2.035
+ $X2=1.395 $Y2=2.035
r174 31 76 28.039 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=5.265 $Y=1.22
+ $X2=5.265 $Y2=1.492
r175 31 33 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.265 $Y=1.22
+ $X2=5.265 $Y2=0.74
r176 28 75 28.039 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=5.205 $Y=1.765
+ $X2=5.205 $Y2=1.492
r177 28 30 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.205 $Y=1.765
+ $X2=5.205 $Y2=2.4
r178 25 74 28.039 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=4.835 $Y=1.22
+ $X2=4.835 $Y2=1.492
r179 25 27 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.835 $Y=1.22
+ $X2=4.835 $Y2=0.74
r180 22 73 28.039 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=4.755 $Y=1.765
+ $X2=4.755 $Y2=1.492
r181 22 24 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.755 $Y=1.765
+ $X2=4.755 $Y2=2.4
r182 19 71 28.039 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=4.37 $Y=1.22
+ $X2=4.37 $Y2=1.492
r183 19 21 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.37 $Y=1.22
+ $X2=4.37 $Y2=0.74
r184 16 70 28.039 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=4.205 $Y=1.765
+ $X2=4.205 $Y2=1.492
r185 16 18 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.205 $Y=1.765
+ $X2=4.205 $Y2=2.4
r186 13 68 28.039 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=3.94 $Y=1.22
+ $X2=3.94 $Y2=1.492
r187 13 15 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.94 $Y=1.22
+ $X2=3.94 $Y2=0.74
r188 10 67 28.039 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=3.755 $Y=1.765
+ $X2=3.755 $Y2=1.492
r189 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.755 $Y=1.765
+ $X2=3.755 $Y2=2.4
r190 3 64 300 $w=1.7e-07 $l=2.47386e-07 $layer=licon1_PDIFF $count=2 $X=2.57
+ $Y=1.935 $X2=2.73 $Y2=2.115
r191 2 62 300 $w=1.7e-07 $l=2.43721e-07 $layer=licon1_PDIFF $count=2 $X=1.08
+ $Y=1.935 $X2=1.23 $Y2=2.115
r192 1 42 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.515
+ $Y=0.625 $X2=2.655 $Y2=0.77
.ends

.subckt PM_SKY130_FD_SC_LS__O21A_4%VPWR 1 2 3 4 5 16 18 24 28 32 36 38 43 44 45
+ 47 59 63 72 75 79
r70 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r71 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r72 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r73 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r74 67 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r75 67 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r76 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r77 64 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.645 $Y=3.33
+ $X2=4.48 $Y2=3.33
r78 64 66 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=4.645 $Y=3.33
+ $X2=5.04 $Y2=3.33
r79 63 78 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=5.315 $Y=3.33
+ $X2=5.537 $Y2=3.33
r80 63 66 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=5.315 $Y=3.33
+ $X2=5.04 $Y2=3.33
r81 62 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r82 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r83 59 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.315 $Y=3.33
+ $X2=4.48 $Y2=3.33
r84 59 61 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=4.315 $Y=3.33
+ $X2=4.08 $Y2=3.33
r85 58 62 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r86 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r87 55 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.395 $Y=3.33
+ $X2=2.23 $Y2=3.33
r88 55 57 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=2.395 $Y=3.33
+ $X2=3.12 $Y2=3.33
r89 54 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r90 53 54 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r91 51 54 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r92 51 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r93 50 53 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=3.33 $X2=1.68
+ $Y2=3.33
r94 50 51 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r95 48 69 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.222 $Y2=3.33
r96 48 50 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.72 $Y2=3.33
r97 47 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.065 $Y=3.33
+ $X2=2.23 $Y2=3.33
r98 47 53 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=2.065 $Y=3.33
+ $X2=1.68 $Y2=3.33
r99 45 58 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=3.12 $Y2=3.33
r100 45 73 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=2.16 $Y2=3.33
r101 43 57 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=3.135 $Y=3.33
+ $X2=3.12 $Y2=3.33
r102 43 44 11.015 $w=1.7e-07 $l=2.4e-07 $layer=LI1_cond $X=3.135 $Y=3.33
+ $X2=3.375 $Y2=3.33
r103 42 61 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=3.615 $Y=3.33
+ $X2=4.08 $Y2=3.33
r104 42 44 11.015 $w=1.7e-07 $l=2.4e-07 $layer=LI1_cond $X=3.615 $Y=3.33
+ $X2=3.375 $Y2=3.33
r105 38 41 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=5.48 $Y=2.115
+ $X2=5.48 $Y2=2.815
r106 36 78 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=5.48 $Y=3.245
+ $X2=5.537 $Y2=3.33
r107 36 41 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=5.48 $Y=3.245
+ $X2=5.48 $Y2=2.815
r108 32 35 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=4.48 $Y=2.145
+ $X2=4.48 $Y2=2.825
r109 30 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.48 $Y=3.245
+ $X2=4.48 $Y2=3.33
r110 30 35 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=4.48 $Y=3.245
+ $X2=4.48 $Y2=2.825
r111 26 44 1.96841 $w=4.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.375 $Y=3.245
+ $X2=3.375 $Y2=3.33
r112 26 28 19.4363 $w=4.78e-07 $l=7.8e-07 $layer=LI1_cond $X=3.375 $Y=3.245
+ $X2=3.375 $Y2=2.465
r113 22 72 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.23 $Y=3.245
+ $X2=2.23 $Y2=3.33
r114 22 24 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=2.23 $Y=3.245
+ $X2=2.23 $Y2=2.455
r115 18 21 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.28 $Y=2.08
+ $X2=0.28 $Y2=2.79
r116 16 69 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.222 $Y2=3.33
r117 16 21 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.28 $Y2=2.79
r118 5 41 400 $w=1.7e-07 $l=1.07034e-06 $layer=licon1_PDIFF $count=1 $X=5.28
+ $Y=1.84 $X2=5.48 $Y2=2.815
r119 5 38 400 $w=1.7e-07 $l=3.61421e-07 $layer=licon1_PDIFF $count=1 $X=5.28
+ $Y=1.84 $X2=5.48 $Y2=2.115
r120 4 35 400 $w=1.7e-07 $l=1.08038e-06 $layer=licon1_PDIFF $count=1 $X=4.28
+ $Y=1.84 $X2=4.48 $Y2=2.825
r121 4 32 400 $w=1.7e-07 $l=3.9246e-07 $layer=licon1_PDIFF $count=1 $X=4.28
+ $Y=1.84 $X2=4.48 $Y2=2.145
r122 3 28 600 $w=1.7e-07 $l=6.4707e-07 $layer=licon1_PDIFF $count=1 $X=3.1
+ $Y=1.935 $X2=3.36 $Y2=2.465
r123 2 24 600 $w=1.7e-07 $l=6.11882e-07 $layer=licon1_PDIFF $count=1 $X=2.03
+ $Y=1.935 $X2=2.23 $Y2=2.455
r124 1 21 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.935 $X2=0.28 $Y2=2.79
r125 1 18 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.935 $X2=0.28 $Y2=2.08
.ends

.subckt PM_SKY130_FD_SC_LS__O21A_4%A_116_387# 1 2 9 13 14 17
r21 15 17 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=1.73 $Y=2.905
+ $X2=1.73 $Y2=2.375
r22 13 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.565 $Y=2.99
+ $X2=1.73 $Y2=2.905
r23 13 14 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.565 $Y=2.99
+ $X2=0.865 $Y2=2.99
r24 9 12 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=0.74 $Y=2.115
+ $X2=0.74 $Y2=2.795
r25 7 14 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.74 $Y=2.905
+ $X2=0.865 $Y2=2.99
r26 7 12 5.07075 $w=2.48e-07 $l=1.1e-07 $layer=LI1_cond $X=0.74 $Y=2.905
+ $X2=0.74 $Y2=2.795
r27 2 17 300 $w=1.7e-07 $l=5.3066e-07 $layer=licon1_PDIFF $count=2 $X=1.53
+ $Y=1.935 $X2=1.73 $Y2=2.375
r28 1 12 400 $w=1.7e-07 $l=9.54777e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.935 $X2=0.78 $Y2=2.795
r29 1 9 400 $w=1.7e-07 $l=2.75681e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.935 $X2=0.78 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_LS__O21A_4%X 1 2 3 4 15 19 21 23 24 25 29 35 38 42 45
r70 41 45 18.7898 $w=2.28e-07 $l=3.75e-07 $layer=LI1_cond $X=5.145 $Y=1.665
+ $X2=5.52 $Y2=1.665
r71 41 42 3.75657 $w=2.3e-07 $l=3.56441e-07 $layer=LI1_cond $X=5.145 $Y=1.665
+ $X2=4.815 $Y2=1.72
r72 38 42 2.39845 $w=1.7e-07 $l=3.08504e-07 $layer=LI1_cond $X=5.05 $Y=1.55
+ $X2=4.815 $Y2=1.72
r73 37 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.05 $Y=1.005
+ $X2=5.05 $Y2=0.92
r74 37 38 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=5.05 $Y=1.005
+ $X2=5.05 $Y2=1.55
r75 33 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.05 $Y=0.835
+ $X2=5.05 $Y2=0.92
r76 33 35 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=5.05 $Y=0.835
+ $X2=5.05 $Y2=0.515
r77 29 31 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=4.98 $Y=1.985
+ $X2=4.98 $Y2=2.815
r78 27 42 2.39845 $w=3.3e-07 $l=2.38642e-07 $layer=LI1_cond $X=4.98 $Y=1.89
+ $X2=4.815 $Y2=1.72
r79 27 29 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=4.98 $Y=1.89
+ $X2=4.98 $Y2=1.985
r80 26 40 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.24 $Y=0.92
+ $X2=4.115 $Y2=0.92
r81 25 44 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.965 $Y=0.92
+ $X2=5.05 $Y2=0.92
r82 25 26 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=4.965 $Y=0.92
+ $X2=4.24 $Y2=0.92
r83 23 42 3.75657 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.815 $Y=1.805
+ $X2=4.815 $Y2=1.72
r84 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.815 $Y=1.805
+ $X2=4.145 $Y2=1.805
r85 19 40 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.115 $Y=0.835
+ $X2=4.115 $Y2=0.92
r86 19 21 15.6732 $w=2.48e-07 $l=3.4e-07 $layer=LI1_cond $X=4.115 $Y=0.835
+ $X2=4.115 $Y2=0.495
r87 15 17 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=3.98 $Y=1.985
+ $X2=3.98 $Y2=2.815
r88 13 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.98 $Y=1.89
+ $X2=4.145 $Y2=1.805
r89 13 15 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=3.98 $Y=1.89
+ $X2=3.98 $Y2=1.985
r90 4 31 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=4.83
+ $Y=1.84 $X2=4.98 $Y2=2.815
r91 4 29 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=4.83
+ $Y=1.84 $X2=4.98 $Y2=1.985
r92 3 17 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=3.83
+ $Y=1.84 $X2=3.98 $Y2=2.815
r93 3 15 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=3.83
+ $Y=1.84 $X2=3.98 $Y2=1.985
r94 2 44 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=4.91
+ $Y=0.37 $X2=5.05 $Y2=0.965
r95 2 35 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=4.91
+ $Y=0.37 $X2=5.05 $Y2=0.515
r96 1 40 182 $w=1.7e-07 $l=6.16036e-07 $layer=licon1_NDIFF $count=1 $X=4.015
+ $Y=0.37 $X2=4.155 $Y2=0.92
r97 1 21 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=4.015
+ $Y=0.37 $X2=4.155 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LS__O21A_4%A_27_125# 1 2 3 4 15 17 18 21 23 28 29 30 33
+ 35
c67 23 0 5.40193e-20 $X=2.06 $Y=1.19
c68 21 0 1.44963e-19 $X=1.215 $Y=0.77
c69 18 0 2.32491e-19 $X=0.445 $Y=1.19
r70 31 33 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.165 $Y=0.435
+ $X2=3.165 $Y2=0.805
r71 29 31 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3 $Y=0.35
+ $X2=3.165 $Y2=0.435
r72 29 30 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=3 $Y=0.35 $X2=2.39
+ $Y2=0.35
r73 26 28 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.225 $Y=1.105
+ $X2=2.225 $Y2=0.77
r74 25 30 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.225 $Y=0.435
+ $X2=2.39 $Y2=0.35
r75 25 28 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.225 $Y=0.435
+ $X2=2.225 $Y2=0.77
r76 24 35 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.38 $Y=1.19
+ $X2=1.255 $Y2=1.19
r77 23 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.06 $Y=1.19
+ $X2=2.225 $Y2=1.105
r78 23 24 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.06 $Y=1.19
+ $X2=1.38 $Y2=1.19
r79 19 35 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.255 $Y=1.105
+ $X2=1.255 $Y2=1.19
r80 19 21 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=1.255 $Y=1.105
+ $X2=1.255 $Y2=0.77
r81 17 35 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.13 $Y=1.19
+ $X2=1.255 $Y2=1.19
r82 17 18 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=1.13 $Y=1.19
+ $X2=0.445 $Y2=1.19
r83 13 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=1.105
+ $X2=0.445 $Y2=1.19
r84 13 15 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.28 $Y=1.105
+ $X2=0.28 $Y2=0.77
r85 4 33 182 $w=1.7e-07 $l=2.96648e-07 $layer=licon1_NDIFF $count=1 $X=2.945
+ $Y=0.625 $X2=3.165 $Y2=0.805
r86 3 28 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.085
+ $Y=0.625 $X2=2.225 $Y2=0.77
r87 2 21 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.075
+ $Y=0.625 $X2=1.215 $Y2=0.77
r88 1 15 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.625 $X2=0.28 $Y2=0.77
.ends

.subckt PM_SKY130_FD_SC_LS__O21A_4%VGND 1 2 3 4 5 18 22 26 30 32 34 36 38 43 48
+ 53 58 64 67 70 73 77
r81 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r82 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r83 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r84 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r85 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r86 62 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r87 62 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.56
+ $Y2=0
r88 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r89 59 73 9.23004 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=4.785 $Y=0 $X2=4.602
+ $Y2=0
r90 59 61 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=4.785 $Y=0 $X2=5.04
+ $Y2=0
r91 58 76 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=5.315 $Y=0 $X2=5.537
+ $Y2=0
r92 58 61 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=5.315 $Y=0 $X2=5.04
+ $Y2=0
r93 57 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r94 57 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r95 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r96 54 70 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.81 $Y=0 $X2=3.685
+ $Y2=0
r97 54 56 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=3.81 $Y=0 $X2=4.08
+ $Y2=0
r98 53 73 9.23004 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=4.42 $Y=0 $X2=4.602
+ $Y2=0
r99 53 56 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=4.42 $Y=0 $X2=4.08
+ $Y2=0
r100 52 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r101 51 52 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r102 49 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.89 $Y=0 $X2=1.725
+ $Y2=0
r103 49 51 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=1.89 $Y=0 $X2=2.16
+ $Y2=0
r104 48 70 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.56 $Y=0 $X2=3.685
+ $Y2=0
r105 48 51 91.3369 $w=1.68e-07 $l=1.4e-06 $layer=LI1_cond $X=3.56 $Y=0 $X2=2.16
+ $Y2=0
r106 47 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r107 47 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r108 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r109 44 64 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=0.95 $Y=0 $X2=0.782
+ $Y2=0
r110 44 46 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.95 $Y=0 $X2=1.2
+ $Y2=0
r111 43 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.56 $Y=0 $X2=1.725
+ $Y2=0
r112 43 46 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=1.56 $Y=0 $X2=1.2
+ $Y2=0
r113 41 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r114 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r115 38 64 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=0.615 $Y=0
+ $X2=0.782 $Y2=0
r116 38 40 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=0
+ $X2=0.24 $Y2=0
r117 36 71 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.88 $Y=0 $X2=3.6
+ $Y2=0
r118 36 52 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.88 $Y=0 $X2=2.16
+ $Y2=0
r119 32 76 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=5.48 $Y=0.085
+ $X2=5.537 $Y2=0
r120 32 34 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=5.48 $Y=0.085
+ $X2=5.48 $Y2=0.515
r121 28 73 1.2012 $w=3.65e-07 $l=8.5e-08 $layer=LI1_cond $X=4.602 $Y=0.085
+ $X2=4.602 $Y2=0
r122 28 30 13.1031 $w=3.63e-07 $l=4.15e-07 $layer=LI1_cond $X=4.602 $Y=0.085
+ $X2=4.602 $Y2=0.5
r123 24 70 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.685 $Y=0.085
+ $X2=3.685 $Y2=0
r124 24 26 19.1306 $w=2.48e-07 $l=4.15e-07 $layer=LI1_cond $X=3.685 $Y=0.085
+ $X2=3.685 $Y2=0.5
r125 20 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.725 $Y=0.085
+ $X2=1.725 $Y2=0
r126 20 22 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=1.725 $Y=0.085
+ $X2=1.725 $Y2=0.77
r127 16 64 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=0.782 $Y=0.085
+ $X2=0.782 $Y2=0
r128 16 18 23.5649 $w=3.33e-07 $l=6.85e-07 $layer=LI1_cond $X=0.782 $Y=0.085
+ $X2=0.782 $Y2=0.77
r129 5 34 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.34
+ $Y=0.37 $X2=5.48 $Y2=0.515
r130 4 30 182 $w=1.7e-07 $l=2.10178e-07 $layer=licon1_NDIFF $count=1 $X=4.445
+ $Y=0.37 $X2=4.6 $Y2=0.5
r131 3 26 91 $w=1.7e-07 $l=1.99687e-07 $layer=licon1_NDIFF $count=2 $X=3.58
+ $Y=0.37 $X2=3.725 $Y2=0.5
r132 2 22 182 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_NDIFF $count=1 $X=1.505
+ $Y=0.625 $X2=1.725 $Y2=0.77
r133 1 18 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.625 $X2=0.78 $Y2=0.77
.ends

