* NGSPICE file created from sky130_fd_sc_ls__o221ai_1.ext - technology: sky130A

.subckt sky130_fd_sc_ls__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
M1000 VPWR C1 Y VPB phighvt w=1.12e+06u l=150000u
+  ad=1.1816e+12p pd=6.59e+06u as=8.008e+11p ps=5.91e+06u
M1001 VGND A2 a_239_74# VNB nshort w=740000u l=150000u
+  ad=4.736e+11p pd=2.76e+06u as=6.808e+11p ps=6.28e+06u
M1002 a_239_74# B2 a_114_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=5.217e+11p ps=4.37e+06u
M1003 a_114_74# B1 a_239_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_522_368# A2 Y VPB phighvt w=1.12e+06u l=150000u
+  ad=4.704e+11p pd=3.08e+06u as=0p ps=0u
M1005 a_239_74# A1 VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR A1 a_522_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y B2 a_324_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.024e+11p ps=2.78e+06u
M1008 a_114_74# C1 Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1009 a_324_368# B1 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

