* File: sky130_fd_sc_ls__decap_4.spice
* Created: Wed Sep  2 10:59:18 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__decap_4.pex.spice"
.subckt sky130_fd_sc_ls__decap_4  VNB VPB VGND VPWR
* 
* VPWR	VPWR
* VGND	VGND
* VPB	VPB
* VNB	VNB
MM1001 N_VGND_M1001_s N_VPWR_M1001_g N_VGND_M1001_s VNB NSHORT L=1 W=0.42
+ AD=0.1176 AS=0.1176 PD=1.4 PS=1.4 NRD=0 NRS=0 M=1 R=0.42 SA=500000 SB=500000
+ A=0.42 P=2.84 MULT=1
MM1000 N_VPWR_M1000_s N_VGND_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=1 W=1 AD=0.28
+ AS=0.28 PD=2.56 PS=2.56 NRD=0 NRS=0 M=1 R=1 SA=500000 SB=500000 A=1 P=4 MULT=1
DX2_noxref VNB VPB NWDIODE A=4.278 P=8.32
*
.include "sky130_fd_sc_ls__decap_4.pxi.spice"
*
.ends
*
*
