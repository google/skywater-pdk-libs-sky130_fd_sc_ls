* NGSPICE file created from sky130_fd_sc_ls__dlrbn_2.ext - technology: sky130A

.subckt sky130_fd_sc_ls__dlrbn_2 D GATE_N RESET_B VGND VNB VPB VPWR Q Q_N
M1000 a_783_508# a_230_74# a_670_74# VPB phighvt w=420000u l=150000u
+  ad=1.995e+11p pd=1.79e+06u as=3.478e+11p ps=2.8e+06u
M1001 a_670_74# a_230_74# a_592_74# VNB nshort w=640000u l=150000u
+  ad=2.44e+11p pd=2.18e+06u as=1.536e+11p ps=1.76e+06u
M1002 a_592_74# a_27_112# VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=1.80345e+12p ps=1.499e+07u
M1003 a_670_74# a_363_74# a_595_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.4e+11p ps=2.48e+06u
M1004 VPWR a_838_48# Q VPB phighvt w=1.12e+06u l=150000u
+  ad=2.8377e+12p pd=2.106e+07u as=3.36e+11p ps=2.84e+06u
M1005 a_1446_368# a_838_48# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.95e+11p pd=2.59e+06u as=0p ps=0u
M1006 a_230_74# GATE_N VPWR VPB phighvt w=840000u l=150000u
+  ad=2.478e+11p pd=2.27e+06u as=0p ps=0u
M1007 a_230_74# GATE_N VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1008 Q_N a_1446_368# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=0p ps=0u
M1009 VGND D a_27_112# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1010 a_790_74# a_363_74# a_670_74# VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1011 a_1446_368# a_838_48# VGND VNB nshort w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=0p ps=0u
M1012 VGND a_838_48# Q VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.072e+11p ps=2.04e+06u
M1013 VPWR D a_27_112# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=2.478e+11p ps=2.27e+06u
M1014 VGND a_1446_368# Q_N VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.368e+11p ps=2.12e+06u
M1015 a_838_48# a_670_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.472e+11p pd=2.86e+06u as=0p ps=0u
M1016 a_595_392# a_27_112# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR RESET_B a_838_48# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR a_1446_368# Q_N VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND a_230_74# a_363_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1020 VGND a_838_48# a_790_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPWR a_838_48# a_783_508# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPWR a_230_74# a_363_74# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=3.83e+11p ps=2.88e+06u
M1023 Q a_838_48# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 Q_N a_1446_368# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_1066_74# a_670_74# a_838_48# VNB nshort w=740000u l=150000u
+  ad=1.776e+11p pd=1.96e+06u as=2.109e+11p ps=2.05e+06u
M1026 VGND RESET_B a_1066_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 Q a_838_48# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

