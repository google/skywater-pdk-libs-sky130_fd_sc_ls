* File: sky130_fd_sc_ls__or4bb_4.spice
* Created: Wed Sep  2 11:26:24 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__or4bb_4.pex.spice"
.subckt sky130_fd_sc_ls__or4bb_4  VNB VPB D_N C_N B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* C_N	C_N
* D_N	D_N
* VPB	VPB
* VNB	VNB
MM1006 N_VGND_M1006_d N_D_N_M1006_g N_A_27_94#_M1006_s VNB NSHORT L=0.15 W=0.64
+ AD=0.137739 AS=0.1824 PD=1.08058 PS=1.85 NRD=13.116 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75003.1 A=0.096 P=1.58 MULT=1
MM1009 N_X_M1009_d N_A_193_277#_M1009_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.159261 PD=1.02 PS=1.24942 NRD=0 NRS=12.156 M=1 R=4.93333
+ SA=75000.7 SB=75002.5 A=0.111 P=1.78 MULT=1
MM1011 N_X_M1009_d N_A_193_277#_M1011_g N_VGND_M1011_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.19035 PD=1.02 PS=1.37 NRD=0 NRS=32.784 M=1 R=4.93333 SA=75001.1
+ SB=75002 A=0.111 P=1.78 MULT=1
MM1016 N_X_M1016_d N_A_193_277#_M1016_g N_VGND_M1011_s VNB NSHORT L=0.15 W=0.74
+ AD=0.24235 AS=0.19035 PD=1.395 PS=1.37 NRD=0 NRS=32.784 M=1 R=4.93333
+ SA=75001.7 SB=75001.4 A=0.111 P=1.78 MULT=1
MM1023 N_X_M1016_d N_A_193_277#_M1023_g N_VGND_M1023_s VNB NSHORT L=0.15 W=0.74
+ AD=0.24235 AS=0.13883 PD=1.395 PS=1.17971 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.5
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1005 N_A_678_368#_M1005_d N_C_N_M1005_g N_VGND_M1023_s VNB NSHORT L=0.15
+ W=0.64 AD=0.1719 AS=0.12007 PD=1.85 PS=1.02029 NRD=0 NRS=15.936 M=1 R=4.26667
+ SA=75003.1 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1010 N_A_193_277#_M1010_d N_A_27_94#_M1010_g N_VGND_M1010_s VNB NSHORT L=0.15
+ W=0.74 AD=0.53465 AS=0.327 PD=2.185 PS=3.11 NRD=0 NRS=62.736 M=1 R=4.93333
+ SA=75000.2 SB=75003.4 A=0.111 P=1.78 MULT=1
MM1020 N_VGND_M1020_d N_A_678_368#_M1020_g N_A_193_277#_M1010_d VNB NSHORT
+ L=0.15 W=0.74 AD=0.18315 AS=0.53465 PD=1.235 PS=2.185 NRD=11.34 NRS=0 M=1
+ R=4.93333 SA=75001.8 SB=75001.8 A=0.111 P=1.78 MULT=1
MM1008 N_A_193_277#_M1008_d N_B_M1008_g N_VGND_M1020_d VNB NSHORT L=0.15 W=0.74
+ AD=0.17205 AS=0.18315 PD=1.205 PS=1.235 NRD=0 NRS=23.508 M=1 R=4.93333
+ SA=75002.5 SB=75001.2 A=0.111 P=1.78 MULT=1
MM1003 N_VGND_M1003_d N_A_M1003_g N_A_193_277#_M1008_d VNB NSHORT L=0.15 W=0.74
+ AD=0.4625 AS=0.17205 PD=2.73 PS=1.205 NRD=0 NRS=30 M=1 R=4.93333 SA=75003.1
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1015 N_VPWR_M1015_d N_D_N_M1015_g N_A_27_94#_M1015_s VPB PHIGHVT L=0.15 W=1
+ AD=0.206226 AS=0.295 PD=1.43396 PS=2.59 NRD=20.6653 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75003 A=0.15 P=2.3 MULT=1
MM1001 N_X_M1001_d N_A_193_277#_M1001_g N_VPWR_M1015_d VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.230974 PD=1.42 PS=1.60604 NRD=1.7533 NRS=3.5066 M=1 R=7.46667
+ SA=75000.7 SB=75002.4 A=0.168 P=2.54 MULT=1
MM1014 N_X_M1001_d N_A_193_277#_M1014_g N_VPWR_M1014_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.2212 PD=1.42 PS=1.515 NRD=1.7533 NRS=9.6727 M=1 R=7.46667
+ SA=75001.2 SB=75002 A=0.168 P=2.54 MULT=1
MM1018 N_X_M1018_d N_A_193_277#_M1018_g N_VPWR_M1014_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3248 AS=0.2212 PD=1.7 PS=1.515 NRD=8.7862 NRS=10.5395 M=1 R=7.46667
+ SA=75001.7 SB=75001.4 A=0.168 P=2.54 MULT=1
MM1021 N_X_M1018_d N_A_193_277#_M1021_g N_VPWR_M1021_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3248 AS=0.222098 PD=1.7 PS=1.59019 NRD=43.9704 NRS=1.7533 M=1 R=7.46667
+ SA=75002.4 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1012 N_A_678_368#_M1012_d N_C_N_M1012_g N_VPWR_M1021_s VPB PHIGHVT L=0.15 W=1
+ AD=0.295 AS=0.198302 PD=2.59 PS=1.41981 NRD=1.9503 NRS=19.6803 M=1 R=6.66667
+ SA=75003 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1000 N_A_791_392#_M1000_d N_A_27_94#_M1000_g N_A_193_277#_M1000_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.295 AS=0.15 PD=2.59 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75001.6 A=0.15 P=2.3 MULT=1
MM1019 N_A_791_392#_M1019_d N_A_27_94#_M1019_g N_A_193_277#_M1000_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75000.7 SB=75001.2 A=0.15 P=2.3 MULT=1
MM1002 N_A_1060_392#_M1002_d N_A_678_368#_M1002_g N_A_791_392#_M1019_d VPB
+ PHIGHVT L=0.15 W=1 AD=0.175 AS=0.15 PD=1.35 PS=1.3 NRD=11.8003 NRS=1.9503 M=1
+ R=6.66667 SA=75001.1 SB=75000.7 A=0.15 P=2.3 MULT=1
MM1007 N_A_1060_392#_M1002_d N_A_678_368#_M1007_g N_A_791_392#_M1007_s VPB
+ PHIGHVT L=0.15 W=1 AD=0.175 AS=0.295 PD=1.35 PS=2.59 NRD=1.9503 NRS=1.9503 M=1
+ R=6.66667 SA=75001.6 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1013 N_A_1060_392#_M1013_d N_B_M1013_g N_A_1273_392#_M1013_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.15 AS=0.295 PD=1.3 PS=2.59 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75001.6 A=0.15 P=2.3 MULT=1
MM1017 N_A_1060_392#_M1013_d N_B_M1017_g N_A_1273_392#_M1017_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75000.7 SB=75001.2 A=0.15 P=2.3 MULT=1
MM1004 N_A_1273_392#_M1017_s N_A_M1004_g N_VPWR_M1004_s VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.175 PD=1.3 PS=1.35 NRD=1.9503 NRS=11.8003 M=1 R=6.66667
+ SA=75001.1 SB=75000.7 A=0.15 P=2.3 MULT=1
MM1022 N_A_1273_392#_M1022_d N_A_M1022_g N_VPWR_M1004_s VPB PHIGHVT L=0.15 W=1
+ AD=0.295 AS=0.175 PD=2.59 PS=1.35 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75001.6 SB=75000.2 A=0.15 P=2.3 MULT=1
DX24_noxref VNB VPB NWDIODE A=16.7772 P=21.76
*
.include "sky130_fd_sc_ls__or4bb_4.pxi.spice"
*
.ends
*
*
