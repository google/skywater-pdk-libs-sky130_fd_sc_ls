* File: sky130_fd_sc_ls__ebufn_1.pxi.spice
* Created: Fri Aug 28 13:22:17 2020
* 
x_PM_SKY130_FD_SC_LS__EBUFN_1%TE_B N_TE_B_c_68_n N_TE_B_M1001_g N_TE_B_M1007_g
+ N_TE_B_c_70_n N_TE_B_c_71_n N_TE_B_c_76_n N_TE_B_M1003_g N_TE_B_c_77_n
+ N_TE_B_c_78_n N_TE_B_c_79_n N_TE_B_c_101_p N_TE_B_c_80_n N_TE_B_c_81_n TE_B
+ PM_SKY130_FD_SC_LS__EBUFN_1%TE_B
x_PM_SKY130_FD_SC_LS__EBUFN_1%A N_A_M1004_g N_A_c_159_n N_A_M1000_g A A
+ N_A_c_161_n PM_SKY130_FD_SC_LS__EBUFN_1%A
x_PM_SKY130_FD_SC_LS__EBUFN_1%A_27_404# N_A_27_404#_M1007_s N_A_27_404#_M1001_s
+ N_A_27_404#_c_194_n N_A_27_404#_c_195_n N_A_27_404#_M1005_g
+ N_A_27_404#_c_196_n N_A_27_404#_c_197_n N_A_27_404#_c_202_n
+ N_A_27_404#_c_198_n N_A_27_404#_c_199_n N_A_27_404#_c_200_n
+ N_A_27_404#_c_201_n PM_SKY130_FD_SC_LS__EBUFN_1%A_27_404#
x_PM_SKY130_FD_SC_LS__EBUFN_1%A_229_74# N_A_229_74#_M1004_d N_A_229_74#_M1000_d
+ N_A_229_74#_M1006_g N_A_229_74#_c_256_n N_A_229_74#_M1002_g
+ N_A_229_74#_c_257_n N_A_229_74#_c_264_n N_A_229_74#_c_258_n
+ N_A_229_74#_c_259_n N_A_229_74#_c_265_n N_A_229_74#_c_260_n
+ N_A_229_74#_c_261_n N_A_229_74#_c_266_n N_A_229_74#_c_267_n
+ N_A_229_74#_c_268_n N_A_229_74#_c_262_n PM_SKY130_FD_SC_LS__EBUFN_1%A_229_74#
x_PM_SKY130_FD_SC_LS__EBUFN_1%VPWR N_VPWR_M1001_d N_VPWR_M1003_s N_VPWR_c_348_n
+ N_VPWR_c_349_n VPWR N_VPWR_c_350_n N_VPWR_c_351_n N_VPWR_c_347_n
+ N_VPWR_c_353_n N_VPWR_c_354_n PM_SKY130_FD_SC_LS__EBUFN_1%VPWR
x_PM_SKY130_FD_SC_LS__EBUFN_1%Z N_Z_M1006_d N_Z_M1002_d N_Z_c_396_n N_Z_c_397_n
+ N_Z_c_394_n Z Z N_Z_c_395_n PM_SKY130_FD_SC_LS__EBUFN_1%Z
x_PM_SKY130_FD_SC_LS__EBUFN_1%VGND N_VGND_M1007_d N_VGND_M1005_s N_VGND_c_419_n
+ N_VGND_c_420_n VGND N_VGND_c_421_n N_VGND_c_422_n N_VGND_c_423_n
+ N_VGND_c_424_n N_VGND_c_425_n PM_SKY130_FD_SC_LS__EBUFN_1%VGND
cc_1 VNB N_TE_B_c_68_n 0.0167472f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.945
cc_2 VNB N_TE_B_M1007_g 0.0507161f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=0.645
cc_3 VNB N_TE_B_c_70_n 0.0118263f $X=-0.19 $Y=-0.245 $X2=2.68 $Y2=1.69
cc_4 VNB N_TE_B_c_71_n 0.0043072f $X=-0.19 $Y=-0.245 $X2=2.195 $Y2=1.69
cc_5 VNB TE_B 0.00341842f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_6 VNB N_A_M1004_g 0.0580975f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.44
cc_7 VNB N_A_c_159_n 0.00846483f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=0.645
cc_8 VNB A 0.00358455f $X=-0.19 $Y=-0.245 $X2=2.195 $Y2=1.69
cc_9 VNB N_A_c_161_n 0.0229517f $X=-0.19 $Y=-0.245 $X2=2.03 $Y2=2.505
cc_10 VNB N_A_27_404#_c_194_n 0.0395168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_27_404#_c_195_n 0.0172236f $X=-0.19 $Y=-0.245 $X2=2.12 $Y2=2.34
cc_12 VNB N_A_27_404#_c_196_n 0.0365396f $X=-0.19 $Y=-0.245 $X2=2.755 $Y2=2.4
cc_13 VNB N_A_27_404#_c_197_n 0.0118865f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_404#_c_198_n 0.0162952f $X=-0.19 $Y=-0.245 $X2=2.03 $Y2=2.505
cc_15 VNB N_A_27_404#_c_199_n 9.95647e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_27_404#_c_200_n 0.0271006f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_27_404#_c_201_n 0.0424548f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.665
cc_18 VNB N_A_229_74#_M1006_g 0.0284822f $X=-0.19 $Y=-0.245 $X2=2.12 $Y2=2.34
cc_19 VNB N_A_229_74#_c_256_n 0.0369877f $X=-0.19 $Y=-0.245 $X2=2.195 $Y2=1.69
cc_20 VNB N_A_229_74#_c_257_n 0.0139199f $X=-0.19 $Y=-0.245 $X2=2.03 $Y2=2.34
cc_21 VNB N_A_229_74#_c_258_n 0.029099f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_229_74#_c_259_n 0.00347683f $X=-0.19 $Y=-0.245 $X2=2.03 $Y2=2.465
cc_23 VNB N_A_229_74#_c_260_n 0.00135177f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_229_74#_c_261_n 0.00449629f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.665
cc_25 VNB N_A_229_74#_c_262_n 0.0147135f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VPWR_c_347_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.665
cc_27 VNB N_Z_c_394_n 0.0252276f $X=-0.19 $Y=-0.245 $X2=2.03 $Y2=2.505
cc_28 VNB N_Z_c_395_n 0.0503455f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_419_n 0.00944084f $X=-0.19 $Y=-0.245 $X2=2.195 $Y2=1.69
cc_30 VNB N_VGND_c_420_n 0.0203845f $X=-0.19 $Y=-0.245 $X2=2.03 $Y2=2.505
cc_31 VNB N_VGND_c_421_n 0.042784f $X=-0.19 $Y=-0.245 $X2=1.865 $Y2=2.505
cc_32 VNB N_VGND_c_422_n 0.033384f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_423_n 0.24203f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.665
cc_34 VNB N_VGND_c_424_n 0.0270337f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.665
cc_35 VNB N_VGND_c_425_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.83
cc_36 VPB N_TE_B_c_68_n 0.0465437f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.945
cc_37 VPB N_TE_B_c_70_n 0.0175721f $X=-0.19 $Y=1.66 $X2=2.68 $Y2=1.69
cc_38 VPB N_TE_B_c_71_n 0.00373927f $X=-0.19 $Y=1.66 $X2=2.195 $Y2=1.69
cc_39 VPB N_TE_B_c_76_n 0.0162967f $X=-0.19 $Y=1.66 $X2=2.755 $Y2=1.765
cc_40 VPB N_TE_B_c_77_n 0.0395776f $X=-0.19 $Y=1.66 $X2=2.03 $Y2=2.34
cc_41 VPB N_TE_B_c_78_n 0.0034088f $X=-0.19 $Y=1.66 $X2=0.75 $Y2=2.42
cc_42 VPB N_TE_B_c_79_n 0.00956627f $X=-0.19 $Y=1.66 $X2=1.865 $Y2=2.505
cc_43 VPB N_TE_B_c_80_n 0.00742537f $X=-0.19 $Y=1.66 $X2=2.03 $Y2=2.505
cc_44 VPB N_TE_B_c_81_n 0.0723932f $X=-0.19 $Y=1.66 $X2=2.03 $Y2=2.505
cc_45 VPB TE_B 0.00363527f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_46 VPB N_A_c_159_n 0.0393247f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=0.645
cc_47 VPB A 0.00240167f $X=-0.19 $Y=1.66 $X2=2.195 $Y2=1.69
cc_48 VPB N_A_c_161_n 0.022161f $X=-0.19 $Y=1.66 $X2=2.03 $Y2=2.505
cc_49 VPB N_A_27_404#_c_202_n 0.0409021f $X=-0.19 $Y=1.66 $X2=2.03 $Y2=2.505
cc_50 VPB N_A_27_404#_c_198_n 0.0159586f $X=-0.19 $Y=1.66 $X2=2.03 $Y2=2.505
cc_51 VPB N_A_229_74#_c_256_n 0.0283379f $X=-0.19 $Y=1.66 $X2=2.195 $Y2=1.69
cc_52 VPB N_A_229_74#_c_264_n 0.00343925f $X=-0.19 $Y=1.66 $X2=0.75 $Y2=2.42
cc_53 VPB N_A_229_74#_c_265_n 0.00833716f $X=-0.19 $Y=1.66 $X2=2.03 $Y2=2.505
cc_54 VPB N_A_229_74#_c_266_n 0.0039456f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_A_229_74#_c_267_n 0.00831023f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.83
cc_56 VPB N_A_229_74#_c_268_n 0.00604866f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_A_229_74#_c_262_n 0.00163226f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_348_n 0.0160797f $X=-0.19 $Y=1.66 $X2=2.195 $Y2=1.69
cc_59 VPB N_VPWR_c_349_n 0.0152717f $X=-0.19 $Y=1.66 $X2=2.03 $Y2=2.505
cc_60 VPB N_VPWR_c_350_n 0.0380943f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_351_n 0.0343749f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.665
cc_62 VPB N_VPWR_c_347_n 0.0878651f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.665
cc_63 VPB N_VPWR_c_353_n 0.02685f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_354_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_Z_c_396_n 0.046779f $X=-0.19 $Y=1.66 $X2=2.12 $Y2=2.34
cc_66 VPB N_Z_c_397_n 0.0202175f $X=-0.19 $Y=1.66 $X2=2.755 $Y2=2.4
cc_67 VPB N_Z_c_394_n 0.00778546f $X=-0.19 $Y=1.66 $X2=2.03 $Y2=2.505
cc_68 N_TE_B_M1007_g N_A_M1004_g 0.0347876f $X=0.62 $Y=0.645 $X2=0 $Y2=0
cc_69 N_TE_B_c_68_n N_A_c_159_n 0.0397137f $X=0.505 $Y=1.945 $X2=0 $Y2=0
cc_70 N_TE_B_c_78_n N_A_c_159_n 0.00943441f $X=0.75 $Y=2.42 $X2=0 $Y2=0
cc_71 N_TE_B_c_79_n N_A_c_159_n 0.0157572f $X=1.865 $Y=2.505 $X2=0 $Y2=0
cc_72 N_TE_B_c_80_n N_A_c_159_n 0.00222065f $X=2.03 $Y=2.505 $X2=0 $Y2=0
cc_73 N_TE_B_c_81_n N_A_c_159_n 0.0105448f $X=2.03 $Y=2.505 $X2=0 $Y2=0
cc_74 TE_B N_A_c_159_n 0.00231785f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_75 N_TE_B_c_68_n A 3.47969e-19 $X=0.505 $Y=1.945 $X2=0 $Y2=0
cc_76 N_TE_B_c_71_n A 0.00172831f $X=2.195 $Y=1.69 $X2=0 $Y2=0
cc_77 N_TE_B_c_79_n A 0.00405436f $X=1.865 $Y=2.505 $X2=0 $Y2=0
cc_78 TE_B A 0.0279811f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_79 N_TE_B_c_71_n N_A_c_161_n 0.00676649f $X=2.195 $Y=1.69 $X2=0 $Y2=0
cc_80 N_TE_B_c_70_n N_A_27_404#_c_194_n 0.0258296f $X=2.68 $Y=1.69 $X2=0 $Y2=0
cc_81 N_TE_B_M1007_g N_A_27_404#_c_196_n 0.0112033f $X=0.62 $Y=0.645 $X2=0 $Y2=0
cc_82 N_TE_B_c_68_n N_A_27_404#_c_197_n 0.00115196f $X=0.505 $Y=1.945 $X2=0
+ $Y2=0
cc_83 TE_B N_A_27_404#_c_197_n 0.00843991f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_84 N_TE_B_c_68_n N_A_27_404#_c_202_n 0.0161858f $X=0.505 $Y=1.945 $X2=0 $Y2=0
cc_85 N_TE_B_c_78_n N_A_27_404#_c_202_n 0.0255666f $X=0.75 $Y=2.42 $X2=0 $Y2=0
cc_86 N_TE_B_c_101_p N_A_27_404#_c_202_n 0.0115776f $X=0.835 $Y=2.505 $X2=0
+ $Y2=0
cc_87 TE_B N_A_27_404#_c_202_n 0.00146231f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_88 N_TE_B_c_68_n N_A_27_404#_c_198_n 0.0102333f $X=0.505 $Y=1.945 $X2=0 $Y2=0
cc_89 N_TE_B_M1007_g N_A_27_404#_c_198_n 0.00389989f $X=0.62 $Y=0.645 $X2=0
+ $Y2=0
cc_90 N_TE_B_c_78_n N_A_27_404#_c_198_n 0.00487266f $X=0.75 $Y=2.42 $X2=0 $Y2=0
cc_91 TE_B N_A_27_404#_c_198_n 0.0252195f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_92 N_TE_B_c_71_n N_A_27_404#_c_199_n 5.97257e-19 $X=2.195 $Y=1.69 $X2=0 $Y2=0
cc_93 N_TE_B_c_68_n N_A_27_404#_c_200_n 5.1855e-19 $X=0.505 $Y=1.945 $X2=0 $Y2=0
cc_94 N_TE_B_M1007_g N_A_27_404#_c_200_n 0.0169119f $X=0.62 $Y=0.645 $X2=0 $Y2=0
cc_95 TE_B N_A_27_404#_c_200_n 0.0224553f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_96 N_TE_B_c_71_n N_A_27_404#_c_201_n 0.0258296f $X=2.195 $Y=1.69 $X2=0 $Y2=0
cc_97 N_TE_B_c_79_n N_A_229_74#_M1000_d 0.00839715f $X=1.865 $Y=2.505 $X2=0
+ $Y2=0
cc_98 N_TE_B_c_70_n N_A_229_74#_c_256_n 0.00768303f $X=2.68 $Y=1.69 $X2=0 $Y2=0
cc_99 N_TE_B_c_76_n N_A_229_74#_c_256_n 0.0575197f $X=2.755 $Y=1.765 $X2=0 $Y2=0
cc_100 N_TE_B_c_78_n N_A_229_74#_c_264_n 0.0110927f $X=0.75 $Y=2.42 $X2=0 $Y2=0
cc_101 N_TE_B_c_79_n N_A_229_74#_c_264_n 0.034259f $X=1.865 $Y=2.505 $X2=0 $Y2=0
cc_102 N_TE_B_c_77_n N_A_229_74#_c_265_n 0.00126228f $X=2.03 $Y=2.34 $X2=0 $Y2=0
cc_103 N_TE_B_c_79_n N_A_229_74#_c_265_n 0.00972763f $X=1.865 $Y=2.505 $X2=0
+ $Y2=0
cc_104 N_TE_B_c_80_n N_A_229_74#_c_265_n 0.0079822f $X=2.03 $Y=2.505 $X2=0 $Y2=0
cc_105 N_TE_B_c_81_n N_A_229_74#_c_265_n 6.96394e-19 $X=2.03 $Y=2.505 $X2=0
+ $Y2=0
cc_106 N_TE_B_c_77_n N_A_229_74#_c_266_n 0.00163127f $X=2.03 $Y=2.34 $X2=0 $Y2=0
cc_107 N_TE_B_c_71_n N_A_229_74#_c_267_n 0.00203925f $X=2.195 $Y=1.69 $X2=0
+ $Y2=0
cc_108 N_TE_B_c_76_n N_A_229_74#_c_267_n 5.96038e-19 $X=2.755 $Y=1.765 $X2=0
+ $Y2=0
cc_109 N_TE_B_c_77_n N_A_229_74#_c_267_n 0.0145621f $X=2.03 $Y=2.34 $X2=0 $Y2=0
cc_110 N_TE_B_c_80_n N_A_229_74#_c_267_n 0.0141324f $X=2.03 $Y=2.505 $X2=0 $Y2=0
cc_111 N_TE_B_c_81_n N_A_229_74#_c_267_n 5.95224e-19 $X=2.03 $Y=2.505 $X2=0
+ $Y2=0
cc_112 N_TE_B_c_70_n N_A_229_74#_c_268_n 0.00771499f $X=2.68 $Y=1.69 $X2=0 $Y2=0
cc_113 N_TE_B_c_71_n N_A_229_74#_c_268_n 0.00114693f $X=2.195 $Y=1.69 $X2=0
+ $Y2=0
cc_114 N_TE_B_c_77_n N_A_229_74#_c_268_n 0.00440865f $X=2.03 $Y=2.34 $X2=0 $Y2=0
cc_115 N_TE_B_c_80_n N_A_229_74#_c_268_n 0.00203003f $X=2.03 $Y=2.505 $X2=0
+ $Y2=0
cc_116 N_TE_B_c_70_n N_A_229_74#_c_262_n 0.0149598f $X=2.68 $Y=1.69 $X2=0 $Y2=0
cc_117 N_TE_B_c_76_n N_A_229_74#_c_262_n 0.011723f $X=2.755 $Y=1.765 $X2=0 $Y2=0
cc_118 N_TE_B_c_78_n N_VPWR_M1001_d 0.0119759f $X=0.75 $Y=2.42 $X2=-0.19
+ $Y2=-0.245
cc_119 N_TE_B_c_79_n N_VPWR_M1001_d 0.00804454f $X=1.865 $Y=2.505 $X2=-0.19
+ $Y2=-0.245
cc_120 N_TE_B_c_101_p N_VPWR_M1001_d 0.00501699f $X=0.835 $Y=2.505 $X2=-0.19
+ $Y2=-0.245
cc_121 N_TE_B_c_68_n N_VPWR_c_348_n 0.00438046f $X=0.505 $Y=1.945 $X2=0 $Y2=0
cc_122 N_TE_B_c_79_n N_VPWR_c_348_n 0.0112732f $X=1.865 $Y=2.505 $X2=0 $Y2=0
cc_123 N_TE_B_c_101_p N_VPWR_c_348_n 0.0146637f $X=0.835 $Y=2.505 $X2=0 $Y2=0
cc_124 N_TE_B_c_70_n N_VPWR_c_349_n 0.00136259f $X=2.68 $Y=1.69 $X2=0 $Y2=0
cc_125 N_TE_B_c_76_n N_VPWR_c_349_n 0.0204486f $X=2.755 $Y=1.765 $X2=0 $Y2=0
cc_126 N_TE_B_c_77_n N_VPWR_c_349_n 0.00444525f $X=2.03 $Y=2.34 $X2=0 $Y2=0
cc_127 N_TE_B_c_80_n N_VPWR_c_349_n 0.0537867f $X=2.03 $Y=2.505 $X2=0 $Y2=0
cc_128 N_TE_B_c_81_n N_VPWR_c_349_n 0.00478718f $X=2.03 $Y=2.505 $X2=0 $Y2=0
cc_129 N_TE_B_c_79_n N_VPWR_c_350_n 0.0117562f $X=1.865 $Y=2.505 $X2=0 $Y2=0
cc_130 N_TE_B_c_80_n N_VPWR_c_350_n 0.015584f $X=2.03 $Y=2.505 $X2=0 $Y2=0
cc_131 N_TE_B_c_81_n N_VPWR_c_350_n 0.00192529f $X=2.03 $Y=2.505 $X2=0 $Y2=0
cc_132 N_TE_B_c_76_n N_VPWR_c_351_n 0.00413917f $X=2.755 $Y=1.765 $X2=0 $Y2=0
cc_133 N_TE_B_c_68_n N_VPWR_c_347_n 0.00514438f $X=0.505 $Y=1.945 $X2=0 $Y2=0
cc_134 N_TE_B_c_76_n N_VPWR_c_347_n 0.00817532f $X=2.755 $Y=1.765 $X2=0 $Y2=0
cc_135 N_TE_B_c_79_n N_VPWR_c_347_n 0.0237096f $X=1.865 $Y=2.505 $X2=0 $Y2=0
cc_136 N_TE_B_c_101_p N_VPWR_c_347_n 7.17789e-19 $X=0.835 $Y=2.505 $X2=0 $Y2=0
cc_137 N_TE_B_c_80_n N_VPWR_c_347_n 0.0120766f $X=2.03 $Y=2.505 $X2=0 $Y2=0
cc_138 N_TE_B_c_68_n N_VPWR_c_353_n 0.00494504f $X=0.505 $Y=1.945 $X2=0 $Y2=0
cc_139 N_TE_B_c_76_n N_Z_c_397_n 0.00353308f $X=2.755 $Y=1.765 $X2=0 $Y2=0
cc_140 N_TE_B_M1007_g N_VGND_c_419_n 0.00408774f $X=0.62 $Y=0.645 $X2=0 $Y2=0
cc_141 N_TE_B_M1007_g N_VGND_c_423_n 0.00911508f $X=0.62 $Y=0.645 $X2=0 $Y2=0
cc_142 N_TE_B_M1007_g N_VGND_c_424_n 0.00461464f $X=0.62 $Y=0.645 $X2=0 $Y2=0
cc_143 N_A_c_159_n N_A_27_404#_c_202_n 8.81476e-19 $X=1.125 $Y=1.945 $X2=0 $Y2=0
cc_144 N_A_M1004_g N_A_27_404#_c_200_n 0.0175221f $X=1.07 $Y=0.645 $X2=0 $Y2=0
cc_145 N_A_c_159_n N_A_27_404#_c_200_n 0.0120221f $X=1.125 $Y=1.945 $X2=0 $Y2=0
cc_146 A N_A_27_404#_c_200_n 0.0568065f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_147 N_A_c_159_n N_A_229_74#_c_264_n 0.00472247f $X=1.125 $Y=1.945 $X2=0 $Y2=0
cc_148 A N_A_229_74#_c_264_n 0.0473241f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_149 N_A_c_161_n N_A_229_74#_c_264_n 0.0103846f $X=1.51 $Y=1.665 $X2=0 $Y2=0
cc_150 N_A_M1004_g N_A_229_74#_c_259_n 0.00357394f $X=1.07 $Y=0.645 $X2=0 $Y2=0
cc_151 A N_A_229_74#_c_267_n 0.0100487f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_152 N_A_c_161_n N_A_229_74#_c_267_n 2.98913e-19 $X=1.51 $Y=1.665 $X2=0 $Y2=0
cc_153 A N_A_229_74#_c_262_n 0.00704617f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_154 N_A_c_159_n N_VPWR_c_348_n 0.00663705f $X=1.125 $Y=1.945 $X2=0 $Y2=0
cc_155 N_A_c_159_n N_VPWR_c_350_n 0.00397762f $X=1.125 $Y=1.945 $X2=0 $Y2=0
cc_156 N_A_c_159_n N_VPWR_c_347_n 0.00514438f $X=1.125 $Y=1.945 $X2=0 $Y2=0
cc_157 N_A_M1004_g N_VGND_c_419_n 0.00405933f $X=1.07 $Y=0.645 $X2=0 $Y2=0
cc_158 N_A_M1004_g N_VGND_c_421_n 0.00461464f $X=1.07 $Y=0.645 $X2=0 $Y2=0
cc_159 N_A_M1004_g N_VGND_c_423_n 0.00912604f $X=1.07 $Y=0.645 $X2=0 $Y2=0
cc_160 N_A_27_404#_c_195_n N_A_229_74#_M1006_g 0.0303584f $X=2.77 $Y=1.185 $X2=0
+ $Y2=0
cc_161 N_A_27_404#_c_194_n N_A_229_74#_c_256_n 0.0303584f $X=2.695 $Y=1.295
+ $X2=0 $Y2=0
cc_162 N_A_27_404#_c_194_n N_A_229_74#_c_258_n 0.00892394f $X=2.695 $Y=1.295
+ $X2=0 $Y2=0
cc_163 N_A_27_404#_c_200_n N_A_229_74#_c_258_n 0.0553447f $X=1.87 $Y=1.245 $X2=0
+ $Y2=0
cc_164 N_A_27_404#_c_201_n N_A_229_74#_c_258_n 0.00808505f $X=2.2 $Y=1.24 $X2=0
+ $Y2=0
cc_165 N_A_27_404#_c_196_n N_A_229_74#_c_259_n 0.00210758f $X=0.405 $Y=0.645
+ $X2=0 $Y2=0
cc_166 N_A_27_404#_c_200_n N_A_229_74#_c_259_n 0.0243942f $X=1.87 $Y=1.245 $X2=0
+ $Y2=0
cc_167 N_A_27_404#_c_199_n N_A_229_74#_c_265_n 0.00244148f $X=2.035 $Y=1.24
+ $X2=0 $Y2=0
cc_168 N_A_27_404#_c_201_n N_A_229_74#_c_265_n 0.0015619f $X=2.2 $Y=1.24 $X2=0
+ $Y2=0
cc_169 N_A_27_404#_c_194_n N_A_229_74#_c_260_n 0.0117554f $X=2.695 $Y=1.295
+ $X2=0 $Y2=0
cc_170 N_A_27_404#_c_195_n N_A_229_74#_c_260_n 0.00393509f $X=2.77 $Y=1.185
+ $X2=0 $Y2=0
cc_171 N_A_27_404#_c_199_n N_A_229_74#_c_260_n 0.00939079f $X=2.035 $Y=1.24
+ $X2=0 $Y2=0
cc_172 N_A_27_404#_c_201_n N_A_229_74#_c_260_n 0.00179597f $X=2.2 $Y=1.24 $X2=0
+ $Y2=0
cc_173 N_A_27_404#_c_199_n N_A_229_74#_c_267_n 0.00701624f $X=2.035 $Y=1.24
+ $X2=0 $Y2=0
cc_174 N_A_27_404#_c_201_n N_A_229_74#_c_267_n 0.00200399f $X=2.2 $Y=1.24 $X2=0
+ $Y2=0
cc_175 N_A_27_404#_c_199_n N_A_229_74#_c_268_n 0.00236052f $X=2.035 $Y=1.24
+ $X2=0 $Y2=0
cc_176 N_A_27_404#_c_201_n N_A_229_74#_c_268_n 0.00164906f $X=2.2 $Y=1.24 $X2=0
+ $Y2=0
cc_177 N_A_27_404#_c_194_n N_A_229_74#_c_262_n 0.0207665f $X=2.695 $Y=1.295
+ $X2=0 $Y2=0
cc_178 N_A_27_404#_c_199_n N_A_229_74#_c_262_n 0.00102519f $X=2.035 $Y=1.24
+ $X2=0 $Y2=0
cc_179 N_A_27_404#_c_202_n N_VPWR_c_348_n 0.00814855f $X=0.28 $Y=2.165 $X2=0
+ $Y2=0
cc_180 N_A_27_404#_c_202_n N_VPWR_c_347_n 0.0123843f $X=0.28 $Y=2.165 $X2=0
+ $Y2=0
cc_181 N_A_27_404#_c_202_n N_VPWR_c_353_n 0.0113277f $X=0.28 $Y=2.165 $X2=0
+ $Y2=0
cc_182 N_A_27_404#_c_195_n N_Z_c_395_n 0.00258266f $X=2.77 $Y=1.185 $X2=0 $Y2=0
cc_183 N_A_27_404#_c_200_n N_VGND_c_419_n 0.0126908f $X=1.87 $Y=1.245 $X2=0
+ $Y2=0
cc_184 N_A_27_404#_c_194_n N_VGND_c_420_n 8.1259e-19 $X=2.695 $Y=1.295 $X2=0
+ $Y2=0
cc_185 N_A_27_404#_c_195_n N_VGND_c_420_n 0.0110763f $X=2.77 $Y=1.185 $X2=0
+ $Y2=0
cc_186 N_A_27_404#_c_195_n N_VGND_c_422_n 0.00383152f $X=2.77 $Y=1.185 $X2=0
+ $Y2=0
cc_187 N_A_27_404#_c_195_n N_VGND_c_423_n 0.0075725f $X=2.77 $Y=1.185 $X2=0
+ $Y2=0
cc_188 N_A_27_404#_c_196_n N_VGND_c_423_n 0.0152899f $X=0.405 $Y=0.645 $X2=0
+ $Y2=0
cc_189 N_A_27_404#_c_196_n N_VGND_c_424_n 0.0129976f $X=0.405 $Y=0.645 $X2=0
+ $Y2=0
cc_190 N_A_229_74#_c_268_n N_VPWR_M1003_s 7.86634e-19 $X=2.46 $Y=1.6 $X2=0 $Y2=0
cc_191 N_A_229_74#_c_262_n N_VPWR_M1003_s 0.00179736f $X=3.065 $Y=1.6 $X2=0
+ $Y2=0
cc_192 N_A_229_74#_c_256_n N_VPWR_c_349_n 0.00322639f $X=3.175 $Y=1.765 $X2=0
+ $Y2=0
cc_193 N_A_229_74#_c_266_n N_VPWR_c_349_n 0.00258243f $X=1.695 $Y=2.125 $X2=0
+ $Y2=0
cc_194 N_A_229_74#_c_267_n N_VPWR_c_349_n 0.00723556f $X=2.05 $Y=1.795 $X2=0
+ $Y2=0
cc_195 N_A_229_74#_c_268_n N_VPWR_c_349_n 0.0232098f $X=2.46 $Y=1.6 $X2=0 $Y2=0
cc_196 N_A_229_74#_c_256_n N_VPWR_c_351_n 0.00445602f $X=3.175 $Y=1.765 $X2=0
+ $Y2=0
cc_197 N_A_229_74#_c_256_n N_VPWR_c_347_n 0.00862073f $X=3.175 $Y=1.765 $X2=0
+ $Y2=0
cc_198 N_A_229_74#_c_262_n A_566_368# 0.0069114f $X=3.065 $Y=1.6 $X2=-0.19
+ $Y2=-0.245
cc_199 N_A_229_74#_c_256_n N_Z_c_396_n 0.0168767f $X=3.175 $Y=1.765 $X2=0 $Y2=0
cc_200 N_A_229_74#_c_256_n N_Z_c_397_n 0.00873641f $X=3.175 $Y=1.765 $X2=0 $Y2=0
cc_201 N_A_229_74#_c_261_n N_Z_c_397_n 0.0150324f $X=3.25 $Y=1.485 $X2=0 $Y2=0
cc_202 N_A_229_74#_c_262_n N_Z_c_397_n 0.00327028f $X=3.065 $Y=1.6 $X2=0 $Y2=0
cc_203 N_A_229_74#_M1006_g N_Z_c_394_n 0.00394404f $X=3.16 $Y=0.74 $X2=0 $Y2=0
cc_204 N_A_229_74#_c_256_n N_Z_c_394_n 0.00462737f $X=3.175 $Y=1.765 $X2=0 $Y2=0
cc_205 N_A_229_74#_c_261_n N_Z_c_394_n 0.0262124f $X=3.25 $Y=1.485 $X2=0 $Y2=0
cc_206 N_A_229_74#_c_262_n N_Z_c_394_n 0.00459995f $X=3.065 $Y=1.6 $X2=0 $Y2=0
cc_207 N_A_229_74#_M1006_g N_Z_c_395_n 0.0164306f $X=3.16 $Y=0.74 $X2=0 $Y2=0
cc_208 N_A_229_74#_c_256_n N_Z_c_395_n 0.00423018f $X=3.175 $Y=1.765 $X2=0 $Y2=0
cc_209 N_A_229_74#_c_260_n N_Z_c_395_n 0.00263651f $X=2.56 $Y=1.32 $X2=0 $Y2=0
cc_210 N_A_229_74#_c_261_n N_Z_c_395_n 0.0157141f $X=3.25 $Y=1.485 $X2=0 $Y2=0
cc_211 N_A_229_74#_c_258_n N_VGND_M1005_s 0.00506875f $X=2.46 $Y=0.895 $X2=0
+ $Y2=0
cc_212 N_A_229_74#_c_260_n N_VGND_M1005_s 0.00433646f $X=2.56 $Y=1.32 $X2=0
+ $Y2=0
cc_213 N_A_229_74#_M1006_g N_VGND_c_420_n 0.00138195f $X=3.16 $Y=0.74 $X2=0
+ $Y2=0
cc_214 N_A_229_74#_c_258_n N_VGND_c_420_n 0.0207988f $X=2.46 $Y=0.895 $X2=0
+ $Y2=0
cc_215 N_A_229_74#_c_257_n N_VGND_c_421_n 0.00811823f $X=1.285 $Y=0.645 $X2=0
+ $Y2=0
cc_216 N_A_229_74#_M1006_g N_VGND_c_422_n 0.00434272f $X=3.16 $Y=0.74 $X2=0
+ $Y2=0
cc_217 N_A_229_74#_M1006_g N_VGND_c_423_n 0.00825123f $X=3.16 $Y=0.74 $X2=0
+ $Y2=0
cc_218 N_A_229_74#_c_257_n N_VGND_c_423_n 0.0100099f $X=1.285 $Y=0.645 $X2=0
+ $Y2=0
cc_219 N_A_229_74#_c_258_n N_VGND_c_423_n 0.0343415f $X=2.46 $Y=0.895 $X2=0
+ $Y2=0
cc_220 N_VPWR_c_351_n N_Z_c_396_n 0.0230718f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_221 N_VPWR_c_347_n N_Z_c_396_n 0.0190639f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_222 N_VPWR_c_349_n N_Z_c_397_n 0.028003f $X=2.53 $Y=2.135 $X2=0 $Y2=0
cc_223 N_Z_c_395_n N_VGND_c_420_n 0.00955365f $X=3.375 $Y=0.515 $X2=0 $Y2=0
cc_224 N_Z_c_395_n N_VGND_c_422_n 0.0241574f $X=3.375 $Y=0.515 $X2=0 $Y2=0
cc_225 N_Z_c_395_n N_VGND_c_423_n 0.019939f $X=3.375 $Y=0.515 $X2=0 $Y2=0
