* NGSPICE file created from sky130_fd_sc_ls__fah_4.ext - technology: sky130A

.subckt sky130_fd_sc_ls__fah_4 A B CI VGND VNB VPB VPWR COUT SUM
M1000 a_200_74# a_586_257# a_528_362# VPB phighvt w=840000u l=150000u
+  ad=7.739e+11p pd=5.79e+06u as=2.562e+11p ps=2.29e+06u
M1001 a_427_362# a_27_74# VGND VNB nshort w=740000u l=150000u
+  ad=4.026e+11p pd=3.94e+06u as=3.15805e+12p ps=2.382e+07u
M1002 a_1378_125# a_536_114# a_1265_379# VPB phighvt w=840000u l=150000u
+  ad=7.451e+11p pd=5.69e+06u as=3.738e+11p ps=2.57e+06u
M1003 SUM a_1278_102# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=6.832e+11p pd=5.7e+06u as=4.77725e+12p ps=2.973e+07u
M1004 a_536_114# B a_200_74# VPB phighvt w=840000u l=150000u
+  ad=2.52e+11p pd=2.28e+06u as=0p ps=0u
M1005 COUT a_1265_379# VGND VNB nshort w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=0p ps=0u
M1006 VGND a_1265_379# COUT VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 COUT a_1265_379# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=6.72e+11p pd=5.68e+06u as=0p ps=0u
M1008 a_1278_102# a_528_362# a_1378_125# VPB phighvt w=840000u l=150000u
+  ad=6.72e+11p pd=3.28e+06u as=0p ps=0u
M1009 VGND a_1265_379# COUT VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR a_1278_102# SUM VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_427_362# a_586_257# a_536_114# VPB phighvt w=840000u l=150000u
+  ad=6.202e+11p pd=5.22e+06u as=0p ps=0u
M1012 a_586_257# B VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=4.0435e+11p pd=3.01e+06u as=0p ps=0u
M1013 VPWR a_1378_125# a_1183_102# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=3.90725e+11p ps=3e+06u
M1014 VPWR a_1265_379# COUT VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND CI a_1378_125# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=3.616e+11p ps=3.69e+06u
M1016 VPWR a_1265_379# COUT VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_536_114# B a_427_362# VNB nshort w=640000u l=150000u
+  ad=1.792e+11p pd=1.84e+06u as=0p ps=0u
M1018 VGND a_1378_125# a_1183_102# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=4.4305e+11p ps=3.95e+06u
M1019 VPWR CI a_1378_125# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 COUT a_1265_379# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_586_257# B VGND VNB nshort w=740000u l=150000u
+  ad=5.59925e+11p pd=5.19e+06u as=0p ps=0u
M1022 a_1278_102# a_528_362# a_1183_102# VNB nshort w=640000u l=150000u
+  ad=2.44125e+11p pd=2.21e+06u as=0p ps=0u
M1023 a_586_257# a_536_114# a_1265_379# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=2.3685e+11p ps=2.18e+06u
M1024 COUT a_1265_379# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 SUM a_1278_102# VGND VNB nshort w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=0p ps=0u
M1026 a_200_74# a_586_257# a_536_114# VNB nshort w=640000u l=150000u
+  ad=4.268e+11p pd=4.01e+06u as=0p ps=0u
M1027 a_528_362# B a_200_74# VNB nshort w=640000u l=150000u
+  ad=2.048e+11p pd=1.92e+06u as=0p ps=0u
M1028 VGND a_1278_102# SUM VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 SUM a_1278_102# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_1183_102# a_536_114# a_1278_102# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VPWR a_1278_102# SUM VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_200_74# A VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_427_362# a_586_257# a_528_362# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 VPWR A a_27_74# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.95e+11p ps=2.59e+06u
M1035 a_427_362# a_27_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_1265_379# a_528_362# a_586_257# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 VGND A a_27_74# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1038 a_200_74# A VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_1378_125# a_536_114# a_1278_102# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1040 a_1265_379# a_528_362# a_1378_125# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1041 SUM a_1278_102# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1042 a_528_362# B a_427_362# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1043 VGND a_1278_102# SUM VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

