* File: sky130_fd_sc_ls__o31ai_4.pex.spice
* Created: Fri Aug 28 13:53:48 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__O31AI_4%A1 3 5 7 8 10 13 15 17 20 22 23 25 26 28 31
+ 33 34 35 36 37
c82 23 0 1.91457e-19 $X=1.5 $Y=1.425
r83 52 53 1.94355 $w=3.72e-07 $l=1.5e-08 $layer=POLY_cond $X=1.41 $Y=1.557
+ $X2=1.425 $Y2=1.557
r84 50 52 18.7876 $w=3.72e-07 $l=1.45e-07 $layer=POLY_cond $X=1.265 $Y=1.557
+ $X2=1.41 $Y2=1.557
r85 50 51 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.265
+ $Y=1.515 $X2=1.265 $Y2=1.515
r86 48 50 34.9839 $w=3.72e-07 $l=2.7e-07 $layer=POLY_cond $X=0.995 $Y=1.557
+ $X2=1.265 $Y2=1.557
r87 47 48 4.53495 $w=3.72e-07 $l=3.5e-08 $layer=POLY_cond $X=0.96 $Y=1.557
+ $X2=0.995 $Y2=1.557
r88 45 47 48.5887 $w=3.72e-07 $l=3.75e-07 $layer=POLY_cond $X=0.585 $Y=1.557
+ $X2=0.96 $Y2=1.557
r89 45 46 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.585
+ $Y=1.515 $X2=0.585 $Y2=1.515
r90 43 45 9.71774 $w=3.72e-07 $l=7.5e-08 $layer=POLY_cond $X=0.51 $Y=1.557
+ $X2=0.585 $Y2=1.557
r91 42 43 1.94355 $w=3.72e-07 $l=1.5e-08 $layer=POLY_cond $X=0.495 $Y=1.557
+ $X2=0.51 $Y2=1.557
r92 37 51 11.1224 $w=4.28e-07 $l=4.15e-07 $layer=LI1_cond $X=1.68 $Y=1.565
+ $X2=1.265 $Y2=1.565
r93 36 51 1.74206 $w=4.28e-07 $l=6.5e-08 $layer=LI1_cond $X=1.2 $Y=1.565
+ $X2=1.265 $Y2=1.565
r94 35 36 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=1.2 $Y2=1.565
r95 35 46 3.61813 $w=4.28e-07 $l=1.35e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=0.585 $Y2=1.565
r96 34 46 9.24634 $w=4.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.24 $Y=1.565
+ $X2=0.585 $Y2=1.565
r97 29 33 18.8402 $w=1.65e-07 $l=8.21584e-08 $layer=POLY_cond $X=1.925 $Y=1.35
+ $X2=1.91 $Y2=1.425
r98 29 31 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=1.925 $Y=1.35
+ $X2=1.925 $Y2=0.78
r99 26 28 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.91 $Y=1.765
+ $X2=1.91 $Y2=2.4
r100 25 26 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.91 $Y=1.675
+ $X2=1.91 $Y2=1.765
r101 24 33 18.8402 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=1.91 $Y=1.5
+ $X2=1.91 $Y2=1.425
r102 24 25 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=1.91 $Y=1.5
+ $X2=1.91 $Y2=1.675
r103 23 53 27.4257 $w=3.72e-07 $l=1.653e-07 $layer=POLY_cond $X=1.5 $Y=1.425
+ $X2=1.425 $Y2=1.557
r104 22 33 6.66866 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=1.82 $Y=1.425
+ $X2=1.91 $Y2=1.425
r105 22 23 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.82 $Y=1.425
+ $X2=1.5 $Y2=1.425
r106 18 53 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.425 $Y=1.35
+ $X2=1.425 $Y2=1.557
r107 18 20 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=1.425 $Y=1.35
+ $X2=1.425 $Y2=0.78
r108 15 52 24.0971 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.41 $Y=1.765
+ $X2=1.41 $Y2=1.557
r109 15 17 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.41 $Y=1.765
+ $X2=1.41 $Y2=2.4
r110 11 48 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.995 $Y=1.35
+ $X2=0.995 $Y2=1.557
r111 11 13 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=0.995 $Y=1.35
+ $X2=0.995 $Y2=0.78
r112 8 47 24.0971 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.96 $Y=1.765
+ $X2=0.96 $Y2=1.557
r113 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.96 $Y=1.765
+ $X2=0.96 $Y2=2.4
r114 5 43 24.0971 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.51 $Y=1.765
+ $X2=0.51 $Y2=1.557
r115 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.51 $Y=1.765
+ $X2=0.51 $Y2=2.4
r116 1 42 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=1.557
r117 1 3 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=0.78
.ends

.subckt PM_SKY130_FD_SC_LS__O31AI_4%A2 3 5 7 8 10 12 15 17 19 22 24 25 28 30 32
+ 35 36 37
c93 30 0 9.50731e-20 $X=4.03 $Y=1.765
c94 28 0 2.00851e-19 $X=4.025 $Y=0.78
c95 25 0 9.74065e-20 $X=3.67 $Y=1.605
c96 17 0 7.17547e-20 $X=3.58 $Y=1.765
r97 49 50 2.00833 $w=3.6e-07 $l=1.5e-08 $layer=POLY_cond $X=3.58 $Y=1.557
+ $X2=3.595 $Y2=1.557
r98 47 49 10.0417 $w=3.6e-07 $l=7.5e-08 $layer=POLY_cond $X=3.505 $Y=1.557
+ $X2=3.58 $Y2=1.557
r99 47 48 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.505
+ $Y=1.515 $X2=3.505 $Y2=1.515
r100 45 47 54.8944 $w=3.6e-07 $l=4.1e-07 $layer=POLY_cond $X=3.095 $Y=1.557
+ $X2=3.505 $Y2=1.557
r101 44 45 31.4639 $w=3.6e-07 $l=2.35e-07 $layer=POLY_cond $X=2.86 $Y=1.557
+ $X2=3.095 $Y2=1.557
r102 42 44 4.68611 $w=3.6e-07 $l=3.5e-08 $layer=POLY_cond $X=2.825 $Y=1.557
+ $X2=2.86 $Y2=1.557
r103 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.825
+ $Y=1.515 $X2=2.825 $Y2=1.515
r104 37 48 2.54609 $w=4.28e-07 $l=9.5e-08 $layer=LI1_cond $X=3.6 $Y=1.565
+ $X2=3.505 $Y2=1.565
r105 36 48 10.3184 $w=4.28e-07 $l=3.85e-07 $layer=LI1_cond $X=3.12 $Y=1.565
+ $X2=3.505 $Y2=1.565
r106 36 43 7.90629 $w=4.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.12 $Y=1.565
+ $X2=2.825 $Y2=1.565
r107 35 43 4.95819 $w=4.28e-07 $l=1.85e-07 $layer=LI1_cond $X=2.64 $Y=1.565
+ $X2=2.825 $Y2=1.565
r108 30 34 48.1959 $w=1.61e-07 $l=1.63951e-07 $layer=POLY_cond $X=4.03 $Y=1.765
+ $X2=4.022 $Y2=1.605
r109 30 32 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.03 $Y=1.765
+ $X2=4.03 $Y2=2.4
r110 26 34 22.7487 $w=1.61e-07 $l=7.64853e-08 $layer=POLY_cond $X=4.025 $Y=1.53
+ $X2=4.022 $Y2=1.605
r111 26 28 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=4.025 $Y=1.53
+ $X2=4.025 $Y2=0.78
r112 25 50 26.8603 $w=3.6e-07 $l=9.60469e-08 $layer=POLY_cond $X=3.67 $Y=1.605
+ $X2=3.595 $Y2=1.557
r113 24 34 4.52116 $w=1.5e-07 $l=8.2e-08 $layer=POLY_cond $X=3.94 $Y=1.605
+ $X2=4.022 $Y2=1.605
r114 24 25 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=3.94 $Y=1.605
+ $X2=3.67 $Y2=1.605
r115 20 50 23.3057 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.595 $Y=1.35
+ $X2=3.595 $Y2=1.557
r116 20 22 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=3.595 $Y=1.35
+ $X2=3.595 $Y2=0.78
r117 17 49 23.3057 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.58 $Y=1.765
+ $X2=3.58 $Y2=1.557
r118 17 19 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.58 $Y=1.765
+ $X2=3.58 $Y2=2.4
r119 13 45 23.3057 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.095 $Y=1.35
+ $X2=3.095 $Y2=1.557
r120 13 15 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=3.095 $Y=1.35
+ $X2=3.095 $Y2=0.78
r121 10 44 23.3057 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.86 $Y=1.765
+ $X2=2.86 $Y2=1.557
r122 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.86 $Y=1.765
+ $X2=2.86 $Y2=2.4
r123 9 33 6.61437 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.45 $Y=1.425 $X2=2.36
+ $Y2=1.425
r124 8 42 38.9103 $w=3.6e-07 $l=2.21371e-07 $layer=POLY_cond $X=2.66 $Y=1.425
+ $X2=2.825 $Y2=1.557
r125 8 9 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=2.66 $Y=1.425
+ $X2=2.45 $Y2=1.425
r126 5 33 94.3029 $w=1.76e-07 $l=3.4e-07 $layer=POLY_cond $X=2.36 $Y=1.765
+ $X2=2.36 $Y2=1.425
r127 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.36 $Y=1.765
+ $X2=2.36 $Y2=2.4
r128 1 33 21.729 $w=1.76e-07 $l=7.74597e-08 $layer=POLY_cond $X=2.355 $Y=1.35
+ $X2=2.36 $Y2=1.425
r129 1 3 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=2.355 $Y=1.35
+ $X2=2.355 $Y2=0.78
.ends

.subckt PM_SKY130_FD_SC_LS__O31AI_4%A3 3 5 6 7 9 12 14 16 19 21 23 24 25 28 30
+ 32 34 35 36
c98 36 0 6.72563e-20 $X=6 $Y=1.665
c99 30 0 5.61847e-20 $X=6.44 $Y=1.765
c100 28 0 1.19111e-20 $X=6.425 $Y=0.78
c101 21 0 1.54703e-20 $X=5.99 $Y=1.765
c102 3 0 1.61283e-19 $X=4.455 $Y=0.78
r103 49 50 22.8534 $w=3.48e-07 $l=1.65e-07 $layer=POLY_cond $X=5.825 $Y=1.557
+ $X2=5.99 $Y2=1.557
r104 47 49 20.0833 $w=3.48e-07 $l=1.45e-07 $layer=POLY_cond $X=5.68 $Y=1.557
+ $X2=5.825 $Y2=1.557
r105 47 48 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=5.68
+ $Y=1.515 $X2=5.68 $Y2=1.515
r106 45 47 19.3908 $w=3.48e-07 $l=1.4e-07 $layer=POLY_cond $X=5.54 $Y=1.557
+ $X2=5.68 $Y2=1.557
r107 44 45 20.0833 $w=3.48e-07 $l=1.45e-07 $layer=POLY_cond $X=5.395 $Y=1.557
+ $X2=5.54 $Y2=1.557
r108 43 44 42.2443 $w=3.48e-07 $l=3.05e-07 $layer=POLY_cond $X=5.09 $Y=1.557
+ $X2=5.395 $Y2=1.557
r109 41 43 12.4655 $w=3.48e-07 $l=9e-08 $layer=POLY_cond $X=5 $Y=1.557 $X2=5.09
+ $Y2=1.557
r110 41 42 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=5
+ $Y=1.515 $X2=5 $Y2=1.515
r111 36 48 8.57632 $w=4.28e-07 $l=3.2e-07 $layer=LI1_cond $X=6 $Y=1.565 $X2=5.68
+ $Y2=1.565
r112 35 48 4.28816 $w=4.28e-07 $l=1.6e-07 $layer=LI1_cond $X=5.52 $Y=1.565
+ $X2=5.68 $Y2=1.565
r113 34 35 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=5.04 $Y=1.565
+ $X2=5.52 $Y2=1.565
r114 34 42 1.07204 $w=4.28e-07 $l=4e-08 $layer=LI1_cond $X=5.04 $Y=1.565 $X2=5
+ $Y2=1.565
r115 30 33 64.4713 $w=1.57e-07 $l=2.13963e-07 $layer=POLY_cond $X=6.44 $Y=1.765
+ $X2=6.432 $Y2=1.555
r116 30 32 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.44 $Y=1.765
+ $X2=6.44 $Y2=2.4
r117 26 33 23.0255 $w=1.57e-07 $l=7.84219e-08 $layer=POLY_cond $X=6.425 $Y=1.48
+ $X2=6.432 $Y2=1.555
r118 26 28 358.936 $w=1.5e-07 $l=7e-07 $layer=POLY_cond $X=6.425 $Y=1.48
+ $X2=6.425 $Y2=0.78
r119 25 50 28.3733 $w=3.48e-07 $l=9.09945e-08 $layer=POLY_cond $X=6.08 $Y=1.555
+ $X2=5.99 $Y2=1.557
r120 24 33 3.92347 $w=1.5e-07 $l=8.2e-08 $layer=POLY_cond $X=6.35 $Y=1.555
+ $X2=6.432 $Y2=1.555
r121 24 25 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=6.35 $Y=1.555
+ $X2=6.08 $Y2=1.555
r122 21 50 22.4912 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=5.99 $Y=1.765
+ $X2=5.99 $Y2=1.557
r123 21 23 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.99 $Y=1.765
+ $X2=5.99 $Y2=2.4
r124 17 49 22.4912 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.825 $Y=1.35
+ $X2=5.825 $Y2=1.557
r125 17 19 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=5.825 $Y=1.35
+ $X2=5.825 $Y2=0.78
r126 14 45 22.4912 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=5.54 $Y=1.765
+ $X2=5.54 $Y2=1.557
r127 14 16 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.54 $Y=1.765
+ $X2=5.54 $Y2=2.4
r128 10 44 22.4912 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.395 $Y=1.35
+ $X2=5.395 $Y2=1.557
r129 10 12 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=5.395 $Y=1.35
+ $X2=5.395 $Y2=0.78
r130 7 43 22.4912 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=5.09 $Y=1.765
+ $X2=5.09 $Y2=1.557
r131 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.09 $Y=1.765
+ $X2=5.09 $Y2=2.4
r132 5 41 38.7612 $w=3.48e-07 $l=2.21371e-07 $layer=POLY_cond $X=4.835 $Y=1.425
+ $X2=5 $Y2=1.557
r133 5 6 156.394 $w=1.5e-07 $l=3.05e-07 $layer=POLY_cond $X=4.835 $Y=1.425
+ $X2=4.53 $Y2=1.425
r134 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.455 $Y=1.35
+ $X2=4.53 $Y2=1.425
r135 1 3 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=4.455 $Y=1.35
+ $X2=4.455 $Y2=0.78
.ends

.subckt PM_SKY130_FD_SC_LS__O31AI_4%B1 3 5 7 10 14 16 17 18 19 20 22 23 25 27 28
+ 29 41
c68 41 0 1.54703e-20 $X=7.625 $Y=1.515
c69 17 0 6.72563e-20 $X=7.79 $Y=1.425
r70 40 42 12.5739 $w=3.45e-07 $l=9e-08 $layer=POLY_cond $X=7.625 $Y=1.557
+ $X2=7.715 $Y2=1.557
r71 40 41 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.625
+ $Y=1.515 $X2=7.625 $Y2=1.515
r72 38 40 47.5014 $w=3.45e-07 $l=3.4e-07 $layer=POLY_cond $X=7.285 $Y=1.557
+ $X2=7.625 $Y2=1.557
r73 36 38 47.5014 $w=3.45e-07 $l=3.4e-07 $layer=POLY_cond $X=6.945 $Y=1.557
+ $X2=7.285 $Y2=1.557
r74 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.945
+ $Y=1.515 $X2=6.945 $Y2=1.515
r75 34 36 0.698551 $w=3.45e-07 $l=5e-09 $layer=POLY_cond $X=6.94 $Y=1.557
+ $X2=6.945 $Y2=1.557
r76 33 34 11.8754 $w=3.45e-07 $l=8.5e-08 $layer=POLY_cond $X=6.855 $Y=1.557
+ $X2=6.94 $Y2=1.557
r77 29 41 4.95819 $w=4.28e-07 $l=1.85e-07 $layer=LI1_cond $X=7.44 $Y=1.565
+ $X2=7.625 $Y2=1.565
r78 28 29 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=6.96 $Y=1.565
+ $X2=7.44 $Y2=1.565
r79 28 37 0.402015 $w=4.28e-07 $l=1.5e-08 $layer=LI1_cond $X=6.96 $Y=1.565
+ $X2=6.945 $Y2=1.565
r80 27 37 12.4625 $w=4.28e-07 $l=4.65e-07 $layer=LI1_cond $X=6.48 $Y=1.565
+ $X2=6.945 $Y2=1.565
r81 23 26 58.0459 $w=1.68e-07 $l=2.04939e-07 $layer=POLY_cond $X=8.145 $Y=1.225
+ $X2=8.135 $Y2=1.425
r82 23 25 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=8.145 $Y=1.225
+ $X2=8.145 $Y2=0.78
r83 20 22 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.135 $Y=1.765
+ $X2=8.135 $Y2=2.4
r84 19 20 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=8.135 $Y=1.675
+ $X2=8.135 $Y2=1.765
r85 18 26 20.3659 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=8.135 $Y=1.5
+ $X2=8.135 $Y2=1.425
r86 18 19 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=8.135 $Y=1.5
+ $X2=8.135 $Y2=1.675
r87 17 42 26.1549 $w=3.45e-07 $l=1.653e-07 $layer=POLY_cond $X=7.79 $Y=1.425
+ $X2=7.715 $Y2=1.557
r88 16 26 5.52526 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=8.045 $Y=1.425
+ $X2=8.135 $Y2=1.425
r89 16 17 130.755 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=8.045 $Y=1.425
+ $X2=7.79 $Y2=1.425
r90 12 42 22.2839 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.715 $Y=1.35
+ $X2=7.715 $Y2=1.557
r91 12 14 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=7.715 $Y=1.35
+ $X2=7.715 $Y2=0.78
r92 8 38 22.2839 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.285 $Y=1.35
+ $X2=7.285 $Y2=1.557
r93 8 10 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=7.285 $Y=1.35
+ $X2=7.285 $Y2=0.78
r94 5 34 22.2839 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=6.94 $Y=1.765
+ $X2=6.94 $Y2=1.557
r95 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.94 $Y=1.765
+ $X2=6.94 $Y2=2.4
r96 1 33 22.2839 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.855 $Y=1.35
+ $X2=6.855 $Y2=1.557
r97 1 3 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=6.855 $Y=1.35
+ $X2=6.855 $Y2=0.78
.ends

.subckt PM_SKY130_FD_SC_LS__O31AI_4%A_28_368# 1 2 3 4 5 16 18 20 24 26 30 32 34
+ 35 36 41 43 46 50
c77 43 0 1.1776e-19 $X=2.135 $Y=1.985
c78 26 0 1.91457e-19 $X=1.97 $Y=2.035
r79 50 53 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=4.305 $Y=2.455
+ $X2=4.305 $Y2=2.55
r80 46 48 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=3.135 $Y=2.455
+ $X2=3.135 $Y2=2.57
r81 37 46 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.3 $Y=2.455
+ $X2=3.135 $Y2=2.455
r82 36 50 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.14 $Y=2.455
+ $X2=4.305 $Y2=2.455
r83 36 37 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=4.14 $Y=2.455
+ $X2=3.3 $Y2=2.455
r84 35 46 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=3.135 $Y=2.37
+ $X2=3.135 $Y2=2.455
r85 34 45 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.135 $Y=2.12
+ $X2=3.135 $Y2=2.035
r86 34 35 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=3.135 $Y=2.12
+ $X2=3.135 $Y2=2.37
r87 33 43 8.61065 $w=1.7e-07 $l=1.94808e-07 $layer=LI1_cond $X=2.3 $Y=2.035
+ $X2=2.135 $Y2=1.97
r88 32 45 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.97 $Y=2.035
+ $X2=3.135 $Y2=2.035
r89 32 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.97 $Y=2.035
+ $X2=2.3 $Y2=2.035
r90 28 43 0.89609 $w=3.3e-07 $l=1.5e-07 $layer=LI1_cond $X=2.135 $Y=2.12
+ $X2=2.135 $Y2=1.97
r91 28 30 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=2.135 $Y=2.12
+ $X2=2.135 $Y2=2.815
r92 27 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.27 $Y=2.035
+ $X2=1.185 $Y2=2.035
r93 26 43 8.61065 $w=1.7e-07 $l=1.94808e-07 $layer=LI1_cond $X=1.97 $Y=2.035
+ $X2=2.135 $Y2=1.97
r94 26 27 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.97 $Y=2.035 $X2=1.27
+ $Y2=2.035
r95 22 41 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=2.12
+ $X2=1.185 $Y2=2.035
r96 22 24 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=1.185 $Y=2.12
+ $X2=1.185 $Y2=2.815
r97 21 39 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.37 $Y=2.035
+ $X2=0.245 $Y2=2.035
r98 20 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=2.035
+ $X2=1.185 $Y2=2.035
r99 20 21 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.1 $Y=2.035
+ $X2=0.37 $Y2=2.035
r100 16 39 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.245 $Y=2.12
+ $X2=0.245 $Y2=2.035
r101 16 18 32.0379 $w=2.48e-07 $l=6.95e-07 $layer=LI1_cond $X=0.245 $Y=2.12
+ $X2=0.245 $Y2=2.815
r102 5 53 600 $w=1.7e-07 $l=8.03803e-07 $layer=licon1_PDIFF $count=1 $X=4.105
+ $Y=1.84 $X2=4.305 $Y2=2.55
r103 4 48 600 $w=1.7e-07 $l=8.23954e-07 $layer=licon1_PDIFF $count=1 $X=2.935
+ $Y=1.84 $X2=3.135 $Y2=2.57
r104 4 45 600 $w=1.7e-07 $l=3.61421e-07 $layer=licon1_PDIFF $count=1 $X=2.935
+ $Y=1.84 $X2=3.135 $Y2=2.115
r105 3 43 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.985
+ $Y=1.84 $X2=2.135 $Y2=1.985
r106 3 30 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.985
+ $Y=1.84 $X2=2.135 $Y2=2.815
r107 2 41 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=1.035
+ $Y=1.84 $X2=1.185 $Y2=2.115
r108 2 24 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.035
+ $Y=1.84 $X2=1.185 $Y2=2.815
r109 1 39 400 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.14
+ $Y=1.84 $X2=0.285 $Y2=2.115
r110 1 18 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.14
+ $Y=1.84 $X2=0.285 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_LS__O31AI_4%VPWR 1 2 3 12 16 18 20 25 30 40 41 44 47 50
r84 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r85 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r86 41 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=7.92 $Y2=3.33
r87 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33 $X2=8.4
+ $Y2=3.33
r88 38 40 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=8.025 $Y=3.33
+ $X2=8.4 $Y2=3.33
r89 37 55 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.92 $Y2=3.33
r90 36 37 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r91 34 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r92 33 36 313.155 $w=1.68e-07 $l=4.8e-06 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=6.96 $Y2=3.33
r93 33 34 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r94 31 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.8 $Y=3.33
+ $X2=1.635 $Y2=3.33
r95 31 33 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=1.8 $Y=3.33 $X2=2.16
+ $Y2=3.33
r96 30 38 11.5506 $w=1.7e-07 $l=4.88e-07 $layer=LI1_cond $X=7.537 $Y=3.33
+ $X2=8.025 $Y2=3.33
r97 30 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r98 30 50 10.9487 $w=9.73e-07 $l=8.75e-07 $layer=LI1_cond $X=7.537 $Y=3.33
+ $X2=7.537 $Y2=2.455
r99 30 36 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=7.05 $Y=3.33 $X2=6.96
+ $Y2=3.33
r100 29 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r101 29 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r102 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r103 26 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.9 $Y=3.33
+ $X2=0.735 $Y2=3.33
r104 26 28 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=0.9 $Y=3.33 $X2=1.2
+ $Y2=3.33
r105 25 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.47 $Y=3.33
+ $X2=1.635 $Y2=3.33
r106 25 28 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=1.47 $Y=3.33 $X2=1.2
+ $Y2=3.33
r107 23 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r108 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r109 20 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.57 $Y=3.33
+ $X2=0.735 $Y2=3.33
r110 20 22 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.57 $Y=3.33
+ $X2=0.24 $Y2=3.33
r111 18 37 0.73586 $w=4.9e-07 $l=2.64e-06 $layer=MET1_cond $X=4.32 $Y=3.33
+ $X2=6.96 $Y2=3.33
r112 18 34 0.602067 $w=4.9e-07 $l=2.16e-06 $layer=MET1_cond $X=4.32 $Y=3.33
+ $X2=2.16 $Y2=3.33
r113 14 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.635 $Y=3.245
+ $X2=1.635 $Y2=3.33
r114 14 16 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=1.635 $Y=3.245
+ $X2=1.635 $Y2=2.455
r115 10 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.735 $Y=3.245
+ $X2=0.735 $Y2=3.33
r116 10 12 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=0.735 $Y=3.245
+ $X2=0.735 $Y2=2.455
r117 3 50 200 $w=1.7e-07 $l=1.16252e-06 $layer=licon1_PDIFF $count=3 $X=7.015
+ $Y=1.84 $X2=7.91 $Y2=2.455
r118 3 50 200 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=3 $X=7.015
+ $Y=1.84 $X2=7.165 $Y2=2.455
r119 2 16 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=1.485
+ $Y=1.84 $X2=1.635 $Y2=2.455
r120 1 12 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.84 $X2=0.735 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_LS__O31AI_4%A_487_368# 1 2 3 4 15 17 18 19 23 25 29 32
+ 36
c59 19 0 7.17547e-20 $X=5.15 $Y=2.99
c60 17 0 7.17547e-20 $X=3.64 $Y=2.99
r61 32 34 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=3.805 $Y=2.805
+ $X2=3.805 $Y2=2.99
r62 27 29 20.744 $w=2.48e-07 $l=4.5e-07 $layer=LI1_cond $X=6.255 $Y=2.905
+ $X2=6.255 $Y2=2.455
r63 26 36 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.4 $Y=2.99
+ $X2=5.275 $Y2=2.99
r64 25 27 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.13 $Y=2.99
+ $X2=6.255 $Y2=2.905
r65 25 26 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=6.13 $Y=2.99 $X2=5.4
+ $Y2=2.99
r66 21 36 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.275 $Y=2.905
+ $X2=5.275 $Y2=2.99
r67 21 23 20.744 $w=2.48e-07 $l=4.5e-07 $layer=LI1_cond $X=5.275 $Y=2.905
+ $X2=5.275 $Y2=2.455
r68 20 34 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.97 $Y=2.99
+ $X2=3.805 $Y2=2.99
r69 19 36 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.15 $Y=2.99
+ $X2=5.275 $Y2=2.99
r70 19 20 76.984 $w=1.68e-07 $l=1.18e-06 $layer=LI1_cond $X=5.15 $Y=2.99
+ $X2=3.97 $Y2=2.99
r71 17 34 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.64 $Y=2.99
+ $X2=3.805 $Y2=2.99
r72 17 18 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=3.64 $Y=2.99 $X2=2.8
+ $Y2=2.99
r73 13 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.635 $Y=2.905
+ $X2=2.8 $Y2=2.99
r74 13 15 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=2.635 $Y=2.905
+ $X2=2.635 $Y2=2.455
r75 4 29 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=6.065
+ $Y=1.84 $X2=6.215 $Y2=2.455
r76 3 23 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=5.165
+ $Y=1.84 $X2=5.315 $Y2=2.455
r77 2 32 600 $w=1.7e-07 $l=1.03729e-06 $layer=licon1_PDIFF $count=1 $X=3.655
+ $Y=1.84 $X2=3.805 $Y2=2.805
r78 1 15 300 $w=1.7e-07 $l=7.07972e-07 $layer=licon1_PDIFF $count=2 $X=2.435
+ $Y=1.84 $X2=2.635 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_LS__O31AI_4%Y 1 2 3 4 5 6 20 22 25 27 28 31 35 37 39 43
+ 45 47 50 52 53 56
c116 53 0 5.61847e-20 $X=6.905 $Y=1.05
c117 28 0 9.74065e-20 $X=4.97 $Y=2.035
c118 22 0 6.10557e-20 $X=4.665 $Y=1.095
r119 56 63 12.7615 $w=4.78e-07 $l=5e-07 $layer=LI1_cond $X=4.08 $Y=1.85 $X2=4.58
+ $Y2=1.85
r120 45 55 3.0656 $w=3.3e-07 $l=1.5e-07 $layer=LI1_cond $X=8.36 $Y=2.12 $X2=8.36
+ $Y2=1.97
r121 45 47 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=8.36 $Y=2.12
+ $X2=8.36 $Y2=2.815
r122 41 43 38.1193 $w=2.58e-07 $l=8.6e-07 $layer=LI1_cond $X=7.07 $Y=1.05
+ $X2=7.93 $Y2=1.05
r123 39 53 7.14225 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=7.035 $Y=1.05
+ $X2=6.905 $Y2=1.05
r124 39 41 1.55137 $w=2.58e-07 $l=3.5e-08 $layer=LI1_cond $X=7.035 $Y=1.05
+ $X2=7.07 $Y2=1.05
r125 38 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.88 $Y=2.035
+ $X2=6.715 $Y2=2.035
r126 37 55 4.70058 $w=1.7e-07 $l=1.94808e-07 $layer=LI1_cond $X=8.195 $Y=2.035
+ $X2=8.36 $Y2=1.97
r127 37 38 85.7914 $w=1.68e-07 $l=1.315e-06 $layer=LI1_cond $X=8.195 $Y=2.035
+ $X2=6.88 $Y2=2.035
r128 33 52 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.715 $Y=2.12
+ $X2=6.715 $Y2=2.035
r129 33 35 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=6.715 $Y=2.12
+ $X2=6.715 $Y2=2.815
r130 32 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.93 $Y=2.035
+ $X2=5.765 $Y2=2.035
r131 31 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.55 $Y=2.035
+ $X2=6.715 $Y2=2.035
r132 31 32 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=6.55 $Y=2.035
+ $X2=5.93 $Y2=2.035
r133 28 66 8.0408 $w=4.78e-07 $l=1.05e-07 $layer=LI1_cond $X=4.97 $Y=2.035
+ $X2=4.865 $Y2=2.035
r134 27 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.6 $Y=2.035
+ $X2=5.765 $Y2=2.035
r135 27 28 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=5.6 $Y=2.035
+ $X2=4.97 $Y2=2.035
r136 23 66 0.76569 $w=4.78e-07 $l=1.29132e-07 $layer=LI1_cond $X=4.835 $Y=2.15
+ $X2=4.865 $Y2=2.035
r137 23 63 6.50837 $w=4.78e-07 $l=4.08044e-07 $layer=LI1_cond $X=4.835 $Y=2.15
+ $X2=4.58 $Y2=1.85
r138 23 25 17.9269 $w=2.68e-07 $l=4.2e-07 $layer=LI1_cond $X=4.835 $Y=2.15
+ $X2=4.835 $Y2=2.57
r139 22 53 146.139 $w=1.68e-07 $l=2.24e-06 $layer=LI1_cond $X=4.665 $Y=1.095
+ $X2=6.905 $Y2=1.095
r140 20 63 6.87511 $w=1.7e-07 $l=3e-07 $layer=LI1_cond $X=4.58 $Y=1.55 $X2=4.58
+ $Y2=1.85
r141 19 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.58 $Y=1.18
+ $X2=4.665 $Y2=1.095
r142 19 20 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=4.58 $Y=1.18
+ $X2=4.58 $Y2=1.55
r143 6 55 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=8.21
+ $Y=1.84 $X2=8.36 $Y2=1.985
r144 6 47 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=8.21
+ $Y=1.84 $X2=8.36 $Y2=2.815
r145 5 52 400 $w=1.7e-07 $l=3.61421e-07 $layer=licon1_PDIFF $count=1 $X=6.515
+ $Y=1.84 $X2=6.715 $Y2=2.115
r146 5 35 400 $w=1.7e-07 $l=1.07034e-06 $layer=licon1_PDIFF $count=1 $X=6.515
+ $Y=1.84 $X2=6.715 $Y2=2.815
r147 4 50 300 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=2 $X=5.615
+ $Y=1.84 $X2=5.765 $Y2=2.115
r148 3 66 600 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=1 $X=4.72
+ $Y=1.84 $X2=4.865 $Y2=2.035
r149 3 25 600 $w=1.7e-07 $l=7.99218e-07 $layer=licon1_PDIFF $count=1 $X=4.72
+ $Y=1.84 $X2=4.865 $Y2=2.57
r150 2 43 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=7.79
+ $Y=0.41 $X2=7.93 $Y2=1.005
r151 1 41 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=6.93
+ $Y=0.41 $X2=7.07 $Y2=1.005
.ends

.subckt PM_SKY130_FD_SC_LS__O31AI_4%A_27_82# 1 2 3 4 5 6 7 8 9 30 32 33 38 40 44
+ 46 50 58 62 66 68 69 73 74 75 83 84
c130 83 0 1.19111e-20 $X=7.335 $Y=0.57
c131 50 0 3.01078e-19 $X=4.24 $Y=0.555
c132 46 0 2.33185e-20 $X=4.155 $Y=1.095
c133 32 0 1.1776e-19 $X=1.975 $Y=1.05
r134 82 84 8.51103 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=7.5 $Y=0.57
+ $X2=7.665 $Y2=0.57
r135 82 83 8.51103 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=7.5 $Y=0.57
+ $X2=7.335 $Y2=0.57
r136 78 79 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=6.64 $Y=0.57
+ $X2=6.64 $Y2=0.665
r137 75 78 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=6.64 $Y=0.475
+ $X2=6.64 $Y2=0.57
r138 72 74 9.22412 $w=4.48e-07 $l=1.65e-07 $layer=LI1_cond $X=5.61 $Y=0.615
+ $X2=5.775 $Y2=0.615
r139 72 73 9.22412 $w=4.48e-07 $l=1.65e-07 $layer=LI1_cond $X=5.61 $Y=0.615
+ $X2=5.445 $Y2=0.615
r140 64 66 0.443247 $w=2.58e-07 $l=1e-08 $layer=LI1_cond $X=8.395 $Y=0.56
+ $X2=8.395 $Y2=0.57
r141 62 64 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=8.265 $Y=0.475
+ $X2=8.395 $Y2=0.56
r142 62 84 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=8.265 $Y=0.475
+ $X2=7.665 $Y2=0.475
r143 61 75 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.805 $Y=0.475
+ $X2=6.64 $Y2=0.475
r144 61 83 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=6.805 $Y=0.475
+ $X2=7.335 $Y2=0.475
r145 58 79 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.475 $Y=0.665
+ $X2=6.64 $Y2=0.665
r146 58 74 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=6.475 $Y=0.665
+ $X2=5.775 $Y2=0.665
r147 57 70 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.325 $Y=0.755
+ $X2=4.24 $Y2=0.755
r148 57 73 73.0695 $w=1.68e-07 $l=1.12e-06 $layer=LI1_cond $X=4.325 $Y=0.755
+ $X2=5.445 $Y2=0.755
r149 53 55 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=4.24 $Y=1.01
+ $X2=4.24 $Y2=1.005
r150 52 70 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.24 $Y=0.84
+ $X2=4.24 $Y2=0.755
r151 52 55 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=4.24 $Y=0.84
+ $X2=4.24 $Y2=1.005
r152 48 70 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.24 $Y=0.67
+ $X2=4.24 $Y2=0.755
r153 48 50 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=4.24 $Y=0.67
+ $X2=4.24 $Y2=0.555
r154 47 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.475 $Y=1.095
+ $X2=3.31 $Y2=1.095
r155 46 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.155 $Y=1.095
+ $X2=4.24 $Y2=1.01
r156 46 47 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.155 $Y=1.095
+ $X2=3.475 $Y2=1.095
r157 42 69 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.31 $Y=1.01
+ $X2=3.31 $Y2=1.095
r158 42 44 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=3.31 $Y=1.01
+ $X2=3.31 $Y2=0.555
r159 41 68 7.25953 $w=2.15e-07 $l=1.86145e-07 $layer=LI1_cond $X=2.305 $Y=1.095
+ $X2=2.14 $Y2=1.05
r160 40 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.145 $Y=1.095
+ $X2=3.31 $Y2=1.095
r161 40 41 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=3.145 $Y=1.095
+ $X2=2.305 $Y2=1.095
r162 36 68 0.144206 $w=3.3e-07 $l=1.3e-07 $layer=LI1_cond $X=2.14 $Y=0.92
+ $X2=2.14 $Y2=1.05
r163 36 38 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=2.14 $Y=0.92
+ $X2=2.14 $Y2=0.555
r164 33 35 33.9084 $w=2.58e-07 $l=7.65e-07 $layer=LI1_cond $X=0.445 $Y=1.05
+ $X2=1.21 $Y2=1.05
r165 32 68 7.25953 $w=2.15e-07 $l=1.65e-07 $layer=LI1_cond $X=1.975 $Y=1.05
+ $X2=2.14 $Y2=1.05
r166 32 35 33.9084 $w=2.58e-07 $l=7.65e-07 $layer=LI1_cond $X=1.975 $Y=1.05
+ $X2=1.21 $Y2=1.05
r167 28 33 6.94204 $w=2.6e-07 $l=2.20624e-07 $layer=LI1_cond $X=0.28 $Y=0.92
+ $X2=0.445 $Y2=1.05
r168 28 30 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=0.28 $Y=0.92
+ $X2=0.28 $Y2=0.555
r169 9 66 91 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=2 $X=8.22
+ $Y=0.41 $X2=8.36 $Y2=0.57
r170 8 82 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=7.36
+ $Y=0.41 $X2=7.5 $Y2=0.57
r171 7 78 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=6.5
+ $Y=0.41 $X2=6.64 $Y2=0.57
r172 6 72 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=5.47
+ $Y=0.41 $X2=5.61 $Y2=0.615
r173 5 55 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=4.1
+ $Y=0.41 $X2=4.24 $Y2=1.005
r174 5 50 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=4.1
+ $Y=0.41 $X2=4.24 $Y2=0.555
r175 4 44 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.17
+ $Y=0.41 $X2=3.31 $Y2=0.555
r176 3 38 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2 $Y=0.41
+ $X2=2.14 $Y2=0.555
r177 2 35 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=1.07
+ $Y=0.41 $X2=1.21 $Y2=1.005
r178 1 30 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.41 $X2=0.28 $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_LS__O31AI_4%VGND 1 2 3 4 5 6 21 25 29 33 35 38 39 40 42
+ 47 52 70 71 74 77 80 85 88 91
r113 91 94 11.016 $w=3.38e-07 $l=3.25e-07 $layer=LI1_cond $X=6.125 $Y=0
+ $X2=6.125 $Y2=0.325
r114 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6 $Y2=0
r115 87 88 10.0584 $w=5.83e-07 $l=1.65e-07 $layer=LI1_cond $X=5.1 $Y=0.207
+ $X2=5.265 $Y2=0.207
r116 84 92 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=6
+ $Y2=0
r117 83 87 1.22675 $w=5.83e-07 $l=6e-08 $layer=LI1_cond $X=5.04 $Y=0.207 $X2=5.1
+ $Y2=0.207
r118 83 85 15.9877 $w=5.83e-07 $l=4.55e-07 $layer=LI1_cond $X=5.04 $Y=0.207
+ $X2=4.585 $Y2=0.207
r119 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r120 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r121 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r122 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r123 70 71 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r124 68 71 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6.48 $Y=0 $X2=8.4
+ $Y2=0
r125 68 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r126 67 70 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=6.48 $Y=0 $X2=8.4
+ $Y2=0
r127 67 68 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r128 65 91 4.80115 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=6.295 $Y=0 $X2=6.125
+ $Y2=0
r129 65 67 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=6.295 $Y=0
+ $X2=6.48 $Y2=0
r130 64 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r131 63 85 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=4.56 $Y=0 $X2=4.585
+ $Y2=0
r132 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r133 60 81 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=2.64
+ $Y2=0
r134 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r135 57 80 10.8012 $w=1.7e-07 $l=2.33e-07 $layer=LI1_cond $X=2.96 $Y=0 $X2=2.727
+ $Y2=0
r136 57 59 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=2.96 $Y=0 $X2=3.6
+ $Y2=0
r137 56 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r138 56 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r139 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r140 53 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.805 $Y=0 $X2=1.64
+ $Y2=0
r141 53 55 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=1.805 $Y=0
+ $X2=2.16 $Y2=0
r142 52 80 10.8012 $w=1.7e-07 $l=2.32e-07 $layer=LI1_cond $X=2.495 $Y=0
+ $X2=2.727 $Y2=0
r143 52 55 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.495 $Y=0
+ $X2=2.16 $Y2=0
r144 51 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r145 51 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r146 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r147 48 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=0.78
+ $Y2=0
r148 48 50 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=1.2
+ $Y2=0
r149 47 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.475 $Y=0 $X2=1.64
+ $Y2=0
r150 47 50 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.475 $Y=0 $X2=1.2
+ $Y2=0
r151 45 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r152 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r153 42 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.78
+ $Y2=0
r154 42 44 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=0
+ $X2=0.24 $Y2=0
r155 40 64 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=0
+ $X2=4.56 $Y2=0
r156 40 60 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=4.32 $Y=0 $X2=3.6
+ $Y2=0
r157 38 59 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=3.645 $Y=0 $X2=3.6
+ $Y2=0
r158 38 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.645 $Y=0 $X2=3.81
+ $Y2=0
r159 37 63 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=3.975 $Y=0
+ $X2=4.56 $Y2=0
r160 37 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.975 $Y=0 $X2=3.81
+ $Y2=0
r161 35 91 4.80115 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=5.955 $Y=0 $X2=6.125
+ $Y2=0
r162 35 88 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.955 $Y=0 $X2=5.265
+ $Y2=0
r163 31 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.81 $Y=0.085
+ $X2=3.81 $Y2=0
r164 31 33 19.9058 $w=3.28e-07 $l=5.7e-07 $layer=LI1_cond $X=3.81 $Y=0.085
+ $X2=3.81 $Y2=0.655
r165 27 80 1.88438 $w=4.65e-07 $l=8.5e-08 $layer=LI1_cond $X=2.727 $Y=0.085
+ $X2=2.727 $Y2=0
r166 27 29 15.0474 $w=4.63e-07 $l=5.85e-07 $layer=LI1_cond $X=2.727 $Y=0.085
+ $X2=2.727 $Y2=0.67
r167 23 77 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.64 $Y=0.085
+ $X2=1.64 $Y2=0
r168 23 25 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=1.64 $Y=0.085
+ $X2=1.64 $Y2=0.57
r169 19 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=0.085
+ $X2=0.78 $Y2=0
r170 19 21 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=0.78 $Y=0.085
+ $X2=0.78 $Y2=0.57
r171 6 94 182 $w=1.7e-07 $l=2.64102e-07 $layer=licon1_NDIFF $count=1 $X=5.9
+ $Y=0.41 $X2=6.125 $Y2=0.325
r172 5 87 91 $w=1.7e-07 $l=6.06341e-07 $layer=licon1_NDIFF $count=2 $X=4.53
+ $Y=0.41 $X2=5.1 $Y2=0.335
r173 4 33 182 $w=1.7e-07 $l=3.07124e-07 $layer=licon1_NDIFF $count=1 $X=3.67
+ $Y=0.41 $X2=3.81 $Y2=0.655
r174 3 29 182 $w=1.7e-07 $l=4.04629e-07 $layer=licon1_NDIFF $count=1 $X=2.43
+ $Y=0.41 $X2=2.725 $Y2=0.67
r175 2 25 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=1.5
+ $Y=0.41 $X2=1.64 $Y2=0.57
r176 1 21 182 $w=1.7e-07 $l=2.78747e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.41 $X2=0.78 $Y2=0.57
.ends

