* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__dfxtp_4 CLK D VGND VNB VPB VPWR Q
M1000 Q a_1226_296# VGND VNB nshort w=740000u l=150000u
+  ad=4.44e+11p pd=4.16e+06u as=1.88282e+12p ps=1.54e+07u
M1001 a_1141_508# a_206_368# a_1034_424# VPB phighvt w=420000u l=150000u
+  ad=1.995e+11p pd=1.79e+06u as=2.856e+11p ps=2.45e+06u
M1002 Q a_1226_296# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=6.72e+11p pd=5.68e+06u as=2.4029e+12p ps=1.958e+07u
M1003 VPWR a_1034_424# a_1226_296# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=2.52e+11p ps=2.28e+06u
M1004 Q a_1226_296# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_696_458# a_544_485# VGND VNB nshort w=550000u l=150000u
+  ad=1.98e+11p pd=1.97e+06u as=0p ps=0u
M1006 a_651_503# a_27_74# a_544_485# VPB phighvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=1.7745e+11p ps=1.79e+06u
M1007 VPWR a_1226_296# Q VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_437_503# D VPWR VPB phighvt w=420000u l=150000u
+  ad=1.7745e+11p pd=1.79e+06u as=0p ps=0u
M1009 VPWR a_696_458# a_651_503# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_544_485# a_206_368# a_437_503# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND a_696_458# a_735_102# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1012 VGND a_1226_296# Q VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 Q a_1226_296# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND a_1226_296# a_1178_124# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.323e+11p ps=1.47e+06u
M1015 VPWR CLK a_27_74# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.304e+11p ps=2.83e+06u
M1016 a_206_368# a_27_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=0p ps=0u
M1017 a_735_102# a_206_368# a_544_485# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.51375e+11p ps=1.66e+06u
M1018 a_1034_424# a_27_74# a_696_458# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=4.452e+11p ps=2.74e+06u
M1019 a_437_503# D VGND VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1020 a_544_485# a_27_74# a_437_503# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_1034_424# a_206_368# a_696_458# VNB nshort w=550000u l=150000u
+  ad=2.152e+11p pd=1.97e+06u as=0p ps=0u
M1022 a_206_368# a_27_74# VGND VNB nshort w=740000u l=150000u
+  ad=2.516e+11p pd=2.16e+06u as=0p ps=0u
M1023 VPWR a_1226_296# a_1141_508# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND a_1034_424# a_1226_296# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1025 VGND CLK a_27_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1026 VPWR a_1226_296# Q VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_696_458# a_544_485# VPWR VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_1178_124# a_27_74# a_1034_424# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_1226_296# a_1034_424# VPWR VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VGND a_1226_296# Q VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
