* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
M1000 VPWR B1 a_84_48# VPB phighvt w=840000u l=150000u
+  ad=9.804e+11p pd=5.95e+06u as=3.748e+11p ps=2.78e+06u
M1001 a_230_94# A3 VGND VNB nshort w=640000u l=150000u
+  ad=4.48e+11p pd=3.96e+06u as=6.755e+11p ps=4.76e+06u
M1002 a_84_48# B1 a_230_94# VNB nshort w=640000u l=150000u
+  ad=2.272e+11p pd=1.99e+06u as=0p ps=0u
M1003 VGND A2 a_230_94# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR a_84_48# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.304e+11p ps=2.83e+06u
M1005 a_340_368# A2 a_256_368# VPB phighvt w=1e+06u l=150000u
+  ad=3.6e+11p pd=2.72e+06u as=2.7e+11p ps=2.54e+06u
M1006 a_84_48# A3 a_340_368# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_230_94# A1 VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND a_84_48# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1009 a_256_368# A1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
