* File: sky130_fd_sc_ls__o22a_2.pxi.spice
* Created: Fri Aug 28 13:48:43 2020
* 
x_PM_SKY130_FD_SC_LS__O22A_2%A_82_48# N_A_82_48#_M1002_d N_A_82_48#_M1004_d
+ N_A_82_48#_M1006_g N_A_82_48#_c_76_n N_A_82_48#_M1000_g N_A_82_48#_M1008_g
+ N_A_82_48#_c_77_n N_A_82_48#_M1003_g N_A_82_48#_c_69_n N_A_82_48#_c_70_n
+ N_A_82_48#_c_83_p N_A_82_48#_c_107_p N_A_82_48#_c_97_p N_A_82_48#_c_79_n
+ N_A_82_48#_c_71_n N_A_82_48#_c_72_n N_A_82_48#_c_73_n N_A_82_48#_c_74_n
+ N_A_82_48#_c_75_n PM_SKY130_FD_SC_LS__O22A_2%A_82_48#
x_PM_SKY130_FD_SC_LS__O22A_2%B1 N_B1_c_159_n N_B1_M1001_g N_B1_M1002_g B1
+ PM_SKY130_FD_SC_LS__O22A_2%B1
x_PM_SKY130_FD_SC_LS__O22A_2%B2 N_B2_c_192_n N_B2_M1004_g N_B2_M1011_g B2
+ N_B2_c_194_n PM_SKY130_FD_SC_LS__O22A_2%B2
x_PM_SKY130_FD_SC_LS__O22A_2%A2 N_A2_c_225_n N_A2_M1005_g N_A2_M1010_g A2
+ PM_SKY130_FD_SC_LS__O22A_2%A2
x_PM_SKY130_FD_SC_LS__O22A_2%A1 N_A1_c_257_n N_A1_M1009_g N_A1_M1007_g A1
+ N_A1_c_259_n PM_SKY130_FD_SC_LS__O22A_2%A1
x_PM_SKY130_FD_SC_LS__O22A_2%VPWR N_VPWR_M1000_d N_VPWR_M1003_d N_VPWR_M1009_d
+ N_VPWR_c_282_n N_VPWR_c_283_n N_VPWR_c_284_n N_VPWR_c_285_n N_VPWR_c_286_n
+ N_VPWR_c_287_n VPWR N_VPWR_c_288_n N_VPWR_c_289_n N_VPWR_c_281_n
+ PM_SKY130_FD_SC_LS__O22A_2%VPWR
x_PM_SKY130_FD_SC_LS__O22A_2%X N_X_M1006_d N_X_M1000_s N_X_c_324_n N_X_c_327_n
+ N_X_c_328_n N_X_c_325_n X PM_SKY130_FD_SC_LS__O22A_2%X
x_PM_SKY130_FD_SC_LS__O22A_2%VGND N_VGND_M1006_s N_VGND_M1008_s N_VGND_M1010_d
+ N_VGND_c_359_n N_VGND_c_360_n N_VGND_c_361_n N_VGND_c_362_n VGND
+ N_VGND_c_363_n N_VGND_c_364_n N_VGND_c_365_n N_VGND_c_366_n N_VGND_c_367_n
+ N_VGND_c_368_n PM_SKY130_FD_SC_LS__O22A_2%VGND
x_PM_SKY130_FD_SC_LS__O22A_2%A_307_74# N_A_307_74#_M1002_s N_A_307_74#_M1011_d
+ N_A_307_74#_M1007_d N_A_307_74#_c_409_n N_A_307_74#_c_410_n
+ N_A_307_74#_c_430_n N_A_307_74#_c_411_n N_A_307_74#_c_412_n
+ N_A_307_74#_c_413_n N_A_307_74#_c_414_n PM_SKY130_FD_SC_LS__O22A_2%A_307_74#
cc_1 VNB N_A_82_48#_M1006_g 0.0338946f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=0.74
cc_2 VNB N_A_82_48#_M1008_g 0.0232514f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=0.74
cc_3 VNB N_A_82_48#_c_69_n 4.10656e-19 $X=-0.19 $Y=-0.245 $X2=1.22 $Y2=1.95
cc_4 VNB N_A_82_48#_c_70_n 0.00178028f $X=-0.19 $Y=-0.245 $X2=1.305 $Y2=1.005
cc_5 VNB N_A_82_48#_c_71_n 0.00319769f $X=-0.19 $Y=-0.245 $X2=1.14 $Y2=1.465
cc_6 VNB N_A_82_48#_c_72_n 0.00341558f $X=-0.19 $Y=-0.245 $X2=1.14 $Y2=1.3
cc_7 VNB N_A_82_48#_c_73_n 0.00372536f $X=-0.19 $Y=-0.245 $X2=2.115 $Y2=0.965
cc_8 VNB N_A_82_48#_c_74_n 0.0223221f $X=-0.19 $Y=-0.245 $X2=2.005 $Y2=0.965
cc_9 VNB N_A_82_48#_c_75_n 0.0806606f $X=-0.19 $Y=-0.245 $X2=1.025 $Y2=1.532
cc_10 VNB N_B1_c_159_n 0.0258166f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=0.37
cc_11 VNB N_B1_M1002_g 0.033506f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB B1 0.0030524f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=0.74
cc_13 VNB N_B2_c_192_n 0.018703f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=0.37
cc_14 VNB N_B2_M1011_g 0.0306575f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_B2_c_194_n 0.00432046f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=2.4
cc_16 VNB N_A2_c_225_n 0.0175712f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=0.37
cc_17 VNB N_A2_M1010_g 0.0311199f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB A2 0.00517424f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=0.74
cc_19 VNB N_A1_c_257_n 0.0607532f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=0.37
cc_20 VNB N_A1_M1007_g 0.0300997f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A1_c_259_n 0.00431187f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=2.4
cc_22 VNB N_VPWR_c_281_n 0.163682f $X=-0.19 $Y=-0.245 $X2=1.14 $Y2=1.532
cc_23 VNB N_X_c_324_n 0.00210995f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=0.74
cc_24 VNB N_X_c_325_n 0.00432789f $X=-0.19 $Y=-0.245 $X2=1.025 $Y2=2.4
cc_25 VNB X 0.00435003f $X=-0.19 $Y=-0.245 $X2=1.025 $Y2=2.4
cc_26 VNB N_VGND_c_359_n 0.0105514f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_360_n 0.0506785f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=2.4
cc_28 VNB N_VGND_c_361_n 0.00898285f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=0.74
cc_29 VNB N_VGND_c_362_n 0.00640205f $X=-0.19 $Y=-0.245 $X2=1.025 $Y2=2.4
cc_30 VNB N_VGND_c_363_n 0.0168951f $X=-0.19 $Y=-0.245 $X2=1.22 $Y2=1.95
cc_31 VNB N_VGND_c_364_n 0.0430142f $X=-0.19 $Y=-0.245 $X2=2.515 $Y2=2.12
cc_32 VNB N_VGND_c_365_n 0.0173909f $X=-0.19 $Y=-0.245 $X2=2.115 $Y2=0.965
cc_33 VNB N_VGND_c_366_n 0.234729f $X=-0.19 $Y=-0.245 $X2=2.005 $Y2=0.965
cc_34 VNB N_VGND_c_367_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=1.532
cc_35 VNB N_VGND_c_368_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_307_74#_c_409_n 0.00296475f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_307_74#_c_410_n 0.00261637f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=2.4
cc_38 VNB N_A_307_74#_c_411_n 0.0128061f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=1.3
cc_39 VNB N_A_307_74#_c_412_n 0.00950245f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=0.74
cc_40 VNB N_A_307_74#_c_413_n 0.0247745f $X=-0.19 $Y=-0.245 $X2=1.025 $Y2=1.765
cc_41 VNB N_A_307_74#_c_414_n 0.00655754f $X=-0.19 $Y=-0.245 $X2=1.025 $Y2=2.4
cc_42 VPB N_A_82_48#_c_76_n 0.0174014f $X=-0.19 $Y=1.66 $X2=0.575 $Y2=1.765
cc_43 VPB N_A_82_48#_c_77_n 0.0174445f $X=-0.19 $Y=1.66 $X2=1.025 $Y2=1.765
cc_44 VPB N_A_82_48#_c_69_n 0.00302398f $X=-0.19 $Y=1.66 $X2=1.22 $Y2=1.95
cc_45 VPB N_A_82_48#_c_79_n 0.00316722f $X=-0.19 $Y=1.66 $X2=2.515 $Y2=2.775
cc_46 VPB N_A_82_48#_c_75_n 0.0170977f $X=-0.19 $Y=1.66 $X2=1.025 $Y2=1.532
cc_47 VPB N_B1_c_159_n 0.0380806f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=0.37
cc_48 VPB B1 0.00205167f $X=-0.19 $Y=1.66 $X2=0.485 $Y2=0.74
cc_49 VPB N_B2_c_192_n 0.0310204f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=0.37
cc_50 VPB N_B2_c_194_n 0.00404989f $X=-0.19 $Y=1.66 $X2=0.575 $Y2=2.4
cc_51 VPB N_A2_c_225_n 0.0329432f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=0.37
cc_52 VPB A2 0.0144733f $X=-0.19 $Y=1.66 $X2=0.485 $Y2=0.74
cc_53 VPB N_A1_c_257_n 0.033885f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=0.37
cc_54 VPB N_A1_c_259_n 0.00745299f $X=-0.19 $Y=1.66 $X2=0.575 $Y2=2.4
cc_55 VPB N_VPWR_c_282_n 0.0128289f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_283_n 0.0679826f $X=-0.19 $Y=1.66 $X2=0.575 $Y2=2.4
cc_57 VPB N_VPWR_c_284_n 0.0186948f $X=-0.19 $Y=1.66 $X2=0.915 $Y2=0.74
cc_58 VPB N_VPWR_c_285_n 0.0109364f $X=-0.19 $Y=1.66 $X2=1.025 $Y2=2.4
cc_59 VPB N_VPWR_c_286_n 0.011929f $X=-0.19 $Y=1.66 $X2=1.22 $Y2=1.3
cc_60 VPB N_VPWR_c_287_n 0.0504241f $X=-0.19 $Y=1.66 $X2=1.22 $Y2=1.95
cc_61 VPB N_VPWR_c_288_n 0.0488009f $X=-0.19 $Y=1.66 $X2=2.515 $Y2=2.775
cc_62 VPB N_VPWR_c_289_n 0.0125729f $X=-0.19 $Y=1.66 $X2=2.515 $Y2=2.035
cc_63 VPB N_VPWR_c_281_n 0.0935613f $X=-0.19 $Y=1.66 $X2=1.14 $Y2=1.532
cc_64 VPB N_X_c_327_n 0.00166049f $X=-0.19 $Y=1.66 $X2=0.915 $Y2=0.74
cc_65 VPB N_X_c_328_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_X_c_325_n 0.00117889f $X=-0.19 $Y=1.66 $X2=1.025 $Y2=2.4
cc_67 N_A_82_48#_c_77_n N_B1_c_159_n 0.00738061f $X=1.025 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_68 N_A_82_48#_c_69_n N_B1_c_159_n 0.00397881f $X=1.22 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_69 N_A_82_48#_c_83_p N_B1_c_159_n 0.0182682f $X=2.35 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_70 N_A_82_48#_c_79_n N_B1_c_159_n 0.00271705f $X=2.515 $Y=2.775 $X2=-0.19
+ $Y2=-0.245
cc_71 N_A_82_48#_c_71_n N_B1_c_159_n 7.6891e-19 $X=1.14 $Y=1.465 $X2=-0.19
+ $Y2=-0.245
cc_72 N_A_82_48#_c_74_n N_B1_c_159_n 0.0017174f $X=2.005 $Y=0.965 $X2=-0.19
+ $Y2=-0.245
cc_73 N_A_82_48#_c_75_n N_B1_c_159_n 0.0139637f $X=1.025 $Y=1.532 $X2=-0.19
+ $Y2=-0.245
cc_74 N_A_82_48#_c_71_n N_B1_M1002_g 6.90513e-19 $X=1.14 $Y=1.465 $X2=0 $Y2=0
cc_75 N_A_82_48#_c_72_n N_B1_M1002_g 0.00407257f $X=1.14 $Y=1.3 $X2=0 $Y2=0
cc_76 N_A_82_48#_c_74_n N_B1_M1002_g 0.0176532f $X=2.005 $Y=0.965 $X2=0 $Y2=0
cc_77 N_A_82_48#_c_75_n N_B1_M1002_g 0.00353902f $X=1.025 $Y=1.532 $X2=0 $Y2=0
cc_78 N_A_82_48#_c_83_p B1 0.0229545f $X=2.35 $Y=2.035 $X2=0 $Y2=0
cc_79 N_A_82_48#_c_71_n B1 0.0201599f $X=1.14 $Y=1.465 $X2=0 $Y2=0
cc_80 N_A_82_48#_c_74_n B1 0.0164979f $X=2.005 $Y=0.965 $X2=0 $Y2=0
cc_81 N_A_82_48#_c_75_n B1 8.54661e-19 $X=1.025 $Y=1.532 $X2=0 $Y2=0
cc_82 N_A_82_48#_c_83_p N_B2_c_192_n 0.0119563f $X=2.35 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_83 N_A_82_48#_c_97_p N_B2_c_192_n 0.00120057f $X=2.515 $Y=2.12 $X2=-0.19
+ $Y2=-0.245
cc_84 N_A_82_48#_c_79_n N_B2_c_192_n 0.0146831f $X=2.515 $Y=2.775 $X2=-0.19
+ $Y2=-0.245
cc_85 N_A_82_48#_c_73_n N_B2_c_192_n 0.00229717f $X=2.115 $Y=0.965 $X2=-0.19
+ $Y2=-0.245
cc_86 N_A_82_48#_c_73_n N_B2_M1011_g 0.00451145f $X=2.115 $Y=0.965 $X2=0 $Y2=0
cc_87 N_A_82_48#_c_83_p N_B2_c_194_n 0.0208355f $X=2.35 $Y=2.035 $X2=0 $Y2=0
cc_88 N_A_82_48#_c_97_p N_B2_c_194_n 0.0102936f $X=2.515 $Y=2.12 $X2=0 $Y2=0
cc_89 N_A_82_48#_c_73_n N_B2_c_194_n 0.0134587f $X=2.115 $Y=0.965 $X2=0 $Y2=0
cc_90 N_A_82_48#_c_79_n N_A2_c_225_n 0.00481807f $X=2.515 $Y=2.775 $X2=-0.19
+ $Y2=-0.245
cc_91 N_A_82_48#_c_69_n N_VPWR_M1003_d 0.00250637f $X=1.22 $Y=1.95 $X2=0 $Y2=0
cc_92 N_A_82_48#_c_83_p N_VPWR_M1003_d 0.0173798f $X=2.35 $Y=2.035 $X2=0 $Y2=0
cc_93 N_A_82_48#_c_107_p N_VPWR_M1003_d 0.00301935f $X=1.305 $Y=2.035 $X2=0
+ $Y2=0
cc_94 N_A_82_48#_c_76_n N_VPWR_c_283_n 0.0261486f $X=0.575 $Y=1.765 $X2=0 $Y2=0
cc_95 N_A_82_48#_c_75_n N_VPWR_c_283_n 0.00255704f $X=1.025 $Y=1.532 $X2=0 $Y2=0
cc_96 N_A_82_48#_c_76_n N_VPWR_c_284_n 0.00445602f $X=0.575 $Y=1.765 $X2=0 $Y2=0
cc_97 N_A_82_48#_c_77_n N_VPWR_c_284_n 0.00445602f $X=1.025 $Y=1.765 $X2=0 $Y2=0
cc_98 N_A_82_48#_c_77_n N_VPWR_c_285_n 0.00300147f $X=1.025 $Y=1.765 $X2=0 $Y2=0
cc_99 N_A_82_48#_c_83_p N_VPWR_c_285_n 0.0345371f $X=2.35 $Y=2.035 $X2=0 $Y2=0
cc_100 N_A_82_48#_c_107_p N_VPWR_c_285_n 0.0132989f $X=1.305 $Y=2.035 $X2=0
+ $Y2=0
cc_101 N_A_82_48#_c_79_n N_VPWR_c_285_n 0.0193064f $X=2.515 $Y=2.775 $X2=0 $Y2=0
cc_102 N_A_82_48#_c_75_n N_VPWR_c_285_n 4.80755e-19 $X=1.025 $Y=1.532 $X2=0
+ $Y2=0
cc_103 N_A_82_48#_c_79_n N_VPWR_c_288_n 0.0125658f $X=2.515 $Y=2.775 $X2=0 $Y2=0
cc_104 N_A_82_48#_c_76_n N_VPWR_c_281_n 0.00860622f $X=0.575 $Y=1.765 $X2=0
+ $Y2=0
cc_105 N_A_82_48#_c_77_n N_VPWR_c_281_n 0.00861719f $X=1.025 $Y=1.765 $X2=0
+ $Y2=0
cc_106 N_A_82_48#_c_79_n N_VPWR_c_281_n 0.011805f $X=2.515 $Y=2.775 $X2=0 $Y2=0
cc_107 N_A_82_48#_M1006_g N_X_c_324_n 0.00563952f $X=0.485 $Y=0.74 $X2=0 $Y2=0
cc_108 N_A_82_48#_M1008_g N_X_c_324_n 2.51515e-19 $X=0.915 $Y=0.74 $X2=0 $Y2=0
cc_109 N_A_82_48#_c_76_n N_X_c_327_n 0.00188635f $X=0.575 $Y=1.765 $X2=0 $Y2=0
cc_110 N_A_82_48#_c_77_n N_X_c_327_n 0.00261226f $X=1.025 $Y=1.765 $X2=0 $Y2=0
cc_111 N_A_82_48#_c_69_n N_X_c_327_n 0.00559275f $X=1.22 $Y=1.95 $X2=0 $Y2=0
cc_112 N_A_82_48#_c_75_n N_X_c_327_n 0.00697862f $X=1.025 $Y=1.532 $X2=0 $Y2=0
cc_113 N_A_82_48#_c_76_n N_X_c_328_n 0.0109216f $X=0.575 $Y=1.765 $X2=0 $Y2=0
cc_114 N_A_82_48#_c_77_n N_X_c_328_n 0.0164541f $X=1.025 $Y=1.765 $X2=0 $Y2=0
cc_115 N_A_82_48#_M1006_g N_X_c_325_n 0.00602646f $X=0.485 $Y=0.74 $X2=0 $Y2=0
cc_116 N_A_82_48#_c_76_n N_X_c_325_n 0.00251865f $X=0.575 $Y=1.765 $X2=0 $Y2=0
cc_117 N_A_82_48#_M1008_g N_X_c_325_n 0.0023958f $X=0.915 $Y=0.74 $X2=0 $Y2=0
cc_118 N_A_82_48#_c_77_n N_X_c_325_n 4.27304e-19 $X=1.025 $Y=1.765 $X2=0 $Y2=0
cc_119 N_A_82_48#_c_69_n N_X_c_325_n 0.00896393f $X=1.22 $Y=1.95 $X2=0 $Y2=0
cc_120 N_A_82_48#_c_71_n N_X_c_325_n 0.0239021f $X=1.14 $Y=1.465 $X2=0 $Y2=0
cc_121 N_A_82_48#_c_72_n N_X_c_325_n 0.00799225f $X=1.14 $Y=1.3 $X2=0 $Y2=0
cc_122 N_A_82_48#_c_75_n N_X_c_325_n 0.0303129f $X=1.025 $Y=1.532 $X2=0 $Y2=0
cc_123 N_A_82_48#_M1006_g X 0.00477711f $X=0.485 $Y=0.74 $X2=0 $Y2=0
cc_124 N_A_82_48#_M1008_g X 0.00776619f $X=0.915 $Y=0.74 $X2=0 $Y2=0
cc_125 N_A_82_48#_c_70_n X 0.0145044f $X=1.305 $Y=1.005 $X2=0 $Y2=0
cc_126 N_A_82_48#_c_83_p A_383_384# 0.0110864f $X=2.35 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_127 N_A_82_48#_c_70_n N_VGND_M1008_s 0.00509051f $X=1.305 $Y=1.005 $X2=0
+ $Y2=0
cc_128 N_A_82_48#_M1006_g N_VGND_c_360_n 0.00478246f $X=0.485 $Y=0.74 $X2=0
+ $Y2=0
cc_129 N_A_82_48#_M1006_g N_VGND_c_361_n 4.28647e-19 $X=0.485 $Y=0.74 $X2=0
+ $Y2=0
cc_130 N_A_82_48#_M1008_g N_VGND_c_361_n 0.00900614f $X=0.915 $Y=0.74 $X2=0
+ $Y2=0
cc_131 N_A_82_48#_c_70_n N_VGND_c_361_n 0.0112419f $X=1.305 $Y=1.005 $X2=0 $Y2=0
cc_132 N_A_82_48#_c_71_n N_VGND_c_361_n 0.00352695f $X=1.14 $Y=1.465 $X2=0 $Y2=0
cc_133 N_A_82_48#_c_75_n N_VGND_c_361_n 0.00118875f $X=1.025 $Y=1.532 $X2=0
+ $Y2=0
cc_134 N_A_82_48#_M1006_g N_VGND_c_363_n 0.00434272f $X=0.485 $Y=0.74 $X2=0
+ $Y2=0
cc_135 N_A_82_48#_M1008_g N_VGND_c_363_n 0.00383152f $X=0.915 $Y=0.74 $X2=0
+ $Y2=0
cc_136 N_A_82_48#_M1006_g N_VGND_c_366_n 0.00823683f $X=0.485 $Y=0.74 $X2=0
+ $Y2=0
cc_137 N_A_82_48#_M1008_g N_VGND_c_366_n 0.00685545f $X=0.915 $Y=0.74 $X2=0
+ $Y2=0
cc_138 N_A_82_48#_c_74_n N_A_307_74#_M1002_s 0.00296342f $X=2.005 $Y=0.965
+ $X2=-0.19 $Y2=-0.245
cc_139 N_A_82_48#_M1002_d N_A_307_74#_c_409_n 0.00262063f $X=1.96 $Y=0.37 $X2=0
+ $Y2=0
cc_140 N_A_82_48#_c_73_n N_A_307_74#_c_409_n 0.0104858f $X=2.115 $Y=0.965 $X2=0
+ $Y2=0
cc_141 N_A_82_48#_c_74_n N_A_307_74#_c_409_n 0.00476112f $X=2.005 $Y=0.965 $X2=0
+ $Y2=0
cc_142 N_A_82_48#_c_73_n N_A_307_74#_c_412_n 0.00799569f $X=2.115 $Y=0.965 $X2=0
+ $Y2=0
cc_143 N_A_82_48#_M1008_g N_A_307_74#_c_414_n 5.23807e-19 $X=0.915 $Y=0.74 $X2=0
+ $Y2=0
cc_144 N_A_82_48#_c_74_n N_A_307_74#_c_414_n 0.021503f $X=2.005 $Y=0.965 $X2=0
+ $Y2=0
cc_145 N_B1_c_159_n N_B2_c_192_n 0.0733289f $X=1.84 $Y=1.845 $X2=-0.19
+ $Y2=-0.245
cc_146 B1 N_B2_c_192_n 2.99285e-19 $X=1.595 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_147 N_B1_M1002_g N_B2_M1011_g 0.0358967f $X=1.885 $Y=0.74 $X2=0 $Y2=0
cc_148 N_B1_c_159_n N_B2_c_194_n 0.00247394f $X=1.84 $Y=1.845 $X2=0 $Y2=0
cc_149 B1 N_B2_c_194_n 0.0283934f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_150 N_B1_c_159_n N_VPWR_c_285_n 0.0173392f $X=1.84 $Y=1.845 $X2=0 $Y2=0
cc_151 N_B1_c_159_n N_VPWR_c_288_n 0.00455951f $X=1.84 $Y=1.845 $X2=0 $Y2=0
cc_152 N_B1_c_159_n N_VPWR_c_281_n 0.00447788f $X=1.84 $Y=1.845 $X2=0 $Y2=0
cc_153 N_B1_M1002_g N_VGND_c_361_n 0.00332629f $X=1.885 $Y=0.74 $X2=0 $Y2=0
cc_154 N_B1_M1002_g N_VGND_c_364_n 0.00292759f $X=1.885 $Y=0.74 $X2=0 $Y2=0
cc_155 N_B1_M1002_g N_VGND_c_366_n 0.00363526f $X=1.885 $Y=0.74 $X2=0 $Y2=0
cc_156 N_B1_M1002_g N_A_307_74#_c_409_n 0.0084546f $X=1.885 $Y=0.74 $X2=0 $Y2=0
cc_157 N_B1_M1002_g N_A_307_74#_c_414_n 0.00558709f $X=1.885 $Y=0.74 $X2=0 $Y2=0
cc_158 N_B2_c_192_n N_A2_c_225_n 0.0453799f $X=2.29 $Y=1.845 $X2=-0.19
+ $Y2=-0.245
cc_159 N_B2_c_194_n N_A2_c_225_n 4.91206e-19 $X=2.335 $Y=1.595 $X2=-0.19
+ $Y2=-0.245
cc_160 N_B2_M1011_g N_A2_M1010_g 0.0286716f $X=2.345 $Y=0.74 $X2=0 $Y2=0
cc_161 N_B2_c_192_n A2 4.34077e-19 $X=2.29 $Y=1.845 $X2=0 $Y2=0
cc_162 N_B2_c_194_n A2 0.0236983f $X=2.335 $Y=1.595 $X2=0 $Y2=0
cc_163 N_B2_c_192_n N_VPWR_c_285_n 0.00246838f $X=2.29 $Y=1.845 $X2=0 $Y2=0
cc_164 N_B2_c_192_n N_VPWR_c_288_n 0.00534256f $X=2.29 $Y=1.845 $X2=0 $Y2=0
cc_165 N_B2_c_192_n N_VPWR_c_281_n 0.00533081f $X=2.29 $Y=1.845 $X2=0 $Y2=0
cc_166 N_B2_M1011_g N_VGND_c_364_n 0.00291649f $X=2.345 $Y=0.74 $X2=0 $Y2=0
cc_167 N_B2_M1011_g N_VGND_c_366_n 0.00360203f $X=2.345 $Y=0.74 $X2=0 $Y2=0
cc_168 N_B2_M1011_g N_A_307_74#_c_409_n 0.014305f $X=2.345 $Y=0.74 $X2=0 $Y2=0
cc_169 N_B2_c_192_n N_A_307_74#_c_412_n 7.565e-19 $X=2.29 $Y=1.845 $X2=0 $Y2=0
cc_170 N_B2_M1011_g N_A_307_74#_c_412_n 9.8635e-19 $X=2.345 $Y=0.74 $X2=0 $Y2=0
cc_171 N_B2_c_194_n N_A_307_74#_c_412_n 0.00194208f $X=2.335 $Y=1.595 $X2=0
+ $Y2=0
cc_172 N_B2_M1011_g N_A_307_74#_c_414_n 6.68686e-19 $X=2.345 $Y=0.74 $X2=0 $Y2=0
cc_173 N_A2_c_225_n N_A1_c_257_n 0.0588053f $X=2.8 $Y=1.845 $X2=-0.19 $Y2=-0.245
cc_174 N_A2_M1010_g N_A1_c_257_n 0.00558036f $X=2.845 $Y=0.74 $X2=-0.19
+ $Y2=-0.245
cc_175 A2 N_A1_c_257_n 0.00287847f $X=3.035 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_176 N_A2_M1010_g N_A1_M1007_g 0.0278115f $X=2.845 $Y=0.74 $X2=0 $Y2=0
cc_177 N_A2_c_225_n N_A1_c_259_n 2.41037e-19 $X=2.8 $Y=1.845 $X2=0 $Y2=0
cc_178 N_A2_M1010_g N_A1_c_259_n 5.8609e-19 $X=2.845 $Y=0.74 $X2=0 $Y2=0
cc_179 A2 N_A1_c_259_n 0.0287241f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_180 N_A2_c_225_n N_VPWR_c_287_n 0.00501236f $X=2.8 $Y=1.845 $X2=0 $Y2=0
cc_181 N_A2_c_225_n N_VPWR_c_288_n 0.00548708f $X=2.8 $Y=1.845 $X2=0 $Y2=0
cc_182 N_A2_c_225_n N_VPWR_c_281_n 0.00533081f $X=2.8 $Y=1.845 $X2=0 $Y2=0
cc_183 N_A2_M1010_g N_VGND_c_362_n 0.00544936f $X=2.845 $Y=0.74 $X2=0 $Y2=0
cc_184 N_A2_M1010_g N_VGND_c_364_n 0.00433139f $X=2.845 $Y=0.74 $X2=0 $Y2=0
cc_185 N_A2_M1010_g N_VGND_c_366_n 0.00817815f $X=2.845 $Y=0.74 $X2=0 $Y2=0
cc_186 N_A2_M1010_g N_A_307_74#_c_410_n 0.00225753f $X=2.845 $Y=0.74 $X2=0 $Y2=0
cc_187 N_A2_M1010_g N_A_307_74#_c_430_n 0.00673645f $X=2.845 $Y=0.74 $X2=0 $Y2=0
cc_188 N_A2_c_225_n N_A_307_74#_c_411_n 0.00245655f $X=2.8 $Y=1.845 $X2=0 $Y2=0
cc_189 N_A2_M1010_g N_A_307_74#_c_411_n 0.0120938f $X=2.845 $Y=0.74 $X2=0 $Y2=0
cc_190 A2 N_A_307_74#_c_411_n 0.0220803f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_191 N_A2_c_225_n N_A_307_74#_c_412_n 0.00146551f $X=2.8 $Y=1.845 $X2=0 $Y2=0
cc_192 N_A2_M1010_g N_A_307_74#_c_412_n 0.00109647f $X=2.845 $Y=0.74 $X2=0 $Y2=0
cc_193 A2 N_A_307_74#_c_412_n 0.00459921f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_194 N_A1_c_257_n N_VPWR_c_287_n 0.0259463f $X=3.34 $Y=1.845 $X2=0 $Y2=0
cc_195 N_A1_c_259_n N_VPWR_c_287_n 0.0262231f $X=3.57 $Y=1.465 $X2=0 $Y2=0
cc_196 N_A1_c_257_n N_VPWR_c_288_n 0.00492531f $X=3.34 $Y=1.845 $X2=0 $Y2=0
cc_197 N_A1_c_257_n N_VPWR_c_281_n 0.00483326f $X=3.34 $Y=1.845 $X2=0 $Y2=0
cc_198 N_A1_M1007_g N_VGND_c_362_n 0.012583f $X=3.345 $Y=0.74 $X2=0 $Y2=0
cc_199 N_A1_M1007_g N_VGND_c_365_n 0.00383152f $X=3.345 $Y=0.74 $X2=0 $Y2=0
cc_200 N_A1_M1007_g N_VGND_c_366_n 0.00761198f $X=3.345 $Y=0.74 $X2=0 $Y2=0
cc_201 N_A1_M1007_g N_A_307_74#_c_430_n 7.30686e-19 $X=3.345 $Y=0.74 $X2=0 $Y2=0
cc_202 N_A1_c_257_n N_A_307_74#_c_411_n 0.00317143f $X=3.34 $Y=1.845 $X2=0 $Y2=0
cc_203 N_A1_M1007_g N_A_307_74#_c_411_n 0.0171242f $X=3.345 $Y=0.74 $X2=0 $Y2=0
cc_204 N_A1_c_259_n N_A_307_74#_c_411_n 0.0270164f $X=3.57 $Y=1.465 $X2=0 $Y2=0
cc_205 N_A1_M1007_g N_A_307_74#_c_413_n 0.00159319f $X=3.345 $Y=0.74 $X2=0 $Y2=0
cc_206 N_VPWR_c_283_n N_X_c_327_n 0.0450694f $X=0.3 $Y=1.985 $X2=0 $Y2=0
cc_207 N_VPWR_c_284_n N_X_c_328_n 0.014552f $X=1.135 $Y=3.33 $X2=0 $Y2=0
cc_208 N_VPWR_c_285_n N_X_c_328_n 0.0267672f $X=1.615 $Y=2.41 $X2=0 $Y2=0
cc_209 N_VPWR_c_281_n N_X_c_328_n 0.0119791f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_210 N_X_c_324_n N_VGND_c_360_n 0.0300732f $X=0.7 $Y=0.515 $X2=0 $Y2=0
cc_211 N_X_c_324_n N_VGND_c_361_n 0.0113761f $X=0.7 $Y=0.515 $X2=0 $Y2=0
cc_212 N_X_c_324_n N_VGND_c_363_n 0.0112174f $X=0.7 $Y=0.515 $X2=0 $Y2=0
cc_213 N_X_c_324_n N_VGND_c_366_n 0.00922837f $X=0.7 $Y=0.515 $X2=0 $Y2=0
cc_214 X N_VGND_c_366_n 0.0025861f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_215 N_VGND_c_364_n N_A_307_74#_c_409_n 0.0247246f $X=2.965 $Y=0 $X2=0 $Y2=0
cc_216 N_VGND_c_366_n N_A_307_74#_c_409_n 0.0209615f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_217 N_VGND_c_362_n N_A_307_74#_c_410_n 0.00795492f $X=3.13 $Y=0.625 $X2=0
+ $Y2=0
cc_218 N_VGND_c_364_n N_A_307_74#_c_410_n 0.0146502f $X=2.965 $Y=0 $X2=0 $Y2=0
cc_219 N_VGND_c_366_n N_A_307_74#_c_410_n 0.0120674f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_220 N_VGND_M1010_d N_A_307_74#_c_411_n 0.00250873f $X=2.92 $Y=0.37 $X2=0
+ $Y2=0
cc_221 N_VGND_c_362_n N_A_307_74#_c_411_n 0.0209867f $X=3.13 $Y=0.625 $X2=0
+ $Y2=0
cc_222 N_VGND_c_362_n N_A_307_74#_c_413_n 0.0164982f $X=3.13 $Y=0.625 $X2=0
+ $Y2=0
cc_223 N_VGND_c_365_n N_A_307_74#_c_413_n 0.011066f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_224 N_VGND_c_366_n N_A_307_74#_c_413_n 0.00915947f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_225 N_VGND_c_361_n N_A_307_74#_c_414_n 0.0208243f $X=1.13 $Y=0.535 $X2=0
+ $Y2=0
cc_226 N_VGND_c_364_n N_A_307_74#_c_414_n 0.0139208f $X=2.965 $Y=0 $X2=0 $Y2=0
cc_227 N_VGND_c_366_n N_A_307_74#_c_414_n 0.0117508f $X=3.6 $Y=0 $X2=0 $Y2=0
