* NGSPICE file created from sky130_fd_sc_ls__a21o_2.ext - technology: sky130A

.subckt sky130_fd_sc_ls__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
M1000 X a_84_244# VGND VNB nshort w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=8.954e+11p ps=6.86e+06u
M1001 a_401_392# A2 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=5.75e+11p pd=5.15e+06u as=9.16e+11p ps=8.18e+06u
M1002 a_84_244# B1 VGND VNB nshort w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1003 X a_84_244# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=0p ps=0u
M1004 VPWR a_84_244# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_401_392# B1 a_84_244# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.75e+11p ps=2.55e+06u
M1006 VGND a_84_244# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND A2 a_484_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.368e+11p ps=2.12e+06u
M1008 a_484_74# A1 a_84_244# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR A1 a_401_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

