* NGSPICE file created from sky130_fd_sc_ls__decaphetap_2.ext - technology: sky130A

.subckt sky130_fd_sc_ls__decaphetap_2 VGND VPB VPWR
R0 VGND VNB short w=0u l=2.03e+06u
M1000 VPWR VGND VPWR VPB pshort w=1.255e+06u l=170000u
+  ad=6.526e+11p pd=6.06e+06u as=0p ps=0u
.ends

