* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
M1000 a_504_392# A2 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=5.75e+11p pd=5.15e+06u as=9.916e+11p ps=8.36e+06u
M1001 X a_187_244# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=0p ps=0u
M1002 a_187_244# a_32_368# VGND VNB nshort w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=9.689e+11p ps=7.11e+06u
M1003 VPWR a_187_244# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 X a_187_244# VGND VNB nshort w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1005 VPWR B1_N a_32_368# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=2.31e+11p ps=2.23e+06u
M1006 VGND A2 a_587_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.368e+11p ps=2.12e+06u
M1007 a_504_392# a_32_368# a_187_244# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.75e+11p ps=2.55e+06u
M1008 VPWR A1 a_504_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND B1_N a_32_368# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=1.4575e+11p ps=1.63e+06u
M1010 a_587_74# A1 a_187_244# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND a_187_244# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
