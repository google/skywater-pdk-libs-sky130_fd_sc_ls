* File: sky130_fd_sc_ls__o211a_1.spice
* Created: Fri Aug 28 13:43:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__o211a_1.pex.spice"
.subckt sky130_fd_sc_ls__o211a_1  VNB VPB A1 A2 B1 C1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* C1	C1
* B1	B1
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1008 N_VGND_M1008_d N_A_83_264#_M1008_g N_X_M1008_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2627 AS=0.2109 PD=2.19 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1003 N_VGND_M1003_d N_A1_M1003_g N_A_257_136#_M1003_s VNB NSHORT L=0.15 W=0.64
+ AD=0.1632 AS=0.2112 PD=1.15 PS=1.94 NRD=10.308 NRS=4.212 M=1 R=4.26667
+ SA=75000.3 SB=75002.3 A=0.096 P=1.58 MULT=1
MM1006 N_A_257_136#_M1006_d N_A2_M1006_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.64
+ AD=0.2352 AS=0.1632 PD=1.375 PS=1.15 NRD=0 NRS=32.808 M=1 R=4.26667 SA=75000.9
+ SB=75001.6 A=0.096 P=1.58 MULT=1
MM1004 A_662_136# N_B1_M1004_g N_A_257_136#_M1006_d VNB NSHORT L=0.15 W=0.64
+ AD=0.104 AS=0.2352 PD=0.965 PS=1.375 NRD=20.148 NRS=0 M=1 R=4.26667 SA=75001.8
+ SB=75000.7 A=0.096 P=1.58 MULT=1
MM1002 N_A_83_264#_M1002_d N_C1_M1002_g A_662_136# VNB NSHORT L=0.15 W=0.64
+ AD=0.2112 AS=0.104 PD=1.94 PS=0.965 NRD=4.212 NRS=20.148 M=1 R=4.26667
+ SA=75002.3 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1005 N_VPWR_M1005_d N_A_83_264#_M1005_g N_X_M1005_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.68246 AS=0.3304 PD=2.51472 PS=2.83 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75003.2 A=0.168 P=2.54 MULT=1
MM1000 A_398_392# N_A1_M1000_g N_VPWR_M1005_d VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.60934 PD=1.27 PS=2.24528 NRD=15.7403 NRS=1.9503 M=1 R=6.66667 SA=75001.6
+ SB=75002.1 A=0.15 P=2.3 MULT=1
MM1007 N_A_83_264#_M1007_d N_A2_M1007_g A_398_392# VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.135 PD=1.3 PS=1.27 NRD=1.9503 NRS=15.7403 M=1 R=6.66667 SA=75002
+ SB=75001.7 A=0.15 P=2.3 MULT=1
MM1001 N_VPWR_M1001_d N_B1_M1001_g N_A_83_264#_M1007_d VPB PHIGHVT L=0.15 W=1
+ AD=0.44 AS=0.15 PD=1.88 PS=1.3 NRD=11.8003 NRS=1.9503 M=1 R=6.66667 SA=75002.5
+ SB=75001.2 A=0.15 P=2.3 MULT=1
MM1009 N_A_83_264#_M1009_d N_C1_M1009_g N_VPWR_M1001_d VPB PHIGHVT L=0.15 W=1
+ AD=0.295 AS=0.44 PD=2.59 PS=1.88 NRD=1.9503 NRS=11.8003 M=1 R=6.66667
+ SA=75003.5 SB=75000.2 A=0.15 P=2.3 MULT=1
DX10_noxref VNB VPB NWDIODE A=8.742 P=13.12
c_35 VNB 0 1.605e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_ls__o211a_1.pxi.spice"
*
.ends
*
*
