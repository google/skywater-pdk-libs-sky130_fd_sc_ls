* NGSPICE file created from sky130_fd_sc_ls__o2bb2ai_1.ext - technology: sky130A

.subckt sky130_fd_sc_ls__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
M1000 a_397_74# B1 VGND VNB nshort w=740000u l=150000u
+  ad=4.699e+11p pd=4.23e+06u as=3.896e+11p ps=3.89e+06u
M1001 a_131_383# A2_N a_114_74# VNB nshort w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=1.536e+11p ps=1.76e+06u
M1002 VPWR B1 a_490_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=1.36223e+12p pd=8.93e+06u as=3.696e+11p ps=2.9e+06u
M1003 Y a_131_383# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=0p ps=0u
M1004 VPWR A2_N a_131_383# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=2.52e+11p ps=2.28e+06u
M1005 VGND B2 a_397_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_490_368# B2 Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_397_74# a_131_383# Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1008 a_131_383# A1_N VPWR VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_114_74# A1_N VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

