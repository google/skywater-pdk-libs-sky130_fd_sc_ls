* NGSPICE file created from sky130_fd_sc_ls__a21oi_2.ext - technology: sky130A

.subckt sky130_fd_sc_ls__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
M1000 VPWR A2 a_131_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=7.392e+11p pd=5.8e+06u as=1.288e+12p ps=1.126e+07u
M1001 a_280_107# A2 VGND VNB nshort w=740000u l=150000u
+  ad=6.5505e+11p pd=6.27e+06u as=5.83425e+11p ps=4.82e+06u
M1002 a_131_368# A2 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VGND A2 a_280_107# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR A1 a_131_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y A1 a_280_107# VNB nshort w=740000u l=150000u
+  ad=4.033e+11p pd=4.05e+06u as=0p ps=0u
M1006 a_131_368# A1 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y B1 a_131_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=0p ps=0u
M1008 Y B1 VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_131_368# B1 Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_280_107# A1 Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

