* File: sky130_fd_sc_ls__a31o_4.pex.spice
* Created: Wed Sep  2 10:52:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__A31O_4%A_83_274# 1 2 3 4 13 15 16 18 19 21 22 24 25
+ 27 28 30 31 33 34 36 37 47 49 50 55 57 61 68 69 71 81
c139 71 0 2.72384e-19 $X=3.405 $Y=1.13
c140 61 0 9.60428e-20 $X=4.585 $Y=0.76
c141 57 0 1.54719e-19 $X=4.42 $Y=1.195
c142 34 0 1.24827e-19 $X=1.955 $Y=1.765
c143 13 0 4.66086e-20 $X=0.505 $Y=1.765
r144 80 81 8.86029 $w=4.08e-07 $l=7.5e-08 $layer=POLY_cond $X=1.88 $Y=1.492
+ $X2=1.955 $Y2=1.492
r145 77 78 9.45098 $w=4.08e-07 $l=8e-08 $layer=POLY_cond $X=1.425 $Y=1.492
+ $X2=1.505 $Y2=1.492
r146 74 75 4.72549 $w=4.08e-07 $l=4e-08 $layer=POLY_cond $X=0.955 $Y=1.492
+ $X2=0.995 $Y2=1.492
r147 73 74 51.3897 $w=4.08e-07 $l=4.35e-07 $layer=POLY_cond $X=0.52 $Y=1.492
+ $X2=0.955 $Y2=1.492
r148 72 73 1.77206 $w=4.08e-07 $l=1.5e-08 $layer=POLY_cond $X=0.505 $Y=1.492
+ $X2=0.52 $Y2=1.492
r149 68 69 7.89515 $w=4.48e-07 $l=1.15e-07 $layer=LI1_cond $X=3.35 $Y=2.085
+ $X2=3.35 $Y2=1.97
r150 65 81 25.3995 $w=4.08e-07 $l=2.15e-07 $layer=POLY_cond $X=2.17 $Y=1.492
+ $X2=1.955 $Y2=1.492
r151 64 65 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.17
+ $Y=1.385 $X2=2.17 $Y2=1.385
r152 59 61 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=4.585 $Y=1.11
+ $X2=4.585 $Y2=0.76
r153 58 71 4.30018 $w=1.7e-07 $l=3.76098e-07 $layer=LI1_cond $X=3.75 $Y=1.195
+ $X2=3.405 $Y2=1.13
r154 57 59 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.42 $Y=1.195
+ $X2=4.585 $Y2=1.11
r155 57 58 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.42 $Y=1.195
+ $X2=3.75 $Y2=1.195
r156 53 71 1.96316 $w=3.3e-07 $l=1.89737e-07 $layer=LI1_cond $X=3.585 $Y=1.11
+ $X2=3.405 $Y2=1.13
r157 53 55 20.7789 $w=3.28e-07 $l=5.95e-07 $layer=LI1_cond $X=3.585 $Y=1.11
+ $X2=3.585 $Y2=0.515
r158 51 71 1.96316 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=3.49 $Y=1.3
+ $X2=3.405 $Y2=1.13
r159 51 69 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.49 $Y=1.3
+ $X2=3.49 $Y2=1.97
r160 49 71 4.30018 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.405 $Y=1.215
+ $X2=3.405 $Y2=1.13
r161 49 50 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=3.405 $Y=1.215
+ $X2=2.74 $Y2=1.215
r162 45 50 7.35534 $w=3e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.615 $Y=1.13
+ $X2=2.74 $Y2=1.215
r163 45 64 18.0967 $w=3e-07 $l=5.39884e-07 $layer=LI1_cond $X=2.615 $Y=1.13
+ $X2=2.17 $Y2=1.34
r164 45 47 28.3501 $w=2.48e-07 $l=6.15e-07 $layer=LI1_cond $X=2.615 $Y=1.13
+ $X2=2.615 $Y2=0.515
r165 44 80 5.90686 $w=4.08e-07 $l=5e-08 $layer=POLY_cond $X=1.83 $Y=1.492
+ $X2=1.88 $Y2=1.492
r166 44 78 38.3946 $w=4.08e-07 $l=3.25e-07 $layer=POLY_cond $X=1.83 $Y=1.492
+ $X2=1.505 $Y2=1.492
r167 43 44 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.83
+ $Y=1.385 $X2=1.83 $Y2=1.385
r168 40 77 32.4877 $w=4.08e-07 $l=2.75e-07 $layer=POLY_cond $X=1.15 $Y=1.492
+ $X2=1.425 $Y2=1.492
r169 40 75 18.3113 $w=4.08e-07 $l=1.55e-07 $layer=POLY_cond $X=1.15 $Y=1.492
+ $X2=0.995 $Y2=1.492
r170 39 43 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.15 $Y=1.385
+ $X2=1.83 $Y2=1.385
r171 39 40 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.15
+ $Y=1.385 $X2=1.15 $Y2=1.385
r172 37 64 10.2918 $w=3.3e-07 $l=2.96648e-07 $layer=LI1_cond $X=1.895 $Y=1.385
+ $X2=2.17 $Y2=1.34
r173 37 43 2.26996 $w=3.28e-07 $l=6.5e-08 $layer=LI1_cond $X=1.895 $Y=1.385
+ $X2=1.83 $Y2=1.385
r174 34 81 26.3468 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=1.955 $Y=1.765
+ $X2=1.955 $Y2=1.492
r175 34 36 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.955 $Y=1.765
+ $X2=1.955 $Y2=2.4
r176 31 80 26.3468 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=1.88 $Y=1.22
+ $X2=1.88 $Y2=1.492
r177 31 33 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.88 $Y=1.22
+ $X2=1.88 $Y2=0.74
r178 28 78 26.3468 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=1.505 $Y=1.765
+ $X2=1.505 $Y2=1.492
r179 28 30 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.505 $Y=1.765
+ $X2=1.505 $Y2=2.4
r180 25 77 26.3468 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=1.425 $Y=1.22
+ $X2=1.425 $Y2=1.492
r181 25 27 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.425 $Y=1.22
+ $X2=1.425 $Y2=0.74
r182 22 75 26.3468 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=0.995 $Y=1.22
+ $X2=0.995 $Y2=1.492
r183 22 24 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.995 $Y=1.22
+ $X2=0.995 $Y2=0.74
r184 19 74 26.3468 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=0.955 $Y=1.765
+ $X2=0.955 $Y2=1.492
r185 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.955 $Y=1.765
+ $X2=0.955 $Y2=2.4
r186 16 73 26.3468 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=0.52 $Y=1.22
+ $X2=0.52 $Y2=1.492
r187 16 18 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.52 $Y=1.22
+ $X2=0.52 $Y2=0.74
r188 13 72 26.3468 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=1.492
r189 13 15 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.4
r190 4 68 300 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=2 $X=3.09
+ $Y=1.96 $X2=3.3 $Y2=2.085
r191 3 61 182 $w=1.7e-07 $l=4.83735e-07 $layer=licon1_NDIFF $count=1 $X=4.375
+ $Y=0.37 $X2=4.585 $Y2=0.76
r192 2 55 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.445
+ $Y=0.37 $X2=3.585 $Y2=0.515
r193 1 47 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=2.51
+ $Y=0.37 $X2=2.655 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__A31O_4%B1 3 5 7 10 12 14 15 22
c62 22 0 7.20501e-20 $X=3.37 $Y=1.677
c63 15 0 1.24827e-19 $X=3.12 $Y=1.665
c64 3 0 9.37482e-20 $X=2.87 $Y=0.69
r65 22 23 24.247 $w=3.28e-07 $l=1.65e-07 $layer=POLY_cond $X=3.37 $Y=1.677
+ $X2=3.535 $Y2=1.677
r66 20 22 44.0854 $w=3.28e-07 $l=3e-07 $layer=POLY_cond $X=3.07 $Y=1.677
+ $X2=3.37 $Y2=1.677
r67 18 20 8.08232 $w=3.28e-07 $l=5.5e-08 $layer=POLY_cond $X=3.015 $Y=1.677
+ $X2=3.07 $Y2=1.677
r68 17 18 21.3079 $w=3.28e-07 $l=1.45e-07 $layer=POLY_cond $X=2.87 $Y=1.677
+ $X2=3.015 $Y2=1.677
r69 15 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.07
+ $Y=1.635 $X2=3.07 $Y2=1.635
r70 12 23 21.0783 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.535 $Y=1.885
+ $X2=3.535 $Y2=1.677
r71 12 14 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.535 $Y=1.885
+ $X2=3.535 $Y2=2.46
r72 8 22 21.0783 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.37 $Y=1.47
+ $X2=3.37 $Y2=1.677
r73 8 10 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=3.37 $Y=1.47 $X2=3.37
+ $Y2=0.69
r74 5 18 21.0783 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.015 $Y=1.885
+ $X2=3.015 $Y2=1.677
r75 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.015 $Y=1.885
+ $X2=3.015 $Y2=2.46
r76 1 17 21.0783 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.87 $Y=1.47
+ $X2=2.87 $Y2=1.677
r77 1 3 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=2.87 $Y=1.47 $X2=2.87
+ $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_LS__A31O_4%A1 1 3 4 5 7 8 10 11 13 14 16 17 18 19 25
r70 25 27 17.0787 $w=3.81e-07 $l=1.35e-07 $layer=POLY_cond $X=4.55 $Y=1.667
+ $X2=4.685 $Y2=1.667
r71 23 25 43.0131 $w=3.81e-07 $l=3.4e-07 $layer=POLY_cond $X=4.21 $Y=1.667
+ $X2=4.55 $Y2=1.667
r72 22 23 9.48819 $w=3.81e-07 $l=7.5e-08 $layer=POLY_cond $X=4.135 $Y=1.667
+ $X2=4.21 $Y2=1.667
r73 19 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.55
+ $Y=1.615 $X2=4.55 $Y2=1.615
r74 18 19 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=4.08 $Y=1.615
+ $X2=4.55 $Y2=1.615
r75 14 27 24.6764 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=4.685 $Y=1.885
+ $X2=4.685 $Y2=1.667
r76 14 16 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=4.685 $Y=1.885
+ $X2=4.685 $Y2=2.46
r77 11 17 13.5877 $w=2.4e-07 $l=1.21861e-07 $layer=POLY_cond $X=4.3 $Y=1.085
+ $X2=4.21 $Y2=1.16
r78 11 13 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=4.3 $Y=1.085
+ $X2=4.3 $Y2=0.69
r79 8 22 24.6764 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=4.135 $Y=1.885
+ $X2=4.135 $Y2=1.667
r80 8 10 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=4.135 $Y=1.885
+ $X2=4.135 $Y2=2.46
r81 7 23 6.23733 $w=3.3e-07 $l=2.17e-07 $layer=POLY_cond $X=4.21 $Y=1.45
+ $X2=4.21 $Y2=1.667
r82 6 17 13.5877 $w=2.4e-07 $l=7.5e-08 $layer=POLY_cond $X=4.21 $Y=1.235
+ $X2=4.21 $Y2=1.16
r83 6 7 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=4.21 $Y=1.235
+ $X2=4.21 $Y2=1.45
r84 4 17 12.1617 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.045 $Y=1.16
+ $X2=4.21 $Y2=1.16
r85 4 5 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=4.045 $Y=1.16
+ $X2=3.875 $Y2=1.16
r86 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.8 $Y=1.085
+ $X2=3.875 $Y2=1.16
r87 1 3 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.8 $Y=1.085 $X2=3.8
+ $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_LS__A31O_4%A2 1 3 5 6 8 10 11 13 16 18 21 23 24 29 30
c71 21 0 9.60428e-20 $X=5.36 $Y=1.16
c72 18 0 1.64432e-19 $X=5.045 $Y=1.6
c73 16 0 1.03588e-19 $X=5.79 $Y=0.69
r74 29 31 10.791 $w=4.02e-07 $l=9e-08 $layer=POLY_cond $X=5.7 $Y=1.667 $X2=5.79
+ $Y2=1.667
r75 29 30 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.7
+ $Y=1.615 $X2=5.7 $Y2=1.615
r76 27 29 0.599503 $w=4.02e-07 $l=5e-09 $layer=POLY_cond $X=5.695 $Y=1.667
+ $X2=5.7 $Y2=1.667
r77 24 30 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=5.52 $Y=1.615
+ $X2=5.7 $Y2=1.615
r78 23 24 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=5.04 $Y=1.615
+ $X2=5.52 $Y2=1.615
r79 19 21 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=5.15 $Y=1.16
+ $X2=5.36 $Y2=1.16
r80 14 31 25.9839 $w=1.5e-07 $l=2.17e-07 $layer=POLY_cond $X=5.79 $Y=1.45
+ $X2=5.79 $Y2=1.667
r81 14 16 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=5.79 $Y=1.45
+ $X2=5.79 $Y2=0.69
r82 11 27 25.9839 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=5.695 $Y=1.885
+ $X2=5.695 $Y2=1.667
r83 11 13 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.695 $Y=1.885
+ $X2=5.695 $Y2=2.46
r84 8 21 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.36 $Y=1.085
+ $X2=5.36 $Y2=1.16
r85 8 10 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=5.36 $Y=1.085
+ $X2=5.36 $Y2=0.69
r86 7 18 5.03009 $w=3.3e-07 $l=1.8735e-07 $layer=POLY_cond $X=5.225 $Y=1.615
+ $X2=5.045 $Y2=1.6
r87 6 27 12.4798 $w=4.02e-07 $l=1.13049e-07 $layer=POLY_cond $X=5.605 $Y=1.615
+ $X2=5.695 $Y2=1.667
r88 6 7 66.4473 $w=3.3e-07 $l=3.8e-07 $layer=POLY_cond $X=5.605 $Y=1.615
+ $X2=5.225 $Y2=1.615
r89 5 18 37.0704 $w=1.5e-07 $l=1.95576e-07 $layer=POLY_cond $X=5.15 $Y=1.45
+ $X2=5.045 $Y2=1.6
r90 4 19 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.15 $Y=1.235
+ $X2=5.15 $Y2=1.16
r91 4 5 110.245 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=5.15 $Y=1.235
+ $X2=5.15 $Y2=1.45
r92 1 18 37.0704 $w=1.5e-07 $l=3.26917e-07 $layer=POLY_cond $X=5.135 $Y=1.885
+ $X2=5.045 $Y2=1.6
r93 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.135 $Y=1.885
+ $X2=5.135 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_LS__A31O_4%A3 1 3 6 10 12 14 15 16 24
r43 24 25 5.63377 $w=3.85e-07 $l=4.5e-08 $layer=POLY_cond $X=6.65 $Y=1.667
+ $X2=6.695 $Y2=1.667
r44 22 24 3.75584 $w=3.85e-07 $l=3e-08 $layer=POLY_cond $X=6.62 $Y=1.667
+ $X2=6.65 $Y2=1.667
r45 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.62
+ $Y=1.615 $X2=6.62 $Y2=1.615
r46 20 22 50.0779 $w=3.85e-07 $l=4e-07 $layer=POLY_cond $X=6.22 $Y=1.667
+ $X2=6.62 $Y2=1.667
r47 19 20 3.12987 $w=3.85e-07 $l=2.5e-08 $layer=POLY_cond $X=6.195 $Y=1.667
+ $X2=6.22 $Y2=1.667
r48 16 23 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=6.96 $Y=1.615
+ $X2=6.62 $Y2=1.615
r49 15 23 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=6.48 $Y=1.615
+ $X2=6.62 $Y2=1.615
r50 12 25 24.9301 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=6.695 $Y=1.885
+ $X2=6.695 $Y2=1.667
r51 12 14 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.695 $Y=1.885
+ $X2=6.695 $Y2=2.46
r52 8 24 24.9301 $w=1.5e-07 $l=2.17e-07 $layer=POLY_cond $X=6.65 $Y=1.45
+ $X2=6.65 $Y2=1.667
r53 8 10 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=6.65 $Y=1.45 $X2=6.65
+ $Y2=0.69
r54 4 20 24.9301 $w=1.5e-07 $l=2.17e-07 $layer=POLY_cond $X=6.22 $Y=1.45
+ $X2=6.22 $Y2=1.667
r55 4 6 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=6.22 $Y=1.45 $X2=6.22
+ $Y2=0.69
r56 1 19 24.9301 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=6.195 $Y=1.885
+ $X2=6.195 $Y2=1.667
r57 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.195 $Y=1.885
+ $X2=6.195 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_LS__A31O_4%VPWR 1 2 3 4 5 6 19 21 27 33 39 43 47 50 51
+ 53 54 55 57 62 77 83 84 90 93 96
r96 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r97 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r98 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r99 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r100 84 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6.48 $Y2=3.33
r101 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r102 81 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.585 $Y=3.33
+ $X2=6.42 $Y2=3.33
r103 81 83 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=6.585 $Y=3.33
+ $X2=6.96 $Y2=3.33
r104 80 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r105 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r106 77 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.255 $Y=3.33
+ $X2=6.42 $Y2=3.33
r107 77 79 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=6.255 $Y=3.33
+ $X2=6 $Y2=3.33
r108 76 80 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33 $X2=6
+ $Y2=3.33
r109 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r110 73 76 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r111 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r112 70 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r113 69 72 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.64 $Y=3.33
+ $X2=4.08 $Y2=3.33
r114 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r115 67 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.395 $Y=3.33
+ $X2=2.23 $Y2=3.33
r116 67 69 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=2.395 $Y=3.33
+ $X2=2.64 $Y2=3.33
r117 66 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r118 66 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r119 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r120 63 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.395 $Y=3.33
+ $X2=1.23 $Y2=3.33
r121 63 65 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.395 $Y=3.33
+ $X2=1.68 $Y2=3.33
r122 62 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.065 $Y=3.33
+ $X2=2.23 $Y2=3.33
r123 62 65 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=2.065 $Y=3.33
+ $X2=1.68 $Y2=3.33
r124 61 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r125 61 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r126 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r127 58 87 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.182 $Y2=3.33
r128 58 60 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.72 $Y2=3.33
r129 57 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.065 $Y=3.33
+ $X2=1.23 $Y2=3.33
r130 57 60 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.065 $Y=3.33
+ $X2=0.72 $Y2=3.33
r131 55 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r132 55 70 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=2.64 $Y2=3.33
r133 53 75 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=5.245 $Y=3.33
+ $X2=5.04 $Y2=3.33
r134 53 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.245 $Y=3.33
+ $X2=5.41 $Y2=3.33
r135 52 79 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=5.575 $Y=3.33
+ $X2=6 $Y2=3.33
r136 52 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.575 $Y=3.33
+ $X2=5.41 $Y2=3.33
r137 50 72 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=4.245 $Y=3.33
+ $X2=4.08 $Y2=3.33
r138 50 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.245 $Y=3.33
+ $X2=4.41 $Y2=3.33
r139 49 75 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=4.575 $Y=3.33
+ $X2=5.04 $Y2=3.33
r140 49 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.575 $Y=3.33
+ $X2=4.41 $Y2=3.33
r141 45 96 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.42 $Y=3.245
+ $X2=6.42 $Y2=3.33
r142 45 47 28.6365 $w=3.28e-07 $l=8.2e-07 $layer=LI1_cond $X=6.42 $Y=3.245
+ $X2=6.42 $Y2=2.425
r143 41 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.41 $Y=3.245
+ $X2=5.41 $Y2=3.33
r144 41 43 28.6365 $w=3.28e-07 $l=8.2e-07 $layer=LI1_cond $X=5.41 $Y=3.245
+ $X2=5.41 $Y2=2.425
r145 37 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.41 $Y=3.245
+ $X2=4.41 $Y2=3.33
r146 37 39 28.6365 $w=3.28e-07 $l=8.2e-07 $layer=LI1_cond $X=4.41 $Y=3.245
+ $X2=4.41 $Y2=2.425
r147 33 36 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=2.23 $Y=1.985
+ $X2=2.23 $Y2=2.815
r148 31 93 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.23 $Y=3.245
+ $X2=2.23 $Y2=3.33
r149 31 36 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.23 $Y=3.245
+ $X2=2.23 $Y2=2.815
r150 27 30 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.23 $Y=2.145
+ $X2=1.23 $Y2=2.825
r151 25 90 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.23 $Y=3.245
+ $X2=1.23 $Y2=3.33
r152 25 30 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=1.23 $Y=3.245
+ $X2=1.23 $Y2=2.825
r153 21 24 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=0.24 $Y=1.985
+ $X2=0.24 $Y2=2.815
r154 19 87 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.182 $Y2=3.33
r155 19 24 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.24 $Y2=2.815
r156 6 47 300 $w=1.7e-07 $l=5.34766e-07 $layer=licon1_PDIFF $count=2 $X=6.27
+ $Y=1.96 $X2=6.42 $Y2=2.425
r157 5 43 300 $w=1.7e-07 $l=5.5608e-07 $layer=licon1_PDIFF $count=2 $X=5.21
+ $Y=1.96 $X2=5.41 $Y2=2.425
r158 4 39 300 $w=1.7e-07 $l=5.5608e-07 $layer=licon1_PDIFF $count=2 $X=4.21
+ $Y=1.96 $X2=4.41 $Y2=2.425
r159 3 36 400 $w=1.7e-07 $l=1.07034e-06 $layer=licon1_PDIFF $count=1 $X=2.03
+ $Y=1.84 $X2=2.23 $Y2=2.815
r160 3 33 400 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=1 $X=2.03
+ $Y=1.84 $X2=2.23 $Y2=1.985
r161 2 30 400 $w=1.7e-07 $l=1.08038e-06 $layer=licon1_PDIFF $count=1 $X=1.03
+ $Y=1.84 $X2=1.23 $Y2=2.825
r162 2 27 400 $w=1.7e-07 $l=3.9246e-07 $layer=licon1_PDIFF $count=1 $X=1.03
+ $Y=1.84 $X2=1.23 $Y2=2.145
r163 1 24 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r164 1 21 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_LS__A31O_4%X 1 2 3 4 15 19 21 25 29 35 36 37 38 54
c57 21 0 1.18659e-19 $X=1.565 $Y=1.805
r58 43 56 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=1.89
+ $X2=0.73 $Y2=1.805
r59 37 38 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.73 $Y=2.405
+ $X2=0.73 $Y2=2.775
r60 36 37 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=0.73 $Y=1.985
+ $X2=0.73 $Y2=2.405
r61 36 43 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=0.73 $Y=1.985
+ $X2=0.73 $Y2=1.89
r62 35 56 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=0.73 $Y=1.665
+ $X2=0.73 $Y2=1.805
r63 35 54 4.72076 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=0.73 $Y=1.665
+ $X2=0.73 $Y2=1.55
r64 29 31 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=1.73 $Y=1.985
+ $X2=1.73 $Y2=2.815
r65 27 29 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=1.73 $Y=1.89
+ $X2=1.73 $Y2=1.985
r66 23 25 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.64 $Y=0.83
+ $X2=1.64 $Y2=0.495
r67 22 56 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=1.805
+ $X2=0.73 $Y2=1.805
r68 21 27 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.565 $Y=1.805
+ $X2=1.73 $Y2=1.89
r69 21 22 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.565 $Y=1.805
+ $X2=0.895 $Y2=1.805
r70 20 34 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.865 $Y=0.915
+ $X2=0.74 $Y2=0.915
r71 19 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.555 $Y=0.915
+ $X2=1.64 $Y2=0.83
r72 19 20 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.555 $Y=0.915
+ $X2=0.865 $Y2=0.915
r73 17 34 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.74 $Y=1 $X2=0.74
+ $Y2=0.915
r74 17 54 25.3537 $w=2.48e-07 $l=5.5e-07 $layer=LI1_cond $X=0.74 $Y=1 $X2=0.74
+ $Y2=1.55
r75 13 34 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.74 $Y=0.83 $X2=0.74
+ $Y2=0.915
r76 13 15 14.5208 $w=2.48e-07 $l=3.15e-07 $layer=LI1_cond $X=0.74 $Y=0.83
+ $X2=0.74 $Y2=0.515
r77 4 31 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.58
+ $Y=1.84 $X2=1.73 $Y2=2.815
r78 4 29 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.58
+ $Y=1.84 $X2=1.73 $Y2=1.985
r79 3 38 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.84 $X2=0.73 $Y2=2.815
r80 3 36 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.84 $X2=0.73 $Y2=1.985
r81 2 25 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.5
+ $Y=0.37 $X2=1.64 $Y2=0.495
r82 1 34 182 $w=1.7e-07 $l=6.81249e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.37 $X2=0.78 $Y2=0.965
r83 1 15 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.37 $X2=0.78 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__A31O_4%A_529_392# 1 2 3 4 5 16 18 20 22 23 24 28 30
+ 34 36 38 40 49 51
c97 49 0 1.54719e-19 $X=4.91 $Y=2.115
c98 36 0 1.47061e-19 $X=6.755 $Y=2.035
c99 22 0 1.78636e-19 $X=3.91 $Y=2.12
r100 38 53 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.92 $Y=2.12 $X2=6.92
+ $Y2=2.035
r101 38 40 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=6.92 $Y=2.12
+ $X2=6.92 $Y2=2.815
r102 37 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.085 $Y=2.035
+ $X2=5.92 $Y2=2.035
r103 36 53 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.755 $Y=2.035
+ $X2=6.92 $Y2=2.035
r104 36 37 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.755 $Y=2.035
+ $X2=6.085 $Y2=2.035
r105 32 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.92 $Y=2.12
+ $X2=5.92 $Y2=2.035
r106 32 34 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=5.92 $Y=2.12
+ $X2=5.92 $Y2=2.815
r107 31 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.075 $Y=2.035
+ $X2=4.91 $Y2=2.035
r108 30 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.755 $Y=2.035
+ $X2=5.92 $Y2=2.035
r109 30 31 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=5.755 $Y=2.035
+ $X2=5.075 $Y2=2.035
r110 26 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.91 $Y=2.12
+ $X2=4.91 $Y2=2.035
r111 26 28 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=4.91 $Y=2.12
+ $X2=4.91 $Y2=2.815
r112 25 45 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.075 $Y=2.035
+ $X2=3.91 $Y2=2.035
r113 24 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.745 $Y=2.035
+ $X2=4.91 $Y2=2.035
r114 24 25 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.745 $Y=2.035
+ $X2=4.075 $Y2=2.035
r115 23 47 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.91 $Y=2.81 $X2=3.91
+ $Y2=2.895
r116 22 45 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.91 $Y=2.12 $X2=3.91
+ $Y2=2.035
r117 22 23 24.0965 $w=3.28e-07 $l=6.9e-07 $layer=LI1_cond $X=3.91 $Y=2.12
+ $X2=3.91 $Y2=2.81
r118 21 43 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.955 $Y=2.895
+ $X2=2.79 $Y2=2.895
r119 20 47 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.745 $Y=2.895
+ $X2=3.91 $Y2=2.895
r120 20 21 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=3.745 $Y=2.895
+ $X2=2.955 $Y2=2.895
r121 16 43 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.79 $Y=2.81 $X2=2.79
+ $Y2=2.895
r122 16 18 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.79 $Y=2.81
+ $X2=2.79 $Y2=2.135
r123 5 53 400 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=1 $X=6.77
+ $Y=1.96 $X2=6.92 $Y2=2.115
r124 5 40 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=6.77
+ $Y=1.96 $X2=6.92 $Y2=2.815
r125 4 51 400 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=1 $X=5.77
+ $Y=1.96 $X2=5.92 $Y2=2.115
r126 4 34 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=5.77
+ $Y=1.96 $X2=5.92 $Y2=2.815
r127 3 49 400 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=1 $X=4.76
+ $Y=1.96 $X2=4.91 $Y2=2.115
r128 3 28 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=4.76
+ $Y=1.96 $X2=4.91 $Y2=2.815
r129 2 47 400 $w=1.7e-07 $l=9.93743e-07 $layer=licon1_PDIFF $count=1 $X=3.61
+ $Y=1.96 $X2=3.91 $Y2=2.815
r130 2 45 400 $w=1.7e-07 $l=3.69459e-07 $layer=licon1_PDIFF $count=1 $X=3.61
+ $Y=1.96 $X2=3.91 $Y2=2.115
r131 1 43 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=2.645
+ $Y=1.96 $X2=2.79 $Y2=2.815
r132 1 18 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=2.645
+ $Y=1.96 $X2=2.79 $Y2=2.135
.ends

.subckt PM_SKY130_FD_SC_LS__A31O_4%VGND 1 2 3 4 5 16 18 22 26 30 34 36 38 43 48
+ 53 63 64 70 73 76 79
r90 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r91 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r92 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r93 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r94 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r95 64 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=6.48
+ $Y2=0
r96 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r97 61 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.6 $Y=0 $X2=6.435
+ $Y2=0
r98 61 63 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=6.6 $Y=0 $X2=6.96
+ $Y2=0
r99 60 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r100 59 60 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6 $Y=0 $X2=6 $Y2=0
r101 56 59 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=3.6 $Y=0 $X2=6
+ $Y2=0
r102 54 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.25 $Y=0 $X2=3.085
+ $Y2=0
r103 54 56 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=3.25 $Y=0 $X2=3.6
+ $Y2=0
r104 53 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.27 $Y=0 $X2=6.435
+ $Y2=0
r105 53 59 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=6.27 $Y=0 $X2=6
+ $Y2=0
r106 52 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r107 52 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r108 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r109 49 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.26 $Y=0 $X2=2.095
+ $Y2=0
r110 49 51 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=2.26 $Y=0 $X2=2.64
+ $Y2=0
r111 48 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.92 $Y=0 $X2=3.085
+ $Y2=0
r112 48 51 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=2.92 $Y=0 $X2=2.64
+ $Y2=0
r113 47 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r114 47 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r115 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r116 44 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.375 $Y=0 $X2=1.21
+ $Y2=0
r117 44 46 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.375 $Y=0
+ $X2=1.68 $Y2=0
r118 43 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.93 $Y=0 $X2=2.095
+ $Y2=0
r119 43 46 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.93 $Y=0 $X2=1.68
+ $Y2=0
r120 42 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r121 42 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r122 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r123 39 67 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=0
+ $X2=0.222 $Y2=0
r124 39 41 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=0
+ $X2=0.72 $Y2=0
r125 38 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.045 $Y=0 $X2=1.21
+ $Y2=0
r126 38 41 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.045 $Y=0
+ $X2=0.72 $Y2=0
r127 36 60 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=3.6 $Y=0 $X2=6
+ $Y2=0
r128 36 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r129 36 56 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r130 32 79 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.435 $Y=0.085
+ $X2=6.435 $Y2=0
r131 32 34 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=6.435 $Y=0.085
+ $X2=6.435 $Y2=0.495
r132 28 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.085 $Y=0.085
+ $X2=3.085 $Y2=0
r133 28 30 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=3.085 $Y=0.085
+ $X2=3.085 $Y2=0.495
r134 24 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.095 $Y=0.085
+ $X2=2.095 $Y2=0
r135 24 26 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.095 $Y=0.085
+ $X2=2.095 $Y2=0.515
r136 20 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.21 $Y=0.085
+ $X2=1.21 $Y2=0
r137 20 22 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=1.21 $Y=0.085
+ $X2=1.21 $Y2=0.565
r138 16 67 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.222 $Y2=0
r139 16 18 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.28 $Y2=0.515
r140 5 34 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=6.295
+ $Y=0.37 $X2=6.435 $Y2=0.495
r141 4 30 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=2.945
+ $Y=0.37 $X2=3.085 $Y2=0.495
r142 3 26 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.955
+ $Y=0.37 $X2=2.095 $Y2=0.515
r143 2 22 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=1.07
+ $Y=0.37 $X2=1.21 $Y2=0.565
r144 1 18 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__A31O_4%A_775_74# 1 2 9 11 12 15
r27 13 15 2.44458 $w=3.28e-07 $l=7e-08 $layer=LI1_cond $X=5.575 $Y=0.425
+ $X2=5.575 $Y2=0.495
r28 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.41 $Y=0.34
+ $X2=5.575 $Y2=0.425
r29 11 12 75.6791 $w=1.68e-07 $l=1.16e-06 $layer=LI1_cond $X=5.41 $Y=0.34
+ $X2=4.25 $Y2=0.34
r30 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.085 $Y=0.425
+ $X2=4.25 $Y2=0.34
r31 7 9 2.44458 $w=3.28e-07 $l=7e-08 $layer=LI1_cond $X=4.085 $Y=0.425 $X2=4.085
+ $Y2=0.495
r32 2 15 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=5.435
+ $Y=0.37 $X2=5.575 $Y2=0.495
r33 1 9 91 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=2 $X=3.875
+ $Y=0.37 $X2=4.085 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LS__A31O_4%A_1000_74# 1 2 3 12 14 15 18 20 24 26
c40 26 0 1.47061e-19 $X=6.005 $Y=1.195
c41 15 0 1.64432e-19 $X=5.23 $Y=1.195
c42 12 0 1.03588e-19 $X=5.145 $Y=0.76
r43 22 24 27.4281 $w=2.48e-07 $l=5.95e-07 $layer=LI1_cond $X=6.905 $Y=1.11
+ $X2=6.905 $Y2=0.515
r44 21 26 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.09 $Y=1.195
+ $X2=6.005 $Y2=1.195
r45 20 22 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.78 $Y=1.195
+ $X2=6.905 $Y2=1.11
r46 20 21 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=6.78 $Y=1.195
+ $X2=6.09 $Y2=1.195
r47 16 26 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.005 $Y=1.11
+ $X2=6.005 $Y2=1.195
r48 16 18 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=6.005 $Y=1.11
+ $X2=6.005 $Y2=0.515
r49 14 26 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.92 $Y=1.195
+ $X2=6.005 $Y2=1.195
r50 14 15 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.92 $Y=1.195
+ $X2=5.23 $Y2=1.195
r51 10 15 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.105 $Y=1.11
+ $X2=5.23 $Y2=1.195
r52 10 12 16.1342 $w=2.48e-07 $l=3.5e-07 $layer=LI1_cond $X=5.105 $Y=1.11
+ $X2=5.105 $Y2=0.76
r53 3 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.725
+ $Y=0.37 $X2=6.865 $Y2=0.515
r54 2 18 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.865
+ $Y=0.37 $X2=6.005 $Y2=0.515
r55 1 12 182 $w=1.7e-07 $l=4.56782e-07 $layer=licon1_NDIFF $count=1 $X=5 $Y=0.37
+ $X2=5.145 $Y2=0.76
.ends

