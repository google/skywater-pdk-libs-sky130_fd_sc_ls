* File: sky130_fd_sc_ls__dfrbp_2.pxi.spice
* Created: Fri Aug 28 13:13:58 2020
* 
x_PM_SKY130_FD_SC_LS__DFRBP_2%D N_D_c_269_n N_D_c_276_n N_D_M1027_g N_D_M1008_g
+ N_D_c_270_n N_D_c_271_n N_D_c_272_n D D N_D_c_274_n
+ PM_SKY130_FD_SC_LS__DFRBP_2%D
x_PM_SKY130_FD_SC_LS__DFRBP_2%A_298_294# N_A_298_294#_M1004_d
+ N_A_298_294#_M1032_s N_A_298_294#_M1001_d N_A_298_294#_c_312_n
+ N_A_298_294#_M1031_g N_A_298_294#_M1034_g N_A_298_294#_c_305_n
+ N_A_298_294#_c_306_n N_A_298_294#_c_307_n N_A_298_294#_c_316_n
+ N_A_298_294#_c_308_n N_A_298_294#_c_318_n N_A_298_294#_c_350_p
+ N_A_298_294#_c_309_n N_A_298_294#_c_310_n N_A_298_294#_c_311_n
+ PM_SKY130_FD_SC_LS__DFRBP_2%A_298_294#
x_PM_SKY130_FD_SC_LS__DFRBP_2%RESET_B N_RESET_B_c_413_n N_RESET_B_M1015_g
+ N_RESET_B_M1009_g N_RESET_B_c_415_n N_RESET_B_c_416_n N_RESET_B_c_430_n
+ N_RESET_B_c_431_n N_RESET_B_M1032_g N_RESET_B_M1025_g N_RESET_B_c_418_n
+ N_RESET_B_M1024_g N_RESET_B_M1019_g N_RESET_B_c_420_n N_RESET_B_c_421_n
+ N_RESET_B_c_422_n N_RESET_B_c_423_n N_RESET_B_c_424_n RESET_B
+ N_RESET_B_c_425_n N_RESET_B_c_426_n N_RESET_B_c_427_n N_RESET_B_c_428_n
+ PM_SKY130_FD_SC_LS__DFRBP_2%RESET_B
x_PM_SKY130_FD_SC_LS__DFRBP_2%A_331_392# N_A_331_392#_M1034_d
+ N_A_331_392#_M1021_d N_A_331_392#_M1031_d N_A_331_392#_M1028_s
+ N_A_331_392#_M1011_g N_A_331_392#_c_613_n N_A_331_392#_c_614_n
+ N_A_331_392#_c_640_n N_A_331_392#_M1022_g N_A_331_392#_c_615_n
+ N_A_331_392#_c_616_n N_A_331_392#_c_617_n N_A_331_392#_c_618_n
+ N_A_331_392#_c_657_n N_A_331_392#_c_642_n N_A_331_392#_c_619_n
+ N_A_331_392#_c_620_n N_A_331_392#_c_621_n N_A_331_392#_c_622_n
+ N_A_331_392#_c_623_n N_A_331_392#_c_624_n N_A_331_392#_c_711_p
+ N_A_331_392#_c_625_n N_A_331_392#_c_626_n N_A_331_392#_c_627_n
+ N_A_331_392#_c_628_n N_A_331_392#_c_629_n N_A_331_392#_c_630_n
+ N_A_331_392#_c_631_n N_A_331_392#_c_632_n N_A_331_392#_c_633_n
+ N_A_331_392#_c_634_n N_A_331_392#_c_635_n N_A_331_392#_c_636_n
+ N_A_331_392#_c_637_n N_A_331_392#_c_638_n
+ PM_SKY130_FD_SC_LS__DFRBP_2%A_331_392#
x_PM_SKY130_FD_SC_LS__DFRBP_2%A_818_418# N_A_818_418#_M1030_s
+ N_A_818_418#_M1029_s N_A_818_418#_c_840_n N_A_818_418#_M1010_g
+ N_A_818_418#_M1035_g N_A_818_418#_c_842_n N_A_818_418#_M1021_g
+ N_A_818_418#_c_843_n N_A_818_418#_c_855_n N_A_818_418#_M1023_g
+ N_A_818_418#_c_844_n N_A_818_418#_c_845_n N_A_818_418#_c_846_n
+ N_A_818_418#_c_857_n N_A_818_418#_c_858_n N_A_818_418#_c_859_n
+ N_A_818_418#_c_860_n N_A_818_418#_c_861_n N_A_818_418#_c_862_n
+ N_A_818_418#_c_847_n N_A_818_418#_c_848_n N_A_818_418#_c_849_n
+ N_A_818_418#_c_850_n N_A_818_418#_c_866_n N_A_818_418#_c_851_n
+ N_A_818_418#_c_852_n PM_SKY130_FD_SC_LS__DFRBP_2%A_818_418#
x_PM_SKY130_FD_SC_LS__DFRBP_2%A_728_331# N_A_728_331#_M1003_d
+ N_A_728_331#_M1007_d N_A_728_331#_c_998_n N_A_728_331#_c_1010_n
+ N_A_728_331#_M1001_g N_A_728_331#_M1004_g N_A_728_331#_c_1000_n
+ N_A_728_331#_c_1001_n N_A_728_331#_M1030_g N_A_728_331#_c_1011_n
+ N_A_728_331#_M1029_g N_A_728_331#_c_1012_n N_A_728_331#_M1013_g
+ N_A_728_331#_c_1014_n N_A_728_331#_M1028_g N_A_728_331#_c_1004_n
+ N_A_728_331#_c_1015_n N_A_728_331#_c_1016_n N_A_728_331#_c_1108_n
+ N_A_728_331#_c_1005_n N_A_728_331#_c_1017_n N_A_728_331#_c_1038_n
+ N_A_728_331#_c_1006_n N_A_728_331#_c_1007_n N_A_728_331#_c_1040_n
+ N_A_728_331#_c_1019_n N_A_728_331#_c_1008_n N_A_728_331#_c_1021_n
+ PM_SKY130_FD_SC_LS__DFRBP_2%A_728_331#
x_PM_SKY130_FD_SC_LS__DFRBP_2%CLK N_CLK_c_1167_n N_CLK_M1003_g N_CLK_c_1168_n
+ N_CLK_M1007_g CLK PM_SKY130_FD_SC_LS__DFRBP_2%CLK
x_PM_SKY130_FD_SC_LS__DFRBP_2%A_1800_291# N_A_1800_291#_M1017_d
+ N_A_1800_291#_M1024_d N_A_1800_291#_c_1206_n N_A_1800_291#_M1018_g
+ N_A_1800_291#_c_1207_n N_A_1800_291#_c_1208_n N_A_1800_291#_M1005_g
+ N_A_1800_291#_c_1209_n N_A_1800_291#_c_1210_n N_A_1800_291#_c_1241_n
+ N_A_1800_291#_c_1245_p N_A_1800_291#_c_1211_n N_A_1800_291#_c_1230_n
+ N_A_1800_291#_c_1216_n N_A_1800_291#_c_1212_n
+ PM_SKY130_FD_SC_LS__DFRBP_2%A_1800_291#
x_PM_SKY130_FD_SC_LS__DFRBP_2%A_1586_149# N_A_1586_149#_M1013_d
+ N_A_1586_149#_M1028_d N_A_1586_149#_M1017_g N_A_1586_149#_c_1294_n
+ N_A_1586_149#_c_1303_n N_A_1586_149#_M1016_g N_A_1586_149#_c_1304_n
+ N_A_1586_149#_M1014_g N_A_1586_149#_c_1295_n N_A_1586_149#_M1006_g
+ N_A_1586_149#_c_1305_n N_A_1586_149#_M1026_g N_A_1586_149#_c_1296_n
+ N_A_1586_149#_M1036_g N_A_1586_149#_c_1306_n N_A_1586_149#_M1002_g
+ N_A_1586_149#_M1020_g N_A_1586_149#_c_1314_n N_A_1586_149#_c_1307_n
+ N_A_1586_149#_c_1298_n N_A_1586_149#_c_1299_n N_A_1586_149#_c_1309_n
+ N_A_1586_149#_c_1300_n N_A_1586_149#_c_1301_n
+ PM_SKY130_FD_SC_LS__DFRBP_2%A_1586_149#
x_PM_SKY130_FD_SC_LS__DFRBP_2%A_2363_352# N_A_2363_352#_M1020_d
+ N_A_2363_352#_M1002_d N_A_2363_352#_c_1437_n N_A_2363_352#_M1000_g
+ N_A_2363_352#_M1012_g N_A_2363_352#_c_1438_n N_A_2363_352#_M1033_g
+ N_A_2363_352#_M1037_g N_A_2363_352#_c_1433_n N_A_2363_352#_c_1440_n
+ N_A_2363_352#_c_1434_n N_A_2363_352#_c_1435_n N_A_2363_352#_c_1436_n
+ PM_SKY130_FD_SC_LS__DFRBP_2%A_2363_352#
x_PM_SKY130_FD_SC_LS__DFRBP_2%VPWR N_VPWR_M1027_s N_VPWR_M1015_d N_VPWR_M1032_d
+ N_VPWR_M1029_d N_VPWR_M1018_d N_VPWR_M1016_d N_VPWR_M1026_s N_VPWR_M1000_d
+ N_VPWR_M1033_d N_VPWR_c_1492_n N_VPWR_c_1493_n N_VPWR_c_1494_n N_VPWR_c_1495_n
+ N_VPWR_c_1496_n N_VPWR_c_1497_n N_VPWR_c_1498_n N_VPWR_c_1499_n
+ N_VPWR_c_1500_n N_VPWR_c_1501_n N_VPWR_c_1502_n N_VPWR_c_1503_n
+ N_VPWR_c_1504_n N_VPWR_c_1505_n N_VPWR_c_1506_n VPWR N_VPWR_c_1507_n
+ N_VPWR_c_1508_n N_VPWR_c_1509_n N_VPWR_c_1510_n N_VPWR_c_1511_n
+ N_VPWR_c_1512_n N_VPWR_c_1513_n N_VPWR_c_1514_n N_VPWR_c_1515_n
+ N_VPWR_c_1491_n PM_SKY130_FD_SC_LS__DFRBP_2%VPWR
x_PM_SKY130_FD_SC_LS__DFRBP_2%A_70_74# N_A_70_74#_M1008_s N_A_70_74#_M1004_s
+ N_A_70_74#_M1027_d N_A_70_74#_M1010_d N_A_70_74#_c_1639_n N_A_70_74#_c_1644_n
+ N_A_70_74#_c_1645_n N_A_70_74#_c_1646_n N_A_70_74#_c_1647_n
+ N_A_70_74#_c_1648_n N_A_70_74#_c_1649_n N_A_70_74#_c_1650_n
+ N_A_70_74#_c_1651_n N_A_70_74#_c_1652_n N_A_70_74#_c_1653_n
+ N_A_70_74#_c_1654_n N_A_70_74#_c_1640_n N_A_70_74#_c_1641_n
+ N_A_70_74#_c_1656_n N_A_70_74#_c_1657_n N_A_70_74#_c_1642_n
+ N_A_70_74#_c_1659_n N_A_70_74#_c_1643_n PM_SKY130_FD_SC_LS__DFRBP_2%A_70_74#
x_PM_SKY130_FD_SC_LS__DFRBP_2%Q_N N_Q_N_M1006_s N_Q_N_M1014_d N_Q_N_c_1793_n
+ N_Q_N_c_1791_n Q_N PM_SKY130_FD_SC_LS__DFRBP_2%Q_N
x_PM_SKY130_FD_SC_LS__DFRBP_2%Q N_Q_M1012_s N_Q_M1000_s N_Q_c_1823_n
+ N_Q_c_1824_n N_Q_c_1820_n Q N_Q_c_1822_n Q PM_SKY130_FD_SC_LS__DFRBP_2%Q
x_PM_SKY130_FD_SC_LS__DFRBP_2%VGND N_VGND_M1009_d N_VGND_M1025_s N_VGND_M1030_d
+ N_VGND_M1005_d N_VGND_M1006_d N_VGND_M1036_d N_VGND_M1012_d N_VGND_M1037_d
+ N_VGND_c_1851_n N_VGND_c_1852_n N_VGND_c_1853_n N_VGND_c_1854_n
+ N_VGND_c_1855_n N_VGND_c_1856_n N_VGND_c_1857_n N_VGND_c_1858_n
+ N_VGND_c_1859_n N_VGND_c_1860_n N_VGND_c_1861_n N_VGND_c_1862_n
+ N_VGND_c_1863_n N_VGND_c_1864_n N_VGND_c_1865_n N_VGND_c_1866_n
+ N_VGND_c_1867_n VGND N_VGND_c_1868_n N_VGND_c_1869_n N_VGND_c_1870_n
+ N_VGND_c_1871_n N_VGND_c_1872_n N_VGND_c_1873_n N_VGND_c_1874_n
+ N_VGND_c_1875_n PM_SKY130_FD_SC_LS__DFRBP_2%VGND
x_PM_SKY130_FD_SC_LS__DFRBP_2%A_614_81# N_A_614_81#_M1011_d N_A_614_81#_M1035_d
+ N_A_614_81#_c_2000_n N_A_614_81#_c_2001_n
+ PM_SKY130_FD_SC_LS__DFRBP_2%A_614_81#
x_PM_SKY130_FD_SC_LS__DFRBP_2%A_1499_149# N_A_1499_149#_M1013_s
+ N_A_1499_149#_M1005_s N_A_1499_149#_c_2024_n N_A_1499_149#_c_2025_n
+ N_A_1499_149#_c_2026_n N_A_1499_149#_c_2027_n
+ PM_SKY130_FD_SC_LS__DFRBP_2%A_1499_149#
cc_1 VNB N_D_c_269_n 0.00700378f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.795
cc_2 VNB N_D_c_270_n 0.0213314f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.9
cc_3 VNB N_D_c_271_n 0.0285408f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.05
cc_4 VNB N_D_c_272_n 0.0321996f $X=-0.19 $Y=-0.245 $X2=0.465 $Y2=1.57
cc_5 VNB D 0.0402073f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_6 VNB N_D_c_274_n 0.0259531f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.065
cc_7 VNB N_A_298_294#_M1034_g 0.0210027f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_8 VNB N_A_298_294#_c_305_n 0.00685435f $X=-0.19 $Y=-0.245 $X2=0.465 $Y2=1.065
cc_9 VNB N_A_298_294#_c_306_n 0.00372798f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=0.925
cc_10 VNB N_A_298_294#_c_307_n 0.0271085f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_298_294#_c_308_n 0.0104447f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_298_294#_c_309_n 0.00334726f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_298_294#_c_310_n 0.00112476f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_298_294#_c_311_n 3.53072e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_RESET_B_c_413_n 0.0209979f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.57
cc_16 VNB N_RESET_B_M1009_g 0.0441018f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=0.58
cc_17 VNB N_RESET_B_c_415_n 0.112144f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=0.58
cc_18 VNB N_RESET_B_c_416_n 0.0121624f $X=-0.19 $Y=-0.245 $X2=0.465 $Y2=1.05
cc_19 VNB N_RESET_B_M1025_g 0.0520604f $X=-0.19 $Y=-0.245 $X2=0.465 $Y2=1.065
cc_20 VNB N_RESET_B_c_418_n 0.0164986f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.065
cc_21 VNB N_RESET_B_M1019_g 0.0431388f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.065
cc_22 VNB N_RESET_B_c_420_n 0.00715114f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_RESET_B_c_421_n 0.00143791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_RESET_B_c_422_n 0.0394685f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_RESET_B_c_423_n 5.88447e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_RESET_B_c_424_n 0.0015362f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_RESET_B_c_425_n 0.00161047f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_RESET_B_c_426_n 0.0180398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_RESET_B_c_427_n 0.00361963f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_RESET_B_c_428_n 0.00386078f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_331_392#_c_613_n 0.0270185f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_331_392#_c_614_n 0.0234715f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.065
cc_33 VNB N_A_331_392#_c_615_n 0.0156643f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_331_392#_c_616_n 0.0113755f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.065
cc_35 VNB N_A_331_392#_c_617_n 0.00229509f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_331_392#_c_618_n 0.0090728f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_331_392#_c_619_n 0.0199884f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_331_392#_c_620_n 0.00387155f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_331_392#_c_621_n 0.0371118f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_331_392#_c_622_n 0.00225927f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_331_392#_c_623_n 0.00311976f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_331_392#_c_624_n 0.00704603f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_331_392#_c_625_n 0.0035579f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_331_392#_c_626_n 0.00153929f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_331_392#_c_627_n 0.0293297f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_331_392#_c_628_n 0.00355388f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_331_392#_c_629_n 0.0273514f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_331_392#_c_630_n 0.0270442f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_331_392#_c_631_n 0.0108619f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_331_392#_c_632_n 0.00314018f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_331_392#_c_633_n 0.00175721f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_331_392#_c_634_n 2.56805e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_331_392#_c_635_n 0.00402758f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_331_392#_c_636_n 4.63774e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_331_392#_c_637_n 0.00230646f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_331_392#_c_638_n 0.0440154f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_818_418#_c_840_n 0.0118362f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=0.58
cc_58 VNB N_A_818_418#_M1035_g 0.040937f $X=-0.19 $Y=-0.245 $X2=0.465 $Y2=1.325
cc_59 VNB N_A_818_418#_c_842_n 0.0204366f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_818_418#_c_843_n 0.00292692f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.065
cc_61 VNB N_A_818_418#_c_844_n 0.0168787f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.295
cc_62 VNB N_A_818_418#_c_845_n 0.0222244f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_818_418#_c_846_n 0.0117883f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_818_418#_c_847_n 6.24838e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_818_418#_c_848_n 0.00117943f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_818_418#_c_849_n 0.0420897f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_818_418#_c_850_n 0.00139432f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_818_418#_c_851_n 0.00520919f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_818_418#_c_852_n 0.0492887f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_728_331#_c_998_n 0.0220127f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=0.58
cc_71 VNB N_A_728_331#_M1004_g 0.0615892f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_72 VNB N_A_728_331#_c_1000_n 0.111851f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_728_331#_c_1001_n 0.0102577f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_728_331#_M1030_g 0.0143554f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=0.925
cc_75 VNB N_A_728_331#_M1013_g 0.0439787f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_728_331#_c_1004_n 0.0147342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_728_331#_c_1005_n 0.00412543f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_728_331#_c_1006_n 0.00496454f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_728_331#_c_1007_n 0.00414255f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_728_331#_c_1008_n 0.0664181f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_CLK_c_1167_n 0.0206637f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.57
cc_82 VNB N_CLK_c_1168_n 0.0389797f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=2.17
cc_83 VNB CLK 0.00912873f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=0.58
cc_84 VNB N_A_1800_291#_c_1206_n 0.0178321f $X=-0.19 $Y=-0.245 $X2=0.705
+ $Y2=0.58
cc_85 VNB N_A_1800_291#_c_1207_n 0.0271658f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.05
cc_86 VNB N_A_1800_291#_c_1208_n 0.0185916f $X=-0.19 $Y=-0.245 $X2=0.465
+ $Y2=1.325
cc_87 VNB N_A_1800_291#_c_1209_n 0.0210915f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_1800_291#_c_1210_n 0.00103268f $X=-0.19 $Y=-0.245 $X2=0.32
+ $Y2=0.925
cc_89 VNB N_A_1800_291#_c_1211_n 0.00794995f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_1800_291#_c_1212_n 0.00950159f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_1586_149#_M1017_g 0.021266f $X=-0.19 $Y=-0.245 $X2=0.465 $Y2=1.05
cc_92 VNB N_A_1586_149#_c_1294_n 0.001735f $X=-0.19 $Y=-0.245 $X2=0.465
+ $Y2=1.325
cc_93 VNB N_A_1586_149#_c_1295_n 0.0164413f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.065
cc_94 VNB N_A_1586_149#_c_1296_n 0.0144188f $X=-0.19 $Y=-0.245 $X2=0.32
+ $Y2=1.295
cc_95 VNB N_A_1586_149#_M1020_g 0.0229039f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_1586_149#_c_1298_n 0.00303624f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_1586_149#_c_1299_n 0.02459f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_A_1586_149#_c_1300_n 0.00358249f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_A_1586_149#_c_1301_n 0.151485f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_A_2363_352#_M1012_g 0.0234349f $X=-0.19 $Y=-0.245 $X2=0.465
+ $Y2=1.325
cc_101 VNB N_A_2363_352#_M1037_g 0.0265988f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.065
cc_102 VNB N_A_2363_352#_c_1433_n 0.00718732f $X=-0.19 $Y=-0.245 $X2=0.32
+ $Y2=0.925
cc_103 VNB N_A_2363_352#_c_1434_n 0.0169817f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_A_2363_352#_c_1435_n 0.0109542f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_A_2363_352#_c_1436_n 0.0860723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_VPWR_c_1491_n 0.581632f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_A_70_74#_c_1639_n 0.0104114f $X=-0.19 $Y=-0.245 $X2=0.465 $Y2=1.57
cc_108 VNB N_A_70_74#_c_1640_n 0.00974934f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_A_70_74#_c_1641_n 0.00594127f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_A_70_74#_c_1642_n 0.00740588f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_A_70_74#_c_1643_n 0.00977141f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_Q_N_c_1791_n 0.00215184f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_113 VNB Q_N 5.1574e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_Q_c_1820_n 0.00335076f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_115 VNB Q 0.00448002f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_Q_c_1822_n 0.00232136f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=0.925
cc_117 VNB N_VGND_c_1851_n 0.0101803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_VGND_c_1852_n 0.0113244f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_VGND_c_1853_n 0.00652305f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_VGND_c_1854_n 0.00396467f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_VGND_c_1855_n 0.00782424f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_VGND_c_1856_n 0.00524489f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB N_VGND_c_1857_n 0.0168886f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_VGND_c_1858_n 0.0103919f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_1859_n 0.0515355f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_1860_n 0.0190288f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_VGND_c_1861_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_1862_n 0.071262f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_1863_n 0.00477852f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_1864_n 0.0835402f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_1865_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_VGND_c_1866_n 0.0311181f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_VGND_c_1867_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_VGND_c_1868_n 0.0337099f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_VGND_c_1869_n 0.0171743f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_VGND_c_1870_n 0.0188091f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_VGND_c_1871_n 0.0189106f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB N_VGND_c_1872_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VNB N_VGND_c_1873_n 0.00632462f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_VGND_c_1874_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_141 VNB N_VGND_c_1875_n 0.736558f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_142 VNB N_A_614_81#_c_2000_n 0.0302536f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=0.58
cc_143 VNB N_A_614_81#_c_2001_n 0.0209611f $X=-0.19 $Y=-0.245 $X2=0.465 $Y2=1.57
cc_144 VNB N_A_1499_149#_c_2024_n 0.00155523f $X=-0.19 $Y=-0.245 $X2=0.465
+ $Y2=1.05
cc_145 VNB N_A_1499_149#_c_2025_n 0.00899648f $X=-0.19 $Y=-0.245 $X2=0.5
+ $Y2=1.05
cc_146 VNB N_A_1499_149#_c_2026_n 0.00304708f $X=-0.19 $Y=-0.245 $X2=0.465
+ $Y2=1.325
cc_147 VNB N_A_1499_149#_c_2027_n 0.00653449f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=0.84
cc_148 VPB N_D_c_269_n 0.0105518f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=1.795
cc_149 VPB N_D_c_276_n 0.0250353f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=1.885
cc_150 VPB N_A_298_294#_c_312_n 0.0179938f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=0.9
cc_151 VPB N_A_298_294#_c_305_n 0.00947655f $X=-0.19 $Y=1.66 $X2=0.465 $Y2=1.065
cc_152 VPB N_A_298_294#_c_306_n 0.0035383f $X=-0.19 $Y=1.66 $X2=0.32 $Y2=0.925
cc_153 VPB N_A_298_294#_c_307_n 0.0224362f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_154 VPB N_A_298_294#_c_316_n 0.0123517f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_155 VPB N_A_298_294#_c_308_n 0.00925129f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_156 VPB N_A_298_294#_c_318_n 0.0135945f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_157 VPB N_RESET_B_c_413_n 0.0340437f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=1.57
cc_158 VPB N_RESET_B_c_430_n 0.0333511f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=1.05
cc_159 VPB N_RESET_B_c_431_n 0.0252042f $X=-0.19 $Y=1.66 $X2=0.465 $Y2=1.325
cc_160 VPB N_RESET_B_c_418_n 0.0358088f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.065
cc_161 VPB N_RESET_B_c_420_n 0.00666344f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_162 VPB N_RESET_B_c_421_n 0.00720642f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_163 VPB N_RESET_B_c_422_n 0.0265356f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_164 VPB N_RESET_B_c_423_n 0.00122693f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_165 VPB N_RESET_B_c_424_n 0.00230825f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_166 VPB N_RESET_B_c_425_n 8.04582e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_167 VPB N_RESET_B_c_426_n 0.00972568f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_168 VPB N_RESET_B_c_427_n 0.00100868f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_169 VPB N_RESET_B_c_428_n 0.00189077f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_170 VPB N_A_331_392#_c_614_n 9.02379e-19 $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.065
cc_171 VPB N_A_331_392#_c_640_n 0.0208595f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.065
cc_172 VPB N_A_331_392#_c_617_n 0.00231184f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_173 VPB N_A_331_392#_c_642_n 0.00186964f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_174 VPB N_A_331_392#_c_633_n 0.0016526f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_175 VPB N_A_331_392#_c_636_n 3.96019e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_176 VPB N_A_331_392#_c_638_n 0.00661599f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_177 VPB N_A_818_418#_c_840_n 0.0221279f $X=-0.19 $Y=1.66 $X2=0.705 $Y2=0.58
cc_178 VPB N_A_818_418#_c_843_n 0.00645031f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.065
cc_179 VPB N_A_818_418#_c_855_n 0.0240905f $X=-0.19 $Y=1.66 $X2=0.32 $Y2=0.925
cc_180 VPB N_A_818_418#_c_846_n 0.00235496f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_181 VPB N_A_818_418#_c_857_n 0.00704052f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_182 VPB N_A_818_418#_c_858_n 0.0130792f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_183 VPB N_A_818_418#_c_859_n 0.012711f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_184 VPB N_A_818_418#_c_860_n 0.00911703f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_185 VPB N_A_818_418#_c_861_n 0.0165779f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_186 VPB N_A_818_418#_c_862_n 0.0053835f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_187 VPB N_A_818_418#_c_847_n 0.0028531f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_188 VPB N_A_818_418#_c_849_n 0.0194541f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_189 VPB N_A_818_418#_c_850_n 0.00504835f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_190 VPB N_A_818_418#_c_866_n 0.00436524f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_191 VPB N_A_728_331#_c_998_n 6.78857e-19 $X=-0.19 $Y=1.66 $X2=0.705 $Y2=0.58
cc_192 VPB N_A_728_331#_c_1010_n 0.0191535f $X=-0.19 $Y=1.66 $X2=0.465 $Y2=1.05
cc_193 VPB N_A_728_331#_c_1011_n 0.0216648f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_194 VPB N_A_728_331#_c_1012_n 0.0206163f $X=-0.19 $Y=1.66 $X2=0.32 $Y2=1.295
cc_195 VPB N_A_728_331#_M1013_g 0.00409839f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_196 VPB N_A_728_331#_c_1014_n 0.0177979f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_197 VPB N_A_728_331#_c_1015_n 0.016648f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_198 VPB N_A_728_331#_c_1016_n 0.00357702f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_199 VPB N_A_728_331#_c_1017_n 0.00529591f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_200 VPB N_A_728_331#_c_1006_n 8.76898e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_201 VPB N_A_728_331#_c_1019_n 0.0017718f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_202 VPB N_A_728_331#_c_1008_n 0.0314894f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_203 VPB N_A_728_331#_c_1021_n 0.0505879f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_204 VPB N_CLK_c_1168_n 0.0352067f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=2.17
cc_205 VPB CLK 0.00114738f $X=-0.19 $Y=1.66 $X2=0.705 $Y2=0.58
cc_206 VPB N_A_1800_291#_c_1206_n 0.0367404f $X=-0.19 $Y=1.66 $X2=0.705 $Y2=0.58
cc_207 VPB N_A_1800_291#_c_1210_n 0.00189897f $X=-0.19 $Y=1.66 $X2=0.32
+ $Y2=0.925
cc_208 VPB N_A_1800_291#_c_1211_n 0.0017906f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_209 VPB N_A_1800_291#_c_1216_n 0.011565f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_210 VPB N_A_1586_149#_c_1294_n 0.00853434f $X=-0.19 $Y=1.66 $X2=0.465
+ $Y2=1.325
cc_211 VPB N_A_1586_149#_c_1303_n 0.0238482f $X=-0.19 $Y=1.66 $X2=0.465 $Y2=1.57
cc_212 VPB N_A_1586_149#_c_1304_n 0.0162194f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_213 VPB N_A_1586_149#_c_1305_n 0.016092f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_214 VPB N_A_1586_149#_c_1306_n 0.0176465f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_215 VPB N_A_1586_149#_c_1307_n 0.00876015f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_216 VPB N_A_1586_149#_c_1298_n 0.00171972f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_217 VPB N_A_1586_149#_c_1309_n 0.00185057f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_218 VPB N_A_1586_149#_c_1301_n 0.0638912f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_219 VPB N_A_2363_352#_c_1437_n 0.0166433f $X=-0.19 $Y=1.66 $X2=0.705 $Y2=0.58
cc_220 VPB N_A_2363_352#_c_1438_n 0.0174014f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=0.84
cc_221 VPB N_A_2363_352#_c_1433_n 0.0138325f $X=-0.19 $Y=1.66 $X2=0.32 $Y2=0.925
cc_222 VPB N_A_2363_352#_c_1440_n 0.01441f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_223 VPB N_A_2363_352#_c_1436_n 0.0176483f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_224 VPB N_VPWR_c_1492_n 0.0213265f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_225 VPB N_VPWR_c_1493_n 0.0551839f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_226 VPB N_VPWR_c_1494_n 0.0105306f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_227 VPB N_VPWR_c_1495_n 0.0722425f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_228 VPB N_VPWR_c_1496_n 0.0599193f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_229 VPB N_VPWR_c_1497_n 0.0301846f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_230 VPB N_VPWR_c_1498_n 0.0169533f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_231 VPB N_VPWR_c_1499_n 0.017438f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_232 VPB N_VPWR_c_1500_n 0.0281699f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_233 VPB N_VPWR_c_1501_n 0.0121909f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_234 VPB N_VPWR_c_1502_n 0.0684963f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_235 VPB N_VPWR_c_1503_n 0.014661f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_236 VPB N_VPWR_c_1504_n 0.00780326f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_237 VPB N_VPWR_c_1505_n 0.0234846f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_238 VPB N_VPWR_c_1506_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_239 VPB N_VPWR_c_1507_n 0.0359407f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_240 VPB N_VPWR_c_1508_n 0.0763132f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_241 VPB N_VPWR_c_1509_n 0.0257899f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_242 VPB N_VPWR_c_1510_n 0.0186948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_243 VPB N_VPWR_c_1511_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_244 VPB N_VPWR_c_1512_n 0.0212004f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_245 VPB N_VPWR_c_1513_n 0.00689862f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_246 VPB N_VPWR_c_1514_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_247 VPB N_VPWR_c_1515_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_248 VPB N_VPWR_c_1491_n 0.218899f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_249 VPB N_A_70_74#_c_1644_n 0.00437214f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_250 VPB N_A_70_74#_c_1645_n 0.00263879f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.065
cc_251 VPB N_A_70_74#_c_1646_n 0.00731839f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_252 VPB N_A_70_74#_c_1647_n 0.00554076f $X=-0.19 $Y=1.66 $X2=0.32 $Y2=1.065
cc_253 VPB N_A_70_74#_c_1648_n 0.0235134f $X=-0.19 $Y=1.66 $X2=0.32 $Y2=1.295
cc_254 VPB N_A_70_74#_c_1649_n 4.20701e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_255 VPB N_A_70_74#_c_1650_n 0.0064597f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_256 VPB N_A_70_74#_c_1651_n 8.66945e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_257 VPB N_A_70_74#_c_1652_n 5.49566e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_258 VPB N_A_70_74#_c_1653_n 0.0123144f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_259 VPB N_A_70_74#_c_1654_n 0.00217659f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_260 VPB N_A_70_74#_c_1641_n 0.00660556f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_261 VPB N_A_70_74#_c_1656_n 0.0117694f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_262 VPB N_A_70_74#_c_1657_n 0.00592749f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_263 VPB N_A_70_74#_c_1642_n 0.00217734f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_264 VPB N_A_70_74#_c_1659_n 0.00118567f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_265 VPB N_Q_N_c_1793_n 0.00441342f $X=-0.19 $Y=1.66 $X2=0.465 $Y2=1.05
cc_266 VPB N_Q_c_1823_n 0.00166049f $X=-0.19 $Y=1.66 $X2=0.465 $Y2=1.05
cc_267 VPB N_Q_c_1824_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=1.05
cc_268 VPB N_Q_c_1820_n 0.00149334f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_269 N_D_c_269_n N_RESET_B_c_413_n 0.00447539f $X=0.62 $Y=1.795 $X2=-0.19
+ $Y2=-0.245
cc_270 N_D_c_276_n N_RESET_B_c_413_n 0.00936496f $X=0.62 $Y=1.885 $X2=-0.19
+ $Y2=-0.245
cc_271 N_D_c_272_n N_RESET_B_c_413_n 0.0171542f $X=0.465 $Y=1.57 $X2=-0.19
+ $Y2=-0.245
cc_272 N_D_c_271_n N_RESET_B_M1009_g 0.0204298f $X=0.5 $Y=1.05 $X2=0 $Y2=0
cc_273 N_D_c_274_n N_RESET_B_M1009_g 0.0141785f $X=0.385 $Y=1.065 $X2=0 $Y2=0
cc_274 N_D_c_270_n N_RESET_B_c_416_n 0.0204298f $X=0.5 $Y=0.9 $X2=0 $Y2=0
cc_275 N_D_c_272_n N_RESET_B_c_425_n 2.85099e-19 $X=0.465 $Y=1.57 $X2=0 $Y2=0
cc_276 N_D_c_276_n N_VPWR_c_1493_n 0.0116836f $X=0.62 $Y=1.885 $X2=0 $Y2=0
cc_277 N_D_c_272_n N_VPWR_c_1493_n 0.00205106f $X=0.465 $Y=1.57 $X2=0 $Y2=0
cc_278 D N_VPWR_c_1493_n 0.0195039f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_279 N_D_c_276_n N_VPWR_c_1503_n 0.00466109f $X=0.62 $Y=1.885 $X2=0 $Y2=0
cc_280 N_D_c_270_n N_A_70_74#_c_1639_n 0.00876622f $X=0.5 $Y=0.9 $X2=0 $Y2=0
cc_281 N_D_c_271_n N_A_70_74#_c_1639_n 0.00462754f $X=0.5 $Y=1.05 $X2=0 $Y2=0
cc_282 D N_A_70_74#_c_1639_n 0.0156724f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_283 N_D_c_276_n N_A_70_74#_c_1644_n 0.00201741f $X=0.62 $Y=1.885 $X2=0 $Y2=0
cc_284 N_D_c_276_n N_A_70_74#_c_1645_n 0.00594681f $X=0.62 $Y=1.885 $X2=0 $Y2=0
cc_285 N_D_c_269_n N_A_70_74#_c_1642_n 0.0104907f $X=0.62 $Y=1.795 $X2=0 $Y2=0
cc_286 N_D_c_276_n N_A_70_74#_c_1642_n 0.00738787f $X=0.62 $Y=1.885 $X2=0 $Y2=0
cc_287 N_D_c_270_n N_A_70_74#_c_1642_n 0.0102779f $X=0.5 $Y=0.9 $X2=0 $Y2=0
cc_288 N_D_c_271_n N_A_70_74#_c_1642_n 0.00579508f $X=0.5 $Y=1.05 $X2=0 $Y2=0
cc_289 N_D_c_272_n N_A_70_74#_c_1642_n 0.00565081f $X=0.465 $Y=1.57 $X2=0 $Y2=0
cc_290 D N_A_70_74#_c_1642_n 0.0551626f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_291 N_D_c_274_n N_A_70_74#_c_1642_n 0.00652495f $X=0.385 $Y=1.065 $X2=0 $Y2=0
cc_292 N_D_c_270_n N_VGND_c_1851_n 0.00115926f $X=0.5 $Y=0.9 $X2=0 $Y2=0
cc_293 N_D_c_270_n N_VGND_c_1868_n 0.00296902f $X=0.5 $Y=0.9 $X2=0 $Y2=0
cc_294 N_D_c_270_n N_VGND_c_1875_n 0.00367837f $X=0.5 $Y=0.9 $X2=0 $Y2=0
cc_295 D N_VGND_c_1875_n 0.00842173f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_296 N_A_298_294#_c_312_n N_RESET_B_c_413_n 0.0189712f $X=1.58 $Y=1.885
+ $X2=-0.19 $Y2=-0.245
cc_297 N_A_298_294#_M1034_g N_RESET_B_c_413_n 0.00107375f $X=1.595 $Y=0.965
+ $X2=-0.19 $Y2=-0.245
cc_298 N_A_298_294#_c_305_n N_RESET_B_c_413_n 0.0237815f $X=1.58 $Y=1.677
+ $X2=-0.19 $Y2=-0.245
cc_299 N_A_298_294#_M1034_g N_RESET_B_M1009_g 0.0247767f $X=1.595 $Y=0.965 $X2=0
+ $Y2=0
cc_300 N_A_298_294#_M1034_g N_RESET_B_c_415_n 0.0101835f $X=1.595 $Y=0.965 $X2=0
+ $Y2=0
cc_301 N_A_298_294#_c_306_n N_RESET_B_c_430_n 0.00477445f $X=1.99 $Y=1.635 $X2=0
+ $Y2=0
cc_302 N_A_298_294#_c_307_n N_RESET_B_c_430_n 0.00105273f $X=1.99 $Y=1.635 $X2=0
+ $Y2=0
cc_303 N_A_298_294#_c_316_n N_RESET_B_c_430_n 0.00856912f $X=2.35 $Y=2.57 $X2=0
+ $Y2=0
cc_304 N_A_298_294#_c_308_n N_RESET_B_c_430_n 0.0184509f $X=3.79 $Y=2.03 $X2=0
+ $Y2=0
cc_305 N_A_298_294#_c_316_n N_RESET_B_c_431_n 0.00254499f $X=2.35 $Y=2.57 $X2=0
+ $Y2=0
cc_306 N_A_298_294#_c_305_n N_RESET_B_c_420_n 3.63e-19 $X=1.58 $Y=1.677 $X2=0
+ $Y2=0
cc_307 N_A_298_294#_c_306_n N_RESET_B_c_420_n 0.0168912f $X=1.99 $Y=1.635 $X2=0
+ $Y2=0
cc_308 N_A_298_294#_c_307_n N_RESET_B_c_420_n 0.00425279f $X=1.99 $Y=1.635 $X2=0
+ $Y2=0
cc_309 N_A_298_294#_c_318_n N_RESET_B_c_420_n 0.0122224f $X=2.435 $Y=2.03 $X2=0
+ $Y2=0
cc_310 N_A_298_294#_c_308_n N_RESET_B_c_422_n 0.0243589f $X=3.79 $Y=2.03 $X2=0
+ $Y2=0
cc_311 N_A_298_294#_c_309_n N_RESET_B_c_422_n 0.0190818f $X=4.002 $Y=1.945 $X2=0
+ $Y2=0
cc_312 N_A_298_294#_c_310_n N_RESET_B_c_422_n 0.00433885f $X=3.955 $Y=2.03 $X2=0
+ $Y2=0
cc_313 N_A_298_294#_c_311_n N_RESET_B_c_422_n 0.00550817f $X=4.05 $Y=1.44 $X2=0
+ $Y2=0
cc_314 N_A_298_294#_c_306_n N_RESET_B_c_423_n 6.49536e-19 $X=1.99 $Y=1.635 $X2=0
+ $Y2=0
cc_315 N_A_298_294#_c_308_n N_RESET_B_c_423_n 0.00789264f $X=3.79 $Y=2.03 $X2=0
+ $Y2=0
cc_316 N_A_298_294#_c_305_n N_RESET_B_c_425_n 8.3331e-19 $X=1.58 $Y=1.677 $X2=0
+ $Y2=0
cc_317 N_A_298_294#_M1034_g N_RESET_B_c_426_n 3.7765e-19 $X=1.595 $Y=0.965 $X2=0
+ $Y2=0
cc_318 N_A_298_294#_c_306_n N_RESET_B_c_426_n 4.89963e-19 $X=1.99 $Y=1.635 $X2=0
+ $Y2=0
cc_319 N_A_298_294#_c_307_n N_RESET_B_c_426_n 0.0184325f $X=1.99 $Y=1.635 $X2=0
+ $Y2=0
cc_320 N_A_298_294#_c_308_n N_RESET_B_c_426_n 8.73334e-19 $X=3.79 $Y=2.03 $X2=0
+ $Y2=0
cc_321 N_A_298_294#_c_318_n N_RESET_B_c_426_n 0.00223986f $X=2.435 $Y=2.03 $X2=0
+ $Y2=0
cc_322 N_A_298_294#_c_306_n N_RESET_B_c_427_n 0.01583f $X=1.99 $Y=1.635 $X2=0
+ $Y2=0
cc_323 N_A_298_294#_c_307_n N_RESET_B_c_427_n 0.00119402f $X=1.99 $Y=1.635 $X2=0
+ $Y2=0
cc_324 N_A_298_294#_c_318_n N_RESET_B_c_427_n 0.0235047f $X=2.435 $Y=2.03 $X2=0
+ $Y2=0
cc_325 N_A_298_294#_c_318_n N_A_331_392#_M1031_d 0.00353399f $X=2.435 $Y=2.03
+ $X2=0 $Y2=0
cc_326 N_A_298_294#_c_308_n N_A_331_392#_c_614_n 0.0132418f $X=3.79 $Y=2.03
+ $X2=0 $Y2=0
cc_327 N_A_298_294#_c_350_p N_A_331_392#_c_614_n 8.15911e-19 $X=3.955 $Y=2.57
+ $X2=0 $Y2=0
cc_328 N_A_298_294#_c_350_p N_A_331_392#_c_640_n 3.92955e-19 $X=3.955 $Y=2.57
+ $X2=0 $Y2=0
cc_329 N_A_298_294#_c_312_n N_A_331_392#_c_617_n 0.009572f $X=1.58 $Y=1.885
+ $X2=0 $Y2=0
cc_330 N_A_298_294#_M1034_g N_A_331_392#_c_617_n 0.015464f $X=1.595 $Y=0.965
+ $X2=0 $Y2=0
cc_331 N_A_298_294#_c_305_n N_A_331_392#_c_617_n 0.0123246f $X=1.58 $Y=1.677
+ $X2=0 $Y2=0
cc_332 N_A_298_294#_c_306_n N_A_331_392#_c_617_n 0.0333362f $X=1.99 $Y=1.635
+ $X2=0 $Y2=0
cc_333 N_A_298_294#_c_316_n N_A_331_392#_c_617_n 0.00575306f $X=2.35 $Y=2.57
+ $X2=0 $Y2=0
cc_334 N_A_298_294#_c_318_n N_A_331_392#_c_617_n 0.013285f $X=2.435 $Y=2.03
+ $X2=0 $Y2=0
cc_335 N_A_298_294#_M1034_g N_A_331_392#_c_618_n 0.0101625f $X=1.595 $Y=0.965
+ $X2=0 $Y2=0
cc_336 N_A_298_294#_c_312_n N_A_331_392#_c_657_n 0.00542396f $X=1.58 $Y=1.885
+ $X2=0 $Y2=0
cc_337 N_A_298_294#_c_307_n N_A_331_392#_c_642_n 0.00366094f $X=1.99 $Y=1.635
+ $X2=0 $Y2=0
cc_338 N_A_298_294#_c_316_n N_A_331_392#_c_642_n 0.0120222f $X=2.35 $Y=2.57
+ $X2=0 $Y2=0
cc_339 N_A_298_294#_c_318_n N_A_331_392#_c_642_n 0.0102734f $X=2.435 $Y=2.03
+ $X2=0 $Y2=0
cc_340 N_A_298_294#_c_306_n N_A_331_392#_c_619_n 0.00825186f $X=1.99 $Y=1.635
+ $X2=0 $Y2=0
cc_341 N_A_298_294#_c_307_n N_A_331_392#_c_619_n 0.00112891f $X=1.99 $Y=1.635
+ $X2=0 $Y2=0
cc_342 N_A_298_294#_M1034_g N_A_331_392#_c_634_n 0.00981844f $X=1.595 $Y=0.965
+ $X2=0 $Y2=0
cc_343 N_A_298_294#_c_306_n N_A_331_392#_c_634_n 0.00744795f $X=1.99 $Y=1.635
+ $X2=0 $Y2=0
cc_344 N_A_298_294#_c_307_n N_A_331_392#_c_634_n 0.00600011f $X=1.99 $Y=1.635
+ $X2=0 $Y2=0
cc_345 N_A_298_294#_c_308_n N_A_331_392#_c_636_n 0.021845f $X=3.79 $Y=2.03 $X2=0
+ $Y2=0
cc_346 N_A_298_294#_c_311_n N_A_331_392#_c_636_n 0.00328107f $X=4.05 $Y=1.44
+ $X2=0 $Y2=0
cc_347 N_A_298_294#_c_308_n N_A_331_392#_c_638_n 0.00855282f $X=3.79 $Y=2.03
+ $X2=0 $Y2=0
cc_348 N_A_298_294#_c_311_n N_A_331_392#_c_638_n 0.00106934f $X=4.05 $Y=1.44
+ $X2=0 $Y2=0
cc_349 N_A_298_294#_c_350_p N_A_818_418#_c_840_n 0.0114334f $X=3.955 $Y=2.57
+ $X2=0 $Y2=0
cc_350 N_A_298_294#_c_310_n N_A_818_418#_c_840_n 0.00148297f $X=3.955 $Y=2.03
+ $X2=0 $Y2=0
cc_351 N_A_298_294#_c_311_n N_A_818_418#_c_840_n 3.65173e-19 $X=4.05 $Y=1.44
+ $X2=0 $Y2=0
cc_352 N_A_298_294#_c_309_n N_A_818_418#_M1035_g 0.00241812f $X=4.002 $Y=1.945
+ $X2=0 $Y2=0
cc_353 N_A_298_294#_c_310_n N_A_818_418#_M1035_g 0.00133552f $X=3.955 $Y=2.03
+ $X2=0 $Y2=0
cc_354 N_A_298_294#_c_308_n N_A_728_331#_c_998_n 0.0129563f $X=3.79 $Y=2.03
+ $X2=0 $Y2=0
cc_355 N_A_298_294#_c_350_p N_A_728_331#_c_998_n 0.00424115f $X=3.955 $Y=2.57
+ $X2=0 $Y2=0
cc_356 N_A_298_294#_c_309_n N_A_728_331#_c_998_n 0.00367203f $X=4.002 $Y=1.945
+ $X2=0 $Y2=0
cc_357 N_A_298_294#_c_310_n N_A_728_331#_c_998_n 0.00312435f $X=3.955 $Y=2.03
+ $X2=0 $Y2=0
cc_358 N_A_298_294#_c_350_p N_A_728_331#_c_1010_n 0.00806344f $X=3.955 $Y=2.57
+ $X2=0 $Y2=0
cc_359 N_A_298_294#_c_309_n N_A_728_331#_M1004_g 0.00100194f $X=4.002 $Y=1.945
+ $X2=0 $Y2=0
cc_360 N_A_298_294#_c_311_n N_A_728_331#_M1004_g 0.00895915f $X=4.05 $Y=1.44
+ $X2=0 $Y2=0
cc_361 N_A_298_294#_c_309_n N_A_728_331#_c_1004_n 0.00470135f $X=4.002 $Y=1.945
+ $X2=0 $Y2=0
cc_362 N_A_298_294#_c_310_n N_A_728_331#_c_1004_n 0.00324895f $X=3.955 $Y=2.03
+ $X2=0 $Y2=0
cc_363 N_A_298_294#_c_312_n N_VPWR_c_1504_n 0.00309988f $X=1.58 $Y=1.885 $X2=0
+ $Y2=0
cc_364 N_A_298_294#_c_312_n N_VPWR_c_1507_n 0.00303904f $X=1.58 $Y=1.885 $X2=0
+ $Y2=0
cc_365 N_A_298_294#_c_312_n N_VPWR_c_1491_n 0.00386627f $X=1.58 $Y=1.885 $X2=0
+ $Y2=0
cc_366 N_A_298_294#_c_312_n N_A_70_74#_c_1644_n 5.17802e-19 $X=1.58 $Y=1.885
+ $X2=0 $Y2=0
cc_367 N_A_298_294#_c_312_n N_A_70_74#_c_1645_n 0.00327344f $X=1.58 $Y=1.885
+ $X2=0 $Y2=0
cc_368 N_A_298_294#_c_312_n N_A_70_74#_c_1646_n 0.00931811f $X=1.58 $Y=1.885
+ $X2=0 $Y2=0
cc_369 N_A_298_294#_c_312_n N_A_70_74#_c_1648_n 0.00102155f $X=1.58 $Y=1.885
+ $X2=0 $Y2=0
cc_370 N_A_298_294#_c_316_n N_A_70_74#_c_1648_n 0.0191246f $X=2.35 $Y=2.57 $X2=0
+ $Y2=0
cc_371 N_A_298_294#_c_316_n N_A_70_74#_c_1649_n 0.0202279f $X=2.35 $Y=2.57 $X2=0
+ $Y2=0
cc_372 N_A_298_294#_c_308_n N_A_70_74#_c_1650_n 0.0555839f $X=3.79 $Y=2.03 $X2=0
+ $Y2=0
cc_373 N_A_298_294#_c_350_p N_A_70_74#_c_1650_n 0.0105082f $X=3.955 $Y=2.57
+ $X2=0 $Y2=0
cc_374 N_A_298_294#_c_316_n N_A_70_74#_c_1651_n 0.0138867f $X=2.35 $Y=2.57 $X2=0
+ $Y2=0
cc_375 N_A_298_294#_c_308_n N_A_70_74#_c_1651_n 0.0133351f $X=3.79 $Y=2.03 $X2=0
+ $Y2=0
cc_376 N_A_298_294#_c_350_p N_A_70_74#_c_1652_n 0.0151127f $X=3.955 $Y=2.57
+ $X2=0 $Y2=0
cc_377 N_A_298_294#_c_350_p N_A_70_74#_c_1653_n 0.0206353f $X=3.955 $Y=2.57
+ $X2=0 $Y2=0
cc_378 N_A_298_294#_c_311_n N_A_70_74#_c_1640_n 0.0169762f $X=4.05 $Y=1.44 $X2=0
+ $Y2=0
cc_379 N_A_298_294#_c_350_p N_A_70_74#_c_1641_n 0.0202223f $X=3.955 $Y=2.57
+ $X2=0 $Y2=0
cc_380 N_A_298_294#_c_309_n N_A_70_74#_c_1641_n 0.0221864f $X=4.002 $Y=1.945
+ $X2=0 $Y2=0
cc_381 N_A_298_294#_c_310_n N_A_70_74#_c_1641_n 0.0127253f $X=3.955 $Y=2.03
+ $X2=0 $Y2=0
cc_382 N_A_298_294#_c_311_n N_A_70_74#_c_1641_n 0.0124256f $X=4.05 $Y=1.44 $X2=0
+ $Y2=0
cc_383 N_A_298_294#_c_350_p N_A_70_74#_c_1656_n 0.0127893f $X=3.955 $Y=2.57
+ $X2=0 $Y2=0
cc_384 N_A_298_294#_c_312_n N_A_70_74#_c_1659_n 0.0183637f $X=1.58 $Y=1.885
+ $X2=0 $Y2=0
cc_385 N_A_298_294#_c_316_n N_A_70_74#_c_1659_n 0.00447891f $X=2.35 $Y=2.57
+ $X2=0 $Y2=0
cc_386 N_A_298_294#_c_308_n N_A_70_74#_c_1643_n 0.00484801f $X=3.79 $Y=2.03
+ $X2=0 $Y2=0
cc_387 N_A_298_294#_M1034_g N_VGND_c_1851_n 0.002225f $X=1.595 $Y=0.965 $X2=0
+ $Y2=0
cc_388 N_A_298_294#_M1034_g N_VGND_c_1852_n 8.31286e-19 $X=1.595 $Y=0.965 $X2=0
+ $Y2=0
cc_389 N_A_298_294#_M1034_g N_VGND_c_1875_n 7.88961e-19 $X=1.595 $Y=0.965 $X2=0
+ $Y2=0
cc_390 N_RESET_B_M1025_g N_A_331_392#_c_613_n 0.0171459f $X=2.605 $Y=0.615 $X2=0
+ $Y2=0
cc_391 N_RESET_B_c_426_n N_A_331_392#_c_613_n 0.00381284f $X=2.55 $Y=1.61 $X2=0
+ $Y2=0
cc_392 N_RESET_B_c_427_n N_A_331_392#_c_613_n 2.21753e-19 $X=2.55 $Y=1.61 $X2=0
+ $Y2=0
cc_393 N_RESET_B_c_430_n N_A_331_392#_c_614_n 0.00526022f $X=2.575 $Y=2.26 $X2=0
+ $Y2=0
cc_394 N_RESET_B_c_431_n N_A_331_392#_c_640_n 0.0128875f $X=2.575 $Y=2.35 $X2=0
+ $Y2=0
cc_395 N_RESET_B_M1025_g N_A_331_392#_c_615_n 0.0348579f $X=2.605 $Y=0.615 $X2=0
+ $Y2=0
cc_396 N_RESET_B_c_413_n N_A_331_392#_c_617_n 0.0032465f $X=1.07 $Y=1.885 $X2=0
+ $Y2=0
cc_397 N_RESET_B_M1009_g N_A_331_392#_c_617_n 0.00141641f $X=1.095 $Y=0.58 $X2=0
+ $Y2=0
cc_398 N_RESET_B_c_420_n N_A_331_392#_c_617_n 0.0232866f $X=2.495 $Y=1.665 $X2=0
+ $Y2=0
cc_399 N_RESET_B_c_421_n N_A_331_392#_c_617_n 0.00266791f $X=1.345 $Y=1.665
+ $X2=0 $Y2=0
cc_400 N_RESET_B_c_425_n N_A_331_392#_c_617_n 0.023733f $X=1.115 $Y=1.615 $X2=0
+ $Y2=0
cc_401 N_RESET_B_M1009_g N_A_331_392#_c_618_n 0.00105701f $X=1.095 $Y=0.58 $X2=0
+ $Y2=0
cc_402 N_RESET_B_c_415_n N_A_331_392#_c_618_n 0.00677421f $X=2.53 $Y=0.18 $X2=0
+ $Y2=0
cc_403 N_RESET_B_M1025_g N_A_331_392#_c_618_n 0.00548205f $X=2.605 $Y=0.615
+ $X2=0 $Y2=0
cc_404 N_RESET_B_c_420_n N_A_331_392#_c_642_n 0.00479833f $X=2.495 $Y=1.665
+ $X2=0 $Y2=0
cc_405 N_RESET_B_M1025_g N_A_331_392#_c_619_n 0.0172211f $X=2.605 $Y=0.615 $X2=0
+ $Y2=0
cc_406 N_RESET_B_c_420_n N_A_331_392#_c_619_n 0.00990898f $X=2.495 $Y=1.665
+ $X2=0 $Y2=0
cc_407 N_RESET_B_c_423_n N_A_331_392#_c_619_n 0.00142776f $X=2.785 $Y=1.665
+ $X2=0 $Y2=0
cc_408 N_RESET_B_c_426_n N_A_331_392#_c_619_n 0.00395315f $X=2.55 $Y=1.61 $X2=0
+ $Y2=0
cc_409 N_RESET_B_c_427_n N_A_331_392#_c_619_n 0.0175537f $X=2.55 $Y=1.61 $X2=0
+ $Y2=0
cc_410 N_RESET_B_M1025_g N_A_331_392#_c_620_n 0.00614625f $X=2.605 $Y=0.615
+ $X2=0 $Y2=0
cc_411 N_RESET_B_M1025_g N_A_331_392#_c_622_n 0.00157742f $X=2.605 $Y=0.615
+ $X2=0 $Y2=0
cc_412 N_RESET_B_M1025_g N_A_331_392#_c_623_n 0.00489643f $X=2.605 $Y=0.615
+ $X2=0 $Y2=0
cc_413 N_RESET_B_c_422_n N_A_331_392#_c_623_n 0.00204418f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_414 N_RESET_B_c_426_n N_A_331_392#_c_623_n 2.34651e-19 $X=2.55 $Y=1.61 $X2=0
+ $Y2=0
cc_415 N_RESET_B_c_427_n N_A_331_392#_c_623_n 0.008544f $X=2.55 $Y=1.61 $X2=0
+ $Y2=0
cc_416 N_RESET_B_c_422_n N_A_331_392#_c_631_n 0.0139858f $X=9.695 $Y=1.665 $X2=0
+ $Y2=0
cc_417 N_RESET_B_c_422_n N_A_331_392#_c_632_n 0.00558182f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_418 N_RESET_B_c_422_n N_A_331_392#_c_633_n 0.0242285f $X=9.695 $Y=1.665 $X2=0
+ $Y2=0
cc_419 N_RESET_B_c_420_n N_A_331_392#_c_634_n 0.00746461f $X=2.495 $Y=1.665
+ $X2=0 $Y2=0
cc_420 N_RESET_B_c_422_n N_A_331_392#_c_635_n 0.00503259f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_421 N_RESET_B_c_423_n N_A_331_392#_c_635_n 0.00118193f $X=2.785 $Y=1.665
+ $X2=0 $Y2=0
cc_422 N_RESET_B_c_422_n N_A_331_392#_c_636_n 0.0217894f $X=9.695 $Y=1.665 $X2=0
+ $Y2=0
cc_423 N_RESET_B_c_423_n N_A_331_392#_c_636_n 0.00230201f $X=2.785 $Y=1.665
+ $X2=0 $Y2=0
cc_424 N_RESET_B_c_426_n N_A_331_392#_c_636_n 3.31881e-19 $X=2.55 $Y=1.61 $X2=0
+ $Y2=0
cc_425 N_RESET_B_c_427_n N_A_331_392#_c_636_n 0.0149803f $X=2.55 $Y=1.61 $X2=0
+ $Y2=0
cc_426 N_RESET_B_c_430_n N_A_331_392#_c_638_n 0.00419637f $X=2.575 $Y=2.26 $X2=0
+ $Y2=0
cc_427 N_RESET_B_c_422_n N_A_331_392#_c_638_n 0.00756058f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_428 N_RESET_B_c_426_n N_A_331_392#_c_638_n 0.0168959f $X=2.55 $Y=1.61 $X2=0
+ $Y2=0
cc_429 N_RESET_B_c_427_n N_A_331_392#_c_638_n 8.2739e-19 $X=2.55 $Y=1.61 $X2=0
+ $Y2=0
cc_430 N_RESET_B_c_422_n N_A_818_418#_c_840_n 0.00175829f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_431 N_RESET_B_c_422_n N_A_818_418#_M1035_g 0.00702513f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_432 N_RESET_B_c_422_n N_A_818_418#_c_843_n 0.00253849f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_433 N_RESET_B_c_422_n N_A_818_418#_c_844_n 0.0108262f $X=9.695 $Y=1.665 $X2=0
+ $Y2=0
cc_434 N_RESET_B_c_422_n N_A_818_418#_c_845_n 0.00323944f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_435 N_RESET_B_c_422_n N_A_818_418#_c_846_n 0.0319081f $X=9.695 $Y=1.665 $X2=0
+ $Y2=0
cc_436 N_RESET_B_c_422_n N_A_818_418#_c_847_n 0.0156071f $X=9.695 $Y=1.665 $X2=0
+ $Y2=0
cc_437 N_RESET_B_c_422_n N_A_818_418#_c_848_n 0.015652f $X=9.695 $Y=1.665 $X2=0
+ $Y2=0
cc_438 N_RESET_B_c_422_n N_A_818_418#_c_850_n 0.0164157f $X=9.695 $Y=1.665 $X2=0
+ $Y2=0
cc_439 N_RESET_B_c_422_n N_A_818_418#_c_851_n 0.0142935f $X=9.695 $Y=1.665 $X2=0
+ $Y2=0
cc_440 N_RESET_B_c_422_n N_A_818_418#_c_852_n 0.0052628f $X=9.695 $Y=1.665 $X2=0
+ $Y2=0
cc_441 N_RESET_B_c_422_n N_A_728_331#_M1004_g 0.00214871f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_442 N_RESET_B_c_422_n N_A_728_331#_c_1012_n 0.00996207f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_443 N_RESET_B_c_422_n N_A_728_331#_M1013_g 0.00279101f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_444 N_RESET_B_c_422_n N_A_728_331#_c_1004_n 0.00419627f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_445 N_RESET_B_c_422_n N_A_728_331#_c_1015_n 0.00829884f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_446 N_RESET_B_c_422_n N_A_728_331#_c_1016_n 0.0132491f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_447 N_RESET_B_c_422_n N_A_728_331#_c_1005_n 6.34002e-19 $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_448 N_RESET_B_c_422_n N_A_728_331#_c_1038_n 0.033043f $X=9.695 $Y=1.665 $X2=0
+ $Y2=0
cc_449 N_RESET_B_c_422_n N_A_728_331#_c_1006_n 0.0200477f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_450 N_RESET_B_c_422_n N_A_728_331#_c_1040_n 0.0405177f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_451 N_RESET_B_c_422_n N_A_728_331#_c_1008_n 0.019344f $X=9.695 $Y=1.665 $X2=0
+ $Y2=0
cc_452 N_RESET_B_c_422_n N_A_728_331#_c_1021_n 0.00622674f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_453 N_RESET_B_c_422_n N_CLK_c_1168_n 0.0122642f $X=9.695 $Y=1.665 $X2=0 $Y2=0
cc_454 N_RESET_B_c_422_n CLK 0.023017f $X=9.695 $Y=1.665 $X2=0 $Y2=0
cc_455 N_RESET_B_c_418_n N_A_1800_291#_c_1206_n 0.0350315f $X=9.77 $Y=1.87 $X2=0
+ $Y2=0
cc_456 N_RESET_B_c_422_n N_A_1800_291#_c_1206_n 0.00447808f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_457 N_RESET_B_c_428_n N_A_1800_291#_c_1206_n 0.00111757f $X=9.705 $Y=1.615
+ $X2=0 $Y2=0
cc_458 N_RESET_B_c_418_n N_A_1800_291#_c_1207_n 2.59732e-19 $X=9.77 $Y=1.87
+ $X2=0 $Y2=0
cc_459 N_RESET_B_M1019_g N_A_1800_291#_c_1207_n 0.0129042f $X=9.795 $Y=0.58
+ $X2=0 $Y2=0
cc_460 N_RESET_B_M1019_g N_A_1800_291#_c_1208_n 0.0189671f $X=9.795 $Y=0.58
+ $X2=0 $Y2=0
cc_461 N_RESET_B_c_418_n N_A_1800_291#_c_1210_n 0.00375536f $X=9.77 $Y=1.87
+ $X2=0 $Y2=0
cc_462 N_RESET_B_c_422_n N_A_1800_291#_c_1210_n 0.0212822f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_463 N_RESET_B_c_424_n N_A_1800_291#_c_1210_n 4.42853e-19 $X=9.84 $Y=1.665
+ $X2=0 $Y2=0
cc_464 N_RESET_B_c_428_n N_A_1800_291#_c_1210_n 0.0185283f $X=9.705 $Y=1.615
+ $X2=0 $Y2=0
cc_465 N_RESET_B_M1019_g N_A_1800_291#_c_1211_n 6.13047e-19 $X=9.795 $Y=0.58
+ $X2=0 $Y2=0
cc_466 N_RESET_B_c_424_n N_A_1800_291#_c_1211_n 0.0057125f $X=9.84 $Y=1.665
+ $X2=0 $Y2=0
cc_467 N_RESET_B_c_428_n N_A_1800_291#_c_1211_n 0.00751959f $X=9.705 $Y=1.615
+ $X2=0 $Y2=0
cc_468 N_RESET_B_c_418_n N_A_1800_291#_c_1230_n 0.0153425f $X=9.77 $Y=1.87 $X2=0
+ $Y2=0
cc_469 N_RESET_B_c_422_n N_A_1800_291#_c_1230_n 0.0101591f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_470 N_RESET_B_c_424_n N_A_1800_291#_c_1230_n 0.00804814f $X=9.84 $Y=1.665
+ $X2=0 $Y2=0
cc_471 N_RESET_B_c_428_n N_A_1800_291#_c_1230_n 0.023488f $X=9.705 $Y=1.615
+ $X2=0 $Y2=0
cc_472 N_RESET_B_c_418_n N_A_1800_291#_c_1216_n 0.00615353f $X=9.77 $Y=1.87
+ $X2=0 $Y2=0
cc_473 N_RESET_B_M1019_g N_A_1800_291#_c_1212_n 0.00122306f $X=9.795 $Y=0.58
+ $X2=0 $Y2=0
cc_474 N_RESET_B_M1019_g N_A_1586_149#_M1017_g 0.0677574f $X=9.795 $Y=0.58 $X2=0
+ $Y2=0
cc_475 N_RESET_B_c_418_n N_A_1586_149#_c_1294_n 0.0112224f $X=9.77 $Y=1.87 $X2=0
+ $Y2=0
cc_476 N_RESET_B_c_418_n N_A_1586_149#_c_1303_n 0.0142317f $X=9.77 $Y=1.87 $X2=0
+ $Y2=0
cc_477 N_RESET_B_c_422_n N_A_1586_149#_c_1314_n 0.0116802f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_478 N_RESET_B_c_422_n N_A_1586_149#_c_1298_n 0.0176982f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_479 N_RESET_B_c_418_n N_A_1586_149#_c_1299_n 0.00417884f $X=9.77 $Y=1.87
+ $X2=0 $Y2=0
cc_480 N_RESET_B_M1019_g N_A_1586_149#_c_1299_n 0.0209819f $X=9.795 $Y=0.58
+ $X2=0 $Y2=0
cc_481 N_RESET_B_c_422_n N_A_1586_149#_c_1299_n 0.017962f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_482 N_RESET_B_c_424_n N_A_1586_149#_c_1299_n 0.00291677f $X=9.84 $Y=1.665
+ $X2=0 $Y2=0
cc_483 N_RESET_B_c_428_n N_A_1586_149#_c_1299_n 0.0280535f $X=9.705 $Y=1.615
+ $X2=0 $Y2=0
cc_484 N_RESET_B_c_422_n N_A_1586_149#_c_1309_n 0.0120089f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_485 N_RESET_B_M1019_g N_A_1586_149#_c_1301_n 0.0112224f $X=9.795 $Y=0.58
+ $X2=0 $Y2=0
cc_486 N_RESET_B_c_424_n N_A_1586_149#_c_1301_n 0.00422176f $X=9.84 $Y=1.665
+ $X2=0 $Y2=0
cc_487 N_RESET_B_c_428_n N_A_1586_149#_c_1301_n 0.00318809f $X=9.705 $Y=1.615
+ $X2=0 $Y2=0
cc_488 N_RESET_B_c_431_n N_VPWR_c_1494_n 0.00109138f $X=2.575 $Y=2.35 $X2=0
+ $Y2=0
cc_489 N_RESET_B_c_418_n N_VPWR_c_1496_n 0.00427005f $X=9.77 $Y=1.87 $X2=0 $Y2=0
cc_490 N_RESET_B_c_422_n N_VPWR_c_1496_n 2.54661e-19 $X=9.695 $Y=1.665 $X2=0
+ $Y2=0
cc_491 N_RESET_B_c_413_n N_VPWR_c_1503_n 2.93609e-19 $X=1.07 $Y=1.885 $X2=0
+ $Y2=0
cc_492 N_RESET_B_c_431_n N_VPWR_c_1507_n 7.53214e-19 $X=2.575 $Y=2.35 $X2=0
+ $Y2=0
cc_493 N_RESET_B_c_418_n N_VPWR_c_1491_n 0.00384901f $X=9.77 $Y=1.87 $X2=0 $Y2=0
cc_494 N_RESET_B_M1009_g N_A_70_74#_c_1639_n 0.001902f $X=1.095 $Y=0.58 $X2=0
+ $Y2=0
cc_495 N_RESET_B_c_413_n N_A_70_74#_c_1644_n 0.00582696f $X=1.07 $Y=1.885 $X2=0
+ $Y2=0
cc_496 N_RESET_B_c_413_n N_A_70_74#_c_1645_n 0.00852752f $X=1.07 $Y=1.885 $X2=0
+ $Y2=0
cc_497 N_RESET_B_c_413_n N_A_70_74#_c_1646_n 0.00592963f $X=1.07 $Y=1.885 $X2=0
+ $Y2=0
cc_498 N_RESET_B_c_431_n N_A_70_74#_c_1648_n 0.0109422f $X=2.575 $Y=2.35 $X2=0
+ $Y2=0
cc_499 N_RESET_B_c_431_n N_A_70_74#_c_1649_n 0.0160525f $X=2.575 $Y=2.35 $X2=0
+ $Y2=0
cc_500 N_RESET_B_c_431_n N_A_70_74#_c_1651_n 0.00667273f $X=2.575 $Y=2.35 $X2=0
+ $Y2=0
cc_501 N_RESET_B_c_422_n N_A_70_74#_c_1640_n 0.0107306f $X=9.695 $Y=1.665 $X2=0
+ $Y2=0
cc_502 N_RESET_B_c_422_n N_A_70_74#_c_1641_n 0.0218579f $X=9.695 $Y=1.665 $X2=0
+ $Y2=0
cc_503 N_RESET_B_c_413_n N_A_70_74#_c_1642_n 0.00404604f $X=1.07 $Y=1.885 $X2=0
+ $Y2=0
cc_504 N_RESET_B_M1009_g N_A_70_74#_c_1642_n 0.00983764f $X=1.095 $Y=0.58 $X2=0
+ $Y2=0
cc_505 N_RESET_B_c_421_n N_A_70_74#_c_1642_n 0.00155586f $X=1.345 $Y=1.665 $X2=0
+ $Y2=0
cc_506 N_RESET_B_c_425_n N_A_70_74#_c_1642_n 0.0230072f $X=1.115 $Y=1.615 $X2=0
+ $Y2=0
cc_507 N_RESET_B_c_422_n N_A_70_74#_c_1643_n 0.0110159f $X=9.695 $Y=1.665 $X2=0
+ $Y2=0
cc_508 N_RESET_B_c_413_n N_VGND_c_1851_n 0.0018485f $X=1.07 $Y=1.885 $X2=0 $Y2=0
cc_509 N_RESET_B_M1009_g N_VGND_c_1851_n 0.0125926f $X=1.095 $Y=0.58 $X2=0 $Y2=0
cc_510 N_RESET_B_c_415_n N_VGND_c_1851_n 0.0185344f $X=2.53 $Y=0.18 $X2=0 $Y2=0
cc_511 N_RESET_B_c_416_n N_VGND_c_1851_n 0.00363087f $X=1.17 $Y=0.18 $X2=0 $Y2=0
cc_512 N_RESET_B_c_425_n N_VGND_c_1851_n 0.00512544f $X=1.115 $Y=1.615 $X2=0
+ $Y2=0
cc_513 N_RESET_B_c_415_n N_VGND_c_1852_n 0.0228038f $X=2.53 $Y=0.18 $X2=0 $Y2=0
cc_514 N_RESET_B_M1025_g N_VGND_c_1852_n 0.00790765f $X=2.605 $Y=0.615 $X2=0
+ $Y2=0
cc_515 N_RESET_B_M1019_g N_VGND_c_1854_n 0.0101946f $X=9.795 $Y=0.58 $X2=0 $Y2=0
cc_516 N_RESET_B_c_415_n N_VGND_c_1860_n 0.0216293f $X=2.53 $Y=0.18 $X2=0 $Y2=0
cc_517 N_RESET_B_c_415_n N_VGND_c_1862_n 0.00564095f $X=2.53 $Y=0.18 $X2=0 $Y2=0
cc_518 N_RESET_B_M1019_g N_VGND_c_1866_n 0.00383152f $X=9.795 $Y=0.58 $X2=0
+ $Y2=0
cc_519 N_RESET_B_c_416_n N_VGND_c_1868_n 0.00486043f $X=1.17 $Y=0.18 $X2=0 $Y2=0
cc_520 N_RESET_B_c_415_n N_VGND_c_1875_n 0.0378561f $X=2.53 $Y=0.18 $X2=0 $Y2=0
cc_521 N_RESET_B_c_416_n N_VGND_c_1875_n 0.00977974f $X=1.17 $Y=0.18 $X2=0 $Y2=0
cc_522 N_RESET_B_M1019_g N_VGND_c_1875_n 0.0075694f $X=9.795 $Y=0.58 $X2=0 $Y2=0
cc_523 N_RESET_B_c_422_n N_A_614_81#_c_2001_n 0.0159116f $X=9.695 $Y=1.665 $X2=0
+ $Y2=0
cc_524 N_RESET_B_c_422_n N_A_1499_149#_c_2024_n 4.58014e-19 $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_525 N_A_331_392#_c_624_n N_A_818_418#_M1030_s 0.00227252f $X=5.15 $Y=0.66
+ $X2=-0.19 $Y2=-0.245
cc_526 N_A_331_392#_c_711_p N_A_818_418#_M1030_s 0.0027085f $X=6.025 $Y=0.745
+ $X2=-0.19 $Y2=-0.245
cc_527 N_A_331_392#_c_625_n N_A_818_418#_M1030_s 0.00199188f $X=5.235 $Y=0.745
+ $X2=-0.19 $Y2=-0.245
cc_528 N_A_331_392#_c_630_n N_A_818_418#_c_842_n 0.0119277f $X=8.615 $Y=0.34
+ $X2=0 $Y2=0
cc_529 N_A_331_392#_c_711_p N_A_818_418#_c_846_n 0.0105363f $X=6.025 $Y=0.745
+ $X2=0 $Y2=0
cc_530 N_A_331_392#_c_625_n N_A_818_418#_c_846_n 0.0124528f $X=5.235 $Y=0.745
+ $X2=0 $Y2=0
cc_531 N_A_331_392#_c_633_n N_A_818_418#_c_859_n 0.0123434f $X=7.795 $Y=2.09
+ $X2=0 $Y2=0
cc_532 N_A_331_392#_c_633_n N_A_818_418#_c_860_n 0.00909366f $X=7.795 $Y=2.09
+ $X2=0 $Y2=0
cc_533 N_A_331_392#_M1028_s N_A_818_418#_c_861_n 0.00410029f $X=7.665 $Y=1.945
+ $X2=0 $Y2=0
cc_534 N_A_331_392#_c_633_n N_A_818_418#_c_861_n 0.012787f $X=7.795 $Y=2.09
+ $X2=0 $Y2=0
cc_535 N_A_331_392#_c_633_n N_A_818_418#_c_847_n 0.0787051f $X=7.795 $Y=2.09
+ $X2=0 $Y2=0
cc_536 N_A_331_392#_c_629_n N_A_818_418#_c_851_n 0.0024581f $X=7.3 $Y=1.355
+ $X2=0 $Y2=0
cc_537 N_A_331_392#_c_631_n N_A_818_418#_c_851_n 0.0147826f $X=7.71 $Y=1.44
+ $X2=0 $Y2=0
cc_538 N_A_331_392#_c_633_n N_A_818_418#_c_851_n 0.00609504f $X=7.795 $Y=2.09
+ $X2=0 $Y2=0
cc_539 N_A_331_392#_c_614_n N_A_728_331#_c_998_n 0.0150517f $X=3.34 $Y=2.26
+ $X2=0 $Y2=0
cc_540 N_A_331_392#_c_640_n N_A_728_331#_c_1010_n 0.0461694f $X=3.34 $Y=2.35
+ $X2=0 $Y2=0
cc_541 N_A_331_392#_c_616_n N_A_728_331#_M1004_g 0.007711f $X=3.012 $Y=1.05
+ $X2=0 $Y2=0
cc_542 N_A_331_392#_c_621_n N_A_728_331#_M1004_g 0.00252325f $X=5.065 $Y=0.34
+ $X2=0 $Y2=0
cc_543 N_A_331_392#_c_623_n N_A_728_331#_M1004_g 7.95442e-19 $X=3.01 $Y=1.555
+ $X2=0 $Y2=0
cc_544 N_A_331_392#_c_636_n N_A_728_331#_M1004_g 2.86655e-19 $X=3.09 $Y=1.68
+ $X2=0 $Y2=0
cc_545 N_A_331_392#_c_638_n N_A_728_331#_M1004_g 0.00556159f $X=3.34 $Y=1.68
+ $X2=0 $Y2=0
cc_546 N_A_331_392#_c_621_n N_A_728_331#_c_1000_n 0.0575563f $X=5.065 $Y=0.34
+ $X2=0 $Y2=0
cc_547 N_A_331_392#_c_711_p N_A_728_331#_c_1000_n 0.00157743f $X=6.025 $Y=0.745
+ $X2=0 $Y2=0
cc_548 N_A_331_392#_c_615_n N_A_728_331#_c_1001_n 0.00720262f $X=3.012 $Y=0.9
+ $X2=0 $Y2=0
cc_549 N_A_331_392#_c_621_n N_A_728_331#_c_1001_n 0.0074164f $X=5.065 $Y=0.34
+ $X2=0 $Y2=0
cc_550 N_A_331_392#_c_621_n N_A_728_331#_M1030_g 2.14932e-19 $X=5.065 $Y=0.34
+ $X2=0 $Y2=0
cc_551 N_A_331_392#_c_624_n N_A_728_331#_M1030_g 0.00722282f $X=5.15 $Y=0.66
+ $X2=0 $Y2=0
cc_552 N_A_331_392#_c_711_p N_A_728_331#_M1030_g 0.0190035f $X=6.025 $Y=0.745
+ $X2=0 $Y2=0
cc_553 N_A_331_392#_c_626_n N_A_728_331#_M1030_g 0.00429098f $X=6.11 $Y=0.66
+ $X2=0 $Y2=0
cc_554 N_A_331_392#_c_633_n N_A_728_331#_c_1012_n 0.00926793f $X=7.795 $Y=2.09
+ $X2=0 $Y2=0
cc_555 N_A_331_392#_c_629_n N_A_728_331#_M1013_g 0.00510454f $X=7.3 $Y=1.355
+ $X2=0 $Y2=0
cc_556 N_A_331_392#_c_630_n N_A_728_331#_M1013_g 9.86678e-19 $X=8.615 $Y=0.34
+ $X2=0 $Y2=0
cc_557 N_A_331_392#_c_631_n N_A_728_331#_M1013_g 0.00939999f $X=7.71 $Y=1.44
+ $X2=0 $Y2=0
cc_558 N_A_331_392#_c_633_n N_A_728_331#_M1013_g 0.00547121f $X=7.795 $Y=2.09
+ $X2=0 $Y2=0
cc_559 N_A_331_392#_c_633_n N_A_728_331#_c_1014_n 0.0045069f $X=7.795 $Y=2.09
+ $X2=0 $Y2=0
cc_560 N_A_331_392#_c_636_n N_A_728_331#_c_1004_n 3.90209e-19 $X=3.09 $Y=1.68
+ $X2=0 $Y2=0
cc_561 N_A_331_392#_c_638_n N_A_728_331#_c_1004_n 0.0150517f $X=3.34 $Y=1.68
+ $X2=0 $Y2=0
cc_562 N_A_331_392#_c_633_n N_A_728_331#_c_1015_n 0.00524491f $X=7.795 $Y=2.09
+ $X2=0 $Y2=0
cc_563 N_A_331_392#_c_631_n N_A_728_331#_c_1017_n 0.00320602f $X=7.71 $Y=1.44
+ $X2=0 $Y2=0
cc_564 N_A_331_392#_c_632_n N_A_728_331#_c_1017_n 0.00513005f $X=7.385 $Y=1.44
+ $X2=0 $Y2=0
cc_565 N_A_331_392#_c_633_n N_A_728_331#_c_1017_n 0.0223244f $X=7.795 $Y=2.09
+ $X2=0 $Y2=0
cc_566 N_A_331_392#_c_711_p N_A_728_331#_c_1038_n 0.0191238f $X=6.025 $Y=0.745
+ $X2=0 $Y2=0
cc_567 N_A_331_392#_c_711_p N_A_728_331#_c_1007_n 0.0151771f $X=6.025 $Y=0.745
+ $X2=0 $Y2=0
cc_568 N_A_331_392#_c_626_n N_A_728_331#_c_1007_n 0.001895f $X=6.11 $Y=0.66
+ $X2=0 $Y2=0
cc_569 N_A_331_392#_c_627_n N_A_728_331#_c_1007_n 0.0322868f $X=7.215 $Y=0.34
+ $X2=0 $Y2=0
cc_570 N_A_331_392#_c_629_n N_A_728_331#_c_1007_n 0.0206296f $X=7.3 $Y=1.355
+ $X2=0 $Y2=0
cc_571 N_A_331_392#_c_633_n N_A_728_331#_c_1019_n 0.00241743f $X=7.795 $Y=2.09
+ $X2=0 $Y2=0
cc_572 N_A_331_392#_c_711_p N_A_728_331#_c_1008_n 0.0116042f $X=6.025 $Y=0.745
+ $X2=0 $Y2=0
cc_573 N_A_331_392#_c_631_n N_A_728_331#_c_1021_n 0.00851598f $X=7.71 $Y=1.44
+ $X2=0 $Y2=0
cc_574 N_A_331_392#_c_632_n N_A_728_331#_c_1021_n 0.00337292f $X=7.385 $Y=1.44
+ $X2=0 $Y2=0
cc_575 N_A_331_392#_c_633_n N_A_728_331#_c_1021_n 0.00109399f $X=7.795 $Y=2.09
+ $X2=0 $Y2=0
cc_576 N_A_331_392#_c_711_p N_CLK_c_1167_n 9.69516e-19 $X=6.025 $Y=0.745
+ $X2=-0.19 $Y2=-0.245
cc_577 N_A_331_392#_c_626_n N_CLK_c_1167_n 0.0063257f $X=6.11 $Y=0.66 $X2=-0.19
+ $Y2=-0.245
cc_578 N_A_331_392#_c_627_n N_CLK_c_1167_n 0.00861985f $X=7.215 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_579 N_A_331_392#_c_629_n N_CLK_c_1167_n 0.0091992f $X=7.3 $Y=1.355 $X2=-0.19
+ $Y2=-0.245
cc_580 N_A_331_392#_c_632_n N_CLK_c_1168_n 0.00108413f $X=7.385 $Y=1.44 $X2=0
+ $Y2=0
cc_581 N_A_331_392#_c_629_n CLK 0.0138701f $X=7.3 $Y=1.355 $X2=0 $Y2=0
cc_582 N_A_331_392#_c_632_n CLK 0.0150422f $X=7.385 $Y=1.44 $X2=0 $Y2=0
cc_583 N_A_331_392#_c_633_n CLK 0.00323555f $X=7.795 $Y=2.09 $X2=0 $Y2=0
cc_584 N_A_331_392#_c_630_n N_A_1800_291#_c_1208_n 0.00175601f $X=8.615 $Y=0.34
+ $X2=0 $Y2=0
cc_585 N_A_331_392#_M1021_d N_A_1586_149#_c_1314_n 0.00571341f $X=8.405 $Y=0.425
+ $X2=0 $Y2=0
cc_586 N_A_331_392#_M1021_d N_A_1586_149#_c_1300_n 0.0013268f $X=8.405 $Y=0.425
+ $X2=0 $Y2=0
cc_587 N_A_331_392#_c_640_n N_VPWR_c_1494_n 0.00376512f $X=3.34 $Y=2.35 $X2=0
+ $Y2=0
cc_588 N_A_331_392#_c_640_n N_VPWR_c_1495_n 0.00355997f $X=3.34 $Y=2.35 $X2=0
+ $Y2=0
cc_589 N_A_331_392#_c_640_n N_VPWR_c_1491_n 0.00339925f $X=3.34 $Y=2.35 $X2=0
+ $Y2=0
cc_590 N_A_331_392#_c_617_n N_A_70_74#_c_1644_n 0.00560278f $X=1.57 $Y=2.285
+ $X2=0 $Y2=0
cc_591 N_A_331_392#_c_657_n N_A_70_74#_c_1646_n 0.00761753f $X=1.655 $Y=2.37
+ $X2=0 $Y2=0
cc_592 N_A_331_392#_M1031_d N_A_70_74#_c_1648_n 0.00346067f $X=1.655 $Y=1.96
+ $X2=0 $Y2=0
cc_593 N_A_331_392#_c_642_n N_A_70_74#_c_1648_n 0.00696584f $X=1.805 $Y=2.37
+ $X2=0 $Y2=0
cc_594 N_A_331_392#_c_640_n N_A_70_74#_c_1649_n 0.00159671f $X=3.34 $Y=2.35
+ $X2=0 $Y2=0
cc_595 N_A_331_392#_c_640_n N_A_70_74#_c_1650_n 0.0139194f $X=3.34 $Y=2.35 $X2=0
+ $Y2=0
cc_596 N_A_331_392#_c_640_n N_A_70_74#_c_1652_n 0.0098205f $X=3.34 $Y=2.35 $X2=0
+ $Y2=0
cc_597 N_A_331_392#_c_640_n N_A_70_74#_c_1654_n 0.00239859f $X=3.34 $Y=2.35
+ $X2=0 $Y2=0
cc_598 N_A_331_392#_c_617_n N_A_70_74#_c_1642_n 0.0107766f $X=1.57 $Y=2.285
+ $X2=0 $Y2=0
cc_599 N_A_331_392#_M1031_d N_A_70_74#_c_1659_n 0.00915137f $X=1.655 $Y=1.96
+ $X2=0 $Y2=0
cc_600 N_A_331_392#_c_657_n N_A_70_74#_c_1659_n 0.00393953f $X=1.655 $Y=2.37
+ $X2=0 $Y2=0
cc_601 N_A_331_392#_c_642_n N_A_70_74#_c_1659_n 0.00487896f $X=1.805 $Y=2.37
+ $X2=0 $Y2=0
cc_602 N_A_331_392#_c_616_n N_A_70_74#_c_1643_n 0.00441246f $X=3.012 $Y=1.05
+ $X2=0 $Y2=0
cc_603 N_A_331_392#_c_620_n N_A_70_74#_c_1643_n 0.00314822f $X=2.79 $Y=1.015
+ $X2=0 $Y2=0
cc_604 N_A_331_392#_c_623_n N_A_70_74#_c_1643_n 0.0114522f $X=3.01 $Y=1.555
+ $X2=0 $Y2=0
cc_605 N_A_331_392#_c_635_n N_A_70_74#_c_1643_n 0.0106126f $X=3.01 $Y=1.1 $X2=0
+ $Y2=0
cc_606 N_A_331_392#_c_638_n N_A_70_74#_c_1643_n 0.00282478f $X=3.34 $Y=1.68
+ $X2=0 $Y2=0
cc_607 N_A_331_392#_c_711_p N_VGND_M1030_d 0.0205914f $X=6.025 $Y=0.745 $X2=0
+ $Y2=0
cc_608 N_A_331_392#_c_626_n N_VGND_M1030_d 0.00621489f $X=6.11 $Y=0.66 $X2=0
+ $Y2=0
cc_609 N_A_331_392#_c_618_n N_VGND_c_1851_n 0.0183123f $X=1.81 $Y=0.76 $X2=0
+ $Y2=0
cc_610 N_A_331_392#_c_615_n N_VGND_c_1852_n 2.1461e-19 $X=3.012 $Y=0.9 $X2=0
+ $Y2=0
cc_611 N_A_331_392#_c_618_n N_VGND_c_1852_n 0.0212369f $X=1.81 $Y=0.76 $X2=0
+ $Y2=0
cc_612 N_A_331_392#_c_619_n N_VGND_c_1852_n 0.0194224f $X=2.705 $Y=1.1 $X2=0
+ $Y2=0
cc_613 N_A_331_392#_c_622_n N_VGND_c_1852_n 0.0133176f $X=2.875 $Y=0.34 $X2=0
+ $Y2=0
cc_614 N_A_331_392#_c_621_n N_VGND_c_1853_n 0.00787195f $X=5.065 $Y=0.34 $X2=0
+ $Y2=0
cc_615 N_A_331_392#_c_624_n N_VGND_c_1853_n 0.00291186f $X=5.15 $Y=0.66 $X2=0
+ $Y2=0
cc_616 N_A_331_392#_c_711_p N_VGND_c_1853_n 0.0190193f $X=6.025 $Y=0.745 $X2=0
+ $Y2=0
cc_617 N_A_331_392#_c_626_n N_VGND_c_1853_n 0.00491053f $X=6.11 $Y=0.66 $X2=0
+ $Y2=0
cc_618 N_A_331_392#_c_628_n N_VGND_c_1853_n 0.0145006f $X=6.195 $Y=0.34 $X2=0
+ $Y2=0
cc_619 N_A_331_392#_c_630_n N_VGND_c_1854_n 0.00292246f $X=8.615 $Y=0.34 $X2=0
+ $Y2=0
cc_620 N_A_331_392#_c_618_n N_VGND_c_1860_n 0.00993789f $X=1.81 $Y=0.76 $X2=0
+ $Y2=0
cc_621 N_A_331_392#_c_615_n N_VGND_c_1862_n 9.15902e-19 $X=3.012 $Y=0.9 $X2=0
+ $Y2=0
cc_622 N_A_331_392#_c_621_n N_VGND_c_1862_n 0.153051f $X=5.065 $Y=0.34 $X2=0
+ $Y2=0
cc_623 N_A_331_392#_c_622_n N_VGND_c_1862_n 0.0121867f $X=2.875 $Y=0.34 $X2=0
+ $Y2=0
cc_624 N_A_331_392#_c_711_p N_VGND_c_1862_n 0.0051071f $X=6.025 $Y=0.745 $X2=0
+ $Y2=0
cc_625 N_A_331_392#_c_711_p N_VGND_c_1864_n 0.00279509f $X=6.025 $Y=0.745 $X2=0
+ $Y2=0
cc_626 N_A_331_392#_c_627_n N_VGND_c_1864_n 0.0656484f $X=7.215 $Y=0.34 $X2=0
+ $Y2=0
cc_627 N_A_331_392#_c_628_n N_VGND_c_1864_n 0.0120335f $X=6.195 $Y=0.34 $X2=0
+ $Y2=0
cc_628 N_A_331_392#_c_630_n N_VGND_c_1864_n 0.0895608f $X=8.615 $Y=0.34 $X2=0
+ $Y2=0
cc_629 N_A_331_392#_c_637_n N_VGND_c_1864_n 0.0121867f $X=7.3 $Y=0.34 $X2=0
+ $Y2=0
cc_630 N_A_331_392#_M1021_d N_VGND_c_1875_n 0.00257669f $X=8.405 $Y=0.425 $X2=0
+ $Y2=0
cc_631 N_A_331_392#_c_618_n N_VGND_c_1875_n 0.00993216f $X=1.81 $Y=0.76 $X2=0
+ $Y2=0
cc_632 N_A_331_392#_c_621_n N_VGND_c_1875_n 0.0889116f $X=5.065 $Y=0.34 $X2=0
+ $Y2=0
cc_633 N_A_331_392#_c_622_n N_VGND_c_1875_n 0.00660921f $X=2.875 $Y=0.34 $X2=0
+ $Y2=0
cc_634 N_A_331_392#_c_711_p N_VGND_c_1875_n 0.0161016f $X=6.025 $Y=0.745 $X2=0
+ $Y2=0
cc_635 N_A_331_392#_c_627_n N_VGND_c_1875_n 0.0383417f $X=7.215 $Y=0.34 $X2=0
+ $Y2=0
cc_636 N_A_331_392#_c_628_n N_VGND_c_1875_n 0.00658039f $X=6.195 $Y=0.34 $X2=0
+ $Y2=0
cc_637 N_A_331_392#_c_630_n N_VGND_c_1875_n 0.052445f $X=8.615 $Y=0.34 $X2=0
+ $Y2=0
cc_638 N_A_331_392#_c_637_n N_VGND_c_1875_n 0.00660921f $X=7.3 $Y=0.34 $X2=0
+ $Y2=0
cc_639 N_A_331_392#_c_620_n A_536_81# 0.00157084f $X=2.79 $Y=1.015 $X2=-0.19
+ $Y2=-0.245
cc_640 N_A_331_392#_c_621_n N_A_614_81#_M1011_d 0.00277417f $X=5.065 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_641 N_A_331_392#_c_615_n N_A_614_81#_c_2000_n 0.00242033f $X=3.012 $Y=0.9
+ $X2=0 $Y2=0
cc_642 N_A_331_392#_c_621_n N_A_614_81#_c_2000_n 0.127151f $X=5.065 $Y=0.34
+ $X2=0 $Y2=0
cc_643 N_A_331_392#_c_624_n N_A_614_81#_c_2000_n 0.00545207f $X=5.15 $Y=0.66
+ $X2=0 $Y2=0
cc_644 N_A_331_392#_c_625_n N_A_614_81#_c_2000_n 0.00983818f $X=5.235 $Y=0.745
+ $X2=0 $Y2=0
cc_645 N_A_331_392#_c_635_n N_A_614_81#_c_2000_n 0.00184287f $X=3.01 $Y=1.1
+ $X2=0 $Y2=0
cc_646 N_A_331_392#_c_625_n N_A_614_81#_c_2001_n 0.00559801f $X=5.235 $Y=0.745
+ $X2=0 $Y2=0
cc_647 N_A_331_392#_c_629_n N_A_1499_149#_c_2024_n 0.0310557f $X=7.3 $Y=1.355
+ $X2=0 $Y2=0
cc_648 N_A_331_392#_c_631_n N_A_1499_149#_c_2024_n 0.0133791f $X=7.71 $Y=1.44
+ $X2=0 $Y2=0
cc_649 N_A_331_392#_M1021_d N_A_1499_149#_c_2025_n 0.00704081f $X=8.405 $Y=0.425
+ $X2=0 $Y2=0
cc_650 N_A_331_392#_c_630_n N_A_1499_149#_c_2025_n 0.0689604f $X=8.615 $Y=0.34
+ $X2=0 $Y2=0
cc_651 N_A_331_392#_c_631_n N_A_1499_149#_c_2025_n 0.00378293f $X=7.71 $Y=1.44
+ $X2=0 $Y2=0
cc_652 N_A_331_392#_c_629_n N_A_1499_149#_c_2026_n 0.0143225f $X=7.3 $Y=1.355
+ $X2=0 $Y2=0
cc_653 N_A_331_392#_c_630_n N_A_1499_149#_c_2026_n 0.0132852f $X=8.615 $Y=0.34
+ $X2=0 $Y2=0
cc_654 N_A_331_392#_c_630_n N_A_1499_149#_c_2027_n 0.00562463f $X=8.615 $Y=0.34
+ $X2=0 $Y2=0
cc_655 N_A_818_418#_c_859_n N_A_728_331#_M1007_d 0.00821329f $X=7.315 $Y=2.51
+ $X2=0 $Y2=0
cc_656 N_A_818_418#_c_840_n N_A_728_331#_c_998_n 0.012312f $X=4.18 $Y=2.35 $X2=0
+ $Y2=0
cc_657 N_A_818_418#_M1035_g N_A_728_331#_c_998_n 0.00720264f $X=4.265 $Y=1.37
+ $X2=0 $Y2=0
cc_658 N_A_818_418#_c_840_n N_A_728_331#_c_1010_n 0.0114096f $X=4.18 $Y=2.35
+ $X2=0 $Y2=0
cc_659 N_A_818_418#_M1035_g N_A_728_331#_M1004_g 0.0191869f $X=4.265 $Y=1.37
+ $X2=0 $Y2=0
cc_660 N_A_818_418#_M1035_g N_A_728_331#_c_1000_n 0.00194711f $X=4.265 $Y=1.37
+ $X2=0 $Y2=0
cc_661 N_A_818_418#_c_846_n N_A_728_331#_c_1000_n 4.78794e-19 $X=5.26 $Y=1.085
+ $X2=0 $Y2=0
cc_662 N_A_818_418#_c_846_n N_A_728_331#_M1030_g 0.0172164f $X=5.26 $Y=1.085
+ $X2=0 $Y2=0
cc_663 N_A_818_418#_c_846_n N_A_728_331#_c_1011_n 0.00148066f $X=5.26 $Y=1.085
+ $X2=0 $Y2=0
cc_664 N_A_818_418#_c_857_n N_A_728_331#_c_1011_n 0.0079437f $X=5.605 $Y=2.425
+ $X2=0 $Y2=0
cc_665 N_A_818_418#_c_858_n N_A_728_331#_c_1011_n 0.0104438f $X=5.62 $Y=2.815
+ $X2=0 $Y2=0
cc_666 N_A_818_418#_c_859_n N_A_728_331#_c_1011_n 0.0147078f $X=7.315 $Y=2.51
+ $X2=0 $Y2=0
cc_667 N_A_818_418#_c_849_n N_A_728_331#_c_1011_n 0.00396352f $X=5.15 $Y=2.075
+ $X2=0 $Y2=0
cc_668 N_A_818_418#_c_850_n N_A_728_331#_c_1011_n 0.00815181f $X=5.62 $Y=2.005
+ $X2=0 $Y2=0
cc_669 N_A_818_418#_c_866_n N_A_728_331#_c_1011_n 2.24111e-19 $X=5.605 $Y=2.51
+ $X2=0 $Y2=0
cc_670 N_A_818_418#_c_842_n N_A_728_331#_M1013_g 0.017713f $X=8.33 $Y=1.275
+ $X2=0 $Y2=0
cc_671 N_A_818_418#_c_843_n N_A_728_331#_M1013_g 0.00179297f $X=8.7 $Y=1.78
+ $X2=0 $Y2=0
cc_672 N_A_818_418#_c_847_n N_A_728_331#_M1013_g 9.47689e-19 $X=8.135 $Y=2.905
+ $X2=0 $Y2=0
cc_673 N_A_818_418#_c_851_n N_A_728_331#_M1013_g 0.0029963f $X=8.455 $Y=1.44
+ $X2=0 $Y2=0
cc_674 N_A_818_418#_c_852_n N_A_728_331#_M1013_g 0.00522227f $X=8.455 $Y=1.44
+ $X2=0 $Y2=0
cc_675 N_A_818_418#_c_855_n N_A_728_331#_c_1014_n 0.00731883f $X=8.7 $Y=1.87
+ $X2=0 $Y2=0
cc_676 N_A_818_418#_c_860_n N_A_728_331#_c_1014_n 0.00265666f $X=7.41 $Y=2.905
+ $X2=0 $Y2=0
cc_677 N_A_818_418#_c_861_n N_A_728_331#_c_1014_n 0.0142322f $X=8.05 $Y=2.99
+ $X2=0 $Y2=0
cc_678 N_A_818_418#_c_847_n N_A_728_331#_c_1014_n 0.0278842f $X=8.135 $Y=2.905
+ $X2=0 $Y2=0
cc_679 N_A_818_418#_c_843_n N_A_728_331#_c_1015_n 0.00285661f $X=8.7 $Y=1.78
+ $X2=0 $Y2=0
cc_680 N_A_818_418#_c_847_n N_A_728_331#_c_1015_n 0.00570974f $X=8.135 $Y=2.905
+ $X2=0 $Y2=0
cc_681 N_A_818_418#_c_851_n N_A_728_331#_c_1015_n 3.54458e-19 $X=8.455 $Y=1.44
+ $X2=0 $Y2=0
cc_682 N_A_818_418#_c_846_n N_A_728_331#_c_1016_n 0.00408573f $X=5.26 $Y=1.085
+ $X2=0 $Y2=0
cc_683 N_A_818_418#_c_859_n N_A_728_331#_c_1108_n 0.00999472f $X=7.315 $Y=2.51
+ $X2=0 $Y2=0
cc_684 N_A_818_418#_c_850_n N_A_728_331#_c_1108_n 0.0180717f $X=5.62 $Y=2.005
+ $X2=0 $Y2=0
cc_685 N_A_818_418#_c_859_n N_A_728_331#_c_1017_n 0.027879f $X=7.315 $Y=2.51
+ $X2=0 $Y2=0
cc_686 N_A_818_418#_c_846_n N_A_728_331#_c_1038_n 0.0251507f $X=5.26 $Y=1.085
+ $X2=0 $Y2=0
cc_687 N_A_818_418#_c_850_n N_A_728_331#_c_1038_n 0.0104702f $X=5.62 $Y=2.005
+ $X2=0 $Y2=0
cc_688 N_A_818_418#_c_859_n N_A_728_331#_c_1040_n 0.0209746f $X=7.315 $Y=2.51
+ $X2=0 $Y2=0
cc_689 N_A_818_418#_c_859_n N_A_728_331#_c_1019_n 0.0212266f $X=7.315 $Y=2.51
+ $X2=0 $Y2=0
cc_690 N_A_818_418#_c_846_n N_A_728_331#_c_1008_n 0.0135309f $X=5.26 $Y=1.085
+ $X2=0 $Y2=0
cc_691 N_A_818_418#_c_850_n N_A_728_331#_c_1008_n 0.00913506f $X=5.62 $Y=2.005
+ $X2=0 $Y2=0
cc_692 N_A_818_418#_c_859_n N_A_728_331#_c_1021_n 0.00761439f $X=7.315 $Y=2.51
+ $X2=0 $Y2=0
cc_693 N_A_818_418#_c_859_n N_CLK_c_1168_n 0.0159755f $X=7.315 $Y=2.51 $X2=0
+ $Y2=0
cc_694 N_A_818_418#_c_860_n N_CLK_c_1168_n 0.00689286f $X=7.41 $Y=2.905 $X2=0
+ $Y2=0
cc_695 N_A_818_418#_c_862_n N_CLK_c_1168_n 0.00449412f $X=7.505 $Y=2.99 $X2=0
+ $Y2=0
cc_696 N_A_818_418#_c_855_n N_A_1800_291#_c_1206_n 0.0322797f $X=8.7 $Y=1.87
+ $X2=0 $Y2=0
cc_697 N_A_818_418#_c_852_n N_A_1800_291#_c_1206_n 0.0212044f $X=8.455 $Y=1.44
+ $X2=0 $Y2=0
cc_698 N_A_818_418#_c_852_n N_A_1800_291#_c_1207_n 0.00528894f $X=8.455 $Y=1.44
+ $X2=0 $Y2=0
cc_699 N_A_818_418#_c_852_n N_A_1800_291#_c_1210_n 4.54987e-19 $X=8.455 $Y=1.44
+ $X2=0 $Y2=0
cc_700 N_A_818_418#_c_855_n N_A_1800_291#_c_1241_n 2.3665e-19 $X=8.7 $Y=1.87
+ $X2=0 $Y2=0
cc_701 N_A_818_418#_c_861_n N_A_1586_149#_M1028_d 0.00180442f $X=8.05 $Y=2.99
+ $X2=0 $Y2=0
cc_702 N_A_818_418#_c_847_n N_A_1586_149#_M1028_d 0.0211819f $X=8.135 $Y=2.905
+ $X2=0 $Y2=0
cc_703 N_A_818_418#_c_842_n N_A_1586_149#_c_1314_n 0.010471f $X=8.33 $Y=1.275
+ $X2=0 $Y2=0
cc_704 N_A_818_418#_c_851_n N_A_1586_149#_c_1314_n 0.0325809f $X=8.455 $Y=1.44
+ $X2=0 $Y2=0
cc_705 N_A_818_418#_c_852_n N_A_1586_149#_c_1314_n 0.0100446f $X=8.455 $Y=1.44
+ $X2=0 $Y2=0
cc_706 N_A_818_418#_c_855_n N_A_1586_149#_c_1307_n 0.00605713f $X=8.7 $Y=1.87
+ $X2=0 $Y2=0
cc_707 N_A_818_418#_c_847_n N_A_1586_149#_c_1307_n 0.0217186f $X=8.135 $Y=2.905
+ $X2=0 $Y2=0
cc_708 N_A_818_418#_c_842_n N_A_1586_149#_c_1298_n 2.62577e-19 $X=8.33 $Y=1.275
+ $X2=0 $Y2=0
cc_709 N_A_818_418#_c_843_n N_A_1586_149#_c_1298_n 0.00380843f $X=8.7 $Y=1.78
+ $X2=0 $Y2=0
cc_710 N_A_818_418#_c_855_n N_A_1586_149#_c_1298_n 0.00434641f $X=8.7 $Y=1.87
+ $X2=0 $Y2=0
cc_711 N_A_818_418#_c_847_n N_A_1586_149#_c_1298_n 0.00840422f $X=8.135 $Y=2.905
+ $X2=0 $Y2=0
cc_712 N_A_818_418#_c_851_n N_A_1586_149#_c_1298_n 0.0242956f $X=8.455 $Y=1.44
+ $X2=0 $Y2=0
cc_713 N_A_818_418#_c_852_n N_A_1586_149#_c_1298_n 0.00983263f $X=8.455 $Y=1.44
+ $X2=0 $Y2=0
cc_714 N_A_818_418#_c_855_n N_A_1586_149#_c_1309_n 0.012081f $X=8.7 $Y=1.87
+ $X2=0 $Y2=0
cc_715 N_A_818_418#_c_847_n N_A_1586_149#_c_1309_n 0.0133994f $X=8.135 $Y=2.905
+ $X2=0 $Y2=0
cc_716 N_A_818_418#_c_851_n N_A_1586_149#_c_1309_n 0.00496924f $X=8.455 $Y=1.44
+ $X2=0 $Y2=0
cc_717 N_A_818_418#_c_852_n N_A_1586_149#_c_1309_n 0.00381709f $X=8.455 $Y=1.44
+ $X2=0 $Y2=0
cc_718 N_A_818_418#_c_842_n N_A_1586_149#_c_1300_n 0.00560477f $X=8.33 $Y=1.275
+ $X2=0 $Y2=0
cc_719 N_A_818_418#_c_859_n N_VPWR_M1029_d 0.0183113f $X=7.315 $Y=2.51 $X2=0
+ $Y2=0
cc_720 N_A_818_418#_c_840_n N_VPWR_c_1495_n 7.35405e-19 $X=4.18 $Y=2.35 $X2=0
+ $Y2=0
cc_721 N_A_818_418#_c_858_n N_VPWR_c_1495_n 0.0159324f $X=5.62 $Y=2.815 $X2=0
+ $Y2=0
cc_722 N_A_818_418#_c_859_n N_VPWR_c_1495_n 0.00237526f $X=7.315 $Y=2.51 $X2=0
+ $Y2=0
cc_723 N_A_818_418#_c_859_n N_VPWR_c_1508_n 0.0108459f $X=7.315 $Y=2.51 $X2=0
+ $Y2=0
cc_724 N_A_818_418#_c_861_n N_VPWR_c_1508_n 0.0467393f $X=8.05 $Y=2.99 $X2=0
+ $Y2=0
cc_725 N_A_818_418#_c_862_n N_VPWR_c_1508_n 0.013574f $X=7.505 $Y=2.99 $X2=0
+ $Y2=0
cc_726 N_A_818_418#_c_858_n N_VPWR_c_1512_n 0.0150806f $X=5.62 $Y=2.815 $X2=0
+ $Y2=0
cc_727 N_A_818_418#_c_859_n N_VPWR_c_1512_n 0.0398389f $X=7.315 $Y=2.51 $X2=0
+ $Y2=0
cc_728 N_A_818_418#_c_855_n N_VPWR_c_1491_n 0.00384901f $X=8.7 $Y=1.87 $X2=0
+ $Y2=0
cc_729 N_A_818_418#_c_858_n N_VPWR_c_1491_n 0.0131546f $X=5.62 $Y=2.815 $X2=0
+ $Y2=0
cc_730 N_A_818_418#_c_859_n N_VPWR_c_1491_n 0.0275274f $X=7.315 $Y=2.51 $X2=0
+ $Y2=0
cc_731 N_A_818_418#_c_861_n N_VPWR_c_1491_n 0.0270012f $X=8.05 $Y=2.99 $X2=0
+ $Y2=0
cc_732 N_A_818_418#_c_862_n N_VPWR_c_1491_n 0.00737799f $X=7.505 $Y=2.99 $X2=0
+ $Y2=0
cc_733 N_A_818_418#_c_840_n N_A_70_74#_c_1653_n 0.0126935f $X=4.18 $Y=2.35 $X2=0
+ $Y2=0
cc_734 N_A_818_418#_M1035_g N_A_70_74#_c_1640_n 0.00741469f $X=4.265 $Y=1.37
+ $X2=0 $Y2=0
cc_735 N_A_818_418#_c_840_n N_A_70_74#_c_1641_n 0.00727448f $X=4.18 $Y=2.35
+ $X2=0 $Y2=0
cc_736 N_A_818_418#_M1035_g N_A_70_74#_c_1641_n 0.0268581f $X=4.265 $Y=1.37
+ $X2=0 $Y2=0
cc_737 N_A_818_418#_c_844_n N_A_70_74#_c_1641_n 5.73127e-19 $X=4.81 $Y=2.075
+ $X2=0 $Y2=0
cc_738 N_A_818_418#_c_845_n N_A_70_74#_c_1641_n 0.0103062f $X=4.645 $Y=2.075
+ $X2=0 $Y2=0
cc_739 N_A_818_418#_c_846_n N_A_70_74#_c_1641_n 0.00560911f $X=5.26 $Y=1.085
+ $X2=0 $Y2=0
cc_740 N_A_818_418#_c_848_n N_A_70_74#_c_1641_n 0.0256551f $X=5.15 $Y=2.075
+ $X2=0 $Y2=0
cc_741 N_A_818_418#_c_850_n N_A_70_74#_c_1641_n 0.00236354f $X=5.62 $Y=2.005
+ $X2=0 $Y2=0
cc_742 N_A_818_418#_c_840_n N_A_70_74#_c_1656_n 0.0116545f $X=4.18 $Y=2.35 $X2=0
+ $Y2=0
cc_743 N_A_818_418#_c_845_n N_A_70_74#_c_1657_n 0.0126159f $X=4.645 $Y=2.075
+ $X2=0 $Y2=0
cc_744 N_A_818_418#_c_858_n N_A_70_74#_c_1657_n 0.00966629f $X=5.62 $Y=2.815
+ $X2=0 $Y2=0
cc_745 N_A_818_418#_c_848_n N_A_70_74#_c_1657_n 0.0185116f $X=5.15 $Y=2.075
+ $X2=0 $Y2=0
cc_746 N_A_818_418#_c_866_n N_A_70_74#_c_1657_n 0.00506182f $X=5.605 $Y=2.51
+ $X2=0 $Y2=0
cc_747 N_A_818_418#_c_842_n N_VGND_c_1864_n 8.63546e-19 $X=8.33 $Y=1.275 $X2=0
+ $Y2=0
cc_748 N_A_818_418#_M1035_g N_A_614_81#_c_2000_n 4.73936e-19 $X=4.265 $Y=1.37
+ $X2=0 $Y2=0
cc_749 N_A_818_418#_M1035_g N_A_614_81#_c_2001_n 0.00301077f $X=4.265 $Y=1.37
+ $X2=0 $Y2=0
cc_750 N_A_818_418#_c_844_n N_A_614_81#_c_2001_n 0.00492069f $X=4.81 $Y=2.075
+ $X2=0 $Y2=0
cc_751 N_A_818_418#_c_846_n N_A_614_81#_c_2001_n 0.0435989f $X=5.26 $Y=1.085
+ $X2=0 $Y2=0
cc_752 N_A_818_418#_c_848_n N_A_614_81#_c_2001_n 0.00853807f $X=5.15 $Y=2.075
+ $X2=0 $Y2=0
cc_753 N_A_818_418#_c_842_n N_A_1499_149#_c_2025_n 0.0127492f $X=8.33 $Y=1.275
+ $X2=0 $Y2=0
cc_754 N_A_818_418#_c_852_n N_A_1499_149#_c_2025_n 5.41815e-19 $X=8.455 $Y=1.44
+ $X2=0 $Y2=0
cc_755 N_A_818_418#_c_842_n N_A_1499_149#_c_2027_n 0.00461776f $X=8.33 $Y=1.275
+ $X2=0 $Y2=0
cc_756 N_A_728_331#_c_1005_n N_CLK_c_1167_n 0.0170252f $X=6.45 $Y=1.34 $X2=-0.19
+ $Y2=-0.245
cc_757 N_A_728_331#_c_1007_n N_CLK_c_1167_n 0.0182609f $X=6.795 $Y=0.8 $X2=-0.19
+ $Y2=-0.245
cc_758 N_A_728_331#_c_1011_n N_CLK_c_1168_n 0.0191733f $X=5.845 $Y=1.765 $X2=0
+ $Y2=0
cc_759 N_A_728_331#_c_1016_n N_CLK_c_1168_n 0.0031001f $X=6.18 $Y=1.84 $X2=0
+ $Y2=0
cc_760 N_A_728_331#_c_1006_n N_CLK_c_1168_n 0.00638468f $X=6.45 $Y=1.505 $X2=0
+ $Y2=0
cc_761 N_A_728_331#_c_1007_n N_CLK_c_1168_n 0.00126299f $X=6.795 $Y=0.8 $X2=0
+ $Y2=0
cc_762 N_A_728_331#_c_1040_n N_CLK_c_1168_n 0.0147725f $X=6.705 $Y=2.047 $X2=0
+ $Y2=0
cc_763 N_A_728_331#_c_1019_n N_CLK_c_1168_n 0.00647792f $X=7.035 $Y=2.047 $X2=0
+ $Y2=0
cc_764 N_A_728_331#_c_1008_n N_CLK_c_1168_n 0.0176885f $X=5.845 $Y=1.552 $X2=0
+ $Y2=0
cc_765 N_A_728_331#_c_1021_n N_CLK_c_1168_n 0.00827568f $X=7.34 $Y=1.795 $X2=0
+ $Y2=0
cc_766 N_A_728_331#_M1003_d CLK 0.00277495f $X=6.655 $Y=0.49 $X2=0 $Y2=0
cc_767 N_A_728_331#_c_1005_n CLK 0.00994406f $X=6.45 $Y=1.34 $X2=0 $Y2=0
cc_768 N_A_728_331#_c_1006_n CLK 0.0259649f $X=6.45 $Y=1.505 $X2=0 $Y2=0
cc_769 N_A_728_331#_c_1007_n CLK 0.0173596f $X=6.795 $Y=0.8 $X2=0 $Y2=0
cc_770 N_A_728_331#_c_1019_n CLK 0.0206641f $X=7.035 $Y=2.047 $X2=0 $Y2=0
cc_771 N_A_728_331#_c_1008_n CLK 2.34167e-19 $X=5.845 $Y=1.552 $X2=0 $Y2=0
cc_772 N_A_728_331#_M1013_g N_A_1586_149#_c_1314_n 0.00269433f $X=7.855 $Y=0.955
+ $X2=0 $Y2=0
cc_773 N_A_728_331#_c_1015_n N_A_1586_149#_c_1314_n 0.00159115f $X=8.02 $Y=1.795
+ $X2=0 $Y2=0
cc_774 N_A_728_331#_c_1014_n N_A_1586_149#_c_1307_n 8.61107e-19 $X=8.02 $Y=1.87
+ $X2=0 $Y2=0
cc_775 N_A_728_331#_c_1014_n N_A_1586_149#_c_1309_n 5.53784e-19 $X=8.02 $Y=1.87
+ $X2=0 $Y2=0
cc_776 N_A_728_331#_c_1108_n N_VPWR_M1029_d 0.00891089f $X=6.265 $Y=2.005 $X2=0
+ $Y2=0
cc_777 N_A_728_331#_c_1040_n N_VPWR_M1029_d 0.00725219f $X=6.705 $Y=2.047 $X2=0
+ $Y2=0
cc_778 N_A_728_331#_c_1010_n N_VPWR_c_1495_n 7.35405e-19 $X=3.73 $Y=2.35 $X2=0
+ $Y2=0
cc_779 N_A_728_331#_c_1011_n N_VPWR_c_1495_n 0.00333203f $X=5.845 $Y=1.765 $X2=0
+ $Y2=0
cc_780 N_A_728_331#_c_1014_n N_VPWR_c_1508_n 0.00301083f $X=8.02 $Y=1.87 $X2=0
+ $Y2=0
cc_781 N_A_728_331#_c_1011_n N_VPWR_c_1512_n 0.00623235f $X=5.845 $Y=1.765 $X2=0
+ $Y2=0
cc_782 N_A_728_331#_c_1011_n N_VPWR_c_1491_n 0.00436423f $X=5.845 $Y=1.765 $X2=0
+ $Y2=0
cc_783 N_A_728_331#_c_1014_n N_VPWR_c_1491_n 0.00378742f $X=8.02 $Y=1.87 $X2=0
+ $Y2=0
cc_784 N_A_728_331#_c_1010_n N_A_70_74#_c_1650_n 0.00137259f $X=3.73 $Y=2.35
+ $X2=0 $Y2=0
cc_785 N_A_728_331#_c_1010_n N_A_70_74#_c_1652_n 0.00551652f $X=3.73 $Y=2.35
+ $X2=0 $Y2=0
cc_786 N_A_728_331#_c_1010_n N_A_70_74#_c_1653_n 0.0116302f $X=3.73 $Y=2.35
+ $X2=0 $Y2=0
cc_787 N_A_728_331#_M1004_g N_A_70_74#_c_1640_n 0.0123257f $X=3.835 $Y=1.37
+ $X2=0 $Y2=0
cc_788 N_A_728_331#_c_1004_n N_A_70_74#_c_1640_n 9.00795e-19 $X=3.775 $Y=1.805
+ $X2=0 $Y2=0
cc_789 N_A_728_331#_M1004_g N_A_70_74#_c_1641_n 7.75671e-19 $X=3.835 $Y=1.37
+ $X2=0 $Y2=0
cc_790 N_A_728_331#_M1004_g N_A_70_74#_c_1643_n 0.00370416f $X=3.835 $Y=1.37
+ $X2=0 $Y2=0
cc_791 N_A_728_331#_c_1004_n N_A_70_74#_c_1643_n 0.00142072f $X=3.775 $Y=1.805
+ $X2=0 $Y2=0
cc_792 N_A_728_331#_c_1005_n N_VGND_M1030_d 0.0103537f $X=6.45 $Y=1.34 $X2=0
+ $Y2=0
cc_793 N_A_728_331#_c_1007_n N_VGND_M1030_d 0.00927667f $X=6.795 $Y=0.8 $X2=0
+ $Y2=0
cc_794 N_A_728_331#_c_1000_n N_VGND_c_1853_n 0.00688197f $X=5.4 $Y=0.34 $X2=0
+ $Y2=0
cc_795 N_A_728_331#_c_1000_n N_VGND_c_1862_n 0.00849616f $X=5.4 $Y=0.34 $X2=0
+ $Y2=0
cc_796 N_A_728_331#_c_1001_n N_VGND_c_1862_n 0.0095216f $X=3.91 $Y=0.34 $X2=0
+ $Y2=0
cc_797 N_A_728_331#_c_1000_n N_VGND_c_1875_n 0.0107407f $X=5.4 $Y=0.34 $X2=0
+ $Y2=0
cc_798 N_A_728_331#_M1004_g N_A_614_81#_c_2000_n 0.0139459f $X=3.835 $Y=1.37
+ $X2=0 $Y2=0
cc_799 N_A_728_331#_c_1000_n N_A_614_81#_c_2000_n 0.00598631f $X=5.4 $Y=0.34
+ $X2=0 $Y2=0
cc_800 N_A_728_331#_M1030_g N_A_614_81#_c_2000_n 5.30126e-19 $X=5.475 $Y=0.86
+ $X2=0 $Y2=0
cc_801 N_A_728_331#_M1030_g N_A_614_81#_c_2001_n 0.00494998f $X=5.475 $Y=0.86
+ $X2=0 $Y2=0
cc_802 N_A_728_331#_c_1012_n N_A_1499_149#_c_2024_n 2.85935e-19 $X=7.78 $Y=1.795
+ $X2=0 $Y2=0
cc_803 N_A_728_331#_M1013_g N_A_1499_149#_c_2024_n 0.0010439f $X=7.855 $Y=0.955
+ $X2=0 $Y2=0
cc_804 N_A_728_331#_M1013_g N_A_1499_149#_c_2025_n 0.0130579f $X=7.855 $Y=0.955
+ $X2=0 $Y2=0
cc_805 N_CLK_c_1168_n N_VPWR_c_1508_n 0.00336577f $X=6.645 $Y=1.765 $X2=0 $Y2=0
cc_806 N_CLK_c_1168_n N_VPWR_c_1512_n 0.0106997f $X=6.645 $Y=1.765 $X2=0 $Y2=0
cc_807 N_CLK_c_1168_n N_VPWR_c_1491_n 0.00445301f $X=6.645 $Y=1.765 $X2=0 $Y2=0
cc_808 N_CLK_c_1167_n N_VGND_c_1853_n 2.58254e-19 $X=6.58 $Y=1.34 $X2=0 $Y2=0
cc_809 N_CLK_c_1167_n N_VGND_c_1864_n 7.26245e-19 $X=6.58 $Y=1.34 $X2=0 $Y2=0
cc_810 N_A_1800_291#_c_1211_n N_A_1586_149#_M1017_g 0.00518619f $X=10.59 $Y=1.95
+ $X2=0 $Y2=0
cc_811 N_A_1800_291#_c_1212_n N_A_1586_149#_M1017_g 0.00799557f $X=10.59
+ $Y=0.557 $X2=0 $Y2=0
cc_812 N_A_1800_291#_c_1211_n N_A_1586_149#_c_1294_n 0.00370178f $X=10.59
+ $Y=1.95 $X2=0 $Y2=0
cc_813 N_A_1800_291#_c_1245_p N_A_1586_149#_c_1303_n 0.0158205f $X=10.505
+ $Y=2.035 $X2=0 $Y2=0
cc_814 N_A_1800_291#_c_1211_n N_A_1586_149#_c_1303_n 0.00163529f $X=10.59
+ $Y=1.95 $X2=0 $Y2=0
cc_815 N_A_1800_291#_c_1216_n N_A_1586_149#_c_1303_n 0.00637605f $X=10.16
+ $Y=2.167 $X2=0 $Y2=0
cc_816 N_A_1800_291#_c_1211_n N_A_1586_149#_c_1304_n 0.0018715f $X=10.59 $Y=1.95
+ $X2=0 $Y2=0
cc_817 N_A_1800_291#_c_1216_n N_A_1586_149#_c_1304_n 5.17071e-19 $X=10.16
+ $Y=2.167 $X2=0 $Y2=0
cc_818 N_A_1800_291#_c_1211_n N_A_1586_149#_c_1295_n 0.00115321f $X=10.59
+ $Y=1.95 $X2=0 $Y2=0
cc_819 N_A_1800_291#_c_1206_n N_A_1586_149#_c_1307_n 0.00117311f $X=9.12 $Y=1.87
+ $X2=0 $Y2=0
cc_820 N_A_1800_291#_c_1241_n N_A_1586_149#_c_1307_n 9.30423e-19 $X=9.33
+ $Y=2.035 $X2=0 $Y2=0
cc_821 N_A_1800_291#_c_1206_n N_A_1586_149#_c_1298_n 0.0025901f $X=9.12 $Y=1.87
+ $X2=0 $Y2=0
cc_822 N_A_1800_291#_c_1207_n N_A_1586_149#_c_1298_n 0.00374138f $X=9.225
+ $Y=1.455 $X2=0 $Y2=0
cc_823 N_A_1800_291#_c_1210_n N_A_1586_149#_c_1298_n 0.0338519f $X=9.165 $Y=1.62
+ $X2=0 $Y2=0
cc_824 N_A_1800_291#_c_1206_n N_A_1586_149#_c_1299_n 0.00342751f $X=9.12 $Y=1.87
+ $X2=0 $Y2=0
cc_825 N_A_1800_291#_c_1207_n N_A_1586_149#_c_1299_n 0.01522f $X=9.225 $Y=1.455
+ $X2=0 $Y2=0
cc_826 N_A_1800_291#_c_1209_n N_A_1586_149#_c_1299_n 0.0167639f $X=9.365 $Y=0.94
+ $X2=0 $Y2=0
cc_827 N_A_1800_291#_c_1210_n N_A_1586_149#_c_1299_n 0.0181585f $X=9.165 $Y=1.62
+ $X2=0 $Y2=0
cc_828 N_A_1800_291#_c_1211_n N_A_1586_149#_c_1299_n 0.0259151f $X=10.59 $Y=1.95
+ $X2=0 $Y2=0
cc_829 N_A_1800_291#_c_1212_n N_A_1586_149#_c_1299_n 0.00784134f $X=10.59
+ $Y=0.557 $X2=0 $Y2=0
cc_830 N_A_1800_291#_c_1206_n N_A_1586_149#_c_1309_n 0.00105515f $X=9.12 $Y=1.87
+ $X2=0 $Y2=0
cc_831 N_A_1800_291#_c_1210_n N_A_1586_149#_c_1309_n 0.00190038f $X=9.165
+ $Y=1.62 $X2=0 $Y2=0
cc_832 N_A_1800_291#_c_1241_n N_A_1586_149#_c_1309_n 0.012306f $X=9.33 $Y=2.035
+ $X2=0 $Y2=0
cc_833 N_A_1800_291#_c_1245_p N_A_1586_149#_c_1301_n 0.00602016f $X=10.505
+ $Y=2.035 $X2=0 $Y2=0
cc_834 N_A_1800_291#_c_1211_n N_A_1586_149#_c_1301_n 0.0343015f $X=10.59 $Y=1.95
+ $X2=0 $Y2=0
cc_835 N_A_1800_291#_c_1216_n N_A_1586_149#_c_1301_n 8.70427e-19 $X=10.16
+ $Y=2.167 $X2=0 $Y2=0
cc_836 N_A_1800_291#_c_1212_n N_A_1586_149#_c_1301_n 0.00667101f $X=10.59
+ $Y=0.557 $X2=0 $Y2=0
cc_837 N_A_1800_291#_c_1241_n N_VPWR_M1018_d 0.00132656f $X=9.33 $Y=2.035 $X2=0
+ $Y2=0
cc_838 N_A_1800_291#_c_1230_n N_VPWR_M1018_d 0.00836353f $X=9.83 $Y=2.167 $X2=0
+ $Y2=0
cc_839 N_A_1800_291#_c_1245_p N_VPWR_M1016_d 0.00665364f $X=10.505 $Y=2.035
+ $X2=0 $Y2=0
cc_840 N_A_1800_291#_c_1211_n N_VPWR_M1016_d 0.00275002f $X=10.59 $Y=1.95 $X2=0
+ $Y2=0
cc_841 N_A_1800_291#_c_1206_n N_VPWR_c_1496_n 0.0050551f $X=9.12 $Y=1.87 $X2=0
+ $Y2=0
cc_842 N_A_1800_291#_c_1241_n N_VPWR_c_1496_n 0.00555396f $X=9.33 $Y=2.035 $X2=0
+ $Y2=0
cc_843 N_A_1800_291#_c_1230_n N_VPWR_c_1496_n 0.0231298f $X=9.83 $Y=2.167 $X2=0
+ $Y2=0
cc_844 N_A_1800_291#_c_1216_n N_VPWR_c_1496_n 0.00641761f $X=10.16 $Y=2.167
+ $X2=0 $Y2=0
cc_845 N_A_1800_291#_c_1245_p N_VPWR_c_1497_n 0.0218664f $X=10.505 $Y=2.035
+ $X2=0 $Y2=0
cc_846 N_A_1800_291#_c_1216_n N_VPWR_c_1497_n 0.00637407f $X=10.16 $Y=2.167
+ $X2=0 $Y2=0
cc_847 N_A_1800_291#_c_1206_n N_VPWR_c_1491_n 0.00384901f $X=9.12 $Y=1.87 $X2=0
+ $Y2=0
cc_848 N_A_1800_291#_c_1211_n N_Q_N_c_1793_n 0.0186743f $X=10.59 $Y=1.95 $X2=0
+ $Y2=0
cc_849 N_A_1800_291#_c_1211_n Q_N 0.0206203f $X=10.59 $Y=1.95 $X2=0 $Y2=0
cc_850 N_A_1800_291#_c_1208_n N_VGND_c_1854_n 0.00904236f $X=9.365 $Y=0.865
+ $X2=0 $Y2=0
cc_851 N_A_1800_291#_c_1212_n N_VGND_c_1854_n 0.0127168f $X=10.59 $Y=0.557 $X2=0
+ $Y2=0
cc_852 N_A_1800_291#_c_1211_n N_VGND_c_1855_n 0.0247783f $X=10.59 $Y=1.95 $X2=0
+ $Y2=0
cc_853 N_A_1800_291#_c_1212_n N_VGND_c_1855_n 0.0333158f $X=10.59 $Y=0.557 $X2=0
+ $Y2=0
cc_854 N_A_1800_291#_c_1208_n N_VGND_c_1864_n 0.00383152f $X=9.365 $Y=0.865
+ $X2=0 $Y2=0
cc_855 N_A_1800_291#_c_1212_n N_VGND_c_1866_n 0.0200848f $X=10.59 $Y=0.557 $X2=0
+ $Y2=0
cc_856 N_A_1800_291#_c_1208_n N_VGND_c_1875_n 0.00762539f $X=9.365 $Y=0.865
+ $X2=0 $Y2=0
cc_857 N_A_1800_291#_c_1209_n N_VGND_c_1875_n 0.00141224f $X=9.365 $Y=0.94 $X2=0
+ $Y2=0
cc_858 N_A_1800_291#_c_1212_n N_VGND_c_1875_n 0.0169453f $X=10.59 $Y=0.557 $X2=0
+ $Y2=0
cc_859 N_A_1800_291#_c_1208_n N_A_1499_149#_c_2027_n 7.31217e-19 $X=9.365
+ $Y=0.865 $X2=0 $Y2=0
cc_860 N_A_1800_291#_c_1209_n N_A_1499_149#_c_2027_n 0.00244996f $X=9.365
+ $Y=0.94 $X2=0 $Y2=0
cc_861 N_A_1586_149#_c_1306_n N_A_2363_352#_c_1433_n 0.00651951f $X=11.74
+ $Y=1.685 $X2=0 $Y2=0
cc_862 N_A_1586_149#_c_1301_n N_A_2363_352#_c_1433_n 0.0211299f $X=11.74 $Y=1.31
+ $X2=0 $Y2=0
cc_863 N_A_1586_149#_c_1306_n N_A_2363_352#_c_1440_n 0.0200384f $X=11.74
+ $Y=1.685 $X2=0 $Y2=0
cc_864 N_A_1586_149#_M1020_g N_A_2363_352#_c_1434_n 0.00874126f $X=12.05 $Y=0.69
+ $X2=0 $Y2=0
cc_865 N_A_1586_149#_c_1301_n N_A_2363_352#_c_1436_n 0.0054628f $X=11.74 $Y=1.31
+ $X2=0 $Y2=0
cc_866 N_A_1586_149#_c_1307_n N_VPWR_c_1496_n 0.00262979f $X=8.475 $Y=2.155
+ $X2=0 $Y2=0
cc_867 N_A_1586_149#_c_1303_n N_VPWR_c_1497_n 0.00394923f $X=10.22 $Y=1.87 $X2=0
+ $Y2=0
cc_868 N_A_1586_149#_c_1304_n N_VPWR_c_1497_n 0.01173f $X=10.755 $Y=1.685 $X2=0
+ $Y2=0
cc_869 N_A_1586_149#_c_1305_n N_VPWR_c_1497_n 5.10325e-19 $X=11.205 $Y=1.685
+ $X2=0 $Y2=0
cc_870 N_A_1586_149#_c_1301_n N_VPWR_c_1497_n 5.87989e-19 $X=11.74 $Y=1.31 $X2=0
+ $Y2=0
cc_871 N_A_1586_149#_c_1304_n N_VPWR_c_1498_n 0.00467292f $X=10.755 $Y=1.685
+ $X2=0 $Y2=0
cc_872 N_A_1586_149#_c_1305_n N_VPWR_c_1498_n 0.00467292f $X=11.205 $Y=1.685
+ $X2=0 $Y2=0
cc_873 N_A_1586_149#_c_1304_n N_VPWR_c_1499_n 6.7751e-19 $X=10.755 $Y=1.685
+ $X2=0 $Y2=0
cc_874 N_A_1586_149#_c_1305_n N_VPWR_c_1499_n 0.017941f $X=11.205 $Y=1.685 $X2=0
+ $Y2=0
cc_875 N_A_1586_149#_c_1306_n N_VPWR_c_1499_n 0.0140731f $X=11.74 $Y=1.685 $X2=0
+ $Y2=0
cc_876 N_A_1586_149#_c_1301_n N_VPWR_c_1499_n 0.00877461f $X=11.74 $Y=1.31 $X2=0
+ $Y2=0
cc_877 N_A_1586_149#_c_1306_n N_VPWR_c_1500_n 0.00348324f $X=11.74 $Y=1.685
+ $X2=0 $Y2=0
cc_878 N_A_1586_149#_c_1306_n N_VPWR_c_1509_n 0.00445514f $X=11.74 $Y=1.685
+ $X2=0 $Y2=0
cc_879 N_A_1586_149#_c_1303_n N_VPWR_c_1491_n 0.00384901f $X=10.22 $Y=1.87 $X2=0
+ $Y2=0
cc_880 N_A_1586_149#_c_1304_n N_VPWR_c_1491_n 0.00471987f $X=10.755 $Y=1.685
+ $X2=0 $Y2=0
cc_881 N_A_1586_149#_c_1305_n N_VPWR_c_1491_n 0.00471987f $X=11.205 $Y=1.685
+ $X2=0 $Y2=0
cc_882 N_A_1586_149#_c_1306_n N_VPWR_c_1491_n 0.00484898f $X=11.74 $Y=1.685
+ $X2=0 $Y2=0
cc_883 N_A_1586_149#_c_1309_n A_1755_389# 0.00367913f $X=8.81 $Y=2.01 $X2=-0.19
+ $Y2=-0.245
cc_884 N_A_1586_149#_c_1304_n N_Q_N_c_1793_n 0.00722149f $X=10.755 $Y=1.685
+ $X2=0 $Y2=0
cc_885 N_A_1586_149#_c_1305_n N_Q_N_c_1793_n 0.00522773f $X=11.205 $Y=1.685
+ $X2=0 $Y2=0
cc_886 N_A_1586_149#_c_1301_n N_Q_N_c_1793_n 0.0113712f $X=11.74 $Y=1.31 $X2=0
+ $Y2=0
cc_887 N_A_1586_149#_c_1295_n N_Q_N_c_1791_n 0.00521369f $X=11.145 $Y=1.185
+ $X2=0 $Y2=0
cc_888 N_A_1586_149#_c_1296_n N_Q_N_c_1791_n 2.74318e-19 $X=11.575 $Y=1.185
+ $X2=0 $Y2=0
cc_889 N_A_1586_149#_c_1295_n Q_N 0.00609559f $X=11.145 $Y=1.185 $X2=0 $Y2=0
cc_890 N_A_1586_149#_c_1296_n Q_N 0.0143409f $X=11.575 $Y=1.185 $X2=0 $Y2=0
cc_891 N_A_1586_149#_M1020_g Q_N 0.00393154f $X=12.05 $Y=0.69 $X2=0 $Y2=0
cc_892 N_A_1586_149#_c_1301_n Q_N 0.0807366f $X=11.74 $Y=1.31 $X2=0 $Y2=0
cc_893 N_A_1586_149#_M1017_g N_VGND_c_1854_n 0.00157764f $X=10.155 $Y=0.58 $X2=0
+ $Y2=0
cc_894 N_A_1586_149#_c_1299_n N_VGND_c_1854_n 0.0192815f $X=10.245 $Y=1.1 $X2=0
+ $Y2=0
cc_895 N_A_1586_149#_M1017_g N_VGND_c_1855_n 0.00300622f $X=10.155 $Y=0.58 $X2=0
+ $Y2=0
cc_896 N_A_1586_149#_c_1295_n N_VGND_c_1855_n 0.00400592f $X=11.145 $Y=1.185
+ $X2=0 $Y2=0
cc_897 N_A_1586_149#_c_1301_n N_VGND_c_1855_n 0.0048246f $X=11.74 $Y=1.31 $X2=0
+ $Y2=0
cc_898 N_A_1586_149#_c_1295_n N_VGND_c_1856_n 4.16356e-19 $X=11.145 $Y=1.185
+ $X2=0 $Y2=0
cc_899 N_A_1586_149#_c_1296_n N_VGND_c_1856_n 0.00689813f $X=11.575 $Y=1.185
+ $X2=0 $Y2=0
cc_900 N_A_1586_149#_M1020_g N_VGND_c_1856_n 0.00197289f $X=12.05 $Y=0.69 $X2=0
+ $Y2=0
cc_901 N_A_1586_149#_c_1301_n N_VGND_c_1856_n 7.47762e-19 $X=11.74 $Y=1.31 $X2=0
+ $Y2=0
cc_902 N_A_1586_149#_M1020_g N_VGND_c_1857_n 0.00293008f $X=12.05 $Y=0.69 $X2=0
+ $Y2=0
cc_903 N_A_1586_149#_M1017_g N_VGND_c_1866_n 0.00433162f $X=10.155 $Y=0.58 $X2=0
+ $Y2=0
cc_904 N_A_1586_149#_c_1295_n N_VGND_c_1869_n 0.00434272f $X=11.145 $Y=1.185
+ $X2=0 $Y2=0
cc_905 N_A_1586_149#_c_1296_n N_VGND_c_1869_n 0.00383152f $X=11.575 $Y=1.185
+ $X2=0 $Y2=0
cc_906 N_A_1586_149#_M1020_g N_VGND_c_1870_n 0.00461464f $X=12.05 $Y=0.69 $X2=0
+ $Y2=0
cc_907 N_A_1586_149#_M1017_g N_VGND_c_1875_n 0.00822018f $X=10.155 $Y=0.58 $X2=0
+ $Y2=0
cc_908 N_A_1586_149#_c_1295_n N_VGND_c_1875_n 0.00825283f $X=11.145 $Y=1.185
+ $X2=0 $Y2=0
cc_909 N_A_1586_149#_c_1296_n N_VGND_c_1875_n 0.0036906f $X=11.575 $Y=1.185
+ $X2=0 $Y2=0
cc_910 N_A_1586_149#_M1020_g N_VGND_c_1875_n 0.00912757f $X=12.05 $Y=0.69 $X2=0
+ $Y2=0
cc_911 N_A_1586_149#_M1013_d N_A_1499_149#_c_2025_n 0.0042087f $X=7.93 $Y=0.745
+ $X2=0 $Y2=0
cc_912 N_A_1586_149#_c_1314_n N_A_1499_149#_c_2025_n 0.0461856f $X=8.725 $Y=1.02
+ $X2=0 $Y2=0
cc_913 N_A_1586_149#_c_1299_n N_A_1499_149#_c_2025_n 0.00709406f $X=10.245
+ $Y=1.1 $X2=0 $Y2=0
cc_914 N_A_1586_149#_c_1300_n N_A_1499_149#_c_2025_n 0.0142962f $X=8.81 $Y=1.1
+ $X2=0 $Y2=0
cc_915 N_A_1586_149#_c_1299_n N_A_1499_149#_c_2027_n 0.0203727f $X=10.245 $Y=1.1
+ $X2=0 $Y2=0
cc_916 N_A_2363_352#_c_1433_n N_VPWR_c_1499_n 0.0110976f $X=12.1 $Y=1.945 $X2=0
+ $Y2=0
cc_917 N_A_2363_352#_c_1440_n N_VPWR_c_1499_n 0.0448464f $X=12.06 $Y=2.615 $X2=0
+ $Y2=0
cc_918 N_A_2363_352#_c_1437_n N_VPWR_c_1500_n 0.0261486f $X=12.915 $Y=1.765
+ $X2=0 $Y2=0
cc_919 N_A_2363_352#_c_1433_n N_VPWR_c_1500_n 0.0106305f $X=12.1 $Y=1.945 $X2=0
+ $Y2=0
cc_920 N_A_2363_352#_c_1440_n N_VPWR_c_1500_n 0.0706467f $X=12.06 $Y=2.615 $X2=0
+ $Y2=0
cc_921 N_A_2363_352#_c_1435_n N_VPWR_c_1500_n 0.0261101f $X=12.8 $Y=1.465 $X2=0
+ $Y2=0
cc_922 N_A_2363_352#_c_1436_n N_VPWR_c_1500_n 0.00389761f $X=13.365 $Y=1.532
+ $X2=0 $Y2=0
cc_923 N_A_2363_352#_c_1438_n N_VPWR_c_1502_n 0.0261486f $X=13.365 $Y=1.765
+ $X2=0 $Y2=0
cc_924 N_A_2363_352#_c_1436_n N_VPWR_c_1502_n 0.00152598f $X=13.365 $Y=1.532
+ $X2=0 $Y2=0
cc_925 N_A_2363_352#_c_1440_n N_VPWR_c_1509_n 0.00996859f $X=12.06 $Y=2.615
+ $X2=0 $Y2=0
cc_926 N_A_2363_352#_c_1437_n N_VPWR_c_1510_n 0.00445602f $X=12.915 $Y=1.765
+ $X2=0 $Y2=0
cc_927 N_A_2363_352#_c_1438_n N_VPWR_c_1510_n 0.00445602f $X=13.365 $Y=1.765
+ $X2=0 $Y2=0
cc_928 N_A_2363_352#_c_1437_n N_VPWR_c_1491_n 0.00861719f $X=12.915 $Y=1.765
+ $X2=0 $Y2=0
cc_929 N_A_2363_352#_c_1438_n N_VPWR_c_1491_n 0.00860566f $X=13.365 $Y=1.765
+ $X2=0 $Y2=0
cc_930 N_A_2363_352#_c_1440_n N_VPWR_c_1491_n 0.0131729f $X=12.06 $Y=2.615 $X2=0
+ $Y2=0
cc_931 N_A_2363_352#_c_1433_n Q_N 0.0130882f $X=12.1 $Y=1.945 $X2=0 $Y2=0
cc_932 N_A_2363_352#_c_1434_n Q_N 0.0259548f $X=12.265 $Y=0.515 $X2=0 $Y2=0
cc_933 N_A_2363_352#_c_1437_n N_Q_c_1823_n 0.00261316f $X=12.915 $Y=1.765 $X2=0
+ $Y2=0
cc_934 N_A_2363_352#_c_1438_n N_Q_c_1823_n 0.00188635f $X=13.365 $Y=1.765 $X2=0
+ $Y2=0
cc_935 N_A_2363_352#_c_1436_n N_Q_c_1823_n 0.00697862f $X=13.365 $Y=1.532 $X2=0
+ $Y2=0
cc_936 N_A_2363_352#_c_1437_n N_Q_c_1824_n 0.0109216f $X=12.915 $Y=1.765 $X2=0
+ $Y2=0
cc_937 N_A_2363_352#_c_1438_n N_Q_c_1824_n 0.0109216f $X=13.365 $Y=1.765 $X2=0
+ $Y2=0
cc_938 N_A_2363_352#_c_1437_n N_Q_c_1820_n 0.00116343f $X=12.915 $Y=1.765 $X2=0
+ $Y2=0
cc_939 N_A_2363_352#_M1012_g N_Q_c_1820_n 0.00405899f $X=13.01 $Y=0.74 $X2=0
+ $Y2=0
cc_940 N_A_2363_352#_c_1438_n N_Q_c_1820_n 0.00251865f $X=13.365 $Y=1.765 $X2=0
+ $Y2=0
cc_941 N_A_2363_352#_M1037_g N_Q_c_1820_n 0.0040077f $X=13.44 $Y=0.74 $X2=0
+ $Y2=0
cc_942 N_A_2363_352#_c_1435_n N_Q_c_1820_n 0.0249855f $X=12.8 $Y=1.465 $X2=0
+ $Y2=0
cc_943 N_A_2363_352#_c_1436_n N_Q_c_1820_n 0.0381787f $X=13.365 $Y=1.532 $X2=0
+ $Y2=0
cc_944 N_A_2363_352#_M1012_g Q 0.00320059f $X=13.01 $Y=0.74 $X2=0 $Y2=0
cc_945 N_A_2363_352#_M1037_g Q 0.00323247f $X=13.44 $Y=0.74 $X2=0 $Y2=0
cc_946 N_A_2363_352#_M1012_g N_Q_c_1822_n 0.00838251f $X=13.01 $Y=0.74 $X2=0
+ $Y2=0
cc_947 N_A_2363_352#_M1037_g N_Q_c_1822_n 0.00821863f $X=13.44 $Y=0.74 $X2=0
+ $Y2=0
cc_948 N_A_2363_352#_c_1434_n N_VGND_c_1856_n 0.00157123f $X=12.265 $Y=0.515
+ $X2=0 $Y2=0
cc_949 N_A_2363_352#_M1012_g N_VGND_c_1857_n 0.00610844f $X=13.01 $Y=0.74 $X2=0
+ $Y2=0
cc_950 N_A_2363_352#_c_1434_n N_VGND_c_1857_n 0.0562664f $X=12.265 $Y=0.515
+ $X2=0 $Y2=0
cc_951 N_A_2363_352#_c_1435_n N_VGND_c_1857_n 0.0209312f $X=12.8 $Y=1.465 $X2=0
+ $Y2=0
cc_952 N_A_2363_352#_c_1436_n N_VGND_c_1857_n 0.00586268f $X=13.365 $Y=1.532
+ $X2=0 $Y2=0
cc_953 N_A_2363_352#_M1037_g N_VGND_c_1859_n 0.00618831f $X=13.44 $Y=0.74 $X2=0
+ $Y2=0
cc_954 N_A_2363_352#_c_1434_n N_VGND_c_1870_n 0.0130739f $X=12.265 $Y=0.515
+ $X2=0 $Y2=0
cc_955 N_A_2363_352#_M1012_g N_VGND_c_1871_n 0.00433834f $X=13.01 $Y=0.74 $X2=0
+ $Y2=0
cc_956 N_A_2363_352#_M1037_g N_VGND_c_1871_n 0.00433834f $X=13.44 $Y=0.74 $X2=0
+ $Y2=0
cc_957 N_A_2363_352#_M1012_g N_VGND_c_1875_n 0.00824977f $X=13.01 $Y=0.74 $X2=0
+ $Y2=0
cc_958 N_A_2363_352#_M1037_g N_VGND_c_1875_n 0.00823359f $X=13.44 $Y=0.74 $X2=0
+ $Y2=0
cc_959 N_A_2363_352#_c_1434_n N_VGND_c_1875_n 0.0108215f $X=12.265 $Y=0.515
+ $X2=0 $Y2=0
cc_960 N_VPWR_c_1493_n N_A_70_74#_c_1644_n 0.036541f $X=0.345 $Y=2.17 $X2=0
+ $Y2=0
cc_961 N_VPWR_M1015_d N_A_70_74#_c_1646_n 0.0108781f $X=0.135 $Y=2.81 $X2=0
+ $Y2=0
cc_962 N_VPWR_c_1503_n N_A_70_74#_c_1646_n 0.0313278f $X=1.21 $Y=3.19 $X2=0
+ $Y2=0
cc_963 N_VPWR_c_1507_n N_A_70_74#_c_1646_n 0.00309506f $X=2.945 $Y=3.33 $X2=0
+ $Y2=0
cc_964 N_VPWR_c_1491_n N_A_70_74#_c_1646_n 0.00707017f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_965 N_VPWR_c_1493_n N_A_70_74#_c_1647_n 0.0152343f $X=0.345 $Y=2.17 $X2=0
+ $Y2=0
cc_966 N_VPWR_c_1503_n N_A_70_74#_c_1647_n 0.0271618f $X=1.21 $Y=3.19 $X2=0
+ $Y2=0
cc_967 N_VPWR_c_1491_n N_A_70_74#_c_1647_n 0.00204634f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_968 N_VPWR_c_1494_n N_A_70_74#_c_1648_n 0.0147095f $X=3.03 $Y=2.79 $X2=0
+ $Y2=0
cc_969 N_VPWR_c_1507_n N_A_70_74#_c_1648_n 0.0656248f $X=2.945 $Y=3.33 $X2=0
+ $Y2=0
cc_970 N_VPWR_c_1491_n N_A_70_74#_c_1648_n 0.0378114f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_971 N_VPWR_M1032_d N_A_70_74#_c_1649_n 0.00466656f $X=2.65 $Y=2.425 $X2=0
+ $Y2=0
cc_972 N_VPWR_c_1494_n N_A_70_74#_c_1649_n 0.0209842f $X=3.03 $Y=2.79 $X2=0
+ $Y2=0
cc_973 N_VPWR_M1032_d N_A_70_74#_c_1650_n 0.0100181f $X=2.65 $Y=2.425 $X2=0
+ $Y2=0
cc_974 N_VPWR_c_1494_n N_A_70_74#_c_1650_n 0.0201769f $X=3.03 $Y=2.79 $X2=0
+ $Y2=0
cc_975 N_VPWR_c_1494_n N_A_70_74#_c_1652_n 0.0203131f $X=3.03 $Y=2.79 $X2=0
+ $Y2=0
cc_976 N_VPWR_c_1495_n N_A_70_74#_c_1653_n 0.0485775f $X=5.99 $Y=3.33 $X2=0
+ $Y2=0
cc_977 N_VPWR_c_1491_n N_A_70_74#_c_1653_n 0.0283783f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_978 N_VPWR_c_1494_n N_A_70_74#_c_1654_n 0.014427f $X=3.03 $Y=2.79 $X2=0 $Y2=0
cc_979 N_VPWR_c_1495_n N_A_70_74#_c_1654_n 0.0121867f $X=5.99 $Y=3.33 $X2=0
+ $Y2=0
cc_980 N_VPWR_c_1491_n N_A_70_74#_c_1654_n 0.00660921f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_981 N_VPWR_c_1495_n N_A_70_74#_c_1656_n 0.0125688f $X=5.99 $Y=3.33 $X2=0
+ $Y2=0
cc_982 N_VPWR_c_1491_n N_A_70_74#_c_1656_n 0.00710542f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_983 N_VPWR_c_1495_n N_A_70_74#_c_1657_n 0.0118092f $X=5.99 $Y=3.33 $X2=0
+ $Y2=0
cc_984 N_VPWR_c_1491_n N_A_70_74#_c_1657_n 0.0155687f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_985 N_VPWR_c_1493_n N_A_70_74#_c_1642_n 7.16836e-19 $X=0.345 $Y=2.17 $X2=0
+ $Y2=0
cc_986 N_VPWR_c_1504_n N_A_70_74#_c_1659_n 0.00879331f $X=1.435 $Y=3.19 $X2=0
+ $Y2=0
cc_987 N_VPWR_c_1507_n N_A_70_74#_c_1659_n 0.0114836f $X=2.945 $Y=3.33 $X2=0
+ $Y2=0
cc_988 N_VPWR_c_1491_n N_A_70_74#_c_1659_n 0.00623473f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_989 N_VPWR_c_1497_n N_Q_N_c_1793_n 0.0397608f $X=10.53 $Y=2.375 $X2=0 $Y2=0
cc_990 N_VPWR_c_1498_n N_Q_N_c_1793_n 0.0056634f $X=11.265 $Y=3.33 $X2=0 $Y2=0
cc_991 N_VPWR_c_1499_n N_Q_N_c_1793_n 0.0756134f $X=11.43 $Y=1.905 $X2=0 $Y2=0
cc_992 N_VPWR_c_1491_n N_Q_N_c_1793_n 0.00589694f $X=13.68 $Y=3.33 $X2=0 $Y2=0
cc_993 N_VPWR_c_1499_n Q_N 0.0257878f $X=11.43 $Y=1.905 $X2=0 $Y2=0
cc_994 N_VPWR_c_1500_n N_Q_c_1823_n 0.0450694f $X=12.64 $Y=1.985 $X2=0 $Y2=0
cc_995 N_VPWR_c_1502_n N_Q_c_1823_n 0.0450694f $X=13.64 $Y=1.985 $X2=0 $Y2=0
cc_996 N_VPWR_c_1510_n N_Q_c_1824_n 0.014552f $X=13.475 $Y=3.33 $X2=0 $Y2=0
cc_997 N_VPWR_c_1491_n N_Q_c_1824_n 0.0119791f $X=13.68 $Y=3.33 $X2=0 $Y2=0
cc_998 N_A_70_74#_c_1650_n A_683_485# 3.02954e-19 $X=3.365 $Y=2.37 $X2=-0.19
+ $Y2=-0.245
cc_999 N_A_70_74#_c_1652_n A_683_485# 0.00394048f $X=3.45 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_1000 N_A_70_74#_c_1639_n A_156_74# 0.00289231f $X=0.685 $Y=0.515 $X2=-0.19
+ $Y2=-0.245
cc_1001 N_A_70_74#_c_1642_n A_156_74# 0.00154524f $X=0.845 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_1002 N_A_70_74#_c_1639_n N_VGND_c_1851_n 0.0134245f $X=0.685 $Y=0.515 $X2=0
+ $Y2=0
cc_1003 N_A_70_74#_c_1642_n N_VGND_c_1851_n 0.00833316f $X=0.845 $Y=1.95 $X2=0
+ $Y2=0
cc_1004 N_A_70_74#_c_1639_n N_VGND_c_1868_n 0.0167633f $X=0.685 $Y=0.515 $X2=0
+ $Y2=0
cc_1005 N_A_70_74#_c_1639_n N_VGND_c_1875_n 0.0179018f $X=0.685 $Y=0.515 $X2=0
+ $Y2=0
cc_1006 N_A_70_74#_c_1641_n N_A_614_81#_M1035_d 0.00447556f $X=4.39 $Y=2.41
+ $X2=0 $Y2=0
cc_1007 N_A_70_74#_c_1640_n N_A_614_81#_c_2000_n 0.0576187f $X=4.305 $Y=1.02
+ $X2=0 $Y2=0
cc_1008 N_A_70_74#_c_1643_n N_A_614_81#_c_2000_n 0.0300095f $X=3.53 $Y=1.02
+ $X2=0 $Y2=0
cc_1009 N_A_70_74#_c_1640_n N_A_614_81#_c_2001_n 0.0147455f $X=4.305 $Y=1.02
+ $X2=0 $Y2=0
cc_1010 N_A_70_74#_c_1641_n N_A_614_81#_c_2001_n 0.0371597f $X=4.39 $Y=2.41
+ $X2=0 $Y2=0
cc_1011 Q_N N_VGND_M1036_d 0.00584895f $X=11.675 $Y=0.84 $X2=0 $Y2=0
cc_1012 N_Q_N_c_1791_n N_VGND_c_1855_n 0.0151654f $X=11.36 $Y=0.515 $X2=0 $Y2=0
cc_1013 Q_N N_VGND_c_1855_n 0.00847611f $X=11.675 $Y=0.84 $X2=0 $Y2=0
cc_1014 N_Q_N_c_1791_n N_VGND_c_1856_n 0.010186f $X=11.36 $Y=0.515 $X2=0 $Y2=0
cc_1015 Q_N N_VGND_c_1856_n 0.0165497f $X=11.675 $Y=0.84 $X2=0 $Y2=0
cc_1016 N_Q_N_c_1791_n N_VGND_c_1869_n 0.0114405f $X=11.36 $Y=0.515 $X2=0 $Y2=0
cc_1017 N_Q_N_c_1791_n N_VGND_c_1875_n 0.00941304f $X=11.36 $Y=0.515 $X2=0 $Y2=0
cc_1018 Q_N N_VGND_c_1875_n 0.00714657f $X=11.675 $Y=0.84 $X2=0 $Y2=0
cc_1019 N_Q_c_1822_n N_VGND_c_1857_n 0.0308594f $X=13.225 $Y=0.495 $X2=0 $Y2=0
cc_1020 N_Q_c_1822_n N_VGND_c_1859_n 0.0323079f $X=13.225 $Y=0.495 $X2=0 $Y2=0
cc_1021 N_Q_c_1822_n N_VGND_c_1871_n 0.0157615f $X=13.225 $Y=0.495 $X2=0 $Y2=0
cc_1022 N_Q_c_1822_n N_VGND_c_1875_n 0.0120285f $X=13.225 $Y=0.495 $X2=0 $Y2=0
cc_1023 N_VGND_c_1864_n N_A_1499_149#_c_2025_n 0.0040788f $X=9.415 $Y=0 $X2=0
+ $Y2=0
cc_1024 N_VGND_c_1875_n N_A_1499_149#_c_2025_n 0.00820175f $X=13.68 $Y=0 $X2=0
+ $Y2=0
cc_1025 N_VGND_c_1854_n N_A_1499_149#_c_2027_n 0.0139893f $X=9.58 $Y=0.555 $X2=0
+ $Y2=0
cc_1026 N_VGND_c_1864_n N_A_1499_149#_c_2027_n 0.0106808f $X=9.415 $Y=0 $X2=0
+ $Y2=0
cc_1027 N_VGND_c_1875_n N_A_1499_149#_c_2027_n 0.00901185f $X=13.68 $Y=0 $X2=0
+ $Y2=0
