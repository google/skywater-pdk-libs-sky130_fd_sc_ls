* NGSPICE file created from sky130_fd_sc_ls__o41a_1.ext - technology: sky130A

.subckt sky130_fd_sc_ls__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
M1000 VPWR A1 a_641_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=1.4016e+12p pd=7.2e+06u as=4.704e+11p ps=3.08e+06u
M1001 a_527_368# A3 a_443_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=4.704e+11p pd=3.08e+06u as=3.024e+11p ps=2.78e+06u
M1002 a_83_270# B1 VPWR VPB phighvt w=840000u l=150000u
+  ad=4.0165e+11p pd=3.01e+06u as=0p ps=0u
M1003 a_641_368# A2 a_527_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND A4 a_326_74# VNB nshort w=640000u l=150000u
+  ad=8.899e+11p pd=6.71e+06u as=6.24e+11p ps=5.79e+06u
M1005 a_326_74# B1 a_83_270# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1006 VPWR a_83_270# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.304e+11p ps=2.83e+06u
M1007 a_443_368# A4 a_83_270# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND A2 a_326_74# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_326_74# A1 VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND a_83_270# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1011 a_326_74# A3 VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

