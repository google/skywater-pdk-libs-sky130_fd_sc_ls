* NGSPICE file created from sky130_fd_sc_ls__a311oi_4.ext - technology: sky130A

.subckt sky130_fd_sc_ls__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
M1000 a_114_368# A3 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=2.688e+12p pd=2.272e+07u as=2.296e+12p ps=1.978e+07u
M1001 a_114_368# B1 a_1213_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=1.6464e+12p ps=1.414e+07u
M1002 a_465_74# A2 a_34_74# VNB nshort w=740000u l=150000u
+  ad=8.288e+11p pd=8.16e+06u as=1.0286e+12p ps=1.018e+07u
M1003 VGND A3 a_34_74# VNB nshort w=740000u l=150000u
+  ad=1.4578e+12p pd=9.86e+06u as=0p ps=0u
M1004 Y C1 VGND VNB nshort w=740000u l=150000u
+  ad=1.0286e+12p pd=1.018e+07u as=0p ps=0u
M1005 VPWR A2 a_114_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR A1 a_114_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_465_74# A1 Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR A3 a_114_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_1213_368# B1 a_114_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND B1 Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_34_74# A2 a_465_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Y A1 a_465_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_114_368# A1 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_114_368# A1 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y C1 a_1213_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=6.72e+11p pd=5.68e+06u as=0p ps=0u
M1016 a_114_368# A2 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR A1 a_114_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND A3 a_34_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 Y B1 VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_114_368# B1 a_1213_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_465_74# A1 Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_1213_368# C1 Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_34_74# A3 VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VPWR A2 a_114_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_1213_368# C1 Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_34_74# A3 VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_1213_368# B1 a_114_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_114_368# A3 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPWR A3 a_114_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VGND C1 Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_114_368# A2 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 Y C1 a_1213_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_465_74# A2 a_34_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_34_74# A2 a_465_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 Y A1 a_465_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

