* File: sky130_fd_sc_ls__einvn_1.spice
* Created: Fri Aug 28 13:23:26 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__einvn_1.pex.spice"
.subckt sky130_fd_sc_ls__einvn_1  VNB VPB TE_B A VPWR Z VGND
* 
* VGND	VGND
* Z	Z
* VPWR	VPWR
* A	A
* TE_B	TE_B
* VPB	VPB
* VNB	VNB
MM1004 N_VGND_M1004_d N_TE_B_M1004_g N_A_22_46#_M1004_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0928345 AS=0.1218 PD=0.854483 PS=1.42 NRD=22.848 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.9 A=0.063 P=1.14 MULT=1
MM1000 A_281_100# N_A_22_46#_M1000_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.74
+ AD=0.0888 AS=0.163566 PD=0.98 PS=1.50552 NRD=10.536 NRS=0 M=1 R=4.93333
+ SA=75000.4 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1002 N_Z_M1002_d N_A_M1002_g A_281_100# VNB NSHORT L=0.15 W=0.74 AD=0.2109
+ AS=0.0888 PD=2.05 PS=0.98 NRD=0 NRS=10.536 M=1 R=4.93333 SA=75000.8 SB=75000.2
+ A=0.111 P=1.78 MULT=1
MM1005 N_VPWR_M1005_d N_TE_B_M1005_g N_A_22_46#_M1005_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.141091 AS=0.1888 PD=1.09455 PS=1.87 NRD=29.2348 NRS=3.0732 M=1
+ R=4.26667 SA=75000.2 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1003 A_278_368# N_TE_B_M1003_g N_VPWR_M1005_d VPB PHIGHVT L=0.15 W=1.12
+ AD=0.1512 AS=0.246909 PD=1.39 PS=1.91545 NRD=14.0658 NRS=1.7533 M=1 R=7.46667
+ SA=75000.5 SB=75000.6 A=0.168 P=2.54 MULT=1
MM1001 N_Z_M1001_d N_A_M1001_g A_278_368# VPB PHIGHVT L=0.15 W=1.12 AD=0.3304
+ AS=0.1512 PD=2.83 PS=1.39 NRD=1.7533 NRS=14.0658 M=1 R=7.46667 SA=75000.9
+ SB=75000.2 A=0.168 P=2.54 MULT=1
DX6_noxref VNB VPB NWDIODE A=5.1708 P=9.28
c_24 VNB 0 9.55478e-20 $X=0 $Y=0
*
.include "sky130_fd_sc_ls__einvn_1.pxi.spice"
*
.ends
*
*
