* File: sky130_fd_sc_ls__xnor2_1.spice
* Created: Fri Aug 28 14:08:39 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__xnor2_1.pex.spice"
.subckt sky130_fd_sc_ls__xnor2_1  VNB VPB B A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* B	B
* VPB	VPB
* VNB	VNB
MM1006 A_112_119# N_A_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.64 AD=0.0672
+ AS=0.176 PD=0.85 PS=1.83 NRD=9.372 NRS=0 M=1 R=4.26667 SA=75000.2 SB=75000.6
+ A=0.096 P=1.58 MULT=1
MM1002 N_A_138_385#_M1002_d N_B_M1002_g A_112_119# VNB NSHORT L=0.15 W=0.64
+ AD=0.176 AS=0.0672 PD=1.83 PS=0.85 NRD=0 NRS=9.372 M=1 R=4.26667 SA=75000.6
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1009 N_VGND_M1009_d N_A_M1009_g N_A_293_74#_M1009_s VNB NSHORT L=0.15 W=0.74
+ AD=0.182 AS=0.2035 PD=1.345 PS=2.03 NRD=12.156 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.2 A=0.111 P=1.78 MULT=1
MM1008 N_A_293_74#_M1008_d N_B_M1008_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.182 PD=1.02 PS=1.345 NRD=0 NRS=12.972 M=1 R=4.93333 SA=75000.8
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1003 N_Y_M1003_d N_A_138_385#_M1003_g N_A_293_74#_M1008_d VNB NSHORT L=0.15
+ W=0.74 AD=0.2294 AS=0.1036 PD=2.1 PS=1.02 NRD=4.044 NRS=0 M=1 R=4.93333
+ SA=75001.2 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1004 N_A_138_385#_M1004_d N_A_M1004_g N_VPWR_M1004_s VPB PHIGHVT L=0.15 W=0.84
+ AD=0.126 AS=0.2898 PD=1.14 PS=2.37 NRD=2.3443 NRS=14.0658 M=1 R=5.6 SA=75000.3
+ SB=75002.4 A=0.126 P=1.98 MULT=1
MM1001 N_VPWR_M1001_d N_B_M1001_g N_A_138_385#_M1004_d VPB PHIGHVT L=0.15 W=0.84
+ AD=0.246707 AS=0.126 PD=1.46571 PS=1.14 NRD=154.783 NRS=0 M=1 R=5.6 SA=75000.7
+ SB=75001.9 A=0.126 P=1.98 MULT=1
MM1000 A_376_368# N_A_M1000_g N_VPWR_M1001_d VPB PHIGHVT L=0.15 W=1.12 AD=0.1512
+ AS=0.328943 PD=1.39 PS=1.95429 NRD=14.0658 NRS=1.7533 M=1 R=7.46667 SA=75001.1
+ SB=75001.2 A=0.168 P=2.54 MULT=1
MM1007 N_Y_M1007_d N_B_M1007_g A_376_368# VPB PHIGHVT L=0.15 W=1.12 AD=0.2352
+ AS=0.1512 PD=1.54 PS=1.39 NRD=14.0658 NRS=14.0658 M=1 R=7.46667 SA=75001.6
+ SB=75000.8 A=0.168 P=2.54 MULT=1
MM1005 N_VPWR_M1005_d N_A_138_385#_M1005_g N_Y_M1007_d VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.2352 PD=2.83 PS=1.54 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75002.1 SB=75000.2 A=0.168 P=2.54 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9564 P=11.2
*
.include "sky130_fd_sc_ls__xnor2_1.pxi.spice"
*
.ends
*
*
