* File: sky130_fd_sc_ls__dlrbp_2.spice
* Created: Fri Aug 28 13:18:19 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__dlrbp_2.pex.spice"
.subckt sky130_fd_sc_ls__dlrbp_2  VNB VPB D GATE RESET_B VPWR Q Q_N VGND
* 
* VGND	VGND
* Q_N	Q_N
* Q	Q
* VPWR	VPWR
* RESET_B	RESET_B
* GATE	GATE
* D	D
* VPB	VPB
* VNB	VNB
MM1012 N_VGND_M1012_d N_D_M1012_g N_A_27_112#_M1012_s VNB NSHORT L=0.15 W=0.55
+ AD=0.129591 AS=0.15675 PD=0.997674 PS=1.67 NRD=18 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75000.8 A=0.0825 P=1.4 MULT=1
MM1009 N_A_230_74#_M1009_d N_GATE_M1009_g N_VGND_M1012_d VNB NSHORT L=0.15
+ W=0.74 AD=0.2109 AS=0.174359 PD=2.05 PS=1.34233 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75000.7 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1000 N_VGND_M1000_d N_A_230_74#_M1000_g N_A_363_82#_M1000_s VNB NSHORT L=0.15
+ W=0.74 AD=0.201864 AS=0.2109 PD=1.51754 PS=2.05 NRD=35.316 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001.6 A=0.111 P=1.78 MULT=1
MM1002 A_569_80# N_A_27_112#_M1002_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.64
+ AD=0.0672 AS=0.174586 PD=0.85 PS=1.31246 NRD=9.372 NRS=16.872 M=1 R=4.26667
+ SA=75000.8 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1022 N_A_641_80#_M1022_d N_A_363_82#_M1022_g A_569_80# VNB NSHORT L=0.15
+ W=0.64 AD=0.162536 AS=0.0672 PD=1.38868 PS=0.85 NRD=21.552 NRS=9.372 M=1
+ R=4.26667 SA=75001.2 SB=75000.9 A=0.096 P=1.58 MULT=1
MM1001 A_773_124# N_A_230_74#_M1001_g N_A_641_80#_M1022_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.106664 PD=0.66 PS=0.911321 NRD=18.564 NRS=32.856 M=1
+ R=2.8 SA=75001.8 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1017 N_VGND_M1017_d N_A_821_98#_M1017_g A_773_124# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75002.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1013 A_1049_74# N_A_641_80#_M1013_g N_A_821_98#_M1013_s VNB NSHORT L=0.15
+ W=0.74 AD=0.0888 AS=0.2109 PD=0.98 PS=2.05 NRD=10.536 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001.6 A=0.111 P=1.78 MULT=1
MM1006 N_VGND_M1006_d N_RESET_B_M1006_g A_1049_74# VNB NSHORT L=0.15 W=0.74
+ AD=0.1443 AS=0.0888 PD=1.13 PS=0.98 NRD=0 NRS=10.536 M=1 R=4.93333 SA=75000.6
+ SB=75001.2 A=0.111 P=1.78 MULT=1
MM1023 N_Q_M1023_d N_A_821_98#_M1023_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1443 PD=1.02 PS=1.13 NRD=0 NRS=17.832 M=1 R=4.93333 SA=75001.1
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1024 N_Q_M1023_d N_A_821_98#_M1024_g N_VGND_M1024_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.2627 PD=1.02 PS=2.19 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.6
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1004 N_VGND_M1004_d N_A_821_98#_M1004_g N_A_1449_368#_M1004_s VNB NSHORT
+ L=0.15 W=0.64 AD=0.136255 AS=0.1824 PD=1.07594 PS=1.85 NRD=13.116 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1007 N_Q_N_M1007_d N_A_1449_368#_M1007_g N_VGND_M1004_d VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.157545 PD=1.02 PS=1.24406 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75000.7 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1014 N_Q_N_M1007_d N_A_1449_368#_M1014_g N_VGND_M1014_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.1 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1019 N_VPWR_M1019_d N_D_M1019_g N_A_27_112#_M1019_s VPB PHIGHVT L=0.15 W=0.84
+ AD=0.22785 AS=0.2478 PD=1.52 PS=2.27 NRD=50.7078 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.9 A=0.126 P=1.98 MULT=1
MM1015 N_A_230_74#_M1015_d N_GATE_M1015_g N_VPWR_M1019_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.2898 AS=0.22785 PD=2.37 PS=1.52 NRD=0 NRS=50.7078 M=1 R=5.6
+ SA=75000.8 SB=75000.3 A=0.126 P=1.98 MULT=1
MM1025 N_VPWR_M1025_d N_A_230_74#_M1025_g N_A_363_82#_M1025_s VPB PHIGHVT L=0.15
+ W=0.84 AD=0.185165 AS=0.2478 PD=1.29652 PS=2.27 NRD=26.9693 NRS=2.3443 M=1
+ R=5.6 SA=75000.2 SB=75002.3 A=0.126 P=1.98 MULT=1
MM1016 A_566_392# N_A_27_112#_M1016_g N_VPWR_M1025_d VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.220435 PD=1.27 PS=1.54348 NRD=15.7403 NRS=5.8903 M=1 R=6.66667
+ SA=75000.7 SB=75002.1 A=0.15 P=2.3 MULT=1
MM1010 N_A_641_80#_M1010_d N_A_230_74#_M1010_g A_566_392# VPB PHIGHVT L=0.15 W=1
+ AD=0.234366 AS=0.135 PD=1.9507 PS=1.27 NRD=1.9503 NRS=15.7403 M=1 R=6.66667
+ SA=75001.1 SB=75001.7 A=0.15 P=2.3 MULT=1
MM1020 A_757_508# N_A_363_82#_M1020_g N_A_641_80#_M1010_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.10605 AS=0.0984338 PD=0.925 PS=0.819296 NRD=92.6294 NRS=46.886 M=1
+ R=2.8 SA=75001.5 SB=75003.1 A=0.063 P=1.14 MULT=1
MM1021 N_VPWR_M1021_d N_A_821_98#_M1021_g A_757_508# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.120464 AS=0.10605 PD=0.943636 PS=0.925 NRD=77.3816 NRS=92.6294 M=1 R=2.8
+ SA=75002.2 SB=75002.5 A=0.063 P=1.14 MULT=1
MM1027 N_A_821_98#_M1027_d N_A_641_80#_M1027_g N_VPWR_M1021_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.196 AS=0.321236 PD=1.47 PS=2.51636 NRD=10.5395 NRS=29.0181 M=1
+ R=7.46667 SA=75001.2 SB=75001.7 A=0.168 P=2.54 MULT=1
MM1005 N_VPWR_M1005_d N_RESET_B_M1005_g N_A_821_98#_M1027_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.2128 AS=0.196 PD=1.5 PS=1.47 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75001.7 SB=75001.2 A=0.168 P=2.54 MULT=1
MM1003 N_VPWR_M1005_d N_A_821_98#_M1003_g N_Q_M1003_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.2128 AS=0.168 PD=1.5 PS=1.42 NRD=7.0329 NRS=1.7533 M=1 R=7.46667
+ SA=75002.3 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1026 N_VPWR_M1026_d N_A_821_98#_M1026_g N_Q_M1003_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.7 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1008 N_VPWR_M1008_d N_A_821_98#_M1008_g N_A_1449_368#_M1008_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.203679 AS=0.295 PD=1.43396 PS=2.59 NRD=11.8003 NRS=1.9503 M=1
+ R=6.66667 SA=75000.2 SB=75001.2 A=0.15 P=2.3 MULT=1
MM1011 N_Q_N_M1011_d N_A_1449_368#_M1011_g N_VPWR_M1008_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.228121 PD=1.42 PS=1.60604 NRD=1.7533 NRS=10.5395 M=1
+ R=7.46667 SA=75000.7 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1018 N_Q_N_M1011_d N_A_1449_368#_M1018_g N_VPWR_M1018_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.2 SB=75000.2 A=0.168 P=2.54 MULT=1
DX28_noxref VNB VPB NWDIODE A=17.67 P=22.72
*
.include "sky130_fd_sc_ls__dlrbp_2.pxi.spice"
*
.ends
*
*
