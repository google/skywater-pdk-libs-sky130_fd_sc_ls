* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__dlrbn_1 D GATE_N RESET_B VGND VNB VPB VPWR Q Q_N
X0 a_1133_74# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X1 VPWR a_1437_112# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X2 a_373_74# a_231_74# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X3 VPWR a_889_92# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X4 a_608_74# a_231_74# a_686_74# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X5 a_611_392# a_373_74# a_686_74# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 a_1437_112# a_889_92# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X7 VPWR GATE_N a_231_74# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X8 VGND a_889_92# Q VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X9 a_686_74# a_231_74# a_802_508# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X10 a_889_92# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X11 VPWR a_27_424# a_611_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 a_686_74# a_373_74# a_841_118# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 VGND a_27_424# a_608_74# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X14 a_841_118# a_889_92# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 a_27_424# D VGND VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X16 a_27_424# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X17 a_802_508# a_889_92# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X18 a_1437_112# a_889_92# VGND VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X19 VPWR a_686_74# a_889_92# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X20 VGND GATE_N a_231_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X21 a_889_92# a_686_74# a_1133_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X22 a_373_74# a_231_74# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X23 VGND a_1437_112# Q_N VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
.ends
