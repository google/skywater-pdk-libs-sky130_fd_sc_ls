* NGSPICE file created from sky130_fd_sc_ls__sdlclkp_4.ext - technology: sky130A

.subckt sky130_fd_sc_ls__sdlclkp_4 CLK GATE SCE VGND VNB VPB VPWR GCLK
M1000 a_792_48# a_634_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=2.6355e+12p ps=1.988e+07u
M1001 VGND a_1289_368# GCLK VNB nshort w=740000u l=150000u
+  ad=1.98545e+12p pd=1.63e+07u as=4.514e+11p ps=4.18e+06u
M1002 a_354_105# a_324_79# VPWR VPB phighvt w=840000u l=150000u
+  ad=4.033e+11p pd=3.02e+06u as=0p ps=0u
M1003 GCLK a_1289_368# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=8.68e+11p pd=6.03e+06u as=0p ps=0u
M1004 a_792_48# a_634_74# VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1005 VGND a_792_48# a_744_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1006 VPWR a_792_48# a_785_455# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1007 a_1292_74# CLK VGND VNB nshort w=740000u l=150000u
+  ad=1.776e+11p pd=1.96e+06u as=0p ps=0u
M1008 a_1289_368# a_792_48# a_1292_74# VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1009 a_116_395# SCE VPWR VPB phighvt w=840000u l=150000u
+  ad=2.268e+11p pd=2.22e+06u as=0p ps=0u
M1010 VPWR a_1289_368# GCLK VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND CLK a_324_79# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1012 a_785_455# a_324_79# a_634_74# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=2.856e+11p ps=2.45e+06u
M1013 GCLK a_1289_368# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_634_74# a_354_105# a_119_143# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=4.956e+11p ps=4.54e+06u
M1015 a_1289_368# CLK VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=5.544e+11p pd=3.23e+06u as=0p ps=0u
M1016 a_744_74# a_354_105# a_634_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=2.1025e+11p ps=1.9e+06u
M1017 a_354_105# a_324_79# VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1018 VPWR a_792_48# a_1289_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_119_143# SCE VGND VNB nshort w=550000u l=150000u
+  ad=5.61e+11p pd=4.24e+06u as=0p ps=0u
M1020 a_119_143# GATE a_116_395# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPWR a_1289_368# GCLK VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_634_74# a_324_79# a_119_143# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VPWR CLK a_324_79# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=2.52e+11p ps=2.28e+06u
M1024 GCLK a_1289_368# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VGND GATE a_119_143# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 GCLK a_1289_368# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VGND a_1289_368# GCLK VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

