* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__ebufn_4 A TE_B VGND VNB VPB VPWR Z
X0 VPWR TE_B a_348_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X1 VPWR TE_B a_348_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X2 a_378_74# a_208_74# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X3 a_348_368# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X4 a_27_368# A VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X5 VPWR TE_B a_208_74# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X6 a_348_368# a_27_368# Z VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X7 Z a_27_368# a_378_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X8 a_348_368# a_27_368# Z VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X9 a_27_368# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X10 Z a_27_368# a_348_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X11 a_348_368# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X12 VGND a_208_74# a_378_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X13 a_378_74# a_208_74# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X14 VGND TE_B a_208_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X15 VGND a_208_74# a_378_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X16 a_378_74# a_27_368# Z VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X17 Z a_27_368# a_348_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X18 Z a_27_368# a_378_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X19 a_378_74# a_27_368# Z VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
.ends
