# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ls__ha_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ls__ha_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.08000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.936000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.455000 1.315000 1.785000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.936000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 1.455000 2.275000 1.785000 ;
    END
  END B
  PIN COUT
    ANTENNADIFFAREA  1.265600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.220000 1.820000 7.555000 2.150000 ;
        RECT 6.350000 0.350000 6.600000 0.880000 ;
        RECT 6.350000 0.880000 7.555000 1.130000 ;
        RECT 7.210000 1.130000 7.555000 1.820000 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  1.470100 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 8.735000 1.920000 9.025000 1.965000 ;
        RECT 8.735000 1.965000 9.985000 2.105000 ;
        RECT 8.735000 2.105000 9.025000 2.150000 ;
        RECT 9.695000 1.920000 9.985000 1.965000 ;
        RECT 9.695000 2.105000 9.985000 2.150000 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.080000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 10.080000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.080000 0.085000 ;
      RECT 0.000000  3.245000 10.080000 3.415000 ;
      RECT 0.105000  1.955000  1.255000 2.125000 ;
      RECT 0.105000  2.125000  0.385000 2.965000 ;
      RECT 0.115000  0.605000  0.365000 1.115000 ;
      RECT 0.115000  1.115000  2.170000 1.285000 ;
      RECT 0.545000  0.085000  0.795000 0.945000 ;
      RECT 0.555000  2.295000  0.805000 3.245000 ;
      RECT 0.980000  0.605000  1.230000 1.115000 ;
      RECT 1.005000  2.125000  1.255000 2.905000 ;
      RECT 1.005000  2.905000  2.235000 3.075000 ;
      RECT 1.410000  0.085000  1.660000 0.945000 ;
      RECT 1.455000  1.955000  3.255000 2.125000 ;
      RECT 1.455000  2.125000  1.735000 2.735000 ;
      RECT 1.840000  0.265000  3.170000 0.435000 ;
      RECT 1.840000  0.435000  2.170000 1.115000 ;
      RECT 1.905000  2.295000  2.235000 2.905000 ;
      RECT 2.340000  0.605000  2.670000 1.285000 ;
      RECT 2.475000  2.405000  2.805000 3.245000 ;
      RECT 2.500000  1.285000  2.670000 1.905000 ;
      RECT 2.500000  1.905000  3.255000 1.955000 ;
      RECT 2.840000  0.435000  3.170000 1.235000 ;
      RECT 2.925000  2.125000  3.255000 2.165000 ;
      RECT 2.925000  2.165000  4.070000 2.235000 ;
      RECT 3.075000  1.405000  4.280000 1.575000 ;
      RECT 3.075000  1.575000  4.070000 1.735000 ;
      RECT 3.085000  2.235000  4.070000 2.320000 ;
      RECT 3.085000  2.320000  7.895000 2.335000 ;
      RECT 3.375000  2.505000  3.705000 3.245000 ;
      RECT 3.520000  0.315000  4.780000 0.485000 ;
      RECT 3.520000  0.485000  3.780000 1.235000 ;
      RECT 3.900000  1.735000  4.070000 1.745000 ;
      RECT 3.900000  1.745000  4.230000 1.820000 ;
      RECT 3.900000  1.820000  6.050000 1.995000 ;
      RECT 3.900000  2.335000  7.895000 2.490000 ;
      RECT 3.950000  0.655000  4.280000 1.405000 ;
      RECT 4.430000  2.660000  4.760000 3.245000 ;
      RECT 4.450000  0.485000  4.780000 1.425000 ;
      RECT 4.450000  1.425000  5.710000 1.595000 ;
      RECT 4.950000  0.085000  5.280000 1.255000 ;
      RECT 4.955000  1.995000  6.050000 2.150000 ;
      RECT 5.460000  0.575000  5.710000 1.425000 ;
      RECT 5.490000  2.660000  5.945000 3.245000 ;
      RECT 5.880000  1.320000  6.955000 1.650000 ;
      RECT 5.880000  1.650000  6.050000 1.820000 ;
      RECT 5.920000  0.085000  6.170000 1.130000 ;
      RECT 6.675000  2.660000  7.005000 3.245000 ;
      RECT 6.780000  0.085000  7.110000 0.710000 ;
      RECT 7.575000  2.660000  7.905000 3.245000 ;
      RECT 7.640000  0.085000  7.970000 0.710000 ;
      RECT 7.725000  1.320000  9.645000 1.650000 ;
      RECT 7.725000  1.650000  7.895000 2.320000 ;
      RECT 8.075000  1.820000  9.995000 2.150000 ;
      RECT 8.075000  2.150000  8.305000 2.980000 ;
      RECT 8.150000  0.350000  8.400000 0.980000 ;
      RECT 8.150000  0.980000  9.995000 1.150000 ;
      RECT 8.475000  2.320000  8.805000 3.245000 ;
      RECT 8.570000  0.085000  8.900000 0.810000 ;
      RECT 9.070000  0.350000  9.400000 0.980000 ;
      RECT 9.075000  2.150000  9.405000 2.980000 ;
      RECT 9.580000  0.085000  9.885000 0.810000 ;
      RECT 9.635000  2.320000  9.965000 3.245000 ;
      RECT 9.825000  1.150000  9.995000 1.820000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  1.950000 8.965000 2.120000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
      RECT 9.275000 -0.085000 9.445000 0.085000 ;
      RECT 9.275000  3.245000 9.445000 3.415000 ;
      RECT 9.755000 -0.085000 9.925000 0.085000 ;
      RECT 9.755000  1.950000 9.925000 2.120000 ;
      RECT 9.755000  3.245000 9.925000 3.415000 ;
  END
END sky130_fd_sc_ls__ha_4
END LIBRARY
