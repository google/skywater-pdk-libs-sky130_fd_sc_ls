* File: sky130_fd_sc_ls__a211oi_1.pxi.spice
* Created: Fri Aug 28 12:49:29 2020
* 
x_PM_SKY130_FD_SC_LS__A211OI_1%A2 N_A2_c_48_n N_A2_M1005_g N_A2_M1003_g A2
+ N_A2_c_50_n PM_SKY130_FD_SC_LS__A211OI_1%A2
x_PM_SKY130_FD_SC_LS__A211OI_1%A1 N_A1_M1001_g N_A1_c_75_n N_A1_M1000_g A1
+ N_A1_c_76_n PM_SKY130_FD_SC_LS__A211OI_1%A1
x_PM_SKY130_FD_SC_LS__A211OI_1%B1 N_B1_M1004_g N_B1_c_107_n N_B1_M1002_g B1
+ N_B1_c_108_n PM_SKY130_FD_SC_LS__A211OI_1%B1
x_PM_SKY130_FD_SC_LS__A211OI_1%C1 N_C1_M1007_g N_C1_c_140_n N_C1_M1006_g
+ N_C1_c_136_n N_C1_c_137_n C1 N_C1_c_139_n PM_SKY130_FD_SC_LS__A211OI_1%C1
x_PM_SKY130_FD_SC_LS__A211OI_1%A_71_368# N_A_71_368#_M1005_s N_A_71_368#_M1000_d
+ N_A_71_368#_c_165_n N_A_71_368#_c_166_n N_A_71_368#_c_171_n
+ N_A_71_368#_c_177_n N_A_71_368#_c_167_n PM_SKY130_FD_SC_LS__A211OI_1%A_71_368#
x_PM_SKY130_FD_SC_LS__A211OI_1%VPWR N_VPWR_M1005_d N_VPWR_c_194_n N_VPWR_c_195_n
+ N_VPWR_c_196_n VPWR N_VPWR_c_197_n N_VPWR_c_193_n
+ PM_SKY130_FD_SC_LS__A211OI_1%VPWR
x_PM_SKY130_FD_SC_LS__A211OI_1%Y N_Y_M1001_d N_Y_M1007_d N_Y_M1006_d N_Y_c_219_n
+ N_Y_c_220_n N_Y_c_225_n N_Y_c_221_n N_Y_c_226_n N_Y_c_222_n Y Y Y N_Y_c_224_n
+ PM_SKY130_FD_SC_LS__A211OI_1%Y
x_PM_SKY130_FD_SC_LS__A211OI_1%VGND N_VGND_M1003_s N_VGND_M1004_d N_VGND_c_270_n
+ N_VGND_c_271_n N_VGND_c_272_n N_VGND_c_273_n VGND N_VGND_c_274_n
+ N_VGND_c_275_n N_VGND_c_276_n N_VGND_c_277_n PM_SKY130_FD_SC_LS__A211OI_1%VGND
cc_1 VNB N_A2_c_48_n 0.034949f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=1.765
cc_2 VNB N_A2_M1003_g 0.03136f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=0.74
cc_3 VNB N_A2_c_50_n 0.0052161f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.515
cc_4 VNB N_A1_M1001_g 0.0248902f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=2.4
cc_5 VNB N_A1_c_75_n 0.0262515f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=0.74
cc_6 VNB N_A1_c_76_n 0.00166449f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.515
cc_7 VNB N_B1_M1004_g 0.0261208f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=2.4
cc_8 VNB N_B1_c_107_n 0.0262555f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=0.74
cc_9 VNB N_B1_c_108_n 0.00166777f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.515
cc_10 VNB N_C1_c_136_n 0.0198581f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_11 VNB N_C1_c_137_n 0.0234756f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB C1 0.0207309f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.515
cc_13 VNB N_C1_c_139_n 0.0638365f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.515
cc_14 VNB N_VPWR_c_193_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_Y_c_219_n 0.00792442f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.515
cc_16 VNB N_Y_c_220_n 0.00317771f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.515
cc_17 VNB N_Y_c_221_n 0.0204378f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_Y_c_222_n 0.00374926f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB Y 0.0086849f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_Y_c_224_n 0.00924258f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_270_n 0.0457851f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_271_n 0.00685406f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.515
cc_23 VNB N_VGND_c_272_n 0.0129628f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_273_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_274_n 0.028216f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_275_n 0.0263115f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_276_n 0.202322f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_277_n 0.0069273f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VPB N_A2_c_48_n 0.0342348f $X=-0.19 $Y=1.66 $X2=0.705 $Y2=1.765
cc_30 VPB N_A2_c_50_n 0.00658929f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.515
cc_31 VPB N_A1_c_75_n 0.0277367f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=0.74
cc_32 VPB N_A1_c_76_n 0.00238178f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.515
cc_33 VPB N_B1_c_107_n 0.026708f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=0.74
cc_34 VPB N_B1_c_108_n 0.00597673f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.515
cc_35 VPB N_C1_c_140_n 0.0207394f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.35
cc_36 VPB N_C1_c_136_n 0.00924193f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_37 VPB N_A_71_368#_c_165_n 0.00880428f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_38 VPB N_A_71_368#_c_166_n 0.0360166f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_39 VPB N_A_71_368#_c_167_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0.65 $Y2=1.665
cc_40 VPB N_VPWR_c_194_n 0.00958771f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=0.74
cc_41 VPB N_VPWR_c_195_n 0.0255159f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_42 VPB N_VPWR_c_196_n 0.00612923f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.515
cc_43 VPB N_VPWR_c_197_n 0.0510638f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_44 VPB N_VPWR_c_193_n 0.0835436f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_45 VPB N_Y_c_225_n 0.0401132f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_Y_c_226_n 0.0141934f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB N_Y_c_222_n 0.00115649f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 N_A2_M1003_g N_A1_M1001_g 0.0426951f $X=0.72 $Y=0.74 $X2=0 $Y2=0
cc_49 N_A2_c_48_n N_A1_c_75_n 0.0713555f $X=0.705 $Y=1.765 $X2=0 $Y2=0
cc_50 N_A2_c_50_n N_A1_c_75_n 0.00214941f $X=0.63 $Y=1.515 $X2=0 $Y2=0
cc_51 N_A2_c_48_n N_A1_c_76_n 7.18891e-19 $X=0.705 $Y=1.765 $X2=0 $Y2=0
cc_52 N_A2_c_50_n N_A1_c_76_n 0.0347535f $X=0.63 $Y=1.515 $X2=0 $Y2=0
cc_53 N_A2_c_48_n N_A_71_368#_c_165_n 0.00123808f $X=0.705 $Y=1.765 $X2=0 $Y2=0
cc_54 N_A2_c_50_n N_A_71_368#_c_165_n 0.0131798f $X=0.63 $Y=1.515 $X2=0 $Y2=0
cc_55 N_A2_c_48_n N_A_71_368#_c_166_n 0.0110297f $X=0.705 $Y=1.765 $X2=0 $Y2=0
cc_56 N_A2_c_48_n N_A_71_368#_c_171_n 0.0124019f $X=0.705 $Y=1.765 $X2=0 $Y2=0
cc_57 N_A2_c_50_n N_A_71_368#_c_171_n 0.012218f $X=0.63 $Y=1.515 $X2=0 $Y2=0
cc_58 N_A2_c_48_n N_A_71_368#_c_167_n 5.94528e-19 $X=0.705 $Y=1.765 $X2=0 $Y2=0
cc_59 N_A2_c_48_n N_VPWR_c_194_n 0.0033519f $X=0.705 $Y=1.765 $X2=0 $Y2=0
cc_60 N_A2_c_48_n N_VPWR_c_195_n 0.00445602f $X=0.705 $Y=1.765 $X2=0 $Y2=0
cc_61 N_A2_c_48_n N_VPWR_c_193_n 0.00861742f $X=0.705 $Y=1.765 $X2=0 $Y2=0
cc_62 N_A2_M1003_g N_Y_c_219_n 0.0012054f $X=0.72 $Y=0.74 $X2=0 $Y2=0
cc_63 N_A2_M1003_g N_Y_c_220_n 0.00134279f $X=0.72 $Y=0.74 $X2=0 $Y2=0
cc_64 N_A2_c_48_n N_VGND_c_270_n 0.00137074f $X=0.705 $Y=1.765 $X2=0 $Y2=0
cc_65 N_A2_M1003_g N_VGND_c_270_n 0.0188126f $X=0.72 $Y=0.74 $X2=0 $Y2=0
cc_66 N_A2_c_50_n N_VGND_c_270_n 0.0143146f $X=0.63 $Y=1.515 $X2=0 $Y2=0
cc_67 N_A2_M1003_g N_VGND_c_274_n 0.00383152f $X=0.72 $Y=0.74 $X2=0 $Y2=0
cc_68 N_A2_M1003_g N_VGND_c_276_n 0.0075694f $X=0.72 $Y=0.74 $X2=0 $Y2=0
cc_69 N_A1_M1001_g N_B1_M1004_g 0.0223185f $X=1.08 $Y=0.74 $X2=0 $Y2=0
cc_70 N_A1_c_75_n N_B1_c_107_n 0.0340611f $X=1.245 $Y=1.765 $X2=0 $Y2=0
cc_71 N_A1_c_76_n N_B1_c_107_n 0.00129529f $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_72 N_A1_c_75_n N_B1_c_108_n 0.00171178f $X=1.245 $Y=1.765 $X2=0 $Y2=0
cc_73 N_A1_c_76_n N_B1_c_108_n 0.0277336f $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_74 N_A1_c_75_n N_A_71_368#_c_166_n 6.65743e-19 $X=1.245 $Y=1.765 $X2=0 $Y2=0
cc_75 N_A1_c_75_n N_A_71_368#_c_171_n 0.013127f $X=1.245 $Y=1.765 $X2=0 $Y2=0
cc_76 N_A1_c_76_n N_A_71_368#_c_171_n 0.020911f $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_77 N_A1_c_75_n N_A_71_368#_c_177_n 4.2644e-19 $X=1.245 $Y=1.765 $X2=0 $Y2=0
cc_78 N_A1_c_76_n N_A_71_368#_c_177_n 0.00179688f $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_79 N_A1_c_75_n N_A_71_368#_c_167_n 0.0106384f $X=1.245 $Y=1.765 $X2=0 $Y2=0
cc_80 N_A1_c_75_n N_VPWR_c_194_n 0.00725721f $X=1.245 $Y=1.765 $X2=0 $Y2=0
cc_81 N_A1_c_75_n N_VPWR_c_197_n 0.00445602f $X=1.245 $Y=1.765 $X2=0 $Y2=0
cc_82 N_A1_c_75_n N_VPWR_c_193_n 0.00857833f $X=1.245 $Y=1.765 $X2=0 $Y2=0
cc_83 N_A1_M1001_g N_Y_c_219_n 0.00897846f $X=1.08 $Y=0.74 $X2=0 $Y2=0
cc_84 N_A1_c_75_n N_Y_c_219_n 0.00140176f $X=1.245 $Y=1.765 $X2=0 $Y2=0
cc_85 N_A1_c_76_n N_Y_c_219_n 0.0211742f $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_86 N_A1_M1001_g N_Y_c_220_n 0.0100683f $X=1.08 $Y=0.74 $X2=0 $Y2=0
cc_87 N_A1_M1001_g N_VGND_c_270_n 0.00263599f $X=1.08 $Y=0.74 $X2=0 $Y2=0
cc_88 N_A1_M1001_g N_VGND_c_271_n 5.90483e-19 $X=1.08 $Y=0.74 $X2=0 $Y2=0
cc_89 N_A1_M1001_g N_VGND_c_274_n 0.00383287f $X=1.08 $Y=0.74 $X2=0 $Y2=0
cc_90 N_A1_M1001_g N_VGND_c_276_n 0.00656608f $X=1.08 $Y=0.74 $X2=0 $Y2=0
cc_91 N_B1_c_107_n N_C1_c_140_n 0.0452034f $X=1.695 $Y=1.765 $X2=0 $Y2=0
cc_92 N_B1_c_107_n N_C1_c_136_n 0.0241625f $X=1.695 $Y=1.765 $X2=0 $Y2=0
cc_93 N_B1_c_108_n N_C1_c_136_n 6.55532e-19 $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_94 N_B1_M1004_g N_C1_c_137_n 0.0248511f $X=1.62 $Y=0.74 $X2=0 $Y2=0
cc_95 N_B1_c_107_n N_A_71_368#_c_177_n 0.00298181f $X=1.695 $Y=1.765 $X2=0 $Y2=0
cc_96 N_B1_c_108_n N_A_71_368#_c_177_n 0.00518699f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_97 N_B1_c_107_n N_A_71_368#_c_167_n 0.0134678f $X=1.695 $Y=1.765 $X2=0 $Y2=0
cc_98 N_B1_c_107_n N_VPWR_c_197_n 0.00445602f $X=1.695 $Y=1.765 $X2=0 $Y2=0
cc_99 N_B1_c_107_n N_VPWR_c_193_n 0.00858782f $X=1.695 $Y=1.765 $X2=0 $Y2=0
cc_100 N_B1_M1004_g N_Y_c_220_n 0.0026934f $X=1.62 $Y=0.74 $X2=0 $Y2=0
cc_101 N_B1_M1004_g N_Y_c_221_n 6.39617e-19 $X=1.62 $Y=0.74 $X2=0 $Y2=0
cc_102 N_B1_M1004_g N_Y_c_222_n 0.00296121f $X=1.62 $Y=0.74 $X2=0 $Y2=0
cc_103 N_B1_c_107_n N_Y_c_222_n 0.00687949f $X=1.695 $Y=1.765 $X2=0 $Y2=0
cc_104 N_B1_c_108_n N_Y_c_222_n 0.0327281f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_105 N_B1_M1004_g N_Y_c_224_n 0.0217865f $X=1.62 $Y=0.74 $X2=0 $Y2=0
cc_106 N_B1_c_107_n N_Y_c_224_n 0.00133088f $X=1.695 $Y=1.765 $X2=0 $Y2=0
cc_107 N_B1_c_108_n N_Y_c_224_n 0.0262137f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_108 N_B1_M1004_g N_VGND_c_271_n 0.00776565f $X=1.62 $Y=0.74 $X2=0 $Y2=0
cc_109 N_B1_M1004_g N_VGND_c_274_n 0.00383152f $X=1.62 $Y=0.74 $X2=0 $Y2=0
cc_110 N_B1_M1004_g N_VGND_c_276_n 0.00378707f $X=1.62 $Y=0.74 $X2=0 $Y2=0
cc_111 N_C1_c_140_n N_A_71_368#_c_167_n 8.51602e-19 $X=2.175 $Y=1.765 $X2=0
+ $Y2=0
cc_112 N_C1_c_140_n N_VPWR_c_197_n 0.00291513f $X=2.175 $Y=1.765 $X2=0 $Y2=0
cc_113 N_C1_c_140_n N_VPWR_c_193_n 0.0036375f $X=2.175 $Y=1.765 $X2=0 $Y2=0
cc_114 N_C1_c_140_n N_Y_c_225_n 0.0207265f $X=2.175 $Y=1.765 $X2=0 $Y2=0
cc_115 N_C1_c_137_n N_Y_c_221_n 0.00733151f $X=2.175 $Y=1.22 $X2=0 $Y2=0
cc_116 N_C1_c_140_n N_Y_c_226_n 0.00732878f $X=2.175 $Y=1.765 $X2=0 $Y2=0
cc_117 N_C1_c_136_n N_Y_c_226_n 7.97465e-19 $X=2.265 $Y=1.385 $X2=0 $Y2=0
cc_118 C1 N_Y_c_226_n 0.00712672f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_119 N_C1_c_139_n N_Y_c_226_n 0.00809123f $X=2.61 $Y=1.385 $X2=0 $Y2=0
cc_120 N_C1_c_140_n N_Y_c_222_n 0.002834f $X=2.175 $Y=1.765 $X2=0 $Y2=0
cc_121 N_C1_c_136_n N_Y_c_222_n 0.022335f $X=2.265 $Y=1.385 $X2=0 $Y2=0
cc_122 N_C1_c_137_n N_Y_c_222_n 9.75292e-19 $X=2.175 $Y=1.22 $X2=0 $Y2=0
cc_123 C1 N_Y_c_222_n 0.0208673f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_124 N_C1_c_137_n Y 0.0214366f $X=2.175 $Y=1.22 $X2=0 $Y2=0
cc_125 C1 Y 0.00830742f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_126 N_C1_c_139_n Y 0.00747729f $X=2.61 $Y=1.385 $X2=0 $Y2=0
cc_127 N_C1_c_137_n N_VGND_c_271_n 0.00493436f $X=2.175 $Y=1.22 $X2=0 $Y2=0
cc_128 N_C1_c_137_n N_VGND_c_275_n 0.00434272f $X=2.175 $Y=1.22 $X2=0 $Y2=0
cc_129 N_C1_c_137_n N_VGND_c_276_n 0.00443636f $X=2.175 $Y=1.22 $X2=0 $Y2=0
cc_130 N_A_71_368#_c_171_n N_VPWR_M1005_d 0.010589f $X=1.305 $Y=2.035 $X2=-0.19
+ $Y2=1.66
cc_131 N_A_71_368#_c_166_n N_VPWR_c_194_n 0.0266773f $X=0.48 $Y=2.815 $X2=0
+ $Y2=0
cc_132 N_A_71_368#_c_171_n N_VPWR_c_194_n 0.022455f $X=1.305 $Y=2.035 $X2=0
+ $Y2=0
cc_133 N_A_71_368#_c_167_n N_VPWR_c_194_n 0.0266773f $X=1.47 $Y=2.815 $X2=0
+ $Y2=0
cc_134 N_A_71_368#_c_166_n N_VPWR_c_195_n 0.0145938f $X=0.48 $Y=2.815 $X2=0
+ $Y2=0
cc_135 N_A_71_368#_c_167_n N_VPWR_c_197_n 0.014552f $X=1.47 $Y=2.815 $X2=0 $Y2=0
cc_136 N_A_71_368#_c_166_n N_VPWR_c_193_n 0.0120466f $X=0.48 $Y=2.815 $X2=0
+ $Y2=0
cc_137 N_A_71_368#_c_167_n N_VPWR_c_193_n 0.0119791f $X=1.47 $Y=2.815 $X2=0
+ $Y2=0
cc_138 N_A_71_368#_c_167_n N_Y_c_225_n 0.0163053f $X=1.47 $Y=2.815 $X2=0 $Y2=0
cc_139 N_VPWR_c_197_n N_Y_c_225_n 0.0226653f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_140 N_VPWR_c_193_n N_Y_c_225_n 0.018408f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_141 N_Y_c_224_n N_VGND_M1004_d 0.00345356f $X=2.045 $Y=0.995 $X2=0 $Y2=0
cc_142 N_Y_c_219_n N_VGND_c_270_n 0.0123945f $X=1.292 $Y=0.81 $X2=0 $Y2=0
cc_143 N_Y_c_220_n N_VGND_c_270_n 0.0170764f $X=1.315 $Y=0.515 $X2=0 $Y2=0
cc_144 N_Y_c_220_n N_VGND_c_271_n 0.0118921f $X=1.315 $Y=0.515 $X2=0 $Y2=0
cc_145 N_Y_c_221_n N_VGND_c_271_n 0.0116858f $X=2.375 $Y=0.515 $X2=0 $Y2=0
cc_146 N_Y_c_224_n N_VGND_c_271_n 0.0249165f $X=2.045 $Y=0.995 $X2=0 $Y2=0
cc_147 N_Y_c_220_n N_VGND_c_274_n 0.0182222f $X=1.315 $Y=0.515 $X2=0 $Y2=0
cc_148 N_Y_c_221_n N_VGND_c_275_n 0.0145369f $X=2.375 $Y=0.515 $X2=0 $Y2=0
cc_149 N_Y_c_220_n N_VGND_c_276_n 0.0149207f $X=1.315 $Y=0.515 $X2=0 $Y2=0
cc_150 N_Y_c_221_n N_VGND_c_276_n 0.0119879f $X=2.375 $Y=0.515 $X2=0 $Y2=0
cc_151 Y N_VGND_c_276_n 0.0057112f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_152 N_Y_c_224_n N_VGND_c_276_n 0.00707419f $X=2.045 $Y=0.995 $X2=0 $Y2=0
