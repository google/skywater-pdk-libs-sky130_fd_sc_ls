* NGSPICE file created from sky130_fd_sc_ls__o211a_4.ext - technology: sky130A

.subckt sky130_fd_sc_ls__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
M1000 a_968_391# A1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=6e+11p pd=5.2e+06u as=2.5064e+12p ps=1.74e+07u
M1001 a_91_48# A2 a_968_391# VPB phighvt w=1e+06u l=150000u
+  ad=8.54e+11p pd=7.26e+06u as=0p ps=0u
M1002 a_510_125# A2 VGND VNB nshort w=640000u l=150000u
+  ad=8.089e+11p pd=7.65e+06u as=1.1032e+12p ps=1.016e+07u
M1003 a_91_48# B1 VPWR VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_91_48# C1 VPWR VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_968_391# A2 a_91_48# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND A1 a_510_125# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_91_48# VGND VNB nshort w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=0p ps=0u
M1008 VPWR a_91_48# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=6.72e+11p ps=5.68e+06u
M1009 VPWR C1 a_91_48# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR B1 a_91_48# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_510_125# B1 a_597_125# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=4.032e+11p ps=3.82e+06u
M1012 X a_91_48# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_597_125# C1 a_91_48# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1014 VPWR A1 a_968_391# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 X a_91_48# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND a_91_48# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 X a_91_48# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_597_125# B1 a_510_125# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND A2 a_510_125# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_510_125# A1 VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_91_48# C1 a_597_125# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPWR a_91_48# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VGND a_91_48# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

