* File: sky130_fd_sc_ls__a221o_1.spice
* Created: Wed Sep  2 10:49:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__a221o_1.pex.spice"
.subckt sky130_fd_sc_ls__a221o_1  VNB VPB A2 A1 B1 B2 C1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* C1	C1
* B2	B2
* B1	B1
* A1	A1
* A2	A2
* VPB	VPB
* VNB	VNB
MM1004 N_VGND_M1004_d N_A_148_260#_M1004_g N_X_M1004_s VNB NSHORT L=0.15 W=0.74
+ AD=0.310465 AS=0.1961 PD=1.7213 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75002.5 A=0.111 P=1.78 MULT=1
MM1002 A_417_79# N_A2_M1002_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.64 AD=0.0672
+ AS=0.26851 PD=0.85 PS=1.4887 NRD=9.372 NRS=0 M=1 R=4.26667 SA=75001.2
+ SB=75001.8 A=0.096 P=1.58 MULT=1
MM1003 N_A_148_260#_M1003_d N_A1_M1003_g A_417_79# VNB NSHORT L=0.15 W=0.64
+ AD=0.1248 AS=0.0672 PD=1.03 PS=0.85 NRD=10.308 NRS=9.372 M=1 R=4.26667
+ SA=75001.6 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1005 A_597_79# N_B1_M1005_g N_A_148_260#_M1003_d VNB NSHORT L=0.15 W=0.64
+ AD=0.0672 AS=0.1248 PD=0.85 PS=1.03 NRD=9.372 NRS=10.308 M=1 R=4.26667
+ SA=75002.1 SB=75000.9 A=0.096 P=1.58 MULT=1
MM1006 N_VGND_M1006_d N_B2_M1006_g A_597_79# VNB NSHORT L=0.15 W=0.64 AD=0.14295
+ AS=0.0672 PD=1.25 PS=0.85 NRD=3.744 NRS=9.372 M=1 R=4.26667 SA=75002.5
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1001 N_A_148_260#_M1001_d N_C1_M1001_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.64
+ AD=0.1696 AS=0.14295 PD=1.81 PS=1.25 NRD=0 NRS=16.872 M=1 R=4.26667 SA=75002
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1007 N_VPWR_M1007_d N_A_148_260#_M1007_g N_X_M1007_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.210264 AS=0.308 PD=1.56906 PS=2.79 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1008 N_A_310_392#_M1008_d N_A2_M1008_g N_VPWR_M1007_d VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.187736 PD=1.3 PS=1.40094 NRD=1.9503 NRS=14.775 M=1 R=6.66667
+ SA=75000.7 SB=75000.6 A=0.15 P=2.3 MULT=1
MM1010 N_VPWR_M1010_d N_A1_M1010_g N_A_310_392#_M1008_d VPB PHIGHVT L=0.15 W=1
+ AD=0.275 AS=0.15 PD=2.55 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75001.2
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1011 N_A_310_392#_M1011_d N_B1_M1011_g N_A_509_392#_M1011_s VPB PHIGHVT L=0.15
+ W=1 AD=0.15 AS=0.275 PD=1.3 PS=2.55 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75001.1 A=0.15 P=2.3 MULT=1
MM1000 N_A_509_392#_M1000_d N_B2_M1000_g N_A_310_392#_M1011_d VPB PHIGHVT L=0.15
+ W=1 AD=0.165 AS=0.15 PD=1.33 PS=1.3 NRD=4.9053 NRS=1.9503 M=1 R=6.66667
+ SA=75000.6 SB=75000.7 A=0.15 P=2.3 MULT=1
MM1009 N_A_148_260#_M1009_d N_C1_M1009_g N_A_509_392#_M1000_d VPB PHIGHVT L=0.15
+ W=1 AD=0.275 AS=0.165 PD=2.55 PS=1.33 NRD=1.9503 NRS=4.9053 M=1 R=6.66667
+ SA=75001.1 SB=75000.2 A=0.15 P=2.3 MULT=1
DX12_noxref VNB VPB NWDIODE A=8.742 P=13.12
*
.include "sky130_fd_sc_ls__a221o_1.pxi.spice"
*
.ends
*
*
