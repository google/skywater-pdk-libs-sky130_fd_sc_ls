* NGSPICE file created from sky130_fd_sc_ls__a2111oi_2.ext - technology: sky130A

.subckt sky130_fd_sc_ls__a2111oi_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
M1000 VGND C1 Y VNB nshort w=740000u l=150000u
+  ad=7.141e+11p pd=6.37e+06u as=6.919e+11p ps=6.31e+06u
M1001 a_722_74# A1 Y VNB nshort w=740000u l=150000u
+  ad=5.994e+11p pd=6.06e+06u as=0p ps=0u
M1002 a_69_368# D1 Y VPB phighvt w=1.12e+06u l=150000u
+  ad=9.52e+11p pd=8.42e+06u as=3.36e+11p ps=2.84e+06u
M1003 VPWR A2 a_533_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=6.72e+11p pd=5.68e+06u as=1.288e+12p ps=1.126e+07u
M1004 a_69_368# C1 a_334_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=6.72e+11p ps=5.68e+06u
M1005 a_533_368# A2 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_334_368# B1 a_533_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_722_74# A2 VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_334_368# C1 a_69_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y D1 VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_533_368# B1 a_334_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Y B1 VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR A1 a_533_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND A2 a_722_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Y A1 a_722_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_533_368# A1 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Y D1 a_69_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

