* NGSPICE file created from sky130_fd_sc_ls__dfstp_1.ext - technology: sky130A

.subckt sky130_fd_sc_ls__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
M1000 VPWR CLK a_224_350# VPB phighvt w=1.12e+06u l=150000u
+  ad=1.8422e+12p pd=1.597e+07u as=3.192e+11p ps=2.81e+06u
M1001 VPWR SET_B a_760_395# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.26e+11p ps=1.44e+06u
M1002 a_1457_508# a_398_74# a_1298_392# VPB phighvt w=420000u l=150000u
+  ad=1.134e+11p pd=1.38e+06u as=5.488e+11p ps=4.68e+06u
M1003 a_1298_392# SET_B VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Q a_1902_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.192e+11p pd=2.81e+06u as=0p ps=0u
M1005 a_1470_48# a_1298_392# VGND VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=1.40335e+12p ps=1.213e+07u
M1006 a_1298_392# a_398_74# a_1215_74# VNB nshort w=640000u l=150000u
+  ad=2.139e+11p pd=2e+06u as=2.4e+11p ps=2.03e+06u
M1007 a_709_463# a_224_350# a_604_74# VPB phighvt w=420000u l=150000u
+  ad=1.134e+11p pd=1.38e+06u as=1.47e+11p ps=1.54e+06u
M1008 VGND SET_B a_1027_118# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1009 a_1027_118# a_604_74# a_760_395# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.176e+11p ps=1.4e+06u
M1010 a_604_74# a_224_350# a_27_74# VNB nshort w=420000u l=150000u
+  ad=2.226e+11p pd=1.9e+06u as=2.9565e+11p ps=3.17e+06u
M1011 a_398_74# a_224_350# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=0p ps=0u
M1012 Q a_1902_74# VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1013 a_1422_74# a_224_350# a_1298_392# VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1014 a_1500_74# a_1470_48# a_1422_74# VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1015 a_398_74# a_224_350# VGND VNB nshort w=740000u l=150000u
+  ad=1.961e+11p pd=2.01e+06u as=0p ps=0u
M1016 a_1470_48# a_1298_392# VPWR VPB phighvt w=420000u l=150000u
+  ad=1.155e+11p pd=1.39e+06u as=0p ps=0u
M1017 VGND a_760_395# a_740_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1018 a_1197_341# a_604_74# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=3.99625e+11p pd=3.22e+06u as=0p ps=0u
M1019 a_1298_392# a_224_350# a_1197_341# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND SET_B a_1500_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPWR D a_27_74# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=2.436e+11p ps=2.84e+06u
M1022 a_740_74# a_398_74# a_604_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VGND a_1298_392# a_1902_74# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1024 VGND D a_27_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPWR a_1470_48# a_1457_508# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VGND CLK a_224_350# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1027 a_604_74# a_398_74# a_27_74# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VPWR a_760_395# a_709_463# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_760_395# a_604_74# VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_1215_74# a_604_74# VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VPWR a_1298_392# a_1902_74# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=2.31e+11p ps=2.23e+06u
.ends

