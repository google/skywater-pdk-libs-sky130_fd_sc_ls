* NGSPICE file created from sky130_fd_sc_ls__sdfxbp_1.ext - technology: sky130A

.subckt sky130_fd_sc_ls__sdfxbp_1 CLK D SCD SCE VGND VNB VPB VPWR Q Q_N
M1000 VPWR SCE a_31_74# VPB phighvt w=640000u l=150000u
+  ad=2.6944e+12p pd=2.048e+07u as=1.888e+11p ps=1.87e+06u
M1001 a_434_74# SCE a_296_74# VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=3.423e+11p ps=3.31e+06u
M1002 VPWR a_1723_48# a_2216_112# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=2.31e+11p ps=2.23e+06u
M1003 a_1157_100# a_828_74# a_1021_100# VNB nshort w=420000u l=150000u
+  ad=1.932e+11p pd=1.76e+06u as=2.226e+11p ps=1.9e+06u
M1004 a_218_74# a_31_74# VGND VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=1.8401e+12p ps=1.538e+07u
M1005 a_296_74# D a_218_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_233_464# SCE VPWR VPB phighvt w=640000u l=150000u
+  ad=1.728e+11p pd=1.82e+06u as=0p ps=0u
M1007 a_828_74# a_612_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1008 VPWR SCD a_407_464# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=2.496e+11p ps=2.06e+06u
M1009 a_1529_74# a_828_74# a_1243_398# VNB nshort w=550000u l=150000u
+  ad=2.887e+11p pd=2.32e+06u as=1.5675e+11p ps=1.67e+06u
M1010 a_1243_398# a_1021_100# VGND VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Q a_1723_48# VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1012 a_1723_48# a_1529_74# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.75e+11p pd=2.55e+06u as=0p ps=0u
M1013 VPWR a_1243_398# a_1180_496# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.386e+11p ps=1.5e+06u
M1014 a_828_74# a_612_74# VGND VNB nshort w=740000u l=150000u
+  ad=1.998e+11p pd=2.02e+06u as=0p ps=0u
M1015 VGND a_1243_398# a_1157_100# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_1021_100# a_828_74# a_296_74# VPB phighvt w=420000u l=150000u
+  ad=1.26e+11p pd=1.44e+06u as=3.096e+11p ps=3.28e+06u
M1017 a_1681_74# a_612_74# a_1529_74# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1018 a_1243_398# a_1021_100# VPWR VPB phighvt w=840000u l=150000u
+  ad=6.468e+11p pd=3.22e+06u as=0p ps=0u
M1019 VGND a_1723_48# a_1681_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_1529_74# a_612_74# a_1243_398# VPB phighvt w=840000u l=150000u
+  ad=2.856e+11p pd=2.45e+06u as=0p ps=0u
M1021 a_612_74# CLK VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1022 a_612_74# CLK VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=0p ps=0u
M1023 VGND SCE a_31_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1024 a_1180_496# a_612_74# a_1021_100# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 Q_N a_2216_112# VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1026 a_296_74# D a_233_464# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VGND SCD a_434_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_1021_100# a_612_74# a_296_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPWR a_1723_48# a_1691_508# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1030 Q a_1723_48# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.08e+11p pd=2.79e+06u as=0p ps=0u
M1031 Q_N a_2216_112# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.192e+11p pd=2.81e+06u as=0p ps=0u
M1032 a_407_464# a_31_74# a_296_74# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VGND a_1723_48# a_2216_112# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1034 a_1691_508# a_828_74# a_1529_74# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_1723_48# a_1529_74# VGND VNB nshort w=550000u l=150000u
+  ad=1.5675e+11p pd=1.67e+06u as=0p ps=0u
.ends

