* File: sky130_fd_sc_ls__clkdlyinv3sd2_1.spice
* Created: Wed Sep  2 10:58:03 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__clkdlyinv3sd2_1.pex.spice"
.subckt sky130_fd_sc_ls__clkdlyinv3sd2_1  VNB VPB A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1001 N_VGND_M1001_d N_A_M1001_g N_A_28_74#_M1001_s VNB NSHORT L=0.15 W=0.42
+ AD=0.14805 AS=0.1113 PD=1.125 PS=1.37 NRD=15.708 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1000 N_A_288_74#_M1000_d N_A_28_74#_M1000_g N_VGND_M1001_d VNB NSHORT L=0.18
+ W=0.42 AD=0.1113 AS=0.14805 PD=1.37 PS=1.125 NRD=0 NRS=105.708 M=1 R=2.33333
+ SA=90001 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1005 N_Y_M1005_d N_A_288_74#_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1002 N_VPWR_M1002_d N_A_M1002_g N_A_28_74#_M1002_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.346989 AS=0.3136 PD=1.84377 PS=2.8 NRD=5.2599 NRS=2.6201 M=1 R=7.46667
+ SA=75000.2 SB=75001 A=0.168 P=2.54 MULT=1
MM1003 N_A_288_74#_M1003_d N_A_28_74#_M1003_g N_VPWR_M1002_d VPB PHIGHVT L=0.25
+ W=1 AD=0.26 AS=0.309811 PD=2.52 PS=1.64623 NRD=0 NRS=62.0353 M=1 R=4 SA=125001
+ SB=125000 A=0.25 P=2.5 MULT=1
MM1004 N_Y_M1004_d N_A_288_74#_M1004_g N_VPWR_M1004_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3136 AS=0.308 PD=2.8 PS=2.79 NRD=2.6201 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.2 A=0.168 P=2.54 MULT=1
DX6_noxref VNB VPB NWDIODE A=6.0636 P=10.24
*
.include "sky130_fd_sc_ls__clkdlyinv3sd2_1.pxi.spice"
*
.ends
*
*
