* NGSPICE file created from sky130_fd_sc_ls__buf_1.ext - technology: sky130A

.subckt sky130_fd_sc_ls__buf_1 A VGND VNB VPB VPWR X
M1000 VPWR A a_27_164# VPB phighvt w=840000u l=150000u
+  ad=4.102e+11p pd=3.04e+06u as=2.478e+11p ps=2.27e+06u
M1001 VGND A a_27_164# VNB nshort w=550000u l=150000u
+  ad=3.0395e+11p pd=2.34e+06u as=2.4915e+11p ps=2.37e+06u
M1002 X a_27_164# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=0p ps=0u
M1003 X a_27_164# VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
.ends

