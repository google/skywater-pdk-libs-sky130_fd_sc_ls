* File: sky130_fd_sc_ls__einvp_2.spice
* Created: Wed Sep  2 11:07:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__einvp_2.pex.spice"
.subckt sky130_fd_sc_ls__einvp_2  VNB VPB A TE Z VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Z	Z
* TE	TE
* A	A
* VPB	VPB
* VNB	VNB
MM1001 N_A_36_74#_M1001_d N_A_M1001_g N_Z_M1001_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.5 A=0.111 P=1.78 MULT=1
MM1008 N_A_36_74#_M1008_d N_A_M1008_g N_Z_M1001_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1003 N_VGND_M1003_d N_TE_M1003_g N_A_36_74#_M1008_d VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1007 N_VGND_M1003_d N_TE_M1007_g N_A_36_74#_M1007_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1009 N_VGND_M1009_d N_TE_M1009_g N_A_263_323#_M1009_s VNB NSHORT L=0.15 W=0.42
+ AD=0.126 AS=0.1197 PD=1.44 PS=1.41 NRD=1.428 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1004 N_Z_M1004_d N_A_M1004_g N_A_27_368#_M1004_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1005 N_Z_M1004_d N_A_M1005_g N_A_27_368#_M1005_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1000 N_A_27_368#_M1005_s N_A_263_323#_M1000_g N_VPWR_M1000_s VPB PHIGHVT
+ L=0.15 W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1
+ R=7.46667 SA=75001.1 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1006 N_A_27_368#_M1006_d N_A_263_323#_M1006_g N_VPWR_M1000_s VPB PHIGHVT
+ L=0.15 W=1.12 AD=0.3248 AS=0.168 PD=2.82 PS=1.42 NRD=1.7533 NRS=1.7533 M=1
+ R=7.46667 SA=75001.6 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1002 N_VPWR_M1002_d N_TE_M1002_g N_A_263_323#_M1002_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1888 AS=0.1856 PD=1.87 PS=1.86 NRD=3.0732 NRS=3.0732 M=1 R=4.26667
+ SA=75000.2 SB=75000.2 A=0.096 P=1.58 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9564 P=11.2
c_43 VNB 0 1.40666e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_ls__einvp_2.pxi.spice"
*
.ends
*
*
