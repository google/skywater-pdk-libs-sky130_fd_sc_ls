* File: sky130_fd_sc_ls__xor3_4.spice
* Created: Fri Aug 28 14:11:10 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__xor3_4.pex.spice"
.subckt sky130_fd_sc_ls__xor3_4  VNB VPB A B C VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* C	C
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1006 N_VGND_M1006_d N_A_74_294#_M1006_g N_A_27_118#_M1006_s VNB NSHORT L=0.15
+ W=0.64 AD=0.24225 AS=0.1824 PD=1.57 PS=1.85 NRD=60.648 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75002.9 A=0.096 P=1.58 MULT=1
MM1024 N_A_74_294#_M1024_d N_A_M1024_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.64
+ AD=0.2208 AS=0.24225 PD=1.33 PS=1.57 NRD=29.988 NRS=60.648 M=1 R=4.26667
+ SA=75000.9 SB=75002.3 A=0.096 P=1.58 MULT=1
MM1017 N_A_416_118#_M1017_d N_B_M1017_g N_A_74_294#_M1024_d VNB NSHORT L=0.15
+ W=0.64 AD=0.125283 AS=0.2208 PD=1.19547 PS=1.33 NRD=0 NRS=46.872 M=1 R=4.26667
+ SA=75001.7 SB=75001.4 A=0.096 P=1.58 MULT=1
MM1020 N_A_27_118#_M1020_d N_A_397_320#_M1020_g N_A_416_118#_M1017_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.0966792 AS=0.082217 PD=0.863774 PS=0.784528 NRD=0
+ NRS=20.712 M=1 R=2.8 SA=75002.2 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1007 N_A_323_392#_M1007_d N_B_M1007_g N_A_27_118#_M1020_d VNB NSHORT L=0.15
+ W=0.64 AD=0.145875 AS=0.147321 PD=1.115 PS=1.31623 NRD=14.988 NRS=31.872 M=1
+ R=4.26667 SA=75001.9 SB=75000.9 A=0.096 P=1.58 MULT=1
MM1026 N_A_74_294#_M1026_d N_A_397_320#_M1026_g N_A_323_392#_M1007_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.2848 AS=0.145875 PD=2.17 PS=1.115 NRD=31.872 NRS=14.988 M=1
+ R=4.26667 SA=75002.5 SB=75000.4 A=0.096 P=1.58 MULT=1
MM1025 N_VGND_M1025_d N_B_M1025_g N_A_397_320#_M1025_s VNB NSHORT L=0.15 W=0.74
+ AD=0.42 AS=0.2072 PD=2.67 PS=2.04 NRD=41.34 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.4 A=0.111 P=1.78 MULT=1
MM1010 N_A_1218_388#_M1010_d N_A_1155_284#_M1010_g N_A_323_392#_M1010_s VNB
+ NSHORT L=0.15 W=0.64 AD=0.1696 AS=0.176 PD=1.17 PS=1.83 NRD=46.872 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75000.9 A=0.096 P=1.58 MULT=1
MM1018 N_A_416_118#_M1018_d N_C_M1018_g N_A_1218_388#_M1010_d VNB NSHORT L=0.15
+ W=0.64 AD=0.1824 AS=0.1696 PD=1.85 PS=1.17 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.9 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1027 N_VGND_M1027_d N_C_M1027_g N_A_1155_284#_M1027_s VNB NSHORT L=0.15 W=0.42
+ AD=0.106521 AS=0.2121 PD=0.847241 PS=1.85 NRD=22.848 NRS=0 M=1 R=2.8
+ SA=75000.4 SB=75002.1 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1027_d N_A_1218_388#_M1003_g N_X_M1003_s VNB NSHORT L=0.15 W=0.74
+ AD=0.187679 AS=0.1036 PD=1.49276 PS=1.02 NRD=5.664 NRS=0 M=1 R=4.93333
+ SA=75000.7 SB=75001.5 A=0.111 P=1.78 MULT=1
MM1011 N_VGND_M1011_d N_A_1218_388#_M1011_g N_X_M1003_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1012 N_VGND_M1011_d N_A_1218_388#_M1012_g N_X_M1012_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.6
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1023 N_VGND_M1023_d N_A_1218_388#_M1023_g N_X_M1012_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2072 AS=0.1036 PD=2.04 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1021 N_VPWR_M1021_d N_A_74_294#_M1021_g N_A_27_118#_M1021_s VPB PHIGHVT L=0.15
+ W=1 AD=0.175 AS=0.295 PD=1.35 PS=2.59 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75002.3 A=0.15 P=2.3 MULT=1
MM1019 N_A_74_294#_M1019_d N_A_M1019_g N_VPWR_M1021_d VPB PHIGHVT L=0.15 W=1
+ AD=0.201413 AS=0.175 PD=1.50543 PS=1.35 NRD=1.9503 NRS=11.8003 M=1 R=6.66667
+ SA=75000.7 SB=75001.8 A=0.15 P=2.3 MULT=1
MM1002 N_A_323_392#_M1002_d N_B_M1002_g N_A_74_294#_M1019_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.173335 AS=0.169187 PD=1.39054 PS=1.26457 NRD=2.3443 NRS=22.655 M=1
+ R=5.6 SA=75001.3 SB=75001.5 A=0.126 P=1.98 MULT=1
MM1000 N_A_27_118#_M1000_d N_A_397_320#_M1000_g N_A_323_392#_M1002_d VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.149875 AS=0.132065 PD=1.215 PS=1.05946 NRD=3.0732
+ NRS=30.0031 M=1 R=4.26667 SA=75001.8 SB=75001.4 A=0.096 P=1.58 MULT=1
MM1004 N_A_416_118#_M1004_d N_B_M1004_g N_A_27_118#_M1000_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.132 AS=0.149875 PD=1.05946 PS=1.215 NRD=29.2348 NRS=47.6937 M=1
+ R=4.26667 SA=75001.9 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1014 N_A_74_294#_M1014_d N_A_397_320#_M1014_g N_A_416_118#_M1004_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.546 AS=0.17325 PD=2.98 PS=1.39054 NRD=75.0373 NRS=2.3443
+ M=1 R=5.6 SA=75001.9 SB=75000.6 A=0.126 P=1.98 MULT=1
MM1009 N_VPWR_M1009_d N_B_M1009_g N_A_397_320#_M1009_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.3304 PD=2.83 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1022 N_A_1218_388#_M1022_d N_A_1155_284#_M1022_g N_A_416_118#_M1022_s VPB
+ PHIGHVT L=0.15 W=0.84 AD=0.2226 AS=0.3822 PD=1.37 PS=2.59 NRD=56.2829
+ NRS=39.8531 M=1 R=5.6 SA=75000.4 SB=75000.9 A=0.126 P=1.98 MULT=1
MM1015 N_A_323_392#_M1015_d N_C_M1015_g N_A_1218_388#_M1022_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.2478 AS=0.2226 PD=2.27 PS=1.37 NRD=2.3443 NRS=2.3443 M=1 R=5.6
+ SA=75001.1 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1016 N_VPWR_M1016_d N_C_M1016_g N_A_1155_284#_M1016_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.291782 AS=0.1888 PD=1.36364 PS=1.87 NRD=123.401 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75002.6 A=0.096 P=1.58 MULT=1
MM1001 N_VPWR_M1016_d N_A_1218_388#_M1001_g N_X_M1001_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.510618 AS=0.168 PD=2.38636 PS=1.42 NRD=66.8224 NRS=1.7533 M=1
+ R=7.46667 SA=75000.9 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1005 N_VPWR_M1005_d N_A_1218_388#_M1005_g N_X_M1001_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.2128 AS=0.168 PD=1.5 PS=1.42 NRD=15.8191 NRS=1.7533 M=1 R=7.46667
+ SA=75001.3 SB=75001.2 A=0.168 P=2.54 MULT=1
MM1008 N_VPWR_M1005_d N_A_1218_388#_M1008_g N_X_M1008_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.2128 AS=0.168 PD=1.5 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.9 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1013 N_VPWR_M1013_d N_A_1218_388#_M1013_g N_X_M1008_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.3 SB=75000.2 A=0.168 P=2.54 MULT=1
DX28_noxref VNB VPB NWDIODE A=20.3484 P=25.6
c_203 VPB 0 1.12299e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_ls__xor3_4.pxi.spice"
*
.ends
*
*
