* NGSPICE file created from sky130_fd_sc_ls__and2_2.ext - technology: sky130A

.subckt sky130_fd_sc_ls__and2_2 A B VGND VNB VPB VPWR X
M1000 VPWR a_31_74# X VPB phighvt w=1.12e+06u l=150000u
+  ad=9.96e+11p pd=8.34e+06u as=3.36e+11p ps=2.84e+06u
M1001 VGND B a_118_74# VNB nshort w=740000u l=150000u
+  ad=5.217e+11p pd=4.37e+06u as=1.776e+11p ps=1.96e+06u
M1002 X a_31_74# VGND VNB nshort w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1003 a_118_74# A a_31_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1004 X a_31_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_31_74# A VPWR VPB phighvt w=1e+06u l=150000u
+  ad=3e+11p pd=2.6e+06u as=0p ps=0u
M1006 VPWR B a_31_74# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND a_31_74# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

