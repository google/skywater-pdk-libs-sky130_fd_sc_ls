* NGSPICE file created from sky130_fd_sc_ls__einvn_8.ext - technology: sky130A

.subckt sky130_fd_sc_ls__einvn_8 A TE_B VGND VNB VPB VPWR Z
M1000 VPWR TE_B a_239_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=2.0104e+12p pd=1.479e+07u as=3.0128e+12p ps=2.554e+07u
M1001 Z A a_239_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=1.4e+12p pd=1.146e+07u as=0p ps=0u
M1002 a_239_368# TE_B VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VGND a_126_74# a_293_74# VNB nshort w=740000u l=150000u
+  ad=1.1433e+12p pd=1.049e+07u as=1.924e+12p ps=1.852e+07u
M1004 Z A a_293_74# VNB nshort w=740000u l=150000u
+  ad=9.324e+11p pd=8.44e+06u as=0p ps=0u
M1005 VGND a_126_74# a_293_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Z A a_239_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Z A a_293_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_239_368# TE_B VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_239_368# A Z VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 Z A a_293_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_239_368# A Z VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR TE_B a_239_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 Z A a_293_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Z A a_239_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_293_74# a_126_74# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND a_126_74# a_293_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_293_74# A Z VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR TE_B a_239_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND a_126_74# a_293_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_126_74# TE_B VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=0p ps=0u
M1021 Z A a_239_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_293_74# A Z VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_239_368# TE_B VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_293_74# A Z VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_239_368# A Z VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_293_74# a_126_74# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_239_368# TE_B VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_239_368# A Z VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_293_74# A Z VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_293_74# a_126_74# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VPWR TE_B a_239_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_126_74# TE_B VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1033 a_293_74# a_126_74# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

