* File: sky130_fd_sc_ls__o2bb2ai_1.pxi.spice
* Created: Wed Sep  2 11:20:53 2020
* 
x_PM_SKY130_FD_SC_LS__O2BB2AI_1%A1_N N_A1_N_M1009_g N_A1_N_c_65_n N_A1_N_c_69_n
+ N_A1_N_M1008_g N_A1_N_c_70_n A1_N N_A1_N_c_67_n
+ PM_SKY130_FD_SC_LS__O2BB2AI_1%A1_N
x_PM_SKY130_FD_SC_LS__O2BB2AI_1%A2_N N_A2_N_c_96_n N_A2_N_M1001_g N_A2_N_c_97_n
+ N_A2_N_c_98_n N_A2_N_c_101_n N_A2_N_M1004_g A2_N N_A2_N_c_99_n
+ PM_SKY130_FD_SC_LS__O2BB2AI_1%A2_N
x_PM_SKY130_FD_SC_LS__O2BB2AI_1%A_131_383# N_A_131_383#_M1001_d
+ N_A_131_383#_M1008_d N_A_131_383#_M1007_g N_A_131_383#_c_144_n
+ N_A_131_383#_M1003_g N_A_131_383#_c_137_n N_A_131_383#_c_138_n
+ N_A_131_383#_c_147_n N_A_131_383#_c_139_n N_A_131_383#_c_140_n
+ N_A_131_383#_c_141_n N_A_131_383#_c_142_n N_A_131_383#_c_143_n
+ PM_SKY130_FD_SC_LS__O2BB2AI_1%A_131_383#
x_PM_SKY130_FD_SC_LS__O2BB2AI_1%B2 N_B2_c_208_n N_B2_M1006_g N_B2_M1005_g B2
+ PM_SKY130_FD_SC_LS__O2BB2AI_1%B2
x_PM_SKY130_FD_SC_LS__O2BB2AI_1%B1 N_B1_M1000_g N_B1_c_244_n N_B1_M1002_g B1
+ N_B1_c_245_n PM_SKY130_FD_SC_LS__O2BB2AI_1%B1
x_PM_SKY130_FD_SC_LS__O2BB2AI_1%VPWR N_VPWR_M1008_s N_VPWR_M1004_d
+ N_VPWR_M1002_d N_VPWR_c_267_n N_VPWR_c_268_n N_VPWR_c_269_n N_VPWR_c_270_n
+ N_VPWR_c_271_n N_VPWR_c_272_n VPWR N_VPWR_c_273_n N_VPWR_c_274_n
+ N_VPWR_c_266_n PM_SKY130_FD_SC_LS__O2BB2AI_1%VPWR
x_PM_SKY130_FD_SC_LS__O2BB2AI_1%Y N_Y_M1007_s N_Y_M1003_d N_Y_c_304_n
+ N_Y_c_305_n N_Y_c_316_n N_Y_c_306_n Y Y PM_SKY130_FD_SC_LS__O2BB2AI_1%Y
x_PM_SKY130_FD_SC_LS__O2BB2AI_1%VGND N_VGND_M1009_s N_VGND_M1005_d
+ N_VGND_c_339_n N_VGND_c_340_n N_VGND_c_341_n N_VGND_c_342_n N_VGND_c_343_n
+ VGND N_VGND_c_344_n N_VGND_c_345_n PM_SKY130_FD_SC_LS__O2BB2AI_1%VGND
x_PM_SKY130_FD_SC_LS__O2BB2AI_1%A_397_74# N_A_397_74#_M1007_d
+ N_A_397_74#_M1000_d N_A_397_74#_c_374_n N_A_397_74#_c_375_n
+ N_A_397_74#_c_376_n PM_SKY130_FD_SC_LS__O2BB2AI_1%A_397_74#
cc_1 VNB N_A1_N_M1009_g 0.0264785f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.69
cc_2 VNB N_A1_N_c_65_n 0.0127045f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.69
cc_3 VNB A1_N 0.00842345f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_A1_N_c_67_n 0.0575593f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.345
cc_5 VNB N_A2_N_c_96_n 0.0213804f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.18
cc_6 VNB N_A2_N_c_97_n 0.0325601f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A2_N_c_98_n 0.0118868f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.51
cc_8 VNB N_A2_N_c_99_n 0.010302f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_131_383#_M1007_g 0.029599f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=2.335
cc_10 VNB N_A_131_383#_c_137_n 0.0320644f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_11 VNB N_A_131_383#_c_138_n 0.0100085f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_131_383#_c_139_n 0.00235188f $X=-0.19 $Y=-0.245 $X2=0.495
+ $Y2=1.345
cc_13 VNB N_A_131_383#_c_140_n 0.00269016f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_131_383#_c_141_n 0.0130007f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_131_383#_c_142_n 0.00978707f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_131_383#_c_143_n 0.00759225f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_B2_c_208_n 0.028427f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.18
cc_18 VNB N_B2_M1005_g 0.0227963f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.69
cc_19 VNB B2 0.00645769f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=2.335
cc_20 VNB N_B1_M1000_g 0.0302424f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.69
cc_21 VNB N_B1_c_244_n 0.0605966f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.51
cc_22 VNB N_B1_c_245_n 0.0051843f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.765
cc_23 VNB N_VPWR_c_266_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_Y_c_304_n 0.00210709f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=2.335
cc_25 VNB N_Y_c_305_n 0.00328206f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_Y_c_306_n 0.00368918f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.345
cc_27 VNB N_VGND_c_339_n 0.0120272f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.84
cc_28 VNB N_VGND_c_340_n 0.0321458f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=2.335
cc_29 VNB N_VGND_c_341_n 0.00799303f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_342_n 0.0583747f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.345
cc_31 VNB N_VGND_c_343_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.345
cc_32 VNB N_VGND_c_344_n 0.0202653f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_345_n 0.223677f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_397_74#_c_374_n 0.0116093f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.84
cc_35 VNB N_A_397_74#_c_375_n 0.02581f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_397_74#_c_376_n 0.00181981f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_37 VPB N_A1_N_c_65_n 0.00246017f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.69
cc_38 VPB N_A1_N_c_69_n 0.016939f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=1.84
cc_39 VPB N_A1_N_c_70_n 0.0207268f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=1.765
cc_40 VPB N_A2_N_c_98_n 0.00485051f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.51
cc_41 VPB N_A2_N_c_101_n 0.025062f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.69
cc_42 VPB N_A_131_383#_c_144_n 0.0175931f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_43 VPB N_A_131_383#_c_137_n 0.0180437f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_44 VPB N_A_131_383#_c_138_n 0.00717278f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_45 VPB N_A_131_383#_c_147_n 0.00356537f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.345
cc_46 VPB N_A_131_383#_c_139_n 0.00223353f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.345
cc_47 VPB N_A_131_383#_c_140_n 3.21295e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 VPB N_A_131_383#_c_142_n 0.00492845f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 VPB N_B2_c_208_n 0.0220556f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.18
cc_50 VPB B2 0.0141211f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=2.335
cc_51 VPB N_B1_c_244_n 0.0269939f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.51
cc_52 VPB N_B1_c_245_n 0.00974946f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=1.765
cc_53 VPB N_VPWR_c_267_n 0.0129883f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.765
cc_54 VPB N_VPWR_c_268_n 0.0618467f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=1.765
cc_55 VPB N_VPWR_c_269_n 0.019533f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_56 VPB N_VPWR_c_270_n 0.0163567f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.345
cc_57 VPB N_VPWR_c_271_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_272_n 0.0496032f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_273_n 0.0379253f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_274_n 0.0105403f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_266_n 0.0815821f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_Y_c_306_n 0.0014009f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.345
cc_63 VPB Y 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 N_A1_N_M1009_g N_A2_N_c_96_n 0.0448844f $X=0.495 $Y=0.69 $X2=-0.19
+ $Y2=-0.245
cc_65 N_A1_N_M1009_g N_A2_N_c_97_n 0.0205752f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_66 N_A1_N_c_70_n N_A2_N_c_98_n 0.00707903f $X=0.58 $Y=1.765 $X2=0 $Y2=0
cc_67 A1_N N_A2_N_c_98_n 2.79582e-19 $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_68 N_A1_N_c_67_n N_A2_N_c_98_n 0.00856416f $X=0.495 $Y=1.345 $X2=0 $Y2=0
cc_69 N_A1_N_c_69_n N_A2_N_c_101_n 0.0146874f $X=0.58 $Y=1.84 $X2=0 $Y2=0
cc_70 N_A1_N_M1009_g N_A2_N_c_99_n 0.0038946f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_71 N_A1_N_c_70_n N_A2_N_c_99_n 0.00162506f $X=0.58 $Y=1.765 $X2=0 $Y2=0
cc_72 A1_N N_A2_N_c_99_n 0.0220973f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_73 N_A1_N_c_69_n N_A_131_383#_c_147_n 0.014408f $X=0.58 $Y=1.84 $X2=0 $Y2=0
cc_74 N_A1_N_c_70_n N_A_131_383#_c_147_n 0.00312821f $X=0.58 $Y=1.765 $X2=0
+ $Y2=0
cc_75 N_A1_N_c_65_n N_A_131_383#_c_140_n 0.00219171f $X=0.495 $Y=1.69 $X2=0
+ $Y2=0
cc_76 N_A1_N_c_70_n N_A_131_383#_c_140_n 0.00639488f $X=0.58 $Y=1.765 $X2=0
+ $Y2=0
cc_77 N_A1_N_M1009_g N_A_131_383#_c_141_n 0.0016931f $X=0.495 $Y=0.69 $X2=0
+ $Y2=0
cc_78 N_A1_N_c_69_n N_VPWR_c_268_n 0.0206887f $X=0.58 $Y=1.84 $X2=0 $Y2=0
cc_79 N_A1_N_c_70_n N_VPWR_c_268_n 0.00241488f $X=0.58 $Y=1.765 $X2=0 $Y2=0
cc_80 A1_N N_VPWR_c_268_n 0.0134833f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_81 N_A1_N_c_67_n N_VPWR_c_268_n 0.00198021f $X=0.495 $Y=1.345 $X2=0 $Y2=0
cc_82 N_A1_N_c_69_n N_VPWR_c_269_n 0.00432667f $X=0.58 $Y=1.84 $X2=0 $Y2=0
cc_83 N_A1_N_c_69_n N_VPWR_c_266_n 0.0048347f $X=0.58 $Y=1.84 $X2=0 $Y2=0
cc_84 N_A1_N_M1009_g N_VGND_c_340_n 0.0157618f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_85 A1_N N_VGND_c_340_n 0.0187971f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_86 N_A1_N_c_67_n N_VGND_c_340_n 0.00211525f $X=0.495 $Y=1.345 $X2=0 $Y2=0
cc_87 N_A1_N_M1009_g N_VGND_c_342_n 0.00383152f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_88 N_A1_N_M1009_g N_VGND_c_345_n 0.0075725f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_89 N_A2_N_c_97_n N_A_131_383#_M1007_g 4.67916e-19 $X=1.03 $Y=1.45 $X2=0 $Y2=0
cc_90 N_A2_N_c_97_n N_A_131_383#_c_137_n 0.0171454f $X=1.03 $Y=1.45 $X2=0 $Y2=0
cc_91 N_A2_N_c_98_n N_A_131_383#_c_138_n 7.37801e-19 $X=1.03 $Y=1.75 $X2=0 $Y2=0
cc_92 N_A2_N_c_101_n N_A_131_383#_c_147_n 0.020113f $X=1.03 $Y=1.84 $X2=0 $Y2=0
cc_93 N_A2_N_c_98_n N_A_131_383#_c_139_n 0.00541749f $X=1.03 $Y=1.75 $X2=0 $Y2=0
cc_94 N_A2_N_c_101_n N_A_131_383#_c_139_n 0.00766035f $X=1.03 $Y=1.84 $X2=0
+ $Y2=0
cc_95 N_A2_N_c_99_n N_A_131_383#_c_139_n 0.00924974f $X=0.945 $Y=1.285 $X2=0
+ $Y2=0
cc_96 N_A2_N_c_97_n N_A_131_383#_c_140_n 0.00424005f $X=1.03 $Y=1.45 $X2=0 $Y2=0
cc_97 N_A2_N_c_98_n N_A_131_383#_c_140_n 0.0023321f $X=1.03 $Y=1.75 $X2=0 $Y2=0
cc_98 N_A2_N_c_101_n N_A_131_383#_c_140_n 5.66671e-19 $X=1.03 $Y=1.84 $X2=0
+ $Y2=0
cc_99 N_A2_N_c_99_n N_A_131_383#_c_140_n 0.0282724f $X=0.945 $Y=1.285 $X2=0
+ $Y2=0
cc_100 N_A2_N_c_96_n N_A_131_383#_c_141_n 0.0109415f $X=0.885 $Y=1.12 $X2=0
+ $Y2=0
cc_101 N_A2_N_c_97_n N_A_131_383#_c_141_n 0.00422317f $X=1.03 $Y=1.45 $X2=0
+ $Y2=0
cc_102 N_A2_N_c_99_n N_A_131_383#_c_141_n 0.01079f $X=0.945 $Y=1.285 $X2=0 $Y2=0
cc_103 N_A2_N_c_98_n N_A_131_383#_c_142_n 0.00312726f $X=1.03 $Y=1.75 $X2=0
+ $Y2=0
cc_104 N_A2_N_c_96_n N_A_131_383#_c_143_n 0.00410973f $X=0.885 $Y=1.12 $X2=0
+ $Y2=0
cc_105 N_A2_N_c_97_n N_A_131_383#_c_143_n 0.0068437f $X=1.03 $Y=1.45 $X2=0 $Y2=0
cc_106 N_A2_N_c_99_n N_A_131_383#_c_143_n 0.0260719f $X=0.945 $Y=1.285 $X2=0
+ $Y2=0
cc_107 N_A2_N_c_101_n N_VPWR_c_269_n 0.00432667f $X=1.03 $Y=1.84 $X2=0 $Y2=0
cc_108 N_A2_N_c_101_n N_VPWR_c_270_n 0.0115748f $X=1.03 $Y=1.84 $X2=0 $Y2=0
cc_109 N_A2_N_c_101_n N_VPWR_c_266_n 0.0048347f $X=1.03 $Y=1.84 $X2=0 $Y2=0
cc_110 N_A2_N_c_96_n N_Y_c_304_n 6.45659e-19 $X=0.885 $Y=1.12 $X2=0 $Y2=0
cc_111 N_A2_N_c_96_n N_VGND_c_340_n 0.00225941f $X=0.885 $Y=1.12 $X2=0 $Y2=0
cc_112 N_A2_N_c_96_n N_VGND_c_342_n 0.00434272f $X=0.885 $Y=1.12 $X2=0 $Y2=0
cc_113 N_A2_N_c_96_n N_VGND_c_345_n 0.00825979f $X=0.885 $Y=1.12 $X2=0 $Y2=0
cc_114 N_A_131_383#_M1007_g N_B2_c_208_n 0.00271721f $X=1.91 $Y=0.74 $X2=-0.19
+ $Y2=-0.245
cc_115 N_A_131_383#_c_144_n N_B2_c_208_n 0.01155f $X=1.925 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_116 N_A_131_383#_c_138_n N_B2_c_208_n 0.0246226f $X=1.925 $Y=1.557 $X2=-0.19
+ $Y2=-0.245
cc_117 N_A_131_383#_M1007_g N_B2_M1005_g 0.0265561f $X=1.91 $Y=0.74 $X2=0 $Y2=0
cc_118 N_A_131_383#_c_138_n B2 8.48581e-19 $X=1.925 $Y=1.557 $X2=0 $Y2=0
cc_119 N_A_131_383#_c_147_n N_VPWR_c_268_n 0.0346007f $X=0.805 $Y=2.06 $X2=0
+ $Y2=0
cc_120 N_A_131_383#_c_147_n N_VPWR_c_269_n 0.0078525f $X=0.805 $Y=2.06 $X2=0
+ $Y2=0
cc_121 N_A_131_383#_c_144_n N_VPWR_c_270_n 0.0244644f $X=1.925 $Y=1.765 $X2=0
+ $Y2=0
cc_122 N_A_131_383#_c_137_n N_VPWR_c_270_n 0.0019796f $X=1.835 $Y=1.515 $X2=0
+ $Y2=0
cc_123 N_A_131_383#_c_147_n N_VPWR_c_270_n 0.0308718f $X=0.805 $Y=2.06 $X2=0
+ $Y2=0
cc_124 N_A_131_383#_c_139_n N_VPWR_c_270_n 0.00914409f $X=1.27 $Y=1.705 $X2=0
+ $Y2=0
cc_125 N_A_131_383#_c_142_n N_VPWR_c_270_n 0.0354246f $X=1.525 $Y=1.515 $X2=0
+ $Y2=0
cc_126 N_A_131_383#_c_144_n N_VPWR_c_273_n 0.00303976f $X=1.925 $Y=1.765 $X2=0
+ $Y2=0
cc_127 N_A_131_383#_c_144_n N_VPWR_c_266_n 0.00404651f $X=1.925 $Y=1.765 $X2=0
+ $Y2=0
cc_128 N_A_131_383#_c_147_n N_VPWR_c_266_n 0.0105202f $X=0.805 $Y=2.06 $X2=0
+ $Y2=0
cc_129 N_A_131_383#_M1007_g N_Y_c_304_n 0.010008f $X=1.91 $Y=0.74 $X2=0 $Y2=0
cc_130 N_A_131_383#_c_141_n N_Y_c_304_n 0.0542827f $X=1.1 $Y=0.515 $X2=0 $Y2=0
cc_131 N_A_131_383#_M1007_g N_Y_c_305_n 0.0118005f $X=1.91 $Y=0.74 $X2=0 $Y2=0
cc_132 N_A_131_383#_c_137_n N_Y_c_305_n 0.00602136f $X=1.835 $Y=1.515 $X2=0
+ $Y2=0
cc_133 N_A_131_383#_c_142_n N_Y_c_305_n 0.00610005f $X=1.525 $Y=1.515 $X2=0
+ $Y2=0
cc_134 N_A_131_383#_c_143_n N_Y_c_305_n 0.0134822f $X=1.48 $Y=1.35 $X2=0 $Y2=0
cc_135 N_A_131_383#_c_144_n N_Y_c_316_n 0.00500881f $X=1.925 $Y=1.765 $X2=0
+ $Y2=0
cc_136 N_A_131_383#_M1007_g N_Y_c_306_n 0.00526729f $X=1.91 $Y=0.74 $X2=0 $Y2=0
cc_137 N_A_131_383#_c_144_n N_Y_c_306_n 0.00899026f $X=1.925 $Y=1.765 $X2=0
+ $Y2=0
cc_138 N_A_131_383#_c_138_n N_Y_c_306_n 0.0127751f $X=1.925 $Y=1.557 $X2=0 $Y2=0
cc_139 N_A_131_383#_c_142_n N_Y_c_306_n 0.0324732f $X=1.525 $Y=1.515 $X2=0 $Y2=0
cc_140 N_A_131_383#_c_143_n N_Y_c_306_n 0.00616212f $X=1.48 $Y=1.35 $X2=0 $Y2=0
cc_141 N_A_131_383#_c_144_n Y 0.0161237f $X=1.925 $Y=1.765 $X2=0 $Y2=0
cc_142 N_A_131_383#_c_141_n N_VGND_c_340_n 0.0196474f $X=1.1 $Y=0.515 $X2=0
+ $Y2=0
cc_143 N_A_131_383#_M1007_g N_VGND_c_342_n 0.00434272f $X=1.91 $Y=0.74 $X2=0
+ $Y2=0
cc_144 N_A_131_383#_c_141_n N_VGND_c_342_n 0.0222387f $X=1.1 $Y=0.515 $X2=0
+ $Y2=0
cc_145 N_A_131_383#_M1007_g N_VGND_c_345_n 0.0082698f $X=1.91 $Y=0.74 $X2=0
+ $Y2=0
cc_146 N_A_131_383#_c_141_n N_VGND_c_345_n 0.0184096f $X=1.1 $Y=0.515 $X2=0
+ $Y2=0
cc_147 N_A_131_383#_M1007_g N_A_397_74#_c_376_n 0.00182405f $X=1.91 $Y=0.74
+ $X2=0 $Y2=0
cc_148 N_B2_M1005_g N_B1_M1000_g 0.0287744f $X=2.41 $Y=0.74 $X2=0 $Y2=0
cc_149 N_B2_c_208_n N_B1_c_244_n 0.0733234f $X=2.375 $Y=1.765 $X2=0 $Y2=0
cc_150 B2 N_B1_c_244_n 0.00419936f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_151 N_B2_c_208_n N_B1_c_245_n 3.23601e-19 $X=2.375 $Y=1.765 $X2=0 $Y2=0
cc_152 B2 N_B1_c_245_n 0.0394472f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_153 N_B2_c_208_n N_VPWR_c_273_n 0.00445602f $X=2.375 $Y=1.765 $X2=0 $Y2=0
cc_154 N_B2_c_208_n N_VPWR_c_266_n 0.00858782f $X=2.375 $Y=1.765 $X2=0 $Y2=0
cc_155 N_B2_M1005_g N_Y_c_304_n 6.44813e-19 $X=2.41 $Y=0.74 $X2=0 $Y2=0
cc_156 N_B2_M1005_g N_Y_c_305_n 0.00118992f $X=2.41 $Y=0.74 $X2=0 $Y2=0
cc_157 N_B2_c_208_n N_Y_c_316_n 0.00471821f $X=2.375 $Y=1.765 $X2=0 $Y2=0
cc_158 B2 N_Y_c_316_n 0.00523276f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_159 N_B2_c_208_n N_Y_c_306_n 0.00276231f $X=2.375 $Y=1.765 $X2=0 $Y2=0
cc_160 N_B2_M1005_g N_Y_c_306_n 0.00217718f $X=2.41 $Y=0.74 $X2=0 $Y2=0
cc_161 B2 N_Y_c_306_n 0.0344158f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_162 N_B2_c_208_n Y 0.0155445f $X=2.375 $Y=1.765 $X2=0 $Y2=0
cc_163 N_B2_M1005_g N_VGND_c_341_n 0.00319142f $X=2.41 $Y=0.74 $X2=0 $Y2=0
cc_164 N_B2_M1005_g N_VGND_c_342_n 0.00424705f $X=2.41 $Y=0.74 $X2=0 $Y2=0
cc_165 N_B2_M1005_g N_VGND_c_345_n 0.00783896f $X=2.41 $Y=0.74 $X2=0 $Y2=0
cc_166 N_B2_c_208_n N_A_397_74#_c_374_n 0.00156944f $X=2.375 $Y=1.765 $X2=0
+ $Y2=0
cc_167 N_B2_M1005_g N_A_397_74#_c_374_n 0.0103661f $X=2.41 $Y=0.74 $X2=0 $Y2=0
cc_168 B2 N_A_397_74#_c_374_n 0.0301911f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_169 N_B2_M1005_g N_A_397_74#_c_375_n 6.28666e-19 $X=2.41 $Y=0.74 $X2=0 $Y2=0
cc_170 N_B2_c_208_n N_A_397_74#_c_376_n 0.0027215f $X=2.375 $Y=1.765 $X2=0 $Y2=0
cc_171 N_B2_M1005_g N_A_397_74#_c_376_n 0.0112613f $X=2.41 $Y=0.74 $X2=0 $Y2=0
cc_172 B2 N_A_397_74#_c_376_n 0.0124003f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_173 N_B1_c_244_n N_VPWR_c_272_n 0.0280207f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_174 N_B1_c_245_n N_VPWR_c_272_n 0.0222392f $X=3.09 $Y=1.465 $X2=0 $Y2=0
cc_175 N_B1_c_244_n N_VPWR_c_273_n 0.00461464f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_176 N_B1_c_244_n N_VPWR_c_266_n 0.00912792f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_177 N_B1_c_244_n N_Y_c_316_n 0.00480438f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_178 N_B1_M1000_g N_VGND_c_341_n 0.00287356f $X=2.84 $Y=0.74 $X2=0 $Y2=0
cc_179 N_B1_M1000_g N_VGND_c_344_n 0.00434272f $X=2.84 $Y=0.74 $X2=0 $Y2=0
cc_180 N_B1_M1000_g N_VGND_c_345_n 0.00824122f $X=2.84 $Y=0.74 $X2=0 $Y2=0
cc_181 N_B1_M1000_g N_A_397_74#_c_374_n 0.0169352f $X=2.84 $Y=0.74 $X2=0 $Y2=0
cc_182 N_B1_c_244_n N_A_397_74#_c_374_n 0.00285817f $X=2.855 $Y=1.765 $X2=0
+ $Y2=0
cc_183 N_B1_c_245_n N_A_397_74#_c_374_n 0.025569f $X=3.09 $Y=1.465 $X2=0 $Y2=0
cc_184 N_B1_M1000_g N_A_397_74#_c_375_n 0.00930389f $X=2.84 $Y=0.74 $X2=0 $Y2=0
cc_185 N_B1_M1000_g N_A_397_74#_c_376_n 6.10655e-19 $X=2.84 $Y=0.74 $X2=0 $Y2=0
cc_186 N_VPWR_c_270_n N_Y_c_316_n 0.0830951f $X=1.415 $Y=2.06 $X2=0 $Y2=0
cc_187 N_VPWR_c_273_n Y 0.0197559f $X=2.995 $Y=3.33 $X2=0 $Y2=0
cc_188 N_VPWR_c_266_n Y 0.0159928f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_189 N_Y_c_304_n N_VGND_c_342_n 0.0109704f $X=1.695 $Y=0.515 $X2=0 $Y2=0
cc_190 N_Y_c_304_n N_VGND_c_345_n 0.00903439f $X=1.695 $Y=0.515 $X2=0 $Y2=0
cc_191 N_Y_c_304_n N_A_397_74#_c_376_n 0.00748774f $X=1.695 $Y=0.515 $X2=0 $Y2=0
cc_192 N_Y_c_305_n N_A_397_74#_c_376_n 0.00622738f $X=1.945 $Y=1.095 $X2=0 $Y2=0
cc_193 N_VGND_M1005_d N_A_397_74#_c_374_n 0.00176461f $X=2.485 $Y=0.37 $X2=0
+ $Y2=0
cc_194 N_VGND_c_341_n N_A_397_74#_c_374_n 0.0135055f $X=2.625 $Y=0.57 $X2=0
+ $Y2=0
cc_195 N_VGND_c_341_n N_A_397_74#_c_375_n 0.0164567f $X=2.625 $Y=0.57 $X2=0
+ $Y2=0
cc_196 N_VGND_c_344_n N_A_397_74#_c_375_n 0.0145639f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_197 N_VGND_c_345_n N_A_397_74#_c_375_n 0.0119984f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_198 N_VGND_c_342_n N_A_397_74#_c_376_n 0.00934777f $X=2.54 $Y=0 $X2=0 $Y2=0
cc_199 N_VGND_c_345_n N_A_397_74#_c_376_n 0.0115074f $X=3.12 $Y=0 $X2=0 $Y2=0
