* File: sky130_fd_sc_ls__o32ai_2.spice
* Created: Fri Aug 28 13:54:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__o32ai_2.pex.spice"
.subckt sky130_fd_sc_ls__o32ai_2  VNB VPB B2 B1 A3 A2 A1 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A1	A1
* A2	A2
* A3	A3
* B1	B1
* B2	B2
* VPB	VPB
* VNB	VNB
MM1015 N_Y_M1015_d N_B2_M1015_g N_A_27_74#_M1015_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75005.5 A=0.111 P=1.78 MULT=1
MM1016 N_Y_M1015_d N_B2_M1016_g N_A_27_74#_M1016_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75000.6
+ SB=75005 A=0.111 P=1.78 MULT=1
MM1009 N_A_27_74#_M1016_s N_B1_M1009_g N_Y_M1009_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1295 AS=0.1295 PD=1.09 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.1
+ SB=75004.5 A=0.111 P=1.78 MULT=1
MM1012 N_A_27_74#_M1012_d N_B1_M1012_g N_Y_M1009_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1295 AS=0.1295 PD=1.09 PS=1.09 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75001.6
+ SB=75004 A=0.111 P=1.78 MULT=1
MM1005 N_VGND_M1005_d N_A3_M1005_g N_A_27_74#_M1012_d VNB NSHORT L=0.15 W=0.74
+ AD=0.2993 AS=0.1295 PD=1.6 PS=1.09 NRD=56.664 NRS=0 M=1 R=4.93333 SA=75002.1
+ SB=75003.5 A=0.111 P=1.78 MULT=1
MM1006 N_VGND_M1005_d N_A3_M1006_g N_A_27_74#_M1006_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2993 AS=0.12765 PD=1.6 PS=1.085 NRD=56.664 NRS=0 M=1 R=4.93333 SA=75003
+ SB=75002.7 A=0.111 P=1.78 MULT=1
MM1013 N_VGND_M1013_d N_A2_M1013_g N_A_27_74#_M1006_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1221 AS=0.12765 PD=1.07 PS=1.085 NRD=0.804 NRS=10.536 M=1 R=4.93333
+ SA=75003.5 SB=75002.2 A=0.111 P=1.78 MULT=1
MM1017 N_VGND_M1013_d N_A2_M1017_g N_A_27_74#_M1017_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1221 AS=0.11285 PD=1.07 PS=1.045 NRD=7.296 NRS=4.044 M=1 R=4.93333
+ SA=75003.9 SB=75001.7 A=0.111 P=1.78 MULT=1
MM1003 N_A_27_74#_M1017_s N_A1_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.74
+ AD=0.11285 AS=0.3367 PD=1.045 PS=1.65 NRD=0 NRS=0 M=1 R=4.93333 SA=75004.4
+ SB=75001.3 A=0.111 P=1.78 MULT=1
MM1010 N_A_27_74#_M1010_d N_A1_M1010_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.3367 PD=2.05 PS=1.65 NRD=0 NRS=0 M=1 R=4.93333 SA=75005.5
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1007 N_Y_M1007_d N_B2_M1007_g N_A_27_368#_M1007_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1008 N_Y_M1007_d N_B2_M1008_g N_A_27_368#_M1008_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1001 N_A_27_368#_M1008_s N_B1_M1001_g N_VPWR_M1001_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1014 N_A_27_368#_M1014_d N_B1_M1014_g N_VPWR_M1001_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.6 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1002 N_Y_M1002_d N_A3_M1002_g N_A_499_368#_M1002_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1004 N_Y_M1002_d N_A3_M1004_g N_A_499_368#_M1004_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1011 N_A_768_368#_M1011_d N_A2_M1011_g N_A_499_368#_M1004_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1019 N_A_768_368#_M1011_d N_A2_M1019_g N_A_499_368#_M1019_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.6 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1000 N_VPWR_M1000_d N_A1_M1000_g N_A_768_368#_M1000_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.3864 AS=0.1708 PD=2.93 PS=1.425 NRD=10.5395 NRS=1.7533 M=1
+ R=7.46667 SA=75000.3 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1018 N_VPWR_M1018_d N_A1_M1018_g N_A_768_368#_M1000_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.3304 AS=0.1708 PD=2.83 PS=1.425 NRD=1.7533 NRS=2.6201 M=1
+ R=7.46667 SA=75000.7 SB=75000.2 A=0.168 P=2.54 MULT=1
DX20_noxref VNB VPB NWDIODE A=12.3132 P=16.96
*
.include "sky130_fd_sc_ls__o32ai_2.pxi.spice"
*
.ends
*
*
