* File: sky130_fd_sc_ls__dfsbp_1.pex.spice
* Created: Wed Sep  2 11:01:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__DFSBP_1%D 2 4 7 9 11 12 13 17 18 21
c33 18 0 8.91633e-20 $X=0.64 $Y=1.175
r34 21 23 39.7991 $w=3.9e-07 $l=1.65e-07 $layer=POLY_cond $X=0.61 $Y=1.855
+ $X2=0.61 $Y2=2.02
r35 21 22 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.64
+ $Y=1.855 $X2=0.64 $Y2=1.855
r36 17 19 45.456 $w=3.9e-07 $l=1.65e-07 $layer=POLY_cond $X=0.61 $Y=1.175
+ $X2=0.61 $Y2=1.01
r37 17 18 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.64
+ $Y=1.175 $X2=0.64 $Y2=1.175
r38 13 22 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=0.64 $Y=1.665
+ $X2=0.64 $Y2=1.855
r39 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.64 $Y=1.295
+ $X2=0.64 $Y2=1.665
r40 12 18 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=0.64 $Y=1.295
+ $X2=0.64 $Y2=1.175
r41 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.505 $Y=2.465
+ $X2=0.505 $Y2=2.75
r42 7 19 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=0.495 $Y=0.61 $X2=0.495
+ $Y2=1.01
r43 4 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.505 $Y=2.375 $X2=0.505
+ $Y2=2.465
r44 4 23 137.992 $w=1.8e-07 $l=3.55e-07 $layer=POLY_cond $X=0.505 $Y=2.375
+ $X2=0.505 $Y2=2.02
r45 2 21 4.27811 $w=3.9e-07 $l=3e-08 $layer=POLY_cond $X=0.61 $Y=1.825 $X2=0.61
+ $Y2=1.855
r46 1 17 4.27811 $w=3.9e-07 $l=3e-08 $layer=POLY_cond $X=0.61 $Y=1.205 $X2=0.61
+ $Y2=1.175
r47 1 2 88.4142 $w=3.9e-07 $l=6.2e-07 $layer=POLY_cond $X=0.61 $Y=1.205 $X2=0.61
+ $Y2=1.825
.ends

.subckt PM_SKY130_FD_SC_LS__DFSBP_1%CLK 1 3 4 6 7
c33 4 0 2.28976e-19 $X=1.515 $Y=1.715
r34 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.465
+ $Y=1.385 $X2=1.465 $Y2=1.385
r35 7 11 6.69663 $w=3.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.68 $Y=1.365
+ $X2=1.465 $Y2=1.365
r36 4 10 67.1335 $w=2.8e-07 $l=3.54119e-07 $layer=POLY_cond $X=1.515 $Y=1.715
+ $X2=1.465 $Y2=1.385
r37 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.515 $Y=1.715
+ $X2=1.515 $Y2=2.35
r38 1 10 38.7299 $w=2.8e-07 $l=1.74714e-07 $layer=POLY_cond $X=1.485 $Y=1.22
+ $X2=1.465 $Y2=1.385
r39 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.485 $Y=1.22 $X2=1.485
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__DFSBP_1%A_398_74# 1 2 7 8 9 11 16 20 21 23 26 30 32
+ 33 34 35 38 45 46 49 50 53 54 55 57 58 59 61 62 63 65 67 68 69 72 73 77 78 81
+ 83 87 91
c296 81 0 1.19048e-19 $X=7.395 $Y=2.185
c297 73 0 1.69669e-19 $X=3.825 $Y=2.25
c298 63 0 2.3488e-20 $X=6.035 $Y=1.705
c299 62 0 1.57368e-19 $X=6.435 $Y=1.705
c300 59 0 1.41158e-19 $X=5.54 $Y=2.21
c301 32 0 8.72473e-20 $X=3.025 $Y=0.34
c302 8 0 1.32821e-19 $X=3.03 $Y=1.94
r303 86 87 16.2455 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=3.665 $Y=1.525
+ $X2=3.59 $Y2=1.525
r304 81 83 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.395 $Y=2.185
+ $X2=7.395 $Y2=2.02
r305 81 82 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.395
+ $Y=2.185 $X2=7.395 $Y2=2.185
r306 78 91 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.715 $Y=1.285
+ $X2=6.715 $Y2=1.12
r307 77 78 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.715
+ $Y=1.285 $X2=6.715 $Y2=1.285
r308 74 77 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=6.52 $Y=1.285
+ $X2=6.715 $Y2=1.285
r309 70 83 104.059 $w=1.68e-07 $l=1.595e-06 $layer=LI1_cond $X=7.475 $Y=0.425
+ $X2=7.475 $Y2=2.02
r310 68 70 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.39 $Y=0.34
+ $X2=7.475 $Y2=0.425
r311 68 69 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=7.39 $Y=0.34
+ $X2=6.605 $Y2=0.34
r312 66 74 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.52 $Y=1.45
+ $X2=6.52 $Y2=1.285
r313 66 67 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=6.52 $Y=1.45
+ $X2=6.52 $Y2=1.62
r314 65 74 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.52 $Y=1.12
+ $X2=6.52 $Y2=1.285
r315 64 69 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.52 $Y=0.425
+ $X2=6.605 $Y2=0.34
r316 64 65 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=6.52 $Y=0.425
+ $X2=6.52 $Y2=1.12
r317 62 67 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.435 $Y=1.705
+ $X2=6.52 $Y2=1.62
r318 62 63 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=6.435 $Y=1.705
+ $X2=6.035 $Y2=1.705
r319 60 63 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.95 $Y=1.79
+ $X2=6.035 $Y2=1.705
r320 60 61 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=5.95 $Y=1.79
+ $X2=5.95 $Y2=2.125
r321 58 61 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.865 $Y=2.21
+ $X2=5.95 $Y2=2.125
r322 58 59 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=5.865 $Y=2.21
+ $X2=5.54 $Y2=2.21
r323 56 59 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.455 $Y=2.295
+ $X2=5.54 $Y2=2.21
r324 56 57 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=5.455 $Y=2.295
+ $X2=5.455 $Y2=2.905
r325 54 57 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.37 $Y=2.99
+ $X2=5.455 $Y2=2.905
r326 54 55 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=5.37 $Y=2.99
+ $X2=4.78 $Y2=2.99
r327 53 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.695 $Y=2.905
+ $X2=4.78 $Y2=2.99
r328 52 53 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=4.695 $Y=2.335
+ $X2=4.695 $Y2=2.905
r329 51 73 2.0246 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=3.945 $Y=2.25
+ $X2=3.825 $Y2=2.25
r330 50 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.61 $Y=2.25
+ $X2=4.695 $Y2=2.335
r331 50 51 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=4.61 $Y=2.25
+ $X2=3.945 $Y2=2.25
r332 48 73 4.40882 $w=2.05e-07 $l=1.00995e-07 $layer=LI1_cond $X=3.79 $Y=2.335
+ $X2=3.825 $Y2=2.25
r333 48 49 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=3.79 $Y=2.335
+ $X2=3.79 $Y2=2.905
r334 46 86 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=3.825 $Y=1.525
+ $X2=3.665 $Y2=1.525
r335 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.825
+ $Y=1.525 $X2=3.825 $Y2=1.525
r336 43 73 4.40882 $w=2.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.825 $Y=2.165
+ $X2=3.825 $Y2=2.25
r337 43 45 30.7318 $w=2.38e-07 $l=6.4e-07 $layer=LI1_cond $X=3.825 $Y=2.165
+ $X2=3.825 $Y2=1.525
r338 41 72 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=3.11 $Y=0.425
+ $X2=3.11 $Y2=1.435
r339 38 72 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.03 $Y=1.6
+ $X2=3.03 $Y2=1.435
r340 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.03
+ $Y=1.6 $X2=3.03 $Y2=1.6
r341 34 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.705 $Y=2.99
+ $X2=3.79 $Y2=2.905
r342 34 35 88.0749 $w=1.68e-07 $l=1.35e-06 $layer=LI1_cond $X=3.705 $Y=2.99
+ $X2=2.355 $Y2=2.99
r343 32 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.025 $Y=0.34
+ $X2=3.11 $Y2=0.425
r344 32 33 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=3.025 $Y=0.34
+ $X2=2.295 $Y2=0.34
r345 28 35 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.23 $Y=2.905
+ $X2=2.355 $Y2=2.99
r346 28 30 15.6732 $w=2.48e-07 $l=3.4e-07 $layer=LI1_cond $X=2.23 $Y=2.905
+ $X2=2.23 $Y2=2.565
r347 24 33 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.17 $Y=0.425
+ $X2=2.295 $Y2=0.34
r348 24 26 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=2.17 $Y=0.425
+ $X2=2.17 $Y2=0.515
r349 21 82 56.7725 $w=3.04e-07 $l=3.24037e-07 $layer=POLY_cond $X=7.51 $Y=2.465
+ $X2=7.415 $Y2=2.185
r350 21 23 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.51 $Y=2.465
+ $X2=7.51 $Y2=2.75
r351 20 91 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=6.725 $Y=0.69
+ $X2=6.725 $Y2=1.12
r352 14 86 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.665 $Y=1.36
+ $X2=3.665 $Y2=1.525
r353 14 16 382.011 $w=1.5e-07 $l=7.45e-07 $layer=POLY_cond $X=3.665 $Y=1.36
+ $X2=3.665 $Y2=0.615
r354 13 39 15.4923 $w=2.55e-07 $l=1.65e-07 $layer=POLY_cond $X=3.195 $Y=1.562
+ $X2=3.03 $Y2=1.562
r355 13 87 96.2149 $w=2.55e-07 $l=3.95e-07 $layer=POLY_cond $X=3.195 $Y=1.562
+ $X2=3.59 $Y2=1.562
r356 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.065 $Y=2.24
+ $X2=3.065 $Y2=2.525
r357 8 9 55.1908 $w=2.62e-07 $l=3.17017e-07 $layer=POLY_cond $X=3.03 $Y=1.94
+ $X2=3.065 $Y2=2.24
r358 7 39 12.0182 $w=3.3e-07 $l=1.28e-07 $layer=POLY_cond $X=3.03 $Y=1.69
+ $X2=3.03 $Y2=1.562
r359 7 8 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=3.03 $Y=1.69 $X2=3.03
+ $Y2=1.94
r360 2 30 600 $w=1.7e-07 $l=8.46685e-07 $layer=licon1_PDIFF $count=1 $X=2.04
+ $Y=1.79 $X2=2.19 $Y2=2.565
r361 1 26 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.99
+ $Y=0.37 $X2=2.13 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__DFSBP_1%A_779_380# 1 2 7 9 10 12 13 15 16 19 21 24
+ 28 31 36 39
c91 36 0 9.58642e-20 $X=4.395 $Y=1.72
c92 21 0 1.31064e-19 $X=4.95 $Y=1.885
c93 7 0 7.37914e-20 $X=3.985 $Y=2.24
r94 36 42 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=4.485 $Y=1.72
+ $X2=4.485 $Y2=1.265
r95 34 42 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.575 $Y=1.1
+ $X2=4.575 $Y2=1.265
r96 34 39 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.575 $Y=1.1 $X2=4.575
+ $Y2=1.01
r97 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.575
+ $Y=1.1 $X2=4.575 $Y2=1.1
r98 31 33 13.3188 $w=4.58e-07 $l=6.09098e-07 $layer=LI1_cond $X=4.817 $Y=0.6
+ $X2=4.575 $Y2=1.1
r99 26 28 23.9708 $w=2.48e-07 $l=5.2e-07 $layer=LI1_cond $X=5.075 $Y=1.995
+ $X2=5.075 $Y2=2.515
r100 24 37 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.395 $Y=1.885
+ $X2=4.395 $Y2=1.975
r101 24 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.395 $Y=1.885
+ $X2=4.395 $Y2=1.72
r102 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.395
+ $Y=1.885 $X2=4.395 $Y2=1.885
r103 21 26 6.85268 $w=2.2e-07 $l=1.71391e-07 $layer=LI1_cond $X=4.95 $Y=1.885
+ $X2=5.075 $Y2=1.995
r104 21 23 29.073 $w=2.18e-07 $l=5.55e-07 $layer=LI1_cond $X=4.95 $Y=1.885
+ $X2=4.395 $Y2=1.885
r105 15 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.41 $Y=1.01
+ $X2=4.575 $Y2=1.01
r106 15 16 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=4.41 $Y=1.01
+ $X2=4.13 $Y2=1.01
r107 14 19 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.075 $Y=1.975
+ $X2=3.985 $Y2=1.975
r108 13 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.23 $Y=1.975
+ $X2=4.395 $Y2=1.975
r109 13 14 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=4.23 $Y=1.975
+ $X2=4.075 $Y2=1.975
r110 10 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.055 $Y=0.935
+ $X2=4.13 $Y2=1.01
r111 10 12 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.055 $Y=0.935
+ $X2=4.055 $Y2=0.615
r112 7 19 105.158 $w=1.8e-07 $l=2.65e-07 $layer=POLY_cond $X=3.985 $Y=2.24
+ $X2=3.985 $Y2=1.975
r113 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.985 $Y=2.24
+ $X2=3.985 $Y2=2.525
r114 2 28 600 $w=1.7e-07 $l=2.64575e-07 $layer=licon1_PDIFF $count=1 $X=4.965
+ $Y=2.315 $X2=5.115 $Y2=2.515
r115 1 31 182 $w=1.7e-07 $l=2.85745e-07 $layer=licon1_NDIFF $count=1 $X=4.89
+ $Y=0.37 $X2=5.015 $Y2=0.6
.ends

.subckt PM_SKY130_FD_SC_LS__DFSBP_1%A_596_81# 1 2 8 9 11 13 16 18 20 21 23 26 30
+ 34 37 38 39 40 41 42 45 46 48 52 61
c162 46 0 7.37914e-20 $X=3.355 $Y=2.295
c163 45 0 1.32821e-19 $X=3.34 $Y=2.515
c164 40 0 9.58642e-20 $X=5.092 $Y=1.29
c165 13 0 1.19393e-19 $X=5.025 $Y=1.57
c166 9 0 4.58062e-20 $X=4.89 $Y=2.24
c167 8 0 9.5352e-20 $X=4.89 $Y=2.15
r168 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.1
+ $Y=1.285 $X2=6.1 $Y2=1.285
r169 52 55 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=6.1 $Y=1.205 $X2=6.1
+ $Y2=1.285
r170 51 61 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=5.115 $Y=1.22
+ $X2=5.23 $Y2=1.22
r171 51 58 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.115 $Y=1.22
+ $X2=5.025 $Y2=1.22
r172 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.115
+ $Y=1.22 $X2=5.115 $Y2=1.22
r173 45 46 10.2717 $w=3.58e-07 $l=2.2e-07 $layer=LI1_cond $X=3.355 $Y=2.515
+ $X2=3.355 $Y2=2.295
r174 43 50 4.42914 $w=1.7e-07 $l=1.58644e-07 $layer=LI1_cond $X=5.235 $Y=1.205
+ $X2=5.092 $Y2=1.172
r175 42 52 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.935 $Y=1.205
+ $X2=6.1 $Y2=1.205
r176 42 43 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=5.935 $Y=1.205
+ $X2=5.235 $Y2=1.205
r177 40 50 2.96953 $w=2.85e-07 $l=1.18e-07 $layer=LI1_cond $X=5.092 $Y=1.29
+ $X2=5.092 $Y2=1.172
r178 40 41 5.86331 $w=2.83e-07 $l=1.45e-07 $layer=LI1_cond $X=5.092 $Y=1.29
+ $X2=5.092 $Y2=1.435
r179 38 41 7.39867 $w=1.7e-07 $l=1.79538e-07 $layer=LI1_cond $X=4.95 $Y=1.52
+ $X2=5.092 $Y2=1.435
r180 38 39 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=4.95 $Y=1.52
+ $X2=4.285 $Y2=1.52
r181 37 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.2 $Y=1.435
+ $X2=4.285 $Y2=1.52
r182 36 37 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=4.2 $Y=1.055
+ $X2=4.2 $Y2=1.435
r183 35 48 2.11342 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.615 $Y=0.97
+ $X2=3.49 $Y2=0.97
r184 34 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.115 $Y=0.97
+ $X2=4.2 $Y2=1.055
r185 34 35 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=4.115 $Y=0.97
+ $X2=3.615 $Y2=0.97
r186 32 48 4.3182 $w=2.1e-07 $l=1.03078e-07 $layer=LI1_cond $X=3.45 $Y=1.055
+ $X2=3.49 $Y2=0.97
r187 32 46 80.8984 $w=1.68e-07 $l=1.24e-06 $layer=LI1_cond $X=3.45 $Y=1.055
+ $X2=3.45 $Y2=2.295
r188 28 48 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.49 $Y=0.885
+ $X2=3.49 $Y2=0.97
r189 28 30 12.4464 $w=2.48e-07 $l=2.7e-07 $layer=LI1_cond $X=3.49 $Y=0.885
+ $X2=3.49 $Y2=0.615
r190 21 56 38.535 $w=3.06e-07 $l=2.14173e-07 $layer=POLY_cond $X=6.235 $Y=1.12
+ $X2=6.122 $Y2=1.285
r191 21 23 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=6.235 $Y=1.12
+ $X2=6.235 $Y2=0.69
r192 18 56 66.888 $w=3.06e-07 $l=3.7975e-07 $layer=POLY_cond $X=6.195 $Y=1.63
+ $X2=6.122 $Y2=1.285
r193 18 20 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.195 $Y=1.63
+ $X2=6.195 $Y2=2.205
r194 14 61 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.23 $Y=1.055
+ $X2=5.23 $Y2=1.22
r195 14 16 243.564 $w=1.5e-07 $l=4.75e-07 $layer=POLY_cond $X=5.23 $Y=1.055
+ $X2=5.23 $Y2=0.58
r196 13 26 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.025 $Y=1.57
+ $X2=5.025 $Y2=1.645
r197 12 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.025 $Y=1.385
+ $X2=5.025 $Y2=1.22
r198 12 13 94.8617 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=5.025 $Y=1.385
+ $X2=5.025 $Y2=1.57
r199 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.89 $Y=2.24 $X2=4.89
+ $Y2=2.525
r200 8 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=4.89 $Y=2.15 $X2=4.89
+ $Y2=2.24
r201 7 26 69.2234 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.89 $Y=1.645
+ $X2=5.025 $Y2=1.645
r202 7 8 167.145 $w=1.8e-07 $l=4.3e-07 $layer=POLY_cond $X=4.89 $Y=1.72 $X2=4.89
+ $Y2=2.15
r203 2 45 600 $w=1.7e-07 $l=2.82843e-07 $layer=licon1_PDIFF $count=1 $X=3.14
+ $Y=2.315 $X2=3.34 $Y2=2.515
r204 1 30 182 $w=1.7e-07 $l=5.65332e-07 $layer=licon1_NDIFF $count=1 $X=2.98
+ $Y=0.405 $X2=3.45 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_LS__DFSBP_1%SET_B 2 3 5 8 12 14 15 16 18 20 21 22 25 27
+ 34 36 40
c148 25 0 1.19393e-19 $X=5.52 $Y=1.665
c149 22 0 1.31064e-19 $X=5.665 $Y=1.665
c150 21 0 1.03271e-19 $X=8.255 $Y=1.665
c151 15 0 2.58188e-20 $X=8.09 $Y=1.3
r152 40 48 8.23174 $w=3.83e-07 $l=2.75e-07 $layer=LI1_cond $X=8.477 $Y=1.39
+ $X2=8.477 $Y2=1.665
r153 39 41 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.505 $Y=1.39
+ $X2=8.505 $Y2=1.555
r154 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.505
+ $Y=1.39 $X2=8.505 $Y2=1.39
r155 36 39 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=8.505 $Y=1.3
+ $X2=8.505 $Y2=1.39
r156 32 34 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.53 $Y=1.79 $X2=5.62
+ $Y2=1.79
r157 29 32 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=5.4 $Y=1.79 $X2=5.53
+ $Y2=1.79
r158 27 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=1.665
+ $X2=8.4 $Y2=1.665
r159 25 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.53
+ $Y=1.79 $X2=5.53 $Y2=1.79
r160 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=1.665
+ $X2=5.52 $Y2=1.665
r161 22 24 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.665 $Y=1.665
+ $X2=5.52 $Y2=1.665
r162 21 27 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.255 $Y=1.665
+ $X2=8.4 $Y2=1.665
r163 21 22 3.20544 $w=1.4e-07 $l=2.59e-06 $layer=MET1_cond $X=8.255 $Y=1.665
+ $X2=5.665 $Y2=1.665
r164 20 41 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=8.415 $Y=2.155
+ $X2=8.415 $Y2=1.555
r165 16 20 79.0582 $w=1.89e-07 $l=3.27032e-07 $layer=POLY_cond $X=8.38 $Y=2.465
+ $X2=8.415 $Y2=2.155
r166 16 18 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=8.38 $Y=2.465
+ $X2=8.38 $Y2=2.75
r167 14 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.34 $Y=1.3
+ $X2=8.505 $Y2=1.3
r168 14 15 128.191 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=8.34 $Y=1.3
+ $X2=8.09 $Y2=1.3
r169 10 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.015 $Y=1.225
+ $X2=8.09 $Y2=1.3
r170 10 12 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=8.015 $Y=1.225
+ $X2=8.015 $Y2=0.58
r171 6 34 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.62 $Y=1.625
+ $X2=5.62 $Y2=1.79
r172 6 8 535.84 $w=1.5e-07 $l=1.045e-06 $layer=POLY_cond $X=5.62 $Y=1.625
+ $X2=5.62 $Y2=0.58
r173 3 5 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=5.4 $Y=2.24 $X2=5.4
+ $Y2=2.525
r174 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.4 $Y=2.15 $X2=5.4
+ $Y2=2.24
r175 1 29 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.4 $Y=1.955
+ $X2=5.4 $Y2=1.79
r176 1 2 75.7984 $w=1.8e-07 $l=1.95e-07 $layer=POLY_cond $X=5.4 $Y=1.955 $X2=5.4
+ $Y2=2.15
.ends

.subckt PM_SKY130_FD_SC_LS__DFSBP_1%A_225_74# 1 2 9 11 13 15 16 18 19 22 24 25
+ 26 28 29 34 35 36 39 43 46 47 48 51 52 53 56 60 64 67
c180 56 0 2.99812e-20 $X=2.025 $Y=1.805
c181 39 0 1.57368e-19 $X=7.235 $Y=0.58
c182 34 0 1.19048e-19 $X=6.7 $Y=2.385
c183 26 0 1.22627e-19 $X=3.565 $Y=2.81
c184 16 0 8.72473e-20 $X=2.83 $Y=1.12
r185 64 66 17.8607 $w=4.58e-07 $l=4.95e-07 $layer=LI1_cond $X=1.205 $Y=0.515
+ $X2=1.205 $Y2=1.01
r186 60 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.19
+ $Y=1.465 $X2=2.19 $Y2=1.465
r187 58 60 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=2.19 $Y=1.72
+ $X2=2.19 $Y2=1.465
r188 56 58 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.025 $Y=1.805
+ $X2=2.19 $Y2=1.72
r189 56 67 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=2.025 $Y=1.805
+ $X2=1.455 $Y2=1.805
r190 53 55 5.57014 $w=2.98e-07 $l=1.45e-07 $layer=LI1_cond $X=1.145 $Y=1.87
+ $X2=1.29 $Y2=1.87
r191 52 67 7.90841 $w=2.98e-07 $l=1.5e-07 $layer=LI1_cond $X=1.305 $Y=1.87
+ $X2=1.455 $Y2=1.87
r192 52 55 0.576222 $w=2.98e-07 $l=1.5e-08 $layer=LI1_cond $X=1.305 $Y=1.87
+ $X2=1.29 $Y2=1.87
r193 51 53 7.51767 $w=3e-07 $l=1.8775e-07 $layer=LI1_cond $X=1.06 $Y=1.72
+ $X2=1.145 $Y2=1.87
r194 51 66 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=1.06 $Y=1.72
+ $X2=1.06 $Y2=1.01
r195 46 61 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=2.41 $Y=1.465
+ $X2=2.19 $Y2=1.465
r196 43 46 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=2.485 $Y=1.12
+ $X2=2.485 $Y2=1.465
r197 42 61 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=2.055 $Y=1.465
+ $X2=2.19 $Y2=1.465
r198 37 39 553.787 $w=1.5e-07 $l=1.08e-06 $layer=POLY_cond $X=7.235 $Y=1.66
+ $X2=7.235 $Y2=0.58
r199 35 37 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.16 $Y=1.735
+ $X2=7.235 $Y2=1.66
r200 35 36 197.415 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=7.16 $Y=1.735
+ $X2=6.775 $Y2=1.735
r201 32 48 76.0046 $w=1.8e-07 $l=1.9e-07 $layer=POLY_cond $X=6.7 $Y=2.96 $X2=6.7
+ $Y2=3.15
r202 32 34 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.7 $Y=2.96 $X2=6.7
+ $Y2=2.385
r203 31 36 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.7 $Y=1.81
+ $X2=6.775 $Y2=1.735
r204 31 34 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.7 $Y=1.81 $X2=6.7
+ $Y2=2.385
r205 30 47 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.655 $Y=3.15
+ $X2=3.565 $Y2=3.15
r206 29 48 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=6.61 $Y=3.15 $X2=6.7
+ $Y2=3.15
r207 29 30 1515.22 $w=1.5e-07 $l=2.955e-06 $layer=POLY_cond $X=6.61 $Y=3.15
+ $X2=3.655 $Y2=3.15
r208 26 28 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.565 $Y=2.81
+ $X2=3.565 $Y2=2.525
r209 25 47 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=3.565 $Y=3.075
+ $X2=3.565 $Y2=3.15
r210 24 26 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.565 $Y=2.9
+ $X2=3.565 $Y2=2.81
r211 24 25 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=3.565 $Y=2.9
+ $X2=3.565 $Y2=3.075
r212 20 22 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.905 $Y=1.045
+ $X2=2.905 $Y2=0.615
r213 18 47 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.475 $Y=3.15
+ $X2=3.565 $Y2=3.15
r214 18 19 469.181 $w=1.5e-07 $l=9.15e-07 $layer=POLY_cond $X=3.475 $Y=3.15
+ $X2=2.56 $Y2=3.15
r215 17 43 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.56 $Y=1.12
+ $X2=2.485 $Y2=1.12
r216 16 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.83 $Y=1.12
+ $X2=2.905 $Y2=1.045
r217 16 17 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.83 $Y=1.12
+ $X2=2.56 $Y2=1.12
r218 15 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.485 $Y=3.075
+ $X2=2.56 $Y2=3.15
r219 14 46 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.485 $Y=1.63
+ $X2=2.485 $Y2=1.465
r220 14 15 740.947 $w=1.5e-07 $l=1.445e-06 $layer=POLY_cond $X=2.485 $Y=1.63
+ $X2=2.485 $Y2=3.075
r221 11 42 65.1975 $w=1.92e-07 $l=2.58844e-07 $layer=POLY_cond $X=1.965 $Y=1.715
+ $X2=1.947 $Y2=1.465
r222 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.965 $Y=1.715
+ $X2=1.965 $Y2=2.35
r223 7 42 43.8589 $w=1.92e-07 $l=1.80291e-07 $layer=POLY_cond $X=1.915 $Y=1.3
+ $X2=1.947 $Y2=1.465
r224 7 9 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.915 $Y=1.3
+ $X2=1.915 $Y2=0.74
r225 2 55 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.145
+ $Y=1.79 $X2=1.29 $Y2=1.935
r226 1 64 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=1.125
+ $Y=0.37 $X2=1.27 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__DFSBP_1%A_1510_48# 1 2 9 12 13 15 18 21 22 25 29 31
+ 33 34 36 37 39
c121 39 0 7.00183e-20 $X=7.93 $Y=1.75
r122 35 36 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=9.65 $Y=1.01
+ $X2=9.65 $Y2=2.39
r123 33 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.565 $Y=2.475
+ $X2=9.65 $Y2=2.39
r124 33 34 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=9.565 $Y=2.475
+ $X2=9.33 $Y2=2.475
r125 32 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.255 $Y=0.925
+ $X2=9.09 $Y2=0.925
r126 31 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.565 $Y=0.925
+ $X2=9.65 $Y2=1.01
r127 31 32 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=9.565 $Y=0.925
+ $X2=9.255 $Y2=0.925
r128 27 34 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.165 $Y=2.56
+ $X2=9.33 $Y2=2.475
r129 27 29 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=9.165 $Y=2.56
+ $X2=9.165 $Y2=2.75
r130 23 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.09 $Y=0.84
+ $X2=9.09 $Y2=0.925
r131 23 25 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=9.09 $Y=0.84
+ $X2=9.09 $Y2=0.58
r132 21 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.925 $Y=0.925
+ $X2=9.09 $Y2=0.925
r133 21 22 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=8.925 $Y=0.925
+ $X2=8.1 $Y2=0.925
r134 19 39 0.934109 $w=2.58e-07 $l=5e-09 $layer=POLY_cond $X=7.935 $Y=1.75
+ $X2=7.93 $Y2=1.75
r135 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.935
+ $Y=1.75 $X2=7.935 $Y2=1.75
r136 16 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.935 $Y=1.01
+ $X2=8.1 $Y2=0.925
r137 16 18 25.8427 $w=3.28e-07 $l=7.4e-07 $layer=LI1_cond $X=7.935 $Y=1.01
+ $X2=7.935 $Y2=1.75
r138 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.93 $Y=2.465
+ $X2=7.93 $Y2=2.75
r139 12 13 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=7.93 $Y=2.375
+ $X2=7.93 $Y2=2.465
r140 11 39 11.2427 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.93 $Y=1.915
+ $X2=7.93 $Y2=1.75
r141 11 12 178.806 $w=1.8e-07 $l=4.6e-07 $layer=POLY_cond $X=7.93 $Y=1.915
+ $X2=7.93 $Y2=2.375
r142 7 39 56.9806 $w=2.58e-07 $l=3.78616e-07 $layer=POLY_cond $X=7.625 $Y=1.585
+ $X2=7.93 $Y2=1.75
r143 7 9 515.33 $w=1.5e-07 $l=1.005e-06 $layer=POLY_cond $X=7.625 $Y=1.585
+ $X2=7.625 $Y2=0.58
r144 2 29 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=9.02
+ $Y=2.54 $X2=9.165 $Y2=2.75
r145 1 25 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=8.95
+ $Y=0.37 $X2=9.09 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_LS__DFSBP_1%A_1355_377# 1 2 3 10 12 14 16 17 19 20 22 23
+ 25 26 27 30 33 34 36 39 41 44 49 50 51 53 56 60 62 64 66 69 74 78 79 80 81
c200 69 0 7.00183e-20 $X=6.885 $Y=1.882
c201 56 0 2.58188e-20 $X=8.44 $Y=2.265
c202 41 0 1.55237e-19 $X=10.925 $Y=1.41
r203 88 89 5.07963 $w=4.27e-07 $l=4.5e-08 $layer=POLY_cond $X=9.935 $Y=1.487
+ $X2=9.98 $Y2=1.487
r204 83 84 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=9.23
+ $Y=2.055 $X2=9.23 $Y2=2.055
r205 79 80 8.9189 $w=4.28e-07 $l=1.7e-07 $layer=LI1_cond $X=7.73 $Y=2.35 $X2=7.9
+ $Y2=2.35
r206 78 79 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=7.45 $Y=2.565
+ $X2=7.73 $Y2=2.565
r207 77 78 8.76046 $w=4.23e-07 $l=1.65e-07 $layer=LI1_cond $X=7.285 $Y=2.692
+ $X2=7.45 $Y2=2.692
r208 72 74 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=6.94 $Y=0.76
+ $X2=7.135 $Y2=0.76
r209 67 85 10.1593 $w=4.27e-07 $l=9e-08 $layer=POLY_cond $X=9.23 $Y=1.487
+ $X2=9.14 $Y2=1.487
r210 66 67 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=9.23
+ $Y=1.375 $X2=9.23 $Y2=1.375
r211 64 83 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.23 $Y=2.05 $X2=9.23
+ $Y2=2.135
r212 64 66 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=9.23 $Y=2.05
+ $X2=9.23 $Y2=1.375
r213 63 81 5.58832 $w=3e-07 $l=2.20624e-07 $layer=LI1_cond $X=8.77 $Y=2.135
+ $X2=8.605 $Y2=2.265
r214 62 83 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.065 $Y=2.135
+ $X2=9.23 $Y2=2.135
r215 62 63 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=9.065 $Y=2.135
+ $X2=8.77 $Y2=2.135
r216 58 81 1.0017 $w=3.3e-07 $l=2.15e-07 $layer=LI1_cond $X=8.605 $Y=2.48
+ $X2=8.605 $Y2=2.265
r217 58 60 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=8.605 $Y=2.48
+ $X2=8.605 $Y2=2.75
r218 56 81 5.58832 $w=3e-07 $l=1.65e-07 $layer=LI1_cond $X=8.44 $Y=2.265
+ $X2=8.605 $Y2=2.265
r219 56 80 14.4725 $w=4.28e-07 $l=5.4e-07 $layer=LI1_cond $X=8.44 $Y=2.265
+ $X2=7.9 $Y2=2.265
r220 53 69 12.249 $w=2.49e-07 $l=3.36155e-07 $layer=LI1_cond $X=7.135 $Y=1.68
+ $X2=6.885 $Y2=1.882
r221 52 74 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.135 $Y=0.925
+ $X2=7.135 $Y2=0.76
r222 52 53 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=7.135 $Y=0.925
+ $X2=7.135 $Y2=1.68
r223 50 77 1.27447 $w=4.23e-07 $l=4.7e-08 $layer=LI1_cond $X=7.238 $Y=2.692
+ $X2=7.285 $Y2=2.692
r224 50 51 6.18252 $w=4.23e-07 $l=2.28e-07 $layer=LI1_cond $X=7.238 $Y=2.692
+ $X2=7.01 $Y2=2.692
r225 47 51 7.42997 $w=4.25e-07 $l=2.6729e-07 $layer=LI1_cond $X=6.885 $Y=2.48
+ $X2=7.01 $Y2=2.692
r226 47 49 10.1415 $w=2.48e-07 $l=2.2e-07 $layer=LI1_cond $X=6.885 $Y=2.48
+ $X2=6.885 $Y2=2.26
r227 46 69 0.692029 $w=2.5e-07 $l=2.03e-07 $layer=LI1_cond $X=6.885 $Y=2.085
+ $X2=6.885 $Y2=1.882
r228 46 49 8.0671 $w=2.48e-07 $l=1.75e-07 $layer=LI1_cond $X=6.885 $Y=2.085
+ $X2=6.885 $Y2=2.26
r229 42 44 33.3298 $w=1.5e-07 $l=6.5e-08 $layer=POLY_cond $X=10.925 $Y=1.865
+ $X2=10.99 $Y2=1.865
r230 37 39 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=8.875 $Y=0.94
+ $X2=9.14 $Y2=0.94
r231 34 44 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.99 $Y=1.94
+ $X2=10.99 $Y2=1.865
r232 34 36 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=10.99 $Y=1.94
+ $X2=10.99 $Y2=2.435
r233 33 42 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.925 $Y=1.79
+ $X2=10.925 $Y2=1.865
r234 32 41 42.0026 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=10.925 $Y=1.61
+ $X2=10.925 $Y2=1.41
r235 32 33 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=10.925 $Y=1.61
+ $X2=10.925 $Y2=1.79
r236 28 41 42.0026 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=10.925 $Y=1.21
+ $X2=10.925 $Y2=1.41
r237 28 30 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=10.925 $Y=1.21
+ $X2=10.925 $Y2=0.645
r238 27 89 10.4161 $w=4.27e-07 $l=1.22597e-07 $layer=POLY_cond $X=10.07 $Y=1.41
+ $X2=9.98 $Y2=1.487
r239 26 41 7.17539 $w=4e-07 $l=7.5e-08 $layer=POLY_cond $X=10.85 $Y=1.41
+ $X2=10.925 $Y2=1.41
r240 26 27 108.45 $w=4e-07 $l=7.8e-07 $layer=POLY_cond $X=10.85 $Y=1.41
+ $X2=10.07 $Y2=1.41
r241 23 89 27.4666 $w=1.5e-07 $l=2.78e-07 $layer=POLY_cond $X=9.98 $Y=1.765
+ $X2=9.98 $Y2=1.487
r242 23 25 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=9.98 $Y=1.765
+ $X2=9.98 $Y2=2.4
r243 20 88 27.4666 $w=1.5e-07 $l=2.77e-07 $layer=POLY_cond $X=9.935 $Y=1.21
+ $X2=9.935 $Y2=1.487
r244 20 22 151.027 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=9.935 $Y=1.21
+ $X2=9.935 $Y2=0.74
r245 17 84 75.3414 $w=3.21e-07 $l=5.20192e-07 $layer=POLY_cond $X=9.475 $Y=2.465
+ $X2=9.225 $Y2=2.055
r246 17 19 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=9.475 $Y=2.465
+ $X2=9.475 $Y2=2.75
r247 16 84 12.0562 $w=4.7e-07 $l=1.04283e-07 $layer=POLY_cond $X=9.3 $Y=1.985
+ $X2=9.225 $Y2=2.055
r248 15 88 71.6792 $w=4.27e-07 $l=6.35e-07 $layer=POLY_cond $X=9.3 $Y=1.487
+ $X2=9.935 $Y2=1.487
r249 15 67 7.90164 $w=4.27e-07 $l=7e-08 $layer=POLY_cond $X=9.3 $Y=1.487
+ $X2=9.23 $Y2=1.487
r250 15 16 44.374 $w=4.7e-07 $l=3.75e-07 $layer=POLY_cond $X=9.3 $Y=1.61 $X2=9.3
+ $Y2=1.985
r251 14 85 27.4666 $w=1.5e-07 $l=2.77e-07 $layer=POLY_cond $X=9.14 $Y=1.21
+ $X2=9.14 $Y2=1.487
r252 13 39 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.14 $Y=1.015
+ $X2=9.14 $Y2=0.94
r253 13 14 99.9894 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=9.14 $Y=1.015
+ $X2=9.14 $Y2=1.21
r254 10 37 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.875 $Y=0.865
+ $X2=8.875 $Y2=0.94
r255 10 12 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=8.875 $Y=0.865
+ $X2=8.875 $Y2=0.58
r256 3 60 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=8.455
+ $Y=2.54 $X2=8.605 $Y2=2.75
r257 2 77 300 $w=1.7e-07 $l=1.08031e-06 $layer=licon1_PDIFF $count=2 $X=6.775
+ $Y=1.885 $X2=7.285 $Y2=2.74
r258 2 49 600 $w=1.7e-07 $l=4.43706e-07 $layer=licon1_PDIFF $count=1 $X=6.775
+ $Y=1.885 $X2=6.925 $Y2=2.26
r259 1 72 182 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_NDIFF $count=1 $X=6.8
+ $Y=0.37 $X2=6.94 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_LS__DFSBP_1%A_2113_74# 1 2 7 9 10 12 15 18 21 25 28 29
c55 18 0 1.55237e-19 $X=10.777 $Y=1.22
r56 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.42
+ $Y=1.385 $X2=11.42 $Y2=1.385
r57 23 29 0.674692 $w=3.3e-07 $l=9.8e-08 $layer=LI1_cond $X=10.875 $Y=1.385
+ $X2=10.777 $Y2=1.385
r58 23 25 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=10.875 $Y=1.385
+ $X2=11.42 $Y2=1.385
r59 19 29 8.18839 $w=1.82e-07 $l=1.70895e-07 $layer=LI1_cond $X=10.765 $Y=1.55
+ $X2=10.777 $Y2=1.385
r60 19 21 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=10.765 $Y=1.55
+ $X2=10.765 $Y2=2.16
r61 18 29 8.18839 $w=1.82e-07 $l=1.65e-07 $layer=LI1_cond $X=10.777 $Y=1.22
+ $X2=10.777 $Y2=1.385
r62 18 28 15.9254 $w=1.93e-07 $l=2.8e-07 $layer=LI1_cond $X=10.777 $Y=1.22
+ $X2=10.777 $Y2=0.94
r63 13 28 7.67512 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=10.71 $Y=0.775
+ $X2=10.71 $Y2=0.94
r64 13 15 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=10.71 $Y=0.775
+ $X2=10.71 $Y2=0.645
r65 10 26 38.9026 $w=2.7e-07 $l=2.03101e-07 $layer=POLY_cond $X=11.505 $Y=1.22
+ $X2=11.42 $Y2=1.385
r66 10 12 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=11.505 $Y=1.22
+ $X2=11.505 $Y2=0.74
r67 7 26 77.2841 $w=2.7e-07 $l=4.15812e-07 $layer=POLY_cond $X=11.495 $Y=1.765
+ $X2=11.42 $Y2=1.385
r68 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=11.495 $Y=1.765
+ $X2=11.495 $Y2=2.4
r69 2 21 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=10.62
+ $Y=2.015 $X2=10.765 $Y2=2.16
r70 1 15 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=10.565
+ $Y=0.37 $X2=10.71 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_LS__DFSBP_1%A_27_80# 1 2 3 4 15 18 21 23 25 28 29 30 31
+ 36
c68 25 0 1.22627e-19 $X=2.525 $Y=2.145
r69 36 38 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.69 $Y=0.68
+ $X2=2.69 $Y2=0.845
r70 31 33 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=1.71 $Y=2.145
+ $X2=1.71 $Y2=2.275
r71 28 38 79.2674 $w=1.68e-07 $l=1.215e-06 $layer=LI1_cond $X=2.61 $Y=2.06
+ $X2=2.61 $Y2=0.845
r72 26 31 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.795 $Y=2.145
+ $X2=1.71 $Y2=2.145
r73 25 41 12.1344 $w=3.72e-07 $l=4.75079e-07 $layer=LI1_cond $X=2.525 $Y=2.145
+ $X2=2.765 $Y2=2.515
r74 25 28 6.42219 $w=3.72e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.525 $Y=2.145
+ $X2=2.61 $Y2=2.06
r75 25 26 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=2.525 $Y=2.145
+ $X2=1.795 $Y2=2.145
r76 24 30 2.11342 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.365 $Y=2.275
+ $X2=0.24 $Y2=2.275
r77 23 33 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.625 $Y=2.275
+ $X2=1.71 $Y2=2.275
r78 23 24 82.2032 $w=1.68e-07 $l=1.26e-06 $layer=LI1_cond $X=1.625 $Y=2.275
+ $X2=0.365 $Y2=2.275
r79 19 30 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.24 $Y=2.36 $X2=0.24
+ $Y2=2.275
r80 19 21 17.9781 $w=2.48e-07 $l=3.9e-07 $layer=LI1_cond $X=0.24 $Y=2.36
+ $X2=0.24 $Y2=2.75
r81 18 30 4.3182 $w=2.1e-07 $l=1.03078e-07 $layer=LI1_cond $X=0.2 $Y=2.19
+ $X2=0.24 $Y2=2.275
r82 18 29 88.0749 $w=1.68e-07 $l=1.35e-06 $layer=LI1_cond $X=0.2 $Y=2.19 $X2=0.2
+ $Y2=0.84
r83 13 29 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=0.24 $Y=0.715
+ $X2=0.24 $Y2=0.84
r84 13 15 4.84026 $w=2.48e-07 $l=1.05e-07 $layer=LI1_cond $X=0.24 $Y=0.715
+ $X2=0.24 $Y2=0.61
r85 4 41 600 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=1 $X=2.695
+ $Y=2.315 $X2=2.84 $Y2=2.515
r86 3 21 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.54 $X2=0.28 $Y2=2.75
r87 2 36 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=2.545
+ $Y=0.405 $X2=2.69 $Y2=0.68
r88 1 15 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.4 $X2=0.28 $Y2=0.61
.ends

.subckt PM_SKY130_FD_SC_LS__DFSBP_1%VPWR 1 2 3 4 5 6 7 24 28 32 36 40 44 48 51
+ 52 53 55 60 65 70 82 89 96 97 100 103 106 109 112 115
c141 28 0 2.99812e-20 $X=1.74 $Y=2.695
c142 4 0 1.03271e-19 $X=5.475 $Y=2.315
r143 115 116 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r144 112 113 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r145 106 107 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r146 103 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r147 100 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r148 97 116 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=11.28 $Y2=3.33
r149 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r150 94 115 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.38 $Y=3.33
+ $X2=11.215 $Y2=3.33
r151 94 96 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=11.38 $Y=3.33
+ $X2=11.76 $Y2=3.33
r152 93 116 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=11.28 $Y2=3.33
r153 93 113 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=9.84 $Y2=3.33
r154 92 93 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r155 90 112 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=9.91 $Y=3.33
+ $X2=9.735 $Y2=3.33
r156 90 92 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=9.91 $Y=3.33
+ $X2=10.8 $Y2=3.33
r157 89 115 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.05 $Y=3.33
+ $X2=11.215 $Y2=3.33
r158 89 92 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=11.05 $Y=3.33
+ $X2=10.8 $Y2=3.33
r159 88 113 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=9.84 $Y2=3.33
r160 87 88 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r161 85 88 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=9.36 $Y2=3.33
r162 84 87 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=8.4 $Y=3.33 $X2=9.36
+ $Y2=3.33
r163 84 85 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r164 82 112 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=9.56 $Y=3.33
+ $X2=9.735 $Y2=3.33
r165 82 87 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=9.56 $Y=3.33 $X2=9.36
+ $Y2=3.33
r166 81 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r167 80 81 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r168 78 109 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=6.05 $Y=3.33
+ $X2=5.88 $Y2=3.33
r169 78 80 122 $w=1.68e-07 $l=1.87e-06 $layer=LI1_cond $X=6.05 $Y=3.33 $X2=7.92
+ $Y2=3.33
r170 76 77 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r171 74 77 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r172 74 107 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r173 73 76 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r174 73 74 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r175 71 106 9.73034 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=4.44 $Y=3.33
+ $X2=4.242 $Y2=3.33
r176 71 73 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=4.44 $Y=3.33
+ $X2=4.56 $Y2=3.33
r177 70 109 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=5.71 $Y=3.33
+ $X2=5.88 $Y2=3.33
r178 70 76 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=5.71 $Y=3.33
+ $X2=5.52 $Y2=3.33
r179 69 107 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=4.08 $Y2=3.33
r180 69 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r181 68 69 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r182 66 103 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.905 $Y=3.33
+ $X2=1.74 $Y2=3.33
r183 66 68 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.905 $Y=3.33
+ $X2=2.16 $Y2=3.33
r184 65 106 9.73034 $w=1.7e-07 $l=1.97e-07 $layer=LI1_cond $X=4.045 $Y=3.33
+ $X2=4.242 $Y2=3.33
r185 65 68 122.979 $w=1.68e-07 $l=1.885e-06 $layer=LI1_cond $X=4.045 $Y=3.33
+ $X2=2.16 $Y2=3.33
r186 64 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r187 64 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r188 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r189 61 100 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=0.73 $Y2=3.33
r190 61 63 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=1.2 $Y2=3.33
r191 60 103 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.575 $Y=3.33
+ $X2=1.74 $Y2=3.33
r192 60 63 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.575 $Y=3.33
+ $X2=1.2 $Y2=3.33
r193 58 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r194 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r195 55 100 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.73 $Y2=3.33
r196 55 57 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.24 $Y2=3.33
r197 53 81 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=7.92 $Y2=3.33
r198 53 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=5.52
+ $Y2=3.33
r199 53 109 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r200 51 80 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=8.07 $Y=3.33
+ $X2=7.92 $Y2=3.33
r201 51 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.07 $Y=3.33
+ $X2=8.155 $Y2=3.33
r202 50 84 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=8.24 $Y=3.33
+ $X2=8.4 $Y2=3.33
r203 50 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.24 $Y=3.33
+ $X2=8.155 $Y2=3.33
r204 46 115 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.215 $Y=3.245
+ $X2=11.215 $Y2=3.33
r205 46 48 37.8909 $w=3.28e-07 $l=1.085e-06 $layer=LI1_cond $X=11.215 $Y=3.245
+ $X2=11.215 $Y2=2.16
r206 42 112 1.07557 $w=3.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.735 $Y=3.245
+ $X2=9.735 $Y2=3.33
r207 42 44 14.1586 $w=3.48e-07 $l=4.3e-07 $layer=LI1_cond $X=9.735 $Y=3.245
+ $X2=9.735 $Y2=2.815
r208 38 52 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.155 $Y=3.245
+ $X2=8.155 $Y2=3.33
r209 38 40 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=8.155 $Y=3.245
+ $X2=8.155 $Y2=2.815
r210 34 109 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=5.88 $Y=3.245
+ $X2=5.88 $Y2=3.33
r211 34 36 20.8457 $w=3.38e-07 $l=6.15e-07 $layer=LI1_cond $X=5.88 $Y=3.245
+ $X2=5.88 $Y2=2.63
r212 30 106 1.43204 $w=3.95e-07 $l=8.5e-08 $layer=LI1_cond $X=4.242 $Y=3.245
+ $X2=4.242 $Y2=3.33
r213 30 32 19.1101 $w=3.93e-07 $l=6.55e-07 $layer=LI1_cond $X=4.242 $Y=3.245
+ $X2=4.242 $Y2=2.59
r214 26 103 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.74 $Y=3.245
+ $X2=1.74 $Y2=3.33
r215 26 28 19.2074 $w=3.28e-07 $l=5.5e-07 $layer=LI1_cond $X=1.74 $Y=3.245
+ $X2=1.74 $Y2=2.695
r216 22 100 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=3.33
r217 22 24 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=2.755
r218 7 48 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=11.065
+ $Y=2.015 $X2=11.215 $Y2=2.16
r219 6 44 600 $w=1.7e-07 $l=3.55668e-07 $layer=licon1_PDIFF $count=1 $X=9.55
+ $Y=2.54 $X2=9.735 $Y2=2.815
r220 5 40 600 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=8.005
+ $Y=2.54 $X2=8.155 $Y2=2.815
r221 4 36 600 $w=1.7e-07 $l=4.98197e-07 $layer=licon1_PDIFF $count=1 $X=5.475
+ $Y=2.315 $X2=5.84 $Y2=2.63
r222 3 32 600 $w=1.7e-07 $l=3.5373e-07 $layer=licon1_PDIFF $count=1 $X=4.06
+ $Y=2.315 $X2=4.24 $Y2=2.59
r223 2 28 600 $w=1.7e-07 $l=9.77126e-07 $layer=licon1_PDIFF $count=1 $X=1.59
+ $Y=1.79 $X2=1.74 $Y2=2.695
r224 1 24 600 $w=1.7e-07 $l=2.80134e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=2.54 $X2=0.73 $Y2=2.755
.ends

.subckt PM_SKY130_FD_SC_LS__DFSBP_1%Q_N 1 2 9 11 12 13 14 15 22 39
r31 22 39 1.62667 $w=3.15e-07 $l=8.54576e-08 $layer=LI1_cond $X=10.277 $Y=1.337
+ $X2=10.21 $Y2=1.295
r32 15 35 1.46342 $w=3.13e-07 $l=4e-08 $layer=LI1_cond $X=10.277 $Y=2.775
+ $X2=10.277 $Y2=2.815
r33 14 15 13.5366 $w=3.13e-07 $l=3.7e-07 $layer=LI1_cond $X=10.277 $Y=2.405
+ $X2=10.277 $Y2=2.775
r34 13 14 13.5366 $w=3.13e-07 $l=3.7e-07 $layer=LI1_cond $X=10.277 $Y=2.035
+ $X2=10.277 $Y2=2.405
r35 13 27 1.82927 $w=3.13e-07 $l=5e-08 $layer=LI1_cond $X=10.277 $Y=2.035
+ $X2=10.277 $Y2=1.985
r36 12 27 11.7074 $w=3.13e-07 $l=3.2e-07 $layer=LI1_cond $X=10.277 $Y=1.665
+ $X2=10.277 $Y2=1.985
r37 11 39 0.88 $w=3.05e-07 $l=2.2e-08 $layer=LI1_cond $X=10.21 $Y=1.273
+ $X2=10.21 $Y2=1.295
r38 11 12 11.2317 $w=3.13e-07 $l=3.07e-07 $layer=LI1_cond $X=10.277 $Y=1.358
+ $X2=10.277 $Y2=1.665
r39 11 22 0.768295 $w=3.13e-07 $l=2.1e-08 $layer=LI1_cond $X=10.277 $Y=1.358
+ $X2=10.277 $Y2=1.337
r40 7 11 11.4767 $w=3.3e-07 $l=3.36666e-07 $layer=LI1_cond $X=10.15 $Y=0.965
+ $X2=10.21 $Y2=1.273
r41 7 9 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=10.15 $Y=0.965
+ $X2=10.15 $Y2=0.515
r42 2 35 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=10.055
+ $Y=1.84 $X2=10.205 $Y2=2.815
r43 2 27 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=10.055
+ $Y=1.84 $X2=10.205 $Y2=1.985
r44 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.01
+ $Y=0.37 $X2=10.15 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__DFSBP_1%Q 1 2 9 13 14 15 16 24 33
r20 15 16 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=11.72 $Y=2.405
+ $X2=11.72 $Y2=2.775
r21 14 24 0.628605 $w=3.28e-07 $l=1.8e-08 $layer=LI1_cond $X=11.72 $Y=1.967
+ $X2=11.72 $Y2=1.985
r22 14 33 7.83357 $w=3.28e-07 $l=1.47e-07 $layer=LI1_cond $X=11.72 $Y=1.967
+ $X2=11.72 $Y2=1.82
r23 14 15 12.3276 $w=3.28e-07 $l=3.53e-07 $layer=LI1_cond $X=11.72 $Y=2.052
+ $X2=11.72 $Y2=2.405
r24 14 24 2.33981 $w=3.28e-07 $l=6.7e-08 $layer=LI1_cond $X=11.72 $Y=2.052
+ $X2=11.72 $Y2=1.985
r25 13 33 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=11.8 $Y=1.05
+ $X2=11.8 $Y2=1.82
r26 7 13 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=11.72 $Y=0.885
+ $X2=11.72 $Y2=1.05
r27 7 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=11.72 $Y=0.885
+ $X2=11.72 $Y2=0.515
r28 2 16 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=11.57
+ $Y=1.84 $X2=11.72 $Y2=2.815
r29 2 24 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=11.57
+ $Y=1.84 $X2=11.72 $Y2=1.985
r30 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=11.58
+ $Y=0.37 $X2=11.72 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__DFSBP_1%VGND 1 2 3 4 5 6 7 24 26 30 34 38 42 46 49
+ 50 52 53 54 56 68 75 87 96 97 100 103 106 110 116
c130 38 0 2.3488e-20 $X=6.02 $Y=0.495
c131 30 0 1.39813e-19 $X=1.7 $Y=0.505
r132 116 117 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r133 110 113 9.62063 $w=6.88e-07 $l=5.55e-07 $layer=LI1_cond $X=8.41 $Y=0
+ $X2=8.41 $Y2=0.555
r134 110 111 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r135 103 104 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0
+ $X2=1.68 $Y2=0
r136 101 104 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0
+ $X2=1.68 $Y2=0
r137 100 101 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0
+ $X2=0.72 $Y2=0
r138 97 117 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=11.28 $Y2=0
r139 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r140 94 116 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.385 $Y=0
+ $X2=11.22 $Y2=0
r141 94 96 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=11.385 $Y=0
+ $X2=11.76 $Y2=0
r142 93 117 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=11.28 $Y2=0
r143 92 93 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.8 $Y=0 $X2=10.8
+ $Y2=0
r144 90 93 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.84 $Y=0 $X2=10.8
+ $Y2=0
r145 89 92 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=9.84 $Y=0 $X2=10.8
+ $Y2=0
r146 89 90 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r147 87 116 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.055 $Y=0
+ $X2=11.22 $Y2=0
r148 87 92 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=11.055 $Y=0
+ $X2=10.8 $Y2=0
r149 86 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0 $X2=9.84
+ $Y2=0
r150 86 111 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.36 $Y=0 $X2=8.4
+ $Y2=0
r151 85 86 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r152 83 110 9.22683 $w=1.7e-07 $l=3.45e-07 $layer=LI1_cond $X=8.755 $Y=0
+ $X2=8.41 $Y2=0
r153 83 85 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=8.755 $Y=0
+ $X2=9.36 $Y2=0
r154 82 111 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.4
+ $Y2=0
r155 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r156 79 82 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=6.48 $Y=0
+ $X2=7.92 $Y2=0
r157 78 81 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=6.48 $Y=0 $X2=7.92
+ $Y2=0
r158 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r159 76 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.185 $Y=0
+ $X2=6.02 $Y2=0
r160 76 78 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=6.185 $Y=0 $X2=6.48
+ $Y2=0
r161 75 110 9.22683 $w=1.7e-07 $l=3.45e-07 $layer=LI1_cond $X=8.065 $Y=0
+ $X2=8.41 $Y2=0
r162 75 81 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=8.065 $Y=0
+ $X2=7.92 $Y2=0
r163 73 74 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r164 71 74 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.52
+ $Y2=0
r165 70 73 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.56 $Y=0 $X2=5.52
+ $Y2=0
r166 70 71 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r167 68 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.855 $Y=0
+ $X2=6.02 $Y2=0
r168 68 73 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=5.855 $Y=0
+ $X2=5.52 $Y2=0
r169 67 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r170 66 67 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r171 64 67 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=4.08 $Y2=0
r172 64 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=1.68 $Y2=0
r173 63 66 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=2.16 $Y=0 $X2=4.08
+ $Y2=0
r174 63 64 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r175 61 103 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.865 $Y=0
+ $X2=1.735 $Y2=0
r176 61 63 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.865 $Y=0 $X2=2.16
+ $Y2=0
r177 59 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0
+ $X2=0.72 $Y2=0
r178 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r179 56 100 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.545 $Y=0
+ $X2=0.67 $Y2=0
r180 56 58 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0
+ $X2=0.24 $Y2=0
r181 54 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r182 54 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.52
+ $Y2=0
r183 54 106 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r184 52 85 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=9.485 $Y=0
+ $X2=9.36 $Y2=0
r185 52 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.485 $Y=0 $X2=9.65
+ $Y2=0
r186 51 89 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=9.815 $Y=0 $X2=9.84
+ $Y2=0
r187 51 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.815 $Y=0 $X2=9.65
+ $Y2=0
r188 49 66 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=4.105 $Y=0 $X2=4.08
+ $Y2=0
r189 49 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.105 $Y=0 $X2=4.27
+ $Y2=0
r190 48 70 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=4.435 $Y=0
+ $X2=4.56 $Y2=0
r191 48 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.435 $Y=0 $X2=4.27
+ $Y2=0
r192 44 116 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.22 $Y=0.085
+ $X2=11.22 $Y2=0
r193 44 46 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=11.22 $Y=0.085
+ $X2=11.22 $Y2=0.495
r194 40 53 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.65 $Y=0.085
+ $X2=9.65 $Y2=0
r195 40 42 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=9.65 $Y=0.085
+ $X2=9.65 $Y2=0.55
r196 36 106 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.02 $Y=0.085
+ $X2=6.02 $Y2=0
r197 36 38 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=6.02 $Y=0.085
+ $X2=6.02 $Y2=0.495
r198 32 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.27 $Y=0.085
+ $X2=4.27 $Y2=0
r199 32 34 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=4.27 $Y=0.085
+ $X2=4.27 $Y2=0.55
r200 28 103 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.735 $Y=0.085
+ $X2=1.735 $Y2=0
r201 28 30 18.6164 $w=2.58e-07 $l=4.2e-07 $layer=LI1_cond $X=1.735 $Y=0.085
+ $X2=1.735 $Y2=0.505
r202 27 100 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.795 $Y=0
+ $X2=0.67 $Y2=0
r203 26 103 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.605 $Y=0
+ $X2=1.735 $Y2=0
r204 26 27 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=1.605 $Y=0
+ $X2=0.795 $Y2=0
r205 22 100 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.67 $Y=0.085
+ $X2=0.67 $Y2=0
r206 22 24 24.2013 $w=2.48e-07 $l=5.25e-07 $layer=LI1_cond $X=0.67 $Y=0.085
+ $X2=0.67 $Y2=0.61
r207 7 46 91 $w=1.7e-07 $l=2.755e-07 $layer=licon1_NDIFF $count=2 $X=11 $Y=0.37
+ $X2=11.22 $Y2=0.495
r208 6 42 182 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_NDIFF $count=1 $X=9.505
+ $Y=0.37 $X2=9.65 $Y2=0.55
r209 5 113 91 $w=1.7e-07 $l=5.85235e-07 $layer=licon1_NDIFF $count=2 $X=8.09
+ $Y=0.37 $X2=8.59 $Y2=0.555
r210 4 38 91 $w=1.7e-07 $l=3.82426e-07 $layer=licon1_NDIFF $count=2 $X=5.695
+ $Y=0.37 $X2=6.02 $Y2=0.495
r211 3 34 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=4.13
+ $Y=0.405 $X2=4.27 $Y2=0.55
r212 2 30 91 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=2 $X=1.56
+ $Y=0.37 $X2=1.7 $Y2=0.505
r213 1 24 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.4 $X2=0.71 $Y2=0.61
.ends

