* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
X0 a_504_392# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 VPWR a_187_244# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X2 VGND a_187_244# X VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X3 a_187_244# A1 a_587_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X4 a_32_368# B1_N VGND VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X5 VPWR A2 a_504_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 X a_187_244# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X7 X a_187_244# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X8 a_32_368# B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X9 a_187_244# a_32_368# a_504_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_587_74# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X11 VGND a_32_368# a_187_244# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
.ends
