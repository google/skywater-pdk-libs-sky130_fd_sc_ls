* File: sky130_fd_sc_ls__nor3b_4.pex.spice
* Created: Wed Sep  2 11:15:16 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__NOR3B_4%B 3 5 7 10 12 14 15 17 20 22 24 27 29 30 31
+ 32 49
c82 15 0 1.9472e-19 $X=1.455 $Y=1.765
c83 10 0 9.05221e-20 $X=0.995 $Y=0.74
r84 49 50 1.96467 $w=3.68e-07 $l=1.5e-08 $layer=POLY_cond $X=1.98 $Y=1.557
+ $X2=1.995 $Y2=1.557
r85 47 49 43.2228 $w=3.68e-07 $l=3.3e-07 $layer=POLY_cond $X=1.65 $Y=1.557
+ $X2=1.98 $Y2=1.557
r86 47 48 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.65
+ $Y=1.515 $X2=1.65 $Y2=1.515
r87 45 47 11.1332 $w=3.68e-07 $l=8.5e-08 $layer=POLY_cond $X=1.565 $Y=1.557
+ $X2=1.65 $Y2=1.557
r88 44 45 14.4076 $w=3.68e-07 $l=1.1e-07 $layer=POLY_cond $X=1.455 $Y=1.557
+ $X2=1.565 $Y2=1.557
r89 43 44 58.9402 $w=3.68e-07 $l=4.5e-07 $layer=POLY_cond $X=1.005 $Y=1.557
+ $X2=1.455 $Y2=1.557
r90 42 43 1.30978 $w=3.68e-07 $l=1e-08 $layer=POLY_cond $X=0.995 $Y=1.557
+ $X2=1.005 $Y2=1.557
r91 40 42 47.8071 $w=3.68e-07 $l=3.65e-07 $layer=POLY_cond $X=0.63 $Y=1.557
+ $X2=0.995 $Y2=1.557
r92 40 41 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.63
+ $Y=1.515 $X2=0.63 $Y2=1.515
r93 38 40 9.82337 $w=3.68e-07 $l=7.5e-08 $layer=POLY_cond $X=0.555 $Y=1.557
+ $X2=0.63 $Y2=1.557
r94 37 38 1.96467 $w=3.68e-07 $l=1.5e-08 $layer=POLY_cond $X=0.54 $Y=1.557
+ $X2=0.555 $Y2=1.557
r95 32 48 0.80403 $w=4.28e-07 $l=3e-08 $layer=LI1_cond $X=1.68 $Y=1.565 $X2=1.65
+ $Y2=1.565
r96 31 48 12.0604 $w=4.28e-07 $l=4.5e-07 $layer=LI1_cond $X=1.2 $Y=1.565
+ $X2=1.65 $Y2=1.565
r97 30 31 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=1.2 $Y2=1.565
r98 30 41 2.41209 $w=4.28e-07 $l=9e-08 $layer=LI1_cond $X=0.72 $Y=1.565 $X2=0.63
+ $Y2=1.565
r99 29 41 10.4524 $w=4.28e-07 $l=3.9e-07 $layer=LI1_cond $X=0.24 $Y=1.565
+ $X2=0.63 $Y2=1.565
r100 25 50 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.995 $Y=1.35
+ $X2=1.995 $Y2=1.557
r101 25 27 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.995 $Y=1.35
+ $X2=1.995 $Y2=0.74
r102 22 49 23.8357 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.98 $Y=1.765
+ $X2=1.98 $Y2=1.557
r103 22 24 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.98 $Y=1.765
+ $X2=1.98 $Y2=2.4
r104 18 45 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.565 $Y=1.35
+ $X2=1.565 $Y2=1.557
r105 18 20 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.565 $Y=1.35
+ $X2=1.565 $Y2=0.74
r106 15 44 23.8357 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.455 $Y=1.765
+ $X2=1.455 $Y2=1.557
r107 15 17 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.455 $Y=1.765
+ $X2=1.455 $Y2=2.4
r108 12 43 23.8357 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.005 $Y=1.765
+ $X2=1.005 $Y2=1.557
r109 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.005 $Y=1.765
+ $X2=1.005 $Y2=2.4
r110 8 42 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.995 $Y=1.35
+ $X2=0.995 $Y2=1.557
r111 8 10 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.995 $Y=1.35
+ $X2=0.995 $Y2=0.74
r112 5 38 23.8357 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.555 $Y=1.765
+ $X2=0.555 $Y2=1.557
r113 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.555 $Y=1.765
+ $X2=0.555 $Y2=2.4
r114 1 37 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.54 $Y=1.35
+ $X2=0.54 $Y2=1.557
r115 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.54 $Y=1.35 $X2=0.54
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__NOR3B_4%A_468_264# 1 2 7 9 12 14 16 19 21 23 26 28
+ 30 33 35 43 49 51 53 54 59 61 70
c149 70 0 2.89644e-19 $X=3.78 $Y=1.542
c150 61 0 1.69815e-19 $X=7.4 $Y=0.5
c151 7 0 8.42778e-20 $X=2.43 $Y=1.765
r152 70 71 9.46335 $w=3.82e-07 $l=7.5e-08 $layer=POLY_cond $X=3.78 $Y=1.542
+ $X2=3.855 $Y2=1.542
r153 67 68 11.9869 $w=3.82e-07 $l=9.5e-08 $layer=POLY_cond $X=3.33 $Y=1.542
+ $X2=3.425 $Y2=1.542
r154 66 67 51.1021 $w=3.82e-07 $l=4.05e-07 $layer=POLY_cond $X=2.925 $Y=1.542
+ $X2=3.33 $Y2=1.542
r155 65 66 5.67801 $w=3.82e-07 $l=4.5e-08 $layer=POLY_cond $X=2.88 $Y=1.542
+ $X2=2.925 $Y2=1.542
r156 62 63 8.20157 $w=3.82e-07 $l=6.5e-08 $layer=POLY_cond $X=2.43 $Y=1.542
+ $X2=2.495 $Y2=1.542
r157 53 61 8.35471 $w=1.7e-07 $l=3.3e-07 $layer=LI1_cond $X=7.48 $Y=1.01
+ $X2=7.48 $Y2=0.68
r158 53 54 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=7.48 $Y=1.01
+ $X2=7.48 $Y2=1.72
r159 52 59 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=7.055 $Y=1.805
+ $X2=6.92 $Y2=1.805
r160 51 54 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.395 $Y=1.805
+ $X2=7.48 $Y2=1.72
r161 51 52 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=7.395 $Y=1.805
+ $X2=7.055 $Y2=1.805
r162 47 59 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.92 $Y=1.89
+ $X2=6.92 $Y2=1.805
r163 47 49 4.05489 $w=2.68e-07 $l=9.5e-08 $layer=LI1_cond $X=6.92 $Y=1.89
+ $X2=6.92 $Y2=1.985
r164 44 57 4.15824 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=4.195 $Y=1.805
+ $X2=4.042 $Y2=1.805
r165 43 59 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=6.785 $Y=1.805
+ $X2=6.92 $Y2=1.805
r166 43 44 168.973 $w=1.68e-07 $l=2.59e-06 $layer=LI1_cond $X=6.785 $Y=1.805
+ $X2=4.195 $Y2=1.805
r167 42 70 1.89267 $w=3.82e-07 $l=1.5e-08 $layer=POLY_cond $X=3.765 $Y=1.542
+ $X2=3.78 $Y2=1.542
r168 42 68 42.9005 $w=3.82e-07 $l=3.4e-07 $layer=POLY_cond $X=3.765 $Y=1.542
+ $X2=3.425 $Y2=1.542
r169 41 42 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.765
+ $Y=1.485 $X2=3.765 $Y2=1.485
r170 38 65 17.034 $w=3.82e-07 $l=1.35e-07 $layer=POLY_cond $X=2.745 $Y=1.542
+ $X2=2.88 $Y2=1.542
r171 38 63 31.5445 $w=3.82e-07 $l=2.5e-07 $layer=POLY_cond $X=2.745 $Y=1.542
+ $X2=2.495 $Y2=1.542
r172 37 41 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=2.745 $Y=1.485
+ $X2=3.765 $Y2=1.485
r173 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.745
+ $Y=1.485 $X2=2.745 $Y2=1.485
r174 35 57 12.0912 $w=3.03e-07 $l=3.2e-07 $layer=LI1_cond $X=4.042 $Y=1.485
+ $X2=4.042 $Y2=1.805
r175 35 41 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=3.89 $Y=1.485
+ $X2=3.765 $Y2=1.485
r176 31 71 24.74 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=3.855 $Y=1.32
+ $X2=3.855 $Y2=1.542
r177 31 33 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.855 $Y=1.32
+ $X2=3.855 $Y2=0.74
r178 28 70 24.74 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=3.78 $Y=1.765
+ $X2=3.78 $Y2=1.542
r179 28 30 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.78 $Y=1.765
+ $X2=3.78 $Y2=2.4
r180 24 68 24.74 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=3.425 $Y=1.32
+ $X2=3.425 $Y2=1.542
r181 24 26 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.425 $Y=1.32
+ $X2=3.425 $Y2=0.74
r182 21 67 24.74 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=3.33 $Y=1.765
+ $X2=3.33 $Y2=1.542
r183 21 23 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.33 $Y=1.765
+ $X2=3.33 $Y2=2.4
r184 17 66 24.74 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=2.925 $Y=1.32
+ $X2=2.925 $Y2=1.542
r185 17 19 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.925 $Y=1.32
+ $X2=2.925 $Y2=0.74
r186 14 65 24.74 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=2.88 $Y=1.765
+ $X2=2.88 $Y2=1.542
r187 14 16 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.88 $Y=1.765
+ $X2=2.88 $Y2=2.4
r188 10 63 24.74 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=2.495 $Y=1.32
+ $X2=2.495 $Y2=1.542
r189 10 12 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.495 $Y=1.32
+ $X2=2.495 $Y2=0.74
r190 7 62 24.74 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=2.43 $Y=1.765
+ $X2=2.43 $Y2=1.542
r191 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.43 $Y=1.765
+ $X2=2.43 $Y2=2.4
r192 2 49 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=6.8
+ $Y=1.84 $X2=6.95 $Y2=1.985
r193 1 61 45.5 $w=1.7e-07 $l=8.32466e-07 $layer=licon1_NDIFF $count=4 $X=6.63
+ $Y=0.37 $X2=7.4 $Y2=0.5
.ends

.subckt PM_SKY130_FD_SC_LS__NOR3B_4%A 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22 24
+ 33 43 46
c89 46 0 1.78853e-19 $X=6.365 $Y=1.365
c90 43 0 1.83401e-19 $X=6.055 $Y=1.492
c91 19 0 1.69815e-19 $X=6.055 $Y=1.22
r92 43 44 10.1915 $w=4.02e-07 $l=8.5e-08 $layer=POLY_cond $X=6.055 $Y=1.492
+ $X2=6.14 $Y2=1.492
r93 40 41 16.1866 $w=4.02e-07 $l=1.35e-07 $layer=POLY_cond $X=5.555 $Y=1.492
+ $X2=5.69 $Y2=1.492
r94 39 40 37.7687 $w=4.02e-07 $l=3.15e-07 $layer=POLY_cond $X=5.24 $Y=1.492
+ $X2=5.555 $Y2=1.492
r95 38 39 46.1617 $w=4.02e-07 $l=3.85e-07 $layer=POLY_cond $X=4.855 $Y=1.492
+ $X2=5.24 $Y2=1.492
r96 37 38 7.79353 $w=4.02e-07 $l=6.5e-08 $layer=POLY_cond $X=4.79 $Y=1.492
+ $X2=4.855 $Y2=1.492
r97 33 46 3.7435 $w=3.68e-07 $l=1.15e-07 $layer=LI1_cond $X=6.48 $Y=1.365
+ $X2=6.365 $Y2=1.365
r98 32 43 10.791 $w=4.02e-07 $l=9e-08 $layer=POLY_cond $X=5.965 $Y=1.492
+ $X2=6.055 $Y2=1.492
r99 32 41 32.9726 $w=4.02e-07 $l=2.75e-07 $layer=POLY_cond $X=5.965 $Y=1.492
+ $X2=5.69 $Y2=1.492
r100 31 46 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=5.965 $Y=1.385
+ $X2=6.365 $Y2=1.385
r101 31 32 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=5.965
+ $Y=1.385 $X2=5.965 $Y2=1.385
r102 28 37 22.1816 $w=4.02e-07 $l=1.85e-07 $layer=POLY_cond $X=4.605 $Y=1.492
+ $X2=4.79 $Y2=1.492
r103 28 35 21.5821 $w=4.02e-07 $l=1.8e-07 $layer=POLY_cond $X=4.605 $Y=1.492
+ $X2=4.425 $Y2=1.492
r104 27 31 47.4946 $w=3.28e-07 $l=1.36e-06 $layer=LI1_cond $X=4.605 $Y=1.385
+ $X2=5.965 $Y2=1.385
r105 27 28 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=4.605
+ $Y=1.385 $X2=4.605 $Y2=1.385
r106 22 44 25.9839 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=6.14 $Y=1.765
+ $X2=6.14 $Y2=1.492
r107 22 24 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.14 $Y=1.765
+ $X2=6.14 $Y2=2.4
r108 19 43 25.9839 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=6.055 $Y=1.22
+ $X2=6.055 $Y2=1.492
r109 19 21 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=6.055 $Y=1.22
+ $X2=6.055 $Y2=0.74
r110 16 41 25.9839 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=5.69 $Y=1.765
+ $X2=5.69 $Y2=1.492
r111 16 18 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.69 $Y=1.765
+ $X2=5.69 $Y2=2.4
r112 13 40 25.9839 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=5.555 $Y=1.22
+ $X2=5.555 $Y2=1.492
r113 13 15 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.555 $Y=1.22
+ $X2=5.555 $Y2=0.74
r114 10 39 25.9839 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=5.24 $Y=1.765
+ $X2=5.24 $Y2=1.492
r115 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.24 $Y=1.765
+ $X2=5.24 $Y2=2.4
r116 7 38 25.9839 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=4.855 $Y=1.22
+ $X2=4.855 $Y2=1.492
r117 7 9 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.855 $Y=1.22
+ $X2=4.855 $Y2=0.74
r118 4 37 25.9839 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=4.79 $Y=1.765
+ $X2=4.79 $Y2=1.492
r119 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.79 $Y=1.765
+ $X2=4.79 $Y2=2.4
r120 1 35 25.9839 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=4.425 $Y=1.22
+ $X2=4.425 $Y2=1.492
r121 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.425 $Y=1.22
+ $X2=4.425 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__NOR3B_4%C_N 1 3 4 6 7 9 10 15
c38 10 0 1.83401e-19 $X=6.96 $Y=1.295
r39 15 17 26.2422 $w=4.5e-07 $l=2.45e-07 $layer=POLY_cond $X=6.93 $Y=1.492
+ $X2=7.175 $Y2=1.492
r40 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.93
+ $Y=1.385 $X2=6.93 $Y2=1.385
r41 13 15 21.9578 $w=4.5e-07 $l=2.05e-07 $layer=POLY_cond $X=6.725 $Y=1.492
+ $X2=6.93 $Y2=1.492
r42 10 16 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=6.93 $Y=1.295 $X2=6.93
+ $Y2=1.385
r43 7 17 28.7666 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=7.175 $Y=1.765
+ $X2=7.175 $Y2=1.492
r44 7 9 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=7.175 $Y=1.765
+ $X2=7.175 $Y2=2.26
r45 4 13 28.7666 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=6.725 $Y=1.765
+ $X2=6.725 $Y2=1.492
r46 4 6 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=6.725 $Y=1.765
+ $X2=6.725 $Y2=2.26
r47 1 13 18.2089 $w=4.5e-07 $l=3.46733e-07 $layer=POLY_cond $X=6.555 $Y=1.22
+ $X2=6.725 $Y2=1.492
r48 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=6.555 $Y=1.22 $X2=6.555
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__NOR3B_4%A_27_368# 1 2 3 4 5 18 22 23 26 28 32 34 35
+ 43 44 45
c66 28 0 8.42778e-20 $X=2.04 $Y=2.99
r67 45 48 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=4.005 $Y=2.665
+ $X2=4.005 $Y2=2.745
r68 42 44 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.105 $Y=2.745
+ $X2=3.27 $Y2=2.745
r69 42 43 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.105 $Y=2.745
+ $X2=2.94 $Y2=2.745
r70 38 39 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=2.205 $Y=2.745
+ $X2=2.205 $Y2=2.99
r71 35 38 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=2.205 $Y=2.665
+ $X2=2.205 $Y2=2.745
r72 32 45 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.84 $Y=2.665
+ $X2=4.005 $Y2=2.665
r73 32 44 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=3.84 $Y=2.665
+ $X2=3.27 $Y2=2.665
r74 31 35 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.37 $Y=2.665
+ $X2=2.205 $Y2=2.665
r75 31 43 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=2.37 $Y=2.665
+ $X2=2.94 $Y2=2.665
r76 29 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.315 $Y=2.99
+ $X2=1.23 $Y2=2.99
r77 28 39 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.04 $Y=2.99
+ $X2=2.205 $Y2=2.99
r78 28 29 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=2.04 $Y=2.99
+ $X2=1.315 $Y2=2.99
r79 24 34 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.23 $Y=2.905
+ $X2=1.23 $Y2=2.99
r80 24 26 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=1.23 $Y=2.905
+ $X2=1.23 $Y2=2.455
r81 22 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.145 $Y=2.99
+ $X2=1.23 $Y2=2.99
r82 22 23 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.145 $Y=2.99
+ $X2=0.445 $Y2=2.99
r83 18 21 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=0.28 $Y=2.115 $X2=0.28
+ $Y2=2.815
r84 16 23 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=2.905
+ $X2=0.445 $Y2=2.99
r85 16 21 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.28 $Y=2.905 $X2=0.28
+ $Y2=2.815
r86 5 48 600 $w=1.7e-07 $l=9.77126e-07 $layer=licon1_PDIFF $count=1 $X=3.855
+ $Y=1.84 $X2=4.005 $Y2=2.745
r87 4 42 600 $w=1.7e-07 $l=9.77126e-07 $layer=licon1_PDIFF $count=1 $X=2.955
+ $Y=1.84 $X2=3.105 $Y2=2.745
r88 3 38 600 $w=1.7e-07 $l=9.77126e-07 $layer=licon1_PDIFF $count=1 $X=2.055
+ $Y=1.84 $X2=2.205 $Y2=2.745
r89 2 26 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=1.08
+ $Y=1.84 $X2=1.23 $Y2=2.455
r90 1 21 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r91 1 18 400 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_LS__NOR3B_4%A_126_368# 1 2 3 4 15 17 21 23 25 27 30 32
+ 35
c68 17 0 1.10791e-19 $X=4.795 $Y=2.325
r69 32 33 10.4675 $w=3.38e-07 $l=2.9e-07 $layer=LI1_cond $X=1.697 $Y=2.035
+ $X2=1.697 $Y2=2.325
r70 25 40 2.81454 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.945 $Y=2.23
+ $X2=5.945 $Y2=2.145
r71 25 27 10.8842 $w=2.68e-07 $l=2.55e-07 $layer=LI1_cond $X=5.945 $Y=2.23
+ $X2=5.945 $Y2=2.485
r72 24 35 4.15824 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=5.1 $Y=2.145
+ $X2=4.947 $Y2=2.145
r73 23 40 4.47015 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.81 $Y=2.145
+ $X2=5.945 $Y2=2.145
r74 23 24 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=5.81 $Y=2.145
+ $X2=5.1 $Y2=2.145
r75 21 38 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=5.015 $Y=2.485
+ $X2=5.015 $Y2=2.41
r76 18 33 4.76605 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=1.87 $Y=2.325
+ $X2=1.697 $Y2=2.325
r77 17 38 5.45178 $w=3.03e-07 $l=8.5e-08 $layer=LI1_cond $X=4.947 $Y=2.325
+ $X2=4.947 $Y2=2.41
r78 17 35 6.8013 $w=3.03e-07 $l=1.8e-07 $layer=LI1_cond $X=4.947 $Y=2.325
+ $X2=4.947 $Y2=2.145
r79 17 18 190.829 $w=1.68e-07 $l=2.925e-06 $layer=LI1_cond $X=4.795 $Y=2.325
+ $X2=1.87 $Y2=2.325
r80 16 30 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=2.035
+ $X2=0.78 $Y2=2.035
r81 15 32 4.76605 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=1.525 $Y=2.035
+ $X2=1.697 $Y2=2.035
r82 15 16 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=1.525 $Y=2.035
+ $X2=0.945 $Y2=2.035
r83 4 40 600 $w=1.7e-07 $l=3.72525e-07 $layer=licon1_PDIFF $count=1 $X=5.765
+ $Y=1.84 $X2=5.915 $Y2=2.145
r84 4 27 300 $w=1.7e-07 $l=7.16083e-07 $layer=licon1_PDIFF $count=2 $X=5.765
+ $Y=1.84 $X2=5.915 $Y2=2.485
r85 3 35 600 $w=1.7e-07 $l=3.72525e-07 $layer=licon1_PDIFF $count=1 $X=4.865
+ $Y=1.84 $X2=5.015 $Y2=2.145
r86 3 21 300 $w=1.7e-07 $l=7.16083e-07 $layer=licon1_PDIFF $count=2 $X=4.865
+ $Y=1.84 $X2=5.015 $Y2=2.485
r87 2 32 300 $w=1.7e-07 $l=2.63106e-07 $layer=licon1_PDIFF $count=2 $X=1.53
+ $Y=1.84 $X2=1.69 $Y2=2.035
r88 1 30 300 $w=1.7e-07 $l=3.00791e-07 $layer=licon1_PDIFF $count=2 $X=0.63
+ $Y=1.84 $X2=0.78 $Y2=2.075
.ends

.subckt PM_SKY130_FD_SC_LS__NOR3B_4%Y 1 2 3 4 5 6 7 8 27 30 33 35 37 41 45 47 51
+ 53 57 59 63 66 69 71 72 73 74
c138 74 0 1.9472e-19 $X=2.16 $Y=1.665
c139 69 0 9.05221e-20 $X=2.275 $Y=1.08
r140 70 74 7.76646 $w=2.28e-07 $l=1.55e-07 $layer=LI1_cond $X=2.16 $Y=1.82
+ $X2=2.16 $Y2=1.665
r141 68 74 24.3015 $w=2.28e-07 $l=4.85e-07 $layer=LI1_cond $X=2.16 $Y=1.18
+ $X2=2.16 $Y2=1.665
r142 68 69 6.65862 $w=1.98e-07 $l=1.15e-07 $layer=LI1_cond $X=2.16 $Y=1.08
+ $X2=2.275 $Y2=1.08
r143 61 63 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=5.77 $Y=0.88
+ $X2=5.77 $Y2=0.515
r144 60 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.805 $Y=0.965
+ $X2=4.64 $Y2=0.965
r145 59 61 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.605 $Y=0.965
+ $X2=5.77 $Y2=0.88
r146 59 60 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=5.605 $Y=0.965
+ $X2=4.805 $Y2=0.965
r147 55 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.64 $Y=0.88
+ $X2=4.64 $Y2=0.965
r148 55 57 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=4.64 $Y=0.88
+ $X2=4.64 $Y2=0.515
r149 54 72 8.61065 $w=1.7e-07 $l=1.88348e-07 $layer=LI1_cond $X=3.805 $Y=0.965
+ $X2=3.64 $Y2=1.015
r150 53 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.475 $Y=0.965
+ $X2=4.64 $Y2=0.965
r151 53 54 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.475 $Y=0.965
+ $X2=3.805 $Y2=0.965
r152 49 72 0.89609 $w=3.3e-07 $l=1.35e-07 $layer=LI1_cond $X=3.64 $Y=0.88
+ $X2=3.64 $Y2=1.015
r153 49 51 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=3.64 $Y=0.88
+ $X2=3.64 $Y2=0.515
r154 48 71 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.795 $Y=1.065
+ $X2=2.71 $Y2=1.065
r155 47 72 8.61065 $w=1.7e-07 $l=1.88348e-07 $layer=LI1_cond $X=3.475 $Y=1.065
+ $X2=3.64 $Y2=1.015
r156 47 48 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.475 $Y=1.065
+ $X2=2.795 $Y2=1.065
r157 43 71 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.71 $Y=0.98
+ $X2=2.71 $Y2=1.065
r158 43 45 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=2.71 $Y=0.98
+ $X2=2.71 $Y2=0.515
r159 39 41 41.4879 $w=2.48e-07 $l=9e-07 $layer=LI1_cond $X=2.655 $Y=1.945
+ $X2=3.555 $Y2=1.945
r160 37 70 6.8319 $w=2.5e-07 $l=1.73205e-07 $layer=LI1_cond $X=2.275 $Y=1.945
+ $X2=2.16 $Y2=1.82
r161 37 39 17.5171 $w=2.48e-07 $l=3.8e-07 $layer=LI1_cond $X=2.275 $Y=1.945
+ $X2=2.655 $Y2=1.945
r162 35 71 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.625 $Y=1.065
+ $X2=2.71 $Y2=1.065
r163 35 69 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=2.625 $Y=1.065
+ $X2=2.275 $Y2=1.065
r164 31 68 21.0727 $w=1.98e-07 $l=3.8e-07 $layer=LI1_cond $X=1.78 $Y=1.08
+ $X2=2.16 $Y2=1.08
r165 31 66 9.43135 $w=1.98e-07 $l=1.65e-07 $layer=LI1_cond $X=1.78 $Y=1.08
+ $X2=1.615 $Y2=1.08
r166 31 33 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=1.78 $Y=0.98
+ $X2=1.78 $Y2=0.515
r167 30 66 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.945 $Y=1.095
+ $X2=1.615 $Y2=1.095
r168 25 30 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.78 $Y=1.01
+ $X2=0.945 $Y2=1.095
r169 25 27 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=0.78 $Y=1.01
+ $X2=0.78 $Y2=0.515
r170 8 41 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=3.405
+ $Y=1.84 $X2=3.555 $Y2=1.985
r171 7 39 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.505
+ $Y=1.84 $X2=2.655 $Y2=1.985
r172 6 63 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.63
+ $Y=0.37 $X2=5.77 $Y2=0.515
r173 5 57 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.5
+ $Y=0.37 $X2=4.64 $Y2=0.515
r174 4 51 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.5
+ $Y=0.37 $X2=3.64 $Y2=0.515
r175 3 45 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.57
+ $Y=0.37 $X2=2.71 $Y2=0.515
r176 2 33 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.64
+ $Y=0.37 $X2=1.78 $Y2=0.515
r177 1 27 91 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=2 $X=0.615
+ $Y=0.37 $X2=0.78 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__NOR3B_4%VPWR 1 2 3 4 15 19 23 27 29 31 33 41 46 51
+ 57 60 63 67
r94 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r95 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r96 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r97 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r98 55 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.44 $Y2=3.33
r99 55 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6.48 $Y2=3.33
r100 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r101 52 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.58 $Y=3.33
+ $X2=6.415 $Y2=3.33
r102 52 54 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=6.58 $Y=3.33
+ $X2=6.96 $Y2=3.33
r103 51 66 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=7.235 $Y=3.33
+ $X2=7.457 $Y2=3.33
r104 51 54 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=7.235 $Y=3.33
+ $X2=6.96 $Y2=3.33
r105 50 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r106 50 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=5.52
+ $Y2=3.33
r107 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r108 47 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.63 $Y=3.33
+ $X2=5.465 $Y2=3.33
r109 47 49 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=5.63 $Y=3.33 $X2=6
+ $Y2=3.33
r110 46 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.25 $Y=3.33
+ $X2=6.415 $Y2=3.33
r111 46 49 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=6.25 $Y=3.33 $X2=6
+ $Y2=3.33
r112 45 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r113 45 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r114 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r115 42 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.73 $Y=3.33
+ $X2=4.565 $Y2=3.33
r116 42 44 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=4.73 $Y=3.33
+ $X2=5.04 $Y2=3.33
r117 41 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.3 $Y=3.33
+ $X2=5.465 $Y2=3.33
r118 41 44 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=5.3 $Y=3.33
+ $X2=5.04 $Y2=3.33
r119 40 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r120 39 40 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r121 35 39 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=4.08 $Y2=3.33
r122 35 36 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r123 33 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.4 $Y=3.33
+ $X2=4.565 $Y2=3.33
r124 33 39 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=4.4 $Y=3.33 $X2=4.08
+ $Y2=3.33
r125 31 40 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=4.08 $Y2=3.33
r126 31 36 1.00344 $w=4.9e-07 $l=3.6e-06 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=0.24 $Y2=3.33
r127 27 66 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=7.4 $Y=3.245
+ $X2=7.457 $Y2=3.33
r128 27 29 37.8909 $w=3.28e-07 $l=1.085e-06 $layer=LI1_cond $X=7.4 $Y=3.245
+ $X2=7.4 $Y2=2.16
r129 23 26 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=6.415 $Y=2.145
+ $X2=6.415 $Y2=2.825
r130 21 63 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.415 $Y=3.245
+ $X2=6.415 $Y2=3.33
r131 21 26 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=6.415 $Y=3.245
+ $X2=6.415 $Y2=2.825
r132 17 60 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.465 $Y=3.245
+ $X2=5.465 $Y2=3.33
r133 17 19 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=5.465 $Y=3.245
+ $X2=5.465 $Y2=2.485
r134 13 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.565 $Y=3.245
+ $X2=4.565 $Y2=3.33
r135 13 15 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=4.565 $Y=3.245
+ $X2=4.565 $Y2=2.745
r136 4 29 300 $w=1.7e-07 $l=3.87814e-07 $layer=licon1_PDIFF $count=2 $X=7.25
+ $Y=1.84 $X2=7.4 $Y2=2.16
r137 3 26 600 $w=1.7e-07 $l=1.08038e-06 $layer=licon1_PDIFF $count=1 $X=6.215
+ $Y=1.84 $X2=6.415 $Y2=2.825
r138 3 23 300 $w=1.7e-07 $l=3.9246e-07 $layer=licon1_PDIFF $count=2 $X=6.215
+ $Y=1.84 $X2=6.415 $Y2=2.145
r139 2 19 300 $w=1.7e-07 $l=7.16083e-07 $layer=licon1_PDIFF $count=2 $X=5.315
+ $Y=1.84 $X2=5.465 $Y2=2.485
r140 1 15 600 $w=1.7e-07 $l=9.74808e-07 $layer=licon1_PDIFF $count=1 $X=4.42
+ $Y=1.84 $X2=4.565 $Y2=2.745
.ends

.subckt PM_SKY130_FD_SC_LS__NOR3B_4%VGND 1 2 3 4 5 6 7 22 24 28 30 34 38 42 44
+ 48 52 55 56 57 59 64 69 82 83 89 92 95 98 101
r109 101 102 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r110 99 102 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0
+ $X2=5.04 $Y2=0
r111 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r112 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r113 92 93 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r114 90 93 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r115 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r116 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r117 82 83 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r118 80 83 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=7.44
+ $Y2=0
r119 79 82 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=6.48 $Y=0 $X2=7.44
+ $Y2=0
r120 79 80 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r121 77 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r122 77 102 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.04
+ $Y2=0
r123 76 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6 $Y2=0
r124 74 101 10.7288 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=5.435 $Y=0
+ $X2=5.205 $Y2=0
r125 74 76 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=5.435 $Y=0 $X2=6
+ $Y2=0
r126 73 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r127 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r128 70 95 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.305 $Y=0 $X2=3.14
+ $Y2=0
r129 70 72 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.305 $Y=0 $X2=3.6
+ $Y2=0
r130 69 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.975 $Y=0 $X2=4.14
+ $Y2=0
r131 69 72 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=3.975 $Y=0 $X2=3.6
+ $Y2=0
r132 68 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r133 68 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r134 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r135 65 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.445 $Y=0 $X2=2.28
+ $Y2=0
r136 65 67 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=2.445 $Y=0
+ $X2=2.64 $Y2=0
r137 64 95 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.975 $Y=0 $X2=3.14
+ $Y2=0
r138 64 67 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.975 $Y=0
+ $X2=2.64 $Y2=0
r139 63 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r140 63 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r141 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r142 60 86 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=0
+ $X2=0.222 $Y2=0
r143 60 62 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=0
+ $X2=0.72 $Y2=0
r144 59 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.115 $Y=0 $X2=1.28
+ $Y2=0
r145 59 62 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.115 $Y=0
+ $X2=0.72 $Y2=0
r146 57 99 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=0
+ $X2=4.08 $Y2=0
r147 57 73 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=0 $X2=3.6
+ $Y2=0
r148 55 76 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=6.105 $Y=0 $X2=6
+ $Y2=0
r149 55 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.105 $Y=0 $X2=6.27
+ $Y2=0
r150 54 79 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=6.435 $Y=0 $X2=6.48
+ $Y2=0
r151 54 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.435 $Y=0 $X2=6.27
+ $Y2=0
r152 50 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.27 $Y=0.085
+ $X2=6.27 $Y2=0
r153 50 52 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=6.27 $Y=0.085
+ $X2=6.27 $Y2=0.515
r154 46 101 1.85547 $w=4.6e-07 $l=8.5e-08 $layer=LI1_cond $X=5.205 $Y=0.085
+ $X2=5.205 $Y2=0
r155 46 48 11.1807 $w=4.58e-07 $l=4.3e-07 $layer=LI1_cond $X=5.205 $Y=0.085
+ $X2=5.205 $Y2=0.515
r156 45 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.305 $Y=0 $X2=4.14
+ $Y2=0
r157 44 101 10.7288 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=4.975 $Y=0
+ $X2=5.205 $Y2=0
r158 44 45 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.975 $Y=0
+ $X2=4.305 $Y2=0
r159 40 98 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.14 $Y=0.085
+ $X2=4.14 $Y2=0
r160 40 42 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=4.14 $Y=0.085
+ $X2=4.14 $Y2=0.53
r161 36 95 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.14 $Y=0.085
+ $X2=3.14 $Y2=0
r162 36 38 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=3.14 $Y=0.085
+ $X2=3.14 $Y2=0.645
r163 32 92 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.28 $Y=0.085
+ $X2=2.28 $Y2=0
r164 32 34 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=2.28 $Y=0.085
+ $X2=2.28 $Y2=0.645
r165 31 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.445 $Y=0 $X2=1.28
+ $Y2=0
r166 30 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.115 $Y=0 $X2=2.28
+ $Y2=0
r167 30 31 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.115 $Y=0
+ $X2=1.445 $Y2=0
r168 26 89 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.28 $Y=0.085
+ $X2=1.28 $Y2=0
r169 26 28 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=1.28 $Y=0.085
+ $X2=1.28 $Y2=0.675
r170 22 86 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.222 $Y2=0
r171 22 24 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.28 $Y2=0.515
r172 7 52 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.13
+ $Y=0.37 $X2=6.27 $Y2=0.515
r173 6 48 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=4.93
+ $Y=0.37 $X2=5.205 $Y2=0.515
r174 5 42 182 $w=1.7e-07 $l=2.78747e-07 $layer=licon1_NDIFF $count=1 $X=3.93
+ $Y=0.37 $X2=4.14 $Y2=0.53
r175 4 38 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=3
+ $Y=0.37 $X2=3.14 $Y2=0.645
r176 3 34 182 $w=1.7e-07 $l=3.65205e-07 $layer=licon1_NDIFF $count=1 $X=2.07
+ $Y=0.37 $X2=2.28 $Y2=0.645
r177 2 28 182 $w=1.7e-07 $l=3.96327e-07 $layer=licon1_NDIFF $count=1 $X=1.07
+ $Y=0.37 $X2=1.28 $Y2=0.675
r178 1 24 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

