* File: sky130_fd_sc_ls__a41oi_1.pxi.spice
* Created: Wed Sep  2 10:53:46 2020
* 
x_PM_SKY130_FD_SC_LS__A41OI_1%B1 N_B1_M1008_g N_B1_c_50_n N_B1_M1007_g B1
+ N_B1_c_51_n PM_SKY130_FD_SC_LS__A41OI_1%B1
x_PM_SKY130_FD_SC_LS__A41OI_1%A4 N_A4_c_76_n N_A4_M1006_g N_A4_M1002_g A4
+ N_A4_c_74_n N_A4_c_75_n PM_SKY130_FD_SC_LS__A41OI_1%A4
x_PM_SKY130_FD_SC_LS__A41OI_1%A3 N_A3_M1003_g N_A3_c_111_n N_A3_M1001_g A3
+ N_A3_c_112_n PM_SKY130_FD_SC_LS__A41OI_1%A3
x_PM_SKY130_FD_SC_LS__A41OI_1%A2 N_A2_M1009_g N_A2_c_139_n N_A2_M1004_g A2
+ PM_SKY130_FD_SC_LS__A41OI_1%A2
x_PM_SKY130_FD_SC_LS__A41OI_1%A1 N_A1_M1000_g N_A1_c_168_n N_A1_M1005_g A1
+ N_A1_c_169_n PM_SKY130_FD_SC_LS__A41OI_1%A1
x_PM_SKY130_FD_SC_LS__A41OI_1%Y N_Y_M1008_s N_Y_M1000_d N_Y_M1007_s N_Y_c_191_n
+ N_Y_c_196_n N_Y_c_192_n N_Y_c_193_n N_Y_c_194_n N_Y_c_197_n Y
+ PM_SKY130_FD_SC_LS__A41OI_1%Y
x_PM_SKY130_FD_SC_LS__A41OI_1%A_116_368# N_A_116_368#_M1007_d
+ N_A_116_368#_M1001_d N_A_116_368#_M1005_d N_A_116_368#_c_249_n
+ N_A_116_368#_c_251_n N_A_116_368#_c_245_n N_A_116_368#_c_246_n
+ N_A_116_368#_c_247_n PM_SKY130_FD_SC_LS__A41OI_1%A_116_368#
x_PM_SKY130_FD_SC_LS__A41OI_1%VPWR N_VPWR_M1006_d N_VPWR_M1004_d N_VPWR_c_282_n
+ VPWR N_VPWR_c_283_n N_VPWR_c_284_n N_VPWR_c_285_n N_VPWR_c_281_n
+ N_VPWR_c_287_n N_VPWR_c_288_n PM_SKY130_FD_SC_LS__A41OI_1%VPWR
x_PM_SKY130_FD_SC_LS__A41OI_1%VGND N_VGND_M1008_d VGND N_VGND_c_318_n
+ N_VGND_c_319_n N_VGND_c_320_n PM_SKY130_FD_SC_LS__A41OI_1%VGND
cc_1 VNB N_B1_M1008_g 0.0333332f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_B1_c_50_n 0.0624499f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_3 VNB N_B1_c_51_n 0.00430714f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_4 VNB N_A4_M1002_g 0.0271041f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_5 VNB N_A4_c_74_n 0.0364966f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_6 VNB N_A4_c_75_n 0.00234054f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_7 VNB N_A3_M1003_g 0.0260165f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_8 VNB N_A3_c_111_n 0.0250772f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_9 VNB N_A3_c_112_n 0.00452292f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_10 VNB N_A2_M1009_g 0.0284012f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_11 VNB N_A2_c_139_n 0.0225726f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_12 VNB A2 0.00682758f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_13 VNB N_A1_M1000_g 0.031841f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_14 VNB N_A1_c_168_n 0.0612826f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_15 VNB N_A1_c_169_n 0.0051843f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_16 VNB N_Y_c_191_n 0.0258829f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_17 VNB N_Y_c_192_n 0.0345375f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_Y_c_193_n 0.0102107f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_Y_c_194_n 0.02581f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB Y 0.0120831f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_VPWR_c_281_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_318_n 0.0412642f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_23 VNB N_VGND_c_319_n 0.0662801f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_24 VNB N_VGND_c_320_n 0.240368f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VPB N_B1_c_50_n 0.0295305f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_26 VPB N_B1_c_51_n 0.00775466f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_27 VPB N_A4_c_76_n 0.0185664f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.3
cc_28 VPB N_A4_c_74_n 0.0162609f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_29 VPB N_A4_c_75_n 0.00327171f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_30 VPB N_A3_c_111_n 0.0285609f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_31 VPB N_A3_c_112_n 0.00384627f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_32 VPB N_A2_c_139_n 0.0274249f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_33 VPB A2 0.005546f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_34 VPB N_A1_c_168_n 0.0300188f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_35 VPB N_A1_c_169_n 0.00775819f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_36 VPB N_Y_c_196_n 0.0354773f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_37 VPB N_Y_c_197_n 0.00719835f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_38 VPB Y 0.00356234f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_39 VPB N_A_116_368#_c_245_n 0.0142315f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_40 VPB N_A_116_368#_c_246_n 0.0289409f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_41 VPB N_A_116_368#_c_247_n 0.00289794f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_42 VPB N_VPWR_c_282_n 0.00912032f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_43 VPB N_VPWR_c_283_n 0.0325002f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_44 VPB N_VPWR_c_284_n 0.0195071f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_45 VPB N_VPWR_c_285_n 0.0191515f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_281_n 0.0704604f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_287_n 0.0223348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_288_n 0.00651392f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 N_B1_c_50_n N_A4_c_76_n 0.0272074f $X=0.505 $Y=1.765 $X2=-0.19 $Y2=-0.245
cc_50 N_B1_M1008_g N_A4_M1002_g 0.0105574f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_51 N_B1_c_50_n N_A4_M1002_g 5.70607e-19 $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_52 N_B1_c_50_n N_A4_c_74_n 0.0137203f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_53 N_B1_M1008_g N_Y_c_191_n 0.0175621f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_54 N_B1_c_50_n N_Y_c_196_n 0.0106511f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_55 N_B1_M1008_g N_Y_c_193_n 0.0179726f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_56 N_B1_c_50_n N_Y_c_193_n 0.00315313f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_57 N_B1_c_51_n N_Y_c_193_n 0.0247471f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_58 N_B1_c_50_n N_Y_c_197_n 0.0181182f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_59 N_B1_c_51_n N_Y_c_197_n 0.0236452f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_60 N_B1_M1008_g Y 0.00516025f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_61 N_B1_c_50_n Y 0.00708613f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_62 N_B1_c_51_n Y 0.0368805f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_63 N_B1_c_50_n N_A_116_368#_c_247_n 0.00283124f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_64 N_B1_c_50_n N_VPWR_c_283_n 0.00445602f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_65 N_B1_c_50_n N_VPWR_c_281_n 0.0086236f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_66 N_B1_M1008_g N_VGND_c_318_n 0.00847491f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_67 N_B1_M1008_g N_VGND_c_320_n 0.00826401f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_68 N_A4_M1002_g N_A3_M1003_g 0.0399236f $X=1.31 $Y=0.74 $X2=0 $Y2=0
cc_69 N_A4_c_76_n N_A3_c_111_n 0.012762f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_70 N_A4_c_74_n N_A3_c_111_n 0.0408635f $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_71 N_A4_c_75_n N_A3_c_111_n 6.52107e-19 $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_72 N_A4_c_74_n N_A3_c_112_n 0.00259287f $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_73 N_A4_c_75_n N_A3_c_112_n 0.0279517f $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_74 N_A4_c_76_n N_Y_c_196_n 4.58902e-19 $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_75 N_A4_M1002_g N_Y_c_192_n 0.0171807f $X=1.31 $Y=0.74 $X2=0 $Y2=0
cc_76 N_A4_c_74_n N_Y_c_192_n 0.0050608f $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_77 N_A4_c_75_n N_Y_c_192_n 0.0204317f $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_78 N_A4_c_76_n N_Y_c_197_n 0.00169696f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_79 N_A4_c_76_n Y 0.00433684f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_80 N_A4_M1002_g Y 0.00420733f $X=1.31 $Y=0.74 $X2=0 $Y2=0
cc_81 N_A4_c_74_n Y 0.00349554f $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_82 N_A4_c_75_n Y 0.0330364f $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_83 N_A4_c_74_n N_A_116_368#_c_249_n 0.00237233f $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_84 N_A4_c_75_n N_A_116_368#_c_249_n 0.00491597f $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_85 N_A4_c_76_n N_A_116_368#_c_251_n 0.0159143f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_86 N_A4_c_74_n N_A_116_368#_c_251_n 9.36874e-19 $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_87 N_A4_c_75_n N_A_116_368#_c_251_n 0.0161156f $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_88 N_A4_c_76_n N_A_116_368#_c_247_n 0.00752062f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_89 N_A4_c_76_n N_VPWR_c_283_n 0.00445602f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_90 N_A4_c_76_n N_VPWR_c_281_n 0.00860009f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_91 N_A4_c_76_n N_VPWR_c_287_n 0.0089138f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_92 N_A4_M1002_g N_VGND_c_318_n 0.0118628f $X=1.31 $Y=0.74 $X2=0 $Y2=0
cc_93 N_A4_M1002_g N_VGND_c_319_n 0.00384553f $X=1.31 $Y=0.74 $X2=0 $Y2=0
cc_94 N_A4_M1002_g N_VGND_c_320_n 0.0075725f $X=1.31 $Y=0.74 $X2=0 $Y2=0
cc_95 N_A3_M1003_g N_A2_M1009_g 0.0373965f $X=1.7 $Y=0.74 $X2=0 $Y2=0
cc_96 N_A3_c_111_n N_A2_c_139_n 0.0599784f $X=1.845 $Y=1.765 $X2=0 $Y2=0
cc_97 N_A3_c_112_n N_A2_c_139_n 7.94787e-19 $X=1.79 $Y=1.515 $X2=0 $Y2=0
cc_98 N_A3_c_111_n A2 0.00160421f $X=1.845 $Y=1.765 $X2=0 $Y2=0
cc_99 N_A3_c_112_n A2 0.0266982f $X=1.79 $Y=1.515 $X2=0 $Y2=0
cc_100 N_A3_M1003_g N_Y_c_192_n 0.0157189f $X=1.7 $Y=0.74 $X2=0 $Y2=0
cc_101 N_A3_c_111_n N_Y_c_192_n 0.00118269f $X=1.845 $Y=1.765 $X2=0 $Y2=0
cc_102 N_A3_c_112_n N_Y_c_192_n 0.024303f $X=1.79 $Y=1.515 $X2=0 $Y2=0
cc_103 N_A3_c_111_n N_A_116_368#_c_249_n 0.0210076f $X=1.845 $Y=1.765 $X2=0
+ $Y2=0
cc_104 N_A3_c_112_n N_A_116_368#_c_249_n 0.0278479f $X=1.79 $Y=1.515 $X2=0 $Y2=0
cc_105 N_A3_c_111_n N_A_116_368#_c_251_n 0.00355759f $X=1.845 $Y=1.765 $X2=0
+ $Y2=0
cc_106 N_A3_c_111_n N_VPWR_c_284_n 0.00413917f $X=1.845 $Y=1.765 $X2=0 $Y2=0
cc_107 N_A3_c_111_n N_VPWR_c_281_n 0.00813195f $X=1.845 $Y=1.765 $X2=0 $Y2=0
cc_108 N_A3_c_111_n N_VPWR_c_287_n 0.0167477f $X=1.845 $Y=1.765 $X2=0 $Y2=0
cc_109 N_A3_M1003_g N_VGND_c_318_n 0.00217763f $X=1.7 $Y=0.74 $X2=0 $Y2=0
cc_110 N_A3_M1003_g N_VGND_c_319_n 0.00461464f $X=1.7 $Y=0.74 $X2=0 $Y2=0
cc_111 N_A3_M1003_g N_VGND_c_320_n 0.0091028f $X=1.7 $Y=0.74 $X2=0 $Y2=0
cc_112 N_A2_M1009_g N_A1_M1000_g 0.0342424f $X=2.27 $Y=0.74 $X2=0 $Y2=0
cc_113 N_A2_c_139_n N_A1_c_168_n 0.0529159f $X=2.295 $Y=1.765 $X2=0 $Y2=0
cc_114 A2 N_A1_c_168_n 0.00401962f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_115 N_A2_M1009_g N_A1_c_169_n 2.13129e-19 $X=2.27 $Y=0.74 $X2=0 $Y2=0
cc_116 N_A2_c_139_n N_A1_c_169_n 2.84133e-19 $X=2.295 $Y=1.765 $X2=0 $Y2=0
cc_117 A2 N_A1_c_169_n 0.0354768f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_118 N_A2_M1009_g N_Y_c_192_n 0.0166695f $X=2.27 $Y=0.74 $X2=0 $Y2=0
cc_119 N_A2_c_139_n N_Y_c_192_n 0.00401243f $X=2.295 $Y=1.765 $X2=0 $Y2=0
cc_120 A2 N_Y_c_192_n 0.0358367f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_121 N_A2_M1009_g N_Y_c_194_n 0.00278148f $X=2.27 $Y=0.74 $X2=0 $Y2=0
cc_122 N_A2_c_139_n N_A_116_368#_c_249_n 0.0199601f $X=2.295 $Y=1.765 $X2=0
+ $Y2=0
cc_123 A2 N_A_116_368#_c_249_n 0.0411687f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_124 N_A2_c_139_n N_A_116_368#_c_246_n 8.68268e-19 $X=2.295 $Y=1.765 $X2=0
+ $Y2=0
cc_125 N_A2_c_139_n N_VPWR_c_282_n 0.00512198f $X=2.295 $Y=1.765 $X2=0 $Y2=0
cc_126 N_A2_c_139_n N_VPWR_c_284_n 0.00461464f $X=2.295 $Y=1.765 $X2=0 $Y2=0
cc_127 N_A2_c_139_n N_VPWR_c_281_n 0.00909345f $X=2.295 $Y=1.765 $X2=0 $Y2=0
cc_128 N_A2_c_139_n N_VPWR_c_287_n 0.00189413f $X=2.295 $Y=1.765 $X2=0 $Y2=0
cc_129 N_A2_M1009_g N_VGND_c_319_n 0.00461464f $X=2.27 $Y=0.74 $X2=0 $Y2=0
cc_130 N_A2_M1009_g N_VGND_c_320_n 0.00911823f $X=2.27 $Y=0.74 $X2=0 $Y2=0
cc_131 N_A1_M1000_g N_Y_c_192_n 0.0176301f $X=2.84 $Y=0.74 $X2=0 $Y2=0
cc_132 N_A1_c_168_n N_Y_c_192_n 0.00285817f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_133 N_A1_c_169_n N_Y_c_192_n 0.025569f $X=3.09 $Y=1.465 $X2=0 $Y2=0
cc_134 N_A1_M1000_g N_Y_c_194_n 0.0142362f $X=2.84 $Y=0.74 $X2=0 $Y2=0
cc_135 N_A1_c_168_n N_A_116_368#_c_249_n 0.0223648f $X=2.855 $Y=1.765 $X2=0
+ $Y2=0
cc_136 N_A1_c_168_n N_A_116_368#_c_245_n 0.00255725f $X=2.855 $Y=1.765 $X2=0
+ $Y2=0
cc_137 N_A1_c_169_n N_A_116_368#_c_245_n 0.025958f $X=3.09 $Y=1.465 $X2=0 $Y2=0
cc_138 N_A1_c_168_n N_A_116_368#_c_246_n 0.00887931f $X=2.855 $Y=1.765 $X2=0
+ $Y2=0
cc_139 N_A1_c_168_n N_VPWR_c_282_n 0.00645753f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_140 N_A1_c_168_n N_VPWR_c_285_n 0.00445602f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_141 N_A1_c_168_n N_VPWR_c_281_n 0.00861394f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_142 N_A1_M1000_g N_VGND_c_319_n 0.00434272f $X=2.84 $Y=0.74 $X2=0 $Y2=0
cc_143 N_A1_M1000_g N_VGND_c_320_n 0.00826262f $X=2.84 $Y=0.74 $X2=0 $Y2=0
cc_144 N_Y_c_197_n N_A_116_368#_M1007_d 0.00506001f $X=0.72 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_145 Y N_A_116_368#_M1007_d 0.00225461f $X=0.635 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_146 N_Y_c_197_n N_A_116_368#_c_251_n 0.0160918f $X=0.72 $Y=1.95 $X2=0 $Y2=0
cc_147 N_Y_c_196_n N_A_116_368#_c_247_n 0.0203021f $X=0.28 $Y=2.815 $X2=0 $Y2=0
cc_148 N_Y_c_196_n N_VPWR_c_283_n 0.0145938f $X=0.28 $Y=2.815 $X2=0 $Y2=0
cc_149 N_Y_c_196_n N_VPWR_c_281_n 0.0120466f $X=0.28 $Y=2.815 $X2=0 $Y2=0
cc_150 N_Y_c_192_n N_VGND_M1008_d 0.00637083f $X=2.89 $Y=1.045 $X2=-0.19
+ $Y2=-0.245
cc_151 N_Y_c_193_n N_VGND_M1008_d 0.0034772f $X=0.835 $Y=1.045 $X2=-0.19
+ $Y2=-0.245
cc_152 N_Y_c_191_n N_VGND_c_318_n 0.0277067f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_153 N_Y_c_193_n N_VGND_c_318_n 0.0321701f $X=0.835 $Y=1.045 $X2=0 $Y2=0
cc_154 N_Y_c_194_n N_VGND_c_319_n 0.0145639f $X=3.055 $Y=0.515 $X2=0 $Y2=0
cc_155 N_Y_c_191_n N_VGND_c_320_n 0.0119539f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_156 N_Y_c_194_n N_VGND_c_320_n 0.0119984f $X=3.055 $Y=0.515 $X2=0 $Y2=0
cc_157 N_Y_c_192_n A_277_74# 0.0048076f $X=2.89 $Y=1.045 $X2=-0.19 $Y2=-0.245
cc_158 N_Y_c_192_n A_355_74# 0.0121704f $X=2.89 $Y=1.045 $X2=-0.19 $Y2=-0.245
cc_159 N_Y_c_192_n A_469_74# 0.0121704f $X=2.89 $Y=1.045 $X2=-0.19 $Y2=-0.245
cc_160 N_A_116_368#_c_249_n N_VPWR_M1006_d 0.0214673f $X=2.915 $Y=2.12 $X2=-0.19
+ $Y2=1.66
cc_161 N_A_116_368#_c_251_n N_VPWR_M1006_d 0.00726186f $X=1.275 $Y=2.12
+ $X2=-0.19 $Y2=1.66
cc_162 N_A_116_368#_c_249_n N_VPWR_M1004_d 0.00717524f $X=2.915 $Y=2.12 $X2=0
+ $Y2=0
cc_163 N_A_116_368#_c_249_n N_VPWR_c_282_n 0.0252617f $X=2.915 $Y=2.12 $X2=0
+ $Y2=0
cc_164 N_A_116_368#_c_246_n N_VPWR_c_282_n 0.0203057f $X=3.08 $Y=2.815 $X2=0
+ $Y2=0
cc_165 N_A_116_368#_c_247_n N_VPWR_c_283_n 0.0146094f $X=0.78 $Y=2.375 $X2=0
+ $Y2=0
cc_166 N_A_116_368#_c_246_n N_VPWR_c_285_n 0.0145938f $X=3.08 $Y=2.815 $X2=0
+ $Y2=0
cc_167 N_A_116_368#_c_246_n N_VPWR_c_281_n 0.0120466f $X=3.08 $Y=2.815 $X2=0
+ $Y2=0
cc_168 N_A_116_368#_c_247_n N_VPWR_c_281_n 0.0120527f $X=0.78 $Y=2.375 $X2=0
+ $Y2=0
cc_169 N_A_116_368#_c_249_n N_VPWR_c_287_n 0.0327457f $X=2.915 $Y=2.12 $X2=0
+ $Y2=0
cc_170 N_A_116_368#_c_251_n N_VPWR_c_287_n 0.0121825f $X=1.275 $Y=2.12 $X2=0
+ $Y2=0
cc_171 N_A_116_368#_c_247_n N_VPWR_c_287_n 0.0197997f $X=0.78 $Y=2.375 $X2=0
+ $Y2=0
