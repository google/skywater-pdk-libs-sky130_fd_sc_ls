* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__nor3_1 A B C VGND VNB VPB VPWR Y
M1000 Y C a_198_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=3.192e+11p pd=2.81e+06u as=4.032e+11p ps=2.96e+06u
M1001 a_198_368# B a_114_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.024e+11p ps=2.78e+06u
M1002 Y C VGND VNB nshort w=740000u l=150000u
+  ad=4.181e+11p pd=4.09e+06u as=4.699e+11p ps=4.23e+06u
M1003 a_114_368# A VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.192e+11p ps=2.81e+06u
M1004 Y A VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND B Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
