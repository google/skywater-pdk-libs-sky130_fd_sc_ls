# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ls__or2b_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ls__or2b_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.035000 1.350000 2.365000 1.780000 ;
    END
  END A
  PIN B_N
    ANTENNAGATEAREA  0.208500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.350000 0.550000 1.780000 ;
    END
  END B_N
  PIN X
    ANTENNADIFFAREA  0.787700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.060000 0.350000 1.390000 1.130000 ;
        RECT 1.060000 1.130000 1.230000 1.820000 ;
        RECT 1.060000 1.820000 1.645000 2.070000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 3.360000 0.085000 ;
        RECT 0.630000  0.085000 0.880000 0.840000 ;
        RECT 1.560000  0.085000 2.235000 0.810000 ;
        RECT 2.915000  0.085000 3.245000 0.810000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 3.360000 3.415000 ;
        RECT 0.650000 2.580000 0.980000 3.245000 ;
        RECT 1.765000 2.580000 2.095000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.115000 1.950000 0.890000 2.240000 ;
      RECT 0.115000 2.240000 2.705000 2.410000 ;
      RECT 0.115000 2.410000 0.445000 2.700000 ;
      RECT 0.120000 0.540000 0.450000 1.010000 ;
      RECT 0.120000 1.010000 0.890000 1.180000 ;
      RECT 0.720000 1.180000 0.890000 1.950000 ;
      RECT 1.465000 1.300000 1.795000 1.630000 ;
      RECT 1.625000 0.980000 3.275000 1.150000 ;
      RECT 1.625000 1.150000 1.795000 1.300000 ;
      RECT 2.405000 0.350000 2.735000 0.980000 ;
      RECT 2.535000 1.320000 2.935000 1.650000 ;
      RECT 2.535000 1.650000 2.705000 2.240000 ;
      RECT 2.875000 1.820000 3.275000 2.860000 ;
      RECT 3.105000 1.150000 3.275000 1.820000 ;
  END
END sky130_fd_sc_ls__or2b_2
