* File: sky130_fd_sc_ls__fah_4.pex.spice
* Created: Fri Aug 28 13:26:06 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__FAH_4%A 3 5 7 10 12 14 15 21 22
c46 5 0 1.1412e-19 $X=0.505 $Y=1.885
c47 3 0 1.40087e-19 $X=0.495 $Y=0.69
r48 21 23 3.23056 $w=3.73e-07 $l=2.5e-08 $layer=POLY_cond $X=0.93 $Y=1.677
+ $X2=0.955 $Y2=1.677
r49 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.93
+ $Y=1.635 $X2=0.93 $Y2=1.635
r50 19 21 0.646113 $w=3.73e-07 $l=5e-09 $layer=POLY_cond $X=0.925 $Y=1.677
+ $X2=0.93 $Y2=1.677
r51 18 19 54.2735 $w=3.73e-07 $l=4.2e-07 $layer=POLY_cond $X=0.505 $Y=1.677
+ $X2=0.925 $Y2=1.677
r52 17 18 1.29223 $w=3.73e-07 $l=1e-08 $layer=POLY_cond $X=0.495 $Y=1.677
+ $X2=0.505 $Y2=1.677
r53 15 22 8.34528 $w=2.88e-07 $l=2.1e-07 $layer=LI1_cond $X=0.72 $Y=1.655
+ $X2=0.93 $Y2=1.655
r54 12 23 24.162 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.955 $Y=1.885
+ $X2=0.955 $Y2=1.677
r55 12 14 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.955 $Y=1.885
+ $X2=0.955 $Y2=2.46
r56 8 19 24.162 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.925 $Y=1.47
+ $X2=0.925 $Y2=1.677
r57 8 10 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=0.925 $Y=1.47
+ $X2=0.925 $Y2=0.69
r58 5 18 24.162 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.505 $Y=1.885
+ $X2=0.505 $Y2=1.677
r59 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.505 $Y=1.885
+ $X2=0.505 $Y2=2.46
r60 1 17 24.162 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.495 $Y=1.47
+ $X2=0.495 $Y2=1.677
r61 1 3 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=0.495 $Y=1.47
+ $X2=0.495 $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_LS__FAH_4%A_27_74# 1 2 7 10 11 13 14 16 17 20 24 26 30
+ 32 33 34 40
c77 40 0 5.85186e-20 $X=1.5 $Y=1.395
r78 38 40 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.5 $Y=1.485 $X2=1.5
+ $Y2=1.395
r79 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.5
+ $Y=1.485 $X2=1.5 $Y2=1.485
r80 34 37 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=1.5 $Y=1.255 $X2=1.5
+ $Y2=1.485
r81 31 32 2.36881 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=0.365 $Y=1.255
+ $X2=0.225 $Y2=1.255
r82 30 34 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.335 $Y=1.255
+ $X2=1.5 $Y2=1.255
r83 30 31 63.2834 $w=1.68e-07 $l=9.7e-07 $layer=LI1_cond $X=1.335 $Y=1.255
+ $X2=0.365 $Y2=1.255
r84 26 28 27.9879 $w=2.78e-07 $l=6.8e-07 $layer=LI1_cond $X=0.225 $Y=2.135
+ $X2=0.225 $Y2=2.815
r85 24 33 7.52792 $w=2.78e-07 $l=1.4e-07 $layer=LI1_cond $X=0.225 $Y=2.11
+ $X2=0.225 $Y2=1.97
r86 24 26 1.02897 $w=2.78e-07 $l=2.5e-08 $layer=LI1_cond $X=0.225 $Y=2.11
+ $X2=0.225 $Y2=2.135
r87 22 32 4.06715 $w=2.25e-07 $l=1.09087e-07 $layer=LI1_cond $X=0.17 $Y=1.34
+ $X2=0.225 $Y2=1.255
r88 22 33 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=0.17 $Y=1.34
+ $X2=0.17 $Y2=1.97
r89 18 32 4.06715 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=0.225 $Y=1.17
+ $X2=0.225 $Y2=1.255
r90 18 20 26.9589 $w=2.78e-07 $l=6.55e-07 $layer=LI1_cond $X=0.225 $Y=1.17
+ $X2=0.225 $Y2=0.515
r91 14 17 18.8402 $w=1.65e-07 $l=9.40744e-08 $layer=POLY_cond $X=2.13 $Y=1.32
+ $X2=2.087 $Y2=1.395
r92 14 16 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.13 $Y=1.32 $X2=2.13
+ $Y2=0.84
r93 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.06 $Y=1.735
+ $X2=2.06 $Y2=2.37
r94 10 11 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.06 $Y=1.645 $X2=2.06
+ $Y2=1.735
r95 9 17 18.8402 $w=1.65e-07 $l=8.74643e-08 $layer=POLY_cond $X=2.06 $Y=1.47
+ $X2=2.087 $Y2=1.395
r96 9 10 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=2.06 $Y=1.47
+ $X2=2.06 $Y2=1.645
r97 8 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.665 $Y=1.395
+ $X2=1.5 $Y2=1.395
r98 7 17 6.66866 $w=1.5e-07 $l=1.17e-07 $layer=POLY_cond $X=1.97 $Y=1.395
+ $X2=2.087 $Y2=1.395
r99 7 8 156.394 $w=1.5e-07 $l=3.05e-07 $layer=POLY_cond $X=1.97 $Y=1.395
+ $X2=1.665 $Y2=1.395
r100 2 28 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.28 $Y2=2.815
r101 2 26 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.28 $Y2=2.135
r102 1 20 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__FAH_4%A_586_257# 1 2 3 10 11 12 14 18 19 20 22 24 25
+ 27 31 34 35 39 41 42 43 44 46 48 50 52
c178 50 0 2.90544e-20 $X=5.94 $Y=2.815
c179 48 0 1.35704e-20 $X=5.94 $Y=2.12
c180 35 0 1.58586e-19 $X=4.385 $Y=0.79
c181 24 0 4.11294e-20 $X=4.015 $Y=0.97
c182 22 0 2.46839e-19 $X=4.015 $Y=1.365
c183 12 0 1.07671e-19 $X=3.02 $Y=1.735
r184 48 54 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.94 $Y=2.12
+ $X2=5.94 $Y2=2.035
r185 48 50 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=5.94 $Y=2.12
+ $X2=5.94 $Y2=2.815
r186 44 46 171.257 $w=1.68e-07 $l=2.625e-06 $layer=LI1_cond $X=5.405 $Y=0.34
+ $X2=8.03 $Y2=0.34
r187 42 54 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.855 $Y=2.035
+ $X2=5.94 $Y2=2.035
r188 42 43 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=5.855 $Y=2.035
+ $X2=5.265 $Y2=2.035
r189 41 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.18 $Y=1.95
+ $X2=5.265 $Y2=2.035
r190 40 52 3.84343 $w=2.4e-07 $l=1.38651e-07 $layer=LI1_cond $X=5.18 $Y=0.92
+ $X2=5.25 $Y2=0.812
r191 40 41 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=5.18 $Y=0.92
+ $X2=5.18 $Y2=1.95
r192 37 52 3.84343 $w=2.4e-07 $l=1.07e-07 $layer=LI1_cond $X=5.25 $Y=0.705
+ $X2=5.25 $Y2=0.812
r193 37 39 7.80687 $w=3.08e-07 $l=2.1e-07 $layer=LI1_cond $X=5.25 $Y=0.705
+ $X2=5.25 $Y2=0.495
r194 36 44 7.59919 $w=1.7e-07 $l=1.92873e-07 $layer=LI1_cond $X=5.25 $Y=0.425
+ $X2=5.405 $Y2=0.34
r195 36 39 2.60229 $w=3.08e-07 $l=7e-08 $layer=LI1_cond $X=5.25 $Y=0.425
+ $X2=5.25 $Y2=0.495
r196 34 52 2.60907 $w=1.7e-07 $l=1.65635e-07 $layer=LI1_cond $X=5.095 $Y=0.79
+ $X2=5.25 $Y2=0.812
r197 34 35 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=5.095 $Y=0.79
+ $X2=4.385 $Y2=0.79
r198 32 58 46.8028 $w=4.45e-07 $l=1.65e-07 $layer=POLY_cond $X=4.162 $Y=0.375
+ $X2=4.162 $Y2=0.54
r199 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.22
+ $Y=0.375 $X2=4.22 $Y2=0.375
r200 29 35 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.22 $Y=0.705
+ $X2=4.385 $Y2=0.79
r201 29 31 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=4.22 $Y=0.705
+ $X2=4.22 $Y2=0.375
r202 25 27 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=4.09 $Y=1.735
+ $X2=4.09 $Y2=2.23
r203 24 58 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=4.015 $Y=0.97
+ $X2=4.015 $Y2=0.54
r204 22 25 87.4216 $w=2.04e-07 $l=4.05771e-07 $layer=POLY_cond $X=4.015 $Y=1.365
+ $X2=4.09 $Y2=1.735
r205 22 24 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=4.015 $Y=1.365
+ $X2=4.015 $Y2=0.97
r206 19 32 21.2463 $w=4.45e-07 $l=1.7e-07 $layer=POLY_cond $X=4.162 $Y=0.205
+ $X2=4.162 $Y2=0.375
r207 19 20 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=3.94 $Y=0.205
+ $X2=3.11 $Y2=0.205
r208 18 28 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.035 $Y=0.89
+ $X2=3.035 $Y2=1.285
r209 15 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.035 $Y=0.28
+ $X2=3.11 $Y2=0.205
r210 15 18 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.035 $Y=0.28
+ $X2=3.035 $Y2=0.89
r211 12 14 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=3.02 $Y=1.735
+ $X2=3.02 $Y2=2.23
r212 11 12 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.02 $Y=1.645
+ $X2=3.02 $Y2=1.735
r213 10 28 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.02 $Y=1.375
+ $X2=3.02 $Y2=1.285
r214 10 11 104.952 $w=1.8e-07 $l=2.7e-07 $layer=POLY_cond $X=3.02 $Y=1.375
+ $X2=3.02 $Y2=1.645
r215 3 54 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=5.79
+ $Y=1.84 $X2=5.94 $Y2=2.115
r216 3 50 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=5.79
+ $Y=1.84 $X2=5.94 $Y2=2.815
r217 2 46 182 $w=1.7e-07 $l=4.92874e-07 $layer=licon1_NDIFF $count=1 $X=7.81
+ $Y=0.735 $X2=8.03 $Y2=0.34
r218 1 39 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=5.1
+ $Y=0.37 $X2=5.24 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LS__FAH_4%B 1 2 6 7 9 11 12 15 17 18 22 23 27 28 30 32
+ 35 37 38 42 43 47 48 49 58
c165 47 0 3.05047e-20 $X=4.8 $Y=2.065
c166 42 0 4.11294e-20 $X=4.8 $Y=1.385
c167 35 0 3.07659e-19 $X=3.64 $Y=1.66
c168 30 0 3.58366e-19 $X=5.715 $Y=1.765
r169 52 59 8.97022 $w=4.65e-07 $l=7.5e-08 $layer=POLY_cond $X=4.867 $Y=1.765
+ $X2=4.867 $Y2=1.69
r170 48 49 9.21977 $w=4.78e-07 $l=3.7e-07 $layer=LI1_cond $X=4.915 $Y=2.405
+ $X2=4.915 $Y2=2.775
r171 48 61 5.60012 $w=4.78e-07 $l=1.15e-07 $layer=LI1_cond $X=4.915 $Y=2.405
+ $X2=4.915 $Y2=2.29
r172 48 55 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.8
+ $Y=2.405 $X2=4.8 $Y2=2.405
r173 47 55 40.665 $w=4.65e-07 $l=3.4e-07 $layer=POLY_cond $X=4.867 $Y=2.065
+ $X2=4.867 $Y2=2.405
r174 47 52 35.8809 $w=4.65e-07 $l=3e-07 $layer=POLY_cond $X=4.867 $Y=2.065
+ $X2=4.867 $Y2=1.765
r175 46 61 10.372 $w=2.48e-07 $l=2.25e-07 $layer=LI1_cond $X=4.8 $Y=2.065
+ $X2=4.8 $Y2=2.29
r176 46 47 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=4.8
+ $Y=2.065 $X2=4.8 $Y2=2.065
r177 43 59 36.4789 $w=4.65e-07 $l=3.05e-07 $layer=POLY_cond $X=4.867 $Y=1.385
+ $X2=4.867 $Y2=1.69
r178 43 58 47.3569 $w=4.65e-07 $l=1.65e-07 $layer=POLY_cond $X=4.867 $Y=1.385
+ $X2=4.867 $Y2=1.22
r179 42 46 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=4.8 $Y=1.385
+ $X2=4.8 $Y2=2.065
r180 42 43 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=4.8
+ $Y=1.385 $X2=4.8 $Y2=1.385
r181 38 55 32.6516 $w=4.65e-07 $l=2.73e-07 $layer=POLY_cond $X=4.867 $Y=2.678
+ $X2=4.867 $Y2=2.405
r182 33 35 48.7128 $w=1.5e-07 $l=9.5e-08 $layer=POLY_cond $X=3.545 $Y=1.66
+ $X2=3.64 $Y2=1.66
r183 30 32 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.715 $Y=1.765
+ $X2=5.715 $Y2=2.4
r184 29 59 29.5843 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=5.1 $Y=1.69
+ $X2=4.867 $Y2=1.69
r185 28 30 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.64 $Y=1.69
+ $X2=5.715 $Y2=1.765
r186 28 29 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=5.64 $Y=1.69
+ $X2=5.1 $Y2=1.69
r187 27 58 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.025 $Y=0.74
+ $X2=5.025 $Y2=1.22
r188 24 37 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.73 $Y=3.095
+ $X2=3.64 $Y2=3.095
r189 23 38 49.4222 $w=4.65e-07 $l=5.20224e-07 $layer=POLY_cond $X=4.635 $Y=3.095
+ $X2=4.867 $Y2=2.678
r190 23 24 464.053 $w=1.5e-07 $l=9.05e-07 $layer=POLY_cond $X=4.635 $Y=3.095
+ $X2=3.73 $Y2=3.095
r191 20 22 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=3.64 $Y=2.725
+ $X2=3.64 $Y2=2.23
r192 19 35 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.64 $Y=1.735
+ $X2=3.64 $Y2=1.66
r193 19 22 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=3.64 $Y=1.735
+ $X2=3.64 $Y2=2.23
r194 18 37 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=3.64 $Y=3.02
+ $X2=3.64 $Y2=3.095
r195 17 20 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.64 $Y=2.815
+ $X2=3.64 $Y2=2.725
r196 17 18 79.6855 $w=1.8e-07 $l=2.05e-07 $layer=POLY_cond $X=3.64 $Y=2.815
+ $X2=3.64 $Y2=3.02
r197 13 33 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.545 $Y=1.585
+ $X2=3.545 $Y2=1.66
r198 13 15 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=3.545 $Y=1.585
+ $X2=3.545 $Y2=0.97
r199 11 37 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.55 $Y=3.095
+ $X2=3.64 $Y2=3.095
r200 11 12 458.926 $w=1.5e-07 $l=8.95e-07 $layer=POLY_cond $X=3.55 $Y=3.095
+ $X2=2.655 $Y2=3.095
r201 7 9 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.605 $Y=1.45
+ $X2=2.605 $Y2=0.89
r202 4 6 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.565 $Y=2.725
+ $X2=2.565 $Y2=2.23
r203 3 7 71.1762 $w=1.93e-07 $l=3.04344e-07 $layer=POLY_cond $X=2.565 $Y=1.735
+ $X2=2.605 $Y2=1.45
r204 3 6 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.565 $Y=1.735
+ $X2=2.565 $Y2=2.23
r205 2 12 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=2.565 $Y=3.02
+ $X2=2.655 $Y2=3.095
r206 1 4 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.565 $Y=2.815
+ $X2=2.565 $Y2=2.725
r207 1 2 79.6855 $w=1.8e-07 $l=2.05e-07 $layer=POLY_cond $X=2.565 $Y=2.815
+ $X2=2.565 $Y2=3.02
.ends

.subckt PM_SKY130_FD_SC_LS__FAH_4%A_528_362# 1 2 7 10 11 12 13 16 17 19 20 21 22
+ 24 29 30 35 39 41 46 47 49 50 51 52 55 59 61 62
c224 62 0 2.03891e-19 $X=5.52 $Y=1.665
c225 59 0 1.58586e-19 $X=4.08 $Y=1.665
c226 41 0 1.84628e-19 $X=3.885 $Y=1.657
c227 30 0 9.38777e-20 $X=6.275 $Y=1.3
c228 17 0 3.0708e-19 $X=6.315 $Y=1.225
c229 13 0 7.42391e-20 $X=6.25 $Y=1.82
c230 12 0 4.0679e-20 $X=6.25 $Y=3.075
r231 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=1.665
+ $X2=5.52 $Y2=1.665
r232 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=1.665
+ $X2=4.08 $Y2=1.665
r233 55 72 14.4306 $w=2.28e-07 $l=2.88e-07 $layer=LI1_cond $X=3.12 $Y=1.665
+ $X2=2.832 $Y2=1.665
r234 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=1.665
+ $X2=3.12 $Y2=1.665
r235 52 58 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.225 $Y=1.665
+ $X2=4.08 $Y2=1.665
r236 51 61 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.375 $Y=1.665
+ $X2=5.52 $Y2=1.665
r237 51 52 1.42326 $w=1.4e-07 $l=1.15e-06 $layer=MET1_cond $X=5.375 $Y=1.665
+ $X2=4.225 $Y2=1.665
r238 50 54 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.265 $Y=1.665
+ $X2=3.12 $Y2=1.665
r239 49 58 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.935 $Y=1.665
+ $X2=4.08 $Y2=1.665
r240 49 50 0.829206 $w=1.4e-07 $l=6.7e-07 $layer=MET1_cond $X=3.935 $Y=1.665
+ $X2=3.265 $Y2=1.665
r241 47 66 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.64 $Y=1.21 $X2=5.64
+ $Y2=1.3
r242 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.64
+ $Y=1.21 $X2=5.64 $Y2=1.21
r243 43 62 16.0818 $w=1.98e-07 $l=2.9e-07 $layer=LI1_cond $X=5.535 $Y=1.375
+ $X2=5.535 $Y2=1.665
r244 42 46 4.24584 $w=2.83e-07 $l=1.05e-07 $layer=LI1_cond $X=5.535 $Y=1.232
+ $X2=5.64 $Y2=1.232
r245 42 43 2.81168 $w=2e-07 $l=1.43e-07 $layer=LI1_cond $X=5.535 $Y=1.232
+ $X2=5.535 $Y2=1.375
r246 41 59 10.4524 $w=2.13e-07 $l=1.95e-07 $layer=LI1_cond $X=3.885 $Y=1.657
+ $X2=4.08 $Y2=1.657
r247 37 41 6.93832 $w=2.15e-07 $l=1.43332e-07 $layer=LI1_cond $X=3.8 $Y=1.55
+ $X2=3.885 $Y2=1.657
r248 37 39 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=3.8 $Y=1.55
+ $X2=3.8 $Y2=0.795
r249 33 72 0.103554 $w=2.55e-07 $l=1.15e-07 $layer=LI1_cond $X=2.832 $Y=1.78
+ $X2=2.832 $Y2=1.665
r250 33 35 7.90892 $w=2.53e-07 $l=1.75e-07 $layer=LI1_cond $X=2.832 $Y=1.78
+ $X2=2.832 $Y2=1.955
r251 27 29 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=7.485 $Y=3.03
+ $X2=7.485 $Y2=2.535
r252 26 32 13.2911 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=7.485 $Y=2.04
+ $X2=7.485 $Y2=1.855
r253 26 29 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=7.485 $Y=2.04
+ $X2=7.485 $Y2=2.535
r254 22 32 49.2255 $w=2.35e-07 $l=3.19374e-07 $layer=POLY_cond $X=7.245 $Y=1.67
+ $X2=7.485 $Y2=1.855
r255 22 24 371.755 $w=1.5e-07 $l=7.25e-07 $layer=POLY_cond $X=7.245 $Y=1.67
+ $X2=7.245 $Y2=0.945
r256 20 27 26.9307 $w=1.5e-07 $l=1.58745e-07 $layer=POLY_cond $X=7.395 $Y=3.15
+ $X2=7.485 $Y2=3.03
r257 20 21 540.968 $w=1.5e-07 $l=1.055e-06 $layer=POLY_cond $X=7.395 $Y=3.15
+ $X2=6.34 $Y2=3.15
r258 17 30 18.8402 $w=1.65e-07 $l=9.28709e-08 $layer=POLY_cond $X=6.315 $Y=1.225
+ $X2=6.275 $Y2=1.3
r259 17 19 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=6.315 $Y=1.225
+ $X2=6.315 $Y2=0.83
r260 14 16 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=6.25 $Y=2.81
+ $X2=6.25 $Y2=2.315
r261 13 16 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=6.25 $Y=1.82
+ $X2=6.25 $Y2=2.315
r262 12 21 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=6.25 $Y=3.075
+ $X2=6.34 $Y2=3.15
r263 11 14 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.25 $Y=2.9 $X2=6.25
+ $Y2=2.81
r264 11 12 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=6.25 $Y=2.9
+ $X2=6.25 $Y2=3.075
r265 10 13 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.25 $Y=1.73 $X2=6.25
+ $Y2=1.82
r266 9 30 18.8402 $w=1.65e-07 $l=8.66025e-08 $layer=POLY_cond $X=6.25 $Y=1.375
+ $X2=6.275 $Y2=1.3
r267 9 10 137.992 $w=1.8e-07 $l=3.55e-07 $layer=POLY_cond $X=6.25 $Y=1.375
+ $X2=6.25 $Y2=1.73
r268 8 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.805 $Y=1.3
+ $X2=5.64 $Y2=1.3
r269 7 30 6.66866 $w=1.5e-07 $l=1.15e-07 $layer=POLY_cond $X=6.16 $Y=1.3
+ $X2=6.275 $Y2=1.3
r270 7 8 182.032 $w=1.5e-07 $l=3.55e-07 $layer=POLY_cond $X=6.16 $Y=1.3
+ $X2=5.805 $Y2=1.3
r271 2 35 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.64
+ $Y=1.81 $X2=2.79 $Y2=1.955
r272 1 39 91 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_NDIFF $count=2 $X=3.62
+ $Y=0.65 $X2=3.8 $Y2=0.795
.ends

.subckt PM_SKY130_FD_SC_LS__FAH_4%A_536_114# 1 2 10 11 13 14 15 19 21 22 23 24
+ 26 29 33 35 36 38 39 40 41 47 52 55
c201 52 0 4.26248e-20 $X=6.795 $Y=1.57
c202 41 0 2.42154e-19 $X=3.745 $Y=2.035
c203 40 0 2.62373e-19 $X=6.815 $Y=2.035
c204 38 0 1.73206e-19 $X=3.46 $Y=1.935
c205 29 0 1.35123e-19 $X=7.89 $Y=1.525
c206 22 0 5.50318e-20 $X=8.36 $Y=1.965
r207 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.795
+ $Y=1.57 $X2=6.795 $Y2=1.57
r208 48 52 12.7592 $w=4.18e-07 $l=4.65e-07 $layer=LI1_cond $X=6.865 $Y=2.035
+ $X2=6.865 $Y2=1.57
r209 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=2.035
+ $X2=6.96 $Y2=2.035
r210 44 55 15.887 $w=1.83e-07 $l=2.65e-07 $layer=LI1_cond $X=3.6 $Y=2.027
+ $X2=3.865 $Y2=2.027
r211 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=2.035
+ $X2=3.6 $Y2=2.035
r212 41 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.745 $Y=2.035
+ $X2=3.6 $Y2=2.035
r213 40 47 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.815 $Y=2.035
+ $X2=6.96 $Y2=2.035
r214 40 41 3.7995 $w=1.4e-07 $l=3.07e-06 $layer=MET1_cond $X=6.815 $Y=2.035
+ $X2=3.745 $Y2=2.035
r215 39 44 3.2973 $w=1.83e-07 $l=5.5e-08 $layer=LI1_cond $X=3.545 $Y=2.027
+ $X2=3.6 $Y2=2.027
r216 38 39 6.83233 $w=1.85e-07 $l=1.27609e-07 $layer=LI1_cond $X=3.46 $Y=1.935
+ $X2=3.545 $Y2=2.027
r217 37 38 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=3.46 $Y=1.38
+ $X2=3.46 $Y2=1.935
r218 35 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.375 $Y=1.295
+ $X2=3.46 $Y2=1.38
r219 35 36 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=3.375 $Y=1.295
+ $X2=2.985 $Y2=1.295
r220 31 36 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.82 $Y=1.21
+ $X2=2.985 $Y2=1.295
r221 31 33 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=2.82 $Y=1.21
+ $X2=2.82 $Y2=0.745
r222 27 29 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=7.735 $Y=1.525
+ $X2=7.89 $Y2=1.525
r223 24 26 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=8.435 $Y=2.04
+ $X2=8.435 $Y2=2.535
r224 22 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.36 $Y=1.965
+ $X2=8.435 $Y2=2.04
r225 22 23 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=8.36 $Y=1.965
+ $X2=7.965 $Y2=1.965
r226 21 23 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.89 $Y=1.89
+ $X2=7.965 $Y2=1.965
r227 20 29 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.89 $Y=1.6
+ $X2=7.89 $Y2=1.525
r228 20 21 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=7.89 $Y=1.6
+ $X2=7.89 $Y2=1.89
r229 17 27 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.735 $Y=1.45
+ $X2=7.735 $Y2=1.525
r230 17 19 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=7.735 $Y=1.45
+ $X2=7.735 $Y2=1.055
r231 16 19 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=7.735 $Y=0.255
+ $X2=7.735 $Y2=1.055
r232 14 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.66 $Y=0.18
+ $X2=7.735 $Y2=0.255
r233 14 15 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=7.66 $Y=0.18
+ $X2=6.89 $Y2=0.18
r234 11 51 52.2586 $w=2.99e-07 $l=2.73861e-07 $layer=POLY_cond $X=6.845 $Y=1.82
+ $X2=6.795 $Y2=1.57
r235 11 13 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=6.845 $Y=1.82
+ $X2=6.845 $Y2=2.315
r236 8 51 38.5562 $w=2.99e-07 $l=1.74714e-07 $layer=POLY_cond $X=6.815 $Y=1.405
+ $X2=6.795 $Y2=1.57
r237 8 10 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=6.815 $Y=1.405
+ $X2=6.815 $Y2=0.945
r238 7 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.815 $Y=0.255
+ $X2=6.89 $Y2=0.18
r239 7 10 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.815 $Y=0.255
+ $X2=6.815 $Y2=0.945
r240 2 55 600 $w=1.7e-07 $l=2.80134e-07 $layer=licon1_PDIFF $count=1 $X=3.715
+ $Y=1.81 $X2=3.865 $Y2=2.025
r241 1 33 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=2.68
+ $Y=0.57 $X2=2.82 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_LS__FAH_4%A_1378_125# 1 2 3 4 13 15 16 18 20 21 22 24 26
+ 28 30 31 32 36 38 39 41 43 46 51 52 54 58 61 62 64 65 66 67 72 73
c225 61 0 1.37274e-19 $X=7.03 $Y=1.11
c226 58 0 1.68117e-19 $X=6.4 $Y=2.065
c227 41 0 1.35123e-19 $X=8.37 $Y=1.485
c228 38 0 1.70833e-19 $X=7.875 $Y=1.565
c229 26 0 1.69806e-19 $X=6.4 $Y=1.98
c230 24 0 4.0679e-20 $X=6.28 $Y=2.905
c231 21 0 2.61071e-20 $X=8.88 $Y=1.485
r232 72 73 6.54147 $w=4.18e-07 $l=8.5e-08 $layer=LI1_cond $X=12.505 $Y=2.035
+ $X2=12.505 $Y2=1.95
r233 67 69 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=8.63 $Y=2.695
+ $X2=8.63 $Y2=2.99
r234 61 62 9.43135 $w=1.98e-07 $l=1.65e-07 $layer=LI1_cond $X=7.03 $Y=1.115
+ $X2=6.865 $Y2=1.115
r235 56 58 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=6.28 $Y=2.065
+ $X2=6.4 $Y2=2.065
r236 52 54 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=12.465 $Y=1.095
+ $X2=12.69 $Y2=1.095
r237 51 75 2.84834 $w=4.2e-07 $l=1.25e-07 $layer=LI1_cond $X=12.505 $Y=2.61
+ $X2=12.505 $Y2=2.735
r238 50 72 3.42989 $w=4.18e-07 $l=1.25e-07 $layer=LI1_cond $X=12.505 $Y=2.16
+ $X2=12.505 $Y2=2.035
r239 50 51 12.3476 $w=4.18e-07 $l=4.5e-07 $layer=LI1_cond $X=12.505 $Y=2.16
+ $X2=12.505 $Y2=2.61
r240 48 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=12.38 $Y=1.18
+ $X2=12.465 $Y2=1.095
r241 48 73 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=12.38 $Y=1.18
+ $X2=12.38 $Y2=1.95
r242 47 67 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.715 $Y=2.695
+ $X2=8.63 $Y2=2.695
r243 46 75 5.69669 $w=1.7e-07 $l=2.29129e-07 $layer=LI1_cond $X=12.295 $Y=2.695
+ $X2=12.505 $Y2=2.735
r244 46 47 233.561 $w=1.68e-07 $l=3.58e-06 $layer=LI1_cond $X=12.295 $Y=2.695
+ $X2=8.715 $Y2=2.695
r245 43 44 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.71
+ $Y=1.485 $X2=8.71 $Y2=1.485
r246 41 66 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=8.37 $Y=1.485
+ $X2=8.205 $Y2=1.485
r247 41 43 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=8.37 $Y=1.485
+ $X2=8.71 $Y2=1.485
r248 40 65 3.58051 $w=2.6e-07 $l=1.25499e-07 $layer=LI1_cond $X=7.875 $Y=2.99
+ $X2=7.79 $Y2=2.9
r249 39 69 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.545 $Y=2.99
+ $X2=8.63 $Y2=2.99
r250 39 40 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.545 $Y=2.99
+ $X2=7.875 $Y2=2.99
r251 38 66 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=7.875 $Y=1.565
+ $X2=8.205 $Y2=1.565
r252 36 65 2.90867 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=7.79 $Y=2.725
+ $X2=7.79 $Y2=2.9
r253 35 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.79 $Y=1.65
+ $X2=7.875 $Y2=1.565
r254 35 36 70.1337 $w=1.68e-07 $l=1.075e-06 $layer=LI1_cond $X=7.79 $Y=1.65
+ $X2=7.79 $Y2=2.725
r255 32 64 8.81775 $w=3.48e-07 $l=1.75e-07 $layer=LI1_cond $X=7.165 $Y=2.9
+ $X2=6.99 $Y2=2.9
r256 32 34 1.31708 $w=3.48e-07 $l=4e-08 $layer=LI1_cond $X=7.165 $Y=2.9
+ $X2=7.205 $Y2=2.9
r257 31 65 3.58051 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=7.705 $Y=2.9
+ $X2=7.79 $Y2=2.9
r258 31 34 16.4635 $w=3.48e-07 $l=5e-07 $layer=LI1_cond $X=7.705 $Y=2.9
+ $X2=7.205 $Y2=2.9
r259 30 62 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=6.485 $Y=1.13
+ $X2=6.865 $Y2=1.13
r260 28 64 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=6.365 $Y=2.99
+ $X2=6.99 $Y2=2.99
r261 26 58 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.4 $Y=1.98 $X2=6.4
+ $Y2=2.065
r262 25 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.4 $Y=1.215
+ $X2=6.485 $Y2=1.13
r263 25 26 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=6.4 $Y=1.215
+ $X2=6.4 $Y2=1.98
r264 24 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.28 $Y=2.905
+ $X2=6.365 $Y2=2.99
r265 23 56 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.28 $Y=2.15
+ $X2=6.28 $Y2=2.065
r266 23 24 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=6.28 $Y=2.15
+ $X2=6.28 $Y2=2.905
r267 21 44 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=8.88 $Y=1.485
+ $X2=8.71 $Y2=1.485
r268 21 22 13.5877 $w=2.4e-07 $l=1.15022e-07 $layer=POLY_cond $X=8.88 $Y=1.485
+ $X2=8.97 $Y2=1.542
r269 18 20 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=9.425 $Y=1.32
+ $X2=9.425 $Y2=0.92
r270 17 22 13.5877 $w=2.4e-07 $l=1.86652e-07 $layer=POLY_cond $X=9.06 $Y=1.395
+ $X2=8.97 $Y2=1.542
r271 16 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.35 $Y=1.395
+ $X2=9.425 $Y2=1.32
r272 16 17 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=9.35 $Y=1.395
+ $X2=9.06 $Y2=1.395
r273 13 22 12.1617 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=8.97 $Y=1.765
+ $X2=8.97 $Y2=1.542
r274 13 15 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=8.97 $Y=1.765
+ $X2=8.97 $Y2=2.34
r275 4 75 400 $w=1.7e-07 $l=9.44722e-07 $layer=licon1_PDIFF $count=1 $X=12.405
+ $Y=1.84 $X2=12.55 $Y2=2.715
r276 4 72 400 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=1 $X=12.405
+ $Y=1.84 $X2=12.55 $Y2=2.035
r277 3 34 600 $w=1.7e-07 $l=1.04785e-06 $layer=licon1_PDIFF $count=1 $X=6.92
+ $Y=1.895 $X2=7.205 $Y2=2.81
r278 2 54 182 $w=1.7e-07 $l=5.6285e-07 $layer=licon1_NDIFF $count=1 $X=12.545
+ $Y=0.6 $X2=12.69 $Y2=1.095
r279 1 61 182 $w=1.7e-07 $l=5.50568e-07 $layer=licon1_NDIFF $count=1 $X=6.89
+ $Y=0.625 $X2=7.03 $Y2=1.11
.ends

.subckt PM_SKY130_FD_SC_LS__FAH_4%A_1265_379# 1 2 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 27 28 30 31 34 35 38 39 40 42 43 44 46 49 52 57 73
c177 31 0 1.8874e-19 $X=7.365 $Y=2.405
r178 73 74 57.7326 $w=3.59e-07 $l=4.3e-07 $layer=POLY_cond $X=11.405 $Y=1.557
+ $X2=11.835 $Y2=1.557
r179 72 73 7.3844 $w=3.59e-07 $l=5.5e-08 $layer=POLY_cond $X=11.35 $Y=1.557
+ $X2=11.405 $Y2=1.557
r180 71 72 60.4178 $w=3.59e-07 $l=4.5e-07 $layer=POLY_cond $X=10.9 $Y=1.557
+ $X2=11.35 $Y2=1.557
r181 70 71 6.04178 $w=3.59e-07 $l=4.5e-08 $layer=POLY_cond $X=10.855 $Y=1.557
+ $X2=10.9 $Y2=1.557
r182 67 68 19.468 $w=3.59e-07 $l=1.45e-07 $layer=POLY_cond $X=10.28 $Y=1.557
+ $X2=10.425 $Y2=1.557
r183 64 67 50.3482 $w=3.59e-07 $l=3.75e-07 $layer=POLY_cond $X=9.905 $Y=1.557
+ $X2=10.28 $Y2=1.557
r184 64 65 10.0696 $w=3.59e-07 $l=7.5e-08 $layer=POLY_cond $X=9.905 $Y=1.557
+ $X2=9.83 $Y2=1.557
r185 63 64 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=9.905
+ $Y=1.515 $X2=9.905 $Y2=1.515
r186 60 61 8.82039 $w=3.18e-07 $l=1.75e-07 $layer=LI1_cond $X=7.525 $Y=1.11
+ $X2=7.525 $Y2=1.285
r187 57 60 3.24125 $w=3.18e-07 $l=9e-08 $layer=LI1_cond $X=7.525 $Y=1.02
+ $X2=7.525 $Y2=1.11
r188 52 55 5.53173 $w=2.48e-07 $l=1.2e-07 $layer=LI1_cond $X=6.66 $Y=2.405
+ $X2=6.66 $Y2=2.525
r189 50 70 36.2507 $w=3.59e-07 $l=2.7e-07 $layer=POLY_cond $X=10.585 $Y=1.557
+ $X2=10.855 $Y2=1.557
r190 50 68 21.4819 $w=3.59e-07 $l=1.6e-07 $layer=POLY_cond $X=10.585 $Y=1.557
+ $X2=10.425 $Y2=1.557
r191 49 50 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=10.585
+ $Y=1.515 $X2=10.585 $Y2=1.515
r192 47 63 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.95 $Y=1.515
+ $X2=9.865 $Y2=1.515
r193 47 49 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=9.95 $Y=1.515
+ $X2=10.585 $Y2=1.515
r194 46 63 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.865 $Y=1.35
+ $X2=9.865 $Y2=1.515
r195 45 46 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=9.865 $Y=1.18
+ $X2=9.865 $Y2=1.35
r196 43 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.78 $Y=1.095
+ $X2=9.865 $Y2=1.18
r197 43 44 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=9.78 $Y=1.095
+ $X2=9.555 $Y2=1.095
r198 42 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.47 $Y=1.01
+ $X2=9.555 $Y2=1.095
r199 41 42 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=9.47 $Y=0.765
+ $X2=9.47 $Y2=1.01
r200 39 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.385 $Y=0.68
+ $X2=9.47 $Y2=0.765
r201 39 40 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=9.385 $Y=0.68
+ $X2=8.875 $Y2=0.68
r202 37 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.79 $Y=0.765
+ $X2=8.875 $Y2=0.68
r203 37 38 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=8.79 $Y=0.765
+ $X2=8.79 $Y2=0.935
r204 36 57 4.44149 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=7.685 $Y=1.02
+ $X2=7.525 $Y2=1.02
r205 35 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.705 $Y=1.02
+ $X2=8.79 $Y2=0.935
r206 35 36 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=8.705 $Y=1.02
+ $X2=7.685 $Y2=1.02
r207 34 61 67.5241 $w=1.68e-07 $l=1.035e-06 $layer=LI1_cond $X=7.45 $Y=2.32
+ $X2=7.45 $Y2=1.285
r208 32 52 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.785 $Y=2.405
+ $X2=6.66 $Y2=2.405
r209 31 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.365 $Y=2.405
+ $X2=7.45 $Y2=2.32
r210 31 32 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=7.365 $Y=2.405
+ $X2=6.785 $Y2=2.405
r211 28 74 23.2387 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=11.835 $Y=1.35
+ $X2=11.835 $Y2=1.557
r212 28 30 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=11.835 $Y=1.35
+ $X2=11.835 $Y2=0.87
r213 25 73 23.2387 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=11.405 $Y=1.35
+ $X2=11.405 $Y2=1.557
r214 25 27 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=11.405 $Y=1.35
+ $X2=11.405 $Y2=0.87
r215 22 72 23.2387 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=11.35 $Y=1.765
+ $X2=11.35 $Y2=1.557
r216 22 24 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=11.35 $Y=1.765
+ $X2=11.35 $Y2=2.4
r217 19 71 23.2387 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=10.9 $Y=1.765
+ $X2=10.9 $Y2=1.557
r218 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=10.9 $Y=1.765
+ $X2=10.9 $Y2=2.4
r219 16 70 23.2387 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=10.855 $Y=1.35
+ $X2=10.855 $Y2=1.557
r220 16 18 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=10.855 $Y=1.35
+ $X2=10.855 $Y2=0.87
r221 13 68 23.2387 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=10.425 $Y=1.35
+ $X2=10.425 $Y2=1.557
r222 13 15 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=10.425 $Y=1.35
+ $X2=10.425 $Y2=0.87
r223 10 67 23.2387 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=10.28 $Y=1.765
+ $X2=10.28 $Y2=1.557
r224 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=10.28 $Y=1.765
+ $X2=10.28 $Y2=2.4
r225 7 65 23.2387 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=9.83 $Y=1.765
+ $X2=9.83 $Y2=1.557
r226 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=9.83 $Y=1.765
+ $X2=9.83 $Y2=2.4
r227 2 55 600 $w=1.7e-07 $l=7.63381e-07 $layer=licon1_PDIFF $count=1 $X=6.325
+ $Y=1.895 $X2=6.62 $Y2=2.525
r228 1 60 182 $w=1.7e-07 $l=5.7639e-07 $layer=licon1_NDIFF $count=1 $X=7.32
+ $Y=0.625 $X2=7.52 $Y2=1.11
.ends

.subckt PM_SKY130_FD_SC_LS__FAH_4%CI 1 3 4 6 7 11
r35 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.815
+ $Y=1.515 $X2=12.815 $Y2=1.515
r36 7 11 5.01062 $w=3.43e-07 $l=1.5e-07 $layer=LI1_cond $X=12.807 $Y=1.665
+ $X2=12.807 $Y2=1.515
r37 4 10 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=12.905 $Y=1.35
+ $X2=12.815 $Y2=1.515
r38 4 6 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=12.905 $Y=1.35
+ $X2=12.905 $Y2=0.92
r39 1 10 52.2586 $w=2.99e-07 $l=2.69258e-07 $layer=POLY_cond $X=12.775 $Y=1.765
+ $X2=12.815 $Y2=1.515
r40 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=12.775 $Y=1.765
+ $X2=12.775 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_LS__FAH_4%A_1278_102# 1 2 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 27 28 30 31 34 35 37 38 40 41 42 44 45 48 49 54 60 62 66 75
c218 62 0 2.61071e-20 $X=8.21 $Y=2.26
c219 19 0 6.40318e-20 $X=14.35 $Y=1.765
c220 16 0 1.44963e-19 $X=13.935 $Y=1.35
r221 75 76 1.97003 $w=3.67e-07 $l=1.5e-08 $layer=POLY_cond $X=14.795 $Y=1.557
+ $X2=14.81 $Y2=1.557
r222 74 75 56.4741 $w=3.67e-07 $l=4.3e-07 $layer=POLY_cond $X=14.365 $Y=1.557
+ $X2=14.795 $Y2=1.557
r223 73 74 1.97003 $w=3.67e-07 $l=1.5e-08 $layer=POLY_cond $X=14.35 $Y=1.557
+ $X2=14.365 $Y2=1.557
r224 70 71 16.4169 $w=3.67e-07 $l=1.25e-07 $layer=POLY_cond $X=13.81 $Y=1.557
+ $X2=13.935 $Y2=1.557
r225 69 70 40.0572 $w=3.67e-07 $l=3.05e-07 $layer=POLY_cond $X=13.505 $Y=1.557
+ $X2=13.81 $Y2=1.557
r226 62 64 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=8.21 $Y=2.26
+ $X2=8.21 $Y2=2.355
r227 58 60 8.79328 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=6.54 $Y=0.72
+ $X2=6.705 $Y2=0.72
r228 55 73 24.9537 $w=3.67e-07 $l=1.9e-07 $layer=POLY_cond $X=14.16 $Y=1.557
+ $X2=14.35 $Y2=1.557
r229 55 71 29.5504 $w=3.67e-07 $l=2.25e-07 $layer=POLY_cond $X=14.16 $Y=1.557
+ $X2=13.935 $Y2=1.557
r230 54 55 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=14.16
+ $Y=1.515 $X2=14.16 $Y2=1.515
r231 52 69 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=13.48 $Y=1.557
+ $X2=13.505 $Y2=1.557
r232 52 67 15.7602 $w=3.67e-07 $l=1.2e-07 $layer=POLY_cond $X=13.48 $Y=1.557
+ $X2=13.36 $Y2=1.557
r233 51 54 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=13.48 $Y=1.515
+ $X2=14.16 $Y2=1.515
r234 51 52 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=13.48
+ $Y=1.515 $X2=13.48 $Y2=1.515
r235 49 51 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=13.385 $Y=1.515
+ $X2=13.48 $Y2=1.515
r236 48 49 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=13.3 $Y=1.35
+ $X2=13.385 $Y2=1.515
r237 47 48 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=13.3 $Y=0.84
+ $X2=13.3 $Y2=1.35
r238 46 66 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.125 $Y=0.755
+ $X2=12.04 $Y2=0.755
r239 45 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=13.215 $Y=0.755
+ $X2=13.3 $Y2=0.84
r240 45 46 71.1123 $w=1.68e-07 $l=1.09e-06 $layer=LI1_cond $X=13.215 $Y=0.755
+ $X2=12.125 $Y2=0.755
r241 43 66 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.04 $Y=0.84
+ $X2=12.04 $Y2=0.755
r242 43 44 93.2941 $w=1.68e-07 $l=1.43e-06 $layer=LI1_cond $X=12.04 $Y=0.84
+ $X2=12.04 $Y2=2.27
r243 41 66 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.955 $Y=0.755
+ $X2=12.04 $Y2=0.755
r244 41 42 134.396 $w=1.68e-07 $l=2.06e-06 $layer=LI1_cond $X=11.955 $Y=0.755
+ $X2=9.895 $Y2=0.755
r245 40 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.81 $Y=0.67
+ $X2=9.895 $Y2=0.755
r246 39 40 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=9.81 $Y=0.425
+ $X2=9.81 $Y2=0.67
r247 37 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.725 $Y=0.34
+ $X2=9.81 $Y2=0.425
r248 37 38 77.6364 $w=1.68e-07 $l=1.19e-06 $layer=LI1_cond $X=9.725 $Y=0.34
+ $X2=8.535 $Y2=0.34
r249 36 64 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.375 $Y=2.355
+ $X2=8.21 $Y2=2.355
r250 35 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.955 $Y=2.355
+ $X2=12.04 $Y2=2.27
r251 35 36 233.561 $w=1.68e-07 $l=3.58e-06 $layer=LI1_cond $X=11.955 $Y=2.355
+ $X2=8.375 $Y2=2.355
r252 33 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.45 $Y=0.425
+ $X2=8.535 $Y2=0.34
r253 33 34 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=8.45 $Y=0.425
+ $X2=8.45 $Y2=0.595
r254 31 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.365 $Y=0.68
+ $X2=8.45 $Y2=0.595
r255 31 60 108.299 $w=1.68e-07 $l=1.66e-06 $layer=LI1_cond $X=8.365 $Y=0.68
+ $X2=6.705 $Y2=0.68
r256 28 76 23.77 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=14.81 $Y=1.765
+ $X2=14.81 $Y2=1.557
r257 28 30 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=14.81 $Y=1.765
+ $X2=14.81 $Y2=2.4
r258 25 75 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=14.795 $Y=1.35
+ $X2=14.795 $Y2=1.557
r259 25 27 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=14.795 $Y=1.35
+ $X2=14.795 $Y2=0.87
r260 22 74 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=14.365 $Y=1.35
+ $X2=14.365 $Y2=1.557
r261 22 24 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=14.365 $Y=1.35
+ $X2=14.365 $Y2=0.87
r262 19 73 23.77 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=14.35 $Y=1.765
+ $X2=14.35 $Y2=1.557
r263 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=14.35 $Y=1.765
+ $X2=14.35 $Y2=2.4
r264 16 71 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=13.935 $Y=1.35
+ $X2=13.935 $Y2=1.557
r265 16 18 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=13.935 $Y=1.35
+ $X2=13.935 $Y2=0.87
r266 13 70 23.77 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=13.81 $Y=1.765
+ $X2=13.81 $Y2=1.557
r267 13 15 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=13.81 $Y=1.765
+ $X2=13.81 $Y2=2.4
r268 10 69 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=13.505 $Y=1.35
+ $X2=13.505 $Y2=1.557
r269 10 12 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=13.505 $Y=1.35
+ $X2=13.505 $Y2=0.87
r270 7 67 23.77 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=13.36 $Y=1.765
+ $X2=13.36 $Y2=1.557
r271 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=13.36 $Y=1.765
+ $X2=13.36 $Y2=2.4
r272 2 62 300 $w=1.7e-07 $l=7.18853e-07 $layer=licon1_PDIFF $count=2 $X=7.56
+ $Y=2.115 $X2=8.21 $Y2=2.26
r273 1 58 182 $w=1.7e-07 $l=2.33238e-07 $layer=licon1_NDIFF $count=1 $X=6.39
+ $Y=0.51 $X2=6.54 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_LS__FAH_4%VPWR 1 2 3 4 5 6 7 8 9 30 36 40 46 48 50 55 58
+ 62 63 64 66 71 76 104 108 114 117 124 129 132 136 139 141 145
r170 144 145 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.12 $Y=3.33
+ $X2=15.12 $Y2=3.33
r171 141 142 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.16 $Y=3.33
+ $X2=14.16 $Y2=3.33
r172 138 139 13.167 $w=4.63e-07 $l=3.15e-07 $layer=LI1_cond $X=11.81 $Y=3.182
+ $X2=12.125 $Y2=3.182
r173 134 138 1.28611 $w=4.63e-07 $l=5e-08 $layer=LI1_cond $X=11.76 $Y=3.182
+ $X2=11.81 $Y2=3.182
r174 134 136 11.8809 $w=4.63e-07 $l=2.65e-07 $layer=LI1_cond $X=11.76 $Y=3.182
+ $X2=11.495 $Y2=3.182
r175 134 135 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r176 131 132 12.3953 $w=4.63e-07 $l=2.85e-07 $layer=LI1_cond $X=9.4 $Y=3.182
+ $X2=9.685 $Y2=3.182
r177 127 131 1.02888 $w=4.63e-07 $l=4e-08 $layer=LI1_cond $X=9.36 $Y=3.182
+ $X2=9.4 $Y2=3.182
r178 127 129 11.3664 $w=4.63e-07 $l=2.45e-07 $layer=LI1_cond $X=9.36 $Y=3.182
+ $X2=9.115 $Y2=3.182
r179 127 128 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r180 124 125 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r181 120 121 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r182 117 120 9.32123 $w=3.38e-07 $l=2.75e-07 $layer=LI1_cond $X=1.745 $Y=3.055
+ $X2=1.745 $Y2=3.33
r183 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r184 112 145 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.64 $Y=3.33
+ $X2=15.12 $Y2=3.33
r185 112 142 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.64 $Y=3.33
+ $X2=14.16 $Y2=3.33
r186 111 112 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.64 $Y=3.33
+ $X2=14.64 $Y2=3.33
r187 109 141 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.25 $Y=3.33
+ $X2=14.085 $Y2=3.33
r188 109 111 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=14.25 $Y=3.33
+ $X2=14.64 $Y2=3.33
r189 108 144 3.9577 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=14.95 $Y=3.33
+ $X2=15.155 $Y2=3.33
r190 108 111 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=14.95 $Y=3.33
+ $X2=14.64 $Y2=3.33
r191 107 142 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=3.33
+ $X2=14.16 $Y2=3.33
r192 106 107 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.68 $Y=3.33
+ $X2=13.68 $Y2=3.33
r193 104 141 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.92 $Y=3.33
+ $X2=14.085 $Y2=3.33
r194 104 106 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=13.92 $Y=3.33
+ $X2=13.68 $Y2=3.33
r195 103 107 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=13.68 $Y2=3.33
r196 103 135 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=11.76 $Y2=3.33
r197 102 139 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=12.72 $Y=3.33
+ $X2=12.125 $Y2=3.33
r198 102 103 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r199 99 135 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=11.76 $Y2=3.33
r200 98 136 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=11.28 $Y=3.33
+ $X2=11.495 $Y2=3.33
r201 98 99 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r202 95 99 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=11.28 $Y2=3.33
r203 95 128 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=9.36 $Y2=3.33
r204 94 132 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=10.32 $Y=3.33
+ $X2=9.685 $Y2=3.33
r205 94 95 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r206 91 128 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=9.36 $Y2=3.33
r207 90 129 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=8.88 $Y=3.33
+ $X2=9.115 $Y2=3.33
r208 90 91 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r209 88 125 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=5.52 $Y2=3.33
r210 87 90 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=6 $Y=3.33 $X2=8.88
+ $Y2=3.33
r211 87 88 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=6 $Y=3.33
+ $X2=6 $Y2=3.33
r212 85 124 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.655 $Y=3.33
+ $X2=5.49 $Y2=3.33
r213 85 87 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=5.655 $Y=3.33 $X2=6
+ $Y2=3.33
r214 83 125 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r215 82 83 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r216 80 83 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=5.04 $Y2=3.33
r217 80 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r218 79 82 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=5.04 $Y2=3.33
r219 79 80 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r220 77 120 4.80115 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=1.915 $Y=3.33
+ $X2=1.745 $Y2=3.33
r221 77 79 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.915 $Y=3.33
+ $X2=2.16 $Y2=3.33
r222 76 124 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.325 $Y=3.33
+ $X2=5.49 $Y2=3.33
r223 76 82 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=5.325 $Y=3.33
+ $X2=5.04 $Y2=3.33
r224 75 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r225 75 115 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r226 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r227 72 114 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.815 $Y=3.33
+ $X2=0.69 $Y2=3.33
r228 72 74 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.815 $Y=3.33
+ $X2=1.2 $Y2=3.33
r229 71 120 4.80115 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=1.575 $Y=3.33
+ $X2=1.745 $Y2=3.33
r230 71 74 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.575 $Y=3.33
+ $X2=1.2 $Y2=3.33
r231 69 115 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r232 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r233 66 114 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.69 $Y2=3.33
r234 66 68 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.24 $Y2=3.33
r235 64 91 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=7.68 $Y=3.33
+ $X2=8.88 $Y2=3.33
r236 64 88 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=7.68 $Y=3.33
+ $X2=6 $Y2=3.33
r237 62 102 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=12.92 $Y=3.33
+ $X2=12.72 $Y2=3.33
r238 62 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.92 $Y=3.33
+ $X2=13.085 $Y2=3.33
r239 61 106 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=13.25 $Y=3.33
+ $X2=13.68 $Y2=3.33
r240 61 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.25 $Y=3.33
+ $X2=13.085 $Y2=3.33
r241 59 98 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=10.755 $Y=3.33
+ $X2=11.28 $Y2=3.33
r242 58 94 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=10.425 $Y=3.33
+ $X2=10.32 $Y2=3.33
r243 57 59 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.59 $Y=3.33
+ $X2=10.755 $Y2=3.33
r244 57 58 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.59 $Y=3.33
+ $X2=10.425 $Y2=3.33
r245 55 57 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=10.59 $Y=3.04
+ $X2=10.59 $Y2=3.33
r246 50 53 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=15.075 $Y=1.985
+ $X2=15.075 $Y2=2.815
r247 48 144 3.18546 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=15.075 $Y=3.245
+ $X2=15.155 $Y2=3.33
r248 48 53 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=15.075 $Y=3.245
+ $X2=15.075 $Y2=2.815
r249 44 141 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=14.085 $Y=3.245
+ $X2=14.085 $Y2=3.33
r250 44 46 31.081 $w=3.28e-07 $l=8.9e-07 $layer=LI1_cond $X=14.085 $Y=3.245
+ $X2=14.085 $Y2=2.355
r251 40 43 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=13.085 $Y=2.035
+ $X2=13.085 $Y2=2.815
r252 38 63 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.085 $Y=3.245
+ $X2=13.085 $Y2=3.33
r253 38 43 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=13.085 $Y=3.245
+ $X2=13.085 $Y2=2.815
r254 34 124 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.49 $Y=3.245
+ $X2=5.49 $Y2=3.33
r255 34 36 30.0334 $w=3.28e-07 $l=8.6e-07 $layer=LI1_cond $X=5.49 $Y=3.245
+ $X2=5.49 $Y2=2.385
r256 30 33 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=0.69 $Y=2.135
+ $X2=0.69 $Y2=2.815
r257 28 114 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=3.245
+ $X2=0.69 $Y2=3.33
r258 28 33 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.69 $Y=3.245
+ $X2=0.69 $Y2=2.815
r259 9 53 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=14.885
+ $Y=1.84 $X2=15.035 $Y2=2.815
r260 9 50 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=14.885
+ $Y=1.84 $X2=15.035 $Y2=1.985
r261 8 46 300 $w=1.7e-07 $l=6.06815e-07 $layer=licon1_PDIFF $count=2 $X=13.885
+ $Y=1.84 $X2=14.085 $Y2=2.355
r262 7 43 600 $w=1.7e-07 $l=1.08616e-06 $layer=licon1_PDIFF $count=1 $X=12.85
+ $Y=1.84 $X2=13.085 $Y2=2.815
r263 7 40 300 $w=1.7e-07 $l=3.17884e-07 $layer=licon1_PDIFF $count=2 $X=12.85
+ $Y=1.84 $X2=13.085 $Y2=2.035
r264 6 138 600 $w=1.7e-07 $l=1.37408e-06 $layer=licon1_PDIFF $count=1 $X=11.425
+ $Y=1.84 $X2=11.81 $Y2=3.035
r265 5 55 600 $w=1.7e-07 $l=1.31225e-06 $layer=licon1_PDIFF $count=1 $X=10.355
+ $Y=1.84 $X2=10.59 $Y2=3.04
r266 4 131 600 $w=1.7e-07 $l=1.36097e-06 $layer=licon1_PDIFF $count=1 $X=9.045
+ $Y=1.84 $X2=9.4 $Y2=3.035
r267 3 36 300 $w=1.7e-07 $l=6.13229e-07 $layer=licon1_PDIFF $count=2 $X=5.345
+ $Y=1.84 $X2=5.49 $Y2=2.385
r268 2 117 600 $w=1.7e-07 $l=1.31787e-06 $layer=licon1_PDIFF $count=1 $X=1.595
+ $Y=1.81 $X2=1.745 $Y2=3.055
r269 1 33 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.96 $X2=0.73 $Y2=2.815
r270 1 30 400 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.96 $X2=0.73 $Y2=2.135
.ends

.subckt PM_SKY130_FD_SC_LS__FAH_4%A_200_74# 1 2 3 4 15 17 19 21 22 23 26 28 29
+ 31 32 35 39 41 42
c115 19 0 5.85186e-20 $X=1.18 $Y=2.135
c116 17 0 1.1412e-19 $X=1.18 $Y=2.63
c117 15 0 1.40087e-19 $X=1.14 $Y=0.515
r118 42 45 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=3.33 $Y=2.715 $X2=3.33
+ $Y2=2.795
r119 39 40 8.26042 $w=1.92e-07 $l=1.3e-07 $layer=LI1_cond $X=1.92 $Y=0.895
+ $X2=2.05 $Y2=0.895
r120 33 35 18.1731 $w=2.58e-07 $l=4.1e-07 $layer=LI1_cond $X=3.285 $Y=0.425
+ $X2=3.285 $Y2=0.835
r121 31 33 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=3.155 $Y=0.34
+ $X2=3.285 $Y2=0.425
r122 31 32 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=3.155 $Y=0.34
+ $X2=2.135 $Y2=0.34
r123 30 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.005 $Y=2.715
+ $X2=1.92 $Y2=2.715
r124 29 42 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.165 $Y=2.715
+ $X2=3.33 $Y2=2.715
r125 29 30 75.6791 $w=1.68e-07 $l=1.16e-06 $layer=LI1_cond $X=3.165 $Y=2.715
+ $X2=2.005 $Y2=2.715
r126 28 40 1.44825 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.05 $Y=0.79
+ $X2=2.05 $Y2=0.895
r127 27 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.05 $Y=0.425
+ $X2=2.135 $Y2=0.34
r128 27 28 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.05 $Y=0.425
+ $X2=2.05 $Y2=0.79
r129 26 41 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.92 $Y=2.63
+ $X2=1.92 $Y2=2.715
r130 25 39 1.44825 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.92 $Y=1 $X2=1.92
+ $Y2=0.895
r131 25 26 106.342 $w=1.68e-07 $l=1.63e-06 $layer=LI1_cond $X=1.92 $Y=1 $X2=1.92
+ $Y2=2.63
r132 24 38 4.60552 $w=1.7e-07 $l=2.05122e-07 $layer=LI1_cond $X=1.345 $Y=2.715
+ $X2=1.18 $Y2=2.805
r133 23 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.835 $Y=2.715
+ $X2=1.92 $Y2=2.715
r134 23 24 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=1.835 $Y=2.715
+ $X2=1.345 $Y2=2.715
r135 21 39 5.05061 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.835 $Y=0.895
+ $X2=1.92 $Y2=0.895
r136 21 22 27.9913 $w=2.08e-07 $l=5.3e-07 $layer=LI1_cond $X=1.835 $Y=0.895
+ $X2=1.305 $Y2=0.895
r137 17 38 3.16065 $w=3.3e-07 $l=1.75e-07 $layer=LI1_cond $X=1.18 $Y=2.63
+ $X2=1.18 $Y2=2.805
r138 17 19 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=1.18 $Y=2.63
+ $X2=1.18 $Y2=2.135
r139 13 22 7.26367 $w=2.1e-07 $l=2.11069e-07 $layer=LI1_cond $X=1.14 $Y=0.79
+ $X2=1.305 $Y2=0.895
r140 13 15 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.14 $Y=0.79
+ $X2=1.14 $Y2=0.515
r141 4 45 600 $w=1.7e-07 $l=1.09622e-06 $layer=licon1_PDIFF $count=1 $X=3.095
+ $Y=1.81 $X2=3.33 $Y2=2.795
r142 3 38 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=1.03
+ $Y=1.96 $X2=1.18 $Y2=2.815
r143 3 19 400 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=1 $X=1.03
+ $Y=1.96 $X2=1.18 $Y2=2.135
r144 2 35 182 $w=1.7e-07 $l=3.27605e-07 $layer=licon1_NDIFF $count=1 $X=3.11
+ $Y=0.57 $X2=3.25 $Y2=0.835
r145 1 15 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1 $Y=0.37
+ $X2=1.14 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__FAH_4%A_427_362# 1 2 3 4 14 16 19 21 22 23 26 33 35
c88 23 0 1.26128e-19 $X=4.367 $Y=2.072
c89 21 0 1.91633e-19 $X=4.23 $Y=2.375
c90 16 0 1.07671e-19 $X=2.34 $Y=1.955
r91 31 33 8.2628 $w=2.63e-07 $l=1.9e-07 $layer=LI1_cond $X=4.23 $Y=1.177
+ $X2=4.42 $Y2=1.177
r92 27 33 3.33486 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=4.42 $Y=1.31
+ $X2=4.42 $Y2=1.177
r93 27 35 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=4.42 $Y=1.31
+ $X2=4.42 $Y2=1.935
r94 24 26 7.96233 $w=2.73e-07 $l=1.9e-07 $layer=LI1_cond $X=4.367 $Y=2.29
+ $X2=4.367 $Y2=2.1
r95 23 35 7.41084 $w=2.73e-07 $l=1.37e-07 $layer=LI1_cond $X=4.367 $Y=2.072
+ $X2=4.367 $Y2=1.935
r96 23 26 1.1734 $w=2.73e-07 $l=2.8e-08 $layer=LI1_cond $X=4.367 $Y=2.072
+ $X2=4.367 $Y2=2.1
r97 21 38 5.44791 $w=2.73e-07 $l=1.3e-07 $layer=LI1_cond $X=4.367 $Y=2.375
+ $X2=4.367 $Y2=2.505
r98 21 24 3.5621 $w=2.73e-07 $l=8.5e-08 $layer=LI1_cond $X=4.367 $Y=2.375
+ $X2=4.367 $Y2=2.29
r99 21 22 112.54 $w=1.68e-07 $l=1.725e-06 $layer=LI1_cond $X=4.23 $Y=2.375
+ $X2=2.505 $Y2=2.375
r100 19 29 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=2.39 $Y=0.895
+ $X2=2.39 $Y2=1.79
r101 16 29 7.72582 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.34 $Y=1.955
+ $X2=2.34 $Y2=1.79
r102 14 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.34 $Y=2.29
+ $X2=2.505 $Y2=2.375
r103 14 16 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.34 $Y=2.29
+ $X2=2.34 $Y2=1.955
r104 4 38 600 $w=1.7e-07 $l=7.66339e-07 $layer=licon1_PDIFF $count=1 $X=4.165
+ $Y=1.81 $X2=4.315 $Y2=2.505
r105 4 26 600 $w=1.7e-07 $l=3.57211e-07 $layer=licon1_PDIFF $count=1 $X=4.165
+ $Y=1.81 $X2=4.315 $Y2=2.1
r106 3 16 300 $w=1.7e-07 $l=2.67862e-07 $layer=licon1_PDIFF $count=2 $X=2.135
+ $Y=1.81 $X2=2.34 $Y2=1.955
r107 2 31 182 $w=1.7e-07 $l=5.50568e-07 $layer=licon1_NDIFF $count=1 $X=4.09
+ $Y=0.65 $X2=4.23 $Y2=1.135
r108 1 19 182 $w=1.7e-07 $l=5.09166e-07 $layer=licon1_NDIFF $count=1 $X=2.205
+ $Y=0.47 $X2=2.39 $Y2=0.895
.ends

.subckt PM_SKY130_FD_SC_LS__FAH_4%A_1183_102# 1 2 3 13 14 20 23 26 27 33 34 38
c109 38 0 1.08608e-19 $X=6.06 $Y=1.665
c110 34 0 5.50318e-20 $X=9.36 $Y=1.665
c111 27 0 7.63717e-20 $X=6.145 $Y=1.665
r112 34 41 14.808 $w=2.76e-07 $l=3.35e-07 $layer=LI1_cond $X=9.215 $Y=1.665
+ $X2=9.215 $Y2=2
r113 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=1.665
+ $X2=9.36 $Y2=1.665
r114 30 38 3.00637 $w=2.28e-07 $l=6e-08 $layer=LI1_cond $X=6 $Y=1.665 $X2=6.06
+ $Y2=1.665
r115 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=1.665 $X2=6
+ $Y2=1.665
r116 27 29 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.145 $Y=1.665
+ $X2=6 $Y2=1.665
r117 26 33 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.215 $Y=1.665
+ $X2=9.36 $Y2=1.665
r118 26 27 3.7995 $w=1.4e-07 $l=3.07e-06 $layer=MET1_cond $X=9.215 $Y=1.665
+ $X2=6.145 $Y2=1.665
r119 23 25 9.50985 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=6.04 $Y=0.68
+ $X2=6.04 $Y2=0.875
r120 18 34 6.87116 $w=2.76e-07 $l=1.51658e-07 $layer=LI1_cond $X=9.13 $Y=1.55
+ $X2=9.215 $Y2=1.665
r121 18 20 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=9.13 $Y=1.55
+ $X2=9.13 $Y2=1.1
r122 14 41 2.62467 $w=2e-07 $l=1.7e-07 $layer=LI1_cond $X=9.045 $Y=2 $X2=9.215
+ $Y2=2
r123 14 16 16.6364 $w=1.98e-07 $l=3e-07 $layer=LI1_cond $X=9.045 $Y=2 $X2=8.745
+ $Y2=2
r124 13 25 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=6.06 $Y=1.02
+ $X2=6.06 $Y2=0.875
r125 11 38 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=6.06 $Y=1.55
+ $X2=6.06 $Y2=1.665
r126 11 13 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=6.06 $Y=1.55
+ $X2=6.06 $Y2=1.02
r127 3 16 600 $w=1.7e-07 $l=2.86793e-07 $layer=licon1_PDIFF $count=1 $X=8.51
+ $Y=2.115 $X2=8.745 $Y2=2
r128 2 20 182 $w=1.7e-07 $l=5.67891e-07 $layer=licon1_NDIFF $count=1 $X=8.985
+ $Y=0.6 $X2=9.13 $Y2=1.1
r129 1 23 182 $w=1.7e-07 $l=2.23942e-07 $layer=licon1_NDIFF $count=1 $X=5.915
+ $Y=0.51 $X2=6.04 $Y2=0.68
r130 1 13 182 $w=1.7e-07 $l=5.77971e-07 $layer=licon1_NDIFF $count=1 $X=5.915
+ $Y=0.51 $X2=6.06 $Y2=1.02
.ends

.subckt PM_SKY130_FD_SC_LS__FAH_4%COUT 1 2 3 4 13 17 23 26 27 30
r46 27 30 4.90119 $w=4.33e-07 $l=1.85e-07 $layer=LI1_cond $X=11.177 $Y=1.85
+ $X2=11.177 $Y2=1.665
r47 27 29 2.73535 $w=4.35e-07 $l=1.25e-07 $layer=LI1_cond $X=11.177 $Y=1.85
+ $X2=11.177 $Y2=1.975
r48 25 30 10.7296 $w=4.33e-07 $l=4.05e-07 $layer=LI1_cond $X=11.177 $Y=1.26
+ $X2=11.177 $Y2=1.665
r49 25 26 1.09397 $w=4.35e-07 $l=1.25e-07 $layer=LI1_cond $X=11.177 $Y=1.26
+ $X2=11.177 $Y2=1.135
r50 21 26 9.00716 $w=2.1e-07 $l=2.18e-07 $layer=LI1_cond $X=11.395 $Y=1.135
+ $X2=11.177 $Y2=1.135
r51 21 23 10.372 $w=2.48e-07 $l=2.25e-07 $layer=LI1_cond $X=11.395 $Y=1.135
+ $X2=11.62 $Y2=1.135
r52 17 26 9.00716 $w=2.1e-07 $l=2.36155e-07 $layer=LI1_cond $X=10.96 $Y=1.095
+ $X2=11.177 $Y2=1.135
r53 17 19 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=10.96 $Y=1.095
+ $X2=10.64 $Y2=1.095
r54 13 29 4.74857 $w=2.5e-07 $l=2.17e-07 $layer=LI1_cond $X=10.96 $Y=1.975
+ $X2=11.177 $Y2=1.975
r55 13 15 41.7184 $w=2.48e-07 $l=9.05e-07 $layer=LI1_cond $X=10.96 $Y=1.975
+ $X2=10.055 $Y2=1.975
r56 4 29 600 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=1 $X=10.975
+ $Y=1.84 $X2=11.125 $Y2=2.015
r57 3 15 600 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=1 $X=9.905
+ $Y=1.84 $X2=10.055 $Y2=2.015
r58 2 23 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=11.48
+ $Y=0.5 $X2=11.62 $Y2=1.095
r59 1 19 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=10.5
+ $Y=0.5 $X2=10.64 $Y2=1.095
.ends

.subckt PM_SKY130_FD_SC_LS__FAH_4%SUM 1 2 3 4 13 15 19 21 23 24 27 30 34 35 36
+ 37 44
c64 35 0 6.40318e-20 $X=14.555 $Y=1.95
c65 19 0 1.44963e-19 $X=13.72 $Y=0.645
r66 42 44 0.516019 $w=3.33e-07 $l=1.5e-08 $layer=LI1_cond $X=14.587 $Y=2.02
+ $X2=14.587 $Y2=2.035
r67 36 37 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=14.587 $Y=2.405
+ $X2=14.587 $Y2=2.775
r68 35 42 3.22182 $w=2.92e-07 $l=8.5e-08 $layer=LI1_cond $X=14.587 $Y=1.935
+ $X2=14.587 $Y2=2.02
r69 35 36 11.5244 $w=3.33e-07 $l=3.35e-07 $layer=LI1_cond $X=14.587 $Y=2.07
+ $X2=14.587 $Y2=2.405
r70 35 44 1.20404 $w=3.33e-07 $l=3.5e-08 $layer=LI1_cond $X=14.587 $Y=2.07
+ $X2=14.587 $Y2=2.035
r71 30 35 3.22182 $w=2.92e-07 $l=1.0015e-07 $layer=LI1_cond $X=14.62 $Y=1.85
+ $X2=14.587 $Y2=1.935
r72 29 34 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=14.62 $Y=1.18
+ $X2=14.62 $Y2=1.095
r73 29 30 30.8855 $w=2.48e-07 $l=6.7e-07 $layer=LI1_cond $X=14.62 $Y=1.18
+ $X2=14.62 $Y2=1.85
r74 25 34 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=14.62 $Y=1.01
+ $X2=14.62 $Y2=1.095
r75 25 27 16.8257 $w=2.48e-07 $l=3.65e-07 $layer=LI1_cond $X=14.62 $Y=1.01
+ $X2=14.62 $Y2=0.645
r76 23 34 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=14.495 $Y=1.095
+ $X2=14.62 $Y2=1.095
r77 23 24 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=14.495 $Y=1.095
+ $X2=13.805 $Y2=1.095
r78 22 32 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.75 $Y=1.935
+ $X2=13.585 $Y2=1.935
r79 21 35 3.35233 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=14.42 $Y=1.935
+ $X2=14.587 $Y2=1.935
r80 21 22 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=14.42 $Y=1.935
+ $X2=13.75 $Y2=1.935
r81 17 24 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=13.68 $Y=1.01
+ $X2=13.805 $Y2=1.095
r82 17 19 16.8257 $w=2.48e-07 $l=3.65e-07 $layer=LI1_cond $X=13.68 $Y=1.01
+ $X2=13.68 $Y2=0.645
r83 13 32 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.585 $Y=2.02
+ $X2=13.585 $Y2=1.935
r84 13 15 27.7634 $w=3.28e-07 $l=7.95e-07 $layer=LI1_cond $X=13.585 $Y=2.02
+ $X2=13.585 $Y2=2.815
r85 4 35 400 $w=1.7e-07 $l=2.42126e-07 $layer=licon1_PDIFF $count=1 $X=14.425
+ $Y=1.84 $X2=14.585 $Y2=2.015
r86 4 37 400 $w=1.7e-07 $l=1.05196e-06 $layer=licon1_PDIFF $count=1 $X=14.425
+ $Y=1.84 $X2=14.585 $Y2=2.815
r87 3 32 400 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=1 $X=13.435
+ $Y=1.84 $X2=13.585 $Y2=2.015
r88 3 15 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=13.435
+ $Y=1.84 $X2=13.585 $Y2=2.815
r89 2 34 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=14.44
+ $Y=0.5 $X2=14.58 $Y2=1.095
r90 2 27 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=14.44
+ $Y=0.5 $X2=14.58 $Y2=0.645
r91 1 19 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=13.58
+ $Y=0.5 $X2=13.72 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_LS__FAH_4%VGND 1 2 3 4 5 6 7 8 9 30 34 38 42 46 50 54 58
+ 60 62 65 66 68 69 71 72 74 75 77 78 79 85 108 112 117 123 126 129 133
r161 132 133 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.12 $Y=0
+ $X2=15.12 $Y2=0
r162 129 130 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.16 $Y=0
+ $X2=14.16 $Y2=0
r163 126 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=0
+ $X2=13.2 $Y2=0
r164 123 124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0
+ $X2=1.68 $Y2=0
r165 121 133 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.64 $Y=0
+ $X2=15.12 $Y2=0
r166 121 130 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.64 $Y=0
+ $X2=14.16 $Y2=0
r167 120 121 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.64 $Y=0
+ $X2=14.64 $Y2=0
r168 118 129 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.315 $Y=0
+ $X2=14.15 $Y2=0
r169 118 120 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=14.315 $Y=0
+ $X2=14.64 $Y2=0
r170 117 132 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=14.915 $Y=0
+ $X2=15.137 $Y2=0
r171 117 120 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=14.915 $Y=0
+ $X2=14.64 $Y2=0
r172 116 130 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=0
+ $X2=14.16 $Y2=0
r173 116 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=0
+ $X2=13.2 $Y2=0
r174 115 116 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=0
+ $X2=13.68 $Y2=0
r175 113 126 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=13.375 $Y=0
+ $X2=13.205 $Y2=0
r176 113 115 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=13.375 $Y=0
+ $X2=13.68 $Y2=0
r177 112 129 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.985 $Y=0
+ $X2=14.15 $Y2=0
r178 112 115 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=13.985 $Y=0
+ $X2=13.68 $Y2=0
r179 111 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=0
+ $X2=13.2 $Y2=0
r180 110 111 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r181 108 126 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=13.035 $Y=0
+ $X2=13.205 $Y2=0
r182 108 110 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=13.035 $Y=0
+ $X2=12.72 $Y2=0
r183 107 111 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=12.72 $Y2=0
r184 106 107 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r185 104 107 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=11.76 $Y2=0
r186 103 104 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.8 $Y=0
+ $X2=10.8 $Y2=0
r187 101 104 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=10.8 $Y2=0
r188 100 101 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=9.84 $Y=0
+ $X2=9.84 $Y2=0
r189 97 100 313.155 $w=1.68e-07 $l=4.8e-06 $layer=LI1_cond $X=5.04 $Y=0 $X2=9.84
+ $Y2=0
r190 97 98 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r191 95 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r192 94 95 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r193 92 95 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=2.16 $Y=0 $X2=4.56
+ $Y2=0
r194 92 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=1.68 $Y2=0
r195 91 94 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=2.16 $Y=0 $X2=4.56
+ $Y2=0
r196 91 92 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r197 89 123 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.795 $Y=0
+ $X2=1.665 $Y2=0
r198 89 91 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.795 $Y=0
+ $X2=2.16 $Y2=0
r199 88 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r200 87 88 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r201 85 123 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.535 $Y=0
+ $X2=1.665 $Y2=0
r202 85 87 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.535 $Y=0 $X2=1.2
+ $Y2=0
r203 83 88 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r204 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r205 79 101 0.602067 $w=4.9e-07 $l=2.16e-06 $layer=MET1_cond $X=7.68 $Y=0
+ $X2=9.84 $Y2=0
r206 79 98 0.73586 $w=4.9e-07 $l=2.64e-06 $layer=MET1_cond $X=7.68 $Y=0 $X2=5.04
+ $Y2=0
r207 77 106 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=11.965 $Y=0
+ $X2=11.76 $Y2=0
r208 77 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.965 $Y=0
+ $X2=12.13 $Y2=0
r209 76 110 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=12.295 $Y=0
+ $X2=12.72 $Y2=0
r210 76 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.295 $Y=0
+ $X2=12.13 $Y2=0
r211 74 103 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=10.965 $Y=0
+ $X2=10.8 $Y2=0
r212 74 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.965 $Y=0
+ $X2=11.13 $Y2=0
r213 73 106 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=11.295 $Y=0
+ $X2=11.76 $Y2=0
r214 73 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.295 $Y=0
+ $X2=11.13 $Y2=0
r215 71 100 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=10.065 $Y=0
+ $X2=9.84 $Y2=0
r216 71 72 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.065 $Y=0
+ $X2=10.19 $Y2=0
r217 70 103 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=10.315 $Y=0
+ $X2=10.8 $Y2=0
r218 70 72 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.315 $Y=0
+ $X2=10.19 $Y2=0
r219 68 94 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=4.585 $Y=0 $X2=4.56
+ $Y2=0
r220 68 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.585 $Y=0 $X2=4.75
+ $Y2=0
r221 67 97 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=4.915 $Y=0
+ $X2=5.04 $Y2=0
r222 67 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.915 $Y=0 $X2=4.75
+ $Y2=0
r223 65 82 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0
+ $X2=0.24 $Y2=0
r224 65 66 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.67
+ $Y2=0
r225 64 87 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=0.795 $Y=0 $X2=1.2
+ $Y2=0
r226 64 66 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.795 $Y=0 $X2=0.67
+ $Y2=0
r227 60 132 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=15.08 $Y=0.085
+ $X2=15.137 $Y2=0
r228 60 62 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=15.08 $Y=0.085
+ $X2=15.08 $Y2=0.645
r229 56 129 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=14.15 $Y=0.085
+ $X2=14.15 $Y2=0
r230 56 58 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=14.15 $Y=0.085
+ $X2=14.15 $Y2=0.7
r231 52 126 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=13.205 $Y=0.085
+ $X2=13.205 $Y2=0
r232 52 54 8.47385 $w=3.38e-07 $l=2.5e-07 $layer=LI1_cond $X=13.205 $Y=0.085
+ $X2=13.205 $Y2=0.335
r233 48 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.13 $Y=0.085
+ $X2=12.13 $Y2=0
r234 48 50 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=12.13 $Y=0.085
+ $X2=12.13 $Y2=0.335
r235 44 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.13 $Y=0.085
+ $X2=11.13 $Y2=0
r236 44 46 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=11.13 $Y=0.085
+ $X2=11.13 $Y2=0.335
r237 40 72 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=10.19 $Y=0.085
+ $X2=10.19 $Y2=0
r238 40 42 11.5244 $w=2.48e-07 $l=2.5e-07 $layer=LI1_cond $X=10.19 $Y=0.085
+ $X2=10.19 $Y2=0.335
r239 36 69 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.75 $Y=0.085
+ $X2=4.75 $Y2=0
r240 36 38 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=4.75 $Y=0.085
+ $X2=4.75 $Y2=0.37
r241 32 123 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.665 $Y=0.085
+ $X2=1.665 $Y2=0
r242 32 34 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=1.665 $Y=0.085
+ $X2=1.665 $Y2=0.455
r243 28 66 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.67 $Y=0.085
+ $X2=0.67 $Y2=0
r244 28 30 18.9001 $w=2.48e-07 $l=4.1e-07 $layer=LI1_cond $X=0.67 $Y=0.085
+ $X2=0.67 $Y2=0.495
r245 9 62 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=14.87
+ $Y=0.5 $X2=15.08 $Y2=0.645
r246 8 58 182 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=1 $X=14.01
+ $Y=0.5 $X2=14.15 $Y2=0.7
r247 7 54 182 $w=1.7e-07 $l=3.60347e-07 $layer=licon1_NDIFF $count=1 $X=12.98
+ $Y=0.6 $X2=13.205 $Y2=0.335
r248 6 50 182 $w=1.7e-07 $l=2.91033e-07 $layer=licon1_NDIFF $count=1 $X=11.91
+ $Y=0.5 $X2=12.13 $Y2=0.335
r249 5 46 182 $w=1.7e-07 $l=2.70185e-07 $layer=licon1_NDIFF $count=1 $X=10.93
+ $Y=0.5 $X2=11.13 $Y2=0.335
r250 4 42 182 $w=1.7e-07 $l=7.712e-07 $layer=licon1_NDIFF $count=1 $X=9.5 $Y=0.6
+ $X2=10.15 $Y2=0.335
r251 3 38 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=4.625
+ $Y=0.225 $X2=4.75 $Y2=0.37
r252 2 34 182 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_NDIFF $count=1 $X=1.555
+ $Y=0.31 $X2=1.705 $Y2=0.455
r253 1 30 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.495
.ends

