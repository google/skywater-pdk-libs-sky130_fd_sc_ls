* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__fa_1 A B CIN VGND VNB VPB VPWR COUT SUM
M1000 a_69_260# CIN a_318_389# VPB phighvt w=1e+06u l=150000u
+  ad=3e+11p pd=2.6e+06u as=3.9175e+11p ps=3.13e+06u
M1001 a_1107_347# B VPWR VPB phighvt w=1e+06u l=150000u
+  ad=7.8e+11p pd=5.56e+06u as=2.2238e+12p ps=1.522e+07u
M1002 VGND CIN a_501_75# VNB nshort w=640000u l=150000u
+  ad=1.65875e+12p pd=1.244e+07u as=4.096e+11p ps=3.84e+06u
M1003 a_509_347# A VPWR VPB phighvt w=1e+06u l=150000u
+  ad=6.9e+11p pd=5.38e+06u as=0p ps=0u
M1004 a_501_75# a_465_249# a_69_260# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=2.496e+11p ps=2.06e+06u
M1005 a_318_389# B a_217_368# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=3.73375e+11p ps=2.92e+06u
M1006 a_509_347# a_465_249# a_69_260# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR CIN a_509_347# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_237_75# A VGND VNB nshort w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1009 a_916_347# A VPWR VPB phighvt w=1e+06u l=150000u
+  ad=3.55e+11p pd=2.71e+06u as=0p ps=0u
M1010 a_465_249# B a_916_347# VPB phighvt w=1e+06u l=150000u
+  ad=3e+11p pd=2.6e+06u as=0p ps=0u
M1011 a_217_368# A VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND B a_501_75# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_1100_75# B VGND VNB nshort w=640000u l=150000u
+  ad=8.888e+11p pd=5.27e+06u as=0p ps=0u
M1014 a_1107_347# CIN a_465_249# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_501_75# A VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_465_249# B a_936_75# VNB nshort w=640000u l=150000u
+  ad=1.792e+11p pd=1.84e+06u as=1.536e+11p ps=1.76e+06u
M1017 COUT a_465_249# VGND VNB nshort w=740000u l=150000u
+  ad=1.998e+11p pd=2.02e+06u as=0p ps=0u
M1018 VGND A a_1100_75# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR B a_509_347# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_1100_75# CIN a_465_249# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPWR a_69_260# SUM VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.192e+11p ps=2.81e+06u
M1022 VPWR A a_1107_347# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 COUT a_465_249# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.192e+11p pd=2.81e+06u as=0p ps=0u
M1024 VGND a_69_260# SUM VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1025 a_315_75# B a_237_75# VNB nshort w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1026 a_69_260# CIN a_315_75# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_936_75# A VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
