* File: sky130_fd_sc_ls__o311ai_1.pxi.spice
* Created: Fri Aug 28 13:51:51 2020
* 
x_PM_SKY130_FD_SC_LS__O311AI_1%A1 N_A1_M1002_g N_A1_c_50_n N_A1_M1003_g A1
+ N_A1_c_51_n PM_SKY130_FD_SC_LS__O311AI_1%A1
x_PM_SKY130_FD_SC_LS__O311AI_1%A2 N_A2_M1007_g N_A2_c_73_n N_A2_M1008_g A2 A2 A2
+ A2 N_A2_c_74_n PM_SKY130_FD_SC_LS__O311AI_1%A2
x_PM_SKY130_FD_SC_LS__O311AI_1%A3 N_A3_c_105_n N_A3_M1001_g N_A3_c_106_n
+ N_A3_M1009_g A3 PM_SKY130_FD_SC_LS__O311AI_1%A3
x_PM_SKY130_FD_SC_LS__O311AI_1%B1 N_B1_c_133_n N_B1_M1006_g N_B1_c_134_n
+ N_B1_M1005_g B1 PM_SKY130_FD_SC_LS__O311AI_1%B1
x_PM_SKY130_FD_SC_LS__O311AI_1%C1 N_C1_c_163_n N_C1_M1000_g N_C1_c_164_n
+ N_C1_M1004_g C1 PM_SKY130_FD_SC_LS__O311AI_1%C1
x_PM_SKY130_FD_SC_LS__O311AI_1%VPWR N_VPWR_M1003_s N_VPWR_M1006_d N_VPWR_c_187_n
+ N_VPWR_c_188_n N_VPWR_c_189_n N_VPWR_c_190_n N_VPWR_c_191_n VPWR
+ N_VPWR_c_192_n N_VPWR_c_186_n PM_SKY130_FD_SC_LS__O311AI_1%VPWR
x_PM_SKY130_FD_SC_LS__O311AI_1%Y N_Y_M1000_d N_Y_M1001_d N_Y_M1004_d N_Y_c_224_n
+ N_Y_c_225_n N_Y_c_226_n N_Y_c_222_n N_Y_c_223_n N_Y_c_228_n Y Y Y N_Y_c_229_n
+ PM_SKY130_FD_SC_LS__O311AI_1%Y
x_PM_SKY130_FD_SC_LS__O311AI_1%VGND N_VGND_M1002_s N_VGND_M1007_d N_VGND_c_270_n
+ N_VGND_c_271_n N_VGND_c_272_n VGND N_VGND_c_273_n N_VGND_c_274_n
+ N_VGND_c_275_n N_VGND_c_276_n PM_SKY130_FD_SC_LS__O311AI_1%VGND
x_PM_SKY130_FD_SC_LS__O311AI_1%A_128_74# N_A_128_74#_M1002_d N_A_128_74#_M1009_d
+ N_A_128_74#_c_305_n N_A_128_74#_c_313_n N_A_128_74#_c_306_n
+ N_A_128_74#_c_321_n N_A_128_74#_c_307_n PM_SKY130_FD_SC_LS__O311AI_1%A_128_74#
cc_1 VNB N_A1_M1002_g 0.0316595f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.74
cc_2 VNB N_A1_c_50_n 0.0290729f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.765
cc_3 VNB N_A1_c_51_n 0.0178902f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.515
cc_4 VNB N_A2_M1007_g 0.0280323f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.74
cc_5 VNB N_A2_c_73_n 0.0251122f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.765
cc_6 VNB N_A2_c_74_n 0.00519747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A3_c_105_n 0.0401467f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.35
cc_8 VNB N_A3_c_106_n 0.020506f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB A3 0.00613168f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=2.4
cc_10 VNB N_B1_c_133_n 0.0378024f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.35
cc_11 VNB N_B1_c_134_n 0.0181734f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB B1 0.00839315f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=2.4
cc_13 VNB N_C1_c_163_n 0.0227334f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.35
cc_14 VNB N_C1_c_164_n 0.0760135f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB C1 0.0124946f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=2.4
cc_16 VNB N_VPWR_c_186_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_Y_c_222_n 0.00413443f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_Y_c_223_n 0.030059f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_VGND_c_270_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=2.4
cc_20 VNB N_VGND_c_271_n 0.0451868f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_272_n 0.0115377f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.565
cc_22 VNB N_VGND_c_273_n 0.018682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_274_n 0.049013f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_275_n 0.214603f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_276_n 0.0107715f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_128_74#_c_305_n 0.00280814f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_128_74#_c_306_n 0.0102186f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.515
cc_28 VNB N_A_128_74#_c_307_n 0.00294871f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VPB N_A1_c_50_n 0.0305878f $X=-0.19 $Y=1.66 $X2=0.615 $Y2=1.765
cc_30 VPB N_A1_c_51_n 0.0132975f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.515
cc_31 VPB N_A2_c_73_n 0.0271021f $X=-0.19 $Y=1.66 $X2=0.615 $Y2=1.765
cc_32 VPB N_A2_c_74_n 0.00249661f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_33 VPB N_A3_c_105_n 0.0263097f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=1.35
cc_34 VPB N_B1_c_133_n 0.0241232f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=1.35
cc_35 VPB N_C1_c_164_n 0.0292377f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_36 VPB N_VPWR_c_187_n 0.0155194f $X=-0.19 $Y=1.66 $X2=0.615 $Y2=2.4
cc_37 VPB N_VPWR_c_188_n 0.0486246f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_38 VPB N_VPWR_c_189_n 0.00976973f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_39 VPB N_VPWR_c_190_n 0.0498591f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_40 VPB N_VPWR_c_191_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_41 VPB N_VPWR_c_192_n 0.0225072f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_42 VPB N_VPWR_c_186_n 0.0846987f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_43 VPB N_Y_c_224_n 0.00299332f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.515
cc_44 VPB N_Y_c_225_n 0.00685577f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.565
cc_45 VPB N_Y_c_226_n 0.0104779f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_Y_c_222_n 7.3943e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB N_Y_c_228_n 0.0109693f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 VPB N_Y_c_229_n 0.0503513f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 N_A1_M1002_g N_A2_M1007_g 0.0181074f $X=0.565 $Y=0.74 $X2=0 $Y2=0
cc_50 N_A1_c_50_n N_A2_c_73_n 0.0801921f $X=0.615 $Y=1.765 $X2=0 $Y2=0
cc_51 N_A1_c_51_n N_A2_c_73_n 0.00154554f $X=0.54 $Y=1.515 $X2=0 $Y2=0
cc_52 N_A1_c_50_n N_A2_c_74_n 0.00476777f $X=0.615 $Y=1.765 $X2=0 $Y2=0
cc_53 N_A1_c_51_n N_A2_c_74_n 0.0259135f $X=0.54 $Y=1.515 $X2=0 $Y2=0
cc_54 N_A1_c_50_n N_VPWR_c_188_n 0.0207617f $X=0.615 $Y=1.765 $X2=0 $Y2=0
cc_55 N_A1_c_51_n N_VPWR_c_188_n 0.0263294f $X=0.54 $Y=1.515 $X2=0 $Y2=0
cc_56 N_A1_c_50_n N_VPWR_c_190_n 0.00413917f $X=0.615 $Y=1.765 $X2=0 $Y2=0
cc_57 N_A1_c_50_n N_VPWR_c_186_n 0.00817532f $X=0.615 $Y=1.765 $X2=0 $Y2=0
cc_58 N_A1_M1002_g N_VGND_c_271_n 0.0184904f $X=0.565 $Y=0.74 $X2=0 $Y2=0
cc_59 N_A1_c_50_n N_VGND_c_271_n 0.00156574f $X=0.615 $Y=1.765 $X2=0 $Y2=0
cc_60 N_A1_c_51_n N_VGND_c_271_n 0.0236882f $X=0.54 $Y=1.515 $X2=0 $Y2=0
cc_61 N_A1_M1002_g N_VGND_c_273_n 0.00434272f $X=0.565 $Y=0.74 $X2=0 $Y2=0
cc_62 N_A1_M1002_g N_VGND_c_275_n 0.0082426f $X=0.565 $Y=0.74 $X2=0 $Y2=0
cc_63 N_A1_M1002_g N_A_128_74#_c_305_n 0.00632535f $X=0.565 $Y=0.74 $X2=0 $Y2=0
cc_64 N_A1_M1002_g N_A_128_74#_c_306_n 0.00375706f $X=0.565 $Y=0.74 $X2=0 $Y2=0
cc_65 N_A1_c_50_n N_A_128_74#_c_306_n 0.0016773f $X=0.615 $Y=1.765 $X2=0 $Y2=0
cc_66 N_A1_c_51_n N_A_128_74#_c_306_n 0.00625586f $X=0.54 $Y=1.515 $X2=0 $Y2=0
cc_67 N_A2_M1007_g N_A3_c_105_n 0.00407278f $X=1.02 $Y=0.74 $X2=-0.19 $Y2=-0.245
cc_68 N_A2_c_73_n N_A3_c_105_n 0.0518845f $X=1.035 $Y=1.765 $X2=-0.19 $Y2=-0.245
cc_69 N_A2_c_74_n N_A3_c_105_n 0.0172184f $X=1.11 $Y=1.515 $X2=-0.19 $Y2=-0.245
cc_70 N_A2_M1007_g N_A3_c_106_n 0.0162896f $X=1.02 $Y=0.74 $X2=0 $Y2=0
cc_71 N_A2_M1007_g A3 0.00151734f $X=1.02 $Y=0.74 $X2=0 $Y2=0
cc_72 N_A2_c_73_n A3 2.36557e-19 $X=1.035 $Y=1.765 $X2=0 $Y2=0
cc_73 N_A2_c_74_n A3 0.0141439f $X=1.11 $Y=1.515 $X2=0 $Y2=0
cc_74 N_A2_c_73_n N_VPWR_c_188_n 0.00195439f $X=1.035 $Y=1.765 $X2=0 $Y2=0
cc_75 N_A2_c_73_n N_VPWR_c_190_n 0.00303293f $X=1.035 $Y=1.765 $X2=0 $Y2=0
cc_76 N_A2_c_74_n N_VPWR_c_190_n 0.0103587f $X=1.11 $Y=1.515 $X2=0 $Y2=0
cc_77 N_A2_c_73_n N_VPWR_c_186_n 0.00372936f $X=1.035 $Y=1.765 $X2=0 $Y2=0
cc_78 N_A2_c_74_n N_VPWR_c_186_n 0.0120835f $X=1.11 $Y=1.515 $X2=0 $Y2=0
cc_79 N_A2_c_74_n A_222_368# 0.0173967f $X=1.11 $Y=1.515 $X2=-0.19 $Y2=-0.245
cc_80 N_A2_c_74_n N_Y_c_224_n 0.0380365f $X=1.11 $Y=1.515 $X2=0 $Y2=0
cc_81 N_A2_c_74_n N_Y_c_226_n 0.00726306f $X=1.11 $Y=1.515 $X2=0 $Y2=0
cc_82 N_A2_M1007_g N_VGND_c_272_n 0.00488678f $X=1.02 $Y=0.74 $X2=0 $Y2=0
cc_83 N_A2_M1007_g N_VGND_c_273_n 0.00461464f $X=1.02 $Y=0.74 $X2=0 $Y2=0
cc_84 N_A2_M1007_g N_VGND_c_275_n 0.00465508f $X=1.02 $Y=0.74 $X2=0 $Y2=0
cc_85 N_A2_M1007_g N_A_128_74#_c_305_n 4.71232e-19 $X=1.02 $Y=0.74 $X2=0 $Y2=0
cc_86 N_A2_M1007_g N_A_128_74#_c_313_n 0.0120154f $X=1.02 $Y=0.74 $X2=0 $Y2=0
cc_87 N_A2_c_73_n N_A_128_74#_c_313_n 9.22877e-19 $X=1.035 $Y=1.765 $X2=0 $Y2=0
cc_88 N_A2_c_74_n N_A_128_74#_c_313_n 0.0155033f $X=1.11 $Y=1.515 $X2=0 $Y2=0
cc_89 N_A2_M1007_g N_A_128_74#_c_306_n 0.00106811f $X=1.02 $Y=0.74 $X2=0 $Y2=0
cc_90 N_A3_c_105_n N_B1_c_133_n 0.0421056f $X=1.605 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_91 A3 N_B1_c_133_n 3.90318e-19 $X=1.595 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_92 N_A3_c_106_n N_B1_c_134_n 0.0200745f $X=1.77 $Y=1.22 $X2=0 $Y2=0
cc_93 N_A3_c_106_n B1 0.00229487f $X=1.77 $Y=1.22 $X2=0 $Y2=0
cc_94 A3 B1 0.0261333f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_95 N_A3_c_105_n N_VPWR_c_190_n 0.00461464f $X=1.605 $Y=1.765 $X2=0 $Y2=0
cc_96 N_A3_c_105_n N_VPWR_c_186_n 0.00911823f $X=1.605 $Y=1.765 $X2=0 $Y2=0
cc_97 N_A3_c_105_n N_Y_c_224_n 0.0149125f $X=1.605 $Y=1.765 $X2=0 $Y2=0
cc_98 N_A3_c_105_n N_Y_c_226_n 0.00283079f $X=1.605 $Y=1.765 $X2=0 $Y2=0
cc_99 A3 N_Y_c_226_n 0.00503923f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_100 N_A3_c_106_n N_VGND_c_272_n 0.00603858f $X=1.77 $Y=1.22 $X2=0 $Y2=0
cc_101 N_A3_c_106_n N_VGND_c_274_n 0.00461464f $X=1.77 $Y=1.22 $X2=0 $Y2=0
cc_102 N_A3_c_106_n N_VGND_c_275_n 0.00465894f $X=1.77 $Y=1.22 $X2=0 $Y2=0
cc_103 N_A3_c_105_n N_A_128_74#_c_313_n 9.99496e-19 $X=1.605 $Y=1.765 $X2=0
+ $Y2=0
cc_104 N_A3_c_106_n N_A_128_74#_c_313_n 0.0134555f $X=1.77 $Y=1.22 $X2=0 $Y2=0
cc_105 A3 N_A_128_74#_c_313_n 0.0228656f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_106 N_A3_c_106_n N_A_128_74#_c_307_n 0.00281817f $X=1.77 $Y=1.22 $X2=0 $Y2=0
cc_107 N_B1_c_134_n N_C1_c_163_n 0.0363339f $X=2.27 $Y=1.22 $X2=-0.19 $Y2=-0.245
cc_108 N_B1_c_133_n N_C1_c_164_n 0.0503808f $X=2.175 $Y=1.765 $X2=0 $Y2=0
cc_109 B1 N_C1_c_164_n 3.61714e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_110 N_B1_c_133_n N_VPWR_c_189_n 0.00899555f $X=2.175 $Y=1.765 $X2=0 $Y2=0
cc_111 N_B1_c_133_n N_VPWR_c_190_n 0.00445602f $X=2.175 $Y=1.765 $X2=0 $Y2=0
cc_112 N_B1_c_133_n N_VPWR_c_186_n 0.00859027f $X=2.175 $Y=1.765 $X2=0 $Y2=0
cc_113 N_B1_c_133_n N_Y_c_224_n 0.0132476f $X=2.175 $Y=1.765 $X2=0 $Y2=0
cc_114 N_B1_c_133_n N_Y_c_225_n 0.0140317f $X=2.175 $Y=1.765 $X2=0 $Y2=0
cc_115 B1 N_Y_c_225_n 0.0221856f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_116 N_B1_c_133_n N_Y_c_226_n 0.00266249f $X=2.175 $Y=1.765 $X2=0 $Y2=0
cc_117 B1 N_Y_c_226_n 0.00592165f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_118 N_B1_c_133_n N_Y_c_222_n 0.00525331f $X=2.175 $Y=1.765 $X2=0 $Y2=0
cc_119 B1 N_Y_c_222_n 0.0282201f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_120 N_B1_c_134_n N_Y_c_223_n 0.00893686f $X=2.27 $Y=1.22 $X2=0 $Y2=0
cc_121 N_B1_c_133_n N_Y_c_229_n 9.55735e-19 $X=2.175 $Y=1.765 $X2=0 $Y2=0
cc_122 N_B1_c_134_n N_VGND_c_274_n 0.00433834f $X=2.27 $Y=1.22 $X2=0 $Y2=0
cc_123 N_B1_c_134_n N_VGND_c_275_n 0.00822046f $X=2.27 $Y=1.22 $X2=0 $Y2=0
cc_124 N_B1_c_133_n N_A_128_74#_c_321_n 6.10824e-19 $X=2.175 $Y=1.765 $X2=0
+ $Y2=0
cc_125 N_B1_c_134_n N_A_128_74#_c_321_n 0.00280745f $X=2.27 $Y=1.22 $X2=0 $Y2=0
cc_126 B1 N_A_128_74#_c_321_n 0.0124978f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_127 N_B1_c_134_n N_A_128_74#_c_307_n 0.00863906f $X=2.27 $Y=1.22 $X2=0 $Y2=0
cc_128 N_C1_c_164_n N_VPWR_c_189_n 0.00868976f $X=2.745 $Y=1.765 $X2=0 $Y2=0
cc_129 N_C1_c_164_n N_VPWR_c_192_n 0.00445602f $X=2.745 $Y=1.765 $X2=0 $Y2=0
cc_130 N_C1_c_164_n N_VPWR_c_186_n 0.00862226f $X=2.745 $Y=1.765 $X2=0 $Y2=0
cc_131 N_C1_c_164_n N_Y_c_224_n 9.39715e-19 $X=2.745 $Y=1.765 $X2=0 $Y2=0
cc_132 N_C1_c_163_n N_Y_c_222_n 0.00786229f $X=2.73 $Y=1.22 $X2=0 $Y2=0
cc_133 N_C1_c_164_n N_Y_c_222_n 0.016326f $X=2.745 $Y=1.765 $X2=0 $Y2=0
cc_134 C1 N_Y_c_222_n 0.0265523f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_135 N_C1_c_163_n N_Y_c_223_n 0.0179308f $X=2.73 $Y=1.22 $X2=0 $Y2=0
cc_136 N_C1_c_164_n N_Y_c_223_n 0.00518195f $X=2.745 $Y=1.765 $X2=0 $Y2=0
cc_137 C1 N_Y_c_223_n 0.0160699f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_138 N_C1_c_164_n N_Y_c_228_n 0.0251189f $X=2.745 $Y=1.765 $X2=0 $Y2=0
cc_139 C1 N_Y_c_228_n 0.0263919f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_140 N_C1_c_164_n N_Y_c_229_n 0.0143516f $X=2.745 $Y=1.765 $X2=0 $Y2=0
cc_141 N_C1_c_163_n N_VGND_c_274_n 0.00291513f $X=2.73 $Y=1.22 $X2=0 $Y2=0
cc_142 N_C1_c_163_n N_VGND_c_275_n 0.00363424f $X=2.73 $Y=1.22 $X2=0 $Y2=0
cc_143 N_C1_c_163_n N_A_128_74#_c_307_n 5.78724e-19 $X=2.73 $Y=1.22 $X2=0 $Y2=0
cc_144 N_VPWR_c_189_n N_Y_c_224_n 0.0353111f $X=2.45 $Y=2.145 $X2=0 $Y2=0
cc_145 N_VPWR_c_190_n N_Y_c_224_n 0.0145938f $X=2.285 $Y=3.33 $X2=0 $Y2=0
cc_146 N_VPWR_c_186_n N_Y_c_224_n 0.0120466f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_147 N_VPWR_M1006_d N_Y_c_225_n 0.00302593f $X=2.25 $Y=1.84 $X2=0 $Y2=0
cc_148 N_VPWR_c_189_n N_Y_c_225_n 0.0225812f $X=2.45 $Y=2.145 $X2=0 $Y2=0
cc_149 N_VPWR_M1006_d N_Y_c_228_n 3.09855e-19 $X=2.25 $Y=1.84 $X2=0 $Y2=0
cc_150 N_VPWR_c_189_n N_Y_c_228_n 0.00252453f $X=2.45 $Y=2.145 $X2=0 $Y2=0
cc_151 N_VPWR_c_189_n N_Y_c_229_n 0.0336136f $X=2.45 $Y=2.145 $X2=0 $Y2=0
cc_152 N_VPWR_c_192_n N_Y_c_229_n 0.0190559f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_153 N_VPWR_c_186_n N_Y_c_229_n 0.0157399f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_154 N_Y_c_223_n N_VGND_c_274_n 0.0228546f $X=2.945 $Y=0.515 $X2=0 $Y2=0
cc_155 N_Y_c_223_n N_VGND_c_275_n 0.0185794f $X=2.945 $Y=0.515 $X2=0 $Y2=0
cc_156 N_Y_c_223_n N_A_128_74#_c_321_n 0.00803923f $X=2.945 $Y=0.515 $X2=0 $Y2=0
cc_157 N_Y_c_223_n N_A_128_74#_c_307_n 0.0219699f $X=2.945 $Y=0.515 $X2=0 $Y2=0
cc_158 N_Y_c_222_n A_469_74# 0.0013188f $X=2.67 $Y=1.72 $X2=-0.19 $Y2=-0.245
cc_159 N_Y_c_223_n A_469_74# 0.00783876f $X=2.945 $Y=0.515 $X2=-0.19 $Y2=-0.245
cc_160 N_VGND_c_271_n N_A_128_74#_c_305_n 0.0191389f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_161 N_VGND_c_272_n N_A_128_74#_c_305_n 0.0132958f $X=1.405 $Y=0.515 $X2=0
+ $Y2=0
cc_162 N_VGND_c_273_n N_A_128_74#_c_305_n 0.0145639f $X=1.115 $Y=0 $X2=0 $Y2=0
cc_163 N_VGND_c_275_n N_A_128_74#_c_305_n 0.0119984f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_164 N_VGND_M1007_d N_A_128_74#_c_313_n 0.0183532f $X=1.095 $Y=0.37 $X2=0
+ $Y2=0
cc_165 N_VGND_c_272_n N_A_128_74#_c_313_n 0.0352958f $X=1.405 $Y=0.515 $X2=0
+ $Y2=0
cc_166 N_VGND_c_275_n N_A_128_74#_c_313_n 0.0130717f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_167 N_VGND_c_271_n N_A_128_74#_c_306_n 0.0124832f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_168 N_VGND_c_272_n N_A_128_74#_c_307_n 0.00286618f $X=1.405 $Y=0.515 $X2=0
+ $Y2=0
cc_169 N_VGND_c_274_n N_A_128_74#_c_307_n 0.0158357f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_170 N_VGND_c_275_n N_A_128_74#_c_307_n 0.0121432f $X=3.12 $Y=0 $X2=0 $Y2=0
