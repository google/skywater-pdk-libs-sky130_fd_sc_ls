* File: sky130_fd_sc_ls__ha_4.pxi.spice
* Created: Fri Aug 28 13:27:46 2020
* 
x_PM_SKY130_FD_SC_LS__HA_4%A_435_99# N_A_435_99#_M1001_s N_A_435_99#_M1012_s
+ N_A_435_99#_M1018_s N_A_435_99#_c_195_n N_A_435_99#_M1022_g
+ N_A_435_99#_c_196_n N_A_435_99#_c_197_n N_A_435_99#_c_198_n
+ N_A_435_99#_M1026_g N_A_435_99#_c_207_n N_A_435_99#_M1009_g
+ N_A_435_99#_c_208_n N_A_435_99#_M1016_g N_A_435_99#_c_209_n
+ N_A_435_99#_M1017_g N_A_435_99#_M1006_g N_A_435_99#_c_210_n
+ N_A_435_99#_M1025_g N_A_435_99#_M1010_g N_A_435_99#_c_211_n
+ N_A_435_99#_M1031_g N_A_435_99#_M1028_g N_A_435_99#_c_212_n
+ N_A_435_99#_M1032_g N_A_435_99#_M1030_g N_A_435_99#_c_203_n
+ N_A_435_99#_c_204_n N_A_435_99#_c_236_p N_A_435_99#_c_215_n
+ N_A_435_99#_c_216_n N_A_435_99#_c_217_n N_A_435_99#_c_205_n
+ N_A_435_99#_c_286_p N_A_435_99#_c_218_n N_A_435_99#_c_219_n
+ N_A_435_99#_c_206_n PM_SKY130_FD_SC_LS__HA_4%A_435_99#
x_PM_SKY130_FD_SC_LS__HA_4%B N_B_M1000_g N_B_c_395_n N_B_M1007_g N_B_M1004_g
+ N_B_c_396_n N_B_M1014_g N_B_c_397_n N_B_c_389_n N_B_c_399_n N_B_c_400_n
+ N_B_c_401_n N_B_c_402_n N_B_c_403_n N_B_c_390_n N_B_M1012_g N_B_M1001_g
+ N_B_c_406_n N_B_c_392_n N_B_M1035_g N_B_c_408_n N_B_M1023_g N_B_c_409_n
+ N_B_c_410_n B B PM_SKY130_FD_SC_LS__HA_4%B
x_PM_SKY130_FD_SC_LS__HA_4%A N_A_M1011_g N_A_c_534_n N_A_M1033_g N_A_M1021_g
+ N_A_c_535_n N_A_M1034_g N_A_c_524_n N_A_c_525_n N_A_c_526_n N_A_c_537_n
+ N_A_M1018_g N_A_M1002_g N_A_c_528_n N_A_c_529_n N_A_M1008_g N_A_c_538_n
+ N_A_M1019_g N_A_c_530_n N_A_c_531_n A A A N_A_c_533_n
+ PM_SKY130_FD_SC_LS__HA_4%A
x_PM_SKY130_FD_SC_LS__HA_4%A_294_392# N_A_294_392#_M1022_d N_A_294_392#_M1007_d
+ N_A_294_392#_M1009_d N_A_294_392#_c_651_n N_A_294_392#_M1005_g
+ N_A_294_392#_M1003_g N_A_294_392#_c_652_n N_A_294_392#_M1013_g
+ N_A_294_392#_M1015_g N_A_294_392#_c_653_n N_A_294_392#_M1020_g
+ N_A_294_392#_M1024_g N_A_294_392#_c_643_n N_A_294_392#_c_644_n
+ N_A_294_392#_M1027_g N_A_294_392#_c_655_n N_A_294_392#_M1029_g
+ N_A_294_392#_c_656_n N_A_294_392#_c_646_n N_A_294_392#_c_647_n
+ N_A_294_392#_c_675_n N_A_294_392#_c_677_n N_A_294_392#_c_680_n
+ N_A_294_392#_c_658_n N_A_294_392#_c_648_n N_A_294_392#_c_782_p
+ N_A_294_392#_c_649_n N_A_294_392#_c_660_n N_A_294_392#_c_650_n
+ N_A_294_392#_c_661_n N_A_294_392#_c_697_n N_A_294_392#_c_702_n
+ PM_SKY130_FD_SC_LS__HA_4%A_294_392#
x_PM_SKY130_FD_SC_LS__HA_4%A_27_392# N_A_27_392#_M1033_s N_A_27_392#_M1034_s
+ N_A_27_392#_M1014_s N_A_27_392#_c_845_n N_A_27_392#_c_846_n
+ N_A_27_392#_c_847_n N_A_27_392#_c_848_n N_A_27_392#_c_866_n
+ N_A_27_392#_c_849_n N_A_27_392#_c_850_n N_A_27_392#_c_851_n
+ PM_SKY130_FD_SC_LS__HA_4%A_27_392#
x_PM_SKY130_FD_SC_LS__HA_4%VPWR N_VPWR_M1033_d N_VPWR_M1009_s N_VPWR_M1016_s
+ N_VPWR_M1023_d N_VPWR_M1019_d N_VPWR_M1025_s N_VPWR_M1032_s N_VPWR_M1013_s
+ N_VPWR_M1029_s N_VPWR_c_890_n N_VPWR_c_891_n N_VPWR_c_892_n N_VPWR_c_893_n
+ N_VPWR_c_894_n N_VPWR_c_895_n N_VPWR_c_896_n N_VPWR_c_897_n N_VPWR_c_898_n
+ N_VPWR_c_899_n N_VPWR_c_900_n N_VPWR_c_901_n N_VPWR_c_902_n N_VPWR_c_903_n
+ N_VPWR_c_904_n N_VPWR_c_905_n N_VPWR_c_906_n VPWR N_VPWR_c_907_n
+ N_VPWR_c_908_n N_VPWR_c_909_n N_VPWR_c_910_n N_VPWR_c_911_n N_VPWR_c_912_n
+ N_VPWR_c_913_n N_VPWR_c_914_n N_VPWR_c_915_n N_VPWR_c_916_n N_VPWR_c_889_n
+ PM_SKY130_FD_SC_LS__HA_4%VPWR
x_PM_SKY130_FD_SC_LS__HA_4%COUT N_COUT_M1006_s N_COUT_M1028_s N_COUT_M1017_d
+ N_COUT_M1031_d N_COUT_c_1049_n N_COUT_c_1046_n N_COUT_c_1047_n N_COUT_c_1048_n
+ N_COUT_c_1066_n COUT COUT COUT N_COUT_c_1075_n PM_SKY130_FD_SC_LS__HA_4%COUT
x_PM_SKY130_FD_SC_LS__HA_4%SUM N_SUM_M1003_s N_SUM_M1024_s N_SUM_M1005_d
+ N_SUM_M1020_d N_SUM_c_1104_n N_SUM_c_1105_n N_SUM_c_1097_n N_SUM_c_1098_n
+ N_SUM_c_1099_n N_SUM_c_1100_n N_SUM_c_1106_n N_SUM_c_1101_n N_SUM_c_1107_n
+ N_SUM_c_1102_n N_SUM_c_1103_n N_SUM_c_1109_n N_SUM_c_1110_n N_SUM_c_1151_n
+ N_SUM_c_1152_n SUM PM_SKY130_FD_SC_LS__HA_4%SUM
x_PM_SKY130_FD_SC_LS__HA_4%A_27_125# N_A_27_125#_M1011_d N_A_27_125#_M1021_d
+ N_A_27_125#_M1004_s N_A_27_125#_M1026_s N_A_27_125#_c_1186_n
+ N_A_27_125#_c_1187_n N_A_27_125#_c_1188_n N_A_27_125#_c_1189_n
+ N_A_27_125#_c_1190_n N_A_27_125#_c_1191_n N_A_27_125#_c_1192_n
+ N_A_27_125#_c_1193_n N_A_27_125#_c_1194_n N_A_27_125#_c_1195_n
+ PM_SKY130_FD_SC_LS__HA_4%A_27_125#
x_PM_SKY130_FD_SC_LS__HA_4%VGND N_VGND_M1011_s N_VGND_M1000_d N_VGND_M1002_d
+ N_VGND_M1006_d N_VGND_M1010_d N_VGND_M1030_d N_VGND_M1015_d N_VGND_M1027_d
+ N_VGND_c_1252_n N_VGND_c_1253_n N_VGND_c_1254_n N_VGND_c_1255_n
+ N_VGND_c_1256_n N_VGND_c_1257_n N_VGND_c_1258_n N_VGND_c_1259_n
+ N_VGND_c_1260_n N_VGND_c_1261_n N_VGND_c_1262_n N_VGND_c_1263_n
+ N_VGND_c_1264_n N_VGND_c_1265_n N_VGND_c_1266_n N_VGND_c_1267_n
+ N_VGND_c_1268_n N_VGND_c_1269_n VGND N_VGND_c_1270_n N_VGND_c_1271_n
+ N_VGND_c_1272_n N_VGND_c_1273_n N_VGND_c_1274_n N_VGND_c_1275_n
+ N_VGND_c_1276_n PM_SKY130_FD_SC_LS__HA_4%VGND
x_PM_SKY130_FD_SC_LS__HA_4%A_707_119# N_A_707_119#_M1001_d N_A_707_119#_M1035_d
+ N_A_707_119#_M1008_s N_A_707_119#_c_1378_n N_A_707_119#_c_1379_n
+ N_A_707_119#_c_1380_n N_A_707_119#_c_1381_n N_A_707_119#_c_1382_n
+ N_A_707_119#_c_1383_n N_A_707_119#_c_1384_n
+ PM_SKY130_FD_SC_LS__HA_4%A_707_119#
cc_1 VNB N_A_435_99#_c_195_n 0.0138943f $X=-0.19 $Y=-0.245 $X2=2.25 $Y2=1.34
cc_2 VNB N_A_435_99#_c_196_n 0.0163286f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=1.415
cc_3 VNB N_A_435_99#_c_197_n 0.00729893f $X=-0.19 $Y=-0.245 $X2=2.325 $Y2=1.415
cc_4 VNB N_A_435_99#_c_198_n 0.0156514f $X=-0.19 $Y=-0.245 $X2=2.72 $Y2=1.34
cc_5 VNB N_A_435_99#_M1006_g 0.0248403f $X=-0.19 $Y=-0.245 $X2=6.3 $Y2=0.74
cc_6 VNB N_A_435_99#_M1010_g 0.0213542f $X=-0.19 $Y=-0.245 $X2=6.73 $Y2=0.74
cc_7 VNB N_A_435_99#_M1028_g 0.0205795f $X=-0.19 $Y=-0.245 $X2=7.16 $Y2=0.74
cc_8 VNB N_A_435_99#_M1030_g 0.0210466f $X=-0.19 $Y=-0.245 $X2=7.59 $Y2=0.74
cc_9 VNB N_A_435_99#_c_203_n 0.00843023f $X=-0.19 $Y=-0.245 $X2=3.9 $Y2=1.57
cc_10 VNB N_A_435_99#_c_204_n 0.0605391f $X=-0.19 $Y=-0.245 $X2=3.24 $Y2=1.57
cc_11 VNB N_A_435_99#_c_205_n 0.00567831f $X=-0.19 $Y=-0.245 $X2=6.05 $Y2=1.485
cc_12 VNB N_A_435_99#_c_206_n 0.12194f $X=-0.19 $Y=-0.245 $X2=7.515 $Y2=1.542
cc_13 VNB N_B_M1000_g 0.0185323f $X=-0.19 $Y=-0.245 $X2=4.895 $Y2=2.05
cc_14 VNB N_B_M1004_g 0.0186662f $X=-0.19 $Y=-0.245 $X2=2.25 $Y2=1.34
cc_15 VNB N_B_c_389_n 0.0268913f $X=-0.19 $Y=-0.245 $X2=2.72 $Y2=0.945
cc_16 VNB N_B_c_390_n 0.00674158f $X=-0.19 $Y=-0.245 $X2=3.315 $Y2=2.315
cc_17 VNB N_B_M1001_g 0.025966f $X=-0.19 $Y=-0.245 $X2=6.3 $Y2=0.74
cc_18 VNB N_B_c_392_n 0.00653496f $X=-0.19 $Y=-0.245 $X2=6.615 $Y2=2.4
cc_19 VNB N_B_M1035_g 0.0231254f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB B 0.0037323f $X=-0.19 $Y=-0.245 $X2=7.515 $Y2=2.4
cc_21 VNB N_A_M1011_g 0.0287386f $X=-0.19 $Y=-0.245 $X2=4.895 $Y2=2.05
cc_22 VNB N_A_M1021_g 0.0316014f $X=-0.19 $Y=-0.245 $X2=2.25 $Y2=0.945
cc_23 VNB N_A_c_524_n 0.283484f $X=-0.19 $Y=-0.245 $X2=2.72 $Y2=1.34
cc_24 VNB N_A_c_525_n 0.0125033f $X=-0.19 $Y=-0.245 $X2=2.72 $Y2=0.945
cc_25 VNB N_A_c_526_n 9.04456e-19 $X=-0.19 $Y=-0.245 $X2=2.865 $Y2=1.82
cc_26 VNB N_A_M1002_g 0.0253437f $X=-0.19 $Y=-0.245 $X2=6.005 $Y2=2.4
cc_27 VNB N_A_c_528_n 0.0242815f $X=-0.19 $Y=-0.245 $X2=6.005 $Y2=2.4
cc_28 VNB N_A_c_529_n 0.0163093f $X=-0.19 $Y=-0.245 $X2=6.3 $Y2=0.74
cc_29 VNB N_A_c_530_n 0.0103242f $X=-0.19 $Y=-0.245 $X2=6.73 $Y2=1.32
cc_30 VNB N_A_c_531_n 0.0159256f $X=-0.19 $Y=-0.245 $X2=6.73 $Y2=0.74
cc_31 VNB A 0.0142582f $X=-0.19 $Y=-0.245 $X2=7.065 $Y2=1.765
cc_32 VNB N_A_c_533_n 0.024547f $X=-0.19 $Y=-0.245 $X2=7.515 $Y2=2.4
cc_33 VNB N_A_294_392#_M1003_g 0.0219202f $X=-0.19 $Y=-0.245 $X2=2.72 $Y2=1.34
cc_34 VNB N_A_294_392#_M1015_g 0.0226903f $X=-0.19 $Y=-0.245 $X2=3.315 $Y2=2.315
cc_35 VNB N_A_294_392#_M1024_g 0.0237211f $X=-0.19 $Y=-0.245 $X2=6.3 $Y2=0.74
cc_36 VNB N_A_294_392#_c_643_n 0.02964f $X=-0.19 $Y=-0.245 $X2=6.615 $Y2=1.765
cc_37 VNB N_A_294_392#_c_644_n 0.0706582f $X=-0.19 $Y=-0.245 $X2=6.615 $Y2=2.4
cc_38 VNB N_A_294_392#_M1027_g 0.0256152f $X=-0.19 $Y=-0.245 $X2=6.73 $Y2=0.74
cc_39 VNB N_A_294_392#_c_646_n 0.00202173f $X=-0.19 $Y=-0.245 $X2=7.515 $Y2=2.4
cc_40 VNB N_A_294_392#_c_647_n 0.00324153f $X=-0.19 $Y=-0.245 $X2=7.59 $Y2=0.74
cc_41 VNB N_A_294_392#_c_648_n 0.00477785f $X=-0.19 $Y=-0.245 $X2=4.115 $Y2=0.74
cc_42 VNB N_A_294_392#_c_649_n 0.0258827f $X=-0.19 $Y=-0.245 $X2=5.12 $Y2=1.985
cc_43 VNB N_A_294_392#_c_650_n 0.00162343f $X=-0.19 $Y=-0.245 $X2=5.965 $Y2=1.82
cc_44 VNB N_VPWR_c_889_n 0.422413f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_COUT_c_1046_n 0.00186123f $X=-0.19 $Y=-0.245 $X2=2.72 $Y2=0.945
cc_46 VNB N_COUT_c_1047_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=2.865 $Y2=2.315
cc_47 VNB N_COUT_c_1048_n 0.00541261f $X=-0.19 $Y=-0.245 $X2=3.315 $Y2=1.82
cc_48 VNB N_SUM_c_1097_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=2.865 $Y2=2.315
cc_49 VNB N_SUM_c_1098_n 0.00307912f $X=-0.19 $Y=-0.245 $X2=3.315 $Y2=1.82
cc_50 VNB N_SUM_c_1099_n 0.00220472f $X=-0.19 $Y=-0.245 $X2=3.315 $Y2=2.315
cc_51 VNB N_SUM_c_1100_n 0.00327315f $X=-0.19 $Y=-0.245 $X2=6.005 $Y2=2.4
cc_52 VNB N_SUM_c_1101_n 0.0154148f $X=-0.19 $Y=-0.245 $X2=6.615 $Y2=1.765
cc_53 VNB N_SUM_c_1102_n 0.0244077f $X=-0.19 $Y=-0.245 $X2=6.73 $Y2=0.74
cc_54 VNB N_SUM_c_1103_n 0.00241905f $X=-0.19 $Y=-0.245 $X2=7.065 $Y2=2.4
cc_55 VNB N_A_27_125#_c_1186_n 0.0221323f $X=-0.19 $Y=-0.245 $X2=2.72 $Y2=1.34
cc_56 VNB N_A_27_125#_c_1187_n 0.0027328f $X=-0.19 $Y=-0.245 $X2=2.72 $Y2=0.945
cc_57 VNB N_A_27_125#_c_1188_n 0.00952244f $X=-0.19 $Y=-0.245 $X2=2.865 $Y2=1.82
cc_58 VNB N_A_27_125#_c_1189_n 0.00244123f $X=-0.19 $Y=-0.245 $X2=3.315 $Y2=1.82
cc_59 VNB N_A_27_125#_c_1190_n 0.00620491f $X=-0.19 $Y=-0.245 $X2=3.315
+ $Y2=2.315
cc_60 VNB N_A_27_125#_c_1191_n 0.00337282f $X=-0.19 $Y=-0.245 $X2=6.3 $Y2=0.74
cc_61 VNB N_A_27_125#_c_1192_n 0.0216937f $X=-0.19 $Y=-0.245 $X2=6.3 $Y2=0.74
cc_62 VNB N_A_27_125#_c_1193_n 0.00432301f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_27_125#_c_1194_n 0.0134046f $X=-0.19 $Y=-0.245 $X2=6.615 $Y2=2.4
cc_64 VNB N_A_27_125#_c_1195_n 0.00207245f $X=-0.19 $Y=-0.245 $X2=6.73 $Y2=0.74
cc_65 VNB N_VGND_c_1252_n 0.0181522f $X=-0.19 $Y=-0.245 $X2=6.3 $Y2=1.32
cc_66 VNB N_VGND_c_1253_n 0.00638216f $X=-0.19 $Y=-0.245 $X2=6.615 $Y2=1.765
cc_67 VNB N_VGND_c_1254_n 0.0151544f $X=-0.19 $Y=-0.245 $X2=6.73 $Y2=0.74
cc_68 VNB N_VGND_c_1255_n 0.0190588f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_1256_n 0.0178645f $X=-0.19 $Y=-0.245 $X2=7.16 $Y2=1.32
cc_70 VNB N_VGND_c_1257_n 0.0026136f $X=-0.19 $Y=-0.245 $X2=7.515 $Y2=1.765
cc_71 VNB N_VGND_c_1258_n 0.002601f $X=-0.19 $Y=-0.245 $X2=7.59 $Y2=0.74
cc_72 VNB N_VGND_c_1259_n 0.00558127f $X=-0.19 $Y=-0.245 $X2=3.24 $Y2=1.57
cc_73 VNB N_VGND_c_1260_n 0.0142878f $X=-0.19 $Y=-0.245 $X2=3.24 $Y2=1.57
cc_74 VNB N_VGND_c_1261_n 0.029743f $X=-0.19 $Y=-0.245 $X2=4.115 $Y2=1.405
cc_75 VNB N_VGND_c_1262_n 0.0183144f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1263_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=4.955 $Y2=1.907
cc_77 VNB N_VGND_c_1264_n 0.0172883f $X=-0.19 $Y=-0.245 $X2=5.88 $Y2=1.985
cc_78 VNB N_VGND_c_1265_n 0.00332923f $X=-0.19 $Y=-0.245 $X2=5.12 $Y2=1.985
cc_79 VNB N_VGND_c_1266_n 0.016486f $X=-0.19 $Y=-0.245 $X2=5.12 $Y2=1.985
cc_80 VNB N_VGND_c_1267_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=5.965 $Y2=1.65
cc_81 VNB N_VGND_c_1268_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=6.05 $Y2=1.485
cc_82 VNB N_VGND_c_1269_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=6.11 $Y2=1.485
cc_83 VNB N_VGND_c_1270_n 0.0807918f $X=-0.19 $Y=-0.245 $X2=4.065 $Y2=1.91
cc_84 VNB N_VGND_c_1271_n 0.0172524f $X=-0.19 $Y=-0.245 $X2=6.11 $Y2=1.542
cc_85 VNB N_VGND_c_1272_n 0.018855f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1273_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1274_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1275_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1276_n 0.527831f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_707_119#_c_1378_n 0.0130452f $X=-0.19 $Y=-0.245 $X2=2.25 $Y2=0.945
cc_91 VNB N_A_707_119#_c_1379_n 0.0106798f $X=-0.19 $Y=-0.245 $X2=2.325
+ $Y2=1.415
cc_92 VNB N_A_707_119#_c_1380_n 0.00422464f $X=-0.19 $Y=-0.245 $X2=2.72 $Y2=1.34
cc_93 VNB N_A_707_119#_c_1381_n 0.00269685f $X=-0.19 $Y=-0.245 $X2=2.865
+ $Y2=2.315
cc_94 VNB N_A_707_119#_c_1382_n 0.00636128f $X=-0.19 $Y=-0.245 $X2=2.865
+ $Y2=2.315
cc_95 VNB N_A_707_119#_c_1383_n 0.00152462f $X=-0.19 $Y=-0.245 $X2=3.315
+ $Y2=1.82
cc_96 VNB N_A_707_119#_c_1384_n 0.0140492f $X=-0.19 $Y=-0.245 $X2=6.005
+ $Y2=1.765
cc_97 VPB N_A_435_99#_c_207_n 0.0131129f $X=-0.19 $Y=1.66 $X2=2.865 $Y2=1.82
cc_98 VPB N_A_435_99#_c_208_n 0.0126735f $X=-0.19 $Y=1.66 $X2=3.315 $Y2=1.82
cc_99 VPB N_A_435_99#_c_209_n 0.0182588f $X=-0.19 $Y=1.66 $X2=6.005 $Y2=1.765
cc_100 VPB N_A_435_99#_c_210_n 0.0160176f $X=-0.19 $Y=1.66 $X2=6.615 $Y2=1.765
cc_101 VPB N_A_435_99#_c_211_n 0.0148707f $X=-0.19 $Y=1.66 $X2=7.065 $Y2=1.765
cc_102 VPB N_A_435_99#_c_212_n 0.014865f $X=-0.19 $Y=1.66 $X2=7.515 $Y2=1.765
cc_103 VPB N_A_435_99#_c_203_n 0.00428654f $X=-0.19 $Y=1.66 $X2=3.9 $Y2=1.57
cc_104 VPB N_A_435_99#_c_204_n 0.0255457f $X=-0.19 $Y=1.66 $X2=3.24 $Y2=1.57
cc_105 VPB N_A_435_99#_c_215_n 0.0103055f $X=-0.19 $Y=1.66 $X2=5.88 $Y2=1.985
cc_106 VPB N_A_435_99#_c_216_n 0.00169914f $X=-0.19 $Y=1.66 $X2=5.12 $Y2=1.985
cc_107 VPB N_A_435_99#_c_217_n 0.00194892f $X=-0.19 $Y=1.66 $X2=5.965 $Y2=1.82
cc_108 VPB N_A_435_99#_c_218_n 0.00391539f $X=-0.19 $Y=1.66 $X2=4.07 $Y2=1.907
cc_109 VPB N_A_435_99#_c_219_n 0.0111012f $X=-0.19 $Y=1.66 $X2=4.955 $Y2=1.985
cc_110 VPB N_A_435_99#_c_206_n 0.0268975f $X=-0.19 $Y=1.66 $X2=7.515 $Y2=1.542
cc_111 VPB N_B_c_395_n 0.0148248f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_B_c_396_n 0.0150115f $X=-0.19 $Y=1.66 $X2=2.25 $Y2=0.945
cc_113 VPB N_B_c_397_n 0.0292803f $X=-0.19 $Y=1.66 $X2=2.72 $Y2=1.34
cc_114 VPB N_B_c_389_n 0.0295206f $X=-0.19 $Y=1.66 $X2=2.72 $Y2=0.945
cc_115 VPB N_B_c_399_n 0.0670697f $X=-0.19 $Y=1.66 $X2=2.865 $Y2=1.82
cc_116 VPB N_B_c_400_n 0.0906391f $X=-0.19 $Y=1.66 $X2=2.865 $Y2=2.315
cc_117 VPB N_B_c_401_n 0.0123718f $X=-0.19 $Y=1.66 $X2=2.865 $Y2=2.315
cc_118 VPB N_B_c_402_n 0.00645803f $X=-0.19 $Y=1.66 $X2=3.315 $Y2=1.82
cc_119 VPB N_B_c_403_n 0.0122415f $X=-0.19 $Y=1.66 $X2=3.315 $Y2=2.315
cc_120 VPB N_B_c_390_n 0.0168261f $X=-0.19 $Y=1.66 $X2=3.315 $Y2=2.315
cc_121 VPB N_B_M1012_g 0.00820227f $X=-0.19 $Y=1.66 $X2=6.005 $Y2=2.4
cc_122 VPB N_B_c_406_n 0.0344138f $X=-0.19 $Y=1.66 $X2=6.615 $Y2=1.765
cc_123 VPB N_B_c_392_n 0.0159362f $X=-0.19 $Y=1.66 $X2=6.615 $Y2=2.4
cc_124 VPB N_B_c_408_n 0.0132794f $X=-0.19 $Y=1.66 $X2=7.065 $Y2=2.4
cc_125 VPB N_B_c_409_n 0.00879521f $X=-0.19 $Y=1.66 $X2=7.16 $Y2=0.74
cc_126 VPB N_B_c_410_n 0.0208791f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_127 VPB B 5.62692e-19 $X=-0.19 $Y=1.66 $X2=7.515 $Y2=2.4
cc_128 VPB N_A_c_534_n 0.0205427f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_129 VPB N_A_c_535_n 0.0151861f $X=-0.19 $Y=1.66 $X2=2.25 $Y2=0.945
cc_130 VPB N_A_c_526_n 0.0166576f $X=-0.19 $Y=1.66 $X2=2.865 $Y2=1.82
cc_131 VPB N_A_c_537_n 0.0216036f $X=-0.19 $Y=1.66 $X2=2.865 $Y2=2.315
cc_132 VPB N_A_c_538_n 0.0172736f $X=-0.19 $Y=1.66 $X2=6.615 $Y2=1.765
cc_133 VPB N_A_c_530_n 0.00127149f $X=-0.19 $Y=1.66 $X2=6.73 $Y2=1.32
cc_134 VPB N_A_c_531_n 0.00753631f $X=-0.19 $Y=1.66 $X2=6.73 $Y2=0.74
cc_135 VPB A 0.012236f $X=-0.19 $Y=1.66 $X2=7.065 $Y2=1.765
cc_136 VPB N_A_c_533_n 0.0353964f $X=-0.19 $Y=1.66 $X2=7.515 $Y2=2.4
cc_137 VPB N_A_294_392#_c_651_n 0.0147853f $X=-0.19 $Y=1.66 $X2=2.25 $Y2=1.34
cc_138 VPB N_A_294_392#_c_652_n 0.0148986f $X=-0.19 $Y=1.66 $X2=2.72 $Y2=0.945
cc_139 VPB N_A_294_392#_c_653_n 0.0166512f $X=-0.19 $Y=1.66 $X2=6.005 $Y2=1.765
cc_140 VPB N_A_294_392#_c_644_n 0.0200339f $X=-0.19 $Y=1.66 $X2=6.615 $Y2=2.4
cc_141 VPB N_A_294_392#_c_655_n 0.0189879f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_142 VPB N_A_294_392#_c_656_n 0.0067261f $X=-0.19 $Y=1.66 $X2=7.16 $Y2=0.74
cc_143 VPB N_A_294_392#_c_647_n 0.00462276f $X=-0.19 $Y=1.66 $X2=7.59 $Y2=0.74
cc_144 VPB N_A_294_392#_c_658_n 0.00105625f $X=-0.19 $Y=1.66 $X2=4.115 $Y2=1.405
cc_145 VPB N_A_294_392#_c_649_n 0.00786705f $X=-0.19 $Y=1.66 $X2=5.12 $Y2=1.985
cc_146 VPB N_A_294_392#_c_660_n 0.00194632f $X=-0.19 $Y=1.66 $X2=5.965 $Y2=1.65
cc_147 VPB N_A_294_392#_c_661_n 5.40493e-19 $X=-0.19 $Y=1.66 $X2=6.05 $Y2=1.485
cc_148 VPB N_A_27_392#_c_845_n 0.0101511f $X=-0.19 $Y=1.66 $X2=2.25 $Y2=1.34
cc_149 VPB N_A_27_392#_c_846_n 0.0340353f $X=-0.19 $Y=1.66 $X2=2.25 $Y2=0.945
cc_150 VPB N_A_27_392#_c_847_n 0.0020579f $X=-0.19 $Y=1.66 $X2=2.325 $Y2=1.415
cc_151 VPB N_A_27_392#_c_848_n 0.00220677f $X=-0.19 $Y=1.66 $X2=2.72 $Y2=0.945
cc_152 VPB N_A_27_392#_c_849_n 0.00664265f $X=-0.19 $Y=1.66 $X2=2.865 $Y2=2.315
cc_153 VPB N_A_27_392#_c_850_n 0.00171072f $X=-0.19 $Y=1.66 $X2=3.315 $Y2=1.82
cc_154 VPB N_A_27_392#_c_851_n 0.00518526f $X=-0.19 $Y=1.66 $X2=6.005 $Y2=1.765
cc_155 VPB N_VPWR_c_890_n 0.00538125f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_156 VPB N_VPWR_c_891_n 0.00907658f $X=-0.19 $Y=1.66 $X2=6.73 $Y2=1.32
cc_157 VPB N_VPWR_c_892_n 0.00328505f $X=-0.19 $Y=1.66 $X2=7.065 $Y2=1.765
cc_158 VPB N_VPWR_c_893_n 0.00490739f $X=-0.19 $Y=1.66 $X2=7.16 $Y2=0.74
cc_159 VPB N_VPWR_c_894_n 0.0231664f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_160 VPB N_VPWR_c_895_n 0.0141169f $X=-0.19 $Y=1.66 $X2=7.59 $Y2=1.32
cc_161 VPB N_VPWR_c_896_n 0.00329129f $X=-0.19 $Y=1.66 $X2=3.9 $Y2=1.57
cc_162 VPB N_VPWR_c_897_n 0.00261791f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_163 VPB N_VPWR_c_898_n 0.00329129f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_164 VPB N_VPWR_c_899_n 0.0120106f $X=-0.19 $Y=1.66 $X2=4.23 $Y2=1.907
cc_165 VPB N_VPWR_c_900_n 0.0345413f $X=-0.19 $Y=1.66 $X2=5.12 $Y2=1.985
cc_166 VPB N_VPWR_c_901_n 0.0228504f $X=-0.19 $Y=1.66 $X2=5.965 $Y2=1.65
cc_167 VPB N_VPWR_c_902_n 0.00601644f $X=-0.19 $Y=1.66 $X2=5.965 $Y2=1.82
cc_168 VPB N_VPWR_c_903_n 0.0177589f $X=-0.19 $Y=1.66 $X2=6.11 $Y2=1.485
cc_169 VPB N_VPWR_c_904_n 0.00601644f $X=-0.19 $Y=1.66 $X2=6.11 $Y2=1.485
cc_170 VPB N_VPWR_c_905_n 0.0159778f $X=-0.19 $Y=1.66 $X2=6.79 $Y2=1.485
cc_171 VPB N_VPWR_c_906_n 0.00601644f $X=-0.19 $Y=1.66 $X2=6.79 $Y2=1.485
cc_172 VPB N_VPWR_c_907_n 0.0175377f $X=-0.19 $Y=1.66 $X2=4.07 $Y2=1.57
cc_173 VPB N_VPWR_c_908_n 0.0400678f $X=-0.19 $Y=1.66 $X2=2.72 $Y2=1.34
cc_174 VPB N_VPWR_c_909_n 0.0159813f $X=-0.19 $Y=1.66 $X2=6.73 $Y2=1.542
cc_175 VPB N_VPWR_c_910_n 0.0209137f $X=-0.19 $Y=1.66 $X2=7.59 $Y2=1.542
cc_176 VPB N_VPWR_c_911_n 0.0234703f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_177 VPB N_VPWR_c_912_n 0.00460249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_178 VPB N_VPWR_c_913_n 0.00436868f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_179 VPB N_VPWR_c_914_n 0.00436868f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_180 VPB N_VPWR_c_915_n 0.00507883f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_181 VPB N_VPWR_c_916_n 0.00854561f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_182 VPB N_VPWR_c_889_n 0.0970882f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_183 VPB N_COUT_c_1049_n 0.00478236f $X=-0.19 $Y=1.66 $X2=2.645 $Y2=1.415
cc_184 VPB COUT 0.00157739f $X=-0.19 $Y=1.66 $X2=6.3 $Y2=0.74
cc_185 VPB N_SUM_c_1104_n 0.00155998f $X=-0.19 $Y=1.66 $X2=2.645 $Y2=1.415
cc_186 VPB N_SUM_c_1105_n 0.00233217f $X=-0.19 $Y=1.66 $X2=2.72 $Y2=1.34
cc_187 VPB N_SUM_c_1106_n 0.00332586f $X=-0.19 $Y=1.66 $X2=6.3 $Y2=0.74
cc_188 VPB N_SUM_c_1107_n 0.00273983f $X=-0.19 $Y=1.66 $X2=6.615 $Y2=2.4
cc_189 VPB N_SUM_c_1102_n 0.0227863f $X=-0.19 $Y=1.66 $X2=6.73 $Y2=0.74
cc_190 VPB N_SUM_c_1109_n 0.00280642f $X=-0.19 $Y=1.66 $X2=7.16 $Y2=1.32
cc_191 VPB N_SUM_c_1110_n 0.0021075f $X=-0.19 $Y=1.66 $X2=7.16 $Y2=0.74
cc_192 VPB SUM 9.18137e-19 $X=-0.19 $Y=1.66 $X2=7.59 $Y2=0.74
cc_193 VPB N_A_707_119#_c_1383_n 0.00305102f $X=-0.19 $Y=1.66 $X2=3.315 $Y2=1.82
cc_194 N_A_435_99#_c_195_n N_B_M1004_g 0.0131498f $X=2.25 $Y=1.34 $X2=0 $Y2=0
cc_195 N_A_435_99#_c_197_n N_B_c_397_n 0.0155157f $X=2.325 $Y=1.415 $X2=0 $Y2=0
cc_196 N_A_435_99#_c_207_n N_B_c_397_n 0.0261776f $X=2.865 $Y=1.82 $X2=0 $Y2=0
cc_197 N_A_435_99#_c_204_n N_B_c_397_n 0.00269064f $X=3.24 $Y=1.57 $X2=0 $Y2=0
cc_198 N_A_435_99#_c_197_n N_B_c_389_n 0.00195768f $X=2.325 $Y=1.415 $X2=0 $Y2=0
cc_199 N_A_435_99#_c_207_n N_B_c_400_n 0.0103562f $X=2.865 $Y=1.82 $X2=0 $Y2=0
cc_200 N_A_435_99#_c_208_n N_B_c_400_n 0.0103562f $X=3.315 $Y=1.82 $X2=0 $Y2=0
cc_201 N_A_435_99#_c_208_n N_B_c_402_n 0.00242326f $X=3.315 $Y=1.82 $X2=0 $Y2=0
cc_202 N_A_435_99#_c_203_n N_B_c_390_n 0.0147823f $X=3.9 $Y=1.57 $X2=0 $Y2=0
cc_203 N_A_435_99#_c_204_n N_B_c_390_n 0.0140234f $X=3.24 $Y=1.57 $X2=0 $Y2=0
cc_204 N_A_435_99#_c_218_n N_B_c_390_n 0.00630158f $X=4.07 $Y=1.907 $X2=0 $Y2=0
cc_205 N_A_435_99#_c_208_n N_B_M1012_g 0.0269826f $X=3.315 $Y=1.82 $X2=0 $Y2=0
cc_206 N_A_435_99#_c_218_n N_B_M1012_g 0.0057445f $X=4.07 $Y=1.907 $X2=0 $Y2=0
cc_207 N_A_435_99#_c_203_n N_B_M1001_g 0.00633468f $X=3.9 $Y=1.57 $X2=0 $Y2=0
cc_208 N_A_435_99#_c_204_n N_B_M1001_g 0.00541031f $X=3.24 $Y=1.57 $X2=0 $Y2=0
cc_209 N_A_435_99#_c_236_p N_B_M1001_g 0.0143629f $X=4.115 $Y=0.74 $X2=0 $Y2=0
cc_210 N_A_435_99#_c_218_n N_B_M1001_g 0.00491066f $X=4.07 $Y=1.907 $X2=0 $Y2=0
cc_211 N_A_435_99#_c_218_n N_B_c_392_n 0.0138324f $X=4.07 $Y=1.907 $X2=0 $Y2=0
cc_212 N_A_435_99#_c_219_n N_B_c_392_n 0.00449678f $X=4.955 $Y=1.985 $X2=0 $Y2=0
cc_213 N_A_435_99#_c_236_p N_B_M1035_g 0.00998427f $X=4.115 $Y=0.74 $X2=0 $Y2=0
cc_214 N_A_435_99#_c_218_n N_B_M1035_g 0.00276031f $X=4.07 $Y=1.907 $X2=0 $Y2=0
cc_215 N_A_435_99#_c_219_n N_B_c_408_n 0.00718914f $X=4.955 $Y=1.985 $X2=0 $Y2=0
cc_216 N_A_435_99#_c_197_n B 0.00706672f $X=2.325 $Y=1.415 $X2=0 $Y2=0
cc_217 N_A_435_99#_c_195_n N_A_c_524_n 0.00737233f $X=2.25 $Y=1.34 $X2=0 $Y2=0
cc_218 N_A_435_99#_c_198_n N_A_c_524_n 0.00737233f $X=2.72 $Y=1.34 $X2=0 $Y2=0
cc_219 N_A_435_99#_c_218_n N_A_c_526_n 0.00238841f $X=4.07 $Y=1.907 $X2=0 $Y2=0
cc_220 N_A_435_99#_c_219_n N_A_c_526_n 0.00637087f $X=4.955 $Y=1.985 $X2=0 $Y2=0
cc_221 N_A_435_99#_c_216_n N_A_c_537_n 0.00502767f $X=5.12 $Y=1.985 $X2=0 $Y2=0
cc_222 N_A_435_99#_c_219_n N_A_c_537_n 0.00843733f $X=4.955 $Y=1.985 $X2=0 $Y2=0
cc_223 N_A_435_99#_c_236_p N_A_M1002_g 2.53475e-19 $X=4.115 $Y=0.74 $X2=0 $Y2=0
cc_224 N_A_435_99#_c_219_n N_A_c_528_n 0.00850337f $X=4.955 $Y=1.985 $X2=0 $Y2=0
cc_225 N_A_435_99#_c_209_n N_A_c_538_n 0.0227273f $X=6.005 $Y=1.765 $X2=0 $Y2=0
cc_226 N_A_435_99#_c_215_n N_A_c_538_n 0.0152441f $X=5.88 $Y=1.985 $X2=0 $Y2=0
cc_227 N_A_435_99#_c_217_n N_A_c_538_n 8.70491e-19 $X=5.965 $Y=1.82 $X2=0 $Y2=0
cc_228 N_A_435_99#_c_218_n N_A_c_530_n 3.08349e-19 $X=4.07 $Y=1.907 $X2=0 $Y2=0
cc_229 N_A_435_99#_c_215_n N_A_c_531_n 8.73915e-19 $X=5.88 $Y=1.985 $X2=0 $Y2=0
cc_230 N_A_435_99#_c_217_n N_A_c_531_n 0.00186939f $X=5.965 $Y=1.82 $X2=0 $Y2=0
cc_231 N_A_435_99#_c_205_n N_A_c_531_n 0.00183083f $X=6.05 $Y=1.485 $X2=0 $Y2=0
cc_232 N_A_435_99#_c_206_n N_A_c_531_n 0.00860065f $X=7.515 $Y=1.542 $X2=0 $Y2=0
cc_233 N_A_435_99#_c_212_n N_A_294_392#_c_651_n 0.0368241f $X=7.515 $Y=1.765
+ $X2=0 $Y2=0
cc_234 N_A_435_99#_M1030_g N_A_294_392#_M1003_g 0.0317962f $X=7.59 $Y=0.74 $X2=0
+ $Y2=0
cc_235 N_A_435_99#_c_206_n N_A_294_392#_c_644_n 0.0233467f $X=7.515 $Y=1.542
+ $X2=0 $Y2=0
cc_236 N_A_435_99#_c_196_n N_A_294_392#_c_656_n 0.00116202f $X=2.645 $Y=1.415
+ $X2=0 $Y2=0
cc_237 N_A_435_99#_c_197_n N_A_294_392#_c_656_n 5.73178e-19 $X=2.325 $Y=1.415
+ $X2=0 $Y2=0
cc_238 N_A_435_99#_c_195_n N_A_294_392#_c_646_n 3.39182e-19 $X=2.25 $Y=1.34
+ $X2=0 $Y2=0
cc_239 N_A_435_99#_c_198_n N_A_294_392#_c_646_n 0.00586917f $X=2.72 $Y=1.34
+ $X2=0 $Y2=0
cc_240 N_A_435_99#_c_195_n N_A_294_392#_c_647_n 0.00113236f $X=2.25 $Y=1.34
+ $X2=0 $Y2=0
cc_241 N_A_435_99#_c_196_n N_A_294_392#_c_647_n 0.00939344f $X=2.645 $Y=1.415
+ $X2=0 $Y2=0
cc_242 N_A_435_99#_c_198_n N_A_294_392#_c_647_n 0.00257225f $X=2.72 $Y=1.34
+ $X2=0 $Y2=0
cc_243 N_A_435_99#_c_207_n N_A_294_392#_c_647_n 0.00192352f $X=2.865 $Y=1.82
+ $X2=0 $Y2=0
cc_244 N_A_435_99#_c_203_n N_A_294_392#_c_647_n 0.0132865f $X=3.9 $Y=1.57 $X2=0
+ $Y2=0
cc_245 N_A_435_99#_c_204_n N_A_294_392#_c_647_n 0.0150559f $X=3.24 $Y=1.57 $X2=0
+ $Y2=0
cc_246 N_A_435_99#_c_207_n N_A_294_392#_c_675_n 0.0158814f $X=2.865 $Y=1.82
+ $X2=0 $Y2=0
cc_247 N_A_435_99#_c_204_n N_A_294_392#_c_675_n 0.00283903f $X=3.24 $Y=1.57
+ $X2=0 $Y2=0
cc_248 N_A_435_99#_M1012_s N_A_294_392#_c_677_n 4.38684e-19 $X=3.84 $Y=1.895
+ $X2=0 $Y2=0
cc_249 N_A_435_99#_c_208_n N_A_294_392#_c_677_n 0.0124791f $X=3.315 $Y=1.82
+ $X2=0 $Y2=0
cc_250 N_A_435_99#_c_203_n N_A_294_392#_c_677_n 0.0207441f $X=3.9 $Y=1.57 $X2=0
+ $Y2=0
cc_251 N_A_435_99#_M1012_s N_A_294_392#_c_680_n 0.004488f $X=3.84 $Y=1.895 $X2=0
+ $Y2=0
cc_252 N_A_435_99#_M1018_s N_A_294_392#_c_680_n 0.00789233f $X=4.895 $Y=2.05
+ $X2=0 $Y2=0
cc_253 N_A_435_99#_c_209_n N_A_294_392#_c_680_n 0.0140661f $X=6.005 $Y=1.765
+ $X2=0 $Y2=0
cc_254 N_A_435_99#_c_210_n N_A_294_392#_c_680_n 0.012771f $X=6.615 $Y=1.765
+ $X2=0 $Y2=0
cc_255 N_A_435_99#_c_211_n N_A_294_392#_c_680_n 0.0120114f $X=7.065 $Y=1.765
+ $X2=0 $Y2=0
cc_256 N_A_435_99#_c_212_n N_A_294_392#_c_680_n 0.0130109f $X=7.515 $Y=1.765
+ $X2=0 $Y2=0
cc_257 N_A_435_99#_c_215_n N_A_294_392#_c_680_n 0.00909891f $X=5.88 $Y=1.985
+ $X2=0 $Y2=0
cc_258 N_A_435_99#_c_216_n N_A_294_392#_c_680_n 0.0606142f $X=5.12 $Y=1.985
+ $X2=0 $Y2=0
cc_259 N_A_435_99#_c_286_p N_A_294_392#_c_680_n 0.0034106f $X=6.79 $Y=1.485
+ $X2=0 $Y2=0
cc_260 N_A_435_99#_c_218_n N_A_294_392#_c_680_n 0.00749389f $X=4.07 $Y=1.907
+ $X2=0 $Y2=0
cc_261 N_A_435_99#_c_219_n N_A_294_392#_c_680_n 0.0267874f $X=4.955 $Y=1.985
+ $X2=0 $Y2=0
cc_262 N_A_435_99#_c_206_n N_A_294_392#_c_680_n 0.00255078f $X=7.515 $Y=1.542
+ $X2=0 $Y2=0
cc_263 N_A_435_99#_c_212_n N_A_294_392#_c_658_n 0.00605309f $X=7.515 $Y=1.765
+ $X2=0 $Y2=0
cc_264 N_A_435_99#_c_206_n N_A_294_392#_c_658_n 7.04585e-19 $X=7.515 $Y=1.542
+ $X2=0 $Y2=0
cc_265 N_A_435_99#_c_206_n N_A_294_392#_c_648_n 0.00279232f $X=7.515 $Y=1.542
+ $X2=0 $Y2=0
cc_266 N_A_435_99#_c_196_n N_A_294_392#_c_650_n 0.00266209f $X=2.645 $Y=1.415
+ $X2=0 $Y2=0
cc_267 N_A_435_99#_c_198_n N_A_294_392#_c_650_n 0.00361003f $X=2.72 $Y=1.34
+ $X2=0 $Y2=0
cc_268 N_A_435_99#_c_207_n N_A_294_392#_c_697_n 0.00622518f $X=2.865 $Y=1.82
+ $X2=0 $Y2=0
cc_269 N_A_435_99#_c_208_n N_A_294_392#_c_697_n 0.00660312f $X=3.315 $Y=1.82
+ $X2=0 $Y2=0
cc_270 N_A_435_99#_c_203_n N_A_294_392#_c_697_n 0.0118485f $X=3.9 $Y=1.57 $X2=0
+ $Y2=0
cc_271 N_A_435_99#_c_204_n N_A_294_392#_c_697_n 0.00663437f $X=3.24 $Y=1.57
+ $X2=0 $Y2=0
cc_272 N_A_435_99#_c_218_n N_A_294_392#_c_697_n 0.00271011f $X=4.07 $Y=1.907
+ $X2=0 $Y2=0
cc_273 N_A_435_99#_M1012_s N_A_294_392#_c_702_n 0.008482f $X=3.84 $Y=1.895 $X2=0
+ $Y2=0
cc_274 N_A_435_99#_c_218_n N_A_294_392#_c_702_n 0.0143157f $X=4.07 $Y=1.907
+ $X2=0 $Y2=0
cc_275 N_A_435_99#_c_215_n N_VPWR_M1019_d 0.00678518f $X=5.88 $Y=1.985 $X2=0
+ $Y2=0
cc_276 N_A_435_99#_c_207_n N_VPWR_c_891_n 0.0100709f $X=2.865 $Y=1.82 $X2=0
+ $Y2=0
cc_277 N_A_435_99#_c_208_n N_VPWR_c_891_n 0.00153805f $X=3.315 $Y=1.82 $X2=0
+ $Y2=0
cc_278 N_A_435_99#_c_207_n N_VPWR_c_892_n 0.00106331f $X=2.865 $Y=1.82 $X2=0
+ $Y2=0
cc_279 N_A_435_99#_c_208_n N_VPWR_c_892_n 0.00820156f $X=3.315 $Y=1.82 $X2=0
+ $Y2=0
cc_280 N_A_435_99#_c_209_n N_VPWR_c_895_n 0.018159f $X=6.005 $Y=1.765 $X2=0
+ $Y2=0
cc_281 N_A_435_99#_c_210_n N_VPWR_c_895_n 0.00189143f $X=6.615 $Y=1.765 $X2=0
+ $Y2=0
cc_282 N_A_435_99#_c_209_n N_VPWR_c_896_n 0.00189741f $X=6.005 $Y=1.765 $X2=0
+ $Y2=0
cc_283 N_A_435_99#_c_210_n N_VPWR_c_896_n 0.0108226f $X=6.615 $Y=1.765 $X2=0
+ $Y2=0
cc_284 N_A_435_99#_c_211_n N_VPWR_c_896_n 0.00963065f $X=7.065 $Y=1.765 $X2=0
+ $Y2=0
cc_285 N_A_435_99#_c_212_n N_VPWR_c_896_n 0.00127141f $X=7.515 $Y=1.765 $X2=0
+ $Y2=0
cc_286 N_A_435_99#_c_211_n N_VPWR_c_897_n 0.00127141f $X=7.065 $Y=1.765 $X2=0
+ $Y2=0
cc_287 N_A_435_99#_c_212_n N_VPWR_c_897_n 0.00959143f $X=7.515 $Y=1.765 $X2=0
+ $Y2=0
cc_288 N_A_435_99#_c_209_n N_VPWR_c_901_n 0.00413917f $X=6.005 $Y=1.765 $X2=0
+ $Y2=0
cc_289 N_A_435_99#_c_210_n N_VPWR_c_901_n 0.00413917f $X=6.615 $Y=1.765 $X2=0
+ $Y2=0
cc_290 N_A_435_99#_c_211_n N_VPWR_c_903_n 0.00413917f $X=7.065 $Y=1.765 $X2=0
+ $Y2=0
cc_291 N_A_435_99#_c_212_n N_VPWR_c_903_n 0.00413917f $X=7.515 $Y=1.765 $X2=0
+ $Y2=0
cc_292 N_A_435_99#_c_207_n N_VPWR_c_889_n 8.51577e-19 $X=2.865 $Y=1.82 $X2=0
+ $Y2=0
cc_293 N_A_435_99#_c_208_n N_VPWR_c_889_n 8.51577e-19 $X=3.315 $Y=1.82 $X2=0
+ $Y2=0
cc_294 N_A_435_99#_c_209_n N_VPWR_c_889_n 0.00415837f $X=6.005 $Y=1.765 $X2=0
+ $Y2=0
cc_295 N_A_435_99#_c_210_n N_VPWR_c_889_n 0.00415837f $X=6.615 $Y=1.765 $X2=0
+ $Y2=0
cc_296 N_A_435_99#_c_211_n N_VPWR_c_889_n 0.00414505f $X=7.065 $Y=1.765 $X2=0
+ $Y2=0
cc_297 N_A_435_99#_c_212_n N_VPWR_c_889_n 0.00414505f $X=7.515 $Y=1.765 $X2=0
+ $Y2=0
cc_298 N_A_435_99#_c_209_n N_COUT_c_1049_n 0.00284052f $X=6.005 $Y=1.765 $X2=0
+ $Y2=0
cc_299 N_A_435_99#_c_210_n N_COUT_c_1049_n 0.0132246f $X=6.615 $Y=1.765 $X2=0
+ $Y2=0
cc_300 N_A_435_99#_c_211_n N_COUT_c_1049_n 0.0182321f $X=7.065 $Y=1.765 $X2=0
+ $Y2=0
cc_301 N_A_435_99#_c_215_n N_COUT_c_1049_n 0.0287017f $X=5.88 $Y=1.985 $X2=0
+ $Y2=0
cc_302 N_A_435_99#_c_286_p N_COUT_c_1049_n 0.057553f $X=6.79 $Y=1.485 $X2=0
+ $Y2=0
cc_303 N_A_435_99#_c_206_n N_COUT_c_1049_n 0.0199091f $X=7.515 $Y=1.542 $X2=0
+ $Y2=0
cc_304 N_A_435_99#_M1006_g N_COUT_c_1046_n 0.00335135f $X=6.3 $Y=0.74 $X2=0
+ $Y2=0
cc_305 N_A_435_99#_c_286_p N_COUT_c_1046_n 0.0192803f $X=6.79 $Y=1.485 $X2=0
+ $Y2=0
cc_306 N_A_435_99#_c_206_n N_COUT_c_1046_n 0.00242376f $X=7.515 $Y=1.542 $X2=0
+ $Y2=0
cc_307 N_A_435_99#_M1006_g N_COUT_c_1047_n 0.0067313f $X=6.3 $Y=0.74 $X2=0 $Y2=0
cc_308 N_A_435_99#_M1010_g N_COUT_c_1047_n 3.97481e-19 $X=6.73 $Y=0.74 $X2=0
+ $Y2=0
cc_309 N_A_435_99#_M1010_g N_COUT_c_1048_n 0.0147737f $X=6.73 $Y=0.74 $X2=0
+ $Y2=0
cc_310 N_A_435_99#_M1028_g N_COUT_c_1048_n 0.0162215f $X=7.16 $Y=0.74 $X2=0
+ $Y2=0
cc_311 N_A_435_99#_c_286_p N_COUT_c_1048_n 0.024649f $X=6.79 $Y=1.485 $X2=0
+ $Y2=0
cc_312 N_A_435_99#_c_206_n N_COUT_c_1048_n 0.00291477f $X=7.515 $Y=1.542 $X2=0
+ $Y2=0
cc_313 N_A_435_99#_M1028_g N_COUT_c_1066_n 0.001989f $X=7.16 $Y=0.74 $X2=0 $Y2=0
cc_314 N_A_435_99#_M1030_g N_COUT_c_1066_n 0.00705268f $X=7.59 $Y=0.74 $X2=0
+ $Y2=0
cc_315 N_A_435_99#_M1010_g COUT 9.18327e-19 $X=6.73 $Y=0.74 $X2=0 $Y2=0
cc_316 N_A_435_99#_c_211_n COUT 0.00146285f $X=7.065 $Y=1.765 $X2=0 $Y2=0
cc_317 N_A_435_99#_M1028_g COUT 0.00571358f $X=7.16 $Y=0.74 $X2=0 $Y2=0
cc_318 N_A_435_99#_c_212_n COUT 0.00136726f $X=7.515 $Y=1.765 $X2=0 $Y2=0
cc_319 N_A_435_99#_M1030_g COUT 0.005924f $X=7.59 $Y=0.74 $X2=0 $Y2=0
cc_320 N_A_435_99#_c_286_p COUT 0.0189686f $X=6.79 $Y=1.485 $X2=0 $Y2=0
cc_321 N_A_435_99#_c_206_n COUT 0.0321032f $X=7.515 $Y=1.542 $X2=0 $Y2=0
cc_322 N_A_435_99#_c_212_n N_COUT_c_1075_n 0.00720355f $X=7.515 $Y=1.765 $X2=0
+ $Y2=0
cc_323 N_A_435_99#_c_195_n N_A_27_125#_c_1191_n 0.00197658f $X=2.25 $Y=1.34
+ $X2=0 $Y2=0
cc_324 N_A_435_99#_c_195_n N_A_27_125#_c_1192_n 0.00371137f $X=2.25 $Y=1.34
+ $X2=0 $Y2=0
cc_325 N_A_435_99#_c_198_n N_A_27_125#_c_1192_n 0.00330783f $X=2.72 $Y=1.34
+ $X2=0 $Y2=0
cc_326 N_A_435_99#_c_198_n N_A_27_125#_c_1194_n 0.0155464f $X=2.72 $Y=1.34 $X2=0
+ $Y2=0
cc_327 N_A_435_99#_c_203_n N_A_27_125#_c_1194_n 0.00783057f $X=3.9 $Y=1.57 $X2=0
+ $Y2=0
cc_328 N_A_435_99#_c_204_n N_A_27_125#_c_1194_n 0.0105914f $X=3.24 $Y=1.57 $X2=0
+ $Y2=0
cc_329 N_A_435_99#_M1006_g N_VGND_c_1256_n 0.00511131f $X=6.3 $Y=0.74 $X2=0
+ $Y2=0
cc_330 N_A_435_99#_c_205_n N_VGND_c_1256_n 0.010681f $X=6.05 $Y=1.485 $X2=0
+ $Y2=0
cc_331 N_A_435_99#_c_286_p N_VGND_c_1256_n 0.00919629f $X=6.79 $Y=1.485 $X2=0
+ $Y2=0
cc_332 N_A_435_99#_c_206_n N_VGND_c_1256_n 0.00381579f $X=7.515 $Y=1.542 $X2=0
+ $Y2=0
cc_333 N_A_435_99#_M1006_g N_VGND_c_1257_n 4.53155e-19 $X=6.3 $Y=0.74 $X2=0
+ $Y2=0
cc_334 N_A_435_99#_M1010_g N_VGND_c_1257_n 0.00813302f $X=6.73 $Y=0.74 $X2=0
+ $Y2=0
cc_335 N_A_435_99#_M1028_g N_VGND_c_1257_n 0.0105568f $X=7.16 $Y=0.74 $X2=0
+ $Y2=0
cc_336 N_A_435_99#_M1030_g N_VGND_c_1257_n 0.00138519f $X=7.59 $Y=0.74 $X2=0
+ $Y2=0
cc_337 N_A_435_99#_M1028_g N_VGND_c_1258_n 0.00138519f $X=7.16 $Y=0.74 $X2=0
+ $Y2=0
cc_338 N_A_435_99#_M1030_g N_VGND_c_1258_n 0.0113816f $X=7.59 $Y=0.74 $X2=0
+ $Y2=0
cc_339 N_A_435_99#_M1028_g N_VGND_c_1266_n 0.00383152f $X=7.16 $Y=0.74 $X2=0
+ $Y2=0
cc_340 N_A_435_99#_M1030_g N_VGND_c_1266_n 0.00383152f $X=7.59 $Y=0.74 $X2=0
+ $Y2=0
cc_341 N_A_435_99#_M1006_g N_VGND_c_1271_n 0.00434272f $X=6.3 $Y=0.74 $X2=0
+ $Y2=0
cc_342 N_A_435_99#_M1010_g N_VGND_c_1271_n 0.00383152f $X=6.73 $Y=0.74 $X2=0
+ $Y2=0
cc_343 N_A_435_99#_M1006_g N_VGND_c_1276_n 0.00825283f $X=6.3 $Y=0.74 $X2=0
+ $Y2=0
cc_344 N_A_435_99#_M1010_g N_VGND_c_1276_n 0.0075754f $X=6.73 $Y=0.74 $X2=0
+ $Y2=0
cc_345 N_A_435_99#_M1028_g N_VGND_c_1276_n 0.0075754f $X=7.16 $Y=0.74 $X2=0
+ $Y2=0
cc_346 N_A_435_99#_M1030_g N_VGND_c_1276_n 0.0075754f $X=7.59 $Y=0.74 $X2=0
+ $Y2=0
cc_347 N_A_435_99#_c_203_n N_A_707_119#_c_1378_n 0.0218973f $X=3.9 $Y=1.57 $X2=0
+ $Y2=0
cc_348 N_A_435_99#_c_236_p N_A_707_119#_c_1379_n 0.0207073f $X=4.115 $Y=0.74
+ $X2=0 $Y2=0
cc_349 N_A_435_99#_c_236_p N_A_707_119#_c_1381_n 0.0351355f $X=4.115 $Y=0.74
+ $X2=0 $Y2=0
cc_350 N_A_435_99#_c_218_n N_A_707_119#_c_1381_n 0.00163629f $X=4.07 $Y=1.907
+ $X2=0 $Y2=0
cc_351 N_A_435_99#_c_215_n N_A_707_119#_c_1382_n 0.0181607f $X=5.88 $Y=1.985
+ $X2=0 $Y2=0
cc_352 N_A_435_99#_c_205_n N_A_707_119#_c_1382_n 0.015926f $X=6.05 $Y=1.485
+ $X2=0 $Y2=0
cc_353 N_A_435_99#_c_219_n N_A_707_119#_c_1382_n 0.0399134f $X=4.955 $Y=1.985
+ $X2=0 $Y2=0
cc_354 N_A_435_99#_c_206_n N_A_707_119#_c_1382_n 6.87859e-19 $X=7.515 $Y=1.542
+ $X2=0 $Y2=0
cc_355 N_A_435_99#_c_218_n N_A_707_119#_c_1383_n 0.0133289f $X=4.07 $Y=1.907
+ $X2=0 $Y2=0
cc_356 N_A_435_99#_c_219_n N_A_707_119#_c_1383_n 0.0224715f $X=4.955 $Y=1.985
+ $X2=0 $Y2=0
cc_357 N_A_435_99#_M1006_g N_A_707_119#_c_1384_n 0.00559358f $X=6.3 $Y=0.74
+ $X2=0 $Y2=0
cc_358 N_A_435_99#_c_205_n N_A_707_119#_c_1384_n 0.00906645f $X=6.05 $Y=1.485
+ $X2=0 $Y2=0
cc_359 N_A_435_99#_c_206_n N_A_707_119#_c_1384_n 3.53737e-19 $X=7.515 $Y=1.542
+ $X2=0 $Y2=0
cc_360 N_B_M1000_g N_A_M1021_g 0.0108461f $X=1.36 $Y=0.945 $X2=0 $Y2=0
cc_361 N_B_c_395_n N_A_c_535_n 0.00888051f $X=1.395 $Y=1.885 $X2=0 $Y2=0
cc_362 N_B_M1000_g N_A_c_524_n 0.00894529f $X=1.36 $Y=0.945 $X2=0 $Y2=0
cc_363 N_B_M1004_g N_A_c_524_n 0.00879826f $X=1.79 $Y=0.945 $X2=0 $Y2=0
cc_364 N_B_M1001_g N_A_c_524_n 0.00880809f $X=3.9 $Y=0.915 $X2=0 $Y2=0
cc_365 N_B_M1035_g N_A_c_524_n 0.00880809f $X=4.33 $Y=0.915 $X2=0 $Y2=0
cc_366 N_B_c_392_n N_A_c_526_n 0.0044794f $X=4.255 $Y=1.605 $X2=0 $Y2=0
cc_367 N_B_c_408_n N_A_c_537_n 0.030511f $X=4.37 $Y=2.965 $X2=0 $Y2=0
cc_368 N_B_c_410_n N_A_c_537_n 0.00242326f $X=4.37 $Y=3.15 $X2=0 $Y2=0
cc_369 N_B_M1035_g N_A_M1002_g 0.0185653f $X=4.33 $Y=0.915 $X2=0 $Y2=0
cc_370 N_B_M1035_g N_A_c_530_n 0.0044794f $X=4.33 $Y=0.915 $X2=0 $Y2=0
cc_371 N_B_c_389_n A 0.01166f $X=1.935 $Y=1.805 $X2=0 $Y2=0
cc_372 B A 0.0204071f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_373 N_B_c_389_n N_A_c_533_n 0.0240678f $X=1.935 $Y=1.805 $X2=0 $Y2=0
cc_374 N_B_c_396_n N_A_294_392#_c_656_n 0.0129792f $X=1.845 $Y=1.885 $X2=0 $Y2=0
cc_375 N_B_c_397_n N_A_294_392#_c_656_n 0.00742923f $X=2.28 $Y=1.805 $X2=0 $Y2=0
cc_376 N_B_c_389_n N_A_294_392#_c_656_n 0.00143098f $X=1.935 $Y=1.805 $X2=0
+ $Y2=0
cc_377 N_B_c_399_n N_A_294_392#_c_656_n 0.016575f $X=2.355 $Y=3.075 $X2=0 $Y2=0
cc_378 B N_A_294_392#_c_656_n 0.0399444f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_379 N_B_M1004_g N_A_294_392#_c_647_n 3.97112e-19 $X=1.79 $Y=0.945 $X2=0 $Y2=0
cc_380 N_B_c_397_n N_A_294_392#_c_647_n 0.00369409f $X=2.28 $Y=1.805 $X2=0 $Y2=0
cc_381 N_B_c_389_n N_A_294_392#_c_647_n 8.30845e-19 $X=1.935 $Y=1.805 $X2=0
+ $Y2=0
cc_382 B N_A_294_392#_c_647_n 0.0222825f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_383 N_B_M1012_g N_A_294_392#_c_677_n 0.0154753f $X=3.765 $Y=2.315 $X2=0 $Y2=0
cc_384 N_B_c_406_n N_A_294_392#_c_680_n 0.00418617f $X=4.28 $Y=3.15 $X2=0 $Y2=0
cc_385 N_B_c_408_n N_A_294_392#_c_680_n 0.012845f $X=4.37 $Y=2.965 $X2=0 $Y2=0
cc_386 N_B_c_395_n N_A_294_392#_c_660_n 0.00917841f $X=1.395 $Y=1.885 $X2=0
+ $Y2=0
cc_387 N_B_c_389_n N_A_294_392#_c_660_n 0.00856402f $X=1.935 $Y=1.805 $X2=0
+ $Y2=0
cc_388 B N_A_294_392#_c_660_n 0.0143348f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_389 N_B_c_397_n N_A_294_392#_c_650_n 6.73123e-19 $X=2.28 $Y=1.805 $X2=0 $Y2=0
cc_390 N_B_c_399_n N_A_294_392#_c_661_n 0.00160313f $X=2.355 $Y=3.075 $X2=0
+ $Y2=0
cc_391 N_B_c_399_n N_A_294_392#_c_697_n 5.06216e-19 $X=2.355 $Y=3.075 $X2=0
+ $Y2=0
cc_392 N_B_M1012_g N_A_294_392#_c_697_n 0.00107405f $X=3.765 $Y=2.315 $X2=0
+ $Y2=0
cc_393 N_B_c_390_n N_A_294_392#_c_702_n 6.2107e-19 $X=3.765 $Y=1.82 $X2=0 $Y2=0
cc_394 N_B_M1012_g N_A_294_392#_c_702_n 0.00450988f $X=3.765 $Y=2.315 $X2=0
+ $Y2=0
cc_395 N_B_c_406_n N_A_294_392#_c_702_n 0.00404757f $X=4.28 $Y=3.15 $X2=0 $Y2=0
cc_396 N_B_c_408_n N_A_294_392#_c_702_n 0.00346968f $X=4.37 $Y=2.965 $X2=0 $Y2=0
cc_397 N_B_c_395_n N_A_27_392#_c_848_n 7.64109e-19 $X=1.395 $Y=1.885 $X2=0 $Y2=0
cc_398 N_B_c_395_n N_A_27_392#_c_849_n 0.0128006f $X=1.395 $Y=1.885 $X2=0 $Y2=0
cc_399 N_B_c_396_n N_A_27_392#_c_849_n 0.0125612f $X=1.845 $Y=1.885 $X2=0 $Y2=0
cc_400 N_B_c_399_n N_A_27_392#_c_849_n 0.00182056f $X=2.355 $Y=3.075 $X2=0 $Y2=0
cc_401 N_B_c_395_n N_A_27_392#_c_851_n 5.92376e-19 $X=1.395 $Y=1.885 $X2=0 $Y2=0
cc_402 N_B_c_396_n N_A_27_392#_c_851_n 0.00807036f $X=1.845 $Y=1.885 $X2=0 $Y2=0
cc_403 N_B_c_399_n N_A_27_392#_c_851_n 0.00805541f $X=2.355 $Y=3.075 $X2=0 $Y2=0
cc_404 N_B_c_399_n N_VPWR_c_891_n 0.00952443f $X=2.355 $Y=3.075 $X2=0 $Y2=0
cc_405 N_B_c_400_n N_VPWR_c_891_n 0.0230431f $X=3.675 $Y=3.15 $X2=0 $Y2=0
cc_406 N_B_c_400_n N_VPWR_c_892_n 0.0171462f $X=3.675 $Y=3.15 $X2=0 $Y2=0
cc_407 N_B_c_402_n N_VPWR_c_892_n 0.00361762f $X=3.765 $Y=2.9 $X2=0 $Y2=0
cc_408 N_B_c_403_n N_VPWR_c_892_n 0.007217f $X=3.765 $Y=3.075 $X2=0 $Y2=0
cc_409 N_B_M1012_g N_VPWR_c_892_n 0.00722471f $X=3.765 $Y=2.315 $X2=0 $Y2=0
cc_410 N_B_c_408_n N_VPWR_c_892_n 0.00200981f $X=4.37 $Y=2.965 $X2=0 $Y2=0
cc_411 N_B_c_409_n N_VPWR_c_892_n 0.00476669f $X=3.765 $Y=3.15 $X2=0 $Y2=0
cc_412 N_B_c_410_n N_VPWR_c_892_n 4.89576e-19 $X=4.37 $Y=3.15 $X2=0 $Y2=0
cc_413 N_B_c_402_n N_VPWR_c_893_n 0.00118913f $X=3.765 $Y=2.9 $X2=0 $Y2=0
cc_414 N_B_M1012_g N_VPWR_c_893_n 6.58575e-19 $X=3.765 $Y=2.315 $X2=0 $Y2=0
cc_415 N_B_c_408_n N_VPWR_c_893_n 0.00718962f $X=4.37 $Y=2.965 $X2=0 $Y2=0
cc_416 N_B_c_410_n N_VPWR_c_893_n 0.012213f $X=4.37 $Y=3.15 $X2=0 $Y2=0
cc_417 N_B_c_395_n N_VPWR_c_908_n 0.00278271f $X=1.395 $Y=1.885 $X2=0 $Y2=0
cc_418 N_B_c_396_n N_VPWR_c_908_n 0.00278257f $X=1.845 $Y=1.885 $X2=0 $Y2=0
cc_419 N_B_c_401_n N_VPWR_c_908_n 0.00757097f $X=2.43 $Y=3.15 $X2=0 $Y2=0
cc_420 N_B_c_400_n N_VPWR_c_909_n 0.0200847f $X=3.675 $Y=3.15 $X2=0 $Y2=0
cc_421 N_B_c_409_n N_VPWR_c_910_n 0.0265807f $X=3.765 $Y=3.15 $X2=0 $Y2=0
cc_422 N_B_c_395_n N_VPWR_c_889_n 0.00353907f $X=1.395 $Y=1.885 $X2=0 $Y2=0
cc_423 N_B_c_396_n N_VPWR_c_889_n 0.0035437f $X=1.845 $Y=1.885 $X2=0 $Y2=0
cc_424 N_B_c_400_n N_VPWR_c_889_n 0.0273473f $X=3.675 $Y=3.15 $X2=0 $Y2=0
cc_425 N_B_c_401_n N_VPWR_c_889_n 0.011411f $X=2.43 $Y=3.15 $X2=0 $Y2=0
cc_426 N_B_c_406_n N_VPWR_c_889_n 0.0136109f $X=4.28 $Y=3.15 $X2=0 $Y2=0
cc_427 N_B_c_409_n N_VPWR_c_889_n 0.00895426f $X=3.765 $Y=3.15 $X2=0 $Y2=0
cc_428 N_B_c_410_n N_VPWR_c_889_n 0.00453024f $X=4.37 $Y=3.15 $X2=0 $Y2=0
cc_429 N_B_M1000_g N_A_27_125#_c_1190_n 0.0159362f $X=1.36 $Y=0.945 $X2=0 $Y2=0
cc_430 N_B_M1004_g N_A_27_125#_c_1190_n 0.0118929f $X=1.79 $Y=0.945 $X2=0 $Y2=0
cc_431 N_B_c_397_n N_A_27_125#_c_1190_n 0.00102984f $X=2.28 $Y=1.805 $X2=0 $Y2=0
cc_432 N_B_c_389_n N_A_27_125#_c_1190_n 0.00442541f $X=1.935 $Y=1.805 $X2=0
+ $Y2=0
cc_433 B N_A_27_125#_c_1190_n 0.0488126f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_434 N_B_M1000_g N_A_27_125#_c_1191_n 6.55263e-19 $X=1.36 $Y=0.945 $X2=0 $Y2=0
cc_435 N_B_M1004_g N_A_27_125#_c_1191_n 0.00945767f $X=1.79 $Y=0.945 $X2=0 $Y2=0
cc_436 N_B_M1001_g N_A_27_125#_c_1194_n 0.00165882f $X=3.9 $Y=0.915 $X2=0 $Y2=0
cc_437 N_B_M1000_g N_VGND_c_1253_n 0.0073425f $X=1.36 $Y=0.945 $X2=0 $Y2=0
cc_438 N_B_M1004_g N_VGND_c_1253_n 9.59856e-19 $X=1.79 $Y=0.945 $X2=0 $Y2=0
cc_439 N_B_M1000_g N_VGND_c_1276_n 7.97988e-19 $X=1.36 $Y=0.945 $X2=0 $Y2=0
cc_440 N_B_M1004_g N_VGND_c_1276_n 7.94319e-19 $X=1.79 $Y=0.945 $X2=0 $Y2=0
cc_441 N_B_c_390_n N_A_707_119#_c_1378_n 5.74615e-19 $X=3.765 $Y=1.82 $X2=0
+ $Y2=0
cc_442 N_B_M1001_g N_A_707_119#_c_1378_n 0.00320107f $X=3.9 $Y=0.915 $X2=0 $Y2=0
cc_443 N_B_M1001_g N_A_707_119#_c_1379_n 0.0076245f $X=3.9 $Y=0.915 $X2=0 $Y2=0
cc_444 N_B_M1035_g N_A_707_119#_c_1379_n 0.00750518f $X=4.33 $Y=0.915 $X2=0
+ $Y2=0
cc_445 N_B_M1035_g N_A_707_119#_c_1381_n 0.00665243f $X=4.33 $Y=0.915 $X2=0
+ $Y2=0
cc_446 N_B_M1035_g N_A_707_119#_c_1383_n 0.0021197f $X=4.33 $Y=0.915 $X2=0 $Y2=0
cc_447 N_A_c_537_n N_A_294_392#_c_680_n 0.0131899f $X=4.82 $Y=1.975 $X2=0 $Y2=0
cc_448 N_A_c_538_n N_A_294_392#_c_680_n 0.0132176f $X=5.345 $Y=1.765 $X2=0 $Y2=0
cc_449 A N_A_27_392#_c_845_n 0.023f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_450 N_A_c_534_n N_A_27_392#_c_847_n 0.0126112f $X=0.495 $Y=1.885 $X2=0 $Y2=0
cc_451 N_A_c_535_n N_A_27_392#_c_847_n 0.0119694f $X=0.945 $Y=1.885 $X2=0 $Y2=0
cc_452 A N_A_27_392#_c_847_n 0.0455407f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_453 N_A_c_533_n N_A_27_392#_c_847_n 0.00799259f $X=0.93 $Y=1.67 $X2=0 $Y2=0
cc_454 N_A_c_535_n N_A_27_392#_c_848_n 3.67482e-19 $X=0.945 $Y=1.885 $X2=0 $Y2=0
cc_455 A N_A_27_392#_c_848_n 0.022047f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_456 N_A_c_534_n N_A_27_392#_c_866_n 4.46154e-19 $X=0.495 $Y=1.885 $X2=0 $Y2=0
cc_457 N_A_c_535_n N_A_27_392#_c_866_n 0.00926981f $X=0.945 $Y=1.885 $X2=0 $Y2=0
cc_458 N_A_c_535_n N_A_27_392#_c_850_n 0.0032261f $X=0.945 $Y=1.885 $X2=0 $Y2=0
cc_459 N_A_c_534_n N_VPWR_c_890_n 0.0134644f $X=0.495 $Y=1.885 $X2=0 $Y2=0
cc_460 N_A_c_535_n N_VPWR_c_890_n 0.0035512f $X=0.945 $Y=1.885 $X2=0 $Y2=0
cc_461 N_A_c_537_n N_VPWR_c_893_n 0.0138383f $X=4.82 $Y=1.975 $X2=0 $Y2=0
cc_462 N_A_c_538_n N_VPWR_c_893_n 6.88497e-19 $X=5.345 $Y=1.765 $X2=0 $Y2=0
cc_463 N_A_c_537_n N_VPWR_c_894_n 0.00473462f $X=4.82 $Y=1.975 $X2=0 $Y2=0
cc_464 N_A_c_538_n N_VPWR_c_894_n 0.00402388f $X=5.345 $Y=1.765 $X2=0 $Y2=0
cc_465 N_A_c_537_n N_VPWR_c_895_n 0.00552528f $X=4.82 $Y=1.975 $X2=0 $Y2=0
cc_466 N_A_c_538_n N_VPWR_c_895_n 0.00465104f $X=5.345 $Y=1.765 $X2=0 $Y2=0
cc_467 N_A_c_534_n N_VPWR_c_907_n 0.00413917f $X=0.495 $Y=1.885 $X2=0 $Y2=0
cc_468 N_A_c_535_n N_VPWR_c_908_n 0.0044313f $X=0.945 $Y=1.885 $X2=0 $Y2=0
cc_469 N_A_c_534_n N_VPWR_c_889_n 0.00821187f $X=0.495 $Y=1.885 $X2=0 $Y2=0
cc_470 N_A_c_535_n N_VPWR_c_889_n 0.00853445f $X=0.945 $Y=1.885 $X2=0 $Y2=0
cc_471 N_A_c_537_n N_VPWR_c_889_n 0.00474795f $X=4.82 $Y=1.975 $X2=0 $Y2=0
cc_472 N_A_c_538_n N_VPWR_c_889_n 0.00462577f $X=5.345 $Y=1.765 $X2=0 $Y2=0
cc_473 N_A_M1011_g N_A_27_125#_c_1186_n 4.43891e-19 $X=0.495 $Y=0.945 $X2=0
+ $Y2=0
cc_474 N_A_M1011_g N_A_27_125#_c_1187_n 0.0124643f $X=0.495 $Y=0.945 $X2=0 $Y2=0
cc_475 N_A_M1021_g N_A_27_125#_c_1187_n 0.0111806f $X=0.93 $Y=0.945 $X2=0 $Y2=0
cc_476 A N_A_27_125#_c_1187_n 0.0452882f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_477 N_A_c_533_n N_A_27_125#_c_1187_n 0.00270935f $X=0.93 $Y=1.67 $X2=0 $Y2=0
cc_478 A N_A_27_125#_c_1188_n 0.0212308f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_479 N_A_M1011_g N_A_27_125#_c_1189_n 5.76881e-19 $X=0.495 $Y=0.945 $X2=0
+ $Y2=0
cc_480 N_A_M1021_g N_A_27_125#_c_1189_n 0.00743339f $X=0.93 $Y=0.945 $X2=0 $Y2=0
cc_481 N_A_c_524_n N_A_27_125#_c_1189_n 0.0026496f $X=4.755 $Y=0.18 $X2=0 $Y2=0
cc_482 A N_A_27_125#_c_1190_n 0.00646543f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_483 N_A_c_524_n N_A_27_125#_c_1192_n 0.0189417f $X=4.755 $Y=0.18 $X2=0 $Y2=0
cc_484 N_A_c_524_n N_A_27_125#_c_1193_n 0.00772631f $X=4.755 $Y=0.18 $X2=0 $Y2=0
cc_485 N_A_M1021_g N_A_27_125#_c_1195_n 9.55648e-19 $X=0.93 $Y=0.945 $X2=0 $Y2=0
cc_486 A N_A_27_125#_c_1195_n 0.0218995f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_487 N_A_M1011_g N_VGND_c_1252_n 0.0104167f $X=0.495 $Y=0.945 $X2=0 $Y2=0
cc_488 N_A_c_525_n N_VGND_c_1252_n 0.013498f $X=1.005 $Y=0.18 $X2=0 $Y2=0
cc_489 N_A_M1021_g N_VGND_c_1253_n 0.00475281f $X=0.93 $Y=0.945 $X2=0 $Y2=0
cc_490 N_A_c_524_n N_VGND_c_1253_n 0.0203576f $X=4.755 $Y=0.18 $X2=0 $Y2=0
cc_491 N_A_c_524_n N_VGND_c_1254_n 0.0164781f $X=4.755 $Y=0.18 $X2=0 $Y2=0
cc_492 N_A_c_528_n N_VGND_c_1254_n 0.00453121f $X=5.255 $Y=1.47 $X2=0 $Y2=0
cc_493 N_A_c_529_n N_VGND_c_1254_n 0.0125021f $X=5.33 $Y=1.31 $X2=0 $Y2=0
cc_494 N_A_c_529_n N_VGND_c_1255_n 0.0035863f $X=5.33 $Y=1.31 $X2=0 $Y2=0
cc_495 N_A_c_529_n N_VGND_c_1256_n 0.00261122f $X=5.33 $Y=1.31 $X2=0 $Y2=0
cc_496 N_A_M1011_g N_VGND_c_1262_n 0.00345209f $X=0.495 $Y=0.945 $X2=0 $Y2=0
cc_497 N_A_c_525_n N_VGND_c_1264_n 0.0177193f $X=1.005 $Y=0.18 $X2=0 $Y2=0
cc_498 N_A_c_524_n N_VGND_c_1270_n 0.0773131f $X=4.755 $Y=0.18 $X2=0 $Y2=0
cc_499 N_A_M1011_g N_VGND_c_1276_n 0.00394323f $X=0.495 $Y=0.945 $X2=0 $Y2=0
cc_500 N_A_c_524_n N_VGND_c_1276_n 0.109515f $X=4.755 $Y=0.18 $X2=0 $Y2=0
cc_501 N_A_c_525_n N_VGND_c_1276_n 0.0106926f $X=1.005 $Y=0.18 $X2=0 $Y2=0
cc_502 N_A_c_529_n N_VGND_c_1276_n 0.00401353f $X=5.33 $Y=1.31 $X2=0 $Y2=0
cc_503 N_A_c_524_n N_A_707_119#_c_1379_n 0.0156098f $X=4.755 $Y=0.18 $X2=0 $Y2=0
cc_504 N_A_M1002_g N_A_707_119#_c_1379_n 0.00599831f $X=4.83 $Y=0.915 $X2=0
+ $Y2=0
cc_505 N_A_c_524_n N_A_707_119#_c_1380_n 0.00626586f $X=4.755 $Y=0.18 $X2=0
+ $Y2=0
cc_506 N_A_M1002_g N_A_707_119#_c_1381_n 0.01109f $X=4.83 $Y=0.915 $X2=0 $Y2=0
cc_507 N_A_c_529_n N_A_707_119#_c_1381_n 4.9686e-19 $X=5.33 $Y=1.31 $X2=0 $Y2=0
cc_508 N_A_c_530_n N_A_707_119#_c_1381_n 0.00685332f $X=4.73 $Y=1.46 $X2=0 $Y2=0
cc_509 N_A_c_528_n N_A_707_119#_c_1382_n 0.0129286f $X=5.255 $Y=1.47 $X2=0 $Y2=0
cc_510 N_A_c_530_n N_A_707_119#_c_1382_n 0.00979406f $X=4.73 $Y=1.46 $X2=0 $Y2=0
cc_511 N_A_c_531_n N_A_707_119#_c_1382_n 0.0141867f $X=5.255 $Y=1.31 $X2=0 $Y2=0
cc_512 N_A_c_530_n N_A_707_119#_c_1383_n 0.00408548f $X=4.73 $Y=1.46 $X2=0 $Y2=0
cc_513 N_A_c_529_n N_A_707_119#_c_1384_n 0.00688907f $X=5.33 $Y=1.31 $X2=0 $Y2=0
cc_514 N_A_294_392#_c_656_n N_A_27_392#_M1014_s 0.00242368f $X=2.5 $Y=2.04 $X2=0
+ $Y2=0
cc_515 N_A_294_392#_c_660_n N_A_27_392#_c_848_n 0.013101f $X=1.62 $Y=2.12 $X2=0
+ $Y2=0
cc_516 N_A_294_392#_c_660_n N_A_27_392#_c_866_n 0.0403355f $X=1.62 $Y=2.12 $X2=0
+ $Y2=0
cc_517 N_A_294_392#_M1007_d N_A_27_392#_c_849_n 0.00197722f $X=1.47 $Y=1.96
+ $X2=0 $Y2=0
cc_518 N_A_294_392#_c_660_n N_A_27_392#_c_849_n 0.0151173f $X=1.62 $Y=2.12 $X2=0
+ $Y2=0
cc_519 N_A_294_392#_c_656_n N_A_27_392#_c_851_n 0.0220233f $X=2.5 $Y=2.04 $X2=0
+ $Y2=0
cc_520 N_A_294_392#_c_675_n N_VPWR_M1009_s 0.00174738f $X=2.925 $Y=2.015 $X2=0
+ $Y2=0
cc_521 N_A_294_392#_c_661_n N_VPWR_M1009_s 0.00228391f $X=2.585 $Y=2.015 $X2=0
+ $Y2=0
cc_522 N_A_294_392#_c_677_n N_VPWR_M1016_s 0.00507752f $X=3.9 $Y=2.25 $X2=0
+ $Y2=0
cc_523 N_A_294_392#_c_680_n N_VPWR_M1023_d 0.00463005f $X=7.725 $Y=2.405 $X2=0
+ $Y2=0
cc_524 N_A_294_392#_c_680_n N_VPWR_M1019_d 0.00990181f $X=7.725 $Y=2.405 $X2=0
+ $Y2=0
cc_525 N_A_294_392#_c_680_n N_VPWR_M1025_s 0.00379251f $X=7.725 $Y=2.405 $X2=0
+ $Y2=0
cc_526 N_A_294_392#_c_680_n N_VPWR_M1032_s 0.00491342f $X=7.725 $Y=2.405 $X2=0
+ $Y2=0
cc_527 N_A_294_392#_c_658_n N_VPWR_M1032_s 0.00447084f $X=7.81 $Y=2.32 $X2=0
+ $Y2=0
cc_528 N_A_294_392#_c_656_n N_VPWR_c_891_n 0.00140427f $X=2.5 $Y=2.04 $X2=0
+ $Y2=0
cc_529 N_A_294_392#_c_675_n N_VPWR_c_891_n 0.00427983f $X=2.925 $Y=2.015 $X2=0
+ $Y2=0
cc_530 N_A_294_392#_c_661_n N_VPWR_c_891_n 0.0105347f $X=2.585 $Y=2.015 $X2=0
+ $Y2=0
cc_531 N_A_294_392#_c_677_n N_VPWR_c_892_n 0.0171814f $X=3.9 $Y=2.25 $X2=0 $Y2=0
cc_532 N_A_294_392#_c_680_n N_VPWR_c_893_n 0.0168032f $X=7.725 $Y=2.405 $X2=0
+ $Y2=0
cc_533 N_A_294_392#_c_680_n N_VPWR_c_895_n 0.0314412f $X=7.725 $Y=2.405 $X2=0
+ $Y2=0
cc_534 N_A_294_392#_c_680_n N_VPWR_c_896_n 0.0168032f $X=7.725 $Y=2.405 $X2=0
+ $Y2=0
cc_535 N_A_294_392#_c_651_n N_VPWR_c_897_n 0.00728862f $X=7.965 $Y=1.765 $X2=0
+ $Y2=0
cc_536 N_A_294_392#_c_652_n N_VPWR_c_897_n 4.09834e-19 $X=8.415 $Y=1.765 $X2=0
+ $Y2=0
cc_537 N_A_294_392#_c_680_n N_VPWR_c_897_n 0.0169636f $X=7.725 $Y=2.405 $X2=0
+ $Y2=0
cc_538 N_A_294_392#_c_651_n N_VPWR_c_898_n 4.98648e-19 $X=7.965 $Y=1.765 $X2=0
+ $Y2=0
cc_539 N_A_294_392#_c_652_n N_VPWR_c_898_n 0.0107727f $X=8.415 $Y=1.765 $X2=0
+ $Y2=0
cc_540 N_A_294_392#_c_653_n N_VPWR_c_898_n 0.0130813f $X=8.865 $Y=1.765 $X2=0
+ $Y2=0
cc_541 N_A_294_392#_c_655_n N_VPWR_c_898_n 6.06284e-19 $X=9.575 $Y=1.765 $X2=0
+ $Y2=0
cc_542 N_A_294_392#_c_653_n N_VPWR_c_900_n 5.86256e-19 $X=8.865 $Y=1.765 $X2=0
+ $Y2=0
cc_543 N_A_294_392#_c_655_n N_VPWR_c_900_n 0.0130652f $X=9.575 $Y=1.765 $X2=0
+ $Y2=0
cc_544 N_A_294_392#_c_651_n N_VPWR_c_905_n 0.00413917f $X=7.965 $Y=1.765 $X2=0
+ $Y2=0
cc_545 N_A_294_392#_c_652_n N_VPWR_c_905_n 0.00413917f $X=8.415 $Y=1.765 $X2=0
+ $Y2=0
cc_546 N_A_294_392#_c_653_n N_VPWR_c_911_n 0.00413917f $X=8.865 $Y=1.765 $X2=0
+ $Y2=0
cc_547 N_A_294_392#_c_655_n N_VPWR_c_911_n 0.00413917f $X=9.575 $Y=1.765 $X2=0
+ $Y2=0
cc_548 N_A_294_392#_c_651_n N_VPWR_c_889_n 0.00817726f $X=7.965 $Y=1.765 $X2=0
+ $Y2=0
cc_549 N_A_294_392#_c_652_n N_VPWR_c_889_n 0.00817726f $X=8.415 $Y=1.765 $X2=0
+ $Y2=0
cc_550 N_A_294_392#_c_653_n N_VPWR_c_889_n 0.00819705f $X=8.865 $Y=1.765 $X2=0
+ $Y2=0
cc_551 N_A_294_392#_c_655_n N_VPWR_c_889_n 0.00819705f $X=9.575 $Y=1.765 $X2=0
+ $Y2=0
cc_552 N_A_294_392#_c_680_n N_VPWR_c_889_n 0.0807447f $X=7.725 $Y=2.405 $X2=0
+ $Y2=0
cc_553 N_A_294_392#_c_702_n N_VPWR_c_889_n 0.00553057f $X=3.985 $Y=2.25 $X2=0
+ $Y2=0
cc_554 N_A_294_392#_c_680_n N_COUT_M1017_d 0.0120222f $X=7.725 $Y=2.405 $X2=0
+ $Y2=0
cc_555 N_A_294_392#_c_680_n N_COUT_M1031_d 0.00556775f $X=7.725 $Y=2.405 $X2=0
+ $Y2=0
cc_556 N_A_294_392#_c_680_n N_COUT_c_1049_n 0.0566155f $X=7.725 $Y=2.405 $X2=0
+ $Y2=0
cc_557 N_A_294_392#_M1003_g N_COUT_c_1066_n 7.75513e-19 $X=8.02 $Y=0.74 $X2=0
+ $Y2=0
cc_558 N_A_294_392#_M1003_g COUT 9.08516e-19 $X=8.02 $Y=0.74 $X2=0 $Y2=0
cc_559 N_A_294_392#_c_644_n COUT 3.86397e-19 $X=9.025 $Y=1.485 $X2=0 $Y2=0
cc_560 N_A_294_392#_c_658_n COUT 0.0127062f $X=7.81 $Y=2.32 $X2=0 $Y2=0
cc_561 N_A_294_392#_c_648_n COUT 0.027912f $X=7.895 $Y=1.485 $X2=0 $Y2=0
cc_562 N_A_294_392#_c_651_n N_COUT_c_1075_n 3.05965e-19 $X=7.965 $Y=1.765 $X2=0
+ $Y2=0
cc_563 N_A_294_392#_c_680_n N_COUT_c_1075_n 0.0227509f $X=7.725 $Y=2.405 $X2=0
+ $Y2=0
cc_564 N_A_294_392#_c_658_n N_COUT_c_1075_n 0.0259639f $X=7.81 $Y=2.32 $X2=0
+ $Y2=0
cc_565 N_A_294_392#_c_644_n N_SUM_c_1104_n 0.00587074f $X=9.025 $Y=1.485 $X2=0
+ $Y2=0
cc_566 N_A_294_392#_c_658_n N_SUM_c_1104_n 0.011581f $X=7.81 $Y=2.32 $X2=0 $Y2=0
cc_567 N_A_294_392#_c_782_p N_SUM_c_1104_n 0.0193967f $X=9.56 $Y=1.485 $X2=0
+ $Y2=0
cc_568 N_A_294_392#_c_651_n N_SUM_c_1105_n 4.08598e-19 $X=7.965 $Y=1.765 $X2=0
+ $Y2=0
cc_569 N_A_294_392#_c_652_n N_SUM_c_1105_n 4.08598e-19 $X=8.415 $Y=1.765 $X2=0
+ $Y2=0
cc_570 N_A_294_392#_M1003_g N_SUM_c_1097_n 3.97481e-19 $X=8.02 $Y=0.74 $X2=0
+ $Y2=0
cc_571 N_A_294_392#_M1015_g N_SUM_c_1097_n 0.00903544f $X=8.45 $Y=0.74 $X2=0
+ $Y2=0
cc_572 N_A_294_392#_M1024_g N_SUM_c_1097_n 6.75677e-19 $X=8.95 $Y=0.74 $X2=0
+ $Y2=0
cc_573 N_A_294_392#_M1015_g N_SUM_c_1098_n 0.0115433f $X=8.45 $Y=0.74 $X2=0
+ $Y2=0
cc_574 N_A_294_392#_M1024_g N_SUM_c_1098_n 0.0153874f $X=8.95 $Y=0.74 $X2=0
+ $Y2=0
cc_575 N_A_294_392#_c_644_n N_SUM_c_1098_n 0.00382577f $X=9.025 $Y=1.485 $X2=0
+ $Y2=0
cc_576 N_A_294_392#_c_782_p N_SUM_c_1098_n 0.0492199f $X=9.56 $Y=1.485 $X2=0
+ $Y2=0
cc_577 N_A_294_392#_M1003_g N_SUM_c_1099_n 6.07621e-19 $X=8.02 $Y=0.74 $X2=0
+ $Y2=0
cc_578 N_A_294_392#_M1015_g N_SUM_c_1099_n 0.00110424f $X=8.45 $Y=0.74 $X2=0
+ $Y2=0
cc_579 N_A_294_392#_c_644_n N_SUM_c_1099_n 0.00232957f $X=9.025 $Y=1.485 $X2=0
+ $Y2=0
cc_580 N_A_294_392#_c_782_p N_SUM_c_1099_n 0.0209731f $X=9.56 $Y=1.485 $X2=0
+ $Y2=0
cc_581 N_A_294_392#_M1024_g N_SUM_c_1100_n 0.00377577f $X=8.95 $Y=0.74 $X2=0
+ $Y2=0
cc_582 N_A_294_392#_M1027_g N_SUM_c_1100_n 5.54424e-19 $X=9.505 $Y=0.74 $X2=0
+ $Y2=0
cc_583 N_A_294_392#_c_653_n N_SUM_c_1106_n 0.0116309f $X=8.865 $Y=1.765 $X2=0
+ $Y2=0
cc_584 N_A_294_392#_c_655_n N_SUM_c_1106_n 0.0120444f $X=9.575 $Y=1.765 $X2=0
+ $Y2=0
cc_585 N_A_294_392#_M1027_g N_SUM_c_1101_n 0.015246f $X=9.505 $Y=0.74 $X2=0
+ $Y2=0
cc_586 N_A_294_392#_c_782_p N_SUM_c_1101_n 0.0177771f $X=9.56 $Y=1.485 $X2=0
+ $Y2=0
cc_587 N_A_294_392#_c_649_n N_SUM_c_1101_n 0.00394214f $X=9.56 $Y=1.485 $X2=0
+ $Y2=0
cc_588 N_A_294_392#_c_643_n N_SUM_c_1107_n 0.00211105f $X=9.43 $Y=1.485 $X2=0
+ $Y2=0
cc_589 N_A_294_392#_c_655_n N_SUM_c_1107_n 0.0265998f $X=9.575 $Y=1.765 $X2=0
+ $Y2=0
cc_590 N_A_294_392#_c_782_p N_SUM_c_1107_n 0.0171428f $X=9.56 $Y=1.485 $X2=0
+ $Y2=0
cc_591 N_A_294_392#_c_649_n N_SUM_c_1107_n 0.00269293f $X=9.56 $Y=1.485 $X2=0
+ $Y2=0
cc_592 N_A_294_392#_M1027_g N_SUM_c_1102_n 0.00533837f $X=9.505 $Y=0.74 $X2=0
+ $Y2=0
cc_593 N_A_294_392#_c_655_n N_SUM_c_1102_n 0.00183882f $X=9.575 $Y=1.765 $X2=0
+ $Y2=0
cc_594 N_A_294_392#_c_782_p N_SUM_c_1102_n 0.0250942f $X=9.56 $Y=1.485 $X2=0
+ $Y2=0
cc_595 N_A_294_392#_c_649_n N_SUM_c_1102_n 0.0135758f $X=9.56 $Y=1.485 $X2=0
+ $Y2=0
cc_596 N_A_294_392#_c_643_n N_SUM_c_1103_n 0.00524152f $X=9.43 $Y=1.485 $X2=0
+ $Y2=0
cc_597 N_A_294_392#_c_782_p N_SUM_c_1103_n 0.0278321f $X=9.56 $Y=1.485 $X2=0
+ $Y2=0
cc_598 N_A_294_392#_c_652_n N_SUM_c_1109_n 0.0176976f $X=8.415 $Y=1.765 $X2=0
+ $Y2=0
cc_599 N_A_294_392#_c_653_n N_SUM_c_1109_n 0.0204453f $X=8.865 $Y=1.765 $X2=0
+ $Y2=0
cc_600 N_A_294_392#_c_644_n N_SUM_c_1109_n 0.0121059f $X=9.025 $Y=1.485 $X2=0
+ $Y2=0
cc_601 N_A_294_392#_c_782_p N_SUM_c_1109_n 0.0577212f $X=9.56 $Y=1.485 $X2=0
+ $Y2=0
cc_602 N_A_294_392#_c_643_n N_SUM_c_1110_n 0.00810171f $X=9.43 $Y=1.485 $X2=0
+ $Y2=0
cc_603 N_A_294_392#_c_782_p N_SUM_c_1110_n 0.0262156f $X=9.56 $Y=1.485 $X2=0
+ $Y2=0
cc_604 N_A_294_392#_c_782_p N_SUM_c_1151_n 0.0032968f $X=9.56 $Y=1.485 $X2=0
+ $Y2=0
cc_605 N_A_294_392#_c_653_n N_SUM_c_1152_n 0.00598214f $X=8.865 $Y=1.765 $X2=0
+ $Y2=0
cc_606 N_A_294_392#_c_782_p N_SUM_c_1152_n 0.00167912f $X=9.56 $Y=1.485 $X2=0
+ $Y2=0
cc_607 N_A_294_392#_c_660_n N_A_27_125#_c_1190_n 0.00344089f $X=1.62 $Y=2.12
+ $X2=0 $Y2=0
cc_608 N_A_294_392#_c_650_n N_A_27_125#_c_1190_n 0.00167954f $X=2.505 $Y=1.285
+ $X2=0 $Y2=0
cc_609 N_A_294_392#_c_646_n N_A_27_125#_c_1191_n 0.00158095f $X=2.505 $Y=0.77
+ $X2=0 $Y2=0
cc_610 N_A_294_392#_c_646_n N_A_27_125#_c_1192_n 0.0258724f $X=2.505 $Y=0.77
+ $X2=0 $Y2=0
cc_611 N_A_294_392#_c_646_n N_A_27_125#_c_1194_n 0.0243921f $X=2.505 $Y=0.77
+ $X2=0 $Y2=0
cc_612 N_A_294_392#_c_675_n N_A_27_125#_c_1194_n 0.00208042f $X=2.925 $Y=2.015
+ $X2=0 $Y2=0
cc_613 N_A_294_392#_c_697_n N_A_27_125#_c_1194_n 0.00363854f $X=3.09 $Y=2.07
+ $X2=0 $Y2=0
cc_614 N_A_294_392#_M1003_g N_VGND_c_1258_n 0.00842225f $X=8.02 $Y=0.74 $X2=0
+ $Y2=0
cc_615 N_A_294_392#_M1015_g N_VGND_c_1258_n 4.51782e-19 $X=8.45 $Y=0.74 $X2=0
+ $Y2=0
cc_616 N_A_294_392#_c_648_n N_VGND_c_1258_n 0.00597123f $X=7.895 $Y=1.485 $X2=0
+ $Y2=0
cc_617 N_A_294_392#_c_782_p N_VGND_c_1258_n 0.00128723f $X=9.56 $Y=1.485 $X2=0
+ $Y2=0
cc_618 N_A_294_392#_M1015_g N_VGND_c_1259_n 0.00408259f $X=8.45 $Y=0.74 $X2=0
+ $Y2=0
cc_619 N_A_294_392#_M1024_g N_VGND_c_1259_n 0.00997407f $X=8.95 $Y=0.74 $X2=0
+ $Y2=0
cc_620 N_A_294_392#_M1027_g N_VGND_c_1259_n 6.10235e-19 $X=9.505 $Y=0.74 $X2=0
+ $Y2=0
cc_621 N_A_294_392#_M1027_g N_VGND_c_1261_n 0.00694336f $X=9.505 $Y=0.74 $X2=0
+ $Y2=0
cc_622 N_A_294_392#_M1003_g N_VGND_c_1268_n 0.00383152f $X=8.02 $Y=0.74 $X2=0
+ $Y2=0
cc_623 N_A_294_392#_M1015_g N_VGND_c_1268_n 0.00434272f $X=8.45 $Y=0.74 $X2=0
+ $Y2=0
cc_624 N_A_294_392#_M1024_g N_VGND_c_1272_n 0.00383152f $X=8.95 $Y=0.74 $X2=0
+ $Y2=0
cc_625 N_A_294_392#_M1027_g N_VGND_c_1272_n 0.00460063f $X=9.505 $Y=0.74 $X2=0
+ $Y2=0
cc_626 N_A_294_392#_M1003_g N_VGND_c_1276_n 0.0075754f $X=8.02 $Y=0.74 $X2=0
+ $Y2=0
cc_627 N_A_294_392#_M1015_g N_VGND_c_1276_n 0.00820718f $X=8.45 $Y=0.74 $X2=0
+ $Y2=0
cc_628 N_A_294_392#_M1024_g N_VGND_c_1276_n 0.00758657f $X=8.95 $Y=0.74 $X2=0
+ $Y2=0
cc_629 N_A_294_392#_M1027_g N_VGND_c_1276_n 0.00912119f $X=9.505 $Y=0.74 $X2=0
+ $Y2=0
cc_630 N_A_27_392#_c_847_n N_VPWR_M1033_d 0.00222494f $X=1.005 $Y=2.04 $X2=-0.19
+ $Y2=1.66
cc_631 N_A_27_392#_c_846_n N_VPWR_c_890_n 0.0242552f $X=0.27 $Y=2.8 $X2=0 $Y2=0
cc_632 N_A_27_392#_c_847_n N_VPWR_c_890_n 0.0154248f $X=1.005 $Y=2.04 $X2=0
+ $Y2=0
cc_633 N_A_27_392#_c_866_n N_VPWR_c_890_n 0.0400325f $X=1.17 $Y=2.815 $X2=0
+ $Y2=0
cc_634 N_A_27_392#_c_850_n N_VPWR_c_890_n 0.012272f $X=1.255 $Y=2.99 $X2=0 $Y2=0
cc_635 N_A_27_392#_c_849_n N_VPWR_c_891_n 0.0117895f $X=1.905 $Y=2.99 $X2=0
+ $Y2=0
cc_636 N_A_27_392#_c_851_n N_VPWR_c_891_n 0.0326488f $X=2.07 $Y=2.38 $X2=0 $Y2=0
cc_637 N_A_27_392#_c_846_n N_VPWR_c_907_n 0.0116996f $X=0.27 $Y=2.8 $X2=0 $Y2=0
cc_638 N_A_27_392#_c_849_n N_VPWR_c_908_n 0.0645908f $X=1.905 $Y=2.99 $X2=0
+ $Y2=0
cc_639 N_A_27_392#_c_850_n N_VPWR_c_908_n 0.017869f $X=1.255 $Y=2.99 $X2=0 $Y2=0
cc_640 N_A_27_392#_c_846_n N_VPWR_c_889_n 0.0101742f $X=0.27 $Y=2.8 $X2=0 $Y2=0
cc_641 N_A_27_392#_c_849_n N_VPWR_c_889_n 0.0358952f $X=1.905 $Y=2.99 $X2=0
+ $Y2=0
cc_642 N_A_27_392#_c_850_n N_VPWR_c_889_n 0.00965079f $X=1.255 $Y=2.99 $X2=0
+ $Y2=0
cc_643 N_A_27_392#_c_845_n N_A_27_125#_c_1188_n 3.57272e-19 $X=0.245 $Y=2.125
+ $X2=0 $Y2=0
cc_644 N_VPWR_M1025_s N_COUT_c_1049_n 0.00202293f $X=6.69 $Y=1.84 $X2=0 $Y2=0
cc_645 N_VPWR_c_897_n N_SUM_c_1105_n 0.0127556f $X=7.74 $Y=2.78 $X2=0 $Y2=0
cc_646 N_VPWR_c_898_n N_SUM_c_1105_n 0.0255132f $X=8.64 $Y=2.405 $X2=0 $Y2=0
cc_647 N_VPWR_c_905_n N_SUM_c_1105_n 0.0101736f $X=8.475 $Y=3.33 $X2=0 $Y2=0
cc_648 N_VPWR_c_889_n N_SUM_c_1105_n 0.0084208f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_649 N_VPWR_c_898_n N_SUM_c_1106_n 0.0359682f $X=8.64 $Y=2.405 $X2=0 $Y2=0
cc_650 N_VPWR_c_900_n N_SUM_c_1106_n 0.0406518f $X=9.8 $Y=2.415 $X2=0 $Y2=0
cc_651 N_VPWR_c_911_n N_SUM_c_1106_n 0.0146357f $X=9.635 $Y=3.33 $X2=0 $Y2=0
cc_652 N_VPWR_c_889_n N_SUM_c_1106_n 0.0121141f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_653 N_VPWR_M1029_s N_SUM_c_1107_n 5.52306e-19 $X=9.65 $Y=1.84 $X2=0 $Y2=0
cc_654 N_VPWR_c_900_n N_SUM_c_1107_n 0.00960525f $X=9.8 $Y=2.415 $X2=0 $Y2=0
cc_655 N_VPWR_M1029_s N_SUM_c_1102_n 0.00253733f $X=9.65 $Y=1.84 $X2=0 $Y2=0
cc_656 N_VPWR_c_900_n N_SUM_c_1102_n 0.0101282f $X=9.8 $Y=2.415 $X2=0 $Y2=0
cc_657 N_VPWR_M1013_s N_SUM_c_1109_n 0.00201799f $X=8.49 $Y=1.84 $X2=0 $Y2=0
cc_658 N_VPWR_c_898_n N_SUM_c_1109_n 0.0188168f $X=8.64 $Y=2.405 $X2=0 $Y2=0
cc_659 N_VPWR_c_900_n N_SUM_c_1151_n 4.38649e-19 $X=9.8 $Y=2.415 $X2=0 $Y2=0
cc_660 N_VPWR_c_898_n N_SUM_c_1152_n 0.00189266f $X=8.64 $Y=2.405 $X2=0 $Y2=0
cc_661 N_VPWR_M1029_s SUM 0.00196766f $X=9.65 $Y=1.84 $X2=0 $Y2=0
cc_662 N_VPWR_c_900_n SUM 0.00488527f $X=9.8 $Y=2.415 $X2=0 $Y2=0
cc_663 N_COUT_c_1066_n N_SUM_c_1099_n 0.00260272f $X=7.382 $Y=1.13 $X2=0 $Y2=0
cc_664 COUT N_SUM_c_1099_n 6.38315e-19 $X=7.355 $Y=1.21 $X2=0 $Y2=0
cc_665 N_COUT_c_1048_n N_VGND_M1010_d 0.00178571f $X=7.21 $Y=1.005 $X2=0 $Y2=0
cc_666 N_COUT_c_1046_n N_VGND_c_1256_n 0.0107873f $X=6.475 $Y=0.88 $X2=0 $Y2=0
cc_667 N_COUT_c_1047_n N_VGND_c_1256_n 0.0188983f $X=6.515 $Y=0.515 $X2=0 $Y2=0
cc_668 N_COUT_c_1047_n N_VGND_c_1257_n 0.0136308f $X=6.515 $Y=0.515 $X2=0 $Y2=0
cc_669 N_COUT_c_1048_n N_VGND_c_1257_n 0.0175375f $X=7.21 $Y=1.005 $X2=0 $Y2=0
cc_670 N_COUT_c_1047_n N_VGND_c_1271_n 0.0109942f $X=6.515 $Y=0.515 $X2=0 $Y2=0
cc_671 N_COUT_c_1047_n N_VGND_c_1276_n 0.00904371f $X=6.515 $Y=0.515 $X2=0 $Y2=0
cc_672 N_SUM_c_1098_n N_VGND_M1015_d 0.00250873f $X=9.07 $Y=1.065 $X2=0 $Y2=0
cc_673 N_SUM_c_1101_n N_VGND_M1027_d 0.00317529f $X=9.825 $Y=1.065 $X2=0 $Y2=0
cc_674 N_SUM_c_1097_n N_VGND_c_1258_n 0.0136308f $X=8.235 $Y=0.515 $X2=0 $Y2=0
cc_675 N_SUM_c_1097_n N_VGND_c_1259_n 0.0173318f $X=8.235 $Y=0.515 $X2=0 $Y2=0
cc_676 N_SUM_c_1098_n N_VGND_c_1259_n 0.0210288f $X=9.07 $Y=1.065 $X2=0 $Y2=0
cc_677 N_SUM_c_1100_n N_VGND_c_1259_n 0.0180508f $X=9.235 $Y=0.515 $X2=0 $Y2=0
cc_678 N_SUM_c_1100_n N_VGND_c_1261_n 0.0157236f $X=9.235 $Y=0.515 $X2=0 $Y2=0
cc_679 N_SUM_c_1101_n N_VGND_c_1261_n 0.0206457f $X=9.825 $Y=1.065 $X2=0 $Y2=0
cc_680 N_SUM_c_1097_n N_VGND_c_1268_n 0.0109942f $X=8.235 $Y=0.515 $X2=0 $Y2=0
cc_681 N_SUM_c_1100_n N_VGND_c_1272_n 0.0146357f $X=9.235 $Y=0.515 $X2=0 $Y2=0
cc_682 N_SUM_c_1097_n N_VGND_c_1276_n 0.00904371f $X=8.235 $Y=0.515 $X2=0 $Y2=0
cc_683 N_SUM_c_1100_n N_VGND_c_1276_n 0.0121141f $X=9.235 $Y=0.515 $X2=0 $Y2=0
cc_684 N_A_27_125#_c_1187_n N_VGND_M1011_s 0.00177524f $X=0.98 $Y=1.2 $X2=-0.19
+ $Y2=-0.245
cc_685 N_A_27_125#_c_1190_n N_VGND_M1000_d 0.00176461f $X=1.84 $Y=1.2 $X2=0
+ $Y2=0
cc_686 N_A_27_125#_c_1186_n N_VGND_c_1252_n 0.0124064f $X=0.28 $Y=0.77 $X2=0
+ $Y2=0
cc_687 N_A_27_125#_c_1187_n N_VGND_c_1252_n 0.015373f $X=0.98 $Y=1.2 $X2=0 $Y2=0
cc_688 N_A_27_125#_c_1189_n N_VGND_c_1252_n 0.0237383f $X=1.145 $Y=0.77 $X2=0
+ $Y2=0
cc_689 N_A_27_125#_c_1189_n N_VGND_c_1253_n 0.0124064f $X=1.145 $Y=0.77 $X2=0
+ $Y2=0
cc_690 N_A_27_125#_c_1190_n N_VGND_c_1253_n 0.0152916f $X=1.84 $Y=1.2 $X2=0
+ $Y2=0
cc_691 N_A_27_125#_c_1191_n N_VGND_c_1253_n 0.0257313f $X=2.005 $Y=0.77 $X2=0
+ $Y2=0
cc_692 N_A_27_125#_c_1193_n N_VGND_c_1253_n 0.0141601f $X=2.17 $Y=0.35 $X2=0
+ $Y2=0
cc_693 N_A_27_125#_c_1186_n N_VGND_c_1262_n 0.00535163f $X=0.28 $Y=0.77 $X2=0
+ $Y2=0
cc_694 N_A_27_125#_c_1189_n N_VGND_c_1264_n 0.00529024f $X=1.145 $Y=0.77 $X2=0
+ $Y2=0
cc_695 N_A_27_125#_c_1192_n N_VGND_c_1270_n 0.0627959f $X=2.84 $Y=0.35 $X2=0
+ $Y2=0
cc_696 N_A_27_125#_c_1193_n N_VGND_c_1270_n 0.0222408f $X=2.17 $Y=0.35 $X2=0
+ $Y2=0
cc_697 N_A_27_125#_c_1186_n N_VGND_c_1276_n 0.00769355f $X=0.28 $Y=0.77 $X2=0
+ $Y2=0
cc_698 N_A_27_125#_c_1189_n N_VGND_c_1276_n 0.00666603f $X=1.145 $Y=0.77 $X2=0
+ $Y2=0
cc_699 N_A_27_125#_c_1192_n N_VGND_c_1276_n 0.0338116f $X=2.84 $Y=0.35 $X2=0
+ $Y2=0
cc_700 N_A_27_125#_c_1193_n N_VGND_c_1276_n 0.0114525f $X=2.17 $Y=0.35 $X2=0
+ $Y2=0
cc_701 N_A_27_125#_c_1194_n N_A_707_119#_c_1378_n 0.0372071f $X=3.005 $Y=0.77
+ $X2=0 $Y2=0
cc_702 N_A_27_125#_c_1192_n N_A_707_119#_c_1380_n 0.00679393f $X=2.84 $Y=0.35
+ $X2=0 $Y2=0
cc_703 N_A_27_125#_c_1194_n N_A_707_119#_c_1380_n 0.00265323f $X=3.005 $Y=0.77
+ $X2=0 $Y2=0
cc_704 N_VGND_c_1254_n N_A_707_119#_c_1379_n 0.0142636f $X=5.115 $Y=0.74 $X2=0
+ $Y2=0
cc_705 N_VGND_c_1270_n N_A_707_119#_c_1379_n 0.048346f $X=4.95 $Y=0 $X2=0 $Y2=0
cc_706 N_VGND_c_1276_n N_A_707_119#_c_1379_n 0.0326371f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_707 N_VGND_c_1270_n N_A_707_119#_c_1380_n 0.0134803f $X=4.95 $Y=0 $X2=0 $Y2=0
cc_708 N_VGND_c_1276_n N_A_707_119#_c_1380_n 0.00875888f $X=9.84 $Y=0 $X2=0
+ $Y2=0
cc_709 N_VGND_c_1254_n N_A_707_119#_c_1381_n 0.0341802f $X=5.115 $Y=0.74 $X2=0
+ $Y2=0
cc_710 N_VGND_c_1254_n N_A_707_119#_c_1382_n 0.0263226f $X=5.115 $Y=0.74 $X2=0
+ $Y2=0
cc_711 N_VGND_c_1254_n N_A_707_119#_c_1384_n 0.025828f $X=5.115 $Y=0.74 $X2=0
+ $Y2=0
cc_712 N_VGND_c_1255_n N_A_707_119#_c_1384_n 0.00571886f $X=5.92 $Y=0 $X2=0
+ $Y2=0
cc_713 N_VGND_c_1256_n N_A_707_119#_c_1384_n 0.0382129f $X=6.085 $Y=0.515 $X2=0
+ $Y2=0
cc_714 N_VGND_c_1276_n N_A_707_119#_c_1384_n 0.00786368f $X=9.84 $Y=0 $X2=0
+ $Y2=0
