* File: sky130_fd_sc_ls__o211a_4.pex.spice
* Created: Wed Sep  2 11:17:26 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__O211A_4%A_91_48# 1 2 3 4 15 17 19 22 24 26 29 31 33
+ 36 38 40 41 50 51 52 55 57 62 63 68 70 75 77 86
c175 86 0 1.89035e-19 $X=1.89 $Y=1.532
c176 77 0 5.28046e-20 $X=5.49 $Y=2.115
c177 57 0 8.88359e-21 $X=3.95 $Y=1.195
c178 36 0 1.6164e-19 $X=1.89 $Y=0.74
r179 86 87 14.2861 $w=3.88e-07 $l=1.15e-07 $layer=POLY_cond $X=1.89 $Y=1.532
+ $X2=2.005 $Y2=1.532
r180 83 84 11.8015 $w=3.88e-07 $l=9.5e-08 $layer=POLY_cond $X=1.46 $Y=1.532
+ $X2=1.555 $Y2=1.532
r181 82 83 56.5232 $w=3.88e-07 $l=4.55e-07 $layer=POLY_cond $X=1.005 $Y=1.532
+ $X2=1.46 $Y2=1.532
r182 81 82 5.59021 $w=3.88e-07 $l=4.5e-08 $layer=POLY_cond $X=0.96 $Y=1.532
+ $X2=1.005 $Y2=1.532
r183 78 79 3.10567 $w=3.88e-07 $l=2.5e-08 $layer=POLY_cond $X=0.53 $Y=1.532
+ $X2=0.555 $Y2=1.532
r184 70 72 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=3.555 $Y=1.105
+ $X2=3.555 $Y2=1.195
r185 64 75 4.30018 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.12 $Y=2.035
+ $X2=3.955 $Y2=2.035
r186 63 77 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.325 $Y=2.035
+ $X2=5.49 $Y2=2.035
r187 63 64 78.615 $w=1.68e-07 $l=1.205e-06 $layer=LI1_cond $X=5.325 $Y=2.035
+ $X2=4.12 $Y2=2.035
r188 62 75 1.96316 $w=1.7e-07 $l=1.18427e-07 $layer=LI1_cond $X=4.035 $Y=1.95
+ $X2=3.955 $Y2=2.035
r189 61 62 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.035 $Y=1.28
+ $X2=4.035 $Y2=1.95
r190 58 72 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.72 $Y=1.195
+ $X2=3.555 $Y2=1.195
r191 57 61 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.95 $Y=1.195
+ $X2=4.035 $Y2=1.28
r192 57 58 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=3.95 $Y=1.195
+ $X2=3.72 $Y2=1.195
r193 56 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.105 $Y=2.035
+ $X2=2.94 $Y2=2.035
r194 55 75 4.30018 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.79 $Y=2.035
+ $X2=3.955 $Y2=2.035
r195 55 56 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=3.79 $Y=2.035
+ $X2=3.105 $Y2=2.035
r196 51 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.775 $Y=2.035
+ $X2=2.94 $Y2=2.035
r197 51 52 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=2.775 $Y=2.035
+ $X2=2.285 $Y2=2.035
r198 50 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.2 $Y=1.95
+ $X2=2.285 $Y2=2.035
r199 49 50 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2.2 $Y=1.63 $X2=2.2
+ $Y2=1.95
r200 48 86 11.1804 $w=3.88e-07 $l=9e-08 $layer=POLY_cond $X=1.8 $Y=1.532
+ $X2=1.89 $Y2=1.532
r201 48 84 30.4356 $w=3.88e-07 $l=2.45e-07 $layer=POLY_cond $X=1.8 $Y=1.532
+ $X2=1.555 $Y2=1.532
r202 47 48 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.8
+ $Y=1.465 $X2=1.8 $Y2=1.465
r203 44 81 22.3608 $w=3.88e-07 $l=1.8e-07 $layer=POLY_cond $X=0.78 $Y=1.532
+ $X2=0.96 $Y2=1.532
r204 44 79 27.951 $w=3.88e-07 $l=2.25e-07 $layer=POLY_cond $X=0.78 $Y=1.532
+ $X2=0.555 $Y2=1.532
r205 43 47 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=0.78 $Y=1.465
+ $X2=1.8 $Y2=1.465
r206 43 44 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.78
+ $Y=1.465 $X2=0.78 $Y2=1.465
r207 41 49 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.115 $Y=1.465
+ $X2=2.2 $Y2=1.63
r208 41 47 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=2.115 $Y=1.465
+ $X2=1.8 $Y2=1.465
r209 38 87 25.1189 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=2.005 $Y=1.765
+ $X2=2.005 $Y2=1.532
r210 38 40 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.005 $Y=1.765
+ $X2=2.005 $Y2=2.4
r211 34 86 25.1189 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=1.89 $Y=1.3
+ $X2=1.89 $Y2=1.532
r212 34 36 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.89 $Y=1.3
+ $X2=1.89 $Y2=0.74
r213 31 84 25.1189 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=1.555 $Y=1.765
+ $X2=1.555 $Y2=1.532
r214 31 33 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.555 $Y=1.765
+ $X2=1.555 $Y2=2.4
r215 27 83 25.1189 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=1.46 $Y=1.3
+ $X2=1.46 $Y2=1.532
r216 27 29 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.46 $Y=1.3
+ $X2=1.46 $Y2=0.74
r217 24 82 25.1189 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=1.005 $Y=1.765
+ $X2=1.005 $Y2=1.532
r218 24 26 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.005 $Y=1.765
+ $X2=1.005 $Y2=2.4
r219 20 81 25.1189 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=0.96 $Y=1.3
+ $X2=0.96 $Y2=1.532
r220 20 22 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.96 $Y=1.3
+ $X2=0.96 $Y2=0.74
r221 17 79 25.1189 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=0.555 $Y=1.765
+ $X2=0.555 $Y2=1.532
r222 17 19 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.555 $Y=1.765
+ $X2=0.555 $Y2=2.4
r223 13 78 25.1189 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=0.53 $Y=1.3
+ $X2=0.53 $Y2=1.532
r224 13 15 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.53 $Y=1.3
+ $X2=0.53 $Y2=0.74
r225 4 77 300 $w=1.7e-07 $l=2.68328e-07 $layer=licon1_PDIFF $count=2 $X=5.29
+ $Y=1.955 $X2=5.49 $Y2=2.115
r226 3 75 300 $w=1.7e-07 $l=2.22711e-07 $layer=licon1_PDIFF $count=2 $X=3.805
+ $Y=1.955 $X2=3.955 $Y2=2.115
r227 2 68 300 $w=1.7e-07 $l=2.22711e-07 $layer=licon1_PDIFF $count=2 $X=2.79
+ $Y=1.955 $X2=2.94 $Y2=2.115
r228 1 70 182 $w=1.7e-07 $l=5.45527e-07 $layer=licon1_NDIFF $count=1 $X=3.415
+ $Y=0.625 $X2=3.555 $Y2=1.105
.ends

.subckt PM_SKY130_FD_SC_LS__O211A_4%C1 1 3 6 8 10 13 15 22
c53 6 0 8.88359e-21 $X=3.34 $Y=0.945
r54 22 23 5.35556 $w=3.6e-07 $l=4e-08 $layer=POLY_cond $X=3.73 $Y=1.665 $X2=3.77
+ $Y2=1.665
r55 20 22 15.3972 $w=3.6e-07 $l=1.15e-07 $layer=POLY_cond $X=3.615 $Y=1.665
+ $X2=3.73 $Y2=1.665
r56 18 20 36.8194 $w=3.6e-07 $l=2.75e-07 $layer=POLY_cond $X=3.34 $Y=1.665
+ $X2=3.615 $Y2=1.665
r57 15 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.615
+ $Y=1.615 $X2=3.615 $Y2=1.615
r58 11 23 23.3057 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=3.77 $Y=1.45
+ $X2=3.77 $Y2=1.665
r59 11 13 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=3.77 $Y=1.45
+ $X2=3.77 $Y2=0.945
r60 8 22 23.3057 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=3.73 $Y=1.88
+ $X2=3.73 $Y2=1.665
r61 8 10 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=3.73 $Y=1.88 $X2=3.73
+ $Y2=2.375
r62 4 18 23.3057 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=3.34 $Y=1.45
+ $X2=3.34 $Y2=1.665
r63 4 6 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=3.34 $Y=1.45 $X2=3.34
+ $Y2=0.945
r64 1 18 23.4306 $w=3.6e-07 $l=2.89569e-07 $layer=POLY_cond $X=3.165 $Y=1.88
+ $X2=3.34 $Y2=1.665
r65 1 3 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=3.165 $Y=1.88
+ $X2=3.165 $Y2=2.375
.ends

.subckt PM_SKY130_FD_SC_LS__O211A_4%B1 2 3 4 5 7 8 10 12 13 15 19 21 22 28
c84 22 0 1.89035e-19 $X=2.64 $Y=1.665
c85 19 0 2.18884e-20 $X=4.27 $Y=0.945
c86 5 0 2.31478e-20 $X=2.715 $Y=1.88
r87 26 28 5.51908 $w=3.93e-07 $l=4.5e-08 $layer=POLY_cond $X=2.67 $Y=1.61
+ $X2=2.715 $Y2=1.61
r88 24 26 33.1145 $w=3.93e-07 $l=2.7e-07 $layer=POLY_cond $X=2.4 $Y=1.61
+ $X2=2.67 $Y2=1.61
r89 22 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.67
+ $Y=1.6 $X2=2.67 $Y2=1.6
r90 20 21 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=4.217 $Y=1.34
+ $X2=4.217 $Y2=1.49
r91 19 20 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=4.27 $Y=0.945
+ $X2=4.27 $Y2=1.34
r92 16 19 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.27 $Y=0.255
+ $X2=4.27 $Y2=0.945
r93 13 15 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=4.18 $Y=1.88
+ $X2=4.18 $Y2=2.375
r94 12 13 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=4.18 $Y=1.79 $X2=4.18
+ $Y2=1.88
r95 12 21 116.613 $w=1.8e-07 $l=3e-07 $layer=POLY_cond $X=4.18 $Y=1.79 $X2=4.18
+ $Y2=1.49
r96 8 28 23.916 $w=3.93e-07 $l=3.5433e-07 $layer=POLY_cond $X=2.91 $Y=1.34
+ $X2=2.715 $Y2=1.61
r97 8 10 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.91 $Y=1.34
+ $X2=2.91 $Y2=0.945
r98 5 28 25.4309 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.715 $Y=1.88
+ $X2=2.715 $Y2=1.61
r99 5 7 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.715 $Y=1.88
+ $X2=2.715 $Y2=2.375
r100 3 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.195 $Y=0.18
+ $X2=4.27 $Y2=0.255
r101 3 4 881.957 $w=1.5e-07 $l=1.72e-06 $layer=POLY_cond $X=4.195 $Y=0.18
+ $X2=2.475 $Y2=0.18
r102 2 24 25.4309 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.4 $Y=1.34 $X2=2.4
+ $Y2=1.61
r103 1 4 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.4 $Y=0.255
+ $X2=2.475 $Y2=0.18
r104 1 2 556.351 $w=1.5e-07 $l=1.085e-06 $layer=POLY_cond $X=2.4 $Y=0.255
+ $X2=2.4 $Y2=1.34
.ends

.subckt PM_SKY130_FD_SC_LS__O211A_4%A2 1 3 6 8 10 13 15 16 23 24
c51 24 0 1.8255e-19 $X=5.715 $Y=1.665
c52 13 0 1.59181e-19 $X=5.725 $Y=0.945
c53 6 0 1.64451e-19 $X=5.24 $Y=0.945
r54 24 25 1.3027 $w=3.7e-07 $l=1e-08 $layer=POLY_cond $X=5.715 $Y=1.665
+ $X2=5.725 $Y2=1.665
r55 22 24 5.86216 $w=3.7e-07 $l=4.5e-08 $layer=POLY_cond $X=5.67 $Y=1.665
+ $X2=5.715 $Y2=1.665
r56 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.67
+ $Y=1.615 $X2=5.67 $Y2=1.615
r57 20 22 56.0162 $w=3.7e-07 $l=4.3e-07 $layer=POLY_cond $X=5.24 $Y=1.665
+ $X2=5.67 $Y2=1.665
r58 19 20 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=5.215 $Y=1.665
+ $X2=5.24 $Y2=1.665
r59 16 23 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=5.52 $Y=1.615
+ $X2=5.67 $Y2=1.615
r60 15 16 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=5.04 $Y=1.615
+ $X2=5.52 $Y2=1.615
r61 11 25 23.9667 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=5.725 $Y=1.45
+ $X2=5.725 $Y2=1.665
r62 11 13 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=5.725 $Y=1.45
+ $X2=5.725 $Y2=0.945
r63 8 24 23.9667 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=5.715 $Y=1.88
+ $X2=5.715 $Y2=1.665
r64 8 10 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.715 $Y=1.88
+ $X2=5.715 $Y2=2.455
r65 4 20 23.9667 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=5.24 $Y=1.45
+ $X2=5.24 $Y2=1.665
r66 4 6 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=5.24 $Y=1.45 $X2=5.24
+ $Y2=0.945
r67 1 19 23.9667 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=5.215 $Y=1.88
+ $X2=5.215 $Y2=1.665
r68 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.215 $Y=1.88
+ $X2=5.215 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_LS__O211A_4%A1 1 2 3 5 9 10 11 12 14 18 20
c65 12 0 5.28046e-20 $X=6.165 $Y=1.88
c66 9 0 1.33941e-19 $X=4.78 $Y=0.945
r67 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.24
+ $Y=1.615 $X2=6.24 $Y2=1.615
r68 20 24 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=6.48 $Y=1.615
+ $X2=6.24 $Y2=1.615
r69 16 23 38.578 $w=2.95e-07 $l=1.72337e-07 $layer=POLY_cond $X=6.225 $Y=1.45
+ $X2=6.24 $Y2=1.615
r70 16 18 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=6.225 $Y=1.45
+ $X2=6.225 $Y2=0.945
r71 15 18 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.225 $Y=0.255
+ $X2=6.225 $Y2=0.945
r72 12 23 54.9169 $w=2.95e-07 $l=3.00167e-07 $layer=POLY_cond $X=6.165 $Y=1.88
+ $X2=6.24 $Y2=1.615
r73 12 14 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.165 $Y=1.88
+ $X2=6.165 $Y2=2.455
r74 10 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.15 $Y=0.18
+ $X2=6.225 $Y2=0.255
r75 10 11 664.032 $w=1.5e-07 $l=1.295e-06 $layer=POLY_cond $X=6.15 $Y=0.18
+ $X2=4.855 $Y2=0.18
r76 9 19 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=4.78 $Y=0.945
+ $X2=4.78 $Y2=1.34
r77 6 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.78 $Y=0.255
+ $X2=4.855 $Y2=0.18
r78 6 9 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.78 $Y=0.255 $X2=4.78
+ $Y2=0.945
r79 3 5 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=4.765 $Y=1.88
+ $X2=4.765 $Y2=2.455
r80 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=4.765 $Y=1.79 $X2=4.765
+ $Y2=1.88
r81 1 19 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=4.765 $Y=1.43 $X2=4.765
+ $Y2=1.34
r82 1 2 139.935 $w=1.8e-07 $l=3.6e-07 $layer=POLY_cond $X=4.765 $Y=1.43
+ $X2=4.765 $Y2=1.79
.ends

.subckt PM_SKY130_FD_SC_LS__O211A_4%VPWR 1 2 3 4 5 6 19 21 25 27 31 37 41 45 47
+ 52 53 54 56 65 69 81 84 87 91
r93 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r94 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r95 84 85 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r96 82 85 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r97 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r98 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r99 76 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r100 75 76 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r101 73 76 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33 $X2=6
+ $Y2=3.33
r102 73 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r103 72 75 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=5.04 $Y=3.33 $X2=6
+ $Y2=3.33
r104 72 73 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r105 70 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.655 $Y=3.33
+ $X2=4.49 $Y2=3.33
r106 70 72 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=4.655 $Y=3.33
+ $X2=5.04 $Y2=3.33
r107 69 90 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=6.275 $Y=3.33
+ $X2=6.497 $Y2=3.33
r108 69 75 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.275 $Y=3.33
+ $X2=6 $Y2=3.33
r109 68 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r110 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r111 65 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.325 $Y=3.33
+ $X2=4.49 $Y2=3.33
r112 65 67 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=4.325 $Y=3.33
+ $X2=4.08 $Y2=3.33
r113 64 85 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.16 $Y2=3.33
r114 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r115 61 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.445 $Y=3.33
+ $X2=2.28 $Y2=3.33
r116 61 63 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=2.445 $Y=3.33
+ $X2=3.12 $Y2=3.33
r117 60 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r118 60 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r119 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r120 57 78 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.222 $Y2=3.33
r121 57 59 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.72 $Y2=3.33
r122 56 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.115 $Y=3.33
+ $X2=1.28 $Y2=3.33
r123 56 59 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.115 $Y=3.33
+ $X2=0.72 $Y2=3.33
r124 54 68 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=4.08 $Y2=3.33
r125 54 64 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=3.12 $Y2=3.33
r126 52 63 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=3.275 $Y=3.33
+ $X2=3.12 $Y2=3.33
r127 52 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.275 $Y=3.33
+ $X2=3.44 $Y2=3.33
r128 51 67 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=3.605 $Y=3.33
+ $X2=4.08 $Y2=3.33
r129 51 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.605 $Y=3.33
+ $X2=3.44 $Y2=3.33
r130 47 50 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=6.44 $Y=2.115
+ $X2=6.44 $Y2=2.81
r131 45 90 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=6.44 $Y=3.245
+ $X2=6.497 $Y2=3.33
r132 45 50 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=6.44 $Y=3.245
+ $X2=6.44 $Y2=2.81
r133 41 44 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=4.49 $Y=2.41 $X2=4.49
+ $Y2=2.81
r134 39 87 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.49 $Y=3.245
+ $X2=4.49 $Y2=3.33
r135 39 44 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=4.49 $Y=3.245
+ $X2=4.49 $Y2=2.81
r136 35 53 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.44 $Y=3.245
+ $X2=3.44 $Y2=3.33
r137 35 37 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=3.44 $Y=3.245
+ $X2=3.44 $Y2=2.455
r138 31 34 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=2.28 $Y=2.405
+ $X2=2.28 $Y2=2.815
r139 29 84 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.28 $Y=3.245
+ $X2=2.28 $Y2=3.33
r140 29 34 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.28 $Y=3.245
+ $X2=2.28 $Y2=2.815
r141 28 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.445 $Y=3.33
+ $X2=1.28 $Y2=3.33
r142 27 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.115 $Y=3.33
+ $X2=2.28 $Y2=3.33
r143 27 28 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.115 $Y=3.33
+ $X2=1.445 $Y2=3.33
r144 23 81 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.28 $Y=3.245
+ $X2=1.28 $Y2=3.33
r145 23 25 32.8272 $w=3.28e-07 $l=9.4e-07 $layer=LI1_cond $X=1.28 $Y=3.245
+ $X2=1.28 $Y2=2.305
r146 19 78 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.222 $Y2=3.33
r147 19 21 32.8272 $w=3.28e-07 $l=9.4e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.28 $Y2=2.305
r148 6 50 400 $w=1.7e-07 $l=9.4975e-07 $layer=licon1_PDIFF $count=1 $X=6.24
+ $Y=1.955 $X2=6.44 $Y2=2.81
r149 6 47 400 $w=1.7e-07 $l=2.68328e-07 $layer=licon1_PDIFF $count=1 $X=6.24
+ $Y=1.955 $X2=6.44 $Y2=2.115
r150 5 44 600 $w=1.7e-07 $l=9.65376e-07 $layer=licon1_PDIFF $count=1 $X=4.255
+ $Y=1.955 $X2=4.49 $Y2=2.81
r151 5 41 600 $w=1.7e-07 $l=5.60312e-07 $layer=licon1_PDIFF $count=1 $X=4.255
+ $Y=1.955 $X2=4.49 $Y2=2.41
r152 4 37 600 $w=1.7e-07 $l=5.91608e-07 $layer=licon1_PDIFF $count=1 $X=3.24
+ $Y=1.955 $X2=3.44 $Y2=2.455
r153 3 34 600 $w=1.7e-07 $l=1.07034e-06 $layer=licon1_PDIFF $count=1 $X=2.08
+ $Y=1.84 $X2=2.28 $Y2=2.815
r154 3 31 600 $w=1.7e-07 $l=6.57438e-07 $layer=licon1_PDIFF $count=1 $X=2.08
+ $Y=1.84 $X2=2.28 $Y2=2.405
r155 2 25 300 $w=1.7e-07 $l=5.5608e-07 $layer=licon1_PDIFF $count=2 $X=1.08
+ $Y=1.84 $X2=1.28 $Y2=2.305
r156 1 21 300 $w=1.7e-07 $l=5.32588e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.305
.ends

.subckt PM_SKY130_FD_SC_LS__O211A_4%X 1 2 3 4 13 14 15 16 19 23 27 29 33 37 43
+ 44 45 46
c79 29 0 2.31478e-20 $X=1.615 $Y=1.885
c80 27 0 1.6164e-19 $X=1.51 $Y=1.045
r81 45 46 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=1.295
+ $X2=0.24 $Y2=1.665
r82 42 46 6.76434 $w=2.28e-07 $l=1.35e-07 $layer=LI1_cond $X=0.24 $Y=1.8
+ $X2=0.24 $Y2=1.665
r83 41 45 8.26753 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.24 $Y=1.13
+ $X2=0.24 $Y2=1.295
r84 37 39 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=1.78 $Y=1.985
+ $X2=1.78 $Y2=2.815
r85 35 37 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=1.78 $Y=1.97
+ $X2=1.78 $Y2=1.985
r86 31 33 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=1.635 $Y=0.96
+ $X2=1.635 $Y2=0.515
r87 30 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=1.885
+ $X2=0.78 $Y2=1.885
r88 29 35 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.615 $Y=1.885
+ $X2=1.78 $Y2=1.97
r89 29 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.615 $Y=1.885
+ $X2=0.945 $Y2=1.885
r90 28 43 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.83 $Y=1.045
+ $X2=0.705 $Y2=1.045
r91 27 31 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.51 $Y=1.045
+ $X2=1.635 $Y2=0.96
r92 27 28 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.51 $Y=1.045
+ $X2=0.83 $Y2=1.045
r93 23 25 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=0.78 $Y=1.985
+ $X2=0.78 $Y2=2.815
r94 21 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=1.97 $X2=0.78
+ $Y2=1.885
r95 21 23 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=0.78 $Y=1.97
+ $X2=0.78 $Y2=1.985
r96 17 43 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=0.96
+ $X2=0.705 $Y2=1.045
r97 17 19 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=0.705 $Y=0.96
+ $X2=0.705 $Y2=0.515
r98 16 42 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.355 $Y=1.885
+ $X2=0.24 $Y2=1.8
r99 15 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=1.885
+ $X2=0.78 $Y2=1.885
r100 15 16 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.615 $Y=1.885
+ $X2=0.355 $Y2=1.885
r101 14 41 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.355 $Y=1.045
+ $X2=0.24 $Y2=1.13
r102 13 43 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.58 $Y=1.045
+ $X2=0.705 $Y2=1.045
r103 13 14 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.58 $Y=1.045
+ $X2=0.355 $Y2=1.045
r104 4 39 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.63
+ $Y=1.84 $X2=1.78 $Y2=2.815
r105 4 37 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.63
+ $Y=1.84 $X2=1.78 $Y2=1.985
r106 3 25 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=0.63
+ $Y=1.84 $X2=0.78 $Y2=2.815
r107 3 23 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=0.63
+ $Y=1.84 $X2=0.78 $Y2=1.985
r108 2 33 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.535
+ $Y=0.37 $X2=1.675 $Y2=0.515
r109 1 19 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.605
+ $Y=0.37 $X2=0.745 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__O211A_4%A_968_391# 1 2 9 11 12 15
r27 15 18 32.0379 $w=2.48e-07 $l=6.95e-07 $layer=LI1_cond $X=5.98 $Y=2.115
+ $X2=5.98 $Y2=2.81
r28 13 18 4.37928 $w=2.48e-07 $l=9.5e-08 $layer=LI1_cond $X=5.98 $Y=2.905
+ $X2=5.98 $Y2=2.81
r29 11 13 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.855 $Y=2.99
+ $X2=5.98 $Y2=2.905
r30 11 12 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=5.855 $Y=2.99
+ $X2=5.155 $Y2=2.99
r31 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.99 $Y=2.905
+ $X2=5.155 $Y2=2.99
r32 7 9 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=4.99 $Y=2.905
+ $X2=4.99 $Y2=2.41
r33 2 18 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=5.79
+ $Y=1.955 $X2=5.94 $Y2=2.81
r34 2 15 400 $w=1.7e-07 $l=2.22711e-07 $layer=licon1_PDIFF $count=1 $X=5.79
+ $Y=1.955 $X2=5.94 $Y2=2.115
r35 1 9 300 $w=1.7e-07 $l=5.24667e-07 $layer=licon1_PDIFF $count=2 $X=4.84
+ $Y=1.955 $X2=4.99 $Y2=2.41
.ends

.subckt PM_SKY130_FD_SC_LS__O211A_4%VGND 1 2 3 4 5 16 18 22 26 30 34 36 38 43 48
+ 56 63 64 70 73 76 79
r88 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r89 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r90 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r91 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r92 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r93 64 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r94 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r95 61 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.105 $Y=0 $X2=5.94
+ $Y2=0
r96 61 63 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=6.105 $Y=0 $X2=6.48
+ $Y2=0
r97 60 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r98 60 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r99 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r100 57 76 8.88104 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=5.175 $Y=0
+ $X2=5.002 $Y2=0
r101 57 59 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=5.175 $Y=0 $X2=5.52
+ $Y2=0
r102 56 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.775 $Y=0 $X2=5.94
+ $Y2=0
r103 56 59 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=5.775 $Y=0
+ $X2=5.52 $Y2=0
r104 55 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r105 54 55 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r106 52 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r107 51 54 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=2.64 $Y=0 $X2=4.56
+ $Y2=0
r108 51 52 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r109 49 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.27 $Y=0 $X2=2.105
+ $Y2=0
r110 49 51 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.27 $Y=0 $X2=2.64
+ $Y2=0
r111 48 76 8.88104 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=4.83 $Y=0 $X2=5.002
+ $Y2=0
r112 48 54 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=4.83 $Y=0 $X2=4.56
+ $Y2=0
r113 47 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r114 47 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r115 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r116 44 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.34 $Y=0 $X2=1.175
+ $Y2=0
r117 44 46 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.34 $Y=0 $X2=1.68
+ $Y2=0
r118 43 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.94 $Y=0 $X2=2.105
+ $Y2=0
r119 43 46 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=1.94 $Y=0 $X2=1.68
+ $Y2=0
r120 42 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r121 42 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r122 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r123 39 67 3.96842 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=0.4 $Y=0 $X2=0.2 $Y2=0
r124 39 41 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.4 $Y=0 $X2=0.72
+ $Y2=0
r125 38 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.01 $Y=0 $X2=1.175
+ $Y2=0
r126 38 41 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.01 $Y=0 $X2=0.72
+ $Y2=0
r127 36 55 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=3.36 $Y=0 $X2=4.56
+ $Y2=0
r128 36 52 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.36 $Y=0 $X2=2.64
+ $Y2=0
r129 32 79 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.94 $Y=0.085
+ $X2=5.94 $Y2=0
r130 32 34 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=5.94 $Y=0.085
+ $X2=5.94 $Y2=0.77
r131 28 76 1.03204 $w=3.45e-07 $l=8.5e-08 $layer=LI1_cond $X=5.002 $Y=0.085
+ $X2=5.002 $Y2=0
r132 28 30 22.8818 $w=3.43e-07 $l=6.85e-07 $layer=LI1_cond $X=5.002 $Y=0.085
+ $X2=5.002 $Y2=0.77
r133 24 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.105 $Y=0.085
+ $X2=2.105 $Y2=0
r134 24 26 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.105 $Y=0.085
+ $X2=2.105 $Y2=0.515
r135 20 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.175 $Y=0.085
+ $X2=1.175 $Y2=0
r136 20 22 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=1.175 $Y=0.085
+ $X2=1.175 $Y2=0.57
r137 16 67 3.17474 $w=2.5e-07 $l=1.16619e-07 $layer=LI1_cond $X=0.275 $Y=0.085
+ $X2=0.2 $Y2=0
r138 16 18 22.3574 $w=2.48e-07 $l=4.85e-07 $layer=LI1_cond $X=0.275 $Y=0.085
+ $X2=0.275 $Y2=0.57
r139 5 34 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=5.8
+ $Y=0.625 $X2=5.94 $Y2=0.77
r140 4 30 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=4.855
+ $Y=0.625 $X2=5 $Y2=0.77
r141 3 26 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.965
+ $Y=0.37 $X2=2.105 $Y2=0.515
r142 2 22 182 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=1 $X=1.035
+ $Y=0.37 $X2=1.175 $Y2=0.57
r143 1 18 182 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_NDIFF $count=1 $X=0.17
+ $Y=0.37 $X2=0.315 $Y2=0.57
.ends

.subckt PM_SKY130_FD_SC_LS__O211A_4%A_510_125# 1 2 3 4 15 17 18 22 23 24 27 29
+ 33 35
c72 27 0 3.23633e-19 $X=5.51 $Y=0.77
c73 24 0 1.33941e-19 $X=4.65 $Y=1.195
c74 23 0 1.8255e-19 $X=5.345 $Y=1.195
r75 31 33 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=6.44 $Y=1.11
+ $X2=6.44 $Y2=0.77
r76 30 35 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.595 $Y=1.195
+ $X2=5.47 $Y2=1.195
r77 29 31 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.275 $Y=1.195
+ $X2=6.44 $Y2=1.11
r78 29 30 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=6.275 $Y=1.195
+ $X2=5.595 $Y2=1.195
r79 25 35 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.47 $Y=1.11
+ $X2=5.47 $Y2=1.195
r80 25 27 15.6732 $w=2.48e-07 $l=3.4e-07 $layer=LI1_cond $X=5.47 $Y=1.11
+ $X2=5.47 $Y2=0.77
r81 23 35 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.345 $Y=1.195
+ $X2=5.47 $Y2=1.195
r82 23 24 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=5.345 $Y=1.195
+ $X2=4.65 $Y2=1.195
r83 20 24 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.525 $Y=1.11
+ $X2=4.65 $Y2=1.195
r84 20 22 15.6732 $w=2.48e-07 $l=3.4e-07 $layer=LI1_cond $X=4.525 $Y=1.11
+ $X2=4.525 $Y2=0.77
r85 19 22 15.9037 $w=2.48e-07 $l=3.45e-07 $layer=LI1_cond $X=4.525 $Y=0.425
+ $X2=4.525 $Y2=0.77
r86 17 19 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.4 $Y=0.34
+ $X2=4.525 $Y2=0.425
r87 17 18 105.69 $w=1.68e-07 $l=1.62e-06 $layer=LI1_cond $X=4.4 $Y=0.34 $X2=2.78
+ $Y2=0.34
r88 13 18 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.655 $Y=0.425
+ $X2=2.78 $Y2=0.34
r89 13 15 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=2.655 $Y=0.425
+ $X2=2.655 $Y2=0.76
r90 4 33 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.3
+ $Y=0.625 $X2=6.44 $Y2=0.77
r91 3 27 91 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_NDIFF $count=2 $X=5.315
+ $Y=0.625 $X2=5.51 $Y2=0.77
r92 2 22 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.345
+ $Y=0.625 $X2=4.485 $Y2=0.77
r93 1 15 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=2.55
+ $Y=0.625 $X2=2.695 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_LS__O211A_4%A_597_125# 1 2 9 11 12 13
c26 11 0 2.18884e-20 $X=3.89 $Y=0.68
r27 13 16 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=4.055 $Y=0.68
+ $X2=4.055 $Y2=0.77
r28 11 13 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.89 $Y=0.68
+ $X2=4.055 $Y2=0.68
r29 11 12 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.89 $Y=0.68
+ $X2=3.21 $Y2=0.68
r30 7 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.125 $Y=0.765
+ $X2=3.21 $Y2=0.68
r31 7 9 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=3.125 $Y=0.765
+ $X2=3.125 $Y2=0.77
r32 2 16 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=3.845
+ $Y=0.625 $X2=4.055 $Y2=0.77
r33 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.985
+ $Y=0.625 $X2=3.125 $Y2=0.77
.ends

