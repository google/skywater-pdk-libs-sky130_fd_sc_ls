* File: sky130_fd_sc_ls__a211o_1.pex.spice
* Created: Fri Aug 28 12:48:55 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__A211O_1%A_81_264# 1 2 3 10 12 15 17 18 19 24 26 28
+ 30 34 39
c80 26 0 3.92783e-20 $X=3.125 $Y=1.18
c81 24 0 1.62677e-19 $X=2.28 $Y=1.195
c82 18 0 1.71301e-19 $X=1.13 $Y=1.485
c83 10 0 1.55122e-19 $X=0.495 $Y=1.765
r84 41 42 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=2.445 $Y=1.18
+ $X2=2.445 $Y2=1.195
r85 39 41 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=2.445 $Y=1.02
+ $X2=2.445 $Y2=1.18
r86 30 32 19.7165 $w=4.13e-07 $l=7.1e-07 $layer=LI1_cond $X=3.332 $Y=2.105
+ $X2=3.332 $Y2=2.815
r87 28 45 2.59301 $w=4.15e-07 $l=1e-07 $layer=LI1_cond $X=3.332 $Y=1.28
+ $X2=3.332 $Y2=1.18
r88 28 30 22.91 $w=4.13e-07 $l=8.25e-07 $layer=LI1_cond $X=3.332 $Y=1.28
+ $X2=3.332 $Y2=2.105
r89 27 41 3.66692 $w=2e-07 $l=1.65e-07 $layer=LI1_cond $X=2.61 $Y=1.18 $X2=2.445
+ $Y2=1.18
r90 26 45 5.36752 $w=2e-07 $l=2.07e-07 $layer=LI1_cond $X=3.125 $Y=1.18
+ $X2=3.332 $Y2=1.18
r91 26 27 28.5591 $w=1.98e-07 $l=5.15e-07 $layer=LI1_cond $X=3.125 $Y=1.18
+ $X2=2.61 $Y2=1.18
r92 25 34 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.415 $Y=1.195
+ $X2=1.33 $Y2=1.195
r93 24 42 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.28 $Y=1.195
+ $X2=2.445 $Y2=1.195
r94 24 25 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=2.28 $Y=1.195
+ $X2=1.415 $Y2=1.195
r95 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.115
+ $Y=1.485 $X2=1.115 $Y2=1.485
r96 19 34 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.33 $Y=1.525
+ $X2=1.33 $Y2=1.195
r97 19 21 5.9927 $w=2.48e-07 $l=1.3e-07 $layer=LI1_cond $X=1.245 $Y=1.525
+ $X2=1.115 $Y2=1.525
r98 18 22 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.13 $Y=1.485
+ $X2=1.115 $Y2=1.485
r99 17 22 92.6765 $w=3.3e-07 $l=5.3e-07 $layer=POLY_cond $X=0.585 $Y=1.485
+ $X2=1.115 $Y2=1.485
r100 13 18 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=1.205 $Y=1.32
+ $X2=1.13 $Y2=1.485
r101 13 15 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.205 $Y=1.32
+ $X2=1.205 $Y2=0.74
r102 10 17 32.1775 $w=3.3e-07 $l=3.2187e-07 $layer=POLY_cond $X=0.495 $Y=1.765
+ $X2=0.585 $Y2=1.485
r103 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.495 $Y=1.765
+ $X2=0.495 $Y2=2.4
r104 3 32 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=3.14
+ $Y=1.96 $X2=3.29 $Y2=2.815
r105 3 30 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=3.14
+ $Y=1.96 $X2=3.29 $Y2=2.105
r106 2 45 182 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_NDIFF $count=1 $X=3.235
+ $Y=0.68 $X2=3.375 $Y2=1.17
r107 1 39 182 $w=1.7e-07 $l=4.0398e-07 $layer=licon1_NDIFF $count=1 $X=2.305
+ $Y=0.68 $X2=2.445 $Y2=1.02
.ends

.subckt PM_SKY130_FD_SC_LS__A211O_1%A2 1 3 6 8
c32 8 0 1.71301e-19 $X=1.68 $Y=1.665
r33 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.67
+ $Y=1.615 $X2=1.67 $Y2=1.615
r34 4 11 38.5916 $w=2.93e-07 $l=2.03101e-07 $layer=POLY_cond $X=1.755 $Y=1.45
+ $X2=1.67 $Y2=1.615
r35 4 6 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=1.755 $Y=1.45
+ $X2=1.755 $Y2=1
r36 1 11 55.8646 $w=2.93e-07 $l=3.05205e-07 $layer=POLY_cond $X=1.745 $Y=1.885
+ $X2=1.67 $Y2=1.615
r37 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.745 $Y=1.885
+ $X2=1.745 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_LS__A211O_1%A1 1 3 6 8 9
c39 6 0 3.92783e-20 $X=2.23 $Y=1
r40 8 9 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=2.16 $Y=1.615 $X2=2.64
+ $Y2=1.615
r41 8 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.21
+ $Y=1.615 $X2=2.21 $Y2=1.615
r42 4 13 38.5916 $w=2.93e-07 $l=1.74714e-07 $layer=POLY_cond $X=2.23 $Y=1.45
+ $X2=2.21 $Y2=1.615
r43 4 6 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=2.23 $Y=1.45 $X2=2.23
+ $Y2=1
r44 1 13 55.8646 $w=2.93e-07 $l=2.77399e-07 $layer=POLY_cond $X=2.225 $Y=1.885
+ $X2=2.21 $Y2=1.615
r45 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.225 $Y=1.885
+ $X2=2.225 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_LS__A211O_1%B1 4 5 6 7 9 13 14 16 24
c47 13 0 1.23467e-19 $X=2.71 $Y=0.405
c48 4 0 3.92096e-20 $X=2.66 $Y=1
r49 16 24 3.89033 $w=4.13e-07 $l=1.15e-07 $layer=LI1_cond $X=2.16 $Y=0.462
+ $X2=2.275 $Y2=0.462
r50 14 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.71 $Y=0.405
+ $X2=2.71 $Y2=0.57
r51 13 24 15.9147 $w=3.13e-07 $l=4.35e-07 $layer=LI1_cond $X=2.71 $Y=0.412
+ $X2=2.275 $Y2=0.412
r52 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.71
+ $Y=0.405 $X2=2.71 $Y2=0.405
r53 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.675 $Y=1.885
+ $X2=2.675 $Y2=2.46
r54 6 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.675 $Y=1.795 $X2=2.675
+ $Y2=1.885
r55 5 10 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.675 $Y=1.485
+ $X2=2.675 $Y2=1.395
r56 5 6 120.5 $w=1.8e-07 $l=3.1e-07 $layer=POLY_cond $X=2.675 $Y=1.485 $X2=2.675
+ $Y2=1.795
r57 4 10 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.66 $Y=1 $X2=2.66
+ $Y2=1.395
r58 4 20 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.66 $Y=1 $X2=2.66
+ $Y2=0.57
.ends

.subckt PM_SKY130_FD_SC_LS__A211O_1%C1 2 3 5 9 11 12 13 16 17
r38 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.55
+ $Y=0.405 $X2=3.55 $Y2=0.405
r39 13 17 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=3.55 $Y=0.555
+ $X2=3.55 $Y2=0.405
r40 12 16 55.0813 $w=3.3e-07 $l=3.15e-07 $layer=POLY_cond $X=3.235 $Y=0.405
+ $X2=3.55 $Y2=0.405
r41 10 11 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=3.105 $Y=1.395
+ $X2=3.105 $Y2=1.545
r42 9 10 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.16 $Y=1 $X2=3.16
+ $Y2=1.395
r43 6 12 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=3.16 $Y=0.57
+ $X2=3.235 $Y2=0.405
r44 6 9 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.16 $Y=0.57 $X2=3.16
+ $Y2=1
r45 3 5 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.065 $Y=1.885
+ $X2=3.065 $Y2=2.46
r46 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.065 $Y=1.795 $X2=3.065
+ $Y2=1.885
r47 2 11 97.1774 $w=1.8e-07 $l=2.5e-07 $layer=POLY_cond $X=3.065 $Y=1.795
+ $X2=3.065 $Y2=1.545
.ends

.subckt PM_SKY130_FD_SC_LS__A211O_1%X 1 2 9 12 13 14 21 30
c21 30 0 1.55122e-19 $X=0.26 $Y=1.82
r22 19 21 1.31708 $w=3.48e-07 $l=4e-08 $layer=LI1_cond $X=0.26 $Y=1.995 $X2=0.26
+ $Y2=2.035
r23 13 14 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.26 $Y=2.405
+ $X2=0.26 $Y2=2.775
r24 12 19 0.75732 $w=3.48e-07 $l=2.3e-08 $layer=LI1_cond $X=0.26 $Y=1.972
+ $X2=0.26 $Y2=1.995
r25 12 30 8.06043 $w=3.48e-07 $l=1.52e-07 $layer=LI1_cond $X=0.26 $Y=1.972
+ $X2=0.26 $Y2=1.82
r26 12 13 11.4586 $w=3.48e-07 $l=3.48e-07 $layer=LI1_cond $X=0.26 $Y=2.057
+ $X2=0.26 $Y2=2.405
r27 12 21 0.724393 $w=3.48e-07 $l=2.2e-08 $layer=LI1_cond $X=0.26 $Y=2.057
+ $X2=0.26 $Y2=2.035
r28 9 11 13.9526 $w=7.17e-07 $l=8.2e-07 $layer=LI1_cond $X=0.17 $Y=0.737
+ $X2=0.99 $Y2=0.737
r29 7 9 9.47984 $w=1.7e-07 $l=3.93e-07 $layer=LI1_cond $X=0.17 $Y=1.13 $X2=0.17
+ $Y2=0.737
r30 7 30 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=0.17 $Y=1.13 $X2=0.17
+ $Y2=1.82
r31 2 12 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.84 $X2=0.27 $Y2=1.985
r32 2 14 400 $w=1.7e-07 $l=1.03562e-06 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.84 $X2=0.27 $Y2=2.815
r33 1 11 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.865
+ $Y=0.37 $X2=0.99 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__A211O_1%VPWR 1 2 9 15 18 19 20 22 35 36 39
r39 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r40 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r41 33 36 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.6 $Y2=3.33
r42 32 35 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=3.6 $Y2=3.33
r43 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r44 30 40 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r45 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r46 27 39 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.885 $Y=3.33
+ $X2=0.76 $Y2=3.33
r47 27 29 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=0.885 $Y=3.33
+ $X2=1.68 $Y2=3.33
r48 25 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r49 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r50 22 39 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.635 $Y=3.33
+ $X2=0.76 $Y2=3.33
r51 22 24 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=0.635 $Y=3.33
+ $X2=0.24 $Y2=3.33
r52 20 33 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.16 $Y2=3.33
r53 20 30 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r54 18 29 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.885 $Y=3.33
+ $X2=1.68 $Y2=3.33
r55 18 19 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=1.885 $Y=3.33 $X2=1.985
+ $Y2=3.33
r56 17 32 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=2.085 $Y=3.33
+ $X2=2.16 $Y2=3.33
r57 17 19 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=2.085 $Y=3.33 $X2=1.985
+ $Y2=3.33
r58 13 19 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=1.985 $Y=3.245
+ $X2=1.985 $Y2=3.33
r59 13 15 43.8091 $w=1.98e-07 $l=7.9e-07 $layer=LI1_cond $X=1.985 $Y=3.245
+ $X2=1.985 $Y2=2.455
r60 9 12 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=0.76 $Y=1.985
+ $X2=0.76 $Y2=2.815
r61 7 39 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.76 $Y=3.245
+ $X2=0.76 $Y2=3.33
r62 7 12 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.76 $Y=3.245 $X2=0.76
+ $Y2=2.815
r63 2 15 300 $w=1.7e-07 $l=5.71577e-07 $layer=licon1_PDIFF $count=2 $X=1.82
+ $Y=1.96 $X2=1.985 $Y2=2.455
r64 1 12 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=0.57
+ $Y=1.84 $X2=0.72 $Y2=2.815
r65 1 9 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=0.57
+ $Y=1.84 $X2=0.72 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_LS__A211O_1%A_279_392# 1 2 7 9 11 13 15
r36 13 20 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.45 $Y=2.12 $X2=2.45
+ $Y2=2.035
r37 13 15 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=2.45 $Y=2.12
+ $X2=2.45 $Y2=2.815
r38 12 18 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.685 $Y=2.035
+ $X2=1.52 $Y2=2.035
r39 11 20 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.285 $Y=2.035
+ $X2=2.45 $Y2=2.035
r40 11 12 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=2.285 $Y=2.035
+ $X2=1.685 $Y2=2.035
r41 7 18 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.52 $Y=2.12 $X2=1.52
+ $Y2=2.035
r42 7 9 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=1.52 $Y=2.12 $X2=1.52
+ $Y2=2.815
r43 2 20 400 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=1 $X=2.3
+ $Y=1.96 $X2=2.45 $Y2=2.115
r44 2 15 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=2.3
+ $Y=1.96 $X2=2.45 $Y2=2.815
r45 1 18 400 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=1 $X=1.395
+ $Y=1.96 $X2=1.52 $Y2=2.115
r46 1 9 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=1.395
+ $Y=1.96 $X2=1.52 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_LS__A211O_1%VGND 1 2 9 13 16 20 22 24 34 35 38 41
r46 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r47 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r48 35 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r49 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r50 32 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.215 $Y=0 $X2=3.13
+ $Y2=0
r51 32 34 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=3.215 $Y=0 $X2=3.6
+ $Y2=0
r52 31 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r53 30 31 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r54 27 31 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r55 26 30 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r56 26 27 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r57 24 38 10.5822 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=1.255 $Y=0 $X2=1.48
+ $Y2=0
r58 24 30 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=1.255 $Y=0 $X2=1.2
+ $Y2=0
r59 22 42 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.92 $Y=0 $X2=3.12
+ $Y2=0
r60 22 39 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r61 18 20 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.945 $Y=0.825
+ $X2=3.13 $Y2=0.825
r62 16 20 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.13 $Y=0.74
+ $X2=3.13 $Y2=0.825
r63 15 41 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.13 $Y=0.085
+ $X2=3.13 $Y2=0
r64 15 16 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=3.13 $Y=0.085
+ $X2=3.13 $Y2=0.74
r65 14 38 10.5822 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=1.705 $Y=0 $X2=1.48
+ $Y2=0
r66 13 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.045 $Y=0 $X2=3.13
+ $Y2=0
r67 13 14 87.4225 $w=1.68e-07 $l=1.34e-06 $layer=LI1_cond $X=3.045 $Y=0
+ $X2=1.705 $Y2=0
r68 9 11 9.03704 $w=4.48e-07 $l=3.4e-07 $layer=LI1_cond $X=1.48 $Y=0.495
+ $X2=1.48 $Y2=0.835
r69 7 38 1.79621 $w=4.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.48 $Y=0.085 $X2=1.48
+ $Y2=0
r70 7 9 10.8976 $w=4.48e-07 $l=4.1e-07 $layer=LI1_cond $X=1.48 $Y=0.085 $X2=1.48
+ $Y2=0.495
r71 2 18 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=2.735
+ $Y=0.68 $X2=2.945 $Y2=0.825
r72 1 11 182 $w=1.7e-07 $l=5.80625e-07 $layer=licon1_NDIFF $count=1 $X=1.28
+ $Y=0.37 $X2=1.54 $Y2=0.835
r73 1 9 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=1.28
+ $Y=0.37 $X2=1.42 $Y2=0.495
.ends

