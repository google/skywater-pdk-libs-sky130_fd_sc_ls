* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__a2bb2oi_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
X0 a_539_368# a_114_392# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X1 VPWR B2 a_539_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X2 a_539_368# a_114_392# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X3 VPWR B2 a_539_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X4 Y a_114_392# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X5 a_29_392# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 Y B2 a_914_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X7 VPWR B1 a_539_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X8 VGND B1 a_914_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X9 a_914_74# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X10 VGND a_114_392# Y VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X11 a_539_368# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X12 a_29_392# A2_N a_114_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 Y a_114_392# a_539_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X14 Y a_114_392# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X15 VGND a_114_392# Y VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X16 a_539_368# B2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X17 a_914_74# B2 Y VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X18 Y a_114_392# a_539_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X19 Y B2 a_914_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X20 a_914_74# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X21 a_914_74# B2 Y VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X22 VGND B1 a_914_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X23 VGND A2_N a_114_392# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X24 VPWR A1_N a_29_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X25 a_114_392# A1_N VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X26 a_114_392# A2_N a_29_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X27 a_539_368# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X28 a_539_368# B2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X29 VPWR B1 a_539_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
.ends
