* File: sky130_fd_sc_ls__dfrtp_1.pex.spice
* Created: Fri Aug 28 13:14:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__DFRTP_1%D 2 4 5 7 10 12 13 14 19 20 23
r35 23 25 40.9207 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=0.402 $Y=1.845
+ $X2=0.402 $Y2=2.01
r36 23 24 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.845 $X2=0.385 $Y2=1.845
r37 19 21 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=0.402 $Y=1.165
+ $X2=0.402 $Y2=1
r38 19 20 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.165 $X2=0.385 $Y2=1.165
r39 14 24 5.61447 $w=3.88e-07 $l=1.9e-07 $layer=LI1_cond $X=0.32 $Y=2.035
+ $X2=0.32 $Y2=1.845
r40 13 24 5.31897 $w=3.88e-07 $l=1.8e-07 $layer=LI1_cond $X=0.32 $Y=1.665
+ $X2=0.32 $Y2=1.845
r41 12 13 10.9334 $w=3.88e-07 $l=3.7e-07 $layer=LI1_cond $X=0.32 $Y=1.295
+ $X2=0.32 $Y2=1.665
r42 12 20 3.84148 $w=3.88e-07 $l=1.3e-07 $layer=LI1_cond $X=0.32 $Y=1.295
+ $X2=0.32 $Y2=1.165
r43 10 21 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=0.51 $Y=0.6 $X2=0.51
+ $Y2=1
r44 5 7 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.495 $Y=2.465
+ $X2=0.495 $Y2=2.75
r45 4 5 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.495 $Y=2.375 $X2=0.495
+ $Y2=2.465
r46 4 25 141.879 $w=1.8e-07 $l=3.65e-07 $layer=POLY_cond $X=0.495 $Y=2.375
+ $X2=0.495 $Y2=2.01
r47 2 23 2.68759 $w=3.65e-07 $l=1.7e-08 $layer=POLY_cond $X=0.402 $Y=1.828
+ $X2=0.402 $Y2=1.845
r48 1 19 2.68759 $w=3.65e-07 $l=1.7e-08 $layer=POLY_cond $X=0.402 $Y=1.182
+ $X2=0.402 $Y2=1.165
r49 1 2 102.129 $w=3.65e-07 $l=6.46e-07 $layer=POLY_cond $X=0.402 $Y=1.182
+ $X2=0.402 $Y2=1.828
.ends

.subckt PM_SKY130_FD_SC_LS__DFRTP_1%CLK 3 7 8 11 13
c48 13 0 2.08211e-19 $X=1.91 $Y=1.435
c49 11 0 3.00326e-19 $X=1.91 $Y=1.61
r50 11 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.91 $Y=1.61
+ $X2=1.91 $Y2=1.775
r51 11 13 47.9601 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=1.91 $Y=1.61
+ $X2=1.91 $Y2=1.435
r52 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.91
+ $Y=1.61 $X2=1.91 $Y2=1.61
r53 8 12 6.53105 $w=4.67e-07 $l=2.5e-07 $layer=LI1_cond $X=2.16 $Y=1.545
+ $X2=1.91 $Y2=1.545
r54 7 13 151.027 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=1.95 $Y=0.965
+ $X2=1.95 $Y2=1.435
r55 3 14 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=1.925 $Y=2.45
+ $X2=1.925 $Y2=1.775
.ends

.subckt PM_SKY130_FD_SC_LS__DFRTP_1%A_490_390# 1 2 7 8 11 12 14 16 18 20 21 22
+ 23 25 26 31 32 34 37 38 39 42 46 49 53 58 59 60 66 69
c202 59 0 2.2444e-20 $X=2.99 $Y=1.345
c203 53 0 9.01765e-20 $X=2.797 $Y=0.415
c204 39 0 1.54738e-19 $X=5.65 $Y=0.34
c205 32 0 8.54071e-20 $X=4.27 $Y=0.415
c206 31 0 6.90861e-20 $X=3.03 $Y=1.56
c207 22 0 1.83796e-19 $X=6.33 $Y=1.27
c208 16 0 9.78499e-20 $X=4.005 $Y=0.9
c209 7 0 8.23352e-20 $X=3.412 $Y=1.985
r210 68 69 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=7.13 $Y=1.18
+ $X2=7.335 $Y2=1.18
r211 66 75 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=6.855 $Y=1.18
+ $X2=6.855 $Y2=1.27
r212 65 68 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=6.855 $Y=1.18
+ $X2=7.13 $Y2=1.18
r213 65 66 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.855
+ $Y=1.18 $X2=6.855 $Y2=1.18
r214 60 62 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=4.355 $Y=0.415
+ $X2=4.355 $Y2=0.65
r215 58 59 6.91466 $w=2.48e-07 $l=1.5e-07 $layer=LI1_cond $X=2.99 $Y=1.195
+ $X2=2.99 $Y2=1.345
r216 57 58 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=2.95 $Y=0.805
+ $X2=2.95 $Y2=1.195
r217 56 57 7.35235 $w=4.73e-07 $l=8.5e-08 $layer=LI1_cond $X=2.797 $Y=0.72
+ $X2=2.797 $Y2=0.805
r218 53 56 7.68008 $w=4.73e-07 $l=3.05e-07 $layer=LI1_cond $X=2.797 $Y=0.415
+ $X2=2.797 $Y2=0.72
r219 52 71 29.2361 $w=3.05e-07 $l=1.85e-07 $layer=POLY_cond $X=3.335 $Y=1.82
+ $X2=3.335 $Y2=1.635
r220 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.335
+ $Y=1.82 $X2=3.335 $Y2=1.82
r221 49 51 10.3649 $w=3.59e-07 $l=3.05e-07 $layer=LI1_cond $X=3.03 $Y=1.882
+ $X2=3.335 $Y2=1.882
r222 48 49 14.273 $w=3.59e-07 $l=4.2e-07 $layer=LI1_cond $X=2.61 $Y=1.882
+ $X2=3.03 $Y2=1.882
r223 46 69 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.335 $Y=1.015
+ $X2=7.335 $Y2=1.18
r224 45 46 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=7.335 $Y=0.425
+ $X2=7.335 $Y2=1.015
r225 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.13
+ $Y=2.14 $X2=7.13 $Y2=2.14
r226 40 68 0.716491 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=7.13 $Y=1.345
+ $X2=7.13 $Y2=1.18
r227 40 42 27.7634 $w=3.28e-07 $l=7.95e-07 $layer=LI1_cond $X=7.13 $Y=1.345
+ $X2=7.13 $Y2=2.14
r228 38 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.25 $Y=0.34
+ $X2=7.335 $Y2=0.425
r229 38 39 104.385 $w=1.68e-07 $l=1.6e-06 $layer=LI1_cond $X=7.25 $Y=0.34
+ $X2=5.65 $Y2=0.34
r230 36 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.565 $Y=0.425
+ $X2=5.65 $Y2=0.34
r231 36 37 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=5.565 $Y=0.425
+ $X2=5.565 $Y2=0.565
r232 35 62 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.44 $Y=0.65
+ $X2=4.355 $Y2=0.65
r233 34 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.48 $Y=0.65
+ $X2=5.565 $Y2=0.565
r234 34 35 67.8503 $w=1.68e-07 $l=1.04e-06 $layer=LI1_cond $X=5.48 $Y=0.65
+ $X2=4.44 $Y2=0.65
r235 33 53 6.83586 $w=1.7e-07 $l=2.38e-07 $layer=LI1_cond $X=3.035 $Y=0.415
+ $X2=2.797 $Y2=0.415
r236 32 60 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.27 $Y=0.415
+ $X2=4.355 $Y2=0.415
r237 32 33 80.5722 $w=1.68e-07 $l=1.235e-06 $layer=LI1_cond $X=4.27 $Y=0.415
+ $X2=3.035 $Y2=0.415
r238 31 49 5.12588 $w=1.7e-07 $l=3.22e-07 $layer=LI1_cond $X=3.03 $Y=1.56
+ $X2=3.03 $Y2=1.882
r239 31 59 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=3.03 $Y=1.56
+ $X2=3.03 $Y2=1.345
r240 23 43 50.5804 $w=3.46e-07 $l=2.97909e-07 $layer=POLY_cond $X=7.265 $Y=2.39
+ $X2=7.16 $Y2=2.14
r241 23 25 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.265 $Y=2.39
+ $X2=7.265 $Y2=2.675
r242 21 75 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.69 $Y=1.27
+ $X2=6.855 $Y2=1.27
r243 21 22 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=6.69 $Y=1.27
+ $X2=6.33 $Y2=1.27
r244 18 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.255 $Y=1.195
+ $X2=6.33 $Y2=1.27
r245 18 20 146.207 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=6.255 $Y=1.195
+ $X2=6.255 $Y2=0.74
r246 14 27 55.5827 $w=2.18e-07 $l=2.62678e-07 $layer=POLY_cond $X=4.005 $Y=1.405
+ $X2=3.935 $Y2=1.635
r247 14 16 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=4.005 $Y=1.405
+ $X2=4.005 $Y2=0.9
r248 13 71 19.3576 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.5 $Y=1.635
+ $X2=3.335 $Y2=1.635
r249 12 27 11.5617 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=3.79 $Y=1.635
+ $X2=3.935 $Y2=1.635
r250 12 13 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=3.79 $Y=1.635
+ $X2=3.5 $Y2=1.635
r251 11 26 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.4 $Y=2.495 $X2=3.4
+ $Y2=2.21
r252 8 26 36.4084 $w=1.75e-07 $l=8.7e-08 $layer=POLY_cond $X=3.412 $Y=2.123
+ $X2=3.412 $Y2=2.21
r253 7 52 34.7586 $w=3.05e-07 $l=1.99825e-07 $layer=POLY_cond $X=3.412 $Y=1.985
+ $X2=3.335 $Y2=1.82
r254 7 8 55.1746 $w=1.75e-07 $l=1.38e-07 $layer=POLY_cond $X=3.412 $Y=1.985
+ $X2=3.412 $Y2=2.123
r255 2 48 600 $w=1.7e-07 $l=2.36854e-07 $layer=licon1_PDIFF $count=1 $X=2.45
+ $Y=1.95 $X2=2.61 $Y2=2.12
r256 1 56 182 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_NDIFF $count=1 $X=2.575
+ $Y=0.595 $X2=2.725 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_LS__DFRTP_1%A_830_359# 1 2 7 9 12 16 19 20 25 28 32
c83 20 0 2.21973e-20 $X=4.445 $Y=0.99
c84 16 0 9.22519e-20 $X=4.355 $Y=1.96
c85 12 0 2.89729e-19 $X=4.395 $Y=0.9
r86 31 32 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=6.065 $Y=1.13
+ $X2=6.065 $Y2=1.865
r87 30 31 7.58911 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=5.985 $Y=0.99
+ $X2=5.985 $Y2=1.13
r88 28 30 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=5.985 $Y=0.855
+ $X2=5.985 $Y2=0.99
r89 25 32 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=6.145 $Y=2.03
+ $X2=6.145 $Y2=1.865
r90 19 30 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.82 $Y=0.99
+ $X2=5.985 $Y2=0.99
r91 19 20 89.7059 $w=1.68e-07 $l=1.375e-06 $layer=LI1_cond $X=5.82 $Y=0.99
+ $X2=4.445 $Y2=0.99
r92 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.355
+ $Y=1.96 $X2=4.355 $Y2=1.96
r93 14 20 6.81835 $w=1.7e-07 $l=1.23386e-07 $layer=LI1_cond $X=4.357 $Y=1.075
+ $X2=4.445 $Y2=0.99
r94 14 16 56.0883 $w=1.73e-07 $l=8.85e-07 $layer=LI1_cond $X=4.357 $Y=1.075
+ $X2=4.357 $Y2=1.96
r95 10 17 38.6069 $w=3.31e-07 $l=1.92678e-07 $layer=POLY_cond $X=4.395 $Y=1.795
+ $X2=4.335 $Y2=1.96
r96 10 12 458.926 $w=1.5e-07 $l=8.95e-07 $layer=POLY_cond $X=4.395 $Y=1.795
+ $X2=4.395 $Y2=0.9
r97 7 17 50.9845 $w=3.31e-07 $l=2.93684e-07 $layer=POLY_cond $X=4.24 $Y=2.21
+ $X2=4.335 $Y2=1.96
r98 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.24 $Y=2.21 $X2=4.24
+ $Y2=2.495
r99 2 25 300 $w=1.7e-07 $l=3.78253e-07 $layer=licon1_PDIFF $count=2 $X=5.955
+ $Y=1.735 $X2=6.145 $Y2=2.03
r100 1 28 182 $w=1.7e-07 $l=6.8057e-07 $layer=licon1_NDIFF $count=1 $X=5.515
+ $Y=0.37 $X2=5.985 $Y2=0.855
.ends

.subckt PM_SKY130_FD_SC_LS__DFRTP_1%RESET_B 4 6 8 11 12 13 17 18 20 22 25 27 29
+ 30 33 35 36 37 38 41 43 46 49 50 53 57 63
c220 50 0 1.18035e-19 $X=1.155 $Y=1.295
c221 49 0 1.16646e-19 $X=1.155 $Y=1.295
c222 37 0 3.91908e-20 $X=7.775 $Y=2.035
c223 33 0 9.22519e-20 $X=4.875 $Y=1.26
c224 17 0 1.54738e-19 $X=4.785 $Y=0.9
c225 12 0 2.21973e-20 $X=4.71 $Y=0.18
r226 62 63 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.18
+ $Y=2.09 $X2=8.18 $Y2=2.09
r227 57 59 32.8941 $w=3.59e-07 $l=2.45e-07 $layer=POLY_cond $X=4.875 $Y=2.002
+ $X2=5.12 $Y2=2.002
r228 56 57 2.01393 $w=3.59e-07 $l=1.5e-08 $layer=POLY_cond $X=4.86 $Y=2.002
+ $X2=4.875 $Y2=2.002
r229 53 55 40.6549 $w=4.95e-07 $l=1.65e-07 $layer=POLY_cond $X=1.072 $Y=1.975
+ $X2=1.072 $Y2=2.14
r230 53 54 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.155
+ $Y=1.975 $X2=1.155 $Y2=1.975
r231 50 54 30.1408 $w=2.58e-07 $l=6.8e-07 $layer=LI1_cond $X=1.155 $Y=1.295
+ $X2=1.155 $Y2=1.975
r232 49 51 46.3954 $w=4.95e-07 $l=1.65e-07 $layer=POLY_cond $X=1.072 $Y=1.295
+ $X2=1.072 $Y2=1.13
r233 49 50 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.155
+ $Y=1.295 $X2=1.155 $Y2=1.295
r234 46 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=2.035
+ $X2=1.2 $Y2=2.035
r235 44 63 8.94433 $w=3.33e-07 $l=2.6e-07 $layer=LI1_cond $X=7.92 $Y=2.087
+ $X2=8.18 $Y2=2.087
r236 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=2.035
+ $X2=7.92 $Y2=2.035
r237 41 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.12
+ $Y=1.96 $X2=5.12 $Y2=1.96
r238 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=2.035
+ $X2=5.04 $Y2=2.035
r239 38 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.185 $Y=2.035
+ $X2=5.04 $Y2=2.035
r240 37 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.775 $Y=2.035
+ $X2=7.92 $Y2=2.035
r241 37 38 3.20544 $w=1.4e-07 $l=2.59e-06 $layer=MET1_cond $X=7.775 $Y=2.035
+ $X2=5.185 $Y2=2.035
r242 36 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.345 $Y=2.035
+ $X2=1.2 $Y2=2.035
r243 35 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.895 $Y=2.035
+ $X2=5.04 $Y2=2.035
r244 35 36 4.39356 $w=1.4e-07 $l=3.55e-06 $layer=MET1_cond $X=4.895 $Y=2.035
+ $X2=1.345 $Y2=2.035
r245 31 33 46.1489 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.785 $Y=1.26
+ $X2=4.875 $Y2=1.26
r246 27 62 61.0536 $w=2.9e-07 $l=3.36749e-07 $layer=POLY_cond $X=8.26 $Y=2.39
+ $X2=8.182 $Y2=2.09
r247 27 29 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=8.26 $Y=2.39
+ $X2=8.26 $Y2=2.675
r248 23 62 38.6157 $w=2.9e-07 $l=1.76125e-07 $layer=POLY_cond $X=8.205 $Y=1.925
+ $X2=8.182 $Y2=2.09
r249 23 25 671.723 $w=1.5e-07 $l=1.31e-06 $layer=POLY_cond $X=8.205 $Y=1.925
+ $X2=8.205 $Y2=0.615
r250 22 57 23.2387 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.875 $Y=1.795
+ $X2=4.875 $Y2=2.002
r251 21 33 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.875 $Y=1.335
+ $X2=4.875 $Y2=1.26
r252 21 22 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=4.875 $Y=1.335
+ $X2=4.875 $Y2=1.795
r253 18 56 23.2387 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=4.86 $Y=2.21
+ $X2=4.86 $Y2=2.002
r254 18 20 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.86 $Y=2.21
+ $X2=4.86 $Y2=2.495
r255 15 31 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.785 $Y=1.185
+ $X2=4.785 $Y2=1.26
r256 15 17 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.785 $Y=1.185
+ $X2=4.785 $Y2=0.9
r257 14 17 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=4.785 $Y=0.255
+ $X2=4.785 $Y2=0.9
r258 12 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.71 $Y=0.18
+ $X2=4.785 $Y2=0.255
r259 12 13 1915.18 $w=1.5e-07 $l=3.735e-06 $layer=POLY_cond $X=4.71 $Y=0.18
+ $X2=0.975 $Y2=0.18
r260 11 30 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.93 $Y=2.75
+ $X2=0.93 $Y2=2.465
r261 8 30 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.945 $Y=2.375
+ $X2=0.945 $Y2=2.465
r262 8 55 91.3468 $w=1.8e-07 $l=2.35e-07 $layer=POLY_cond $X=0.945 $Y=2.375
+ $X2=0.945 $Y2=2.14
r263 6 53 8.86311 $w=4.95e-07 $l=8.2e-08 $layer=POLY_cond $X=1.072 $Y=1.893
+ $X2=1.072 $Y2=1.975
r264 5 49 8.86311 $w=4.95e-07 $l=8.2e-08 $layer=POLY_cond $X=1.072 $Y=1.377
+ $X2=1.072 $Y2=1.295
r265 5 6 55.7728 $w=4.95e-07 $l=5.16e-07 $layer=POLY_cond $X=1.072 $Y=1.377
+ $X2=1.072 $Y2=1.893
r266 4 51 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.9 $Y=0.6 $X2=0.9
+ $Y2=1.13
r267 1 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.9 $Y=0.255
+ $X2=0.975 $Y2=0.18
r268 1 4 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=0.9 $Y=0.255 $X2=0.9
+ $Y2=0.6
.ends

.subckt PM_SKY130_FD_SC_LS__DFRTP_1%A_695_457# 1 2 3 12 14 16 22 23 26 27 29 30
+ 34 39 42 43 44
c126 43 0 1.48228e-19 $X=4.215 $Y=2.562
c127 42 0 8.46396e-20 $X=3.93 $Y=2.562
c128 39 0 9.01498e-20 $X=4.015 $Y=0.86
c129 22 0 1.23481e-19 $X=4.015 $Y=2.4
r130 37 39 6.82368 $w=3.78e-07 $l=2.25e-07 $layer=LI1_cond $X=3.79 $Y=0.86
+ $X2=4.015 $Y2=0.86
r131 32 44 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=4.785 $Y=2.445
+ $X2=4.7 $Y2=2.445
r132 32 34 13.8293 $w=2.48e-07 $l=3e-07 $layer=LI1_cond $X=4.785 $Y=2.445
+ $X2=5.085 $Y2=2.445
r133 30 47 72.1174 $w=2.64e-07 $l=3.95e-07 $layer=POLY_cond $X=5.485 $Y=1.452
+ $X2=5.88 $Y2=1.452
r134 30 45 8.21591 $w=2.64e-07 $l=4.5e-08 $layer=POLY_cond $X=5.485 $Y=1.452
+ $X2=5.44 $Y2=1.452
r135 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.485
+ $Y=1.41 $X2=5.485 $Y2=1.41
r136 27 29 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=4.785 $Y=1.41
+ $X2=5.485 $Y2=1.41
r137 26 44 2.11342 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.7 $Y=2.32 $X2=4.7
+ $Y2=2.445
r138 25 27 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.7 $Y=1.575
+ $X2=4.785 $Y2=1.41
r139 25 26 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=4.7 $Y=1.575
+ $X2=4.7 $Y2=2.32
r140 23 44 4.3182 $w=2.1e-07 $l=1.03078e-07 $layer=LI1_cond $X=4.615 $Y=2.485
+ $X2=4.7 $Y2=2.445
r141 23 43 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=4.615 $Y=2.485
+ $X2=4.215 $Y2=2.485
r142 22 43 9.70126 $w=3.23e-07 $l=2e-07 $layer=LI1_cond $X=4.015 $Y=2.562
+ $X2=4.215 $Y2=2.562
r143 22 42 4.01401 $w=3.23e-07 $l=8.5e-08 $layer=LI1_cond $X=4.015 $Y=2.562
+ $X2=3.93 $Y2=2.562
r144 21 39 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.015 $Y=1.05
+ $X2=4.015 $Y2=0.86
r145 21 22 88.0749 $w=1.68e-07 $l=1.35e-06 $layer=LI1_cond $X=4.015 $Y=1.05
+ $X2=4.015 $Y2=2.4
r146 19 42 15.2824 $w=2.28e-07 $l=3.05e-07 $layer=LI1_cond $X=3.625 $Y=2.61
+ $X2=3.93 $Y2=2.61
r147 14 47 15.9823 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=5.88 $Y=1.66
+ $X2=5.88 $Y2=1.452
r148 14 16 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.88 $Y=1.66
+ $X2=5.88 $Y2=2.235
r149 10 45 15.9823 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.44 $Y=1.245
+ $X2=5.44 $Y2=1.452
r150 10 12 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=5.44 $Y=1.245
+ $X2=5.44 $Y2=0.74
r151 3 34 600 $w=1.7e-07 $l=2.64575e-07 $layer=licon1_PDIFF $count=1 $X=4.935
+ $Y=2.285 $X2=5.085 $Y2=2.485
r152 2 19 600 $w=1.7e-07 $l=3.62319e-07 $layer=licon1_PDIFF $count=1 $X=3.475
+ $Y=2.285 $X2=3.625 $Y2=2.58
r153 1 37 182 $w=1.7e-07 $l=2.82489e-07 $layer=licon1_NDIFF $count=1 $X=3.58
+ $Y=0.69 $X2=3.79 $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_LS__DFRTP_1%A_306_96# 1 2 9 11 13 15 16 17 18 19 20 22
+ 25 27 32 33 34 37 39 40 44 47 48 52 53 57 59
c189 59 0 1.84578e-19 $X=2.61 $Y=1.49
c190 57 0 8.23352e-20 $X=2.61 $Y=1.61
c191 52 0 1.16646e-19 $X=1.647 $Y=1.055
c192 27 0 1.48228e-19 $X=6.295 $Y=3.15
c193 25 0 1.33086e-19 $X=3.85 $Y=2.495
c194 20 0 2.2444e-20 $X=3.505 $Y=1.2
c195 19 0 9.84449e-20 $X=3.095 $Y=1.275
c196 18 0 1.23481e-19 $X=3.43 $Y=1.275
c197 15 0 8.46396e-20 $X=2.885 $Y=3.075
c198 11 0 1.54493e-19 $X=2.5 $Y=1.41
c199 9 0 1.95608e-19 $X=2.375 $Y=2.45
r200 58 64 36.7175 $w=3.61e-07 $l=2.75e-07 $layer=POLY_cond $X=2.61 $Y=1.487
+ $X2=2.885 $Y2=1.487
r201 57 59 4.89537 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=2.61 $Y=1.61
+ $X2=2.61 $Y2=1.49
r202 57 58 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.61
+ $Y=1.61 $X2=2.61 $Y2=1.61
r203 53 55 7.83936 $w=2.49e-07 $l=1.6e-07 $layer=LI1_cond $X=1.54 $Y=2.092
+ $X2=1.7 $Y2=2.092
r204 50 59 16.1342 $w=2.48e-07 $l=3.5e-07 $layer=LI1_cond $X=2.57 $Y=1.14
+ $X2=2.57 $Y2=1.49
r205 49 52 3.15366 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=1.84 $Y=1.055
+ $X2=1.647 $Y2=1.055
r206 48 50 10.7448 $w=1.39e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.445 $Y=1.055
+ $X2=2.57 $Y2=1.14
r207 48 49 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=2.445 $Y=1.055
+ $X2=1.84 $Y2=1.055
r208 47 53 2.97181 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=1.54 $Y=1.945
+ $X2=1.54 $Y2=2.092
r209 46 52 3.37808 $w=2.77e-07 $l=1.43332e-07 $layer=LI1_cond $X=1.54 $Y=1.14
+ $X2=1.647 $Y2=1.055
r210 46 47 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=1.54 $Y=1.14
+ $X2=1.54 $Y2=1.945
r211 42 52 3.37808 $w=2.77e-07 $l=8.5e-08 $layer=LI1_cond $X=1.647 $Y=0.97
+ $X2=1.647 $Y2=1.055
r212 42 44 10.3271 $w=3.83e-07 $l=3.45e-07 $layer=LI1_cond $X=1.647 $Y=0.97
+ $X2=1.647 $Y2=0.625
r213 35 37 497.383 $w=1.5e-07 $l=9.7e-07 $layer=POLY_cond $X=7.305 $Y=1.585
+ $X2=7.305 $Y2=0.615
r214 33 35 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.23 $Y=1.66
+ $X2=7.305 $Y2=1.585
r215 33 34 387.138 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=7.23 $Y=1.66
+ $X2=6.475 $Y2=1.66
r216 30 40 76.0046 $w=1.8e-07 $l=1.9e-07 $layer=POLY_cond $X=6.385 $Y=2.96
+ $X2=6.385 $Y2=3.15
r217 30 32 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.385 $Y=2.96
+ $X2=6.385 $Y2=2.385
r218 29 34 26.9307 $w=1.5e-07 $l=1.89737e-07 $layer=POLY_cond $X=6.385 $Y=1.81
+ $X2=6.475 $Y2=1.66
r219 29 32 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.385 $Y=1.81
+ $X2=6.385 $Y2=2.385
r220 28 39 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.925 $Y=3.15
+ $X2=3.85 $Y2=3.15
r221 27 40 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=6.295 $Y=3.15
+ $X2=6.385 $Y2=3.15
r222 27 28 1215.26 $w=1.5e-07 $l=2.37e-06 $layer=POLY_cond $X=6.295 $Y=3.15
+ $X2=3.925 $Y2=3.15
r223 23 39 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.85 $Y=3.075
+ $X2=3.85 $Y2=3.15
r224 23 25 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.85 $Y=3.075
+ $X2=3.85 $Y2=2.495
r225 20 22 96.4 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=3.505 $Y=1.2 $X2=3.505
+ $Y2=0.9
r226 19 64 44.9323 $w=3.61e-07 $l=2.99105e-07 $layer=POLY_cond $X=3.095 $Y=1.275
+ $X2=2.885 $Y2=1.487
r227 18 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.43 $Y=1.275
+ $X2=3.505 $Y2=1.2
r228 18 19 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=3.43 $Y=1.275
+ $X2=3.095 $Y2=1.275
r229 16 39 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.775 $Y=3.15
+ $X2=3.85 $Y2=3.15
r230 16 17 417.904 $w=1.5e-07 $l=8.15e-07 $layer=POLY_cond $X=3.775 $Y=3.15
+ $X2=2.96 $Y2=3.15
r231 15 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.885 $Y=3.075
+ $X2=2.96 $Y2=3.15
r232 14 64 23.3725 $w=1.5e-07 $l=2.88e-07 $layer=POLY_cond $X=2.885 $Y=1.775
+ $X2=2.885 $Y2=1.487
r233 14 15 666.596 $w=1.5e-07 $l=1.3e-06 $layer=POLY_cond $X=2.885 $Y=1.775
+ $X2=2.885 $Y2=3.075
r234 11 58 14.687 $w=3.61e-07 $l=1.1e-07 $layer=POLY_cond $X=2.5 $Y=1.487
+ $X2=2.61 $Y2=1.487
r235 11 61 16.6898 $w=3.61e-07 $l=1.25e-07 $layer=POLY_cond $X=2.5 $Y=1.487
+ $X2=2.375 $Y2=1.487
r236 11 13 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.5 $Y=1.41
+ $X2=2.5 $Y2=0.965
r237 7 61 23.3725 $w=1.5e-07 $l=2.88e-07 $layer=POLY_cond $X=2.375 $Y=1.775
+ $X2=2.375 $Y2=1.487
r238 7 9 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=2.375 $Y=1.775
+ $X2=2.375 $Y2=2.45
r239 2 55 600 $w=1.7e-07 $l=2.13542e-07 $layer=licon1_PDIFF $count=1 $X=1.54
+ $Y=1.95 $X2=1.7 $Y2=2.075
r240 1 44 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=1.53
+ $Y=0.48 $X2=1.675 $Y2=0.625
.ends

.subckt PM_SKY130_FD_SC_LS__DFRTP_1%A_1518_203# 1 2 9 10 11 13 16 18 19 25 27 28
+ 30 31 35 38 39 42
r119 38 39 10.5766 $w=3.63e-07 $l=2.3e-07 $layer=LI1_cond $X=8.502 $Y=2.675
+ $X2=8.502 $Y2=2.445
r120 35 46 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.755 $Y=1.18
+ $X2=7.755 $Y2=1.345
r121 35 45 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.755 $Y=1.18
+ $X2=7.755 $Y2=1.015
r122 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.755
+ $Y=1.18 $X2=7.755 $Y2=1.18
r123 31 34 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=7.755 $Y=1.1 $X2=7.755
+ $Y2=1.18
r124 29 42 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.105 $Y=1.185
+ $X2=9.105 $Y2=1.1
r125 29 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.105 $Y=1.185
+ $X2=9.105 $Y2=1.855
r126 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.02 $Y=1.94
+ $X2=9.105 $Y2=1.855
r127 27 28 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=9.02 $Y=1.94
+ $X2=8.685 $Y2=1.94
r128 23 42 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=8.78 $Y=1.1
+ $X2=9.105 $Y2=1.1
r129 23 25 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=8.78 $Y=1.015 $X2=8.78
+ $Y2=0.615
r130 21 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.6 $Y=2.025
+ $X2=8.685 $Y2=1.94
r131 21 39 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=8.6 $Y=2.025
+ $X2=8.6 $Y2=2.445
r132 20 31 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.92 $Y=1.1
+ $X2=7.755 $Y2=1.1
r133 19 23 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=8.615 $Y=1.1
+ $X2=8.78 $Y2=1.1
r134 19 20 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=8.615 $Y=1.1
+ $X2=7.92 $Y2=1.1
r135 18 46 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=7.67 $Y=1.745
+ $X2=7.67 $Y2=1.345
r136 16 45 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=7.695 $Y=0.615
+ $X2=7.695 $Y2=1.015
r137 11 13 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.685 $Y=2.39
+ $X2=7.685 $Y2=2.675
r138 10 11 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=7.685 $Y=2.3
+ $X2=7.685 $Y2=2.39
r139 9 18 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=7.685 $Y=1.835
+ $X2=7.685 $Y2=1.745
r140 9 10 180.75 $w=1.8e-07 $l=4.65e-07 $layer=POLY_cond $X=7.685 $Y=1.835
+ $X2=7.685 $Y2=2.3
r141 2 38 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=8.335
+ $Y=2.465 $X2=8.485 $Y2=2.675
r142 1 25 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=8.64
+ $Y=0.405 $X2=8.78 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_LS__DFRTP_1%A_1266_74# 1 2 9 12 13 15 16 17 19 21 22 24
+ 25 26 27 29 30 31 32 34 37 39 40 44 45 46 51 54
c161 51 0 1.44605e-19 $X=6.565 $Y=1.6
c162 46 0 1.4888e-19 $X=7.635 $Y=1.6
c163 45 0 3.23044e-20 $X=8.52 $Y=1.6
c164 44 0 1.01622e-19 $X=7.55 $Y=2.475
r165 55 61 3.86218 $w=3.12e-07 $l=2.5e-08 $layer=POLY_cond $X=8.685 $Y=1.52
+ $X2=8.71 $Y2=1.52
r166 55 59 18.5385 $w=3.12e-07 $l=1.2e-07 $layer=POLY_cond $X=8.685 $Y=1.52
+ $X2=8.565 $Y2=1.52
r167 54 57 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=8.685 $Y=1.52
+ $X2=8.685 $Y2=1.6
r168 54 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.685
+ $Y=1.52 $X2=8.685 $Y2=1.52
r169 49 51 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=6.405 $Y=1.6
+ $X2=6.565 $Y2=1.6
r170 45 57 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.52 $Y=1.6
+ $X2=8.685 $Y2=1.6
r171 45 46 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=8.52 $Y=1.6
+ $X2=7.635 $Y2=1.6
r172 43 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.55 $Y=1.685
+ $X2=7.635 $Y2=1.6
r173 43 44 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=7.55 $Y=1.685
+ $X2=7.55 $Y2=2.475
r174 40 42 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=6.65 $Y=2.64
+ $X2=7.04 $Y2=2.64
r175 39 44 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.465 $Y=2.64
+ $X2=7.55 $Y2=2.475
r176 39 42 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=7.465 $Y=2.64
+ $X2=7.04 $Y2=2.64
r177 35 48 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.49 $Y=0.72
+ $X2=6.405 $Y2=0.72
r178 35 37 19.5915 $w=2.48e-07 $l=4.25e-07 $layer=LI1_cond $X=6.49 $Y=0.72
+ $X2=6.915 $Y2=0.72
r179 34 40 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.565 $Y=2.475
+ $X2=6.65 $Y2=2.64
r180 33 51 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.565 $Y=1.685
+ $X2=6.565 $Y2=1.6
r181 33 34 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=6.565 $Y=1.685
+ $X2=6.565 $Y2=2.475
r182 32 49 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.405 $Y=1.515
+ $X2=6.405 $Y2=1.6
r183 31 48 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.405 $Y=0.845
+ $X2=6.405 $Y2=0.72
r184 31 32 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.405 $Y=0.845
+ $X2=6.405 $Y2=1.515
r185 27 29 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=9.555 $Y=0.995
+ $X2=9.555 $Y2=0.645
r186 25 27 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.48 $Y=1.07
+ $X2=9.555 $Y2=0.995
r187 25 26 89.734 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=9.48 $Y=1.07
+ $X2=9.305 $Y2=1.07
r188 22 24 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=9.245 $Y=1.97
+ $X2=9.245 $Y2=2.465
r189 21 22 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=9.245 $Y=1.88
+ $X2=9.245 $Y2=1.97
r190 20 30 34.7346 $w=1.65e-07 $l=1.65e-07 $layer=POLY_cond $X=9.245 $Y=1.685
+ $X2=9.245 $Y2=1.52
r191 20 21 75.7984 $w=1.8e-07 $l=1.95e-07 $layer=POLY_cond $X=9.245 $Y=1.685
+ $X2=9.245 $Y2=1.88
r192 19 30 34.7346 $w=1.65e-07 $l=1.72337e-07 $layer=POLY_cond $X=9.23 $Y=1.355
+ $X2=9.245 $Y2=1.52
r193 18 26 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.23 $Y=1.145
+ $X2=9.305 $Y2=1.07
r194 18 19 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=9.23 $Y=1.145
+ $X2=9.23 $Y2=1.355
r195 17 61 13.3422 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=8.8 $Y=1.52 $X2=8.71
+ $Y2=1.52
r196 16 30 3.90195 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=9.155 $Y=1.52
+ $X2=9.245 $Y2=1.52
r197 16 17 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=9.155 $Y=1.52
+ $X2=8.8 $Y2=1.52
r198 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=8.71 $Y=2.39
+ $X2=8.71 $Y2=2.675
r199 12 13 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=8.71 $Y=2.3 $X2=8.71
+ $Y2=2.39
r200 11 61 15.628 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=8.71 $Y=1.685
+ $X2=8.71 $Y2=1.52
r201 11 12 239.056 $w=1.8e-07 $l=6.15e-07 $layer=POLY_cond $X=8.71 $Y=1.685
+ $X2=8.71 $Y2=2.3
r202 7 59 19.893 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.565 $Y=1.355
+ $X2=8.565 $Y2=1.52
r203 7 9 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=8.565 $Y=1.355
+ $X2=8.565 $Y2=0.615
r204 2 42 300 $w=1.7e-07 $l=1.00395e-06 $layer=licon1_PDIFF $count=2 $X=6.46
+ $Y=1.885 $X2=7.04 $Y2=2.64
r205 1 48 182 $w=1.7e-07 $l=3.79671e-07 $layer=licon1_NDIFF $count=1 $X=6.33
+ $Y=0.37 $X2=6.485 $Y2=0.68
r206 1 37 182 $w=1.7e-07 $l=7.23585e-07 $layer=licon1_NDIFF $count=1 $X=6.33
+ $Y=0.37 $X2=6.915 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_LS__DFRTP_1%A_1864_409# 1 2 7 9 12 14 15 18 22 27
r54 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.77
+ $Y=1.55 $X2=9.77 $Y2=1.55
r55 24 27 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=9.47 $Y=1.55 $X2=9.77
+ $Y2=1.55
r56 20 27 0.716491 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=9.77 $Y=1.385
+ $X2=9.77 $Y2=1.55
r57 20 22 25.8427 $w=3.28e-07 $l=7.4e-07 $layer=LI1_cond $X=9.77 $Y=1.385
+ $X2=9.77 $Y2=0.645
r58 16 24 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.47 $Y=1.715
+ $X2=9.47 $Y2=1.55
r59 16 18 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=9.47 $Y=1.715
+ $X2=9.47 $Y2=2.19
r60 14 28 117.157 $w=3.3e-07 $l=6.7e-07 $layer=POLY_cond $X=10.44 $Y=1.55
+ $X2=9.77 $Y2=1.55
r61 14 15 5.03009 $w=3.3e-07 $l=1.01735e-07 $layer=POLY_cond $X=10.44 $Y=1.55
+ $X2=10.53 $Y2=1.575
r62 10 15 37.0704 $w=1.5e-07 $l=1.97358e-07 $layer=POLY_cond $X=10.545 $Y=1.385
+ $X2=10.53 $Y2=1.575
r63 10 12 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=10.545 $Y=1.385
+ $X2=10.545 $Y2=0.74
r64 7 15 37.0704 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=10.53 $Y=1.765
+ $X2=10.53 $Y2=1.575
r65 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=10.53 $Y=1.765
+ $X2=10.53 $Y2=2.4
r66 2 18 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=9.32
+ $Y=2.045 $X2=9.47 $Y2=2.19
r67 1 22 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=9.63
+ $Y=0.37 $X2=9.77 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_LS__DFRTP_1%VPWR 1 2 3 4 5 6 7 8 25 27 31 35 39 41 45 51
+ 53 57 59 61 65 67 72 77 85 93 105 108 111 114 117 120 124
r149 123 124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r150 120 121 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r151 118 121 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.88 $Y2=3.33
r152 117 118 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r153 111 112 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r154 108 109 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r155 105 106 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r156 102 103 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r157 100 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=10.8 $Y2=3.33
r158 99 100 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r159 97 100 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=10.32 $Y2=3.33
r160 97 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=8.88 $Y2=3.33
r161 96 99 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=9.36 $Y=3.33
+ $X2=10.32 $Y2=3.33
r162 96 97 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r163 94 120 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.185 $Y=3.33
+ $X2=9.02 $Y2=3.33
r164 94 96 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=9.185 $Y=3.33
+ $X2=9.36 $Y2=3.33
r165 93 123 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=10.595 $Y=3.33
+ $X2=10.817 $Y2=3.33
r166 93 99 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=10.595 $Y=3.33
+ $X2=10.32 $Y2=3.33
r167 92 118 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r168 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r169 89 92 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=7.44 $Y2=3.33
r170 88 91 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=6 $Y=3.33 $X2=7.44
+ $Y2=3.33
r171 88 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r172 86 114 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.81 $Y=3.33
+ $X2=5.645 $Y2=3.33
r173 86 88 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=5.81 $Y=3.33 $X2=6
+ $Y2=3.33
r174 85 117 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.805 $Y=3.33
+ $X2=7.97 $Y2=3.33
r175 85 91 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=7.805 $Y=3.33
+ $X2=7.44 $Y2=3.33
r176 84 112 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r177 83 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r178 81 84 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=4.08 $Y2=3.33
r179 81 109 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r180 80 83 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.64 $Y=3.33
+ $X2=4.08 $Y2=3.33
r181 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r182 78 108 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.315 $Y=3.33
+ $X2=2.15 $Y2=3.33
r183 78 80 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.315 $Y=3.33
+ $X2=2.64 $Y2=3.33
r184 77 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.385 $Y=3.33
+ $X2=4.55 $Y2=3.33
r185 77 83 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.385 $Y=3.33
+ $X2=4.08 $Y2=3.33
r186 76 109 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r187 76 106 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r188 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r189 73 105 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.31 $Y=3.33
+ $X2=1.145 $Y2=3.33
r190 73 75 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.31 $Y=3.33
+ $X2=1.68 $Y2=3.33
r191 72 108 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.985 $Y=3.33
+ $X2=2.15 $Y2=3.33
r192 72 75 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.985 $Y=3.33
+ $X2=1.68 $Y2=3.33
r193 71 106 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r194 71 103 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r195 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r196 68 102 4.02368 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=0.355 $Y=3.33
+ $X2=0.177 $Y2=3.33
r197 68 70 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.355 $Y=3.33
+ $X2=0.72 $Y2=3.33
r198 67 105 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.98 $Y=3.33
+ $X2=1.145 $Y2=3.33
r199 67 70 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.98 $Y=3.33
+ $X2=0.72 $Y2=3.33
r200 65 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33 $X2=6
+ $Y2=3.33
r201 65 112 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=4.56 $Y2=3.33
r202 65 114 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r203 61 64 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=10.76 $Y=1.985
+ $X2=10.76 $Y2=2.815
r204 59 123 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=10.76 $Y=3.245
+ $X2=10.817 $Y2=3.33
r205 59 64 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=10.76 $Y=3.245
+ $X2=10.76 $Y2=2.815
r206 55 120 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.02 $Y=3.245
+ $X2=9.02 $Y2=3.33
r207 55 57 30.9064 $w=3.28e-07 $l=8.85e-07 $layer=LI1_cond $X=9.02 $Y=3.245
+ $X2=9.02 $Y2=2.36
r208 54 117 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.135 $Y=3.33
+ $X2=7.97 $Y2=3.33
r209 53 120 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.855 $Y=3.33
+ $X2=9.02 $Y2=3.33
r210 53 54 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=8.855 $Y=3.33
+ $X2=8.135 $Y2=3.33
r211 49 117 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.97 $Y=3.245
+ $X2=7.97 $Y2=3.33
r212 49 51 19.9058 $w=3.28e-07 $l=5.7e-07 $layer=LI1_cond $X=7.97 $Y=3.245
+ $X2=7.97 $Y2=2.675
r213 45 48 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=5.645 $Y=1.91
+ $X2=5.645 $Y2=2.59
r214 43 114 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.645 $Y=3.245
+ $X2=5.645 $Y2=3.33
r215 43 48 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=5.645 $Y=3.245
+ $X2=5.645 $Y2=2.59
r216 42 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.715 $Y=3.33
+ $X2=4.55 $Y2=3.33
r217 41 114 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.48 $Y=3.33
+ $X2=5.645 $Y2=3.33
r218 41 42 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=5.48 $Y=3.33
+ $X2=4.715 $Y2=3.33
r219 37 111 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.55 $Y=3.245
+ $X2=4.55 $Y2=3.33
r220 37 39 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=4.55 $Y=3.245
+ $X2=4.55 $Y2=2.825
r221 33 108 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.15 $Y=3.245
+ $X2=2.15 $Y2=3.33
r222 33 35 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=2.15 $Y=3.245
+ $X2=2.15 $Y2=2.825
r223 29 105 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.145 $Y=3.245
+ $X2=1.145 $Y2=3.33
r224 29 31 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=1.145 $Y=3.245
+ $X2=1.145 $Y2=2.815
r225 25 102 3.11948 $w=2.5e-07 $l=1.08305e-07 $layer=LI1_cond $X=0.23 $Y=3.245
+ $X2=0.177 $Y2=3.33
r226 25 27 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=0.23 $Y=3.245
+ $X2=0.23 $Y2=2.75
r227 8 64 400 $w=1.7e-07 $l=1.04964e-06 $layer=licon1_PDIFF $count=1 $X=10.605
+ $Y=1.84 $X2=10.76 $Y2=2.815
r228 8 61 400 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=1 $X=10.605
+ $Y=1.84 $X2=10.76 $Y2=1.985
r229 7 57 300 $w=1.7e-07 $l=2.82666e-07 $layer=licon1_PDIFF $count=2 $X=8.785
+ $Y=2.465 $X2=9.02 $Y2=2.36
r230 6 51 600 $w=1.7e-07 $l=2.96985e-07 $layer=licon1_PDIFF $count=1 $X=7.76
+ $Y=2.465 $X2=7.97 $Y2=2.675
r231 5 48 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=5.5
+ $Y=1.735 $X2=5.645 $Y2=2.59
r232 5 45 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=5.5
+ $Y=1.735 $X2=5.645 $Y2=1.91
r233 4 39 600 $w=1.7e-07 $l=6.46916e-07 $layer=licon1_PDIFF $count=1 $X=4.315
+ $Y=2.285 $X2=4.55 $Y2=2.825
r234 3 35 600 $w=1.7e-07 $l=9.47035e-07 $layer=licon1_PDIFF $count=1 $X=2
+ $Y=1.95 $X2=2.15 $Y2=2.825
r235 2 31 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=1.005
+ $Y=2.54 $X2=1.145 $Y2=2.815
r236 1 27 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.54 $X2=0.27 $Y2=2.75
.ends

.subckt PM_SKY130_FD_SC_LS__DFRTP_1%A_30_78# 1 2 3 4 13 17 20 21 23 25 28 29 32
+ 34 38 40 44 49
c133 44 0 9.78499e-20 $X=3.29 $Y=0.88
c134 40 0 2.31531e-19 $X=3.172 $Y=2.472
c135 25 0 1.15748e-19 $X=3.01 $Y=2.472
c136 23 0 1.95608e-19 $X=1.835 $Y=2.51
r137 47 49 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.37 $Y=1.305
+ $X2=3.675 $Y2=1.305
r138 44 46 8.79328 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=3.33 $Y=0.88
+ $X2=3.33 $Y2=1.045
r139 40 42 0.998577 $w=2.81e-07 $l=2.3e-08 $layer=LI1_cond $X=3.172 $Y=2.472
+ $X2=3.172 $Y2=2.495
r140 39 40 10.0726 $w=2.81e-07 $l=2.32e-07 $layer=LI1_cond $X=3.172 $Y=2.24
+ $X2=3.172 $Y2=2.472
r141 34 36 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=0.295 $Y=0.6
+ $X2=0.295 $Y2=0.745
r142 31 49 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.675 $Y=1.39
+ $X2=3.675 $Y2=1.305
r143 31 32 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=3.675 $Y=1.39
+ $X2=3.675 $Y2=2.155
r144 30 39 3.67734 $w=1.7e-07 $l=1.63e-07 $layer=LI1_cond $X=3.335 $Y=2.24
+ $X2=3.172 $Y2=2.24
r145 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.59 $Y=2.24
+ $X2=3.675 $Y2=2.155
r146 29 30 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=3.59 $Y=2.24
+ $X2=3.335 $Y2=2.24
r147 28 47 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.37 $Y=1.22
+ $X2=3.37 $Y2=1.305
r148 28 46 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.37 $Y=1.22
+ $X2=3.37 $Y2=1.045
r149 25 40 2.89855 $w=1.95e-07 $l=1.62e-07 $layer=LI1_cond $X=3.01 $Y=2.472
+ $X2=3.172 $Y2=2.472
r150 25 26 61.711 $w=1.93e-07 $l=1.085e-06 $layer=LI1_cond $X=3.01 $Y=2.472
+ $X2=1.925 $Y2=2.472
r151 23 26 5.46269 $w=2.01e-07 $l=1.07331e-07 $layer=LI1_cond $X=1.835 $Y=2.51
+ $X2=1.925 $Y2=2.472
r152 23 24 16.9136 $w=1.98e-07 $l=3.05e-07 $layer=LI1_cond $X=1.835 $Y=2.51
+ $X2=1.53 $Y2=2.51
r153 22 38 0.764409 $w=2.5e-07 $l=3.44891e-07 $layer=LI1_cond $X=0.86 $Y=2.435
+ $X2=0.555 $Y2=2.52
r154 21 24 6.00394 $w=2.54e-07 $l=1.58114e-07 $layer=LI1_cond $X=1.405 $Y=2.435
+ $X2=1.53 $Y2=2.51
r155 21 22 25.1233 $w=2.48e-07 $l=5.45e-07 $layer=LI1_cond $X=1.405 $Y=2.435
+ $X2=0.86 $Y2=2.435
r156 20 38 5.90115 $w=2.12e-07 $l=3.02283e-07 $layer=LI1_cond $X=0.77 $Y=2.31
+ $X2=0.555 $Y2=2.52
r157 19 20 96.5562 $w=1.68e-07 $l=1.48e-06 $layer=LI1_cond $X=0.77 $Y=0.83
+ $X2=0.77 $Y2=2.31
r158 15 38 5.90115 $w=2.12e-07 $l=1.77113e-07 $layer=LI1_cond $X=0.682 $Y=2.64
+ $X2=0.555 $Y2=2.52
r159 15 17 4.97132 $w=2.53e-07 $l=1.1e-07 $layer=LI1_cond $X=0.682 $Y=2.64
+ $X2=0.682 $Y2=2.75
r160 14 36 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.46 $Y=0.745
+ $X2=0.295 $Y2=0.745
r161 13 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.685 $Y=0.745
+ $X2=0.77 $Y2=0.83
r162 13 14 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.685 $Y=0.745
+ $X2=0.46 $Y2=0.745
r163 4 42 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=3.035
+ $Y=2.285 $X2=3.175 $Y2=2.495
r164 3 17 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=0.57
+ $Y=2.54 $X2=0.715 $Y2=2.75
r165 2 44 182 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_NDIFF $count=1 $X=3.145
+ $Y=0.69 $X2=3.29 $Y2=0.88
r166 1 34 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.15
+ $Y=0.39 $X2=0.295 $Y2=0.6
.ends

.subckt PM_SKY130_FD_SC_LS__DFRTP_1%Q 1 2 9 13 14 15 16 29
r29 20 32 3.16106 $w=6.98e-07 $l=1.85e-07 $layer=LI1_cond $X=10.075 $Y=2.235
+ $X2=10.075 $Y2=2.05
r30 16 26 0.683473 $w=6.98e-07 $l=4e-08 $layer=LI1_cond $X=10.075 $Y=2.775
+ $X2=10.075 $Y2=2.815
r31 15 16 6.32213 $w=6.98e-07 $l=3.7e-07 $layer=LI1_cond $X=10.075 $Y=2.405
+ $X2=10.075 $Y2=2.775
r32 15 20 2.90476 $w=6.98e-07 $l=1.7e-07 $layer=LI1_cond $X=10.075 $Y=2.405
+ $X2=10.075 $Y2=2.235
r33 14 32 0.256303 $w=6.98e-07 $l=1.5e-08 $layer=LI1_cond $X=10.075 $Y=2.035
+ $X2=10.075 $Y2=2.05
r34 14 29 7.51816 $w=6.98e-07 $l=1.5e-07 $layer=LI1_cond $X=10.075 $Y=2.035
+ $X2=10.075 $Y2=1.885
r35 13 29 33.4652 $w=2.58e-07 $l=7.55e-07 $layer=LI1_cond $X=10.295 $Y=1.13
+ $X2=10.295 $Y2=1.885
r36 7 13 6.31279 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=10.33 $Y=0.965
+ $X2=10.33 $Y2=1.13
r37 7 9 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=10.33 $Y=0.965
+ $X2=10.33 $Y2=0.515
r38 2 32 400 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=10.115
+ $Y=1.84 $X2=10.26 $Y2=2.05
r39 2 26 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=10.115
+ $Y=1.84 $X2=10.26 $Y2=2.815
r40 1 9 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=10.185
+ $Y=0.37 $X2=10.33 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__DFRTP_1%VGND 1 2 3 4 5 6 21 25 29 33 35 37 40 41 42
+ 48 52 60 68 73 79 89 92 96
c104 96 0 1.99579e-19 $X=10.8 $Y=0
c105 29 0 3.23044e-20 $X=7.91 $Y=0.615
r106 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=0 $X2=10.8
+ $Y2=0
r107 92 93 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r108 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r109 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r110 77 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=10.8 $Y2=0
r111 77 93 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=9.36 $Y2=0
r112 76 77 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r113 74 92 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.425 $Y=0 $X2=9.3
+ $Y2=0
r114 74 76 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=9.425 $Y=0
+ $X2=10.32 $Y2=0
r115 73 95 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=10.675 $Y=0
+ $X2=10.857 $Y2=0
r116 73 76 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=10.675 $Y=0
+ $X2=10.32 $Y2=0
r117 72 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=9.36
+ $Y2=0
r118 72 90 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=7.92
+ $Y2=0
r119 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r120 69 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.075 $Y=0 $X2=7.91
+ $Y2=0
r121 69 71 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=8.075 $Y=0
+ $X2=8.88 $Y2=0
r122 68 92 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.175 $Y=0 $X2=9.3
+ $Y2=0
r123 68 71 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=9.175 $Y=0 $X2=8.88
+ $Y2=0
r124 67 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=7.92
+ $Y2=0
r125 66 67 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r126 63 66 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=5.52 $Y=0 $X2=7.44
+ $Y2=0
r127 61 63 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=5.31 $Y=0 $X2=5.52
+ $Y2=0
r128 60 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.745 $Y=0 $X2=7.91
+ $Y2=0
r129 60 66 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7.745 $Y=0
+ $X2=7.44 $Y2=0
r130 59 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r131 58 59 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r132 56 59 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=4.56 $Y2=0
r133 56 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r134 55 58 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=2.64 $Y=0 $X2=4.56
+ $Y2=0
r135 55 56 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r136 53 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.39 $Y=0 $X2=2.225
+ $Y2=0
r137 53 55 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.39 $Y=0 $X2=2.64
+ $Y2=0
r138 52 86 9.04449 $w=3.93e-07 $l=3.1e-07 $layer=LI1_cond $X=5.112 $Y=0
+ $X2=5.112 $Y2=0.31
r139 52 61 5.70203 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=5.112 $Y=0 $X2=5.31
+ $Y2=0
r140 52 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r141 52 58 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=4.915 $Y=0
+ $X2=4.56 $Y2=0
r142 51 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r143 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r144 48 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.06 $Y=0 $X2=2.225
+ $Y2=0
r145 48 50 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=2.06 $Y=0 $X2=1.68
+ $Y2=0
r146 46 51 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r147 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r148 42 67 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=5.52 $Y=0
+ $X2=7.44 $Y2=0
r149 42 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r150 42 63 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r151 40 45 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1.03 $Y=0 $X2=0.72
+ $Y2=0
r152 40 41 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.03 $Y=0 $X2=1.155
+ $Y2=0
r153 39 50 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=1.28 $Y=0 $X2=1.68
+ $Y2=0
r154 39 41 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.28 $Y=0 $X2=1.155
+ $Y2=0
r155 35 95 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=10.8 $Y=0.085
+ $X2=10.857 $Y2=0
r156 35 37 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=10.8 $Y=0.085
+ $X2=10.8 $Y2=0.515
r157 31 92 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.3 $Y=0.085
+ $X2=9.3 $Y2=0
r158 31 33 23.5098 $w=2.48e-07 $l=5.1e-07 $layer=LI1_cond $X=9.3 $Y=0.085
+ $X2=9.3 $Y2=0.595
r159 27 89 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.91 $Y=0.085
+ $X2=7.91 $Y2=0
r160 27 29 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=7.91 $Y=0.085
+ $X2=7.91 $Y2=0.615
r161 23 79 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.225 $Y=0.085
+ $X2=2.225 $Y2=0
r162 23 25 22.0012 $w=3.28e-07 $l=6.3e-07 $layer=LI1_cond $X=2.225 $Y=0.085
+ $X2=2.225 $Y2=0.715
r163 19 41 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.155 $Y=0.085
+ $X2=1.155 $Y2=0
r164 19 21 23.7403 $w=2.48e-07 $l=5.15e-07 $layer=LI1_cond $X=1.155 $Y=0.085
+ $X2=1.155 $Y2=0.6
r165 6 37 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.62
+ $Y=0.37 $X2=10.76 $Y2=0.515
r166 5 33 182 $w=1.7e-07 $l=2.88531e-07 $layer=licon1_NDIFF $count=1 $X=9.195
+ $Y=0.37 $X2=9.34 $Y2=0.595
r167 4 29 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=7.77
+ $Y=0.405 $X2=7.91 $Y2=0.615
r168 3 86 182 $w=1.7e-07 $l=4.89285e-07 $layer=licon1_NDIFF $count=1 $X=4.86
+ $Y=0.69 $X2=5.11 $Y2=0.31
r169 2 25 182 $w=1.7e-07 $l=2.52982e-07 $layer=licon1_NDIFF $count=1 $X=2.025
+ $Y=0.595 $X2=2.225 $Y2=0.715
r170 1 21 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.975
+ $Y=0.39 $X2=1.115 $Y2=0.6
.ends

