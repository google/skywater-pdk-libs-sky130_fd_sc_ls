* File: sky130_fd_sc_ls__diode_2.pxi.spice
* Created: Wed Sep  2 11:02:40 2020
* 
x_PM_SKY130_FD_SC_LS__DIODE_2%DIODE N_DIODE_D0_noxref_neg DIODE DIODE DIODE
+ DIODE DIODE DIODE DIODE N_DIODE_c_7_n PM_SKY130_FD_SC_LS__DIODE_2%DIODE
x_PM_SKY130_FD_SC_LS__DIODE_2%VGND VGND VGND PM_SKY130_FD_SC_LS__DIODE_2%VGND
x_PM_SKY130_FD_SC_LS__DIODE_2%VPWR VPWR VPWR PM_SKY130_FD_SC_LS__DIODE_2%VPWR
cc_1 VNB N_DIODE_c_7_n 0.135211f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=0.445
cc_2 VNB VGND 0.122102f $X=-0.19 $Y=-0.245 $X2=0.135 $Y2=0.32
cc_3 VNB VPWR 0.0442671f $X=-0.19 $Y=-0.245 $X2=0.135 $Y2=0.32
cc_4 VPB N_DIODE_c_7_n 0.160044f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=0.445
cc_5 VPB VPWR 0.0500209f $X=-0.19 $Y=1.66 $X2=0.135 $Y2=0.32
cc_6 VPB VPWR 0.027814f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_7 N_DIODE_c_7_n VGND 0.0814983f $X=0.28 $Y=0.445 $X2=-0.19 $Y2=-0.245
cc_8 N_DIODE_c_7_n VPWR 0.0297164f $X=0.28 $Y=0.445 $X2=-0.19 $Y2=-0.245
cc_9 N_DIODE_c_7_n VPWR 0.051782f $X=0.28 $Y=0.445 $X2=0 $Y2=0
