# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ls__or2b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_ls__or2b_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.232500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.035000 1.350000 2.365000 1.780000 ;
    END
  END A
  PIN B_N
    ANTENNAGATEAREA  0.208500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.180000 0.455000 1.550000 ;
    END
  END B_N
  PIN X
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.755000 1.820000 3.275000 2.980000 ;
        RECT 2.875000 0.350000 3.275000 1.130000 ;
        RECT 3.105000 1.130000 3.275000 1.820000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.115000  0.680000 0.830000 1.010000 ;
      RECT 0.115000  1.760000 0.830000 1.930000 ;
      RECT 0.115000  1.930000 0.445000 2.980000 ;
      RECT 0.615000  2.100000 0.945000 3.245000 ;
      RECT 0.660000  1.010000 0.830000 1.300000 ;
      RECT 0.660000  1.300000 1.525000 1.630000 ;
      RECT 0.660000  1.630000 0.830000 1.760000 ;
      RECT 1.000000  0.085000 1.525000 1.130000 ;
      RECT 1.300000  1.820000 1.865000 1.990000 ;
      RECT 1.300000  1.990000 1.630000 2.860000 ;
      RECT 1.695000  0.540000 2.045000 1.010000 ;
      RECT 1.695000  1.010000 2.705000 1.180000 ;
      RECT 1.695000  1.180000 1.865000 1.820000 ;
      RECT 2.255000  1.950000 2.585000 3.245000 ;
      RECT 2.265000  0.085000 2.680000 0.840000 ;
      RECT 2.535000  1.180000 2.705000 1.300000 ;
      RECT 2.535000  1.300000 2.935000 1.630000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_ls__or2b_1
END LIBRARY
