* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__dlxtn_2 D GATE_N VGND VNB VPB VPWR Q
M1000 a_658_79# a_27_120# VGND VNB nshort w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=1.54015e+12p ps=1.207e+07u
M1001 a_232_82# GATE_N VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1002 VGND a_842_405# a_875_139# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1003 VPWR a_842_405# Q VPB phighvt w=1.12e+06u l=150000u
+  ad=2.00335e+12p pd=1.509e+07u as=3.864e+11p ps=2.93e+06u
M1004 VPWR a_842_405# a_791_503# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1005 VGND a_232_82# a_369_392# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1006 VPWR a_232_82# a_369_392# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=2.478e+11p ps=2.27e+06u
M1007 a_791_503# a_232_82# a_669_392# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=4.05175e+11p ps=2.92e+06u
M1008 VGND a_842_405# Q VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.516e+11p ps=2.16e+06u
M1009 a_842_405# a_669_392# VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1010 a_875_139# a_369_392# a_669_392# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=2.803e+11p ps=2.53e+06u
M1011 a_669_392# a_369_392# a_585_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1012 a_585_392# a_27_120# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR D a_27_120# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=2.478e+11p ps=2.27e+06u
M1014 VGND D a_27_120# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1015 a_842_405# a_669_392# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=0p ps=0u
M1016 Q a_842_405# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_232_82# GATE_N VPWR VPB phighvt w=840000u l=150000u
+  ad=2.478e+11p pd=2.27e+06u as=0p ps=0u
M1018 Q a_842_405# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_669_392# a_232_82# a_658_79# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
