* File: sky130_fd_sc_ls__sedfxtp_2.pxi.spice
* Created: Fri Aug 28 14:07:33 2020
* 
x_PM_SKY130_FD_SC_LS__SEDFXTP_2%D N_D_c_339_n N_D_c_340_n N_D_M1009_g
+ N_D_M1005_g D D N_D_c_336_n N_D_c_337_n N_D_c_338_n N_D_c_343_n
+ PM_SKY130_FD_SC_LS__SEDFXTP_2%D
x_PM_SKY130_FD_SC_LS__SEDFXTP_2%A_180_290# N_A_180_290#_M1013_s
+ N_A_180_290#_M1038_s N_A_180_290#_c_385_n N_A_180_290#_M1034_g
+ N_A_180_290#_M1015_g N_A_180_290#_c_386_n N_A_180_290#_c_378_n
+ N_A_180_290#_c_379_n N_A_180_290#_c_380_n N_A_180_290#_c_381_n
+ N_A_180_290#_c_388_n N_A_180_290#_c_389_n N_A_180_290#_c_382_n
+ N_A_180_290#_c_390_n N_A_180_290#_c_391_n N_A_180_290#_c_383_n
+ N_A_180_290#_c_384_n PM_SKY130_FD_SC_LS__SEDFXTP_2%A_180_290#
x_PM_SKY130_FD_SC_LS__SEDFXTP_2%DE N_DE_M1029_g N_DE_c_485_n N_DE_c_486_n
+ N_DE_c_487_n N_DE_c_493_n N_DE_c_494_n N_DE_c_488_n N_DE_M1013_g N_DE_c_495_n
+ N_DE_M1038_g N_DE_c_496_n N_DE_c_497_n N_DE_M1014_g N_DE_c_489_n N_DE_c_498_n
+ DE N_DE_c_490_n N_DE_c_499_n N_DE_c_491_n PM_SKY130_FD_SC_LS__SEDFXTP_2%DE
x_PM_SKY130_FD_SC_LS__SEDFXTP_2%A_548_87# N_A_548_87#_M1023_d
+ N_A_548_87#_M1035_d N_A_548_87#_M1025_g N_A_548_87#_c_590_n
+ N_A_548_87#_c_591_n N_A_548_87#_M1032_g N_A_548_87#_c_578_n
+ N_A_548_87#_M1021_g N_A_548_87#_c_579_n N_A_548_87#_c_580_n
+ N_A_548_87#_c_592_n N_A_548_87#_M1037_g N_A_548_87#_c_581_n
+ N_A_548_87#_c_594_n N_A_548_87#_c_582_n N_A_548_87#_c_583_n
+ N_A_548_87#_c_595_n N_A_548_87#_c_596_n N_A_548_87#_c_584_n
+ N_A_548_87#_c_597_n N_A_548_87#_c_598_n N_A_548_87#_c_585_n
+ N_A_548_87#_c_586_n N_A_548_87#_c_601_n N_A_548_87#_c_587_n
+ N_A_548_87#_c_588_n N_A_548_87#_c_589_n
+ PM_SKY130_FD_SC_LS__SEDFXTP_2%A_548_87#
x_PM_SKY130_FD_SC_LS__SEDFXTP_2%A_663_87# N_A_663_87#_M1031_s
+ N_A_663_87#_M1003_s N_A_663_87#_c_829_n N_A_663_87#_M1026_g
+ N_A_663_87#_c_830_n N_A_663_87#_c_831_n N_A_663_87#_c_839_n
+ N_A_663_87#_M1010_g N_A_663_87#_c_832_n N_A_663_87#_c_840_n
+ N_A_663_87#_c_833_n N_A_663_87#_c_834_n N_A_663_87#_c_849_n
+ N_A_663_87#_c_835_n N_A_663_87#_c_842_n N_A_663_87#_c_843_n
+ N_A_663_87#_c_836_n N_A_663_87#_c_837_n N_A_663_87#_c_838_n
+ N_A_663_87#_c_845_n N_A_663_87#_c_846_n
+ PM_SKY130_FD_SC_LS__SEDFXTP_2%A_663_87#
x_PM_SKY130_FD_SC_LS__SEDFXTP_2%SCD N_SCD_M1041_g N_SCD_c_942_n N_SCD_c_943_n
+ N_SCD_M1018_g SCD N_SCD_c_941_n PM_SKY130_FD_SC_LS__SEDFXTP_2%SCD
x_PM_SKY130_FD_SC_LS__SEDFXTP_2%SCE N_SCE_c_989_n N_SCE_M1002_g N_SCE_c_990_n
+ N_SCE_c_991_n N_SCE_c_982_n N_SCE_c_993_n N_SCE_M1003_g N_SCE_M1031_g
+ N_SCE_c_984_n N_SCE_c_985_n N_SCE_M1004_g SCE N_SCE_c_987_n N_SCE_c_988_n
+ PM_SKY130_FD_SC_LS__SEDFXTP_2%SCE
x_PM_SKY130_FD_SC_LS__SEDFXTP_2%CLK N_CLK_c_1067_n N_CLK_M1042_g N_CLK_c_1068_n
+ N_CLK_M1011_g CLK PM_SKY130_FD_SC_LS__SEDFXTP_2%CLK
x_PM_SKY130_FD_SC_LS__SEDFXTP_2%A_1538_74# N_A_1538_74#_M1024_d
+ N_A_1538_74#_M1033_d N_A_1538_74#_c_1126_n N_A_1538_74#_M1000_g
+ N_A_1538_74#_c_1101_n N_A_1538_74#_M1016_g N_A_1538_74#_M1040_g
+ N_A_1538_74#_c_1103_n N_A_1538_74#_c_1128_n N_A_1538_74#_M1006_g
+ N_A_1538_74#_c_1104_n N_A_1538_74#_c_1105_n N_A_1538_74#_c_1106_n
+ N_A_1538_74#_c_1129_n N_A_1538_74#_c_1107_n N_A_1538_74#_c_1108_n
+ N_A_1538_74#_c_1109_n N_A_1538_74#_c_1208_p N_A_1538_74#_c_1110_n
+ N_A_1538_74#_c_1111_n N_A_1538_74#_c_1112_n N_A_1538_74#_c_1113_n
+ N_A_1538_74#_c_1114_n N_A_1538_74#_c_1115_n N_A_1538_74#_c_1116_n
+ N_A_1538_74#_c_1117_n N_A_1538_74#_c_1118_n N_A_1538_74#_c_1119_n
+ N_A_1538_74#_c_1133_n N_A_1538_74#_c_1134_n N_A_1538_74#_c_1120_n
+ N_A_1538_74#_c_1121_n N_A_1538_74#_c_1122_n N_A_1538_74#_c_1123_n
+ N_A_1538_74#_c_1124_n N_A_1538_74#_c_1125_n
+ PM_SKY130_FD_SC_LS__SEDFXTP_2%A_1538_74#
x_PM_SKY130_FD_SC_LS__SEDFXTP_2%A_1340_74# N_A_1340_74#_M1042_d
+ N_A_1340_74#_M1011_d N_A_1340_74#_M1024_g N_A_1340_74#_c_1339_n
+ N_A_1340_74#_c_1354_n N_A_1340_74#_M1033_g N_A_1340_74#_c_1340_n
+ N_A_1340_74#_M1012_g N_A_1340_74#_c_1342_n N_A_1340_74#_c_1357_n
+ N_A_1340_74#_c_1358_n N_A_1340_74#_M1007_g N_A_1340_74#_c_1343_n
+ N_A_1340_74#_M1043_g N_A_1340_74#_M1020_g N_A_1340_74#_c_1345_n
+ N_A_1340_74#_c_1346_n N_A_1340_74#_c_1347_n N_A_1340_74#_c_1348_n
+ N_A_1340_74#_c_1362_n N_A_1340_74#_c_1363_n N_A_1340_74#_c_1349_n
+ N_A_1340_74#_c_1350_n N_A_1340_74#_c_1351_n N_A_1340_74#_c_1366_n
+ N_A_1340_74#_c_1352_n PM_SKY130_FD_SC_LS__SEDFXTP_2%A_1340_74#
x_PM_SKY130_FD_SC_LS__SEDFXTP_2%A_1979_71# N_A_1979_71#_M1017_d
+ N_A_1979_71#_M1030_d N_A_1979_71#_M1019_g N_A_1979_71#_c_1527_n
+ N_A_1979_71#_c_1540_n N_A_1979_71#_M1001_g N_A_1979_71#_c_1528_n
+ N_A_1979_71#_c_1529_n N_A_1979_71#_c_1542_n N_A_1979_71#_M1028_g
+ N_A_1979_71#_c_1530_n N_A_1979_71#_M1039_g N_A_1979_71#_c_1531_n
+ N_A_1979_71#_c_1532_n N_A_1979_71#_c_1533_n N_A_1979_71#_c_1534_n
+ N_A_1979_71#_c_1535_n N_A_1979_71#_c_1536_n N_A_1979_71#_c_1544_n
+ N_A_1979_71#_c_1537_n N_A_1979_71#_c_1538_n
+ PM_SKY130_FD_SC_LS__SEDFXTP_2%A_1979_71#
x_PM_SKY130_FD_SC_LS__SEDFXTP_2%A_1736_97# N_A_1736_97#_M1012_d
+ N_A_1736_97#_M1000_d N_A_1736_97#_c_1632_n N_A_1736_97#_M1030_g
+ N_A_1736_97#_M1017_g N_A_1736_97#_c_1634_n N_A_1736_97#_c_1636_n
+ N_A_1736_97#_c_1637_n N_A_1736_97#_c_1638_n N_A_1736_97#_c_1639_n
+ N_A_1736_97#_c_1640_n PM_SKY130_FD_SC_LS__SEDFXTP_2%A_1736_97#
x_PM_SKY130_FD_SC_LS__SEDFXTP_2%A_2474_74# N_A_2474_74#_M1040_d
+ N_A_2474_74#_M1043_d N_A_2474_74#_M1023_g N_A_2474_74#_c_1729_n
+ N_A_2474_74#_M1035_g N_A_2474_74#_c_1718_n N_A_2474_74#_M1008_g
+ N_A_2474_74#_c_1730_n N_A_2474_74#_M1022_g N_A_2474_74#_M1036_g
+ N_A_2474_74#_c_1731_n N_A_2474_74#_M1027_g N_A_2474_74#_c_1721_n
+ N_A_2474_74#_c_1732_n N_A_2474_74#_c_1722_n N_A_2474_74#_c_1723_n
+ N_A_2474_74#_c_1724_n N_A_2474_74#_c_1725_n N_A_2474_74#_c_1734_n
+ N_A_2474_74#_c_1735_n N_A_2474_74#_c_1736_n N_A_2474_74#_c_1726_n
+ N_A_2474_74#_c_1738_n N_A_2474_74#_c_1739_n N_A_2474_74#_c_1727_n
+ N_A_2474_74#_c_1728_n PM_SKY130_FD_SC_LS__SEDFXTP_2%A_2474_74#
x_PM_SKY130_FD_SC_LS__SEDFXTP_2%A_40_464# N_A_40_464#_M1005_s
+ N_A_40_464#_M1025_d N_A_40_464#_M1009_s N_A_40_464#_M1032_d
+ N_A_40_464#_c_1885_n N_A_40_464#_c_1892_n N_A_40_464#_c_1893_n
+ N_A_40_464#_c_1894_n N_A_40_464#_c_1895_n N_A_40_464#_c_1896_n
+ N_A_40_464#_c_1928_n N_A_40_464#_c_1897_n N_A_40_464#_c_1898_n
+ N_A_40_464#_c_1886_n N_A_40_464#_c_1899_n N_A_40_464#_c_1887_n
+ N_A_40_464#_c_1888_n N_A_40_464#_c_1901_n N_A_40_464#_c_1889_n
+ N_A_40_464#_c_1890_n N_A_40_464#_c_1902_n
+ PM_SKY130_FD_SC_LS__SEDFXTP_2%A_40_464#
x_PM_SKY130_FD_SC_LS__SEDFXTP_2%VPWR N_VPWR_M1034_d N_VPWR_M1038_d
+ N_VPWR_M1003_d N_VPWR_M1011_s N_VPWR_M1033_s N_VPWR_M1001_d N_VPWR_M1028_s
+ N_VPWR_M1037_d N_VPWR_M1022_d N_VPWR_M1027_d N_VPWR_c_2014_n N_VPWR_c_2015_n
+ N_VPWR_c_2016_n N_VPWR_c_2017_n N_VPWR_c_2018_n N_VPWR_c_2019_n
+ N_VPWR_c_2020_n N_VPWR_c_2021_n N_VPWR_c_2022_n N_VPWR_c_2023_n
+ N_VPWR_c_2024_n N_VPWR_c_2025_n N_VPWR_c_2026_n N_VPWR_c_2027_n
+ N_VPWR_c_2028_n VPWR N_VPWR_c_2029_n N_VPWR_c_2030_n N_VPWR_c_2031_n
+ N_VPWR_c_2032_n N_VPWR_c_2033_n N_VPWR_c_2034_n N_VPWR_c_2035_n
+ N_VPWR_c_2036_n N_VPWR_c_2037_n N_VPWR_c_2038_n N_VPWR_c_2039_n
+ N_VPWR_c_2040_n N_VPWR_c_2041_n N_VPWR_c_2042_n N_VPWR_c_2043_n
+ N_VPWR_c_2013_n PM_SKY130_FD_SC_LS__SEDFXTP_2%VPWR
x_PM_SKY130_FD_SC_LS__SEDFXTP_2%A_693_113# N_A_693_113#_M1026_d
+ N_A_693_113#_M1004_d N_A_693_113#_M1012_s N_A_693_113#_M1002_d
+ N_A_693_113#_M1010_d N_A_693_113#_M1000_s N_A_693_113#_c_2204_n
+ N_A_693_113#_c_2260_n N_A_693_113#_c_2205_n N_A_693_113#_c_2216_n
+ N_A_693_113#_c_2228_n N_A_693_113#_c_2206_n N_A_693_113#_c_2207_n
+ N_A_693_113#_c_2208_n N_A_693_113#_c_2209_n N_A_693_113#_c_2197_n
+ N_A_693_113#_c_2198_n N_A_693_113#_c_2284_n N_A_693_113#_c_2199_n
+ N_A_693_113#_c_2210_n N_A_693_113#_c_2211_n N_A_693_113#_c_2200_n
+ N_A_693_113#_c_2201_n N_A_693_113#_c_2202_n N_A_693_113#_c_2203_n
+ N_A_693_113#_c_2214_n N_A_693_113#_c_2357_n N_A_693_113#_c_2294_n
+ PM_SKY130_FD_SC_LS__SEDFXTP_2%A_693_113#
x_PM_SKY130_FD_SC_LS__SEDFXTP_2%Q N_Q_M1008_d N_Q_M1022_s N_Q_c_2373_n
+ N_Q_c_2374_n N_Q_c_2377_n N_Q_c_2375_n Q Q PM_SKY130_FD_SC_LS__SEDFXTP_2%Q
x_PM_SKY130_FD_SC_LS__SEDFXTP_2%VGND N_VGND_M1029_d N_VGND_M1013_d
+ N_VGND_M1031_d N_VGND_M1042_s N_VGND_M1024_s N_VGND_M1019_d N_VGND_M1039_s
+ N_VGND_M1021_d N_VGND_M1008_s N_VGND_M1036_s N_VGND_c_2406_n N_VGND_c_2407_n
+ N_VGND_c_2408_n N_VGND_c_2409_n N_VGND_c_2410_n N_VGND_c_2411_n
+ N_VGND_c_2412_n N_VGND_c_2413_n N_VGND_c_2414_n N_VGND_c_2415_n
+ N_VGND_c_2416_n N_VGND_c_2417_n VGND N_VGND_c_2418_n N_VGND_c_2419_n
+ N_VGND_c_2420_n N_VGND_c_2421_n N_VGND_c_2422_n N_VGND_c_2423_n
+ N_VGND_c_2424_n N_VGND_c_2425_n N_VGND_c_2426_n N_VGND_c_2427_n
+ N_VGND_c_2428_n N_VGND_c_2429_n N_VGND_c_2430_n N_VGND_c_2431_n
+ N_VGND_c_2432_n N_VGND_c_2433_n N_VGND_c_2434_n N_VGND_c_2435_n
+ PM_SKY130_FD_SC_LS__SEDFXTP_2%VGND
cc_1 VNB N_D_M1005_g 0.0260114f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=0.58
cc_2 VNB N_D_c_336_n 0.0165369f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.145
cc_3 VNB N_D_c_337_n 0.010567f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.145
cc_4 VNB N_D_c_338_n 0.0397312f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.825
cc_5 VNB N_A_180_290#_M1015_g 0.040638f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_6 VNB N_A_180_290#_c_378_n 0.0035874f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.145
cc_7 VNB N_A_180_290#_c_379_n 0.0223828f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.145
cc_8 VNB N_A_180_290#_c_380_n 0.00932288f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.825
cc_9 VNB N_A_180_290#_c_381_n 0.00210868f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.825
cc_10 VNB N_A_180_290#_c_382_n 0.00790857f $X=-0.19 $Y=-0.245 $X2=0.615
+ $Y2=1.295
cc_11 VNB N_A_180_290#_c_383_n 0.00433271f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_180_290#_c_384_n 0.0190488f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_DE_M1029_g 0.0296573f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=2.245
cc_14 VNB N_DE_c_485_n 0.0291452f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=2.64
cc_15 VNB N_DE_c_486_n 0.00716237f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=0.98
cc_16 VNB N_DE_c_487_n 3.94837e-19 $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.145
cc_17 VNB N_DE_c_488_n 0.0158293f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_18 VNB N_DE_c_489_n 0.0326795f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_DE_c_490_n 0.023491f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_DE_c_491_n 0.0164279f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_548_87#_M1025_g 0.0426392f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_548_87#_c_578_n 0.0186115f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.825
cc_23 VNB N_A_548_87#_c_579_n 0.0394088f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.145
cc_24 VNB N_A_548_87#_c_580_n 0.00644191f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.825
cc_25 VNB N_A_548_87#_c_581_n 0.0348273f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_548_87#_c_582_n 0.0121241f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.825
cc_27 VNB N_A_548_87#_c_583_n 0.00158358f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_548_87#_c_584_n 0.00864587f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_548_87#_c_585_n 0.0651529f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_548_87#_c_586_n 0.00204689f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_548_87#_c_587_n 2.18259e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_548_87#_c_588_n 0.00744674f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_548_87#_c_589_n 0.025642f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_663_87#_c_829_n 0.0171115f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=0.58
cc_35 VNB N_A_663_87#_c_830_n 0.033708f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.145
cc_36 VNB N_A_663_87#_c_831_n 0.00938744f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=0.98
cc_37 VNB N_A_663_87#_c_832_n 0.00866805f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.145
cc_38 VNB N_A_663_87#_c_833_n 0.00203688f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.825
cc_39 VNB N_A_663_87#_c_834_n 0.0784723f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.825
cc_40 VNB N_A_663_87#_c_835_n 0.0342598f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.665
cc_41 VNB N_A_663_87#_c_836_n 0.00315597f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_663_87#_c_837_n 0.0267328f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_663_87#_c_838_n 0.00709414f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_SCD_M1041_g 0.0304223f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=2.245
cc_45 VNB SCD 0.0124313f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.145
cc_46 VNB N_SCD_c_941_n 0.0208697f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_47 VNB N_SCE_c_982_n 0.00807656f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=0.58
cc_48 VNB N_SCE_M1031_g 0.0319157f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_SCE_c_984_n 0.0616487f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.825
cc_50 VNB N_SCE_c_985_n 0.012806f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.145
cc_51 VNB N_SCE_M1004_g 0.0386896f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.825
cc_52 VNB N_SCE_c_987_n 0.031307f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_SCE_c_988_n 0.00275365f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.295
cc_54 VNB N_CLK_c_1067_n 0.0210376f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.99
cc_55 VNB N_CLK_c_1068_n 0.0560825f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=2.64
cc_56 VNB CLK 0.00751673f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=0.58
cc_57 VNB N_A_1538_74#_c_1101_n 0.018902f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.145
cc_58 VNB N_A_1538_74#_M1040_g 0.0352219f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_1538_74#_c_1103_n 0.00362656f $X=-0.19 $Y=-0.245 $X2=0.525
+ $Y2=1.145
cc_60 VNB N_A_1538_74#_c_1104_n 0.0099863f $X=-0.19 $Y=-0.245 $X2=0.615
+ $Y2=1.145
cc_61 VNB N_A_1538_74#_c_1105_n 0.0189124f $X=-0.19 $Y=-0.245 $X2=0.615
+ $Y2=1.295
cc_62 VNB N_A_1538_74#_c_1106_n 0.00279267f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_1538_74#_c_1107_n 0.00587229f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_1538_74#_c_1108_n 0.0176487f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_1538_74#_c_1109_n 0.00896906f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_1538_74#_c_1110_n 0.0113155f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_1538_74#_c_1111_n 0.0020311f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_1538_74#_c_1112_n 0.00981814f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_1538_74#_c_1113_n 0.00520534f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_1538_74#_c_1114_n 0.00320136f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_1538_74#_c_1115_n 0.0030334f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_1538_74#_c_1116_n 7.65667e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_1538_74#_c_1117_n 0.0175898f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_1538_74#_c_1118_n 0.0117094f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_1538_74#_c_1119_n 0.00123754f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_1538_74#_c_1120_n 0.00236228f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_1538_74#_c_1121_n 6.44577e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_1538_74#_c_1122_n 0.0452835f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_1538_74#_c_1123_n 0.0015664f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_1538_74#_c_1124_n 0.00361396f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_1538_74#_c_1125_n 0.0309263f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_1340_74#_M1024_g 0.0447807f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=0.98
cc_83 VNB N_A_1340_74#_c_1339_n 0.0127601f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_84 VNB N_A_1340_74#_c_1340_n 0.00990482f $X=-0.19 $Y=-0.245 $X2=0.525
+ $Y2=1.145
cc_85 VNB N_A_1340_74#_M1012_g 0.0513349f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.825
cc_86 VNB N_A_1340_74#_c_1342_n 0.0277393f $X=-0.19 $Y=-0.245 $X2=0.615
+ $Y2=1.145
cc_87 VNB N_A_1340_74#_c_1343_n 0.0157309f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_1340_74#_M1020_g 0.0508942f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_1340_74#_c_1345_n 0.00611157f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_1340_74#_c_1346_n 0.00382845f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_1340_74#_c_1347_n 0.00788613f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_1340_74#_c_1348_n 0.0117619f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_1340_74#_c_1349_n 0.0019697f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_1340_74#_c_1350_n 0.00991103f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_1340_74#_c_1351_n 0.0171048f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_1340_74#_c_1352_n 0.00213748f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_1979_71#_M1019_g 0.029864f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_A_1979_71#_c_1527_n 0.0108759f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_99 VNB N_A_1979_71#_c_1528_n 0.0319705f $X=-0.19 $Y=-0.245 $X2=0.525
+ $Y2=1.145
cc_100 VNB N_A_1979_71#_c_1529_n 0.00906352f $X=-0.19 $Y=-0.245 $X2=0.525
+ $Y2=1.145
cc_101 VNB N_A_1979_71#_c_1530_n 0.0203438f $X=-0.19 $Y=-0.245 $X2=0.525
+ $Y2=1.99
cc_102 VNB N_A_1979_71#_c_1531_n 0.00977398f $X=-0.19 $Y=-0.245 $X2=0.615
+ $Y2=1.295
cc_103 VNB N_A_1979_71#_c_1532_n 0.0100358f $X=-0.19 $Y=-0.245 $X2=0.615
+ $Y2=1.825
cc_104 VNB N_A_1979_71#_c_1533_n 0.00246868f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_A_1979_71#_c_1534_n 0.00200186f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_A_1979_71#_c_1535_n 0.0591256f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_A_1979_71#_c_1536_n 0.00167554f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_A_1979_71#_c_1537_n 0.00289677f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_A_1979_71#_c_1538_n 0.0392121f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_A_1736_97#_c_1632_n 0.0181373f $X=-0.19 $Y=-0.245 $X2=0.615
+ $Y2=0.58
cc_111 VNB N_A_1736_97#_M1017_g 0.0430138f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_112 VNB N_A_1736_97#_c_1634_n 0.0190396f $X=-0.19 $Y=-0.245 $X2=0.525
+ $Y2=1.825
cc_113 VNB N_A_2474_74#_M1023_g 0.0525498f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_A_2474_74#_c_1718_n 0.0682933f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_A_2474_74#_M1008_g 0.0273344f $X=-0.19 $Y=-0.245 $X2=0.525
+ $Y2=1.145
cc_116 VNB N_A_2474_74#_M1036_g 0.030592f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_A_2474_74#_c_1721_n 0.0161401f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_A_2474_74#_c_1722_n 0.0505973f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_A_2474_74#_c_1723_n 0.00286116f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_A_2474_74#_c_1724_n 0.0162708f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_A_2474_74#_c_1725_n 0.00250462f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_A_2474_74#_c_1726_n 0.00931714f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB N_A_2474_74#_c_1727_n 0.0044313f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_A_2474_74#_c_1728_n 0.00407735f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_A_40_464#_c_1885_n 0.040464f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_A_40_464#_c_1886_n 0.00249806f $X=-0.19 $Y=-0.245 $X2=0.615
+ $Y2=1.825
cc_127 VNB N_A_40_464#_c_1887_n 0.00686598f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_A_40_464#_c_1888_n 0.0307549f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_A_40_464#_c_1889_n 0.00290645f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_A_40_464#_c_1890_n 0.00466982f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_VPWR_c_2013_n 0.681144f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_A_693_113#_c_2197_n 0.00684236f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_A_693_113#_c_2198_n 0.00395819f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_A_693_113#_c_2199_n 0.0169765f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_A_693_113#_c_2200_n 0.0086414f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_A_693_113#_c_2201_n 0.008346f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_A_693_113#_c_2202_n 0.0230602f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB N_A_693_113#_c_2203_n 0.0138055f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VNB N_Q_c_2373_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_Q_c_2374_n 0.0021782f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_141 VNB N_Q_c_2375_n 0.00244365f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.145
cc_142 VNB Q 0.00910163f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.145
cc_143 VNB N_VGND_c_2406_n 0.0134339f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_144 VNB N_VGND_c_2407_n 0.0186543f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_145 VNB N_VGND_c_2408_n 0.00748215f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_146 VNB N_VGND_c_2409_n 0.0145323f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_147 VNB N_VGND_c_2410_n 0.0177254f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_148 VNB N_VGND_c_2411_n 0.0109527f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_149 VNB N_VGND_c_2412_n 0.00590394f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_150 VNB N_VGND_c_2413_n 0.0149399f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_151 VNB N_VGND_c_2414_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_152 VNB N_VGND_c_2415_n 0.0463778f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_153 VNB N_VGND_c_2416_n 0.0297887f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_154 VNB N_VGND_c_2417_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_155 VNB N_VGND_c_2418_n 0.0318151f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_156 VNB N_VGND_c_2419_n 0.0196191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_157 VNB N_VGND_c_2420_n 0.0701939f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_158 VNB N_VGND_c_2421_n 0.0204536f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_159 VNB N_VGND_c_2422_n 0.0658283f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_160 VNB N_VGND_c_2423_n 0.0314465f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_161 VNB N_VGND_c_2424_n 0.0206041f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_162 VNB N_VGND_c_2425_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_163 VNB N_VGND_c_2426_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_164 VNB N_VGND_c_2427_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_165 VNB N_VGND_c_2428_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_166 VNB N_VGND_c_2429_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_167 VNB N_VGND_c_2430_n 0.00509721f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_168 VNB N_VGND_c_2431_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_169 VNB N_VGND_c_2432_n 0.0392213f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_170 VNB N_VGND_c_2433_n 0.030707f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_171 VNB N_VGND_c_2434_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_172 VNB N_VGND_c_2435_n 0.887438f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_173 VPB N_D_c_339_n 0.00981639f $X=-0.19 $Y=1.66 $X2=0.57 $Y2=2.155
cc_174 VPB N_D_c_340_n 0.0256345f $X=-0.19 $Y=1.66 $X2=0.57 $Y2=2.245
cc_175 VPB N_D_c_337_n 0.00427155f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=1.145
cc_176 VPB N_D_c_338_n 0.0112525f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=1.825
cc_177 VPB N_D_c_343_n 0.0156029f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=1.99
cc_178 VPB N_A_180_290#_c_385_n 0.0184393f $X=-0.19 $Y=1.66 $X2=0.615 $Y2=0.58
cc_179 VPB N_A_180_290#_c_386_n 0.0312105f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_180 VPB N_A_180_290#_c_379_n 0.0211145f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=1.145
cc_181 VPB N_A_180_290#_c_388_n 0.0120947f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=1.825
cc_182 VPB N_A_180_290#_c_389_n 0.00210347f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=1.99
cc_183 VPB N_A_180_290#_c_390_n 0.00254697f $X=-0.19 $Y=1.66 $X2=0.615 $Y2=1.825
cc_184 VPB N_A_180_290#_c_391_n 0.01375f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_185 VPB N_A_180_290#_c_383_n 0.00545274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_186 VPB N_A_180_290#_c_384_n 0.0210867f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_187 VPB N_DE_c_487_n 0.0236617f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=1.145
cc_188 VPB N_DE_c_493_n 0.0165624f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=0.98
cc_189 VPB N_DE_c_494_n 0.0118692f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_190 VPB N_DE_c_495_n 0.0183363f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=1.825
cc_191 VPB N_DE_c_496_n 0.0349079f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=1.145
cc_192 VPB N_DE_c_497_n 0.0161255f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=1.825
cc_193 VPB N_DE_c_498_n 0.00428187f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_194 VPB N_DE_c_499_n 0.00316864f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_195 VPB N_A_548_87#_c_590_n 0.0255862f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_196 VPB N_A_548_87#_c_591_n 0.0212328f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_197 VPB N_A_548_87#_c_592_n 0.054811f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=1.825
cc_198 VPB N_A_548_87#_c_581_n 0.0190144f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_199 VPB N_A_548_87#_c_594_n 0.00545435f $X=-0.19 $Y=1.66 $X2=0.615 $Y2=1.295
cc_200 VPB N_A_548_87#_c_595_n 0.0115835f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_201 VPB N_A_548_87#_c_596_n 0.00289649f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_202 VPB N_A_548_87#_c_597_n 0.0107564f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_203 VPB N_A_548_87#_c_598_n 5.2388e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_204 VPB N_A_548_87#_c_585_n 0.0711649f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_205 VPB N_A_548_87#_c_586_n 5.99535e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_206 VPB N_A_548_87#_c_601_n 0.00219825f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_207 VPB N_A_548_87#_c_587_n 0.0090202f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_208 VPB N_A_548_87#_c_588_n 0.00243538f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_209 VPB N_A_548_87#_c_589_n 0.0269046f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_210 VPB N_A_663_87#_c_839_n 0.0175717f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_211 VPB N_A_663_87#_c_840_n 0.0231189f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=1.145
cc_212 VPB N_A_663_87#_c_835_n 0.0334036f $X=-0.19 $Y=1.66 $X2=0.615 $Y2=1.665
cc_213 VPB N_A_663_87#_c_842_n 0.00470336f $X=-0.19 $Y=1.66 $X2=0.615 $Y2=1.825
cc_214 VPB N_A_663_87#_c_843_n 0.01966f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_215 VPB N_A_663_87#_c_837_n 0.0191866f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_216 VPB N_A_663_87#_c_845_n 0.00599833f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_217 VPB N_A_663_87#_c_846_n 0.00872009f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_218 VPB N_SCD_c_942_n 0.020419f $X=-0.19 $Y=1.66 $X2=0.615 $Y2=0.98
cc_219 VPB N_SCD_c_943_n 0.0218708f $X=-0.19 $Y=1.66 $X2=0.615 $Y2=0.58
cc_220 VPB SCD 0.00336543f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=1.145
cc_221 VPB N_SCD_c_941_n 0.00959716f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_222 VPB N_SCE_c_989_n 0.0185503f $X=-0.19 $Y=1.66 $X2=0.57 $Y2=1.99
cc_223 VPB N_SCE_c_990_n 0.0824846f $X=-0.19 $Y=1.66 $X2=0.57 $Y2=2.64
cc_224 VPB N_SCE_c_991_n 0.0132883f $X=-0.19 $Y=1.66 $X2=0.57 $Y2=2.64
cc_225 VPB N_SCE_c_982_n 0.0277783f $X=-0.19 $Y=1.66 $X2=0.615 $Y2=0.58
cc_226 VPB N_SCE_c_993_n 0.00747999f $X=-0.19 $Y=1.66 $X2=0.615 $Y2=0.58
cc_227 VPB N_SCE_M1003_g 0.00951438f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=0.98
cc_228 VPB N_CLK_c_1068_n 0.0287024f $X=-0.19 $Y=1.66 $X2=0.57 $Y2=2.64
cc_229 VPB N_A_1538_74#_c_1126_n 0.0194459f $X=-0.19 $Y=1.66 $X2=0.615 $Y2=0.58
cc_230 VPB N_A_1538_74#_c_1103_n 0.0377235f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=1.145
cc_231 VPB N_A_1538_74#_c_1128_n 0.0220217f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=1.145
cc_232 VPB N_A_1538_74#_c_1129_n 0.00348725f $X=-0.19 $Y=1.66 $X2=0.615
+ $Y2=1.665
cc_233 VPB N_A_1538_74#_c_1107_n 0.00101962f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_234 VPB N_A_1538_74#_c_1116_n 0.00531976f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_235 VPB N_A_1538_74#_c_1117_n 0.0182276f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_236 VPB N_A_1538_74#_c_1133_n 0.00925755f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_237 VPB N_A_1538_74#_c_1134_n 0.057484f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_238 VPB N_A_1340_74#_c_1339_n 0.0101509f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_239 VPB N_A_1340_74#_c_1354_n 0.0211204f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_240 VPB N_A_1340_74#_c_1340_n 0.00853083f $X=-0.19 $Y=1.66 $X2=0.525
+ $Y2=1.145
cc_241 VPB N_A_1340_74#_c_1342_n 0.0269179f $X=-0.19 $Y=1.66 $X2=0.615 $Y2=1.145
cc_242 VPB N_A_1340_74#_c_1357_n 0.0156382f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_243 VPB N_A_1340_74#_c_1358_n 0.0583143f $X=-0.19 $Y=1.66 $X2=0.615 $Y2=1.665
cc_244 VPB N_A_1340_74#_c_1343_n 0.0440313f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_245 VPB N_A_1340_74#_c_1345_n 0.00167153f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_246 VPB N_A_1340_74#_c_1346_n 0.00543223f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_247 VPB N_A_1340_74#_c_1362_n 0.0178838f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_248 VPB N_A_1340_74#_c_1363_n 0.00578836f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_249 VPB N_A_1340_74#_c_1350_n 0.00460109f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_250 VPB N_A_1340_74#_c_1351_n 0.0534049f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_251 VPB N_A_1340_74#_c_1366_n 0.00799871f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_252 VPB N_A_1340_74#_c_1352_n 0.0016284f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_253 VPB N_A_1979_71#_c_1527_n 0.0410266f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_254 VPB N_A_1979_71#_c_1540_n 0.0231982f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_255 VPB N_A_1979_71#_c_1529_n 0.00873471f $X=-0.19 $Y=1.66 $X2=0.525
+ $Y2=1.145
cc_256 VPB N_A_1979_71#_c_1542_n 0.0330378f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=1.825
cc_257 VPB N_A_1979_71#_c_1533_n 0.00941663f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_258 VPB N_A_1979_71#_c_1544_n 0.00355131f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_259 VPB N_A_1736_97#_c_1632_n 0.0419806f $X=-0.19 $Y=1.66 $X2=0.615 $Y2=0.58
cc_260 VPB N_A_1736_97#_c_1636_n 0.0169703f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=1.825
cc_261 VPB N_A_1736_97#_c_1637_n 0.00322281f $X=-0.19 $Y=1.66 $X2=0.525
+ $Y2=1.825
cc_262 VPB N_A_1736_97#_c_1638_n 0.0086284f $X=-0.19 $Y=1.66 $X2=0.615 $Y2=1.295
cc_263 VPB N_A_1736_97#_c_1639_n 0.00920798f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_264 VPB N_A_1736_97#_c_1640_n 0.00223518f $X=-0.19 $Y=1.66 $X2=0.615
+ $Y2=1.825
cc_265 VPB N_A_2474_74#_c_1729_n 0.0189516f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=0.98
cc_266 VPB N_A_2474_74#_c_1730_n 0.0177175f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=1.825
cc_267 VPB N_A_2474_74#_c_1731_n 0.0174832f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_268 VPB N_A_2474_74#_c_1732_n 0.0269336f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_269 VPB N_A_2474_74#_c_1722_n 0.0159257f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_270 VPB N_A_2474_74#_c_1734_n 0.00225496f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_271 VPB N_A_2474_74#_c_1735_n 0.0104172f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_272 VPB N_A_2474_74#_c_1736_n 0.00414133f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_273 VPB N_A_2474_74#_c_1726_n 0.00116664f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_274 VPB N_A_2474_74#_c_1738_n 0.00543964f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_275 VPB N_A_2474_74#_c_1739_n 4.15279e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_276 VPB N_A_2474_74#_c_1727_n 0.00158659f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_277 VPB N_A_2474_74#_c_1728_n 0.0223927f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_278 VPB N_A_40_464#_c_1885_n 0.0302944f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_279 VPB N_A_40_464#_c_1892_n 0.0257246f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=1.145
cc_280 VPB N_A_40_464#_c_1893_n 0.0160391f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=1.145
cc_281 VPB N_A_40_464#_c_1894_n 0.00998336f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=1.825
cc_282 VPB N_A_40_464#_c_1895_n 0.00788509f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=1.99
cc_283 VPB N_A_40_464#_c_1896_n 0.00349119f $X=-0.19 $Y=1.66 $X2=0.615 $Y2=1.145
cc_284 VPB N_A_40_464#_c_1897_n 0.00539904f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_285 VPB N_A_40_464#_c_1898_n 8.46064e-19 $X=-0.19 $Y=1.66 $X2=0.615 $Y2=1.665
cc_286 VPB N_A_40_464#_c_1899_n 0.00216571f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_287 VPB N_A_40_464#_c_1887_n 0.0127153f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_288 VPB N_A_40_464#_c_1901_n 0.0134314f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_289 VPB N_A_40_464#_c_1902_n 0.00125429f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_290 VPB N_VPWR_c_2014_n 0.00600898f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_291 VPB N_VPWR_c_2015_n 0.00554607f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_292 VPB N_VPWR_c_2016_n 0.00745483f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_293 VPB N_VPWR_c_2017_n 0.0114885f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_294 VPB N_VPWR_c_2018_n 0.0197665f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_295 VPB N_VPWR_c_2019_n 0.0114729f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_296 VPB N_VPWR_c_2020_n 0.0139022f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_297 VPB N_VPWR_c_2021_n 0.00880467f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_298 VPB N_VPWR_c_2022_n 0.0152675f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_299 VPB N_VPWR_c_2023_n 0.0120106f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_300 VPB N_VPWR_c_2024_n 0.0342038f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_301 VPB N_VPWR_c_2025_n 0.0242802f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_302 VPB N_VPWR_c_2026_n 0.00633387f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_303 VPB N_VPWR_c_2027_n 0.0618187f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_304 VPB N_VPWR_c_2028_n 0.0101806f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_305 VPB N_VPWR_c_2029_n 0.0320939f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_306 VPB N_VPWR_c_2030_n 0.0296515f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_307 VPB N_VPWR_c_2031_n 0.0586722f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_308 VPB N_VPWR_c_2032_n 0.0325948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_309 VPB N_VPWR_c_2033_n 0.0336414f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_310 VPB N_VPWR_c_2034_n 0.0604054f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_311 VPB N_VPWR_c_2035_n 0.0204479f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_312 VPB N_VPWR_c_2036_n 0.0163251f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_313 VPB N_VPWR_c_2037_n 0.00460249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_314 VPB N_VPWR_c_2038_n 0.00463855f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_315 VPB N_VPWR_c_2039_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_316 VPB N_VPWR_c_2040_n 0.00638292f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_317 VPB N_VPWR_c_2041_n 0.00614248f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_318 VPB N_VPWR_c_2042_n 0.00614151f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_319 VPB N_VPWR_c_2043_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_320 VPB N_VPWR_c_2013_n 0.210496f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_321 VPB N_A_693_113#_c_2204_n 0.0023497f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=1.825
cc_322 VPB N_A_693_113#_c_2205_n 0.00747967f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_323 VPB N_A_693_113#_c_2206_n 0.013184f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_324 VPB N_A_693_113#_c_2207_n 0.00104828f $X=-0.19 $Y=1.66 $X2=0.615
+ $Y2=1.825
cc_325 VPB N_A_693_113#_c_2208_n 0.0305569f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_326 VPB N_A_693_113#_c_2209_n 0.00111746f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_327 VPB N_A_693_113#_c_2210_n 0.00888537f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_328 VPB N_A_693_113#_c_2211_n 0.00664178f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_329 VPB N_A_693_113#_c_2201_n 0.010433f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_330 VPB N_A_693_113#_c_2203_n 0.0141093f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_331 VPB N_A_693_113#_c_2214_n 0.0075629f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_332 VPB N_Q_c_2377_n 0.00247218f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_333 VPB Q 0.0222499f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=1.145
cc_334 N_D_c_340_n N_A_180_290#_c_385_n 0.0383515f $X=0.57 $Y=2.245 $X2=0 $Y2=0
cc_335 N_D_c_339_n N_A_180_290#_c_386_n 0.0143143f $X=0.57 $Y=2.155 $X2=0 $Y2=0
cc_336 N_D_c_343_n N_A_180_290#_c_386_n 0.0169395f $X=0.525 $Y=1.99 $X2=0 $Y2=0
cc_337 N_D_c_337_n N_A_180_290#_c_378_n 0.0649021f $X=0.525 $Y=1.145 $X2=0 $Y2=0
cc_338 N_D_c_338_n N_A_180_290#_c_378_n 0.00183375f $X=0.525 $Y=1.825 $X2=0
+ $Y2=0
cc_339 N_D_c_337_n N_A_180_290#_c_379_n 0.00368273f $X=0.525 $Y=1.145 $X2=0
+ $Y2=0
cc_340 N_D_c_338_n N_A_180_290#_c_379_n 0.0169395f $X=0.525 $Y=1.825 $X2=0 $Y2=0
cc_341 N_D_c_337_n N_A_180_290#_c_381_n 0.0143758f $X=0.525 $Y=1.145 $X2=0 $Y2=0
cc_342 N_D_c_339_n N_A_180_290#_c_389_n 7.16047e-19 $X=0.57 $Y=2.155 $X2=0 $Y2=0
cc_343 N_D_c_337_n N_A_180_290#_c_389_n 0.00339233f $X=0.525 $Y=1.145 $X2=0
+ $Y2=0
cc_344 N_D_M1005_g N_DE_M1029_g 0.0249654f $X=0.615 $Y=0.58 $X2=0 $Y2=0
cc_345 N_D_c_337_n N_DE_M1029_g 0.00159522f $X=0.525 $Y=1.145 $X2=0 $Y2=0
cc_346 N_D_c_336_n N_DE_c_486_n 0.0249654f $X=0.525 $Y=1.145 $X2=0 $Y2=0
cc_347 N_D_c_339_n N_A_40_464#_c_1885_n 0.00836819f $X=0.57 $Y=2.155 $X2=0 $Y2=0
cc_348 N_D_c_340_n N_A_40_464#_c_1885_n 0.00139731f $X=0.57 $Y=2.245 $X2=0 $Y2=0
cc_349 N_D_M1005_g N_A_40_464#_c_1885_n 0.00513151f $X=0.615 $Y=0.58 $X2=0 $Y2=0
cc_350 N_D_c_336_n N_A_40_464#_c_1885_n 0.024408f $X=0.525 $Y=1.145 $X2=0 $Y2=0
cc_351 N_D_c_337_n N_A_40_464#_c_1885_n 0.0766522f $X=0.525 $Y=1.145 $X2=0 $Y2=0
cc_352 N_D_c_340_n N_A_40_464#_c_1892_n 0.00947726f $X=0.57 $Y=2.245 $X2=0 $Y2=0
cc_353 N_D_c_340_n N_A_40_464#_c_1893_n 0.0127112f $X=0.57 $Y=2.245 $X2=0 $Y2=0
cc_354 N_D_c_337_n N_A_40_464#_c_1893_n 0.0153217f $X=0.525 $Y=1.145 $X2=0 $Y2=0
cc_355 N_D_M1005_g N_A_40_464#_c_1888_n 0.00972913f $X=0.615 $Y=0.58 $X2=0 $Y2=0
cc_356 N_D_c_336_n N_A_40_464#_c_1888_n 0.00389045f $X=0.525 $Y=1.145 $X2=0
+ $Y2=0
cc_357 N_D_c_337_n N_A_40_464#_c_1888_n 0.0118563f $X=0.525 $Y=1.145 $X2=0 $Y2=0
cc_358 N_D_c_340_n N_A_40_464#_c_1901_n 0.00164304f $X=0.57 $Y=2.245 $X2=0 $Y2=0
cc_359 N_D_c_337_n N_A_40_464#_c_1901_n 0.00482473f $X=0.525 $Y=1.145 $X2=0
+ $Y2=0
cc_360 N_D_c_343_n N_A_40_464#_c_1901_n 0.00315876f $X=0.525 $Y=1.99 $X2=0 $Y2=0
cc_361 N_D_c_340_n N_VPWR_c_2014_n 0.001556f $X=0.57 $Y=2.245 $X2=0 $Y2=0
cc_362 N_D_c_340_n N_VPWR_c_2029_n 0.00445602f $X=0.57 $Y=2.245 $X2=0 $Y2=0
cc_363 N_D_c_340_n N_VPWR_c_2013_n 0.00861848f $X=0.57 $Y=2.245 $X2=0 $Y2=0
cc_364 N_D_M1005_g N_VGND_c_2406_n 0.00186675f $X=0.615 $Y=0.58 $X2=0 $Y2=0
cc_365 N_D_M1005_g N_VGND_c_2418_n 0.00433162f $X=0.615 $Y=0.58 $X2=0 $Y2=0
cc_366 N_D_M1005_g N_VGND_c_2435_n 0.00821332f $X=0.615 $Y=0.58 $X2=0 $Y2=0
cc_367 N_A_180_290#_c_381_n N_DE_M1029_g 0.00767961f $X=1.305 $Y=1.065 $X2=0
+ $Y2=0
cc_368 N_A_180_290#_c_382_n N_DE_M1029_g 0.00465695f $X=1.78 $Y=0.775 $X2=0
+ $Y2=0
cc_369 N_A_180_290#_c_378_n N_DE_c_485_n 0.0063489f $X=1.14 $Y=1.615 $X2=0 $Y2=0
cc_370 N_A_180_290#_c_380_n N_DE_c_485_n 0.012769f $X=1.615 $Y=1.065 $X2=0 $Y2=0
cc_371 N_A_180_290#_c_381_n N_DE_c_485_n 0.00402704f $X=1.305 $Y=1.065 $X2=0
+ $Y2=0
cc_372 N_A_180_290#_c_378_n N_DE_c_486_n 0.00199694f $X=1.14 $Y=1.615 $X2=0
+ $Y2=0
cc_373 N_A_180_290#_c_379_n N_DE_c_486_n 0.0215668f $X=1.14 $Y=1.615 $X2=0 $Y2=0
cc_374 N_A_180_290#_c_381_n N_DE_c_486_n 0.001395f $X=1.305 $Y=1.065 $X2=0 $Y2=0
cc_375 N_A_180_290#_c_378_n N_DE_c_487_n 0.00113204f $X=1.14 $Y=1.615 $X2=0
+ $Y2=0
cc_376 N_A_180_290#_c_379_n N_DE_c_487_n 0.00793894f $X=1.14 $Y=1.615 $X2=0
+ $Y2=0
cc_377 N_A_180_290#_c_388_n N_DE_c_487_n 0.00579788f $X=1.81 $Y=2.035 $X2=0
+ $Y2=0
cc_378 N_A_180_290#_c_391_n N_DE_c_487_n 0.00331704f $X=2.22 $Y=1.95 $X2=0 $Y2=0
cc_379 N_A_180_290#_c_383_n N_DE_c_487_n 0.00405247f $X=2.22 $Y=1.685 $X2=0
+ $Y2=0
cc_380 N_A_180_290#_c_384_n N_DE_c_487_n 0.0110148f $X=2.425 $Y=1.685 $X2=0
+ $Y2=0
cc_381 N_A_180_290#_c_390_n N_DE_c_493_n 0.0113241f $X=1.895 $Y=2.515 $X2=0
+ $Y2=0
cc_382 N_A_180_290#_c_391_n N_DE_c_493_n 0.00730631f $X=2.22 $Y=1.95 $X2=0 $Y2=0
cc_383 N_A_180_290#_c_386_n N_DE_c_494_n 0.0114968f $X=1.102 $Y=1.918 $X2=0
+ $Y2=0
cc_384 N_A_180_290#_c_388_n N_DE_c_494_n 0.00629372f $X=1.81 $Y=2.035 $X2=0
+ $Y2=0
cc_385 N_A_180_290#_c_390_n N_DE_c_494_n 0.00464691f $X=1.895 $Y=2.515 $X2=0
+ $Y2=0
cc_386 N_A_180_290#_M1015_g N_DE_c_488_n 0.0188666f $X=2.425 $Y=0.775 $X2=0
+ $Y2=0
cc_387 N_A_180_290#_c_380_n N_DE_c_488_n 0.00310065f $X=1.615 $Y=1.065 $X2=0
+ $Y2=0
cc_388 N_A_180_290#_c_382_n N_DE_c_488_n 9.22767e-19 $X=1.78 $Y=0.775 $X2=0
+ $Y2=0
cc_389 N_A_180_290#_c_390_n N_DE_c_495_n 0.00415054f $X=1.895 $Y=2.515 $X2=0
+ $Y2=0
cc_390 N_A_180_290#_c_391_n N_DE_c_496_n 0.00514267f $X=2.22 $Y=1.95 $X2=0 $Y2=0
cc_391 N_A_180_290#_c_380_n N_DE_c_489_n 0.0165235f $X=1.615 $Y=1.065 $X2=0
+ $Y2=0
cc_392 N_A_180_290#_c_384_n N_DE_c_489_n 6.31753e-19 $X=2.425 $Y=1.685 $X2=0
+ $Y2=0
cc_393 N_A_180_290#_c_391_n N_DE_c_498_n 0.00669704f $X=2.22 $Y=1.95 $X2=0 $Y2=0
cc_394 N_A_180_290#_c_383_n N_DE_c_498_n 3.19241e-19 $X=2.22 $Y=1.685 $X2=0
+ $Y2=0
cc_395 N_A_180_290#_c_384_n N_DE_c_498_n 0.0251598f $X=2.425 $Y=1.685 $X2=0
+ $Y2=0
cc_396 N_A_180_290#_M1015_g N_DE_c_490_n 0.00863509f $X=2.425 $Y=0.775 $X2=0
+ $Y2=0
cc_397 N_A_180_290#_c_378_n N_DE_c_490_n 0.00782514f $X=1.14 $Y=1.615 $X2=0
+ $Y2=0
cc_398 N_A_180_290#_c_379_n N_DE_c_490_n 0.0123493f $X=1.14 $Y=1.615 $X2=0 $Y2=0
cc_399 N_A_180_290#_M1015_g N_DE_c_499_n 0.00106172f $X=2.425 $Y=0.775 $X2=0
+ $Y2=0
cc_400 N_A_180_290#_c_378_n N_DE_c_499_n 0.0302117f $X=1.14 $Y=1.615 $X2=0 $Y2=0
cc_401 N_A_180_290#_c_379_n N_DE_c_499_n 0.00172549f $X=1.14 $Y=1.615 $X2=0
+ $Y2=0
cc_402 N_A_180_290#_c_380_n N_DE_c_499_n 0.0259217f $X=1.615 $Y=1.065 $X2=0
+ $Y2=0
cc_403 N_A_180_290#_c_388_n N_DE_c_499_n 0.0255862f $X=1.81 $Y=2.035 $X2=0 $Y2=0
cc_404 N_A_180_290#_c_383_n N_DE_c_499_n 0.0170229f $X=2.22 $Y=1.685 $X2=0 $Y2=0
cc_405 N_A_180_290#_c_384_n N_DE_c_499_n 0.00129966f $X=2.425 $Y=1.685 $X2=0
+ $Y2=0
cc_406 N_A_180_290#_c_388_n N_DE_c_491_n 7.51173e-19 $X=1.81 $Y=2.035 $X2=0
+ $Y2=0
cc_407 N_A_180_290#_c_383_n N_DE_c_491_n 4.52778e-19 $X=2.22 $Y=1.685 $X2=0
+ $Y2=0
cc_408 N_A_180_290#_c_384_n N_DE_c_491_n 0.00810547f $X=2.425 $Y=1.685 $X2=0
+ $Y2=0
cc_409 N_A_180_290#_M1015_g N_A_548_87#_M1025_g 0.0382648f $X=2.425 $Y=0.775
+ $X2=0 $Y2=0
cc_410 N_A_180_290#_c_383_n N_A_548_87#_c_586_n 0.00678737f $X=2.22 $Y=1.685
+ $X2=0 $Y2=0
cc_411 N_A_180_290#_c_384_n N_A_548_87#_c_586_n 0.00348757f $X=2.425 $Y=1.685
+ $X2=0 $Y2=0
cc_412 N_A_180_290#_M1015_g N_A_548_87#_c_588_n 0.00234571f $X=2.425 $Y=0.775
+ $X2=0 $Y2=0
cc_413 N_A_180_290#_c_383_n N_A_548_87#_c_588_n 0.0230712f $X=2.22 $Y=1.685
+ $X2=0 $Y2=0
cc_414 N_A_180_290#_c_383_n N_A_548_87#_c_589_n 2.4687e-19 $X=2.22 $Y=1.685
+ $X2=0 $Y2=0
cc_415 N_A_180_290#_c_384_n N_A_548_87#_c_589_n 0.0382648f $X=2.425 $Y=1.685
+ $X2=0 $Y2=0
cc_416 N_A_180_290#_c_385_n N_A_40_464#_c_1892_n 0.00181946f $X=0.99 $Y=2.245
+ $X2=0 $Y2=0
cc_417 N_A_180_290#_c_385_n N_A_40_464#_c_1893_n 0.0180284f $X=0.99 $Y=2.245
+ $X2=0 $Y2=0
cc_418 N_A_180_290#_c_386_n N_A_40_464#_c_1893_n 0.00273833f $X=1.102 $Y=1.918
+ $X2=0 $Y2=0
cc_419 N_A_180_290#_c_388_n N_A_40_464#_c_1893_n 0.0267076f $X=1.81 $Y=2.035
+ $X2=0 $Y2=0
cc_420 N_A_180_290#_c_389_n N_A_40_464#_c_1893_n 0.0259512f $X=1.305 $Y=2.035
+ $X2=0 $Y2=0
cc_421 N_A_180_290#_c_390_n N_A_40_464#_c_1893_n 0.0141649f $X=1.895 $Y=2.515
+ $X2=0 $Y2=0
cc_422 N_A_180_290#_c_385_n N_A_40_464#_c_1894_n 0.00426176f $X=0.99 $Y=2.245
+ $X2=0 $Y2=0
cc_423 N_A_180_290#_c_390_n N_A_40_464#_c_1894_n 0.0203028f $X=1.895 $Y=2.515
+ $X2=0 $Y2=0
cc_424 N_A_180_290#_M1038_s N_A_40_464#_c_1895_n 0.00320543f $X=1.75 $Y=2.315
+ $X2=0 $Y2=0
cc_425 N_A_180_290#_c_390_n N_A_40_464#_c_1895_n 0.0126885f $X=1.895 $Y=2.515
+ $X2=0 $Y2=0
cc_426 N_A_180_290#_c_385_n N_A_40_464#_c_1896_n 6.5162e-19 $X=0.99 $Y=2.245
+ $X2=0 $Y2=0
cc_427 N_A_180_290#_c_390_n N_A_40_464#_c_1928_n 0.0192722f $X=1.895 $Y=2.515
+ $X2=0 $Y2=0
cc_428 N_A_180_290#_c_391_n N_A_40_464#_c_1897_n 0.00461079f $X=2.22 $Y=1.95
+ $X2=0 $Y2=0
cc_429 N_A_180_290#_c_390_n N_A_40_464#_c_1898_n 0.0133944f $X=1.895 $Y=2.515
+ $X2=0 $Y2=0
cc_430 N_A_180_290#_c_391_n N_A_40_464#_c_1898_n 0.0134805f $X=2.22 $Y=1.95
+ $X2=0 $Y2=0
cc_431 N_A_180_290#_M1015_g N_A_40_464#_c_1889_n 9.2741e-19 $X=2.425 $Y=0.775
+ $X2=0 $Y2=0
cc_432 N_A_180_290#_c_385_n N_VPWR_c_2014_n 0.0107235f $X=0.99 $Y=2.245 $X2=0
+ $Y2=0
cc_433 N_A_180_290#_c_385_n N_VPWR_c_2029_n 0.00413917f $X=0.99 $Y=2.245 $X2=0
+ $Y2=0
cc_434 N_A_180_290#_c_385_n N_VPWR_c_2013_n 0.00817532f $X=0.99 $Y=2.245 $X2=0
+ $Y2=0
cc_435 N_A_180_290#_c_380_n N_VGND_c_2406_n 0.00663369f $X=1.615 $Y=1.065 $X2=0
+ $Y2=0
cc_436 N_A_180_290#_c_381_n N_VGND_c_2406_n 0.0231121f $X=1.305 $Y=1.065 $X2=0
+ $Y2=0
cc_437 N_A_180_290#_c_382_n N_VGND_c_2406_n 0.0174982f $X=1.78 $Y=0.775 $X2=0
+ $Y2=0
cc_438 N_A_180_290#_M1015_g N_VGND_c_2407_n 0.0130041f $X=2.425 $Y=0.775 $X2=0
+ $Y2=0
cc_439 N_A_180_290#_c_380_n N_VGND_c_2407_n 0.00175056f $X=1.615 $Y=1.065 $X2=0
+ $Y2=0
cc_440 N_A_180_290#_c_382_n N_VGND_c_2407_n 0.0163189f $X=1.78 $Y=0.775 $X2=0
+ $Y2=0
cc_441 N_A_180_290#_c_383_n N_VGND_c_2407_n 0.0117414f $X=2.22 $Y=1.685 $X2=0
+ $Y2=0
cc_442 N_A_180_290#_c_384_n N_VGND_c_2407_n 0.00187021f $X=2.425 $Y=1.685 $X2=0
+ $Y2=0
cc_443 N_A_180_290#_c_382_n N_VGND_c_2419_n 0.00607888f $X=1.78 $Y=0.775 $X2=0
+ $Y2=0
cc_444 N_A_180_290#_M1015_g N_VGND_c_2420_n 0.00372658f $X=2.425 $Y=0.775 $X2=0
+ $Y2=0
cc_445 N_A_180_290#_M1015_g N_VGND_c_2435_n 0.00408518f $X=2.425 $Y=0.775 $X2=0
+ $Y2=0
cc_446 N_A_180_290#_c_382_n N_VGND_c_2435_n 0.00799492f $X=1.78 $Y=0.775 $X2=0
+ $Y2=0
cc_447 N_DE_c_496_n N_A_548_87#_c_590_n 0.0106312f $X=2.725 $Y=2.165 $X2=0 $Y2=0
cc_448 N_DE_c_497_n N_A_548_87#_c_591_n 0.0437219f $X=2.8 $Y=2.24 $X2=0 $Y2=0
cc_449 N_DE_c_496_n N_A_548_87#_c_586_n 0.00118486f $X=2.725 $Y=2.165 $X2=0
+ $Y2=0
cc_450 N_DE_c_496_n N_A_548_87#_c_588_n 0.00522508f $X=2.725 $Y=2.165 $X2=0
+ $Y2=0
cc_451 N_DE_c_496_n N_A_548_87#_c_589_n 0.00880655f $X=2.725 $Y=2.165 $X2=0
+ $Y2=0
cc_452 N_DE_c_495_n N_A_40_464#_c_1894_n 0.00326422f $X=2.12 $Y=2.24 $X2=0 $Y2=0
cc_453 N_DE_c_493_n N_A_40_464#_c_1895_n 7.52982e-19 $X=2.045 $Y=2.165 $X2=0
+ $Y2=0
cc_454 N_DE_c_494_n N_A_40_464#_c_1895_n 0.00408551f $X=1.815 $Y=2.165 $X2=0
+ $Y2=0
cc_455 N_DE_c_495_n N_A_40_464#_c_1895_n 0.0134964f $X=2.12 $Y=2.24 $X2=0 $Y2=0
cc_456 N_DE_c_497_n N_A_40_464#_c_1895_n 4.28313e-19 $X=2.8 $Y=2.24 $X2=0 $Y2=0
cc_457 N_DE_c_495_n N_A_40_464#_c_1928_n 0.0118088f $X=2.12 $Y=2.24 $X2=0 $Y2=0
cc_458 N_DE_c_497_n N_A_40_464#_c_1928_n 0.00283455f $X=2.8 $Y=2.24 $X2=0 $Y2=0
cc_459 N_DE_c_496_n N_A_40_464#_c_1897_n 0.0105127f $X=2.725 $Y=2.165 $X2=0
+ $Y2=0
cc_460 N_DE_c_497_n N_A_40_464#_c_1897_n 0.0155117f $X=2.8 $Y=2.24 $X2=0 $Y2=0
cc_461 N_DE_c_495_n N_A_40_464#_c_1898_n 0.00584584f $X=2.12 $Y=2.24 $X2=0 $Y2=0
cc_462 N_DE_c_496_n N_A_40_464#_c_1898_n 8.1141e-19 $X=2.725 $Y=2.165 $X2=0
+ $Y2=0
cc_463 N_DE_c_497_n N_A_40_464#_c_1899_n 0.00179485f $X=2.8 $Y=2.24 $X2=0 $Y2=0
cc_464 N_DE_M1029_g N_A_40_464#_c_1888_n 0.00129488f $X=1.005 $Y=0.58 $X2=0
+ $Y2=0
cc_465 N_DE_c_495_n N_VPWR_c_2015_n 0.00153478f $X=2.12 $Y=2.24 $X2=0 $Y2=0
cc_466 N_DE_c_497_n N_VPWR_c_2015_n 0.00967911f $X=2.8 $Y=2.24 $X2=0 $Y2=0
cc_467 N_DE_c_495_n N_VPWR_c_2030_n 0.00275664f $X=2.12 $Y=2.24 $X2=0 $Y2=0
cc_468 N_DE_c_497_n N_VPWR_c_2031_n 0.00410286f $X=2.8 $Y=2.24 $X2=0 $Y2=0
cc_469 N_DE_c_495_n N_VPWR_c_2013_n 0.00544287f $X=2.12 $Y=2.24 $X2=0 $Y2=0
cc_470 N_DE_c_497_n N_VPWR_c_2013_n 0.00493487f $X=2.8 $Y=2.24 $X2=0 $Y2=0
cc_471 N_DE_M1029_g N_VGND_c_2406_n 0.014051f $X=1.005 $Y=0.58 $X2=0 $Y2=0
cc_472 N_DE_c_485_n N_VGND_c_2406_n 0.00140716f $X=1.515 $Y=1.135 $X2=0 $Y2=0
cc_473 N_DE_c_488_n N_VGND_c_2406_n 0.00221288f $X=1.995 $Y=1.06 $X2=0 $Y2=0
cc_474 N_DE_c_488_n N_VGND_c_2407_n 0.0108147f $X=1.995 $Y=1.06 $X2=0 $Y2=0
cc_475 N_DE_M1029_g N_VGND_c_2418_n 0.00383152f $X=1.005 $Y=0.58 $X2=0 $Y2=0
cc_476 N_DE_c_488_n N_VGND_c_2419_n 0.00372658f $X=1.995 $Y=1.06 $X2=0 $Y2=0
cc_477 N_DE_M1029_g N_VGND_c_2435_n 0.0075725f $X=1.005 $Y=0.58 $X2=0 $Y2=0
cc_478 N_DE_c_488_n N_VGND_c_2435_n 0.00408518f $X=1.995 $Y=1.06 $X2=0 $Y2=0
cc_479 N_A_548_87#_M1025_g N_A_663_87#_c_829_n 0.0208346f $X=2.815 $Y=0.775
+ $X2=0 $Y2=0
cc_480 N_A_548_87#_c_585_n N_A_663_87#_c_830_n 0.0063913f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_481 N_A_548_87#_c_585_n N_A_663_87#_c_849_n 0.0235991f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_482 N_A_548_87#_c_585_n N_A_663_87#_c_835_n 0.00602768f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_483 N_A_548_87#_c_589_n N_A_663_87#_c_835_n 0.00503886f $X=3.19 $Y=1.68 $X2=0
+ $Y2=0
cc_484 N_A_548_87#_c_585_n N_A_663_87#_c_843_n 0.0363111f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_485 N_A_548_87#_c_585_n N_A_663_87#_c_836_n 0.0165193f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_486 N_A_548_87#_c_585_n N_A_663_87#_c_837_n 0.0039757f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_487 N_A_548_87#_c_585_n N_A_663_87#_c_838_n 0.00669559f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_488 N_A_548_87#_c_585_n N_A_663_87#_c_846_n 3.9432e-19 $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_489 N_A_548_87#_c_585_n SCD 0.0315857f $X=14.975 $Y=1.665 $X2=0 $Y2=0
cc_490 N_A_548_87#_c_585_n N_SCD_c_941_n 6.94548e-19 $X=14.975 $Y=1.665 $X2=0
+ $Y2=0
cc_491 N_A_548_87#_c_591_n N_SCE_c_989_n 0.0074134f $X=3.19 $Y=2.24 $X2=-0.19
+ $Y2=-0.245
cc_492 N_A_548_87#_c_585_n N_SCE_c_989_n 0.00250527f $X=14.975 $Y=1.665
+ $X2=-0.19 $Y2=-0.245
cc_493 N_A_548_87#_c_591_n N_SCE_c_991_n 0.00288121f $X=3.19 $Y=2.24 $X2=0 $Y2=0
cc_494 N_A_548_87#_c_585_n N_SCE_c_982_n 0.00598741f $X=14.975 $Y=1.665 $X2=0
+ $Y2=0
cc_495 N_A_548_87#_c_585_n N_SCE_M1004_g 0.00168364f $X=14.975 $Y=1.665 $X2=0
+ $Y2=0
cc_496 N_A_548_87#_c_585_n N_SCE_c_987_n 0.00436451f $X=14.975 $Y=1.665 $X2=0
+ $Y2=0
cc_497 N_A_548_87#_c_585_n N_SCE_c_988_n 0.00949212f $X=14.975 $Y=1.665 $X2=0
+ $Y2=0
cc_498 N_A_548_87#_c_585_n N_CLK_c_1068_n 0.0130241f $X=14.975 $Y=1.665 $X2=0
+ $Y2=0
cc_499 N_A_548_87#_c_585_n CLK 0.0168623f $X=14.975 $Y=1.665 $X2=0 $Y2=0
cc_500 N_A_548_87#_c_592_n N_A_1538_74#_c_1103_n 0.0196577f $X=13.63 $Y=2.465
+ $X2=0 $Y2=0
cc_501 N_A_548_87#_c_581_n N_A_1538_74#_c_1103_n 0.0141746f $X=13.765 $Y=2.05
+ $X2=0 $Y2=0
cc_502 N_A_548_87#_c_596_n N_A_1538_74#_c_1103_n 9.24008e-19 $X=13.675 $Y=2.215
+ $X2=0 $Y2=0
cc_503 N_A_548_87#_c_585_n N_A_1538_74#_c_1103_n 0.00571827f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_504 N_A_548_87#_c_592_n N_A_1538_74#_c_1128_n 0.0317522f $X=13.63 $Y=2.465
+ $X2=0 $Y2=0
cc_505 N_A_548_87#_c_596_n N_A_1538_74#_c_1128_n 5.62571e-19 $X=13.675 $Y=2.215
+ $X2=0 $Y2=0
cc_506 N_A_548_87#_c_585_n N_A_1538_74#_c_1104_n 0.00797831f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_507 N_A_548_87#_c_585_n N_A_1538_74#_c_1129_n 0.015081f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_508 N_A_548_87#_c_585_n N_A_1538_74#_c_1107_n 0.0205755f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_509 N_A_548_87#_c_585_n N_A_1538_74#_c_1109_n 0.0059249f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_510 N_A_548_87#_c_585_n N_A_1538_74#_c_1113_n 0.00739409f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_511 N_A_548_87#_c_585_n N_A_1538_74#_c_1116_n 0.041172f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_512 N_A_548_87#_c_585_n N_A_1538_74#_c_1117_n 0.00147662f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_513 N_A_548_87#_c_580_n N_A_1538_74#_c_1118_n 2.40283e-19 $X=13.235 $Y=0.94
+ $X2=0 $Y2=0
cc_514 N_A_548_87#_c_585_n N_A_1538_74#_c_1118_n 0.01616f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_515 N_A_548_87#_c_585_n N_A_1538_74#_c_1133_n 0.00623863f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_516 N_A_548_87#_c_585_n N_A_1538_74#_c_1120_n 0.00832911f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_517 N_A_548_87#_c_585_n N_A_1538_74#_c_1122_n 0.00151598f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_518 N_A_548_87#_c_580_n N_A_1538_74#_c_1124_n 0.0011337f $X=13.235 $Y=0.94
+ $X2=0 $Y2=0
cc_519 N_A_548_87#_c_581_n N_A_1538_74#_c_1124_n 7.75578e-19 $X=13.765 $Y=2.05
+ $X2=0 $Y2=0
cc_520 N_A_548_87#_c_585_n N_A_1538_74#_c_1124_n 0.00932399f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_521 N_A_548_87#_c_580_n N_A_1538_74#_c_1125_n 0.0181563f $X=13.235 $Y=0.94
+ $X2=0 $Y2=0
cc_522 N_A_548_87#_c_581_n N_A_1538_74#_c_1125_n 0.0173139f $X=13.765 $Y=2.05
+ $X2=0 $Y2=0
cc_523 N_A_548_87#_c_585_n N_A_1340_74#_c_1339_n 0.010523f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_524 N_A_548_87#_c_585_n N_A_1340_74#_c_1340_n 0.00452786f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_525 N_A_548_87#_c_585_n N_A_1340_74#_c_1342_n 0.00377856f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_526 N_A_548_87#_c_585_n N_A_1340_74#_c_1343_n 6.94548e-19 $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_527 N_A_548_87#_c_578_n N_A_1340_74#_M1020_g 0.04003f $X=13.16 $Y=0.865 $X2=0
+ $Y2=0
cc_528 N_A_548_87#_c_585_n N_A_1340_74#_c_1345_n 0.00567161f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_529 N_A_548_87#_c_585_n N_A_1340_74#_c_1346_n 0.00559008f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_530 N_A_548_87#_c_585_n N_A_1340_74#_c_1348_n 0.00152612f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_531 N_A_548_87#_c_585_n N_A_1340_74#_c_1363_n 0.00308541f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_532 N_A_548_87#_c_585_n N_A_1340_74#_c_1349_n 0.00574496f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_533 N_A_548_87#_c_585_n N_A_1340_74#_c_1350_n 0.0705059f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_534 N_A_548_87#_c_585_n N_A_1340_74#_c_1351_n 0.00518971f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_535 N_A_548_87#_c_585_n N_A_1340_74#_c_1366_n 0.00220897f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_536 N_A_548_87#_c_585_n N_A_1340_74#_c_1352_n 0.0238337f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_537 N_A_548_87#_c_585_n N_A_1979_71#_c_1527_n 0.0023931f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_538 N_A_548_87#_c_585_n N_A_1979_71#_c_1528_n 0.00494526f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_539 N_A_548_87#_c_585_n N_A_1979_71#_c_1529_n 0.0127614f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_540 N_A_548_87#_c_585_n N_A_1979_71#_c_1531_n 0.0109985f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_541 N_A_548_87#_c_585_n N_A_1979_71#_c_1533_n 0.0201256f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_542 N_A_548_87#_c_585_n N_A_1979_71#_c_1534_n 0.0327997f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_543 N_A_548_87#_c_585_n N_A_1979_71#_c_1535_n 0.0129863f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_544 N_A_548_87#_c_585_n N_A_1979_71#_c_1536_n 0.00824337f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_545 N_A_548_87#_c_585_n N_A_1979_71#_c_1544_n 0.00737978f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_546 N_A_548_87#_c_585_n N_A_1979_71#_c_1537_n 0.00395024f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_547 N_A_548_87#_c_585_n N_A_1979_71#_c_1538_n 0.00488722f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_548 N_A_548_87#_c_585_n N_A_1736_97#_c_1632_n 0.0033031f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_549 N_A_548_87#_c_585_n N_A_1736_97#_c_1634_n 0.0126985f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_550 N_A_548_87#_c_585_n N_A_1736_97#_c_1636_n 0.0542375f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_551 N_A_548_87#_c_585_n N_A_1736_97#_c_1637_n 0.0125798f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_552 N_A_548_87#_c_585_n N_A_1736_97#_c_1639_n 0.00120832f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_553 N_A_548_87#_c_585_n N_A_1736_97#_c_1640_n 0.0253166f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_554 N_A_548_87#_c_579_n N_A_2474_74#_M1023_g 0.00999105f $X=13.69 $Y=0.94
+ $X2=0 $Y2=0
cc_555 N_A_548_87#_c_582_n N_A_2474_74#_M1023_g 0.0236141f $X=14.48 $Y=0.58
+ $X2=0 $Y2=0
cc_556 N_A_548_87#_c_583_n N_A_2474_74#_M1023_g 0.00219123f $X=14.665 $Y=1.55
+ $X2=0 $Y2=0
cc_557 N_A_548_87#_c_584_n N_A_2474_74#_M1023_g 0.00703637f $X=14.532 $Y=1.29
+ $X2=0 $Y2=0
cc_558 N_A_548_87#_c_592_n N_A_2474_74#_c_1729_n 0.0152899f $X=13.63 $Y=2.465
+ $X2=0 $Y2=0
cc_559 N_A_548_87#_c_594_n N_A_2474_74#_c_1729_n 0.00978681f $X=14.4 $Y=2.385
+ $X2=0 $Y2=0
cc_560 N_A_548_87#_c_595_n N_A_2474_74#_c_1729_n 0.0018588f $X=14.665 $Y=2.3
+ $X2=0 $Y2=0
cc_561 N_A_548_87#_c_596_n N_A_2474_74#_c_1729_n 4.3236e-19 $X=13.675 $Y=2.215
+ $X2=0 $Y2=0
cc_562 N_A_548_87#_c_597_n N_A_2474_74#_c_1729_n 0.00856906f $X=14.565 $Y=2.465
+ $X2=0 $Y2=0
cc_563 N_A_548_87#_c_583_n N_A_2474_74#_c_1718_n 0.0202084f $X=14.665 $Y=1.55
+ $X2=0 $Y2=0
cc_564 N_A_548_87#_c_584_n N_A_2474_74#_c_1718_n 0.0072045f $X=14.532 $Y=1.29
+ $X2=0 $Y2=0
cc_565 N_A_548_87#_c_597_n N_A_2474_74#_c_1718_n 0.00295373f $X=14.565 $Y=2.465
+ $X2=0 $Y2=0
cc_566 N_A_548_87#_c_598_n N_A_2474_74#_c_1718_n 0.00586175f $X=14.665 $Y=1.665
+ $X2=0 $Y2=0
cc_567 N_A_548_87#_c_585_n N_A_2474_74#_c_1718_n 0.00289525f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_568 N_A_548_87#_c_601_n N_A_2474_74#_c_1718_n 0.00525975f $X=15.12 $Y=1.665
+ $X2=0 $Y2=0
cc_569 N_A_548_87#_c_587_n N_A_2474_74#_c_1718_n 0.022941f $X=15.12 $Y=1.665
+ $X2=0 $Y2=0
cc_570 N_A_548_87#_c_582_n N_A_2474_74#_M1008_g 0.00493039f $X=14.48 $Y=0.58
+ $X2=0 $Y2=0
cc_571 N_A_548_87#_c_584_n N_A_2474_74#_M1008_g 0.00618705f $X=14.532 $Y=1.29
+ $X2=0 $Y2=0
cc_572 N_A_548_87#_c_595_n N_A_2474_74#_c_1730_n 0.00272083f $X=14.665 $Y=2.3
+ $X2=0 $Y2=0
cc_573 N_A_548_87#_c_597_n N_A_2474_74#_c_1730_n 8.92646e-19 $X=14.565 $Y=2.465
+ $X2=0 $Y2=0
cc_574 N_A_548_87#_c_601_n N_A_2474_74#_c_1730_n 3.812e-19 $X=15.12 $Y=1.665
+ $X2=0 $Y2=0
cc_575 N_A_548_87#_c_587_n N_A_2474_74#_c_1730_n 3.05685e-19 $X=15.12 $Y=1.665
+ $X2=0 $Y2=0
cc_576 N_A_548_87#_c_581_n N_A_2474_74#_c_1721_n 0.0286462f $X=13.765 $Y=2.05
+ $X2=0 $Y2=0
cc_577 N_A_548_87#_c_585_n N_A_2474_74#_c_1721_n 3.04627e-19 $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_578 N_A_548_87#_c_592_n N_A_2474_74#_c_1732_n 0.00374141f $X=13.63 $Y=2.465
+ $X2=0 $Y2=0
cc_579 N_A_548_87#_c_594_n N_A_2474_74#_c_1732_n 0.00162878f $X=14.4 $Y=2.385
+ $X2=0 $Y2=0
cc_580 N_A_548_87#_c_596_n N_A_2474_74#_c_1732_n 8.00821e-19 $X=13.675 $Y=2.215
+ $X2=0 $Y2=0
cc_581 N_A_548_87#_c_597_n N_A_2474_74#_c_1732_n 8.17456e-19 $X=14.565 $Y=2.465
+ $X2=0 $Y2=0
cc_582 N_A_548_87#_c_601_n N_A_2474_74#_c_1722_n 0.00515183f $X=15.12 $Y=1.665
+ $X2=0 $Y2=0
cc_583 N_A_548_87#_c_587_n N_A_2474_74#_c_1722_n 0.00336166f $X=15.12 $Y=1.665
+ $X2=0 $Y2=0
cc_584 N_A_548_87#_c_578_n N_A_2474_74#_c_1723_n 0.00177547f $X=13.16 $Y=0.865
+ $X2=0 $Y2=0
cc_585 N_A_548_87#_c_578_n N_A_2474_74#_c_1724_n 0.00387158f $X=13.16 $Y=0.865
+ $X2=0 $Y2=0
cc_586 N_A_548_87#_c_579_n N_A_2474_74#_c_1724_n 0.0220102f $X=13.69 $Y=0.94
+ $X2=0 $Y2=0
cc_587 N_A_548_87#_c_580_n N_A_2474_74#_c_1724_n 0.00439386f $X=13.235 $Y=0.94
+ $X2=0 $Y2=0
cc_588 N_A_548_87#_c_582_n N_A_2474_74#_c_1724_n 0.00542813f $X=14.48 $Y=0.58
+ $X2=0 $Y2=0
cc_589 N_A_548_87#_c_585_n N_A_2474_74#_c_1724_n 0.00608858f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_590 N_A_548_87#_c_592_n N_A_2474_74#_c_1734_n 0.00317561f $X=13.63 $Y=2.465
+ $X2=0 $Y2=0
cc_591 N_A_548_87#_c_596_n N_A_2474_74#_c_1734_n 0.0201628f $X=13.675 $Y=2.215
+ $X2=0 $Y2=0
cc_592 N_A_548_87#_c_592_n N_A_2474_74#_c_1735_n 0.00289846f $X=13.63 $Y=2.465
+ $X2=0 $Y2=0
cc_593 N_A_548_87#_c_596_n N_A_2474_74#_c_1735_n 0.00780014f $X=13.675 $Y=2.215
+ $X2=0 $Y2=0
cc_594 N_A_548_87#_c_585_n N_A_2474_74#_c_1735_n 0.0147772f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_595 N_A_548_87#_c_592_n N_A_2474_74#_c_1736_n 3.01282e-19 $X=13.63 $Y=2.465
+ $X2=0 $Y2=0
cc_596 N_A_548_87#_c_581_n N_A_2474_74#_c_1736_n 6.57788e-19 $X=13.765 $Y=2.05
+ $X2=0 $Y2=0
cc_597 N_A_548_87#_c_596_n N_A_2474_74#_c_1736_n 2.69369e-19 $X=13.675 $Y=2.215
+ $X2=0 $Y2=0
cc_598 N_A_548_87#_c_585_n N_A_2474_74#_c_1736_n 0.0105856f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_599 N_A_548_87#_c_581_n N_A_2474_74#_c_1726_n 0.0210794f $X=13.765 $Y=2.05
+ $X2=0 $Y2=0
cc_600 N_A_548_87#_c_582_n N_A_2474_74#_c_1726_n 0.00774336f $X=14.48 $Y=0.58
+ $X2=0 $Y2=0
cc_601 N_A_548_87#_c_585_n N_A_2474_74#_c_1726_n 0.0191547f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_602 N_A_548_87#_c_581_n N_A_2474_74#_c_1738_n 0.00383999f $X=13.765 $Y=2.05
+ $X2=0 $Y2=0
cc_603 N_A_548_87#_c_594_n N_A_2474_74#_c_1738_n 0.00906073f $X=14.4 $Y=2.385
+ $X2=0 $Y2=0
cc_604 N_A_548_87#_c_596_n N_A_2474_74#_c_1738_n 0.00330635f $X=13.675 $Y=2.215
+ $X2=0 $Y2=0
cc_605 N_A_548_87#_c_585_n N_A_2474_74#_c_1738_n 0.0149659f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_606 N_A_548_87#_c_592_n N_A_2474_74#_c_1739_n 0.00200719f $X=13.63 $Y=2.465
+ $X2=0 $Y2=0
cc_607 N_A_548_87#_c_581_n N_A_2474_74#_c_1739_n 0.00560273f $X=13.765 $Y=2.05
+ $X2=0 $Y2=0
cc_608 N_A_548_87#_c_596_n N_A_2474_74#_c_1739_n 0.013301f $X=13.675 $Y=2.215
+ $X2=0 $Y2=0
cc_609 N_A_548_87#_c_581_n N_A_2474_74#_c_1727_n 0.00238202f $X=13.765 $Y=2.05
+ $X2=0 $Y2=0
cc_610 N_A_548_87#_c_594_n N_A_2474_74#_c_1727_n 0.024293f $X=14.4 $Y=2.385
+ $X2=0 $Y2=0
cc_611 N_A_548_87#_c_583_n N_A_2474_74#_c_1727_n 0.00639324f $X=14.665 $Y=1.55
+ $X2=0 $Y2=0
cc_612 N_A_548_87#_c_595_n N_A_2474_74#_c_1727_n 0.026229f $X=14.665 $Y=2.3
+ $X2=0 $Y2=0
cc_613 N_A_548_87#_c_596_n N_A_2474_74#_c_1727_n 0.00199397f $X=13.675 $Y=2.215
+ $X2=0 $Y2=0
cc_614 N_A_548_87#_c_584_n N_A_2474_74#_c_1727_n 0.00761289f $X=14.532 $Y=1.29
+ $X2=0 $Y2=0
cc_615 N_A_548_87#_c_597_n N_A_2474_74#_c_1727_n 7.40414e-19 $X=14.565 $Y=2.465
+ $X2=0 $Y2=0
cc_616 N_A_548_87#_c_598_n N_A_2474_74#_c_1727_n 0.0169075f $X=14.665 $Y=1.665
+ $X2=0 $Y2=0
cc_617 N_A_548_87#_c_585_n N_A_2474_74#_c_1727_n 0.0263253f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_618 N_A_548_87#_c_601_n N_A_2474_74#_c_1727_n 2.89456e-19 $X=15.12 $Y=1.665
+ $X2=0 $Y2=0
cc_619 N_A_548_87#_c_592_n N_A_2474_74#_c_1728_n 0.0186552f $X=13.63 $Y=2.465
+ $X2=0 $Y2=0
cc_620 N_A_548_87#_c_595_n N_A_2474_74#_c_1728_n 0.0122157f $X=14.665 $Y=2.3
+ $X2=0 $Y2=0
cc_621 N_A_548_87#_c_598_n N_A_2474_74#_c_1728_n 0.00327333f $X=14.665 $Y=1.665
+ $X2=0 $Y2=0
cc_622 N_A_548_87#_c_585_n N_A_2474_74#_c_1728_n 0.0030092f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_623 N_A_548_87#_c_591_n N_A_40_464#_c_1897_n 0.0133663f $X=3.19 $Y=2.24 $X2=0
+ $Y2=0
cc_624 N_A_548_87#_c_585_n N_A_40_464#_c_1897_n 0.00615181f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_625 N_A_548_87#_c_586_n N_A_40_464#_c_1897_n 0.00338869f $X=2.785 $Y=1.665
+ $X2=0 $Y2=0
cc_626 N_A_548_87#_c_588_n N_A_40_464#_c_1897_n 0.015783f $X=2.905 $Y=1.68 $X2=0
+ $Y2=0
cc_627 N_A_548_87#_c_589_n N_A_40_464#_c_1897_n 0.00459904f $X=3.19 $Y=1.68
+ $X2=0 $Y2=0
cc_628 N_A_548_87#_M1025_g N_A_40_464#_c_1886_n 0.00328556f $X=2.815 $Y=0.775
+ $X2=0 $Y2=0
cc_629 N_A_548_87#_c_591_n N_A_40_464#_c_1899_n 0.00870642f $X=3.19 $Y=2.24
+ $X2=0 $Y2=0
cc_630 N_A_548_87#_M1025_g N_A_40_464#_c_1887_n 0.00436523f $X=2.815 $Y=0.775
+ $X2=0 $Y2=0
cc_631 N_A_548_87#_c_591_n N_A_40_464#_c_1887_n 0.00116727f $X=3.19 $Y=2.24
+ $X2=0 $Y2=0
cc_632 N_A_548_87#_c_585_n N_A_40_464#_c_1887_n 0.0171118f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_633 N_A_548_87#_c_586_n N_A_40_464#_c_1887_n 3.84274e-19 $X=2.785 $Y=1.665
+ $X2=0 $Y2=0
cc_634 N_A_548_87#_c_588_n N_A_40_464#_c_1887_n 0.0163955f $X=2.905 $Y=1.68
+ $X2=0 $Y2=0
cc_635 N_A_548_87#_c_589_n N_A_40_464#_c_1887_n 0.0185455f $X=3.19 $Y=1.68 $X2=0
+ $Y2=0
cc_636 N_A_548_87#_M1025_g N_A_40_464#_c_1889_n 0.0118478f $X=2.815 $Y=0.775
+ $X2=0 $Y2=0
cc_637 N_A_548_87#_c_585_n N_A_40_464#_c_1889_n 0.00423042f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_638 N_A_548_87#_c_588_n N_A_40_464#_c_1889_n 0.00559384f $X=2.905 $Y=1.68
+ $X2=0 $Y2=0
cc_639 N_A_548_87#_c_589_n N_A_40_464#_c_1889_n 0.00624078f $X=3.19 $Y=1.68
+ $X2=0 $Y2=0
cc_640 N_A_548_87#_M1025_g N_A_40_464#_c_1890_n 0.00517201f $X=2.815 $Y=0.775
+ $X2=0 $Y2=0
cc_641 N_A_548_87#_c_585_n N_A_40_464#_c_1890_n 0.00699364f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_642 N_A_548_87#_c_589_n N_A_40_464#_c_1890_n 0.00456568f $X=3.19 $Y=1.68
+ $X2=0 $Y2=0
cc_643 N_A_548_87#_c_591_n N_A_40_464#_c_1902_n 0.00166465f $X=3.19 $Y=2.24
+ $X2=0 $Y2=0
cc_644 N_A_548_87#_c_585_n N_A_40_464#_c_1902_n 0.00276825f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_645 N_A_548_87#_c_594_n N_VPWR_M1037_d 0.00278057f $X=14.4 $Y=2.385 $X2=0
+ $Y2=0
cc_646 N_A_548_87#_c_591_n N_VPWR_c_2015_n 0.00150486f $X=3.19 $Y=2.24 $X2=0
+ $Y2=0
cc_647 N_A_548_87#_c_592_n N_VPWR_c_2021_n 0.0161132f $X=13.63 $Y=2.465 $X2=0
+ $Y2=0
cc_648 N_A_548_87#_c_594_n N_VPWR_c_2021_n 0.0282015f $X=14.4 $Y=2.385 $X2=0
+ $Y2=0
cc_649 N_A_548_87#_c_596_n N_VPWR_c_2021_n 0.00959871f $X=13.675 $Y=2.215 $X2=0
+ $Y2=0
cc_650 N_A_548_87#_c_597_n N_VPWR_c_2021_n 0.013346f $X=14.565 $Y=2.465 $X2=0
+ $Y2=0
cc_651 N_A_548_87#_c_595_n N_VPWR_c_2022_n 0.0238978f $X=14.665 $Y=2.3 $X2=0
+ $Y2=0
cc_652 N_A_548_87#_c_597_n N_VPWR_c_2022_n 0.0497073f $X=14.565 $Y=2.465 $X2=0
+ $Y2=0
cc_653 N_A_548_87#_c_601_n N_VPWR_c_2022_n 0.00903602f $X=15.12 $Y=1.665 $X2=0
+ $Y2=0
cc_654 N_A_548_87#_c_587_n N_VPWR_c_2022_n 0.0192745f $X=15.12 $Y=1.665 $X2=0
+ $Y2=0
cc_655 N_A_548_87#_c_592_n N_VPWR_c_2027_n 0.00413917f $X=13.63 $Y=2.465 $X2=0
+ $Y2=0
cc_656 N_A_548_87#_c_591_n N_VPWR_c_2031_n 0.0044174f $X=3.19 $Y=2.24 $X2=0
+ $Y2=0
cc_657 N_A_548_87#_c_597_n N_VPWR_c_2035_n 0.0154862f $X=14.565 $Y=2.465 $X2=0
+ $Y2=0
cc_658 N_A_548_87#_c_591_n N_VPWR_c_2013_n 0.00544287f $X=3.19 $Y=2.24 $X2=0
+ $Y2=0
cc_659 N_A_548_87#_c_592_n N_VPWR_c_2013_n 0.00418596f $X=13.63 $Y=2.465 $X2=0
+ $Y2=0
cc_660 N_A_548_87#_c_594_n N_VPWR_c_2013_n 0.00607335f $X=14.4 $Y=2.385 $X2=0
+ $Y2=0
cc_661 N_A_548_87#_c_596_n N_VPWR_c_2013_n 0.00607203f $X=13.675 $Y=2.215 $X2=0
+ $Y2=0
cc_662 N_A_548_87#_c_597_n N_VPWR_c_2013_n 0.0127853f $X=14.565 $Y=2.465 $X2=0
+ $Y2=0
cc_663 N_A_548_87#_c_585_n N_A_693_113#_c_2204_n 0.00396843f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_664 N_A_548_87#_c_591_n N_A_693_113#_c_2216_n 5.18926e-19 $X=3.19 $Y=2.24
+ $X2=0 $Y2=0
cc_665 N_A_548_87#_c_585_n N_A_693_113#_c_2206_n 0.00719012f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_666 N_A_548_87#_c_585_n N_A_693_113#_c_2209_n 0.0135215f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_667 N_A_548_87#_c_585_n N_A_693_113#_c_2197_n 0.0284899f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_668 N_A_548_87#_c_585_n N_A_693_113#_c_2198_n 0.00557586f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_669 N_A_548_87#_c_585_n N_A_693_113#_c_2200_n 0.00539994f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_670 N_A_548_87#_c_585_n N_A_693_113#_c_2201_n 0.0179309f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_671 N_A_548_87#_c_585_n N_A_693_113#_c_2202_n 0.0069318f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_672 N_A_548_87#_c_585_n N_A_693_113#_c_2203_n 0.0256048f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_673 N_A_548_87#_c_584_n N_Q_c_2375_n 3.0226e-19 $X=14.532 $Y=1.29 $X2=0 $Y2=0
cc_674 N_A_548_87#_c_601_n Q 0.00658326f $X=15.12 $Y=1.665 $X2=0 $Y2=0
cc_675 N_A_548_87#_c_587_n Q 0.0123872f $X=15.12 $Y=1.665 $X2=0 $Y2=0
cc_676 N_A_548_87#_M1025_g N_VGND_c_2407_n 0.00212753f $X=2.815 $Y=0.775 $X2=0
+ $Y2=0
cc_677 N_A_548_87#_c_585_n N_VGND_c_2408_n 0.00348115f $X=14.975 $Y=1.665 $X2=0
+ $Y2=0
cc_678 N_A_548_87#_c_585_n N_VGND_c_2410_n 0.00182967f $X=14.975 $Y=1.665 $X2=0
+ $Y2=0
cc_679 N_A_548_87#_c_582_n N_VGND_c_2413_n 0.0404514f $X=14.48 $Y=0.58 $X2=0
+ $Y2=0
cc_680 N_A_548_87#_c_601_n N_VGND_c_2413_n 0.00427042f $X=15.12 $Y=1.665 $X2=0
+ $Y2=0
cc_681 N_A_548_87#_c_587_n N_VGND_c_2413_n 0.00642692f $X=15.12 $Y=1.665 $X2=0
+ $Y2=0
cc_682 N_A_548_87#_M1025_g N_VGND_c_2420_n 0.00431664f $X=2.815 $Y=0.775 $X2=0
+ $Y2=0
cc_683 N_A_548_87#_c_582_n N_VGND_c_2424_n 0.0145639f $X=14.48 $Y=0.58 $X2=0
+ $Y2=0
cc_684 N_A_548_87#_c_578_n N_VGND_c_2432_n 0.00383152f $X=13.16 $Y=0.865 $X2=0
+ $Y2=0
cc_685 N_A_548_87#_c_578_n N_VGND_c_2433_n 0.0115585f $X=13.16 $Y=0.865 $X2=0
+ $Y2=0
cc_686 N_A_548_87#_c_579_n N_VGND_c_2433_n 0.00645873f $X=13.69 $Y=0.94 $X2=0
+ $Y2=0
cc_687 N_A_548_87#_c_582_n N_VGND_c_2433_n 0.0132893f $X=14.48 $Y=0.58 $X2=0
+ $Y2=0
cc_688 N_A_548_87#_M1025_g N_VGND_c_2435_n 0.00486331f $X=2.815 $Y=0.775 $X2=0
+ $Y2=0
cc_689 N_A_548_87#_c_578_n N_VGND_c_2435_n 0.00384101f $X=13.16 $Y=0.865 $X2=0
+ $Y2=0
cc_690 N_A_548_87#_c_582_n N_VGND_c_2435_n 0.0119984f $X=14.48 $Y=0.58 $X2=0
+ $Y2=0
cc_691 N_A_663_87#_c_840_n N_SCD_c_942_n 0.0283165f $X=5.785 $Y=1.92 $X2=0 $Y2=0
cc_692 N_A_663_87#_c_843_n N_SCD_c_942_n 0.01197f $X=5.62 $Y=2 $X2=0 $Y2=0
cc_693 N_A_663_87#_c_839_n N_SCD_c_943_n 0.0385396f $X=5.74 $Y=2.2 $X2=0 $Y2=0
cc_694 N_A_663_87#_c_849_n SCD 0.00443615f $X=4.13 $Y=1.78 $X2=0 $Y2=0
cc_695 N_A_663_87#_c_843_n SCD 0.0325296f $X=5.62 $Y=2 $X2=0 $Y2=0
cc_696 N_A_663_87#_c_836_n SCD 0.0193736f $X=5.785 $Y=1.58 $X2=0 $Y2=0
cc_697 N_A_663_87#_c_837_n SCD 0.00113825f $X=5.785 $Y=1.58 $X2=0 $Y2=0
cc_698 N_A_663_87#_c_843_n N_SCD_c_941_n 0.00105366f $X=5.62 $Y=2 $X2=0 $Y2=0
cc_699 N_A_663_87#_c_836_n N_SCD_c_941_n 0.00227865f $X=5.785 $Y=1.58 $X2=0
+ $Y2=0
cc_700 N_A_663_87#_c_837_n N_SCD_c_941_n 0.0217422f $X=5.785 $Y=1.58 $X2=0 $Y2=0
cc_701 N_A_663_87#_c_842_n N_SCE_c_989_n 3.49329e-19 $X=4.21 $Y=2.255 $X2=-0.19
+ $Y2=-0.245
cc_702 N_A_663_87#_c_846_n N_SCE_c_989_n 0.00103127f $X=4.415 $Y=2.495 $X2=-0.19
+ $Y2=-0.245
cc_703 N_A_663_87#_c_846_n N_SCE_c_990_n 0.00213313f $X=4.415 $Y=2.495 $X2=0
+ $Y2=0
cc_704 N_A_663_87#_c_849_n N_SCE_c_982_n 0.00221467f $X=4.13 $Y=1.78 $X2=0 $Y2=0
cc_705 N_A_663_87#_c_835_n N_SCE_c_982_n 0.0232065f $X=4.13 $Y=1.78 $X2=0 $Y2=0
cc_706 N_A_663_87#_c_842_n N_SCE_c_982_n 0.00363753f $X=4.21 $Y=2.255 $X2=0
+ $Y2=0
cc_707 N_A_663_87#_c_843_n N_SCE_c_982_n 0.0189248f $X=5.62 $Y=2 $X2=0 $Y2=0
cc_708 N_A_663_87#_c_842_n N_SCE_M1003_g 0.00167654f $X=4.21 $Y=2.255 $X2=0
+ $Y2=0
cc_709 N_A_663_87#_c_846_n N_SCE_M1003_g 0.00322271f $X=4.415 $Y=2.495 $X2=0
+ $Y2=0
cc_710 N_A_663_87#_c_833_n N_SCE_M1031_g 0.00135337f $X=4.13 $Y=0.42 $X2=0 $Y2=0
cc_711 N_A_663_87#_c_834_n N_SCE_M1031_g 0.0220325f $X=4.13 $Y=0.42 $X2=0 $Y2=0
cc_712 N_A_663_87#_c_849_n N_SCE_M1031_g 9.75671e-19 $X=4.13 $Y=1.78 $X2=0 $Y2=0
cc_713 N_A_663_87#_c_838_n N_SCE_M1031_g 0.00545163f $X=4.55 $Y=0.805 $X2=0
+ $Y2=0
cc_714 N_A_663_87#_c_836_n N_SCE_M1004_g 5.1902e-19 $X=5.785 $Y=1.58 $X2=0 $Y2=0
cc_715 N_A_663_87#_c_837_n N_SCE_M1004_g 0.00456126f $X=5.785 $Y=1.58 $X2=0
+ $Y2=0
cc_716 N_A_663_87#_c_832_n N_SCE_c_987_n 0.0207308f $X=4.13 $Y=1.135 $X2=0 $Y2=0
cc_717 N_A_663_87#_c_849_n N_SCE_c_987_n 3.77471e-19 $X=4.13 $Y=1.78 $X2=0 $Y2=0
cc_718 N_A_663_87#_c_843_n N_SCE_c_987_n 0.00383649f $X=5.62 $Y=2 $X2=0 $Y2=0
cc_719 N_A_663_87#_c_838_n N_SCE_c_987_n 0.00463638f $X=4.55 $Y=0.805 $X2=0
+ $Y2=0
cc_720 N_A_663_87#_c_832_n N_SCE_c_988_n 0.00185703f $X=4.13 $Y=1.135 $X2=0
+ $Y2=0
cc_721 N_A_663_87#_c_849_n N_SCE_c_988_n 0.025711f $X=4.13 $Y=1.78 $X2=0 $Y2=0
cc_722 N_A_663_87#_c_843_n N_SCE_c_988_n 0.00594157f $X=5.62 $Y=2 $X2=0 $Y2=0
cc_723 N_A_663_87#_c_838_n N_SCE_c_988_n 0.0170506f $X=4.55 $Y=0.805 $X2=0 $Y2=0
cc_724 N_A_663_87#_c_837_n N_CLK_c_1068_n 0.00535178f $X=5.785 $Y=1.58 $X2=0
+ $Y2=0
cc_725 N_A_663_87#_c_829_n N_A_40_464#_c_1886_n 0.00146461f $X=3.39 $Y=1.06
+ $X2=0 $Y2=0
cc_726 N_A_663_87#_c_831_n N_A_40_464#_c_1886_n 0.00376733f $X=3.465 $Y=1.135
+ $X2=0 $Y2=0
cc_727 N_A_663_87#_c_831_n N_A_40_464#_c_1887_n 9.15581e-19 $X=3.465 $Y=1.135
+ $X2=0 $Y2=0
cc_728 N_A_663_87#_c_829_n N_A_40_464#_c_1889_n 0.00925923f $X=3.39 $Y=1.06
+ $X2=0 $Y2=0
cc_729 N_A_663_87#_c_830_n N_A_40_464#_c_1890_n 0.00265188f $X=3.965 $Y=1.135
+ $X2=0 $Y2=0
cc_730 N_A_663_87#_c_831_n N_A_40_464#_c_1890_n 0.00898456f $X=3.465 $Y=1.135
+ $X2=0 $Y2=0
cc_731 N_A_663_87#_c_839_n N_VPWR_c_2016_n 0.00151367f $X=5.74 $Y=2.2 $X2=0
+ $Y2=0
cc_732 N_A_663_87#_c_839_n N_VPWR_c_2017_n 0.00319238f $X=5.74 $Y=2.2 $X2=0
+ $Y2=0
cc_733 N_A_663_87#_c_839_n N_VPWR_c_2032_n 0.00530811f $X=5.74 $Y=2.2 $X2=0
+ $Y2=0
cc_734 N_A_663_87#_c_839_n N_VPWR_c_2013_n 0.005315f $X=5.74 $Y=2.2 $X2=0 $Y2=0
cc_735 N_A_663_87#_c_846_n N_A_693_113#_c_2204_n 0.035221f $X=4.415 $Y=2.495
+ $X2=0 $Y2=0
cc_736 N_A_663_87#_M1003_s N_A_693_113#_c_2205_n 0.00270287f $X=4.275 $Y=2.275
+ $X2=0 $Y2=0
cc_737 N_A_663_87#_c_846_n N_A_693_113#_c_2205_n 0.0280635f $X=4.415 $Y=2.495
+ $X2=0 $Y2=0
cc_738 N_A_663_87#_c_846_n N_A_693_113#_c_2228_n 0.0231836f $X=4.415 $Y=2.495
+ $X2=0 $Y2=0
cc_739 N_A_663_87#_c_839_n N_A_693_113#_c_2206_n 0.0155481f $X=5.74 $Y=2.2 $X2=0
+ $Y2=0
cc_740 N_A_663_87#_c_840_n N_A_693_113#_c_2206_n 0.00465705f $X=5.785 $Y=1.92
+ $X2=0 $Y2=0
cc_741 N_A_663_87#_c_843_n N_A_693_113#_c_2206_n 0.0761498f $X=5.62 $Y=2 $X2=0
+ $Y2=0
cc_742 N_A_663_87#_c_843_n N_A_693_113#_c_2207_n 0.0134263f $X=5.62 $Y=2 $X2=0
+ $Y2=0
cc_743 N_A_663_87#_c_846_n N_A_693_113#_c_2207_n 0.0141567f $X=4.415 $Y=2.495
+ $X2=0 $Y2=0
cc_744 N_A_663_87#_c_829_n N_A_693_113#_c_2200_n 0.00373895f $X=3.39 $Y=1.06
+ $X2=0 $Y2=0
cc_745 N_A_663_87#_c_830_n N_A_693_113#_c_2200_n 0.00505284f $X=3.965 $Y=1.135
+ $X2=0 $Y2=0
cc_746 N_A_663_87#_c_833_n N_A_693_113#_c_2200_n 0.00469807f $X=4.13 $Y=0.42
+ $X2=0 $Y2=0
cc_747 N_A_663_87#_c_834_n N_A_693_113#_c_2200_n 0.00512646f $X=4.13 $Y=0.42
+ $X2=0 $Y2=0
cc_748 N_A_663_87#_c_838_n N_A_693_113#_c_2200_n 0.0338556f $X=4.55 $Y=0.805
+ $X2=0 $Y2=0
cc_749 N_A_663_87#_c_829_n N_A_693_113#_c_2201_n 4.79113e-19 $X=3.39 $Y=1.06
+ $X2=0 $Y2=0
cc_750 N_A_663_87#_c_830_n N_A_693_113#_c_2201_n 0.0149913f $X=3.965 $Y=1.135
+ $X2=0 $Y2=0
cc_751 N_A_663_87#_c_849_n N_A_693_113#_c_2201_n 0.0656831f $X=4.13 $Y=1.78
+ $X2=0 $Y2=0
cc_752 N_A_663_87#_c_835_n N_A_693_113#_c_2201_n 0.0117795f $X=4.13 $Y=1.78
+ $X2=0 $Y2=0
cc_753 N_A_663_87#_c_842_n N_A_693_113#_c_2201_n 0.00891632f $X=4.21 $Y=2.255
+ $X2=0 $Y2=0
cc_754 N_A_663_87#_c_845_n N_A_693_113#_c_2201_n 0.0142218f $X=4.152 $Y=2 $X2=0
+ $Y2=0
cc_755 N_A_663_87#_c_846_n N_A_693_113#_c_2201_n 0.00216189f $X=4.415 $Y=2.495
+ $X2=0 $Y2=0
cc_756 N_A_663_87#_c_836_n N_A_693_113#_c_2202_n 0.00897337f $X=5.785 $Y=1.58
+ $X2=0 $Y2=0
cc_757 N_A_663_87#_c_837_n N_A_693_113#_c_2202_n 0.00375671f $X=5.785 $Y=1.58
+ $X2=0 $Y2=0
cc_758 N_A_663_87#_c_840_n N_A_693_113#_c_2203_n 0.00378886f $X=5.785 $Y=1.92
+ $X2=0 $Y2=0
cc_759 N_A_663_87#_c_843_n N_A_693_113#_c_2203_n 0.0135425f $X=5.62 $Y=2 $X2=0
+ $Y2=0
cc_760 N_A_663_87#_c_836_n N_A_693_113#_c_2203_n 0.0360687f $X=5.785 $Y=1.58
+ $X2=0 $Y2=0
cc_761 N_A_663_87#_c_837_n N_A_693_113#_c_2203_n 0.0114743f $X=5.785 $Y=1.58
+ $X2=0 $Y2=0
cc_762 N_A_663_87#_c_839_n N_A_693_113#_c_2214_n 0.00721931f $X=5.74 $Y=2.2
+ $X2=0 $Y2=0
cc_763 N_A_663_87#_c_833_n N_VGND_c_2408_n 0.0106324f $X=4.13 $Y=0.42 $X2=0
+ $Y2=0
cc_764 N_A_663_87#_c_838_n N_VGND_c_2408_n 0.0178216f $X=4.55 $Y=0.805 $X2=0
+ $Y2=0
cc_765 N_A_663_87#_c_829_n N_VGND_c_2420_n 0.00431664f $X=3.39 $Y=1.06 $X2=0
+ $Y2=0
cc_766 N_A_663_87#_c_833_n N_VGND_c_2420_n 0.0184034f $X=4.13 $Y=0.42 $X2=0
+ $Y2=0
cc_767 N_A_663_87#_c_834_n N_VGND_c_2420_n 0.00356704f $X=4.13 $Y=0.42 $X2=0
+ $Y2=0
cc_768 N_A_663_87#_c_838_n N_VGND_c_2420_n 0.00867058f $X=4.55 $Y=0.805 $X2=0
+ $Y2=0
cc_769 N_A_663_87#_c_829_n N_VGND_c_2435_n 0.00486331f $X=3.39 $Y=1.06 $X2=0
+ $Y2=0
cc_770 N_A_663_87#_c_833_n N_VGND_c_2435_n 0.0106565f $X=4.13 $Y=0.42 $X2=0
+ $Y2=0
cc_771 N_A_663_87#_c_834_n N_VGND_c_2435_n 0.00169532f $X=4.13 $Y=0.42 $X2=0
+ $Y2=0
cc_772 N_A_663_87#_c_838_n N_VGND_c_2435_n 0.0126496f $X=4.55 $Y=0.805 $X2=0
+ $Y2=0
cc_773 N_SCD_c_943_n N_SCE_c_990_n 0.00100522f $X=5.32 $Y=2.2 $X2=0 $Y2=0
cc_774 N_SCD_c_942_n N_SCE_c_982_n 0.00601231f $X=5.32 $Y=2.11 $X2=0 $Y2=0
cc_775 SCD N_SCE_c_982_n 0.00228345f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_776 N_SCD_c_941_n N_SCE_c_982_n 0.00803162f $X=5.245 $Y=1.58 $X2=0 $Y2=0
cc_777 N_SCD_c_943_n N_SCE_c_993_n 0.00601231f $X=5.32 $Y=2.2 $X2=0 $Y2=0
cc_778 N_SCD_c_943_n N_SCE_M1003_g 0.0111767f $X=5.32 $Y=2.2 $X2=0 $Y2=0
cc_779 N_SCD_M1041_g N_SCE_M1031_g 0.0231737f $X=5.265 $Y=0.835 $X2=0 $Y2=0
cc_780 N_SCD_M1041_g N_SCE_c_984_n 0.00894529f $X=5.265 $Y=0.835 $X2=0 $Y2=0
cc_781 N_SCD_M1041_g N_SCE_M1004_g 0.040291f $X=5.265 $Y=0.835 $X2=0 $Y2=0
cc_782 SCD N_SCE_c_987_n 0.0026706f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_783 N_SCD_c_941_n N_SCE_c_987_n 0.00496971f $X=5.245 $Y=1.58 $X2=0 $Y2=0
cc_784 SCD N_SCE_c_988_n 0.0267067f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_785 N_SCD_c_943_n N_VPWR_c_2016_n 0.00985948f $X=5.32 $Y=2.2 $X2=0 $Y2=0
cc_786 N_SCD_c_943_n N_VPWR_c_2032_n 0.00489294f $X=5.32 $Y=2.2 $X2=0 $Y2=0
cc_787 N_SCD_c_943_n N_VPWR_c_2013_n 0.00481893f $X=5.32 $Y=2.2 $X2=0 $Y2=0
cc_788 N_SCD_c_943_n N_A_693_113#_c_2205_n 3.76568e-19 $X=5.32 $Y=2.2 $X2=0
+ $Y2=0
cc_789 N_SCD_c_943_n N_A_693_113#_c_2228_n 0.00283455f $X=5.32 $Y=2.2 $X2=0
+ $Y2=0
cc_790 N_SCD_c_943_n N_A_693_113#_c_2206_n 0.0181248f $X=5.32 $Y=2.2 $X2=0 $Y2=0
cc_791 N_SCD_M1041_g N_A_693_113#_c_2202_n 0.00137701f $X=5.265 $Y=0.835 $X2=0
+ $Y2=0
cc_792 SCD N_A_693_113#_c_2203_n 0.00754501f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_793 N_SCD_M1041_g N_VGND_c_2408_n 0.010608f $X=5.265 $Y=0.835 $X2=0 $Y2=0
cc_794 SCD N_VGND_c_2408_n 0.0201937f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_795 N_SCD_c_941_n N_VGND_c_2408_n 4.02357e-19 $X=5.245 $Y=1.58 $X2=0 $Y2=0
cc_796 N_SCD_M1041_g N_VGND_c_2435_n 7.97988e-19 $X=5.265 $Y=0.835 $X2=0 $Y2=0
cc_797 N_SCE_c_989_n N_A_40_464#_c_1899_n 0.00161473f $X=3.64 $Y=3.03 $X2=0
+ $Y2=0
cc_798 N_SCE_c_989_n N_A_40_464#_c_1887_n 7.32247e-19 $X=3.64 $Y=3.03 $X2=0
+ $Y2=0
cc_799 N_SCE_c_989_n N_A_40_464#_c_1902_n 7.52181e-19 $X=3.64 $Y=3.03 $X2=0
+ $Y2=0
cc_800 N_SCE_c_990_n N_VPWR_c_2016_n 0.00310923f $X=4.55 $Y=3.105 $X2=0 $Y2=0
cc_801 N_SCE_M1003_g N_VPWR_c_2016_n 0.00117443f $X=4.64 $Y=2.595 $X2=0 $Y2=0
cc_802 N_SCE_c_991_n N_VPWR_c_2031_n 0.0245206f $X=3.715 $Y=3.105 $X2=0 $Y2=0
cc_803 N_SCE_c_990_n N_VPWR_c_2013_n 0.0258055f $X=4.55 $Y=3.105 $X2=0 $Y2=0
cc_804 N_SCE_c_991_n N_VPWR_c_2013_n 0.0100661f $X=3.715 $Y=3.105 $X2=0 $Y2=0
cc_805 N_SCE_c_989_n N_A_693_113#_c_2204_n 0.00196983f $X=3.64 $Y=3.03 $X2=0
+ $Y2=0
cc_806 N_SCE_M1003_g N_A_693_113#_c_2204_n 0.00440072f $X=4.64 $Y=2.595 $X2=0
+ $Y2=0
cc_807 N_SCE_c_989_n N_A_693_113#_c_2260_n 0.00538071f $X=3.64 $Y=3.03 $X2=0
+ $Y2=0
cc_808 N_SCE_c_990_n N_A_693_113#_c_2205_n 0.0224452f $X=4.55 $Y=3.105 $X2=0
+ $Y2=0
cc_809 N_SCE_M1003_g N_A_693_113#_c_2205_n 0.00872278f $X=4.64 $Y=2.595 $X2=0
+ $Y2=0
cc_810 N_SCE_c_989_n N_A_693_113#_c_2216_n 0.00373701f $X=3.64 $Y=3.03 $X2=0
+ $Y2=0
cc_811 N_SCE_c_990_n N_A_693_113#_c_2216_n 0.00837949f $X=4.55 $Y=3.105 $X2=0
+ $Y2=0
cc_812 N_SCE_c_991_n N_A_693_113#_c_2216_n 0.0013142f $X=3.715 $Y=3.105 $X2=0
+ $Y2=0
cc_813 N_SCE_M1003_g N_A_693_113#_c_2228_n 0.0162802f $X=4.64 $Y=2.595 $X2=0
+ $Y2=0
cc_814 N_SCE_c_993_n N_A_693_113#_c_2207_n 4.69291e-19 $X=4.64 $Y=2.2 $X2=0
+ $Y2=0
cc_815 N_SCE_M1003_g N_A_693_113#_c_2207_n 0.00578626f $X=4.64 $Y=2.595 $X2=0
+ $Y2=0
cc_816 N_SCE_c_989_n N_A_693_113#_c_2201_n 0.00415211f $X=3.64 $Y=3.03 $X2=0
+ $Y2=0
cc_817 N_SCE_M1004_g N_A_693_113#_c_2202_n 0.00981231f $X=5.625 $Y=0.835 $X2=0
+ $Y2=0
cc_818 N_SCE_M1004_g N_A_693_113#_c_2203_n 0.00168744f $X=5.625 $Y=0.835 $X2=0
+ $Y2=0
cc_819 N_SCE_M1031_g N_VGND_c_2408_n 0.00828092f $X=4.765 $Y=0.835 $X2=0 $Y2=0
cc_820 N_SCE_c_984_n N_VGND_c_2408_n 0.0240275f $X=5.55 $Y=0.18 $X2=0 $Y2=0
cc_821 N_SCE_M1004_g N_VGND_c_2408_n 0.00701307f $X=5.625 $Y=0.835 $X2=0 $Y2=0
cc_822 N_SCE_c_984_n N_VGND_c_2409_n 0.0111527f $X=5.55 $Y=0.18 $X2=0 $Y2=0
cc_823 N_SCE_c_984_n N_VGND_c_2416_n 0.0177004f $X=5.55 $Y=0.18 $X2=0 $Y2=0
cc_824 N_SCE_c_985_n N_VGND_c_2420_n 0.00729633f $X=4.84 $Y=0.18 $X2=0 $Y2=0
cc_825 N_SCE_c_984_n N_VGND_c_2435_n 0.0293095f $X=5.55 $Y=0.18 $X2=0 $Y2=0
cc_826 N_SCE_c_985_n N_VGND_c_2435_n 0.0106185f $X=4.84 $Y=0.18 $X2=0 $Y2=0
cc_827 N_CLK_c_1068_n N_A_1340_74#_M1024_g 0.00318552f $X=6.755 $Y=1.745 $X2=0
+ $Y2=0
cc_828 N_CLK_c_1067_n N_A_1340_74#_c_1347_n 0.00765331f $X=6.625 $Y=1.22 $X2=0
+ $Y2=0
cc_829 N_CLK_c_1067_n N_A_1340_74#_c_1348_n 0.00256256f $X=6.625 $Y=1.22 $X2=0
+ $Y2=0
cc_830 N_CLK_c_1068_n N_A_1340_74#_c_1348_n 0.00441194f $X=6.755 $Y=1.745 $X2=0
+ $Y2=0
cc_831 CLK N_A_1340_74#_c_1348_n 0.0264662f $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_832 N_CLK_c_1067_n N_A_1340_74#_c_1349_n 0.00414863f $X=6.625 $Y=1.22 $X2=0
+ $Y2=0
cc_833 N_CLK_c_1068_n N_A_1340_74#_c_1349_n 0.00477883f $X=6.755 $Y=1.745 $X2=0
+ $Y2=0
cc_834 CLK N_A_1340_74#_c_1349_n 0.00287256f $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_835 N_CLK_c_1068_n N_A_1340_74#_c_1350_n 0.00928281f $X=6.755 $Y=1.745 $X2=0
+ $Y2=0
cc_836 CLK N_A_1340_74#_c_1350_n 0.00160974f $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_837 N_CLK_c_1068_n N_A_1340_74#_c_1351_n 0.0112794f $X=6.755 $Y=1.745 $X2=0
+ $Y2=0
cc_838 N_CLK_c_1068_n N_VPWR_c_2017_n 0.0184615f $X=6.755 $Y=1.745 $X2=0 $Y2=0
cc_839 N_CLK_c_1068_n N_VPWR_c_2033_n 0.00505726f $X=6.755 $Y=1.745 $X2=0 $Y2=0
cc_840 N_CLK_c_1068_n N_VPWR_c_2013_n 0.00489105f $X=6.755 $Y=1.745 $X2=0 $Y2=0
cc_841 N_CLK_c_1068_n N_A_693_113#_c_2206_n 4.24902e-19 $X=6.755 $Y=1.745 $X2=0
+ $Y2=0
cc_842 N_CLK_c_1068_n N_A_693_113#_c_2208_n 0.0199322f $X=6.755 $Y=1.745 $X2=0
+ $Y2=0
cc_843 N_CLK_c_1067_n N_A_693_113#_c_2202_n 0.006603f $X=6.625 $Y=1.22 $X2=0
+ $Y2=0
cc_844 N_CLK_c_1067_n N_A_693_113#_c_2203_n 0.00256104f $X=6.625 $Y=1.22 $X2=0
+ $Y2=0
cc_845 N_CLK_c_1068_n N_A_693_113#_c_2203_n 0.0197522f $X=6.755 $Y=1.745 $X2=0
+ $Y2=0
cc_846 CLK N_A_693_113#_c_2203_n 0.0279729f $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_847 N_CLK_c_1068_n N_A_693_113#_c_2214_n 0.00297827f $X=6.755 $Y=1.745 $X2=0
+ $Y2=0
cc_848 N_CLK_c_1067_n N_VGND_c_2409_n 0.00490233f $X=6.625 $Y=1.22 $X2=0 $Y2=0
cc_849 N_CLK_c_1068_n N_VGND_c_2409_n 6.09068e-19 $X=6.755 $Y=1.745 $X2=0 $Y2=0
cc_850 CLK N_VGND_c_2409_n 0.00393057f $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_851 N_CLK_c_1067_n N_VGND_c_2410_n 0.00354158f $X=6.625 $Y=1.22 $X2=0 $Y2=0
cc_852 N_CLK_c_1067_n N_VGND_c_2421_n 0.00434272f $X=6.625 $Y=1.22 $X2=0 $Y2=0
cc_853 N_CLK_c_1067_n N_VGND_c_2435_n 0.00830282f $X=6.625 $Y=1.22 $X2=0 $Y2=0
cc_854 N_A_1538_74#_c_1104_n N_A_1340_74#_M1024_g 0.0098853f $X=7.83 $Y=0.515
+ $X2=0 $Y2=0
cc_855 N_A_1538_74#_c_1106_n N_A_1340_74#_M1024_g 0.00474255f $X=7.995 $Y=0.34
+ $X2=0 $Y2=0
cc_856 N_A_1538_74#_c_1104_n N_A_1340_74#_c_1339_n 0.0036247f $X=7.83 $Y=0.515
+ $X2=0 $Y2=0
cc_857 N_A_1538_74#_c_1129_n N_A_1340_74#_c_1354_n 0.00445689f $X=8.645 $Y=2.01
+ $X2=0 $Y2=0
cc_858 N_A_1538_74#_c_1107_n N_A_1340_74#_c_1354_n 9.25721e-19 $X=8.73 $Y=1.82
+ $X2=0 $Y2=0
cc_859 N_A_1538_74#_c_1133_n N_A_1340_74#_c_1354_n 0.00122318f $X=8.73 $Y=2.085
+ $X2=0 $Y2=0
cc_860 N_A_1538_74#_c_1134_n N_A_1340_74#_c_1354_n 0.00526331f $X=8.84 $Y=2.185
+ $X2=0 $Y2=0
cc_861 N_A_1538_74#_c_1129_n N_A_1340_74#_c_1340_n 0.012852f $X=8.645 $Y=2.01
+ $X2=0 $Y2=0
cc_862 N_A_1538_74#_c_1101_n N_A_1340_74#_M1012_g 0.0135328f $X=9.285 $Y=1.015
+ $X2=0 $Y2=0
cc_863 N_A_1538_74#_c_1104_n N_A_1340_74#_M1012_g 0.00327787f $X=7.83 $Y=0.515
+ $X2=0 $Y2=0
cc_864 N_A_1538_74#_c_1105_n N_A_1340_74#_M1012_g 0.00929412f $X=8.645 $Y=0.34
+ $X2=0 $Y2=0
cc_865 N_A_1538_74#_c_1107_n N_A_1340_74#_M1012_g 0.0287338f $X=8.73 $Y=1.82
+ $X2=0 $Y2=0
cc_866 N_A_1538_74#_c_1119_n N_A_1340_74#_M1012_g 0.00206916f $X=8.73 $Y=0.34
+ $X2=0 $Y2=0
cc_867 N_A_1538_74#_c_1121_n N_A_1340_74#_M1012_g 2.72689e-19 $X=9.49 $Y=0.85
+ $X2=0 $Y2=0
cc_868 N_A_1538_74#_c_1107_n N_A_1340_74#_c_1342_n 0.0078182f $X=8.73 $Y=1.82
+ $X2=0 $Y2=0
cc_869 N_A_1538_74#_c_1133_n N_A_1340_74#_c_1342_n 0.00111269f $X=8.73 $Y=2.085
+ $X2=0 $Y2=0
cc_870 N_A_1538_74#_c_1134_n N_A_1340_74#_c_1342_n 0.0058857f $X=8.84 $Y=2.185
+ $X2=0 $Y2=0
cc_871 N_A_1538_74#_c_1120_n N_A_1340_74#_c_1342_n 9.90768e-19 $X=9.49 $Y=0.935
+ $X2=0 $Y2=0
cc_872 N_A_1538_74#_c_1122_n N_A_1340_74#_c_1342_n 0.0227493f $X=9.49 $Y=1.18
+ $X2=0 $Y2=0
cc_873 N_A_1538_74#_c_1133_n N_A_1340_74#_c_1357_n 5.0577e-19 $X=8.73 $Y=2.085
+ $X2=0 $Y2=0
cc_874 N_A_1538_74#_c_1126_n N_A_1340_74#_c_1358_n 0.0101282f $X=9.155 $Y=2.465
+ $X2=0 $Y2=0
cc_875 N_A_1538_74#_c_1134_n N_A_1340_74#_c_1358_n 0.0153672f $X=8.84 $Y=2.185
+ $X2=0 $Y2=0
cc_876 N_A_1538_74#_c_1103_n N_A_1340_74#_c_1343_n 0.0182136f $X=13.21 $Y=2.375
+ $X2=0 $Y2=0
cc_877 N_A_1538_74#_c_1128_n N_A_1340_74#_c_1343_n 0.011586f $X=13.21 $Y=2.465
+ $X2=0 $Y2=0
cc_878 N_A_1538_74#_c_1116_n N_A_1340_74#_c_1343_n 8.48635e-19 $X=12.205
+ $Y=1.635 $X2=0 $Y2=0
cc_879 N_A_1538_74#_c_1117_n N_A_1340_74#_c_1343_n 0.0217312f $X=12.205 $Y=1.635
+ $X2=0 $Y2=0
cc_880 N_A_1538_74#_c_1118_n N_A_1340_74#_c_1343_n 0.0047697f $X=13.12 $Y=1.275
+ $X2=0 $Y2=0
cc_881 N_A_1538_74#_c_1124_n N_A_1340_74#_c_1343_n 5.03473e-19 $X=13.285
+ $Y=1.275 $X2=0 $Y2=0
cc_882 N_A_1538_74#_c_1125_n N_A_1340_74#_c_1343_n 0.02153f $X=13.285 $Y=1.42
+ $X2=0 $Y2=0
cc_883 N_A_1538_74#_M1040_g N_A_1340_74#_M1020_g 0.0311612f $X=12.295 $Y=0.69
+ $X2=0 $Y2=0
cc_884 N_A_1538_74#_c_1116_n N_A_1340_74#_M1020_g 6.57068e-19 $X=12.205 $Y=1.635
+ $X2=0 $Y2=0
cc_885 N_A_1538_74#_c_1118_n N_A_1340_74#_M1020_g 0.0110881f $X=13.12 $Y=1.275
+ $X2=0 $Y2=0
cc_886 N_A_1538_74#_c_1124_n N_A_1340_74#_M1020_g 0.001f $X=13.285 $Y=1.275
+ $X2=0 $Y2=0
cc_887 N_A_1538_74#_c_1125_n N_A_1340_74#_M1020_g 0.0101758f $X=13.285 $Y=1.42
+ $X2=0 $Y2=0
cc_888 N_A_1538_74#_c_1107_n N_A_1340_74#_c_1346_n 0.00619439f $X=8.73 $Y=1.82
+ $X2=0 $Y2=0
cc_889 N_A_1538_74#_c_1134_n N_A_1340_74#_c_1346_n 0.0160713f $X=8.84 $Y=2.185
+ $X2=0 $Y2=0
cc_890 N_A_1538_74#_c_1116_n N_A_1340_74#_c_1362_n 0.00959834f $X=12.205
+ $Y=1.635 $X2=0 $Y2=0
cc_891 N_A_1538_74#_c_1117_n N_A_1340_74#_c_1362_n 0.00166902f $X=12.205
+ $Y=1.635 $X2=0 $Y2=0
cc_892 N_A_1538_74#_c_1103_n N_A_1340_74#_c_1363_n 6.13746e-19 $X=13.21 $Y=2.375
+ $X2=0 $Y2=0
cc_893 N_A_1538_74#_c_1116_n N_A_1340_74#_c_1363_n 0.00311056f $X=12.205
+ $Y=1.635 $X2=0 $Y2=0
cc_894 N_A_1538_74#_c_1117_n N_A_1340_74#_c_1363_n 2.38342e-19 $X=12.205
+ $Y=1.635 $X2=0 $Y2=0
cc_895 N_A_1538_74#_c_1116_n N_A_1340_74#_c_1352_n 0.0147071f $X=12.205 $Y=1.635
+ $X2=0 $Y2=0
cc_896 N_A_1538_74#_c_1117_n N_A_1340_74#_c_1352_n 0.00105244f $X=12.205
+ $Y=1.635 $X2=0 $Y2=0
cc_897 N_A_1538_74#_c_1118_n N_A_1340_74#_c_1352_n 0.0230085f $X=13.12 $Y=1.275
+ $X2=0 $Y2=0
cc_898 N_A_1538_74#_c_1124_n N_A_1340_74#_c_1352_n 0.00345228f $X=13.285
+ $Y=1.275 $X2=0 $Y2=0
cc_899 N_A_1538_74#_c_1125_n N_A_1340_74#_c_1352_n 0.0019234f $X=13.285 $Y=1.42
+ $X2=0 $Y2=0
cc_900 N_A_1538_74#_c_1110_n N_A_1979_71#_M1017_d 0.00273752f $X=11.295 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_901 N_A_1538_74#_c_1101_n N_A_1979_71#_M1019_g 0.0109283f $X=9.285 $Y=1.015
+ $X2=0 $Y2=0
cc_902 N_A_1538_74#_c_1108_n N_A_1979_71#_M1019_g 6.9823e-19 $X=9.325 $Y=0.34
+ $X2=0 $Y2=0
cc_903 N_A_1538_74#_c_1109_n N_A_1979_71#_M1019_g 0.0136736f $X=10.535 $Y=0.935
+ $X2=0 $Y2=0
cc_904 N_A_1538_74#_c_1208_p N_A_1979_71#_M1019_g 0.00304387f $X=10.62 $Y=0.85
+ $X2=0 $Y2=0
cc_905 N_A_1538_74#_c_1120_n N_A_1979_71#_M1019_g 0.00191779f $X=9.49 $Y=0.935
+ $X2=0 $Y2=0
cc_906 N_A_1538_74#_c_1121_n N_A_1979_71#_M1019_g 0.00504823f $X=9.49 $Y=0.85
+ $X2=0 $Y2=0
cc_907 N_A_1538_74#_c_1122_n N_A_1979_71#_M1019_g 0.0183448f $X=9.49 $Y=1.18
+ $X2=0 $Y2=0
cc_908 N_A_1538_74#_M1040_g N_A_1979_71#_c_1528_n 0.00541818f $X=12.295 $Y=0.69
+ $X2=0 $Y2=0
cc_909 N_A_1538_74#_c_1116_n N_A_1979_71#_c_1528_n 0.00290016f $X=12.205
+ $Y=1.635 $X2=0 $Y2=0
cc_910 N_A_1538_74#_c_1117_n N_A_1979_71#_c_1528_n 0.019026f $X=12.205 $Y=1.635
+ $X2=0 $Y2=0
cc_911 N_A_1538_74#_c_1123_n N_A_1979_71#_c_1528_n 0.00122173f $X=12.205
+ $Y=1.275 $X2=0 $Y2=0
cc_912 N_A_1538_74#_M1040_g N_A_1979_71#_c_1530_n 0.0598858f $X=12.295 $Y=0.69
+ $X2=0 $Y2=0
cc_913 N_A_1538_74#_c_1110_n N_A_1979_71#_c_1530_n 6.63977e-19 $X=11.295 $Y=0.34
+ $X2=0 $Y2=0
cc_914 N_A_1538_74#_c_1112_n N_A_1979_71#_c_1530_n 0.004173f $X=11.38 $Y=0.85
+ $X2=0 $Y2=0
cc_915 N_A_1538_74#_c_1113_n N_A_1979_71#_c_1530_n 0.013812f $X=12.04 $Y=0.935
+ $X2=0 $Y2=0
cc_916 N_A_1538_74#_c_1115_n N_A_1979_71#_c_1530_n 0.00409215f $X=12.125 $Y=1.19
+ $X2=0 $Y2=0
cc_917 N_A_1538_74#_c_1109_n N_A_1979_71#_c_1531_n 0.0136568f $X=10.535 $Y=0.935
+ $X2=0 $Y2=0
cc_918 N_A_1538_74#_c_1109_n N_A_1979_71#_c_1532_n 0.00752165f $X=10.535
+ $Y=0.935 $X2=0 $Y2=0
cc_919 N_A_1538_74#_c_1110_n N_A_1979_71#_c_1532_n 0.0188549f $X=11.295 $Y=0.34
+ $X2=0 $Y2=0
cc_920 N_A_1538_74#_c_1112_n N_A_1979_71#_c_1532_n 0.0197429f $X=11.38 $Y=0.85
+ $X2=0 $Y2=0
cc_921 N_A_1538_74#_c_1114_n N_A_1979_71#_c_1532_n 0.0147457f $X=11.465 $Y=0.935
+ $X2=0 $Y2=0
cc_922 N_A_1538_74#_M1040_g N_A_1979_71#_c_1534_n 2.58966e-19 $X=12.295 $Y=0.69
+ $X2=0 $Y2=0
cc_923 N_A_1538_74#_c_1113_n N_A_1979_71#_c_1534_n 0.0244256f $X=12.04 $Y=0.935
+ $X2=0 $Y2=0
cc_924 N_A_1538_74#_c_1114_n N_A_1979_71#_c_1534_n 0.0139155f $X=11.465 $Y=0.935
+ $X2=0 $Y2=0
cc_925 N_A_1538_74#_c_1116_n N_A_1979_71#_c_1534_n 0.010054f $X=12.205 $Y=1.635
+ $X2=0 $Y2=0
cc_926 N_A_1538_74#_c_1123_n N_A_1979_71#_c_1534_n 0.0116173f $X=12.205 $Y=1.275
+ $X2=0 $Y2=0
cc_927 N_A_1538_74#_c_1110_n N_A_1979_71#_c_1535_n 0.00373856f $X=11.295 $Y=0.34
+ $X2=0 $Y2=0
cc_928 N_A_1538_74#_c_1113_n N_A_1979_71#_c_1535_n 0.0114193f $X=12.04 $Y=0.935
+ $X2=0 $Y2=0
cc_929 N_A_1538_74#_c_1114_n N_A_1979_71#_c_1535_n 0.00455553f $X=11.465
+ $Y=0.935 $X2=0 $Y2=0
cc_930 N_A_1538_74#_c_1109_n N_A_1979_71#_c_1536_n 0.0446734f $X=10.535 $Y=0.935
+ $X2=0 $Y2=0
cc_931 N_A_1538_74#_c_1120_n N_A_1979_71#_c_1536_n 0.00873996f $X=9.49 $Y=0.935
+ $X2=0 $Y2=0
cc_932 N_A_1538_74#_c_1122_n N_A_1979_71#_c_1536_n 5.80651e-19 $X=9.49 $Y=1.18
+ $X2=0 $Y2=0
cc_933 N_A_1538_74#_c_1109_n N_A_1979_71#_c_1538_n 0.00528445f $X=10.535
+ $Y=0.935 $X2=0 $Y2=0
cc_934 N_A_1538_74#_c_1107_n N_A_1736_97#_M1012_d 0.0043242f $X=8.73 $Y=1.82
+ $X2=-0.19 $Y2=-0.245
cc_935 N_A_1538_74#_c_1109_n N_A_1736_97#_M1017_g 0.00580245f $X=10.535 $Y=0.935
+ $X2=0 $Y2=0
cc_936 N_A_1538_74#_c_1208_p N_A_1736_97#_M1017_g 0.0119684f $X=10.62 $Y=0.85
+ $X2=0 $Y2=0
cc_937 N_A_1538_74#_c_1110_n N_A_1736_97#_M1017_g 0.0113672f $X=11.295 $Y=0.34
+ $X2=0 $Y2=0
cc_938 N_A_1538_74#_c_1111_n N_A_1736_97#_M1017_g 0.00333597f $X=10.705 $Y=0.34
+ $X2=0 $Y2=0
cc_939 N_A_1538_74#_c_1112_n N_A_1736_97#_M1017_g 0.00304194f $X=11.38 $Y=0.85
+ $X2=0 $Y2=0
cc_940 N_A_1538_74#_c_1101_n N_A_1736_97#_c_1634_n 0.00503807f $X=9.285 $Y=1.015
+ $X2=0 $Y2=0
cc_941 N_A_1538_74#_c_1107_n N_A_1736_97#_c_1634_n 0.0788002f $X=8.73 $Y=1.82
+ $X2=0 $Y2=0
cc_942 N_A_1538_74#_c_1108_n N_A_1736_97#_c_1634_n 0.012971f $X=9.325 $Y=0.34
+ $X2=0 $Y2=0
cc_943 N_A_1538_74#_c_1121_n N_A_1736_97#_c_1634_n 0.0436611f $X=9.49 $Y=0.85
+ $X2=0 $Y2=0
cc_944 N_A_1538_74#_c_1109_n N_A_1736_97#_c_1636_n 0.00408713f $X=10.535
+ $Y=0.935 $X2=0 $Y2=0
cc_945 N_A_1538_74#_c_1107_n N_A_1736_97#_c_1637_n 0.0117546f $X=8.73 $Y=1.82
+ $X2=0 $Y2=0
cc_946 N_A_1538_74#_c_1133_n N_A_1736_97#_c_1637_n 0.00210558f $X=8.73 $Y=2.085
+ $X2=0 $Y2=0
cc_947 N_A_1538_74#_c_1134_n N_A_1736_97#_c_1637_n 0.0034213f $X=8.84 $Y=2.185
+ $X2=0 $Y2=0
cc_948 N_A_1538_74#_c_1120_n N_A_1736_97#_c_1637_n 0.0104166f $X=9.49 $Y=0.935
+ $X2=0 $Y2=0
cc_949 N_A_1538_74#_c_1122_n N_A_1736_97#_c_1637_n 0.00184141f $X=9.49 $Y=1.18
+ $X2=0 $Y2=0
cc_950 N_A_1538_74#_c_1126_n N_A_1736_97#_c_1638_n 0.00682633f $X=9.155 $Y=2.465
+ $X2=0 $Y2=0
cc_951 N_A_1538_74#_c_1126_n N_A_1736_97#_c_1639_n 0.00260822f $X=9.155 $Y=2.465
+ $X2=0 $Y2=0
cc_952 N_A_1538_74#_c_1133_n N_A_1736_97#_c_1639_n 0.0333974f $X=8.73 $Y=2.085
+ $X2=0 $Y2=0
cc_953 N_A_1538_74#_c_1134_n N_A_1736_97#_c_1639_n 0.0114168f $X=8.84 $Y=2.185
+ $X2=0 $Y2=0
cc_954 N_A_1538_74#_M1040_g N_A_2474_74#_c_1723_n 7.35604e-19 $X=12.295 $Y=0.69
+ $X2=0 $Y2=0
cc_955 N_A_1538_74#_c_1118_n N_A_2474_74#_c_1724_n 0.028365f $X=13.12 $Y=1.275
+ $X2=0 $Y2=0
cc_956 N_A_1538_74#_c_1124_n N_A_2474_74#_c_1724_n 0.02584f $X=13.285 $Y=1.275
+ $X2=0 $Y2=0
cc_957 N_A_1538_74#_c_1125_n N_A_2474_74#_c_1724_n 8.40831e-19 $X=13.285 $Y=1.42
+ $X2=0 $Y2=0
cc_958 N_A_1538_74#_M1040_g N_A_2474_74#_c_1725_n 9.17078e-19 $X=12.295 $Y=0.69
+ $X2=0 $Y2=0
cc_959 N_A_1538_74#_c_1113_n N_A_2474_74#_c_1725_n 8.0891e-19 $X=12.04 $Y=0.935
+ $X2=0 $Y2=0
cc_960 N_A_1538_74#_c_1118_n N_A_2474_74#_c_1725_n 0.0268237f $X=13.12 $Y=1.275
+ $X2=0 $Y2=0
cc_961 N_A_1538_74#_c_1103_n N_A_2474_74#_c_1734_n 0.00842885f $X=13.21 $Y=2.375
+ $X2=0 $Y2=0
cc_962 N_A_1538_74#_c_1128_n N_A_2474_74#_c_1734_n 0.017419f $X=13.21 $Y=2.465
+ $X2=0 $Y2=0
cc_963 N_A_1538_74#_c_1103_n N_A_2474_74#_c_1735_n 0.00607654f $X=13.21 $Y=2.375
+ $X2=0 $Y2=0
cc_964 N_A_1538_74#_c_1124_n N_A_2474_74#_c_1735_n 0.0116579f $X=13.285 $Y=1.275
+ $X2=0 $Y2=0
cc_965 N_A_1538_74#_c_1125_n N_A_2474_74#_c_1735_n 0.00105037f $X=13.285 $Y=1.42
+ $X2=0 $Y2=0
cc_966 N_A_1538_74#_c_1103_n N_A_2474_74#_c_1736_n 0.0114833f $X=13.21 $Y=2.375
+ $X2=0 $Y2=0
cc_967 N_A_1538_74#_c_1118_n N_A_2474_74#_c_1736_n 0.00352142f $X=13.12 $Y=1.275
+ $X2=0 $Y2=0
cc_968 N_A_1538_74#_c_1124_n N_A_2474_74#_c_1736_n 0.00816138f $X=13.285
+ $Y=1.275 $X2=0 $Y2=0
cc_969 N_A_1538_74#_c_1103_n N_A_2474_74#_c_1726_n 0.00234444f $X=13.21 $Y=2.375
+ $X2=0 $Y2=0
cc_970 N_A_1538_74#_c_1124_n N_A_2474_74#_c_1726_n 0.0299545f $X=13.285 $Y=1.275
+ $X2=0 $Y2=0
cc_971 N_A_1538_74#_c_1125_n N_A_2474_74#_c_1726_n 0.00187211f $X=13.285 $Y=1.42
+ $X2=0 $Y2=0
cc_972 N_A_1538_74#_c_1128_n N_VPWR_c_2021_n 0.00144848f $X=13.21 $Y=2.465 $X2=0
+ $Y2=0
cc_973 N_A_1538_74#_c_1128_n N_VPWR_c_2027_n 0.00332301f $X=13.21 $Y=2.465 $X2=0
+ $Y2=0
cc_974 N_A_1538_74#_c_1126_n N_VPWR_c_2034_n 0.00411612f $X=9.155 $Y=2.465 $X2=0
+ $Y2=0
cc_975 N_A_1538_74#_c_1126_n N_VPWR_c_2013_n 0.00753176f $X=9.155 $Y=2.465 $X2=0
+ $Y2=0
cc_976 N_A_1538_74#_c_1128_n N_VPWR_c_2013_n 0.00529948f $X=13.21 $Y=2.465 $X2=0
+ $Y2=0
cc_977 N_A_1538_74#_c_1134_n N_VPWR_c_2013_n 3.25067e-19 $X=8.84 $Y=2.185 $X2=0
+ $Y2=0
cc_978 N_A_1538_74#_c_1129_n N_A_693_113#_c_2209_n 0.0164655f $X=8.645 $Y=2.01
+ $X2=0 $Y2=0
cc_979 N_A_1538_74#_c_1107_n N_A_693_113#_c_2209_n 0.00324754f $X=8.73 $Y=1.82
+ $X2=0 $Y2=0
cc_980 N_A_1538_74#_c_1129_n N_A_693_113#_c_2197_n 0.0178882f $X=8.645 $Y=2.01
+ $X2=0 $Y2=0
cc_981 N_A_1538_74#_c_1107_n N_A_693_113#_c_2197_n 0.0125466f $X=8.73 $Y=1.82
+ $X2=0 $Y2=0
cc_982 N_A_1538_74#_c_1104_n N_A_693_113#_c_2198_n 0.00624344f $X=7.83 $Y=0.515
+ $X2=0 $Y2=0
cc_983 N_A_1538_74#_c_1129_n N_A_693_113#_c_2284_n 0.00104513f $X=8.645 $Y=2.01
+ $X2=0 $Y2=0
cc_984 N_A_1538_74#_c_1104_n N_A_693_113#_c_2199_n 0.0353265f $X=7.83 $Y=0.515
+ $X2=0 $Y2=0
cc_985 N_A_1538_74#_c_1105_n N_A_693_113#_c_2199_n 0.0191962f $X=8.645 $Y=0.34
+ $X2=0 $Y2=0
cc_986 N_A_1538_74#_c_1107_n N_A_693_113#_c_2199_n 0.0528515f $X=8.73 $Y=1.82
+ $X2=0 $Y2=0
cc_987 N_A_1538_74#_M1033_d N_A_693_113#_c_2210_n 0.00410007f $X=8.22 $Y=1.84
+ $X2=0 $Y2=0
cc_988 N_A_1538_74#_c_1126_n N_A_693_113#_c_2210_n 0.00127808f $X=9.155 $Y=2.465
+ $X2=0 $Y2=0
cc_989 N_A_1538_74#_c_1129_n N_A_693_113#_c_2210_n 0.0110685f $X=8.645 $Y=2.01
+ $X2=0 $Y2=0
cc_990 N_A_1538_74#_c_1133_n N_A_693_113#_c_2210_n 0.0296089f $X=8.73 $Y=2.085
+ $X2=0 $Y2=0
cc_991 N_A_1538_74#_c_1134_n N_A_693_113#_c_2210_n 0.00285137f $X=8.84 $Y=2.185
+ $X2=0 $Y2=0
cc_992 N_A_1538_74#_c_1126_n N_A_693_113#_c_2211_n 0.00152236f $X=9.155 $Y=2.465
+ $X2=0 $Y2=0
cc_993 N_A_1538_74#_M1033_d N_A_693_113#_c_2294_n 0.00763764f $X=8.22 $Y=1.84
+ $X2=0 $Y2=0
cc_994 N_A_1538_74#_c_1126_n N_A_693_113#_c_2294_n 0.00115318f $X=9.155 $Y=2.465
+ $X2=0 $Y2=0
cc_995 N_A_1538_74#_c_1129_n N_A_693_113#_c_2294_n 0.0119472f $X=8.645 $Y=2.01
+ $X2=0 $Y2=0
cc_996 N_A_1538_74#_c_1134_n N_A_693_113#_c_2294_n 0.00204278f $X=8.84 $Y=2.185
+ $X2=0 $Y2=0
cc_997 N_A_1538_74#_c_1109_n N_VGND_M1019_d 0.00739508f $X=10.535 $Y=0.935 $X2=0
+ $Y2=0
cc_998 N_A_1538_74#_c_1208_p N_VGND_M1019_d 0.00497836f $X=10.62 $Y=0.85 $X2=0
+ $Y2=0
cc_999 N_A_1538_74#_c_1111_n N_VGND_M1019_d 5.40435e-19 $X=10.705 $Y=0.34 $X2=0
+ $Y2=0
cc_1000 N_A_1538_74#_c_1113_n N_VGND_M1039_s 0.00391333f $X=12.04 $Y=0.935 $X2=0
+ $Y2=0
cc_1001 N_A_1538_74#_c_1104_n N_VGND_c_2410_n 0.0259603f $X=7.83 $Y=0.515 $X2=0
+ $Y2=0
cc_1002 N_A_1538_74#_c_1106_n N_VGND_c_2410_n 0.0112234f $X=7.995 $Y=0.34 $X2=0
+ $Y2=0
cc_1003 N_A_1538_74#_c_1108_n N_VGND_c_2411_n 0.00608133f $X=9.325 $Y=0.34 $X2=0
+ $Y2=0
cc_1004 N_A_1538_74#_c_1109_n N_VGND_c_2411_n 0.0208664f $X=10.535 $Y=0.935
+ $X2=0 $Y2=0
cc_1005 N_A_1538_74#_c_1208_p N_VGND_c_2411_n 0.0191216f $X=10.62 $Y=0.85 $X2=0
+ $Y2=0
cc_1006 N_A_1538_74#_c_1111_n N_VGND_c_2411_n 0.014628f $X=10.705 $Y=0.34 $X2=0
+ $Y2=0
cc_1007 N_A_1538_74#_c_1121_n N_VGND_c_2411_n 0.0046174f $X=9.49 $Y=0.85 $X2=0
+ $Y2=0
cc_1008 N_A_1538_74#_M1040_g N_VGND_c_2412_n 0.00149332f $X=12.295 $Y=0.69 $X2=0
+ $Y2=0
cc_1009 N_A_1538_74#_c_1110_n N_VGND_c_2412_n 0.0146661f $X=11.295 $Y=0.34 $X2=0
+ $Y2=0
cc_1010 N_A_1538_74#_c_1112_n N_VGND_c_2412_n 0.0193741f $X=11.38 $Y=0.85 $X2=0
+ $Y2=0
cc_1011 N_A_1538_74#_c_1113_n N_VGND_c_2412_n 0.015048f $X=12.04 $Y=0.935 $X2=0
+ $Y2=0
cc_1012 N_A_1538_74#_c_1101_n N_VGND_c_2422_n 7.53287e-19 $X=9.285 $Y=1.015
+ $X2=0 $Y2=0
cc_1013 N_A_1538_74#_c_1105_n N_VGND_c_2422_n 0.0418136f $X=8.645 $Y=0.34 $X2=0
+ $Y2=0
cc_1014 N_A_1538_74#_c_1106_n N_VGND_c_2422_n 0.0235688f $X=7.995 $Y=0.34 $X2=0
+ $Y2=0
cc_1015 N_A_1538_74#_c_1108_n N_VGND_c_2422_n 0.0449818f $X=9.325 $Y=0.34 $X2=0
+ $Y2=0
cc_1016 N_A_1538_74#_c_1119_n N_VGND_c_2422_n 0.0121867f $X=8.73 $Y=0.34 $X2=0
+ $Y2=0
cc_1017 N_A_1538_74#_c_1110_n N_VGND_c_2423_n 0.0498034f $X=11.295 $Y=0.34 $X2=0
+ $Y2=0
cc_1018 N_A_1538_74#_c_1111_n N_VGND_c_2423_n 0.0120637f $X=10.705 $Y=0.34 $X2=0
+ $Y2=0
cc_1019 N_A_1538_74#_M1040_g N_VGND_c_2432_n 0.00461464f $X=12.295 $Y=0.69 $X2=0
+ $Y2=0
cc_1020 N_A_1538_74#_M1040_g N_VGND_c_2435_n 0.0090922f $X=12.295 $Y=0.69 $X2=0
+ $Y2=0
cc_1021 N_A_1538_74#_c_1105_n N_VGND_c_2435_n 0.0244305f $X=8.645 $Y=0.34 $X2=0
+ $Y2=0
cc_1022 N_A_1538_74#_c_1106_n N_VGND_c_2435_n 0.0127152f $X=7.995 $Y=0.34 $X2=0
+ $Y2=0
cc_1023 N_A_1538_74#_c_1108_n N_VGND_c_2435_n 0.025776f $X=9.325 $Y=0.34 $X2=0
+ $Y2=0
cc_1024 N_A_1538_74#_c_1109_n N_VGND_c_2435_n 0.0214463f $X=10.535 $Y=0.935
+ $X2=0 $Y2=0
cc_1025 N_A_1538_74#_c_1110_n N_VGND_c_2435_n 0.0282611f $X=11.295 $Y=0.34 $X2=0
+ $Y2=0
cc_1026 N_A_1538_74#_c_1111_n N_VGND_c_2435_n 0.00644906f $X=10.705 $Y=0.34
+ $X2=0 $Y2=0
cc_1027 N_A_1538_74#_c_1113_n N_VGND_c_2435_n 0.0176914f $X=12.04 $Y=0.935 $X2=0
+ $Y2=0
cc_1028 N_A_1538_74#_c_1119_n N_VGND_c_2435_n 0.00660921f $X=8.73 $Y=0.34 $X2=0
+ $Y2=0
cc_1029 N_A_1538_74#_c_1120_n N_VGND_c_2435_n 0.00602284f $X=9.49 $Y=0.935 $X2=0
+ $Y2=0
cc_1030 N_A_1538_74#_c_1109_n A_1872_97# 0.0038466f $X=10.535 $Y=0.935 $X2=-0.19
+ $Y2=-0.245
cc_1031 N_A_1538_74#_c_1120_n A_1872_97# 0.00379972f $X=9.49 $Y=0.935 $X2=-0.19
+ $Y2=-0.245
cc_1032 N_A_1538_74#_c_1121_n A_1872_97# 0.00547066f $X=9.49 $Y=0.85 $X2=-0.19
+ $Y2=-0.245
cc_1033 N_A_1538_74#_c_1113_n A_2402_74# 0.00229931f $X=12.04 $Y=0.935 $X2=-0.19
+ $Y2=-0.245
cc_1034 N_A_1340_74#_c_1362_n N_A_1979_71#_M1030_d 0.0081007f $X=12.56 $Y=2.475
+ $X2=0 $Y2=0
cc_1035 N_A_1340_74#_c_1342_n N_A_1979_71#_c_1527_n 0.0129715f $X=9.505 $Y=1.69
+ $X2=0 $Y2=0
cc_1036 N_A_1340_74#_c_1358_n N_A_1979_71#_c_1527_n 0.022808f $X=9.605 $Y=2.465
+ $X2=0 $Y2=0
cc_1037 N_A_1340_74#_c_1366_n N_A_1979_71#_c_1527_n 0.00847136f $X=9.69 $Y=2.185
+ $X2=0 $Y2=0
cc_1038 N_A_1340_74#_c_1358_n N_A_1979_71#_c_1540_n 0.0178226f $X=9.605 $Y=2.465
+ $X2=0 $Y2=0
cc_1039 N_A_1340_74#_c_1362_n N_A_1979_71#_c_1540_n 0.0156192f $X=12.56 $Y=2.475
+ $X2=0 $Y2=0
cc_1040 N_A_1340_74#_c_1362_n N_A_1979_71#_c_1542_n 0.0202137f $X=12.56 $Y=2.475
+ $X2=0 $Y2=0
cc_1041 N_A_1340_74#_c_1362_n N_A_1979_71#_c_1544_n 0.0231265f $X=12.56 $Y=2.475
+ $X2=0 $Y2=0
cc_1042 N_A_1340_74#_c_1362_n N_A_1736_97#_c_1632_n 0.0164119f $X=12.56 $Y=2.475
+ $X2=0 $Y2=0
cc_1043 N_A_1340_74#_M1012_g N_A_1736_97#_c_1634_n 0.00341647f $X=8.605 $Y=0.695
+ $X2=0 $Y2=0
cc_1044 N_A_1340_74#_c_1342_n N_A_1736_97#_c_1634_n 0.00613057f $X=9.505 $Y=1.69
+ $X2=0 $Y2=0
cc_1045 N_A_1340_74#_c_1342_n N_A_1736_97#_c_1636_n 0.00686717f $X=9.505 $Y=1.69
+ $X2=0 $Y2=0
cc_1046 N_A_1340_74#_c_1357_n N_A_1736_97#_c_1636_n 0.0060253f $X=9.58 $Y=2.02
+ $X2=0 $Y2=0
cc_1047 N_A_1340_74#_c_1358_n N_A_1736_97#_c_1636_n 0.00137373f $X=9.605
+ $Y=2.465 $X2=0 $Y2=0
cc_1048 N_A_1340_74#_c_1362_n N_A_1736_97#_c_1636_n 0.0172473f $X=12.56 $Y=2.475
+ $X2=0 $Y2=0
cc_1049 N_A_1340_74#_c_1366_n N_A_1736_97#_c_1636_n 0.0228253f $X=9.69 $Y=2.185
+ $X2=0 $Y2=0
cc_1050 N_A_1340_74#_c_1342_n N_A_1736_97#_c_1637_n 0.0115003f $X=9.505 $Y=1.69
+ $X2=0 $Y2=0
cc_1051 N_A_1340_74#_c_1358_n N_A_1736_97#_c_1638_n 0.0109297f $X=9.605 $Y=2.465
+ $X2=0 $Y2=0
cc_1052 N_A_1340_74#_c_1366_n N_A_1736_97#_c_1638_n 0.00391347f $X=9.69 $Y=2.185
+ $X2=0 $Y2=0
cc_1053 N_A_1340_74#_c_1342_n N_A_1736_97#_c_1639_n 0.00106527f $X=9.505 $Y=1.69
+ $X2=0 $Y2=0
cc_1054 N_A_1340_74#_c_1357_n N_A_1736_97#_c_1639_n 0.00921692f $X=9.58 $Y=2.02
+ $X2=0 $Y2=0
cc_1055 N_A_1340_74#_c_1358_n N_A_1736_97#_c_1639_n 0.00131685f $X=9.605
+ $Y=2.465 $X2=0 $Y2=0
cc_1056 N_A_1340_74#_c_1366_n N_A_1736_97#_c_1639_n 0.0333545f $X=9.69 $Y=2.185
+ $X2=0 $Y2=0
cc_1057 N_A_1340_74#_c_1362_n N_A_1736_97#_c_1640_n 0.00733642f $X=12.56
+ $Y=2.475 $X2=0 $Y2=0
cc_1058 N_A_1340_74#_M1020_g N_A_2474_74#_c_1723_n 0.00995617f $X=12.77 $Y=0.58
+ $X2=0 $Y2=0
cc_1059 N_A_1340_74#_M1020_g N_A_2474_74#_c_1724_n 0.00821531f $X=12.77 $Y=0.58
+ $X2=0 $Y2=0
cc_1060 N_A_1340_74#_M1020_g N_A_2474_74#_c_1725_n 0.00270117f $X=12.77 $Y=0.58
+ $X2=0 $Y2=0
cc_1061 N_A_1340_74#_c_1343_n N_A_2474_74#_c_1734_n 0.0139495f $X=12.67 $Y=1.885
+ $X2=0 $Y2=0
cc_1062 N_A_1340_74#_c_1362_n N_A_2474_74#_c_1734_n 0.0140691f $X=12.56 $Y=2.475
+ $X2=0 $Y2=0
cc_1063 N_A_1340_74#_c_1363_n N_A_2474_74#_c_1734_n 0.0214863f $X=12.645 $Y=2.39
+ $X2=0 $Y2=0
cc_1064 N_A_1340_74#_c_1343_n N_A_2474_74#_c_1736_n 0.00284371f $X=12.67
+ $Y=1.885 $X2=0 $Y2=0
cc_1065 N_A_1340_74#_c_1363_n N_A_2474_74#_c_1736_n 0.0211419f $X=12.645 $Y=2.39
+ $X2=0 $Y2=0
cc_1066 N_A_1340_74#_c_1352_n N_A_2474_74#_c_1736_n 7.37738e-19 $X=12.745
+ $Y=1.635 $X2=0 $Y2=0
cc_1067 N_A_1340_74#_c_1362_n N_VPWR_M1001_d 0.00672263f $X=12.56 $Y=2.475 $X2=0
+ $Y2=0
cc_1068 N_A_1340_74#_c_1362_n N_VPWR_M1028_s 0.0132092f $X=12.56 $Y=2.475 $X2=0
+ $Y2=0
cc_1069 N_A_1340_74#_c_1354_n N_VPWR_c_2018_n 0.0191632f $X=8.145 $Y=1.765 $X2=0
+ $Y2=0
cc_1070 N_A_1340_74#_c_1358_n N_VPWR_c_2019_n 0.00127838f $X=9.605 $Y=2.465
+ $X2=0 $Y2=0
cc_1071 N_A_1340_74#_c_1362_n N_VPWR_c_2019_n 0.0213202f $X=12.56 $Y=2.475 $X2=0
+ $Y2=0
cc_1072 N_A_1340_74#_c_1362_n N_VPWR_c_2020_n 0.0221685f $X=12.56 $Y=2.475 $X2=0
+ $Y2=0
cc_1073 N_A_1340_74#_c_1343_n N_VPWR_c_2027_n 0.00461464f $X=12.67 $Y=1.885
+ $X2=0 $Y2=0
cc_1074 N_A_1340_74#_c_1354_n N_VPWR_c_2034_n 0.00413917f $X=8.145 $Y=1.765
+ $X2=0 $Y2=0
cc_1075 N_A_1340_74#_c_1358_n N_VPWR_c_2034_n 0.00445602f $X=9.605 $Y=2.465
+ $X2=0 $Y2=0
cc_1076 N_A_1340_74#_c_1354_n N_VPWR_c_2013_n 0.00407982f $X=8.145 $Y=1.765
+ $X2=0 $Y2=0
cc_1077 N_A_1340_74#_c_1358_n N_VPWR_c_2013_n 0.00894404f $X=9.605 $Y=2.465
+ $X2=0 $Y2=0
cc_1078 N_A_1340_74#_c_1343_n N_VPWR_c_2013_n 0.00499117f $X=12.67 $Y=1.885
+ $X2=0 $Y2=0
cc_1079 N_A_1340_74#_c_1362_n N_VPWR_c_2013_n 0.0797366f $X=12.56 $Y=2.475 $X2=0
+ $Y2=0
cc_1080 N_A_1340_74#_c_1366_n N_VPWR_c_2013_n 0.00697075f $X=9.69 $Y=2.185 $X2=0
+ $Y2=0
cc_1081 N_A_1340_74#_M1011_d N_A_693_113#_c_2208_n 0.00839555f $X=6.83 $Y=1.82
+ $X2=0 $Y2=0
cc_1082 N_A_1340_74#_c_1339_n N_A_693_113#_c_2208_n 0.0019256f $X=8.07 $Y=1.655
+ $X2=0 $Y2=0
cc_1083 N_A_1340_74#_c_1350_n N_A_693_113#_c_2208_n 0.058258f $X=7.45 $Y=1.695
+ $X2=0 $Y2=0
cc_1084 N_A_1340_74#_c_1351_n N_A_693_113#_c_2208_n 0.0117116f $X=7.45 $Y=1.695
+ $X2=0 $Y2=0
cc_1085 N_A_1340_74#_c_1339_n N_A_693_113#_c_2209_n 0.00845418f $X=8.07 $Y=1.655
+ $X2=0 $Y2=0
cc_1086 N_A_1340_74#_c_1354_n N_A_693_113#_c_2209_n 0.00634674f $X=8.145
+ $Y=1.765 $X2=0 $Y2=0
cc_1087 N_A_1340_74#_c_1350_n N_A_693_113#_c_2209_n 0.030781f $X=7.45 $Y=1.695
+ $X2=0 $Y2=0
cc_1088 N_A_1340_74#_c_1351_n N_A_693_113#_c_2209_n 0.00370578f $X=7.45 $Y=1.695
+ $X2=0 $Y2=0
cc_1089 N_A_1340_74#_c_1339_n N_A_693_113#_c_2197_n 0.00162422f $X=8.07 $Y=1.655
+ $X2=0 $Y2=0
cc_1090 N_A_1340_74#_c_1340_n N_A_693_113#_c_2197_n 0.0102855f $X=8.53 $Y=1.655
+ $X2=0 $Y2=0
cc_1091 N_A_1340_74#_M1012_g N_A_693_113#_c_2197_n 0.00146886f $X=8.605 $Y=0.695
+ $X2=0 $Y2=0
cc_1092 N_A_1340_74#_c_1345_n N_A_693_113#_c_2197_n 0.00713545f $X=8.145
+ $Y=1.655 $X2=0 $Y2=0
cc_1093 N_A_1340_74#_M1024_g N_A_693_113#_c_2198_n 0.00238026f $X=7.615 $Y=0.74
+ $X2=0 $Y2=0
cc_1094 N_A_1340_74#_c_1339_n N_A_693_113#_c_2198_n 0.00577896f $X=8.07 $Y=1.655
+ $X2=0 $Y2=0
cc_1095 N_A_1340_74#_c_1350_n N_A_693_113#_c_2198_n 0.00638169f $X=7.45 $Y=1.695
+ $X2=0 $Y2=0
cc_1096 N_A_1340_74#_c_1354_n N_A_693_113#_c_2284_n 0.0182322f $X=8.145 $Y=1.765
+ $X2=0 $Y2=0
cc_1097 N_A_1340_74#_M1024_g N_A_693_113#_c_2199_n 0.00960169f $X=7.615 $Y=0.74
+ $X2=0 $Y2=0
cc_1098 N_A_1340_74#_M1012_g N_A_693_113#_c_2199_n 0.0127542f $X=8.605 $Y=0.695
+ $X2=0 $Y2=0
cc_1099 N_A_1340_74#_c_1354_n N_A_693_113#_c_2211_n 0.00701557f $X=8.145
+ $Y=1.765 $X2=0 $Y2=0
cc_1100 N_A_1340_74#_c_1347_n N_A_693_113#_c_2202_n 0.00605527f $X=6.84 $Y=0.515
+ $X2=0 $Y2=0
cc_1101 N_A_1340_74#_c_1348_n N_A_693_113#_c_2202_n 0.00163551f $X=6.98 $Y=1.53
+ $X2=0 $Y2=0
cc_1102 N_A_1340_74#_c_1349_n N_A_693_113#_c_2202_n 0.00465443f $X=6.87 $Y=1.01
+ $X2=0 $Y2=0
cc_1103 N_A_1340_74#_c_1348_n N_A_693_113#_c_2203_n 0.00336942f $X=6.98 $Y=1.53
+ $X2=0 $Y2=0
cc_1104 N_A_1340_74#_c_1350_n N_A_693_113#_c_2203_n 0.0176968f $X=7.45 $Y=1.695
+ $X2=0 $Y2=0
cc_1105 N_A_1340_74#_c_1362_n A_1936_508# 0.00258756f $X=12.56 $Y=2.475
+ $X2=-0.19 $Y2=-0.245
cc_1106 N_A_1340_74#_c_1366_n A_1936_508# 0.00337569f $X=9.69 $Y=2.185 $X2=-0.19
+ $Y2=-0.245
cc_1107 N_A_1340_74#_c_1362_n A_2357_392# 0.0369361f $X=12.56 $Y=2.475 $X2=-0.19
+ $Y2=-0.245
cc_1108 N_A_1340_74#_c_1347_n N_VGND_c_2409_n 0.0128662f $X=6.84 $Y=0.515 $X2=0
+ $Y2=0
cc_1109 N_A_1340_74#_M1024_g N_VGND_c_2410_n 0.00473533f $X=7.615 $Y=0.74 $X2=0
+ $Y2=0
cc_1110 N_A_1340_74#_c_1347_n N_VGND_c_2410_n 0.0637571f $X=6.84 $Y=0.515 $X2=0
+ $Y2=0
cc_1111 N_A_1340_74#_c_1350_n N_VGND_c_2410_n 0.00966282f $X=7.45 $Y=1.695 $X2=0
+ $Y2=0
cc_1112 N_A_1340_74#_c_1351_n N_VGND_c_2410_n 0.00456957f $X=7.45 $Y=1.695 $X2=0
+ $Y2=0
cc_1113 N_A_1340_74#_c_1347_n N_VGND_c_2421_n 0.0172202f $X=6.84 $Y=0.515 $X2=0
+ $Y2=0
cc_1114 N_A_1340_74#_M1024_g N_VGND_c_2422_n 0.00430908f $X=7.615 $Y=0.74 $X2=0
+ $Y2=0
cc_1115 N_A_1340_74#_M1012_g N_VGND_c_2422_n 7.53287e-19 $X=8.605 $Y=0.695 $X2=0
+ $Y2=0
cc_1116 N_A_1340_74#_M1020_g N_VGND_c_2432_n 0.00434272f $X=12.77 $Y=0.58 $X2=0
+ $Y2=0
cc_1117 N_A_1340_74#_M1020_g N_VGND_c_2433_n 0.00148617f $X=12.77 $Y=0.58 $X2=0
+ $Y2=0
cc_1118 N_A_1340_74#_M1024_g N_VGND_c_2435_n 0.0082568f $X=7.615 $Y=0.74 $X2=0
+ $Y2=0
cc_1119 N_A_1340_74#_M1020_g N_VGND_c_2435_n 0.00448332f $X=12.77 $Y=0.58 $X2=0
+ $Y2=0
cc_1120 N_A_1340_74#_c_1347_n N_VGND_c_2435_n 0.0142062f $X=6.84 $Y=0.515 $X2=0
+ $Y2=0
cc_1121 N_A_1979_71#_c_1527_n N_A_1736_97#_c_1632_n 0.0240099f $X=10.155
+ $Y=2.375 $X2=0 $Y2=0
cc_1122 N_A_1979_71#_c_1540_n N_A_1736_97#_c_1632_n 0.00966501f $X=10.155
+ $Y=2.465 $X2=0 $Y2=0
cc_1123 N_A_1979_71#_c_1531_n N_A_1736_97#_c_1632_n 0.00524691f $X=10.875
+ $Y=1.275 $X2=0 $Y2=0
cc_1124 N_A_1979_71#_c_1533_n N_A_1736_97#_c_1632_n 0.0131636f $X=11.04 $Y=2.05
+ $X2=0 $Y2=0
cc_1125 N_A_1979_71#_c_1544_n N_A_1736_97#_c_1632_n 0.00363374f $X=11.04
+ $Y=2.135 $X2=0 $Y2=0
cc_1126 N_A_1979_71#_c_1538_n N_A_1736_97#_c_1632_n 0.0219807f $X=10.155 $Y=1.34
+ $X2=0 $Y2=0
cc_1127 N_A_1979_71#_M1019_g N_A_1736_97#_M1017_g 0.0116773f $X=9.97 $Y=0.695
+ $X2=0 $Y2=0
cc_1128 N_A_1979_71#_c_1531_n N_A_1736_97#_M1017_g 0.0147655f $X=10.875 $Y=1.275
+ $X2=0 $Y2=0
cc_1129 N_A_1979_71#_c_1532_n N_A_1736_97#_M1017_g 0.00642025f $X=10.96 $Y=0.81
+ $X2=0 $Y2=0
cc_1130 N_A_1979_71#_c_1535_n N_A_1736_97#_M1017_g 0.0152227f $X=11.635 $Y=1.355
+ $X2=0 $Y2=0
cc_1131 N_A_1979_71#_c_1536_n N_A_1736_97#_M1017_g 7.29242e-19 $X=10.245 $Y=1.34
+ $X2=0 $Y2=0
cc_1132 N_A_1979_71#_c_1537_n N_A_1736_97#_M1017_g 0.00466193f $X=10.875 $Y=1.19
+ $X2=0 $Y2=0
cc_1133 N_A_1979_71#_c_1538_n N_A_1736_97#_M1017_g 0.00830579f $X=10.155 $Y=1.34
+ $X2=0 $Y2=0
cc_1134 N_A_1979_71#_c_1527_n N_A_1736_97#_c_1636_n 0.0130754f $X=10.155
+ $Y=2.375 $X2=0 $Y2=0
cc_1135 N_A_1979_71#_c_1531_n N_A_1736_97#_c_1636_n 0.00764905f $X=10.875
+ $Y=1.275 $X2=0 $Y2=0
cc_1136 N_A_1979_71#_c_1536_n N_A_1736_97#_c_1636_n 0.0207638f $X=10.245 $Y=1.34
+ $X2=0 $Y2=0
cc_1137 N_A_1979_71#_c_1538_n N_A_1736_97#_c_1636_n 0.00447738f $X=10.155
+ $Y=1.34 $X2=0 $Y2=0
cc_1138 N_A_1979_71#_c_1540_n N_A_1736_97#_c_1638_n 0.00156791f $X=10.155
+ $Y=2.465 $X2=0 $Y2=0
cc_1139 N_A_1979_71#_c_1527_n N_A_1736_97#_c_1640_n 0.0012697f $X=10.155
+ $Y=2.375 $X2=0 $Y2=0
cc_1140 N_A_1979_71#_c_1531_n N_A_1736_97#_c_1640_n 0.0222299f $X=10.875
+ $Y=1.275 $X2=0 $Y2=0
cc_1141 N_A_1979_71#_c_1533_n N_A_1736_97#_c_1640_n 0.0215301f $X=11.04 $Y=2.05
+ $X2=0 $Y2=0
cc_1142 N_A_1979_71#_c_1544_n N_A_1736_97#_c_1640_n 0.00133552f $X=11.04
+ $Y=2.135 $X2=0 $Y2=0
cc_1143 N_A_1979_71#_c_1540_n N_VPWR_c_2019_n 0.0101378f $X=10.155 $Y=2.465
+ $X2=0 $Y2=0
cc_1144 N_A_1979_71#_c_1542_n N_VPWR_c_2020_n 0.0183827f $X=11.71 $Y=1.885 $X2=0
+ $Y2=0
cc_1145 N_A_1979_71#_c_1542_n N_VPWR_c_2027_n 0.00413917f $X=11.71 $Y=1.885
+ $X2=0 $Y2=0
cc_1146 N_A_1979_71#_c_1540_n N_VPWR_c_2034_n 0.00413917f $X=10.155 $Y=2.465
+ $X2=0 $Y2=0
cc_1147 N_A_1979_71#_c_1540_n N_VPWR_c_2013_n 0.00399549f $X=10.155 $Y=2.465
+ $X2=0 $Y2=0
cc_1148 N_A_1979_71#_c_1542_n N_VPWR_c_2013_n 0.00403443f $X=11.71 $Y=1.885
+ $X2=0 $Y2=0
cc_1149 N_A_1979_71#_M1019_g N_VGND_c_2411_n 0.00381481f $X=9.97 $Y=0.695 $X2=0
+ $Y2=0
cc_1150 N_A_1979_71#_c_1530_n N_VGND_c_2412_n 0.010644f $X=11.935 $Y=1.11 $X2=0
+ $Y2=0
cc_1151 N_A_1979_71#_M1019_g N_VGND_c_2422_n 0.00497279f $X=9.97 $Y=0.695 $X2=0
+ $Y2=0
cc_1152 N_A_1979_71#_c_1530_n N_VGND_c_2432_n 0.00383152f $X=11.935 $Y=1.11
+ $X2=0 $Y2=0
cc_1153 N_A_1979_71#_M1019_g N_VGND_c_2435_n 0.00509887f $X=9.97 $Y=0.695 $X2=0
+ $Y2=0
cc_1154 N_A_1979_71#_c_1530_n N_VGND_c_2435_n 0.00385458f $X=11.935 $Y=1.11
+ $X2=0 $Y2=0
cc_1155 N_A_1736_97#_c_1632_n N_VPWR_c_2019_n 0.00641581f $X=10.69 $Y=1.915
+ $X2=0 $Y2=0
cc_1156 N_A_1736_97#_c_1638_n N_VPWR_c_2019_n 0.00599853f $X=9.38 $Y=2.75 $X2=0
+ $Y2=0
cc_1157 N_A_1736_97#_c_1632_n N_VPWR_c_2020_n 0.00578989f $X=10.69 $Y=1.915
+ $X2=0 $Y2=0
cc_1158 N_A_1736_97#_c_1632_n N_VPWR_c_2025_n 0.00487664f $X=10.69 $Y=1.915
+ $X2=0 $Y2=0
cc_1159 N_A_1736_97#_c_1638_n N_VPWR_c_2034_n 0.015569f $X=9.38 $Y=2.75 $X2=0
+ $Y2=0
cc_1160 N_A_1736_97#_c_1632_n N_VPWR_c_2013_n 0.00505379f $X=10.69 $Y=1.915
+ $X2=0 $Y2=0
cc_1161 N_A_1736_97#_c_1638_n N_VPWR_c_2013_n 0.0128526f $X=9.38 $Y=2.75 $X2=0
+ $Y2=0
cc_1162 N_A_1736_97#_c_1638_n N_A_693_113#_c_2210_n 0.0140012f $X=9.38 $Y=2.75
+ $X2=0 $Y2=0
cc_1163 N_A_1736_97#_c_1638_n N_A_693_113#_c_2211_n 0.0221746f $X=9.38 $Y=2.75
+ $X2=0 $Y2=0
cc_1164 N_A_1736_97#_M1017_g N_VGND_c_2411_n 0.00195433f $X=10.745 $Y=0.69 $X2=0
+ $Y2=0
cc_1165 N_A_1736_97#_M1017_g N_VGND_c_2423_n 0.00278237f $X=10.745 $Y=0.69 $X2=0
+ $Y2=0
cc_1166 N_A_1736_97#_M1017_g N_VGND_c_2435_n 0.00363424f $X=10.745 $Y=0.69 $X2=0
+ $Y2=0
cc_1167 N_A_2474_74#_c_1729_n N_VPWR_c_2021_n 0.00634677f $X=14.34 $Y=2.245
+ $X2=0 $Y2=0
cc_1168 N_A_2474_74#_c_1734_n N_VPWR_c_2021_n 0.0119691f $X=12.985 $Y=2.75 $X2=0
+ $Y2=0
cc_1169 N_A_2474_74#_c_1729_n N_VPWR_c_2022_n 0.00385791f $X=14.34 $Y=2.245
+ $X2=0 $Y2=0
cc_1170 N_A_2474_74#_c_1718_n N_VPWR_c_2022_n 0.00141722f $X=15.25 $Y=1.485
+ $X2=0 $Y2=0
cc_1171 N_A_2474_74#_c_1730_n N_VPWR_c_2022_n 0.0153862f $X=15.35 $Y=1.765 $X2=0
+ $Y2=0
cc_1172 N_A_2474_74#_c_1731_n N_VPWR_c_2022_n 5.40159e-19 $X=15.815 $Y=1.765
+ $X2=0 $Y2=0
cc_1173 N_A_2474_74#_c_1730_n N_VPWR_c_2024_n 4.94953e-19 $X=15.35 $Y=1.765
+ $X2=0 $Y2=0
cc_1174 N_A_2474_74#_c_1731_n N_VPWR_c_2024_n 0.0117128f $X=15.815 $Y=1.765
+ $X2=0 $Y2=0
cc_1175 N_A_2474_74#_c_1734_n N_VPWR_c_2027_n 0.0151873f $X=12.985 $Y=2.75 $X2=0
+ $Y2=0
cc_1176 N_A_2474_74#_c_1729_n N_VPWR_c_2035_n 0.00445602f $X=14.34 $Y=2.245
+ $X2=0 $Y2=0
cc_1177 N_A_2474_74#_c_1730_n N_VPWR_c_2036_n 0.00413917f $X=15.35 $Y=1.765
+ $X2=0 $Y2=0
cc_1178 N_A_2474_74#_c_1731_n N_VPWR_c_2036_n 0.00413917f $X=15.815 $Y=1.765
+ $X2=0 $Y2=0
cc_1179 N_A_2474_74#_c_1729_n N_VPWR_c_2013_n 0.00463274f $X=14.34 $Y=2.245
+ $X2=0 $Y2=0
cc_1180 N_A_2474_74#_c_1730_n N_VPWR_c_2013_n 0.00817869f $X=15.35 $Y=1.765
+ $X2=0 $Y2=0
cc_1181 N_A_2474_74#_c_1731_n N_VPWR_c_2013_n 0.00817869f $X=15.815 $Y=1.765
+ $X2=0 $Y2=0
cc_1182 N_A_2474_74#_c_1734_n N_VPWR_c_2013_n 0.0123029f $X=12.985 $Y=2.75 $X2=0
+ $Y2=0
cc_1183 N_A_2474_74#_M1008_g N_Q_c_2373_n 0.00818596f $X=15.325 $Y=0.74 $X2=0
+ $Y2=0
cc_1184 N_A_2474_74#_M1036_g N_Q_c_2373_n 0.00772833f $X=15.755 $Y=0.74 $X2=0
+ $Y2=0
cc_1185 N_A_2474_74#_M1008_g N_Q_c_2374_n 0.00582381f $X=15.325 $Y=0.74 $X2=0
+ $Y2=0
cc_1186 N_A_2474_74#_M1036_g N_Q_c_2374_n 0.0116235f $X=15.755 $Y=0.74 $X2=0
+ $Y2=0
cc_1187 N_A_2474_74#_c_1722_n N_Q_c_2374_n 0.0239602f $X=15.755 $Y=1.562 $X2=0
+ $Y2=0
cc_1188 N_A_2474_74#_c_1730_n N_Q_c_2377_n 4.00259e-19 $X=15.35 $Y=1.765 $X2=0
+ $Y2=0
cc_1189 N_A_2474_74#_c_1731_n N_Q_c_2377_n 4.00259e-19 $X=15.815 $Y=1.765 $X2=0
+ $Y2=0
cc_1190 N_A_2474_74#_c_1722_n N_Q_c_2377_n 5.15401e-19 $X=15.755 $Y=1.562 $X2=0
+ $Y2=0
cc_1191 N_A_2474_74#_M1008_g N_Q_c_2375_n 0.00840716f $X=15.325 $Y=0.74 $X2=0
+ $Y2=0
cc_1192 N_A_2474_74#_M1036_g N_Q_c_2375_n 0.00198651f $X=15.755 $Y=0.74 $X2=0
+ $Y2=0
cc_1193 N_A_2474_74#_c_1730_n Q 0.00211524f $X=15.35 $Y=1.765 $X2=0 $Y2=0
cc_1194 N_A_2474_74#_c_1731_n Q 0.0210093f $X=15.815 $Y=1.765 $X2=0 $Y2=0
cc_1195 N_A_2474_74#_c_1722_n Q 0.0297277f $X=15.755 $Y=1.562 $X2=0 $Y2=0
cc_1196 N_A_2474_74#_c_1723_n N_VGND_c_2412_n 0.0052468f $X=12.555 $Y=0.58 $X2=0
+ $Y2=0
cc_1197 N_A_2474_74#_M1023_g N_VGND_c_2413_n 0.00423534f $X=14.265 $Y=0.58 $X2=0
+ $Y2=0
cc_1198 N_A_2474_74#_c_1718_n N_VGND_c_2413_n 0.00588403f $X=15.25 $Y=1.485
+ $X2=0 $Y2=0
cc_1199 N_A_2474_74#_M1008_g N_VGND_c_2413_n 0.0149418f $X=15.325 $Y=0.74 $X2=0
+ $Y2=0
cc_1200 N_A_2474_74#_M1036_g N_VGND_c_2415_n 0.0184907f $X=15.755 $Y=0.74 $X2=0
+ $Y2=0
cc_1201 N_A_2474_74#_c_1722_n N_VGND_c_2415_n 6.84561e-19 $X=15.755 $Y=1.562
+ $X2=0 $Y2=0
cc_1202 N_A_2474_74#_M1023_g N_VGND_c_2424_n 0.00434272f $X=14.265 $Y=0.58 $X2=0
+ $Y2=0
cc_1203 N_A_2474_74#_M1008_g N_VGND_c_2425_n 0.00434272f $X=15.325 $Y=0.74 $X2=0
+ $Y2=0
cc_1204 N_A_2474_74#_M1036_g N_VGND_c_2425_n 0.00434272f $X=15.755 $Y=0.74 $X2=0
+ $Y2=0
cc_1205 N_A_2474_74#_c_1723_n N_VGND_c_2432_n 0.0145482f $X=12.555 $Y=0.58 $X2=0
+ $Y2=0
cc_1206 N_A_2474_74#_M1023_g N_VGND_c_2433_n 0.0115871f $X=14.265 $Y=0.58 $X2=0
+ $Y2=0
cc_1207 N_A_2474_74#_c_1723_n N_VGND_c_2433_n 0.0110541f $X=12.555 $Y=0.58 $X2=0
+ $Y2=0
cc_1208 N_A_2474_74#_c_1724_n N_VGND_c_2433_n 0.0454208f $X=13.62 $Y=0.935 $X2=0
+ $Y2=0
cc_1209 N_A_2474_74#_M1023_g N_VGND_c_2435_n 0.00830035f $X=14.265 $Y=0.58 $X2=0
+ $Y2=0
cc_1210 N_A_2474_74#_M1008_g N_VGND_c_2435_n 0.00825059f $X=15.325 $Y=0.74 $X2=0
+ $Y2=0
cc_1211 N_A_2474_74#_M1036_g N_VGND_c_2435_n 0.00823934f $X=15.755 $Y=0.74 $X2=0
+ $Y2=0
cc_1212 N_A_2474_74#_c_1723_n N_VGND_c_2435_n 0.0119922f $X=12.555 $Y=0.58 $X2=0
+ $Y2=0
cc_1213 N_A_2474_74#_c_1724_n N_VGND_c_2435_n 0.0168873f $X=13.62 $Y=0.935 $X2=0
+ $Y2=0
cc_1214 N_A_40_464#_c_1893_n A_129_464# 0.00595227f $X=1.47 $Y=2.375 $X2=-0.19
+ $Y2=-0.245
cc_1215 N_A_40_464#_c_1893_n N_VPWR_M1034_d 0.00509381f $X=1.47 $Y=2.375
+ $X2=-0.19 $Y2=-0.245
cc_1216 N_A_40_464#_c_1895_n N_VPWR_M1038_d 4.76982e-19 $X=2.15 $Y=2.99 $X2=0
+ $Y2=0
cc_1217 N_A_40_464#_c_1928_n N_VPWR_M1038_d 0.00490162f $X=2.235 $Y=2.905 $X2=0
+ $Y2=0
cc_1218 N_A_40_464#_c_1897_n N_VPWR_M1038_d 0.00972296f $X=3.25 $Y=2.375 $X2=0
+ $Y2=0
cc_1219 N_A_40_464#_c_1892_n N_VPWR_c_2014_n 0.010167f $X=0.345 $Y=2.465 $X2=0
+ $Y2=0
cc_1220 N_A_40_464#_c_1893_n N_VPWR_c_2014_n 0.0154248f $X=1.47 $Y=2.375 $X2=0
+ $Y2=0
cc_1221 N_A_40_464#_c_1894_n N_VPWR_c_2014_n 0.0208967f $X=1.555 $Y=2.905 $X2=0
+ $Y2=0
cc_1222 N_A_40_464#_c_1896_n N_VPWR_c_2014_n 0.0146662f $X=1.64 $Y=2.99 $X2=0
+ $Y2=0
cc_1223 N_A_40_464#_c_1895_n N_VPWR_c_2015_n 0.0145842f $X=2.15 $Y=2.99 $X2=0
+ $Y2=0
cc_1224 N_A_40_464#_c_1928_n N_VPWR_c_2015_n 0.0205316f $X=2.235 $Y=2.905 $X2=0
+ $Y2=0
cc_1225 N_A_40_464#_c_1897_n N_VPWR_c_2015_n 0.0154248f $X=3.25 $Y=2.375 $X2=0
+ $Y2=0
cc_1226 N_A_40_464#_c_1899_n N_VPWR_c_2015_n 0.0101141f $X=3.415 $Y=2.46 $X2=0
+ $Y2=0
cc_1227 N_A_40_464#_c_1892_n N_VPWR_c_2029_n 0.0188448f $X=0.345 $Y=2.465 $X2=0
+ $Y2=0
cc_1228 N_A_40_464#_c_1895_n N_VPWR_c_2030_n 0.0445209f $X=2.15 $Y=2.99 $X2=0
+ $Y2=0
cc_1229 N_A_40_464#_c_1896_n N_VPWR_c_2030_n 0.0121867f $X=1.64 $Y=2.99 $X2=0
+ $Y2=0
cc_1230 N_A_40_464#_c_1899_n N_VPWR_c_2031_n 0.0108086f $X=3.415 $Y=2.46 $X2=0
+ $Y2=0
cc_1231 N_A_40_464#_c_1892_n N_VPWR_c_2013_n 0.01556f $X=0.345 $Y=2.465 $X2=0
+ $Y2=0
cc_1232 N_A_40_464#_c_1895_n N_VPWR_c_2013_n 0.0250929f $X=2.15 $Y=2.99 $X2=0
+ $Y2=0
cc_1233 N_A_40_464#_c_1896_n N_VPWR_c_2013_n 0.00660921f $X=1.64 $Y=2.99 $X2=0
+ $Y2=0
cc_1234 N_A_40_464#_c_1899_n N_VPWR_c_2013_n 0.00906495f $X=3.415 $Y=2.46 $X2=0
+ $Y2=0
cc_1235 N_A_40_464#_c_1897_n A_575_463# 0.0048076f $X=3.25 $Y=2.375 $X2=-0.19
+ $Y2=-0.245
cc_1236 N_A_40_464#_c_1899_n N_A_693_113#_c_2260_n 0.033328f $X=3.415 $Y=2.46
+ $X2=0 $Y2=0
cc_1237 N_A_40_464#_c_1899_n N_A_693_113#_c_2216_n 0.00568204f $X=3.415 $Y=2.46
+ $X2=0 $Y2=0
cc_1238 N_A_40_464#_c_1889_n N_A_693_113#_c_2200_n 0.0138346f $X=3.255 $Y=0.84
+ $X2=0 $Y2=0
cc_1239 N_A_40_464#_c_1886_n N_A_693_113#_c_2201_n 0.00694013f $X=3.255 $Y=1.175
+ $X2=0 $Y2=0
cc_1240 N_A_40_464#_c_1887_n N_A_693_113#_c_2201_n 0.0700565f $X=3.415 $Y=2.29
+ $X2=0 $Y2=0
cc_1241 N_A_40_464#_c_1890_n N_A_693_113#_c_2201_n 0.0131144f $X=3.415 $Y=1.26
+ $X2=0 $Y2=0
cc_1242 N_A_40_464#_c_1902_n N_A_693_113#_c_2201_n 0.0138383f $X=3.375 $Y=2.375
+ $X2=0 $Y2=0
cc_1243 N_A_40_464#_c_1888_n N_VGND_c_2406_n 0.0149691f $X=0.4 $Y=0.58 $X2=0
+ $Y2=0
cc_1244 N_A_40_464#_c_1889_n N_VGND_c_2407_n 0.0107115f $X=3.255 $Y=0.84 $X2=0
+ $Y2=0
cc_1245 N_A_40_464#_c_1888_n N_VGND_c_2418_n 0.0206634f $X=0.4 $Y=0.58 $X2=0
+ $Y2=0
cc_1246 N_A_40_464#_c_1889_n N_VGND_c_2420_n 0.00699844f $X=3.255 $Y=0.84 $X2=0
+ $Y2=0
cc_1247 N_A_40_464#_c_1888_n N_VGND_c_2435_n 0.0173659f $X=0.4 $Y=0.58 $X2=0
+ $Y2=0
cc_1248 N_A_40_464#_c_1889_n N_VGND_c_2435_n 0.0134667f $X=3.255 $Y=0.84 $X2=0
+ $Y2=0
cc_1249 N_VPWR_c_2016_n N_A_693_113#_c_2205_n 0.0147124f $X=5.095 $Y=2.765 $X2=0
+ $Y2=0
cc_1250 N_VPWR_c_2031_n N_A_693_113#_c_2205_n 0.0561824f $X=5.01 $Y=3.33 $X2=0
+ $Y2=0
cc_1251 N_VPWR_c_2013_n N_A_693_113#_c_2205_n 0.0300887f $X=16.08 $Y=3.33 $X2=0
+ $Y2=0
cc_1252 N_VPWR_c_2031_n N_A_693_113#_c_2216_n 0.0190556f $X=5.01 $Y=3.33 $X2=0
+ $Y2=0
cc_1253 N_VPWR_c_2013_n N_A_693_113#_c_2216_n 0.00957028f $X=16.08 $Y=3.33 $X2=0
+ $Y2=0
cc_1254 N_VPWR_M1003_d N_A_693_113#_c_2228_n 0.00522241f $X=4.715 $Y=2.275 $X2=0
+ $Y2=0
cc_1255 N_VPWR_c_2016_n N_A_693_113#_c_2228_n 0.0231493f $X=5.095 $Y=2.765 $X2=0
+ $Y2=0
cc_1256 N_VPWR_M1003_d N_A_693_113#_c_2206_n 0.00977001f $X=4.715 $Y=2.275 $X2=0
+ $Y2=0
cc_1257 N_VPWR_c_2016_n N_A_693_113#_c_2206_n 0.0154248f $X=5.095 $Y=2.765 $X2=0
+ $Y2=0
cc_1258 N_VPWR_c_2013_n N_A_693_113#_c_2206_n 0.00387372f $X=16.08 $Y=3.33 $X2=0
+ $Y2=0
cc_1259 N_VPWR_M1011_s N_A_693_113#_c_2208_n 0.012925f $X=6.38 $Y=1.82 $X2=0
+ $Y2=0
cc_1260 N_VPWR_M1033_s N_A_693_113#_c_2208_n 0.00335285f $X=7.775 $Y=1.84 $X2=0
+ $Y2=0
cc_1261 N_VPWR_c_2017_n N_A_693_113#_c_2208_n 0.0218718f $X=6.525 $Y=2.795 $X2=0
+ $Y2=0
cc_1262 N_VPWR_c_2018_n N_A_693_113#_c_2208_n 0.008683f $X=7.92 $Y=2.805 $X2=0
+ $Y2=0
cc_1263 N_VPWR_c_2013_n N_A_693_113#_c_2208_n 0.0443221f $X=16.08 $Y=3.33 $X2=0
+ $Y2=0
cc_1264 N_VPWR_M1033_s N_A_693_113#_c_2209_n 0.012189f $X=7.775 $Y=1.84 $X2=0
+ $Y2=0
cc_1265 N_VPWR_c_2018_n N_A_693_113#_c_2284_n 9.99205e-19 $X=7.92 $Y=2.805 $X2=0
+ $Y2=0
cc_1266 N_VPWR_c_2013_n N_A_693_113#_c_2284_n 0.00535256f $X=16.08 $Y=3.33 $X2=0
+ $Y2=0
cc_1267 N_VPWR_c_2034_n N_A_693_113#_c_2210_n 0.0060566f $X=10.215 $Y=3.33 $X2=0
+ $Y2=0
cc_1268 N_VPWR_c_2013_n N_A_693_113#_c_2210_n 0.00967159f $X=16.08 $Y=3.33 $X2=0
+ $Y2=0
cc_1269 N_VPWR_c_2034_n N_A_693_113#_c_2211_n 0.0107588f $X=10.215 $Y=3.33 $X2=0
+ $Y2=0
cc_1270 N_VPWR_c_2013_n N_A_693_113#_c_2211_n 0.00904147f $X=16.08 $Y=3.33 $X2=0
+ $Y2=0
cc_1271 N_VPWR_c_2016_n N_A_693_113#_c_2214_n 0.00968143f $X=5.095 $Y=2.765
+ $X2=0 $Y2=0
cc_1272 N_VPWR_c_2017_n N_A_693_113#_c_2214_n 0.0151865f $X=6.525 $Y=2.795 $X2=0
+ $Y2=0
cc_1273 N_VPWR_c_2032_n N_A_693_113#_c_2214_n 0.0123502f $X=6.36 $Y=3.33 $X2=0
+ $Y2=0
cc_1274 N_VPWR_c_2013_n N_A_693_113#_c_2214_n 0.0117672f $X=16.08 $Y=3.33 $X2=0
+ $Y2=0
cc_1275 N_VPWR_M1033_s N_A_693_113#_c_2357_n 0.00183306f $X=7.775 $Y=1.84 $X2=0
+ $Y2=0
cc_1276 N_VPWR_c_2018_n N_A_693_113#_c_2357_n 0.0129485f $X=7.92 $Y=2.805 $X2=0
+ $Y2=0
cc_1277 N_VPWR_c_2013_n N_A_693_113#_c_2357_n 6.63299e-19 $X=16.08 $Y=3.33 $X2=0
+ $Y2=0
cc_1278 N_VPWR_c_2034_n N_A_693_113#_c_2294_n 0.0028606f $X=10.215 $Y=3.33 $X2=0
+ $Y2=0
cc_1279 N_VPWR_c_2013_n N_A_693_113#_c_2294_n 0.00491103f $X=16.08 $Y=3.33 $X2=0
+ $Y2=0
cc_1280 N_VPWR_c_2022_n N_Q_c_2377_n 0.0318992f $X=15.125 $Y=2.035 $X2=0 $Y2=0
cc_1281 N_VPWR_c_2024_n N_Q_c_2377_n 0.0255204f $X=16.04 $Y=2.405 $X2=0 $Y2=0
cc_1282 N_VPWR_c_2036_n N_Q_c_2377_n 0.0108429f $X=15.875 $Y=3.33 $X2=0 $Y2=0
cc_1283 N_VPWR_c_2013_n N_Q_c_2377_n 0.0089748f $X=16.08 $Y=3.33 $X2=0 $Y2=0
cc_1284 N_VPWR_M1027_d Q 0.00450961f $X=15.89 $Y=1.84 $X2=0 $Y2=0
cc_1285 N_VPWR_c_2024_n Q 0.0232122f $X=16.04 $Y=2.405 $X2=0 $Y2=0
cc_1286 N_A_693_113#_c_2206_n A_1079_455# 0.00595227f $X=5.8 $Y=2.34 $X2=-0.19
+ $Y2=-0.245
cc_1287 N_A_693_113#_c_2202_n N_VGND_c_2408_n 0.0137378f $X=5.84 $Y=0.835 $X2=0
+ $Y2=0
cc_1288 N_A_693_113#_c_2202_n N_VGND_c_2409_n 0.00498408f $X=5.84 $Y=0.835 $X2=0
+ $Y2=0
cc_1289 N_A_693_113#_c_2202_n N_VGND_c_2416_n 0.006859f $X=5.84 $Y=0.835 $X2=0
+ $Y2=0
cc_1290 N_A_693_113#_c_2200_n N_VGND_c_2420_n 0.00799869f $X=3.675 $Y=0.775
+ $X2=0 $Y2=0
cc_1291 N_A_693_113#_c_2200_n N_VGND_c_2435_n 0.0105426f $X=3.675 $Y=0.775 $X2=0
+ $Y2=0
cc_1292 N_A_693_113#_c_2202_n N_VGND_c_2435_n 0.00993188f $X=5.84 $Y=0.835 $X2=0
+ $Y2=0
cc_1293 N_Q_c_2373_n N_VGND_c_2413_n 0.0233039f $X=15.54 $Y=0.515 $X2=0 $Y2=0
cc_1294 N_Q_c_2373_n N_VGND_c_2415_n 0.0308109f $X=15.54 $Y=0.515 $X2=0 $Y2=0
cc_1295 Q N_VGND_c_2415_n 0.0156089f $X=15.995 $Y=1.58 $X2=0 $Y2=0
cc_1296 N_Q_c_2373_n N_VGND_c_2425_n 0.0144922f $X=15.54 $Y=0.515 $X2=0 $Y2=0
cc_1297 N_Q_c_2373_n N_VGND_c_2435_n 0.0118826f $X=15.54 $Y=0.515 $X2=0 $Y2=0
