* NGSPICE file created from sky130_fd_sc_ls__sdfxtp_4.ext - technology: sky130A

.subckt sky130_fd_sc_ls__sdfxtp_4 CLK D SCD SCE VGND VNB VPB VPWR Q
M1000 a_1026_100# a_828_74# a_301_74# VPB phighvt w=420000u l=150000u
+  ad=1.26e+11p pd=1.44e+06u as=3.159e+11p ps=3.31e+06u
M1001 a_630_74# CLK VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=1.77695e+12p ps=1.604e+07u
M1002 VPWR a_1814_48# Q VPB phighvt w=1.12e+06u l=150000u
+  ad=3.01978e+12p pd=2.28e+07u as=6.72e+11p ps=5.68e+06u
M1003 VGND a_1814_48# Q VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=4.773e+11p ps=4.25e+06u
M1004 a_1257_74# a_1026_100# VPWR VPB phighvt w=840000u l=150000u
+  ad=7.56e+11p pd=3.48e+06u as=0p ps=0u
M1005 a_1764_476# a_828_74# a_1587_74# VPB phighvt w=420000u l=150000u
+  ad=1.134e+11p pd=1.38e+06u as=2.898e+11p ps=2.46e+06u
M1006 VPWR a_1814_48# Q VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_301_74# D a_238_464# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1008 VGND SCD a_452_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1009 a_452_74# SCE a_301_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=3.738e+11p ps=3.46e+06u
M1010 a_1814_48# a_1587_74# VPWR VPB phighvt w=840000u l=150000u
+  ad=2.52e+11p pd=2.28e+06u as=0p ps=0u
M1011 a_1214_506# a_630_74# a_1026_100# VPB phighvt w=420000u l=150000u
+  ad=1.638e+11p pd=1.62e+06u as=0p ps=0u
M1012 a_1162_100# a_828_74# a_1026_100# VNB nshort w=420000u l=150000u
+  ad=1.995e+11p pd=1.79e+06u as=2.226e+11p ps=1.9e+06u
M1013 Q a_1814_48# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND a_1814_48# a_1766_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1015 Q a_1814_48# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_412_464# a_36_74# a_301_74# VPB phighvt w=640000u l=150000u
+  ad=2.496e+11p pd=2.06e+06u as=0p ps=0u
M1017 a_828_74# a_630_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=0p ps=0u
M1018 a_1766_74# a_630_74# a_1587_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=4e+11p ps=2.59e+06u
M1019 a_828_74# a_630_74# VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1020 a_223_74# a_36_74# VGND VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1021 a_301_74# D a_223_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_1587_74# a_630_74# a_1257_74# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_630_74# CLK VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=0p ps=0u
M1024 VPWR SCE a_36_74# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.888e+11p ps=1.87e+06u
M1025 a_1026_100# a_630_74# a_301_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VPWR a_1257_74# a_1214_506# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VGND a_1587_74# a_1814_48# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1028 VGND a_1814_48# Q VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPWR SCD a_412_464# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_1587_74# a_828_74# a_1257_74# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=2.365e+11p ps=1.96e+06u
M1031 a_238_464# SCE VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 Q a_1814_48# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 Q a_1814_48# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 VGND a_1257_74# a_1162_100# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_1257_74# a_1026_100# VGND VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 VGND SCE a_36_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1037 VPWR a_1814_48# a_1764_476# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 VPWR a_1587_74# a_1814_48# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

