* File: sky130_fd_sc_ls__or4bb_2.spice
* Created: Fri Aug 28 14:01:06 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__or4bb_2.pex.spice"
.subckt sky130_fd_sc_ls__or4bb_2  VNB VPB D_N B A C_N VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* C_N	C_N
* A	A
* B	B
* D_N	D_N
* VPB	VPB
* VNB	VNB
MM1004 N_VGND_M1004_d N_D_N_M1004_g N_A_27_424#_M1004_s VNB NSHORT L=0.15 W=0.55
+ AD=0.109083 AS=0.15675 PD=0.942248 PS=1.67 NRD=31.272 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75003.8 A=0.0825 P=1.4 MULT=1
MM1002 N_X_M1002_d N_A_182_270#_M1002_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.146767 PD=1.02 PS=1.26775 NRD=0 NRS=0.804 M=1 R=4.93333
+ SA=75000.6 SB=75002.7 A=0.111 P=1.78 MULT=1
MM1003 N_X_M1002_d N_A_182_270#_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.214171 PD=1.02 PS=1.42101 NRD=0 NRS=25.944 M=1 R=4.93333
+ SA=75001 SB=75002.3 A=0.111 P=1.78 MULT=1
MM1011 N_A_182_270#_M1011_d N_A_27_424#_M1011_g N_VGND_M1003_s VNB NSHORT L=0.15
+ W=0.64 AD=0.1668 AS=0.185229 PD=1.205 PS=1.22899 NRD=14.988 NRS=27.18 M=1
+ R=4.26667 SA=75001.8 SB=75001.9 A=0.096 P=1.58 MULT=1
MM1014 N_VGND_M1014_d N_A_548_110#_M1014_g N_A_182_270#_M1011_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.1248 AS=0.1668 PD=1.03 PS=1.205 NRD=0 NRS=23.904 M=1
+ R=4.26667 SA=75002.2 SB=75001.4 A=0.096 P=1.58 MULT=1
MM1000 N_A_182_270#_M1000_d N_B_M1000_g N_VGND_M1014_d VNB NSHORT L=0.15 W=0.64
+ AD=0.0928 AS=0.1248 PD=0.93 PS=1.03 NRD=0 NRS=20.616 M=1 R=4.26667 SA=75002.8
+ SB=75000.9 A=0.096 P=1.58 MULT=1
MM1012 N_VGND_M1012_d N_A_M1012_g N_A_182_270#_M1000_d VNB NSHORT L=0.15 W=0.64
+ AD=0.139765 AS=0.0928 PD=1.31765 PS=0.93 NRD=30.624 NRS=0 M=1 R=4.26667
+ SA=75003.2 SB=75000.5 A=0.096 P=1.58 MULT=1
MM1007 N_A_548_110#_M1007_d N_C_N_M1007_g N_VGND_M1012_d VNB NSHORT L=0.15
+ W=0.55 AD=0.15675 AS=0.12011 PD=1.67 PS=1.13235 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75002.4 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1010 N_VPWR_M1010_d N_D_N_M1010_g N_A_27_424#_M1010_s VPB PHIGHVT L=0.15
+ W=0.84 AD=0.1596 AS=0.2394 PD=1.26429 PS=2.25 NRD=14.0658 NRS=2.3443 M=1 R=5.6
+ SA=75000.2 SB=75001.2 A=0.126 P=1.98 MULT=1
MM1008 N_X_M1008_d N_A_182_270#_M1008_g N_VPWR_M1010_d VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.2128 PD=1.42 PS=1.68571 NRD=1.7533 NRS=2.6201 M=1 R=7.46667
+ SA=75000.6 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1013 N_X_M1008_d N_A_182_270#_M1013_g N_VPWR_M1013_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.3192 PD=1.42 PS=2.81 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1009 A_503_392# N_A_27_424#_M1009_g N_A_182_270#_M1009_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.285 PD=1.27 PS=2.57 NRD=15.7403 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75002 A=0.15 P=2.3 MULT=1
MM1005 A_587_392# N_A_548_110#_M1005_g A_503_392# VPB PHIGHVT L=0.15 W=1 AD=0.18
+ AS=0.135 PD=1.36 PS=1.27 NRD=24.6053 NRS=15.7403 M=1 R=6.66667 SA=75000.6
+ SB=75001.6 A=0.15 P=2.3 MULT=1
MM1006 A_689_392# N_B_M1006_g A_587_392# VPB PHIGHVT L=0.15 W=1 AD=0.12 AS=0.18
+ PD=1.24 PS=1.36 NRD=12.7853 NRS=24.6053 M=1 R=6.66667 SA=75001.1 SB=75001.1
+ A=0.15 P=2.3 MULT=1
MM1015 N_VPWR_M1015_d N_A_M1015_g A_689_392# VPB PHIGHVT L=0.15 W=1 AD=0.203696
+ AS=0.12 PD=1.51087 PS=1.24 NRD=1.9503 NRS=12.7853 M=1 R=6.66667 SA=75001.5
+ SB=75000.7 A=0.15 P=2.3 MULT=1
MM1001 N_A_548_110#_M1001_d N_C_N_M1001_g N_VPWR_M1015_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.2436 AS=0.171104 PD=2.26 PS=1.26913 NRD=2.3443 NRS=24.034 M=1
+ R=5.6 SA=75002.1 SB=75000.2 A=0.126 P=1.98 MULT=1
DX16_noxref VNB VPB NWDIODE A=9.6348 P=14.08
c_607 A_587_392# 0 1.16141e-19 $X=2.935 $Y=1.96
*
.include "sky130_fd_sc_ls__or4bb_2.pxi.spice"
*
.ends
*
*
