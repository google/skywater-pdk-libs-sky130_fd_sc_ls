* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__dfxtp_2 CLK D VGND VNB VPB VPWR Q
X0 Q a_1217_314# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X1 VPWR D a_431_508# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 a_1125_508# a_1217_314# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 a_1019_424# a_27_74# a_1172_124# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_1217_314# a_1019_424# VGND VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X5 VGND D a_431_508# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_538_429# a_27_74# a_644_504# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 a_1217_314# a_1019_424# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 a_695_459# a_206_368# a_1019_424# VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X9 a_1019_424# a_206_368# a_1125_508# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X10 a_27_74# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X11 VPWR a_538_429# a_695_459# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X12 a_1172_124# a_1217_314# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 VGND a_27_74# a_206_368# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X14 a_431_508# a_27_74# a_538_429# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 a_538_429# a_206_368# a_708_101# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 VPWR a_1217_314# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X17 a_644_504# a_695_459# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X18 a_431_508# a_206_368# a_538_429# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X19 VGND a_1217_314# Q VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X20 Q a_1217_314# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X21 VPWR a_27_74# a_206_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X22 a_27_74# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X23 a_695_459# a_27_74# a_1019_424# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X24 VGND a_538_429# a_695_459# VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X25 a_708_101# a_695_459# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
