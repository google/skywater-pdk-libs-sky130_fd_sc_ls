* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__dfxbp_2 CLK D VGND VNB VPB VPWR Q Q_N
X0 VPWR a_1835_368# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X1 a_702_445# a_753_284# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 VGND a_1290_102# Q VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X3 VGND a_27_74# a_206_368# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X4 a_1208_479# a_1290_102# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 a_1248_128# a_1290_102# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 Q a_1290_102# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X7 VPWR a_558_445# a_753_284# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X8 a_558_445# a_27_74# a_702_445# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X9 a_717_102# a_753_284# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_451_503# a_27_74# a_558_445# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 a_1290_102# a_1000_424# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X12 a_1000_424# a_27_74# a_1248_128# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 Q a_1290_102# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X14 a_1290_102# a_1000_424# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X15 VPWR a_1000_424# a_1290_102# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X16 VPWR a_1290_102# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X17 a_451_503# a_206_368# a_558_445# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X18 a_1835_368# a_1290_102# VGND VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X19 a_27_74# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X20 Q_N a_1835_368# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X21 a_1000_424# a_206_368# a_1208_479# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X22 a_753_284# a_27_74# a_1000_424# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X23 VPWR D a_451_503# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X24 VPWR a_27_74# a_206_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X25 a_27_74# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X26 a_1835_368# a_1290_102# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X27 VGND a_558_445# a_753_284# VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X28 VGND D a_451_503# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X29 a_558_445# a_206_368# a_717_102# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X30 Q_N a_1835_368# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X31 a_753_284# a_206_368# a_1000_424# VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X32 VGND a_1835_368# Q_N VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
.ends
