* File: sky130_fd_sc_ls__nand4_1.spice
* Created: Fri Aug 28 13:34:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__nand4_1.pex.spice"
.subckt sky130_fd_sc_ls__nand4_1  VNB VPB D C B A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* B	B
* C	C
* D	D
* VPB	VPB
* VNB	VNB
MM1000 A_181_74# N_D_M1000_g N_VGND_M1000_s VNB NSHORT L=0.15 W=0.74 AD=0.0888
+ AS=0.2923 PD=0.98 PS=2.72 NRD=10.536 NRS=0 M=1 R=4.93333 SA=75000.3 SB=75001.7
+ A=0.111 P=1.78 MULT=1
MM1001 A_259_74# N_C_M1001_g A_181_74# VNB NSHORT L=0.15 W=0.74 AD=0.1554
+ AS=0.0888 PD=1.16 PS=0.98 NRD=25.128 NRS=10.536 M=1 R=4.93333 SA=75000.7
+ SB=75001.3 A=0.111 P=1.78 MULT=1
MM1002 A_373_74# N_B_M1002_g A_259_74# VNB NSHORT L=0.15 W=0.74 AD=0.1554
+ AS=0.1554 PD=1.16 PS=1.16 NRD=25.128 NRS=25.128 M=1 R=4.93333 SA=75001.3
+ SB=75000.8 A=0.111 P=1.78 MULT=1
MM1007 N_Y_M1007_d N_A_M1007_g A_373_74# VNB NSHORT L=0.15 W=0.74 AD=0.2085
+ AS=0.1554 PD=2.05 PS=1.16 NRD=0 NRS=25.128 M=1 R=4.93333 SA=75001.8 SB=75000.2
+ A=0.111 P=1.78 MULT=1
MM1003 N_Y_M1003_d N_D_M1003_g N_VPWR_M1003_s VPB PHIGHVT L=0.15 W=1.12 AD=0.168
+ AS=0.3864 PD=1.42 PS=2.93 NRD=1.7533 NRS=10.5395 M=1 R=7.46667 SA=75000.3
+ SB=75001.8 A=0.168 P=2.54 MULT=1
MM1005 N_VPWR_M1005_d N_C_M1005_g N_Y_M1003_d VPB PHIGHVT L=0.15 W=1.12
+ AD=0.2576 AS=0.168 PD=1.58 PS=1.42 NRD=14.9326 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75001.3 A=0.168 P=2.54 MULT=1
MM1004 N_Y_M1004_d N_B_M1004_g N_VPWR_M1005_d VPB PHIGHVT L=0.15 W=1.12 AD=0.196
+ AS=0.2576 PD=1.47 PS=1.58 NRD=1.7533 NRS=16.7056 M=1 R=7.46667 SA=75001.3
+ SB=75000.7 A=0.168 P=2.54 MULT=1
MM1006 N_VPWR_M1006_d N_A_M1006_g N_Y_M1004_d VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.196 PD=2.83 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75001.8 SB=75000.2 A=0.168 P=2.54 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.0636 P=10.24
*
.include "sky130_fd_sc_ls__nand4_1.pxi.spice"
*
.ends
*
*
