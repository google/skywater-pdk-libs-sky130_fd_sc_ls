* File: sky130_fd_sc_ls__dfrtn_1.pxi.spice
* Created: Fri Aug 28 13:14:06 2020
* 
x_PM_SKY130_FD_SC_LS__DFRTN_1%D N_D_c_240_n N_D_c_247_n N_D_c_248_n N_D_c_249_n
+ N_D_M1023_g N_D_M1029_g N_D_c_242_n N_D_c_243_n D D D N_D_c_244_n N_D_c_245_n
+ PM_SKY130_FD_SC_LS__DFRTN_1%D
x_PM_SKY130_FD_SC_LS__DFRTN_1%CLK_N N_CLK_N_M1027_g N_CLK_N_M1007_g CLK_N
+ N_CLK_N_c_279_n N_CLK_N_c_280_n N_CLK_N_c_283_n
+ PM_SKY130_FD_SC_LS__DFRTN_1%CLK_N
x_PM_SKY130_FD_SC_LS__DFRTN_1%A_507_347# N_A_507_347#_M1005_d
+ N_A_507_347#_M1017_d N_A_507_347#_c_321_n N_A_507_347#_M1013_g
+ N_A_507_347#_c_322_n N_A_507_347#_c_342_n N_A_507_347#_c_343_n
+ N_A_507_347#_M1018_g N_A_507_347#_c_323_n N_A_507_347#_c_345_n
+ N_A_507_347#_M1002_g N_A_507_347#_c_324_n N_A_507_347#_c_325_n
+ N_A_507_347#_c_326_n N_A_507_347#_M1022_g N_A_507_347#_c_327_n
+ N_A_507_347#_c_346_n N_A_507_347#_c_328_n N_A_507_347#_c_329_n
+ N_A_507_347#_c_330_n N_A_507_347#_c_331_n N_A_507_347#_c_332_n
+ N_A_507_347#_c_360_p N_A_507_347#_c_354_p N_A_507_347#_c_333_n
+ N_A_507_347#_c_334_n N_A_507_347#_c_335_n N_A_507_347#_c_336_n
+ N_A_507_347#_c_378_p N_A_507_347#_c_379_p N_A_507_347#_c_337_n
+ N_A_507_347#_c_338_n N_A_507_347#_c_339_n N_A_507_347#_c_340_n
+ N_A_507_347#_c_341_n PM_SKY130_FD_SC_LS__DFRTN_1%A_507_347#
x_PM_SKY130_FD_SC_LS__DFRTN_1%A_841_288# N_A_841_288#_M1020_d
+ N_A_841_288#_M1008_d N_A_841_288#_c_506_n N_A_841_288#_M1031_g
+ N_A_841_288#_M1026_g N_A_841_288#_c_507_n N_A_841_288#_c_500_n
+ N_A_841_288#_c_501_n N_A_841_288#_c_502_n N_A_841_288#_c_503_n
+ N_A_841_288#_c_504_n N_A_841_288#_c_510_n N_A_841_288#_c_539_p
+ N_A_841_288#_c_540_p N_A_841_288#_c_505_n
+ PM_SKY130_FD_SC_LS__DFRTN_1%A_841_288#
x_PM_SKY130_FD_SC_LS__DFRTN_1%RESET_B N_RESET_B_M1025_g N_RESET_B_c_606_n
+ N_RESET_B_c_607_n N_RESET_B_M1024_g N_RESET_B_c_609_n N_RESET_B_c_610_n
+ N_RESET_B_M1016_g N_RESET_B_c_592_n N_RESET_B_c_611_n N_RESET_B_M1009_g
+ N_RESET_B_M1010_g N_RESET_B_c_613_n N_RESET_B_c_614_n N_RESET_B_M1019_g
+ N_RESET_B_c_594_n N_RESET_B_c_615_n N_RESET_B_c_595_n N_RESET_B_c_596_n
+ N_RESET_B_c_597_n N_RESET_B_c_598_n N_RESET_B_c_599_n N_RESET_B_c_600_n
+ RESET_B N_RESET_B_c_601_n N_RESET_B_c_602_n N_RESET_B_c_603_n
+ N_RESET_B_c_682_n N_RESET_B_c_604_n N_RESET_B_c_605_n
+ PM_SKY130_FD_SC_LS__DFRTN_1%RESET_B
x_PM_SKY130_FD_SC_LS__DFRTN_1%A_714_127# N_A_714_127#_M1013_d
+ N_A_714_127#_M1011_d N_A_714_127#_M1009_d N_A_714_127#_M1020_g
+ N_A_714_127#_c_823_n N_A_714_127#_M1008_g N_A_714_127#_c_824_n
+ N_A_714_127#_c_825_n N_A_714_127#_c_830_n N_A_714_127#_c_831_n
+ N_A_714_127#_c_832_n N_A_714_127#_c_833_n N_A_714_127#_c_826_n
+ PM_SKY130_FD_SC_LS__DFRTN_1%A_714_127#
x_PM_SKY130_FD_SC_LS__DFRTN_1%A_300_74# N_A_300_74#_M1027_d N_A_300_74#_M1007_d
+ N_A_300_74#_c_938_n N_A_300_74#_M1017_g N_A_300_74#_M1005_g
+ N_A_300_74#_c_924_n N_A_300_74#_c_925_n N_A_300_74#_c_926_n
+ N_A_300_74#_c_940_n N_A_300_74#_c_941_n N_A_300_74#_c_942_n
+ N_A_300_74#_c_943_n N_A_300_74#_M1011_g N_A_300_74#_M1030_g
+ N_A_300_74#_c_928_n N_A_300_74#_M1006_g N_A_300_74#_c_944_n
+ N_A_300_74#_M1012_g N_A_300_74#_c_930_n N_A_300_74#_c_931_n
+ N_A_300_74#_c_932_n N_A_300_74#_c_947_n N_A_300_74#_c_948_n
+ N_A_300_74#_c_933_n N_A_300_74#_c_934_n N_A_300_74#_c_951_n
+ N_A_300_74#_c_952_n N_A_300_74#_c_935_n N_A_300_74#_c_936_n
+ N_A_300_74#_c_937_n PM_SKY130_FD_SC_LS__DFRTN_1%A_300_74#
x_PM_SKY130_FD_SC_LS__DFRTN_1%A_1598_93# N_A_1598_93#_M1001_d
+ N_A_1598_93#_M1019_d N_A_1598_93#_M1000_g N_A_1598_93#_c_1122_n
+ N_A_1598_93#_M1003_g N_A_1598_93#_c_1123_n N_A_1598_93#_c_1124_n
+ N_A_1598_93#_c_1125_n N_A_1598_93#_c_1119_n N_A_1598_93#_c_1127_n
+ N_A_1598_93#_c_1120_n PM_SKY130_FD_SC_LS__DFRTN_1%A_1598_93#
x_PM_SKY130_FD_SC_LS__DFRTN_1%A_1266_119# N_A_1266_119#_M1006_d
+ N_A_1266_119#_M1002_d N_A_1266_119#_c_1207_n N_A_1266_119#_M1001_g
+ N_A_1266_119#_c_1208_n N_A_1266_119#_c_1218_n N_A_1266_119#_c_1219_n
+ N_A_1266_119#_M1014_g N_A_1266_119#_c_1209_n N_A_1266_119#_c_1220_n
+ N_A_1266_119#_c_1210_n N_A_1266_119#_M1021_g N_A_1266_119#_c_1221_n
+ N_A_1266_119#_M1015_g N_A_1266_119#_c_1211_n N_A_1266_119#_c_1229_n
+ N_A_1266_119#_c_1222_n N_A_1266_119#_c_1212_n N_A_1266_119#_c_1213_n
+ N_A_1266_119#_c_1214_n N_A_1266_119#_c_1224_n N_A_1266_119#_c_1237_n
+ N_A_1266_119#_c_1215_n N_A_1266_119#_c_1216_n
+ PM_SKY130_FD_SC_LS__DFRTN_1%A_1266_119#
x_PM_SKY130_FD_SC_LS__DFRTN_1%A_1934_94# N_A_1934_94#_M1021_s
+ N_A_1934_94#_M1015_s N_A_1934_94#_c_1345_n N_A_1934_94#_M1028_g
+ N_A_1934_94#_c_1346_n N_A_1934_94#_M1004_g N_A_1934_94#_c_1352_n
+ N_A_1934_94#_c_1353_n N_A_1934_94#_c_1347_n N_A_1934_94#_c_1348_n
+ N_A_1934_94#_c_1349_n N_A_1934_94#_c_1350_n
+ PM_SKY130_FD_SC_LS__DFRTN_1%A_1934_94#
x_PM_SKY130_FD_SC_LS__DFRTN_1%VPWR N_VPWR_M1023_s N_VPWR_M1024_d N_VPWR_M1017_s
+ N_VPWR_M1031_d N_VPWR_M1008_s N_VPWR_M1003_d N_VPWR_M1014_d N_VPWR_M1015_d
+ N_VPWR_c_1406_n N_VPWR_c_1407_n N_VPWR_c_1408_n N_VPWR_c_1409_n
+ N_VPWR_c_1410_n N_VPWR_c_1411_n N_VPWR_c_1412_n N_VPWR_c_1413_n
+ N_VPWR_c_1414_n N_VPWR_c_1415_n N_VPWR_c_1416_n N_VPWR_c_1417_n
+ N_VPWR_c_1418_n N_VPWR_c_1419_n VPWR N_VPWR_c_1420_n N_VPWR_c_1421_n
+ N_VPWR_c_1422_n N_VPWR_c_1423_n N_VPWR_c_1424_n N_VPWR_c_1405_n
+ N_VPWR_c_1426_n N_VPWR_c_1427_n N_VPWR_c_1428_n N_VPWR_c_1429_n
+ N_VPWR_c_1430_n PM_SKY130_FD_SC_LS__DFRTN_1%VPWR
x_PM_SKY130_FD_SC_LS__DFRTN_1%A_33_74# N_A_33_74#_M1029_s N_A_33_74#_M1013_s
+ N_A_33_74#_M1023_d N_A_33_74#_M1011_s N_A_33_74#_c_1537_n N_A_33_74#_c_1543_n
+ N_A_33_74#_c_1544_n N_A_33_74#_c_1598_n N_A_33_74#_c_1538_n
+ N_A_33_74#_c_1546_n N_A_33_74#_c_1539_n N_A_33_74#_c_1540_n
+ N_A_33_74#_c_1547_n N_A_33_74#_c_1541_n N_A_33_74#_c_1548_n
+ N_A_33_74#_c_1618_n PM_SKY130_FD_SC_LS__DFRTN_1%A_33_74#
x_PM_SKY130_FD_SC_LS__DFRTN_1%Q N_Q_M1028_d N_Q_M1004_d N_Q_c_1642_n
+ N_Q_c_1643_n Q Q Q Q N_Q_c_1644_n PM_SKY130_FD_SC_LS__DFRTN_1%Q
x_PM_SKY130_FD_SC_LS__DFRTN_1%VGND N_VGND_M1025_d N_VGND_M1005_s N_VGND_M1016_d
+ N_VGND_M1000_d N_VGND_M1021_d N_VGND_c_1670_n N_VGND_c_1671_n N_VGND_c_1672_n
+ N_VGND_c_1673_n N_VGND_c_1674_n VGND N_VGND_c_1675_n N_VGND_c_1676_n
+ N_VGND_c_1677_n N_VGND_c_1678_n N_VGND_c_1679_n N_VGND_c_1680_n
+ N_VGND_c_1681_n N_VGND_c_1682_n N_VGND_c_1683_n N_VGND_c_1684_n
+ N_VGND_c_1685_n N_VGND_c_1686_n PM_SKY130_FD_SC_LS__DFRTN_1%VGND
cc_1 VNB N_D_c_240_n 0.00193067f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=1.92
cc_2 VNB N_D_M1029_g 0.027501f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=0.58
cc_3 VNB N_D_c_242_n 0.0345854f $X=-0.19 $Y=-0.245 $X2=0.352 $Y2=1.11
cc_4 VNB N_D_c_243_n 0.0230272f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.63
cc_5 VNB N_D_c_244_n 0.0384016f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.125
cc_6 VNB N_D_c_245_n 0.00478024f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.125
cc_7 VNB CLK_N 0.00476718f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.75
cc_8 VNB N_CLK_N_c_279_n 0.0300365f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=0.58
cc_9 VNB N_CLK_N_c_280_n 0.0183832f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.11
cc_10 VNB N_A_507_347#_c_321_n 0.0153846f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.75
cc_11 VNB N_A_507_347#_c_322_n 0.0127269f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_507_347#_c_323_n 0.0165317f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_507_347#_c_324_n 0.0171653f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_14 VNB N_A_507_347#_c_325_n 0.0191633f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_507_347#_c_326_n 0.0231425f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_507_347#_c_327_n 0.0278721f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_507_347#_c_328_n 0.00466045f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_507_347#_c_329_n 0.00927063f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_507_347#_c_330_n 0.0218387f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_507_347#_c_331_n 0.00899291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_507_347#_c_332_n 0.00201735f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_507_347#_c_333_n 0.0039155f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_507_347#_c_334_n 0.0193653f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_507_347#_c_335_n 0.00260538f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_507_347#_c_336_n 0.00739636f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_507_347#_c_337_n 0.00166696f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_507_347#_c_338_n 0.0294493f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_507_347#_c_339_n 0.00628108f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_507_347#_c_340_n 0.0185091f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_507_347#_c_341_n 0.0169284f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_841_288#_M1026_g 0.0269266f $X=-0.19 $Y=-0.245 $X2=0.352 $Y2=1.11
cc_32 VNB N_A_841_288#_c_500_n 0.00386614f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.995
cc_33 VNB N_A_841_288#_c_501_n 0.0239207f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_841_288#_c_502_n 0.013115f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_35 VNB N_A_841_288#_c_503_n 0.00513663f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_36 VNB N_A_841_288#_c_504_n 0.00112198f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_841_288#_c_505_n 0.0021497f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_RESET_B_M1025_g 0.0343992f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.07
cc_39 VNB N_RESET_B_c_592_n 0.00905845f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.63
cc_40 VNB N_RESET_B_M1010_g 0.034399f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_RESET_B_c_594_n 0.0147263f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_RESET_B_c_595_n 0.00379793f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_RESET_B_c_596_n 0.00230496f $X=-0.19 $Y=-0.245 $X2=0.237 $Y2=2.035
cc_44 VNB N_RESET_B_c_597_n 0.0136272f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_RESET_B_c_598_n 4.82544e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_RESET_B_c_599_n 6.54175e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_RESET_B_c_600_n 0.00357755f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_RESET_B_c_601_n 0.0365981f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_RESET_B_c_602_n 0.00380174f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_RESET_B_c_603_n 0.0157849f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_RESET_B_c_604_n 0.0153888f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_RESET_B_c_605_n 0.0154637f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_714_127#_M1020_g 0.018017f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.11
cc_54 VNB N_A_714_127#_c_823_n 0.00936981f $X=-0.19 $Y=-0.245 $X2=0.352 $Y2=1.11
cc_55 VNB N_A_714_127#_c_824_n 0.0201987f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_714_127#_c_825_n 0.0103252f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_57 VNB N_A_714_127#_c_826_n 0.00434299f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_300_74#_M1005_g 0.0109841f $X=-0.19 $Y=-0.245 $X2=0.352 $Y2=0.96
cc_59 VNB N_A_300_74#_c_924_n 0.109169f $X=-0.19 $Y=-0.245 $X2=0.352 $Y2=1.11
cc_60 VNB N_A_300_74#_c_925_n 0.0125115f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_61 VNB N_A_300_74#_c_926_n 0.0509496f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.63
cc_62 VNB N_A_300_74#_M1030_g 0.0379845f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.125
cc_63 VNB N_A_300_74#_c_928_n 0.148495f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.125
cc_64 VNB N_A_300_74#_M1006_g 0.030044f $X=-0.19 $Y=-0.245 $X2=0.237 $Y2=1.665
cc_65 VNB N_A_300_74#_c_930_n 0.0404677f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_300_74#_c_931_n 0.00646948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_300_74#_c_932_n 0.00749069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_300_74#_c_933_n 0.00283216f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_300_74#_c_934_n 0.00454971f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_300_74#_c_935_n 0.015793f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_300_74#_c_936_n 0.00265148f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_300_74#_c_937_n 0.018162f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_1598_93#_M1000_g 0.0473326f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=0.58
cc_74 VNB N_A_1598_93#_c_1119_n 0.0107986f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_1598_93#_c_1120_n 0.0121095f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_1266_119#_c_1207_n 0.0202606f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.75
cc_77 VNB N_A_1266_119#_c_1208_n 0.00226217f $X=-0.19 $Y=-0.245 $X2=0.525
+ $Y2=0.58
cc_78 VNB N_A_1266_119#_c_1209_n 0.0586053f $X=-0.19 $Y=-0.245 $X2=0.27
+ $Y2=1.465
cc_79 VNB N_A_1266_119#_c_1210_n 0.0219742f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.995
cc_80 VNB N_A_1266_119#_c_1211_n 0.00948676f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_1266_119#_c_1212_n 0.00100139f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_1266_119#_c_1213_n 0.0107396f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_1266_119#_c_1214_n 0.0235899f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_1266_119#_c_1215_n 5.53899e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_1266_119#_c_1216_n 0.024655f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_1934_94#_c_1345_n 0.0213736f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.75
cc_87 VNB N_A_1934_94#_c_1346_n 0.0409762f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=0.58
cc_88 VNB N_A_1934_94#_c_1347_n 0.00180273f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.995
cc_89 VNB N_A_1934_94#_c_1348_n 2.65185e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_1934_94#_c_1349_n 0.0106069f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.125
cc_91 VNB N_A_1934_94#_c_1350_n 0.00429191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_VPWR_c_1405_n 0.462217f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_33_74#_c_1537_n 0.0118682f $X=-0.19 $Y=-0.245 $X2=0.352 $Y2=1.11
cc_94 VNB N_A_33_74#_c_1538_n 6.12392e-19 $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_95 VNB N_A_33_74#_c_1539_n 0.00943902f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_33_74#_c_1540_n 0.00638058f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.125
cc_97 VNB N_A_33_74#_c_1541_n 0.0216357f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_Q_c_1642_n 0.0243417f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=0.58
cc_99 VNB N_Q_c_1643_n 0.00719696f $X=-0.19 $Y=-0.245 $X2=0.352 $Y2=0.96
cc_100 VNB N_Q_c_1644_n 0.0236409f $X=-0.19 $Y=-0.245 $X2=0.237 $Y2=1.295
cc_101 VNB N_VGND_c_1670_n 0.00928007f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_VGND_c_1671_n 0.00636257f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_103 VNB N_VGND_c_1672_n 0.00664093f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_VGND_c_1673_n 0.0246564f $X=-0.19 $Y=-0.245 $X2=0.237 $Y2=1.125
cc_105 VNB N_VGND_c_1674_n 0.017712f $X=-0.19 $Y=-0.245 $X2=0.237 $Y2=1.665
cc_106 VNB N_VGND_c_1675_n 0.0309922f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_VGND_c_1676_n 0.0195319f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_VGND_c_1677_n 0.0684194f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_VGND_c_1678_n 0.0716605f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_1679_n 0.0470737f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_1680_n 0.0198148f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_1681_n 0.597513f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_1682_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_1683_n 0.0044892f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_VGND_c_1684_n 0.0043699f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_VGND_c_1685_n 0.00846329f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_VGND_c_1686_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VPB N_D_c_240_n 0.0176231f $X=-0.19 $Y=1.66 $X2=0.36 $Y2=1.92
cc_119 VPB N_D_c_247_n 0.0220469f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=2.07
cc_120 VPB N_D_c_248_n 0.0223644f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=2.375
cc_121 VPB N_D_c_249_n 0.0276505f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=2.465
cc_122 VPB N_D_c_245_n 0.0217648f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.125
cc_123 VPB CLK_N 6.29912e-19 $X=-0.19 $Y=1.66 $X2=0.5 $Y2=2.75
cc_124 VPB N_CLK_N_c_279_n 0.0133601f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=0.58
cc_125 VPB N_CLK_N_c_283_n 0.016043f $X=-0.19 $Y=1.66 $X2=0.352 $Y2=0.96
cc_126 VPB N_A_507_347#_c_342_n 0.0126039f $X=-0.19 $Y=1.66 $X2=0.352 $Y2=0.96
cc_127 VPB N_A_507_347#_c_343_n 0.0129604f $X=-0.19 $Y=1.66 $X2=0.352 $Y2=1.11
cc_128 VPB N_A_507_347#_c_323_n 0.00582876f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_129 VPB N_A_507_347#_c_345_n 0.0310581f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=1.995
cc_130 VPB N_A_507_347#_c_346_n 0.013403f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_A_507_347#_c_329_n 0.00602251f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_A_507_347#_c_340_n 0.0254664f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_A_841_288#_c_506_n 0.0130943f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=0.96
cc_134 VPB N_A_841_288#_c_507_n 0.0247999f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.63
cc_135 VPB N_A_841_288#_c_500_n 8.82777e-19 $X=-0.19 $Y=1.66 $X2=0.5 $Y2=1.995
cc_136 VPB N_A_841_288#_c_501_n 0.0175338f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_A_841_288#_c_510_n 0.00690074f $X=-0.19 $Y=1.66 $X2=0.237 $Y2=1.295
cc_138 VPB N_A_841_288#_c_505_n 0.00306186f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_RESET_B_c_606_n 0.0294946f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=2.75
cc_140 VPB N_RESET_B_c_607_n 0.00535616f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=2.75
cc_141 VPB N_RESET_B_M1024_g 0.0222714f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=0.58
cc_142 VPB N_RESET_B_c_609_n 0.315603f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_143 VPB N_RESET_B_c_610_n 0.0123638f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.11
cc_144 VPB N_RESET_B_c_611_n 0.0209255f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=1.995
cc_145 VPB N_RESET_B_M1009_g 0.0265476f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.95
cc_146 VPB N_RESET_B_c_613_n 0.0283395f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.125
cc_147 VPB N_RESET_B_c_614_n 0.0223436f $X=-0.19 $Y=1.66 $X2=0.237 $Y2=1.125
cc_148 VPB N_RESET_B_c_615_n 0.010471f $X=-0.19 $Y=1.66 $X2=0.237 $Y2=1.665
cc_149 VPB N_RESET_B_c_595_n 0.0046103f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_150 VPB N_RESET_B_c_596_n 8.51761e-19 $X=-0.19 $Y=1.66 $X2=0.237 $Y2=2.035
cc_151 VPB N_RESET_B_c_597_n 0.00642192f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_152 VPB N_RESET_B_c_598_n 4.71639e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_153 VPB N_RESET_B_c_599_n 6.35107e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_154 VPB N_RESET_B_c_600_n 0.00257552f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_155 VPB N_RESET_B_c_601_n 0.00784665f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_156 VPB N_RESET_B_c_602_n 0.00172327f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_157 VPB N_RESET_B_c_603_n 0.0104353f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_158 VPB N_RESET_B_c_605_n 0.0112707f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_159 VPB N_A_714_127#_c_823_n 0.0340257f $X=-0.19 $Y=1.66 $X2=0.352 $Y2=1.11
cc_160 VPB N_A_714_127#_c_824_n 0.0166419f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_161 VPB N_A_714_127#_c_825_n 0.00241618f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_162 VPB N_A_714_127#_c_830_n 0.0153919f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.95
cc_163 VPB N_A_714_127#_c_831_n 0.00270356f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_164 VPB N_A_714_127#_c_832_n 0.0115736f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.125
cc_165 VPB N_A_714_127#_c_833_n 0.0125069f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.125
cc_166 VPB N_A_714_127#_c_826_n 0.00401148f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_167 VPB N_A_300_74#_c_938_n 0.0191333f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=2.75
cc_168 VPB N_A_300_74#_c_926_n 0.0177294f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.63
cc_169 VPB N_A_300_74#_c_940_n 0.0235678f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=1.995
cc_170 VPB N_A_300_74#_c_941_n 0.0270943f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_171 VPB N_A_300_74#_c_942_n 0.0100929f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_172 VPB N_A_300_74#_c_943_n 0.0171049f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_173 VPB N_A_300_74#_c_944_n 0.0178649f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_174 VPB N_A_300_74#_c_930_n 0.0209755f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_175 VPB N_A_300_74#_c_931_n 0.00183868f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_176 VPB N_A_300_74#_c_947_n 0.0322371f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_177 VPB N_A_300_74#_c_948_n 0.00523806f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_178 VPB N_A_300_74#_c_933_n 0.00188302f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_179 VPB N_A_300_74#_c_934_n 0.0168815f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_180 VPB N_A_300_74#_c_951_n 0.00232654f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_181 VPB N_A_300_74#_c_952_n 0.0463369f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_182 VPB N_A_300_74#_c_936_n 0.00280482f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_183 VPB N_A_300_74#_c_937_n 0.0167017f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_184 VPB N_A_1598_93#_M1000_g 0.01871f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=0.58
cc_185 VPB N_A_1598_93#_c_1122_n 0.0544767f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_186 VPB N_A_1598_93#_c_1123_n 0.00706063f $X=-0.19 $Y=1.66 $X2=0.352 $Y2=1.11
cc_187 VPB N_A_1598_93#_c_1124_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_188 VPB N_A_1598_93#_c_1125_n 0.00961486f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.95
cc_189 VPB N_A_1598_93#_c_1119_n 0.00471733f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_190 VPB N_A_1598_93#_c_1127_n 0.00400474f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.125
cc_191 VPB N_A_1266_119#_c_1208_n 0.023609f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=0.58
cc_192 VPB N_A_1266_119#_c_1218_n 0.0201446f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_193 VPB N_A_1266_119#_c_1219_n 0.0231244f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.11
cc_194 VPB N_A_1266_119#_c_1220_n 0.059564f $X=-0.19 $Y=1.66 $X2=0.36 $Y2=1.995
cc_195 VPB N_A_1266_119#_c_1221_n 0.0184812f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_196 VPB N_A_1266_119#_c_1222_n 0.00674641f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_197 VPB N_A_1266_119#_c_1213_n 0.0132664f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_198 VPB N_A_1266_119#_c_1224_n 0.00103675f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_199 VPB N_A_1266_119#_c_1215_n 5.52803e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_200 VPB N_A_1934_94#_c_1346_n 0.0302218f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=0.58
cc_201 VPB N_A_1934_94#_c_1352_n 0.00268013f $X=-0.19 $Y=1.66 $X2=0.352 $Y2=0.96
cc_202 VPB N_A_1934_94#_c_1353_n 0.00754272f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_203 VPB N_A_1934_94#_c_1348_n 0.0059282f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_204 VPB N_VPWR_c_1406_n 0.0117486f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_205 VPB N_VPWR_c_1407_n 0.0301196f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.125
cc_206 VPB N_VPWR_c_1408_n 0.0115905f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_207 VPB N_VPWR_c_1409_n 0.0222401f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_208 VPB N_VPWR_c_1410_n 0.0147806f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_209 VPB N_VPWR_c_1411_n 0.0195713f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_210 VPB N_VPWR_c_1412_n 0.0144237f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_211 VPB N_VPWR_c_1413_n 0.00931072f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_212 VPB N_VPWR_c_1414_n 0.0161288f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_213 VPB N_VPWR_c_1415_n 0.00977211f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_214 VPB N_VPWR_c_1416_n 0.0619705f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_215 VPB N_VPWR_c_1417_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_216 VPB N_VPWR_c_1418_n 0.0193312f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_217 VPB N_VPWR_c_1419_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_218 VPB N_VPWR_c_1420_n 0.0160436f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_219 VPB N_VPWR_c_1421_n 0.0201182f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_220 VPB N_VPWR_c_1422_n 0.0599998f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_221 VPB N_VPWR_c_1423_n 0.0209223f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_222 VPB N_VPWR_c_1424_n 0.0197908f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_223 VPB N_VPWR_c_1405_n 0.1054f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_224 VPB N_VPWR_c_1426_n 0.00436868f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_225 VPB N_VPWR_c_1427_n 0.00436868f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_226 VPB N_VPWR_c_1428_n 0.00436868f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_227 VPB N_VPWR_c_1429_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_228 VPB N_VPWR_c_1430_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_229 VPB N_A_33_74#_c_1537_n 0.00638316f $X=-0.19 $Y=1.66 $X2=0.352 $Y2=1.11
cc_230 VPB N_A_33_74#_c_1543_n 0.00584297f $X=-0.19 $Y=1.66 $X2=0.36 $Y2=1.995
cc_231 VPB N_A_33_74#_c_1544_n 0.0143135f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=1.995
cc_232 VPB N_A_33_74#_c_1538_n 2.52696e-19 $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_233 VPB N_A_33_74#_c_1546_n 0.0099755f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.95
cc_234 VPB N_A_33_74#_c_1547_n 0.00810438f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_235 VPB N_A_33_74#_c_1548_n 0.00688265f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_236 VPB Q 0.00930674f $X=-0.19 $Y=1.66 $X2=0.352 $Y2=1.11
cc_237 VPB Q 0.0416636f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.95
cc_238 VPB N_Q_c_1644_n 0.00772285f $X=-0.19 $Y=1.66 $X2=0.237 $Y2=1.295
cc_239 N_D_M1029_g N_RESET_B_M1025_g 0.0435282f $X=0.525 $Y=0.58 $X2=0 $Y2=0
cc_240 N_D_c_244_n N_RESET_B_M1025_g 0.00161151f $X=0.27 $Y=1.125 $X2=0 $Y2=0
cc_241 N_D_c_240_n N_RESET_B_c_606_n 0.00501286f $X=0.36 $Y=1.92 $X2=0 $Y2=0
cc_242 N_D_c_247_n N_RESET_B_c_606_n 0.00699779f $X=0.5 $Y=2.07 $X2=0 $Y2=0
cc_243 N_D_c_248_n N_RESET_B_c_607_n 0.00699779f $X=0.5 $Y=2.375 $X2=0 $Y2=0
cc_244 N_D_c_248_n N_RESET_B_M1024_g 0.00877322f $X=0.5 $Y=2.375 $X2=0 $Y2=0
cc_245 N_D_c_249_n N_RESET_B_M1024_g 0.00816466f $X=0.5 $Y=2.465 $X2=0 $Y2=0
cc_246 N_D_c_244_n N_RESET_B_c_601_n 0.0122082f $X=0.27 $Y=1.125 $X2=0 $Y2=0
cc_247 N_D_c_247_n N_VPWR_c_1407_n 0.00199186f $X=0.5 $Y=2.07 $X2=0 $Y2=0
cc_248 N_D_c_249_n N_VPWR_c_1407_n 0.0120556f $X=0.5 $Y=2.465 $X2=0 $Y2=0
cc_249 N_D_c_245_n N_VPWR_c_1407_n 0.0140568f $X=0.27 $Y=1.125 $X2=0 $Y2=0
cc_250 N_D_c_249_n N_VPWR_c_1420_n 0.00413917f $X=0.5 $Y=2.465 $X2=0 $Y2=0
cc_251 N_D_c_249_n N_VPWR_c_1405_n 0.00853987f $X=0.5 $Y=2.465 $X2=0 $Y2=0
cc_252 N_D_c_247_n N_A_33_74#_c_1537_n 0.00493271f $X=0.5 $Y=2.07 $X2=0 $Y2=0
cc_253 N_D_c_248_n N_A_33_74#_c_1537_n 0.00297569f $X=0.5 $Y=2.375 $X2=0 $Y2=0
cc_254 N_D_M1029_g N_A_33_74#_c_1537_n 0.00857134f $X=0.525 $Y=0.58 $X2=0 $Y2=0
cc_255 N_D_c_242_n N_A_33_74#_c_1537_n 0.00517676f $X=0.352 $Y=1.11 $X2=0 $Y2=0
cc_256 N_D_c_244_n N_A_33_74#_c_1537_n 0.00664601f $X=0.27 $Y=1.125 $X2=0 $Y2=0
cc_257 N_D_c_245_n N_A_33_74#_c_1537_n 0.0866708f $X=0.27 $Y=1.125 $X2=0 $Y2=0
cc_258 N_D_c_248_n N_A_33_74#_c_1543_n 0.0029291f $X=0.5 $Y=2.375 $X2=0 $Y2=0
cc_259 N_D_c_249_n N_A_33_74#_c_1543_n 0.00324529f $X=0.5 $Y=2.465 $X2=0 $Y2=0
cc_260 N_D_M1029_g N_A_33_74#_c_1541_n 0.0152419f $X=0.525 $Y=0.58 $X2=0 $Y2=0
cc_261 N_D_c_242_n N_A_33_74#_c_1541_n 0.0040449f $X=0.352 $Y=1.11 $X2=0 $Y2=0
cc_262 N_D_c_245_n N_A_33_74#_c_1541_n 0.0188861f $X=0.27 $Y=1.125 $X2=0 $Y2=0
cc_263 N_D_c_248_n N_A_33_74#_c_1548_n 0.0128528f $X=0.5 $Y=2.375 $X2=0 $Y2=0
cc_264 N_D_M1029_g N_VGND_c_1675_n 0.00291649f $X=0.525 $Y=0.58 $X2=0 $Y2=0
cc_265 N_D_M1029_g N_VGND_c_1681_n 0.00362587f $X=0.525 $Y=0.58 $X2=0 $Y2=0
cc_266 N_CLK_N_c_280_n N_RESET_B_M1025_g 0.0216977f $X=1.527 $Y=1.185 $X2=0
+ $Y2=0
cc_267 N_CLK_N_c_283_n N_RESET_B_c_606_n 0.0210883f $X=1.527 $Y=1.66 $X2=0 $Y2=0
cc_268 N_CLK_N_c_283_n N_RESET_B_M1024_g 0.0142048f $X=1.527 $Y=1.66 $X2=0 $Y2=0
cc_269 N_CLK_N_c_283_n N_RESET_B_c_609_n 0.0104164f $X=1.527 $Y=1.66 $X2=0 $Y2=0
cc_270 CLK_N N_RESET_B_c_595_n 0.0113341f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_271 N_CLK_N_c_279_n N_RESET_B_c_595_n 0.00659523f $X=1.54 $Y=1.41 $X2=0 $Y2=0
cc_272 N_CLK_N_c_283_n N_RESET_B_c_595_n 0.0033227f $X=1.527 $Y=1.66 $X2=0 $Y2=0
cc_273 CLK_N N_RESET_B_c_596_n 0.00137295f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_274 N_CLK_N_c_279_n N_RESET_B_c_596_n 7.75208e-19 $X=1.54 $Y=1.41 $X2=0 $Y2=0
cc_275 N_CLK_N_c_283_n N_RESET_B_c_596_n 7.78161e-19 $X=1.527 $Y=1.66 $X2=0
+ $Y2=0
cc_276 CLK_N N_RESET_B_c_601_n 6.88904e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_277 N_CLK_N_c_279_n N_RESET_B_c_601_n 0.0301644f $X=1.54 $Y=1.41 $X2=0 $Y2=0
cc_278 CLK_N N_RESET_B_c_602_n 0.0312595f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_279 N_CLK_N_c_279_n N_RESET_B_c_602_n 0.00290042f $X=1.54 $Y=1.41 $X2=0 $Y2=0
cc_280 N_CLK_N_c_283_n N_RESET_B_c_602_n 0.00137593f $X=1.527 $Y=1.66 $X2=0
+ $Y2=0
cc_281 N_CLK_N_c_279_n N_A_300_74#_M1005_g 2.43084e-19 $X=1.54 $Y=1.41 $X2=0
+ $Y2=0
cc_282 CLK_N N_A_300_74#_c_930_n 0.00273214f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_283 N_CLK_N_c_279_n N_A_300_74#_c_930_n 0.0299497f $X=1.54 $Y=1.41 $X2=0
+ $Y2=0
cc_284 CLK_N N_A_300_74#_c_948_n 0.0139359f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_285 N_CLK_N_c_279_n N_A_300_74#_c_948_n 0.00303239f $X=1.54 $Y=1.41 $X2=0
+ $Y2=0
cc_286 N_CLK_N_c_283_n N_A_300_74#_c_948_n 0.00411882f $X=1.527 $Y=1.66 $X2=0
+ $Y2=0
cc_287 CLK_N N_A_300_74#_c_933_n 0.035677f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_288 N_CLK_N_c_279_n N_A_300_74#_c_933_n 6.47976e-19 $X=1.54 $Y=1.41 $X2=0
+ $Y2=0
cc_289 N_CLK_N_c_280_n N_A_300_74#_c_933_n 0.00329654f $X=1.527 $Y=1.185 $X2=0
+ $Y2=0
cc_290 N_CLK_N_c_283_n N_A_300_74#_c_933_n 0.00168547f $X=1.527 $Y=1.66 $X2=0
+ $Y2=0
cc_291 CLK_N N_A_300_74#_c_935_n 0.0224579f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_292 N_CLK_N_c_279_n N_A_300_74#_c_935_n 0.00141168f $X=1.54 $Y=1.41 $X2=0
+ $Y2=0
cc_293 N_CLK_N_c_280_n N_A_300_74#_c_935_n 0.010507f $X=1.527 $Y=1.185 $X2=0
+ $Y2=0
cc_294 N_CLK_N_c_283_n N_VPWR_c_1408_n 0.00506115f $X=1.527 $Y=1.66 $X2=0 $Y2=0
cc_295 N_CLK_N_c_283_n N_VPWR_c_1409_n 0.00869604f $X=1.527 $Y=1.66 $X2=0 $Y2=0
cc_296 N_CLK_N_c_283_n N_VPWR_c_1405_n 9.39239e-19 $X=1.527 $Y=1.66 $X2=0 $Y2=0
cc_297 CLK_N N_A_33_74#_c_1544_n 8.57372e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_298 N_CLK_N_c_283_n N_A_33_74#_c_1544_n 0.0182985f $X=1.527 $Y=1.66 $X2=0
+ $Y2=0
cc_299 N_CLK_N_c_280_n N_VGND_c_1670_n 0.00334184f $X=1.527 $Y=1.185 $X2=0 $Y2=0
cc_300 N_CLK_N_c_280_n N_VGND_c_1671_n 0.00288682f $X=1.527 $Y=1.185 $X2=0 $Y2=0
cc_301 N_CLK_N_c_280_n N_VGND_c_1676_n 0.00433139f $X=1.527 $Y=1.185 $X2=0 $Y2=0
cc_302 N_CLK_N_c_280_n N_VGND_c_1681_n 0.00822407f $X=1.527 $Y=1.185 $X2=0 $Y2=0
cc_303 N_A_507_347#_c_342_n N_A_841_288#_c_506_n 0.00743758f $X=3.92 $Y=2.09
+ $X2=0 $Y2=0
cc_304 N_A_507_347#_c_346_n N_A_841_288#_c_506_n 0.0195543f $X=4.01 $Y=2.165
+ $X2=0 $Y2=0
cc_305 N_A_507_347#_c_327_n N_A_841_288#_M1026_g 0.00338587f $X=3.795 $Y=1.215
+ $X2=0 $Y2=0
cc_306 N_A_507_347#_c_330_n N_A_841_288#_M1026_g 0.00226261f $X=4.685 $Y=0.36
+ $X2=0 $Y2=0
cc_307 N_A_507_347#_c_332_n N_A_841_288#_M1026_g 0.00460805f $X=4.77 $Y=0.79
+ $X2=0 $Y2=0
cc_308 N_A_507_347#_c_354_p N_A_841_288#_M1026_g 0.00240852f $X=4.855 $Y=0.875
+ $X2=0 $Y2=0
cc_309 N_A_507_347#_c_343_n N_A_841_288#_c_507_n 0.0195543f $X=4.01 $Y=2.24
+ $X2=0 $Y2=0
cc_310 N_A_507_347#_c_340_n N_A_841_288#_c_500_n 2.98915e-19 $X=3.92 $Y=1.715
+ $X2=0 $Y2=0
cc_311 N_A_507_347#_c_322_n N_A_841_288#_c_501_n 0.00353124f $X=3.795 $Y=1.55
+ $X2=0 $Y2=0
cc_312 N_A_507_347#_c_340_n N_A_841_288#_c_501_n 0.0215924f $X=3.92 $Y=1.715
+ $X2=0 $Y2=0
cc_313 N_A_507_347#_c_330_n N_A_841_288#_c_502_n 8.56224e-19 $X=4.685 $Y=0.36
+ $X2=0 $Y2=0
cc_314 N_A_507_347#_c_360_p N_A_841_288#_c_502_n 0.0587678f $X=5.525 $Y=0.875
+ $X2=0 $Y2=0
cc_315 N_A_507_347#_c_354_p N_A_841_288#_c_502_n 0.0112104f $X=4.855 $Y=0.875
+ $X2=0 $Y2=0
cc_316 N_A_507_347#_c_330_n N_A_841_288#_c_503_n 0.0117521f $X=4.685 $Y=0.36
+ $X2=0 $Y2=0
cc_317 N_A_507_347#_c_334_n N_A_841_288#_c_504_n 0.0206843f $X=6.365 $Y=0.34
+ $X2=0 $Y2=0
cc_318 N_A_507_347#_c_345_n N_A_841_288#_c_510_n 9.21729e-19 $X=6.81 $Y=1.885
+ $X2=0 $Y2=0
cc_319 N_A_507_347#_c_345_n N_A_841_288#_c_505_n 0.00175018f $X=6.81 $Y=1.885
+ $X2=0 $Y2=0
cc_320 N_A_507_347#_c_343_n N_RESET_B_c_609_n 0.00976827f $X=4.01 $Y=2.24 $X2=0
+ $Y2=0
cc_321 N_A_507_347#_c_360_p N_RESET_B_c_592_n 0.00211559f $X=5.525 $Y=0.875
+ $X2=0 $Y2=0
cc_322 N_A_507_347#_c_332_n N_RESET_B_c_594_n 0.00708744f $X=4.77 $Y=0.79 $X2=0
+ $Y2=0
cc_323 N_A_507_347#_c_360_p N_RESET_B_c_594_n 0.0084462f $X=5.525 $Y=0.875 $X2=0
+ $Y2=0
cc_324 N_A_507_347#_c_354_p N_RESET_B_c_594_n 0.00195216f $X=4.855 $Y=0.875
+ $X2=0 $Y2=0
cc_325 N_A_507_347#_c_333_n N_RESET_B_c_594_n 0.00267306f $X=5.61 $Y=0.79 $X2=0
+ $Y2=0
cc_326 N_A_507_347#_M1017_d N_RESET_B_c_595_n 0.00154568f $X=2.535 $Y=1.735
+ $X2=0 $Y2=0
cc_327 N_A_507_347#_c_328_n N_RESET_B_c_595_n 7.90984e-19 $X=2.76 $Y=0.99 $X2=0
+ $Y2=0
cc_328 N_A_507_347#_c_329_n N_RESET_B_c_595_n 0.0621753f $X=3.62 $Y=1.245 $X2=0
+ $Y2=0
cc_329 N_A_507_347#_c_340_n N_RESET_B_c_595_n 0.00788426f $X=3.92 $Y=1.715 $X2=0
+ $Y2=0
cc_330 N_A_507_347#_c_323_n N_RESET_B_c_597_n 0.00221676f $X=6.81 $Y=1.795 $X2=0
+ $Y2=0
cc_331 N_A_507_347#_c_325_n N_RESET_B_c_597_n 0.00405791f $X=7.6 $Y=1.2 $X2=0
+ $Y2=0
cc_332 N_A_507_347#_c_378_p N_RESET_B_c_597_n 0.00155657f $X=6.535 $Y=1.21 $X2=0
+ $Y2=0
cc_333 N_A_507_347#_c_379_p N_RESET_B_c_597_n 0.0169144f $X=7.08 $Y=1.29 $X2=0
+ $Y2=0
cc_334 N_A_507_347#_c_338_n N_RESET_B_c_597_n 0.011489f $X=7.255 $Y=1.29 $X2=0
+ $Y2=0
cc_335 N_A_507_347#_c_339_n N_RESET_B_c_597_n 0.00501712f $X=6.75 $Y=1.29 $X2=0
+ $Y2=0
cc_336 N_A_507_347#_c_329_n N_A_714_127#_M1013_d 0.00383506f $X=3.62 $Y=1.245
+ $X2=-0.19 $Y2=-0.245
cc_337 N_A_507_347#_c_333_n N_A_714_127#_M1020_g 0.00745398f $X=5.61 $Y=0.79
+ $X2=0 $Y2=0
cc_338 N_A_507_347#_c_334_n N_A_714_127#_M1020_g 0.00330666f $X=6.365 $Y=0.34
+ $X2=0 $Y2=0
cc_339 N_A_507_347#_c_321_n N_A_714_127#_c_825_n 0.00141765f $X=3.495 $Y=1.14
+ $X2=0 $Y2=0
cc_340 N_A_507_347#_c_342_n N_A_714_127#_c_825_n 0.00205943f $X=3.92 $Y=2.09
+ $X2=0 $Y2=0
cc_341 N_A_507_347#_c_327_n N_A_714_127#_c_825_n 0.00513222f $X=3.795 $Y=1.215
+ $X2=0 $Y2=0
cc_342 N_A_507_347#_c_329_n N_A_714_127#_c_825_n 0.101833f $X=3.62 $Y=1.245
+ $X2=0 $Y2=0
cc_343 N_A_507_347#_c_330_n N_A_714_127#_c_825_n 0.0144559f $X=4.685 $Y=0.36
+ $X2=0 $Y2=0
cc_344 N_A_507_347#_c_340_n N_A_714_127#_c_825_n 0.0115203f $X=3.92 $Y=1.715
+ $X2=0 $Y2=0
cc_345 N_A_507_347#_c_346_n N_A_714_127#_c_830_n 0.00109218f $X=4.01 $Y=2.165
+ $X2=0 $Y2=0
cc_346 N_A_507_347#_c_342_n N_A_714_127#_c_831_n 0.00485719f $X=3.92 $Y=2.09
+ $X2=0 $Y2=0
cc_347 N_A_507_347#_c_343_n N_A_714_127#_c_831_n 0.0146858f $X=4.01 $Y=2.24
+ $X2=0 $Y2=0
cc_348 N_A_507_347#_c_346_n N_A_714_127#_c_831_n 0.0108788f $X=4.01 $Y=2.165
+ $X2=0 $Y2=0
cc_349 N_A_507_347#_c_329_n N_A_714_127#_c_831_n 0.0108998f $X=3.62 $Y=1.245
+ $X2=0 $Y2=0
cc_350 N_A_507_347#_c_340_n N_A_714_127#_c_831_n 0.00608099f $X=3.92 $Y=1.715
+ $X2=0 $Y2=0
cc_351 N_A_507_347#_c_329_n N_A_300_74#_c_938_n 0.00301668f $X=3.62 $Y=1.245
+ $X2=0 $Y2=0
cc_352 N_A_507_347#_c_328_n N_A_300_74#_M1005_g 0.00601889f $X=2.76 $Y=0.99
+ $X2=0 $Y2=0
cc_353 N_A_507_347#_c_321_n N_A_300_74#_c_924_n 0.00850225f $X=3.495 $Y=1.14
+ $X2=0 $Y2=0
cc_354 N_A_507_347#_c_330_n N_A_300_74#_c_924_n 0.0072068f $X=4.685 $Y=0.36
+ $X2=0 $Y2=0
cc_355 N_A_507_347#_c_331_n N_A_300_74#_c_924_n 0.00363979f $X=3.705 $Y=0.36
+ $X2=0 $Y2=0
cc_356 N_A_507_347#_c_322_n N_A_300_74#_c_926_n 0.00122112f $X=3.795 $Y=1.55
+ $X2=0 $Y2=0
cc_357 N_A_507_347#_c_327_n N_A_300_74#_c_926_n 0.00486442f $X=3.795 $Y=1.215
+ $X2=0 $Y2=0
cc_358 N_A_507_347#_c_328_n N_A_300_74#_c_926_n 0.00844965f $X=2.76 $Y=0.99
+ $X2=0 $Y2=0
cc_359 N_A_507_347#_c_329_n N_A_300_74#_c_926_n 0.0423425f $X=3.62 $Y=1.245
+ $X2=0 $Y2=0
cc_360 N_A_507_347#_c_340_n N_A_300_74#_c_926_n 0.0214165f $X=3.92 $Y=1.715
+ $X2=0 $Y2=0
cc_361 N_A_507_347#_c_342_n N_A_300_74#_c_940_n 0.00281124f $X=3.92 $Y=2.09
+ $X2=0 $Y2=0
cc_362 N_A_507_347#_c_329_n N_A_300_74#_c_940_n 0.0169164f $X=3.62 $Y=1.245
+ $X2=0 $Y2=0
cc_363 N_A_507_347#_c_346_n N_A_300_74#_c_941_n 0.0101142f $X=4.01 $Y=2.165
+ $X2=0 $Y2=0
cc_364 N_A_507_347#_c_329_n N_A_300_74#_c_941_n 0.0110426f $X=3.62 $Y=1.245
+ $X2=0 $Y2=0
cc_365 N_A_507_347#_c_340_n N_A_300_74#_c_941_n 0.0147787f $X=3.92 $Y=1.715
+ $X2=0 $Y2=0
cc_366 N_A_507_347#_c_343_n N_A_300_74#_c_943_n 0.010856f $X=4.01 $Y=2.24 $X2=0
+ $Y2=0
cc_367 N_A_507_347#_c_321_n N_A_300_74#_M1030_g 0.00726508f $X=3.495 $Y=1.14
+ $X2=0 $Y2=0
cc_368 N_A_507_347#_c_327_n N_A_300_74#_M1030_g 0.00224969f $X=3.795 $Y=1.215
+ $X2=0 $Y2=0
cc_369 N_A_507_347#_c_329_n N_A_300_74#_M1030_g 0.00406678f $X=3.62 $Y=1.245
+ $X2=0 $Y2=0
cc_370 N_A_507_347#_c_330_n N_A_300_74#_M1030_g 0.0206665f $X=4.685 $Y=0.36
+ $X2=0 $Y2=0
cc_371 N_A_507_347#_c_332_n N_A_300_74#_M1030_g 0.00146995f $X=4.77 $Y=0.79
+ $X2=0 $Y2=0
cc_372 N_A_507_347#_c_330_n N_A_300_74#_c_928_n 0.00937668f $X=4.685 $Y=0.36
+ $X2=0 $Y2=0
cc_373 N_A_507_347#_c_360_p N_A_300_74#_c_928_n 0.00549731f $X=5.525 $Y=0.875
+ $X2=0 $Y2=0
cc_374 N_A_507_347#_c_334_n N_A_300_74#_c_928_n 0.00676815f $X=6.365 $Y=0.34
+ $X2=0 $Y2=0
cc_375 N_A_507_347#_c_335_n N_A_300_74#_c_928_n 0.0041995f $X=5.695 $Y=0.34
+ $X2=0 $Y2=0
cc_376 N_A_507_347#_c_324_n N_A_300_74#_M1006_g 0.00954257f $X=6.9 $Y=1.29 $X2=0
+ $Y2=0
cc_377 N_A_507_347#_c_333_n N_A_300_74#_M1006_g 8.97611e-19 $X=5.61 $Y=0.79
+ $X2=0 $Y2=0
cc_378 N_A_507_347#_c_334_n N_A_300_74#_M1006_g 0.0169375f $X=6.365 $Y=0.34
+ $X2=0 $Y2=0
cc_379 N_A_507_347#_c_336_n N_A_300_74#_M1006_g 0.0152469f $X=6.45 $Y=1.125
+ $X2=0 $Y2=0
cc_380 N_A_507_347#_c_379_p N_A_300_74#_M1006_g 8.5704e-19 $X=7.08 $Y=1.29 $X2=0
+ $Y2=0
cc_381 N_A_507_347#_c_345_n N_A_300_74#_c_944_n 0.00540267f $X=6.81 $Y=1.885
+ $X2=0 $Y2=0
cc_382 N_A_507_347#_c_345_n N_A_300_74#_c_947_n 0.00223241f $X=6.81 $Y=1.885
+ $X2=0 $Y2=0
cc_383 N_A_507_347#_c_323_n N_A_300_74#_c_934_n 0.00883406f $X=6.81 $Y=1.795
+ $X2=0 $Y2=0
cc_384 N_A_507_347#_c_345_n N_A_300_74#_c_934_n 0.00783008f $X=6.81 $Y=1.885
+ $X2=0 $Y2=0
cc_385 N_A_507_347#_c_325_n N_A_300_74#_c_934_n 0.00107089f $X=7.6 $Y=1.2 $X2=0
+ $Y2=0
cc_386 N_A_507_347#_c_378_p N_A_300_74#_c_934_n 8.672e-19 $X=6.535 $Y=1.21 $X2=0
+ $Y2=0
cc_387 N_A_507_347#_c_379_p N_A_300_74#_c_934_n 0.0348735f $X=7.08 $Y=1.29 $X2=0
+ $Y2=0
cc_388 N_A_507_347#_c_337_n N_A_300_74#_c_934_n 0.00717074f $X=7.255 $Y=1.29
+ $X2=0 $Y2=0
cc_389 N_A_507_347#_c_338_n N_A_300_74#_c_934_n 0.00892364f $X=7.255 $Y=1.29
+ $X2=0 $Y2=0
cc_390 N_A_507_347#_c_339_n N_A_300_74#_c_934_n 0.00691585f $X=6.75 $Y=1.29
+ $X2=0 $Y2=0
cc_391 N_A_507_347#_c_341_n N_A_300_74#_c_934_n 6.09268e-19 $X=7.42 $Y=1.29
+ $X2=0 $Y2=0
cc_392 N_A_507_347#_c_345_n N_A_300_74#_c_951_n 0.00250118f $X=6.81 $Y=1.885
+ $X2=0 $Y2=0
cc_393 N_A_507_347#_c_323_n N_A_300_74#_c_952_n 0.00562911f $X=6.81 $Y=1.795
+ $X2=0 $Y2=0
cc_394 N_A_507_347#_c_345_n N_A_300_74#_c_952_n 0.0130552f $X=6.81 $Y=1.885
+ $X2=0 $Y2=0
cc_395 N_A_507_347#_c_325_n N_A_300_74#_c_952_n 0.00873909f $X=7.6 $Y=1.2 $X2=0
+ $Y2=0
cc_396 N_A_507_347#_c_341_n N_A_300_74#_c_952_n 0.00582183f $X=7.42 $Y=1.29
+ $X2=0 $Y2=0
cc_397 N_A_507_347#_c_323_n N_A_300_74#_c_936_n 0.00134609f $X=6.81 $Y=1.795
+ $X2=0 $Y2=0
cc_398 N_A_507_347#_c_378_p N_A_300_74#_c_936_n 0.00994746f $X=6.535 $Y=1.21
+ $X2=0 $Y2=0
cc_399 N_A_507_347#_c_323_n N_A_300_74#_c_937_n 0.0215527f $X=6.81 $Y=1.795
+ $X2=0 $Y2=0
cc_400 N_A_507_347#_c_378_p N_A_300_74#_c_937_n 0.00106755f $X=6.535 $Y=1.21
+ $X2=0 $Y2=0
cc_401 N_A_507_347#_c_326_n N_A_1598_93#_M1000_g 0.0413341f $X=7.675 $Y=1.125
+ $X2=0 $Y2=0
cc_402 N_A_507_347#_c_341_n N_A_1598_93#_M1000_g 0.00246675f $X=7.42 $Y=1.29
+ $X2=0 $Y2=0
cc_403 N_A_507_347#_c_336_n N_A_1266_119#_M1006_d 0.0153989f $X=6.45 $Y=1.125
+ $X2=-0.19 $Y2=-0.245
cc_404 N_A_507_347#_c_378_p N_A_1266_119#_M1006_d 0.00269935f $X=6.535 $Y=1.21
+ $X2=-0.19 $Y2=-0.245
cc_405 N_A_507_347#_c_339_n N_A_1266_119#_M1006_d 0.0025788f $X=6.75 $Y=1.29
+ $X2=-0.19 $Y2=-0.245
cc_406 N_A_507_347#_c_324_n N_A_1266_119#_c_1229_n 0.0198469f $X=6.9 $Y=1.29
+ $X2=0 $Y2=0
cc_407 N_A_507_347#_c_326_n N_A_1266_119#_c_1229_n 0.0148493f $X=7.675 $Y=1.125
+ $X2=0 $Y2=0
cc_408 N_A_507_347#_c_336_n N_A_1266_119#_c_1229_n 0.0266855f $X=6.45 $Y=1.125
+ $X2=0 $Y2=0
cc_409 N_A_507_347#_c_339_n N_A_1266_119#_c_1229_n 0.0553581f $X=6.75 $Y=1.29
+ $X2=0 $Y2=0
cc_410 N_A_507_347#_c_345_n N_A_1266_119#_c_1222_n 0.00416251f $X=6.81 $Y=1.885
+ $X2=0 $Y2=0
cc_411 N_A_507_347#_c_326_n N_A_1266_119#_c_1212_n 0.00779099f $X=7.675 $Y=1.125
+ $X2=0 $Y2=0
cc_412 N_A_507_347#_c_337_n N_A_1266_119#_c_1213_n 0.0080525f $X=7.255 $Y=1.29
+ $X2=0 $Y2=0
cc_413 N_A_507_347#_c_341_n N_A_1266_119#_c_1213_n 6.25344e-19 $X=7.42 $Y=1.29
+ $X2=0 $Y2=0
cc_414 N_A_507_347#_c_325_n N_A_1266_119#_c_1237_n 0.00534427f $X=7.6 $Y=1.2
+ $X2=0 $Y2=0
cc_415 N_A_507_347#_c_337_n N_A_1266_119#_c_1237_n 0.00890259f $X=7.255 $Y=1.29
+ $X2=0 $Y2=0
cc_416 N_A_507_347#_c_343_n N_VPWR_c_1410_n 0.00174644f $X=4.01 $Y=2.24 $X2=0
+ $Y2=0
cc_417 N_A_507_347#_c_345_n N_VPWR_c_1416_n 0.00445972f $X=6.81 $Y=1.885 $X2=0
+ $Y2=0
cc_418 N_A_507_347#_c_343_n N_VPWR_c_1405_n 9.39239e-19 $X=4.01 $Y=2.24 $X2=0
+ $Y2=0
cc_419 N_A_507_347#_c_345_n N_VPWR_c_1405_n 0.00863862f $X=6.81 $Y=1.885 $X2=0
+ $Y2=0
cc_420 N_A_507_347#_c_328_n N_A_33_74#_c_1538_n 0.0305218f $X=2.76 $Y=0.99 $X2=0
+ $Y2=0
cc_421 N_A_507_347#_c_329_n N_A_33_74#_c_1538_n 0.0577149f $X=3.62 $Y=1.245
+ $X2=0 $Y2=0
cc_422 N_A_507_347#_M1017_d N_A_33_74#_c_1546_n 0.0170633f $X=2.535 $Y=1.735
+ $X2=0 $Y2=0
cc_423 N_A_507_347#_c_329_n N_A_33_74#_c_1546_n 0.0590222f $X=3.62 $Y=1.245
+ $X2=0 $Y2=0
cc_424 N_A_507_347#_M1005_d N_A_33_74#_c_1539_n 0.00768358f $X=2.55 $Y=0.395
+ $X2=0 $Y2=0
cc_425 N_A_507_347#_c_321_n N_A_33_74#_c_1539_n 0.00337435f $X=3.495 $Y=1.14
+ $X2=0 $Y2=0
cc_426 N_A_507_347#_c_328_n N_A_33_74#_c_1539_n 0.0201664f $X=2.76 $Y=0.99 $X2=0
+ $Y2=0
cc_427 N_A_507_347#_c_329_n N_A_33_74#_c_1539_n 0.018223f $X=3.62 $Y=1.245 $X2=0
+ $Y2=0
cc_428 N_A_507_347#_c_321_n N_A_33_74#_c_1540_n 6.3235e-19 $X=3.495 $Y=1.14
+ $X2=0 $Y2=0
cc_429 N_A_507_347#_c_328_n N_A_33_74#_c_1540_n 0.0196428f $X=2.76 $Y=0.99 $X2=0
+ $Y2=0
cc_430 N_A_507_347#_c_329_n N_A_33_74#_c_1540_n 0.0368142f $X=3.62 $Y=1.245
+ $X2=0 $Y2=0
cc_431 N_A_507_347#_c_360_p N_VGND_M1016_d 0.0157496f $X=5.525 $Y=0.875 $X2=0
+ $Y2=0
cc_432 N_A_507_347#_c_333_n N_VGND_M1016_d 0.00476888f $X=5.61 $Y=0.79 $X2=0
+ $Y2=0
cc_433 N_A_507_347#_c_330_n N_VGND_c_1672_n 0.0185769f $X=4.685 $Y=0.36 $X2=0
+ $Y2=0
cc_434 N_A_507_347#_c_332_n N_VGND_c_1672_n 0.0118158f $X=4.77 $Y=0.79 $X2=0
+ $Y2=0
cc_435 N_A_507_347#_c_360_p N_VGND_c_1672_n 0.0260579f $X=5.525 $Y=0.875 $X2=0
+ $Y2=0
cc_436 N_A_507_347#_c_333_n N_VGND_c_1672_n 0.0153511f $X=5.61 $Y=0.79 $X2=0
+ $Y2=0
cc_437 N_A_507_347#_c_335_n N_VGND_c_1672_n 0.0150385f $X=5.695 $Y=0.34 $X2=0
+ $Y2=0
cc_438 N_A_507_347#_c_326_n N_VGND_c_1673_n 0.00102171f $X=7.675 $Y=1.125 $X2=0
+ $Y2=0
cc_439 N_A_507_347#_c_330_n N_VGND_c_1677_n 0.0751579f $X=4.685 $Y=0.36 $X2=0
+ $Y2=0
cc_440 N_A_507_347#_c_331_n N_VGND_c_1677_n 0.0115893f $X=3.705 $Y=0.36 $X2=0
+ $Y2=0
cc_441 N_A_507_347#_c_326_n N_VGND_c_1678_n 0.00332223f $X=7.675 $Y=1.125 $X2=0
+ $Y2=0
cc_442 N_A_507_347#_c_334_n N_VGND_c_1678_n 0.0548435f $X=6.365 $Y=0.34 $X2=0
+ $Y2=0
cc_443 N_A_507_347#_c_335_n N_VGND_c_1678_n 0.0116199f $X=5.695 $Y=0.34 $X2=0
+ $Y2=0
cc_444 N_A_507_347#_c_321_n N_VGND_c_1681_n 7.33403e-19 $X=3.495 $Y=1.14 $X2=0
+ $Y2=0
cc_445 N_A_507_347#_c_326_n N_VGND_c_1681_n 0.00477801f $X=7.675 $Y=1.125 $X2=0
+ $Y2=0
cc_446 N_A_507_347#_c_330_n N_VGND_c_1681_n 0.0387929f $X=4.685 $Y=0.36 $X2=0
+ $Y2=0
cc_447 N_A_507_347#_c_331_n N_VGND_c_1681_n 0.00583135f $X=3.705 $Y=0.36 $X2=0
+ $Y2=0
cc_448 N_A_507_347#_c_360_p N_VGND_c_1681_n 0.011753f $X=5.525 $Y=0.875 $X2=0
+ $Y2=0
cc_449 N_A_507_347#_c_334_n N_VGND_c_1681_n 0.0291469f $X=6.365 $Y=0.34 $X2=0
+ $Y2=0
cc_450 N_A_507_347#_c_335_n N_VGND_c_1681_n 0.00583764f $X=5.695 $Y=0.34 $X2=0
+ $Y2=0
cc_451 N_A_507_347#_c_332_n A_922_127# 0.00212931f $X=4.77 $Y=0.79 $X2=-0.19
+ $Y2=-0.245
cc_452 N_A_507_347#_c_354_p A_922_127# 0.00332183f $X=4.855 $Y=0.875 $X2=-0.19
+ $Y2=-0.245
cc_453 N_A_841_288#_c_507_n N_RESET_B_c_609_n 0.0103562f $X=4.467 $Y=2.24 $X2=0
+ $Y2=0
cc_454 N_A_841_288#_c_501_n N_RESET_B_c_592_n 0.0276001f $X=4.37 $Y=1.61 $X2=0
+ $Y2=0
cc_455 N_A_841_288#_c_502_n N_RESET_B_c_592_n 0.00845009f $X=5.865 $Y=1.215
+ $X2=0 $Y2=0
cc_456 N_A_841_288#_c_507_n N_RESET_B_c_611_n 0.0276001f $X=4.467 $Y=2.24 $X2=0
+ $Y2=0
cc_457 N_A_841_288#_c_507_n N_RESET_B_M1009_g 0.00779205f $X=4.467 $Y=2.24 $X2=0
+ $Y2=0
cc_458 N_A_841_288#_M1026_g N_RESET_B_c_594_n 0.0276001f $X=4.535 $Y=0.845 $X2=0
+ $Y2=0
cc_459 N_A_841_288#_c_500_n N_RESET_B_c_595_n 0.0318831f $X=4.37 $Y=1.61 $X2=0
+ $Y2=0
cc_460 N_A_841_288#_c_501_n N_RESET_B_c_595_n 0.00297425f $X=4.37 $Y=1.61 $X2=0
+ $Y2=0
cc_461 N_A_841_288#_c_502_n N_RESET_B_c_595_n 0.00550332f $X=5.865 $Y=1.215
+ $X2=0 $Y2=0
cc_462 N_A_841_288#_c_502_n N_RESET_B_c_597_n 0.0118991f $X=5.865 $Y=1.215 $X2=0
+ $Y2=0
cc_463 N_A_841_288#_c_539_p N_RESET_B_c_597_n 0.00468242f $X=6.03 $Y=1.215 $X2=0
+ $Y2=0
cc_464 N_A_841_288#_c_540_p N_RESET_B_c_597_n 0.00919057f $X=6.11 $Y=2.135 $X2=0
+ $Y2=0
cc_465 N_A_841_288#_c_505_n N_RESET_B_c_597_n 0.0226321f $X=6.282 $Y=1.97 $X2=0
+ $Y2=0
cc_466 N_A_841_288#_c_500_n N_RESET_B_c_598_n 6.10351e-19 $X=4.37 $Y=1.61 $X2=0
+ $Y2=0
cc_467 N_A_841_288#_c_502_n N_RESET_B_c_598_n 0.00242896f $X=5.865 $Y=1.215
+ $X2=0 $Y2=0
cc_468 N_A_841_288#_c_506_n N_RESET_B_c_603_n 0.0276001f $X=4.467 $Y=2.098 $X2=0
+ $Y2=0
cc_469 N_A_841_288#_c_502_n N_RESET_B_c_603_n 0.0025155f $X=5.865 $Y=1.215 $X2=0
+ $Y2=0
cc_470 N_A_841_288#_c_500_n N_RESET_B_c_682_n 0.0190798f $X=4.37 $Y=1.61 $X2=0
+ $Y2=0
cc_471 N_A_841_288#_c_501_n N_RESET_B_c_682_n 5.77947e-19 $X=4.37 $Y=1.61 $X2=0
+ $Y2=0
cc_472 N_A_841_288#_c_502_n N_RESET_B_c_682_n 0.0201627f $X=5.865 $Y=1.215 $X2=0
+ $Y2=0
cc_473 N_A_841_288#_c_500_n N_RESET_B_c_604_n 0.00571075f $X=4.37 $Y=1.61 $X2=0
+ $Y2=0
cc_474 N_A_841_288#_c_502_n N_RESET_B_c_604_n 0.00623435f $X=5.865 $Y=1.215
+ $X2=0 $Y2=0
cc_475 N_A_841_288#_c_502_n N_A_714_127#_M1020_g 0.0128664f $X=5.865 $Y=1.215
+ $X2=0 $Y2=0
cc_476 N_A_841_288#_c_504_n N_A_714_127#_M1020_g 0.011387f $X=6.03 $Y=0.76 $X2=0
+ $Y2=0
cc_477 N_A_841_288#_c_539_p N_A_714_127#_M1020_g 3.84191e-19 $X=6.03 $Y=1.215
+ $X2=0 $Y2=0
cc_478 N_A_841_288#_c_505_n N_A_714_127#_M1020_g 0.00824116f $X=6.282 $Y=1.97
+ $X2=0 $Y2=0
cc_479 N_A_841_288#_c_510_n N_A_714_127#_c_823_n 4.6813e-19 $X=6.11 $Y=2.815
+ $X2=0 $Y2=0
cc_480 N_A_841_288#_c_540_p N_A_714_127#_c_823_n 0.00709683f $X=6.11 $Y=2.135
+ $X2=0 $Y2=0
cc_481 N_A_841_288#_c_505_n N_A_714_127#_c_823_n 0.0157335f $X=6.282 $Y=1.97
+ $X2=0 $Y2=0
cc_482 N_A_841_288#_c_502_n N_A_714_127#_c_824_n 0.00222478f $X=5.865 $Y=1.215
+ $X2=0 $Y2=0
cc_483 N_A_841_288#_c_506_n N_A_714_127#_c_825_n 0.00181217f $X=4.467 $Y=2.098
+ $X2=0 $Y2=0
cc_484 N_A_841_288#_M1026_g N_A_714_127#_c_825_n 7.05398e-19 $X=4.535 $Y=0.845
+ $X2=0 $Y2=0
cc_485 N_A_841_288#_c_500_n N_A_714_127#_c_825_n 0.0314133f $X=4.37 $Y=1.61
+ $X2=0 $Y2=0
cc_486 N_A_841_288#_c_501_n N_A_714_127#_c_825_n 0.00445995f $X=4.37 $Y=1.61
+ $X2=0 $Y2=0
cc_487 N_A_841_288#_c_503_n N_A_714_127#_c_825_n 0.0129398f $X=4.655 $Y=1.215
+ $X2=0 $Y2=0
cc_488 N_A_841_288#_c_506_n N_A_714_127#_c_830_n 0.0102406f $X=4.467 $Y=2.098
+ $X2=0 $Y2=0
cc_489 N_A_841_288#_c_507_n N_A_714_127#_c_830_n 0.00915247f $X=4.467 $Y=2.24
+ $X2=0 $Y2=0
cc_490 N_A_841_288#_c_500_n N_A_714_127#_c_830_n 0.0237981f $X=4.37 $Y=1.61
+ $X2=0 $Y2=0
cc_491 N_A_841_288#_c_501_n N_A_714_127#_c_830_n 0.00431321f $X=4.37 $Y=1.61
+ $X2=0 $Y2=0
cc_492 N_A_841_288#_c_502_n N_A_714_127#_c_830_n 0.00409967f $X=5.865 $Y=1.215
+ $X2=0 $Y2=0
cc_493 N_A_841_288#_c_507_n N_A_714_127#_c_831_n 0.0025681f $X=4.467 $Y=2.24
+ $X2=0 $Y2=0
cc_494 N_A_841_288#_c_507_n N_A_714_127#_c_832_n 5.05233e-19 $X=4.467 $Y=2.24
+ $X2=0 $Y2=0
cc_495 N_A_841_288#_c_540_p N_A_714_127#_c_833_n 0.0146166f $X=6.11 $Y=2.135
+ $X2=0 $Y2=0
cc_496 N_A_841_288#_c_502_n N_A_714_127#_c_826_n 0.0256509f $X=5.865 $Y=1.215
+ $X2=0 $Y2=0
cc_497 N_A_841_288#_c_505_n N_A_714_127#_c_826_n 0.0360167f $X=6.282 $Y=1.97
+ $X2=0 $Y2=0
cc_498 N_A_841_288#_M1026_g N_A_300_74#_M1030_g 0.0406821f $X=4.535 $Y=0.845
+ $X2=0 $Y2=0
cc_499 N_A_841_288#_c_501_n N_A_300_74#_M1030_g 0.00294835f $X=4.37 $Y=1.61
+ $X2=0 $Y2=0
cc_500 N_A_841_288#_c_503_n N_A_300_74#_M1030_g 4.53579e-19 $X=4.655 $Y=1.215
+ $X2=0 $Y2=0
cc_501 N_A_841_288#_M1026_g N_A_300_74#_c_928_n 0.00695615f $X=4.535 $Y=0.845
+ $X2=0 $Y2=0
cc_502 N_A_841_288#_c_504_n N_A_300_74#_M1006_g 0.00547135f $X=6.03 $Y=0.76
+ $X2=0 $Y2=0
cc_503 N_A_841_288#_c_539_p N_A_300_74#_M1006_g 0.00198105f $X=6.03 $Y=1.215
+ $X2=0 $Y2=0
cc_504 N_A_841_288#_c_505_n N_A_300_74#_M1006_g 0.00421803f $X=6.282 $Y=1.97
+ $X2=0 $Y2=0
cc_505 N_A_841_288#_c_540_p N_A_300_74#_c_934_n 0.013462f $X=6.11 $Y=2.135 $X2=0
+ $Y2=0
cc_506 N_A_841_288#_c_540_p N_A_300_74#_c_936_n 0.0229541f $X=6.11 $Y=2.135
+ $X2=0 $Y2=0
cc_507 N_A_841_288#_c_505_n N_A_300_74#_c_936_n 0.0236964f $X=6.282 $Y=1.97
+ $X2=0 $Y2=0
cc_508 N_A_841_288#_c_540_p N_A_300_74#_c_937_n 0.00343033f $X=6.11 $Y=2.135
+ $X2=0 $Y2=0
cc_509 N_A_841_288#_c_507_n N_VPWR_c_1410_n 0.0146807f $X=4.467 $Y=2.24 $X2=0
+ $Y2=0
cc_510 N_A_841_288#_c_510_n N_VPWR_c_1412_n 0.0241513f $X=6.11 $Y=2.815 $X2=0
+ $Y2=0
cc_511 N_A_841_288#_c_510_n N_VPWR_c_1416_n 0.0315916f $X=6.11 $Y=2.815 $X2=0
+ $Y2=0
cc_512 N_A_841_288#_c_507_n N_VPWR_c_1405_n 8.51577e-19 $X=4.467 $Y=2.24 $X2=0
+ $Y2=0
cc_513 N_A_841_288#_c_510_n N_VPWR_c_1405_n 0.0261488f $X=6.11 $Y=2.815 $X2=0
+ $Y2=0
cc_514 N_A_841_288#_c_502_n N_VGND_M1016_d 0.00417413f $X=5.865 $Y=1.215 $X2=0
+ $Y2=0
cc_515 N_RESET_B_c_592_n N_A_714_127#_M1020_g 0.0056249f $X=4.937 $Y=1.247 $X2=0
+ $Y2=0
cc_516 N_RESET_B_c_597_n N_A_714_127#_c_823_n 0.00611789f $X=8.255 $Y=1.665
+ $X2=0 $Y2=0
cc_517 N_RESET_B_c_597_n N_A_714_127#_c_824_n 0.00200601f $X=8.255 $Y=1.665
+ $X2=0 $Y2=0
cc_518 N_RESET_B_c_603_n N_A_714_127#_c_824_n 0.0219651f $X=5 $Y=1.635 $X2=0
+ $Y2=0
cc_519 N_RESET_B_c_682_n N_A_714_127#_c_824_n 5.06483e-19 $X=5 $Y=1.635 $X2=0
+ $Y2=0
cc_520 N_RESET_B_c_595_n N_A_714_127#_c_825_n 0.0251047f $X=4.895 $Y=1.665 $X2=0
+ $Y2=0
cc_521 N_RESET_B_c_611_n N_A_714_127#_c_830_n 0.00589641f $X=4.937 $Y=2.123
+ $X2=0 $Y2=0
cc_522 N_RESET_B_c_615_n N_A_714_127#_c_830_n 0.00695901f $X=4.937 $Y=2.24 $X2=0
+ $Y2=0
cc_523 N_RESET_B_c_595_n N_A_714_127#_c_830_n 0.0167174f $X=4.895 $Y=1.665 $X2=0
+ $Y2=0
cc_524 N_RESET_B_c_598_n N_A_714_127#_c_830_n 0.00180322f $X=5.185 $Y=1.665
+ $X2=0 $Y2=0
cc_525 N_RESET_B_c_682_n N_A_714_127#_c_830_n 0.01988f $X=5 $Y=1.635 $X2=0 $Y2=0
cc_526 N_RESET_B_c_609_n N_A_714_127#_c_831_n 0.00569293f $X=4.82 $Y=3.15 $X2=0
+ $Y2=0
cc_527 N_RESET_B_c_595_n N_A_714_127#_c_831_n 0.0064065f $X=4.895 $Y=1.665 $X2=0
+ $Y2=0
cc_528 N_RESET_B_M1009_g N_A_714_127#_c_832_n 0.00403916f $X=4.895 $Y=2.525
+ $X2=0 $Y2=0
cc_529 N_RESET_B_c_615_n N_A_714_127#_c_832_n 0.0064209f $X=4.937 $Y=2.24 $X2=0
+ $Y2=0
cc_530 N_RESET_B_c_611_n N_A_714_127#_c_833_n 0.00587984f $X=4.937 $Y=2.123
+ $X2=0 $Y2=0
cc_531 N_RESET_B_c_615_n N_A_714_127#_c_833_n 7.68935e-19 $X=4.937 $Y=2.24 $X2=0
+ $Y2=0
cc_532 N_RESET_B_c_597_n N_A_714_127#_c_833_n 0.00584063f $X=8.255 $Y=1.665
+ $X2=0 $Y2=0
cc_533 N_RESET_B_c_598_n N_A_714_127#_c_833_n 9.59006e-19 $X=5.185 $Y=1.665
+ $X2=0 $Y2=0
cc_534 N_RESET_B_c_603_n N_A_714_127#_c_833_n 0.0025155f $X=5 $Y=1.635 $X2=0
+ $Y2=0
cc_535 N_RESET_B_c_611_n N_A_714_127#_c_826_n 0.00592612f $X=4.937 $Y=2.123
+ $X2=0 $Y2=0
cc_536 N_RESET_B_c_597_n N_A_714_127#_c_826_n 0.017441f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_537 N_RESET_B_c_598_n N_A_714_127#_c_826_n 0.00269227f $X=5.185 $Y=1.665
+ $X2=0 $Y2=0
cc_538 N_RESET_B_c_603_n N_A_714_127#_c_826_n 0.00166642f $X=5 $Y=1.635 $X2=0
+ $Y2=0
cc_539 N_RESET_B_c_682_n N_A_714_127#_c_826_n 0.0222275f $X=5 $Y=1.635 $X2=0
+ $Y2=0
cc_540 N_RESET_B_c_595_n N_A_300_74#_M1007_d 0.00212136f $X=4.895 $Y=1.665 $X2=0
+ $Y2=0
cc_541 N_RESET_B_c_609_n N_A_300_74#_c_938_n 0.0103562f $X=4.82 $Y=3.15 $X2=0
+ $Y2=0
cc_542 N_RESET_B_c_595_n N_A_300_74#_c_938_n 0.0010986f $X=4.895 $Y=1.665 $X2=0
+ $Y2=0
cc_543 N_RESET_B_c_595_n N_A_300_74#_c_926_n 0.00503591f $X=4.895 $Y=1.665 $X2=0
+ $Y2=0
cc_544 N_RESET_B_c_609_n N_A_300_74#_c_943_n 0.0103469f $X=4.82 $Y=3.15 $X2=0
+ $Y2=0
cc_545 N_RESET_B_c_595_n N_A_300_74#_M1030_g 0.00277153f $X=4.895 $Y=1.665 $X2=0
+ $Y2=0
cc_546 N_RESET_B_c_594_n N_A_300_74#_c_928_n 0.00809285f $X=4.937 $Y=1.13 $X2=0
+ $Y2=0
cc_547 N_RESET_B_c_595_n N_A_300_74#_c_930_n 0.00870077f $X=4.895 $Y=1.665 $X2=0
+ $Y2=0
cc_548 N_RESET_B_c_595_n N_A_300_74#_c_931_n 0.00189004f $X=4.895 $Y=1.665 $X2=0
+ $Y2=0
cc_549 N_RESET_B_c_597_n N_A_300_74#_c_947_n 2.3419e-19 $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_550 N_RESET_B_c_606_n N_A_300_74#_c_948_n 8.89268e-19 $X=0.95 $Y=2.15 $X2=0
+ $Y2=0
cc_551 N_RESET_B_c_595_n N_A_300_74#_c_948_n 0.0153372f $X=4.895 $Y=1.665 $X2=0
+ $Y2=0
cc_552 N_RESET_B_c_595_n N_A_300_74#_c_933_n 0.02346f $X=4.895 $Y=1.665 $X2=0
+ $Y2=0
cc_553 N_RESET_B_c_596_n N_A_300_74#_c_933_n 0.00100473f $X=1.345 $Y=1.665 $X2=0
+ $Y2=0
cc_554 N_RESET_B_c_602_n N_A_300_74#_c_933_n 0.00195266f $X=0.975 $Y=1.41 $X2=0
+ $Y2=0
cc_555 N_RESET_B_c_597_n N_A_300_74#_c_934_n 0.0603286f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_556 N_RESET_B_c_597_n N_A_300_74#_c_952_n 0.00727375f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_557 N_RESET_B_M1025_g N_A_300_74#_c_935_n 0.00104425f $X=0.915 $Y=0.58 $X2=0
+ $Y2=0
cc_558 N_RESET_B_c_595_n N_A_300_74#_c_935_n 0.00676127f $X=4.895 $Y=1.665 $X2=0
+ $Y2=0
cc_559 N_RESET_B_c_597_n N_A_300_74#_c_936_n 0.0194318f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_560 N_RESET_B_c_597_n N_A_300_74#_c_937_n 0.00169661f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_561 N_RESET_B_M1010_g N_A_1598_93#_M1000_g 0.0206165f $X=8.605 $Y=0.805 $X2=0
+ $Y2=0
cc_562 N_RESET_B_c_613_n N_A_1598_93#_M1000_g 0.0068596f $X=8.62 $Y=2.375 $X2=0
+ $Y2=0
cc_563 N_RESET_B_c_597_n N_A_1598_93#_M1000_g 0.00903792f $X=8.255 $Y=1.665
+ $X2=0 $Y2=0
cc_564 N_RESET_B_c_599_n N_A_1598_93#_M1000_g 0.00140024f $X=8.4 $Y=1.665 $X2=0
+ $Y2=0
cc_565 N_RESET_B_c_600_n N_A_1598_93#_M1000_g 0.00248623f $X=8.4 $Y=1.665 $X2=0
+ $Y2=0
cc_566 N_RESET_B_c_605_n N_A_1598_93#_M1000_g 0.0174849f $X=8.545 $Y=1.63 $X2=0
+ $Y2=0
cc_567 N_RESET_B_c_613_n N_A_1598_93#_c_1122_n 0.0255241f $X=8.62 $Y=2.375 $X2=0
+ $Y2=0
cc_568 N_RESET_B_c_614_n N_A_1598_93#_c_1122_n 0.0102544f $X=8.62 $Y=2.465 $X2=0
+ $Y2=0
cc_569 N_RESET_B_c_600_n N_A_1598_93#_c_1122_n 2.32727e-19 $X=8.4 $Y=1.665 $X2=0
+ $Y2=0
cc_570 N_RESET_B_c_613_n N_A_1598_93#_c_1123_n 0.0179198f $X=8.62 $Y=2.375 $X2=0
+ $Y2=0
cc_571 N_RESET_B_c_597_n N_A_1598_93#_c_1123_n 0.00534563f $X=8.255 $Y=1.665
+ $X2=0 $Y2=0
cc_572 N_RESET_B_c_599_n N_A_1598_93#_c_1123_n 0.00307024f $X=8.4 $Y=1.665 $X2=0
+ $Y2=0
cc_573 N_RESET_B_c_600_n N_A_1598_93#_c_1123_n 0.0292669f $X=8.4 $Y=1.665 $X2=0
+ $Y2=0
cc_574 N_RESET_B_c_605_n N_A_1598_93#_c_1123_n 0.00342754f $X=8.545 $Y=1.63
+ $X2=0 $Y2=0
cc_575 N_RESET_B_c_613_n N_A_1598_93#_c_1124_n 0.00121111f $X=8.62 $Y=2.375
+ $X2=0 $Y2=0
cc_576 N_RESET_B_c_614_n N_A_1598_93#_c_1124_n 0.0107743f $X=8.62 $Y=2.465 $X2=0
+ $Y2=0
cc_577 N_RESET_B_c_613_n N_A_1598_93#_c_1119_n 2.15799e-19 $X=8.62 $Y=2.375
+ $X2=0 $Y2=0
cc_578 N_RESET_B_c_605_n N_A_1598_93#_c_1119_n 0.00106075f $X=8.545 $Y=1.63
+ $X2=0 $Y2=0
cc_579 N_RESET_B_c_613_n N_A_1598_93#_c_1127_n 0.00567658f $X=8.62 $Y=2.375
+ $X2=0 $Y2=0
cc_580 N_RESET_B_c_600_n N_A_1598_93#_c_1127_n 0.00239474f $X=8.4 $Y=1.665 $X2=0
+ $Y2=0
cc_581 N_RESET_B_M1010_g N_A_1598_93#_c_1120_n 0.00117144f $X=8.605 $Y=0.805
+ $X2=0 $Y2=0
cc_582 N_RESET_B_M1010_g N_A_1266_119#_c_1207_n 0.0535388f $X=8.605 $Y=0.805
+ $X2=0 $Y2=0
cc_583 N_RESET_B_c_613_n N_A_1266_119#_c_1208_n 0.0166298f $X=8.62 $Y=2.375
+ $X2=0 $Y2=0
cc_584 N_RESET_B_c_614_n N_A_1266_119#_c_1218_n 0.0166298f $X=8.62 $Y=2.465
+ $X2=0 $Y2=0
cc_585 N_RESET_B_c_614_n N_A_1266_119#_c_1219_n 0.00943438f $X=8.62 $Y=2.465
+ $X2=0 $Y2=0
cc_586 N_RESET_B_c_597_n N_A_1266_119#_c_1213_n 0.0247374f $X=8.255 $Y=1.665
+ $X2=0 $Y2=0
cc_587 N_RESET_B_c_599_n N_A_1266_119#_c_1213_n 0.00232289f $X=8.4 $Y=1.665
+ $X2=0 $Y2=0
cc_588 N_RESET_B_c_600_n N_A_1266_119#_c_1213_n 0.0115131f $X=8.4 $Y=1.665 $X2=0
+ $Y2=0
cc_589 N_RESET_B_M1010_g N_A_1266_119#_c_1214_n 0.0144298f $X=8.605 $Y=0.805
+ $X2=0 $Y2=0
cc_590 N_RESET_B_c_597_n N_A_1266_119#_c_1214_n 0.0108617f $X=8.255 $Y=1.665
+ $X2=0 $Y2=0
cc_591 N_RESET_B_c_599_n N_A_1266_119#_c_1214_n 0.0025054f $X=8.4 $Y=1.665 $X2=0
+ $Y2=0
cc_592 N_RESET_B_c_600_n N_A_1266_119#_c_1214_n 0.0302597f $X=8.4 $Y=1.665 $X2=0
+ $Y2=0
cc_593 N_RESET_B_c_605_n N_A_1266_119#_c_1214_n 0.0041539f $X=8.545 $Y=1.63
+ $X2=0 $Y2=0
cc_594 N_RESET_B_M1010_g N_A_1266_119#_c_1215_n 0.00109666f $X=8.605 $Y=0.805
+ $X2=0 $Y2=0
cc_595 N_RESET_B_c_599_n N_A_1266_119#_c_1215_n 0.00111187f $X=8.4 $Y=1.665
+ $X2=0 $Y2=0
cc_596 N_RESET_B_c_600_n N_A_1266_119#_c_1215_n 0.0199249f $X=8.4 $Y=1.665 $X2=0
+ $Y2=0
cc_597 N_RESET_B_c_605_n N_A_1266_119#_c_1215_n 4.14158e-19 $X=8.545 $Y=1.63
+ $X2=0 $Y2=0
cc_598 N_RESET_B_c_600_n N_A_1266_119#_c_1216_n 0.0011399f $X=8.4 $Y=1.665 $X2=0
+ $Y2=0
cc_599 N_RESET_B_c_605_n N_A_1266_119#_c_1216_n 0.0207482f $X=8.545 $Y=1.63
+ $X2=0 $Y2=0
cc_600 N_RESET_B_c_595_n N_VPWR_M1024_d 3.75379e-19 $X=4.895 $Y=1.665 $X2=0
+ $Y2=0
cc_601 N_RESET_B_c_596_n N_VPWR_M1024_d 0.0031457f $X=1.345 $Y=1.665 $X2=0 $Y2=0
cc_602 N_RESET_B_c_602_n N_VPWR_M1024_d 0.0022453f $X=0.975 $Y=1.41 $X2=0 $Y2=0
cc_603 N_RESET_B_c_595_n N_VPWR_M1017_s 0.0018769f $X=4.895 $Y=1.665 $X2=0 $Y2=0
cc_604 N_RESET_B_M1024_g N_VPWR_c_1407_n 4.78696e-19 $X=0.95 $Y=2.75 $X2=0 $Y2=0
cc_605 N_RESET_B_c_610_n N_VPWR_c_1407_n 0.00177402f $X=1.025 $Y=3.15 $X2=0
+ $Y2=0
cc_606 N_RESET_B_M1024_g N_VPWR_c_1408_n 0.00510234f $X=0.95 $Y=2.75 $X2=0 $Y2=0
cc_607 N_RESET_B_c_609_n N_VPWR_c_1408_n 0.0222198f $X=4.82 $Y=3.15 $X2=0 $Y2=0
cc_608 N_RESET_B_c_609_n N_VPWR_c_1409_n 0.0255937f $X=4.82 $Y=3.15 $X2=0 $Y2=0
cc_609 N_RESET_B_c_609_n N_VPWR_c_1410_n 0.0239371f $X=4.82 $Y=3.15 $X2=0 $Y2=0
cc_610 N_RESET_B_M1009_g N_VPWR_c_1410_n 0.0130384f $X=4.895 $Y=2.525 $X2=0
+ $Y2=0
cc_611 N_RESET_B_c_609_n N_VPWR_c_1411_n 0.00698559f $X=4.82 $Y=3.15 $X2=0 $Y2=0
cc_612 N_RESET_B_M1009_g N_VPWR_c_1412_n 0.0119399f $X=4.895 $Y=2.525 $X2=0
+ $Y2=0
cc_613 N_RESET_B_c_614_n N_VPWR_c_1413_n 0.00722976f $X=8.62 $Y=2.465 $X2=0
+ $Y2=0
cc_614 N_RESET_B_c_610_n N_VPWR_c_1420_n 0.0064002f $X=1.025 $Y=3.15 $X2=0 $Y2=0
cc_615 N_RESET_B_c_609_n N_VPWR_c_1421_n 0.0246736f $X=4.82 $Y=3.15 $X2=0 $Y2=0
cc_616 N_RESET_B_c_609_n N_VPWR_c_1422_n 0.0648783f $X=4.82 $Y=3.15 $X2=0 $Y2=0
cc_617 N_RESET_B_c_614_n N_VPWR_c_1423_n 0.00445602f $X=8.62 $Y=2.465 $X2=0
+ $Y2=0
cc_618 N_RESET_B_c_609_n N_VPWR_c_1405_n 0.13137f $X=4.82 $Y=3.15 $X2=0 $Y2=0
cc_619 N_RESET_B_c_610_n N_VPWR_c_1405_n 0.011325f $X=1.025 $Y=3.15 $X2=0 $Y2=0
cc_620 N_RESET_B_c_614_n N_VPWR_c_1405_n 0.00896557f $X=8.62 $Y=2.465 $X2=0
+ $Y2=0
cc_621 N_RESET_B_M1025_g N_A_33_74#_c_1537_n 0.00825329f $X=0.915 $Y=0.58 $X2=0
+ $Y2=0
cc_622 N_RESET_B_c_606_n N_A_33_74#_c_1537_n 0.00959854f $X=0.95 $Y=2.15 $X2=0
+ $Y2=0
cc_623 N_RESET_B_c_596_n N_A_33_74#_c_1537_n 0.00112473f $X=1.345 $Y=1.665 $X2=0
+ $Y2=0
cc_624 N_RESET_B_c_601_n N_A_33_74#_c_1537_n 0.00498535f $X=0.975 $Y=1.41 $X2=0
+ $Y2=0
cc_625 N_RESET_B_c_602_n N_A_33_74#_c_1537_n 0.0397689f $X=0.975 $Y=1.41 $X2=0
+ $Y2=0
cc_626 N_RESET_B_M1024_g N_A_33_74#_c_1543_n 0.00505633f $X=0.95 $Y=2.75 $X2=0
+ $Y2=0
cc_627 N_RESET_B_c_607_n N_A_33_74#_c_1544_n 0.00590946f $X=0.95 $Y=2.24 $X2=0
+ $Y2=0
cc_628 N_RESET_B_M1024_g N_A_33_74#_c_1544_n 0.0109584f $X=0.95 $Y=2.75 $X2=0
+ $Y2=0
cc_629 N_RESET_B_c_595_n N_A_33_74#_c_1544_n 0.0119937f $X=4.895 $Y=1.665 $X2=0
+ $Y2=0
cc_630 N_RESET_B_c_596_n N_A_33_74#_c_1544_n 0.00388391f $X=1.345 $Y=1.665 $X2=0
+ $Y2=0
cc_631 N_RESET_B_c_601_n N_A_33_74#_c_1544_n 4.69904e-19 $X=0.975 $Y=1.41 $X2=0
+ $Y2=0
cc_632 N_RESET_B_c_602_n N_A_33_74#_c_1544_n 0.0127196f $X=0.975 $Y=1.41 $X2=0
+ $Y2=0
cc_633 N_RESET_B_c_595_n N_A_33_74#_c_1538_n 0.0232099f $X=4.895 $Y=1.665 $X2=0
+ $Y2=0
cc_634 N_RESET_B_c_595_n N_A_33_74#_c_1546_n 0.00885572f $X=4.895 $Y=1.665 $X2=0
+ $Y2=0
cc_635 N_RESET_B_c_595_n N_A_33_74#_c_1540_n 0.00104731f $X=4.895 $Y=1.665 $X2=0
+ $Y2=0
cc_636 N_RESET_B_c_609_n N_A_33_74#_c_1547_n 0.00487673f $X=4.82 $Y=3.15 $X2=0
+ $Y2=0
cc_637 N_RESET_B_M1025_g N_A_33_74#_c_1541_n 0.00390091f $X=0.915 $Y=0.58 $X2=0
+ $Y2=0
cc_638 N_RESET_B_c_607_n N_A_33_74#_c_1548_n 0.00150754f $X=0.95 $Y=2.24 $X2=0
+ $Y2=0
cc_639 N_RESET_B_c_601_n N_A_33_74#_c_1548_n 0.00163166f $X=0.975 $Y=1.41 $X2=0
+ $Y2=0
cc_640 N_RESET_B_M1025_g N_VGND_c_1670_n 0.00554804f $X=0.915 $Y=0.58 $X2=0
+ $Y2=0
cc_641 N_RESET_B_c_601_n N_VGND_c_1670_n 0.00211787f $X=0.975 $Y=1.41 $X2=0
+ $Y2=0
cc_642 N_RESET_B_c_602_n N_VGND_c_1670_n 0.0105404f $X=0.975 $Y=1.41 $X2=0 $Y2=0
cc_643 N_RESET_B_c_594_n N_VGND_c_1672_n 0.00257506f $X=4.937 $Y=1.13 $X2=0
+ $Y2=0
cc_644 N_RESET_B_M1010_g N_VGND_c_1673_n 0.0103576f $X=8.605 $Y=0.805 $X2=0
+ $Y2=0
cc_645 N_RESET_B_M1025_g N_VGND_c_1675_n 0.00461464f $X=0.915 $Y=0.58 $X2=0
+ $Y2=0
cc_646 N_RESET_B_M1010_g N_VGND_c_1679_n 0.0035863f $X=8.605 $Y=0.805 $X2=0
+ $Y2=0
cc_647 N_RESET_B_M1025_g N_VGND_c_1681_n 0.00908835f $X=0.915 $Y=0.58 $X2=0
+ $Y2=0
cc_648 N_RESET_B_M1010_g N_VGND_c_1681_n 0.00401353f $X=8.605 $Y=0.805 $X2=0
+ $Y2=0
cc_649 N_RESET_B_c_594_n N_VGND_c_1681_n 7.33403e-19 $X=4.937 $Y=1.13 $X2=0
+ $Y2=0
cc_650 N_A_714_127#_c_831_n N_A_300_74#_c_940_n 3.88968e-19 $X=4.075 $Y=2.055
+ $X2=0 $Y2=0
cc_651 N_A_714_127#_c_831_n N_A_300_74#_c_941_n 0.00229506f $X=4.075 $Y=2.055
+ $X2=0 $Y2=0
cc_652 N_A_714_127#_c_831_n N_A_300_74#_c_943_n 0.0069401f $X=4.075 $Y=2.055
+ $X2=0 $Y2=0
cc_653 N_A_714_127#_c_825_n N_A_300_74#_M1030_g 0.00280137f $X=3.96 $Y=0.855
+ $X2=0 $Y2=0
cc_654 N_A_714_127#_M1020_g N_A_300_74#_c_928_n 0.00882199f $X=5.815 $Y=0.965
+ $X2=0 $Y2=0
cc_655 N_A_714_127#_M1020_g N_A_300_74#_M1006_g 0.0106687f $X=5.815 $Y=0.965
+ $X2=0 $Y2=0
cc_656 N_A_714_127#_c_823_n N_A_300_74#_c_936_n 4.20525e-19 $X=5.88 $Y=1.885
+ $X2=0 $Y2=0
cc_657 N_A_714_127#_c_823_n N_A_300_74#_c_937_n 0.0214064f $X=5.88 $Y=1.885
+ $X2=0 $Y2=0
cc_658 N_A_714_127#_c_833_n N_VPWR_M1008_s 0.00513921f $X=5.515 $Y=1.97 $X2=0
+ $Y2=0
cc_659 N_A_714_127#_c_826_n N_VPWR_M1008_s 5.6908e-19 $X=5.54 $Y=1.635 $X2=0
+ $Y2=0
cc_660 N_A_714_127#_c_830_n N_VPWR_c_1410_n 0.0262693f $X=4.97 $Y=2.055 $X2=0
+ $Y2=0
cc_661 N_A_714_127#_c_831_n N_VPWR_c_1410_n 0.0169789f $X=4.075 $Y=2.055 $X2=0
+ $Y2=0
cc_662 N_A_714_127#_c_832_n N_VPWR_c_1410_n 0.0155034f $X=5.135 $Y=2.55 $X2=0
+ $Y2=0
cc_663 N_A_714_127#_c_832_n N_VPWR_c_1411_n 0.00632461f $X=5.135 $Y=2.55 $X2=0
+ $Y2=0
cc_664 N_A_714_127#_c_823_n N_VPWR_c_1412_n 0.0143441f $X=5.88 $Y=1.885 $X2=0
+ $Y2=0
cc_665 N_A_714_127#_c_824_n N_VPWR_c_1412_n 0.00226809f $X=5.74 $Y=1.635 $X2=0
+ $Y2=0
cc_666 N_A_714_127#_c_832_n N_VPWR_c_1412_n 0.028876f $X=5.135 $Y=2.55 $X2=0
+ $Y2=0
cc_667 N_A_714_127#_c_833_n N_VPWR_c_1412_n 0.0138008f $X=5.515 $Y=1.97 $X2=0
+ $Y2=0
cc_668 N_A_714_127#_c_823_n N_VPWR_c_1416_n 0.00413917f $X=5.88 $Y=1.885 $X2=0
+ $Y2=0
cc_669 N_A_714_127#_c_831_n N_VPWR_c_1422_n 0.00813378f $X=4.075 $Y=2.055 $X2=0
+ $Y2=0
cc_670 N_A_714_127#_c_823_n N_VPWR_c_1405_n 0.00822528f $X=5.88 $Y=1.885 $X2=0
+ $Y2=0
cc_671 N_A_714_127#_c_831_n N_VPWR_c_1405_n 0.0121384f $X=4.075 $Y=2.055 $X2=0
+ $Y2=0
cc_672 N_A_714_127#_c_832_n N_VPWR_c_1405_n 0.010188f $X=5.135 $Y=2.55 $X2=0
+ $Y2=0
cc_673 N_A_714_127#_c_831_n N_A_33_74#_c_1546_n 0.0126499f $X=4.075 $Y=2.055
+ $X2=0 $Y2=0
cc_674 N_A_714_127#_c_831_n N_A_33_74#_c_1547_n 0.0265303f $X=4.075 $Y=2.055
+ $X2=0 $Y2=0
cc_675 N_A_300_74#_c_952_n N_A_1598_93#_M1000_g 0.0139991f $X=7.475 $Y=1.86
+ $X2=0 $Y2=0
cc_676 N_A_300_74#_c_944_n N_A_1598_93#_c_1122_n 0.0275569f $X=7.66 $Y=2.465
+ $X2=0 $Y2=0
cc_677 N_A_300_74#_c_947_n N_A_1598_93#_c_1122_n 0.0185966f $X=7.515 $Y=2.16
+ $X2=0 $Y2=0
cc_678 N_A_300_74#_c_934_n N_A_1266_119#_c_1229_n 0.00277079f $X=7.31 $Y=1.715
+ $X2=0 $Y2=0
cc_679 N_A_300_74#_c_947_n N_A_1266_119#_c_1222_n 9.05598e-19 $X=7.515 $Y=2.16
+ $X2=0 $Y2=0
cc_680 N_A_300_74#_c_951_n N_A_1266_119#_c_1222_n 0.0103637f $X=7.475 $Y=1.86
+ $X2=0 $Y2=0
cc_681 N_A_300_74#_c_944_n N_A_1266_119#_c_1213_n 0.00314472f $X=7.66 $Y=2.465
+ $X2=0 $Y2=0
cc_682 N_A_300_74#_c_947_n N_A_1266_119#_c_1213_n 0.0046061f $X=7.515 $Y=2.16
+ $X2=0 $Y2=0
cc_683 N_A_300_74#_c_934_n N_A_1266_119#_c_1213_n 0.01265f $X=7.31 $Y=1.715
+ $X2=0 $Y2=0
cc_684 N_A_300_74#_c_951_n N_A_1266_119#_c_1213_n 0.0415019f $X=7.475 $Y=1.86
+ $X2=0 $Y2=0
cc_685 N_A_300_74#_c_952_n N_A_1266_119#_c_1213_n 0.0057575f $X=7.475 $Y=1.86
+ $X2=0 $Y2=0
cc_686 N_A_300_74#_c_944_n N_A_1266_119#_c_1224_n 0.0157277f $X=7.66 $Y=2.465
+ $X2=0 $Y2=0
cc_687 N_A_300_74#_c_947_n N_A_1266_119#_c_1224_n 0.00213739f $X=7.515 $Y=2.16
+ $X2=0 $Y2=0
cc_688 N_A_300_74#_c_951_n N_A_1266_119#_c_1224_n 0.010457f $X=7.475 $Y=1.86
+ $X2=0 $Y2=0
cc_689 N_A_300_74#_c_948_n N_VPWR_M1017_s 0.00319186f $X=1.935 $Y=1.915 $X2=0
+ $Y2=0
cc_690 N_A_300_74#_c_933_n N_VPWR_M1017_s 7.22503e-19 $X=2.08 $Y=1.41 $X2=0
+ $Y2=0
cc_691 N_A_300_74#_c_938_n N_VPWR_c_1409_n 0.0176245f $X=2.46 $Y=1.66 $X2=0
+ $Y2=0
cc_692 N_A_300_74#_c_944_n N_VPWR_c_1413_n 0.00171173f $X=7.66 $Y=2.465 $X2=0
+ $Y2=0
cc_693 N_A_300_74#_c_944_n N_VPWR_c_1416_n 0.00323148f $X=7.66 $Y=2.465 $X2=0
+ $Y2=0
cc_694 N_A_300_74#_c_938_n N_VPWR_c_1405_n 8.51577e-19 $X=2.46 $Y=1.66 $X2=0
+ $Y2=0
cc_695 N_A_300_74#_c_943_n N_VPWR_c_1405_n 9.39239e-19 $X=3.56 $Y=2.24 $X2=0
+ $Y2=0
cc_696 N_A_300_74#_c_944_n N_VPWR_c_1405_n 0.00410412f $X=7.66 $Y=2.465 $X2=0
+ $Y2=0
cc_697 N_A_300_74#_M1007_d N_A_33_74#_c_1544_n 0.0121929f $X=1.53 $Y=1.735 $X2=0
+ $Y2=0
cc_698 N_A_300_74#_c_930_n N_A_33_74#_c_1544_n 0.00417404f $X=2.385 $Y=1.435
+ $X2=0 $Y2=0
cc_699 N_A_300_74#_c_948_n N_A_33_74#_c_1544_n 0.0440268f $X=1.935 $Y=1.915
+ $X2=0 $Y2=0
cc_700 N_A_300_74#_M1005_g N_A_33_74#_c_1598_n 0.0166858f $X=2.475 $Y=0.765
+ $X2=0 $Y2=0
cc_701 N_A_300_74#_c_935_n N_A_33_74#_c_1598_n 0.0090012f $X=1.64 $Y=0.515 $X2=0
+ $Y2=0
cc_702 N_A_300_74#_c_938_n N_A_33_74#_c_1538_n 0.0179363f $X=2.46 $Y=1.66 $X2=0
+ $Y2=0
cc_703 N_A_300_74#_M1005_g N_A_33_74#_c_1538_n 0.0167373f $X=2.475 $Y=0.765
+ $X2=0 $Y2=0
cc_704 N_A_300_74#_c_940_n N_A_33_74#_c_1538_n 0.00124925f $X=3.115 $Y=2.09
+ $X2=0 $Y2=0
cc_705 N_A_300_74#_c_930_n N_A_33_74#_c_1538_n 0.00989881f $X=2.385 $Y=1.435
+ $X2=0 $Y2=0
cc_706 N_A_300_74#_c_931_n N_A_33_74#_c_1538_n 0.0111237f $X=2.467 $Y=1.435
+ $X2=0 $Y2=0
cc_707 N_A_300_74#_c_933_n N_A_33_74#_c_1538_n 0.0544606f $X=2.08 $Y=1.41 $X2=0
+ $Y2=0
cc_708 N_A_300_74#_c_935_n N_A_33_74#_c_1538_n 0.0231781f $X=1.64 $Y=0.515 $X2=0
+ $Y2=0
cc_709 N_A_300_74#_c_938_n N_A_33_74#_c_1546_n 0.00597687f $X=2.46 $Y=1.66 $X2=0
+ $Y2=0
cc_710 N_A_300_74#_c_926_n N_A_33_74#_c_1546_n 0.00193439f $X=3.04 $Y=1.435
+ $X2=0 $Y2=0
cc_711 N_A_300_74#_c_941_n N_A_33_74#_c_1546_n 0.00898602f $X=3.485 $Y=2.165
+ $X2=0 $Y2=0
cc_712 N_A_300_74#_c_942_n N_A_33_74#_c_1546_n 0.00647124f $X=3.19 $Y=2.165
+ $X2=0 $Y2=0
cc_713 N_A_300_74#_c_943_n N_A_33_74#_c_1546_n 0.00254756f $X=3.56 $Y=2.24 $X2=0
+ $Y2=0
cc_714 N_A_300_74#_c_924_n N_A_33_74#_c_1539_n 0.0148765f $X=4.1 $Y=0.18 $X2=0
+ $Y2=0
cc_715 N_A_300_74#_c_926_n N_A_33_74#_c_1539_n 0.00656358f $X=3.04 $Y=1.435
+ $X2=0 $Y2=0
cc_716 N_A_300_74#_M1005_g N_A_33_74#_c_1540_n 0.00235195f $X=2.475 $Y=0.765
+ $X2=0 $Y2=0
cc_717 N_A_300_74#_c_926_n N_A_33_74#_c_1540_n 0.00209068f $X=3.04 $Y=1.435
+ $X2=0 $Y2=0
cc_718 N_A_300_74#_c_938_n N_A_33_74#_c_1547_n 0.00852038f $X=2.46 $Y=1.66 $X2=0
+ $Y2=0
cc_719 N_A_300_74#_c_943_n N_A_33_74#_c_1547_n 0.00141256f $X=3.56 $Y=2.24 $X2=0
+ $Y2=0
cc_720 N_A_300_74#_c_938_n N_A_33_74#_c_1618_n 0.0113559f $X=2.46 $Y=1.66 $X2=0
+ $Y2=0
cc_721 N_A_300_74#_c_933_n N_VGND_M1005_s 0.00119788f $X=2.08 $Y=1.41 $X2=0
+ $Y2=0
cc_722 N_A_300_74#_c_935_n N_VGND_M1005_s 0.00674215f $X=1.64 $Y=0.515 $X2=0
+ $Y2=0
cc_723 N_A_300_74#_c_935_n N_VGND_c_1670_n 0.0179276f $X=1.64 $Y=0.515 $X2=0
+ $Y2=0
cc_724 N_A_300_74#_c_925_n N_VGND_c_1671_n 0.0132299f $X=2.55 $Y=0.18 $X2=0
+ $Y2=0
cc_725 N_A_300_74#_c_935_n N_VGND_c_1671_n 0.0185934f $X=1.64 $Y=0.515 $X2=0
+ $Y2=0
cc_726 N_A_300_74#_c_928_n N_VGND_c_1672_n 0.0251635f $X=6.18 $Y=0.18 $X2=0
+ $Y2=0
cc_727 N_A_300_74#_c_935_n N_VGND_c_1676_n 0.0185803f $X=1.64 $Y=0.515 $X2=0
+ $Y2=0
cc_728 N_A_300_74#_c_925_n N_VGND_c_1677_n 0.0628542f $X=2.55 $Y=0.18 $X2=0
+ $Y2=0
cc_729 N_A_300_74#_c_928_n N_VGND_c_1678_n 0.0230598f $X=6.18 $Y=0.18 $X2=0
+ $Y2=0
cc_730 N_A_300_74#_c_924_n N_VGND_c_1681_n 0.0403945f $X=4.1 $Y=0.18 $X2=0 $Y2=0
cc_731 N_A_300_74#_c_925_n N_VGND_c_1681_n 0.00634026f $X=2.55 $Y=0.18 $X2=0
+ $Y2=0
cc_732 N_A_300_74#_c_928_n N_VGND_c_1681_n 0.0449069f $X=6.18 $Y=0.18 $X2=0
+ $Y2=0
cc_733 N_A_300_74#_c_932_n N_VGND_c_1681_n 0.00370846f $X=4.175 $Y=0.18 $X2=0
+ $Y2=0
cc_734 N_A_300_74#_c_935_n N_VGND_c_1681_n 0.0191168f $X=1.64 $Y=0.515 $X2=0
+ $Y2=0
cc_735 N_A_1598_93#_c_1119_n N_A_1266_119#_c_1207_n 0.0048734f $X=9.475 $Y=1.965
+ $X2=0 $Y2=0
cc_736 N_A_1598_93#_c_1120_n N_A_1266_119#_c_1207_n 0.00750942f $X=9.475
+ $Y=0.765 $X2=0 $Y2=0
cc_737 N_A_1598_93#_c_1125_n N_A_1266_119#_c_1208_n 0.00514416f $X=9.39 $Y=2.05
+ $X2=0 $Y2=0
cc_738 N_A_1598_93#_c_1127_n N_A_1266_119#_c_1208_n 0.00291268f $X=8.865 $Y=2.15
+ $X2=0 $Y2=0
cc_739 N_A_1598_93#_c_1124_n N_A_1266_119#_c_1218_n 0.00130111f $X=8.845 $Y=2.75
+ $X2=0 $Y2=0
cc_740 N_A_1598_93#_c_1125_n N_A_1266_119#_c_1218_n 0.00755711f $X=9.39 $Y=2.05
+ $X2=0 $Y2=0
cc_741 N_A_1598_93#_c_1127_n N_A_1266_119#_c_1218_n 0.015254f $X=8.865 $Y=2.15
+ $X2=0 $Y2=0
cc_742 N_A_1598_93#_c_1124_n N_A_1266_119#_c_1219_n 0.0111813f $X=8.845 $Y=2.75
+ $X2=0 $Y2=0
cc_743 N_A_1598_93#_c_1125_n N_A_1266_119#_c_1209_n 6.15368e-19 $X=9.39 $Y=2.05
+ $X2=0 $Y2=0
cc_744 N_A_1598_93#_c_1119_n N_A_1266_119#_c_1209_n 0.0128412f $X=9.475 $Y=1.965
+ $X2=0 $Y2=0
cc_745 N_A_1598_93#_c_1120_n N_A_1266_119#_c_1209_n 8.36802e-19 $X=9.475
+ $Y=0.765 $X2=0 $Y2=0
cc_746 N_A_1598_93#_c_1125_n N_A_1266_119#_c_1220_n 0.0109475f $X=9.39 $Y=2.05
+ $X2=0 $Y2=0
cc_747 N_A_1598_93#_c_1119_n N_A_1266_119#_c_1220_n 0.00680794f $X=9.475
+ $Y=1.965 $X2=0 $Y2=0
cc_748 N_A_1598_93#_c_1119_n N_A_1266_119#_c_1210_n 7.21124e-19 $X=9.475
+ $Y=1.965 $X2=0 $Y2=0
cc_749 N_A_1598_93#_c_1120_n N_A_1266_119#_c_1210_n 7.36949e-19 $X=9.475
+ $Y=0.765 $X2=0 $Y2=0
cc_750 N_A_1598_93#_c_1125_n N_A_1266_119#_c_1221_n 3.81375e-19 $X=9.39 $Y=2.05
+ $X2=0 $Y2=0
cc_751 N_A_1598_93#_c_1120_n N_A_1266_119#_c_1211_n 0.0071021f $X=9.475 $Y=0.765
+ $X2=0 $Y2=0
cc_752 N_A_1598_93#_M1000_g N_A_1266_119#_c_1229_n 0.00369318f $X=8.065 $Y=0.805
+ $X2=0 $Y2=0
cc_753 N_A_1598_93#_M1000_g N_A_1266_119#_c_1212_n 0.00375809f $X=8.065 $Y=0.805
+ $X2=0 $Y2=0
cc_754 N_A_1598_93#_M1000_g N_A_1266_119#_c_1213_n 0.0199131f $X=8.065 $Y=0.805
+ $X2=0 $Y2=0
cc_755 N_A_1598_93#_c_1122_n N_A_1266_119#_c_1213_n 0.00132521f $X=8.08 $Y=2.465
+ $X2=0 $Y2=0
cc_756 N_A_1598_93#_c_1123_n N_A_1266_119#_c_1213_n 0.0293641f $X=8.68 $Y=2.15
+ $X2=0 $Y2=0
cc_757 N_A_1598_93#_M1000_g N_A_1266_119#_c_1214_n 0.0157592f $X=8.065 $Y=0.805
+ $X2=0 $Y2=0
cc_758 N_A_1598_93#_c_1123_n N_A_1266_119#_c_1214_n 0.0023008f $X=8.68 $Y=2.15
+ $X2=0 $Y2=0
cc_759 N_A_1598_93#_c_1127_n N_A_1266_119#_c_1214_n 0.00676946f $X=8.865 $Y=2.15
+ $X2=0 $Y2=0
cc_760 N_A_1598_93#_c_1122_n N_A_1266_119#_c_1224_n 0.00189609f $X=8.08 $Y=2.465
+ $X2=0 $Y2=0
cc_761 N_A_1598_93#_c_1125_n N_A_1266_119#_c_1215_n 0.0128235f $X=9.39 $Y=2.05
+ $X2=0 $Y2=0
cc_762 N_A_1598_93#_c_1119_n N_A_1266_119#_c_1215_n 0.0502151f $X=9.475 $Y=1.965
+ $X2=0 $Y2=0
cc_763 N_A_1598_93#_c_1127_n N_A_1266_119#_c_1215_n 0.0110236f $X=8.865 $Y=2.15
+ $X2=0 $Y2=0
cc_764 N_A_1598_93#_c_1120_n N_A_1266_119#_c_1215_n 0.0121056f $X=9.475 $Y=0.765
+ $X2=0 $Y2=0
cc_765 N_A_1598_93#_c_1119_n N_A_1266_119#_c_1216_n 0.0103445f $X=9.475 $Y=1.965
+ $X2=0 $Y2=0
cc_766 N_A_1598_93#_c_1124_n N_A_1934_94#_c_1352_n 0.00529924f $X=8.845 $Y=2.75
+ $X2=0 $Y2=0
cc_767 N_A_1598_93#_c_1127_n N_A_1934_94#_c_1352_n 9.63229e-19 $X=8.865 $Y=2.15
+ $X2=0 $Y2=0
cc_768 N_A_1598_93#_c_1119_n N_A_1934_94#_c_1347_n 0.0270211f $X=9.475 $Y=1.965
+ $X2=0 $Y2=0
cc_769 N_A_1598_93#_c_1120_n N_A_1934_94#_c_1347_n 0.0315201f $X=9.475 $Y=0.765
+ $X2=0 $Y2=0
cc_770 N_A_1598_93#_c_1125_n N_A_1934_94#_c_1348_n 0.0140451f $X=9.39 $Y=2.05
+ $X2=0 $Y2=0
cc_771 N_A_1598_93#_c_1119_n N_A_1934_94#_c_1348_n 0.0238206f $X=9.475 $Y=1.965
+ $X2=0 $Y2=0
cc_772 N_A_1598_93#_c_1119_n N_A_1934_94#_c_1350_n 0.0278717f $X=9.475 $Y=1.965
+ $X2=0 $Y2=0
cc_773 N_A_1598_93#_c_1122_n N_VPWR_c_1413_n 0.0154036f $X=8.08 $Y=2.465 $X2=0
+ $Y2=0
cc_774 N_A_1598_93#_c_1123_n N_VPWR_c_1413_n 0.0267292f $X=8.68 $Y=2.15 $X2=0
+ $Y2=0
cc_775 N_A_1598_93#_c_1124_n N_VPWR_c_1413_n 0.0304142f $X=8.845 $Y=2.75 $X2=0
+ $Y2=0
cc_776 N_A_1598_93#_c_1124_n N_VPWR_c_1414_n 0.0309026f $X=8.845 $Y=2.75 $X2=0
+ $Y2=0
cc_777 N_A_1598_93#_c_1125_n N_VPWR_c_1414_n 0.0121819f $X=9.39 $Y=2.05 $X2=0
+ $Y2=0
cc_778 N_A_1598_93#_c_1122_n N_VPWR_c_1416_n 0.00413917f $X=8.08 $Y=2.465 $X2=0
+ $Y2=0
cc_779 N_A_1598_93#_c_1124_n N_VPWR_c_1423_n 0.014552f $X=8.845 $Y=2.75 $X2=0
+ $Y2=0
cc_780 N_A_1598_93#_c_1122_n N_VPWR_c_1405_n 0.0085536f $X=8.08 $Y=2.465 $X2=0
+ $Y2=0
cc_781 N_A_1598_93#_c_1124_n N_VPWR_c_1405_n 0.0119791f $X=8.845 $Y=2.75 $X2=0
+ $Y2=0
cc_782 N_A_1598_93#_M1000_g N_VGND_c_1673_n 0.00889071f $X=8.065 $Y=0.805 $X2=0
+ $Y2=0
cc_783 N_A_1598_93#_c_1120_n N_VGND_c_1673_n 0.0110474f $X=9.475 $Y=0.765 $X2=0
+ $Y2=0
cc_784 N_A_1598_93#_M1000_g N_VGND_c_1678_n 0.0035863f $X=8.065 $Y=0.805 $X2=0
+ $Y2=0
cc_785 N_A_1598_93#_c_1120_n N_VGND_c_1679_n 0.0112924f $X=9.475 $Y=0.765 $X2=0
+ $Y2=0
cc_786 N_A_1598_93#_M1000_g N_VGND_c_1681_n 0.00401353f $X=8.065 $Y=0.805 $X2=0
+ $Y2=0
cc_787 N_A_1598_93#_c_1120_n N_VGND_c_1681_n 0.0158807f $X=9.475 $Y=0.765 $X2=0
+ $Y2=0
cc_788 N_A_1266_119#_c_1210_n N_A_1934_94#_c_1345_n 0.0160558f $X=10.03 $Y=1.125
+ $X2=0 $Y2=0
cc_789 N_A_1266_119#_c_1220_n N_A_1934_94#_c_1346_n 0.00551483f $X=9.965 $Y=1.97
+ $X2=0 $Y2=0
cc_790 N_A_1266_119#_c_1221_n N_A_1934_94#_c_1346_n 0.0170234f $X=10.04 $Y=2.045
+ $X2=0 $Y2=0
cc_791 N_A_1266_119#_c_1218_n N_A_1934_94#_c_1352_n 0.00273194f $X=9.07 $Y=2.375
+ $X2=0 $Y2=0
cc_792 N_A_1266_119#_c_1219_n N_A_1934_94#_c_1352_n 0.0015885f $X=9.07 $Y=2.465
+ $X2=0 $Y2=0
cc_793 N_A_1266_119#_c_1220_n N_A_1934_94#_c_1352_n 0.00292339f $X=9.965 $Y=1.97
+ $X2=0 $Y2=0
cc_794 N_A_1266_119#_c_1221_n N_A_1934_94#_c_1352_n 0.00167606f $X=10.04
+ $Y=2.045 $X2=0 $Y2=0
cc_795 N_A_1266_119#_c_1221_n N_A_1934_94#_c_1353_n 0.00842612f $X=10.04
+ $Y=2.045 $X2=0 $Y2=0
cc_796 N_A_1266_119#_c_1207_n N_A_1934_94#_c_1347_n 0.00140435f $X=8.995
+ $Y=1.125 $X2=0 $Y2=0
cc_797 N_A_1266_119#_c_1209_n N_A_1934_94#_c_1347_n 0.0161335f $X=9.955 $Y=1.2
+ $X2=0 $Y2=0
cc_798 N_A_1266_119#_c_1210_n N_A_1934_94#_c_1347_n 0.010444f $X=10.03 $Y=1.125
+ $X2=0 $Y2=0
cc_799 N_A_1266_119#_c_1218_n N_A_1934_94#_c_1348_n 0.00438224f $X=9.07 $Y=2.375
+ $X2=0 $Y2=0
cc_800 N_A_1266_119#_c_1220_n N_A_1934_94#_c_1348_n 0.0166743f $X=9.965 $Y=1.97
+ $X2=0 $Y2=0
cc_801 N_A_1266_119#_c_1221_n N_A_1934_94#_c_1348_n 0.00434926f $X=10.04
+ $Y=2.045 $X2=0 $Y2=0
cc_802 N_A_1266_119#_c_1209_n N_A_1934_94#_c_1349_n 0.00434645f $X=9.955 $Y=1.2
+ $X2=0 $Y2=0
cc_803 N_A_1266_119#_c_1220_n N_A_1934_94#_c_1349_n 0.00425121f $X=9.965 $Y=1.97
+ $X2=0 $Y2=0
cc_804 N_A_1266_119#_c_1213_n N_VPWR_c_1413_n 8.41136e-19 $X=7.815 $Y=2.535
+ $X2=0 $Y2=0
cc_805 N_A_1266_119#_c_1224_n N_VPWR_c_1413_n 0.0157089f $X=7.435 $Y=2.7 $X2=0
+ $Y2=0
cc_806 N_A_1266_119#_c_1219_n N_VPWR_c_1414_n 0.00729942f $X=9.07 $Y=2.465 $X2=0
+ $Y2=0
cc_807 N_A_1266_119#_c_1220_n N_VPWR_c_1414_n 0.00128121f $X=9.965 $Y=1.97 $X2=0
+ $Y2=0
cc_808 N_A_1266_119#_c_1221_n N_VPWR_c_1414_n 0.00366284f $X=10.04 $Y=2.045
+ $X2=0 $Y2=0
cc_809 N_A_1266_119#_c_1221_n N_VPWR_c_1415_n 0.00784561f $X=10.04 $Y=2.045
+ $X2=0 $Y2=0
cc_810 N_A_1266_119#_c_1222_n N_VPWR_c_1416_n 0.0150066f $X=7.435 $Y=2.7 $X2=0
+ $Y2=0
cc_811 N_A_1266_119#_c_1224_n N_VPWR_c_1416_n 0.00884848f $X=7.435 $Y=2.7 $X2=0
+ $Y2=0
cc_812 N_A_1266_119#_c_1221_n N_VPWR_c_1418_n 0.00445602f $X=10.04 $Y=2.045
+ $X2=0 $Y2=0
cc_813 N_A_1266_119#_c_1219_n N_VPWR_c_1423_n 0.00445602f $X=9.07 $Y=2.465 $X2=0
+ $Y2=0
cc_814 N_A_1266_119#_c_1219_n N_VPWR_c_1405_n 0.00900303f $X=9.07 $Y=2.465 $X2=0
+ $Y2=0
cc_815 N_A_1266_119#_c_1221_n N_VPWR_c_1405_n 0.00862274f $X=10.04 $Y=2.045
+ $X2=0 $Y2=0
cc_816 N_A_1266_119#_c_1222_n N_VPWR_c_1405_n 0.0187253f $X=7.435 $Y=2.7 $X2=0
+ $Y2=0
cc_817 N_A_1266_119#_c_1224_n N_VPWR_c_1405_n 0.013677f $X=7.435 $Y=2.7 $X2=0
+ $Y2=0
cc_818 N_A_1266_119#_c_1224_n A_1547_508# 0.00356592f $X=7.435 $Y=2.7 $X2=-0.19
+ $Y2=-0.245
cc_819 N_A_1266_119#_c_1209_n N_Q_c_1642_n 2.48707e-19 $X=9.955 $Y=1.2 $X2=0
+ $Y2=0
cc_820 N_A_1266_119#_c_1220_n Q 6.01794e-19 $X=9.965 $Y=1.97 $X2=0 $Y2=0
cc_821 N_A_1266_119#_c_1221_n Q 4.02579e-19 $X=10.04 $Y=2.045 $X2=0 $Y2=0
cc_822 N_A_1266_119#_c_1207_n N_VGND_c_1673_n 0.00147671f $X=8.995 $Y=1.125
+ $X2=0 $Y2=0
cc_823 N_A_1266_119#_c_1229_n N_VGND_c_1673_n 0.0196844f $X=7.73 $Y=0.79 $X2=0
+ $Y2=0
cc_824 N_A_1266_119#_c_1214_n N_VGND_c_1673_n 0.0254301f $X=8.92 $Y=1.21 $X2=0
+ $Y2=0
cc_825 N_A_1266_119#_c_1210_n N_VGND_c_1674_n 0.0072589f $X=10.03 $Y=1.125 $X2=0
+ $Y2=0
cc_826 N_A_1266_119#_c_1229_n N_VGND_c_1678_n 0.0212446f $X=7.73 $Y=0.79 $X2=0
+ $Y2=0
cc_827 N_A_1266_119#_c_1207_n N_VGND_c_1679_n 0.00414396f $X=8.995 $Y=1.125
+ $X2=0 $Y2=0
cc_828 N_A_1266_119#_c_1210_n N_VGND_c_1679_n 0.00486718f $X=10.03 $Y=1.125
+ $X2=0 $Y2=0
cc_829 N_A_1266_119#_c_1207_n N_VGND_c_1681_n 0.00477801f $X=8.995 $Y=1.125
+ $X2=0 $Y2=0
cc_830 N_A_1266_119#_c_1210_n N_VGND_c_1681_n 0.00514438f $X=10.03 $Y=1.125
+ $X2=0 $Y2=0
cc_831 N_A_1266_119#_c_1229_n N_VGND_c_1681_n 0.0353228f $X=7.73 $Y=0.79 $X2=0
+ $Y2=0
cc_832 N_A_1266_119#_c_1229_n A_1550_119# 0.00494929f $X=7.73 $Y=0.79 $X2=-0.19
+ $Y2=-0.245
cc_833 N_A_1266_119#_c_1212_n A_1550_119# 6.55526e-19 $X=7.815 $Y=1.125
+ $X2=-0.19 $Y2=-0.245
cc_834 N_A_1934_94#_c_1353_n N_VPWR_c_1414_n 0.0346921f $X=9.815 $Y=2.815 $X2=0
+ $Y2=0
cc_835 N_A_1934_94#_c_1346_n N_VPWR_c_1415_n 0.00845898f $X=10.545 $Y=1.765
+ $X2=0 $Y2=0
cc_836 N_A_1934_94#_c_1348_n N_VPWR_c_1415_n 0.0341417f $X=9.815 $Y=2.27 $X2=0
+ $Y2=0
cc_837 N_A_1934_94#_c_1349_n N_VPWR_c_1415_n 0.0104409f $X=10.48 $Y=1.485 $X2=0
+ $Y2=0
cc_838 N_A_1934_94#_c_1353_n N_VPWR_c_1418_n 0.0145919f $X=9.815 $Y=2.815 $X2=0
+ $Y2=0
cc_839 N_A_1934_94#_c_1346_n N_VPWR_c_1424_n 0.00445602f $X=10.545 $Y=1.765
+ $X2=0 $Y2=0
cc_840 N_A_1934_94#_c_1346_n N_VPWR_c_1405_n 0.00861717f $X=10.545 $Y=1.765
+ $X2=0 $Y2=0
cc_841 N_A_1934_94#_c_1353_n N_VPWR_c_1405_n 0.0120459f $X=9.815 $Y=2.815 $X2=0
+ $Y2=0
cc_842 N_A_1934_94#_c_1345_n N_Q_c_1642_n 0.00640271f $X=10.54 $Y=1.32 $X2=0
+ $Y2=0
cc_843 N_A_1934_94#_c_1345_n N_Q_c_1643_n 0.00241276f $X=10.54 $Y=1.32 $X2=0
+ $Y2=0
cc_844 N_A_1934_94#_c_1347_n N_Q_c_1643_n 5.13862e-19 $X=9.815 $Y=0.745 $X2=0
+ $Y2=0
cc_845 N_A_1934_94#_c_1349_n N_Q_c_1643_n 0.00188005f $X=10.48 $Y=1.485 $X2=0
+ $Y2=0
cc_846 N_A_1934_94#_c_1346_n Q 0.0049232f $X=10.545 $Y=1.765 $X2=0 $Y2=0
cc_847 N_A_1934_94#_c_1348_n Q 0.0072771f $X=9.815 $Y=2.27 $X2=0 $Y2=0
cc_848 N_A_1934_94#_c_1349_n Q 7.18422e-19 $X=10.48 $Y=1.485 $X2=0 $Y2=0
cc_849 N_A_1934_94#_c_1346_n Q 0.0126267f $X=10.545 $Y=1.765 $X2=0 $Y2=0
cc_850 N_A_1934_94#_c_1345_n N_Q_c_1644_n 0.0040915f $X=10.54 $Y=1.32 $X2=0
+ $Y2=0
cc_851 N_A_1934_94#_c_1346_n N_Q_c_1644_n 0.0119541f $X=10.545 $Y=1.765 $X2=0
+ $Y2=0
cc_852 N_A_1934_94#_c_1349_n N_Q_c_1644_n 0.0262114f $X=10.48 $Y=1.485 $X2=0
+ $Y2=0
cc_853 N_A_1934_94#_c_1345_n N_VGND_c_1674_n 0.00292117f $X=10.54 $Y=1.32 $X2=0
+ $Y2=0
cc_854 N_A_1934_94#_c_1346_n N_VGND_c_1674_n 0.00216466f $X=10.545 $Y=1.765
+ $X2=0 $Y2=0
cc_855 N_A_1934_94#_c_1347_n N_VGND_c_1674_n 0.024751f $X=9.815 $Y=0.745 $X2=0
+ $Y2=0
cc_856 N_A_1934_94#_c_1349_n N_VGND_c_1674_n 0.0194281f $X=10.48 $Y=1.485 $X2=0
+ $Y2=0
cc_857 N_A_1934_94#_c_1347_n N_VGND_c_1679_n 0.00541117f $X=9.815 $Y=0.745 $X2=0
+ $Y2=0
cc_858 N_A_1934_94#_c_1345_n N_VGND_c_1680_n 0.00485341f $X=10.54 $Y=1.32 $X2=0
+ $Y2=0
cc_859 N_A_1934_94#_c_1345_n N_VGND_c_1681_n 0.00514438f $X=10.54 $Y=1.32 $X2=0
+ $Y2=0
cc_860 N_A_1934_94#_c_1347_n N_VGND_c_1681_n 0.00809617f $X=9.815 $Y=0.745 $X2=0
+ $Y2=0
cc_861 N_VPWR_c_1407_n N_A_33_74#_c_1543_n 0.0307071f $X=0.275 $Y=2.75 $X2=0
+ $Y2=0
cc_862 N_VPWR_c_1408_n N_A_33_74#_c_1543_n 0.00307778f $X=1.18 $Y=2.685 $X2=0
+ $Y2=0
cc_863 N_VPWR_c_1420_n N_A_33_74#_c_1543_n 0.0101736f $X=1.04 $Y=3.33 $X2=0
+ $Y2=0
cc_864 N_VPWR_c_1405_n N_A_33_74#_c_1543_n 0.0084208f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_865 N_VPWR_M1024_d N_A_33_74#_c_1544_n 0.00534841f $X=1.025 $Y=2.54 $X2=0
+ $Y2=0
cc_866 N_VPWR_M1017_s N_A_33_74#_c_1544_n 0.00545122f $X=2.09 $Y=1.735 $X2=0
+ $Y2=0
cc_867 N_VPWR_c_1408_n N_A_33_74#_c_1544_n 0.0231726f $X=1.18 $Y=2.685 $X2=0
+ $Y2=0
cc_868 N_VPWR_c_1409_n N_A_33_74#_c_1544_n 0.0209681f $X=2.235 $Y=2.605 $X2=0
+ $Y2=0
cc_869 N_VPWR_c_1422_n N_A_33_74#_c_1547_n 0.00516451f $X=4.46 $Y=3.33 $X2=0
+ $Y2=0
cc_870 N_VPWR_c_1405_n N_A_33_74#_c_1547_n 0.00669853f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_871 N_VPWR_c_1409_n N_A_33_74#_c_1618_n 0.00114279f $X=2.235 $Y=2.605 $X2=0
+ $Y2=0
cc_872 N_VPWR_c_1415_n Q 0.0581843f $X=10.315 $Y=2.265 $X2=0 $Y2=0
cc_873 N_VPWR_c_1424_n Q 0.0154862f $X=10.8 $Y=3.33 $X2=0 $Y2=0
cc_874 N_VPWR_c_1405_n Q 0.0127853f $X=10.8 $Y=3.33 $X2=0 $Y2=0
cc_875 N_A_33_74#_c_1541_n A_120_74# 0.00489958f $X=0.625 $Y=0.57 $X2=-0.19
+ $Y2=-0.245
cc_876 N_A_33_74#_c_1598_n N_VGND_M1005_s 0.00155908f $X=2.42 $Y=0.725 $X2=0
+ $Y2=0
cc_877 N_A_33_74#_c_1538_n N_VGND_M1005_s 0.00435099f $X=2.42 $Y=2.18 $X2=0
+ $Y2=0
cc_878 N_A_33_74#_c_1537_n N_VGND_c_1670_n 9.42187e-19 $X=0.625 $Y=2.18 $X2=0
+ $Y2=0
cc_879 N_A_33_74#_c_1541_n N_VGND_c_1670_n 0.0120647f $X=0.625 $Y=0.57 $X2=0
+ $Y2=0
cc_880 N_A_33_74#_c_1541_n N_VGND_c_1675_n 0.0239076f $X=0.625 $Y=0.57 $X2=0
+ $Y2=0
cc_881 N_A_33_74#_c_1598_n N_VGND_c_1677_n 0.00442729f $X=2.42 $Y=0.725 $X2=0
+ $Y2=0
cc_882 N_A_33_74#_c_1539_n N_VGND_c_1677_n 0.0205725f $X=3.115 $Y=0.57 $X2=0
+ $Y2=0
cc_883 N_A_33_74#_c_1598_n N_VGND_c_1681_n 0.00690817f $X=2.42 $Y=0.725 $X2=0
+ $Y2=0
cc_884 N_A_33_74#_c_1539_n N_VGND_c_1681_n 0.022547f $X=3.115 $Y=0.57 $X2=0
+ $Y2=0
cc_885 N_A_33_74#_c_1541_n N_VGND_c_1681_n 0.0198316f $X=0.625 $Y=0.57 $X2=0
+ $Y2=0
cc_886 N_Q_c_1642_n N_VGND_c_1674_n 0.0261897f $X=10.755 $Y=0.605 $X2=0 $Y2=0
cc_887 N_Q_c_1642_n N_VGND_c_1680_n 0.0118258f $X=10.755 $Y=0.605 $X2=0 $Y2=0
cc_888 N_Q_c_1642_n N_VGND_c_1681_n 0.0126447f $X=10.755 $Y=0.605 $X2=0 $Y2=0
