* File: sky130_fd_sc_ls__or4b_1.pex.spice
* Created: Fri Aug 28 14:00:11 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__OR4B_1%D_N 3 5 6 7 9 10 14
r37 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.405
+ $Y=1.615 $X2=0.405 $Y2=1.615
r38 10 14 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.24 $Y=1.615
+ $X2=0.405 $Y2=1.615
r39 7 9 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.51 $Y=2.045 $X2=0.51
+ $Y2=2.54
r40 6 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.51 $Y=1.955 $X2=0.51
+ $Y2=2.045
r41 5 13 34.0194 $w=3.43e-07 $l=2.05122e-07 $layer=POLY_cond $X=0.51 $Y=1.78
+ $X2=0.42 $Y2=1.615
r42 5 6 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=0.51 $Y=1.78 $X2=0.51
+ $Y2=1.955
r43 1 13 38.7084 $w=3.43e-07 $l=1.98997e-07 $layer=POLY_cond $X=0.495 $Y=1.45
+ $X2=0.42 $Y2=1.615
r44 1 3 412.777 $w=1.5e-07 $l=8.05e-07 $layer=POLY_cond $X=0.495 $Y=1.45
+ $X2=0.495 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_LS__OR4B_1%A_27_74# 1 2 9 11 13 15 18 22 24 25 26 27 29
+ 31 34
c72 13 0 1.1364e-19 $X=1.705 $Y=1.765
r73 34 35 36.5941 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=0.975 $Y=1.69
+ $X2=0.975 $Y2=1.58
r74 32 34 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=0.975 $Y=1.745
+ $X2=0.975 $Y2=1.69
r75 31 33 13.2509 $w=2.67e-07 $l=2.9e-07 $layer=LI1_cond $X=0.975 $Y=1.745
+ $X2=0.975 $Y2=2.035
r76 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.975
+ $Y=1.745 $X2=0.975 $Y2=1.745
r77 29 31 9.14344 $w=2.67e-07 $l=2.0106e-07 $layer=LI1_cond $X=0.895 $Y=1.58
+ $X2=0.975 $Y2=1.745
r78 28 29 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=0.895 $Y=1.28
+ $X2=0.895 $Y2=1.58
r79 26 33 3.37873 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.81 $Y=2.035
+ $X2=0.975 $Y2=2.035
r80 26 27 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=0.81 $Y=2.035
+ $X2=0.45 $Y2=2.035
r81 24 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.81 $Y=1.195
+ $X2=0.895 $Y2=1.28
r82 24 25 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.81 $Y=1.195
+ $X2=0.445 $Y2=1.195
r83 20 27 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.285 $Y=2.12
+ $X2=0.45 $Y2=2.035
r84 20 22 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=0.285 $Y=2.12
+ $X2=0.285 $Y2=2.265
r85 16 25 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=1.11
+ $X2=0.445 $Y2=1.195
r86 16 18 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=0.28 $Y=1.11
+ $X2=0.28 $Y2=0.645
r87 13 15 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.705 $Y=1.765
+ $X2=1.705 $Y2=2.34
r88 12 34 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.14 $Y=1.69
+ $X2=0.975 $Y2=1.69
r89 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.63 $Y=1.69
+ $X2=1.705 $Y2=1.765
r90 11 12 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=1.63 $Y=1.69
+ $X2=1.14 $Y2=1.69
r91 9 35 479.436 $w=1.5e-07 $l=9.35e-07 $layer=POLY_cond $X=1.065 $Y=0.645
+ $X2=1.065 $Y2=1.58
r92 2 22 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.14
+ $Y=2.12 $X2=0.285 $Y2=2.265
r93 1 18 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_LS__OR4B_1%C 2 3 5 8 9 10 14 15 16
c37 15 0 1.65595e-19 $X=2.05 $Y=1.21
c38 3 0 4.38706e-20 $X=2.125 $Y=1.765
r39 14 17 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.05 $Y=1.21
+ $X2=2.05 $Y2=1.375
r40 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.05 $Y=1.21
+ $X2=2.05 $Y2=1.045
r41 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.05
+ $Y=1.21 $X2=2.05 $Y2=1.21
r42 9 10 10.9334 $w=3.88e-07 $l=3.7e-07 $layer=LI1_cond $X=2.08 $Y=1.295
+ $X2=2.08 $Y2=1.665
r43 9 15 2.51173 $w=3.88e-07 $l=8.5e-08 $layer=LI1_cond $X=2.08 $Y=1.295
+ $X2=2.08 $Y2=1.21
r44 8 16 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.14 $Y=0.645 $X2=2.14
+ $Y2=1.045
r45 3 5 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.125 $Y=1.765
+ $X2=2.125 $Y2=2.34
r46 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.125 $Y=1.675 $X2=2.125
+ $Y2=1.765
r47 2 17 116.613 $w=1.8e-07 $l=3e-07 $layer=POLY_cond $X=2.125 $Y=1.675
+ $X2=2.125 $Y2=1.375
.ends

.subckt PM_SKY130_FD_SC_LS__OR4B_1%B 2 3 5 8 10 11 15
c36 10 0 4.38706e-20 $X=2.64 $Y=1.295
c37 3 0 9.28485e-20 $X=2.545 $Y=1.765
r38 15 18 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.62 $Y=1.345
+ $X2=2.62 $Y2=1.51
r39 15 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.62 $Y=1.345
+ $X2=2.62 $Y2=1.18
r40 10 11 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.62 $Y=1.295
+ $X2=2.62 $Y2=1.665
r41 10 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.62
+ $Y=1.345 $X2=2.62 $Y2=1.345
r42 8 17 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=2.71 $Y=0.645
+ $X2=2.71 $Y2=1.18
r43 3 5 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.545 $Y=1.765
+ $X2=2.545 $Y2=2.34
r44 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.545 $Y=1.675 $X2=2.545
+ $Y2=1.765
r45 2 18 64.1371 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.545 $Y=1.675
+ $X2=2.545 $Y2=1.51
.ends

.subckt PM_SKY130_FD_SC_LS__OR4B_1%A 1 3 6 8 12
c39 12 0 4.08937e-20 $X=3.16 $Y=1.515
c40 6 0 7.34258e-20 $X=3.14 $Y=0.645
c41 1 0 1.19108e-19 $X=3.085 $Y=1.765
r42 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.16
+ $Y=1.515 $X2=3.16 $Y2=1.515
r43 8 12 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=3.16 $Y=1.665
+ $X2=3.16 $Y2=1.515
r44 4 11 38.5562 $w=2.99e-07 $l=1.74714e-07 $layer=POLY_cond $X=3.14 $Y=1.35
+ $X2=3.16 $Y2=1.515
r45 4 6 361.5 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=3.14 $Y=1.35 $X2=3.14
+ $Y2=0.645
r46 1 11 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=3.085 $Y=1.765
+ $X2=3.16 $Y2=1.515
r47 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.085 $Y=1.765
+ $X2=3.085 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_LS__OR4B_1%A_228_74# 1 2 3 10 12 15 17 18 21 25 27 29 32
+ 34 35 39
r100 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.73
+ $Y=1.465 $X2=3.73 $Y2=1.465
r101 34 43 9.00568 $w=2.92e-07 $l=2.14942e-07 $layer=LI1_cond $X=3.58 $Y=1.63
+ $X2=3.695 $Y2=1.465
r102 34 35 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=3.58 $Y=1.63
+ $X2=3.58 $Y2=1.95
r103 33 40 3.08766 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=3.125 $Y=1.095
+ $X2=2.955 $Y2=1.095
r104 32 43 15.4589 $w=2.92e-07 $l=4.59238e-07 $layer=LI1_cond $X=3.495 $Y=1.095
+ $X2=3.695 $Y2=1.465
r105 32 33 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.495 $Y=1.095
+ $X2=3.125 $Y2=1.095
r106 29 40 12.4049 $w=3.65e-07 $l=3.43439e-07 $layer=LI1_cond $X=2.942 $Y=0.758
+ $X2=2.955 $Y2=1.095
r107 29 31 3.77699 $w=3.65e-07 $l=1.13e-07 $layer=LI1_cond $X=2.942 $Y=0.758
+ $X2=2.942 $Y2=0.645
r108 28 39 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.645 $Y=2.035
+ $X2=1.48 $Y2=2.035
r109 27 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.495 $Y=2.035
+ $X2=3.58 $Y2=1.95
r110 27 28 120.695 $w=1.68e-07 $l=1.85e-06 $layer=LI1_cond $X=3.495 $Y=2.035
+ $X2=1.645 $Y2=2.035
r111 23 37 3.40825 $w=3.3e-07 $l=2.65e-07 $layer=LI1_cond $X=1.645 $Y=0.71
+ $X2=1.38 $Y2=0.71
r112 23 25 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=1.645 $Y=0.71
+ $X2=1.925 $Y2=0.71
r113 19 39 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.48 $Y=2.12
+ $X2=1.48 $Y2=2.035
r114 19 21 20.0804 $w=3.28e-07 $l=5.75e-07 $layer=LI1_cond $X=1.48 $Y=2.12
+ $X2=1.48 $Y2=2.695
r115 18 39 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.48 $Y=1.95
+ $X2=1.48 $Y2=2.035
r116 17 37 3.40825 $w=3.3e-07 $l=2.09105e-07 $layer=LI1_cond $X=1.48 $Y=0.875
+ $X2=1.38 $Y2=0.71
r117 17 18 37.5417 $w=3.28e-07 $l=1.075e-06 $layer=LI1_cond $X=1.48 $Y=0.875
+ $X2=1.48 $Y2=1.95
r118 13 44 38.6549 $w=2.86e-07 $l=1.90526e-07 $layer=POLY_cond $X=3.785 $Y=1.3
+ $X2=3.73 $Y2=1.465
r119 13 15 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.785 $Y=1.3
+ $X2=3.785 $Y2=0.74
r120 10 44 61.4066 $w=2.86e-07 $l=3.21714e-07 $layer=POLY_cond $X=3.775 $Y=1.765
+ $X2=3.73 $Y2=1.465
r121 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.775 $Y=1.765
+ $X2=3.775 $Y2=2.4
r122 3 39 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.335
+ $Y=1.84 $X2=1.48 $Y2=1.985
r123 3 21 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.335
+ $Y=1.84 $X2=1.48 $Y2=2.695
r124 2 31 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=2.785
+ $Y=0.37 $X2=2.925 $Y2=0.645
r125 1 37 182 $w=1.7e-07 $l=4.0398e-07 $layer=licon1_NDIFF $count=1 $X=1.14
+ $Y=0.37 $X2=1.28 $Y2=0.71
r126 1 25 182 $w=1.7e-07 $l=9.39747e-07 $layer=licon1_NDIFF $count=1 $X=1.14
+ $Y=0.37 $X2=1.925 $Y2=0.71
.ends

.subckt PM_SKY130_FD_SC_LS__OR4B_1%VPWR 1 2 9 13 18 19 20 22 35 36 39
r41 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r42 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r43 33 36 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r44 32 33 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r45 30 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r46 29 32 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=3.12 $Y2=3.33
r47 29 30 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r48 27 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.95 $Y=3.33
+ $X2=0.785 $Y2=3.33
r49 27 29 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.95 $Y=3.33 $X2=1.2
+ $Y2=3.33
r50 25 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r51 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r52 22 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.62 $Y=3.33
+ $X2=0.785 $Y2=3.33
r53 22 24 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=0.62 $Y=3.33
+ $X2=0.24 $Y2=3.33
r54 20 33 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r55 20 30 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.2 $Y2=3.33
r56 18 32 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=3.335 $Y=3.33
+ $X2=3.12 $Y2=3.33
r57 18 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.335 $Y=3.33
+ $X2=3.5 $Y2=3.33
r58 17 35 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=3.665 $Y=3.33
+ $X2=4.08 $Y2=3.33
r59 17 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.665 $Y=3.33
+ $X2=3.5 $Y2=3.33
r60 13 16 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=3.5 $Y=2.455 $X2=3.5
+ $Y2=2.815
r61 11 19 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.5 $Y=3.245 $X2=3.5
+ $Y2=3.33
r62 11 16 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.5 $Y=3.245 $X2=3.5
+ $Y2=2.815
r63 7 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.785 $Y=3.245
+ $X2=0.785 $Y2=3.33
r64 7 9 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=0.785 $Y=3.245
+ $X2=0.785 $Y2=2.455
r65 2 16 600 $w=1.7e-07 $l=1.13231e-06 $layer=licon1_PDIFF $count=1 $X=3.16
+ $Y=1.84 $X2=3.5 $Y2=2.815
r66 2 13 600 $w=1.7e-07 $l=7.66371e-07 $layer=licon1_PDIFF $count=1 $X=3.16
+ $Y=1.84 $X2=3.5 $Y2=2.455
r67 1 9 300 $w=1.7e-07 $l=4.2335e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=2.12 $X2=0.785 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_LS__OR4B_1%X 1 2 9 13 14 15 16 23 33
c26 14 0 1.19108e-19 $X=3.995 $Y=1.95
c27 13 0 7.34258e-20 $X=4.035 $Y=1.13
r28 21 23 0.432166 $w=3.98e-07 $l=1.5e-08 $layer=LI1_cond $X=4.035 $Y=2.02
+ $X2=4.035 $Y2=2.035
r29 15 16 10.6601 $w=3.98e-07 $l=3.7e-07 $layer=LI1_cond $X=4.035 $Y=2.405
+ $X2=4.035 $Y2=2.775
r30 14 21 1.00839 $w=3.98e-07 $l=3.5e-08 $layer=LI1_cond $X=4.035 $Y=1.985
+ $X2=4.035 $Y2=2.02
r31 14 33 8.64761 $w=3.98e-07 $l=1.65e-07 $layer=LI1_cond $X=4.035 $Y=1.985
+ $X2=4.035 $Y2=1.82
r32 14 15 9.65171 $w=3.98e-07 $l=3.35e-07 $layer=LI1_cond $X=4.035 $Y=2.07
+ $X2=4.035 $Y2=2.405
r33 14 23 1.00839 $w=3.98e-07 $l=3.5e-08 $layer=LI1_cond $X=4.035 $Y=2.07
+ $X2=4.035 $Y2=2.035
r34 13 33 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.15 $Y=1.13 $X2=4.15
+ $Y2=1.82
r35 7 13 9.656 $w=3.98e-07 $l=2e-07 $layer=LI1_cond $X=4.035 $Y=0.93 $X2=4.035
+ $Y2=1.13
r36 7 9 11.9566 $w=3.98e-07 $l=4.15e-07 $layer=LI1_cond $X=4.035 $Y=0.93
+ $X2=4.035 $Y2=0.515
r37 2 14 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=3.85
+ $Y=1.84 $X2=4 $Y2=1.985
r38 2 16 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=3.85
+ $Y=1.84 $X2=4 $Y2=2.815
r39 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.86
+ $Y=0.37 $X2=4 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__OR4B_1%VGND 1 2 3 12 16 20 23 24 26 27 28 30 46 47
+ 50
r54 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r55 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r56 44 47 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r57 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r58 38 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r59 37 40 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r60 37 38 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r61 35 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=0.78
+ $Y2=0
r62 35 37 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=1.2
+ $Y2=0
r63 33 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r64 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r65 30 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.78
+ $Y2=0
r66 30 32 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.24
+ $Y2=0
r67 28 44 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r68 28 38 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.2
+ $Y2=0
r69 28 40 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r70 26 43 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.295 $Y=0 $X2=3.12
+ $Y2=0
r71 26 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.295 $Y=0 $X2=3.46
+ $Y2=0
r72 25 46 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=3.625 $Y=0 $X2=4.08
+ $Y2=0
r73 25 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.625 $Y=0 $X2=3.46
+ $Y2=0
r74 23 40 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=2.26 $Y=0 $X2=2.16
+ $Y2=0
r75 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.26 $Y=0 $X2=2.425
+ $Y2=0
r76 22 43 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=2.59 $Y=0 $X2=3.12
+ $Y2=0
r77 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.59 $Y=0 $X2=2.425
+ $Y2=0
r78 18 27 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.46 $Y=0.085
+ $X2=3.46 $Y2=0
r79 18 20 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=3.46 $Y=0.085
+ $X2=3.46 $Y2=0.595
r80 14 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.425 $Y=0.085
+ $X2=2.425 $Y2=0
r81 14 16 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=2.425 $Y=0.085
+ $X2=2.425 $Y2=0.61
r82 10 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=0.085
+ $X2=0.78 $Y2=0
r83 10 12 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=0.78 $Y=0.085
+ $X2=0.78 $Y2=0.645
r84 3 20 182 $w=1.7e-07 $l=3.39338e-07 $layer=licon1_NDIFF $count=1 $X=3.215
+ $Y=0.37 $X2=3.46 $Y2=0.595
r85 2 16 182 $w=1.7e-07 $l=3.28634e-07 $layer=licon1_NDIFF $count=1 $X=2.215
+ $Y=0.37 $X2=2.425 $Y2=0.61
r86 1 12 182 $w=1.7e-07 $l=3.65205e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.78 $Y2=0.645
.ends

