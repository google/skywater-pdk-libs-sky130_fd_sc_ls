* NGSPICE file created from sky130_fd_sc_ls__diode_2.ext - technology: sky130A

.subckt sky130_fd_sc_ls__diode_2 DIODE VGND VNB VPB VPWR
D0 VNB DIODE ndiode p=7.32e+06u a=6.417e+11p
.ends

