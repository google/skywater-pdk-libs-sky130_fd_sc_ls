* File: sky130_fd_sc_ls__and2_4.pex.spice
* Created: Fri Aug 28 13:02:54 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__AND2_4%A_83_269# 1 2 3 10 12 13 15 16 18 19 21 22 24
+ 25 27 28 30 31 33 34 43 44 45 48 50 54 56 57 59 62 64 65 74
c147 74 0 1.03487e-19 $X=1.875 $Y=1.555
c148 34 0 9.81068e-20 $X=1.885 $Y=1.51
c149 31 0 4.21777e-20 $X=1.935 $Y=1.345
c150 28 0 4.53088e-20 $X=1.875 $Y=1.765
r151 74 75 7.81622 $w=3.7e-07 $l=6e-08 $layer=POLY_cond $X=1.875 $Y=1.555
+ $X2=1.935 $Y2=1.555
r152 71 72 6.51351 $w=3.7e-07 $l=5e-08 $layer=POLY_cond $X=1.355 $Y=1.555
+ $X2=1.405 $Y2=1.555
r153 68 69 3.90811 $w=3.7e-07 $l=3e-08 $layer=POLY_cond $X=0.925 $Y=1.555
+ $X2=0.955 $Y2=1.555
r154 67 68 54.7135 $w=3.7e-07 $l=4.2e-07 $layer=POLY_cond $X=0.505 $Y=1.555
+ $X2=0.925 $Y2=1.555
r155 66 67 1.3027 $w=3.7e-07 $l=1e-08 $layer=POLY_cond $X=0.495 $Y=1.555
+ $X2=0.505 $Y2=1.555
r156 60 65 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.585 $Y=2.12
+ $X2=3.585 $Y2=2.035
r157 60 62 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=3.585 $Y=2.12
+ $X2=3.585 $Y2=2.19
r158 59 65 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.585 $Y=1.95
+ $X2=3.585 $Y2=2.035
r159 58 59 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.585 $Y=1.28
+ $X2=3.585 $Y2=1.95
r160 56 58 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.5 $Y=1.195
+ $X2=3.585 $Y2=1.28
r161 56 57 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.5 $Y=1.195
+ $X2=3.325 $Y2=1.195
r162 52 57 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.16 $Y=1.11
+ $X2=3.325 $Y2=1.195
r163 52 54 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=3.16 $Y=1.11
+ $X2=3.16 $Y2=0.72
r164 51 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.8 $Y=2.035
+ $X2=2.635 $Y2=2.035
r165 50 65 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.5 $Y=2.035
+ $X2=3.585 $Y2=2.035
r166 50 51 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=3.5 $Y=2.035 $X2=2.8
+ $Y2=2.035
r167 46 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.635 $Y=2.12
+ $X2=2.635 $Y2=2.035
r168 46 48 2.44458 $w=3.28e-07 $l=7e-08 $layer=LI1_cond $X=2.635 $Y=2.12
+ $X2=2.635 $Y2=2.19
r169 44 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.47 $Y=2.035
+ $X2=2.635 $Y2=2.035
r170 44 45 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=2.47 $Y=2.035
+ $X2=2.055 $Y2=2.035
r171 43 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.97 $Y=1.95
+ $X2=2.055 $Y2=2.035
r172 42 43 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.97 $Y=1.675
+ $X2=1.97 $Y2=1.95
r173 41 74 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=1.85 $Y=1.555
+ $X2=1.875 $Y2=1.555
r174 41 72 57.9703 $w=3.7e-07 $l=4.45e-07 $layer=POLY_cond $X=1.85 $Y=1.555
+ $X2=1.405 $Y2=1.555
r175 40 41 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.85
+ $Y=1.51 $X2=1.85 $Y2=1.51
r176 37 71 24.1 $w=3.7e-07 $l=1.85e-07 $layer=POLY_cond $X=1.17 $Y=1.555
+ $X2=1.355 $Y2=1.555
r177 37 69 28.0081 $w=3.7e-07 $l=2.15e-07 $layer=POLY_cond $X=1.17 $Y=1.555
+ $X2=0.955 $Y2=1.555
r178 36 40 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.17 $Y=1.51
+ $X2=1.85 $Y2=1.51
r179 36 37 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.17
+ $Y=1.51 $X2=1.17 $Y2=1.51
r180 34 42 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.885 $Y=1.51
+ $X2=1.97 $Y2=1.675
r181 34 40 1.22229 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=1.885 $Y=1.51
+ $X2=1.85 $Y2=1.51
r182 31 75 23.9667 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=1.935 $Y=1.345
+ $X2=1.935 $Y2=1.555
r183 31 33 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.935 $Y=1.345
+ $X2=1.935 $Y2=0.865
r184 28 74 23.9667 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=1.875 $Y=1.765
+ $X2=1.875 $Y2=1.555
r185 28 30 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.875 $Y=1.765
+ $X2=1.875 $Y2=2.4
r186 25 72 23.9667 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=1.405 $Y=1.765
+ $X2=1.405 $Y2=1.555
r187 25 27 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.405 $Y=1.765
+ $X2=1.405 $Y2=2.4
r188 22 71 23.9667 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=1.355 $Y=1.345
+ $X2=1.355 $Y2=1.555
r189 22 24 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.355 $Y=1.345
+ $X2=1.355 $Y2=0.865
r190 19 69 23.9667 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=0.955 $Y=1.765
+ $X2=0.955 $Y2=1.555
r191 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.955 $Y=1.765
+ $X2=0.955 $Y2=2.4
r192 16 68 23.9667 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=0.925 $Y=1.345
+ $X2=0.925 $Y2=1.555
r193 16 18 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.925 $Y=1.345
+ $X2=0.925 $Y2=0.865
r194 13 67 23.9667 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=1.555
r195 13 15 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.4
r196 10 66 23.9667 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=0.495 $Y=1.345
+ $X2=0.495 $Y2=1.555
r197 10 12 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.495 $Y=1.345
+ $X2=0.495 $Y2=0.865
r198 3 62 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=3.435
+ $Y=2.045 $X2=3.585 $Y2=2.19
r199 2 48 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=2.485
+ $Y=2.045 $X2=2.635 $Y2=2.19
r200 1 54 91 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=2 $X=2.975
+ $Y=0.595 $X2=3.16 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_LS__AND2_4%A 1 3 6 8 10 13 15 22
c48 15 0 2.42266e-19 $X=3.12 $Y=1.665
r49 22 23 1.46061 $w=4.95e-07 $l=1.5e-08 $layer=POLY_cond $X=3.36 $Y=1.71
+ $X2=3.375 $Y2=1.71
r50 20 22 26.2909 $w=4.95e-07 $l=2.7e-07 $layer=POLY_cond $X=3.09 $Y=1.71
+ $X2=3.36 $Y2=1.71
r51 18 20 18.501 $w=4.95e-07 $l=1.9e-07 $layer=POLY_cond $X=2.9 $Y=1.71 $X2=3.09
+ $Y2=1.71
r52 17 18 1.46061 $w=4.95e-07 $l=1.5e-08 $layer=POLY_cond $X=2.885 $Y=1.71
+ $X2=2.9 $Y2=1.71
r53 15 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.09
+ $Y=1.615 $X2=3.09 $Y2=1.615
r54 11 23 31.1543 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=3.375 $Y=1.45
+ $X2=3.375 $Y2=1.71
r55 11 13 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=3.375 $Y=1.45
+ $X2=3.375 $Y2=0.915
r56 8 22 31.1543 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=3.36 $Y=1.97 $X2=3.36
+ $Y2=1.71
r57 8 10 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=3.36 $Y=1.97 $X2=3.36
+ $Y2=2.465
r58 4 18 31.1543 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=2.9 $Y=1.45 $X2=2.9
+ $Y2=1.71
r59 4 6 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=2.9 $Y=1.45 $X2=2.9
+ $Y2=0.915
r60 1 17 31.1543 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=2.885 $Y=1.97
+ $X2=2.885 $Y2=1.71
r61 1 3 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.885 $Y=1.97
+ $X2=2.885 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LS__AND2_4%B 2 3 5 9 10 11 12 13 14 16 20 22 25
c75 25 0 1.68219e-19 $X=2.42 $Y=1.51
c76 22 0 4.53088e-20 $X=2.64 $Y=1.665
c77 2 0 7.40463e-20 $X=2.41 $Y=1.88
r78 25 28 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.42 $Y=1.51
+ $X2=2.42 $Y2=1.675
r79 25 27 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.42 $Y=1.51
+ $X2=2.42 $Y2=1.345
r80 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.42
+ $Y=1.51 $X2=2.42 $Y2=1.51
r81 22 26 5.82845 $w=4.33e-07 $l=2.2e-07 $layer=LI1_cond $X=2.64 $Y=1.562
+ $X2=2.42 $Y2=1.562
r82 20 21 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.825 $Y=0.915
+ $X2=3.825 $Y2=1.31
r83 17 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.825 $Y=0.255
+ $X2=3.825 $Y2=0.915
r84 14 16 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=3.81 $Y=1.97
+ $X2=3.81 $Y2=2.465
r85 13 14 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.81 $Y=1.88 $X2=3.81
+ $Y2=1.97
r86 12 21 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.81 $Y=1.4 $X2=3.81
+ $Y2=1.31
r87 12 13 186.581 $w=1.8e-07 $l=4.8e-07 $layer=POLY_cond $X=3.81 $Y=1.4 $X2=3.81
+ $Y2=1.88
r88 10 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.75 $Y=0.18
+ $X2=3.825 $Y2=0.255
r89 10 11 630.702 $w=1.5e-07 $l=1.23e-06 $layer=POLY_cond $X=3.75 $Y=0.18
+ $X2=2.52 $Y2=0.18
r90 9 27 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.445 $Y=0.915
+ $X2=2.445 $Y2=1.345
r91 6 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.445 $Y=0.255
+ $X2=2.52 $Y2=0.18
r92 6 9 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.445 $Y=0.255
+ $X2=2.445 $Y2=0.915
r93 3 5 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.41 $Y=1.97 $X2=2.41
+ $Y2=2.465
r94 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.41 $Y=1.88 $X2=2.41
+ $Y2=1.97
r95 2 28 79.6855 $w=1.8e-07 $l=2.05e-07 $layer=POLY_cond $X=2.41 $Y=1.88
+ $X2=2.41 $Y2=1.675
.ends

.subckt PM_SKY130_FD_SC_LS__AND2_4%VPWR 1 2 3 4 5 16 18 24 28 34 36 38 41 42 43
+ 49 53 58 67 70 74
c73 28 0 1.03487e-19 $X=2.1 $Y=2.455
r74 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r75 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r76 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r77 62 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r78 62 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r79 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r80 59 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.3 $Y=3.33
+ $X2=3.135 $Y2=3.33
r81 59 61 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=3.3 $Y=3.33 $X2=3.6
+ $Y2=3.33
r82 58 73 4.72267 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=3.87 $Y=3.33
+ $X2=4.095 $Y2=3.33
r83 58 61 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=3.87 $Y=3.33 $X2=3.6
+ $Y2=3.33
r84 57 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r85 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r86 54 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.265 $Y=3.33
+ $X2=2.1 $Y2=3.33
r87 54 56 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=2.265 $Y=3.33
+ $X2=2.64 $Y2=3.33
r88 53 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.97 $Y=3.33
+ $X2=3.135 $Y2=3.33
r89 53 56 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.97 $Y=3.33
+ $X2=2.64 $Y2=3.33
r90 51 52 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r91 49 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.935 $Y=3.33
+ $X2=2.1 $Y2=3.33
r92 49 51 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.935 $Y=3.33
+ $X2=1.68 $Y2=3.33
r93 48 52 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r94 48 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r95 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r96 45 64 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.182 $Y2=3.33
r97 45 47 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.72 $Y2=3.33
r98 43 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r99 43 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r100 43 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r101 41 47 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.015 $Y=3.33
+ $X2=0.72 $Y2=3.33
r102 41 42 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.015 $Y=3.33
+ $X2=1.14 $Y2=3.33
r103 40 51 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=1.265 $Y=3.33
+ $X2=1.68 $Y2=3.33
r104 40 42 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.265 $Y=3.33
+ $X2=1.14 $Y2=3.33
r105 36 73 3.0435 $w=3.3e-07 $l=1.11018e-07 $layer=LI1_cond $X=4.035 $Y=3.245
+ $X2=4.095 $Y2=3.33
r106 36 38 36.8433 $w=3.28e-07 $l=1.055e-06 $layer=LI1_cond $X=4.035 $Y=3.245
+ $X2=4.035 $Y2=2.19
r107 32 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.135 $Y=3.245
+ $X2=3.135 $Y2=3.33
r108 32 34 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=3.135 $Y=3.245
+ $X2=3.135 $Y2=2.415
r109 28 31 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=2.1 $Y=2.455
+ $X2=2.1 $Y2=2.815
r110 26 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.1 $Y=3.245 $X2=2.1
+ $Y2=3.33
r111 26 31 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.1 $Y=3.245
+ $X2=2.1 $Y2=2.815
r112 22 42 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=3.245
+ $X2=1.14 $Y2=3.33
r113 22 24 41.2575 $w=2.48e-07 $l=8.95e-07 $layer=LI1_cond $X=1.14 $Y=3.245
+ $X2=1.14 $Y2=2.35
r114 18 21 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=0.24 $Y=1.985
+ $X2=0.24 $Y2=2.815
r115 16 64 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.182 $Y2=3.33
r116 16 21 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.24 $Y2=2.815
r117 5 38 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=3.885
+ $Y=2.045 $X2=4.035 $Y2=2.19
r118 4 34 300 $w=1.7e-07 $l=4.49055e-07 $layer=licon1_PDIFF $count=2 $X=2.96
+ $Y=2.045 $X2=3.135 $Y2=2.415
r119 3 31 600 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.95
+ $Y=1.84 $X2=2.1 $Y2=2.815
r120 3 28 600 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=1 $X=1.95
+ $Y=1.84 $X2=2.1 $Y2=2.455
r121 2 24 300 $w=1.7e-07 $l=5.80172e-07 $layer=licon1_PDIFF $count=2 $X=1.03
+ $Y=1.84 $X2=1.18 $Y2=2.35
r122 1 21 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r123 1 18 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_LS__AND2_4%X 1 2 3 4 15 21 23 25 27 29 33 36 39 42 48 50
c64 42 0 1.92991e-19 $X=0.635 $Y=1.58
r65 45 50 1.19218 $w=2.88e-07 $l=3e-08 $layer=LI1_cond $X=0.69 $Y=1.695 $X2=0.69
+ $Y2=1.665
r66 42 50 1.1127 $w=2.88e-07 $l=2.8e-08 $layer=LI1_cond $X=0.69 $Y=1.637
+ $X2=0.69 $Y2=1.665
r67 42 48 3.7084 $w=2.88e-07 $l=8.7e-08 $layer=LI1_cond $X=0.69 $Y=1.637
+ $X2=0.69 $Y2=1.55
r68 42 45 1.07296 $w=2.88e-07 $l=2.7e-08 $layer=LI1_cond $X=0.69 $Y=1.722
+ $X2=0.69 $Y2=1.695
r69 37 42 4.88795 $w=2.88e-07 $l=1.23e-07 $layer=LI1_cond $X=0.69 $Y=1.845
+ $X2=0.69 $Y2=1.722
r70 37 39 3.351 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=1.845 $X2=0.69
+ $Y2=1.93
r71 31 33 16.8257 $w=2.48e-07 $l=3.65e-07 $layer=LI1_cond $X=1.6 $Y=1.005
+ $X2=1.6 $Y2=0.64
r72 27 41 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.59 $Y=2.015
+ $X2=1.59 $Y2=1.93
r73 27 29 36.8782 $w=2.48e-07 $l=8e-07 $layer=LI1_cond $X=1.59 $Y=2.015 $X2=1.59
+ $Y2=2.815
r74 26 39 3.18746 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=0.835 $Y=1.93
+ $X2=0.69 $Y2=1.93
r75 25 41 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.465 $Y=1.93
+ $X2=1.59 $Y2=1.93
r76 25 26 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=1.465 $Y=1.93
+ $X2=0.835 $Y2=1.93
r77 24 36 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.795 $Y=1.09
+ $X2=0.67 $Y2=1.09
r78 23 31 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.475 $Y=1.09
+ $X2=1.6 $Y2=1.005
r79 23 24 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.475 $Y=1.09
+ $X2=0.795 $Y2=1.09
r80 19 39 3.351 $w=2.8e-07 $l=8.9861e-08 $layer=LI1_cond $X=0.68 $Y=2.015
+ $X2=0.69 $Y2=1.93
r81 19 21 34.1465 $w=2.68e-07 $l=8e-07 $layer=LI1_cond $X=0.68 $Y=2.015 $X2=0.68
+ $Y2=2.815
r82 17 36 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.67 $Y=1.175
+ $X2=0.67 $Y2=1.09
r83 17 48 17.2866 $w=2.48e-07 $l=3.75e-07 $layer=LI1_cond $X=0.67 $Y=1.175
+ $X2=0.67 $Y2=1.55
r84 13 36 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.67 $Y=1.005
+ $X2=0.67 $Y2=1.09
r85 13 15 16.8257 $w=2.48e-07 $l=3.65e-07 $layer=LI1_cond $X=0.67 $Y=1.005
+ $X2=0.67 $Y2=0.64
r86 4 41 400 $w=1.7e-07 $l=2.33238e-07 $layer=licon1_PDIFF $count=1 $X=1.48
+ $Y=1.84 $X2=1.63 $Y2=2.01
r87 4 29 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.48
+ $Y=1.84 $X2=1.63 $Y2=2.815
r88 3 39 400 $w=1.7e-07 $l=2.33238e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.84 $X2=0.73 $Y2=2.01
r89 3 21 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.84 $X2=0.73 $Y2=2.815
r90 2 33 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=1.43
+ $Y=0.495 $X2=1.64 $Y2=0.64
r91 1 36 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.495 $X2=0.71 $Y2=1.09
r92 1 15 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.495 $X2=0.71 $Y2=0.64
.ends

.subckt PM_SKY130_FD_SC_LS__AND2_4%VGND 1 2 3 4 13 15 19 23 25 27 29 31 36 41 53
+ 56 60
r60 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r61 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r62 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r63 48 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r64 47 48 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r65 45 48 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r66 44 47 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r67 44 45 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r68 42 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.315 $Y=0 $X2=2.15
+ $Y2=0
r69 42 44 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.315 $Y=0 $X2=2.64
+ $Y2=0
r70 41 59 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=3.875 $Y=0 $X2=4.097
+ $Y2=0
r71 41 47 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3.875 $Y=0 $X2=3.6
+ $Y2=0
r72 40 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r73 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r74 37 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.305 $Y=0 $X2=1.14
+ $Y2=0
r75 37 39 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.305 $Y=0 $X2=1.68
+ $Y2=0
r76 36 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.985 $Y=0 $X2=2.15
+ $Y2=0
r77 36 39 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.985 $Y=0 $X2=1.68
+ $Y2=0
r78 35 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r79 35 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r80 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r81 32 50 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=0 $X2=0.182
+ $Y2=0
r82 32 34 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=0 $X2=0.72
+ $Y2=0
r83 31 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.975 $Y=0 $X2=1.14
+ $Y2=0
r84 31 34 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.975 $Y=0 $X2=0.72
+ $Y2=0
r85 29 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r86 29 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r87 29 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r88 25 59 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=4.04 $Y=0.085
+ $X2=4.097 $Y2=0
r89 25 27 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=4.04 $Y=0.085
+ $X2=4.04 $Y2=0.74
r90 21 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.15 $Y=0.085
+ $X2=2.15 $Y2=0
r91 21 23 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=2.15 $Y=0.085
+ $X2=2.15 $Y2=0.7
r92 17 53 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=0.085
+ $X2=1.14 $Y2=0
r93 17 19 20.4297 $w=3.28e-07 $l=5.85e-07 $layer=LI1_cond $X=1.14 $Y=0.085
+ $X2=1.14 $Y2=0.67
r94 13 50 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.182 $Y2=0
r95 13 15 25.5842 $w=2.48e-07 $l=5.55e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.24 $Y2=0.64
r96 4 27 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.9
+ $Y=0.595 $X2=4.04 $Y2=0.74
r97 3 23 91 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=2 $X=2.01
+ $Y=0.495 $X2=2.15 $Y2=0.7
r98 2 19 182 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=1 $X=1
+ $Y=0.495 $X2=1.14 $Y2=0.67
r99 1 15 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.495 $X2=0.28 $Y2=0.64
.ends

.subckt PM_SKY130_FD_SC_LS__AND2_4%A_504_119# 1 2 9 11 12 15
c29 12 0 4.21777e-20 $X=2.825 $Y=0.34
r30 13 15 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=3.59 $Y=0.425
+ $X2=3.59 $Y2=0.755
r31 11 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.505 $Y=0.34
+ $X2=3.59 $Y2=0.425
r32 11 12 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.505 $Y=0.34
+ $X2=2.825 $Y2=0.34
r33 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.66 $Y=0.425
+ $X2=2.825 $Y2=0.34
r34 7 9 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.66 $Y=0.425
+ $X2=2.66 $Y2=0.72
r35 2 15 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=3.45
+ $Y=0.595 $X2=3.59 $Y2=0.755
r36 1 9 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=2.52
+ $Y=0.595 $X2=2.66 $Y2=0.72
.ends

