* File: sky130_fd_sc_ls__o2bb2a_1.spice
* Created: Fri Aug 28 13:49:51 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__o2bb2a_1.pex.spice"
.subckt sky130_fd_sc_ls__o2bb2a_1  VNB VPB A1_N A2_N B2 B1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* B1	B1
* B2	B2
* A2_N	A2_N
* A1_N	A1_N
* VPB	VPB
* VNB	VNB
MM1002 N_VGND_M1002_d N_A_83_260#_M1002_g N_X_M1002_s VNB NSHORT L=0.15 W=0.74
+ AD=0.202642 AS=0.2109 PD=1.36739 PS=2.05 NRD=19.044 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1003 A_253_94# N_A1_N_M1003_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.64
+ AD=0.0768 AS=0.175258 PD=0.88 PS=1.18261 NRD=12.18 NRS=26.244 M=1 R=4.26667
+ SA=75000.9 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1004 N_A_233_384#_M1004_d N_A2_N_M1004_g A_253_94# VNB NSHORT L=0.15 W=0.64
+ AD=0.1824 AS=0.0768 PD=1.85 PS=0.88 NRD=0 NRS=12.18 M=1 R=4.26667 SA=75001.3
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1005 N_A_588_74#_M1005_d N_A_233_384#_M1005_g N_A_83_260#_M1005_s VNB NSHORT
+ L=0.15 W=0.64 AD=0.0896 AS=0.1824 PD=0.92 PS=1.85 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1011 N_VGND_M1011_d N_B2_M1011_g N_A_588_74#_M1005_d VNB NSHORT L=0.15 W=0.64
+ AD=0.1216 AS=0.0896 PD=1.02 PS=0.92 NRD=13.116 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75000.7 A=0.096 P=1.58 MULT=1
MM1010 N_A_588_74#_M1010_d N_B1_M1010_g N_VGND_M1011_d VNB NSHORT L=0.15 W=0.64
+ AD=0.1824 AS=0.1216 PD=1.85 PS=1.02 NRD=0 NRS=5.616 M=1 R=4.26667 SA=75001.2
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1007 N_VPWR_M1007_d N_A_83_260#_M1007_g N_X_M1007_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.260343 AS=0.3304 PD=1.77714 PS=2.83 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75002.7 A=0.168 P=2.54 MULT=1
MM1000 N_A_233_384#_M1000_d N_A1_N_M1000_g N_VPWR_M1007_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.1491 AS=0.195257 PD=1.195 PS=1.33286 NRD=2.3443 NRS=22.655 M=1
+ R=5.6 SA=75000.8 SB=75002.9 A=0.126 P=1.98 MULT=1
MM1001 N_VPWR_M1001_d N_A2_N_M1001_g N_A_233_384#_M1000_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.4767 AS=0.1491 PD=1.975 PS=1.195 NRD=2.3443 NRS=15.2281 M=1 R=5.6
+ SA=75001.3 SB=75002.4 A=0.126 P=1.98 MULT=1
MM1008 N_A_83_260#_M1008_d N_A_233_384#_M1008_g N_VPWR_M1001_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.157409 AS=0.4767 PD=1.24174 PS=1.975 NRD=14.0658 NRS=2.3443
+ M=1 R=5.6 SA=75002.6 SB=75001.1 A=0.126 P=1.98 MULT=1
MM1009 A_693_384# N_B2_M1009_g N_A_83_260#_M1008_d VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.187391 PD=1.27 PS=1.47826 NRD=15.7403 NRS=3.9203 M=1 R=6.66667
+ SA=75002.6 SB=75000.6 A=0.15 P=2.3 MULT=1
MM1006 N_VPWR_M1006_d N_B1_M1006_g A_693_384# VPB PHIGHVT L=0.15 W=1 AD=0.295
+ AS=0.135 PD=2.59 PS=1.27 NRD=1.9503 NRS=15.7403 M=1 R=6.66667 SA=75003.1
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX12_noxref VNB VPB NWDIODE A=8.742 P=13.12
*
.include "sky130_fd_sc_ls__o2bb2a_1.pxi.spice"
*
.ends
*
*
