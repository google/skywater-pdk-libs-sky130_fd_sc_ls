* File: sky130_fd_sc_ls__sdfrtp_2.spice
* Created: Fri Aug 28 14:03:15 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__sdfrtp_2.pex.spice"
.subckt sky130_fd_sc_ls__sdfrtp_2  VNB VPB SCE D SCD CLK RESET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* RESET_B	RESET_B
* CLK	CLK
* SCD	SCD
* D	D
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1031 N_VGND_M1031_d N_SCE_M1031_g N_A_27_74#_M1031_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.1197 PD=1.41 PS=1.41 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1005 noxref_25 N_A_27_74#_M1005_g N_noxref_24_M1005_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.3 A=0.063 P=1.14 MULT=1
MM1006 N_A_390_81#_M1006_d N_D_M1006_g noxref_25 VNB NSHORT L=0.15 W=0.42
+ AD=0.13125 AS=0.0504 PD=1.045 PS=0.66 NRD=98.568 NRS=18.564 M=1 R=2.8
+ SA=75000.6 SB=75001.9 A=0.063 P=1.14 MULT=1
MM1026 noxref_26 N_SCE_M1026_g N_A_390_81#_M1006_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.13125 PD=0.66 PS=1.045 NRD=18.564 NRS=0 M=1 R=2.8 SA=75001.4
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1011 N_noxref_24_M1011_d N_SCD_M1011_g noxref_26 VNB NSHORT L=0.15 W=0.42
+ AD=0.0651 AS=0.0504 PD=0.73 PS=0.66 NRD=5.712 NRS=18.564 M=1 R=2.8 SA=75001.8
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1036 N_VGND_M1036_d N_RESET_B_M1036_g N_noxref_24_M1011_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1386 AS=0.0651 PD=1.5 PS=0.73 NRD=12.852 NRS=2.856 M=1 R=2.8
+ SA=75002.2 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1029 N_VGND_M1029_d N_CLK_M1029_g N_A_835_98#_M1029_s VNB NSHORT L=0.15 W=0.74
+ AD=0.166125 AS=0.2619 PD=1.285 PS=2.38 NRD=10.536 NRS=10.536 M=1 R=4.93333
+ SA=75000.2 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1032 N_A_1034_392#_M1032_d N_A_835_98#_M1032_g N_VGND_M1029_d VNB NSHORT
+ L=0.15 W=0.74 AD=0.1961 AS=0.166125 PD=2.01 PS=1.285 NRD=0 NRS=10.536 M=1
+ R=4.93333 SA=75000.8 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1034 N_A_1234_119#_M1034_d N_A_835_98#_M1034_g N_A_390_81#_M1034_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75004.3 A=0.063 P=1.14 MULT=1
MM1000 A_1320_119# N_A_1034_392#_M1000_g N_A_1234_119#_M1034_d VNB NSHORT L=0.15
+ W=0.42 AD=0.04935 AS=0.0588 PD=0.655 PS=0.7 NRD=17.856 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75003.8 A=0.063 P=1.14 MULT=1
MM1019 A_1397_119# N_A_1367_93#_M1019_g A_1320_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.04935 PD=0.66 PS=0.655 NRD=18.564 NRS=17.856 M=1 R=2.8 SA=75001
+ SB=75003.5 A=0.063 P=1.14 MULT=1
MM1009 N_VGND_M1009_d N_RESET_B_M1009_g A_1397_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.276584 AS=0.0504 PD=1.46276 PS=0.66 NRD=172.428 NRS=18.564 M=1 R=2.8
+ SA=75001.4 SB=75003.1 A=0.063 P=1.14 MULT=1
MM1035 N_A_1367_93#_M1035_d N_A_1234_119#_M1035_g N_VGND_M1009_d VNB NSHORT
+ L=0.15 W=0.74 AD=0.13135 AS=0.487316 PD=1.095 PS=2.57724 NRD=0 NRS=97.86 M=1
+ R=4.93333 SA=75001.8 SB=75002.1 A=0.111 P=1.78 MULT=1
MM1016 N_A_1824_74#_M1016_d N_A_1034_392#_M1016_g N_A_1367_93#_M1035_d VNB
+ NSHORT L=0.15 W=0.74 AD=0.351117 AS=0.13135 PD=2.3731 PS=1.095 NRD=54.324
+ NRS=12.156 M=1 R=4.93333 SA=75002.3 SB=75001.6 A=0.111 P=1.78 MULT=1
MM1002 A_2078_74# N_A_835_98#_M1002_g N_A_1824_74#_M1016_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.199283 PD=0.66 PS=1.3469 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75003.5 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_A_2082_446#_M1003_g A_2078_74# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0504 PD=0.7 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75003.9
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1014 A_2242_74# N_RESET_B_M1014_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75004.3
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1007 N_A_2082_446#_M1007_d N_A_1824_74#_M1007_g A_2242_74# VNB NSHORT L=0.15
+ W=0.42 AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8
+ SA=75004.7 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1021 N_A_2492_392#_M1021_d N_A_1824_74#_M1021_g N_VGND_M1021_s VNB NSHORT
+ L=0.15 W=0.64 AD=0.1824 AS=0.1824 PD=1.85 PS=1.85 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1023 N_VGND_M1023_d N_A_2492_392#_M1023_g N_Q_M1023_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1041 N_VGND_M1041_d N_A_2492_392#_M1041_g N_Q_M1023_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1022 N_VPWR_M1022_d N_SCE_M1022_g N_A_27_74#_M1022_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.3104 AS=0.1888 PD=1.61 PS=1.87 NRD=18.4589 NRS=3.0732 M=1 R=4.26667
+ SA=75000.2 SB=75003.3 A=0.096 P=1.58 MULT=1
MM1025 A_340_464# N_SCE_M1025_g N_VPWR_M1022_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0864 AS=0.3104 PD=0.91 PS=1.61 NRD=24.625 NRS=3.0732 M=1 R=4.26667
+ SA=75001.3 SB=75002.2 A=0.096 P=1.58 MULT=1
MM1004 N_A_390_81#_M1004_d N_D_M1004_g A_340_464# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0928 AS=0.0864 PD=0.93 PS=0.91 NRD=0 NRS=24.625 M=1 R=4.26667 SA=75001.8
+ SB=75001.8 A=0.096 P=1.58 MULT=1
MM1017 A_512_464# N_A_27_74#_M1017_g N_A_390_81#_M1004_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.128 AS=0.0928 PD=1.04 PS=0.93 NRD=44.6205 NRS=3.0732 M=1 R=4.26667
+ SA=75002.2 SB=75001.3 A=0.096 P=1.58 MULT=1
MM1027 N_VPWR_M1027_d N_SCD_M1027_g A_512_464# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1344 AS=0.128 PD=1.06 PS=1.04 NRD=3.0732 NRS=44.6205 M=1 R=4.26667
+ SA=75002.8 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1039 N_A_390_81#_M1039_d N_RESET_B_M1039_g N_VPWR_M1027_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1888 AS=0.1344 PD=1.87 PS=1.06 NRD=3.0732 NRS=40.0107 M=1
+ R=4.26667 SA=75003.3 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1028 N_VPWR_M1028_d N_CLK_M1028_g N_A_835_98#_M1028_s VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.295 PD=1.3 PS=2.59 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75000.2
+ SB=75000.7 A=0.15 P=2.3 MULT=1
MM1030 N_A_1034_392#_M1030_d N_A_835_98#_M1030_g N_VPWR_M1028_d VPB PHIGHVT
+ L=0.15 W=1 AD=0.295 AS=0.15 PD=2.59 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75000.7 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1040 N_A_1234_119#_M1040_d N_A_1034_392#_M1040_g N_A_390_81#_M1040_s VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.063 AS=0.1239 PD=0.72 PS=1.43 NRD=4.6886 NRS=4.6886
+ M=1 R=2.8 SA=75000.2 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1008 A_1332_457# N_A_835_98#_M1008_g N_A_1234_119#_M1040_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.063 PD=0.63 PS=0.72 NRD=23.443 NRS=4.6886 M=1 R=2.8
+ SA=75000.7 SB=75001 A=0.063 P=1.14 MULT=1
MM1033 N_VPWR_M1033_d N_A_1367_93#_M1033_g A_1332_457# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.063 AS=0.0441 PD=0.72 PS=0.63 NRD=4.6886 NRS=23.443 M=1 R=2.8 SA=75001
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1001 N_A_1234_119#_M1001_d N_RESET_B_M1001_g N_VPWR_M1033_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1239 AS=0.063 PD=1.43 PS=0.72 NRD=4.6886 NRS=4.6886 M=1 R=2.8
+ SA=75001.5 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1015 N_A_1367_93#_M1015_d N_A_1234_119#_M1015_g N_VPWR_M1015_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.248775 AS=0.295 PD=1.565 PS=2.59 NRD=18.715 NRS=1.9503 M=1
+ R=6.66667 SA=75000.2 SB=75001.4 A=0.15 P=2.3 MULT=1
MM1018 N_A_1824_74#_M1018_d N_A_835_98#_M1018_g N_A_1367_93#_M1015_d VPB PHIGHVT
+ L=0.15 W=1 AD=0.314965 AS=0.248775 PD=2.57746 PS=1.565 NRD=1.9503 NRS=19.0302
+ M=1 R=6.66667 SA=75000.8 SB=75001.1 A=0.15 P=2.3 MULT=1
MM1037 A_2037_508# N_A_1034_392#_M1037_g N_A_1824_74#_M1018_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0504 AS=0.132285 PD=0.66 PS=1.08254 NRD=30.4759 NRS=4.6886 M=1
+ R=2.8 SA=75001.1 SB=75002.5 A=0.063 P=1.14 MULT=1
MM1038 N_VPWR_M1038_d N_A_2082_446#_M1038_g A_2037_508# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.147 AS=0.0504 PD=1.12 PS=0.66 NRD=4.6886 NRS=30.4759 M=1 R=2.8
+ SA=75001.5 SB=75002.1 A=0.063 P=1.14 MULT=1
MM1013 N_A_2082_446#_M1013_d N_RESET_B_M1013_g N_VPWR_M1038_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.063 AS=0.147 PD=0.72 PS=1.12 NRD=4.6886 NRS=28.1316 M=1 R=2.8
+ SA=75002.4 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1024 N_VPWR_M1024_d N_A_1824_74#_M1024_g N_A_2082_446#_M1013_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.113223 AS=0.063 PD=0.848873 PS=0.72 NRD=44.5417 NRS=4.6886
+ M=1 R=2.8 SA=75002.8 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1010 N_A_2492_392#_M1010_d N_A_1824_74#_M1010_g N_VPWR_M1024_d VPB PHIGHVT
+ L=0.15 W=1 AD=0.295 AS=0.269577 PD=2.59 PS=2.02113 NRD=1.9503 NRS=11.8003 M=1
+ R=6.66667 SA=75001.6 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1012 N_Q_M1012_d N_A_2492_392#_M1012_g N_VPWR_M1012_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1020 N_Q_M1012_d N_A_2492_392#_M1020_g N_VPWR_M1020_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.3864 PD=1.42 PS=2.93 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75000.7 SB=75000.3 A=0.168 P=2.54 MULT=1
DX42_noxref VNB VPB NWDIODE A=27.6463 P=33.52
c_150 VNB 0 1.61901e-19 $X=0 $Y=0
c_282 VPB 0 2.86164e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_ls__sdfrtp_2.pxi.spice"
*
.ends
*
*
