* File: sky130_fd_sc_ls__nor2b_2.pex.spice
* Created: Fri Aug 28 13:37:50 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__NOR2B_2%B_N 1 3 6 8 12
c34 8 0 1.67585e-19 $X=0.72 $Y=1.665
r35 12 14 18.075 $w=3.6e-07 $l=1.35e-07 $layer=POLY_cond $X=0.695 $Y=1.677
+ $X2=0.83 $Y2=1.677
r36 10 12 26.1083 $w=3.6e-07 $l=1.95e-07 $layer=POLY_cond $X=0.5 $Y=1.677
+ $X2=0.695 $Y2=1.677
r37 8 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.695
+ $Y=1.635 $X2=0.695 $Y2=1.635
r38 4 14 23.3057 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.83 $Y=1.47
+ $X2=0.83 $Y2=1.677
r39 4 6 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=0.83 $Y=1.47 $X2=0.83
+ $Y2=0.79
r40 1 10 23.3057 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.5 $Y=1.885 $X2=0.5
+ $Y2=1.677
r41 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.5 $Y=1.885 $X2=0.5
+ $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_LS__NOR2B_2%A_27_392# 1 2 7 9 10 12 13 15 16 18 21 25 29
+ 31 32 41
c79 16 0 1.40477e-19 $X=1.96 $Y=1.765
c80 13 0 1.68904e-19 $X=1.915 $Y=1.22
c81 10 0 1.67585e-19 $X=1.51 $Y=1.765
r82 41 42 4.85235 $w=4.47e-07 $l=4.5e-08 $layer=POLY_cond $X=1.915 $Y=1.492
+ $X2=1.96 $Y2=1.492
r83 40 41 43.6711 $w=4.47e-07 $l=4.05e-07 $layer=POLY_cond $X=1.51 $Y=1.492
+ $X2=1.915 $Y2=1.492
r84 39 40 8.08725 $w=4.47e-07 $l=7.5e-08 $layer=POLY_cond $X=1.435 $Y=1.492
+ $X2=1.51 $Y2=1.492
r85 36 39 13.4787 $w=4.47e-07 $l=1.25e-07 $layer=POLY_cond $X=1.31 $Y=1.492
+ $X2=1.435 $Y2=1.492
r86 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.31
+ $Y=1.385 $X2=1.31 $Y2=1.385
r87 32 35 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=1.31 $Y=1.215
+ $X2=1.31 $Y2=1.385
r88 30 31 5.07913 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=0.78 $Y=1.215
+ $X2=0.445 $Y2=1.215
r89 29 32 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.145 $Y=1.215
+ $X2=1.31 $Y2=1.215
r90 29 30 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.145 $Y=1.215
+ $X2=0.78 $Y2=1.215
r91 25 27 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=0.235 $Y=2.105
+ $X2=0.235 $Y2=2.815
r92 23 31 2.1225 $w=4.6e-07 $l=2.48898e-07 $layer=LI1_cond $X=0.235 $Y=1.3
+ $X2=0.445 $Y2=1.215
r93 23 25 37.1087 $w=2.48e-07 $l=8.05e-07 $layer=LI1_cond $X=0.235 $Y=1.3
+ $X2=0.235 $Y2=2.105
r94 19 31 2.1225 $w=4.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.445 $Y=1.13
+ $X2=0.445 $Y2=1.215
r95 19 21 9.19374 $w=6.68e-07 $l=5.15e-07 $layer=LI1_cond $X=0.445 $Y=1.13
+ $X2=0.445 $Y2=0.615
r96 16 42 28.6003 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=1.96 $Y=1.765
+ $X2=1.96 $Y2=1.492
r97 16 18 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.96 $Y=1.765
+ $X2=1.96 $Y2=2.4
r98 13 41 28.6003 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=1.915 $Y=1.22
+ $X2=1.915 $Y2=1.492
r99 13 15 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.915 $Y=1.22
+ $X2=1.915 $Y2=0.74
r100 10 40 28.6003 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=1.51 $Y=1.765
+ $X2=1.51 $Y2=1.492
r101 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.51 $Y=1.765
+ $X2=1.51 $Y2=2.4
r102 7 39 28.6003 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=1.435 $Y=1.22
+ $X2=1.435 $Y2=1.492
r103 7 9 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.435 $Y=1.22
+ $X2=1.435 $Y2=0.74
r104 2 27 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.275 $Y2=2.815
r105 2 25 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.275 $Y2=2.105
r106 1 21 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.47
+ $Y=0.47 $X2=0.615 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_LS__NOR2B_2%A 3 5 7 10 12 14 15 16 24
c51 24 0 1.64401e-19 $X=2.845 $Y=1.557
c52 16 0 1.40477e-19 $X=2.64 $Y=1.665
c53 12 0 1.02086e-19 $X=2.86 $Y=1.765
c54 3 0 3.68458e-20 $X=2.365 $Y=0.74
r55 24 25 1.95935 $w=3.69e-07 $l=1.5e-08 $layer=POLY_cond $X=2.845 $Y=1.557
+ $X2=2.86 $Y2=1.557
r56 22 24 50.9431 $w=3.69e-07 $l=3.9e-07 $layer=POLY_cond $X=2.455 $Y=1.557
+ $X2=2.845 $Y2=1.557
r57 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.455
+ $Y=1.515 $X2=2.455 $Y2=1.515
r58 20 22 5.87805 $w=3.69e-07 $l=4.5e-08 $layer=POLY_cond $X=2.41 $Y=1.557
+ $X2=2.455 $Y2=1.557
r59 19 20 5.87805 $w=3.69e-07 $l=4.5e-08 $layer=POLY_cond $X=2.365 $Y=1.557
+ $X2=2.41 $Y2=1.557
r60 16 23 4.95819 $w=4.28e-07 $l=1.85e-07 $layer=LI1_cond $X=2.64 $Y=1.565
+ $X2=2.455 $Y2=1.565
r61 15 23 7.90629 $w=4.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.16 $Y=1.565
+ $X2=2.455 $Y2=1.565
r62 12 25 23.9013 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.86 $Y=1.765
+ $X2=2.86 $Y2=1.557
r63 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.86 $Y=1.765
+ $X2=2.86 $Y2=2.4
r64 8 24 23.9013 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.845 $Y=1.35
+ $X2=2.845 $Y2=1.557
r65 8 10 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.845 $Y=1.35
+ $X2=2.845 $Y2=0.74
r66 5 20 23.9013 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.41 $Y=1.765
+ $X2=2.41 $Y2=1.557
r67 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.41 $Y=1.765
+ $X2=2.41 $Y2=2.4
r68 1 19 23.9013 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.365 $Y=1.35
+ $X2=2.365 $Y2=1.557
r69 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.365 $Y=1.35
+ $X2=2.365 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__NOR2B_2%VPWR 1 2 9 15 17 19 24 34 35 38 41
r42 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r43 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r44 35 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r45 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r46 32 41 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.8 $Y=3.33
+ $X2=2.675 $Y2=3.33
r47 32 34 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2.8 $Y=3.33 $X2=3.12
+ $Y2=3.33
r48 31 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r49 30 31 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r50 28 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r51 27 30 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r52 27 28 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r53 25 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.89 $Y=3.33
+ $X2=0.725 $Y2=3.33
r54 25 27 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.89 $Y=3.33 $X2=1.2
+ $Y2=3.33
r55 24 41 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.55 $Y=3.33
+ $X2=2.675 $Y2=3.33
r56 24 30 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=2.55 $Y=3.33
+ $X2=2.16 $Y2=3.33
r57 22 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r58 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r59 19 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.56 $Y=3.33
+ $X2=0.725 $Y2=3.33
r60 19 21 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.56 $Y=3.33 $X2=0.24
+ $Y2=3.33
r61 17 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r62 17 28 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r63 13 41 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.675 $Y=3.245
+ $X2=2.675 $Y2=3.33
r64 13 15 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=2.675 $Y=3.245
+ $X2=2.675 $Y2=2.455
r65 9 12 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.725 $Y=2.135
+ $X2=0.725 $Y2=2.815
r66 7 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.725 $Y=3.245
+ $X2=0.725 $Y2=3.33
r67 7 12 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.725 $Y=3.245
+ $X2=0.725 $Y2=2.815
r68 2 15 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=2.485
+ $Y=1.84 $X2=2.635 $Y2=2.455
r69 1 12 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=0.575
+ $Y=1.96 $X2=0.725 $Y2=2.815
r70 1 9 400 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=1 $X=0.575
+ $Y=1.96 $X2=0.725 $Y2=2.135
.ends

.subckt PM_SKY130_FD_SC_LS__NOR2B_2%A_228_368# 1 2 3 12 16 17 18 21 22 24 26
c49 24 0 1.67113e-19 $X=3.125 $Y=2.12
c50 16 0 1.02086e-19 $X=2.02 $Y=2.99
r51 24 31 3.1514 $w=2.5e-07 $l=1.5e-07 $layer=LI1_cond $X=3.125 $Y=2.12
+ $X2=3.125 $Y2=1.97
r52 24 26 12.9074 $w=2.48e-07 $l=2.8e-07 $layer=LI1_cond $X=3.125 $Y=2.12
+ $X2=3.125 $Y2=2.4
r53 23 29 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.35 $Y=2.035
+ $X2=2.185 $Y2=2.035
r54 22 31 3.99177 $w=1.7e-07 $l=1.5411e-07 $layer=LI1_cond $X=3 $Y=2.035
+ $X2=3.125 $Y2=1.97
r55 22 23 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=3 $Y=2.035 $X2=2.35
+ $Y2=2.035
r56 19 21 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=2.185 $Y=2.905
+ $X2=2.185 $Y2=2.815
r57 18 29 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.185 $Y=2.12
+ $X2=2.185 $Y2=2.035
r58 18 21 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=2.185 $Y=2.12
+ $X2=2.185 $Y2=2.815
r59 16 19 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.02 $Y=2.99
+ $X2=2.185 $Y2=2.905
r60 16 17 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=2.02 $Y=2.99
+ $X2=1.45 $Y2=2.99
r61 12 15 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=1.285 $Y=1.985
+ $X2=1.285 $Y2=2.815
r62 10 17 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.285 $Y=2.905
+ $X2=1.45 $Y2=2.99
r63 10 15 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=1.285 $Y=2.905
+ $X2=1.285 $Y2=2.815
r64 3 31 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.935
+ $Y=1.84 $X2=3.085 $Y2=1.985
r65 3 26 300 $w=1.7e-07 $l=6.30555e-07 $layer=licon1_PDIFF $count=2 $X=2.935
+ $Y=1.84 $X2=3.085 $Y2=2.4
r66 2 29 400 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=2.035
+ $Y=1.84 $X2=2.185 $Y2=2.035
r67 2 21 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.035
+ $Y=1.84 $X2=2.185 $Y2=2.815
r68 1 15 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=1.14
+ $Y=1.84 $X2=1.285 $Y2=2.815
r69 1 12 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.14
+ $Y=1.84 $X2=1.285 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_LS__NOR2B_2%Y 1 2 3 12 14 16 18 22 24 27 28 30
c54 30 0 3.68458e-20 $X=3.12 $Y=1.095
c55 24 0 1.67113e-19 $X=3.005 $Y=1.095
c56 16 0 1.64401e-19 $X=1.735 $Y=1.985
c57 12 0 1.68904e-19 $X=1.65 $Y=0.515
r58 28 30 10.0212 $w=2.28e-07 $l=2e-07 $layer=LI1_cond $X=3.12 $Y=1.295 $X2=3.12
+ $Y2=1.095
r59 25 27 6.31926 $w=1.95e-07 $l=1.36931e-07 $layer=LI1_cond $X=2.745 $Y=1.095
+ $X2=2.62 $Y2=1.07
r60 24 30 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=3.005 $Y=1.095
+ $X2=3.12 $Y2=1.095
r61 24 25 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=3.005 $Y=1.095
+ $X2=2.745 $Y2=1.095
r62 20 27 0.465126 $w=2.5e-07 $l=1.1e-07 $layer=LI1_cond $X=2.62 $Y=0.96
+ $X2=2.62 $Y2=1.07
r63 20 22 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=2.62 $Y=0.96
+ $X2=2.62 $Y2=0.515
r64 19 26 1.26644 $w=2.2e-07 $l=1.68e-07 $layer=LI1_cond $X=1.82 $Y=1.07
+ $X2=1.652 $Y2=1.07
r65 18 27 6.31926 $w=1.95e-07 $l=1.25e-07 $layer=LI1_cond $X=2.495 $Y=1.07
+ $X2=2.62 $Y2=1.07
r66 18 19 35.359 $w=2.18e-07 $l=6.75e-07 $layer=LI1_cond $X=2.495 $Y=1.07
+ $X2=1.82 $Y2=1.07
r67 14 26 6.50489 $w=2.41e-07 $l=1.44568e-07 $layer=LI1_cond $X=1.732 $Y=1.18
+ $X2=1.652 $Y2=1.07
r68 14 16 51.0182 $w=1.73e-07 $l=8.05e-07 $layer=LI1_cond $X=1.732 $Y=1.18
+ $X2=1.732 $Y2=1.985
r69 10 26 11.0766 $w=3.3e-07 $l=2.75998e-07 $layer=LI1_cond $X=1.65 $Y=0.795
+ $X2=1.652 $Y2=1.07
r70 10 12 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=1.65 $Y=0.795
+ $X2=1.65 $Y2=0.515
r71 3 16 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=1.585
+ $Y=1.84 $X2=1.735 $Y2=1.985
r72 2 22 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.44
+ $Y=0.37 $X2=2.58 $Y2=0.515
r73 1 12 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.51
+ $Y=0.37 $X2=1.65 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__NOR2B_2%VGND 1 2 3 12 16 18 20 22 24 29 34 40 43 47
r48 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r49 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r50 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r51 38 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r52 38 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r53 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r54 35 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.315 $Y=0 $X2=2.15
+ $Y2=0
r55 35 37 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.315 $Y=0 $X2=2.64
+ $Y2=0
r56 34 46 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=2.915 $Y=0 $X2=3.137
+ $Y2=0
r57 34 37 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.915 $Y=0 $X2=2.64
+ $Y2=0
r58 30 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.315 $Y=0 $X2=1.15
+ $Y2=0
r59 30 32 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.315 $Y=0 $X2=1.68
+ $Y2=0
r60 29 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.985 $Y=0 $X2=2.15
+ $Y2=0
r61 29 32 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.985 $Y=0 $X2=1.68
+ $Y2=0
r62 27 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r63 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r64 24 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.985 $Y=0 $X2=1.15
+ $Y2=0
r65 24 26 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.985 $Y=0 $X2=0.72
+ $Y2=0
r66 22 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r67 22 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r68 22 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r69 18 46 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=3.08 $Y=0.085
+ $X2=3.137 $Y2=0
r70 18 20 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=3.08 $Y=0.085
+ $X2=3.08 $Y2=0.675
r71 14 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.15 $Y=0.085
+ $X2=2.15 $Y2=0
r72 14 16 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=2.15 $Y=0.085
+ $X2=2.15 $Y2=0.625
r73 10 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.15 $Y=0.085
+ $X2=1.15 $Y2=0
r74 10 12 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=1.15 $Y=0.085
+ $X2=1.15 $Y2=0.535
r75 3 20 182 $w=1.7e-07 $l=3.76597e-07 $layer=licon1_NDIFF $count=1 $X=2.92
+ $Y=0.37 $X2=3.08 $Y2=0.675
r76 2 16 182 $w=1.7e-07 $l=3.25308e-07 $layer=licon1_NDIFF $count=1 $X=1.99
+ $Y=0.37 $X2=2.15 $Y2=0.625
r77 1 12 91 $w=1.7e-07 $l=2.7559e-07 $layer=licon1_NDIFF $count=2 $X=0.905
+ $Y=0.47 $X2=1.15 $Y2=0.535
.ends

