# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ls__o221a_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ls__o221a_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.680000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.925000 1.350000 5.320000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.365000 1.445000 4.695000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005000 1.445000 4.195000 1.780000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.445000 2.755000 1.780000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.445000 0.890000 1.780000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  1.235700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.735000 0.475000 5.985000 1.010000 ;
        RECT 5.735000 1.010000 7.065000 1.180000 ;
        RECT 5.830000 1.850000 7.115000 2.020000 ;
        RECT 5.830000 2.020000 6.160000 2.980000 ;
        RECT 6.735000 0.475000 7.065000 1.010000 ;
        RECT 6.785000 1.180000 7.065000 1.550000 ;
        RECT 6.785000 1.550000 7.555000 1.780000 ;
        RECT 6.785000 1.780000 7.115000 1.850000 ;
        RECT 6.785000 2.020000 7.115000 2.980000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 7.680000 0.085000 ;
        RECT 3.430000  0.085000 3.760000 0.935000 ;
        RECT 4.295000  0.085000 4.625000 0.840000 ;
        RECT 5.235000  0.085000 5.565000 1.180000 ;
        RECT 6.165000  0.085000 6.565000 0.805000 ;
        RECT 7.235000  0.085000 7.565000 1.255000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
        RECT 6.395000 -0.085000 6.565000 0.085000 ;
        RECT 6.875000 -0.085000 7.045000 0.085000 ;
        RECT 7.355000 -0.085000 7.525000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.680000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 7.680000 3.415000 ;
        RECT 0.115000 1.950000 0.365000 3.245000 ;
        RECT 1.095000 2.290000 1.345000 3.245000 ;
        RECT 2.915000 2.290000 3.630000 3.245000 ;
        RECT 5.300000 2.290000 5.630000 3.245000 ;
        RECT 6.360000 2.190000 6.610000 3.245000 ;
        RECT 7.315000 1.950000 7.565000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
        RECT 6.395000 3.245000 6.565000 3.415000 ;
        RECT 6.875000 3.245000 7.045000 3.415000 ;
        RECT 7.355000 3.245000 7.525000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 7.680000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.115000 0.265000 2.305000 0.285000 ;
      RECT 0.115000 0.285000 3.170000 0.435000 ;
      RECT 0.115000 0.435000 0.365000 1.275000 ;
      RECT 0.545000 0.605000 0.795000 1.105000 ;
      RECT 0.545000 1.105000 1.230000 1.275000 ;
      RECT 0.565000 1.950000 5.660000 2.120000 ;
      RECT 0.565000 2.120000 0.895000 2.955000 ;
      RECT 0.975000 0.435000 1.305000 0.935000 ;
      RECT 1.060000 1.275000 1.230000 1.950000 ;
      RECT 1.475000 0.605000 1.805000 1.025000 ;
      RECT 1.475000 1.025000 2.740000 1.105000 ;
      RECT 1.475000 1.105000 5.055000 1.180000 ;
      RECT 1.475000 1.180000 4.115000 1.275000 ;
      RECT 1.475000 1.275000 1.805000 1.285000 ;
      RECT 1.515000 2.290000 1.845000 2.905000 ;
      RECT 1.515000 2.905000 2.745000 3.075000 ;
      RECT 1.975000 0.435000 3.170000 0.455000 ;
      RECT 1.975000 0.455000 2.305000 0.855000 ;
      RECT 2.045000 2.120000 2.215000 2.735000 ;
      RECT 2.415000 2.290000 2.745000 2.905000 ;
      RECT 2.475000 0.635000 2.670000 1.025000 ;
      RECT 2.840000 0.455000 3.170000 0.855000 ;
      RECT 3.800000 2.290000 4.130000 2.905000 ;
      RECT 3.800000 2.905000 5.130000 3.075000 ;
      RECT 3.940000 0.585000 4.115000 1.010000 ;
      RECT 3.940000 1.010000 5.055000 1.105000 ;
      RECT 4.300000 2.120000 4.630000 2.735000 ;
      RECT 4.800000 2.290000 5.130000 2.905000 ;
      RECT 4.805000 0.590000 5.055000 1.010000 ;
      RECT 5.490000 1.350000 6.615000 1.680000 ;
      RECT 5.490000 1.680000 5.660000 1.950000 ;
  END
END sky130_fd_sc_ls__o221a_4
