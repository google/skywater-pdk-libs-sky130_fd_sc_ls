* File: sky130_fd_sc_ls__decaphe_4.spice
* Created: Wed Sep  2 10:59:54 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__decaphe_4.pex.spice"
.subckt sky130_fd_sc_ls__decaphe_4  VNB VPB VGND VPWR
* 
* VPWR	VPWR
* VGND	VGND
* VPB	VPB
* VNB	VNB
MM1000 N_VGND_M1000_s N_VPWR_M1000_g N_VGND_M1000_s VNB NSHORT L=1.13 W=0.775
+ AD=0.2015 AS=0.2015 PD=2.07 PS=2.07 NRD=0 NRS=0 M=1 R=0.685841 SA=565000
+ SB=565000 A=0.87575 P=3.81 MULT=1
MM1001 N_VPWR_M1001_s N_VGND_M1001_g N_VPWR_M1001_s VPB PSHORT L=1.13 W=1.255
+ AD=0.3263 AS=0.3263 PD=3.03 PS=3.03 NRD=0 NRS=0 M=1 R=1.11062 SA=565000
+ SB=565000 A=1.41815 P=4.77 MULT=1
DX2_noxref VNB VPB NWDIODE A=4.278 P=8.32
*
.include "sky130_fd_sc_ls__decaphe_4.pxi.spice"
*
.ends
*
*
