* File: sky130_fd_sc_ls__a2111oi_1.spice
* Created: Fri Aug 28 12:48:11 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__a2111oi_1.pex.spice"
.subckt sky130_fd_sc_ls__a2111oi_1  VNB VPB D1 C1 B1 A1 A2 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A2	A2
* A1	A1
* B1	B1
* C1	C1
* D1	D1
* VPB	VPB
* VNB	VNB
MM1003 N_Y_M1003_d N_D1_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1961 PD=1.02 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75002.2 A=0.111 P=1.78 MULT=1
MM1006 N_VGND_M1006_d N_C1_M1006_g N_Y_M1003_d VNB NSHORT L=0.15 W=0.74 AD=0.185
+ AS=0.1036 PD=1.24 PS=1.02 NRD=17.832 NRS=0 M=1 R=4.93333 SA=75000.6 SB=75001.8
+ A=0.111 P=1.78 MULT=1
MM1008 N_Y_M1008_d N_B1_M1008_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.185 PD=1.02 PS=1.24 NRD=0 NRS=17.832 M=1 R=4.93333 SA=75001.3
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1002 A_461_74# N_A1_M1002_g N_Y_M1008_d VNB NSHORT L=0.15 W=0.74 AD=0.1184
+ AS=0.1036 PD=1.06 PS=1.02 NRD=17.016 NRS=0 M=1 R=4.93333 SA=75001.7 SB=75000.7
+ A=0.111 P=1.78 MULT=1
MM1001 N_VGND_M1001_d N_A2_M1001_g A_461_74# VNB NSHORT L=0.15 W=0.74 AD=0.2109
+ AS=0.1184 PD=2.05 PS=1.06 NRD=0 NRS=17.016 M=1 R=4.93333 SA=75002.2 SB=75000.2
+ A=0.111 P=1.78 MULT=1
MM1007 A_156_368# N_D1_M1007_g N_Y_M1007_s VPB PHIGHVT L=0.15 W=1.12 AD=0.1344
+ AS=0.308 PD=1.36 PS=2.79 NRD=11.426 NRS=1.7533 M=1 R=7.46667 SA=75000.2
+ SB=75002.2 A=0.168 P=2.54 MULT=1
MM1000 A_234_368# N_C1_M1000_g A_156_368# VPB PHIGHVT L=0.15 W=1.12 AD=0.2184
+ AS=0.1344 PD=1.51 PS=1.36 NRD=24.6053 NRS=11.426 M=1 R=7.46667 SA=75000.6
+ SB=75001.8 A=0.168 P=2.54 MULT=1
MM1005 N_A_342_368#_M1005_d N_B1_M1005_g A_234_368# VPB PHIGHVT L=0.15 W=1.12
+ AD=0.2184 AS=0.2184 PD=1.51 PS=1.51 NRD=5.2599 NRS=24.6053 M=1 R=7.46667
+ SA=75001.1 SB=75001.3 A=0.168 P=2.54 MULT=1
MM1009 N_VPWR_M1009_d N_A1_M1009_g N_A_342_368#_M1005_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.2184 AS=0.2184 PD=1.51 PS=1.51 NRD=5.2599 NRS=14.0658 M=1
+ R=7.46667 SA=75001.7 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1004 N_A_342_368#_M1004_d N_A2_M1004_g N_VPWR_M1009_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.308 AS=0.2184 PD=2.79 PS=1.51 NRD=1.7533 NRS=14.0658 M=1 R=7.46667
+ SA=75002.2 SB=75000.2 A=0.168 P=2.54 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9564 P=11.2
*
.include "sky130_fd_sc_ls__a2111oi_1.pxi.spice"
*
.ends
*
*
