* File: sky130_fd_sc_ls__or3b_2.pxi.spice
* Created: Fri Aug 28 13:59:01 2020
* 
x_PM_SKY130_FD_SC_LS__OR3B_2%C_N N_C_N_c_68_n N_C_N_M1007_g N_C_N_M1004_g C_N
+ N_C_N_c_70_n PM_SKY130_FD_SC_LS__OR3B_2%C_N
x_PM_SKY130_FD_SC_LS__OR3B_2%A_190_260# N_A_190_260#_M1006_d
+ N_A_190_260#_M1011_d N_A_190_260#_M1002_d N_A_190_260#_c_94_n
+ N_A_190_260#_c_109_n N_A_190_260#_M1000_g N_A_190_260#_M1003_g
+ N_A_190_260#_c_96_n N_A_190_260#_c_97_n N_A_190_260#_M1009_g
+ N_A_190_260#_M1008_g N_A_190_260#_c_99_n N_A_190_260#_c_100_n
+ N_A_190_260#_c_101_n N_A_190_260#_c_102_n N_A_190_260#_c_103_n
+ N_A_190_260#_c_104_n N_A_190_260#_c_105_n N_A_190_260#_c_111_n
+ N_A_190_260#_c_106_n N_A_190_260#_c_107_n
+ PM_SKY130_FD_SC_LS__OR3B_2%A_190_260#
x_PM_SKY130_FD_SC_LS__OR3B_2%A N_A_c_208_n N_A_M1001_g N_A_M1006_g A A
+ N_A_c_210_n PM_SKY130_FD_SC_LS__OR3B_2%A
x_PM_SKY130_FD_SC_LS__OR3B_2%B N_B_c_242_n N_B_M1010_g N_B_M1005_g B N_B_c_244_n
+ PM_SKY130_FD_SC_LS__OR3B_2%B
x_PM_SKY130_FD_SC_LS__OR3B_2%A_27_368# N_A_27_368#_M1004_s N_A_27_368#_M1007_s
+ N_A_27_368#_c_277_n N_A_27_368#_M1002_g N_A_27_368#_M1011_g
+ N_A_27_368#_c_279_n N_A_27_368#_c_306_n N_A_27_368#_c_309_n
+ N_A_27_368#_c_310_n N_A_27_368#_c_322_n N_A_27_368#_c_280_n
+ N_A_27_368#_c_285_n N_A_27_368#_c_281_n PM_SKY130_FD_SC_LS__OR3B_2%A_27_368#
x_PM_SKY130_FD_SC_LS__OR3B_2%VPWR N_VPWR_M1007_d N_VPWR_M1009_d N_VPWR_c_365_n
+ N_VPWR_c_366_n N_VPWR_c_367_n VPWR N_VPWR_c_368_n N_VPWR_c_364_n
+ N_VPWR_c_370_n N_VPWR_c_371_n PM_SKY130_FD_SC_LS__OR3B_2%VPWR
x_PM_SKY130_FD_SC_LS__OR3B_2%X N_X_M1003_d N_X_M1000_s N_X_c_403_n N_X_c_404_n
+ N_X_c_405_n X X PM_SKY130_FD_SC_LS__OR3B_2%X
x_PM_SKY130_FD_SC_LS__OR3B_2%VGND N_VGND_M1004_d N_VGND_M1008_s N_VGND_M1005_d
+ N_VGND_c_446_n N_VGND_c_447_n N_VGND_c_448_n N_VGND_c_449_n N_VGND_c_450_n
+ N_VGND_c_451_n N_VGND_c_452_n N_VGND_c_453_n VGND N_VGND_c_454_n
+ N_VGND_c_455_n N_VGND_c_456_n PM_SKY130_FD_SC_LS__OR3B_2%VGND
cc_1 VNB N_C_N_c_68_n 0.0647682f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_2 VNB N_C_N_M1004_g 0.029568f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.835
cc_3 VNB N_C_N_c_70_n 0.00652172f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_4 VNB N_A_190_260#_c_94_n 0.0113917f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_5 VNB N_A_190_260#_M1003_g 0.0217342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_A_190_260#_c_96_n 0.00863897f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_190_260#_c_97_n 0.0295183f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_190_260#_M1008_g 0.0236017f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_190_260#_c_99_n 0.00904656f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_190_260#_c_100_n 0.0089459f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_190_260#_c_101_n 0.00897658f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_190_260#_c_102_n 0.00328996f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_190_260#_c_103_n 0.00951425f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_190_260#_c_104_n 0.0272219f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_190_260#_c_105_n 0.00761269f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_190_260#_c_106_n 0.0226504f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_190_260#_c_107_n 0.0149819f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_c_208_n 0.0268186f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_19 VNB N_A_M1006_g 0.0271057f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.835
cc_20 VNB N_A_c_210_n 0.0016809f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_B_c_242_n 0.0266197f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_22 VNB N_B_M1005_g 0.0258186f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.835
cc_23 VNB N_B_c_244_n 0.0016559f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_24 VNB N_A_27_368#_c_277_n 0.0289634f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_27_368#_M1011_g 0.0311299f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_26 VNB N_A_27_368#_c_279_n 0.00523497f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.665
cc_27 VNB N_A_27_368#_c_280_n 0.00167078f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_27_368#_c_281_n 0.0293174f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VPWR_c_364_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_X_c_403_n 0.00273546f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_31 VNB N_X_c_404_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_32 VNB N_X_c_405_n 0.00422231f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_446_n 0.0111927f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_34 VNB N_VGND_c_447_n 0.019013f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_448_n 0.0166983f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_449_n 0.018099f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_450_n 0.024548f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_451_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_452_n 0.0205837f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_453_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_454_n 0.020559f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_455_n 0.247561f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_456_n 0.00980973f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VPB N_C_N_c_68_n 0.0292535f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_45 VPB N_C_N_c_70_n 0.00775819f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_46 VPB N_A_190_260#_c_94_n 7.63079e-19 $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_47 VPB N_A_190_260#_c_109_n 0.022733f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_48 VPB N_A_190_260#_c_97_n 0.0240562f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 VPB N_A_190_260#_c_111_n 0.0337914f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_A_190_260#_c_106_n 0.0300549f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_51 VPB N_A_c_208_n 0.0274487f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_52 VPB N_A_c_210_n 0.00268239f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_B_c_242_n 0.0262759f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_54 VPB N_B_c_244_n 0.00302461f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_55 VPB N_A_27_368#_c_277_n 0.0325861f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_A_27_368#_c_279_n 0.00320306f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.665
cc_57 VPB N_A_27_368#_c_280_n 0.00191406f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_A_27_368#_c_285_n 0.0346865f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_365_n 0.0165272f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_60 VPB N_VPWR_c_366_n 0.0206218f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_61 VPB N_VPWR_c_367_n 0.0148287f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_368_n 0.0552717f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_364_n 0.0885823f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_370_n 0.0274851f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_371_n 0.00834123f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_X_c_403_n 0.00152627f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_67 VPB X 0.0061934f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 N_C_N_c_68_n N_A_190_260#_c_94_n 0.00574427f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_69 N_C_N_c_68_n N_A_190_260#_c_109_n 0.0268815f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_70 N_C_N_M1004_g N_A_190_260#_M1003_g 0.0195624f $X=0.565 $Y=0.835 $X2=0
+ $Y2=0
cc_71 N_C_N_c_68_n N_A_190_260#_c_99_n 0.00597962f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_72 N_C_N_c_68_n N_A_27_368#_c_279_n 0.00959112f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_73 N_C_N_M1004_g N_A_27_368#_c_279_n 0.00652595f $X=0.565 $Y=0.835 $X2=0
+ $Y2=0
cc_74 N_C_N_c_70_n N_A_27_368#_c_279_n 0.0354724f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_75 N_C_N_c_68_n N_A_27_368#_c_285_n 0.0307333f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_76 N_C_N_c_70_n N_A_27_368#_c_285_n 0.025958f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_77 N_C_N_c_68_n N_A_27_368#_c_281_n 0.00464704f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_78 N_C_N_M1004_g N_A_27_368#_c_281_n 0.024675f $X=0.565 $Y=0.835 $X2=0 $Y2=0
cc_79 N_C_N_c_70_n N_A_27_368#_c_281_n 0.0214092f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_80 N_C_N_c_68_n N_VPWR_c_365_n 0.00343137f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_81 N_C_N_c_68_n N_VPWR_c_364_n 0.00462577f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_82 N_C_N_c_68_n N_VPWR_c_370_n 0.00393265f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_83 N_C_N_c_68_n N_X_c_403_n 5.81109e-19 $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_84 N_C_N_M1004_g N_X_c_404_n 5.95409e-19 $X=0.565 $Y=0.835 $X2=0 $Y2=0
cc_85 N_C_N_M1004_g N_X_c_405_n 2.34935e-19 $X=0.565 $Y=0.835 $X2=0 $Y2=0
cc_86 N_C_N_M1004_g N_VGND_c_446_n 0.00417177f $X=0.565 $Y=0.835 $X2=0 $Y2=0
cc_87 N_C_N_M1004_g N_VGND_c_450_n 0.00366404f $X=0.565 $Y=0.835 $X2=0 $Y2=0
cc_88 N_C_N_M1004_g N_VGND_c_455_n 0.00487769f $X=0.565 $Y=0.835 $X2=0 $Y2=0
cc_89 N_A_190_260#_c_97_n N_A_c_208_n 0.0385188f $X=1.49 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_90 N_A_190_260#_c_100_n N_A_c_208_n 0.00126003f $X=2.35 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_91 N_A_190_260#_c_101_n N_A_c_208_n 0.00172393f $X=1.795 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_92 N_A_190_260#_c_97_n N_A_M1006_g 0.00119833f $X=1.49 $Y=1.765 $X2=0 $Y2=0
cc_93 N_A_190_260#_M1008_g N_A_M1006_g 0.0147478f $X=1.505 $Y=0.74 $X2=0 $Y2=0
cc_94 N_A_190_260#_c_100_n N_A_M1006_g 0.0162422f $X=2.35 $Y=1.095 $X2=0 $Y2=0
cc_95 N_A_190_260#_c_101_n N_A_M1006_g 0.00325729f $X=1.795 $Y=1.095 $X2=0 $Y2=0
cc_96 N_A_190_260#_c_102_n N_A_M1006_g 0.00299701f $X=2.515 $Y=0.615 $X2=0 $Y2=0
cc_97 N_A_190_260#_c_97_n N_A_c_210_n 0.00424632f $X=1.49 $Y=1.765 $X2=0 $Y2=0
cc_98 N_A_190_260#_c_100_n N_A_c_210_n 0.0256551f $X=2.35 $Y=1.095 $X2=0 $Y2=0
cc_99 N_A_190_260#_c_101_n N_A_c_210_n 0.0216131f $X=1.795 $Y=1.095 $X2=0 $Y2=0
cc_100 N_A_190_260#_c_103_n N_B_c_242_n 2.7493e-19 $X=3.35 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_101 N_A_190_260#_c_105_n N_B_c_242_n 0.00109075f $X=2.515 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_102 N_A_190_260#_c_111_n N_B_c_242_n 0.00227754f $X=3.4 $Y=2.375 $X2=-0.19
+ $Y2=-0.245
cc_103 N_A_190_260#_c_102_n N_B_M1005_g 0.00798791f $X=2.515 $Y=0.615 $X2=0
+ $Y2=0
cc_104 N_A_190_260#_c_103_n N_B_M1005_g 0.0116271f $X=3.35 $Y=1.095 $X2=0 $Y2=0
cc_105 N_A_190_260#_c_104_n N_B_M1005_g 6.07993e-19 $X=3.515 $Y=0.615 $X2=0
+ $Y2=0
cc_106 N_A_190_260#_c_105_n N_B_M1005_g 0.00171282f $X=2.515 $Y=1.095 $X2=0
+ $Y2=0
cc_107 N_A_190_260#_c_103_n N_B_c_244_n 0.0121392f $X=3.35 $Y=1.095 $X2=0 $Y2=0
cc_108 N_A_190_260#_c_105_n N_B_c_244_n 0.0140411f $X=2.515 $Y=1.095 $X2=0 $Y2=0
cc_109 N_A_190_260#_c_103_n N_A_27_368#_c_277_n 9.67719e-19 $X=3.35 $Y=1.095
+ $X2=0 $Y2=0
cc_110 N_A_190_260#_c_111_n N_A_27_368#_c_277_n 0.0123558f $X=3.4 $Y=2.375 $X2=0
+ $Y2=0
cc_111 N_A_190_260#_c_106_n N_A_27_368#_c_277_n 0.0129105f $X=3.495 $Y=2.29
+ $X2=0 $Y2=0
cc_112 N_A_190_260#_c_107_n N_A_27_368#_c_277_n 3.08066e-19 $X=3.552 $Y=1.095
+ $X2=0 $Y2=0
cc_113 N_A_190_260#_c_102_n N_A_27_368#_M1011_g 6.0898e-19 $X=2.515 $Y=0.615
+ $X2=0 $Y2=0
cc_114 N_A_190_260#_c_103_n N_A_27_368#_M1011_g 0.0116271f $X=3.35 $Y=1.095
+ $X2=0 $Y2=0
cc_115 N_A_190_260#_c_104_n N_A_27_368#_M1011_g 0.00816329f $X=3.515 $Y=0.615
+ $X2=0 $Y2=0
cc_116 N_A_190_260#_c_106_n N_A_27_368#_M1011_g 0.00391901f $X=3.495 $Y=2.29
+ $X2=0 $Y2=0
cc_117 N_A_190_260#_c_107_n N_A_27_368#_M1011_g 0.00221813f $X=3.552 $Y=1.095
+ $X2=0 $Y2=0
cc_118 N_A_190_260#_c_109_n N_A_27_368#_c_279_n 0.00147603f $X=1.04 $Y=1.765
+ $X2=0 $Y2=0
cc_119 N_A_190_260#_M1003_g N_A_27_368#_c_279_n 0.00123682f $X=1.075 $Y=0.74
+ $X2=0 $Y2=0
cc_120 N_A_190_260#_c_99_n N_A_27_368#_c_279_n 0.00383029f $X=1.05 $Y=1.375
+ $X2=0 $Y2=0
cc_121 N_A_190_260#_c_109_n N_A_27_368#_c_306_n 0.0154275f $X=1.04 $Y=1.765
+ $X2=0 $Y2=0
cc_122 N_A_190_260#_c_97_n N_A_27_368#_c_306_n 0.0131964f $X=1.49 $Y=1.765 $X2=0
+ $Y2=0
cc_123 N_A_190_260#_c_111_n N_A_27_368#_c_306_n 0.00500371f $X=3.4 $Y=2.375
+ $X2=0 $Y2=0
cc_124 N_A_190_260#_c_111_n N_A_27_368#_c_309_n 7.83292e-19 $X=3.4 $Y=2.375
+ $X2=0 $Y2=0
cc_125 N_A_190_260#_M1002_d N_A_27_368#_c_310_n 0.00306998f $X=3.25 $Y=1.84
+ $X2=0 $Y2=0
cc_126 N_A_190_260#_c_111_n N_A_27_368#_c_310_n 0.0106948f $X=3.4 $Y=2.375 $X2=0
+ $Y2=0
cc_127 N_A_190_260#_c_106_n N_A_27_368#_c_310_n 0.0140566f $X=3.495 $Y=2.29
+ $X2=0 $Y2=0
cc_128 N_A_190_260#_M1002_d N_A_27_368#_c_280_n 0.00118548f $X=3.25 $Y=1.84
+ $X2=0 $Y2=0
cc_129 N_A_190_260#_c_103_n N_A_27_368#_c_280_n 0.0205962f $X=3.35 $Y=1.095
+ $X2=0 $Y2=0
cc_130 N_A_190_260#_c_106_n N_A_27_368#_c_280_n 0.0458137f $X=3.495 $Y=2.29
+ $X2=0 $Y2=0
cc_131 N_A_190_260#_c_107_n N_A_27_368#_c_280_n 0.0055933f $X=3.552 $Y=1.095
+ $X2=0 $Y2=0
cc_132 N_A_190_260#_c_109_n N_A_27_368#_c_285_n 0.00705234f $X=1.04 $Y=1.765
+ $X2=0 $Y2=0
cc_133 N_A_190_260#_M1003_g N_A_27_368#_c_281_n 0.00203846f $X=1.075 $Y=0.74
+ $X2=0 $Y2=0
cc_134 N_A_190_260#_c_109_n N_VPWR_c_365_n 0.0111655f $X=1.04 $Y=1.765 $X2=0
+ $Y2=0
cc_135 N_A_190_260#_c_97_n N_VPWR_c_365_n 0.00131191f $X=1.49 $Y=1.765 $X2=0
+ $Y2=0
cc_136 N_A_190_260#_c_109_n N_VPWR_c_366_n 0.00413917f $X=1.04 $Y=1.765 $X2=0
+ $Y2=0
cc_137 N_A_190_260#_c_97_n N_VPWR_c_366_n 0.00461464f $X=1.49 $Y=1.765 $X2=0
+ $Y2=0
cc_138 N_A_190_260#_c_97_n N_VPWR_c_367_n 0.00903582f $X=1.49 $Y=1.765 $X2=0
+ $Y2=0
cc_139 N_A_190_260#_c_111_n N_VPWR_c_368_n 0.0153632f $X=3.4 $Y=2.375 $X2=0
+ $Y2=0
cc_140 N_A_190_260#_c_109_n N_VPWR_c_364_n 0.00414505f $X=1.04 $Y=1.765 $X2=0
+ $Y2=0
cc_141 N_A_190_260#_c_97_n N_VPWR_c_364_n 0.00469135f $X=1.49 $Y=1.765 $X2=0
+ $Y2=0
cc_142 N_A_190_260#_c_111_n N_VPWR_c_364_n 0.0175967f $X=3.4 $Y=2.375 $X2=0
+ $Y2=0
cc_143 N_A_190_260#_c_94_n N_X_c_403_n 0.005054f $X=1.04 $Y=1.675 $X2=0 $Y2=0
cc_144 N_A_190_260#_c_109_n N_X_c_403_n 0.00932545f $X=1.04 $Y=1.765 $X2=0 $Y2=0
cc_145 N_A_190_260#_M1003_g N_X_c_403_n 0.00382206f $X=1.075 $Y=0.74 $X2=0 $Y2=0
cc_146 N_A_190_260#_c_96_n N_X_c_403_n 0.00355252f $X=1.4 $Y=1.375 $X2=0 $Y2=0
cc_147 N_A_190_260#_c_97_n N_X_c_403_n 0.00502985f $X=1.49 $Y=1.765 $X2=0 $Y2=0
cc_148 N_A_190_260#_M1008_g N_X_c_403_n 0.00127735f $X=1.505 $Y=0.74 $X2=0 $Y2=0
cc_149 N_A_190_260#_c_99_n N_X_c_403_n 0.00275812f $X=1.05 $Y=1.375 $X2=0 $Y2=0
cc_150 N_A_190_260#_c_101_n N_X_c_403_n 0.0321078f $X=1.795 $Y=1.095 $X2=0 $Y2=0
cc_151 N_A_190_260#_M1003_g N_X_c_404_n 0.00881022f $X=1.075 $Y=0.74 $X2=0 $Y2=0
cc_152 N_A_190_260#_M1008_g N_X_c_404_n 0.0135262f $X=1.505 $Y=0.74 $X2=0 $Y2=0
cc_153 N_A_190_260#_M1003_g N_X_c_405_n 0.00618144f $X=1.075 $Y=0.74 $X2=0 $Y2=0
cc_154 N_A_190_260#_c_96_n N_X_c_405_n 0.00432913f $X=1.4 $Y=1.375 $X2=0 $Y2=0
cc_155 N_A_190_260#_M1008_g N_X_c_405_n 0.00405854f $X=1.505 $Y=0.74 $X2=0 $Y2=0
cc_156 N_A_190_260#_c_101_n N_X_c_405_n 0.00957189f $X=1.795 $Y=1.095 $X2=0
+ $Y2=0
cc_157 N_A_190_260#_c_96_n X 0.00226301f $X=1.4 $Y=1.375 $X2=0 $Y2=0
cc_158 N_A_190_260#_c_97_n X 0.0160122f $X=1.49 $Y=1.765 $X2=0 $Y2=0
cc_159 N_A_190_260#_c_101_n X 0.0287603f $X=1.795 $Y=1.095 $X2=0 $Y2=0
cc_160 N_A_190_260#_c_100_n N_VGND_M1008_s 0.00464866f $X=2.35 $Y=1.095 $X2=0
+ $Y2=0
cc_161 N_A_190_260#_c_101_n N_VGND_M1008_s 0.002869f $X=1.795 $Y=1.095 $X2=0
+ $Y2=0
cc_162 N_A_190_260#_c_103_n N_VGND_M1005_d 0.00358162f $X=3.35 $Y=1.095 $X2=0
+ $Y2=0
cc_163 N_A_190_260#_M1003_g N_VGND_c_446_n 0.00490645f $X=1.075 $Y=0.74 $X2=0
+ $Y2=0
cc_164 N_A_190_260#_M1003_g N_VGND_c_447_n 0.00434272f $X=1.075 $Y=0.74 $X2=0
+ $Y2=0
cc_165 N_A_190_260#_M1008_g N_VGND_c_447_n 0.00434272f $X=1.505 $Y=0.74 $X2=0
+ $Y2=0
cc_166 N_A_190_260#_c_97_n N_VGND_c_448_n 4.47758e-19 $X=1.49 $Y=1.765 $X2=0
+ $Y2=0
cc_167 N_A_190_260#_M1008_g N_VGND_c_448_n 0.00820727f $X=1.505 $Y=0.74 $X2=0
+ $Y2=0
cc_168 N_A_190_260#_c_100_n N_VGND_c_448_n 0.0196678f $X=2.35 $Y=1.095 $X2=0
+ $Y2=0
cc_169 N_A_190_260#_c_101_n N_VGND_c_448_n 0.0112912f $X=1.795 $Y=1.095 $X2=0
+ $Y2=0
cc_170 N_A_190_260#_c_102_n N_VGND_c_448_n 0.00138617f $X=2.515 $Y=0.615 $X2=0
+ $Y2=0
cc_171 N_A_190_260#_c_102_n N_VGND_c_449_n 0.0154242f $X=2.515 $Y=0.615 $X2=0
+ $Y2=0
cc_172 N_A_190_260#_c_103_n N_VGND_c_449_n 0.0248957f $X=3.35 $Y=1.095 $X2=0
+ $Y2=0
cc_173 N_A_190_260#_c_104_n N_VGND_c_449_n 0.01589f $X=3.515 $Y=0.615 $X2=0
+ $Y2=0
cc_174 N_A_190_260#_c_102_n N_VGND_c_452_n 0.0103491f $X=2.515 $Y=0.615 $X2=0
+ $Y2=0
cc_175 N_A_190_260#_c_104_n N_VGND_c_454_n 0.0127299f $X=3.515 $Y=0.615 $X2=0
+ $Y2=0
cc_176 N_A_190_260#_M1003_g N_VGND_c_455_n 0.00825283f $X=1.075 $Y=0.74 $X2=0
+ $Y2=0
cc_177 N_A_190_260#_M1008_g N_VGND_c_455_n 0.00825059f $X=1.505 $Y=0.74 $X2=0
+ $Y2=0
cc_178 N_A_190_260#_c_102_n N_VGND_c_455_n 0.0113354f $X=2.515 $Y=0.615 $X2=0
+ $Y2=0
cc_179 N_A_190_260#_c_104_n N_VGND_c_455_n 0.0139328f $X=3.515 $Y=0.615 $X2=0
+ $Y2=0
cc_180 N_A_c_208_n N_B_c_242_n 0.0810179f $X=2.215 $Y=1.765 $X2=-0.19 $Y2=-0.245
cc_181 N_A_c_210_n N_B_c_242_n 0.00285666f $X=2.14 $Y=1.515 $X2=-0.19 $Y2=-0.245
cc_182 N_A_M1006_g N_B_M1005_g 0.021941f $X=2.23 $Y=0.79 $X2=0 $Y2=0
cc_183 N_A_c_208_n N_B_c_244_n 0.00168387f $X=2.215 $Y=1.765 $X2=0 $Y2=0
cc_184 N_A_c_210_n N_B_c_244_n 0.0277335f $X=2.14 $Y=1.515 $X2=0 $Y2=0
cc_185 N_A_c_208_n N_A_27_368#_c_306_n 0.0132649f $X=2.215 $Y=1.765 $X2=0 $Y2=0
cc_186 N_A_c_210_n N_A_27_368#_c_306_n 0.0201317f $X=2.14 $Y=1.515 $X2=0 $Y2=0
cc_187 N_A_c_208_n N_A_27_368#_c_309_n 0.00350556f $X=2.215 $Y=1.765 $X2=0 $Y2=0
cc_188 N_A_c_208_n N_A_27_368#_c_322_n 6.55039e-19 $X=2.215 $Y=1.765 $X2=0 $Y2=0
cc_189 N_A_c_210_n N_VPWR_M1009_d 0.00414144f $X=2.14 $Y=1.515 $X2=0 $Y2=0
cc_190 N_A_c_208_n N_VPWR_c_367_n 0.0097414f $X=2.215 $Y=1.765 $X2=0 $Y2=0
cc_191 N_A_c_208_n N_VPWR_c_368_n 0.0049405f $X=2.215 $Y=1.765 $X2=0 $Y2=0
cc_192 N_A_c_208_n N_VPWR_c_364_n 0.00508379f $X=2.215 $Y=1.765 $X2=0 $Y2=0
cc_193 N_A_c_208_n X 0.00108439f $X=2.215 $Y=1.765 $X2=0 $Y2=0
cc_194 N_A_c_210_n X 0.026828f $X=2.14 $Y=1.515 $X2=0 $Y2=0
cc_195 N_A_M1006_g N_VGND_c_448_n 0.00658658f $X=2.23 $Y=0.79 $X2=0 $Y2=0
cc_196 N_A_M1006_g N_VGND_c_452_n 0.00507111f $X=2.23 $Y=0.79 $X2=0 $Y2=0
cc_197 N_A_M1006_g N_VGND_c_455_n 0.00514438f $X=2.23 $Y=0.79 $X2=0 $Y2=0
cc_198 N_B_c_242_n N_A_27_368#_c_277_n 0.0565457f $X=2.635 $Y=1.765 $X2=0 $Y2=0
cc_199 N_B_c_244_n N_A_27_368#_c_277_n 0.00188135f $X=2.68 $Y=1.515 $X2=0 $Y2=0
cc_200 N_B_M1005_g N_A_27_368#_M1011_g 0.0240664f $X=2.73 $Y=0.79 $X2=0 $Y2=0
cc_201 N_B_c_242_n N_A_27_368#_c_306_n 0.00803895f $X=2.635 $Y=1.765 $X2=0 $Y2=0
cc_202 N_B_c_242_n N_A_27_368#_c_309_n 0.00565434f $X=2.635 $Y=1.765 $X2=0 $Y2=0
cc_203 N_B_c_242_n N_A_27_368#_c_310_n 0.00780984f $X=2.635 $Y=1.765 $X2=0 $Y2=0
cc_204 N_B_c_244_n N_A_27_368#_c_310_n 0.0133767f $X=2.68 $Y=1.515 $X2=0 $Y2=0
cc_205 N_B_c_242_n N_A_27_368#_c_322_n 0.00350007f $X=2.635 $Y=1.765 $X2=0 $Y2=0
cc_206 N_B_c_244_n N_A_27_368#_c_322_n 0.00875303f $X=2.68 $Y=1.515 $X2=0 $Y2=0
cc_207 N_B_c_242_n N_A_27_368#_c_280_n 0.00283175f $X=2.635 $Y=1.765 $X2=0 $Y2=0
cc_208 N_B_c_244_n N_A_27_368#_c_280_n 0.0249838f $X=2.68 $Y=1.515 $X2=0 $Y2=0
cc_209 N_B_c_242_n N_VPWR_c_368_n 0.0049405f $X=2.635 $Y=1.765 $X2=0 $Y2=0
cc_210 N_B_c_242_n N_VPWR_c_364_n 0.00508379f $X=2.635 $Y=1.765 $X2=0 $Y2=0
cc_211 N_B_M1005_g N_VGND_c_449_n 0.00564618f $X=2.73 $Y=0.79 $X2=0 $Y2=0
cc_212 N_B_M1005_g N_VGND_c_452_n 0.00485498f $X=2.73 $Y=0.79 $X2=0 $Y2=0
cc_213 N_B_M1005_g N_VGND_c_455_n 0.00514438f $X=2.73 $Y=0.79 $X2=0 $Y2=0
cc_214 N_A_27_368#_c_279_n N_VPWR_M1007_d 0.00124681f $X=0.69 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_215 N_A_27_368#_c_306_n N_VPWR_M1007_d 0.00650439f $X=2.475 $Y=2.405
+ $X2=-0.19 $Y2=-0.245
cc_216 N_A_27_368#_c_285_n N_VPWR_M1007_d 0.00664477f $X=0.28 $Y=2.115 $X2=-0.19
+ $Y2=-0.245
cc_217 N_A_27_368#_c_306_n N_VPWR_M1009_d 0.0168222f $X=2.475 $Y=2.405 $X2=0
+ $Y2=0
cc_218 N_A_27_368#_c_306_n N_VPWR_c_365_n 0.0115499f $X=2.475 $Y=2.405 $X2=0
+ $Y2=0
cc_219 N_A_27_368#_c_285_n N_VPWR_c_365_n 0.0135988f $X=0.28 $Y=2.115 $X2=0
+ $Y2=0
cc_220 N_A_27_368#_c_306_n N_VPWR_c_367_n 0.0344564f $X=2.475 $Y=2.405 $X2=0
+ $Y2=0
cc_221 N_A_27_368#_c_277_n N_VPWR_c_368_n 0.00481995f $X=3.175 $Y=1.765 $X2=0
+ $Y2=0
cc_222 N_A_27_368#_c_277_n N_VPWR_c_364_n 0.00508379f $X=3.175 $Y=1.765 $X2=0
+ $Y2=0
cc_223 N_A_27_368#_c_306_n N_VPWR_c_364_n 0.0424245f $X=2.475 $Y=2.405 $X2=0
+ $Y2=0
cc_224 N_A_27_368#_c_285_n N_VPWR_c_364_n 0.0179459f $X=0.28 $Y=2.115 $X2=0
+ $Y2=0
cc_225 N_A_27_368#_c_285_n N_VPWR_c_370_n 0.00671799f $X=0.28 $Y=2.115 $X2=0
+ $Y2=0
cc_226 N_A_27_368#_c_306_n N_X_M1000_s 0.00571991f $X=2.475 $Y=2.405 $X2=0 $Y2=0
cc_227 N_A_27_368#_c_279_n N_X_c_403_n 0.0403465f $X=0.69 $Y=1.95 $X2=0 $Y2=0
cc_228 N_A_27_368#_c_306_n N_X_c_403_n 0.0088501f $X=2.475 $Y=2.405 $X2=0 $Y2=0
cc_229 N_A_27_368#_c_285_n N_X_c_403_n 0.0115377f $X=0.28 $Y=2.115 $X2=0 $Y2=0
cc_230 N_A_27_368#_c_281_n N_X_c_404_n 0.00520473f $X=0.35 $Y=0.835 $X2=0 $Y2=0
cc_231 N_A_27_368#_c_281_n N_X_c_405_n 0.00935177f $X=0.35 $Y=0.835 $X2=0 $Y2=0
cc_232 N_A_27_368#_c_306_n X 0.0332551f $X=2.475 $Y=2.405 $X2=0 $Y2=0
cc_233 N_A_27_368#_c_306_n A_458_368# 0.00804595f $X=2.475 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_234 N_A_27_368#_c_309_n A_458_368# 0.00222425f $X=2.56 $Y=2.32 $X2=-0.19
+ $Y2=-0.245
cc_235 N_A_27_368#_c_322_n A_458_368# 0.00271734f $X=2.645 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_236 N_A_27_368#_c_310_n A_542_368# 0.0190705f $X=3.085 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_237 N_A_27_368#_c_281_n N_VGND_M1004_d 0.00517204f $X=0.35 $Y=0.835 $X2=-0.19
+ $Y2=-0.245
cc_238 N_A_27_368#_c_281_n N_VGND_c_446_n 0.0189052f $X=0.35 $Y=0.835 $X2=0
+ $Y2=0
cc_239 N_A_27_368#_M1011_g N_VGND_c_449_n 0.00564618f $X=3.3 $Y=0.79 $X2=0 $Y2=0
cc_240 N_A_27_368#_c_281_n N_VGND_c_450_n 0.0101249f $X=0.35 $Y=0.835 $X2=0
+ $Y2=0
cc_241 N_A_27_368#_M1011_g N_VGND_c_454_n 0.00485498f $X=3.3 $Y=0.79 $X2=0 $Y2=0
cc_242 N_A_27_368#_M1011_g N_VGND_c_455_n 0.00514438f $X=3.3 $Y=0.79 $X2=0 $Y2=0
cc_243 N_A_27_368#_c_281_n N_VGND_c_455_n 0.0134471f $X=0.35 $Y=0.835 $X2=0
+ $Y2=0
cc_244 N_VPWR_M1009_d X 0.0056818f $X=1.565 $Y=1.84 $X2=0 $Y2=0
cc_245 N_X_c_404_n N_VGND_c_446_n 0.0164567f $X=1.29 $Y=0.515 $X2=0 $Y2=0
cc_246 N_X_c_404_n N_VGND_c_447_n 0.0144922f $X=1.29 $Y=0.515 $X2=0 $Y2=0
cc_247 N_X_c_404_n N_VGND_c_448_n 0.0169789f $X=1.29 $Y=0.515 $X2=0 $Y2=0
cc_248 N_X_c_404_n N_VGND_c_455_n 0.0118826f $X=1.29 $Y=0.515 $X2=0 $Y2=0
