* NGSPICE file created from sky130_fd_sc_ls__nor3b_1.ext - technology: sky130A

.subckt sky130_fd_sc_ls__nor3b_1 A B C_N VGND VNB VPB VPWR Y
M1000 Y a_27_112# a_344_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=4.704e+11p ps=3.08e+06u
M1001 a_344_368# B a_260_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.024e+11p ps=2.78e+06u
M1002 a_260_368# A VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=4.354e+11p ps=3.08e+06u
M1003 VPWR C_N a_27_112# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=2.478e+11p ps=2.27e+06u
M1004 VGND C_N a_27_112# VNB nshort w=550000u l=150000u
+  ad=5.8515e+11p pd=4.58e+06u as=2.695e+11p ps=2.08e+06u
M1005 VGND B Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=4.477e+11p ps=4.17e+06u
M1006 Y A VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y a_27_112# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

