* File: sky130_fd_sc_ls__decaphe_6.spice
* Created: Fri Aug 28 13:12:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__decaphe_6.pex.spice"
.subckt sky130_fd_sc_ls__decaphe_6  VNB VPB VGND VPWR
* 
* VPWR	VPWR
* VGND	VGND
* VPB	VPB
* VNB	VNB
MM1000 N_VGND_M1000_s N_VPWR_M1000_g N_VGND_M1000_s VNB NSHORT L=2.09 W=0.775
+ AD=0.2015 AS=0.2015 PD=2.07 PS=2.07 NRD=0 NRS=0 M=1 R=0.370813 SA=1.045e+06
+ SB=1.045e+06 A=1.61975 P=5.73 MULT=1
MM1001 N_VPWR_M1001_s N_VGND_M1001_g N_VPWR_M1001_s VPB PSHORT L=2.09 W=1.255
+ AD=0.3263 AS=0.3263 PD=3.03 PS=3.03 NRD=0 NRS=0 M=1 R=0.600478 SA=1.045e+06
+ SB=1.045e+06 A=2.62295 P=6.69 MULT=1
DX2_noxref VNB VPB NWDIODE A=6.0636 P=10.24
*
.include "sky130_fd_sc_ls__decaphe_6.pxi.spice"
*
.ends
*
*
