# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ls__sdfrbp_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ls__sdfrbp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  14.88000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 0.810000 2.090000 1.190000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 14.055000 0.350000 14.325000 2.980000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.030000 0.915000 12.465000 1.085000 ;
        RECT 12.030000 1.085000 12.360000 2.980000 ;
        RECT 12.135000 0.350000 12.465000 0.915000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.411000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  3.785000 1.820000  4.165000 2.150000 ;
        RECT  7.720000 1.795000  8.020000 2.150000 ;
        RECT 10.715000 1.820000 11.395000 2.150000 ;
      LAYER mcon ;
        RECT  3.995000 1.950000  4.165000 2.120000 ;
        RECT  7.835000 1.950000  8.005000 2.120000 ;
        RECT 10.715000 1.950000 10.885000 2.120000 ;
      LAYER met1 ;
        RECT  3.935000 1.920000  4.225000 1.965000 ;
        RECT  3.935000 1.965000 10.945000 2.105000 ;
        RECT  3.935000 2.105000  4.225000 2.150000 ;
        RECT  7.775000 1.920000  8.065000 1.965000 ;
        RECT  7.775000 2.105000  8.065000 2.150000 ;
        RECT 10.655000 1.920000 10.945000 1.965000 ;
        RECT 10.655000 2.105000 10.945000 2.150000 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.945000 1.440000 3.275000 2.150000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.540000 1.820000 1.795000 2.150000 ;
        RECT 1.625000 1.360000 2.735000 1.620000 ;
        RECT 1.625000 1.620000 1.795000 1.820000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.905000 1.180000 4.235000 1.550000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 14.880000 0.085000 ;
        RECT  0.545000  0.085000  0.875000 0.835000 ;
        RECT  3.640000  0.085000  3.970000 0.835000 ;
        RECT  4.750000  0.085000  4.920000 1.130000 ;
        RECT  7.450000  0.085000  7.985000 0.410000 ;
        RECT 10.335000  0.085000 10.665000 0.810000 ;
        RECT 11.645000  0.085000 11.895000 0.535000 ;
        RECT 12.635000  0.085000 12.895000 1.050000 ;
        RECT 13.670000  0.085000 13.840000 1.130000 ;
        RECT 14.495000  0.085000 14.780000 1.130000 ;
      LAYER mcon ;
        RECT  0.155000 -0.085000  0.325000 0.085000 ;
        RECT  0.635000 -0.085000  0.805000 0.085000 ;
        RECT  1.115000 -0.085000  1.285000 0.085000 ;
        RECT  1.595000 -0.085000  1.765000 0.085000 ;
        RECT  2.075000 -0.085000  2.245000 0.085000 ;
        RECT  2.555000 -0.085000  2.725000 0.085000 ;
        RECT  3.035000 -0.085000  3.205000 0.085000 ;
        RECT  3.515000 -0.085000  3.685000 0.085000 ;
        RECT  3.995000 -0.085000  4.165000 0.085000 ;
        RECT  4.475000 -0.085000  4.645000 0.085000 ;
        RECT  4.955000 -0.085000  5.125000 0.085000 ;
        RECT  5.435000 -0.085000  5.605000 0.085000 ;
        RECT  5.915000 -0.085000  6.085000 0.085000 ;
        RECT  6.395000 -0.085000  6.565000 0.085000 ;
        RECT  6.875000 -0.085000  7.045000 0.085000 ;
        RECT  7.355000 -0.085000  7.525000 0.085000 ;
        RECT  7.835000 -0.085000  8.005000 0.085000 ;
        RECT  8.315000 -0.085000  8.485000 0.085000 ;
        RECT  8.795000 -0.085000  8.965000 0.085000 ;
        RECT  9.275000 -0.085000  9.445000 0.085000 ;
        RECT  9.755000 -0.085000  9.925000 0.085000 ;
        RECT 10.235000 -0.085000 10.405000 0.085000 ;
        RECT 10.715000 -0.085000 10.885000 0.085000 ;
        RECT 11.195000 -0.085000 11.365000 0.085000 ;
        RECT 11.675000 -0.085000 11.845000 0.085000 ;
        RECT 12.155000 -0.085000 12.325000 0.085000 ;
        RECT 12.635000 -0.085000 12.805000 0.085000 ;
        RECT 13.115000 -0.085000 13.285000 0.085000 ;
        RECT 13.595000 -0.085000 13.765000 0.085000 ;
        RECT 14.075000 -0.085000 14.245000 0.085000 ;
        RECT 14.555000 -0.085000 14.725000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 14.880000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 3.245000 14.880000 3.415000 ;
        RECT  0.615000 2.730000  1.400000 3.245000 ;
        RECT  3.115000 2.660000  3.445000 3.245000 ;
        RECT  4.705000 2.750000  5.035000 3.245000 ;
        RECT  7.070000 2.680000  7.320000 3.245000 ;
        RECT  8.190000 1.745000  8.440000 3.245000 ;
        RECT 10.265000 2.660000 10.860000 3.245000 ;
        RECT 11.600000 1.820000 11.850000 3.245000 ;
        RECT 12.540000 1.920000 12.830000 3.245000 ;
        RECT 13.545000 1.820000 13.875000 3.245000 ;
        RECT 14.495000 1.820000 14.775000 3.245000 ;
      LAYER mcon ;
        RECT  0.155000 3.245000  0.325000 3.415000 ;
        RECT  0.635000 3.245000  0.805000 3.415000 ;
        RECT  1.115000 3.245000  1.285000 3.415000 ;
        RECT  1.595000 3.245000  1.765000 3.415000 ;
        RECT  2.075000 3.245000  2.245000 3.415000 ;
        RECT  2.555000 3.245000  2.725000 3.415000 ;
        RECT  3.035000 3.245000  3.205000 3.415000 ;
        RECT  3.515000 3.245000  3.685000 3.415000 ;
        RECT  3.995000 3.245000  4.165000 3.415000 ;
        RECT  4.475000 3.245000  4.645000 3.415000 ;
        RECT  4.955000 3.245000  5.125000 3.415000 ;
        RECT  5.435000 3.245000  5.605000 3.415000 ;
        RECT  5.915000 3.245000  6.085000 3.415000 ;
        RECT  6.395000 3.245000  6.565000 3.415000 ;
        RECT  6.875000 3.245000  7.045000 3.415000 ;
        RECT  7.355000 3.245000  7.525000 3.415000 ;
        RECT  7.835000 3.245000  8.005000 3.415000 ;
        RECT  8.315000 3.245000  8.485000 3.415000 ;
        RECT  8.795000 3.245000  8.965000 3.415000 ;
        RECT  9.275000 3.245000  9.445000 3.415000 ;
        RECT  9.755000 3.245000  9.925000 3.415000 ;
        RECT 10.235000 3.245000 10.405000 3.415000 ;
        RECT 10.715000 3.245000 10.885000 3.415000 ;
        RECT 11.195000 3.245000 11.365000 3.415000 ;
        RECT 11.675000 3.245000 11.845000 3.415000 ;
        RECT 12.155000 3.245000 12.325000 3.415000 ;
        RECT 12.635000 3.245000 12.805000 3.415000 ;
        RECT 13.115000 3.245000 13.285000 3.415000 ;
        RECT 13.595000 3.245000 13.765000 3.415000 ;
        RECT 14.075000 3.245000 14.245000 3.415000 ;
        RECT 14.555000 3.245000 14.725000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 14.880000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.115000 0.375000  0.365000 1.250000 ;
      RECT  0.115000 1.250000  1.395000 1.580000 ;
      RECT  0.115000 1.580000  0.285000 2.320000 ;
      RECT  0.115000 2.320000  2.605000 2.490000 ;
      RECT  0.115000 2.490000  0.445000 2.980000 ;
      RECT  1.095000 0.255000  3.430000 0.425000 ;
      RECT  1.095000 0.425000  1.345000 0.835000 ;
      RECT  1.940000 2.660000  2.945000 2.910000 ;
      RECT  2.260000 0.595000  2.610000 1.005000 ;
      RECT  2.260000 1.005000  3.615000 1.175000 ;
      RECT  2.275000 1.830000  2.605000 2.320000 ;
      RECT  2.775000 2.320000  3.995000 2.420000 ;
      RECT  2.775000 2.420000  5.985000 2.490000 ;
      RECT  2.775000 2.490000  2.945000 2.660000 ;
      RECT  3.100000 0.425000  3.430000 0.835000 ;
      RECT  3.445000 1.175000  3.615000 2.320000 ;
      RECT  3.615000 2.490000  5.985000 2.580000 ;
      RECT  3.615000 2.580000  4.645000 2.590000 ;
      RECT  3.615000 2.590000  3.995000 2.980000 ;
      RECT  4.240000 0.595000  4.575000 1.010000 ;
      RECT  4.335000 1.820000  4.985000 1.990000 ;
      RECT  4.335000 1.990000  4.505000 2.250000 ;
      RECT  4.405000 1.010000  4.575000 1.445000 ;
      RECT  4.405000 1.445000  5.305000 1.775000 ;
      RECT  4.405000 1.775000  4.985000 1.820000 ;
      RECT  4.570000 2.410000  5.985000 2.420000 ;
      RECT  5.100000 0.310000  7.170000 0.480000 ;
      RECT  5.100000 0.480000  5.430000 0.990000 ;
      RECT  5.100000 0.990000  5.645000 1.275000 ;
      RECT  5.155000 1.945000  6.150000 1.985000 ;
      RECT  5.155000 1.985000  5.675000 2.030000 ;
      RECT  5.155000 2.030000  5.630000 2.240000 ;
      RECT  5.430000 1.900000  6.150000 1.945000 ;
      RECT  5.475000 1.275000  5.645000 1.500000 ;
      RECT  5.475000 1.500000  6.150000 1.900000 ;
      RECT  5.660000 0.650000  5.990000 0.820000 ;
      RECT  5.710000 2.580000  5.985000 2.725000 ;
      RECT  5.800000 2.155000  6.490000 2.325000 ;
      RECT  5.800000 2.325000  5.985000 2.410000 ;
      RECT  5.820000 0.820000  5.990000 1.120000 ;
      RECT  5.820000 1.120000  6.490000 1.290000 ;
      RECT  6.160000 0.650000  6.830000 0.950000 ;
      RECT  6.160000 2.495000  7.915000 2.510000 ;
      RECT  6.160000 2.510000  6.900000 2.725000 ;
      RECT  6.320000 1.290000  6.490000 2.155000 ;
      RECT  6.660000 0.950000  6.830000 2.340000 ;
      RECT  6.660000 2.340000  7.915000 2.495000 ;
      RECT  7.000000 0.480000  7.170000 0.580000 ;
      RECT  7.000000 0.580000  8.325000 0.750000 ;
      RECT  7.000000 0.920000  8.930000 1.090000 ;
      RECT  7.000000 1.090000  7.210000 1.780000 ;
      RECT  7.380000 1.260000  8.590000 1.575000 ;
      RECT  7.380000 1.575000  7.550000 2.320000 ;
      RECT  7.380000 2.320000  7.915000 2.340000 ;
      RECT  7.550000 2.510000  7.915000 2.725000 ;
      RECT  8.155000 0.255000  9.270000 0.425000 ;
      RECT  8.155000 0.425000  8.325000 0.580000 ;
      RECT  8.495000 0.595000  8.930000 0.920000 ;
      RECT  8.640000 1.745000  8.930000 2.755000 ;
      RECT  8.760000 1.090000  8.930000 1.745000 ;
      RECT  9.100000 0.425000  9.270000 0.905000 ;
      RECT  9.100000 0.905000  9.640000 1.235000 ;
      RECT  9.100000 2.365000 10.095000 2.695000 ;
      RECT  9.310000 1.235000  9.640000 1.865000 ;
      RECT  9.310000 1.865000  9.755000 2.195000 ;
      RECT  9.440000 0.405000 10.095000 0.735000 ;
      RECT  9.925000 0.735000 10.095000 1.045000 ;
      RECT  9.925000 1.045000 11.520000 1.310000 ;
      RECT  9.925000 1.310000 10.095000 2.365000 ;
      RECT 10.265000 1.480000 11.860000 1.650000 ;
      RECT 10.265000 1.650000 10.545000 2.320000 ;
      RECT 10.265000 2.320000 11.395000 2.490000 ;
      RECT 11.065000 2.490000 11.395000 2.795000 ;
      RECT 11.125000 0.350000 11.455000 0.705000 ;
      RECT 11.125000 0.705000 11.860000 0.875000 ;
      RECT 11.690000 0.875000 11.860000 1.480000 ;
      RECT 13.065000 0.350000 13.325000 1.300000 ;
      RECT 13.065000 1.300000 13.885000 1.630000 ;
      RECT 13.065000 1.630000 13.325000 2.980000 ;
  END
END sky130_fd_sc_ls__sdfrbp_2
