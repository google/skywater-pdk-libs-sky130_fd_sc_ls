* File: sky130_fd_sc_ls__decaphe_8.spice
* Created: Fri Aug 28 13:12:50 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__decaphe_8.pex.spice"
.subckt sky130_fd_sc_ls__decaphe_8  VNB VPB VGND VPWR
* 
* VPWR	VPWR
* VGND	VGND
* VPB	VPB
* VNB	VNB
MM1000 N_VGND_M1000_s N_VPWR_M1000_g N_VGND_M1000_s VNB NSHORT L=3.05 W=0.775
+ AD=0.2015 AS=0.2015 PD=2.07 PS=2.07 NRD=0 NRS=0 M=1 R=0.254098 SA=1.525e+06
+ SB=1.525e+06 A=2.36375 P=7.65 MULT=1
MM1001 N_VPWR_M1001_s N_VGND_M1001_g N_VPWR_M1001_s VPB PSHORT L=3.05 W=1.255
+ AD=0.3263 AS=0.3263 PD=3.03 PS=3.03 NRD=0 NRS=0 M=1 R=0.411475 SA=1.525e+06
+ SB=1.525e+06 A=3.82775 P=8.61 MULT=1
DX2_noxref VNB VPB NWDIODE A=7.8492 P=12.16
*
.include "sky130_fd_sc_ls__decaphe_8.pxi.spice"
*
.ends
*
*
