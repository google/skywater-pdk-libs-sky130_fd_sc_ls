* File: sky130_fd_sc_ls__nor4_1.pex.spice
* Created: Fri Aug 28 13:39:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__NOR4_1%A 1 3 6 8 9 10 14
r25 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.375
+ $Y=1.385 $X2=0.375 $Y2=1.385
r26 10 14 4.20486 $w=3.68e-07 $l=1.35e-07 $layer=LI1_cond $X=0.24 $Y=1.365
+ $X2=0.375 $Y2=1.365
r27 8 13 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=0.555 $Y=1.385
+ $X2=0.375 $Y2=1.385
r28 8 9 66.2869 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.645 $Y=1.385
+ $X2=0.645 $Y2=1.22
r29 6 9 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.66 $Y=0.74 $X2=0.66
+ $Y2=1.22
r30 1 8 149.859 $w=1.8e-07 $l=3.8e-07 $layer=POLY_cond $X=0.645 $Y=1.765
+ $X2=0.645 $Y2=1.385
r31 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.645 $Y=1.765
+ $X2=0.645 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__NOR4_1%B 1 3 6 8 9 10 11 18
r37 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.14
+ $Y=1.515 $X2=1.14 $Y2=1.515
r38 10 11 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=1.145 $Y=2.405
+ $X2=1.145 $Y2=2.775
r39 9 10 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=1.145 $Y=2.035
+ $X2=1.145 $Y2=2.405
r40 8 9 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=1.145 $Y=1.665
+ $X2=1.145 $Y2=2.035
r41 8 18 5.08431 $w=3.38e-07 $l=1.5e-07 $layer=LI1_cond $X=1.145 $Y=1.665
+ $X2=1.145 $Y2=1.515
r42 4 17 38.5562 $w=2.99e-07 $l=1.88348e-07 $layer=POLY_cond $X=1.09 $Y=1.35
+ $X2=1.14 $Y2=1.515
r43 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.09 $Y=1.35 $X2=1.09
+ $Y2=0.74
r44 1 17 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=1.065 $Y=1.765
+ $X2=1.14 $Y2=1.515
r45 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.065 $Y=1.765
+ $X2=1.065 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__NOR4_1%C 1 3 6 8 9 14
r31 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.71
+ $Y=1.515 $X2=1.71 $Y2=1.515
r32 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.71 $Y=1.665 $X2=1.71
+ $Y2=2.035
r33 8 14 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.71 $Y=1.665
+ $X2=1.71 $Y2=1.515
r34 4 13 38.5562 $w=2.99e-07 $l=1.88348e-07 $layer=POLY_cond $X=1.76 $Y=1.35
+ $X2=1.71 $Y2=1.515
r35 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.76 $Y=1.35 $X2=1.76
+ $Y2=0.74
r36 1 13 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=1.635 $Y=1.765
+ $X2=1.71 $Y2=1.515
r37 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.635 $Y=1.765
+ $X2=1.635 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__NOR4_1%D 3 5 7 8 12
r27 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.28
+ $Y=1.515 $X2=2.28 $Y2=1.515
r28 8 12 4.32166 $w=3.98e-07 $l=1.5e-07 $layer=LI1_cond $X=2.245 $Y=1.665
+ $X2=2.245 $Y2=1.515
r29 5 11 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=2.205 $Y=1.765
+ $X2=2.28 $Y2=1.515
r30 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.205 $Y=1.765
+ $X2=2.205 $Y2=2.4
r31 1 11 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=2.19 $Y=1.35
+ $X2=2.28 $Y2=1.515
r32 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.19 $Y=1.35 $X2=2.19
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__NOR4_1%VPWR 1 4 6 10 17 18
r22 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r23 17 18 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r24 15 22 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r25 14 17 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.72 $Y=3.33
+ $X2=2.64 $Y2=3.33
r26 14 15 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r27 12 21 4.49701 $w=1.7e-07 $l=2.93e-07 $layer=LI1_cond $X=0.585 $Y=3.33
+ $X2=0.292 $Y2=3.33
r28 12 14 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=0.585 $Y=3.33
+ $X2=0.72 $Y2=3.33
r29 10 18 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=2.64 $Y2=3.33
r30 10 15 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=0.72 $Y2=3.33
r31 6 9 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=0.42 $Y=1.985 $X2=0.42
+ $Y2=2.815
r32 4 21 3.26916 $w=3.3e-07 $l=1.65118e-07 $layer=LI1_cond $X=0.42 $Y=3.245
+ $X2=0.292 $Y2=3.33
r33 4 9 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.42 $Y=3.245 $X2=0.42
+ $Y2=2.815
r34 1 9 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.275
+ $Y=1.84 $X2=0.42 $Y2=2.815
r35 1 6 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.275
+ $Y=1.84 $X2=0.42 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_LS__NOR4_1%Y 1 2 3 12 14 15 18 20 24 27 28 29
r56 29 34 0.92006 $w=5.18e-07 $l=4e-08 $layer=LI1_cond $X=2.525 $Y=2.775
+ $X2=2.525 $Y2=2.815
r57 27 28 9.6413 $w=5.18e-07 $l=1.65e-07 $layer=LI1_cond $X=2.525 $Y=2.115
+ $X2=2.525 $Y2=1.95
r58 25 29 12.9959 $w=5.18e-07 $l=5.65e-07 $layer=LI1_cond $X=2.525 $Y=2.21
+ $X2=2.525 $Y2=2.775
r59 25 27 2.18514 $w=5.18e-07 $l=9.5e-08 $layer=LI1_cond $X=2.525 $Y=2.21
+ $X2=2.525 $Y2=2.115
r60 22 28 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=2.7 $Y=1.18 $X2=2.7
+ $Y2=1.95
r61 21 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.14 $Y=1.095
+ $X2=1.975 $Y2=1.095
r62 20 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.615 $Y=1.095
+ $X2=2.7 $Y2=1.18
r63 20 21 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=2.615 $Y=1.095
+ $X2=2.14 $Y2=1.095
r64 16 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.975 $Y=1.01
+ $X2=1.975 $Y2=1.095
r65 16 18 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=1.975 $Y=1.01
+ $X2=1.975 $Y2=0.515
r66 14 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.81 $Y=1.095
+ $X2=1.975 $Y2=1.095
r67 14 15 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.81 $Y=1.095
+ $X2=1.04 $Y2=1.095
r68 10 15 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.91 $Y=1.01
+ $X2=1.04 $Y2=1.095
r69 10 12 21.9407 $w=2.58e-07 $l=4.95e-07 $layer=LI1_cond $X=0.91 $Y=1.01
+ $X2=0.91 $Y2=0.515
r70 3 34 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.28
+ $Y=1.84 $X2=2.43 $Y2=2.815
r71 3 27 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=2.28
+ $Y=1.84 $X2=2.43 $Y2=2.115
r72 2 18 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.835
+ $Y=0.37 $X2=1.975 $Y2=0.515
r73 1 12 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.735
+ $Y=0.37 $X2=0.875 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__NOR4_1%VGND 1 2 3 10 12 16 18 20 23 24 25 31 40
r36 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r37 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r38 34 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r39 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r40 31 39 4.51706 $w=1.7e-07 $l=2.85e-07 $layer=LI1_cond $X=2.31 $Y=0 $X2=2.595
+ $Y2=0
r41 31 33 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=2.31 $Y=0 $X2=2.16
+ $Y2=0
r42 30 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.24
+ $Y2=0
r43 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r44 27 36 5.15784 $w=1.7e-07 $l=3.05e-07 $layer=LI1_cond $X=0.61 $Y=0 $X2=0.305
+ $Y2=0
r45 27 29 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=0.61 $Y=0 $X2=1.2
+ $Y2=0
r46 25 34 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=2.16
+ $Y2=0
r47 25 30 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.2
+ $Y2=0
r48 23 29 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=1.21 $Y=0 $X2=1.2
+ $Y2=0
r49 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.21 $Y=0 $X2=1.375
+ $Y2=0
r50 22 33 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=1.54 $Y=0 $X2=2.16
+ $Y2=0
r51 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.54 $Y=0 $X2=1.375
+ $Y2=0
r52 18 39 3.24911 $w=3.3e-07 $l=1.56844e-07 $layer=LI1_cond $X=2.475 $Y=0.085
+ $X2=2.595 $Y2=0
r53 18 20 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=2.475 $Y=0.085
+ $X2=2.475 $Y2=0.675
r54 14 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.375 $Y=0.085
+ $X2=1.375 $Y2=0
r55 14 16 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=1.375 $Y=0.085
+ $X2=1.375 $Y2=0.675
r56 10 36 3.21308 $w=4e-07 $l=1.41244e-07 $layer=LI1_cond $X=0.41 $Y=0.085
+ $X2=0.305 $Y2=0
r57 10 12 12.3888 $w=3.98e-07 $l=4.3e-07 $layer=LI1_cond $X=0.41 $Y=0.085
+ $X2=0.41 $Y2=0.515
r58 3 20 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=2.265
+ $Y=0.37 $X2=2.405 $Y2=0.675
r59 2 16 182 $w=1.7e-07 $l=3.96327e-07 $layer=licon1_NDIFF $count=1 $X=1.165
+ $Y=0.37 $X2=1.375 $Y2=0.675
r60 1 12 91 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_NDIFF $count=2 $X=0.23
+ $Y=0.37 $X2=0.445 $Y2=0.515
.ends

