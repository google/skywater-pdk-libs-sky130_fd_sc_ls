* NGSPICE file created from sky130_fd_sc_ls__a222oi_1.ext - technology: sky130A

.subckt sky130_fd_sc_ls__a222oi_1 A1 A2 B1 B2 C1 C2 VGND VNB VPB VPWR Y
M1000 a_461_74# B2 VGND VNB nshort w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=9.312e+11p ps=5.47e+06u
M1001 a_116_392# B2 a_369_392# VPB phighvt w=1e+06u l=150000u
+  ad=7e+11p pd=5.4e+06u as=9.4e+11p ps=7.88e+06u
M1002 a_119_74# C1 Y VNB nshort w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=5.92e+11p ps=4.41e+06u
M1003 Y B1 a_461_74# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_369_392# B1 a_116_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_697_74# A1 Y VNB nshort w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1006 VGND A2 a_697_74# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR A1 a_369_392# VPB phighvt w=1e+06u l=150000u
+  ad=4.5e+11p pd=2.9e+06u as=0p ps=0u
M1008 Y C2 a_116_392# VPB phighvt w=1e+06u l=150000u
+  ad=6.4e+11p pd=5.28e+06u as=0p ps=0u
M1009 a_116_392# C1 Y VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_369_392# A2 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND C2 a_119_74# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

