* File: sky130_fd_sc_ls__a31o_1.pxi.spice
* Created: Fri Aug 28 12:58:36 2020
* 
x_PM_SKY130_FD_SC_LS__A31O_1%A_81_270# N_A_81_270#_M1009_d N_A_81_270#_M1004_d
+ N_A_81_270#_c_57_n N_A_81_270#_M1006_g N_A_81_270#_c_58_n N_A_81_270#_M1005_g
+ N_A_81_270#_c_59_n N_A_81_270#_c_91_p N_A_81_270#_c_60_n N_A_81_270#_c_61_n
+ N_A_81_270#_c_62_n N_A_81_270#_c_63_n PM_SKY130_FD_SC_LS__A31O_1%A_81_270#
x_PM_SKY130_FD_SC_LS__A31O_1%A3 N_A3_c_130_n N_A3_M1002_g N_A3_M1008_g A3
+ PM_SKY130_FD_SC_LS__A31O_1%A3
x_PM_SKY130_FD_SC_LS__A31O_1%A2 N_A2_M1003_g N_A2_c_163_n N_A2_M1007_g A2
+ PM_SKY130_FD_SC_LS__A31O_1%A2
x_PM_SKY130_FD_SC_LS__A31O_1%A1 N_A1_M1009_g N_A1_c_193_n N_A1_M1001_g A1
+ PM_SKY130_FD_SC_LS__A31O_1%A1
x_PM_SKY130_FD_SC_LS__A31O_1%B1 N_B1_c_225_n N_B1_c_231_n N_B1_M1004_g
+ N_B1_M1000_g N_B1_c_227_n B1 B1 B1 N_B1_c_228_n N_B1_c_229_n
+ PM_SKY130_FD_SC_LS__A31O_1%B1
x_PM_SKY130_FD_SC_LS__A31O_1%X N_X_M1005_s N_X_M1006_s N_X_c_266_n N_X_c_267_n X
+ X X X N_X_c_268_n PM_SKY130_FD_SC_LS__A31O_1%X
x_PM_SKY130_FD_SC_LS__A31O_1%VPWR N_VPWR_M1006_d N_VPWR_M1007_d N_VPWR_c_289_n
+ N_VPWR_c_290_n N_VPWR_c_291_n N_VPWR_c_292_n VPWR N_VPWR_c_293_n
+ N_VPWR_c_294_n N_VPWR_c_288_n N_VPWR_c_296_n PM_SKY130_FD_SC_LS__A31O_1%VPWR
x_PM_SKY130_FD_SC_LS__A31O_1%A_250_392# N_A_250_392#_M1002_d
+ N_A_250_392#_M1001_d N_A_250_392#_c_330_n N_A_250_392#_c_328_n
+ N_A_250_392#_c_331_n N_A_250_392#_c_332_n N_A_250_392#_c_329_n
+ PM_SKY130_FD_SC_LS__A31O_1%A_250_392#
x_PM_SKY130_FD_SC_LS__A31O_1%VGND N_VGND_M1005_d N_VGND_M1000_d N_VGND_c_362_n
+ N_VGND_c_363_n N_VGND_c_364_n N_VGND_c_365_n VGND N_VGND_c_366_n
+ N_VGND_c_367_n N_VGND_c_368_n N_VGND_c_369_n PM_SKY130_FD_SC_LS__A31O_1%VGND
cc_1 VNB N_A_81_270#_c_57_n 0.0289684f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.765
cc_2 VNB N_A_81_270#_c_58_n 0.0221308f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.35
cc_3 VNB N_A_81_270#_c_59_n 0.0121926f $X=-0.19 $Y=-0.245 $X2=2.28 $Y2=1.235
cc_4 VNB N_A_81_270#_c_60_n 0.0088318f $X=-0.19 $Y=-0.245 $X2=2.845 $Y2=1.235
cc_5 VNB N_A_81_270#_c_61_n 0.0173236f $X=-0.19 $Y=-0.245 $X2=2.93 $Y2=2.105
cc_6 VNB N_A_81_270#_c_62_n 0.00531266f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.235
cc_7 VNB N_A_81_270#_c_63_n 0.00437417f $X=-0.19 $Y=-0.245 $X2=2.445 $Y2=1.235
cc_8 VNB N_A3_c_130_n 0.0155191f $X=-0.19 $Y=-0.245 $X2=2.225 $Y2=0.615
cc_9 VNB N_A3_M1008_g 0.0237957f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB A3 0.0021755f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_11 VNB N_A2_M1003_g 0.0226062f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A2_c_163_n 0.0173059f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A1_M1009_g 0.0235943f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A1_c_193_n 0.0153134f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB A1 0.00279888f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_16 VNB N_B1_c_225_n 0.0042235f $X=-0.19 $Y=-0.245 $X2=2.78 $Y2=1.96
cc_17 VNB N_B1_M1000_g 0.0179075f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_18 VNB N_B1_c_227_n 0.011517f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.87
cc_19 VNB N_B1_c_228_n 0.0473693f $X=-0.19 $Y=-0.245 $X2=2.845 $Y2=1.235
cc_20 VNB N_B1_c_229_n 0.0142364f $X=-0.19 $Y=-0.245 $X2=2.61 $Y2=1.235
cc_21 VNB N_X_c_266_n 0.0248845f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_22 VNB N_X_c_267_n 0.00743257f $X=-0.19 $Y=-0.245 $X2=2.28 $Y2=1.235
cc_23 VNB N_X_c_268_n 0.0221277f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.515
cc_24 VNB N_VPWR_c_288_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_362_n 0.0209501f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_26 VNB N_VGND_c_363_n 0.0120067f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.87
cc_27 VNB N_VGND_c_364_n 0.0295961f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.87
cc_28 VNB N_VGND_c_365_n 0.00921063f $X=-0.19 $Y=-0.245 $X2=2.445 $Y2=0.955
cc_29 VNB N_VGND_c_366_n 0.0196766f $X=-0.19 $Y=-0.245 $X2=2.61 $Y2=1.235
cc_30 VNB N_VGND_c_367_n 0.0448011f $X=-0.19 $Y=-0.245 $X2=2.93 $Y2=2.815
cc_31 VNB N_VGND_c_368_n 0.0111562f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_369_n 0.219881f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VPB N_A_81_270#_c_57_n 0.0349277f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.765
cc_34 VPB N_A_81_270#_c_61_n 0.0568318f $X=-0.19 $Y=1.66 $X2=2.93 $Y2=2.105
cc_35 VPB N_A_81_270#_c_62_n 0.00341417f $X=-0.19 $Y=1.66 $X2=0.625 $Y2=1.235
cc_36 VPB N_A3_c_130_n 0.0373158f $X=-0.19 $Y=1.66 $X2=2.225 $Y2=0.615
cc_37 VPB A3 0.00257381f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_38 VPB N_A2_c_163_n 0.0372541f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_39 VPB A2 0.00138051f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_40 VPB N_A1_c_193_n 0.0350146f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_41 VPB A1 0.00235147f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_42 VPB N_B1_c_225_n 0.00764796f $X=-0.19 $Y=1.66 $X2=2.78 $Y2=1.96
cc_43 VPB N_B1_c_231_n 0.0258306f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_44 VPB X 0.00695105f $X=-0.19 $Y=1.66 $X2=0.825 $Y2=1.235
cc_45 VPB X 0.0408286f $X=-0.19 $Y=1.66 $X2=2.93 $Y2=2.105
cc_46 VPB N_X_c_268_n 0.00911725f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=1.515
cc_47 VPB N_VPWR_c_289_n 0.010418f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_48 VPB N_VPWR_c_290_n 0.0098755f $X=-0.19 $Y=1.66 $X2=2.445 $Y2=1.15
cc_49 VPB N_VPWR_c_291_n 0.0186948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_292_n 0.00786036f $X=-0.19 $Y=1.66 $X2=2.845 $Y2=1.235
cc_51 VPB N_VPWR_c_293_n 0.018677f $X=-0.19 $Y=1.66 $X2=2.97 $Y2=2.105
cc_52 VPB N_VPWR_c_294_n 0.0363074f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_288_n 0.0679086f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_296_n 0.0088221f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_A_250_392#_c_328_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_56 VPB N_A_250_392#_c_329_n 0.00257348f $X=-0.19 $Y=1.66 $X2=2.445 $Y2=1.15
cc_57 N_A_81_270#_c_57_n N_A3_c_130_n 0.0334861f $X=0.495 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_58 N_A_81_270#_c_59_n N_A3_c_130_n 0.00445011f $X=2.28 $Y=1.235 $X2=-0.19
+ $Y2=-0.245
cc_59 N_A_81_270#_c_62_n N_A3_c_130_n 0.00117732f $X=0.625 $Y=1.235 $X2=-0.19
+ $Y2=-0.245
cc_60 N_A_81_270#_c_57_n N_A3_M1008_g 0.00287123f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_61 N_A_81_270#_c_58_n N_A3_M1008_g 0.00806675f $X=0.51 $Y=1.35 $X2=0 $Y2=0
cc_62 N_A_81_270#_c_59_n N_A3_M1008_g 0.0149586f $X=2.28 $Y=1.235 $X2=0 $Y2=0
cc_63 N_A_81_270#_c_62_n N_A3_M1008_g 0.00309045f $X=0.625 $Y=1.235 $X2=0 $Y2=0
cc_64 N_A_81_270#_c_57_n A3 8.94439e-19 $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_65 N_A_81_270#_c_59_n A3 0.0241217f $X=2.28 $Y=1.235 $X2=0 $Y2=0
cc_66 N_A_81_270#_c_62_n A3 0.0153381f $X=0.625 $Y=1.235 $X2=0 $Y2=0
cc_67 N_A_81_270#_c_59_n N_A2_M1003_g 0.0127685f $X=2.28 $Y=1.235 $X2=0 $Y2=0
cc_68 N_A_81_270#_c_59_n N_A2_c_163_n 0.00421126f $X=2.28 $Y=1.235 $X2=0 $Y2=0
cc_69 N_A_81_270#_c_59_n A2 0.024098f $X=2.28 $Y=1.235 $X2=0 $Y2=0
cc_70 N_A_81_270#_c_59_n N_A1_M1009_g 0.0134426f $X=2.28 $Y=1.235 $X2=0 $Y2=0
cc_71 N_A_81_270#_c_59_n N_A1_c_193_n 0.00148156f $X=2.28 $Y=1.235 $X2=0 $Y2=0
cc_72 N_A_81_270#_c_63_n N_A1_c_193_n 0.00317136f $X=2.445 $Y=1.235 $X2=0 $Y2=0
cc_73 N_A_81_270#_c_59_n A1 0.0171013f $X=2.28 $Y=1.235 $X2=0 $Y2=0
cc_74 N_A_81_270#_c_61_n A1 0.0117728f $X=2.93 $Y=2.105 $X2=0 $Y2=0
cc_75 N_A_81_270#_c_63_n A1 0.0102517f $X=2.445 $Y=1.235 $X2=0 $Y2=0
cc_76 N_A_81_270#_c_61_n N_B1_c_225_n 0.00934319f $X=2.93 $Y=2.105 $X2=0 $Y2=0
cc_77 N_A_81_270#_c_61_n N_B1_c_231_n 0.00706625f $X=2.93 $Y=2.105 $X2=0 $Y2=0
cc_78 N_A_81_270#_c_60_n N_B1_M1000_g 0.0184208f $X=2.845 $Y=1.235 $X2=0 $Y2=0
cc_79 N_A_81_270#_c_61_n N_B1_M1000_g 0.00983966f $X=2.93 $Y=2.105 $X2=0 $Y2=0
cc_80 N_A_81_270#_c_60_n N_B1_c_227_n 0.00184241f $X=2.845 $Y=1.235 $X2=0 $Y2=0
cc_81 N_A_81_270#_c_91_p N_B1_c_228_n 6.83819e-19 $X=2.445 $Y=0.955 $X2=0 $Y2=0
cc_82 N_A_81_270#_M1009_d N_B1_c_229_n 0.00355368f $X=2.225 $Y=0.615 $X2=0 $Y2=0
cc_83 N_A_81_270#_c_59_n N_B1_c_229_n 0.0174185f $X=2.28 $Y=1.235 $X2=0 $Y2=0
cc_84 N_A_81_270#_c_91_p N_B1_c_229_n 0.0266869f $X=2.445 $Y=0.955 $X2=0 $Y2=0
cc_85 N_A_81_270#_c_60_n N_B1_c_229_n 0.00368593f $X=2.845 $Y=1.235 $X2=0 $Y2=0
cc_86 N_A_81_270#_c_58_n N_X_c_266_n 0.00629257f $X=0.51 $Y=1.35 $X2=0 $Y2=0
cc_87 N_A_81_270#_c_58_n N_X_c_267_n 0.00702486f $X=0.51 $Y=1.35 $X2=0 $Y2=0
cc_88 N_A_81_270#_c_62_n N_X_c_267_n 0.00146264f $X=0.625 $Y=1.235 $X2=0 $Y2=0
cc_89 N_A_81_270#_c_57_n X 0.00322907f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_90 N_A_81_270#_c_62_n X 7.22171e-19 $X=0.625 $Y=1.235 $X2=0 $Y2=0
cc_91 N_A_81_270#_c_57_n X 0.0102397f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_92 N_A_81_270#_c_57_n N_X_c_268_n 0.0118864f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_93 N_A_81_270#_c_58_n N_X_c_268_n 0.00249972f $X=0.51 $Y=1.35 $X2=0 $Y2=0
cc_94 N_A_81_270#_c_62_n N_X_c_268_n 0.0307829f $X=0.625 $Y=1.235 $X2=0 $Y2=0
cc_95 N_A_81_270#_c_57_n N_VPWR_c_289_n 0.0122001f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_96 N_A_81_270#_c_59_n N_VPWR_c_289_n 0.00527561f $X=2.28 $Y=1.235 $X2=0 $Y2=0
cc_97 N_A_81_270#_c_62_n N_VPWR_c_289_n 0.0120968f $X=0.625 $Y=1.235 $X2=0 $Y2=0
cc_98 N_A_81_270#_c_57_n N_VPWR_c_293_n 0.00445602f $X=0.495 $Y=1.765 $X2=0
+ $Y2=0
cc_99 N_A_81_270#_c_61_n N_VPWR_c_294_n 0.011066f $X=2.93 $Y=2.105 $X2=0 $Y2=0
cc_100 N_A_81_270#_c_57_n N_VPWR_c_288_n 0.00862155f $X=0.495 $Y=1.765 $X2=0
+ $Y2=0
cc_101 N_A_81_270#_c_61_n N_VPWR_c_288_n 0.00915947f $X=2.93 $Y=2.105 $X2=0
+ $Y2=0
cc_102 N_A_81_270#_c_59_n N_A_250_392#_c_330_n 0.00586046f $X=2.28 $Y=1.235
+ $X2=0 $Y2=0
cc_103 N_A_81_270#_c_59_n N_A_250_392#_c_331_n 0.00507286f $X=2.28 $Y=1.235
+ $X2=0 $Y2=0
cc_104 N_A_81_270#_c_60_n N_A_250_392#_c_332_n 6.87169e-19 $X=2.845 $Y=1.235
+ $X2=0 $Y2=0
cc_105 N_A_81_270#_c_61_n N_A_250_392#_c_332_n 0.0121024f $X=2.93 $Y=2.105 $X2=0
+ $Y2=0
cc_106 N_A_81_270#_c_63_n N_A_250_392#_c_332_n 0.00633471f $X=2.445 $Y=1.235
+ $X2=0 $Y2=0
cc_107 N_A_81_270#_c_61_n N_A_250_392#_c_329_n 0.0563195f $X=2.93 $Y=2.105 $X2=0
+ $Y2=0
cc_108 N_A_81_270#_c_59_n N_VGND_M1005_d 0.00351422f $X=2.28 $Y=1.235 $X2=-0.19
+ $Y2=-0.245
cc_109 N_A_81_270#_c_62_n N_VGND_M1005_d 0.00221237f $X=0.625 $Y=1.235 $X2=-0.19
+ $Y2=-0.245
cc_110 N_A_81_270#_c_60_n N_VGND_M1000_d 0.00280144f $X=2.845 $Y=1.235 $X2=0
+ $Y2=0
cc_111 N_A_81_270#_c_57_n N_VGND_c_362_n 6.25171e-19 $X=0.495 $Y=1.765 $X2=0
+ $Y2=0
cc_112 N_A_81_270#_c_58_n N_VGND_c_362_n 0.00650193f $X=0.51 $Y=1.35 $X2=0 $Y2=0
cc_113 N_A_81_270#_c_59_n N_VGND_c_362_n 0.0255877f $X=2.28 $Y=1.235 $X2=0 $Y2=0
cc_114 N_A_81_270#_c_62_n N_VGND_c_362_n 0.0162002f $X=0.625 $Y=1.235 $X2=0
+ $Y2=0
cc_115 N_A_81_270#_c_60_n N_VGND_c_365_n 0.0198501f $X=2.845 $Y=1.235 $X2=0
+ $Y2=0
cc_116 N_A_81_270#_c_58_n N_VGND_c_366_n 0.00475875f $X=0.51 $Y=1.35 $X2=0 $Y2=0
cc_117 N_A_81_270#_c_58_n N_VGND_c_369_n 0.00505379f $X=0.51 $Y=1.35 $X2=0 $Y2=0
cc_118 N_A_81_270#_c_59_n A_265_120# 0.00366293f $X=2.28 $Y=1.235 $X2=-0.19
+ $Y2=-0.245
cc_119 N_A_81_270#_c_59_n A_337_120# 0.00521091f $X=2.28 $Y=1.235 $X2=-0.19
+ $Y2=-0.245
cc_120 N_A3_M1008_g N_A2_M1003_g 0.0416465f $X=1.25 $Y=0.92 $X2=0 $Y2=0
cc_121 N_A3_c_130_n N_A2_c_163_n 0.0548505f $X=1.175 $Y=1.885 $X2=0 $Y2=0
cc_122 A3 N_A2_c_163_n 0.0010743f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_123 N_A3_c_130_n A2 3.89032e-19 $X=1.175 $Y=1.885 $X2=0 $Y2=0
cc_124 A3 A2 0.0196026f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_125 N_A3_M1008_g N_B1_c_229_n 5.34903e-19 $X=1.25 $Y=0.92 $X2=0 $Y2=0
cc_126 N_A3_c_130_n X 6.62132e-19 $X=1.175 $Y=1.885 $X2=0 $Y2=0
cc_127 N_A3_c_130_n N_VPWR_c_289_n 0.0112253f $X=1.175 $Y=1.885 $X2=0 $Y2=0
cc_128 A3 N_VPWR_c_289_n 0.00473079f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_129 N_A3_c_130_n N_VPWR_c_291_n 0.00445602f $X=1.175 $Y=1.885 $X2=0 $Y2=0
cc_130 N_A3_c_130_n N_VPWR_c_288_n 0.00858778f $X=1.175 $Y=1.885 $X2=0 $Y2=0
cc_131 N_A3_c_130_n N_A_250_392#_c_330_n 0.00337298f $X=1.175 $Y=1.885 $X2=0
+ $Y2=0
cc_132 A3 N_A_250_392#_c_330_n 0.0047583f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_133 N_A3_c_130_n N_A_250_392#_c_328_n 0.0085477f $X=1.175 $Y=1.885 $X2=0
+ $Y2=0
cc_134 N_A3_M1008_g N_VGND_c_362_n 0.013823f $X=1.25 $Y=0.92 $X2=0 $Y2=0
cc_135 N_A3_M1008_g N_VGND_c_367_n 0.00356352f $X=1.25 $Y=0.92 $X2=0 $Y2=0
cc_136 N_A3_M1008_g N_VGND_c_369_n 0.00400172f $X=1.25 $Y=0.92 $X2=0 $Y2=0
cc_137 N_A2_M1003_g N_A1_M1009_g 0.0326149f $X=1.61 $Y=0.92 $X2=0 $Y2=0
cc_138 N_A2_c_163_n N_A1_c_193_n 0.0455825f $X=1.625 $Y=1.885 $X2=0 $Y2=0
cc_139 A2 N_A1_c_193_n 3.63175e-19 $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_140 N_A2_c_163_n A1 0.00175997f $X=1.625 $Y=1.885 $X2=0 $Y2=0
cc_141 A2 A1 0.0236226f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_142 N_A2_M1003_g N_B1_c_229_n 0.0115129f $X=1.61 $Y=0.92 $X2=0 $Y2=0
cc_143 N_A2_c_163_n N_VPWR_c_290_n 0.00667156f $X=1.625 $Y=1.885 $X2=0 $Y2=0
cc_144 N_A2_c_163_n N_VPWR_c_291_n 0.00445602f $X=1.625 $Y=1.885 $X2=0 $Y2=0
cc_145 N_A2_c_163_n N_VPWR_c_288_n 0.00858468f $X=1.625 $Y=1.885 $X2=0 $Y2=0
cc_146 N_A2_c_163_n N_A_250_392#_c_330_n 4.2644e-19 $X=1.625 $Y=1.885 $X2=0
+ $Y2=0
cc_147 A2 N_A_250_392#_c_330_n 0.0016817f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_148 N_A2_c_163_n N_A_250_392#_c_328_n 0.0103402f $X=1.625 $Y=1.885 $X2=0
+ $Y2=0
cc_149 N_A2_c_163_n N_A_250_392#_c_331_n 0.0137172f $X=1.625 $Y=1.885 $X2=0
+ $Y2=0
cc_150 A2 N_A_250_392#_c_331_n 0.0196417f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_151 N_A2_c_163_n N_A_250_392#_c_329_n 8.5062e-19 $X=1.625 $Y=1.885 $X2=0
+ $Y2=0
cc_152 N_A2_M1003_g N_VGND_c_362_n 0.00212757f $X=1.61 $Y=0.92 $X2=0 $Y2=0
cc_153 N_A2_M1003_g N_VGND_c_367_n 0.0013085f $X=1.61 $Y=0.92 $X2=0 $Y2=0
cc_154 N_A2_M1003_g N_VGND_c_369_n 9.5279e-19 $X=1.61 $Y=0.92 $X2=0 $Y2=0
cc_155 N_A1_c_193_n N_B1_c_231_n 0.0130041f $X=2.255 $Y=1.885 $X2=0 $Y2=0
cc_156 N_A1_M1009_g N_B1_M1000_g 0.0223483f $X=2.15 $Y=0.935 $X2=0 $Y2=0
cc_157 N_A1_M1009_g N_B1_c_227_n 0.00117875f $X=2.15 $Y=0.935 $X2=0 $Y2=0
cc_158 N_A1_c_193_n N_B1_c_227_n 0.0200275f $X=2.255 $Y=1.885 $X2=0 $Y2=0
cc_159 A1 N_B1_c_227_n 0.00114125f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_160 N_A1_M1009_g N_B1_c_228_n 9.92136e-19 $X=2.15 $Y=0.935 $X2=0 $Y2=0
cc_161 N_A1_M1009_g N_B1_c_229_n 0.013629f $X=2.15 $Y=0.935 $X2=0 $Y2=0
cc_162 N_A1_c_193_n N_VPWR_c_290_n 0.00812936f $X=2.255 $Y=1.885 $X2=0 $Y2=0
cc_163 N_A1_c_193_n N_VPWR_c_294_n 0.00445602f $X=2.255 $Y=1.885 $X2=0 $Y2=0
cc_164 N_A1_c_193_n N_VPWR_c_288_n 0.00858468f $X=2.255 $Y=1.885 $X2=0 $Y2=0
cc_165 N_A1_c_193_n N_A_250_392#_c_328_n 8.5062e-19 $X=2.255 $Y=1.885 $X2=0
+ $Y2=0
cc_166 N_A1_c_193_n N_A_250_392#_c_331_n 0.0150443f $X=2.255 $Y=1.885 $X2=0
+ $Y2=0
cc_167 A1 N_A_250_392#_c_331_n 0.0175308f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_168 N_A1_c_193_n N_A_250_392#_c_332_n 0.00169682f $X=2.255 $Y=1.885 $X2=0
+ $Y2=0
cc_169 A1 N_A_250_392#_c_332_n 0.0047583f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_170 N_A1_c_193_n N_A_250_392#_c_329_n 0.0103402f $X=2.255 $Y=1.885 $X2=0
+ $Y2=0
cc_171 N_A1_M1009_g N_VGND_c_367_n 5.46057e-19 $X=2.15 $Y=0.935 $X2=0 $Y2=0
cc_172 N_B1_c_231_n N_VPWR_c_294_n 0.00445602f $X=2.705 $Y=1.885 $X2=0 $Y2=0
cc_173 N_B1_c_231_n N_VPWR_c_288_n 0.0086233f $X=2.705 $Y=1.885 $X2=0 $Y2=0
cc_174 N_B1_c_231_n N_A_250_392#_c_332_n 0.00219514f $X=2.705 $Y=1.885 $X2=0
+ $Y2=0
cc_175 N_B1_c_231_n N_A_250_392#_c_329_n 0.00938763f $X=2.705 $Y=1.885 $X2=0
+ $Y2=0
cc_176 N_B1_c_229_n N_VGND_c_362_n 0.0192005f $X=2.65 $Y=0.34 $X2=0 $Y2=0
cc_177 N_B1_M1000_g N_VGND_c_364_n 0.00399579f $X=2.74 $Y=0.935 $X2=0 $Y2=0
cc_178 N_B1_c_228_n N_VGND_c_364_n 0.00511411f $X=2.65 $Y=0.34 $X2=0 $Y2=0
cc_179 N_B1_c_229_n N_VGND_c_364_n 0.0305341f $X=2.65 $Y=0.34 $X2=0 $Y2=0
cc_180 N_B1_M1000_g N_VGND_c_365_n 0.00244045f $X=2.74 $Y=0.935 $X2=0 $Y2=0
cc_181 N_B1_c_229_n N_VGND_c_365_n 0.00172851f $X=2.65 $Y=0.34 $X2=0 $Y2=0
cc_182 N_B1_c_228_n N_VGND_c_367_n 0.00659816f $X=2.65 $Y=0.34 $X2=0 $Y2=0
cc_183 N_B1_c_229_n N_VGND_c_367_n 0.084256f $X=2.65 $Y=0.34 $X2=0 $Y2=0
cc_184 N_B1_c_228_n N_VGND_c_369_n 0.0102618f $X=2.65 $Y=0.34 $X2=0 $Y2=0
cc_185 N_B1_c_229_n N_VGND_c_369_n 0.0463662f $X=2.65 $Y=0.34 $X2=0 $Y2=0
cc_186 N_B1_c_229_n A_337_120# 0.00524643f $X=2.65 $Y=0.34 $X2=-0.19 $Y2=-0.245
cc_187 X N_VPWR_c_289_n 0.0390338f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_188 X N_VPWR_c_293_n 0.0154862f $X=0.24 $Y=2.035 $X2=0 $Y2=0
cc_189 X N_VPWR_c_288_n 0.0127853f $X=0.24 $Y=2.035 $X2=0 $Y2=0
cc_190 N_X_c_266_n N_VGND_c_362_n 0.0199137f $X=0.295 $Y=0.645 $X2=0 $Y2=0
cc_191 N_X_c_266_n N_VGND_c_366_n 0.0105642f $X=0.295 $Y=0.645 $X2=0 $Y2=0
cc_192 N_X_c_266_n N_VGND_c_369_n 0.0123086f $X=0.295 $Y=0.645 $X2=0 $Y2=0
cc_193 N_VPWR_c_289_n N_A_250_392#_c_328_n 0.0323125f $X=0.835 $Y=2.135 $X2=0
+ $Y2=0
cc_194 N_VPWR_c_290_n N_A_250_392#_c_328_n 0.0259568f $X=1.94 $Y=2.42 $X2=0
+ $Y2=0
cc_195 N_VPWR_c_291_n N_A_250_392#_c_328_n 0.014552f $X=1.735 $Y=3.33 $X2=0
+ $Y2=0
cc_196 N_VPWR_c_288_n N_A_250_392#_c_328_n 0.0119791f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_197 N_VPWR_M1007_d N_A_250_392#_c_331_n 0.0103211f $X=1.7 $Y=1.96 $X2=0 $Y2=0
cc_198 N_VPWR_c_290_n N_A_250_392#_c_331_n 0.0297772f $X=1.94 $Y=2.42 $X2=0
+ $Y2=0
cc_199 N_VPWR_c_290_n N_A_250_392#_c_329_n 0.0259568f $X=1.94 $Y=2.42 $X2=0
+ $Y2=0
cc_200 N_VPWR_c_294_n N_A_250_392#_c_329_n 0.014552f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_201 N_VPWR_c_288_n N_A_250_392#_c_329_n 0.0119791f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
