* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__ha_4 A B VGND VNB VPB VPWR COUT SUM
M1000 VGND B a_27_125# VNB nshort w=640000u l=150000u
+  ad=1.6734e+12p pd=1.601e+07u as=7.744e+11p ps=7.54e+06u
M1001 a_707_119# B a_435_99# VNB nshort w=640000u l=150000u
+  ad=5.856e+11p pd=5.67e+06u as=1.792e+11p ps=1.84e+06u
M1002 VGND A a_707_119# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VGND a_294_392# SUM VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=5.069e+11p ps=4.33e+06u
M1004 a_27_125# B VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 SUM a_294_392# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=9.632e+11p pd=6.2e+06u as=2.9278e+12p ps=2.402e+07u
M1006 VGND a_435_99# COUT VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=4.144e+11p ps=4.08e+06u
M1007 a_294_392# B a_27_392# VPB phighvt w=1e+06u l=150000u
+  ad=5.52e+11p pd=4.88e+06u as=8.7e+11p ps=7.74e+06u
M1008 a_707_119# A VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_294_392# a_435_99# VPWR VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND a_435_99# COUT VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_27_125# A VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR B a_435_99# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=7.96825e+11p ps=6.01e+06u
M1013 VPWR a_294_392# SUM VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_27_392# B a_294_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 SUM a_294_392# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR a_435_99# a_294_392# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 COUT a_435_99# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=8.512e+11p pd=6e+06u as=0p ps=0u
M1018 VPWR A a_435_99# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_435_99# A VPWR VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 SUM a_294_392# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND A a_27_125# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_294_392# a_435_99# a_27_125# VNB nshort w=640000u l=150000u
+  ad=2.048e+11p pd=1.92e+06u as=0p ps=0u
M1023 a_435_99# B VPWR VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 SUM a_294_392# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 COUT a_435_99# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_27_125# a_435_99# a_294_392# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VGND a_294_392# SUM VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 COUT a_435_99# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPWR a_294_392# SUM VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 COUT a_435_99# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VPWR a_435_99# COUT VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 VPWR a_435_99# COUT VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VPWR A a_27_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_27_392# A VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_435_99# B a_707_119# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
