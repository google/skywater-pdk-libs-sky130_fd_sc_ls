* File: sky130_fd_sc_ls__nor3_1.pex.spice
* Created: Fri Aug 28 13:38:10 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__NOR3_1%A 1 3 4 6 7 8
r28 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.385 $X2=0.27 $Y2=1.385
r29 8 13 12.6543 $w=2.53e-07 $l=2.8e-07 $layer=LI1_cond $X=0.232 $Y=1.665
+ $X2=0.232 $Y2=1.385
r30 7 13 4.06745 $w=2.53e-07 $l=9e-08 $layer=LI1_cond $X=0.232 $Y=1.295
+ $X2=0.232 $Y2=1.385
r31 4 12 67.6304 $w=3.61e-07 $l=4.48776e-07 $layer=POLY_cond $X=0.495 $Y=1.765
+ $X2=0.345 $Y2=1.385
r32 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.495 $Y=1.765
+ $X2=0.495 $Y2=2.4
r33 1 12 38.924 $w=3.61e-07 $l=2.2798e-07 $layer=POLY_cond $X=0.495 $Y=1.22
+ $X2=0.345 $Y2=1.385
r34 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.495 $Y=1.22 $X2=0.495
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__NOR3_1%B 1 3 6 8
r33 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.96
+ $Y=1.465 $X2=0.96 $Y2=1.465
r34 8 12 5.98039 $w=4.78e-07 $l=2.4e-07 $layer=LI1_cond $X=1.2 $Y=1.54 $X2=0.96
+ $Y2=1.54
r35 4 11 38.6549 $w=2.86e-07 $l=1.81659e-07 $layer=POLY_cond $X=0.925 $Y=1.3
+ $X2=0.96 $Y2=1.465
r36 4 6 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.925 $Y=1.3 $X2=0.925
+ $Y2=0.74
r37 1 11 61.4066 $w=2.86e-07 $l=3.21714e-07 $layer=POLY_cond $X=0.915 $Y=1.765
+ $X2=0.96 $Y2=1.465
r38 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.915 $Y=1.765
+ $X2=0.915 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__NOR3_1%C 3 5 7 8 12
r21 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.65
+ $Y=1.465 $X2=1.65 $Y2=1.465
r22 8 12 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=1.65 $Y=1.665 $X2=1.65
+ $Y2=1.465
r23 5 11 56.0318 $w=3.92e-07 $l=3.67423e-07 $layer=POLY_cond $X=1.425 $Y=1.765
+ $X2=1.575 $Y2=1.465
r24 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.425 $Y=1.765
+ $X2=1.425 $Y2=2.4
r25 1 11 39.4323 $w=3.92e-07 $l=2.2798e-07 $layer=POLY_cond $X=1.425 $Y=1.3
+ $X2=1.575 $Y2=1.465
r26 1 3 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.425 $Y=1.3 $X2=1.425
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__NOR3_1%VPWR 1 6 9 11 13 20 21
r24 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r25 20 21 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r26 18 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r27 17 20 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=3.33 $X2=1.68
+ $Y2=3.33
r28 17 18 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r29 15 24 4.75569 $w=1.7e-07 $l=2.18e-07 $layer=LI1_cond $X=0.435 $Y=3.33
+ $X2=0.217 $Y2=3.33
r30 15 17 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.435 $Y=3.33
+ $X2=0.72 $Y2=3.33
r31 13 21 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=1.68 $Y2=3.33
r32 13 18 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=0.72 $Y2=3.33
r33 11 12 5.24459 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=0.27 $Y=2.455
+ $X2=0.27 $Y2=2.325
r34 9 24 3.01048 $w=3.3e-07 $l=1.08305e-07 $layer=LI1_cond $X=0.27 $Y=3.245
+ $X2=0.217 $Y2=3.33
r35 8 11 1.22229 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=0.27 $Y=2.49 $X2=0.27
+ $Y2=2.455
r36 8 9 26.3665 $w=3.28e-07 $l=7.55e-07 $layer=LI1_cond $X=0.27 $Y=2.49 $X2=0.27
+ $Y2=3.245
r37 6 12 9.68052 $w=2.48e-07 $l=2.1e-07 $layer=LI1_cond $X=0.23 $Y=2.115
+ $X2=0.23 $Y2=2.325
r38 1 11 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.84 $X2=0.27 $Y2=2.455
r39 1 6 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.27 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_LS__NOR3_1%Y 1 2 3 11 14 16 20 23 24 25 26 33
r48 31 33 0.236893 $w=1.028e-06 $l=2e-08 $layer=LI1_cond $X=0.7 $Y=2.465
+ $X2=0.72 $Y2=2.465
r49 26 38 0.35534 $w=1.028e-06 $l=3e-08 $layer=LI1_cond $X=1.68 $Y=2.465
+ $X2=1.65 $Y2=2.465
r50 25 38 5.3301 $w=1.028e-06 $l=4.5e-07 $layer=LI1_cond $X=1.2 $Y=2.465
+ $X2=1.65 $Y2=2.465
r51 24 31 1.83245 $w=1.03e-06 $l=8.5e-08 $layer=LI1_cond $X=0.615 $Y=2.465
+ $X2=0.7 $Y2=2.465
r52 24 25 5.30641 $w=1.028e-06 $l=4.48e-07 $layer=LI1_cond $X=0.752 $Y=2.465
+ $X2=1.2 $Y2=2.465
r53 24 33 0.379029 $w=1.028e-06 $l=3.2e-08 $layer=LI1_cond $X=0.752 $Y=2.465
+ $X2=0.72 $Y2=2.465
r54 18 20 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=1.64 $Y=0.88
+ $X2=1.64 $Y2=0.515
r55 17 23 0.191034 $w=2.5e-07 $l=1.38e-07 $layer=LI1_cond $X=0.805 $Y=1.005
+ $X2=0.667 $Y2=1.005
r56 16 18 6.98653 $w=2.5e-07 $l=2.18746e-07 $layer=LI1_cond $X=1.475 $Y=1.005
+ $X2=1.64 $Y2=0.88
r57 16 17 30.8855 $w=2.48e-07 $l=6.7e-07 $layer=LI1_cond $X=1.475 $Y=1.005
+ $X2=0.805 $Y2=1.005
r58 12 23 6.72674 $w=1.8e-07 $l=1.44914e-07 $layer=LI1_cond $X=0.71 $Y=0.88
+ $X2=0.667 $Y2=1.005
r59 12 14 20.4306 $w=1.88e-07 $l=3.5e-07 $layer=LI1_cond $X=0.71 $Y=0.88
+ $X2=0.71 $Y2=0.53
r60 11 24 11.1025 $w=1.7e-07 $l=5.15e-07 $layer=LI1_cond $X=0.615 $Y=1.95
+ $X2=0.615 $Y2=2.465
r61 10 23 6.72674 $w=1.8e-07 $l=1.48745e-07 $layer=LI1_cond $X=0.615 $Y=1.13
+ $X2=0.667 $Y2=1.005
r62 10 11 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=0.615 $Y=1.13
+ $X2=0.615 $Y2=1.95
r63 3 38 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.5
+ $Y=1.84 $X2=1.65 $Y2=2.815
r64 3 38 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=1.5
+ $Y=1.84 $X2=1.65 $Y2=2.115
r65 2 20 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.5
+ $Y=0.37 $X2=1.64 $Y2=0.515
r66 1 23 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.965
r67 1 14 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.53
.ends

.subckt PM_SKY130_FD_SC_LS__NOR3_1%VGND 1 2 7 10 13 17 19 20 22 29 30 36
r34 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r35 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r36 30 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r37 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r38 27 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.305 $Y=0 $X2=1.14
+ $Y2=0
r39 27 29 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.305 $Y=0 $X2=1.68
+ $Y2=0
r40 26 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r41 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r42 23 33 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.222
+ $Y2=0
r43 23 25 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.72
+ $Y2=0
r44 22 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.975 $Y=0 $X2=1.14
+ $Y2=0
r45 22 25 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.975 $Y=0 $X2=0.72
+ $Y2=0
r46 20 37 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=1.2
+ $Y2=0
r47 20 26 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=0.72
+ $Y2=0
r48 15 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=0.085
+ $X2=1.14 $Y2=0
r49 15 17 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=1.14 $Y=0.085
+ $X2=1.14 $Y2=0.53
r50 13 19 6.3502 $w=2.43e-07 $l=1.35e-07 $layer=LI1_cond $X=0.237 $Y=0.845
+ $X2=0.237 $Y2=0.71
r51 8 19 6.55101 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.28 $Y=0.545
+ $X2=0.28 $Y2=0.71
r52 8 10 1.3969 $w=3.28e-07 $l=4e-08 $layer=LI1_cond $X=0.28 $Y=0.545 $X2=0.28
+ $Y2=0.505
r53 7 33 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.222 $Y2=0
r54 7 10 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.28 $Y2=0.505
r55 2 17 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=1 $Y=0.37
+ $X2=1.14 $Y2=0.53
r56 1 13 182 $w=1.7e-07 $l=5.40486e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.275 $Y2=0.845
r57 1 10 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.505
.ends

