* File: sky130_fd_sc_ls__and4_1.pex.spice
* Created: Wed Sep  2 10:55:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__AND4_1%A 2 3 5 8 10 11 13 14 15 19 20
c40 2 0 8.64864e-20 $X=0.555 $Y=1.955
r41 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.59
+ $Y=1.285 $X2=0.59 $Y2=1.285
r42 14 15 10.9334 $w=3.88e-07 $l=3.7e-07 $layer=LI1_cond $X=0.62 $Y=1.295
+ $X2=0.62 $Y2=1.665
r43 14 20 0.295498 $w=3.88e-07 $l=1e-08 $layer=LI1_cond $X=0.62 $Y=1.295
+ $X2=0.62 $Y2=1.285
r44 12 19 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.59 $Y=1.625
+ $X2=0.59 $Y2=1.285
r45 12 13 36.5727 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.59 $Y=1.625
+ $X2=0.59 $Y2=1.79
r46 11 19 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=0.59 $Y=1.235 $X2=0.59
+ $Y2=1.285
r47 10 11 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=0.66 $Y=1.085
+ $X2=0.66 $Y2=1.235
r48 8 10 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.82 $Y=0.69
+ $X2=0.82 $Y2=1.085
r49 3 5 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.555 $Y=2.045
+ $X2=0.555 $Y2=2.54
r50 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.555 $Y=1.955 $X2=0.555
+ $Y2=2.045
r51 2 13 64.1371 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.555 $Y=1.955
+ $X2=0.555 $Y2=1.79
.ends

.subckt PM_SKY130_FD_SC_LS__AND4_1%B 2 3 5 8 10 11 12 13 19
c42 10 0 1.73901e-19 $X=1.2 $Y=0.555
r43 19 22 40.7727 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.14 $Y=1.64
+ $X2=1.14 $Y2=1.805
r44 19 21 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.14 $Y=1.64
+ $X2=1.14 $Y2=1.475
r45 13 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.15
+ $Y=1.64 $X2=1.15 $Y2=1.64
r46 12 13 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=1.15 $Y=1.295
+ $X2=1.15 $Y2=1.64
r47 11 12 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.15 $Y=0.925
+ $X2=1.15 $Y2=1.295
r48 10 11 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.15 $Y=0.555
+ $X2=1.15 $Y2=0.925
r49 8 21 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=1.21 $Y=0.69
+ $X2=1.21 $Y2=1.475
r50 3 5 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.055 $Y=2.045
+ $X2=1.055 $Y2=2.54
r51 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.055 $Y=1.955 $X2=1.055
+ $Y2=2.045
r52 2 22 58.3064 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=1.055 $Y=1.955
+ $X2=1.055 $Y2=1.805
.ends

.subckt PM_SKY130_FD_SC_LS__AND4_1%C 3 5 6 8 10 11 12 13 14 15 16 22
c44 13 0 1.66221e-19 $X=1.68 $Y=0.555
c45 5 0 8.74143e-20 $X=1.765 $Y=1.955
r46 15 16 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=1.69 $Y=1.285
+ $X2=1.69 $Y2=1.665
r47 15 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.69
+ $Y=1.285 $X2=1.69 $Y2=1.285
r48 14 15 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=1.69 $Y=0.925
+ $X2=1.69 $Y2=1.285
r49 13 14 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.69 $Y=0.555
+ $X2=1.69 $Y2=0.925
r50 11 22 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.69 $Y=1.625
+ $X2=1.69 $Y2=1.285
r51 11 12 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.69 $Y=1.625
+ $X2=1.69 $Y2=1.79
r52 10 22 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.69 $Y=1.12
+ $X2=1.69 $Y2=1.285
r53 6 8 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.765 $Y=2.045
+ $X2=1.765 $Y2=2.54
r54 5 6 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.765 $Y=1.955 $X2=1.765
+ $Y2=2.045
r55 5 12 64.1371 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.765 $Y=1.955
+ $X2=1.765 $Y2=1.79
r56 3 10 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.6 $Y=0.69 $X2=1.6
+ $Y2=1.12
.ends

.subckt PM_SKY130_FD_SC_LS__AND4_1%D 3 6 7 9 10 13 14
c46 7 0 8.35939e-20 $X=2.265 $Y=2.045
c47 6 0 1.66221e-19 $X=2.265 $Y=1.955
r48 13 16 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.23 $Y=1.515
+ $X2=2.23 $Y2=1.68
r49 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.23 $Y=1.515
+ $X2=2.23 $Y2=1.35
r50 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.23
+ $Y=1.515 $X2=2.23 $Y2=1.515
r51 10 14 4.93904 $w=3.48e-07 $l=1.5e-07 $layer=LI1_cond $X=2.22 $Y=1.665
+ $X2=2.22 $Y2=1.515
r52 7 9 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.265 $Y=2.045
+ $X2=2.265 $Y2=2.54
r53 6 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.265 $Y=1.955 $X2=2.265
+ $Y2=2.045
r54 6 16 106.895 $w=1.8e-07 $l=2.75e-07 $layer=POLY_cond $X=2.265 $Y=1.955
+ $X2=2.265 $Y2=1.68
r55 3 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.17 $Y=0.69 $X2=2.17
+ $Y2=1.35
.ends

.subckt PM_SKY130_FD_SC_LS__AND4_1%A_96_74# 1 2 3 12 14 16 18 19 20 23 25 29 31
+ 34 38 40 41 45
r96 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.77
+ $Y=1.485 $X2=2.77 $Y2=1.485
r97 42 45 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=2.655 $Y=1.485
+ $X2=2.77 $Y2=1.485
r98 35 38 8.74444 $w=5.93e-07 $l=4.35e-07 $layer=LI1_cond $X=0.17 $Y=0.652
+ $X2=0.605 $Y2=0.652
r99 33 42 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.655 $Y=1.65
+ $X2=2.655 $Y2=1.485
r100 33 34 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=2.655 $Y=1.65
+ $X2=2.655 $Y2=1.96
r101 32 41 8.61065 $w=1.7e-07 $l=1.68464e-07 $layer=LI1_cond $X=2.205 $Y=2.045
+ $X2=2.04 $Y2=2.052
r102 31 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.57 $Y=2.045
+ $X2=2.655 $Y2=1.96
r103 31 32 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.57 $Y=2.045
+ $X2=2.205 $Y2=2.045
r104 27 41 0.89609 $w=3.3e-07 $l=9.3e-08 $layer=LI1_cond $X=2.04 $Y=2.145
+ $X2=2.04 $Y2=2.052
r105 27 29 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=2.04 $Y=2.145
+ $X2=2.04 $Y2=2.28
r106 26 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=2.06
+ $X2=0.78 $Y2=2.06
r107 25 41 8.61065 $w=1.7e-07 $l=1.68953e-07 $layer=LI1_cond $X=1.875 $Y=2.06
+ $X2=2.04 $Y2=2.052
r108 25 26 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=1.875 $Y=2.06
+ $X2=0.945 $Y2=2.06
r109 21 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=2.145
+ $X2=0.78 $Y2=2.06
r110 21 23 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=0.78 $Y=2.145
+ $X2=0.78 $Y2=2.28
r111 19 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=2.06
+ $X2=0.78 $Y2=2.06
r112 19 20 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=0.615 $Y=2.06
+ $X2=0.255 $Y2=2.06
r113 18 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.17 $Y=1.975
+ $X2=0.255 $Y2=2.06
r114 17 35 8.26286 $w=1.7e-07 $l=2.98e-07 $layer=LI1_cond $X=0.17 $Y=0.95
+ $X2=0.17 $Y2=0.652
r115 17 18 66.8717 $w=1.68e-07 $l=1.025e-06 $layer=LI1_cond $X=0.17 $Y=0.95
+ $X2=0.17 $Y2=1.975
r116 14 46 57.4383 $w=2.94e-07 $l=3.16607e-07 $layer=POLY_cond $X=2.85 $Y=1.765
+ $X2=2.772 $Y2=1.485
r117 14 16 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.85 $Y=1.765
+ $X2=2.85 $Y2=2.4
r118 10 46 38.5845 $w=2.94e-07 $l=2.05925e-07 $layer=POLY_cond $X=2.68 $Y=1.32
+ $X2=2.772 $Y2=1.485
r119 10 12 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.68 $Y=1.32
+ $X2=2.68 $Y2=0.74
r120 3 29 300 $w=1.7e-07 $l=2.68328e-07 $layer=licon1_PDIFF $count=2 $X=1.84
+ $Y=2.12 $X2=2.04 $Y2=2.28
r121 2 23 300 $w=1.7e-07 $l=2.22711e-07 $layer=licon1_PDIFF $count=2 $X=0.63
+ $Y=2.12 $X2=0.78 $Y2=2.28
r122 1 38 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.48
+ $Y=0.37 $X2=0.605 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__AND4_1%VPWR 1 2 3 10 12 16 20 22 24 29 36 37 43 46
r48 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r49 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r50 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r51 37 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r52 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r53 34 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.74 $Y=3.33
+ $X2=2.575 $Y2=3.33
r54 34 36 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=2.74 $Y=3.33
+ $X2=3.12 $Y2=3.33
r55 33 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r56 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r57 30 43 12.4404 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=1.705 $Y=3.33
+ $X2=1.41 $Y2=3.33
r58 30 32 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=1.705 $Y=3.33
+ $X2=2.16 $Y2=3.33
r59 29 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.41 $Y=3.33
+ $X2=2.575 $Y2=3.33
r60 29 32 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.41 $Y=3.33
+ $X2=2.16 $Y2=3.33
r61 28 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r62 28 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r63 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r64 25 40 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.222 $Y2=3.33
r65 25 27 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.72 $Y2=3.33
r66 24 43 12.4404 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=1.115 $Y=3.33
+ $X2=1.41 $Y2=3.33
r67 24 27 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.115 $Y=3.33
+ $X2=0.72 $Y2=3.33
r68 22 33 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r69 22 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r70 18 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.575 $Y=3.245
+ $X2=2.575 $Y2=3.33
r71 18 20 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=2.575 $Y=3.245
+ $X2=2.575 $Y2=2.465
r72 14 43 2.48142 $w=5.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.41 $Y=3.245
+ $X2=1.41 $Y2=3.33
r73 14 16 16.4207 $w=5.88e-07 $l=8.1e-07 $layer=LI1_cond $X=1.41 $Y=3.245
+ $X2=1.41 $Y2=2.435
r74 10 40 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.222 $Y2=3.33
r75 10 12 28.2872 $w=3.28e-07 $l=8.1e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.28 $Y2=2.435
r76 3 20 300 $w=1.7e-07 $l=4.47325e-07 $layer=licon1_PDIFF $count=2 $X=2.34
+ $Y=2.12 $X2=2.575 $Y2=2.465
r77 2 16 300 $w=1.7e-07 $l=4.32926e-07 $layer=licon1_PDIFF $count=2 $X=1.13
+ $Y=2.12 $X2=1.41 $Y2=2.435
r78 1 12 300 $w=1.7e-07 $l=3.80657e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.12 $X2=0.28 $Y2=2.435
.ends

.subckt PM_SKY130_FD_SC_LS__AND4_1%X 1 2 9 14 15 16 17 21
c24 14 0 8.35939e-20 $X=3.075 $Y=1.985
r25 17 27 10.6778 $w=5.43e-07 $l=2.05e-07 $layer=LI1_cond $X=3.002 $Y=0.925
+ $X2=3.002 $Y2=1.13
r26 16 17 8.12016 $w=5.43e-07 $l=3.7e-07 $layer=LI1_cond $X=3.002 $Y=0.555
+ $X2=3.002 $Y2=0.925
r27 16 21 0.877856 $w=5.43e-07 $l=4e-08 $layer=LI1_cond $X=3.002 $Y=0.555
+ $X2=3.002 $Y2=0.515
r28 15 27 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.19 $Y=1.82 $X2=3.19
+ $Y2=1.13
r29 14 15 8.52431 $w=3.63e-07 $l=1.65e-07 $layer=LI1_cond $X=3.092 $Y=1.985
+ $X2=3.092 $Y2=1.82
r30 7 14 0.536754 $w=3.63e-07 $l=1.7e-08 $layer=LI1_cond $X=3.092 $Y=2.002
+ $X2=3.092 $Y2=1.985
r31 7 9 25.6695 $w=3.63e-07 $l=8.13e-07 $layer=LI1_cond $X=3.092 $Y=2.002
+ $X2=3.092 $Y2=2.815
r32 2 14 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.925
+ $Y=1.84 $X2=3.075 $Y2=1.985
r33 2 9 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.925
+ $Y=1.84 $X2=3.075 $Y2=2.815
r34 1 21 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.755
+ $Y=0.37 $X2=2.895 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__AND4_1%VGND 1 6 9 10 11 21 22
r30 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r31 19 22 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r32 18 19 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r33 14 18 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=2.16
+ $Y2=0
r34 14 15 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r35 11 19 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r36 11 15 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.24
+ $Y2=0
r37 9 18 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=2.22 $Y=0 $X2=2.16
+ $Y2=0
r38 9 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.22 $Y=0 $X2=2.385
+ $Y2=0
r39 8 21 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=2.55 $Y=0 $X2=3.12
+ $Y2=0
r40 8 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.55 $Y=0 $X2=2.385
+ $Y2=0
r41 4 10 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.385 $Y=0.085
+ $X2=2.385 $Y2=0
r42 4 6 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.385 $Y=0.085
+ $X2=2.385 $Y2=0.515
r43 1 6 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.245
+ $Y=0.37 $X2=2.385 $Y2=0.515
.ends

