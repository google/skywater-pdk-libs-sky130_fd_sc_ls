* NGSPICE file created from sky130_fd_sc_ls__and3_2.ext - technology: sky130A

.subckt sky130_fd_sc_ls__and3_2 A B C VGND VNB VPB VPWR X
M1000 VPWR A a_41_384# VPB phighvt w=840000u l=150000u
+  ad=1.3306e+12p pd=8.87e+06u as=4.998e+11p ps=4.55e+06u
M1001 X a_41_384# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=0p ps=0u
M1002 VPWR C a_41_384# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VGND C a_247_136# VNB nshort w=640000u l=150000u
+  ad=6.9565e+11p pd=5.12e+06u as=1.536e+11p ps=1.76e+06u
M1004 VPWR a_41_384# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_247_136# B a_133_136# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=2.688e+11p ps=2.12e+06u
M1006 a_133_136# A a_41_384# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1007 VGND a_41_384# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.368e+11p ps=2.12e+06u
M1008 a_41_384# B VPWR VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 X a_41_384# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

