* NGSPICE file created from sky130_fd_sc_ls__a22oi_2.ext - technology: sky130A

.subckt sky130_fd_sc_ls__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
M1000 a_148_74# A2 VGND VNB nshort w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=4.662e+11p ps=4.22e+06u
M1001 Y A1 a_148_74# VNB nshort w=740000u l=150000u
+  ad=7.918e+11p pd=6.58e+06u as=0p ps=0u
M1002 VPWR A1 a_66_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=1.0192e+12p pd=6.3e+06u as=1.624e+12p ps=1.41e+07u
M1003 VGND A2 a_148_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_558_74# B1 Y VNB nshort w=740000u l=150000u
+  ad=4.958e+11p pd=4.3e+06u as=0p ps=0u
M1005 a_66_368# A2 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_66_368# B2 Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=7.056e+11p ps=5.74e+06u
M1007 Y B1 a_558_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_66_368# A1 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND B2 a_558_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR A2 a_66_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Y B2 a_66_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Y B1 a_66_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_66_368# B1 Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_148_74# A1 Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_558_74# B2 VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

