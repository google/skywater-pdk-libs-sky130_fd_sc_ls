* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__sdfbbp_1 CLK D RESET_B SCD SCE SET_B VGND VNB VPB VPWR Q
+ Q_N
X0 a_2037_442# a_1625_93# a_2271_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X1 VGND a_2037_442# Q_N VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X2 a_1250_231# a_1625_93# a_1418_125# VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X3 VPWR a_2881_74# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X4 a_1766_379# a_622_98# a_1878_420# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X5 a_1878_420# a_877_98# a_1986_504# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 a_1986_504# a_2037_442# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 a_1580_379# a_1625_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X8 a_2881_74# a_2037_442# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X9 a_197_119# a_341_93# a_27_464# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X10 a_1880_119# a_877_98# a_1878_420# VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X11 a_197_119# a_877_98# a_1092_96# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X12 VGND SCD a_119_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 a_622_98# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X14 a_1250_231# a_1092_96# a_1580_379# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X15 a_622_98# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X16 a_27_464# SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X17 VPWR SET_B a_1250_231# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X18 VGND a_1250_231# a_1880_119# VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X19 a_2384_392# a_1625_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X20 VGND a_2881_74# Q VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X21 a_1878_420# a_622_98# a_2061_74# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X22 a_2881_74# a_2037_442# VGND VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X23 a_197_119# D a_299_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X24 VPWR a_1250_231# a_1766_379# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X25 a_1092_96# a_877_98# a_1192_96# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X26 VPWR a_2037_442# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X27 VPWR SCE a_218_464# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X28 a_1221_419# a_1250_231# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X29 VGND SET_B a_2271_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X30 a_119_119# SCE a_197_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X31 a_1192_96# a_1250_231# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X32 VGND SET_B a_1418_125# VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X33 a_1092_96# a_622_98# a_1221_419# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X34 VGND SCE a_341_93# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X35 a_1418_125# a_1092_96# a_1250_231# VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X36 a_2061_74# a_2037_442# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X37 a_1625_93# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X38 a_218_464# D a_197_119# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X39 VPWR SCE a_341_93# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X40 VGND a_622_98# a_877_98# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X41 VPWR a_622_98# a_877_98# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X42 a_299_119# a_341_93# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X43 a_197_119# a_622_98# a_1092_96# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X44 VPWR SET_B a_2037_442# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X45 a_2037_442# a_1878_420# a_2384_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X46 a_1625_93# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X47 a_2271_74# a_1878_420# a_2037_442# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
.ends
