* File: sky130_fd_sc_ls__o2111a_1.pex.spice
* Created: Wed Sep  2 11:16:27 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__O2111A_1%A_82_48# 1 2 3 10 12 13 15 17 18 20 21 24
+ 28 32 39 41
c74 32 0 1.4602e-19 $X=0.61 $Y=1.295
c75 24 0 1.39983e-20 $X=1.245 $Y=0.515
c76 18 0 1.10157e-19 $X=1.08 $Y=1.295
r77 35 37 8.48848 $w=3.48e-07 $l=1.65e-07 $layer=LI1_cond $X=0.61 $Y=1.385
+ $X2=0.61 $Y2=1.55
r78 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.6
+ $Y=1.385 $X2=0.6 $Y2=1.385
r79 32 35 2.96342 $w=3.48e-07 $l=9e-08 $layer=LI1_cond $X=0.61 $Y=1.295 $X2=0.61
+ $Y2=1.385
r80 29 39 8.52281 $w=1.72e-07 $l=1.65e-07 $layer=LI1_cond $X=1.525 $Y=2.157
+ $X2=1.36 $Y2=2.157
r81 28 41 4.91184 $w=1.75e-07 $l=1.70895e-07 $layer=LI1_cond $X=2.535 $Y=2.157
+ $X2=2.7 $Y2=2.145
r82 28 29 64.0104 $w=1.73e-07 $l=1.01e-06 $layer=LI1_cond $X=2.535 $Y=2.157
+ $X2=1.525 $Y2=2.157
r83 22 24 32.0379 $w=2.48e-07 $l=6.95e-07 $layer=LI1_cond $X=1.205 $Y=1.21
+ $X2=1.205 $Y2=0.515
r84 20 39 8.52281 $w=1.72e-07 $l=1.65997e-07 $layer=LI1_cond $X=1.195 $Y=2.155
+ $X2=1.36 $Y2=2.157
r85 20 21 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=1.195 $Y=2.155
+ $X2=0.785 $Y2=2.155
r86 19 32 4.974 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=0.785 $Y=1.295
+ $X2=0.61 $Y2=1.295
r87 18 22 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.08 $Y=1.295
+ $X2=1.205 $Y2=1.21
r88 18 19 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.08 $Y=1.295
+ $X2=0.785 $Y2=1.295
r89 17 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.7 $Y=2.07
+ $X2=0.785 $Y2=2.155
r90 17 37 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.7 $Y=2.07 $X2=0.7
+ $Y2=1.55
r91 13 36 75.0274 $w=2.85e-07 $l=4.18999e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.587 $Y2=1.385
r92 13 15 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.4
r93 10 36 38.666 $w=2.85e-07 $l=2.09893e-07 $layer=POLY_cond $X=0.485 $Y=1.22
+ $X2=0.587 $Y2=1.385
r94 10 12 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.485 $Y=1.22
+ $X2=0.485 $Y2=0.74
r95 3 41 300 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=2 $X=2.465
+ $Y=2.065 $X2=2.7 $Y2=2.21
r96 2 39 300 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=2 $X=1.21
+ $Y=2.065 $X2=1.36 $Y2=2.24
r97 1 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.105
+ $Y=0.37 $X2=1.245 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__O2111A_1%D1 1 3 5 6 8 11 13
c40 13 0 1.71808e-20 $X=1.2 $Y=1.665
c41 11 0 1.4602e-19 $X=1.53 $Y=1.26
c42 1 0 1.59935e-20 $X=1.135 $Y=1.99
r43 13 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.17
+ $Y=1.715 $X2=1.17 $Y2=1.715
r44 9 11 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=1.26 $Y=1.26 $X2=1.53
+ $Y2=1.26
r45 6 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.53 $Y=1.185
+ $X2=1.53 $Y2=1.26
r46 6 8 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.53 $Y=1.185
+ $X2=1.53 $Y2=0.74
r47 5 16 38.5991 $w=2.92e-07 $l=2.05122e-07 $layer=POLY_cond $X=1.26 $Y=1.55
+ $X2=1.17 $Y2=1.715
r48 4 9 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.26 $Y=1.335 $X2=1.26
+ $Y2=1.26
r49 4 5 110.245 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=1.26 $Y=1.335
+ $X2=1.26 $Y2=1.55
r50 1 16 56.7567 $w=2.92e-07 $l=2.91976e-07 $layer=POLY_cond $X=1.135 $Y=1.99
+ $X2=1.17 $Y2=1.715
r51 1 3 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.135 $Y=1.99
+ $X2=1.135 $Y2=2.485
.ends

.subckt PM_SKY130_FD_SC_LS__O2111A_1%C1 1 3 6 8 9 10 11
c38 6 0 1.41336e-19 $X=1.89 $Y=0.74
r39 11 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.71
+ $Y=1.735 $X2=1.71 $Y2=1.735
r40 10 11 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.71 $Y=1.295
+ $X2=1.71 $Y2=1.665
r41 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.71 $Y=0.925
+ $X2=1.71 $Y2=1.295
r42 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.71 $Y=0.555 $X2=1.71
+ $Y2=0.925
r43 4 17 39.0253 $w=3.68e-07 $l=2.22486e-07 $layer=POLY_cond $X=1.89 $Y=1.57
+ $X2=1.755 $Y2=1.735
r44 4 6 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=1.89 $Y=1.57 $X2=1.89
+ $Y2=0.74
r45 1 17 50.8133 $w=3.68e-07 $l=3.09233e-07 $layer=POLY_cond $X=1.635 $Y=1.99
+ $X2=1.755 $Y2=1.735
r46 1 3 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.635 $Y=1.99
+ $X2=1.635 $Y2=2.485
.ends

.subckt PM_SKY130_FD_SC_LS__O2111A_1%B1 3 6 7 9 10 13 14
c36 6 0 1.33536e-19 $X=2.39 $Y=1.9
r37 13 16 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.34 $Y=1.58
+ $X2=2.34 $Y2=1.745
r38 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.34 $Y=1.58
+ $X2=2.34 $Y2=1.415
r39 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.34
+ $Y=1.58 $X2=2.34 $Y2=1.58
r40 10 14 5.68328 $w=3.63e-07 $l=1.8e-07 $layer=LI1_cond $X=2.16 $Y=1.597
+ $X2=2.34 $Y2=1.597
r41 7 9 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.39 $Y=1.99 $X2=2.39
+ $Y2=2.485
r42 6 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.39 $Y=1.9 $X2=2.39
+ $Y2=1.99
r43 6 16 60.25 $w=1.8e-07 $l=1.55e-07 $layer=POLY_cond $X=2.39 $Y=1.9 $X2=2.39
+ $Y2=1.745
r44 3 15 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=2.28 $Y=0.74
+ $X2=2.28 $Y2=1.415
.ends

.subckt PM_SKY130_FD_SC_LS__O2111A_1%A2 3 5 7 8
c31 8 0 1.33536e-19 $X=3.12 $Y=1.665
r32 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.88
+ $Y=1.58 $X2=2.88 $Y2=1.58
r33 8 12 7.57771 $w=3.63e-07 $l=2.4e-07 $layer=LI1_cond $X=3.12 $Y=1.597
+ $X2=2.88 $Y2=1.597
r34 5 11 52.2586 $w=2.99e-07 $l=2.7157e-07 $layer=POLY_cond $X=2.925 $Y=1.83
+ $X2=2.88 $Y2=1.58
r35 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.925 $Y=1.83
+ $X2=2.925 $Y2=2.405
r36 1 11 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=2.79 $Y=1.415
+ $X2=2.88 $Y2=1.58
r37 1 3 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=2.79 $Y=1.415
+ $X2=2.79 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__O2111A_1%A1 3 5 7 8 12
r23 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.57
+ $Y=1.465 $X2=3.57 $Y2=1.465
r24 8 12 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=3.57 $Y=1.665 $X2=3.57
+ $Y2=1.465
r25 5 11 65.3342 $w=3.66e-07 $l=4.33561e-07 $layer=POLY_cond $X=3.345 $Y=1.83
+ $X2=3.495 $Y2=1.465
r26 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.345 $Y=1.83
+ $X2=3.345 $Y2=2.405
r27 1 11 38.9954 $w=3.66e-07 $l=2.33345e-07 $layer=POLY_cond $X=3.33 $Y=1.3
+ $X2=3.495 $Y2=1.465
r28 1 3 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.33 $Y=1.3 $X2=3.33
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__O2111A_1%X 1 2 9 13 14 15 16 23 32
c22 14 0 1.59935e-20 $X=0.155 $Y=1.95
r23 21 23 1.31708 $w=3.48e-07 $l=4e-08 $layer=LI1_cond $X=0.27 $Y=1.995 $X2=0.27
+ $Y2=2.035
r24 15 16 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.27 $Y=2.405
+ $X2=0.27 $Y2=2.775
r25 14 21 0.75732 $w=3.48e-07 $l=2.3e-08 $layer=LI1_cond $X=0.27 $Y=1.972
+ $X2=0.27 $Y2=1.995
r26 14 32 8.06043 $w=3.48e-07 $l=1.52e-07 $layer=LI1_cond $X=0.27 $Y=1.972
+ $X2=0.27 $Y2=1.82
r27 14 15 11.4586 $w=3.48e-07 $l=3.48e-07 $layer=LI1_cond $X=0.27 $Y=2.057
+ $X2=0.27 $Y2=2.405
r28 14 23 0.724393 $w=3.48e-07 $l=2.2e-08 $layer=LI1_cond $X=0.27 $Y=2.057
+ $X2=0.27 $Y2=2.035
r29 13 32 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=0.18 $Y=1.04
+ $X2=0.18 $Y2=1.82
r30 7 13 7.14225 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=0.225 $Y=0.91
+ $X2=0.225 $Y2=1.04
r31 7 9 17.5083 $w=2.58e-07 $l=3.95e-07 $layer=LI1_cond $X=0.225 $Y=0.91
+ $X2=0.225 $Y2=0.515
r32 2 14 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
r33 2 16 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r34 1 9 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.27 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__O2111A_1%VPWR 1 2 3 12 16 18 20 24 26 31 36 42 45 49
r48 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r49 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r50 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r51 40 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r52 40 46 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.16 $Y2=3.33
r53 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r54 37 45 11.9488 $w=1.7e-07 $l=2.75e-07 $layer=LI1_cond $X=2.29 $Y=3.33
+ $X2=2.015 $Y2=3.33
r55 37 39 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=2.29 $Y=3.33
+ $X2=3.12 $Y2=3.33
r56 36 48 4.76062 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=3.405 $Y=3.33
+ $X2=3.622 $Y2=3.33
r57 36 39 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=3.405 $Y=3.33
+ $X2=3.12 $Y2=3.33
r58 35 43 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r59 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r60 32 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=0.78 $Y2=3.33
r61 32 34 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=1.68 $Y2=3.33
r62 31 45 11.9488 $w=1.7e-07 $l=2.75e-07 $layer=LI1_cond $X=1.74 $Y=3.33
+ $X2=2.015 $Y2=3.33
r63 31 34 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=1.74 $Y=3.33 $X2=1.68
+ $Y2=3.33
r64 29 43 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r65 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r66 26 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.78 $Y2=3.33
r67 26 28 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.24 $Y2=3.33
r68 24 46 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.16 $Y2=3.33
r69 24 35 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r70 20 23 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=3.57 $Y=2.08
+ $X2=3.57 $Y2=2.76
r71 18 48 3.00555 $w=3.3e-07 $l=1.07912e-07 $layer=LI1_cond $X=3.57 $Y=3.245
+ $X2=3.622 $Y2=3.33
r72 18 23 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=3.57 $Y=3.245
+ $X2=3.57 $Y2=2.76
r73 14 45 2.31338 $w=5.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.015 $Y=3.245
+ $X2=2.015 $Y2=3.33
r74 14 16 13.5918 $w=5.48e-07 $l=6.25e-07 $layer=LI1_cond $X=2.015 $Y=3.245
+ $X2=2.015 $Y2=2.62
r75 10 42 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=3.245
+ $X2=0.78 $Y2=3.33
r76 10 12 26.1919 $w=3.28e-07 $l=7.5e-07 $layer=LI1_cond $X=0.78 $Y=3.245
+ $X2=0.78 $Y2=2.495
r77 3 23 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=3.42
+ $Y=1.905 $X2=3.57 $Y2=2.76
r78 3 20 400 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=1 $X=3.42
+ $Y=1.905 $X2=3.57 $Y2=2.08
r79 2 16 600 $w=1.7e-07 $l=6.90869e-07 $layer=licon1_PDIFF $count=1 $X=1.71
+ $Y=2.065 $X2=2.015 $Y2=2.62
r80 1 12 300 $w=1.7e-07 $l=7.48348e-07 $layer=licon1_PDIFF $count=2 $X=0.58
+ $Y=1.84 $X2=0.78 $Y2=2.495
.ends

.subckt PM_SKY130_FD_SC_LS__O2111A_1%VGND 1 2 9 13 15 17 22 32 33 36 39
r43 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r44 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r45 33 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r46 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r47 30 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.21 $Y=0 $X2=3.045
+ $Y2=0
r48 30 32 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=3.21 $Y=0 $X2=3.6
+ $Y2=0
r49 29 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r50 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r51 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r52 25 28 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r53 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r54 23 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.865 $Y=0 $X2=0.7
+ $Y2=0
r55 23 25 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.865 $Y=0 $X2=1.2
+ $Y2=0
r56 22 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.88 $Y=0 $X2=3.045
+ $Y2=0
r57 22 28 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=2.88 $Y=0 $X2=2.64
+ $Y2=0
r58 20 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r59 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r60 17 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.535 $Y=0 $X2=0.7
+ $Y2=0
r61 17 19 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.535 $Y=0 $X2=0.24
+ $Y2=0
r62 15 29 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.64
+ $Y2=0
r63 15 26 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.2
+ $Y2=0
r64 11 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.045 $Y=0.085
+ $X2=3.045 $Y2=0
r65 11 13 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=3.045 $Y=0.085
+ $X2=3.045 $Y2=0.57
r66 7 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.7 $Y=0.085 $X2=0.7
+ $Y2=0
r67 7 9 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.7 $Y=0.085 $X2=0.7
+ $Y2=0.515
r68 2 13 182 $w=1.7e-07 $l=2.75681e-07 $layer=licon1_NDIFF $count=1 $X=2.865
+ $Y=0.37 $X2=3.045 $Y2=0.57
r69 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.56
+ $Y=0.37 $X2=0.7 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__O2111A_1%A_471_74# 1 2 9 11 12 15
r26 13 15 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=3.545 $Y=0.96
+ $X2=3.545 $Y2=0.515
r27 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.38 $Y=1.045
+ $X2=3.545 $Y2=0.96
r28 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.38 $Y=1.045
+ $X2=2.71 $Y2=1.045
r29 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.545 $Y=0.96
+ $X2=2.71 $Y2=1.045
r30 7 9 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=2.545 $Y=0.96
+ $X2=2.545 $Y2=0.515
r31 2 15 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.405
+ $Y=0.37 $X2=3.545 $Y2=0.515
r32 1 9 91 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_NDIFF $count=2 $X=2.355
+ $Y=0.37 $X2=2.545 $Y2=0.515
.ends

