* File: sky130_fd_sc_ls__o41ai_4.spice
* Created: Wed Sep  2 11:23:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__o41ai_4.pex.spice"
.subckt sky130_fd_sc_ls__o41ai_4  VNB VPB B1 A4 A3 A2 A1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A1	A1
* A2	A2
* A3	A3
* A4	A4
* B1	B1
* VPB	VPB
* VNB	VNB
MM1010 N_A_27_74#_M1010_d N_B1_M1010_g N_Y_M1010_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75009.3 A=0.111 P=1.78 MULT=1
MM1012 N_A_27_74#_M1012_d N_B1_M1012_g N_Y_M1010_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75008.9 A=0.111 P=1.78 MULT=1
MM1027 N_A_27_74#_M1012_d N_B1_M1027_g N_Y_M1027_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.1
+ SB=75008.4 A=0.111 P=1.78 MULT=1
MM1028 N_A_27_74#_M1028_d N_B1_M1028_g N_Y_M1027_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1295 AS=0.1295 PD=1.09 PS=1.09 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75001.6
+ SB=75007.9 A=0.111 P=1.78 MULT=1
MM1008 N_VGND_M1008_d N_A4_M1008_g N_A_27_74#_M1028_d VNB NSHORT L=0.15 W=0.74
+ AD=0.2146 AS=0.1295 PD=1.32 PS=1.09 NRD=25.944 NRS=0 M=1 R=4.93333 SA=75002.1
+ SB=75007.4 A=0.111 P=1.78 MULT=1
MM1014 N_VGND_M1008_d N_A4_M1014_g N_A_27_74#_M1014_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2146 AS=0.11285 PD=1.32 PS=1.045 NRD=22.692 NRS=4.044 M=1 R=4.93333
+ SA=75002.8 SB=75006.7 A=0.111 P=1.78 MULT=1
MM1019 N_VGND_M1019_d N_A4_M1019_g N_A_27_74#_M1014_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.11285 PD=1.02 PS=1.045 NRD=0 NRS=0 M=1 R=4.93333 SA=75003.3
+ SB=75006.3 A=0.111 P=1.78 MULT=1
MM1036 N_VGND_M1019_d N_A4_M1036_g N_A_27_74#_M1036_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75003.7
+ SB=75005.8 A=0.111 P=1.78 MULT=1
MM1029 N_A_27_74#_M1036_s N_A3_M1029_g N_VGND_M1029_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75004.1
+ SB=75005.4 A=0.111 P=1.78 MULT=1
MM1033 N_A_27_74#_M1033_d N_A3_M1033_g N_VGND_M1029_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75004.6
+ SB=75004.9 A=0.111 P=1.78 MULT=1
MM1034 N_A_27_74#_M1033_d N_A3_M1034_g N_VGND_M1034_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75005
+ SB=75004.5 A=0.111 P=1.78 MULT=1
MM1037 N_A_27_74#_M1037_d N_A3_M1037_g N_VGND_M1034_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75005.5
+ SB=75004 A=0.111 P=1.78 MULT=1
MM1001 N_A_27_74#_M1037_d N_A2_M1001_g N_VGND_M1001_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75006
+ SB=75003.5 A=0.111 P=1.78 MULT=1
MM1013 N_A_27_74#_M1013_d N_A2_M1013_g N_VGND_M1001_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75006.5
+ SB=75003 A=0.111 P=1.78 MULT=1
MM1017 N_A_27_74#_M1013_d N_A2_M1017_g N_VGND_M1017_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.11655 PD=1.02 PS=1.055 NRD=0 NRS=0 M=1 R=4.93333 SA=75006.9
+ SB=75002.6 A=0.111 P=1.78 MULT=1
MM1024 N_A_27_74#_M1024_d N_A2_M1024_g N_VGND_M1017_s VNB NSHORT L=0.15 W=0.74
+ AD=0.12395 AS=0.11655 PD=1.075 PS=1.055 NRD=0 NRS=5.664 M=1 R=4.93333
+ SA=75007.4 SB=75002.1 A=0.111 P=1.78 MULT=1
MM1002 N_A_27_74#_M1024_d N_A1_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.74
+ AD=0.12395 AS=0.13505 PD=1.075 PS=1.105 NRD=8.916 NRS=2.424 M=1 R=4.93333
+ SA=75007.9 SB=75001.7 A=0.111 P=1.78 MULT=1
MM1004 N_A_27_74#_M1004_d N_A1_M1004_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.13505 PD=1.02 PS=1.105 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75008.4
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1030 N_A_27_74#_M1004_d N_A1_M1030_g N_VGND_M1030_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75008.8
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1031 N_A_27_74#_M1031_d N_A1_M1031_g N_VGND_M1030_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.1295 PD=2.05 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75009.3
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1018 N_VPWR_M1018_d N_B1_M1018_g N_Y_M1018_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.224 PD=2.83 PS=1.52 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75000.2 SB=75000.8 A=0.168 P=2.54 MULT=1
MM1020 N_VPWR_M1020_d N_B1_M1020_g N_Y_M1018_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.224 PD=2.83 PS=1.52 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75000.8 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1000 N_A_339_368#_M1000_d N_A4_M1000_g N_Y_M1000_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75003.5 A=0.168 P=2.54 MULT=1
MM1007 N_A_339_368#_M1007_d N_A4_M1007_g N_Y_M1000_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75003 A=0.168 P=2.54 MULT=1
MM1015 N_A_339_368#_M1007_d N_A4_M1015_g N_Y_M1015_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75002.6 A=0.168 P=2.54 MULT=1
MM1025 N_A_339_368#_M1025_d N_A4_M1025_g N_Y_M1015_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.6 SB=75002.1 A=0.168 P=2.54 MULT=1
MM1003 N_A_788_368#_M1003_d N_A3_M1003_g N_A_339_368#_M1025_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.224 AS=0.168 PD=1.52 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75002 SB=75001.7 A=0.168 P=2.54 MULT=1
MM1005 N_A_788_368#_M1003_d N_A3_M1005_g N_A_339_368#_M1005_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.224 AS=0.168 PD=1.52 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75002.6 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1022 N_A_788_368#_M1022_d N_A3_M1022_g N_A_339_368#_M1005_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75003 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1032 N_A_788_368#_M1022_d N_A3_M1032_g N_A_339_368#_M1032_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75003.5 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1009 N_A_788_368#_M1009_d N_A2_M1009_g N_A_1191_368#_M1009_s VPB PHIGHVT
+ L=0.15 W=1.12 AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1
+ R=7.46667 SA=75000.2 SB=75003.5 A=0.168 P=2.54 MULT=1
MM1016 N_A_788_368#_M1009_d N_A2_M1016_g N_A_1191_368#_M1016_s VPB PHIGHVT
+ L=0.15 W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1
+ R=7.46667 SA=75000.7 SB=75003 A=0.168 P=2.54 MULT=1
MM1023 N_A_788_368#_M1023_d N_A2_M1023_g N_A_1191_368#_M1016_s VPB PHIGHVT
+ L=0.15 W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1
+ R=7.46667 SA=75001.1 SB=75002.6 A=0.168 P=2.54 MULT=1
MM1035 N_A_788_368#_M1023_d N_A2_M1035_g N_A_1191_368#_M1035_s VPB PHIGHVT
+ L=0.15 W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1
+ R=7.46667 SA=75001.6 SB=75002.1 A=0.168 P=2.54 MULT=1
MM1006 N_VPWR_M1006_d N_A1_M1006_g N_A_1191_368#_M1035_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.196 AS=0.168 PD=1.47 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002 SB=75001.7 A=0.168 P=2.54 MULT=1
MM1011 N_VPWR_M1006_d N_A1_M1011_g N_A_1191_368#_M1011_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.196 AS=0.168 PD=1.47 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75002.5 SB=75001.2 A=0.168 P=2.54 MULT=1
MM1021 N_VPWR_M1021_d N_A1_M1021_g N_A_1191_368#_M1011_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.196 AS=0.168 PD=1.47 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75003 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1026 N_VPWR_M1021_d N_A1_M1026_g N_A_1191_368#_M1026_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.196 AS=0.3304 PD=1.47 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75003.5 SB=75000.2 A=0.168 P=2.54 MULT=1
DX38_noxref VNB VPB NWDIODE A=19.4556 P=24.64
*
.include "sky130_fd_sc_ls__o41ai_4.pxi.spice"
*
.ends
*
*
