* NGSPICE file created from sky130_fd_sc_ls__o22a_4.ext - technology: sky130A

.subckt sky130_fd_sc_ls__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
M1000 X a_206_392# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=7.112e+11p pd=5.75e+06u as=2.1626e+12p ps=1.475e+07u
M1001 a_27_136# B1 a_206_392# VNB nshort w=640000u l=150000u
+  ad=1.0112e+12p pd=9.56e+06u as=3.616e+11p ps=3.69e+06u
M1002 VGND a_206_392# X VNB nshort w=740000u l=150000u
+  ad=1.1945e+12p pd=1.055e+07u as=4.144e+11p ps=4.08e+06u
M1003 VPWR A1 a_116_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=6.5e+11p ps=5.3e+06u
M1004 VGND a_206_392# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_516_392# B1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=6.5e+11p pd=5.3e+06u as=0p ps=0u
M1006 a_206_392# B2 a_27_136# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_206_392# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR a_206_392# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 X a_206_392# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_206_392# B2 a_516_392# VPB phighvt w=1e+06u l=150000u
+  ad=7e+11p pd=5.4e+06u as=0p ps=0u
M1011 a_27_136# B2 a_206_392# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_27_136# A2 VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR a_206_392# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND A2 a_27_136# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND A1 a_27_136# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_27_136# A1 VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_206_392# A2 a_116_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_116_392# A1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_516_392# B2 a_206_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 X a_206_392# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_206_392# B1 a_27_136# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_116_392# A2 a_206_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VPWR B1 a_516_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

