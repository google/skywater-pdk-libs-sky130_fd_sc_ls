* File: sky130_fd_sc_ls__sedfxtp_4.pex.spice
* Created: Wed Sep  2 11:29:38 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__SEDFXTP_4%D 2 3 5 8 12 13 18 19 21 23
c42 23 0 2.17154e-19 $X=0.51 $Y=1.99
c43 18 0 1.43045e-19 $X=0.51 $Y=1.145
r44 21 23 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.51 $Y=1.825
+ $X2=0.51 $Y2=1.99
r45 21 22 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.51
+ $Y=1.825 $X2=0.51 $Y2=1.825
r46 18 21 118.906 $w=3.3e-07 $l=6.8e-07 $layer=POLY_cond $X=0.51 $Y=1.145
+ $X2=0.51 $Y2=1.825
r47 18 19 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.51
+ $Y=1.145 $X2=0.51 $Y2=1.145
r48 13 22 4.60977 $w=3.98e-07 $l=1.6e-07 $layer=LI1_cond $X=0.625 $Y=1.665
+ $X2=0.625 $Y2=1.825
r49 12 13 10.6601 $w=3.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.625 $Y=1.295
+ $X2=0.625 $Y2=1.665
r50 12 19 4.32166 $w=3.98e-07 $l=1.5e-07 $layer=LI1_cond $X=0.625 $Y=1.295
+ $X2=0.625 $Y2=1.145
r51 11 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.51 $Y=0.98
+ $X2=0.51 $Y2=1.145
r52 8 11 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=0.6 $Y=0.58 $X2=0.6
+ $Y2=0.98
r53 3 5 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.555 $Y=2.245
+ $X2=0.555 $Y2=2.64
r54 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.555 $Y=2.155 $X2=0.555
+ $Y2=2.245
r55 2 23 64.1371 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.555 $Y=2.155
+ $X2=0.555 $Y2=1.99
.ends

.subckt PM_SKY130_FD_SC_LS__SEDFXTP_4%A_177_290# 1 2 7 9 12 14 18 19 20 21 22 23
+ 26 30 32 34 44
c108 32 0 7.47378e-20 $X=2.24 $Y=1.95
c109 23 0 3.15633e-20 $X=1.325 $Y=2.035
c110 21 0 1.43045e-19 $X=1.325 $Y=1.065
c111 19 0 1.82239e-19 $X=1.16 $Y=1.615
r112 35 44 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=2.24 $Y=1.685
+ $X2=2.41 $Y2=1.685
r113 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.24
+ $Y=1.685 $X2=2.24 $Y2=1.685
r114 32 37 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=2.24 $Y=2.035
+ $X2=1.88 $Y2=2.035
r115 32 34 12.2159 $w=2.48e-07 $l=2.65e-07 $layer=LI1_cond $X=2.24 $Y=1.95
+ $X2=2.24 $Y2=1.685
r116 28 37 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.88 $Y=2.12
+ $X2=1.88 $Y2=2.035
r117 28 30 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.88 $Y=2.12
+ $X2=1.88 $Y2=2.515
r118 24 26 9.45003 $w=2.48e-07 $l=2.05e-07 $layer=LI1_cond $X=1.725 $Y=0.98
+ $X2=1.725 $Y2=0.775
r119 22 37 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.795 $Y=2.035
+ $X2=1.88 $Y2=2.035
r120 22 23 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=1.795 $Y=2.035
+ $X2=1.325 $Y2=2.035
r121 20 24 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.6 $Y=1.065
+ $X2=1.725 $Y2=0.98
r122 20 21 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.6 $Y=1.065
+ $X2=1.325 $Y2=1.065
r123 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.16
+ $Y=1.615 $X2=1.16 $Y2=1.615
r124 16 23 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.16 $Y=1.95
+ $X2=1.325 $Y2=2.035
r125 16 18 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.16 $Y=1.95
+ $X2=1.16 $Y2=1.615
r126 15 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.16 $Y=1.15
+ $X2=1.325 $Y2=1.065
r127 15 18 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=1.16 $Y=1.15
+ $X2=1.16 $Y2=1.615
r128 14 19 36.0236 $w=4.4e-07 $l=2.85e-07 $layer=POLY_cond $X=1.105 $Y=1.9
+ $X2=1.105 $Y2=1.615
r129 10 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.41 $Y=1.52
+ $X2=2.41 $Y2=1.685
r130 10 12 382.011 $w=1.5e-07 $l=7.45e-07 $layer=POLY_cond $X=2.41 $Y=1.52
+ $X2=2.41 $Y2=0.775
r131 7 14 48.2 $w=3.45e-07 $l=4.04815e-07 $layer=POLY_cond $X=0.975 $Y=2.245
+ $X2=1.105 $Y2=1.9
r132 7 9 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.975 $Y=2.245
+ $X2=0.975 $Y2=2.64
r133 2 30 600 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=1 $X=1.735
+ $Y=2.315 $X2=1.88 $Y2=2.515
r134 1 26 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=1.62
+ $Y=0.565 $X2=1.765 $Y2=0.775
.ends

.subckt PM_SKY130_FD_SC_LS__SEDFXTP_4%DE 3 5 6 10 11 12 13 15 16 18 19 21 23 24
+ 25 26 29 30 31
c93 31 0 7.47378e-20 $X=1.7 $Y=1.65
c94 30 0 1.36415e-19 $X=1.7 $Y=1.485
r95 29 31 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.7 $Y=1.485
+ $X2=1.7 $Y2=1.65
r96 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.7
+ $Y=1.485 $X2=1.7 $Y2=1.485
r97 26 30 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=1.7 $Y=1.665 $X2=1.7
+ $Y2=1.485
r98 21 23 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.785 $Y=2.24
+ $X2=2.785 $Y2=2.635
r99 20 25 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.18 $Y=2.165
+ $X2=2.105 $Y2=2.165
r100 19 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.71 $Y=2.165
+ $X2=2.785 $Y2=2.24
r101 19 20 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.71 $Y=2.165
+ $X2=2.18 $Y2=2.165
r102 16 25 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.105 $Y=2.24
+ $X2=2.105 $Y2=2.165
r103 16 18 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.105 $Y=2.24
+ $X2=2.105 $Y2=2.635
r104 13 24 13.5877 $w=2.4e-07 $l=2.19317e-07 $layer=POLY_cond $X=1.98 $Y=1.06
+ $X2=1.795 $Y2=1.135
r105 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.98 $Y=1.06
+ $X2=1.98 $Y2=0.775
r106 11 25 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.03 $Y=2.165
+ $X2=2.105 $Y2=2.165
r107 11 12 99.9894 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=2.03 $Y=2.165
+ $X2=1.835 $Y2=2.165
r108 10 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.76 $Y=2.09
+ $X2=1.835 $Y2=2.165
r109 10 31 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=1.76 $Y=2.09
+ $X2=1.76 $Y2=1.65
r110 7 24 13.5877 $w=2.4e-07 $l=1.27083e-07 $layer=POLY_cond $X=1.7 $Y=1.21
+ $X2=1.795 $Y2=1.135
r111 7 29 48.0869 $w=3.3e-07 $l=2.75e-07 $layer=POLY_cond $X=1.7 $Y=1.21 $X2=1.7
+ $Y2=1.485
r112 5 24 12.1617 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=1.535 $Y=1.135
+ $X2=1.795 $Y2=1.135
r113 5 6 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=1.535 $Y=1.135 $X2=1.065
+ $Y2=1.135
r114 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.99 $Y=1.06
+ $X2=1.065 $Y2=1.135
r115 1 3 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.99 $Y=1.06 $X2=0.99
+ $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_LS__SEDFXTP_4%A_545_87# 1 2 9 12 13 15 16 18 19 20 21 23
+ 25 26 30 33 35 40 42 45 47 48 49 55 56 62 63
c241 55 0 1.04115e-19 $X=14.64 $Y=1.665
c242 48 0 5.67286e-20 $X=14.495 $Y=1.665
c243 25 0 5.64986e-20 $X=13.41 $Y=2.05
c244 13 0 1.85697e-19 $X=3.175 $Y=2.24
r245 61 63 49.8355 $w=3.3e-07 $l=2.85e-07 $layer=POLY_cond $X=2.89 $Y=1.685
+ $X2=3.175 $Y2=1.685
r246 61 62 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.89
+ $Y=1.685 $X2=2.89 $Y2=1.685
r247 58 61 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.8 $Y=1.685 $X2=2.89
+ $Y2=1.685
r248 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.64 $Y=1.665
+ $X2=14.64 $Y2=1.665
r249 52 62 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=2.64 $Y=1.685
+ $X2=2.89 $Y2=1.685
r250 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=1.665
+ $X2=2.64 $Y2=1.665
r251 49 51 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.785 $Y=1.665
+ $X2=2.64 $Y2=1.665
r252 48 55 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=14.495 $Y=1.665
+ $X2=14.64 $Y2=1.665
r253 48 49 14.4925 $w=1.4e-07 $l=1.171e-05 $layer=MET1_cond $X=14.495 $Y=1.665
+ $X2=2.785 $Y2=1.665
r254 46 56 12.276 $w=2.28e-07 $l=2.45e-07 $layer=LI1_cond $X=14.395 $Y=1.665
+ $X2=14.64 $Y2=1.665
r255 46 47 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=14.395 $Y=1.665
+ $X2=14.31 $Y2=1.665
r256 42 44 10.5284 $w=3.88e-07 $l=2.3e-07 $layer=LI1_cond $X=14.2 $Y=0.58
+ $X2=14.2 $Y2=0.81
r257 37 40 8.74048 $w=2.53e-07 $l=1.65e-07 $layer=LI1_cond $X=13.32 $Y=2.222
+ $X2=13.485 $Y2=2.222
r258 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.32
+ $Y=2.215 $X2=13.32 $Y2=2.215
r259 35 45 3.58051 $w=2.6e-07 $l=1.25499e-07 $layer=LI1_cond $X=14.31 $Y=2.18
+ $X2=14.22 $Y2=2.265
r260 34 47 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=14.31 $Y=1.78
+ $X2=14.31 $Y2=1.665
r261 34 35 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=14.31 $Y=1.78
+ $X2=14.31 $Y2=2.18
r262 33 47 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=14.31 $Y=1.55
+ $X2=14.31 $Y2=1.665
r263 33 44 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=14.31 $Y=1.55
+ $X2=14.31 $Y2=0.81
r264 28 45 3.58051 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=14.22 $Y=2.35
+ $X2=14.22 $Y2=2.265
r265 28 30 3.7866 $w=3.48e-07 $l=1.15e-07 $layer=LI1_cond $X=14.22 $Y=2.35
+ $X2=14.22 $Y2=2.465
r266 26 45 2.90867 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=14.045 $Y=2.265
+ $X2=14.22 $Y2=2.265
r267 26 40 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=14.045 $Y=2.265
+ $X2=13.485 $Y2=2.265
r268 25 38 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=13.41 $Y=2.05
+ $X2=13.32 $Y2=2.215
r269 24 25 530.713 $w=1.5e-07 $l=1.035e-06 $layer=POLY_cond $X=13.41 $Y=1.015
+ $X2=13.41 $Y2=2.05
r270 21 38 52.2586 $w=2.99e-07 $l=2.7157e-07 $layer=POLY_cond $X=13.275 $Y=2.465
+ $X2=13.32 $Y2=2.215
r271 21 23 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=13.275 $Y=2.465
+ $X2=13.275 $Y2=2.75
r272 19 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=13.335 $Y=0.94
+ $X2=13.41 $Y2=1.015
r273 19 20 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=13.335 $Y=0.94
+ $X2=12.88 $Y2=0.94
r274 16 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=12.805 $Y=0.865
+ $X2=12.88 $Y2=0.94
r275 16 18 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=12.805 $Y=0.865
+ $X2=12.805 $Y2=0.58
r276 13 15 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.175 $Y=2.24
+ $X2=3.175 $Y2=2.635
r277 12 13 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.175 $Y=2.15
+ $X2=3.175 $Y2=2.24
r278 11 63 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.175 $Y=1.85
+ $X2=3.175 $Y2=1.685
r279 11 12 116.613 $w=1.8e-07 $l=3e-07 $layer=POLY_cond $X=3.175 $Y=1.85
+ $X2=3.175 $Y2=2.15
r280 7 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.8 $Y=1.52 $X2=2.8
+ $Y2=1.685
r281 7 9 382.011 $w=1.5e-07 $l=7.45e-07 $layer=POLY_cond $X=2.8 $Y=1.52 $X2=2.8
+ $Y2=0.775
r282 2 30 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=14.06
+ $Y=2.32 $X2=14.21 $Y2=2.465
r283 1 42 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=14.03
+ $Y=0.37 $X2=14.17 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_LS__SEDFXTP_4%A_631_87# 1 2 7 9 10 11 12 14 17 18 21 22
+ 27 28 30 31 35 36 41 43 47
r115 44 47 4.60989 $w=4.78e-07 $l=1.85e-07 $layer=LI1_cond $X=4.19 $Y=2.495
+ $X2=4.375 $Y2=2.495
r116 35 36 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.745
+ $Y=1.58 $X2=5.745 $Y2=1.58
r117 33 35 13.7882 $w=2.78e-07 $l=3.35e-07 $layer=LI1_cond $X=5.72 $Y=1.915
+ $X2=5.72 $Y2=1.58
r118 32 43 2.36881 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=4.275 $Y=2 $X2=4.135
+ $Y2=2
r119 31 33 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=5.58 $Y=2
+ $X2=5.72 $Y2=1.915
r120 31 32 85.139 $w=1.68e-07 $l=1.305e-06 $layer=LI1_cond $X=5.58 $Y=2
+ $X2=4.275 $Y2=2
r121 30 44 6.90116 $w=1.7e-07 $l=2.4e-07 $layer=LI1_cond $X=4.19 $Y=2.255
+ $X2=4.19 $Y2=2.495
r122 29 43 4.06715 $w=2.25e-07 $l=1.09087e-07 $layer=LI1_cond $X=4.19 $Y=2.085
+ $X2=4.135 $Y2=2
r123 29 30 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.19 $Y=2.085
+ $X2=4.19 $Y2=2.255
r124 27 28 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=4.08
+ $Y=1.78 $X2=4.08 $Y2=1.78
r125 25 43 4.06715 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=4.135 $Y=1.915
+ $X2=4.135 $Y2=2
r126 25 27 5.55642 $w=2.78e-07 $l=1.35e-07 $layer=LI1_cond $X=4.135 $Y=1.915
+ $X2=4.135 $Y2=1.78
r127 24 27 31.6922 $w=2.78e-07 $l=7.7e-07 $layer=LI1_cond $X=4.135 $Y=1.01
+ $X2=4.135 $Y2=1.78
r128 21 22 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=4.08
+ $Y=0.42 $X2=4.08 $Y2=0.42
r129 19 41 10.3862 $w=4.03e-07 $l=3.65e-07 $layer=LI1_cond $X=4.135 $Y=0.807
+ $X2=4.5 $Y2=0.807
r130 19 24 2.89865 $w=2.8e-07 $l=2.03e-07 $layer=LI1_cond $X=4.135 $Y=0.807
+ $X2=4.135 $Y2=1.01
r131 19 21 7.61436 $w=2.78e-07 $l=1.85e-07 $layer=LI1_cond $X=4.135 $Y=0.605
+ $X2=4.135 $Y2=0.42
r132 18 36 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=5.745 $Y=1.92
+ $X2=5.745 $Y2=1.58
r133 16 28 99.6709 $w=3.3e-07 $l=5.7e-07 $layer=POLY_cond $X=4.08 $Y=1.21
+ $X2=4.08 $Y2=1.78
r134 16 17 10.1687 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.08 $Y=1.21
+ $X2=4.08 $Y2=1.135
r135 15 22 111.911 $w=3.3e-07 $l=6.4e-07 $layer=POLY_cond $X=4.08 $Y=1.06
+ $X2=4.08 $Y2=0.42
r136 15 17 10.1687 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.08 $Y=1.06
+ $X2=4.08 $Y2=1.135
r137 12 18 50.3582 $w=2.68e-07 $l=3.15278e-07 $layer=POLY_cond $X=5.67 $Y=2.2
+ $X2=5.745 $Y2=1.92
r138 12 14 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=5.67 $Y=2.2
+ $X2=5.67 $Y2=2.595
r139 10 17 16.9349 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.915 $Y=1.135
+ $X2=4.08 $Y2=1.135
r140 10 11 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.915 $Y=1.135
+ $X2=3.305 $Y2=1.135
r141 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.23 $Y=1.06
+ $X2=3.305 $Y2=1.135
r142 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.23 $Y=1.06 $X2=3.23
+ $Y2=0.775
r143 2 47 600 $w=1.7e-07 $l=2.77489e-07 $layer=licon1_PDIFF $count=1 $X=4.245
+ $Y=2.275 $X2=4.375 $Y2=2.495
r144 1 41 182 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_NDIFF $count=1 $X=4.355
+ $Y=0.625 $X2=4.5 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LS__SEDFXTP_4%SCD 3 6 7 9 10 13
c46 13 0 1.01011e-19 $X=5.205 $Y=1.58
r47 13 16 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.205 $Y=1.58
+ $X2=5.205 $Y2=1.745
r48 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.205 $Y=1.58
+ $X2=5.205 $Y2=1.415
r49 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.205
+ $Y=1.58 $X2=5.205 $Y2=1.58
r50 10 14 7.91437 $w=4.13e-07 $l=2.85e-07 $layer=LI1_cond $X=5.162 $Y=1.295
+ $X2=5.162 $Y2=1.58
r51 7 9 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=5.28 $Y=2.2 $X2=5.28
+ $Y2=2.595
r52 6 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.28 $Y=2.11 $X2=5.28
+ $Y2=2.2
r53 6 16 141.879 $w=1.8e-07 $l=3.65e-07 $layer=POLY_cond $X=5.28 $Y=2.11
+ $X2=5.28 $Y2=1.745
r54 3 15 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=5.145 $Y=0.835
+ $X2=5.145 $Y2=1.415
.ends

.subckt PM_SKY130_FD_SC_LS__SEDFXTP_4%SCE 1 3 4 5 7 8 11 15 16 17 20 22 25
c88 22 0 1.01011e-19 $X=4.56 $Y=1.295
r89 25 28 40.6969 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=4.622 $Y=1.345
+ $X2=4.622 $Y2=1.51
r90 25 27 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=4.622 $Y=1.345
+ $X2=4.622 $Y2=1.18
r91 22 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.62
+ $Y=1.345 $X2=4.62 $Y2=1.345
r92 18 20 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=5.505 $Y=0.255
+ $X2=5.505 $Y2=0.835
r93 16 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.43 $Y=0.18
+ $X2=5.505 $Y2=0.255
r94 16 17 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=5.43 $Y=0.18 $X2=4.79
+ $Y2=0.18
r95 15 27 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=4.715 $Y=0.835
+ $X2=4.715 $Y2=1.18
r96 12 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.715 $Y=0.255
+ $X2=4.79 $Y2=0.18
r97 12 15 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=4.715 $Y=0.255
+ $X2=4.715 $Y2=0.835
r98 9 11 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=4.6 $Y=2.99 $X2=4.6
+ $Y2=2.595
r99 8 11 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=4.6 $Y=2.2 $X2=4.6
+ $Y2=2.595
r100 7 8 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=4.6 $Y=2.11 $X2=4.6
+ $Y2=2.2
r101 7 28 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=4.6 $Y=2.11 $X2=4.6
+ $Y2=1.51
r102 4 9 26.9307 $w=1.5e-07 $l=1.53542e-07 $layer=POLY_cond $X=4.51 $Y=3.105
+ $X2=4.6 $Y2=2.99
r103 4 5 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=4.51 $Y=3.105 $X2=3.7
+ $Y2=3.105
r104 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.625 $Y=3.03
+ $X2=3.7 $Y2=3.105
r105 1 3 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.625 $Y=3.03
+ $X2=3.625 $Y2=2.635
.ends

.subckt PM_SKY130_FD_SC_LS__SEDFXTP_4%CLK 1 3 4 6 7
r35 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.58
+ $Y=1.385 $X2=6.58 $Y2=1.385
r36 7 11 11.8359 $w=3.68e-07 $l=3.8e-07 $layer=LI1_cond $X=6.96 $Y=1.365
+ $X2=6.58 $Y2=1.365
r37 4 10 70.0964 $w=2.77e-07 $l=3.78385e-07 $layer=POLY_cond $X=6.65 $Y=1.73
+ $X2=6.58 $Y2=1.385
r38 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.65 $Y=1.73 $X2=6.65
+ $Y2=2.365
r39 1 10 38.7751 $w=2.77e-07 $l=2.05122e-07 $layer=POLY_cond $X=6.49 $Y=1.22
+ $X2=6.58 $Y2=1.385
r40 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=6.49 $Y=1.22 $X2=6.49
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__SEDFXTP_4%A_1510_74# 1 2 7 9 10 12 15 18 19 21 24 26
+ 27 28 33 34 37 38 41 42 43 45 46 47 49 52 53 55 57 58 61 62 65 67 68 72
c227 72 0 2.65373e-20 $X=12.93 $Y=1.42
c228 65 0 1.91272e-19 $X=9.34 $Y=1.09
c229 62 0 6.82068e-20 $X=9.34 $Y=0.945
c230 61 0 1.60056e-19 $X=8.675 $Y=2.17
c231 33 0 1.55586e-19 $X=8.58 $Y=1.82
c232 19 0 1.1504e-19 $X=12.855 $Y=2.465
r233 72 85 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=12.93 $Y=1.42
+ $X2=12.93 $Y2=1.585
r234 71 72 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.93
+ $Y=1.42 $X2=12.93 $Y2=1.42
r235 68 71 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=12.93 $Y=1.275
+ $X2=12.93 $Y2=1.42
r236 65 76 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=9.34 $Y=1.09
+ $X2=9.215 $Y2=1.09
r237 64 65 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.34
+ $Y=1.09 $X2=9.34 $Y2=1.09
r238 62 64 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=9.34 $Y=0.945
+ $X2=9.34 $Y2=1.09
r239 61 75 47.3967 $w=3e-07 $l=2.95e-07 $layer=POLY_cond $X=8.675 $Y=2.235
+ $X2=8.97 $Y2=2.235
r240 60 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.675
+ $Y=2.17 $X2=8.675 $Y2=2.17
r241 58 60 2.70794 $w=4.28e-07 $l=9.5e-08 $layer=LI1_cond $X=8.58 $Y=2.077
+ $X2=8.675 $Y2=2.077
r242 56 67 2.28545 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=11.955 $Y=1.275
+ $X2=11.82 $Y2=1.275
r243 55 68 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.765 $Y=1.275
+ $X2=12.93 $Y2=1.275
r244 55 56 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=12.765 $Y=1.275
+ $X2=11.955 $Y2=1.275
r245 53 81 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=11.85 $Y=1.635
+ $X2=11.85 $Y2=1.47
r246 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.85
+ $Y=1.635 $X2=11.85 $Y2=1.635
r247 50 67 4.14756 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=11.82 $Y=1.36
+ $X2=11.82 $Y2=1.275
r248 50 52 11.7378 $w=2.68e-07 $l=2.75e-07 $layer=LI1_cond $X=11.82 $Y=1.36
+ $X2=11.82 $Y2=1.635
r249 49 67 4.14756 $w=2.2e-07 $l=1.07121e-07 $layer=LI1_cond $X=11.77 $Y=1.19
+ $X2=11.82 $Y2=1.275
r250 48 49 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=11.77 $Y=1.03
+ $X2=11.77 $Y2=1.19
r251 46 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.685 $Y=0.945
+ $X2=11.77 $Y2=1.03
r252 46 47 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=11.685 $Y=0.945
+ $X2=11.11 $Y2=0.945
r253 45 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.025 $Y=0.86
+ $X2=11.11 $Y2=0.945
r254 44 45 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=11.025 $Y=0.425
+ $X2=11.025 $Y2=0.86
r255 42 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.94 $Y=0.34
+ $X2=11.025 $Y2=0.425
r256 42 43 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=10.94 $Y=0.34
+ $X2=10.43 $Y2=0.34
r257 40 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.345 $Y=0.425
+ $X2=10.43 $Y2=0.34
r258 40 41 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=10.345 $Y=0.425
+ $X2=10.345 $Y2=0.86
r259 39 62 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.505 $Y=0.945
+ $X2=9.34 $Y2=0.945
r260 38 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.26 $Y=0.945
+ $X2=10.345 $Y2=0.86
r261 38 39 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=10.26 $Y=0.945
+ $X2=9.505 $Y2=0.945
r262 37 62 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=9.34 $Y=0.86
+ $X2=9.34 $Y2=0.945
r263 36 37 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=9.34 $Y=0.425
+ $X2=9.34 $Y2=0.86
r264 35 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.665 $Y=0.34
+ $X2=8.58 $Y2=0.34
r265 34 36 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.175 $Y=0.34
+ $X2=9.34 $Y2=0.425
r266 34 35 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=9.175 $Y=0.34
+ $X2=8.665 $Y2=0.34
r267 33 58 6.19161 $w=1.7e-07 $l=2.57e-07 $layer=LI1_cond $X=8.58 $Y=1.82
+ $X2=8.58 $Y2=2.077
r268 32 57 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.58 $Y=0.425
+ $X2=8.58 $Y2=0.34
r269 32 33 91.0107 $w=1.68e-07 $l=1.395e-06 $layer=LI1_cond $X=8.58 $Y=0.425
+ $X2=8.58 $Y2=1.82
r270 28 58 2.91725 $w=4.28e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.495 $Y=1.992
+ $X2=8.58 $Y2=2.077
r271 28 30 9.01912 $w=3.43e-07 $l=2.7e-07 $layer=LI1_cond $X=8.495 $Y=1.992
+ $X2=8.225 $Y2=1.992
r272 26 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.495 $Y=0.34
+ $X2=8.58 $Y2=0.34
r273 26 27 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=8.495 $Y=0.34
+ $X2=7.855 $Y2=0.34
r274 22 27 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=7.73 $Y=0.425
+ $X2=7.855 $Y2=0.34
r275 22 24 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=7.73 $Y=0.425
+ $X2=7.73 $Y2=0.515
r276 19 21 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=12.855 $Y=2.465
+ $X2=12.855 $Y2=2.75
r277 18 19 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=12.855 $Y=2.375
+ $X2=12.855 $Y2=2.465
r278 18 85 307.081 $w=1.8e-07 $l=7.9e-07 $layer=POLY_cond $X=12.855 $Y=2.375
+ $X2=12.855 $Y2=1.585
r279 15 81 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=11.94 $Y=0.69
+ $X2=11.94 $Y2=1.47
r280 10 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.215 $Y=0.925
+ $X2=9.215 $Y2=1.09
r281 10 12 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=9.215 $Y=0.925
+ $X2=9.215 $Y2=0.605
r282 7 75 18.9685 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=8.97 $Y=2.465
+ $X2=8.97 $Y2=2.235
r283 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=8.97 $Y=2.465 $X2=8.97
+ $Y2=2.75
r284 2 30 600 $w=1.7e-07 $l=2.12132e-07 $layer=licon1_PDIFF $count=1 $X=8.075
+ $Y=1.84 $X2=8.225 $Y2=1.99
r285 1 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.55
+ $Y=0.37 $X2=7.69 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__SEDFXTP_4%A_1313_74# 1 2 9 11 13 15 16 20 22 25 26
+ 28 29 31 34 36 37 40 42 46 47 49 50 53 58 64 67
c191 58 0 1.29864e-19 $X=9.435 $Y=2.165
c192 50 0 1.1504e-19 $X=12.125 $Y=2.475
c193 25 0 1.55586e-19 $X=9.345 $Y=2
r194 67 68 32.6217 $w=3.9e-07 $l=7.5e-08 $layer=POLY_cond $X=7.355 $Y=1.69
+ $X2=7.355 $Y2=1.615
r195 64 65 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.39
+ $Y=1.635 $X2=12.39 $Y2=1.635
r196 61 64 9.21954 $w=2.23e-07 $l=1.8e-07 $layer=LI1_cond $X=12.21 $Y=1.642
+ $X2=12.39 $Y2=1.642
r197 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.435
+ $Y=2.165 $X2=9.435 $Y2=2.165
r198 56 67 37.0769 $w=3.9e-07 $l=2.6e-07 $layer=POLY_cond $X=7.355 $Y=1.95
+ $X2=7.355 $Y2=1.69
r199 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.325
+ $Y=1.95 $X2=7.325 $Y2=1.95
r200 52 61 2.38091 $w=1.7e-07 $l=1.13e-07 $layer=LI1_cond $X=12.21 $Y=1.755
+ $X2=12.21 $Y2=1.642
r201 52 53 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=12.21 $Y=1.755
+ $X2=12.21 $Y2=2.39
r202 51 58 13.4591 $w=2.81e-07 $l=3.89743e-07 $layer=LI1_cond $X=9.7 $Y=2.475
+ $X2=9.52 $Y2=2.165
r203 50 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=12.125 $Y=2.475
+ $X2=12.21 $Y2=2.39
r204 50 51 158.209 $w=1.68e-07 $l=2.425e-06 $layer=LI1_cond $X=12.125 $Y=2.475
+ $X2=9.7 $Y2=2.475
r205 49 55 5.33137 $w=1.7e-07 $l=2.07678e-07 $layer=LI1_cond $X=7.33 $Y=1.785
+ $X2=7.367 $Y2=1.975
r206 48 49 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=7.33 $Y=1.01
+ $X2=7.33 $Y2=1.785
r207 46 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.245 $Y=0.925
+ $X2=7.33 $Y2=1.01
r208 46 47 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=7.245 $Y=0.925
+ $X2=6.87 $Y2=0.925
r209 42 55 2.86532 $w=3.8e-07 $l=1.22e-07 $layer=LI1_cond $X=7.245 $Y=1.975
+ $X2=7.367 $Y2=1.975
r210 42 44 11.2212 $w=3.78e-07 $l=3.7e-07 $layer=LI1_cond $X=7.245 $Y=1.975
+ $X2=6.875 $Y2=1.975
r211 38 47 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.705 $Y=0.84
+ $X2=6.87 $Y2=0.925
r212 38 40 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=6.705 $Y=0.84
+ $X2=6.705 $Y2=0.515
r213 32 65 38.5562 $w=2.99e-07 $l=1.77059e-07 $layer=POLY_cond $X=12.415 $Y=1.47
+ $X2=12.39 $Y2=1.635
r214 32 34 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=12.415 $Y=1.47
+ $X2=12.415 $Y2=0.58
r215 29 65 52.2586 $w=2.99e-07 $l=2.7157e-07 $layer=POLY_cond $X=12.345 $Y=1.885
+ $X2=12.39 $Y2=1.635
r216 29 31 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=12.345 $Y=1.885
+ $X2=12.345 $Y2=2.46
r217 26 59 61.4066 $w=2.86e-07 $l=3.07409e-07 $layer=POLY_cond $X=9.42 $Y=2.465
+ $X2=9.435 $Y2=2.165
r218 26 28 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=9.42 $Y=2.465
+ $X2=9.42 $Y2=2.75
r219 25 59 38.6549 $w=2.86e-07 $l=2.05122e-07 $layer=POLY_cond $X=9.345 $Y=2
+ $X2=9.435 $Y2=2.165
r220 24 25 120.5 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=9.345 $Y=1.765
+ $X2=9.345 $Y2=2
r221 23 37 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.78 $Y=1.69
+ $X2=8.705 $Y2=1.69
r222 22 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.27 $Y=1.69
+ $X2=9.345 $Y2=1.765
r223 22 23 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=9.27 $Y=1.69
+ $X2=8.78 $Y2=1.69
r224 18 37 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.705 $Y=1.615
+ $X2=8.705 $Y2=1.69
r225 18 20 471.745 $w=1.5e-07 $l=9.2e-07 $layer=POLY_cond $X=8.705 $Y=1.615
+ $X2=8.705 $Y2=0.695
r226 17 36 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.075 $Y=1.69 $X2=8
+ $Y2=1.69
r227 16 37 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.63 $Y=1.69
+ $X2=8.705 $Y2=1.69
r228 16 17 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=8.63 $Y=1.69
+ $X2=8.075 $Y2=1.69
r229 13 36 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8 $Y=1.765 $X2=8
+ $Y2=1.69
r230 13 15 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8 $Y=1.765 $X2=8
+ $Y2=2.4
r231 12 67 25.2441 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=7.55 $Y=1.69
+ $X2=7.355 $Y2=1.69
r232 11 36 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.925 $Y=1.69 $X2=8
+ $Y2=1.69
r233 11 12 192.287 $w=1.5e-07 $l=3.75e-07 $layer=POLY_cond $X=7.925 $Y=1.69
+ $X2=7.55 $Y2=1.69
r234 9 68 448.67 $w=1.5e-07 $l=8.75e-07 $layer=POLY_cond $X=7.475 $Y=0.74
+ $X2=7.475 $Y2=1.615
r235 2 44 600 $w=1.7e-07 $l=2.33238e-07 $layer=licon1_PDIFF $count=1 $X=6.725
+ $Y=1.805 $X2=6.875 $Y2=1.975
r236 1 40 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.565
+ $Y=0.37 $X2=6.705 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__SEDFXTP_4%A_1943_53# 1 2 9 12 13 15 17 18 20 21 23
+ 24 26 32 35 36 38 43 45 52
c106 45 0 1.91272e-19 $X=10.045 $Y=1.302
c107 43 0 6.82068e-20 $X=9.88 $Y=1.315
r108 46 47 7.47431 $w=2.53e-07 $l=1.55e-07 $layer=LI1_cond $X=10.685 $Y=1.365
+ $X2=10.84 $Y2=1.365
r109 43 50 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.88 $Y=1.315
+ $X2=9.88 $Y2=1.48
r110 43 49 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.88 $Y=1.315
+ $X2=9.88 $Y2=1.15
r111 42 45 9.2829 $w=2.03e-07 $l=1.65e-07 $layer=LI1_cond $X=9.88 $Y=1.302
+ $X2=10.045 $Y2=1.302
r112 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.88
+ $Y=1.315 $X2=9.88 $Y2=1.315
r113 39 52 11.1574 $w=3.24e-07 $l=7.5e-08 $layer=POLY_cond $X=11.31 $Y=1.32
+ $X2=11.385 $Y2=1.32
r114 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.31
+ $Y=1.365 $X2=11.31 $Y2=1.365
r115 36 47 3.83738 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.925 $Y=1.365
+ $X2=10.84 $Y2=1.365
r116 36 38 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=10.925 $Y=1.365
+ $X2=11.31 $Y2=1.365
r117 34 47 3.06467 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.84 $Y=1.53
+ $X2=10.84 $Y2=1.365
r118 34 35 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=10.84 $Y=1.53
+ $X2=10.84 $Y2=1.97
r119 30 46 3.06467 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.685 $Y=1.2
+ $X2=10.685 $Y2=1.365
r120 30 32 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=10.685 $Y=1.2
+ $X2=10.685 $Y2=0.825
r121 26 35 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=10.755 $Y=2.095
+ $X2=10.84 $Y2=1.97
r122 26 28 5.30124 $w=2.48e-07 $l=1.15e-07 $layer=LI1_cond $X=10.755 $Y=2.095
+ $X2=10.64 $Y2=2.095
r123 24 46 5.41671 $w=2.53e-07 $l=1.18427e-07 $layer=LI1_cond $X=10.6 $Y=1.285
+ $X2=10.685 $Y2=1.365
r124 24 45 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=10.6 $Y=1.285
+ $X2=10.045 $Y2=1.285
r125 21 52 29.0093 $w=3.24e-07 $l=2.91633e-07 $layer=POLY_cond $X=11.58 $Y=1.11
+ $X2=11.385 $Y2=1.32
r126 21 23 134.96 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=11.58 $Y=1.11
+ $X2=11.58 $Y2=0.69
r127 18 20 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=11.385 $Y=1.885
+ $X2=11.385 $Y2=2.46
r128 17 18 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=11.385 $Y=1.795
+ $X2=11.385 $Y2=1.885
r129 16 52 16.5046 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=11.385 $Y=1.53
+ $X2=11.385 $Y2=1.32
r130 16 17 103.008 $w=1.8e-07 $l=2.65e-07 $layer=POLY_cond $X=11.385 $Y=1.53
+ $X2=11.385 $Y2=1.795
r131 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=9.9 $Y=2.465 $X2=9.9
+ $Y2=2.75
r132 12 13 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=9.9 $Y=2.375 $X2=9.9
+ $Y2=2.465
r133 12 50 347.895 $w=1.8e-07 $l=8.95e-07 $layer=POLY_cond $X=9.9 $Y=2.375
+ $X2=9.9 $Y2=1.48
r134 9 49 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=9.79 $Y=0.605
+ $X2=9.79 $Y2=1.15
r135 2 28 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=10.49
+ $Y=1.99 $X2=10.64 $Y2=2.135
r136 1 32 182 $w=1.7e-07 $l=4.95076e-07 $layer=licon1_NDIFF $count=1 $X=10.545
+ $Y=0.395 $X2=10.685 $Y2=0.825
.ends

.subckt PM_SKY130_FD_SC_LS__SEDFXTP_4%A_1756_97# 1 2 7 9 12 16 21 26 27 30 32
r88 30 32 8.69362 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=10.42 $Y=1.67
+ $X2=10.255 $Y2=1.67
r89 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.42
+ $Y=1.655 $X2=10.42 $Y2=1.655
r90 26 27 10.5918 $w=3.58e-07 $l=2.3e-07 $layer=LI1_cond $X=9.18 $Y=2.75
+ $X2=9.18 $Y2=2.52
r91 22 24 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=8.92 $Y=1.715
+ $X2=9.085 $Y2=1.715
r92 21 24 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=9.17 $Y=1.715
+ $X2=9.085 $Y2=1.715
r93 21 32 70.7861 $w=1.68e-07 $l=1.085e-06 $layer=LI1_cond $X=9.17 $Y=1.715
+ $X2=10.255 $Y2=1.715
r94 18 24 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.085 $Y=1.8
+ $X2=9.085 $Y2=1.715
r95 18 27 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=9.085 $Y=1.8
+ $X2=9.085 $Y2=2.52
r96 14 22 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.92 $Y=1.63
+ $X2=8.92 $Y2=1.715
r97 14 16 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=8.92 $Y=1.63
+ $X2=8.92 $Y2=0.76
r98 10 31 38.5718 $w=2.96e-07 $l=1.88348e-07 $layer=POLY_cond $X=10.47 $Y=1.49
+ $X2=10.42 $Y2=1.655
r99 10 12 397.394 $w=1.5e-07 $l=7.75e-07 $layer=POLY_cond $X=10.47 $Y=1.49
+ $X2=10.47 $Y2=0.715
r100 7 31 54.0414 $w=2.96e-07 $l=2.62488e-07 $layer=POLY_cond $X=10.415 $Y=1.915
+ $X2=10.42 $Y2=1.655
r101 7 9 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=10.415 $Y=1.915
+ $X2=10.415 $Y2=2.41
r102 2 26 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=9.045
+ $Y=2.54 $X2=9.195 $Y2=2.75
r103 1 16 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=8.78
+ $Y=0.485 $X2=8.92 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_LS__SEDFXTP_4%A_2403_74# 1 2 8 11 14 15 17 18 20 22 23
+ 25 26 28 29 31 32 34 35 37 38 40 41 43 50 54 56 57 60 62 63 65 67 68 75
c185 65 0 1.04115e-19 $X=13.66 $Y=1.755
c186 56 0 5.64986e-20 $X=13.265 $Y=0.935
r187 72 77 40.7727 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=13.9 $Y=1.825
+ $X2=13.9 $Y2=1.99
r188 72 75 47.4823 $w=3.5e-07 $l=2.88e-07 $layer=POLY_cond $X=13.9 $Y=1.825
+ $X2=13.9 $Y2=1.537
r189 71 72 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=13.89
+ $Y=1.825 $X2=13.89 $Y2=1.825
r190 68 74 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=13.9 $Y=1.145
+ $X2=13.9 $Y2=0.98
r191 67 68 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=13.89
+ $Y=1.145 $X2=13.89 $Y2=1.145
r192 65 71 2.45986 $w=7.9e-07 $l=1.17e-07 $layer=LI1_cond $X=13.66 $Y=1.755
+ $X2=13.66 $Y2=1.872
r193 65 67 9.23554 $w=7.88e-07 $l=6.1e-07 $layer=LI1_cond $X=13.66 $Y=1.755
+ $X2=13.66 $Y2=1.145
r194 64 67 1.89253 $w=7.88e-07 $l=1.25e-07 $layer=LI1_cond $X=13.66 $Y=1.02
+ $X2=13.66 $Y2=1.145
r195 62 71 8.97743 $w=1.7e-07 $l=4.10688e-07 $layer=LI1_cond $X=13.265 $Y=1.84
+ $X2=13.66 $Y2=1.872
r196 62 63 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=13.265 $Y=1.84
+ $X2=12.895 $Y2=1.84
r197 58 63 11.2112 $w=2.82e-07 $l=2.63116e-07 $layer=LI1_cond $X=12.68 $Y=1.947
+ $X2=12.895 $Y2=1.84
r198 58 60 16.3486 $w=4.28e-07 $l=6.1e-07 $layer=LI1_cond $X=12.68 $Y=2.14
+ $X2=12.68 $Y2=2.75
r199 56 64 140.512 $w=3.9e-08 $l=4.35431e-07 $layer=LI1_cond $X=13.265 $Y=0.935
+ $X2=13.66 $Y2=1.02
r200 56 57 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=13.265 $Y=0.935
+ $X2=12.365 $Y2=0.935
r201 52 57 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=12.2 $Y=0.85
+ $X2=12.365 $Y2=0.935
r202 52 54 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=12.2 $Y=0.85
+ $X2=12.2 $Y2=0.58
r203 50 51 2.22462 $w=3.25e-07 $l=1.5e-08 $layer=POLY_cond $X=16.305 $Y=1.58
+ $X2=16.32 $Y2=1.58
r204 49 50 63.7723 $w=3.25e-07 $l=4.3e-07 $layer=POLY_cond $X=15.875 $Y=1.58
+ $X2=16.305 $Y2=1.58
r205 48 49 2.96615 $w=3.25e-07 $l=2e-08 $layer=POLY_cond $X=15.855 $Y=1.58
+ $X2=15.875 $Y2=1.58
r206 47 48 66.7385 $w=3.25e-07 $l=4.5e-07 $layer=POLY_cond $X=15.405 $Y=1.58
+ $X2=15.855 $Y2=1.58
r207 46 47 4.44923 $w=3.25e-07 $l=3e-08 $layer=POLY_cond $X=15.375 $Y=1.58
+ $X2=15.405 $Y2=1.58
r208 45 46 62.2892 $w=3.25e-07 $l=4.2e-07 $layer=POLY_cond $X=14.955 $Y=1.58
+ $X2=15.375 $Y2=1.58
r209 44 45 1.48308 $w=3.25e-07 $l=1e-08 $layer=POLY_cond $X=14.945 $Y=1.58
+ $X2=14.955 $Y2=1.58
r210 41 51 20.86 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=16.32 $Y=1.395
+ $X2=16.32 $Y2=1.58
r211 41 43 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=16.32 $Y=1.395
+ $X2=16.32 $Y2=0.95
r212 38 50 20.86 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=16.305 $Y=1.765
+ $X2=16.305 $Y2=1.58
r213 38 40 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=16.305 $Y=1.765
+ $X2=16.305 $Y2=2.4
r214 35 49 20.86 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=15.875 $Y=1.395
+ $X2=15.875 $Y2=1.58
r215 35 37 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=15.875 $Y=1.395
+ $X2=15.875 $Y2=0.95
r216 32 48 20.86 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=15.855 $Y=1.765
+ $X2=15.855 $Y2=1.58
r217 32 34 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=15.855 $Y=1.765
+ $X2=15.855 $Y2=2.4
r218 29 47 20.86 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=15.405 $Y=1.765
+ $X2=15.405 $Y2=1.58
r219 29 31 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=15.405 $Y=1.765
+ $X2=15.405 $Y2=2.4
r220 26 46 20.86 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=15.375 $Y=1.395
+ $X2=15.375 $Y2=1.58
r221 26 28 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=15.375 $Y=1.395
+ $X2=15.375 $Y2=0.95
r222 23 45 20.86 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=14.955 $Y=1.765
+ $X2=14.955 $Y2=1.58
r223 23 25 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=14.955 $Y=1.765
+ $X2=14.955 $Y2=2.4
r224 20 44 20.86 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=14.945 $Y=1.395
+ $X2=14.945 $Y2=1.58
r225 20 22 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=14.945 $Y=1.395
+ $X2=14.945 $Y2=0.95
r226 19 75 7.74396 $w=2.85e-07 $l=1.75e-07 $layer=POLY_cond $X=14.075 $Y=1.537
+ $X2=13.9 $Y2=1.537
r227 18 44 12.7189 $w=3.25e-07 $l=9.91968e-08 $layer=POLY_cond $X=14.865
+ $Y=1.537 $X2=14.945 $Y2=1.58
r228 18 19 166.279 $w=2.85e-07 $l=7.9e-07 $layer=POLY_cond $X=14.865 $Y=1.537
+ $X2=14.075 $Y2=1.537
r229 15 17 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=13.985 $Y=2.245
+ $X2=13.985 $Y2=2.64
r230 14 15 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=13.985 $Y=2.155
+ $X2=13.985 $Y2=2.245
r231 14 77 64.1371 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=13.985 $Y=2.155
+ $X2=13.985 $Y2=1.99
r232 11 74 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=13.955 $Y=0.58
+ $X2=13.955 $Y2=0.98
r233 8 75 23.4114 $w=3.5e-07 $l=1.42e-07 $layer=POLY_cond $X=13.9 $Y=1.395
+ $X2=13.9 $Y2=1.537
r234 7 68 1.64869 $w=3.5e-07 $l=1e-08 $layer=POLY_cond $X=13.9 $Y=1.155 $X2=13.9
+ $Y2=1.145
r235 7 8 39.5686 $w=3.5e-07 $l=2.4e-07 $layer=POLY_cond $X=13.9 $Y=1.155
+ $X2=13.9 $Y2=1.395
r236 2 60 600 $w=1.7e-07 $l=8.88819e-07 $layer=licon1_PDIFF $count=1 $X=12.42
+ $Y=1.96 $X2=12.63 $Y2=2.75
r237 1 54 182 $w=1.7e-07 $l=2.8801e-07 $layer=licon1_NDIFF $count=1 $X=12.015
+ $Y=0.37 $X2=12.2 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_LS__SEDFXTP_4%A_37_464# 1 2 3 4 14 17 19 22 23 24 26 27
+ 28 31 35 38 42 44 47 49
c124 19 0 1.8559e-19 $X=1.455 $Y=2.375
r125 39 42 5.47142 $w=4.68e-07 $l=2.15e-07 $layer=LI1_cond $X=0.17 $Y=0.575
+ $X2=0.385 $Y2=0.575
r126 38 49 4.3182 $w=2.1e-07 $l=1.03078e-07 $layer=LI1_cond $X=3.4 $Y=2.29
+ $X2=3.36 $Y2=2.375
r127 37 47 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.4 $Y=1.345
+ $X2=3.4 $Y2=1.26
r128 37 38 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=3.4 $Y=1.345
+ $X2=3.4 $Y2=2.29
r129 35 49 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.36 $Y=2.46 $X2=3.36
+ $Y2=2.375
r130 29 47 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=3.015 $Y=1.26
+ $X2=3.4 $Y2=1.26
r131 29 31 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=3.015 $Y=1.175
+ $X2=3.015 $Y2=0.775
r132 27 49 2.11342 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.235 $Y=2.375
+ $X2=3.36 $Y2=2.375
r133 27 28 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=3.235 $Y=2.375
+ $X2=2.305 $Y2=2.375
r134 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.22 $Y=2.46
+ $X2=2.305 $Y2=2.375
r135 25 26 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=2.22 $Y=2.46
+ $X2=2.22 $Y2=2.905
r136 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.135 $Y=2.99
+ $X2=2.22 $Y2=2.905
r137 23 24 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=2.135 $Y=2.99
+ $X2=1.625 $Y2=2.99
r138 22 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.54 $Y=2.905
+ $X2=1.625 $Y2=2.99
r139 21 22 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=1.54 $Y=2.46
+ $X2=1.54 $Y2=2.905
r140 20 44 3.3199 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=0.495 $Y=2.375
+ $X2=0.29 $Y2=2.375
r141 19 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.455 $Y=2.375
+ $X2=1.54 $Y2=2.46
r142 19 20 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.455 $Y=2.375
+ $X2=0.495 $Y2=2.375
r143 15 44 3.24686 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.29 $Y=2.46
+ $X2=0.29 $Y2=2.375
r144 15 17 0.140542 $w=4.08e-07 $l=5e-09 $layer=LI1_cond $X=0.29 $Y=2.46
+ $X2=0.29 $Y2=2.465
r145 14 44 3.24686 $w=2.9e-07 $l=1.56844e-07 $layer=LI1_cond $X=0.17 $Y=2.29
+ $X2=0.29 $Y2=2.375
r146 13 39 6.76998 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=0.17 $Y=0.81
+ $X2=0.17 $Y2=0.575
r147 13 14 96.5562 $w=1.68e-07 $l=1.48e-06 $layer=LI1_cond $X=0.17 $Y=0.81
+ $X2=0.17 $Y2=2.29
r148 4 35 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=3.25
+ $Y=2.315 $X2=3.4 $Y2=2.46
r149 3 17 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.185
+ $Y=2.32 $X2=0.33 $Y2=2.465
r150 2 31 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.875
+ $Y=0.565 $X2=3.015 $Y2=0.775
r151 1 42 182 $w=1.7e-07 $l=2.67862e-07 $layer=licon1_NDIFF $count=1 $X=0.24
+ $Y=0.37 $X2=0.385 $Y2=0.575
.ends

.subckt PM_SKY130_FD_SC_LS__SEDFXTP_4%VPWR 1 2 3 4 5 6 7 8 9 10 11 36 40 44 48
+ 52 56 60 64 66 70 76 78 80 83 84 85 87 92 97 102 107 116 120 125 130 136 139
+ 142 145 148 151 154 157 160 164
c195 3 0 9.53964e-20 $X=4.675 $Y=2.275
r196 163 164 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=16.56 $Y=3.33
+ $X2=16.56 $Y2=3.33
r197 160 161 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.6 $Y=3.33
+ $X2=15.6 $Y2=3.33
r198 157 158 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=14.64 $Y=3.33
+ $X2=14.64 $Y2=3.33
r199 155 158 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=13.68 $Y=3.33
+ $X2=14.64 $Y2=3.33
r200 154 155 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=3.33
+ $X2=13.68 $Y2=3.33
r201 151 152 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r202 148 149 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r203 145 146 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r204 142 143 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r205 139 140 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r206 136 137 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r207 134 164 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=16.08 $Y=3.33
+ $X2=16.56 $Y2=3.33
r208 134 161 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=16.08 $Y=3.33
+ $X2=15.6 $Y2=3.33
r209 133 134 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=16.08 $Y=3.33
+ $X2=16.08 $Y2=3.33
r210 131 160 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=15.795 $Y=3.33
+ $X2=15.63 $Y2=3.33
r211 131 133 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=15.795 $Y=3.33
+ $X2=16.08 $Y2=3.33
r212 130 163 4.76062 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=16.365 $Y=3.33
+ $X2=16.582 $Y2=3.33
r213 130 133 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=16.365 $Y=3.33
+ $X2=16.08 $Y2=3.33
r214 129 161 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=15.12 $Y=3.33
+ $X2=15.6 $Y2=3.33
r215 129 158 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=15.12 $Y=3.33
+ $X2=14.64 $Y2=3.33
r216 128 129 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.12 $Y=3.33
+ $X2=15.12 $Y2=3.33
r217 126 157 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.895 $Y=3.33
+ $X2=14.73 $Y2=3.33
r218 126 128 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=14.895 $Y=3.33
+ $X2=15.12 $Y2=3.33
r219 125 160 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=15.465 $Y=3.33
+ $X2=15.63 $Y2=3.33
r220 125 128 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=15.465 $Y=3.33
+ $X2=15.12 $Y2=3.33
r221 124 155 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=3.33
+ $X2=13.68 $Y2=3.33
r222 124 152 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=13.2 $Y=3.33
+ $X2=11.28 $Y2=3.33
r223 123 124 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=13.2 $Y=3.33
+ $X2=13.2 $Y2=3.33
r224 121 151 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.325 $Y=3.33
+ $X2=11.16 $Y2=3.33
r225 121 123 122.326 $w=1.68e-07 $l=1.875e-06 $layer=LI1_cond $X=11.325 $Y=3.33
+ $X2=13.2 $Y2=3.33
r226 120 154 11.8214 $w=1.7e-07 $l=2.7e-07 $layer=LI1_cond $X=13.335 $Y=3.33
+ $X2=13.605 $Y2=3.33
r227 120 123 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=13.335 $Y=3.33
+ $X2=13.2 $Y2=3.33
r228 119 152 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=11.28 $Y2=3.33
r229 118 119 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r230 116 151 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.995 $Y=3.33
+ $X2=11.16 $Y2=3.33
r231 116 118 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=10.995 $Y=3.33
+ $X2=10.8 $Y2=3.33
r232 115 119 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=10.8 $Y2=3.33
r233 114 115 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r234 112 148 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.94 $Y=3.33
+ $X2=7.775 $Y2=3.33
r235 112 114 123.957 $w=1.68e-07 $l=1.9e-06 $layer=LI1_cond $X=7.94 $Y=3.33
+ $X2=9.84 $Y2=3.33
r236 111 149 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r237 111 146 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6.48 $Y2=3.33
r238 110 111 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r239 108 145 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.59 $Y=3.33
+ $X2=6.425 $Y2=3.33
r240 108 110 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=6.59 $Y=3.33
+ $X2=7.44 $Y2=3.33
r241 107 148 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.61 $Y=3.33
+ $X2=7.775 $Y2=3.33
r242 107 110 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=7.61 $Y=3.33
+ $X2=7.44 $Y2=3.33
r243 106 146 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=6.48 $Y2=3.33
r244 106 143 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=5.04 $Y2=3.33
r245 105 106 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r246 103 142 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.22 $Y=3.33
+ $X2=5.095 $Y2=3.33
r247 103 105 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=5.22 $Y=3.33
+ $X2=6 $Y2=3.33
r248 102 145 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.26 $Y=3.33
+ $X2=6.425 $Y2=3.33
r249 102 105 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=6.26 $Y=3.33
+ $X2=6 $Y2=3.33
r250 101 143 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=5.04 $Y2=3.33
r251 101 140 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r252 100 101 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r253 98 139 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.725 $Y=3.33
+ $X2=2.6 $Y2=3.33
r254 98 100 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=2.725 $Y=3.33
+ $X2=3.12 $Y2=3.33
r255 97 142 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.97 $Y=3.33
+ $X2=5.095 $Y2=3.33
r256 97 100 120.695 $w=1.68e-07 $l=1.85e-06 $layer=LI1_cond $X=4.97 $Y=3.33
+ $X2=3.12 $Y2=3.33
r257 96 140 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r258 96 137 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.2 $Y2=3.33
r259 95 96 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r260 93 136 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.285 $Y=3.33
+ $X2=1.16 $Y2=3.33
r261 93 95 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=1.285 $Y=3.33
+ $X2=2.16 $Y2=3.33
r262 92 139 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.475 $Y=3.33
+ $X2=2.6 $Y2=3.33
r263 92 95 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.475 $Y=3.33
+ $X2=2.16 $Y2=3.33
r264 90 137 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r265 89 90 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r266 87 136 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.035 $Y=3.33
+ $X2=1.16 $Y2=3.33
r267 87 89 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.035 $Y=3.33
+ $X2=0.72 $Y2=3.33
r268 85 115 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=9.84 $Y2=3.33
r269 85 149 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=7.92 $Y2=3.33
r270 83 114 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=9.96 $Y=3.33
+ $X2=9.84 $Y2=3.33
r271 83 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.96 $Y=3.33
+ $X2=10.125 $Y2=3.33
r272 82 118 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=10.29 $Y=3.33
+ $X2=10.8 $Y2=3.33
r273 82 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.29 $Y=3.33
+ $X2=10.125 $Y2=3.33
r274 78 163 3.00555 $w=3.3e-07 $l=1.07912e-07 $layer=LI1_cond $X=16.53 $Y=3.245
+ $X2=16.582 $Y2=3.33
r275 78 80 29.3349 $w=3.28e-07 $l=8.4e-07 $layer=LI1_cond $X=16.53 $Y=3.245
+ $X2=16.53 $Y2=2.405
r276 74 160 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=15.63 $Y=3.245
+ $X2=15.63 $Y2=3.33
r277 74 76 29.3349 $w=3.28e-07 $l=8.4e-07 $layer=LI1_cond $X=15.63 $Y=3.245
+ $X2=15.63 $Y2=2.405
r278 70 73 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=14.73 $Y=2.035
+ $X2=14.73 $Y2=2.815
r279 68 157 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=14.73 $Y=3.245
+ $X2=14.73 $Y2=3.33
r280 68 73 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=14.73 $Y=3.245
+ $X2=14.73 $Y2=2.815
r281 67 154 11.8214 $w=1.7e-07 $l=2.7e-07 $layer=LI1_cond $X=13.875 $Y=3.33
+ $X2=13.605 $Y2=3.33
r282 66 157 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.565 $Y=3.33
+ $X2=14.73 $Y2=3.33
r283 66 67 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=14.565 $Y=3.33
+ $X2=13.875 $Y2=3.33
r284 62 154 2.26835 $w=5.4e-07 $l=8.5e-08 $layer=LI1_cond $X=13.605 $Y=3.245
+ $X2=13.605 $Y2=3.33
r285 62 64 9.52433 $w=5.38e-07 $l=4.3e-07 $layer=LI1_cond $X=13.605 $Y=3.245
+ $X2=13.605 $Y2=2.815
r286 58 151 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.16 $Y=3.245
+ $X2=11.16 $Y2=3.33
r287 58 60 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=11.16 $Y=3.245
+ $X2=11.16 $Y2=2.815
r288 54 84 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.125 $Y=3.245
+ $X2=10.125 $Y2=3.33
r289 54 56 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=10.125 $Y=3.245
+ $X2=10.125 $Y2=2.815
r290 50 148 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.775 $Y=3.245
+ $X2=7.775 $Y2=3.33
r291 50 52 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=7.775 $Y=3.245
+ $X2=7.775 $Y2=2.785
r292 46 145 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.425 $Y=3.245
+ $X2=6.425 $Y2=3.33
r293 46 48 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=6.425 $Y=3.245
+ $X2=6.425 $Y2=2.77
r294 42 142 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.095 $Y=3.245
+ $X2=5.095 $Y2=3.33
r295 42 44 22.1269 $w=2.48e-07 $l=4.8e-07 $layer=LI1_cond $X=5.095 $Y=3.245
+ $X2=5.095 $Y2=2.765
r296 38 139 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.6 $Y=3.245
+ $X2=2.6 $Y2=3.33
r297 38 40 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=2.6 $Y=3.245
+ $X2=2.6 $Y2=2.8
r298 34 136 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.16 $Y=3.245
+ $X2=1.16 $Y2=3.33
r299 34 36 20.283 $w=2.48e-07 $l=4.4e-07 $layer=LI1_cond $X=1.16 $Y=3.245
+ $X2=1.16 $Y2=2.805
r300 11 80 300 $w=1.7e-07 $l=6.3559e-07 $layer=licon1_PDIFF $count=2 $X=16.38
+ $Y=1.84 $X2=16.53 $Y2=2.405
r301 10 76 300 $w=1.7e-07 $l=6.3559e-07 $layer=licon1_PDIFF $count=2 $X=15.48
+ $Y=1.84 $X2=15.63 $Y2=2.405
r302 9 73 400 $w=1.7e-07 $l=1.03562e-06 $layer=licon1_PDIFF $count=1 $X=14.605
+ $Y=1.84 $X2=14.73 $Y2=2.815
r303 9 70 400 $w=1.7e-07 $l=2.498e-07 $layer=licon1_PDIFF $count=1 $X=14.605
+ $Y=1.84 $X2=14.73 $Y2=2.035
r304 8 64 600 $w=1.7e-07 $l=3.81772e-07 $layer=licon1_PDIFF $count=1 $X=13.35
+ $Y=2.54 $X2=13.605 $Y2=2.815
r305 7 60 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=11.035
+ $Y=1.96 $X2=11.16 $Y2=2.815
r306 6 56 600 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=9.975
+ $Y=2.54 $X2=10.125 $Y2=2.815
r307 5 52 600 $w=1.7e-07 $l=1.00556e-06 $layer=licon1_PDIFF $count=1 $X=7.65
+ $Y=1.84 $X2=7.775 $Y2=2.785
r308 4 48 600 $w=1.7e-07 $l=1.02795e-06 $layer=licon1_PDIFF $count=1 $X=6.295
+ $Y=1.805 $X2=6.425 $Y2=2.77
r309 3 44 600 $w=1.7e-07 $l=6.52917e-07 $layer=licon1_PDIFF $count=1 $X=4.675
+ $Y=2.275 $X2=5.055 $Y2=2.765
r310 2 40 600 $w=1.7e-07 $l=6.47708e-07 $layer=licon1_PDIFF $count=1 $X=2.18
+ $Y=2.315 $X2=2.56 $Y2=2.8
r311 1 36 600 $w=1.7e-07 $l=5.54955e-07 $layer=licon1_PDIFF $count=1 $X=1.05
+ $Y=2.32 $X2=1.2 $Y2=2.805
.ends

.subckt PM_SKY130_FD_SC_LS__SEDFXTP_4%A_661_113# 1 2 3 4 5 6 21 24 25 26 28 30
+ 33 38 39 42 43 44 45 49 54 56 59 62 63 65 66
c177 56 0 1.85697e-19 $X=3.795 $Y=2.295
c178 25 0 9.53964e-20 $X=4.63 $Y=2.99
r179 64 65 5.10546 $w=2.48e-07 $l=8.5e-08 $layer=LI1_cond $X=6.115 $Y=2.38
+ $X2=6.2 $Y2=2.38
r180 62 64 10.1415 $w=2.48e-07 $l=2.2e-07 $layer=LI1_cond $X=5.895 $Y=2.38
+ $X2=6.115 $Y2=2.38
r181 62 63 8.79328 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=5.895 $Y=2.38
+ $X2=5.73 $Y2=2.38
r182 52 54 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=3.585 $Y=0.84
+ $X2=3.74 $Y2=0.84
r183 47 49 33.1904 $w=2.48e-07 $l=7.2e-07 $layer=LI1_cond $X=8.2 $Y=1.48 $X2=8.2
+ $Y2=0.76
r184 46 66 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.89 $Y=2.42
+ $X2=7.805 $Y2=2.42
r185 45 68 19.844 $w=5.17e-07 $l=6.9852e-07 $layer=LI1_cond $X=8.155 $Y=2.42
+ $X2=8.745 $Y2=2.657
r186 45 46 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=8.155 $Y=2.42
+ $X2=7.89 $Y2=2.42
r187 43 47 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=8.075 $Y=1.565
+ $X2=8.2 $Y2=1.48
r188 43 44 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=8.075 $Y=1.565
+ $X2=7.89 $Y2=1.565
r189 42 66 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.805 $Y=2.335
+ $X2=7.805 $Y2=2.42
r190 41 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.805 $Y=1.65
+ $X2=7.89 $Y2=1.565
r191 41 42 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=7.805 $Y=1.65
+ $X2=7.805 $Y2=2.335
r192 39 66 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.72 $Y=2.42
+ $X2=7.805 $Y2=2.42
r193 39 65 99.1658 $w=1.68e-07 $l=1.52e-06 $layer=LI1_cond $X=7.72 $Y=2.42
+ $X2=6.2 $Y2=2.42
r194 38 64 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.115 $Y=2.255
+ $X2=6.115 $Y2=2.38
r195 37 59 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.115 $Y=1.245
+ $X2=6.115 $Y2=1.16
r196 37 38 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=6.115 $Y=1.245
+ $X2=6.115 $Y2=2.255
r197 31 59 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=5.72 $Y=1.16
+ $X2=6.115 $Y2=1.16
r198 31 33 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=5.72 $Y=1.075
+ $X2=5.72 $Y2=0.835
r199 30 63 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=4.8 $Y=2.34
+ $X2=5.73 $Y2=2.34
r200 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.715 $Y=2.425
+ $X2=4.8 $Y2=2.34
r201 27 28 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=4.715 $Y=2.425
+ $X2=4.715 $Y2=2.905
r202 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.63 $Y=2.99
+ $X2=4.715 $Y2=2.905
r203 25 26 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=4.63 $Y=2.99
+ $X2=3.935 $Y2=2.99
r204 22 26 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=3.795 $Y=2.905
+ $X2=3.935 $Y2=2.99
r205 22 24 18.3156 $w=2.78e-07 $l=4.45e-07 $layer=LI1_cond $X=3.795 $Y=2.905
+ $X2=3.795 $Y2=2.46
r206 21 56 7.52792 $w=2.78e-07 $l=1.4e-07 $layer=LI1_cond $X=3.795 $Y=2.435
+ $X2=3.795 $Y2=2.295
r207 21 24 1.02897 $w=2.78e-07 $l=2.5e-08 $layer=LI1_cond $X=3.795 $Y=2.435
+ $X2=3.795 $Y2=2.46
r208 19 54 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.74 $Y=1.005
+ $X2=3.74 $Y2=0.84
r209 19 56 84.1604 $w=1.68e-07 $l=1.29e-06 $layer=LI1_cond $X=3.74 $Y=1.005
+ $X2=3.74 $Y2=2.295
r210 6 68 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=8.62
+ $Y=2.54 $X2=8.745 $Y2=2.75
r211 5 62 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=5.745
+ $Y=2.275 $X2=5.895 $Y2=2.42
r212 4 24 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=3.7
+ $Y=2.315 $X2=3.85 $Y2=2.46
r213 3 49 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=8.1
+ $Y=0.485 $X2=8.24 $Y2=0.76
r214 2 33 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=5.58
+ $Y=0.625 $X2=5.72 $Y2=0.835
r215 1 52 182 $w=1.7e-07 $l=3.94208e-07 $layer=licon1_NDIFF $count=1 $X=3.305
+ $Y=0.565 $X2=3.585 $Y2=0.84
.ends

.subckt PM_SKY130_FD_SC_LS__SEDFXTP_4%Q 1 2 3 4 15 19 23 27 29
r52 41 43 0.178016 $w=1.028e-06 $l=1.5e-08 $layer=LI1_cond $X=16.08 $Y=1.62
+ $X2=16.095 $Y2=1.62
r53 39 41 0.0356031 $w=1.028e-06 $l=3e-09 $layer=LI1_cond $X=16.077 $Y=1.62
+ $X2=16.08 $Y2=1.62
r54 38 39 10.408 $w=1.028e-06 $l=8.77e-07 $layer=LI1_cond $X=15.2 $Y=1.62
+ $X2=16.077 $Y2=1.62
r55 37 38 0.237354 $w=1.028e-06 $l=2e-08 $layer=LI1_cond $X=15.18 $Y=1.62
+ $X2=15.2 $Y2=1.62
r56 35 37 0.0593385 $w=1.028e-06 $l=5e-09 $layer=LI1_cond $X=15.175 $Y=1.62
+ $X2=15.18 $Y2=1.62
r57 29 43 5.51848 $w=1.028e-06 $l=4.65e-07 $layer=LI1_cond $X=16.56 $Y=1.62
+ $X2=16.095 $Y2=1.62
r58 25 43 10.6424 $w=2.05e-07 $l=5.30999e-07 $layer=LI1_cond $X=16.097 $Y=1.09
+ $X2=16.095 $Y2=1.62
r59 25 27 18.9357 $w=2.03e-07 $l=3.5e-07 $layer=LI1_cond $X=16.097 $Y=1.09
+ $X2=16.097 $Y2=0.74
r60 21 39 10.3216 $w=2.15e-07 $l=5.3e-07 $layer=LI1_cond $X=16.077 $Y=2.15
+ $X2=16.077 $Y2=1.62
r61 21 23 15.8126 $w=2.13e-07 $l=2.95e-07 $layer=LI1_cond $X=16.077 $Y=2.15
+ $X2=16.077 $Y2=2.445
r62 17 38 9.31248 $w=2.5e-07 $l=5.3e-07 $layer=LI1_cond $X=15.2 $Y=1.09 $X2=15.2
+ $Y2=1.62
r63 17 19 16.8257 $w=2.48e-07 $l=3.65e-07 $layer=LI1_cond $X=15.2 $Y=1.09
+ $X2=15.2 $Y2=0.725
r64 13 35 10.1615 $w=2.2e-07 $l=5.3e-07 $layer=LI1_cond $X=15.175 $Y=2.15
+ $X2=15.175 $Y2=1.62
r65 13 15 15.4532 $w=2.18e-07 $l=2.95e-07 $layer=LI1_cond $X=15.175 $Y=2.15
+ $X2=15.175 $Y2=2.445
r66 4 41 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=15.93
+ $Y=1.84 $X2=16.08 $Y2=1.985
r67 4 23 300 $w=1.7e-07 $l=6.75851e-07 $layer=licon1_PDIFF $count=2 $X=15.93
+ $Y=1.84 $X2=16.08 $Y2=2.445
r68 3 37 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=15.03
+ $Y=1.84 $X2=15.18 $Y2=1.985
r69 3 15 300 $w=1.7e-07 $l=6.75851e-07 $layer=licon1_PDIFF $count=2 $X=15.03
+ $Y=1.84 $X2=15.18 $Y2=2.445
r70 2 43 182 $w=1.7e-07 $l=6.63551e-07 $layer=licon1_NDIFF $count=1 $X=15.95
+ $Y=0.58 $X2=16.095 $Y2=1.175
r71 2 27 182 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=1 $X=15.95
+ $Y=0.58 $X2=16.095 $Y2=0.74
r72 1 19 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=15.02
+ $Y=0.58 $X2=15.16 $Y2=0.725
.ends

.subckt PM_SKY130_FD_SC_LS__SEDFXTP_4%VGND 1 2 3 4 5 6 7 8 9 10 11 36 40 44 48
+ 52 56 60 62 66 70 72 74 77 78 80 81 82 84 89 94 109 113 126 131 137 140 143
+ 146 149 153 157 159 162 166
c210 36 0 1.82239e-19 $X=1.205 $Y=0.58
r211 165 166 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=16.56 $Y=0
+ $X2=16.56 $Y2=0
r212 162 163 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.6 $Y=0
+ $X2=15.6 $Y2=0
r213 159 160 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=14.64 $Y=0
+ $X2=14.64 $Y2=0
r214 156 160 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=13.68 $Y=0
+ $X2=14.64 $Y2=0
r215 155 157 11.0607 $w=7.63e-07 $l=1.55e-07 $layer=LI1_cond $X=13.68 $Y=0.297
+ $X2=13.835 $Y2=0.297
r216 155 156 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.68 $Y=0
+ $X2=13.68 $Y2=0
r217 152 155 0.15635 $w=7.63e-07 $l=1e-08 $layer=LI1_cond $X=13.67 $Y=0.297
+ $X2=13.68 $Y2=0.297
r218 152 153 21.3798 $w=7.63e-07 $l=8.15e-07 $layer=LI1_cond $X=13.67 $Y=0.297
+ $X2=12.855 $Y2=0.297
r219 149 150 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r220 146 147 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=9.84 $Y=0
+ $X2=9.84 $Y2=0
r221 143 144 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r222 140 141 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r223 137 138 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r224 135 166 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=16.08 $Y=0
+ $X2=16.56 $Y2=0
r225 135 163 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=16.08 $Y=0
+ $X2=15.6 $Y2=0
r226 134 135 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=16.08 $Y=0
+ $X2=16.08 $Y2=0
r227 132 162 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=15.825 $Y=0
+ $X2=15.66 $Y2=0
r228 132 134 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=15.825 $Y=0
+ $X2=16.08 $Y2=0
r229 131 165 4.77065 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=16.37 $Y=0
+ $X2=16.585 $Y2=0
r230 131 134 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=16.37 $Y=0
+ $X2=16.08 $Y2=0
r231 130 163 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=15.12 $Y=0
+ $X2=15.6 $Y2=0
r232 130 160 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=15.12 $Y=0
+ $X2=14.64 $Y2=0
r233 129 130 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.12 $Y=0
+ $X2=15.12 $Y2=0
r234 127 159 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.895 $Y=0
+ $X2=14.73 $Y2=0
r235 127 129 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=14.895 $Y=0
+ $X2=15.12 $Y2=0
r236 126 162 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=15.495 $Y=0
+ $X2=15.66 $Y2=0
r237 126 129 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=15.495 $Y=0
+ $X2=15.12 $Y2=0
r238 125 156 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=12.72 $Y=0
+ $X2=13.68 $Y2=0
r239 124 153 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=12.72 $Y=0
+ $X2=12.855 $Y2=0
r240 124 125 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r241 122 125 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=12.72 $Y2=0
r242 122 150 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=11.28 $Y2=0
r243 121 124 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=11.76 $Y=0
+ $X2=12.72 $Y2=0
r244 121 122 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r245 119 149 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.53 $Y=0
+ $X2=11.405 $Y2=0
r246 119 121 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=11.53 $Y=0
+ $X2=11.76 $Y2=0
r247 117 150 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=11.28 $Y2=0
r248 117 147 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=9.84 $Y2=0
r249 116 117 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r250 114 146 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.09 $Y=0
+ $X2=9.965 $Y2=0
r251 114 116 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=10.09 $Y=0
+ $X2=10.32 $Y2=0
r252 113 149 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.28 $Y=0
+ $X2=11.405 $Y2=0
r253 113 116 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=11.28 $Y=0
+ $X2=10.32 $Y2=0
r254 111 112 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r255 109 146 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.84 $Y=0
+ $X2=9.965 $Y2=0
r256 109 111 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=9.84 $Y=0
+ $X2=7.44 $Y2=0
r257 108 112 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0
+ $X2=7.44 $Y2=0
r258 107 108 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r259 105 108 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.96
+ $Y2=0
r260 105 144 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.04
+ $Y2=0
r261 104 105 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6
+ $Y2=0
r262 102 143 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.095 $Y=0
+ $X2=4.93 $Y2=0
r263 102 104 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=5.095 $Y=0 $X2=6
+ $Y2=0
r264 101 144 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0
+ $X2=5.04 $Y2=0
r265 100 101 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r266 98 101 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=4.56 $Y2=0
r267 98 141 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=2.16 $Y2=0
r268 97 100 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=2.64 $Y=0
+ $X2=4.56 $Y2=0
r269 97 98 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r270 95 140 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.36 $Y=0
+ $X2=2.195 $Y2=0
r271 95 97 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=2.36 $Y=0 $X2=2.64
+ $Y2=0
r272 94 143 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.765 $Y=0
+ $X2=4.93 $Y2=0
r273 94 100 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=4.765 $Y=0
+ $X2=4.56 $Y2=0
r274 93 141 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0
+ $X2=2.16 $Y2=0
r275 93 138 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r276 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r277 90 137 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.37 $Y=0
+ $X2=1.205 $Y2=0
r278 90 92 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1.37 $Y=0 $X2=1.68
+ $Y2=0
r279 89 140 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.03 $Y=0
+ $X2=2.195 $Y2=0
r280 89 92 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=2.03 $Y=0 $X2=1.68
+ $Y2=0
r281 87 138 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r282 86 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r283 84 137 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.04 $Y=0
+ $X2=1.205 $Y2=0
r284 84 86 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.04 $Y=0 $X2=0.72
+ $Y2=0
r285 82 147 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=8.4 $Y=0
+ $X2=9.84 $Y2=0
r286 82 112 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=7.44
+ $Y2=0
r287 80 107 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=7.095 $Y=0
+ $X2=6.96 $Y2=0
r288 80 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.095 $Y=0 $X2=7.26
+ $Y2=0
r289 79 111 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=7.425 $Y=0
+ $X2=7.44 $Y2=0
r290 79 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.425 $Y=0 $X2=7.26
+ $Y2=0
r291 77 104 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=6.11 $Y=0 $X2=6
+ $Y2=0
r292 77 78 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.11 $Y=0 $X2=6.235
+ $Y2=0
r293 76 107 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=6.36 $Y=0 $X2=6.96
+ $Y2=0
r294 76 78 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.36 $Y=0 $X2=6.235
+ $Y2=0
r295 72 165 2.99552 $w=3.3e-07 $l=1.07121e-07 $layer=LI1_cond $X=16.535 $Y=0.085
+ $X2=16.585 $Y2=0
r296 72 74 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=16.535 $Y=0.085
+ $X2=16.535 $Y2=0.74
r297 68 162 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=15.66 $Y=0.085
+ $X2=15.66 $Y2=0
r298 68 70 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=15.66 $Y=0.085
+ $X2=15.66 $Y2=0.74
r299 64 159 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=14.73 $Y=0.085
+ $X2=14.73 $Y2=0
r300 64 66 22.3504 $w=3.28e-07 $l=6.4e-07 $layer=LI1_cond $X=14.73 $Y=0.085
+ $X2=14.73 $Y2=0.725
r301 62 159 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.565 $Y=0
+ $X2=14.73 $Y2=0
r302 62 157 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=14.565 $Y=0
+ $X2=13.835 $Y2=0
r303 58 149 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=11.405 $Y=0.085
+ $X2=11.405 $Y2=0
r304 58 60 20.0525 $w=2.48e-07 $l=4.35e-07 $layer=LI1_cond $X=11.405 $Y=0.085
+ $X2=11.405 $Y2=0.52
r305 54 146 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.965 $Y=0.085
+ $X2=9.965 $Y2=0
r306 54 56 20.283 $w=2.48e-07 $l=4.4e-07 $layer=LI1_cond $X=9.965 $Y=0.085
+ $X2=9.965 $Y2=0.525
r307 50 81 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.26 $Y=0.085
+ $X2=7.26 $Y2=0
r308 50 52 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=7.26 $Y=0.085
+ $X2=7.26 $Y2=0.55
r309 46 78 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.235 $Y=0.085
+ $X2=6.235 $Y2=0
r310 46 48 24.6623 $w=2.48e-07 $l=5.35e-07 $layer=LI1_cond $X=6.235 $Y=0.085
+ $X2=6.235 $Y2=0.62
r311 42 143 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.93 $Y=0.085
+ $X2=4.93 $Y2=0
r312 42 44 25.1442 $w=3.28e-07 $l=7.2e-07 $layer=LI1_cond $X=4.93 $Y=0.085
+ $X2=4.93 $Y2=0.805
r313 38 140 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.195 $Y=0.085
+ $X2=2.195 $Y2=0
r314 38 40 24.0965 $w=3.28e-07 $l=6.9e-07 $layer=LI1_cond $X=2.195 $Y=0.085
+ $X2=2.195 $Y2=0.775
r315 34 137 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=0.085
+ $X2=1.205 $Y2=0
r316 34 36 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=1.205 $Y=0.085
+ $X2=1.205 $Y2=0.58
r317 11 74 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=16.395
+ $Y=0.58 $X2=16.535 $Y2=0.74
r318 10 70 182 $w=1.7e-07 $l=2.78747e-07 $layer=licon1_NDIFF $count=1 $X=15.45
+ $Y=0.58 $X2=15.66 $Y2=0.74
r319 9 66 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=14.585
+ $Y=0.58 $X2=14.73 $Y2=0.725
r320 8 152 91 $w=1.7e-07 $l=8.59448e-07 $layer=licon1_NDIFF $count=2 $X=12.88
+ $Y=0.37 $X2=13.67 $Y2=0.515
r321 7 60 182 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_NDIFF $count=1 $X=11.22
+ $Y=0.37 $X2=11.365 $Y2=0.52
r322 6 56 182 $w=1.7e-07 $l=1.94422e-07 $layer=licon1_NDIFF $count=1 $X=9.865
+ $Y=0.395 $X2=10.005 $Y2=0.525
r323 5 52 182 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_NDIFF $count=1 $X=7.115
+ $Y=0.37 $X2=7.26 $Y2=0.55
r324 4 48 182 $w=1.7e-07 $l=3.14245e-07 $layer=licon1_NDIFF $count=1 $X=6.13
+ $Y=0.37 $X2=6.275 $Y2=0.62
r325 3 44 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=4.79
+ $Y=0.625 $X2=4.93 $Y2=0.805
r326 2 40 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.055
+ $Y=0.565 $X2=2.195 $Y2=0.775
r327 1 36 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.065
+ $Y=0.37 $X2=1.205 $Y2=0.58
.ends

