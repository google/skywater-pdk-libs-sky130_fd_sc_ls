* File: sky130_fd_sc_ls__nand3_4.spice
* Created: Fri Aug 28 13:33:38 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__nand3_4.pex.spice"
.subckt sky130_fd_sc_ls__nand3_4  VNB VPB A B C VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* C	C
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1005 N_Y_M1005_d N_A_M1005_g N_A_27_82#_M1005_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.19525 PD=1.02 PS=2.03 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75003.2 A=0.111 P=1.78 MULT=1
MM1012 N_Y_M1005_d N_A_M1012_g N_A_27_82#_M1012_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75002.8 A=0.111 P=1.78 MULT=1
MM1013 N_Y_M1013_d N_A_M1013_g N_A_27_82#_M1012_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001
+ SB=75002.3 A=0.111 P=1.78 MULT=1
MM1016 N_Y_M1013_d N_A_M1016_g N_A_27_82#_M1016_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75001.9 A=0.111 P=1.78 MULT=1
MM1003 N_A_27_82#_M1016_s N_B_M1003_g N_A_456_82#_M1003_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.9 SB=75001.5 A=0.111 P=1.78 MULT=1
MM1004 N_A_27_82#_M1004_d N_B_M1004_g N_A_456_82#_M1003_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75002.3 SB=75001 A=0.111 P=1.78 MULT=1
MM1009 N_A_27_82#_M1004_d N_B_M1009_g N_A_456_82#_M1009_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75002.8 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1015 N_A_27_82#_M1015_d N_B_M1015_g N_A_456_82#_M1009_s VNB NSHORT L=0.15
+ W=0.74 AD=0.19525 AS=0.1036 PD=2.03 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75003.2 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1000 N_A_456_82#_M1000_d N_C_M1000_g N_VGND_M1000_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.2035 PD=1.02 PS=2.03 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.5 A=0.111 P=1.78 MULT=1
MM1001 N_A_456_82#_M1000_d N_C_M1001_g N_VGND_M1001_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1007 N_A_456_82#_M1007_d N_C_M1007_g N_VGND_M1001_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1010 N_A_456_82#_M1007_d N_C_M1010_g N_VGND_M1010_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.2035 PD=1.02 PS=2.03 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1006 N_VPWR_M1006_d N_A_M1006_g N_Y_M1006_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.4592 PD=2.83 PS=1.94 NRD=1.7533 NRS=2.6201 M=1 R=7.46667
+ SA=75000.2 SB=75005.1 A=0.168 P=2.54 MULT=1
MM1011 N_VPWR_M1011_d N_A_M1011_g N_Y_M1006_s VPB PHIGHVT L=0.15 W=1.12 AD=0.196
+ AS=0.4592 PD=1.47 PS=1.94 NRD=1.7533 NRS=2.6201 M=1 R=7.46667 SA=75001.2
+ SB=75004.1 A=0.168 P=2.54 MULT=1
MM1008 N_Y_M1008_d N_B_M1008_g N_VPWR_M1011_d VPB PHIGHVT L=0.15 W=1.12 AD=0.168
+ AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667 SA=75001.7
+ SB=75003.6 A=0.168 P=2.54 MULT=1
MM1014 N_Y_M1008_d N_B_M1014_g N_VPWR_M1014_s VPB PHIGHVT L=0.15 W=1.12 AD=0.168
+ AS=0.742 PD=1.42 PS=2.445 NRD=1.7533 NRS=2.6201 M=1 R=7.46667 SA=75002.1
+ SB=75003.2 A=0.168 P=2.54 MULT=1
MM1002 N_VPWR_M1014_s N_C_M1002_g N_Y_M1002_s VPB PHIGHVT L=0.15 W=1.12 AD=0.742
+ AS=0.168 PD=2.445 PS=1.42 NRD=2.6201 NRS=1.7533 M=1 R=7.46667 SA=75003.6
+ SB=75001.7 A=0.168 P=2.54 MULT=1
MM1017 N_VPWR_M1017_d N_C_M1017_g N_Y_M1002_s VPB PHIGHVT L=0.15 W=1.12 AD=1.484
+ AS=0.168 PD=4.89 PS=1.42 NRD=2.6201 NRS=1.7533 M=1 R=7.46667 SA=75004.1
+ SB=75001.2 A=0.168 P=2.54 MULT=1
DX18_noxref VNB VPB NWDIODE A=12.3132 P=16.96
*
.include "sky130_fd_sc_ls__nand3_4.pxi.spice"
*
.ends
*
*
