* File: sky130_fd_sc_ls__decaphe_8.pxi.spice
* Created: Wed Sep  2 11:00:08 2020
* 
x_PM_SKY130_FD_SC_LS__DECAPHE_8%VGND N_VGND_M1000_s VGND N_VGND_M1001_g
+ N_VGND_c_12_n N_VGND_c_13_n PM_SKY130_FD_SC_LS__DECAPHE_8%VGND
x_PM_SKY130_FD_SC_LS__DECAPHE_8%VPWR N_VPWR_M1001_s N_VPWR_c_21_n N_VPWR_c_22_n
+ N_VPWR_M1000_g VPWR N_VPWR_c_24_n VPWR PM_SKY130_FD_SC_LS__DECAPHE_8%VPWR
cc_1 VNB N_VGND_M1001_g 0.0884661f $X=-0.19 $Y=-0.245 $X2=1.92 $Y2=2.467
cc_2 VNB N_VGND_c_12_n 0.174462f $X=-0.19 $Y=-0.245 $X2=3.58 $Y2=0.38
cc_3 VNB N_VGND_c_13_n 0.206277f $X=-0.19 $Y=-0.245 $X2=3.6 $Y2=0
cc_4 VNB N_VPWR_c_21_n 0.172799f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_5 VNB N_VPWR_c_22_n 0.145486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB VPWR 0.163682f $X=-0.19 $Y=-0.245 $X2=0.765 $Y2=1.515
cc_7 VNB N_VPWR_c_24_n 0.028581f $X=-0.19 $Y=-0.245 $X2=3.58 $Y2=0.38
cc_8 VPB N_VGND_M1001_g 0.230199f $X=-0.19 $Y=1.66 $X2=1.92 $Y2=2.467
cc_9 VPB VPWR 0.0425959f $X=-0.19 $Y=1.66 $X2=0.765 $Y2=1.515
cc_10 VPB N_VPWR_c_24_n 0.187292f $X=-0.19 $Y=1.66 $X2=3.58 $Y2=0.38
cc_11 N_VGND_M1001_g N_VPWR_c_21_n 0.0923543f $X=1.92 $Y=2.467 $X2=0 $Y2=0
cc_12 N_VGND_c_12_n N_VPWR_c_21_n 0.227804f $X=3.58 $Y=0.38 $X2=0 $Y2=0
cc_13 N_VGND_M1001_g N_VPWR_c_22_n 0.100861f $X=1.92 $Y=2.467 $X2=0 $Y2=0
cc_14 N_VGND_c_12_n N_VPWR_c_22_n 0.199723f $X=3.58 $Y=0.38 $X2=0 $Y2=0
cc_15 N_VGND_M1001_g N_VPWR_c_24_n 0.569394f $X=1.92 $Y=2.467 $X2=0 $Y2=0
cc_16 N_VGND_c_12_n N_VPWR_c_24_n 0.366433f $X=3.58 $Y=0.38 $X2=0 $Y2=0
