* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__or2b_4 A B_N VGND VNB VPB VPWR X
X0 a_81_296# A VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X1 VPWR a_81_296# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X2 X a_81_296# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X3 VPWR A a_489_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 VPWR a_81_296# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X5 X a_81_296# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X6 a_489_392# a_676_48# a_81_296# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 VGND B_N a_676_48# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X8 X a_81_296# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X9 a_489_392# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 X a_81_296# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X11 VPWR B_N a_676_48# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 VGND a_676_48# a_81_296# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X13 VGND a_81_296# X VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X14 VGND A a_81_296# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X15 a_81_296# a_676_48# VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X16 VGND a_81_296# X VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X17 a_81_296# a_676_48# a_489_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends
