* File: sky130_fd_sc_ls__o22ai_1.spice
* Created: Wed Sep  2 11:20:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__o22ai_1.pex.spice"
.subckt sky130_fd_sc_ls__o22ai_1  VNB VPB B1 B2 A2 A1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A1	A1
* A2	A2
* B2	B2
* B1	B1
* VPB	VPB
* VNB	VNB
MM1007 N_Y_M1007_d N_B1_M1007_g N_A_27_74#_M1007_s VNB NSHORT L=0.15 W=0.74
+ AD=0.21275 AS=0.2109 PD=1.315 PS=2.05 NRD=23.508 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75002 A=0.111 P=1.78 MULT=1
MM1002 N_A_27_74#_M1002_d N_B2_M1002_g N_Y_M1007_d VNB NSHORT L=0.15 W=0.74
+ AD=0.1295 AS=0.21275 PD=1.09 PS=1.315 NRD=11.34 NRS=24.324 M=1 R=4.93333
+ SA=75000.9 SB=75001.3 A=0.111 P=1.78 MULT=1
MM1001 N_VGND_M1001_d N_A2_M1001_g N_A_27_74#_M1002_d VNB NSHORT L=0.15 W=0.74
+ AD=0.1554 AS=0.1295 PD=1.16 PS=1.09 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75001.4
+ SB=75000.8 A=0.111 P=1.78 MULT=1
MM1003 N_A_27_74#_M1003_d N_A1_M1003_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.1554 PD=2.05 PS=1.16 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75002
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1000 A_142_368# N_B1_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.1512 AS=0.4648 PD=1.39 PS=3.07 NRD=14.0658 NRS=22.852 M=1 R=7.46667
+ SA=75000.3 SB=75001.8 A=0.168 P=2.54 MULT=1
MM1005 N_Y_M1005_d N_B2_M1005_g A_142_368# VPB PHIGHVT L=0.15 W=1.12 AD=0.2352
+ AS=0.1512 PD=1.54 PS=1.39 NRD=11.426 NRS=14.0658 M=1 R=7.46667 SA=75000.8
+ SB=75001.4 A=0.168 P=2.54 MULT=1
MM1006 A_340_368# N_A2_M1006_g N_Y_M1005_d VPB PHIGHVT L=0.15 W=1.12 AD=0.2352
+ AS=0.2352 PD=1.54 PS=1.54 NRD=27.2451 NRS=13.1793 M=1 R=7.46667 SA=75001.3
+ SB=75000.8 A=0.168 P=2.54 MULT=1
MM1004 N_VPWR_M1004_d N_A1_M1004_g A_340_368# VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.2352 PD=2.83 PS=1.54 NRD=1.7533 NRS=27.2451 M=1 R=7.46667
+ SA=75001.9 SB=75000.2 A=0.168 P=2.54 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.0636 P=10.24
*
.include "sky130_fd_sc_ls__o22ai_1.pxi.spice"
*
.ends
*
*
