* File: sky130_fd_sc_ls__xnor3_4.spice
* Created: Wed Sep  2 11:30:46 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__xnor3_4.pex.spice"
.subckt sky130_fd_sc_ls__xnor3_4  VNB VPB A B C VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* C	C
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1012 N_VGND_M1012_d N_A_75_227#_M1012_g N_A_27_373#_M1012_s VNB NSHORT L=0.15
+ W=0.64 AD=0.112 AS=0.1824 PD=0.99 PS=1.85 NRD=13.116 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75002.2 A=0.096 P=1.58 MULT=1
MM1000 N_A_75_227#_M1000_d N_A_M1000_g N_VGND_M1012_d VNB NSHORT L=0.15 W=0.64
+ AD=0.1072 AS=0.112 PD=0.975 PS=0.99 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.7
+ SB=75001.7 A=0.096 P=1.58 MULT=1
MM1024 N_A_321_77#_M1024_d N_B_M1024_g N_A_75_227#_M1000_d VNB NSHORT L=0.15
+ W=0.64 AD=0.115623 AS=0.1072 PD=1.16528 PS=0.975 NRD=8.436 NRS=10.308 M=1
+ R=4.26667 SA=75001.2 SB=75001.3 A=0.096 P=1.58 MULT=1
MM1003 N_A_27_373#_M1003_d N_A_386_23#_M1003_g N_A_321_77#_M1024_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.111379 AS=0.0758774 PD=0.87566 PS=0.764717 NRD=60.048 NRS=0
+ M=1 R=2.8 SA=75001.7 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1002 N_A_324_373#_M1002_d N_B_M1002_g N_A_27_373#_M1003_d VNB NSHORT L=0.15
+ W=0.64 AD=0.096 AS=0.169721 PD=0.94 PS=1.33434 NRD=1.872 NRS=19.68 M=1
+ R=4.26667 SA=75001.6 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1004 N_A_75_227#_M1004_d N_A_386_23#_M1004_g N_A_324_373#_M1002_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.3467 AS=0.096 PD=2.79 PS=0.94 NRD=91.248 NRS=1.872 M=1
+ R=4.26667 SA=75002.1 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1021 N_VGND_M1021_d N_B_M1021_g N_A_386_23#_M1021_s VNB NSHORT L=0.15 W=0.74
+ AD=0.3368 AS=0.2109 PD=2.67 PS=2.05 NRD=64.884 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1026 N_A_1057_74#_M1026_d N_A_1024_300#_M1026_g N_A_321_77#_M1026_s VNB NSHORT
+ L=0.15 W=0.64 AD=0.1296 AS=0.1824 PD=1.045 PS=1.85 NRD=13.116 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1005 N_A_324_373#_M1005_d N_C_M1005_g N_A_1057_74#_M1026_d VNB NSHORT L=0.15
+ W=0.64 AD=0.192 AS=0.1296 PD=1.88 PS=1.045 NRD=2.808 NRS=10.308 M=1 R=4.26667
+ SA=75000.8 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1013 N_VGND_M1013_d N_C_M1013_g N_A_1024_300#_M1013_s VNB NSHORT L=0.15 W=0.42
+ AD=0.497211 AS=0.1197 PD=1.75603 PS=1.41 NRD=312.852 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75003 A=0.063 P=1.14 MULT=1
MM1001 N_X_M1001_d N_A_1057_74#_M1001_g N_VGND_M1013_d VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.876039 PD=1.02 PS=3.09397 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75001.5 A=0.111 P=1.78 MULT=1
MM1006 N_X_M1001_d N_A_1057_74#_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.9
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1009 N_X_M1009_d N_A_1057_74#_M1009_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.4
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1027 N_X_M1009_d N_A_1057_74#_M1027_g N_VGND_M1027_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.8
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1011 N_VPWR_M1011_d N_A_75_227#_M1011_g N_A_27_373#_M1011_s VPB PHIGHVT L=0.15
+ W=1 AD=0.175 AS=0.295 PD=1.35 PS=2.59 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75002.3 A=0.15 P=2.3 MULT=1
MM1010 N_A_75_227#_M1010_d N_A_M1010_g N_VPWR_M1011_d VPB PHIGHVT L=0.15 W=1
+ AD=0.203696 AS=0.175 PD=1.51087 PS=1.35 NRD=1.9503 NRS=11.8003 M=1 R=6.66667
+ SA=75000.7 SB=75001.8 A=0.15 P=2.3 MULT=1
MM1022 N_A_324_373#_M1022_d N_B_M1022_g N_A_75_227#_M1010_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.229865 AS=0.171104 PD=1.57784 PS=1.26913 NRD=60.9715 NRS=23.837
+ M=1 R=5.6 SA=75001.3 SB=75001.5 A=0.126 P=1.98 MULT=1
MM1007 N_A_27_373#_M1007_d N_A_386_23#_M1007_g N_A_324_373#_M1022_d VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.096 AS=0.175135 PD=0.94 PS=1.20216 NRD=3.0732 NRS=3.0732
+ M=1 R=4.26667 SA=75002 SB=75001.3 A=0.096 P=1.58 MULT=1
MM1015 N_A_321_77#_M1015_d N_B_M1015_g N_A_27_373#_M1007_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.122551 AS=0.096 PD=1.03784 PS=0.94 NRD=21.5321 NRS=3.0732 M=1
+ R=4.26667 SA=75002.4 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1017 N_A_75_227#_M1017_d N_A_386_23#_M1017_g N_A_321_77#_M1015_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.38735 AS=0.160849 PD=2.91 PS=1.36216 NRD=95.2298 NRS=2.3443
+ M=1 R=5.6 SA=75002.3 SB=75000.3 A=0.126 P=1.98 MULT=1
MM1014 N_VPWR_M1014_d N_B_M1014_g N_A_386_23#_M1014_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.3304 PD=2.83 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1025 N_A_1057_74#_M1025_d N_A_1024_300#_M1025_g N_A_324_373#_M1025_s VPB
+ PHIGHVT L=0.15 W=0.84 AD=0.22785 AS=0.2478 PD=1.52 PS=2.27 NRD=50.7078 NRS=0
+ M=1 R=5.6 SA=75000.2 SB=75000.8 A=0.126 P=1.98 MULT=1
MM1020 N_A_321_77#_M1020_d N_C_M1020_g N_A_1057_74#_M1025_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.2478 AS=0.22785 PD=2.27 PS=1.52 NRD=0 NRS=50.7078 M=1 R=5.6
+ SA=75000.8 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1018 N_VPWR_M1018_d N_C_M1018_g N_A_1024_300#_M1018_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.386618 AS=0.1888 PD=1.57818 PS=1.87 NRD=164.672 NRS=3.0732 M=1
+ R=4.26667 SA=75000.2 SB=75002.8 A=0.096 P=1.58 MULT=1
MM1008 N_X_M1008_d N_A_1057_74#_M1008_g N_VPWR_M1018_d VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.676582 PD=1.42 PS=2.76182 NRD=1.7533 NRS=21.5321 M=1 R=7.46667
+ SA=75001.1 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1016 N_X_M1008_d N_A_1057_74#_M1016_g N_VPWR_M1016_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.6 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1019 N_X_M1019_d N_A_1057_74#_M1019_g N_VPWR_M1016_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75002
+ SB=75000.7 A=0.168 P=2.54 MULT=1
MM1023 N_X_M1019_d N_A_1057_74#_M1023_g N_VPWR_M1023_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.5 SB=75000.2 A=0.168 P=2.54 MULT=1
DX28_noxref VNB VPB NWDIODE A=19.4556 P=24.64
c_98 VNB 0 1.89638e-19 $X=0 $Y=0
c_189 VPB 0 1.87651e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_ls__xnor3_4.pxi.spice"
*
.ends
*
*
