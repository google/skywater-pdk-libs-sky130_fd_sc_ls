* File: sky130_fd_sc_ls__o41ai_1.spice
* Created: Wed Sep  2 11:23:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__o41ai_1.pex.spice"
.subckt sky130_fd_sc_ls__o41ai_1  VNB VPB B1 A4 A3 A2 A1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A1	A1
* A2	A2
* A3	A3
* A4	A4
* B1	B1
* VPB	VPB
* VNB	VNB
MM1008 N_A_157_74#_M1008_d N_B1_M1008_g N_Y_M1008_s VNB NSHORT L=0.15 W=0.74
+ AD=0.14615 AS=0.2109 PD=1.135 PS=2.05 NRD=18.648 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75002.3 A=0.111 P=1.78 MULT=1
MM1007 N_VGND_M1007_d N_A4_M1007_g N_A_157_74#_M1008_d VNB NSHORT L=0.15 W=0.74
+ AD=0.16095 AS=0.14615 PD=1.175 PS=1.135 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75000.8 SB=75001.8 A=0.111 P=1.78 MULT=1
MM1002 N_A_157_74#_M1002_d N_A3_M1002_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.16095 PD=1.02 PS=1.175 NRD=0 NRS=13.776 M=1 R=4.93333
+ SA=75001.3 SB=75001.2 A=0.111 P=1.78 MULT=1
MM1006 N_VGND_M1006_d N_A2_M1006_g N_A_157_74#_M1002_d VNB NSHORT L=0.15 W=0.74
+ AD=0.1554 AS=0.1036 PD=1.16 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75001.8
+ SB=75000.8 A=0.111 P=1.78 MULT=1
MM1000 N_A_157_74#_M1000_d N_A1_M1000_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.1554 PD=2.05 PS=1.16 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75002.3
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1001 N_Y_M1001_d N_B1_M1001_g N_VPWR_M1001_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.196 AS=0.5768 PD=1.47 PS=3.27 NRD=10.5395 NRS=7.3284 M=1 R=7.46667
+ SA=75000.4 SB=75002.3 A=0.168 P=2.54 MULT=1
MM1003 A_260_368# N_A4_M1003_g N_Y_M1001_d VPB PHIGHVT L=0.15 W=1.12 AD=0.1904
+ AS=0.196 PD=1.46 PS=1.47 NRD=20.2122 NRS=1.7533 M=1 R=7.46667 SA=75000.9
+ SB=75001.8 A=0.168 P=2.54 MULT=1
MM1009 A_358_368# N_A3_M1009_g A_260_368# VPB PHIGHVT L=0.15 W=1.12 AD=0.2352
+ AS=0.1904 PD=1.54 PS=1.46 NRD=27.2451 NRS=20.2122 M=1 R=7.46667 SA=75001.4
+ SB=75001.4 A=0.168 P=2.54 MULT=1
MM1005 A_472_368# N_A2_M1005_g A_358_368# VPB PHIGHVT L=0.15 W=1.12 AD=0.2352
+ AS=0.2352 PD=1.54 PS=1.54 NRD=27.2451 NRS=27.2451 M=1 R=7.46667 SA=75002
+ SB=75000.8 A=0.168 P=2.54 MULT=1
MM1004 N_VPWR_M1004_d N_A1_M1004_g A_472_368# VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.2352 PD=2.83 PS=1.54 NRD=1.7533 NRS=27.2451 M=1 R=7.46667
+ SA=75002.6 SB=75000.2 A=0.168 P=2.54 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9564 P=11.2
*
.include "sky130_fd_sc_ls__o41ai_1.pxi.spice"
*
.ends
*
*
