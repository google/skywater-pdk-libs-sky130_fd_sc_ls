* NGSPICE file created from sky130_fd_sc_ls__and2_4.ext - technology: sky130A

.subckt sky130_fd_sc_ls__and2_4 A B VGND VNB VPB VPWR X
M1000 X a_83_269# VGND VNB nshort w=740000u l=150000u
+  ad=5.254e+11p pd=4.38e+06u as=8.594e+11p ps=8.14e+06u
M1001 a_83_269# A a_504_119# VNB nshort w=640000u l=150000u
+  ad=2.08e+11p pd=1.93e+06u as=3.872e+11p ps=3.77e+06u
M1002 VGND a_83_269# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_504_119# B VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR A a_83_269# VPB phighvt w=840000u l=150000u
+  ad=1.58705e+12p pd=1.328e+07u as=5.25e+11p ps=4.61e+06u
M1005 VPWR B a_83_269# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_504_119# A a_83_269# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND B a_504_119# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR a_83_269# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=6.944e+11p ps=5.72e+06u
M1009 a_83_269# B VPWR VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 X a_83_269# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 X a_83_269# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR a_83_269# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 X a_83_269# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_83_269# A VPWR VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND a_83_269# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

