* NGSPICE file created from sky130_fd_sc_ls__o32ai_1.ext - technology: sky130A

.subckt sky130_fd_sc_ls__o32ai_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
M1000 VPWR A1 a_456_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=7.056e+11p pd=5.74e+06u as=4.704e+11p ps=3.08e+06u
M1001 VGND A3 a_27_74# VNB nshort w=740000u l=150000u
+  ad=5.439e+11p pd=4.43e+06u as=6.771e+11p ps=6.27e+06u
M1002 a_456_368# A2 a_342_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=4.704e+11p ps=3.08e+06u
M1003 VGND A1 a_27_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_27_74# B2 Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=4.329e+11p ps=2.65e+06u
M1005 a_128_368# B1 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1006 a_342_368# A3 Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=5.6e+11p ps=3.24e+06u
M1007 a_27_74# A2 VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y B1 a_27_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y B2 a_128_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

