* File: sky130_fd_sc_ls__a311o_1.pex.spice
* Created: Wed Sep  2 10:51:29 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__A311O_1%A_89_270# 1 2 3 10 12 13 15 16 17 18 22 26
+ 35 41 42 43
c96 35 0 1.72877e-19 $X=2.405 $Y=1.005
c97 18 0 1.06923e-19 $X=3.245 $Y=1.53
c98 16 0 4.83091e-20 $X=2.24 $Y=1.195
r99 41 42 5.27442 $w=4.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.34 $Y=2.105
+ $X2=3.34 $Y2=1.94
r100 37 38 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.405 $Y=1.195
+ $X2=2.405 $Y2=1.53
r101 35 37 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=2.405 $Y=1.005
+ $X2=2.405 $Y2=1.195
r102 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.645
+ $Y=1.515 $X2=0.645 $Y2=1.515
r103 28 43 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.41 $Y=1.615
+ $X2=3.41 $Y2=1.53
r104 28 42 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=3.41 $Y=1.615
+ $X2=3.41 $Y2=1.94
r105 24 43 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.41 $Y=1.445
+ $X2=3.41 $Y2=1.53
r106 24 26 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=3.41 $Y=1.445
+ $X2=3.41 $Y2=1.105
r107 20 41 1.78139 $w=4.68e-07 $l=7e-08 $layer=LI1_cond $X=3.34 $Y=2.175
+ $X2=3.34 $Y2=2.105
r108 20 22 16.287 $w=4.68e-07 $l=6.4e-07 $layer=LI1_cond $X=3.34 $Y=2.175
+ $X2=3.34 $Y2=2.815
r109 19 38 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.57 $Y=1.53
+ $X2=2.405 $Y2=1.53
r110 18 43 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.245 $Y=1.53
+ $X2=3.41 $Y2=1.53
r111 18 19 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=3.245 $Y=1.53
+ $X2=2.57 $Y2=1.53
r112 17 32 11.4824 $w=3.4e-07 $l=4.20666e-07 $layer=LI1_cond $X=0.945 $Y=1.195
+ $X2=0.712 $Y2=1.515
r113 16 37 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.24 $Y=1.195
+ $X2=2.405 $Y2=1.195
r114 16 17 84.4866 $w=1.68e-07 $l=1.295e-06 $layer=LI1_cond $X=2.24 $Y=1.195
+ $X2=0.945 $Y2=1.195
r115 13 33 38.5818 $w=3.27e-07 $l=2.12238e-07 $layer=POLY_cond $X=0.735 $Y=1.35
+ $X2=0.627 $Y2=1.515
r116 13 15 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.735 $Y=1.35
+ $X2=0.735 $Y2=0.87
r117 10 33 51.1109 $w=3.27e-07 $l=2.92404e-07 $layer=POLY_cond $X=0.535 $Y=1.765
+ $X2=0.627 $Y2=1.515
r118 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.535 $Y=1.765
+ $X2=0.535 $Y2=2.4
r119 3 41 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=3.12
+ $Y=1.96 $X2=3.27 $Y2=2.105
r120 3 22 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=3.12
+ $Y=1.96 $X2=3.27 $Y2=2.815
r121 2 26 182 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_NDIFF $count=1 $X=3.27
+ $Y=0.615 $X2=3.41 $Y2=1.105
r122 1 35 182 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_NDIFF $count=1 $X=2.265
+ $Y=0.615 $X2=2.405 $Y2=1.005
.ends

.subckt PM_SKY130_FD_SC_LS__A311O_1%A3 1 3 6 8
c30 6 0 1.5978e-19 $X=1.245 $Y=0.92
r31 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.2
+ $Y=1.615 $X2=1.2 $Y2=1.615
r32 4 11 38.5916 $w=2.93e-07 $l=1.86145e-07 $layer=POLY_cond $X=1.245 $Y=1.45
+ $X2=1.2 $Y2=1.615
r33 4 6 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.245 $Y=1.45
+ $X2=1.245 $Y2=0.92
r34 1 11 55.8646 $w=2.93e-07 $l=2.77399e-07 $layer=POLY_cond $X=1.215 $Y=1.885
+ $X2=1.2 $Y2=1.615
r35 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.215 $Y=1.885
+ $X2=1.215 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_LS__A311O_1%A2 1 3 6 8
c31 6 0 1.69592e-19 $X=1.72 $Y=0.935
c32 1 0 2.18517e-19 $X=1.665 $Y=1.885
r33 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.74
+ $Y=1.615 $X2=1.74 $Y2=1.615
r34 4 11 38.5916 $w=2.93e-07 $l=1.74714e-07 $layer=POLY_cond $X=1.72 $Y=1.45
+ $X2=1.74 $Y2=1.615
r35 4 6 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=1.72 $Y=1.45 $X2=1.72
+ $Y2=0.935
r36 1 11 55.8646 $w=2.93e-07 $l=3.05205e-07 $layer=POLY_cond $X=1.665 $Y=1.885
+ $X2=1.74 $Y2=1.615
r37 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.665 $Y=1.885
+ $X2=1.665 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_LS__A311O_1%A1 4 5 6 7 9 11 12 16 17 20
c52 17 0 1.83039e-19 $X=2.17 $Y=0.34
c53 16 0 1.46334e-19 $X=2.17 $Y=0.34
c54 6 0 1.06923e-19 $X=2.205 $Y=1.795
r55 16 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.17 $Y=0.34
+ $X2=2.17 $Y2=0.505
r56 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.17
+ $Y=0.34 $X2=2.17 $Y2=0.34
r57 12 17 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=2.17 $Y=0.555
+ $X2=2.17 $Y2=0.34
r58 12 20 2.85155 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=2.17 $Y=0.555
+ $X2=2.005 $Y2=0.555
r59 11 20 16.2845 $w=2.28e-07 $l=3.25e-07 $layer=LI1_cond $X=1.68 $Y=0.555
+ $X2=2.005 $Y2=0.555
r60 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.205 $Y=1.885
+ $X2=2.205 $Y2=2.46
r61 6 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.205 $Y=1.795 $X2=2.205
+ $Y2=1.885
r62 5 10 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.205 $Y=1.42 $X2=2.205
+ $Y2=1.33
r63 5 6 145.766 $w=1.8e-07 $l=3.75e-07 $layer=POLY_cond $X=2.205 $Y=1.42
+ $X2=2.205 $Y2=1.795
r64 4 10 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.19 $Y=0.935
+ $X2=2.19 $Y2=1.33
r65 4 19 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.19 $Y=0.935
+ $X2=2.19 $Y2=0.505
.ends

.subckt PM_SKY130_FD_SC_LS__A311O_1%B1 4 6 7 9 11 12 15
c44 11 0 1.12525e-19 $X=2.645 $Y=1.48
c45 4 0 4.83091e-20 $X=2.62 $Y=0.935
r46 15 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.71 $Y=0.34
+ $X2=2.71 $Y2=0.505
r47 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.71
+ $Y=0.34 $X2=2.71 $Y2=0.34
r48 12 16 9.04483 $w=2.9e-07 $l=2.15e-07 $layer=LI1_cond $X=2.7 $Y=0.555 $X2=2.7
+ $Y2=0.34
r49 10 11 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=2.645 $Y=1.33
+ $X2=2.645 $Y2=1.48
r50 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.655 $Y=1.885
+ $X2=2.655 $Y2=2.46
r51 6 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.655 $Y=1.795 $X2=2.655
+ $Y2=1.885
r52 6 11 122.444 $w=1.8e-07 $l=3.15e-07 $layer=POLY_cond $X=2.655 $Y=1.795
+ $X2=2.655 $Y2=1.48
r53 4 10 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.62 $Y=0.935
+ $X2=2.62 $Y2=1.33
r54 4 18 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.62 $Y=0.935
+ $X2=2.62 $Y2=0.505
.ends

.subckt PM_SKY130_FD_SC_LS__A311O_1%C1 2 3 5 9 12 14 15 18 19
r43 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.55
+ $Y=0.34 $X2=3.55 $Y2=0.34
r44 15 19 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=3.55 $Y=0.555
+ $X2=3.55 $Y2=0.34
r45 14 18 48.9612 $w=3.3e-07 $l=2.8e-07 $layer=POLY_cond $X=3.27 $Y=0.34
+ $X2=3.55 $Y2=0.34
r46 7 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.195 $Y=1.33
+ $X2=3.195 $Y2=1.405
r47 7 9 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.195 $Y=1.33
+ $X2=3.195 $Y2=0.935
r48 6 14 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=3.195 $Y=0.505
+ $X2=3.27 $Y2=0.34
r49 6 9 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.195 $Y=0.505
+ $X2=3.195 $Y2=0.935
r50 3 5 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.045 $Y=1.885
+ $X2=3.045 $Y2=2.46
r51 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.045 $Y=1.795 $X2=3.045
+ $Y2=1.885
r52 1 12 76.9149 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=3.045 $Y=1.405
+ $X2=3.195 $Y2=1.405
r53 1 2 122.444 $w=1.8e-07 $l=3.15e-07 $layer=POLY_cond $X=3.045 $Y=1.48
+ $X2=3.045 $Y2=1.795
.ends

.subckt PM_SKY130_FD_SC_LS__A311O_1%X 1 2 9 11 17 18 19 26 35
r21 24 26 0.329269 $w=3.48e-07 $l=1e-08 $layer=LI1_cond $X=0.3 $Y=2.025 $X2=0.3
+ $Y2=2.035
r22 18 19 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.3 $Y=2.405 $X2=0.3
+ $Y2=2.775
r23 17 24 1.25122 $w=3.48e-07 $l=3.8e-08 $layer=LI1_cond $X=0.3 $Y=1.987 $X2=0.3
+ $Y2=2.025
r24 17 35 7.56653 $w=3.48e-07 $l=1.37e-07 $layer=LI1_cond $X=0.3 $Y=1.987
+ $X2=0.3 $Y2=1.85
r25 17 18 10.9647 $w=3.48e-07 $l=3.33e-07 $layer=LI1_cond $X=0.3 $Y=2.072
+ $X2=0.3 $Y2=2.405
r26 17 26 1.2183 $w=3.48e-07 $l=3.7e-08 $layer=LI1_cond $X=0.3 $Y=2.072 $X2=0.3
+ $Y2=2.035
r27 9 13 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.48 $Y=1.095 $X2=0.21
+ $Y2=1.095
r28 9 11 16.8257 $w=2.48e-07 $l=3.65e-07 $layer=LI1_cond $X=0.48 $Y=1.01
+ $X2=0.48 $Y2=0.645
r29 7 13 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.21 $Y=1.18 $X2=0.21
+ $Y2=1.095
r30 7 35 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.21 $Y=1.18 $X2=0.21
+ $Y2=1.85
r31 2 17 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.185
+ $Y=1.84 $X2=0.31 $Y2=2.015
r32 2 19 400 $w=1.7e-07 $l=1.03562e-06 $layer=licon1_PDIFF $count=1 $X=0.185
+ $Y=1.84 $X2=0.31 $Y2=2.815
r33 1 11 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.395
+ $Y=0.5 $X2=0.52 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_LS__A311O_1%VPWR 1 2 11 17 20 21 22 32 33 36
r41 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r42 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r43 30 33 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.6 $Y2=3.33
r44 29 32 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=3.6 $Y2=3.33
r45 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r46 27 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r47 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r48 24 36 10.7288 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=1.105 $Y=3.33
+ $X2=0.875 $Y2=3.33
r49 24 26 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=1.105 $Y=3.33
+ $X2=1.68 $Y2=3.33
r50 22 30 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.16 $Y2=3.33
r51 22 27 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r52 20 26 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=1.805 $Y=3.33
+ $X2=1.68 $Y2=3.33
r53 20 21 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=1.805 $Y=3.33
+ $X2=1.95 $Y2=3.33
r54 19 29 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=2.095 $Y=3.33
+ $X2=2.16 $Y2=3.33
r55 19 21 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=2.095 $Y=3.33
+ $X2=1.95 $Y2=3.33
r56 15 21 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.95 $Y=3.245
+ $X2=1.95 $Y2=3.33
r57 15 17 31.3941 $w=2.88e-07 $l=7.9e-07 $layer=LI1_cond $X=1.95 $Y=3.245
+ $X2=1.95 $Y2=2.455
r58 11 14 18.2012 $w=4.58e-07 $l=7e-07 $layer=LI1_cond $X=0.875 $Y=2.115
+ $X2=0.875 $Y2=2.815
r59 9 36 1.85547 $w=4.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.875 $Y=3.245
+ $X2=0.875 $Y2=3.33
r60 9 14 11.1807 $w=4.58e-07 $l=4.3e-07 $layer=LI1_cond $X=0.875 $Y=3.245
+ $X2=0.875 $Y2=2.815
r61 2 17 300 $w=1.7e-07 $l=5.73738e-07 $layer=licon1_PDIFF $count=2 $X=1.74
+ $Y=1.96 $X2=1.91 $Y2=2.455
r62 1 14 400 $w=1.7e-07 $l=1.09955e-06 $layer=licon1_PDIFF $count=1 $X=0.61
+ $Y=1.84 $X2=0.875 $Y2=2.815
r63 1 11 400 $w=1.7e-07 $l=3.85357e-07 $layer=licon1_PDIFF $count=1 $X=0.61
+ $Y=1.84 $X2=0.875 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_LS__A311O_1%A_258_392# 1 2 7 9 11 13 15
c39 13 0 1.58165e-19 $X=2.43 $Y=2.12
r40 13 20 2.68829 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=2.43 $Y=2.12 $X2=2.43
+ $Y2=2.03
r41 13 15 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=2.43 $Y=2.12
+ $X2=2.43 $Y2=2.815
r42 12 18 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.605 $Y=2.035
+ $X2=1.44 $Y2=2.035
r43 11 20 5.07788 $w=1.7e-07 $l=1.67481e-07 $layer=LI1_cond $X=2.265 $Y=2.035
+ $X2=2.43 $Y2=2.03
r44 11 12 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=2.265 $Y=2.035
+ $X2=1.605 $Y2=2.035
r45 7 18 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.44 $Y=2.12 $X2=1.44
+ $Y2=2.035
r46 7 9 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=1.44 $Y=2.12 $X2=1.44
+ $Y2=2.815
r47 2 20 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.28
+ $Y=1.96 $X2=2.43 $Y2=2.105
r48 2 15 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=2.28
+ $Y=1.96 $X2=2.43 $Y2=2.815
r49 1 18 400 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=1 $X=1.29
+ $Y=1.96 $X2=1.44 $Y2=2.115
r50 1 9 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=1.29
+ $Y=1.96 $X2=1.44 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_LS__A311O_1%VGND 1 2 9 12 14 15 18 24 30 31 34
r48 34 35 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r49 31 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r50 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r51 28 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.215 $Y=0 $X2=3.13
+ $Y2=0
r52 28 30 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=3.215 $Y=0 $X2=3.6
+ $Y2=0
r53 26 27 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r54 24 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.045 $Y=0 $X2=3.13
+ $Y2=0
r55 24 26 120.369 $w=1.68e-07 $l=1.845e-06 $layer=LI1_cond $X=3.045 $Y=0 $X2=1.2
+ $Y2=0
r56 22 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r57 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r58 18 35 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.92 $Y=0 $X2=3.12
+ $Y2=0
r59 18 27 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.2
+ $Y2=0
r60 14 21 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=0.785 $Y=0 $X2=0.72
+ $Y2=0
r61 14 15 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.785 $Y=0 $X2=0.95
+ $Y2=0
r62 13 26 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.115 $Y=0 $X2=1.2
+ $Y2=0
r63 13 15 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.115 $Y=0 $X2=0.95
+ $Y2=0
r64 12 17 15.8187 $w=3.2e-07 $l=4.12414e-07 $layer=LI1_cond $X=3.13 $Y=0.675
+ $X2=2.982 $Y2=1.02
r65 11 34 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.13 $Y=0.085
+ $X2=3.13 $Y2=0
r66 11 12 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=3.13 $Y=0.085
+ $X2=3.13 $Y2=0.675
r67 7 15 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.95 $Y=0.085 $X2=0.95
+ $Y2=0
r68 7 9 24.0965 $w=3.28e-07 $l=6.9e-07 $layer=LI1_cond $X=0.95 $Y=0.085 $X2=0.95
+ $Y2=0.775
r69 2 17 182 $w=1.7e-07 $l=5.03115e-07 $layer=licon1_NDIFF $count=1 $X=2.695
+ $Y=0.615 $X2=2.915 $Y2=1.02
r70 1 9 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=0.81
+ $Y=0.5 $X2=0.95 $Y2=0.775
.ends

