* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__o311a_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
M1000 a_83_244# A3 a_1034_392# VPB phighvt w=1e+06u l=150000u
+  ad=1.09e+12p pd=8.18e+06u as=1.075e+12p ps=8.15e+06u
M1001 a_1338_392# A2 a_1034_392# VPB phighvt w=1e+06u l=150000u
+  ad=7.4e+11p pd=5.48e+06u as=0p ps=0u
M1002 a_564_78# A1 VGND VNB nshort w=640000u l=150000u
+  ad=1.02922e+12p pd=9.63e+06u as=1.5521e+12p ps=1.276e+07u
M1003 a_651_78# B1 a_564_78# VNB nshort w=640000u l=150000u
+  ad=6.88e+11p pd=4.71e+06u as=0p ps=0u
M1004 X a_83_244# VGND VNB nshort w=740000u l=150000u
+  ad=4.662e+11p pd=4.22e+06u as=0p ps=0u
M1005 VGND a_83_244# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_564_78# A2 VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_83_244# C1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.4192e+12p ps=1.734e+07u
M1008 a_83_244# C1 a_651_78# VNB nshort w=640000u l=150000u
+  ad=3.4395e+11p pd=2.59e+06u as=0p ps=0u
M1009 X a_83_244# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=8.792e+11p pd=6.05e+06u as=0p ps=0u
M1010 VPWR a_83_244# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR B1 a_83_244# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_564_78# A3 VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR a_83_244# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND A2 a_564_78# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR C1 a_83_244# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR A1 a_1338_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_651_78# C1 a_83_244# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND A3 a_564_78# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 X a_83_244# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_1034_392# A2 a_1338_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND a_83_244# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_83_244# B1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_1034_392# A3 a_83_244# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_564_78# B1 a_651_78# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VGND A1 a_564_78# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 X a_83_244# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_1338_392# A1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
