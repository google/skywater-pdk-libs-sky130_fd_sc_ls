# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ls__nand4bb_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ls__nand4bb_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.720000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A_N
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.435000 1.300000 0.835000 1.780000 ;
    END
  END A_N
  PIN B_N
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005000 1.180000 1.335000 1.510000 ;
    END
  END B_N
  PIN C
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445000 1.350000 5.385000 1.780000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.625000 1.350000 6.595000 1.680000 ;
        RECT 6.365000 1.680000 6.595000 1.780000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  1.614500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.345000 0.670000 2.855000 0.840000 ;
        RECT 2.345000 1.820000 2.675000 1.850000 ;
        RECT 2.345000 1.850000 4.195000 1.950000 ;
        RECT 2.345000 1.950000 6.105000 2.020000 ;
        RECT 2.345000 2.020000 2.675000 2.980000 ;
        RECT 2.685000 0.840000 2.855000 1.090000 ;
        RECT 2.685000 1.090000 4.195000 1.260000 ;
        RECT 3.345000 2.020000 6.105000 2.120000 ;
        RECT 3.345000 2.120000 3.675000 2.980000 ;
        RECT 3.965000 1.260000 4.195000 1.850000 ;
        RECT 4.775000 2.120000 5.105000 2.980000 ;
        RECT 5.775000 1.850000 6.105000 1.950000 ;
        RECT 5.775000 2.120000 6.105000 2.980000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.720000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 6.720000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.720000 0.085000 ;
      RECT 0.000000  3.245000 6.720000 3.415000 ;
      RECT 0.095000  0.350000 0.460000 1.030000 ;
      RECT 0.095000  1.030000 0.265000 1.950000 ;
      RECT 0.095000  1.950000 0.445000 2.240000 ;
      RECT 0.095000  2.240000 2.175000 2.410000 ;
      RECT 0.095000  2.410000 0.445000 2.860000 ;
      RECT 0.630000  0.085000 0.960000 1.010000 ;
      RECT 0.650000  2.580000 0.980000 3.245000 ;
      RECT 1.130000  0.350000 1.675000 1.010000 ;
      RECT 1.185000  1.820000 1.675000 2.070000 ;
      RECT 1.505000  1.010000 2.515000 1.180000 ;
      RECT 1.505000  1.180000 1.675000 1.820000 ;
      RECT 1.845000  0.330000 3.195000 0.500000 ;
      RECT 1.845000  0.500000 2.175000 0.840000 ;
      RECT 1.845000  1.350000 2.175000 2.240000 ;
      RECT 1.845000  2.580000 2.175000 3.245000 ;
      RECT 2.345000  1.180000 2.515000 1.430000 ;
      RECT 2.345000  1.430000 3.795000 1.600000 ;
      RECT 2.845000  2.190000 3.175000 3.245000 ;
      RECT 3.025000  0.500000 3.195000 0.750000 ;
      RECT 3.025000  0.750000 4.180000 0.920000 ;
      RECT 3.125000  1.600000 3.795000 1.680000 ;
      RECT 3.365000  0.255000 5.240000 0.425000 ;
      RECT 3.365000  0.425000 3.695000 0.580000 ;
      RECT 3.845000  2.290000 4.605000 3.245000 ;
      RECT 4.410000  0.620000 4.740000 1.010000 ;
      RECT 4.410000  1.010000 6.600000 1.180000 ;
      RECT 4.910000  0.425000 5.240000 0.815000 ;
      RECT 5.275000  2.290000 5.605000 3.245000 ;
      RECT 5.420000  0.350000 5.670000 1.010000 ;
      RECT 5.840000  0.085000 6.170000 0.815000 ;
      RECT 6.275000  1.950000 6.605000 3.245000 ;
      RECT 6.350000  0.350000 6.600000 1.010000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
  END
END sky130_fd_sc_ls__nand4bb_2
END LIBRARY
