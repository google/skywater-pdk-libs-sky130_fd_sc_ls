* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__maj3_4 A B C VGND VNB VPB VPWR X
X0 a_114_125# A VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X1 a_219_392# B a_501_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 VGND A a_114_125# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X3 X a_219_392# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X4 VGND A a_906_78# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X5 a_219_392# C a_905_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 X a_219_392# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X7 a_219_392# B a_119_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 a_501_392# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 VGND C a_504_125# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X10 a_504_125# C VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X11 VPWR C a_501_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 VPWR A a_905_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 X a_219_392# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X14 a_905_392# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 a_114_125# B a_219_392# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X16 VGND a_219_392# X VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X17 VPWR a_219_392# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X18 a_219_392# B a_504_125# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X19 a_219_392# C a_906_78# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X20 VPWR a_219_392# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X21 VPWR A a_119_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X22 a_119_392# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X23 a_906_78# C a_219_392# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X24 a_501_392# B a_219_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X25 a_219_392# B a_114_125# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X26 VGND a_219_392# X VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X27 X a_219_392# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X28 a_119_392# B a_219_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X29 a_504_125# B a_219_392# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X30 a_905_392# C a_219_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X31 a_906_78# A VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
.ends
