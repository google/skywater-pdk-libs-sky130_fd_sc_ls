* File: sky130_fd_sc_ls__einvp_4.spice
* Created: Wed Sep  2 11:07:18 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__einvp_4.pex.spice"
.subckt sky130_fd_sc_ls__einvp_4  VNB VPB A TE Z VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Z	Z
* TE	TE
* A	A
* VPB	VPB
* VNB	VNB
MM1002 N_A_27_74#_M1002_d N_A_M1002_g N_Z_M1002_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.1295 PD=2.05 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75000.2
+ SB=75003.8 A=0.111 P=1.78 MULT=1
MM1005 N_A_27_74#_M1005_d N_A_M1005_g N_Z_M1002_s VNB NSHORT L=0.15 W=0.74
+ AD=0.13875 AS=0.1295 PD=1.115 PS=1.09 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.7
+ SB=75003.3 A=0.111 P=1.78 MULT=1
MM1014 N_A_27_74#_M1005_d N_A_M1014_g N_Z_M1014_s VNB NSHORT L=0.15 W=0.74
+ AD=0.13875 AS=0.12025 PD=1.115 PS=1.065 NRD=4.044 NRS=7.296 M=1 R=4.93333
+ SA=75001.2 SB=75002.8 A=0.111 P=1.78 MULT=1
MM1016 N_A_27_74#_M1016_d N_A_M1016_g N_Z_M1014_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1295 AS=0.12025 PD=1.09 PS=1.065 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75001.7
+ SB=75002.3 A=0.111 P=1.78 MULT=1
MM1001 N_VGND_M1001_d N_TE_M1001_g N_A_27_74#_M1016_d VNB NSHORT L=0.15 W=0.74
+ AD=0.1554 AS=0.1295 PD=1.16 PS=1.09 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75002.2
+ SB=75001.8 A=0.111 P=1.78 MULT=1
MM1006 N_VGND_M1001_d N_TE_M1006_g N_A_27_74#_M1006_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1554 AS=0.1036 PD=1.16 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75002.8
+ SB=75001.2 A=0.111 P=1.78 MULT=1
MM1010 N_VGND_M1010_d N_TE_M1010_g N_A_27_74#_M1006_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1554 AS=0.1036 PD=1.16 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75003.2
+ SB=75000.8 A=0.111 P=1.78 MULT=1
MM1017 N_VGND_M1010_d N_TE_M1017_g N_A_27_74#_M1017_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1554 AS=0.2109 PD=1.16 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75003.8
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1015 N_VGND_M1015_d N_TE_M1015_g N_A_473_323#_M1015_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2627 AS=0.2109 PD=2.19 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1000 N_A_27_368#_M1000_d N_A_M1000_g N_Z_M1000_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.336 AS=0.1932 PD=2.84 PS=1.465 NRD=2.6201 NRS=9.6727 M=1 R=7.46667
+ SA=75000.2 SB=75003.6 A=0.168 P=2.54 MULT=1
MM1008 N_A_27_368#_M1008_d N_A_M1008_g N_Z_M1000_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.196 AS=0.1932 PD=1.47 PS=1.465 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75003.1 A=0.168 P=2.54 MULT=1
MM1009 N_A_27_368#_M1008_d N_A_M1009_g N_Z_M1009_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.196 AS=0.168 PD=1.47 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.2 SB=75002.6 A=0.168 P=2.54 MULT=1
MM1013 N_A_27_368#_M1013_d N_A_M1013_g N_Z_M1009_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.196 AS=0.168 PD=1.47 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75001.7 SB=75002.1 A=0.168 P=2.54 MULT=1
MM1003 N_VPWR_M1003_d N_A_473_323#_M1003_g N_A_27_368#_M1013_d VPB PHIGHVT
+ L=0.15 W=1.12 AD=0.196 AS=0.196 PD=1.47 PS=1.47 NRD=10.5395 NRS=1.7533 M=1
+ R=7.46667 SA=75002.2 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1007 N_VPWR_M1003_d N_A_473_323#_M1007_g N_A_27_368#_M1007_s VPB PHIGHVT
+ L=0.15 W=1.12 AD=0.196 AS=0.168 PD=1.47 PS=1.42 NRD=1.7533 NRS=1.7533 M=1
+ R=7.46667 SA=75002.7 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1011 N_VPWR_M1011_d N_A_473_323#_M1011_g N_A_27_368#_M1007_s VPB PHIGHVT
+ L=0.15 W=1.12 AD=0.1736 AS=0.168 PD=1.43 PS=1.42 NRD=2.6201 NRS=1.7533 M=1
+ R=7.46667 SA=75003.1 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1012 N_VPWR_M1011_d N_A_473_323#_M1012_g N_A_27_368#_M1012_s VPB PHIGHVT
+ L=0.15 W=1.12 AD=0.1736 AS=0.3304 PD=1.43 PS=2.83 NRD=2.6201 NRS=1.7533 M=1
+ R=7.46667 SA=75003.6 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1004 N_VPWR_M1004_d N_TE_M1004_g N_A_473_323#_M1004_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.3304 AS=0.3304 PD=2.83 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.2 A=0.168 P=2.54 MULT=1
DX18_noxref VNB VPB NWDIODE A=11.4204 P=16
*
.include "sky130_fd_sc_ls__einvp_4.pxi.spice"
*
.ends
*
*
