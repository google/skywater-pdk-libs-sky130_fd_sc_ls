# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ls__and4bb_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_ls__and4bb_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.120000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A_N
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005000 1.450000 1.335000 1.780000 ;
    END
  END A_N
  PIN B_N
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.450000 0.835000 1.780000 ;
    END
  END B_N
  PIN C
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.965000 1.450000 6.115000 1.780000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.365000 1.350000 6.875000 1.780000 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  1.116000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.240000 0.350000 7.570000 0.980000 ;
        RECT 7.240000 0.980000 8.995000 1.150000 ;
        RECT 7.405000 1.820000 8.995000 2.150000 ;
        RECT 7.405000 2.150000 7.575000 2.980000 ;
        RECT 8.240000 0.770000 8.995000 0.980000 ;
        RECT 8.765000 1.150000 8.995000 1.820000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 9.120000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 9.120000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.120000 0.085000 ;
      RECT 0.000000  3.245000 9.120000 3.415000 ;
      RECT 0.115000  0.350000 0.365000 1.110000 ;
      RECT 0.115000  1.110000 1.870000 1.280000 ;
      RECT 0.115000  1.950000 1.675000 2.120000 ;
      RECT 0.115000  2.120000 0.445000 2.980000 ;
      RECT 0.545000  0.085000 0.875000 0.940000 ;
      RECT 0.615000  2.290000 0.945000 3.245000 ;
      RECT 1.045000  0.255000 1.690000 0.585000 ;
      RECT 1.045000  0.585000 1.530000 0.940000 ;
      RECT 1.115000  2.290000 2.260000 2.460000 ;
      RECT 1.115000  2.460000 1.445000 2.980000 ;
      RECT 1.505000  1.280000 1.675000 1.950000 ;
      RECT 1.700000  0.755000 2.030000 0.925000 ;
      RECT 1.700000  0.925000 1.870000 1.110000 ;
      RECT 1.860000  0.255000 3.605000 0.585000 ;
      RECT 1.860000  0.585000 2.030000 0.755000 ;
      RECT 1.890000  2.630000 2.225000 3.245000 ;
      RECT 1.930000  1.450000 2.260000 2.290000 ;
      RECT 2.040000  1.095000 2.370000 1.280000 ;
      RECT 2.200000  0.755000 3.220000 0.925000 ;
      RECT 2.200000  0.925000 2.370000 1.095000 ;
      RECT 2.430000  1.595000 4.795000 1.765000 ;
      RECT 2.430000  1.765000 2.760000 2.960000 ;
      RECT 2.540000  1.095000 2.870000 1.360000 ;
      RECT 2.540000  1.360000 2.760000 1.595000 ;
      RECT 2.965000  1.935000 3.295000 3.245000 ;
      RECT 3.050000  0.925000 3.220000 1.255000 ;
      RECT 3.050000  1.255000 4.160000 1.425000 ;
      RECT 3.400000  0.755000 5.220000 0.925000 ;
      RECT 3.400000  0.925000 3.650000 1.085000 ;
      RECT 3.465000  1.765000 3.795000 2.960000 ;
      RECT 3.830000  1.095000 4.160000 1.255000 ;
      RECT 3.965000  1.935000 4.295000 3.245000 ;
      RECT 4.390000  1.095000 4.720000 1.110000 ;
      RECT 4.390000  1.110000 6.560000 1.180000 ;
      RECT 4.390000  1.180000 5.650000 1.280000 ;
      RECT 4.390000  1.280000 4.720000 1.345000 ;
      RECT 4.465000  1.765000 4.795000 1.950000 ;
      RECT 4.465000  1.950000 7.235000 2.120000 ;
      RECT 4.465000  2.120000 4.795000 2.960000 ;
      RECT 4.890000  0.665000 5.220000 0.755000 ;
      RECT 4.890000  0.925000 5.220000 0.940000 ;
      RECT 4.965000  2.290000 6.165000 3.245000 ;
      RECT 5.400000  0.665000 5.650000 1.010000 ;
      RECT 5.400000  1.010000 6.560000 1.110000 ;
      RECT 5.880000  0.085000 6.130000 0.840000 ;
      RECT 6.310000  0.450000 6.560000 1.010000 ;
      RECT 6.335000  2.120000 6.665000 2.860000 ;
      RECT 6.740000  0.085000 7.070000 1.130000 ;
      RECT 6.875000  2.290000 7.205000 3.245000 ;
      RECT 7.065000  1.320000 8.565000 1.650000 ;
      RECT 7.065000  1.650000 7.235000 1.950000 ;
      RECT 7.740000  0.085000 8.070000 0.810000 ;
      RECT 7.775000  2.320000 8.105000 3.245000 ;
      RECT 8.670000  0.085000 9.005000 0.600000 ;
      RECT 8.675000  2.320000 9.005000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
  END
END sky130_fd_sc_ls__and4bb_4
END LIBRARY
