* File: sky130_fd_sc_ls__a222oi_1.pxi.spice
* Created: Fri Aug 28 12:54:21 2020
* 
x_PM_SKY130_FD_SC_LS__A222OI_1%C1 N_C1_c_70_n N_C1_c_75_n N_C1_M1009_g
+ N_C1_M1002_g C1 N_C1_c_71_n N_C1_c_72_n N_C1_c_73_n
+ PM_SKY130_FD_SC_LS__A222OI_1%C1
x_PM_SKY130_FD_SC_LS__A222OI_1%C2 N_C2_c_102_n N_C2_M1011_g N_C2_c_103_n
+ N_C2_M1008_g C2 C2 PM_SKY130_FD_SC_LS__A222OI_1%C2
x_PM_SKY130_FD_SC_LS__A222OI_1%B2 N_B2_c_140_n N_B2_M1001_g N_B2_M1000_g
+ N_B2_c_136_n N_B2_c_137_n B2 B2 N_B2_c_139_n PM_SKY130_FD_SC_LS__A222OI_1%B2
x_PM_SKY130_FD_SC_LS__A222OI_1%B1 N_B1_M1003_g N_B1_c_178_n N_B1_M1004_g
+ N_B1_c_174_n N_B1_c_175_n B1 B1 N_B1_c_177_n PM_SKY130_FD_SC_LS__A222OI_1%B1
x_PM_SKY130_FD_SC_LS__A222OI_1%A1 N_A1_c_212_n N_A1_c_217_n N_A1_M1007_g
+ N_A1_M1005_g A1 A1 N_A1_c_213_n N_A1_c_214_n N_A1_c_215_n
+ PM_SKY130_FD_SC_LS__A222OI_1%A1
x_PM_SKY130_FD_SC_LS__A222OI_1%A2 N_A2_M1006_g N_A2_c_250_n N_A2_c_254_n
+ N_A2_M1010_g A2 A2 N_A2_c_252_n PM_SKY130_FD_SC_LS__A222OI_1%A2
x_PM_SKY130_FD_SC_LS__A222OI_1%Y N_Y_M1002_s N_Y_M1003_d N_Y_M1009_s N_Y_M1008_d
+ N_Y_c_283_n N_Y_c_284_n N_Y_c_278_n N_Y_c_293_n N_Y_c_295_n N_Y_c_279_n
+ N_Y_c_285_n N_Y_c_286_n N_Y_c_280_n N_Y_c_318_n Y Y Y Y
+ PM_SKY130_FD_SC_LS__A222OI_1%Y
x_PM_SKY130_FD_SC_LS__A222OI_1%A_116_392# N_A_116_392#_M1009_d
+ N_A_116_392#_M1001_d N_A_116_392#_c_361_n N_A_116_392#_c_358_n
+ N_A_116_392#_c_359_n N_A_116_392#_c_366_n
+ PM_SKY130_FD_SC_LS__A222OI_1%A_116_392#
x_PM_SKY130_FD_SC_LS__A222OI_1%A_369_392# N_A_369_392#_M1001_s
+ N_A_369_392#_M1004_d N_A_369_392#_M1010_d N_A_369_392#_c_388_n
+ N_A_369_392#_c_383_n N_A_369_392#_c_401_n N_A_369_392#_c_384_n
+ N_A_369_392#_c_385_n N_A_369_392#_c_386_n N_A_369_392#_c_387_n
+ PM_SKY130_FD_SC_LS__A222OI_1%A_369_392#
x_PM_SKY130_FD_SC_LS__A222OI_1%VPWR N_VPWR_M1007_d N_VPWR_c_427_n N_VPWR_c_428_n
+ N_VPWR_c_429_n VPWR N_VPWR_c_430_n N_VPWR_c_426_n
+ PM_SKY130_FD_SC_LS__A222OI_1%VPWR
x_PM_SKY130_FD_SC_LS__A222OI_1%VGND N_VGND_M1011_d N_VGND_M1006_d N_VGND_c_462_n
+ N_VGND_c_463_n VGND N_VGND_c_464_n N_VGND_c_465_n N_VGND_c_466_n
+ N_VGND_c_467_n PM_SKY130_FD_SC_LS__A222OI_1%VGND
cc_1 VNB N_C1_c_70_n 0.0124041f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.795
cc_2 VNB N_C1_c_71_n 0.0334751f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.285
cc_3 VNB N_C1_c_72_n 0.0274553f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.285
cc_4 VNB N_C1_c_73_n 0.023864f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.12
cc_5 VNB N_C2_c_102_n 0.0197172f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.45
cc_6 VNB N_C2_c_103_n 0.0628469f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.46
cc_7 VNB C2 0.0030793f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.69
cc_8 VNB N_B2_c_136_n 0.0194107f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.69
cc_9 VNB N_B2_c_137_n 0.0308246f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_10 VNB B2 0.00168047f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_B2_c_139_n 0.0187447f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.45
cc_12 VNB N_B1_c_174_n 0.0196919f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.69
cc_13 VNB N_B1_c_175_n 0.0242061f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_14 VNB B1 0.00551108f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_B1_c_177_n 0.0158166f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.45
cc_16 VNB N_A1_c_212_n 0.0243798f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.795
cc_17 VNB N_A1_c_213_n 0.018178f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.12
cc_18 VNB N_A1_c_214_n 0.0152451f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.45
cc_19 VNB N_A1_c_215_n 0.0199469f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.455
cc_20 VNB N_A2_M1006_g 0.0265625f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.885
cc_21 VNB N_A2_c_250_n 0.00970738f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.12
cc_22 VNB A2 0.0100538f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A2_c_252_n 0.0590063f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_Y_c_278_n 0.0189692f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.455
cc_25 VNB N_Y_c_279_n 0.0072208f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_Y_c_280_n 0.00618121f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB Y 0.0158532f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB Y 8.17974e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VPWR_c_426_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_462_n 0.0128247f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.69
cc_31 VNB N_VGND_c_463_n 0.0321458f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_32 VNB N_VGND_c_464_n 0.0459918f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_465_n 0.0299712f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_466_n 0.0355947f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_467_n 0.253868f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VPB N_C1_c_70_n 0.00799152f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.795
cc_37 VPB N_C1_c_75_n 0.0304076f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.885
cc_38 VPB N_C1_c_72_n 0.00936426f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.285
cc_39 VPB N_C2_c_103_n 0.0461427f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.46
cc_40 VPB C2 0.0020523f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=0.69
cc_41 VPB N_B2_c_140_n 0.0179951f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.45
cc_42 VPB N_B2_c_137_n 0.0222178f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_43 VPB B2 0.00139606f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_44 VPB N_B1_c_178_n 0.016408f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.46
cc_45 VPB N_B1_c_175_n 0.019203f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_46 VPB B1 0.00245553f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB N_A1_c_212_n 0.0208295f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.795
cc_48 VPB N_A1_c_217_n 0.0175131f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.885
cc_49 VPB N_A1_c_214_n 0.00483286f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.45
cc_50 VPB N_A2_c_250_n 0.00893127f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.12
cc_51 VPB N_A2_c_254_n 0.0313345f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=0.69
cc_52 VPB A2 0.00812361f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_Y_c_283_n 0.00956607f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.285
cc_54 VPB N_Y_c_284_n 0.0350163f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.45
cc_55 VPB N_Y_c_285_n 0.00527344f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_Y_c_286_n 0.0220994f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB Y 0.0084656f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_A_116_392#_c_358_n 0.0220555f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.285
cc_59 VPB N_A_116_392#_c_359_n 0.00395905f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.285
cc_60 VPB N_A_369_392#_c_383_n 0.00289633f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.455
cc_61 VPB N_A_369_392#_c_384_n 0.00892105f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_A_369_392#_c_385_n 0.0350163f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_A_369_392#_c_386_n 0.0147117f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_A_369_392#_c_387_n 0.00867752f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_427_n 0.0097742f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.12
cc_66 VPB N_VPWR_c_428_n 0.083223f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_67 VPB N_VPWR_c_429_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_430_n 0.0207426f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_426_n 0.0737932f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 N_C1_c_73_n N_C2_c_102_n 0.041753f $X=0.43 $Y=1.12 $X2=-0.19 $Y2=-0.245
cc_71 N_C1_c_70_n N_C2_c_103_n 0.00437412f $X=0.505 $Y=1.795 $X2=0 $Y2=0
cc_72 N_C1_c_75_n N_C2_c_103_n 0.025963f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_73 N_C1_c_71_n N_C2_c_103_n 0.041753f $X=0.43 $Y=1.285 $X2=0 $Y2=0
cc_74 N_C1_c_72_n N_C2_c_103_n 0.00286882f $X=0.43 $Y=1.285 $X2=0 $Y2=0
cc_75 N_C1_c_71_n C2 6.88337e-19 $X=0.43 $Y=1.285 $X2=0 $Y2=0
cc_76 N_C1_c_72_n C2 0.0264482f $X=0.43 $Y=1.285 $X2=0 $Y2=0
cc_77 N_C1_c_75_n N_Y_c_283_n 4.27055e-19 $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_78 N_C1_c_71_n N_Y_c_283_n 5.12337e-19 $X=0.43 $Y=1.285 $X2=0 $Y2=0
cc_79 N_C1_c_72_n N_Y_c_283_n 0.0264916f $X=0.43 $Y=1.285 $X2=0 $Y2=0
cc_80 N_C1_c_75_n N_Y_c_284_n 0.0102668f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_81 N_C1_c_73_n N_Y_c_278_n 0.00793201f $X=0.43 $Y=1.12 $X2=0 $Y2=0
cc_82 N_C1_c_75_n N_Y_c_293_n 0.01222f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_83 N_C1_c_72_n N_Y_c_293_n 0.010813f $X=0.43 $Y=1.285 $X2=0 $Y2=0
cc_84 N_C1_c_72_n N_Y_c_295_n 0.00942884f $X=0.43 $Y=1.285 $X2=0 $Y2=0
cc_85 N_C1_c_73_n N_Y_c_295_n 0.00806212f $X=0.43 $Y=1.12 $X2=0 $Y2=0
cc_86 N_C1_c_71_n N_Y_c_279_n 0.00412259f $X=0.43 $Y=1.285 $X2=0 $Y2=0
cc_87 N_C1_c_72_n N_Y_c_279_n 0.026382f $X=0.43 $Y=1.285 $X2=0 $Y2=0
cc_88 N_C1_c_73_n N_Y_c_279_n 7.15802e-19 $X=0.43 $Y=1.12 $X2=0 $Y2=0
cc_89 N_C1_c_75_n N_A_116_392#_c_359_n 0.00364659f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_90 N_C1_c_75_n N_VPWR_c_428_n 0.00445602f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_91 N_C1_c_75_n N_VPWR_c_426_n 0.0086236f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_92 N_C1_c_73_n N_VGND_c_465_n 0.00434272f $X=0.43 $Y=1.12 $X2=0 $Y2=0
cc_93 N_C1_c_73_n N_VGND_c_466_n 0.00126064f $X=0.43 $Y=1.12 $X2=0 $Y2=0
cc_94 N_C1_c_73_n N_VGND_c_467_n 0.00437003f $X=0.43 $Y=1.12 $X2=0 $Y2=0
cc_95 N_C2_c_103_n N_B2_c_139_n 0.00733596f $X=1.005 $Y=1.885 $X2=0 $Y2=0
cc_96 N_C2_c_103_n N_Y_c_284_n 6.19367e-19 $X=1.005 $Y=1.885 $X2=0 $Y2=0
cc_97 N_C2_c_102_n N_Y_c_278_n 0.00159871f $X=0.91 $Y=1.12 $X2=0 $Y2=0
cc_98 N_C2_c_103_n N_Y_c_293_n 0.021152f $X=1.005 $Y=1.885 $X2=0 $Y2=0
cc_99 C2 N_Y_c_293_n 0.00862258f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_100 N_C2_c_102_n N_Y_c_295_n 0.0178302f $X=0.91 $Y=1.12 $X2=0 $Y2=0
cc_101 N_C2_c_103_n N_Y_c_295_n 0.00216104f $X=1.005 $Y=1.885 $X2=0 $Y2=0
cc_102 C2 N_Y_c_295_n 0.0237068f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_103 N_C2_c_103_n N_Y_c_285_n 0.00460586f $X=1.005 $Y=1.885 $X2=0 $Y2=0
cc_104 N_C2_c_103_n N_Y_c_286_n 0.00149128f $X=1.005 $Y=1.885 $X2=0 $Y2=0
cc_105 C2 N_Y_c_286_n 0.0163828f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_106 N_C2_c_102_n Y 0.00440102f $X=0.91 $Y=1.12 $X2=0 $Y2=0
cc_107 N_C2_c_103_n Y 0.00765712f $X=1.005 $Y=1.885 $X2=0 $Y2=0
cc_108 C2 Y 0.0526461f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_109 N_C2_c_103_n N_A_116_392#_c_361_n 0.0117097f $X=1.005 $Y=1.885 $X2=0
+ $Y2=0
cc_110 N_C2_c_103_n N_A_116_392#_c_358_n 0.012762f $X=1.005 $Y=1.885 $X2=0 $Y2=0
cc_111 N_C2_c_103_n N_A_116_392#_c_359_n 0.00169686f $X=1.005 $Y=1.885 $X2=0
+ $Y2=0
cc_112 N_C2_c_103_n N_VPWR_c_428_n 0.00278257f $X=1.005 $Y=1.885 $X2=0 $Y2=0
cc_113 N_C2_c_103_n N_VPWR_c_426_n 0.00359138f $X=1.005 $Y=1.885 $X2=0 $Y2=0
cc_114 N_C2_c_102_n N_VGND_c_465_n 0.00383152f $X=0.91 $Y=1.12 $X2=0 $Y2=0
cc_115 N_C2_c_102_n N_VGND_c_466_n 0.0102512f $X=0.91 $Y=1.12 $X2=0 $Y2=0
cc_116 N_C2_c_102_n N_VGND_c_467_n 0.00369533f $X=0.91 $Y=1.12 $X2=0 $Y2=0
cc_117 N_B2_c_140_n N_B1_c_178_n 0.0266842f $X=2.215 $Y=1.885 $X2=0 $Y2=0
cc_118 N_B2_c_136_n N_B1_c_174_n 0.0273469f $X=2.14 $Y=1.12 $X2=0 $Y2=0
cc_119 N_B2_c_137_n N_B1_c_175_n 0.0317442f $X=2.14 $Y=1.625 $X2=0 $Y2=0
cc_120 B2 B1 0.0438819f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_121 N_B2_c_139_n B1 0.00410205f $X=2.14 $Y=1.285 $X2=0 $Y2=0
cc_122 B2 N_B1_c_177_n 8.23261e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_123 N_B2_c_139_n N_B1_c_177_n 0.0273469f $X=2.14 $Y=1.285 $X2=0 $Y2=0
cc_124 N_B2_c_140_n N_Y_c_285_n 0.00180785f $X=2.215 $Y=1.885 $X2=0 $Y2=0
cc_125 N_B2_c_137_n N_Y_c_285_n 0.00251131f $X=2.14 $Y=1.625 $X2=0 $Y2=0
cc_126 B2 N_Y_c_285_n 4.44645e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_127 N_B2_c_140_n N_Y_c_286_n 0.00109537f $X=2.215 $Y=1.885 $X2=0 $Y2=0
cc_128 N_B2_c_136_n N_Y_c_280_n 0.0013851f $X=2.14 $Y=1.12 $X2=0 $Y2=0
cc_129 N_B2_c_136_n N_Y_c_318_n 0.0132291f $X=2.14 $Y=1.12 $X2=0 $Y2=0
cc_130 B2 N_Y_c_318_n 0.0233092f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_131 N_B2_c_139_n N_Y_c_318_n 0.00112191f $X=2.14 $Y=1.285 $X2=0 $Y2=0
cc_132 N_B2_c_136_n Y 0.00508329f $X=2.14 $Y=1.12 $X2=0 $Y2=0
cc_133 B2 Y 0.0496775f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_134 N_B2_c_139_n Y 0.00350374f $X=2.14 $Y=1.285 $X2=0 $Y2=0
cc_135 N_B2_c_137_n Y 0.00350374f $X=2.14 $Y=1.625 $X2=0 $Y2=0
cc_136 N_B2_c_140_n N_A_116_392#_c_358_n 0.0157136f $X=2.215 $Y=1.885 $X2=0
+ $Y2=0
cc_137 N_B2_c_140_n N_A_369_392#_c_388_n 0.0122144f $X=2.215 $Y=1.885 $X2=0
+ $Y2=0
cc_138 B2 N_A_369_392#_c_388_n 0.0108252f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_139 N_B2_c_140_n N_A_369_392#_c_386_n 0.00914301f $X=2.215 $Y=1.885 $X2=0
+ $Y2=0
cc_140 N_B2_c_137_n N_A_369_392#_c_386_n 0.00103923f $X=2.14 $Y=1.625 $X2=0
+ $Y2=0
cc_141 B2 N_A_369_392#_c_386_n 0.0129752f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_142 N_B2_c_140_n N_VPWR_c_428_n 0.00278271f $X=2.215 $Y=1.885 $X2=0 $Y2=0
cc_143 N_B2_c_140_n N_VPWR_c_426_n 0.00359139f $X=2.215 $Y=1.885 $X2=0 $Y2=0
cc_144 N_B2_c_136_n N_VGND_c_464_n 0.00383152f $X=2.14 $Y=1.12 $X2=0 $Y2=0
cc_145 N_B2_c_136_n N_VGND_c_466_n 0.00946983f $X=2.14 $Y=1.12 $X2=0 $Y2=0
cc_146 N_B2_c_136_n N_VGND_c_467_n 0.00369533f $X=2.14 $Y=1.12 $X2=0 $Y2=0
cc_147 N_B1_c_175_n N_A1_c_212_n 0.021061f $X=2.71 $Y=1.625 $X2=0 $Y2=0
cc_148 N_B1_c_178_n N_A1_c_217_n 0.0204794f $X=2.715 $Y=1.885 $X2=0 $Y2=0
cc_149 B1 N_A1_c_213_n 0.00258451f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_150 N_B1_c_177_n N_A1_c_213_n 0.0166638f $X=2.71 $Y=1.285 $X2=0 $Y2=0
cc_151 B1 N_A1_c_214_n 0.0352122f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_152 N_B1_c_177_n N_A1_c_214_n 0.00237949f $X=2.71 $Y=1.285 $X2=0 $Y2=0
cc_153 N_B1_c_174_n N_A1_c_215_n 0.00516683f $X=2.71 $Y=1.12 $X2=0 $Y2=0
cc_154 N_B1_c_174_n N_Y_c_280_n 0.0157946f $X=2.71 $Y=1.12 $X2=0 $Y2=0
cc_155 B1 N_Y_c_280_n 0.0262962f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_156 N_B1_c_177_n N_Y_c_280_n 0.00121333f $X=2.71 $Y=1.285 $X2=0 $Y2=0
cc_157 N_B1_c_178_n N_A_116_392#_c_358_n 0.00422861f $X=2.715 $Y=1.885 $X2=0
+ $Y2=0
cc_158 N_B1_c_178_n N_A_116_392#_c_366_n 0.00594533f $X=2.715 $Y=1.885 $X2=0
+ $Y2=0
cc_159 N_B1_c_178_n N_A_369_392#_c_388_n 0.0153046f $X=2.715 $Y=1.885 $X2=0
+ $Y2=0
cc_160 N_B1_c_175_n N_A_369_392#_c_388_n 4.64784e-19 $X=2.71 $Y=1.625 $X2=0
+ $Y2=0
cc_161 B1 N_A_369_392#_c_388_n 0.0198394f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_162 N_B1_c_178_n N_A_369_392#_c_383_n 0.00458691f $X=2.715 $Y=1.885 $X2=0
+ $Y2=0
cc_163 N_B1_c_178_n N_A_369_392#_c_386_n 4.54023e-19 $X=2.715 $Y=1.885 $X2=0
+ $Y2=0
cc_164 N_B1_c_175_n N_A_369_392#_c_387_n 3.16946e-19 $X=2.71 $Y=1.625 $X2=0
+ $Y2=0
cc_165 B1 N_A_369_392#_c_387_n 0.00328641f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_166 N_B1_c_178_n N_VPWR_c_428_n 0.0044313f $X=2.715 $Y=1.885 $X2=0 $Y2=0
cc_167 N_B1_c_178_n N_VPWR_c_426_n 0.00855151f $X=2.715 $Y=1.885 $X2=0 $Y2=0
cc_168 N_B1_c_174_n N_VGND_c_464_n 0.00288916f $X=2.71 $Y=1.12 $X2=0 $Y2=0
cc_169 N_B1_c_174_n N_VGND_c_466_n 7.41728e-19 $X=2.71 $Y=1.12 $X2=0 $Y2=0
cc_170 N_B1_c_174_n N_VGND_c_467_n 0.00359465f $X=2.71 $Y=1.12 $X2=0 $Y2=0
cc_171 N_A1_c_214_n N_A2_M1006_g 0.0074729f $X=3.32 $Y=1.285 $X2=0 $Y2=0
cc_172 N_A1_c_215_n N_A2_M1006_g 0.0263949f $X=3.305 $Y=1.12 $X2=0 $Y2=0
cc_173 N_A1_c_212_n N_A2_c_250_n 0.0298121f $X=3.305 $Y=1.61 $X2=0 $Y2=0
cc_174 N_A1_c_217_n N_A2_c_254_n 0.0238571f $X=3.215 $Y=1.885 $X2=0 $Y2=0
cc_175 N_A1_c_213_n A2 4.05463e-19 $X=3.32 $Y=1.285 $X2=0 $Y2=0
cc_176 N_A1_c_214_n A2 0.0495144f $X=3.32 $Y=1.285 $X2=0 $Y2=0
cc_177 N_A1_c_213_n N_A2_c_252_n 0.0263949f $X=3.32 $Y=1.285 $X2=0 $Y2=0
cc_178 N_A1_c_213_n N_Y_c_280_n 0.00268566f $X=3.32 $Y=1.285 $X2=0 $Y2=0
cc_179 N_A1_c_214_n N_Y_c_280_n 0.0149686f $X=3.32 $Y=1.285 $X2=0 $Y2=0
cc_180 N_A1_c_215_n N_Y_c_280_n 0.0116062f $X=3.305 $Y=1.12 $X2=0 $Y2=0
cc_181 N_A1_c_217_n N_A_116_392#_c_358_n 3.17734e-19 $X=3.215 $Y=1.885 $X2=0
+ $Y2=0
cc_182 N_A1_c_217_n N_A_369_392#_c_383_n 0.0103347f $X=3.215 $Y=1.885 $X2=0
+ $Y2=0
cc_183 N_A1_c_212_n N_A_369_392#_c_401_n 0.00116058f $X=3.305 $Y=1.61 $X2=0
+ $Y2=0
cc_184 N_A1_c_217_n N_A_369_392#_c_401_n 0.0126488f $X=3.215 $Y=1.885 $X2=0
+ $Y2=0
cc_185 N_A1_c_214_n N_A_369_392#_c_401_n 0.0413061f $X=3.32 $Y=1.285 $X2=0 $Y2=0
cc_186 N_A1_c_217_n N_A_369_392#_c_385_n 9.06108e-19 $X=3.215 $Y=1.885 $X2=0
+ $Y2=0
cc_187 N_A1_c_217_n N_A_369_392#_c_387_n 9.50925e-19 $X=3.215 $Y=1.885 $X2=0
+ $Y2=0
cc_188 N_A1_c_217_n N_VPWR_c_427_n 0.00658062f $X=3.215 $Y=1.885 $X2=0 $Y2=0
cc_189 N_A1_c_217_n N_VPWR_c_428_n 0.00445602f $X=3.215 $Y=1.885 $X2=0 $Y2=0
cc_190 N_A1_c_217_n N_VPWR_c_426_n 0.00858698f $X=3.215 $Y=1.885 $X2=0 $Y2=0
cc_191 N_A1_c_215_n N_VGND_c_463_n 0.00222027f $X=3.305 $Y=1.12 $X2=0 $Y2=0
cc_192 N_A1_c_215_n N_VGND_c_464_n 0.00432706f $X=3.305 $Y=1.12 $X2=0 $Y2=0
cc_193 N_A1_c_215_n N_VGND_c_467_n 0.00819572f $X=3.305 $Y=1.12 $X2=0 $Y2=0
cc_194 N_A2_M1006_g N_Y_c_280_n 0.00174219f $X=3.8 $Y=0.69 $X2=0 $Y2=0
cc_195 N_A2_c_254_n N_A_369_392#_c_383_n 8.72447e-19 $X=3.815 $Y=1.885 $X2=0
+ $Y2=0
cc_196 N_A2_c_254_n N_A_369_392#_c_401_n 0.0167469f $X=3.815 $Y=1.885 $X2=0
+ $Y2=0
cc_197 N_A2_c_254_n N_A_369_392#_c_384_n 7.95179e-19 $X=3.815 $Y=1.885 $X2=0
+ $Y2=0
cc_198 A2 N_A_369_392#_c_384_n 0.0252928f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_199 N_A2_c_252_n N_A_369_392#_c_384_n 0.00123847f $X=4.05 $Y=1.345 $X2=0
+ $Y2=0
cc_200 N_A2_c_254_n N_A_369_392#_c_385_n 0.0113134f $X=3.815 $Y=1.885 $X2=0
+ $Y2=0
cc_201 N_A2_c_254_n N_VPWR_c_427_n 0.00970855f $X=3.815 $Y=1.885 $X2=0 $Y2=0
cc_202 N_A2_c_254_n N_VPWR_c_430_n 0.00445602f $X=3.815 $Y=1.885 $X2=0 $Y2=0
cc_203 N_A2_c_254_n N_VPWR_c_426_n 0.00862798f $X=3.815 $Y=1.885 $X2=0 $Y2=0
cc_204 N_A2_M1006_g N_VGND_c_463_n 0.0161695f $X=3.8 $Y=0.69 $X2=0 $Y2=0
cc_205 A2 N_VGND_c_463_n 0.0184523f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_206 N_A2_c_252_n N_VGND_c_463_n 0.00206912f $X=4.05 $Y=1.345 $X2=0 $Y2=0
cc_207 N_A2_M1006_g N_VGND_c_464_n 0.00383152f $X=3.8 $Y=0.69 $X2=0 $Y2=0
cc_208 N_A2_M1006_g N_VGND_c_467_n 0.0075725f $X=3.8 $Y=0.69 $X2=0 $Y2=0
cc_209 N_Y_c_293_n N_A_116_392#_M1009_d 0.0105043f $X=1.115 $Y=2.045 $X2=-0.19
+ $Y2=-0.245
cc_210 N_Y_c_293_n N_A_116_392#_c_361_n 0.0202249f $X=1.115 $Y=2.045 $X2=0 $Y2=0
cc_211 N_Y_M1008_d N_A_116_392#_c_358_n 0.00355467f $X=1.08 $Y=1.96 $X2=0 $Y2=0
cc_212 N_Y_c_286_n N_A_116_392#_c_358_n 0.0400134f $X=1.28 $Y=2.125 $X2=0 $Y2=0
cc_213 N_Y_c_284_n N_A_116_392#_c_359_n 0.00371331f $X=0.28 $Y=2.815 $X2=0 $Y2=0
cc_214 N_Y_c_286_n N_A_369_392#_c_386_n 0.0681654f $X=1.28 $Y=2.125 $X2=0 $Y2=0
cc_215 N_Y_c_284_n N_VPWR_c_428_n 0.0145938f $X=0.28 $Y=2.815 $X2=0 $Y2=0
cc_216 N_Y_c_284_n N_VPWR_c_426_n 0.0120466f $X=0.28 $Y=2.815 $X2=0 $Y2=0
cc_217 N_Y_c_295_n A_119_74# 0.0072096f $X=1.485 $Y=0.865 $X2=-0.19 $Y2=-0.245
cc_218 N_Y_c_295_n N_VGND_M1011_d 0.0162958f $X=1.485 $Y=0.865 $X2=-0.19
+ $Y2=-0.245
cc_219 N_Y_c_318_n N_VGND_M1011_d 0.0126943f $X=2.525 $Y=0.64 $X2=-0.19
+ $Y2=-0.245
cc_220 Y N_VGND_M1011_d 0.00918472f $X=1.595 $Y=0.84 $X2=-0.19 $Y2=-0.245
cc_221 N_Y_c_280_n N_VGND_c_463_n 0.0207642f $X=3.195 $Y=0.495 $X2=0 $Y2=0
cc_222 N_Y_c_280_n N_VGND_c_464_n 0.0395123f $X=3.195 $Y=0.495 $X2=0 $Y2=0
cc_223 N_Y_c_278_n N_VGND_c_465_n 0.0144324f $X=0.305 $Y=0.515 $X2=0 $Y2=0
cc_224 N_Y_c_278_n N_VGND_c_466_n 0.00836615f $X=0.305 $Y=0.515 $X2=0 $Y2=0
cc_225 N_Y_c_295_n N_VGND_c_466_n 0.0349649f $X=1.485 $Y=0.865 $X2=0 $Y2=0
cc_226 N_Y_c_280_n N_VGND_c_466_n 0.00748454f $X=3.195 $Y=0.495 $X2=0 $Y2=0
cc_227 N_Y_c_318_n N_VGND_c_466_n 0.024446f $X=2.525 $Y=0.64 $X2=0 $Y2=0
cc_228 Y N_VGND_c_466_n 0.0257144f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_229 N_Y_c_278_n N_VGND_c_467_n 0.0119472f $X=0.305 $Y=0.515 $X2=0 $Y2=0
cc_230 N_Y_c_295_n N_VGND_c_467_n 0.0179064f $X=1.485 $Y=0.865 $X2=0 $Y2=0
cc_231 N_Y_c_280_n N_VGND_c_467_n 0.0302537f $X=3.195 $Y=0.495 $X2=0 $Y2=0
cc_232 N_Y_c_318_n N_VGND_c_467_n 0.0130236f $X=2.525 $Y=0.64 $X2=0 $Y2=0
cc_233 Y N_VGND_c_467_n 0.00127411f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_234 N_Y_c_318_n A_461_74# 0.0072096f $X=2.525 $Y=0.64 $X2=-0.19 $Y2=-0.245
cc_235 N_A_116_392#_c_358_n N_A_369_392#_M1001_s 0.00287371f $X=2.325 $Y=2.99
+ $X2=-0.19 $Y2=1.66
cc_236 N_A_116_392#_M1001_d N_A_369_392#_c_388_n 0.00985787f $X=2.29 $Y=1.96
+ $X2=0 $Y2=0
cc_237 N_A_116_392#_c_366_n N_A_369_392#_c_388_n 0.0202249f $X=2.49 $Y=2.465
+ $X2=0 $Y2=0
cc_238 N_A_116_392#_c_358_n N_A_369_392#_c_383_n 0.00395311f $X=2.325 $Y=2.99
+ $X2=0 $Y2=0
cc_239 N_A_116_392#_c_358_n N_A_369_392#_c_386_n 0.0205764f $X=2.325 $Y=2.99
+ $X2=0 $Y2=0
cc_240 N_A_116_392#_c_358_n N_VPWR_c_427_n 0.0027524f $X=2.325 $Y=2.99 $X2=0
+ $Y2=0
cc_241 N_A_116_392#_c_358_n N_VPWR_c_428_n 0.111616f $X=2.325 $Y=2.99 $X2=0
+ $Y2=0
cc_242 N_A_116_392#_c_359_n N_VPWR_c_428_n 0.0236039f $X=0.945 $Y=2.99 $X2=0
+ $Y2=0
cc_243 N_A_116_392#_c_358_n N_VPWR_c_426_n 0.0633416f $X=2.325 $Y=2.99 $X2=0
+ $Y2=0
cc_244 N_A_116_392#_c_359_n N_VPWR_c_426_n 0.012761f $X=0.945 $Y=2.99 $X2=0
+ $Y2=0
cc_245 N_A_369_392#_c_401_n N_VPWR_M1007_d 0.00841922f $X=3.875 $Y=2.045
+ $X2=-0.19 $Y2=1.66
cc_246 N_A_369_392#_c_383_n N_VPWR_c_427_n 0.0263057f $X=2.99 $Y=2.815 $X2=0
+ $Y2=0
cc_247 N_A_369_392#_c_401_n N_VPWR_c_427_n 0.0249771f $X=3.875 $Y=2.045 $X2=0
+ $Y2=0
cc_248 N_A_369_392#_c_385_n N_VPWR_c_427_n 0.0433294f $X=4.04 $Y=2.815 $X2=0
+ $Y2=0
cc_249 N_A_369_392#_c_383_n N_VPWR_c_428_n 0.0145938f $X=2.99 $Y=2.815 $X2=0
+ $Y2=0
cc_250 N_A_369_392#_c_385_n N_VPWR_c_430_n 0.0145938f $X=4.04 $Y=2.815 $X2=0
+ $Y2=0
cc_251 N_A_369_392#_c_383_n N_VPWR_c_426_n 0.0120466f $X=2.99 $Y=2.815 $X2=0
+ $Y2=0
cc_252 N_A_369_392#_c_385_n N_VPWR_c_426_n 0.0120466f $X=4.04 $Y=2.815 $X2=0
+ $Y2=0
