# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_ls__a21o_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.760000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485000 1.450000 4.195000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445000 1.260000 4.905000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.425000 1.435000 2.755000 1.780000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  1.086400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.960000 1.690000 1.130000 ;
        RECT 0.125000 1.130000 0.355000 1.800000 ;
        RECT 0.125000 1.800000 1.835000 1.970000 ;
        RECT 0.660000 0.350000 0.830000 0.960000 ;
        RECT 0.685000 1.970000 0.855000 2.980000 ;
        RECT 1.440000 0.350000 1.690000 0.960000 ;
        RECT 1.505000 1.970000 1.835000 2.980000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.760000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.760000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.760000 0.085000 ;
      RECT 0.000000  3.245000 5.760000 3.415000 ;
      RECT 0.150000  0.085000 0.480000 0.790000 ;
      RECT 0.155000  2.140000 0.485000 3.245000 ;
      RECT 0.635000  1.300000 2.205000 1.630000 ;
      RECT 1.010000  0.085000 1.260000 0.790000 ;
      RECT 1.055000  2.140000 1.305000 3.245000 ;
      RECT 1.870000  0.085000 2.120000 0.925000 ;
      RECT 1.870000  1.095000 3.255000 1.110000 ;
      RECT 1.870000  1.110000 4.220000 1.265000 ;
      RECT 1.870000  1.265000 2.205000 1.300000 ;
      RECT 2.035000  1.950000 2.285000 3.245000 ;
      RECT 2.360000  0.450000 2.610000 1.095000 ;
      RECT 2.475000  1.950000 2.725000 2.905000 ;
      RECT 2.475000  2.905000 3.625000 3.075000 ;
      RECT 2.790000  0.085000 3.120000 0.925000 ;
      RECT 2.925000  1.265000 4.220000 1.280000 ;
      RECT 2.925000  1.280000 3.255000 2.735000 ;
      RECT 3.455000  1.950000 5.505000 2.120000 ;
      RECT 3.455000  2.120000 3.625000 2.905000 ;
      RECT 3.460000  0.255000 4.570000 0.425000 ;
      RECT 3.460000  0.425000 3.790000 0.940000 ;
      RECT 3.825000  2.290000 4.075000 3.245000 ;
      RECT 3.960000  0.595000 4.220000 1.110000 ;
      RECT 4.275000  2.120000 4.525000 2.980000 ;
      RECT 4.400000  0.425000 4.570000 0.920000 ;
      RECT 4.400000  0.920000 5.510000 1.090000 ;
      RECT 4.725000  2.290000 5.055000 3.245000 ;
      RECT 4.750000  0.085000 5.080000 0.750000 ;
      RECT 5.255000  1.940000 5.505000 1.950000 ;
      RECT 5.255000  2.120000 5.505000 2.980000 ;
      RECT 5.260000  0.350000 5.510000 0.920000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
  END
END sky130_fd_sc_ls__a21o_4
END LIBRARY
