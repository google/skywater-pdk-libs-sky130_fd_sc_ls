* File: sky130_fd_sc_ls__dlygate4sd3_1.pxi.spice
* Created: Wed Sep  2 11:05:23 2020
* 
x_PM_SKY130_FD_SC_LS__DLYGATE4SD3_1%A N_A_M1005_g N_A_c_61_n N_A_c_65_n
+ N_A_M1002_g A A N_A_c_63_n PM_SKY130_FD_SC_LS__DLYGATE4SD3_1%A
x_PM_SKY130_FD_SC_LS__DLYGATE4SD3_1%A_28_74# N_A_28_74#_M1005_s
+ N_A_28_74#_M1002_s N_A_28_74#_c_94_n N_A_28_74#_c_98_n N_A_28_74#_c_99_n
+ N_A_28_74#_c_100_n N_A_28_74#_c_95_n N_A_28_74#_c_96_n N_A_28_74#_c_114_n
+ N_A_28_74#_M1007_g N_A_28_74#_M1003_g
+ PM_SKY130_FD_SC_LS__DLYGATE4SD3_1%A_28_74#
x_PM_SKY130_FD_SC_LS__DLYGATE4SD3_1%A_289_74# N_A_289_74#_M1007_d
+ N_A_289_74#_M1003_d N_A_289_74#_M1000_g N_A_289_74#_M1001_g
+ N_A_289_74#_c_150_n N_A_289_74#_c_151_n N_A_289_74#_c_152_n
+ N_A_289_74#_c_153_n N_A_289_74#_c_157_n N_A_289_74#_c_154_n
+ N_A_289_74#_c_155_n PM_SKY130_FD_SC_LS__DLYGATE4SD3_1%A_289_74#
x_PM_SKY130_FD_SC_LS__DLYGATE4SD3_1%A_405_138# N_A_405_138#_M1000_s
+ N_A_405_138#_M1001_s N_A_405_138#_M1006_g N_A_405_138#_c_202_n
+ N_A_405_138#_M1004_g N_A_405_138#_c_203_n N_A_405_138#_c_208_n
+ N_A_405_138#_c_204_n N_A_405_138#_c_205_n N_A_405_138#_c_206_n
+ N_A_405_138#_c_210_n PM_SKY130_FD_SC_LS__DLYGATE4SD3_1%A_405_138#
x_PM_SKY130_FD_SC_LS__DLYGATE4SD3_1%VPWR N_VPWR_M1002_d N_VPWR_M1001_d
+ N_VPWR_c_257_n N_VPWR_c_258_n N_VPWR_c_259_n N_VPWR_c_260_n VPWR
+ N_VPWR_c_261_n N_VPWR_c_262_n N_VPWR_c_256_n N_VPWR_c_264_n
+ PM_SKY130_FD_SC_LS__DLYGATE4SD3_1%VPWR
x_PM_SKY130_FD_SC_LS__DLYGATE4SD3_1%X N_X_M1006_d N_X_M1004_d X X X X X X X
+ N_X_c_289_n X X N_X_c_293_n PM_SKY130_FD_SC_LS__DLYGATE4SD3_1%X
x_PM_SKY130_FD_SC_LS__DLYGATE4SD3_1%VGND N_VGND_M1005_d N_VGND_M1000_d
+ N_VGND_c_309_n N_VGND_c_310_n N_VGND_c_311_n N_VGND_c_312_n VGND
+ N_VGND_c_313_n N_VGND_c_314_n N_VGND_c_315_n N_VGND_c_316_n
+ PM_SKY130_FD_SC_LS__DLYGATE4SD3_1%VGND
cc_1 VNB N_A_M1005_g 0.0437392f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=0.58
cc_2 VNB N_A_c_61_n 0.00890285f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.17
cc_3 VNB A 0.0265853f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_A_c_63_n 0.0358668f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.355
cc_5 VNB N_A_28_74#_c_94_n 0.0226356f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.545
cc_6 VNB N_A_28_74#_c_95_n 0.0126015f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.19
cc_7 VNB N_A_28_74#_c_96_n 0.0121635f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.52
cc_8 VNB N_A_28_74#_M1007_g 0.117704f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_289_74#_M1000_g 0.0495228f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.545
cc_10 VNB N_A_289_74#_M1001_g 0.00313542f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_289_74#_c_150_n 0.013071f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.355
cc_12 VNB N_A_289_74#_c_151_n 0.0161413f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.355
cc_13 VNB N_A_289_74#_c_152_n 0.0219379f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_289_74#_c_153_n 0.0495392f $X=-0.19 $Y=-0.245 $X2=0.415 $Y2=1.355
cc_15 VNB N_A_289_74#_c_154_n 0.00135856f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_289_74#_c_155_n 0.00336402f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_405_138#_M1006_g 0.0275176f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.545
cc_18 VNB N_A_405_138#_c_202_n 0.0358021f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_19 VNB N_A_405_138#_c_203_n 0.00175453f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.355
cc_20 VNB N_A_405_138#_c_204_n 0.00323188f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.52
cc_21 VNB N_A_405_138#_c_205_n 2.9305e-19 $X=-0.19 $Y=-0.245 $X2=0.415 $Y2=1.295
cc_22 VNB N_A_405_138#_c_206_n 0.00790239f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VPWR_c_256_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB X 0.0286532f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.545
cc_25 VNB N_X_c_289_n 0.029118f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB X 0.0145768f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_309_n 0.00961213f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.545
cc_28 VNB N_VGND_c_310_n 0.0187989f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_311_n 0.0567418f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.355
cc_30 VNB N_VGND_c_312_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.19
cc_31 VNB N_VGND_c_313_n 0.0180717f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_314_n 0.0205885f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_315_n 0.243362f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_316_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VPB N_A_c_61_n 0.0368635f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.17
cc_36 VPB N_A_c_65_n 0.0270096f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.26
cc_37 VPB A 0.0145994f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_38 VPB N_A_28_74#_c_98_n 0.0222081f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_39 VPB N_A_28_74#_c_99_n 0.00180999f $X=-0.19 $Y=1.66 $X2=0.57 $Y2=1.355
cc_40 VPB N_A_28_74#_c_100_n 0.0109668f $X=-0.19 $Y=1.66 $X2=0.57 $Y2=1.355
cc_41 VPB N_A_28_74#_M1007_g 0.0637558f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_42 VPB N_A_289_74#_M1001_g 0.0499439f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_43 VPB N_A_289_74#_c_157_n 0.00516643f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_44 VPB N_A_289_74#_c_154_n 0.0129551f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_45 VPB N_A_405_138#_c_202_n 0.0265074f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_46 VPB N_A_405_138#_c_208_n 0.00175644f $X=-0.19 $Y=1.66 $X2=0.57 $Y2=1.355
cc_47 VPB N_A_405_138#_c_205_n 0.00160201f $X=-0.19 $Y=1.66 $X2=0.415 $Y2=1.295
cc_48 VPB N_A_405_138#_c_210_n 0.00745707f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_257_n 0.0183719f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.545
cc_50 VPB N_VPWR_c_258_n 0.0111617f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_259_n 0.0596029f $X=-0.19 $Y=1.66 $X2=0.57 $Y2=1.52
cc_52 VPB N_VPWR_c_260_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0.415 $Y2=1.295
cc_53 VPB N_VPWR_c_261_n 0.018958f $X=-0.19 $Y=1.66 $X2=0.415 $Y2=1.355
cc_54 VPB N_VPWR_c_262_n 0.0200102f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_256_n 0.0940165f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_264_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB X 0.00819691f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.545
cc_58 VPB X 0.0507685f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_X_c_293_n 0.0146297f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 N_A_M1005_g N_A_28_74#_c_94_n 0.00873346f $X=0.48 $Y=0.58 $X2=0 $Y2=0
cc_61 N_A_c_65_n N_A_28_74#_c_98_n 0.00624408f $X=0.495 $Y=2.26 $X2=0 $Y2=0
cc_62 N_A_c_61_n N_A_28_74#_c_99_n 0.00956435f $X=0.495 $Y=2.17 $X2=0 $Y2=0
cc_63 N_A_c_65_n N_A_28_74#_c_99_n 0.00925083f $X=0.495 $Y=2.26 $X2=0 $Y2=0
cc_64 A N_A_28_74#_c_99_n 0.0262324f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_65 N_A_c_63_n N_A_28_74#_c_99_n 6.49888e-19 $X=0.57 $Y=1.355 $X2=0 $Y2=0
cc_66 A N_A_28_74#_c_100_n 0.0280303f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_67 N_A_M1005_g N_A_28_74#_c_95_n 0.0109614f $X=0.48 $Y=0.58 $X2=0 $Y2=0
cc_68 A N_A_28_74#_c_95_n 0.0251751f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_69 N_A_c_63_n N_A_28_74#_c_95_n 0.00146766f $X=0.57 $Y=1.355 $X2=0 $Y2=0
cc_70 N_A_M1005_g N_A_28_74#_c_96_n 0.00415005f $X=0.48 $Y=0.58 $X2=0 $Y2=0
cc_71 A N_A_28_74#_c_96_n 0.0289843f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_72 N_A_M1005_g N_A_28_74#_c_114_n 9.24862e-19 $X=0.48 $Y=0.58 $X2=0 $Y2=0
cc_73 N_A_c_61_n N_A_28_74#_c_114_n 0.0013064f $X=0.495 $Y=2.17 $X2=0 $Y2=0
cc_74 A N_A_28_74#_c_114_n 0.0410693f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_75 N_A_c_63_n N_A_28_74#_c_114_n 0.00110303f $X=0.57 $Y=1.355 $X2=0 $Y2=0
cc_76 N_A_M1005_g N_A_28_74#_M1007_g 0.0170485f $X=0.48 $Y=0.58 $X2=0 $Y2=0
cc_77 N_A_c_61_n N_A_28_74#_M1007_g 0.0251826f $X=0.495 $Y=2.17 $X2=0 $Y2=0
cc_78 N_A_c_65_n N_A_28_74#_M1007_g 0.012328f $X=0.495 $Y=2.26 $X2=0 $Y2=0
cc_79 A N_A_28_74#_M1007_g 0.0042554f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_80 N_A_c_63_n N_A_28_74#_M1007_g 0.0208886f $X=0.57 $Y=1.355 $X2=0 $Y2=0
cc_81 N_A_c_65_n N_VPWR_c_257_n 0.00399172f $X=0.495 $Y=2.26 $X2=0 $Y2=0
cc_82 N_A_c_65_n N_VPWR_c_261_n 0.00442668f $X=0.495 $Y=2.26 $X2=0 $Y2=0
cc_83 N_A_c_65_n N_VPWR_c_256_n 0.0048347f $X=0.495 $Y=2.26 $X2=0 $Y2=0
cc_84 N_A_M1005_g N_VGND_c_309_n 0.00249326f $X=0.48 $Y=0.58 $X2=0 $Y2=0
cc_85 N_A_M1005_g N_VGND_c_313_n 0.00456766f $X=0.48 $Y=0.58 $X2=0 $Y2=0
cc_86 N_A_M1005_g N_VGND_c_315_n 0.00454604f $X=0.48 $Y=0.58 $X2=0 $Y2=0
cc_87 N_A_28_74#_M1007_g N_A_289_74#_c_150_n 0.0114617f $X=1.195 $Y=0.58 $X2=0
+ $Y2=0
cc_88 N_A_28_74#_c_95_n N_A_289_74#_c_151_n 0.0164121f $X=0.975 $Y=0.92 $X2=0
+ $Y2=0
cc_89 N_A_28_74#_c_114_n N_A_289_74#_c_151_n 0.0277479f $X=1.14 $Y=1.295 $X2=0
+ $Y2=0
cc_90 N_A_28_74#_M1007_g N_A_289_74#_c_151_n 0.0169212f $X=1.195 $Y=0.58 $X2=0
+ $Y2=0
cc_91 N_A_28_74#_M1007_g N_A_289_74#_c_153_n 0.00416224f $X=1.195 $Y=0.58 $X2=0
+ $Y2=0
cc_92 N_A_28_74#_M1007_g N_A_289_74#_c_157_n 0.0102218f $X=1.195 $Y=0.58 $X2=0
+ $Y2=0
cc_93 N_A_28_74#_c_114_n N_A_289_74#_c_154_n 0.0295618f $X=1.14 $Y=1.295 $X2=0
+ $Y2=0
cc_94 N_A_28_74#_M1007_g N_A_289_74#_c_154_n 0.0203813f $X=1.195 $Y=0.58 $X2=0
+ $Y2=0
cc_95 N_A_28_74#_c_114_n N_A_289_74#_c_155_n 0.0193935f $X=1.14 $Y=1.295 $X2=0
+ $Y2=0
cc_96 N_A_28_74#_M1007_g N_A_289_74#_c_155_n 0.00352926f $X=1.195 $Y=0.58 $X2=0
+ $Y2=0
cc_97 N_A_28_74#_c_99_n N_VPWR_M1002_d 0.00835292f $X=0.975 $Y=2.117 $X2=-0.19
+ $Y2=-0.245
cc_98 N_A_28_74#_c_99_n N_VPWR_c_257_n 0.0227744f $X=0.975 $Y=2.117 $X2=0 $Y2=0
cc_99 N_A_28_74#_M1007_g N_VPWR_c_257_n 0.0119144f $X=1.195 $Y=0.58 $X2=0 $Y2=0
cc_100 N_A_28_74#_M1007_g N_VPWR_c_259_n 0.0151141f $X=1.195 $Y=0.58 $X2=0 $Y2=0
cc_101 N_A_28_74#_c_98_n N_VPWR_c_261_n 0.00593336f $X=0.265 $Y=2.56 $X2=0 $Y2=0
cc_102 N_A_28_74#_c_98_n N_VPWR_c_256_n 0.00940928f $X=0.265 $Y=2.56 $X2=0 $Y2=0
cc_103 N_A_28_74#_M1007_g N_VPWR_c_256_n 0.0292865f $X=1.195 $Y=0.58 $X2=0 $Y2=0
cc_104 N_A_28_74#_c_94_n N_VGND_c_309_n 0.0151665f $X=0.265 $Y=0.58 $X2=0 $Y2=0
cc_105 N_A_28_74#_c_95_n N_VGND_c_309_n 0.0244282f $X=0.975 $Y=0.92 $X2=0 $Y2=0
cc_106 N_A_28_74#_M1007_g N_VGND_c_309_n 0.00305775f $X=1.195 $Y=0.58 $X2=0
+ $Y2=0
cc_107 N_A_28_74#_M1007_g N_VGND_c_311_n 0.0150298f $X=1.195 $Y=0.58 $X2=0 $Y2=0
cc_108 N_A_28_74#_c_94_n N_VGND_c_313_n 0.0170785f $X=0.265 $Y=0.58 $X2=0 $Y2=0
cc_109 N_A_28_74#_c_94_n N_VGND_c_315_n 0.0118627f $X=0.265 $Y=0.58 $X2=0 $Y2=0
cc_110 N_A_28_74#_c_95_n N_VGND_c_315_n 0.018948f $X=0.975 $Y=0.92 $X2=0 $Y2=0
cc_111 N_A_28_74#_M1007_g N_VGND_c_315_n 0.0183085f $X=1.195 $Y=0.58 $X2=0 $Y2=0
cc_112 N_A_289_74#_M1000_g N_A_405_138#_M1006_g 0.021259f $X=2.535 $Y=0.9 $X2=0
+ $Y2=0
cc_113 N_A_289_74#_M1000_g N_A_405_138#_c_202_n 2.80094e-19 $X=2.535 $Y=0.9
+ $X2=0 $Y2=0
cc_114 N_A_289_74#_M1001_g N_A_405_138#_c_202_n 0.0313737f $X=2.535 $Y=2.34
+ $X2=0 $Y2=0
cc_115 N_A_289_74#_c_152_n N_A_405_138#_c_202_n 2.17534e-19 $X=2.575 $Y=1.465
+ $X2=0 $Y2=0
cc_116 N_A_289_74#_c_153_n N_A_405_138#_c_202_n 0.0215648f $X=2.575 $Y=1.465
+ $X2=0 $Y2=0
cc_117 N_A_289_74#_M1000_g N_A_405_138#_c_203_n 0.0347882f $X=2.535 $Y=0.9 $X2=0
+ $Y2=0
cc_118 N_A_289_74#_c_152_n N_A_405_138#_c_203_n 0.02741f $X=2.575 $Y=1.465 $X2=0
+ $Y2=0
cc_119 N_A_289_74#_M1001_g N_A_405_138#_c_208_n 0.0366973f $X=2.535 $Y=2.34
+ $X2=0 $Y2=0
cc_120 N_A_289_74#_c_152_n N_A_405_138#_c_208_n 0.0227169f $X=2.575 $Y=1.465
+ $X2=0 $Y2=0
cc_121 N_A_289_74#_M1000_g N_A_405_138#_c_204_n 0.00230419f $X=2.535 $Y=0.9
+ $X2=0 $Y2=0
cc_122 N_A_289_74#_c_152_n N_A_405_138#_c_204_n 0.0193923f $X=2.575 $Y=1.465
+ $X2=0 $Y2=0
cc_123 N_A_289_74#_c_153_n N_A_405_138#_c_204_n 0.00410963f $X=2.575 $Y=1.465
+ $X2=0 $Y2=0
cc_124 N_A_289_74#_M1001_g N_A_405_138#_c_205_n 0.00496065f $X=2.535 $Y=2.34
+ $X2=0 $Y2=0
cc_125 N_A_289_74#_M1000_g N_A_405_138#_c_206_n 0.0191803f $X=2.535 $Y=0.9 $X2=0
+ $Y2=0
cc_126 N_A_289_74#_c_151_n N_A_405_138#_c_206_n 0.0301027f $X=1.597 $Y=1.38
+ $X2=0 $Y2=0
cc_127 N_A_289_74#_c_152_n N_A_405_138#_c_206_n 0.0287835f $X=2.575 $Y=1.465
+ $X2=0 $Y2=0
cc_128 N_A_289_74#_c_153_n N_A_405_138#_c_206_n 0.00545878f $X=2.575 $Y=1.465
+ $X2=0 $Y2=0
cc_129 N_A_289_74#_M1001_g N_A_405_138#_c_210_n 0.0147779f $X=2.535 $Y=2.34
+ $X2=0 $Y2=0
cc_130 N_A_289_74#_c_152_n N_A_405_138#_c_210_n 0.0235446f $X=2.575 $Y=1.465
+ $X2=0 $Y2=0
cc_131 N_A_289_74#_c_153_n N_A_405_138#_c_210_n 0.00490082f $X=2.575 $Y=1.465
+ $X2=0 $Y2=0
cc_132 N_A_289_74#_c_154_n N_A_405_138#_c_210_n 0.021975f $X=1.567 $Y=2.395
+ $X2=0 $Y2=0
cc_133 N_A_289_74#_M1001_g N_VPWR_c_258_n 0.00865052f $X=2.535 $Y=2.34 $X2=0
+ $Y2=0
cc_134 N_A_289_74#_M1001_g N_VPWR_c_259_n 0.0164683f $X=2.535 $Y=2.34 $X2=0
+ $Y2=0
cc_135 N_A_289_74#_c_157_n N_VPWR_c_259_n 0.00561205f $X=1.58 $Y=2.56 $X2=0
+ $Y2=0
cc_136 N_A_289_74#_M1001_g N_VPWR_c_256_n 0.016946f $X=2.535 $Y=2.34 $X2=0 $Y2=0
cc_137 N_A_289_74#_c_157_n N_VPWR_c_256_n 0.00918412f $X=1.58 $Y=2.56 $X2=0
+ $Y2=0
cc_138 N_A_289_74#_c_150_n N_VGND_c_309_n 0.00634199f $X=1.597 $Y=0.635 $X2=0
+ $Y2=0
cc_139 N_A_289_74#_M1000_g N_VGND_c_310_n 0.00512562f $X=2.535 $Y=0.9 $X2=0
+ $Y2=0
cc_140 N_A_289_74#_M1000_g N_VGND_c_311_n 0.0124333f $X=2.535 $Y=0.9 $X2=0 $Y2=0
cc_141 N_A_289_74#_c_150_n N_VGND_c_311_n 0.0163385f $X=1.597 $Y=0.635 $X2=0
+ $Y2=0
cc_142 N_A_289_74#_M1000_g N_VGND_c_315_n 0.0150611f $X=2.535 $Y=0.9 $X2=0 $Y2=0
cc_143 N_A_289_74#_c_150_n N_VGND_c_315_n 0.0113715f $X=1.597 $Y=0.635 $X2=0
+ $Y2=0
cc_144 N_A_405_138#_c_208_n N_VPWR_M1001_d 0.00262668f $X=2.91 $Y=1.91 $X2=0
+ $Y2=0
cc_145 N_A_405_138#_c_202_n N_VPWR_c_258_n 0.0153694f $X=3.215 $Y=1.765 $X2=0
+ $Y2=0
cc_146 N_A_405_138#_c_208_n N_VPWR_c_258_n 0.0222367f $X=2.91 $Y=1.91 $X2=0
+ $Y2=0
cc_147 N_A_405_138#_c_202_n N_VPWR_c_262_n 0.00413917f $X=3.215 $Y=1.765 $X2=0
+ $Y2=0
cc_148 N_A_405_138#_c_202_n N_VPWR_c_256_n 0.00821556f $X=3.215 $Y=1.765 $X2=0
+ $Y2=0
cc_149 N_A_405_138#_M1006_g X 0.00260428f $X=3.205 $Y=0.74 $X2=0 $Y2=0
cc_150 N_A_405_138#_c_202_n X 0.0110819f $X=3.215 $Y=1.765 $X2=0 $Y2=0
cc_151 N_A_405_138#_c_204_n X 0.0327059f $X=3.032 $Y=1.625 $X2=0 $Y2=0
cc_152 N_A_405_138#_c_205_n X 0.00709928f $X=3.032 $Y=1.825 $X2=0 $Y2=0
cc_153 N_A_405_138#_M1006_g N_X_c_289_n 0.00143568f $X=3.205 $Y=0.74 $X2=0 $Y2=0
cc_154 N_A_405_138#_c_204_n X 0.0037592f $X=3.032 $Y=1.625 $X2=0 $Y2=0
cc_155 N_A_405_138#_c_202_n N_X_c_293_n 0.00396238f $X=3.215 $Y=1.765 $X2=0
+ $Y2=0
cc_156 N_A_405_138#_c_208_n N_X_c_293_n 0.00776663f $X=2.91 $Y=1.91 $X2=0 $Y2=0
cc_157 N_A_405_138#_c_205_n N_X_c_293_n 7.53348e-19 $X=3.032 $Y=1.825 $X2=0
+ $Y2=0
cc_158 N_A_405_138#_c_203_n N_VGND_M1000_d 7.12223e-19 $X=2.91 $Y=1.125 $X2=0
+ $Y2=0
cc_159 N_A_405_138#_c_204_n N_VGND_M1000_d 0.0018038f $X=3.032 $Y=1.625 $X2=0
+ $Y2=0
cc_160 N_A_405_138#_M1006_g N_VGND_c_310_n 0.0156117f $X=3.205 $Y=0.74 $X2=0
+ $Y2=0
cc_161 N_A_405_138#_c_202_n N_VGND_c_310_n 4.77198e-19 $X=3.215 $Y=1.765 $X2=0
+ $Y2=0
cc_162 N_A_405_138#_c_203_n N_VGND_c_310_n 0.00549591f $X=2.91 $Y=1.125 $X2=0
+ $Y2=0
cc_163 N_A_405_138#_c_204_n N_VGND_c_310_n 0.016728f $X=3.032 $Y=1.625 $X2=0
+ $Y2=0
cc_164 N_A_405_138#_c_206_n N_VGND_c_311_n 0.00526925f $X=2.15 $Y=0.875 $X2=0
+ $Y2=0
cc_165 N_A_405_138#_M1006_g N_VGND_c_314_n 0.00383152f $X=3.205 $Y=0.74 $X2=0
+ $Y2=0
cc_166 N_A_405_138#_M1006_g N_VGND_c_315_n 0.00761589f $X=3.205 $Y=0.74 $X2=0
+ $Y2=0
cc_167 N_A_405_138#_c_206_n N_VGND_c_315_n 0.0100411f $X=2.15 $Y=0.875 $X2=0
+ $Y2=0
cc_168 N_VPWR_c_258_n X 0.0378466f $X=2.99 $Y=2.27 $X2=0 $Y2=0
cc_169 N_VPWR_c_262_n X 0.0270407f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_170 N_VPWR_c_256_n X 0.0159412f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_171 N_X_c_289_n N_VGND_c_310_n 0.019927f $X=3.42 $Y=0.52 $X2=0 $Y2=0
cc_172 N_X_c_289_n N_VGND_c_314_n 0.0180659f $X=3.42 $Y=0.52 $X2=0 $Y2=0
cc_173 N_X_c_289_n N_VGND_c_315_n 0.0152075f $X=3.42 $Y=0.52 $X2=0 $Y2=0
