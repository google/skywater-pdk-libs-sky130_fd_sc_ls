* File: sky130_fd_sc_ls__xnor2_1.pex.spice
* Created: Fri Aug 28 14:08:39 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__XNOR2_1%B 1 3 4 6 7 9 12 15 16 17 19 23 26 36
c82 36 0 1.14536e-19 $X=1.26 $Y=1.607
c83 16 0 6.8969e-20 $X=2.015 $Y=2.035
r84 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.11
+ $Y=1.6 $X2=1.11 $Y2=1.6
r85 26 36 2.00425 $w=3.43e-07 $l=6e-08 $layer=LI1_cond $X=1.2 $Y=1.607 $X2=1.26
+ $Y2=1.607
r86 26 30 3.00637 $w=3.43e-07 $l=9e-08 $layer=LI1_cond $X=1.2 $Y=1.607 $X2=1.11
+ $Y2=1.607
r87 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.3
+ $Y=1.515 $X2=2.3 $Y2=1.515
r88 20 23 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=2.1 $Y=1.515 $X2=2.3
+ $Y2=1.515
r89 18 20 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.1 $Y=1.68 $X2=2.1
+ $Y2=1.515
r90 18 19 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=2.1 $Y=1.68 $X2=2.1
+ $Y2=1.95
r91 16 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.015 $Y=2.035
+ $X2=2.1 $Y2=1.95
r92 16 17 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.015 $Y=2.035
+ $X2=1.345 $Y2=2.035
r93 15 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.26 $Y=1.95
+ $X2=1.345 $Y2=2.035
r94 14 36 4.88813 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=1.26 $Y=1.78
+ $X2=1.26 $Y2=1.607
r95 14 15 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.26 $Y=1.78
+ $X2=1.26 $Y2=1.95
r96 10 24 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=2.39 $Y=1.35
+ $X2=2.3 $Y2=1.515
r97 10 12 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.39 $Y=1.35
+ $X2=2.39 $Y2=0.74
r98 7 24 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=2.225 $Y=1.765
+ $X2=2.3 $Y2=1.515
r99 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.225 $Y=1.765
+ $X2=2.225 $Y2=2.4
r100 4 29 50.3854 $w=3.55e-07 $l=2.70647e-07 $layer=POLY_cond $X=1.065 $Y=1.85
+ $X2=1.022 $Y2=1.6
r101 4 6 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.065 $Y=1.85
+ $X2=1.065 $Y2=2.345
r102 1 29 55.8164 $w=3.55e-07 $l=3.68008e-07 $layer=POLY_cond $X=0.845 $Y=1.31
+ $X2=1.022 $Y2=1.6
r103 1 3 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.845 $Y=1.31
+ $X2=0.845 $Y2=0.915
.ends

.subckt PM_SKY130_FD_SC_LS__XNOR2_1%A 4 5 7 8 9 10 12 16 19 21 25
c62 19 0 1.14536e-19 $X=0.615 $Y=1.775
r63 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.68
+ $Y=1.515 $X2=1.68 $Y2=1.515
r64 21 25 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.68 $Y=1.665
+ $X2=1.68 $Y2=1.515
r65 17 19 66.6596 $w=1.5e-07 $l=1.3e-07 $layer=POLY_cond $X=0.485 $Y=1.775
+ $X2=0.615 $Y2=1.775
r66 14 24 38.6704 $w=3.39e-07 $l=2.13014e-07 $layer=POLY_cond $X=1.815 $Y=1.35
+ $X2=1.705 $Y2=1.515
r67 14 16 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.815 $Y=1.35
+ $X2=1.815 $Y2=0.74
r68 13 16 248.691 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=1.815 $Y=0.255
+ $X2=1.815 $Y2=0.74
r69 10 24 50.756 $w=3.39e-07 $l=2.95804e-07 $layer=POLY_cond $X=1.805 $Y=1.765
+ $X2=1.705 $Y2=1.515
r70 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.805 $Y=1.765
+ $X2=1.805 $Y2=2.4
r71 8 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.74 $Y=0.18
+ $X2=1.815 $Y2=0.255
r72 8 9 605.064 $w=1.5e-07 $l=1.18e-06 $layer=POLY_cond $X=1.74 $Y=0.18 $X2=0.56
+ $Y2=0.18
r73 5 19 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.615 $Y=1.85
+ $X2=0.615 $Y2=1.775
r74 5 7 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.615 $Y=1.85
+ $X2=0.615 $Y2=2.345
r75 2 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.485 $Y=1.7
+ $X2=0.485 $Y2=1.775
r76 2 4 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=0.485 $Y=1.7
+ $X2=0.485 $Y2=0.915
r77 1 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.485 $Y=0.255
+ $X2=0.56 $Y2=0.18
r78 1 4 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.485 $Y=0.255
+ $X2=0.485 $Y2=0.915
.ends

.subckt PM_SKY130_FD_SC_LS__XNOR2_1%A_138_385# 1 2 7 9 12 20 22 23 27 28 30
c82 7 0 2.58324e-19 $X=2.795 $Y=1.765
r83 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.84
+ $Y=1.465 $X2=2.84 $Y2=1.465
r84 30 32 18.887 $w=2.39e-07 $l=3.7e-07 $layer=LI1_cond $X=2.785 $Y=1.095
+ $X2=2.785 $Y2=1.465
r85 27 28 8.64761 $w=3.98e-07 $l=1.65e-07 $layer=LI1_cond $X=0.805 $Y=2.115
+ $X2=0.805 $Y2=1.95
r86 22 30 2.73298 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=2.635 $Y=1.095
+ $X2=2.785 $Y2=1.095
r87 22 23 91.9893 $w=1.68e-07 $l=1.41e-06 $layer=LI1_cond $X=2.635 $Y=1.095
+ $X2=1.225 $Y2=1.095
r88 18 23 10.0923 $w=2.09e-07 $l=1.82565e-07 $layer=LI1_cond $X=1.06 $Y=1.132
+ $X2=1.225 $Y2=1.095
r89 18 24 21.5981 $w=2.09e-07 $l=3.7e-07 $layer=LI1_cond $X=1.06 $Y=1.132
+ $X2=0.69 $Y2=1.132
r90 18 20 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=1.06 $Y=1.01
+ $X2=1.06 $Y2=0.74
r91 14 24 1.94907 $w=1.7e-07 $l=1.23e-07 $layer=LI1_cond $X=0.69 $Y=1.255
+ $X2=0.69 $Y2=1.132
r92 14 28 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=0.69 $Y=1.255
+ $X2=0.69 $Y2=1.95
r93 10 33 38.6549 $w=2.86e-07 $l=1.74714e-07 $layer=POLY_cond $X=2.82 $Y=1.3
+ $X2=2.84 $Y2=1.465
r94 10 12 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.82 $Y=1.3 $X2=2.82
+ $Y2=0.74
r95 7 33 61.4066 $w=2.86e-07 $l=3.21714e-07 $layer=POLY_cond $X=2.795 $Y=1.765
+ $X2=2.84 $Y2=1.465
r96 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.795 $Y=1.765
+ $X2=2.795 $Y2=2.4
r97 2 27 300 $w=1.7e-07 $l=2.54165e-07 $layer=licon1_PDIFF $count=2 $X=0.69
+ $Y=1.925 $X2=0.84 $Y2=2.115
r98 1 20 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.92
+ $Y=0.595 $X2=1.06 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__XNOR2_1%VPWR 1 2 3 12 14 15 17 20 24 26 29 31 36 45
+ 49
c48 3 0 1.38916e-19 $X=2.87 $Y=1.84
r49 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r50 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r51 40 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r52 39 40 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r53 37 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.745 $Y=3.33
+ $X2=1.58 $Y2=3.33
r54 37 39 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=1.745 $Y=3.33
+ $X2=2.64 $Y2=3.33
r55 36 48 4.61575 $w=1.7e-07 $l=2.52e-07 $layer=LI1_cond $X=2.855 $Y=3.33
+ $X2=3.107 $Y2=3.33
r56 36 39 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.855 $Y=3.33
+ $X2=2.64 $Y2=3.33
r57 35 43 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.24 $Y2=3.33
r58 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r59 32 42 4.61231 $w=1.7e-07 $l=2.53e-07 $layer=LI1_cond $X=0.505 $Y=3.33
+ $X2=0.252 $Y2=3.33
r60 32 34 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=0.505 $Y=3.33
+ $X2=1.2 $Y2=3.33
r61 31 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.415 $Y=3.33
+ $X2=1.58 $Y2=3.33
r62 31 34 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.415 $Y=3.33
+ $X2=1.2 $Y2=3.33
r63 29 40 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r64 29 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r65 29 45 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r66 24 48 3.15043 $w=3.3e-07 $l=1.22327e-07 $layer=LI1_cond $X=3.02 $Y=3.245
+ $X2=3.107 $Y2=3.33
r67 24 26 33.0018 $w=3.28e-07 $l=9.45e-07 $layer=LI1_cond $X=3.02 $Y=3.245
+ $X2=3.02 $Y2=2.3
r68 20 23 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=1.58 $Y=2.415 $X2=1.58
+ $Y2=2.815
r69 18 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.58 $Y=3.245
+ $X2=1.58 $Y2=3.33
r70 18 23 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=1.58 $Y=3.245
+ $X2=1.58 $Y2=2.815
r71 15 42 3.15387 $w=3.3e-07 $l=1.23386e-07 $layer=LI1_cond $X=0.34 $Y=3.245
+ $X2=0.252 $Y2=3.33
r72 15 17 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.34 $Y=3.245
+ $X2=0.34 $Y2=2.535
r73 14 28 6.46688 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.34 $Y=2.455
+ $X2=0.34 $Y2=2.29
r74 14 17 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=0.34 $Y=2.455 $X2=0.34
+ $Y2=2.535
r75 12 28 10.1415 $w=2.48e-07 $l=2.2e-07 $layer=LI1_cond $X=0.3 $Y=2.07 $X2=0.3
+ $Y2=2.29
r76 3 26 300 $w=1.7e-07 $l=5.29717e-07 $layer=licon1_PDIFF $count=2 $X=2.87
+ $Y=1.84 $X2=3.02 $Y2=2.3
r77 2 23 600 $w=1.7e-07 $l=1.08798e-06 $layer=licon1_PDIFF $count=1 $X=1.14
+ $Y=1.925 $X2=1.58 $Y2=2.815
r78 2 20 600 $w=1.7e-07 $l=6.75056e-07 $layer=licon1_PDIFF $count=1 $X=1.14
+ $Y=1.925 $X2=1.58 $Y2=2.415
r79 1 17 600 $w=1.7e-07 $l=6.78638e-07 $layer=licon1_PDIFF $count=1 $X=0.195
+ $Y=1.925 $X2=0.34 $Y2=2.535
r80 1 12 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.195
+ $Y=1.925 $X2=0.34 $Y2=2.07
.ends

.subckt PM_SKY130_FD_SC_LS__XNOR2_1%Y 1 2 7 9 13 16 19 20 26
c34 16 0 1.38916e-19 $X=3.19 $Y=1.85
r35 20 26 6.24041 $w=6.88e-07 $l=3.6e-07 $layer=LI1_cond $X=2.16 $Y=2.635
+ $X2=2.52 $Y2=2.635
r36 16 19 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=3.19 $Y=1.85
+ $X2=3.19 $Y2=1.13
r37 11 19 7.90841 $w=2.98e-07 $l=1.5e-07 $layer=LI1_cond $X=3.125 $Y=0.98
+ $X2=3.125 $Y2=1.13
r38 11 13 17.8629 $w=2.98e-07 $l=4.65e-07 $layer=LI1_cond $X=3.125 $Y=0.98
+ $X2=3.125 $Y2=0.515
r39 10 18 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.685 $Y=1.935
+ $X2=2.52 $Y2=1.935
r40 9 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.105 $Y=1.935
+ $X2=3.19 $Y2=1.85
r41 9 10 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=3.105 $Y=1.935
+ $X2=2.685 $Y2=1.935
r42 8 26 5.06645 $w=3.3e-07 $l=3.45e-07 $layer=LI1_cond $X=2.52 $Y=2.29 $X2=2.52
+ $Y2=2.635
r43 7 18 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.52 $Y=2.02 $X2=2.52
+ $Y2=1.935
r44 7 8 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=2.52 $Y=2.02 $X2=2.52
+ $Y2=2.29
r45 2 26 300 $w=1.7e-07 $l=6.7611e-07 $layer=licon1_PDIFF $count=2 $X=2.3
+ $Y=1.84 $X2=2.52 $Y2=2.415
r46 2 18 600 $w=1.7e-07 $l=2.94788e-07 $layer=licon1_PDIFF $count=1 $X=2.3
+ $Y=1.84 $X2=2.52 $Y2=2.015
r47 1 13 91 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=2 $X=2.895
+ $Y=0.37 $X2=3.06 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__XNOR2_1%VGND 1 2 7 9 13 15 17 27 28 34
r37 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r38 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r39 28 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.16
+ $Y2=0
r40 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r41 25 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.265 $Y=0 $X2=2.1
+ $Y2=0
r42 25 27 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=2.265 $Y=0 $X2=3.12
+ $Y2=0
r43 21 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r44 20 23 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r45 20 21 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r46 18 31 4.75569 $w=1.7e-07 $l=2.18e-07 $layer=LI1_cond $X=0.435 $Y=0 $X2=0.217
+ $Y2=0
r47 18 20 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.435 $Y=0 $X2=0.72
+ $Y2=0
r48 17 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.935 $Y=0 $X2=2.1
+ $Y2=0
r49 17 23 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.935 $Y=0 $X2=1.68
+ $Y2=0
r50 15 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r51 15 21 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r52 15 23 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r53 11 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.1 $Y=0.085 $X2=2.1
+ $Y2=0
r54 11 13 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=2.1 $Y=0.085
+ $X2=2.1 $Y2=0.37
r55 7 31 3.01048 $w=3.3e-07 $l=1.08305e-07 $layer=LI1_cond $X=0.27 $Y=0.085
+ $X2=0.217 $Y2=0
r56 7 9 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=0.27 $Y=0.085
+ $X2=0.27 $Y2=0.74
r57 2 13 182 $w=1.7e-07 $l=2.1e-07 $layer=licon1_NDIFF $count=1 $X=1.89 $Y=0.37
+ $X2=2.1 $Y2=0.37
r58 1 9 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.595 $X2=0.27 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__XNOR2_1%A_293_74# 1 2 7 10 15
c28 15 0 1.89355e-19 $X=2.605 $Y=0.675
r29 15 17 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=2.605 $Y=0.675
+ $X2=2.605 $Y2=0.755
r30 10 12 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=1.6 $Y=0.675 $X2=1.6
+ $Y2=0.755
r31 8 12 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.765 $Y=0.755
+ $X2=1.6 $Y2=0.755
r32 7 17 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.44 $Y=0.755
+ $X2=2.605 $Y2=0.755
r33 7 8 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=2.44 $Y=0.755
+ $X2=1.765 $Y2=0.755
r34 2 15 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=2.465
+ $Y=0.37 $X2=2.605 $Y2=0.675
r35 1 10 182 $w=1.7e-07 $l=3.66333e-07 $layer=licon1_NDIFF $count=1 $X=1.465
+ $Y=0.37 $X2=1.6 $Y2=0.675
.ends

