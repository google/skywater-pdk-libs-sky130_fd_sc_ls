* File: sky130_fd_sc_ls__o2111ai_4.pex.spice
* Created: Wed Sep  2 11:17:04 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__O2111AI_4%D1 1 3 4 6 7 9 10 12 13 15 16 18 19 20 21
+ 35
c60 16 0 2.41904e-19 $X=1.855 $Y=1.185
r61 35 36 4.32934 $w=5.01e-07 $l=4.5e-08 $layer=POLY_cond $X=1.81 $Y=1.475
+ $X2=1.855 $Y2=1.475
r62 34 35 37.0399 $w=5.01e-07 $l=3.85e-07 $layer=POLY_cond $X=1.425 $Y=1.475
+ $X2=1.81 $Y2=1.475
r63 33 34 15.8743 $w=5.01e-07 $l=1.65e-07 $layer=POLY_cond $X=1.26 $Y=1.475
+ $X2=1.425 $Y2=1.475
r64 31 33 7.21557 $w=5.01e-07 $l=7.5e-08 $layer=POLY_cond $X=1.185 $Y=1.475
+ $X2=1.26 $Y2=1.475
r65 31 32 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.185
+ $Y=1.515 $X2=1.185 $Y2=1.515
r66 29 31 18.2794 $w=5.01e-07 $l=1.9e-07 $layer=POLY_cond $X=0.995 $Y=1.475
+ $X2=1.185 $Y2=1.475
r67 27 29 47.1417 $w=5.01e-07 $l=4.9e-07 $layer=POLY_cond $X=0.505 $Y=1.475
+ $X2=0.995 $Y2=1.475
r68 27 28 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.505
+ $Y=1.515 $X2=0.505 $Y2=1.515
r69 25 27 0.962076 $w=5.01e-07 $l=1e-08 $layer=POLY_cond $X=0.495 $Y=1.475
+ $X2=0.505 $Y2=1.475
r70 21 32 0.402015 $w=4.28e-07 $l=1.5e-08 $layer=LI1_cond $X=1.2 $Y=1.565
+ $X2=1.185 $Y2=1.565
r71 20 32 12.4625 $w=4.28e-07 $l=4.65e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=1.185 $Y2=1.565
r72 20 28 5.76222 $w=4.28e-07 $l=2.15e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=0.505 $Y2=1.565
r73 19 28 7.10226 $w=4.28e-07 $l=2.65e-07 $layer=LI1_cond $X=0.24 $Y=1.565
+ $X2=0.505 $Y2=1.565
r74 16 36 31.4585 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=1.855 $Y=1.185
+ $X2=1.855 $Y2=1.475
r75 16 18 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.855 $Y=1.185
+ $X2=1.855 $Y2=0.74
r76 13 35 31.4585 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=1.81 $Y=1.765
+ $X2=1.81 $Y2=1.475
r77 13 15 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.81 $Y=1.765
+ $X2=1.81 $Y2=2.4
r78 10 34 31.4585 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=1.425 $Y=1.185
+ $X2=1.425 $Y2=1.475
r79 10 12 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.425 $Y=1.185
+ $X2=1.425 $Y2=0.74
r80 7 33 31.4585 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=1.26 $Y=1.765
+ $X2=1.26 $Y2=1.475
r81 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.26 $Y=1.765
+ $X2=1.26 $Y2=2.4
r82 4 29 31.4585 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=0.995 $Y=1.185
+ $X2=0.995 $Y2=1.475
r83 4 6 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=0.995 $Y=1.185
+ $X2=0.995 $Y2=0.74
r84 1 25 31.4585 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=0.495 $Y=1.185
+ $X2=0.495 $Y2=1.475
r85 1 3 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=0.495 $Y=1.185
+ $X2=0.495 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__O2111AI_4%C1 1 3 4 6 7 9 10 12 13 15 16 17 18 20 29
+ 39
c76 16 0 6.98451e-20 $X=3.5 $Y=1.26
c77 4 0 2.84156e-19 $X=2.285 $Y=1.185
r78 36 37 1.34387 $w=5.38e-07 $l=1.5e-08 $layer=POLY_cond $X=3.13 $Y=1.475
+ $X2=3.145 $Y2=1.475
r79 31 32 2.23978 $w=5.38e-07 $l=2.5e-08 $layer=POLY_cond $X=2.26 $Y=1.475
+ $X2=2.285 $Y2=1.475
r80 29 39 4.04332 $w=4.78e-07 $l=1.15e-07 $layer=LI1_cond $X=4.08 $Y=1.54
+ $X2=3.965 $Y2=1.54
r81 28 36 6.71933 $w=5.38e-07 $l=7.5e-08 $layer=POLY_cond $X=3.055 $Y=1.475
+ $X2=3.13 $Y2=1.475
r82 28 34 30.461 $w=5.38e-07 $l=3.4e-07 $layer=POLY_cond $X=3.055 $Y=1.475
+ $X2=2.715 $Y2=1.475
r83 27 39 31.7795 $w=3.28e-07 $l=9.1e-07 $layer=LI1_cond $X=3.055 $Y=1.465
+ $X2=3.965 $Y2=1.465
r84 27 28 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.055
+ $Y=1.465 $X2=3.055 $Y2=1.465
r85 24 34 30.461 $w=5.38e-07 $l=3.4e-07 $layer=POLY_cond $X=2.375 $Y=1.475
+ $X2=2.715 $Y2=1.475
r86 24 32 8.0632 $w=5.38e-07 $l=9e-08 $layer=POLY_cond $X=2.375 $Y=1.475
+ $X2=2.285 $Y2=1.475
r87 23 27 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=2.375 $Y=1.465
+ $X2=3.055 $Y2=1.465
r88 23 24 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.375
+ $Y=1.465 $X2=2.375 $Y2=1.465
r89 18 20 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=3.575 $Y=1.185
+ $X2=3.575 $Y2=0.74
r90 17 37 34.859 $w=5.38e-07 $l=2.497e-07 $layer=POLY_cond $X=3.22 $Y=1.26
+ $X2=3.145 $Y2=1.475
r91 16 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.5 $Y=1.26
+ $X2=3.575 $Y2=1.185
r92 16 17 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.5 $Y=1.26 $X2=3.22
+ $Y2=1.26
r93 13 37 33.2685 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=3.145 $Y=1.185
+ $X2=3.145 $Y2=1.475
r94 13 15 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=3.145 $Y=1.185
+ $X2=3.145 $Y2=0.74
r95 10 36 33.2685 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=3.13 $Y=1.765
+ $X2=3.13 $Y2=1.475
r96 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.13 $Y=1.765
+ $X2=3.13 $Y2=2.4
r97 7 34 33.2685 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.715 $Y=1.185
+ $X2=2.715 $Y2=1.475
r98 7 9 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.715 $Y=1.185
+ $X2=2.715 $Y2=0.74
r99 4 32 33.2685 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.285 $Y=1.185
+ $X2=2.285 $Y2=1.475
r100 4 6 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.285 $Y=1.185
+ $X2=2.285 $Y2=0.74
r101 1 31 33.2685 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.26 $Y=1.765
+ $X2=2.26 $Y2=1.475
r102 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.26 $Y=1.765
+ $X2=2.26 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__O2111AI_4%B1 1 3 4 5 6 8 13 17 21 23 25 27 28 29 30
+ 31 37
c88 37 0 1.99442e-19 $X=4.49 $Y=1.537
c89 17 0 3.32178e-19 $X=4.995 $Y=0.74
c90 1 0 2.47931e-20 $X=3.58 $Y=1.765
r91 44 45 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.675
+ $Y=1.515 $X2=5.675 $Y2=1.515
r92 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.655
+ $Y=1.515 $X2=4.655 $Y2=1.515
r93 31 45 8.71033 $w=4.28e-07 $l=3.25e-07 $layer=LI1_cond $X=6 $Y=1.565
+ $X2=5.675 $Y2=1.565
r94 30 45 4.15415 $w=4.28e-07 $l=1.55e-07 $layer=LI1_cond $X=5.52 $Y=1.565
+ $X2=5.675 $Y2=1.565
r95 29 30 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=5.04 $Y=1.565
+ $X2=5.52 $Y2=1.565
r96 29 40 10.3184 $w=4.28e-07 $l=3.85e-07 $layer=LI1_cond $X=5.04 $Y=1.565
+ $X2=4.655 $Y2=1.565
r97 28 40 2.54609 $w=4.28e-07 $l=9.5e-08 $layer=LI1_cond $X=4.56 $Y=1.565
+ $X2=4.655 $Y2=1.565
r98 23 44 26.6954 $w=3.75e-07 $l=1.8e-07 $layer=POLY_cond $X=5.855 $Y=1.537
+ $X2=5.675 $Y2=1.537
r99 23 25 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.855 $Y=1.35
+ $X2=5.855 $Y2=0.74
r100 19 44 37.0769 $w=3.75e-07 $l=2.5e-07 $layer=POLY_cond $X=5.425 $Y=1.537
+ $X2=5.675 $Y2=1.537
r101 19 21 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.425 $Y=1.35
+ $X2=5.425 $Y2=0.74
r102 15 19 63.7723 $w=3.75e-07 $l=4.3e-07 $layer=POLY_cond $X=4.995 $Y=1.537
+ $X2=5.425 $Y2=1.537
r103 15 39 50.4246 $w=3.75e-07 $l=3.4e-07 $layer=POLY_cond $X=4.995 $Y=1.537
+ $X2=4.655 $Y2=1.537
r104 15 17 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.995 $Y=1.35
+ $X2=4.995 $Y2=0.74
r105 11 39 13.3477 $w=3.75e-07 $l=9e-08 $layer=POLY_cond $X=4.565 $Y=1.537
+ $X2=4.655 $Y2=1.537
r106 11 37 31.8081 $w=3.75e-07 $l=7.5e-08 $layer=POLY_cond $X=4.565 $Y=1.537
+ $X2=4.49 $Y2=1.537
r107 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.565 $Y=1.35
+ $X2=4.565 $Y2=0.74
r108 10 27 20.4101 $w=1.5e-07 $l=9.94987e-08 $layer=POLY_cond $X=4.22 $Y=1.65
+ $X2=4.13 $Y2=1.67
r109 10 37 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=4.22 $Y=1.65
+ $X2=4.49 $Y2=1.65
r110 6 27 5.30422 $w=1.5e-07 $l=9.5e-08 $layer=POLY_cond $X=4.13 $Y=1.765
+ $X2=4.13 $Y2=1.67
r111 6 8 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.13 $Y=1.765
+ $X2=4.13 $Y2=2.4
r112 4 27 20.4101 $w=1.5e-07 $l=9.94987e-08 $layer=POLY_cond $X=4.04 $Y=1.65
+ $X2=4.13 $Y2=1.67
r113 4 5 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=4.04 $Y=1.65 $X2=3.67
+ $Y2=1.65
r114 1 5 26.9307 $w=1.5e-07 $l=1.53542e-07 $layer=POLY_cond $X=3.58 $Y=1.765
+ $X2=3.67 $Y2=1.65
r115 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.58 $Y=1.765
+ $X2=3.58 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__O2111AI_4%A1 1 3 6 8 10 13 15 17 20 22 24 27 29 30
+ 31 46 47
c87 46 0 1.08803e-20 $X=7.47 $Y=1.515
c88 22 0 1.03312e-19 $X=7.625 $Y=1.765
c89 13 0 1.61888e-19 $X=6.855 $Y=0.74
c90 6 0 8.45991e-20 $X=6.355 $Y=0.74
r91 47 48 11.1804 $w=3.88e-07 $l=9e-08 $layer=POLY_cond $X=7.625 $Y=1.542
+ $X2=7.715 $Y2=1.542
r92 45 47 19.2552 $w=3.88e-07 $l=1.55e-07 $layer=POLY_cond $X=7.47 $Y=1.542
+ $X2=7.625 $Y2=1.542
r93 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.47
+ $Y=1.515 $X2=7.47 $Y2=1.515
r94 43 45 22.982 $w=3.88e-07 $l=1.85e-07 $layer=POLY_cond $X=7.285 $Y=1.542
+ $X2=7.47 $Y2=1.542
r95 42 43 13.6649 $w=3.88e-07 $l=1.1e-07 $layer=POLY_cond $X=7.175 $Y=1.542
+ $X2=7.285 $Y2=1.542
r96 41 42 39.7526 $w=3.88e-07 $l=3.2e-07 $layer=POLY_cond $X=6.855 $Y=1.542
+ $X2=7.175 $Y2=1.542
r97 40 41 16.1495 $w=3.88e-07 $l=1.3e-07 $layer=POLY_cond $X=6.725 $Y=1.542
+ $X2=6.855 $Y2=1.542
r98 38 40 34.1624 $w=3.88e-07 $l=2.75e-07 $layer=POLY_cond $X=6.45 $Y=1.542
+ $X2=6.725 $Y2=1.542
r99 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.45
+ $Y=1.515 $X2=6.45 $Y2=1.515
r100 36 38 11.8015 $w=3.88e-07 $l=9.5e-08 $layer=POLY_cond $X=6.355 $Y=1.542
+ $X2=6.45 $Y2=1.542
r101 35 36 11.8015 $w=3.88e-07 $l=9.5e-08 $layer=POLY_cond $X=6.26 $Y=1.542
+ $X2=6.355 $Y2=1.542
r102 31 46 0.80403 $w=4.28e-07 $l=3e-08 $layer=LI1_cond $X=7.44 $Y=1.565
+ $X2=7.47 $Y2=1.565
r103 30 31 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=6.96 $Y=1.565
+ $X2=7.44 $Y2=1.565
r104 29 30 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=6.48 $Y=1.565
+ $X2=6.96 $Y2=1.565
r105 29 39 0.80403 $w=4.28e-07 $l=3e-08 $layer=LI1_cond $X=6.48 $Y=1.565
+ $X2=6.45 $Y2=1.565
r106 25 48 25.1189 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=7.715 $Y=1.32
+ $X2=7.715 $Y2=1.542
r107 25 27 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=7.715 $Y=1.32
+ $X2=7.715 $Y2=0.74
r108 22 47 25.1189 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=7.625 $Y=1.765
+ $X2=7.625 $Y2=1.542
r109 22 24 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.625 $Y=1.765
+ $X2=7.625 $Y2=2.4
r110 18 43 25.1189 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=7.285 $Y=1.32
+ $X2=7.285 $Y2=1.542
r111 18 20 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=7.285 $Y=1.32
+ $X2=7.285 $Y2=0.74
r112 15 42 25.1189 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=7.175 $Y=1.765
+ $X2=7.175 $Y2=1.542
r113 15 17 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.175 $Y=1.765
+ $X2=7.175 $Y2=2.4
r114 11 41 25.1189 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=6.855 $Y=1.32
+ $X2=6.855 $Y2=1.542
r115 11 13 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.855 $Y=1.32
+ $X2=6.855 $Y2=0.74
r116 8 40 25.1189 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=6.725 $Y=1.765
+ $X2=6.725 $Y2=1.542
r117 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.725 $Y=1.765
+ $X2=6.725 $Y2=2.4
r118 4 36 25.1189 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=6.355 $Y=1.32
+ $X2=6.355 $Y2=1.542
r119 4 6 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.355 $Y=1.32
+ $X2=6.355 $Y2=0.74
r120 1 35 25.1189 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=6.26 $Y=1.765
+ $X2=6.26 $Y2=1.542
r121 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.26 $Y=1.765
+ $X2=6.26 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__O2111AI_4%A2 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 26 27 28 44 45
c83 44 0 1.03312e-19 $X=9.405 $Y=1.515
c84 1 0 1.08803e-20 $X=8.09 $Y=1.765
r85 45 46 0.95069 $w=5.07e-07 $l=1e-08 $layer=POLY_cond $X=9.575 $Y=1.495
+ $X2=9.585 $Y2=1.495
r86 43 45 16.1617 $w=5.07e-07 $l=1.7e-07 $layer=POLY_cond $X=9.405 $Y=1.495
+ $X2=9.575 $Y2=1.495
r87 43 44 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.405
+ $Y=1.515 $X2=9.405 $Y2=1.515
r88 41 43 23.7673 $w=5.07e-07 $l=2.5e-07 $layer=POLY_cond $X=9.155 $Y=1.495
+ $X2=9.405 $Y2=1.495
r89 40 41 7.60552 $w=5.07e-07 $l=8e-08 $layer=POLY_cond $X=9.075 $Y=1.495
+ $X2=9.155 $Y2=1.495
r90 39 40 40.8797 $w=5.07e-07 $l=4.3e-07 $layer=POLY_cond $X=8.645 $Y=1.495
+ $X2=9.075 $Y2=1.495
r91 38 39 6.65483 $w=5.07e-07 $l=7e-08 $layer=POLY_cond $X=8.575 $Y=1.495
+ $X2=8.645 $Y2=1.495
r92 36 38 18.0631 $w=5.07e-07 $l=1.9e-07 $layer=POLY_cond $X=8.385 $Y=1.495
+ $X2=8.575 $Y2=1.495
r93 36 37 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.385
+ $Y=1.515 $X2=8.385 $Y2=1.515
r94 34 36 22.8166 $w=5.07e-07 $l=2.4e-07 $layer=POLY_cond $X=8.145 $Y=1.495
+ $X2=8.385 $Y2=1.495
r95 33 34 5.2288 $w=5.07e-07 $l=5.5e-08 $layer=POLY_cond $X=8.09 $Y=1.495
+ $X2=8.145 $Y2=1.495
r96 28 44 1.20605 $w=4.28e-07 $l=4.5e-08 $layer=LI1_cond $X=9.36 $Y=1.565
+ $X2=9.405 $Y2=1.565
r97 27 28 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=8.88 $Y=1.565
+ $X2=9.36 $Y2=1.565
r98 26 27 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=8.4 $Y=1.565
+ $X2=8.88 $Y2=1.565
r99 26 37 0.402015 $w=4.28e-07 $l=1.5e-08 $layer=LI1_cond $X=8.4 $Y=1.565
+ $X2=8.385 $Y2=1.565
r100 25 37 12.4625 $w=4.28e-07 $l=4.65e-07 $layer=LI1_cond $X=7.92 $Y=1.565
+ $X2=8.385 $Y2=1.565
r101 22 46 31.7597 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=9.585 $Y=1.225
+ $X2=9.585 $Y2=1.495
r102 22 24 155.847 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=9.585 $Y=1.225
+ $X2=9.585 $Y2=0.74
r103 19 45 31.7597 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=9.575 $Y=1.765
+ $X2=9.575 $Y2=1.495
r104 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=9.575 $Y=1.765
+ $X2=9.575 $Y2=2.4
r105 16 41 31.7597 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=9.155 $Y=1.225
+ $X2=9.155 $Y2=1.495
r106 16 18 155.847 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=9.155 $Y=1.225
+ $X2=9.155 $Y2=0.74
r107 13 40 31.7597 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=9.075 $Y=1.765
+ $X2=9.075 $Y2=1.495
r108 13 15 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=9.075 $Y=1.765
+ $X2=9.075 $Y2=2.4
r109 10 39 31.7597 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=8.645 $Y=1.225
+ $X2=8.645 $Y2=1.495
r110 10 12 155.847 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=8.645 $Y=1.225
+ $X2=8.645 $Y2=0.74
r111 7 38 31.7597 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=8.575 $Y=1.765
+ $X2=8.575 $Y2=1.495
r112 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.575 $Y=1.765
+ $X2=8.575 $Y2=2.4
r113 4 34 31.7597 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=8.145 $Y=1.225
+ $X2=8.145 $Y2=1.495
r114 4 6 155.847 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=8.145 $Y=1.225
+ $X2=8.145 $Y2=0.74
r115 1 33 31.7597 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=8.09 $Y=1.765
+ $X2=8.09 $Y2=1.495
r116 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.09 $Y=1.765
+ $X2=8.09 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__O2111AI_4%Y 1 2 3 4 5 6 7 8 25 29 31 32 35 37 38 41
+ 43 47 49 53 65 68 74 76 78 79
c134 43 0 6.98451e-20 $X=4.19 $Y=2.035
c135 37 0 2.47931e-20 $X=3.19 $Y=1.885
c136 31 0 9.95308e-20 $X=1.685 $Y=1.13
r137 71 72 1.74613 $w=3.28e-07 $l=5e-08 $layer=LI1_cond $X=3.355 $Y=1.985
+ $X2=3.355 $Y2=2.035
r138 68 71 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=3.355 $Y=1.885
+ $X2=3.355 $Y2=1.985
r139 64 65 13.0168 $w=1.028e-06 $l=1.65e-07 $layer=LI1_cond $X=1.035 $Y=2.465
+ $X2=1.2 $Y2=2.465
r140 61 64 4.50097 $w=1.028e-06 $l=3.8e-07 $layer=LI1_cond $X=0.655 $Y=2.465
+ $X2=1.035 $Y2=2.465
r141 58 61 4.44175 $w=1.028e-06 $l=3.75e-07 $layer=LI1_cond $X=0.28 $Y=2.465
+ $X2=0.655 $Y2=2.465
r142 54 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.515 $Y=2.035
+ $X2=8.35 $Y2=2.035
r143 53 78 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.185 $Y=2.035
+ $X2=9.35 $Y2=2.035
r144 53 54 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.185 $Y=2.035
+ $X2=8.515 $Y2=2.035
r145 50 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.52 $Y=2.035
+ $X2=4.355 $Y2=2.035
r146 49 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.185 $Y=2.035
+ $X2=8.35 $Y2=2.035
r147 49 50 239.107 $w=1.68e-07 $l=3.665e-06 $layer=LI1_cond $X=8.185 $Y=2.035
+ $X2=4.52 $Y2=2.035
r148 45 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.355 $Y=2.12
+ $X2=4.355 $Y2=2.035
r149 45 47 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=4.355 $Y=2.12
+ $X2=4.355 $Y2=2.815
r150 44 72 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.52 $Y=2.035
+ $X2=3.355 $Y2=2.035
r151 43 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.19 $Y=2.035
+ $X2=4.355 $Y2=2.035
r152 43 44 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.19 $Y=2.035
+ $X2=3.52 $Y2=2.035
r153 39 72 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=3.355 $Y=2.12
+ $X2=3.355 $Y2=2.035
r154 39 41 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=3.355 $Y=2.12
+ $X2=3.355 $Y2=2.815
r155 38 85 8.97309 $w=3.43e-07 $l=1.88348e-07 $layer=LI1_cond $X=2.2 $Y=1.885
+ $X2=2.035 $Y2=1.835
r156 37 68 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.19 $Y=1.885
+ $X2=3.355 $Y2=1.885
r157 37 38 64.5882 $w=1.68e-07 $l=9.9e-07 $layer=LI1_cond $X=3.19 $Y=1.885
+ $X2=2.2 $Y2=1.885
r158 33 85 0.950996 $w=3.3e-07 $l=2.85e-07 $layer=LI1_cond $X=2.035 $Y=2.12
+ $X2=2.035 $Y2=1.835
r159 33 35 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=2.035 $Y=2.12
+ $X2=2.035 $Y2=2.815
r160 32 85 12.449 $w=3.43e-07 $l=4.71434e-07 $layer=LI1_cond $X=1.685 $Y=1.55
+ $X2=2.035 $Y2=1.835
r161 32 79 0.177843 $w=3.43e-07 $l=1.17473e-07 $layer=LI1_cond $X=1.685 $Y=1.55
+ $X2=1.68 $Y2=1.665
r162 31 67 4.30634 $w=2.4e-07 $l=1.8e-07 $layer=LI1_cond $X=1.685 $Y=1.13
+ $X2=1.685 $Y2=0.95
r163 31 32 20.1678 $w=2.38e-07 $l=4.2e-07 $layer=LI1_cond $X=1.685 $Y=1.13
+ $X2=1.685 $Y2=1.55
r164 29 79 9.8623 $w=3.43e-07 $l=4.55192e-07 $layer=LI1_cond $X=1.87 $Y=2.035
+ $X2=1.68 $Y2=1.665
r165 29 65 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.87 $Y=2.035
+ $X2=1.2 $Y2=2.035
r166 25 67 2.87089 $w=3.6e-07 $l=1.2e-07 $layer=LI1_cond $X=1.565 $Y=0.95
+ $X2=1.685 $Y2=0.95
r167 25 27 25.1297 $w=3.58e-07 $l=7.85e-07 $layer=LI1_cond $X=1.565 $Y=0.95
+ $X2=0.78 $Y2=0.95
r168 8 78 300 $w=1.7e-07 $l=3.61421e-07 $layer=licon1_PDIFF $count=2 $X=9.15
+ $Y=1.84 $X2=9.35 $Y2=2.115
r169 7 76 300 $w=1.7e-07 $l=3.55668e-07 $layer=licon1_PDIFF $count=2 $X=8.165
+ $Y=1.84 $X2=8.35 $Y2=2.115
r170 6 74 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=4.205
+ $Y=1.84 $X2=4.355 $Y2=2.115
r171 6 47 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=4.205
+ $Y=1.84 $X2=4.355 $Y2=2.815
r172 5 71 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=3.205
+ $Y=1.84 $X2=3.355 $Y2=1.985
r173 5 41 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=3.205
+ $Y=1.84 $X2=3.355 $Y2=2.815
r174 4 85 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.885
+ $Y=1.84 $X2=2.035 $Y2=1.985
r175 4 35 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.885
+ $Y=1.84 $X2=2.035 $Y2=2.815
r176 3 64 266.667 $w=1.7e-07 $l=1.1463e-06 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.84 $X2=1.035 $Y2=2.4
r177 3 61 266.667 $w=1.7e-07 $l=1.20732e-06 $layer=licon1_PDIFF $count=2
+ $X=0.135 $Y=1.84 $X2=0.655 $Y2=2.815
r178 3 61 266.667 $w=1.7e-07 $l=6.09754e-07 $layer=licon1_PDIFF $count=2
+ $X=0.135 $Y=1.84 $X2=0.655 $Y2=2.035
r179 3 58 266.667 $w=1.7e-07 $l=6.28331e-07 $layer=licon1_PDIFF $count=2
+ $X=0.135 $Y=1.84 $X2=0.28 $Y2=2.4
r180 2 67 182 $w=1.7e-07 $l=6.0597e-07 $layer=licon1_NDIFF $count=1 $X=1.5
+ $Y=0.37 $X2=1.64 $Y2=0.91
r181 1 27 182 $w=1.7e-07 $l=6.76905e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.78 $Y2=0.95
.ends

.subckt PM_SKY130_FD_SC_LS__O2111AI_4%VPWR 1 2 3 4 5 18 22 26 30 34 37 38 40 41
+ 42 51 59 66 73 74 77 80 83
r99 83 84 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r100 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r101 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r102 74 84 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=7.44 $Y2=3.33
r103 73 74 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r104 71 83 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.485 $Y=3.33
+ $X2=7.4 $Y2=3.33
r105 71 73 153.642 $w=1.68e-07 $l=2.355e-06 $layer=LI1_cond $X=7.485 $Y=3.33
+ $X2=9.84 $Y2=3.33
r106 70 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.44 $Y2=3.33
r107 70 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6.48 $Y2=3.33
r108 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r109 67 80 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.585 $Y=3.33
+ $X2=6.46 $Y2=3.33
r110 67 69 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=6.585 $Y=3.33
+ $X2=6.96 $Y2=3.33
r111 66 83 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.315 $Y=3.33
+ $X2=7.4 $Y2=3.33
r112 66 69 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=7.315 $Y=3.33
+ $X2=6.96 $Y2=3.33
r113 65 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r114 64 65 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r115 61 64 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.08 $Y=3.33 $X2=6
+ $Y2=3.33
r116 61 62 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r117 59 80 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.335 $Y=3.33
+ $X2=6.46 $Y2=3.33
r118 59 64 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=6.335 $Y=3.33
+ $X2=6 $Y2=3.33
r119 58 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r120 58 78 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=2.64 $Y2=3.33
r121 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r122 55 77 13.1282 $w=1.7e-07 $l=3.25e-07 $layer=LI1_cond $X=3.02 $Y=3.33
+ $X2=2.695 $Y2=3.33
r123 55 57 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=3.02 $Y=3.33
+ $X2=3.6 $Y2=3.33
r124 54 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r125 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r126 51 77 13.1282 $w=1.7e-07 $l=3.25e-07 $layer=LI1_cond $X=2.37 $Y=3.33
+ $X2=2.695 $Y2=3.33
r127 51 53 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=2.37 $Y=3.33
+ $X2=2.16 $Y2=3.33
r128 50 54 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r129 49 50 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r130 46 50 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r131 45 49 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=3.33 $X2=1.2
+ $Y2=3.33
r132 45 46 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r133 42 65 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33 $X2=6
+ $Y2=3.33
r134 42 62 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.08 $Y2=3.33
r135 40 57 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=3.69 $Y=3.33 $X2=3.6
+ $Y2=3.33
r136 40 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.69 $Y=3.33
+ $X2=3.855 $Y2=3.33
r137 39 61 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=4.02 $Y=3.33 $X2=4.08
+ $Y2=3.33
r138 39 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.02 $Y=3.33
+ $X2=3.855 $Y2=3.33
r139 37 49 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.37 $Y=3.33
+ $X2=1.2 $Y2=3.33
r140 37 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.37 $Y=3.33
+ $X2=1.535 $Y2=3.33
r141 36 53 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=1.7 $Y=3.33
+ $X2=2.16 $Y2=3.33
r142 36 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.7 $Y=3.33
+ $X2=1.535 $Y2=3.33
r143 32 83 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.4 $Y=3.245 $X2=7.4
+ $Y2=3.33
r144 32 34 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=7.4 $Y=3.245
+ $X2=7.4 $Y2=2.805
r145 28 80 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.46 $Y=3.245
+ $X2=6.46 $Y2=3.33
r146 28 30 20.283 $w=2.48e-07 $l=4.4e-07 $layer=LI1_cond $X=6.46 $Y=3.245
+ $X2=6.46 $Y2=2.805
r147 24 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.855 $Y=3.245
+ $X2=3.855 $Y2=3.33
r148 24 26 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=3.855 $Y=3.245
+ $X2=3.855 $Y2=2.455
r149 20 77 2.7021 $w=6.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.695 $Y=3.245
+ $X2=2.695 $Y2=3.33
r150 20 22 17.2971 $w=6.48e-07 $l=9.4e-07 $layer=LI1_cond $X=2.695 $Y=3.245
+ $X2=2.695 $Y2=2.305
r151 16 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.535 $Y=3.245
+ $X2=1.535 $Y2=3.33
r152 16 18 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=1.535 $Y=3.245
+ $X2=1.535 $Y2=2.455
r153 5 34 600 $w=1.7e-07 $l=1.03729e-06 $layer=licon1_PDIFF $count=1 $X=7.25
+ $Y=1.84 $X2=7.4 $Y2=2.805
r154 4 30 600 $w=1.7e-07 $l=1.04425e-06 $layer=licon1_PDIFF $count=1 $X=6.335
+ $Y=1.84 $X2=6.5 $Y2=2.805
r155 3 26 300 $w=1.7e-07 $l=7.07972e-07 $layer=licon1_PDIFF $count=2 $X=3.655
+ $Y=1.84 $X2=3.855 $Y2=2.455
r156 2 22 150 $w=1.7e-07 $l=7.68082e-07 $layer=licon1_PDIFF $count=4 $X=2.335
+ $Y=1.84 $X2=2.905 $Y2=2.305
r157 1 18 300 $w=1.7e-07 $l=7.07972e-07 $layer=licon1_PDIFF $count=2 $X=1.335
+ $Y=1.84 $X2=1.535 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_LS__O2111AI_4%A_954_368# 1 2 3 4 5 16 22 26 28 29 30 31
+ 34 36 40 46 48 51
r68 45 46 10.2208 $w=6.88e-07 $l=1.35e-07 $layer=LI1_cond $X=6.03 $Y=2.635
+ $X2=6.165 $Y2=2.635
r69 40 43 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=9.84 $Y=1.985
+ $X2=9.84 $Y2=2.815
r70 38 43 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=9.84 $Y=2.905 $X2=9.84
+ $Y2=2.815
r71 37 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.015 $Y=2.99
+ $X2=8.85 $Y2=2.99
r72 36 38 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=9.715 $Y=2.99
+ $X2=9.84 $Y2=2.905
r73 36 37 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=9.715 $Y=2.99
+ $X2=9.015 $Y2=2.99
r74 32 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.85 $Y=2.905
+ $X2=8.85 $Y2=2.99
r75 32 34 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=8.85 $Y=2.905
+ $X2=8.85 $Y2=2.455
r76 30 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.685 $Y=2.99
+ $X2=8.85 $Y2=2.99
r77 30 31 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.685 $Y=2.99
+ $X2=8.015 $Y2=2.99
r78 29 31 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.85 $Y=2.905
+ $X2=8.015 $Y2=2.99
r79 28 50 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.85 $Y=2.46 $X2=7.85
+ $Y2=2.375
r80 28 29 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=7.85 $Y=2.46
+ $X2=7.85 $Y2=2.905
r81 27 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.115 $Y=2.375
+ $X2=6.95 $Y2=2.375
r82 26 50 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.685 $Y=2.375
+ $X2=7.85 $Y2=2.375
r83 26 27 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=7.685 $Y=2.375
+ $X2=7.115 $Y2=2.375
r84 22 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.785 $Y=2.375
+ $X2=6.95 $Y2=2.375
r85 22 46 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=6.785 $Y=2.375
+ $X2=6.165 $Y2=2.375
r86 18 21 12.5675 $w=6.88e-07 $l=7.25e-07 $layer=LI1_cond $X=4.945 $Y=2.635
+ $X2=5.67 $Y2=2.635
r87 16 45 3.64024 $w=6.88e-07 $l=2.1e-07 $layer=LI1_cond $X=5.82 $Y=2.635
+ $X2=6.03 $Y2=2.635
r88 16 21 2.60017 $w=6.88e-07 $l=1.5e-07 $layer=LI1_cond $X=5.82 $Y=2.635
+ $X2=5.67 $Y2=2.635
r89 5 43 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=9.65
+ $Y=1.84 $X2=9.8 $Y2=2.815
r90 5 40 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=9.65
+ $Y=1.84 $X2=9.8 $Y2=1.985
r91 4 34 300 $w=1.7e-07 $l=7.07972e-07 $layer=licon1_PDIFF $count=2 $X=8.65
+ $Y=1.84 $X2=8.85 $Y2=2.455
r92 3 50 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=7.7
+ $Y=1.84 $X2=7.85 $Y2=2.455
r93 2 48 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=6.8
+ $Y=1.84 $X2=6.95 $Y2=2.455
r94 1 45 300 $w=1.7e-07 $l=1.50389e-06 $layer=licon1_PDIFF $count=2 $X=4.77
+ $Y=1.84 $X2=6.03 $Y2=2.375
r95 1 21 200 $w=1.7e-07 $l=1.13644e-06 $layer=licon1_PDIFF $count=3 $X=4.77
+ $Y=1.84 $X2=5.67 $Y2=2.375
r96 1 18 200 $w=1.7e-07 $l=6.1632e-07 $layer=licon1_PDIFF $count=3 $X=4.77
+ $Y=1.84 $X2=4.945 $Y2=2.375
.ends

.subckt PM_SKY130_FD_SC_LS__O2111AI_4%A_27_74# 1 2 3 4 5 18 22 23 28 31
c47 23 0 1.61246e-19 $X=2.07 $Y=0.815
c48 22 0 1.84625e-19 $X=2.07 $Y=0.6
r49 26 28 31.4635 $w=3.13e-07 $l=8.6e-07 $layer=LI1_cond $X=2.93 $Y=0.972
+ $X2=3.79 $Y2=0.972
r50 24 35 2.68365 $w=3.15e-07 $l=8.5e-08 $layer=LI1_cond $X=2.155 $Y=0.972
+ $X2=2.07 $Y2=0.972
r51 24 26 28.3538 $w=3.13e-07 $l=7.75e-07 $layer=LI1_cond $X=2.155 $Y=0.972
+ $X2=2.93 $Y2=0.972
r52 23 35 4.95685 $w=1.7e-07 $l=1.57e-07 $layer=LI1_cond $X=2.07 $Y=0.815
+ $X2=2.07 $Y2=0.972
r53 22 33 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.07 $Y=0.6 $X2=2.07
+ $Y2=0.475
r54 22 23 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.07 $Y=0.6
+ $X2=2.07 $Y2=0.815
r55 19 31 3.97509 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=0.445 $Y=0.475
+ $X2=0.28 $Y2=0.475
r56 19 21 35.2648 $w=2.48e-07 $l=7.65e-07 $layer=LI1_cond $X=0.445 $Y=0.475
+ $X2=1.21 $Y2=0.475
r57 18 33 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.985 $Y=0.475
+ $X2=2.07 $Y2=0.475
r58 18 21 35.7257 $w=2.48e-07 $l=7.75e-07 $layer=LI1_cond $X=1.985 $Y=0.475
+ $X2=1.21 $Y2=0.475
r59 5 28 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=3.65
+ $Y=0.37 $X2=3.79 $Y2=0.95
r60 4 26 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=2.79
+ $Y=0.37 $X2=2.93 $Y2=0.95
r61 3 35 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=1.93
+ $Y=0.37 $X2=2.07 $Y2=0.965
r62 3 33 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1.93
+ $Y=0.37 $X2=2.07 $Y2=0.515
r63 2 21 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1.07
+ $Y=0.37 $X2=1.21 $Y2=0.515
r64 1 31 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__O2111AI_4%A_472_74# 1 2 3 4 22 23
c28 23 0 8.0658e-20 $X=5.475 $Y=0.515
c29 22 0 2.50688e-19 $X=5.64 $Y=0.515
r30 22 23 5.91831 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=5.64 $Y=0.515
+ $X2=5.475 $Y2=0.515
r31 20 23 27.1508 $w=2.93e-07 $l=6.95e-07 $layer=LI1_cond $X=4.78 $Y=0.497
+ $X2=5.475 $Y2=0.497
r32 18 20 55.4735 $w=2.93e-07 $l=1.42e-06 $layer=LI1_cond $X=3.36 $Y=0.497
+ $X2=4.78 $Y2=0.497
r33 15 18 33.5966 $w=2.93e-07 $l=8.6e-07 $layer=LI1_cond $X=2.5 $Y=0.497
+ $X2=3.36 $Y2=0.497
r34 4 22 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=5.5
+ $Y=0.37 $X2=5.64 $Y2=0.515
r35 3 20 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=4.64
+ $Y=0.37 $X2=4.78 $Y2=0.515
r36 2 18 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.22
+ $Y=0.37 $X2=3.36 $Y2=0.515
r37 1 15 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.36
+ $Y=0.37 $X2=2.5 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__O2111AI_4%A_841_74# 1 2 3 4 5 6 7 24 27 30 32 36 38
+ 42 44 48 50 54 59 60 62 63 64 65
c108 59 0 3.65531e-19 $X=4.515 $Y=0.972
c109 30 0 1.61888e-19 $X=6.14 $Y=0.515
r110 59 60 21.8141 $w=2.78e-07 $l=5.3e-07 $layer=LI1_cond $X=4.515 $Y=0.99
+ $X2=5.045 $Y2=0.99
r111 57 59 6.20639 $w=3.13e-07 $l=1.65e-07 $layer=LI1_cond $X=4.35 $Y=0.972
+ $X2=4.515 $Y2=0.972
r112 52 54 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=9.84 $Y=1.01
+ $X2=9.84 $Y2=0.515
r113 51 65 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.025 $Y=1.095
+ $X2=8.9 $Y2=1.095
r114 50 52 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=9.715 $Y=1.095
+ $X2=9.84 $Y2=1.01
r115 50 51 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=9.715 $Y=1.095
+ $X2=9.025 $Y2=1.095
r116 46 65 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.9 $Y=1.01
+ $X2=8.9 $Y2=1.095
r117 46 48 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=8.9 $Y=1.01
+ $X2=8.9 $Y2=0.515
r118 45 64 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.095 $Y=1.095
+ $X2=7.97 $Y2=1.095
r119 44 65 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.775 $Y=1.095
+ $X2=8.9 $Y2=1.095
r120 44 45 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=8.775 $Y=1.095
+ $X2=8.095 $Y2=1.095
r121 40 64 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.97 $Y=1.01
+ $X2=7.97 $Y2=1.095
r122 40 42 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=7.97 $Y=1.01
+ $X2=7.97 $Y2=0.515
r123 39 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.155 $Y=1.095
+ $X2=7.07 $Y2=1.095
r124 38 64 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.845 $Y=1.095
+ $X2=7.97 $Y2=1.095
r125 38 39 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=7.845 $Y=1.095
+ $X2=7.155 $Y2=1.095
r126 34 63 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.07 $Y=1.01
+ $X2=7.07 $Y2=1.095
r127 34 36 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=7.07 $Y=1.01
+ $X2=7.07 $Y2=0.515
r128 33 62 6.46576 $w=2.5e-07 $l=2.0106e-07 $layer=LI1_cond $X=6.305 $Y=1.095
+ $X2=6.14 $Y2=1.015
r129 32 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.985 $Y=1.095
+ $X2=7.07 $Y2=1.095
r130 32 33 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=6.985 $Y=1.095
+ $X2=6.305 $Y2=1.095
r131 28 62 0.364692 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=6.14 $Y=0.85
+ $X2=6.14 $Y2=1.015
r132 28 30 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=6.14 $Y=0.85
+ $X2=6.14 $Y2=0.515
r133 27 60 6.05995 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=5.21 $Y=1.015
+ $X2=5.045 $Y2=1.015
r134 24 62 6.46576 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=5.975 $Y=1.015
+ $X2=6.14 $Y2=1.015
r135 24 27 26.7157 $w=3.28e-07 $l=7.65e-07 $layer=LI1_cond $X=5.975 $Y=1.015
+ $X2=5.21 $Y2=1.015
r136 7 54 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.66
+ $Y=0.37 $X2=9.8 $Y2=0.515
r137 6 48 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.72
+ $Y=0.37 $X2=8.86 $Y2=0.515
r138 5 42 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.79
+ $Y=0.37 $X2=7.93 $Y2=0.515
r139 4 36 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.93
+ $Y=0.37 $X2=7.07 $Y2=0.515
r140 3 62 182 $w=1.7e-07 $l=6.9208e-07 $layer=licon1_NDIFF $count=1 $X=5.93
+ $Y=0.37 $X2=6.14 $Y2=0.965
r141 3 30 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=5.93
+ $Y=0.37 $X2=6.14 $Y2=0.515
r142 2 27 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=5.07
+ $Y=0.37 $X2=5.21 $Y2=0.95
r143 1 57 182 $w=1.7e-07 $l=6.4846e-07 $layer=licon1_NDIFF $count=1 $X=4.205
+ $Y=0.37 $X2=4.35 $Y2=0.95
.ends

.subckt PM_SKY130_FD_SC_LS__O2111AI_4%VGND 1 2 3 4 15 19 23 27 29 31 36 41 46 53
+ 54 57 60 63 66
r103 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r104 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r105 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r106 57 58 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r107 54 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0 $X2=9.36
+ $Y2=0
r108 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r109 51 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.535 $Y=0 $X2=9.37
+ $Y2=0
r110 51 53 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=9.535 $Y=0
+ $X2=9.84 $Y2=0
r111 50 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=9.36
+ $Y2=0
r112 50 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=8.4
+ $Y2=0
r113 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r114 47 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.595 $Y=0 $X2=8.43
+ $Y2=0
r115 47 49 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=8.595 $Y=0
+ $X2=8.88 $Y2=0
r116 46 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.205 $Y=0 $X2=9.37
+ $Y2=0
r117 46 49 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=9.205 $Y=0
+ $X2=8.88 $Y2=0
r118 45 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.4
+ $Y2=0
r119 45 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=7.44
+ $Y2=0
r120 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r121 42 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.665 $Y=0 $X2=7.5
+ $Y2=0
r122 42 44 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=7.665 $Y=0
+ $X2=7.92 $Y2=0
r123 41 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.265 $Y=0 $X2=8.43
+ $Y2=0
r124 41 44 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=8.265 $Y=0 $X2=7.92
+ $Y2=0
r125 40 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r126 40 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=6.48
+ $Y2=0
r127 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r128 37 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.805 $Y=0 $X2=6.64
+ $Y2=0
r129 37 39 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=6.805 $Y=0
+ $X2=6.96 $Y2=0
r130 36 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.335 $Y=0 $X2=7.5
+ $Y2=0
r131 36 39 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=7.335 $Y=0
+ $X2=6.96 $Y2=0
r132 33 34 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r133 31 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.475 $Y=0 $X2=6.64
+ $Y2=0
r134 31 33 406.775 $w=1.68e-07 $l=6.235e-06 $layer=LI1_cond $X=6.475 $Y=0
+ $X2=0.24 $Y2=0
r135 29 58 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=6.48 $Y2=0
r136 29 34 1.33793 $w=4.9e-07 $l=4.8e-06 $layer=MET1_cond $X=5.04 $Y=0 $X2=0.24
+ $Y2=0
r137 25 66 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.37 $Y=0.085
+ $X2=9.37 $Y2=0
r138 25 27 19.9058 $w=3.28e-07 $l=5.7e-07 $layer=LI1_cond $X=9.37 $Y=0.085
+ $X2=9.37 $Y2=0.655
r139 21 63 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.43 $Y=0.085
+ $X2=8.43 $Y2=0
r140 21 23 19.9058 $w=3.28e-07 $l=5.7e-07 $layer=LI1_cond $X=8.43 $Y=0.085
+ $X2=8.43 $Y2=0.655
r141 17 60 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.5 $Y=0.085 $X2=7.5
+ $Y2=0
r142 17 19 19.9058 $w=3.28e-07 $l=5.7e-07 $layer=LI1_cond $X=7.5 $Y=0.085
+ $X2=7.5 $Y2=0.655
r143 13 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.64 $Y=0.085
+ $X2=6.64 $Y2=0
r144 13 15 19.9058 $w=3.28e-07 $l=5.7e-07 $layer=LI1_cond $X=6.64 $Y=0.085
+ $X2=6.64 $Y2=0.655
r145 4 27 182 $w=1.7e-07 $l=3.4803e-07 $layer=licon1_NDIFF $count=1 $X=9.23
+ $Y=0.37 $X2=9.37 $Y2=0.655
r146 3 23 182 $w=1.7e-07 $l=3.756e-07 $layer=licon1_NDIFF $count=1 $X=8.22
+ $Y=0.37 $X2=8.43 $Y2=0.655
r147 2 19 182 $w=1.7e-07 $l=3.4803e-07 $layer=licon1_NDIFF $count=1 $X=7.36
+ $Y=0.37 $X2=7.5 $Y2=0.655
r148 1 15 182 $w=1.7e-07 $l=3.756e-07 $layer=licon1_NDIFF $count=1 $X=6.43
+ $Y=0.37 $X2=6.64 $Y2=0.655
.ends

