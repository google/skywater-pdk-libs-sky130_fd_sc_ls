* File: sky130_fd_sc_ls__sdfstp_1.spice
* Created: Wed Sep  2 11:27:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__sdfstp_1.pex.spice"
.subckt sky130_fd_sc_ls__sdfstp_1  VNB VPB SCE D SCD CLK SET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* SET_B	SET_B
* CLK	CLK
* SCD	SCD
* D	D
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1020 N_VGND_M1020_d N_SCE_M1020_g N_A_27_464#_M1020_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0819 AS=0.1197 PD=0.81 PS=1.41 NRD=19.992 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1001 A_238_74# N_A_27_464#_M1001_g N_VGND_M1020_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0819 PD=0.66 PS=0.81 NRD=18.564 NRS=11.424 M=1 R=2.8 SA=75000.7
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1025 N_A_289_464#_M1025_d N_D_M1025_g A_238_74# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0504 PD=0.7 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.1
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1002 A_402_74# N_SCE_M1002_g N_A_289_464#_M1025_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0588 PD=0.66 PS=0.7 NRD=18.564 NRS=0 M=1 R=2.8 SA=75001.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1000 N_VGND_M1000_d N_SCD_M1000_g A_402_74# VNB NSHORT L=0.15 W=0.42 AD=0.1197
+ AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75002 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_CLK_M1003_g N_A_599_74#_M1003_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1554 AS=0.2109 PD=1.16 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.8 A=0.111 P=1.78 MULT=1
MM1015 N_A_800_74#_M1015_d N_A_599_74#_M1015_g N_VGND_M1003_d VNB NSHORT L=0.15
+ W=0.74 AD=0.2109 AS=0.1554 PD=2.05 PS=1.16 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75000.8 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1014 N_A_998_81#_M1014_d N_A_599_74#_M1014_g N_A_289_464#_M1014_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.1281 AS=0.1197 PD=1.03 PS=1.41 NRD=94.284 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1012 A_1150_81# N_A_800_74#_M1012_g N_A_998_81#_M1014_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.1281 PD=0.66 PS=1.03 NRD=18.564 NRS=0 M=1 R=2.8 SA=75001
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1010 N_VGND_M1010_d N_A_1198_55#_M1010_g A_1150_81# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1023 A_1426_118# N_A_998_81#_M1023_g N_A_1198_55#_M1023_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75003.3 A=0.063 P=1.14 MULT=1
MM1013 N_VGND_M1013_d N_SET_B_M1013_g A_1426_118# VNB NSHORT L=0.15 W=0.42
+ AD=0.186187 AS=0.0504 PD=1.10943 PS=0.66 NRD=12.132 NRS=18.564 M=1 R=2.8
+ SA=75000.6 SB=75002.9 A=0.063 P=1.14 MULT=1
MM1038 A_1686_74# N_A_998_81#_M1038_g N_VGND_M1013_d VNB NSHORT L=0.15 W=0.64
+ AD=0.0768 AS=0.283713 PD=0.88 PS=1.69057 NRD=12.18 NRS=0 M=1 R=4.26667
+ SA=75001.2 SB=75002.4 A=0.096 P=1.58 MULT=1
MM1039 N_A_1764_74#_M1039_d N_A_800_74#_M1039_g A_1686_74# VNB NSHORT L=0.15
+ W=0.64 AD=0.214158 AS=0.0768 PD=1.47321 PS=0.88 NRD=20.616 NRS=12.18 M=1
+ R=4.26667 SA=75001.6 SB=75002 A=0.096 P=1.58 MULT=1
MM1031 A_1910_74# N_A_599_74#_M1031_g N_A_1764_74#_M1039_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.140542 PD=0.66 PS=0.966792 NRD=18.564 NRS=54.996 M=1
+ R=2.8 SA=75002.2 SB=75002.1 A=0.063 P=1.14 MULT=1
MM1006 A_1988_74# N_A_1958_48#_M1006_g A_1910_74# VNB NSHORT L=0.15 W=0.42
+ AD=0.1596 AS=0.0504 PD=1.18 PS=0.66 NRD=92.856 NRS=18.564 M=1 R=2.8 SA=75002.5
+ SB=75001.7 A=0.063 P=1.14 MULT=1
MM1018 N_VGND_M1018_d N_SET_B_M1018_g A_1988_74# VNB NSHORT L=0.15 W=0.42
+ AD=0.0882 AS=0.1596 PD=0.84 PS=1.18 NRD=0 NRS=92.856 M=1 R=2.8 SA=75003.5
+ SB=75000.8 A=0.063 P=1.14 MULT=1
MM1033 N_A_1958_48#_M1033_d N_A_1764_74#_M1033_g N_VGND_M1018_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.1197 AS=0.0882 PD=1.41 PS=0.84 NRD=0 NRS=39.996 M=1 R=2.8
+ SA=75004 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1029 N_VGND_M1029_d N_A_1764_74#_M1029_g N_A_2395_112#_M1029_s VNB NSHORT
+ L=0.15 W=0.55 AD=0.129591 AS=0.385 PD=0.997674 PS=2.5 NRD=18 NRS=140.724 M=1
+ R=3.66667 SA=75000.6 SB=75000.8 A=0.0825 P=1.4 MULT=1
MM1019 N_Q_M1019_d N_A_2395_112#_M1019_g N_VGND_M1029_d VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.174359 PD=2.05 PS=1.34233 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75001 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1026 N_VPWR_M1026_d N_SCE_M1026_g N_A_27_464#_M1026_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.096 AS=0.1856 PD=0.94 PS=1.86 NRD=3.0732 NRS=3.0732 M=1 R=4.26667
+ SA=75000.2 SB=75002.2 A=0.096 P=1.58 MULT=1
MM1027 A_205_464# N_SCE_M1027_g N_VPWR_M1026_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0864 AS=0.096 PD=0.91 PS=0.94 NRD=24.625 NRS=3.0732 M=1 R=4.26667
+ SA=75000.7 SB=75001.8 A=0.096 P=1.58 MULT=1
MM1021 N_A_289_464#_M1021_d N_D_M1021_g A_205_464# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1536 AS=0.0864 PD=1.12 PS=0.91 NRD=30.7714 NRS=24.625 M=1 R=4.26667
+ SA=75001.1 SB=75001.4 A=0.096 P=1.58 MULT=1
MM1005 A_415_464# N_A_27_464#_M1005_g N_A_289_464#_M1021_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0864 AS=0.1536 PD=0.91 PS=1.12 NRD=24.625 NRS=30.7714 M=1
+ R=4.26667 SA=75001.7 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1035 N_VPWR_M1035_d N_SCD_M1035_g A_415_464# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.2954 AS=0.0864 PD=2.4 PS=0.91 NRD=30.7714 NRS=24.625 M=1 R=4.26667
+ SA=75002.1 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1017 N_VPWR_M1017_d N_CLK_M1017_g N_A_599_74#_M1017_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.6 A=0.168 P=2.54 MULT=1
MM1024 N_A_800_74#_M1024_d N_A_599_74#_M1024_g N_VPWR_M1017_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.3076 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1030 N_A_998_81#_M1030_d N_A_800_74#_M1030_g N_A_289_464#_M1030_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0735 AS=0.1239 PD=0.77 PS=1.43 NRD=28.1316 NRS=4.6886 M=1
+ R=2.8 SA=75000.2 SB=75003.1 A=0.063 P=1.14 MULT=1
MM1032 A_1128_457# N_A_599_74#_M1032_g N_A_998_81#_M1030_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.07665 AS=0.0735 PD=0.785 PS=0.77 NRD=59.7895 NRS=4.6886 M=1 R=2.8
+ SA=75000.7 SB=75002.6 A=0.063 P=1.14 MULT=1
MM1007 N_VPWR_M1007_d N_A_1198_55#_M1007_g A_1128_457# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1649 AS=0.07665 PD=1.295 PS=0.785 NRD=158.349 NRS=59.7895 M=1 R=2.8
+ SA=75001.2 SB=75002.1 A=0.063 P=1.14 MULT=1
MM1022 N_A_1198_55#_M1022_d N_A_998_81#_M1022_g N_VPWR_M1007_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0693 AS=0.1649 PD=0.75 PS=1.295 NRD=18.7544 NRS=158.349 M=1
+ R=2.8 SA=75002 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1011 N_VPWR_M1011_d N_SET_B_M1011_g N_A_1198_55#_M1022_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.0693 PD=0.90507 PS=0.75 NRD=112.566 NRS=4.6886 M=1 R=2.8
+ SA=75002.4 SB=75000.9 A=0.063 P=1.14 MULT=1
MM1008 N_A_1610_341#_M1008_d N_A_998_81#_M1008_g N_VPWR_M1011_d VPB PHIGHVT
+ L=0.15 W=1 AD=0.285 AS=0.265 PD=2.57 PS=2.15493 NRD=1.9503 NRS=1.9503 M=1
+ R=6.66667 SA=75001.4 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1036 N_A_1764_74#_M1036_d N_A_800_74#_M1036_g N_A_1721_374#_M1036_s VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.096393 AS=0.2584 PD=0.834085 PS=3.07 NRD=53.9386
+ NRS=262.778 M=1 R=2.8 SA=75000.2 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1037 N_A_1610_341#_M1037_d N_A_599_74#_M1037_g N_A_1764_74#_M1036_d VPB
+ PHIGHVT L=0.15 W=1 AD=0.28 AS=0.229507 PD=2.56 PS=1.98592 NRD=1.9503
+ NRS=2.9353 M=1 R=6.66667 SA=75000.4 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1009 N_VPWR_M1009_d N_A_1958_48#_M1009_g N_A_1721_374#_M1009_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.063 AS=0.1197 PD=0.72 PS=1.41 NRD=4.6886 NRS=4.6886 M=1
+ R=2.8 SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1016 N_A_1764_74#_M1016_d N_SET_B_M1016_g N_VPWR_M1009_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1197 AS=0.063 PD=1.41 PS=0.72 NRD=4.6886 NRS=4.6886 M=1 R=2.8
+ SA=75000.7 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1034 N_VPWR_M1034_d N_A_1764_74#_M1034_g N_A_1958_48#_M1034_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.1197 AS=0.1197 PD=1.41 PS=1.41 NRD=4.6886 NRS=4.6886 M=1
+ R=2.8 SA=75000.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1004 N_VPWR_M1004_d N_A_1764_74#_M1004_g N_A_2395_112#_M1004_s VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.1596 AS=0.2394 PD=1.26429 PS=2.25 NRD=14.0658 NRS=2.3443
+ M=1 R=5.6 SA=75000.2 SB=75000.7 A=0.126 P=1.98 MULT=1
MM1028 N_Q_M1028_d N_A_2395_112#_M1028_g N_VPWR_M1004_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.3192 AS=0.2128 PD=2.81 PS=1.68571 NRD=1.7533 NRS=2.6201 M=1
+ R=7.46667 SA=75000.6 SB=75000.2 A=0.168 P=2.54 MULT=1
DX40_noxref VNB VPB NWDIODE A=26.7411 P=32.59
*
.include "sky130_fd_sc_ls__sdfstp_1.pxi.spice"
*
.ends
*
*
