* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__mux2_4 A0 A1 S VGND VNB VPB VPWR X
M1000 a_937_119# a_27_368# VGND VNB nshort w=640000u l=150000u
+  ad=3.712e+11p pd=3.72e+06u as=1.76805e+12p ps=1.249e+07u
M1001 X a_193_241# VGND VNB nshort w=740000u l=150000u
+  ad=4.44e+11p pd=4.16e+06u as=0p ps=0u
M1002 VGND a_27_368# a_937_119# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPWR S a_722_391# VPB phighvt w=1e+06u l=150000u
+  ad=2.49868e+12p pd=1.636e+07u as=6e+11p ps=5.2e+06u
M1004 VPWR a_27_368# a_936_391# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=6e+11p ps=5.2e+06u
M1005 a_193_241# A1 a_936_391# VPB phighvt w=1e+06u l=150000u
+  ad=9.85e+11p pd=7.97e+06u as=0p ps=0u
M1006 VPWR a_193_241# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=1.13255e+12p ps=6.91e+06u
M1007 a_936_391# a_27_368# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND a_193_241# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_193_241# A1 a_709_119# VNB nshort w=640000u l=150000u
+  ad=9.216e+11p pd=6.72e+06u as=4.224e+11p ps=3.88e+06u
M1010 X a_193_241# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 X a_193_241# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR S a_27_368# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.95e+11p ps=2.59e+06u
M1013 a_937_119# A0 a_193_241# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR a_193_241# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_722_391# A0 a_193_241# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND a_193_241# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_193_241# A0 a_937_119# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 X a_193_241# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_722_391# S VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND S a_709_119# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_709_119# A1 a_193_241# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_193_241# A0 a_722_391# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_709_119# S VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_936_391# A1 a_193_241# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VGND S a_27_368# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
.ends
