# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ls__o2bb2ai_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ls__o2bb2ai_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.08000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1_N
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.350000 1.935000 1.780000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.225000 1.350000 3.235000 1.780000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.150000 1.350000 9.955000 1.780000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.885000 1.350000 7.640000 1.780000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  1.758400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.155000 1.800000 5.715000 1.950000 ;
        RECT 4.155000 1.950000 7.725000 1.970000 ;
        RECT 4.155000 1.970000 4.485000 2.980000 ;
        RECT 4.695000 0.595000 5.025000 0.960000 ;
        RECT 4.695000 0.960000 5.885000 1.130000 ;
        RECT 5.055000 1.970000 7.725000 2.120000 ;
        RECT 5.055000 2.120000 5.635000 2.150000 ;
        RECT 5.055000 2.150000 5.305000 2.980000 ;
        RECT 5.545000 0.595000 5.885000 0.960000 ;
        RECT 5.545000 1.130000 5.715000 1.800000 ;
        RECT 6.495000 2.120000 6.825000 2.735000 ;
        RECT 7.395000 2.120000 7.725000 2.735000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 10.080000 0.085000 ;
        RECT 0.545000  0.085000  0.875000 0.840000 ;
        RECT 1.415000  0.085000  1.745000 0.840000 ;
        RECT 6.415000  0.085000  6.745000 0.830000 ;
        RECT 7.345000  0.085000  7.675000 0.830000 ;
        RECT 8.275000  0.085000  8.605000 0.830000 ;
        RECT 9.205000  0.085000  9.535000 0.830000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
        RECT 6.395000 -0.085000 6.565000 0.085000 ;
        RECT 6.875000 -0.085000 7.045000 0.085000 ;
        RECT 7.355000 -0.085000 7.525000 0.085000 ;
        RECT 7.835000 -0.085000 8.005000 0.085000 ;
        RECT 8.315000 -0.085000 8.485000 0.085000 ;
        RECT 8.795000 -0.085000 8.965000 0.085000 ;
        RECT 9.275000 -0.085000 9.445000 0.085000 ;
        RECT 9.755000 -0.085000 9.925000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.080000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 10.080000 3.415000 ;
        RECT 0.105000 1.950000  0.355000 3.245000 ;
        RECT 1.085000 2.290000  1.255000 3.245000 ;
        RECT 1.985000 2.290000  2.155000 3.245000 ;
        RECT 2.885000 2.290000  3.055000 3.245000 ;
        RECT 3.785000 1.820000  3.955000 3.245000 ;
        RECT 4.685000 2.140000  4.855000 3.245000 ;
        RECT 5.505000 2.320000  5.835000 3.245000 ;
        RECT 8.295000 2.290000  8.560000 3.245000 ;
        RECT 9.260000 2.290000  9.465000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
        RECT 6.395000 3.245000 6.565000 3.415000 ;
        RECT 6.875000 3.245000 7.045000 3.415000 ;
        RECT 7.355000 3.245000 7.525000 3.415000 ;
        RECT 7.835000 3.245000 8.005000 3.415000 ;
        RECT 8.315000 3.245000 8.485000 3.415000 ;
        RECT 8.795000 3.245000 8.965000 3.415000 ;
        RECT 9.275000 3.245000 9.445000 3.415000 ;
        RECT 9.755000 3.245000 9.925000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 10.080000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.115000 0.350000 0.365000 1.010000 ;
      RECT 0.115000 1.010000 2.095000 1.180000 ;
      RECT 0.555000 1.950000 3.585000 2.120000 ;
      RECT 0.555000 2.120000 0.885000 2.980000 ;
      RECT 1.055000 0.350000 1.235000 1.010000 ;
      RECT 1.455000 2.120000 1.785000 2.980000 ;
      RECT 1.925000 0.255000 4.035000 0.425000 ;
      RECT 1.925000 0.425000 2.095000 1.010000 ;
      RECT 2.275000 0.595000 2.605000 1.010000 ;
      RECT 2.275000 1.010000 3.605000 1.180000 ;
      RECT 2.355000 2.120000 2.685000 2.980000 ;
      RECT 2.775000 0.425000 3.105000 0.840000 ;
      RECT 3.255000 2.120000 3.585000 2.980000 ;
      RECT 3.275000 0.595000 3.605000 1.010000 ;
      RECT 3.415000 1.180000 3.605000 1.300000 ;
      RECT 3.415000 1.300000 5.375000 1.630000 ;
      RECT 3.415000 1.630000 3.585000 1.950000 ;
      RECT 3.785000 0.425000 4.035000 1.130000 ;
      RECT 4.265000 0.255000 6.235000 0.425000 ;
      RECT 4.265000 0.425000 4.515000 1.130000 ;
      RECT 5.205000 0.425000 5.375000 0.790000 ;
      RECT 6.045000 2.290000 6.310000 2.905000 ;
      RECT 6.045000 2.905000 8.110000 3.075000 ;
      RECT 6.065000 0.425000 6.235000 1.010000 ;
      RECT 6.065000 1.010000 9.965000 1.180000 ;
      RECT 6.915000 0.350000 7.165000 1.010000 ;
      RECT 7.010000 2.290000 7.210000 2.905000 ;
      RECT 7.845000 0.350000 8.095000 1.010000 ;
      RECT 7.910000 1.950000 9.975000 2.120000 ;
      RECT 7.910000 2.120000 8.110000 2.905000 ;
      RECT 8.745000 2.120000 9.075000 2.980000 ;
      RECT 8.785000 0.350000 9.035000 1.010000 ;
      RECT 9.645000 2.120000 9.975000 2.980000 ;
      RECT 9.715000 0.350000 9.965000 1.010000 ;
  END
END sky130_fd_sc_ls__o2bb2ai_4
