* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__nand3_4 A B C VGND VNB VPB VPWR Y
M1000 a_456_82# C VGND VNB nshort w=740000u l=150000u
+  ad=8.288e+11p pd=8.16e+06u as=6.142e+11p ps=6.1e+06u
M1001 VGND C a_456_82# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 VPWR C Y VPB phighvt w=1.12e+06u l=150000u
+  ad=3.6904e+12p pd=1.555e+07u as=1.5904e+12p ps=9.56e+06u
M1003 a_27_82# B a_456_82# VNB nshort w=740000u l=150000u
+  ad=1.0121e+12p pd=1.018e+07u as=0p ps=0u
M1004 a_456_82# B a_27_82# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y A a_27_82# VNB nshort w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=0p ps=0u
M1006 VPWR A Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND C a_456_82# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y B VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_27_82# B a_456_82# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_456_82# C VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Y A VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_27_82# A Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 Y A a_27_82# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR B Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_456_82# B a_27_82# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_27_82# A Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 Y C VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
