# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ls__and2_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_ls__and2_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.444000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.925000 1.450000 3.255000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.444000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.255000 1.345000 2.755000 1.780000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  1.219800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545000 0.475000 0.795000 1.005000 ;
        RECT 0.545000 1.005000 1.725000 1.175000 ;
        RECT 0.545000 1.175000 0.795000 1.550000 ;
        RECT 0.545000 1.550000 0.835000 1.845000 ;
        RECT 0.545000 1.845000 1.715000 2.015000 ;
        RECT 0.545000 2.015000 0.815000 2.980000 ;
        RECT 1.465000 2.015000 1.715000 2.980000 ;
        RECT 1.475000 0.475000 1.725000 1.005000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.115000  0.085000 0.365000 1.255000 ;
      RECT 0.115000  1.820000 0.365000 3.245000 ;
      RECT 0.975000  0.085000 1.305000 0.835000 ;
      RECT 1.005000  1.345000 2.055000 1.675000 ;
      RECT 1.015000  2.185000 1.265000 3.245000 ;
      RECT 1.885000  1.675000 2.055000 1.950000 ;
      RECT 1.885000  1.950000 3.670000 2.120000 ;
      RECT 1.935000  2.290000 2.265000 3.245000 ;
      RECT 1.985000  0.085000 2.315000 1.175000 ;
      RECT 2.470000  2.120000 2.800000 2.905000 ;
      RECT 2.495000  0.255000 3.675000 0.425000 ;
      RECT 2.495000  0.425000 2.825000 1.175000 ;
      RECT 2.970000  2.290000 3.300000 3.245000 ;
      RECT 2.995000  0.595000 3.325000 1.110000 ;
      RECT 2.995000  1.110000 3.670000 1.280000 ;
      RECT 3.500000  1.280000 3.670000 1.950000 ;
      RECT 3.500000  2.120000 3.670000 2.905000 ;
      RECT 3.505000  0.425000 3.675000 0.940000 ;
      RECT 3.870000  2.025000 4.200000 3.245000 ;
      RECT 3.875000  0.085000 4.205000 1.255000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_ls__and2_4
END LIBRARY
