* File: sky130_fd_sc_ls__decaphe_18.pex.spice
* Created: Fri Aug 28 13:11:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__DECAPHE_18%VPWR 1 8 12 13 15 23 24 28 29 44 48 53
r24 48 53 1.0564 $w=4.9e-07 $l=3.79e-06 $layer=MET1_cond $X=8.4 $Y=3.33 $X2=4.61
+ $Y2=3.33
r25 47 48 1.03333 $w=1.7e-07 $l=1.53e-06 $layer=mcon $count=9 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r26 44 47 0.136925 $w=1.782e-06 $l=2e-08 $layer=LI1_cond $X=8.38 $Y=2.332
+ $X2=8.4 $Y2=2.332
r27 34 37 0.136925 $w=1.782e-06 $l=2e-08 $layer=LI1_cond $X=0.24 $Y=2.332
+ $X2=0.26 $Y2=2.332
r28 34 35 1.03333 $w=1.7e-07 $l=1.53e-06 $layer=mcon $count=9 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r29 32 44 8.62626 $w=1.782e-06 $l=1.26e-06 $layer=LI1_cond $X=7.12 $Y=2.332
+ $X2=8.38 $Y2=2.332
r30 31 32 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.12
+ $Y=1.335 $X2=7.12 $Y2=1.335
r31 27 32 12.0494 $w=1.782e-06 $l=1.76e-06 $layer=LI1_cond $X=5.36 $Y=2.332
+ $X2=7.12 $Y2=2.332
r32 26 29 9.23771 $w=1.395e-06 $l=1.65e-07 $layer=POLY_cond $X=5.36 $Y=0.802
+ $X2=5.525 $Y2=0.802
r33 26 28 21.2799 $w=1.395e-06 $l=5.05e-07 $layer=POLY_cond $X=5.36 $Y=0.802
+ $X2=4.855 $Y2=0.802
r34 26 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.36
+ $Y=1.335 $X2=5.36 $Y2=1.335
r35 22 27 12.0494 $w=1.782e-06 $l=1.76e-06 $layer=LI1_cond $X=3.6 $Y=2.332
+ $X2=5.36 $Y2=2.332
r36 21 24 9.23771 $w=1.395e-06 $l=1.65e-07 $layer=POLY_cond $X=3.6 $Y=0.802
+ $X2=3.765 $Y2=0.802
r37 21 23 21.2799 $w=1.395e-06 $l=5.05e-07 $layer=POLY_cond $X=3.6 $Y=0.802
+ $X2=3.095 $Y2=0.802
r38 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.6
+ $Y=1.335 $X2=3.6 $Y2=1.335
r39 19 22 12.0494 $w=1.782e-06 $l=1.76e-06 $layer=LI1_cond $X=1.84 $Y=2.332
+ $X2=3.6 $Y2=2.332
r40 19 37 10.8171 $w=1.782e-06 $l=1.58e-06 $layer=LI1_cond $X=1.84 $Y=2.332
+ $X2=0.26 $Y2=2.332
r41 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.84
+ $Y=1.335 $X2=1.84 $Y2=1.335
r42 15 53 0.0808331 $w=4.9e-07 $l=2.9e-07 $layer=MET1_cond $X=4.32 $Y=3.33
+ $X2=4.61 $Y2=3.33
r43 15 35 1.13724 $w=4.9e-07 $l=4.08e-06 $layer=MET1_cond $X=4.32 $Y=3.33
+ $X2=0.24 $Y2=3.33
r44 13 31 21.4636 $w=1.182e-06 $l=5.88154e-07 $layer=POLY_cond $X=6.615 $Y=0.622
+ $X2=7.12 $Y2=0.802
r45 13 29 54.1495 $w=1.035e-06 $l=1.09e-06 $layer=POLY_cond $X=6.615 $Y=0.622
+ $X2=5.525 $Y2=0.622
r46 12 28 26.578 $w=1.035e-06 $l=5.35e-07 $layer=POLY_cond $X=4.32 $Y=0.622
+ $X2=4.855 $Y2=0.622
r47 12 24 27.5715 $w=1.035e-06 $l=5.55e-07 $layer=POLY_cond $X=4.32 $Y=0.622
+ $X2=3.765 $Y2=0.622
r48 8 18 7.60645 $w=1.184e-06 $l=2.49199e-07 $layer=POLY_cond $X=2.005 $Y=0.622
+ $X2=1.84 $Y2=0.802
r49 8 23 54.1495 $w=1.035e-06 $l=1.09e-06 $layer=POLY_cond $X=2.005 $Y=0.622
+ $X2=3.095 $Y2=0.622
r50 1 44 400 $w=1.7e-07 $l=1.17556e-06 $layer=licon1_PDIFF $count=1 $X=8.245
+ $Y=1.84 $X2=8.38 $Y2=2.95
r51 1 44 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=8.245
+ $Y=1.84 $X2=8.38 $Y2=1.985
r52 1 37 400 $w=1.7e-07 $l=1.17083e-06 $layer=licon1_PDIFF $count=1 $X=8.245
+ $Y=1.84 $X2=0.26 $Y2=2.95
r53 1 37 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=8.245
+ $Y=1.84 $X2=0.26 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_LS__DECAPHE_18%VGND 1 7 16 21 40 43 49
r18 43 49 1.04247 $w=4.9e-07 $l=3.74e-06 $layer=MET1_cond $X=8.4 $Y=0 $X2=4.66
+ $Y2=0
r19 42 43 1.09412 $w=1.7e-07 $l=1.445e-06 $layer=mcon $count=8 $X=8.4 $Y=0
+ $X2=8.4 $Y2=0
r20 40 42 0.174535 $w=1.398e-06 $l=2e-08 $layer=LI1_cond $X=8.38 $Y=0.757
+ $X2=8.4 $Y2=0.757
r21 32 33 1.09412 $w=1.7e-07 $l=1.445e-06 $layer=mcon $count=8 $X=0.72 $Y=0
+ $X2=0.72 $Y2=0
r22 30 32 4.01431 $w=1.398e-06 $l=4.6e-07 $layer=LI1_cond $X=0.26 $Y=0.757
+ $X2=0.72 $Y2=0.757
r23 28 33 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r24 27 30 0.174535 $w=1.398e-06 $l=2e-08 $layer=LI1_cond $X=0.24 $Y=0.757
+ $X2=0.26 $Y2=0.757
r25 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r26 25 40 3.31617 $w=1.398e-06 $l=3.8e-07 $layer=LI1_cond $X=8 $Y=0.757 $X2=8.38
+ $Y2=0.757
r27 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8 $Y=1.515
+ $X2=8 $Y2=1.515
r28 22 25 15.3591 $w=1.398e-06 $l=1.76e-06 $layer=LI1_cond $X=6.24 $Y=0.757
+ $X2=8 $Y2=0.757
r29 21 24 50.646 $w=1.675e-06 $l=1.76e-06 $layer=POLY_cond $X=6.24 $Y=2.287
+ $X2=8 $Y2=2.287
r30 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.24
+ $Y=1.515 $X2=6.24 $Y2=1.515
r31 19 22 15.3591 $w=1.398e-06 $l=1.76e-06 $layer=LI1_cond $X=4.48 $Y=0.757
+ $X2=6.24 $Y2=0.757
r32 18 21 50.646 $w=1.675e-06 $l=1.76e-06 $layer=POLY_cond $X=4.48 $Y=2.287
+ $X2=6.24 $Y2=2.287
r33 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.48
+ $Y=1.515 $X2=4.48 $Y2=1.515
r34 16 18 4.60418 $w=1.675e-06 $l=1.6e-07 $layer=POLY_cond $X=4.32 $Y=2.287
+ $X2=4.48 $Y2=2.287
r35 14 19 15.3591 $w=1.398e-06 $l=1.76e-06 $layer=LI1_cond $X=2.72 $Y=0.757
+ $X2=4.48 $Y2=0.757
r36 13 16 46.0418 $w=1.675e-06 $l=1.6e-06 $layer=POLY_cond $X=2.72 $Y=2.287
+ $X2=4.32 $Y2=2.287
r37 13 14 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.72
+ $Y=1.515 $X2=2.72 $Y2=1.515
r38 11 14 15.3591 $w=1.398e-06 $l=1.76e-06 $layer=LI1_cond $X=0.96 $Y=0.757
+ $X2=2.72 $Y2=0.757
r39 11 32 2.09442 $w=1.398e-06 $l=2.4e-07 $layer=LI1_cond $X=0.96 $Y=0.757
+ $X2=0.72 $Y2=0.757
r40 10 13 50.646 $w=1.675e-06 $l=1.76e-06 $layer=POLY_cond $X=0.96 $Y=2.287
+ $X2=2.72 $Y2=2.287
r41 10 11 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.96
+ $Y=1.515 $X2=0.96 $Y2=1.515
r42 7 49 0.0947698 $w=4.9e-07 $l=3.4e-07 $layer=MET1_cond $X=4.32 $Y=0 $X2=4.66
+ $Y2=0
r43 7 33 1.00344 $w=4.9e-07 $l=3.6e-06 $layer=MET1_cond $X=4.32 $Y=0 $X2=0.72
+ $Y2=0
r44 1 40 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=8.245
+ $Y=0.235 $X2=8.38 $Y2=0.38
r45 1 30 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=8.245
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

