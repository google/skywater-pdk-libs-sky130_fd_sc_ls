# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ls__bufinv_16
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ls__bufinv_16 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  12.00000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.837000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.350000 1.430000 1.780000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  4.390400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 4.660000 1.920000 11.400000 2.150000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 12.000000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 12.000000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 12.000000 0.085000 ;
      RECT  0.000000  3.245000 12.000000 3.415000 ;
      RECT  0.115000  0.350000  0.365000 1.010000 ;
      RECT  0.115000  1.010000  1.770000 1.180000 ;
      RECT  0.120000  1.950000  1.770000 2.120000 ;
      RECT  0.120000  2.120000  0.450000 2.980000 ;
      RECT  0.545000  0.085000  0.875000 0.840000 ;
      RECT  0.650000  2.290000  0.820000 3.245000 ;
      RECT  1.020000  2.120000  1.350000 2.980000 ;
      RECT  1.115000  0.350000  1.285000 1.010000 ;
      RECT  1.465000  0.085000  1.795000 0.840000 ;
      RECT  1.550000  2.290000  1.720000 3.245000 ;
      RECT  1.600000  1.180000  1.770000 1.300000 ;
      RECT  1.600000  1.300000  3.460000 1.630000 ;
      RECT  1.600000  1.630000  1.770000 1.950000 ;
      RECT  1.940000  1.800000  4.070000 1.970000 ;
      RECT  1.940000  1.970000  2.270000 2.980000 ;
      RECT  1.975000  0.350000  2.145000 0.960000 ;
      RECT  1.975000  0.960000  3.935000 1.130000 ;
      RECT  2.325000  0.085000  2.575000 0.790000 ;
      RECT  2.470000  2.140000  2.640000 3.245000 ;
      RECT  2.755000  0.350000  3.005000 0.960000 ;
      RECT  2.840000  1.970000  3.170000 2.980000 ;
      RECT  3.185000  0.085000  3.515000 0.790000 ;
      RECT  3.370000  2.140000  3.540000 3.245000 ;
      RECT  3.685000  0.350000  3.935000 0.960000 ;
      RECT  3.685000  1.130000  3.935000 1.300000 ;
      RECT  3.740000  1.300000  4.435000 1.750000 ;
      RECT  3.740000  1.750000  4.070000 1.800000 ;
      RECT  3.740000  1.970000  4.070000 2.980000 ;
      RECT  4.115000  0.085000  4.445000 1.130000 ;
      RECT  4.270000  1.920000  4.440000 3.245000 ;
      RECT  4.615000  0.350000  4.865000 1.920000 ;
      RECT  4.615000  1.920000  4.970000 2.020000 ;
      RECT  4.640000  2.020000  4.970000 2.980000 ;
      RECT  5.035000  1.300000  5.305000 1.750000 ;
      RECT  5.045000  0.085000  5.295000 1.105000 ;
      RECT  5.170000  1.920000  5.340000 3.245000 ;
      RECT  5.510000  0.350000  5.725000 1.920000 ;
      RECT  5.510000  1.920000  5.870000 2.020000 ;
      RECT  5.540000  2.020000  5.870000 2.980000 ;
      RECT  5.900000  1.300000  6.230000 1.750000 ;
      RECT  5.905000  0.085000  6.235000 1.105000 ;
      RECT  6.070000  1.920000  6.240000 3.245000 ;
      RECT  6.420000  0.350000  6.655000 1.920000 ;
      RECT  6.420000  1.920000  6.770000 2.020000 ;
      RECT  6.440000  2.020000  6.770000 2.980000 ;
      RECT  6.835000  0.085000  7.165000 1.105000 ;
      RECT  6.840000  1.300000  7.170000 1.750000 ;
      RECT  6.970000  1.920000  7.140000 3.245000 ;
      RECT  7.340000  0.350000  7.585000 1.920000 ;
      RECT  7.340000  1.920000  7.670000 2.980000 ;
      RECT  7.760000  1.300000  8.090000 1.750000 ;
      RECT  7.765000  0.085000  8.095000 1.105000 ;
      RECT  7.870000  1.920000  8.040000 3.245000 ;
      RECT  8.240000  2.020000  8.570000 2.980000 ;
      RECT  8.265000  0.350000  8.515000 1.920000 ;
      RECT  8.265000  1.920000  8.570000 2.020000 ;
      RECT  8.685000  1.300000  9.015000 1.750000 ;
      RECT  8.695000  0.085000  9.025000 1.105000 ;
      RECT  8.770000  1.920000  8.995000 3.245000 ;
      RECT  9.190000  2.020000  9.520000 2.980000 ;
      RECT  9.195000  0.350000  9.445000 1.920000 ;
      RECT  9.195000  1.920000  9.520000 2.020000 ;
      RECT  9.615000  1.300000  9.945000 1.750000 ;
      RECT  9.625000  0.085000  9.955000 1.105000 ;
      RECT  9.720000  1.920000  9.955000 3.245000 ;
      RECT 10.125000  0.350000 10.375000 1.920000 ;
      RECT 10.125000  1.920000 10.470000 2.020000 ;
      RECT 10.140000  2.020000 10.470000 2.980000 ;
      RECT 10.545000  1.300000 10.875000 1.750000 ;
      RECT 10.555000  0.085000 10.885000 1.105000 ;
      RECT 10.670000  1.920000 10.885000 3.245000 ;
      RECT 11.055000  0.350000 11.385000 1.790000 ;
      RECT 11.055000  1.790000 11.420000 2.020000 ;
      RECT 11.090000  2.020000 11.420000 2.980000 ;
      RECT 11.555000  0.085000 11.885000 1.130000 ;
      RECT 11.620000  1.820000 11.870000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.225000  1.580000  4.395000 1.750000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.730000  1.950000  4.900000 2.120000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.090000  1.580000  5.260000 1.750000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.620000  1.950000  5.790000 2.120000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  5.980000  1.580000  6.150000 1.750000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.520000  1.950000  6.690000 2.120000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  6.920000  1.580000  7.090000 1.750000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.420000  1.950000  7.590000 2.120000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  1.580000  8.005000 1.750000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.320000  1.950000  8.490000 2.120000 ;
      RECT  8.765000  1.580000  8.935000 1.750000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.270000  1.950000  9.440000 2.120000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.690000  1.580000  9.860000 1.750000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.220000  1.950000 10.390000 2.120000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.625000  1.580000 10.795000 1.750000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.170000  1.950000 11.340000 2.120000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
    LAYER met1 ;
      RECT 4.155000 1.550000 10.855000 1.780000 ;
  END
END sky130_fd_sc_ls__bufinv_16
END LIBRARY
