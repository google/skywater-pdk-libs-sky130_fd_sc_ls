* File: sky130_fd_sc_ls__a221oi_1.pxi.spice
* Created: Fri Aug 28 12:53:17 2020
* 
x_PM_SKY130_FD_SC_LS__A221OI_1%C1 N_C1_c_56_n N_C1_M1006_g N_C1_M1003_g C1
+ N_C1_c_54_n N_C1_c_55_n PM_SKY130_FD_SC_LS__A221OI_1%C1
x_PM_SKY130_FD_SC_LS__A221OI_1%B2 N_B2_c_80_n N_B2_M1009_g N_B2_M1007_g B2 B2
+ PM_SKY130_FD_SC_LS__A221OI_1%B2
x_PM_SKY130_FD_SC_LS__A221OI_1%B1 N_B1_M1002_g N_B1_c_111_n N_B1_M1001_g B1
+ N_B1_c_112_n PM_SKY130_FD_SC_LS__A221OI_1%B1
x_PM_SKY130_FD_SC_LS__A221OI_1%A1 N_A1_c_141_n N_A1_M1008_g N_A1_M1004_g A1
+ N_A1_c_143_n PM_SKY130_FD_SC_LS__A221OI_1%A1
x_PM_SKY130_FD_SC_LS__A221OI_1%A2 N_A2_c_172_n N_A2_M1005_g N_A2_c_173_n
+ N_A2_M1000_g A2 A2 PM_SKY130_FD_SC_LS__A221OI_1%A2
x_PM_SKY130_FD_SC_LS__A221OI_1%Y N_Y_M1003_s N_Y_M1002_d N_Y_M1006_s N_Y_c_194_n
+ N_Y_c_195_n Y Y Y Y Y Y N_Y_c_197_n PM_SKY130_FD_SC_LS__A221OI_1%Y
x_PM_SKY130_FD_SC_LS__A221OI_1%A_118_368# N_A_118_368#_M1006_d
+ N_A_118_368#_M1009_d N_A_118_368#_c_233_n N_A_118_368#_c_234_n
+ N_A_118_368#_c_235_n N_A_118_368#_c_242_n
+ PM_SKY130_FD_SC_LS__A221OI_1%A_118_368#
x_PM_SKY130_FD_SC_LS__A221OI_1%A_263_368# N_A_263_368#_M1009_s
+ N_A_263_368#_M1001_d N_A_263_368#_M1000_d N_A_263_368#_c_261_n
+ N_A_263_368#_c_262_n N_A_263_368#_c_268_n N_A_263_368#_c_263_n
+ N_A_263_368#_c_276_n N_A_263_368#_c_264_n N_A_263_368#_c_265_n
+ N_A_263_368#_c_273_n PM_SKY130_FD_SC_LS__A221OI_1%A_263_368#
x_PM_SKY130_FD_SC_LS__A221OI_1%VPWR N_VPWR_M1008_d N_VPWR_c_302_n N_VPWR_c_303_n
+ N_VPWR_c_304_n VPWR N_VPWR_c_305_n N_VPWR_c_301_n
+ PM_SKY130_FD_SC_LS__A221OI_1%VPWR
x_PM_SKY130_FD_SC_LS__A221OI_1%VGND N_VGND_M1003_d N_VGND_M1005_d N_VGND_c_334_n
+ N_VGND_c_335_n N_VGND_c_336_n N_VGND_c_337_n N_VGND_c_338_n N_VGND_c_339_n
+ VGND N_VGND_c_340_n N_VGND_c_341_n PM_SKY130_FD_SC_LS__A221OI_1%VGND
cc_1 VNB N_C1_M1003_g 0.031956f $X=-0.19 $Y=-0.245 $X2=1.14 $Y2=0.74
cc_2 VNB N_C1_c_54_n 0.0539437f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.515
cc_3 VNB N_C1_c_55_n 0.00305603f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.515
cc_4 VNB N_B2_c_80_n 0.0215337f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.765
cc_5 VNB N_B2_M1007_g 0.0236982f $X=-0.19 $Y=-0.245 $X2=1.14 $Y2=0.74
cc_6 VNB B2 0.00423229f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_B1_M1002_g 0.0264675f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=2.4
cc_8 VNB N_B1_c_111_n 0.0262387f $X=-0.19 $Y=-0.245 $X2=1.14 $Y2=0.74
cc_9 VNB N_B1_c_112_n 0.00166531f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.515
cc_10 VNB N_A1_c_141_n 0.0262687f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.765
cc_11 VNB N_A1_M1004_g 0.0272859f $X=-0.19 $Y=-0.245 $X2=1.14 $Y2=0.74
cc_12 VNB N_A1_c_143_n 0.00487854f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.515
cc_13 VNB N_A2_c_172_n 0.0204958f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.765
cc_14 VNB N_A2_c_173_n 0.0424977f $X=-0.19 $Y=-0.245 $X2=1.14 $Y2=1.35
cc_15 VNB A2 0.0422683f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_16 VNB N_Y_c_194_n 0.0208183f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.557
cc_17 VNB N_Y_c_195_n 0.00420435f $X=-0.19 $Y=-0.245 $X2=1.14 $Y2=1.557
cc_18 VNB Y 0.0267465f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_Y_c_197_n 0.0616195f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_VPWR_c_301_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_334_n 0.00685096f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_335_n 0.0351314f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.515
cc_23 VNB N_VGND_c_336_n 0.0347153f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_337_n 0.0069273f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.665
cc_25 VNB N_VGND_c_338_n 0.0453999f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_339_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_340_n 0.0129628f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_341_n 0.255119f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VPB N_C1_c_56_n 0.0225683f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=1.765
cc_30 VPB N_C1_c_54_n 0.0305215f $X=-0.19 $Y=1.66 $X2=0.71 $Y2=1.515
cc_31 VPB N_C1_c_55_n 0.00363032f $X=-0.19 $Y=1.66 $X2=0.71 $Y2=1.515
cc_32 VPB N_B2_c_80_n 0.0304193f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=1.765
cc_33 VPB B2 0.0124171f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_34 VPB N_B1_c_111_n 0.0261546f $X=-0.19 $Y=1.66 $X2=1.14 $Y2=0.74
cc_35 VPB N_B1_c_112_n 0.00293322f $X=-0.19 $Y=1.66 $X2=0.71 $Y2=1.515
cc_36 VPB N_A1_c_141_n 0.0281677f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=1.765
cc_37 VPB N_A1_c_143_n 0.00283747f $X=-0.19 $Y=1.66 $X2=0.71 $Y2=1.515
cc_38 VPB N_A2_c_173_n 0.0316663f $X=-0.19 $Y=1.66 $X2=1.14 $Y2=1.35
cc_39 VPB Y 0.054467f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_40 VPB N_A_118_368#_c_233_n 0.0127217f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_41 VPB N_A_118_368#_c_234_n 0.0230644f $X=-0.19 $Y=1.66 $X2=0.71 $Y2=1.515
cc_42 VPB N_A_118_368#_c_235_n 0.00294869f $X=-0.19 $Y=1.66 $X2=1.14 $Y2=1.557
cc_43 VPB N_A_263_368#_c_261_n 0.00242573f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=1.557
cc_44 VPB N_A_263_368#_c_262_n 0.00759638f $X=-0.19 $Y=1.66 $X2=0.71 $Y2=1.515
cc_45 VPB N_A_263_368#_c_263_n 0.00254209f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_A_263_368#_c_264_n 0.0151999f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB N_A_263_368#_c_265_n 0.0360166f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_302_n 0.00993371f $X=-0.19 $Y=1.66 $X2=1.14 $Y2=0.74
cc_49 VPB N_VPWR_c_303_n 0.0690385f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_304_n 0.00670627f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=1.557
cc_51 VPB N_VPWR_c_305_n 0.0255159f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_301_n 0.0783071f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 N_C1_c_54_n N_B2_c_80_n 0.0205274f $X=0.71 $Y=1.515 $X2=-0.19 $Y2=-0.245
cc_54 N_C1_M1003_g N_B2_M1007_g 0.026363f $X=1.14 $Y=0.74 $X2=0 $Y2=0
cc_55 N_C1_c_54_n B2 0.0162492f $X=0.71 $Y=1.515 $X2=0 $Y2=0
cc_56 N_C1_c_55_n B2 0.0298996f $X=0.71 $Y=1.515 $X2=0 $Y2=0
cc_57 N_C1_M1003_g N_Y_c_194_n 0.0116701f $X=1.14 $Y=0.74 $X2=0 $Y2=0
cc_58 N_C1_c_56_n Y 0.00993465f $X=0.515 $Y=1.765 $X2=0 $Y2=0
cc_59 N_C1_M1003_g Y 0.00356034f $X=1.14 $Y=0.74 $X2=0 $Y2=0
cc_60 N_C1_c_54_n Y 0.012015f $X=0.71 $Y=1.515 $X2=0 $Y2=0
cc_61 N_C1_c_55_n Y 0.033251f $X=0.71 $Y=1.515 $X2=0 $Y2=0
cc_62 N_C1_M1003_g N_Y_c_197_n 0.0140845f $X=1.14 $Y=0.74 $X2=0 $Y2=0
cc_63 N_C1_c_54_n N_Y_c_197_n 0.0168196f $X=0.71 $Y=1.515 $X2=0 $Y2=0
cc_64 N_C1_c_55_n N_Y_c_197_n 0.0281815f $X=0.71 $Y=1.515 $X2=0 $Y2=0
cc_65 N_C1_c_56_n N_A_118_368#_c_233_n 0.0104363f $X=0.515 $Y=1.765 $X2=0 $Y2=0
cc_66 N_C1_c_54_n N_A_118_368#_c_233_n 0.00267593f $X=0.71 $Y=1.515 $X2=0 $Y2=0
cc_67 N_C1_c_55_n N_A_118_368#_c_233_n 0.023771f $X=0.71 $Y=1.515 $X2=0 $Y2=0
cc_68 N_C1_c_56_n N_A_118_368#_c_235_n 0.00803572f $X=0.515 $Y=1.765 $X2=0 $Y2=0
cc_69 N_C1_c_56_n N_VPWR_c_303_n 0.0044313f $X=0.515 $Y=1.765 $X2=0 $Y2=0
cc_70 N_C1_c_56_n N_VPWR_c_301_n 0.00862451f $X=0.515 $Y=1.765 $X2=0 $Y2=0
cc_71 N_C1_M1003_g N_VGND_c_334_n 0.00601099f $X=1.14 $Y=0.74 $X2=0 $Y2=0
cc_72 N_C1_M1003_g N_VGND_c_336_n 0.00433162f $X=1.14 $Y=0.74 $X2=0 $Y2=0
cc_73 N_C1_M1003_g N_VGND_c_341_n 0.00822437f $X=1.14 $Y=0.74 $X2=0 $Y2=0
cc_74 N_B2_M1007_g N_B1_M1002_g 0.0441025f $X=1.68 $Y=0.74 $X2=0 $Y2=0
cc_75 N_B2_c_80_n N_B1_c_111_n 0.0744247f $X=1.665 $Y=1.765 $X2=0 $Y2=0
cc_76 B2 N_B1_c_111_n 0.00235456f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_77 N_B2_c_80_n N_B1_c_112_n 6.89489e-19 $X=1.665 $Y=1.765 $X2=0 $Y2=0
cc_78 B2 N_B1_c_112_n 0.0366307f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_79 N_B2_c_80_n N_Y_c_194_n 0.00411108f $X=1.665 $Y=1.765 $X2=0 $Y2=0
cc_80 N_B2_M1007_g N_Y_c_194_n 0.0143728f $X=1.68 $Y=0.74 $X2=0 $Y2=0
cc_81 N_B2_M1007_g N_Y_c_197_n 9.00978e-19 $X=1.68 $Y=0.74 $X2=0 $Y2=0
cc_82 B2 N_Y_c_197_n 0.0544896f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_83 N_B2_c_80_n N_A_118_368#_c_233_n 0.00469763f $X=1.665 $Y=1.765 $X2=0 $Y2=0
cc_84 N_B2_c_80_n N_A_118_368#_c_234_n 0.0144793f $X=1.665 $Y=1.765 $X2=0 $Y2=0
cc_85 N_B2_c_80_n N_A_118_368#_c_242_n 0.0124846f $X=1.665 $Y=1.765 $X2=0 $Y2=0
cc_86 N_B2_c_80_n N_A_263_368#_c_261_n 7.09603e-19 $X=1.665 $Y=1.765 $X2=0 $Y2=0
cc_87 B2 N_A_263_368#_c_261_n 0.0233995f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_88 N_B2_c_80_n N_A_263_368#_c_268_n 0.0126342f $X=1.665 $Y=1.765 $X2=0 $Y2=0
cc_89 B2 N_A_263_368#_c_268_n 0.0152441f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_90 N_B2_c_80_n N_VPWR_c_303_n 0.00278257f $X=1.665 $Y=1.765 $X2=0 $Y2=0
cc_91 N_B2_c_80_n N_VPWR_c_301_n 0.00358707f $X=1.665 $Y=1.765 $X2=0 $Y2=0
cc_92 N_B2_M1007_g N_VGND_c_334_n 0.0141323f $X=1.68 $Y=0.74 $X2=0 $Y2=0
cc_93 N_B2_M1007_g N_VGND_c_338_n 0.00383152f $X=1.68 $Y=0.74 $X2=0 $Y2=0
cc_94 N_B2_M1007_g N_VGND_c_341_n 0.0075694f $X=1.68 $Y=0.74 $X2=0 $Y2=0
cc_95 N_B1_c_111_n N_A1_c_141_n 0.0312135f $X=2.115 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_96 N_B1_c_112_n N_A1_c_141_n 0.00173907f $X=2.13 $Y=1.515 $X2=-0.19
+ $Y2=-0.245
cc_97 N_B1_M1002_g N_A1_M1004_g 0.0173199f $X=2.04 $Y=0.74 $X2=0 $Y2=0
cc_98 N_B1_c_111_n N_A1_c_143_n 0.00128912f $X=2.115 $Y=1.765 $X2=0 $Y2=0
cc_99 N_B1_c_112_n N_A1_c_143_n 0.0277336f $X=2.13 $Y=1.515 $X2=0 $Y2=0
cc_100 N_B1_M1002_g N_Y_c_194_n 0.0154892f $X=2.04 $Y=0.74 $X2=0 $Y2=0
cc_101 N_B1_c_111_n N_Y_c_194_n 0.00136813f $X=2.115 $Y=1.765 $X2=0 $Y2=0
cc_102 N_B1_c_112_n N_Y_c_194_n 0.0259226f $X=2.13 $Y=1.515 $X2=0 $Y2=0
cc_103 N_B1_M1002_g N_Y_c_195_n 0.00528753f $X=2.04 $Y=0.74 $X2=0 $Y2=0
cc_104 N_B1_c_111_n N_A_118_368#_c_234_n 0.00401993f $X=2.115 $Y=1.765 $X2=0
+ $Y2=0
cc_105 N_B1_c_111_n N_A_118_368#_c_242_n 0.00701365f $X=2.115 $Y=1.765 $X2=0
+ $Y2=0
cc_106 N_B1_c_111_n N_A_263_368#_c_268_n 0.0130645f $X=2.115 $Y=1.765 $X2=0
+ $Y2=0
cc_107 N_B1_c_112_n N_A_263_368#_c_268_n 0.0178949f $X=2.13 $Y=1.515 $X2=0 $Y2=0
cc_108 N_B1_c_111_n N_A_263_368#_c_263_n 0.00613504f $X=2.115 $Y=1.765 $X2=0
+ $Y2=0
cc_109 N_B1_c_111_n N_A_263_368#_c_273_n 2.39865e-19 $X=2.115 $Y=1.765 $X2=0
+ $Y2=0
cc_110 N_B1_c_112_n N_A_263_368#_c_273_n 0.00346357f $X=2.13 $Y=1.515 $X2=0
+ $Y2=0
cc_111 N_B1_c_111_n N_VPWR_c_303_n 0.0044313f $X=2.115 $Y=1.765 $X2=0 $Y2=0
cc_112 N_B1_c_111_n N_VPWR_c_301_n 0.00854553f $X=2.115 $Y=1.765 $X2=0 $Y2=0
cc_113 N_B1_M1002_g N_VGND_c_334_n 0.00191029f $X=2.04 $Y=0.74 $X2=0 $Y2=0
cc_114 N_B1_M1002_g N_VGND_c_338_n 0.00461464f $X=2.04 $Y=0.74 $X2=0 $Y2=0
cc_115 N_B1_M1002_g N_VGND_c_341_n 0.00910921f $X=2.04 $Y=0.74 $X2=0 $Y2=0
cc_116 N_A1_M1004_g N_A2_c_172_n 0.0432957f $X=2.76 $Y=0.74 $X2=-0.19 $Y2=-0.245
cc_117 N_A1_c_141_n N_A2_c_173_n 0.0707565f $X=2.595 $Y=1.765 $X2=0 $Y2=0
cc_118 N_A1_c_143_n N_A2_c_173_n 0.00344439f $X=2.67 $Y=1.515 $X2=0 $Y2=0
cc_119 N_A1_M1004_g A2 0.00572702f $X=2.76 $Y=0.74 $X2=0 $Y2=0
cc_120 N_A1_c_143_n A2 0.0168427f $X=2.67 $Y=1.515 $X2=0 $Y2=0
cc_121 N_A1_c_141_n N_Y_c_194_n 5.40529e-19 $X=2.595 $Y=1.765 $X2=0 $Y2=0
cc_122 N_A1_M1004_g N_Y_c_194_n 0.00555347f $X=2.76 $Y=0.74 $X2=0 $Y2=0
cc_123 N_A1_c_143_n N_Y_c_194_n 0.00595492f $X=2.67 $Y=1.515 $X2=0 $Y2=0
cc_124 N_A1_M1004_g N_Y_c_195_n 0.0103902f $X=2.76 $Y=0.74 $X2=0 $Y2=0
cc_125 N_A1_c_141_n N_A_118_368#_c_234_n 3.07234e-19 $X=2.595 $Y=1.765 $X2=0
+ $Y2=0
cc_126 N_A1_c_141_n N_A_263_368#_c_263_n 2.47509e-19 $X=2.595 $Y=1.765 $X2=0
+ $Y2=0
cc_127 N_A1_c_141_n N_A_263_368#_c_276_n 0.0142324f $X=2.595 $Y=1.765 $X2=0
+ $Y2=0
cc_128 N_A1_c_143_n N_A_263_368#_c_276_n 0.0226207f $X=2.67 $Y=1.515 $X2=0 $Y2=0
cc_129 N_A1_c_141_n N_A_263_368#_c_264_n 5.93323e-19 $X=2.595 $Y=1.765 $X2=0
+ $Y2=0
cc_130 N_A1_c_141_n N_A_263_368#_c_265_n 7.14599e-19 $X=2.595 $Y=1.765 $X2=0
+ $Y2=0
cc_131 N_A1_c_141_n N_VPWR_c_302_n 0.00252449f $X=2.595 $Y=1.765 $X2=0 $Y2=0
cc_132 N_A1_c_141_n N_VPWR_c_303_n 0.00461464f $X=2.595 $Y=1.765 $X2=0 $Y2=0
cc_133 N_A1_c_141_n N_VPWR_c_301_n 0.00908785f $X=2.595 $Y=1.765 $X2=0 $Y2=0
cc_134 N_A1_M1004_g N_VGND_c_335_n 0.00249753f $X=2.76 $Y=0.74 $X2=0 $Y2=0
cc_135 N_A1_M1004_g N_VGND_c_338_n 0.00461464f $X=2.76 $Y=0.74 $X2=0 $Y2=0
cc_136 N_A1_M1004_g N_VGND_c_341_n 0.00910921f $X=2.76 $Y=0.74 $X2=0 $Y2=0
cc_137 N_A2_c_173_n N_A_263_368#_c_276_n 0.0135061f $X=3.135 $Y=1.765 $X2=0
+ $Y2=0
cc_138 A2 N_A_263_368#_c_276_n 0.00609203f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_139 N_A2_c_173_n N_A_263_368#_c_264_n 0.0071736f $X=3.135 $Y=1.765 $X2=0
+ $Y2=0
cc_140 A2 N_A_263_368#_c_264_n 0.0204504f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_141 N_A2_c_173_n N_A_263_368#_c_265_n 0.0114033f $X=3.135 $Y=1.765 $X2=0
+ $Y2=0
cc_142 N_A2_c_173_n N_VPWR_c_302_n 0.00731029f $X=3.135 $Y=1.765 $X2=0 $Y2=0
cc_143 N_A2_c_173_n N_VPWR_c_305_n 0.00445602f $X=3.135 $Y=1.765 $X2=0 $Y2=0
cc_144 N_A2_c_173_n N_VPWR_c_301_n 0.00861742f $X=3.135 $Y=1.765 $X2=0 $Y2=0
cc_145 N_A2_c_172_n N_VGND_c_335_n 0.017286f $X=3.12 $Y=1.22 $X2=0 $Y2=0
cc_146 N_A2_c_173_n N_VGND_c_335_n 0.00111834f $X=3.135 $Y=1.765 $X2=0 $Y2=0
cc_147 A2 N_VGND_c_335_n 0.0259761f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_148 N_A2_c_172_n N_VGND_c_338_n 0.00383152f $X=3.12 $Y=1.22 $X2=0 $Y2=0
cc_149 N_A2_c_172_n N_VGND_c_341_n 0.0075694f $X=3.12 $Y=1.22 $X2=0 $Y2=0
cc_150 Y N_A_118_368#_c_233_n 0.0640009f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_151 Y N_A_118_368#_c_235_n 0.00536881f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_152 Y N_VPWR_c_303_n 0.011066f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_153 Y N_VPWR_c_301_n 0.00915947f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_154 N_Y_c_194_n N_VGND_M1003_d 0.00320495f $X=2.16 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_155 N_Y_c_194_n N_VGND_c_334_n 0.0227484f $X=2.16 $Y=1.095 $X2=0 $Y2=0
cc_156 N_Y_c_195_n N_VGND_c_334_n 0.00751247f $X=2.375 $Y=0.495 $X2=0 $Y2=0
cc_157 N_Y_c_197_n N_VGND_c_334_n 0.020732f $X=1.09 $Y=0.765 $X2=0 $Y2=0
cc_158 N_Y_c_195_n N_VGND_c_335_n 0.0194588f $X=2.375 $Y=0.495 $X2=0 $Y2=0
cc_159 N_Y_c_197_n N_VGND_c_336_n 0.0428125f $X=1.09 $Y=0.765 $X2=0 $Y2=0
cc_160 N_Y_c_195_n N_VGND_c_338_n 0.0184284f $X=2.375 $Y=0.495 $X2=0 $Y2=0
cc_161 N_Y_c_195_n N_VGND_c_341_n 0.0152535f $X=2.375 $Y=0.495 $X2=0 $Y2=0
cc_162 N_Y_c_197_n N_VGND_c_341_n 0.0354986f $X=1.09 $Y=0.765 $X2=0 $Y2=0
cc_163 N_Y_c_194_n A_351_74# 0.00366293f $X=2.16 $Y=1.095 $X2=-0.19 $Y2=-0.245
cc_164 N_A_118_368#_c_234_n N_A_263_368#_M1009_s 0.00260133f $X=1.725 $Y=2.99
+ $X2=-0.19 $Y2=1.66
cc_165 N_A_118_368#_c_233_n N_A_263_368#_c_261_n 0.00876529f $X=0.74 $Y=2.115
+ $X2=0 $Y2=0
cc_166 N_A_118_368#_c_233_n N_A_263_368#_c_262_n 0.0294466f $X=0.74 $Y=2.115
+ $X2=0 $Y2=0
cc_167 N_A_118_368#_c_234_n N_A_263_368#_c_262_n 0.0196739f $X=1.725 $Y=2.99
+ $X2=0 $Y2=0
cc_168 N_A_118_368#_M1009_d N_A_263_368#_c_268_n 0.00857291f $X=1.74 $Y=1.84
+ $X2=0 $Y2=0
cc_169 N_A_118_368#_c_242_n N_A_263_368#_c_268_n 0.0171814f $X=1.89 $Y=2.4 $X2=0
+ $Y2=0
cc_170 N_A_118_368#_c_234_n N_A_263_368#_c_263_n 0.00536881f $X=1.725 $Y=2.99
+ $X2=0 $Y2=0
cc_171 N_A_118_368#_c_242_n N_A_263_368#_c_263_n 0.0412035f $X=1.89 $Y=2.4 $X2=0
+ $Y2=0
cc_172 N_A_118_368#_c_234_n N_VPWR_c_302_n 0.00295634f $X=1.725 $Y=2.99 $X2=0
+ $Y2=0
cc_173 N_A_118_368#_c_234_n N_VPWR_c_303_n 0.0759258f $X=1.725 $Y=2.99 $X2=0
+ $Y2=0
cc_174 N_A_118_368#_c_235_n N_VPWR_c_303_n 0.0236039f $X=0.905 $Y=2.99 $X2=0
+ $Y2=0
cc_175 N_A_118_368#_c_234_n N_VPWR_c_301_n 0.0429008f $X=1.725 $Y=2.99 $X2=0
+ $Y2=0
cc_176 N_A_118_368#_c_235_n N_VPWR_c_301_n 0.012761f $X=0.905 $Y=2.99 $X2=0
+ $Y2=0
cc_177 N_A_263_368#_c_276_n N_VPWR_M1008_d 0.010589f $X=3.195 $Y=2.035 $X2=-0.19
+ $Y2=1.66
cc_178 N_A_263_368#_c_263_n N_VPWR_c_302_n 0.00155548f $X=2.34 $Y=2.44 $X2=0
+ $Y2=0
cc_179 N_A_263_368#_c_276_n N_VPWR_c_302_n 0.022455f $X=3.195 $Y=2.035 $X2=0
+ $Y2=0
cc_180 N_A_263_368#_c_265_n N_VPWR_c_302_n 0.026688f $X=3.36 $Y=2.815 $X2=0
+ $Y2=0
cc_181 N_A_263_368#_c_263_n N_VPWR_c_303_n 0.011066f $X=2.34 $Y=2.44 $X2=0 $Y2=0
cc_182 N_A_263_368#_c_265_n N_VPWR_c_305_n 0.0145938f $X=3.36 $Y=2.815 $X2=0
+ $Y2=0
cc_183 N_A_263_368#_c_263_n N_VPWR_c_301_n 0.00915947f $X=2.34 $Y=2.44 $X2=0
+ $Y2=0
cc_184 N_A_263_368#_c_265_n N_VPWR_c_301_n 0.0120466f $X=3.36 $Y=2.815 $X2=0
+ $Y2=0
