* File: sky130_fd_sc_ls__or4b_1.spice
* Created: Fri Aug 28 14:00:11 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__or4b_1.pex.spice"
.subckt sky130_fd_sc_ls__or4b_1  VNB VPB D_N C B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* C	C
* D_N	D_N
* VPB	VPB
* VNB	VNB
MM1008 N_VGND_M1008_d N_D_N_M1008_g N_A_27_74#_M1008_s VNB NSHORT L=0.15 W=0.55
+ AD=0.1155 AS=0.15675 PD=0.97 PS=1.67 NRD=15.264 NRS=0 M=1 R=3.66667 SA=75000.2
+ SB=75003.5 A=0.0825 P=1.4 MULT=1
MM1010 N_A_228_74#_M1010_d N_A_27_74#_M1010_g N_VGND_M1008_d VNB NSHORT L=0.15
+ W=0.55 AD=0.254375 AS=0.1155 PD=1.475 PS=0.97 NRD=0 NRS=15.264 M=1 R=3.66667
+ SA=75000.8 SB=75002.9 A=0.0825 P=1.4 MULT=1
MM1000 N_VGND_M1000_d N_C_M1000_g N_A_228_74#_M1010_d VNB NSHORT L=0.15 W=0.55
+ AD=0.1155 AS=0.254375 PD=0.97 PS=1.475 NRD=15.264 NRS=0 M=1 R=3.66667
+ SA=75001.9 SB=75001.9 A=0.0825 P=1.4 MULT=1
MM1007 N_A_228_74#_M1007_d N_B_M1007_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.55
+ AD=0.077 AS=0.1155 PD=0.83 PS=0.97 NRD=0 NRS=15.264 M=1 R=3.66667 SA=75002.4
+ SB=75001.3 A=0.0825 P=1.4 MULT=1
MM1011 N_VGND_M1011_d N_A_M1011_g N_A_228_74#_M1007_d VNB NSHORT L=0.15 W=0.55
+ AD=0.136328 AS=0.077 PD=1.0531 PS=0.83 NRD=22.908 NRS=0 M=1 R=3.66667
+ SA=75002.9 SB=75000.9 A=0.0825 P=1.4 MULT=1
MM1004 N_X_M1004_d N_A_228_74#_M1004_g N_VGND_M1011_d VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.183422 PD=2.05 PS=1.4169 NRD=0 NRS=17.832 M=1 R=4.93333
+ SA=75002.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1006 N_VPWR_M1006_d N_D_N_M1006_g N_A_27_74#_M1006_s VPB PHIGHVT L=0.15 W=0.84
+ AD=0.2898 AS=0.2478 PD=2.37 PS=2.27 NRD=14.0658 NRS=2.3443 M=1 R=5.6
+ SA=75000.2 SB=75000.3 A=0.126 P=1.98 MULT=1
MM1001 A_356_368# N_A_27_74#_M1001_g N_A_228_74#_M1001_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.295 PD=1.27 PS=2.59 NRD=15.7403 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75002.3 A=0.15 P=2.3 MULT=1
MM1009 A_440_368# N_C_M1009_g A_356_368# VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=15.7403 NRS=15.7403 M=1 R=6.66667 SA=75000.6
+ SB=75001.9 A=0.15 P=2.3 MULT=1
MM1003 A_524_368# N_B_M1003_g A_440_368# VPB PHIGHVT L=0.15 W=1 AD=0.195
+ AS=0.135 PD=1.39 PS=1.27 NRD=27.5603 NRS=15.7403 M=1 R=6.66667 SA=75001.1
+ SB=75001.4 A=0.15 P=2.3 MULT=1
MM1002 N_VPWR_M1002_d N_A_M1002_g A_524_368# VPB PHIGHVT L=0.15 W=1 AD=0.274245
+ AS=0.195 PD=1.56604 PS=1.39 NRD=39.8728 NRS=27.5603 M=1 R=6.66667 SA=75001.6
+ SB=75000.9 A=0.15 P=2.3 MULT=1
MM1005 N_X_M1005_d N_A_228_74#_M1005_g N_VPWR_M1002_d VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.307155 PD=2.83 PS=1.75396 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75002.1 SB=75000.2 A=0.168 P=2.54 MULT=1
DX12_noxref VNB VPB NWDIODE A=8.742 P=13.12
*
.include "sky130_fd_sc_ls__or4b_1.pxi.spice"
*
.ends
*
*
