* NGSPICE file created from sky130_fd_sc_ls__fill_diode_4.ext - technology: sky130A

.subckt sky130_fd_sc_ls__fill_diode_4 VGND VNB VPB VPWR
.ends

