# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_ls__and4bb_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_ls__and4bb_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.280000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A_N
    ANTENNAGATEAREA  0.208500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.450000 0.550000 1.780000 ;
    END
  END A_N
  PIN B_N
    ANTENNAGATEAREA  0.208500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.825000 1.180000 5.155000 1.590000 ;
    END
  END B_N
  PIN C
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.310000 1.420000 2.755000 1.780000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.925000 1.420000 3.255000 1.780000 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.815000 0.920000 4.195000 1.170000 ;
        RECT 3.835000 1.840000 4.195000 2.980000 ;
        RECT 4.025000 1.170000 4.195000 1.840000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.280000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000000 0.000000 5.280000 0.245000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.660000 5.470000 3.520000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.280000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.280000 0.085000 ;
      RECT 0.000000  3.245000 5.280000 3.415000 ;
      RECT 0.115000  0.350000 0.365000 1.110000 ;
      RECT 0.115000  1.110000 0.935000 1.280000 ;
      RECT 0.210000  1.950000 0.935000 2.120000 ;
      RECT 0.210000  2.120000 0.540000 2.820000 ;
      RECT 0.545000  0.085000 0.875000 0.940000 ;
      RECT 0.765000  1.280000 0.935000 1.340000 ;
      RECT 0.765000  1.340000 1.260000 1.670000 ;
      RECT 0.765000  1.670000 0.935000 1.950000 ;
      RECT 0.780000  2.290000 1.110000 3.245000 ;
      RECT 1.105000  0.390000 1.600000 1.170000 ;
      RECT 1.430000  1.170000 1.600000 1.940000 ;
      RECT 1.430000  1.940000 1.760000 1.950000 ;
      RECT 1.430000  1.950000 3.665000 2.120000 ;
      RECT 1.430000  2.120000 1.760000 2.980000 ;
      RECT 1.770000  1.000000 3.645000 1.170000 ;
      RECT 1.770000  1.170000 2.100000 1.590000 ;
      RECT 2.065000  2.290000 2.395000 3.245000 ;
      RECT 2.610000  2.120000 2.940000 2.980000 ;
      RECT 2.975000  0.085000 3.305000 0.830000 ;
      RECT 3.200000  2.290000 3.530000 3.245000 ;
      RECT 3.475000  0.580000 5.165000 0.750000 ;
      RECT 3.475000  0.750000 3.645000 1.000000 ;
      RECT 3.495000  1.340000 3.855000 1.670000 ;
      RECT 3.495000  1.670000 3.665000 1.950000 ;
      RECT 4.325000  0.085000 4.655000 0.410000 ;
      RECT 4.365000  0.750000 4.535000 1.760000 ;
      RECT 4.365000  1.760000 5.165000 1.930000 ;
      RECT 4.365000  2.100000 4.615000 3.245000 ;
      RECT 4.820000  1.930000 5.165000 2.700000 ;
      RECT 4.835000  0.750000 5.165000 1.010000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
  END
END sky130_fd_sc_ls__and4bb_2
END LIBRARY
