* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__sdfbbn_2 CLK_N D RESET_B SCD SCE SET_B VGND VNB VPB VPWR
+ Q Q_N
M1000 a_197_119# D a_206_464# VPB phighvt w=640000u l=150000u
+  ad=4.128e+11p pd=3.85e+06u as=1.536e+11p ps=1.76e+06u
M1001 VPWR a_3272_94# Q VPB phighvt w=1.12e+06u l=150000u
+  ad=4.12873e+12p pd=3.022e+07u as=3.36e+11p ps=2.84e+06u
M1002 a_2452_74# SET_B VGND VNB nshort w=740000u l=150000u
+  ad=5.7435e+11p pd=4.64e+06u as=2.86405e+12p ps=2.37e+07u
M1003 VGND a_2216_410# Q_N VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.072e+11p ps=2.04e+06u
M1004 a_119_119# SCD VGND VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1005 VGND RESET_B a_1643_257# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.176e+11p ps=1.4e+06u
M1006 a_197_119# a_868_368# a_1154_464# VNB nshort w=420000u l=150000u
+  ad=4.347e+11p pd=3.75e+06u as=1.281e+11p ps=1.45e+06u
M1007 a_2452_74# a_1997_82# a_2216_410# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.072e+11p ps=2.04e+06u
M1008 VPWR a_2216_410# a_2171_508# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1009 a_1986_424# a_1007_366# VPWR VPB phighvt w=840000u l=150000u
+  ad=2.016e+11p pd=2.16e+06u as=0p ps=0u
M1010 a_1997_82# a_868_368# a_1986_424# VPB phighvt w=840000u l=150000u
+  ad=2.856e+11p pd=2.45e+06u as=0p ps=0u
M1011 VPWR SET_B a_2216_410# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=5.9e+11p ps=5.18e+06u
M1012 a_2247_82# a_868_368# a_1997_82# VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=4.945e+11p ps=3.3e+06u
M1013 a_197_119# a_688_98# a_1154_464# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=2.266e+11p ps=2.05e+06u
M1014 a_2556_392# a_1643_257# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1015 a_27_464# a_341_410# a_197_119# VPB phighvt w=640000u l=150000u
+  ad=3.776e+11p pd=3.74e+06u as=0p ps=0u
M1016 a_1154_464# a_688_98# a_1185_125# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1017 a_1007_366# a_1154_464# a_1473_73# VNB nshort w=550000u l=150000u
+  ad=1.54e+11p pd=1.66e+06u as=6.0335e+11p ps=4.55e+06u
M1018 a_1473_73# a_1643_257# a_1007_366# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND a_2216_410# a_3272_94# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1020 a_1997_82# a_688_98# a_1902_125# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=2.16375e+11p ps=2.18e+06u
M1021 Q_N a_2216_410# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 Q a_3272_94# VGND VNB nshort w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1023 Q_N a_2216_410# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=0p ps=0u
M1024 a_341_410# SCE VPWR VPB phighvt w=640000u l=150000u
+  ad=1.888e+11p pd=1.87e+06u as=0p ps=0u
M1025 VGND a_341_410# a_363_119# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1026 VPWR RESET_B a_1643_257# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.888e+11p ps=1.87e+06u
M1027 a_1185_125# a_1007_366# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VPWR SCD a_27_464# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_206_464# SCE VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VPWR a_1643_257# a_1592_424# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=2.268e+11p ps=2.22e+06u
M1031 a_2171_508# a_688_98# a_1997_82# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_197_119# SCE a_119_119# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VPWR a_2216_410# Q_N VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_1592_424# a_1154_464# a_1007_366# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=9.954e+11p ps=5.73e+06u
M1035 VGND CLK_N a_688_98# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1036 VPWR CLK_N a_688_98# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.304e+11p ps=2.83e+06u
M1037 a_341_410# SCE VGND VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1038 a_2216_410# a_1643_257# a_2452_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_1154_464# a_868_368# a_1070_464# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1040 Q a_3272_94# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1041 VGND a_3272_94# Q VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1042 a_363_119# D a_197_119# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1043 a_868_368# a_688_98# VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1044 VGND a_2216_410# a_2247_82# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1045 a_1070_464# a_1007_366# VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1046 a_1902_125# a_1007_366# VGND VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1047 VGND SET_B a_1473_73# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1048 a_868_368# a_688_98# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=0p ps=0u
M1049 a_1007_366# SET_B VPWR VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1050 VPWR a_2216_410# a_3272_94# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1051 a_2216_410# a_1997_82# a_2556_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
