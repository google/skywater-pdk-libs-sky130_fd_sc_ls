* File: sky130_fd_sc_ls__sdfbbn_2.pex.spice
* Created: Fri Aug 28 14:01:53 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__SDFBBN_2%SCD 2 3 5 8 9 10 14 15 16
r29 18 19 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.97 $X2=0.385 $Y2=1.97
r30 14 16 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.407 $Y=1.29
+ $X2=0.407 $Y2=1.125
r31 14 15 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.29 $X2=0.385 $Y2=1.29
r32 10 19 8.27047 $w=4.23e-07 $l=3.05e-07 $layer=LI1_cond $X=0.337 $Y=1.665
+ $X2=0.337 $Y2=1.97
r33 9 10 10.033 $w=4.23e-07 $l=3.7e-07 $layer=LI1_cond $X=0.337 $Y=1.295
+ $X2=0.337 $Y2=1.665
r34 9 15 0.135582 $w=4.23e-07 $l=5e-09 $layer=LI1_cond $X=0.337 $Y=1.295
+ $X2=0.337 $Y2=1.29
r35 8 16 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.52 $Y=0.805
+ $X2=0.52 $Y2=1.125
r36 3 18 56.1009 $w=3.02e-07 $l=3.20273e-07 $layer=POLY_cond $X=0.505 $Y=2.245
+ $X2=0.407 $Y2=1.97
r37 3 5 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.505 $Y=2.245
+ $X2=0.505 $Y2=2.64
r38 2 18 4.79453 $w=3.75e-07 $l=2.2e-08 $layer=POLY_cond $X=0.407 $Y=1.948
+ $X2=0.407 $Y2=1.97
r39 1 14 3.26277 $w=3.75e-07 $l=2.2e-08 $layer=POLY_cond $X=0.407 $Y=1.312
+ $X2=0.407 $Y2=1.29
r40 1 2 94.3237 $w=3.75e-07 $l=6.36e-07 $layer=POLY_cond $X=0.407 $Y=1.312
+ $X2=0.407 $Y2=1.948
.ends

.subckt PM_SKY130_FD_SC_LS__SDFBBN_2%D 1 3 5 8 10 12 19
c59 12 0 1.16605e-19 $X=1.68 $Y=1.665
r60 17 19 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.65 $Y=1.625 $X2=1.74
+ $Y2=1.625
r61 14 17 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=1.42 $Y=1.625
+ $X2=1.65 $Y2=1.625
r62 12 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.65
+ $Y=1.625 $X2=1.65 $Y2=1.625
r63 10 11 18.5385 $w=1.95e-07 $l=7.5e-08 $layer=POLY_cond $X=1.345 $Y=2.14
+ $X2=1.42 $Y2=2.14
r64 6 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.74 $Y=1.46
+ $X2=1.74 $Y2=1.625
r65 6 8 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=1.74 $Y=1.46 $X2=1.74
+ $Y2=0.805
r66 5 11 8.99251 $w=1.5e-07 $l=1.05e-07 $layer=POLY_cond $X=1.42 $Y=2.035
+ $X2=1.42 $Y2=2.14
r67 4 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.42 $Y=1.79
+ $X2=1.42 $Y2=1.625
r68 4 5 125.628 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=1.42 $Y=1.79 $X2=1.42
+ $Y2=2.035
r69 1 10 8.99251 $w=1.5e-07 $l=1.05e-07 $layer=POLY_cond $X=1.345 $Y=2.245
+ $X2=1.345 $Y2=2.14
r70 1 3 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.345 $Y=2.245
+ $X2=1.345 $Y2=2.64
.ends

.subckt PM_SKY130_FD_SC_LS__SDFBBN_2%A_341_410# 1 2 7 9 10 11 14 17 18 20 21 24
+ 28 32 34
c82 34 0 2.50597e-19 $X=3.067 $Y=1.645
c83 28 0 1.21362e-19 $X=3.025 $Y=0.815
c84 24 0 3.52871e-20 $X=2.77 $Y=1.645
c85 21 0 3.06618e-19 $X=2.94 $Y=1.645
c86 11 0 1.16605e-19 $X=1.885 $Y=2.125
r87 30 34 6.41553 $w=2.52e-07 $l=1.66493e-07 $layer=LI1_cond $X=3.07 $Y=1.81
+ $X2=3.067 $Y2=1.645
r88 30 32 30.194 $w=2.48e-07 $l=6.55e-07 $layer=LI1_cond $X=3.07 $Y=1.81
+ $X2=3.07 $Y2=2.465
r89 26 34 6.41553 $w=2.52e-07 $l=1.65e-07 $layer=LI1_cond $X=3.067 $Y=1.48
+ $X2=3.067 $Y2=1.645
r90 26 28 30.0539 $w=2.53e-07 $l=6.65e-07 $layer=LI1_cond $X=3.067 $Y=1.48
+ $X2=3.067 $Y2=0.815
r91 24 37 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.77 $Y=1.645 $X2=2.77
+ $Y2=1.735
r92 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.77
+ $Y=1.645 $X2=2.77 $Y2=1.645
r93 21 34 0.398883 $w=3.3e-07 $l=1.27e-07 $layer=LI1_cond $X=2.94 $Y=1.645
+ $X2=3.067 $Y2=1.645
r94 21 23 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=2.94 $Y=1.645
+ $X2=2.77 $Y2=1.645
r95 19 20 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.205 $Y=1.735
+ $X2=2.13 $Y2=1.735
r96 18 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.605 $Y=1.735
+ $X2=2.77 $Y2=1.735
r97 18 19 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.605 $Y=1.735
+ $X2=2.205 $Y2=1.735
r98 16 20 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.13 $Y=1.81
+ $X2=2.13 $Y2=1.735
r99 16 17 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=2.13 $Y=1.81
+ $X2=2.13 $Y2=2.05
r100 12 20 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.13 $Y=1.66
+ $X2=2.13 $Y2=1.735
r101 12 14 438.415 $w=1.5e-07 $l=8.55e-07 $layer=POLY_cond $X=2.13 $Y=1.66
+ $X2=2.13 $Y2=0.805
r102 10 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.055 $Y=2.125
+ $X2=2.13 $Y2=2.05
r103 10 11 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=2.055 $Y=2.125
+ $X2=1.885 $Y2=2.125
r104 7 11 26.9307 $w=1.5e-07 $l=1.58745e-07 $layer=POLY_cond $X=1.795 $Y=2.245
+ $X2=1.885 $Y2=2.125
r105 7 9 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.795 $Y=2.245
+ $X2=1.795 $Y2=2.64
r106 2 32 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=2.88
+ $Y=2.32 $X2=3.03 $Y2=2.465
r107 1 28 182 $w=1.7e-07 $l=2.81425e-07 $layer=licon1_NDIFF $count=1 $X=2.885
+ $Y=0.595 $X2=3.025 $Y2=0.815
.ends

.subckt PM_SKY130_FD_SC_LS__SDFBBN_2%SCE 4 6 7 9 10 11 12 14 18 19 20 21 22 24
+ 27 28 29 30 34 35
c104 21 0 3.4396e-19 $X=3.175 $Y=2.125
c105 19 0 1.53309e-19 $X=3.175 $Y=1.165
c106 7 0 2.32704e-19 $X=0.955 $Y=2.245
c107 4 0 1.01507e-19 $X=0.91 $Y=0.805
r108 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.97
+ $Y=1.29 $X2=0.97 $Y2=1.29
r109 29 30 8.67743 $w=5.08e-07 $l=3.7e-07 $layer=LI1_cond $X=1.06 $Y=1.295
+ $X2=1.06 $Y2=1.665
r110 29 35 0.117263 $w=5.08e-07 $l=5e-09 $layer=LI1_cond $X=1.06 $Y=1.295
+ $X2=1.06 $Y2=1.29
r111 27 34 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.97 $Y=1.63
+ $X2=0.97 $Y2=1.29
r112 27 28 35.4289 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.97 $Y=1.63
+ $X2=0.97 $Y2=1.795
r113 26 34 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.97 $Y=1.125
+ $X2=0.97 $Y2=1.29
r114 23 24 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=3.25 $Y=1.24
+ $X2=3.25 $Y2=2.05
r115 21 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.175 $Y=2.125
+ $X2=3.25 $Y2=2.05
r116 21 22 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.175 $Y=2.125
+ $X2=2.895 $Y2=2.125
r117 19 23 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.175 $Y=1.165
+ $X2=3.25 $Y2=1.24
r118 19 20 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=3.175 $Y=1.165
+ $X2=2.885 $Y2=1.165
r119 16 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.81 $Y=1.09
+ $X2=2.885 $Y2=1.165
r120 16 18 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.81 $Y=1.09
+ $X2=2.81 $Y2=0.805
r121 15 18 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.81 $Y=0.255
+ $X2=2.81 $Y2=0.805
r122 12 22 26.9307 $w=1.5e-07 $l=1.58745e-07 $layer=POLY_cond $X=2.805 $Y=2.245
+ $X2=2.895 $Y2=2.125
r123 12 14 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.805 $Y=2.245
+ $X2=2.805 $Y2=2.64
r124 10 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.735 $Y=0.18
+ $X2=2.81 $Y2=0.255
r125 10 11 897.34 $w=1.5e-07 $l=1.75e-06 $layer=POLY_cond $X=2.735 $Y=0.18
+ $X2=0.985 $Y2=0.18
r126 7 9 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.955 $Y=2.245
+ $X2=0.955 $Y2=2.64
r127 6 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.955 $Y=2.155
+ $X2=0.955 $Y2=2.245
r128 6 28 139.935 $w=1.8e-07 $l=3.6e-07 $layer=POLY_cond $X=0.955 $Y=2.155
+ $X2=0.955 $Y2=1.795
r129 4 26 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.91 $Y=0.805
+ $X2=0.91 $Y2=1.125
r130 1 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.91 $Y=0.255
+ $X2=0.985 $Y2=0.18
r131 1 4 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.91 $Y=0.255
+ $X2=0.91 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LS__SDFBBN_2%CLK_N 1 3 4 6 7 11
c40 11 0 4.09367e-20 $X=3.73 $Y=1.515
c41 4 0 1.21362e-19 $X=3.815 $Y=1.765
r42 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.73
+ $Y=1.515 $X2=3.73 $Y2=1.515
r43 7 11 4.21625 $w=4.08e-07 $l=1.5e-07 $layer=LI1_cond $X=3.69 $Y=1.665
+ $X2=3.69 $Y2=1.515
r44 4 10 51.8789 $w=3.07e-07 $l=2.87228e-07 $layer=POLY_cond $X=3.815 $Y=1.765
+ $X2=3.735 $Y2=1.515
r45 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.815 $Y=1.765
+ $X2=3.815 $Y2=2.4
r46 1 10 38.5336 $w=3.07e-07 $l=1.94808e-07 $layer=POLY_cond $X=3.8 $Y=1.35
+ $X2=3.735 $Y2=1.515
r47 1 3 157.453 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=3.8 $Y=1.35 $X2=3.8
+ $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_LS__SDFBBN_2%A_1007_366# 1 2 3 10 12 14 15 16 17 19 22
+ 24 26 28 30 31 32 34 36 39 41 45 49 50 53 56 58 61 62 63 67
c198 53 0 3.62521e-20 $X=5.2 $Y=1.995
c199 49 0 1.46444e-19 $X=9.78 $Y=1.745
c200 22 0 8.54043e-20 $X=9.435 $Y=0.9
c201 15 0 8.01569e-20 $X=5.775 $Y=1.195
c202 10 0 1.26757e-20 $X=5.275 $Y=2.245
r203 65 67 1.92074 $w=3.28e-07 $l=5.5e-08 $layer=LI1_cond $X=9.07 $Y=2.21
+ $X2=9.07 $Y2=2.265
r204 63 65 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=9.07 $Y=2.035
+ $X2=9.07 $Y2=2.21
r205 60 61 8.63679 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=8.077 $Y=0.945
+ $X2=8.077 $Y2=1.115
r206 58 59 14.878 $w=2.46e-07 $l=3e-07 $layer=LI1_cond $X=7.66 $Y=2.9 $X2=7.96
+ $Y2=2.9
r207 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.2
+ $Y=1.995 $X2=5.2 $Y2=1.995
r208 50 71 9.74394 $w=3.71e-07 $l=7.5e-08 $layer=POLY_cond $X=9.78 $Y=1.812
+ $X2=9.855 $Y2=1.812
r209 50 69 44.8221 $w=3.71e-07 $l=3.45e-07 $layer=POLY_cond $X=9.78 $Y=1.812
+ $X2=9.435 $Y2=1.812
r210 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.78
+ $Y=1.745 $X2=9.78 $Y2=1.745
r211 47 49 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=9.78 $Y=1.95
+ $X2=9.78 $Y2=1.745
r212 46 63 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.235 $Y=2.035
+ $X2=9.07 $Y2=2.035
r213 45 47 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.615 $Y=2.035
+ $X2=9.78 $Y2=1.95
r214 45 46 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=9.615 $Y=2.035
+ $X2=9.235 $Y2=2.035
r215 42 62 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.045 $Y=2.21
+ $X2=7.96 $Y2=2.21
r216 41 65 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.905 $Y=2.21
+ $X2=9.07 $Y2=2.21
r217 41 42 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=8.905 $Y=2.21
+ $X2=8.045 $Y2=2.21
r218 39 60 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=8.115 $Y=0.86
+ $X2=8.115 $Y2=0.945
r219 36 59 2.90119 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=7.96 $Y=2.73
+ $X2=7.96 $Y2=2.9
r220 35 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.96 $Y=2.295
+ $X2=7.96 $Y2=2.21
r221 35 36 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=7.96 $Y=2.295
+ $X2=7.96 $Y2=2.73
r222 34 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.96 $Y=2.125
+ $X2=7.96 $Y2=2.21
r223 34 61 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=7.96 $Y=2.125
+ $X2=7.96 $Y2=1.115
r224 32 56 8.71323 $w=3.43e-07 $l=1.72e-07 $layer=LI1_cond $X=7.072 $Y=2.902
+ $X2=6.9 $Y2=2.902
r225 31 58 1.26986 $w=3.45e-07 $l=7.93725e-09 $layer=LI1_cond $X=7.653 $Y=2.902
+ $X2=7.66 $Y2=2.9
r226 31 32 19.4078 $w=3.43e-07 $l=5.81e-07 $layer=LI1_cond $X=7.653 $Y=2.902
+ $X2=7.072 $Y2=2.902
r227 30 56 87.7487 $w=1.68e-07 $l=1.345e-06 $layer=LI1_cond $X=5.555 $Y=2.99
+ $X2=6.9 $Y2=2.99
r228 28 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.47 $Y=2.905
+ $X2=5.555 $Y2=2.99
r229 27 53 11.5986 $w=2.84e-07 $l=3.46627e-07 $layer=LI1_cond $X=5.47 $Y=2.18
+ $X2=5.2 $Y2=2.005
r230 27 28 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=5.47 $Y=2.18
+ $X2=5.47 $Y2=2.905
r231 24 71 24.032 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=9.855 $Y=2.045
+ $X2=9.855 $Y2=1.812
r232 24 26 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=9.855 $Y=2.045
+ $X2=9.855 $Y2=2.54
r233 20 69 24.032 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=9.435 $Y=1.58
+ $X2=9.435 $Y2=1.812
r234 20 22 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=9.435 $Y=1.58
+ $X2=9.435 $Y2=0.9
r235 17 19 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=5.85 $Y=1.12
+ $X2=5.85 $Y2=0.835
r236 15 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.775 $Y=1.195
+ $X2=5.85 $Y2=1.12
r237 15 16 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=5.775 $Y=1.195
+ $X2=5.355 $Y2=1.195
r238 14 54 38.5562 $w=2.99e-07 $l=2.0106e-07 $layer=POLY_cond $X=5.28 $Y=1.83
+ $X2=5.2 $Y2=1.995
r239 13 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.28 $Y=1.27
+ $X2=5.355 $Y2=1.195
r240 13 14 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=5.28 $Y=1.27
+ $X2=5.28 $Y2=1.83
r241 10 54 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=5.275 $Y=2.245
+ $X2=5.2 $Y2=1.995
r242 10 12 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=5.275 $Y=2.245
+ $X2=5.275 $Y2=2.53
r243 3 67 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=8.92
+ $Y=2.12 $X2=9.07 $Y2=2.265
r244 2 58 300 $w=1.7e-07 $l=1.03049e-06 $layer=licon1_PDIFF $count=2 $X=6.92
+ $Y=2.12 $X2=7.66 $Y2=2.815
r245 1 39 182 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=1 $X=7.975
+ $Y=0.625 $X2=8.115 $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_LS__SDFBBN_2%A_868_368# 1 2 8 9 11 14 17 18 20 23 27 33
+ 35 41 42 45 46 47 49 50 51 53 54 60 61 64 72 79
c210 79 0 1.26757e-20 $X=5.855 $Y=1.265
c211 72 0 1.62439e-20 $X=10.32 $Y=1.59
c212 64 0 1.15277e-19 $X=5.76 $Y=1.675
c213 54 0 1.27085e-19 $X=6.145 $Y=1.295
c214 53 0 6.70526e-20 $X=10.175 $Y=1.295
c215 49 0 9.35685e-20 $X=6.66 $Y=1.69
c216 23 0 1.08678e-19 $X=11.16 $Y=0.62
r217 73 87 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=10.32 $Y=1.59
+ $X2=10.32 $Y2=1.43
r218 72 75 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.32 $Y=1.59
+ $X2=10.32 $Y2=1.755
r219 72 73 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.32
+ $Y=1.59 $X2=10.32 $Y2=1.59
r220 65 83 0.161011 $w=5.18e-07 $l=7e-09 $layer=LI1_cond $X=5.855 $Y=1.675
+ $X2=5.855 $Y2=1.682
r221 64 67 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.76 $Y=1.675
+ $X2=5.76 $Y2=1.84
r222 64 65 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.76
+ $Y=1.675 $X2=5.76 $Y2=1.675
r223 61 87 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=10.32 $Y=1.295
+ $X2=10.32 $Y2=1.43
r224 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=1.295
+ $X2=10.32 $Y2=1.295
r225 57 65 8.74057 $w=5.18e-07 $l=3.8e-07 $layer=LI1_cond $X=5.855 $Y=1.295
+ $X2=5.855 $Y2=1.675
r226 57 79 0.690045 $w=5.18e-07 $l=3e-08 $layer=LI1_cond $X=5.855 $Y=1.295
+ $X2=5.855 $Y2=1.265
r227 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=1.295 $X2=6
+ $Y2=1.295
r228 54 56 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.145 $Y=1.295
+ $X2=6 $Y2=1.295
r229 53 60 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=10.175 $Y=1.295
+ $X2=10.32 $Y2=1.295
r230 53 54 4.98761 $w=1.4e-07 $l=4.03e-06 $layer=MET1_cond $X=10.175 $Y=1.295
+ $X2=6.145 $Y2=1.295
r231 50 69 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.66 $Y=1.69
+ $X2=6.66 $Y2=1.525
r232 49 51 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=6.66 $Y=1.69
+ $X2=6.495 $Y2=1.69
r233 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.66
+ $Y=1.69 $X2=6.66 $Y2=1.69
r234 45 46 8.5712 $w=3.78e-07 $l=1.65e-07 $layer=LI1_cond $X=4.595 $Y=2.005
+ $X2=4.595 $Y2=1.84
r235 42 77 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=11.22 $Y=1.43
+ $X2=11.22 $Y2=1.265
r236 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.22
+ $Y=1.43 $X2=11.22 $Y2=1.43
r237 39 87 1.29116 $w=3e-07 $l=1.65e-07 $layer=LI1_cond $X=10.485 $Y=1.43
+ $X2=10.32 $Y2=1.43
r238 39 41 28.2349 $w=2.98e-07 $l=7.35e-07 $layer=LI1_cond $X=10.485 $Y=1.43
+ $X2=11.22 $Y2=1.43
r239 38 83 3.68146 $w=3.15e-07 $l=2.6e-07 $layer=LI1_cond $X=6.115 $Y=1.682
+ $X2=5.855 $Y2=1.682
r240 38 51 13.9025 $w=3.13e-07 $l=3.8e-07 $layer=LI1_cond $X=6.115 $Y=1.682
+ $X2=6.495 $Y2=1.682
r241 36 47 2.11342 $w=1.7e-07 $l=1.63e-07 $layer=LI1_cond $X=4.94 $Y=1.265
+ $X2=4.777 $Y2=1.265
r242 35 79 7.40362 $w=1.7e-07 $l=2.6e-07 $layer=LI1_cond $X=5.595 $Y=1.265
+ $X2=5.855 $Y2=1.265
r243 35 36 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=5.595 $Y=1.265
+ $X2=4.94 $Y2=1.265
r244 31 47 4.3182 $w=2.1e-07 $l=1.0225e-07 $layer=LI1_cond $X=4.815 $Y=1.18
+ $X2=4.777 $Y2=1.265
r245 31 33 19.361 $w=2.48e-07 $l=4.2e-07 $layer=LI1_cond $X=4.815 $Y=1.18
+ $X2=4.815 $Y2=0.76
r246 29 47 4.3182 $w=2.1e-07 $l=1.17346e-07 $layer=LI1_cond $X=4.7 $Y=1.35
+ $X2=4.777 $Y2=1.265
r247 29 46 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=4.7 $Y=1.35 $X2=4.7
+ $Y2=1.84
r248 25 45 0.758186 $w=3.78e-07 $l=2.5e-08 $layer=LI1_cond $X=4.595 $Y=2.03
+ $X2=4.595 $Y2=2.005
r249 25 27 23.807 $w=3.78e-07 $l=7.85e-07 $layer=LI1_cond $X=4.595 $Y=2.03
+ $X2=4.595 $Y2=2.815
r250 23 77 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=11.16 $Y=0.62
+ $X2=11.16 $Y2=1.265
r251 18 20 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=10.245 $Y=2.045
+ $X2=10.245 $Y2=2.54
r252 17 18 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=10.245 $Y=1.955
+ $X2=10.245 $Y2=2.045
r253 17 75 77.7419 $w=1.8e-07 $l=2e-07 $layer=POLY_cond $X=10.245 $Y=1.955
+ $X2=10.245 $Y2=1.755
r254 14 69 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.665 $Y=0.835
+ $X2=6.665 $Y2=1.525
r255 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=5.695 $Y=2.245
+ $X2=5.695 $Y2=2.53
r256 8 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.695 $Y=2.155
+ $X2=5.695 $Y2=2.245
r257 8 67 122.444 $w=1.8e-07 $l=3.15e-07 $layer=POLY_cond $X=5.695 $Y=2.155
+ $X2=5.695 $Y2=1.84
r258 2 45 400 $w=1.7e-07 $l=2.2798e-07 $layer=licon1_PDIFF $count=1 $X=4.34
+ $Y=1.84 $X2=4.49 $Y2=2.005
r259 2 27 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=4.34
+ $Y=1.84 $X2=4.49 $Y2=2.815
r260 1 33 91 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_NDIFF $count=2 $X=4.715
+ $Y=0.49 $X2=4.855 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_LS__SDFBBN_2%A_1154_464# 1 2 7 8 10 11 13 14 16 18 21 23
+ 24 27 29 30 34 35
c102 30 0 8.01569e-20 $X=6.615 $Y=1.27
c103 27 0 1.27085e-19 $X=6.45 $Y=0.835
c104 8 0 6.70526e-20 $X=7.365 $Y=1.36
r105 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.2
+ $Y=1.45 $X2=7.2 $Y2=1.45
r106 32 34 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=7.2 $Y=2.04 $X2=7.2
+ $Y2=1.45
r107 31 34 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=7.2 $Y=1.355
+ $X2=7.2 $Y2=1.45
r108 29 31 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.035 $Y=1.27
+ $X2=7.2 $Y2=1.355
r109 29 30 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=7.035 $Y=1.27
+ $X2=6.615 $Y2=1.27
r110 25 30 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.45 $Y=1.185
+ $X2=6.615 $Y2=1.27
r111 25 27 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=6.45 $Y=1.185
+ $X2=6.45 $Y2=0.835
r112 23 32 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.035 $Y=2.125
+ $X2=7.2 $Y2=2.04
r113 23 24 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=7.035 $Y=2.125
+ $X2=6.17 $Y2=2.125
r114 19 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.005 $Y=2.21
+ $X2=6.17 $Y2=2.125
r115 19 21 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=6.005 $Y=2.21
+ $X2=6.005 $Y2=2.515
r116 17 35 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=7.2 $Y=1.435
+ $X2=7.2 $Y2=1.45
r117 14 18 18.8402 $w=1.65e-07 $l=8.21584e-08 $layer=POLY_cond $X=7.9 $Y=1.285
+ $X2=7.885 $Y2=1.36
r118 14 16 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=7.9 $Y=1.285
+ $X2=7.9 $Y2=0.9
r119 11 13 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=7.885 $Y=2.045
+ $X2=7.885 $Y2=2.54
r120 10 11 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=7.885 $Y=1.955
+ $X2=7.885 $Y2=2.045
r121 9 18 18.8402 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=7.885 $Y=1.435
+ $X2=7.885 $Y2=1.36
r122 9 10 202.129 $w=1.8e-07 $l=5.2e-07 $layer=POLY_cond $X=7.885 $Y=1.435
+ $X2=7.885 $Y2=1.955
r123 8 17 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=7.365 $Y=1.36
+ $X2=7.2 $Y2=1.435
r124 7 18 6.66866 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=7.795 $Y=1.36
+ $X2=7.885 $Y2=1.36
r125 7 8 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=7.795 $Y=1.36
+ $X2=7.365 $Y2=1.36
r126 2 21 600 $w=1.7e-07 $l=3.17884e-07 $layer=licon1_PDIFF $count=1 $X=5.77
+ $Y=2.32 $X2=6.005 $Y2=2.515
r127 1 27 182 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_NDIFF $count=1 $X=6.285
+ $Y=0.625 $X2=6.45 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_LS__SDFBBN_2%A_1643_257# 1 2 7 9 12 14 17 18 20 22 23 26
+ 29 30 31 33 34 35 36 40 43 46 50 51 52 56 57 60 62 66 70
c205 70 0 1.11129e-19 $X=12.66 $Y=1.22
c206 57 0 1.91513e-19 $X=12.66 $Y=1.13
c207 56 0 1.28025e-19 $X=12.66 $Y=1.215
c208 31 0 7.74904e-20 $X=9.725 $Y=0.345
r209 63 66 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=13.69 $Y=2.17
+ $X2=13.91 $Y2=2.17
r210 60 71 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=12.66 $Y=1.385
+ $X2=12.66 $Y2=1.55
r211 60 70 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=12.66 $Y=1.385
+ $X2=12.66 $Y2=1.22
r212 59 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.66
+ $Y=1.385 $X2=12.66 $Y2=1.385
r213 56 59 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=12.66 $Y=1.215
+ $X2=12.66 $Y2=1.385
r214 56 57 5.66838 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=12.66 $Y=1.215
+ $X2=12.66 $Y2=1.13
r215 52 54 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=11.98 $Y=0.685
+ $X2=11.98 $Y2=0.855
r216 50 51 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.38
+ $Y=1.45 $X2=8.38 $Y2=1.45
r217 44 62 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=13.775 $Y=1.17
+ $X2=13.69 $Y2=1.17
r218 44 46 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=13.775 $Y=1.17
+ $X2=13.985 $Y2=1.17
r219 43 63 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.69 $Y=2.005
+ $X2=13.69 $Y2=2.17
r220 42 62 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.69 $Y=1.335
+ $X2=13.69 $Y2=1.17
r221 42 43 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=13.69 $Y=1.335
+ $X2=13.69 $Y2=2.005
r222 41 56 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.825 $Y=1.215
+ $X2=12.66 $Y2=1.215
r223 40 62 3.70735 $w=2.5e-07 $l=1.05119e-07 $layer=LI1_cond $X=13.605 $Y=1.215
+ $X2=13.69 $Y2=1.17
r224 40 41 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=13.605 $Y=1.215
+ $X2=12.825 $Y2=1.215
r225 38 57 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=12.58 $Y=0.94
+ $X2=12.58 $Y2=1.13
r226 37 54 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.065 $Y=0.855
+ $X2=11.98 $Y2=0.855
r227 36 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=12.495 $Y=0.855
+ $X2=12.58 $Y2=0.94
r228 36 37 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=12.495 $Y=0.855
+ $X2=12.065 $Y2=0.855
r229 34 52 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.895 $Y=0.685
+ $X2=11.98 $Y2=0.685
r230 34 35 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=11.895 $Y=0.685
+ $X2=11.51 $Y2=0.685
r231 33 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.425 $Y=0.6
+ $X2=11.51 $Y2=0.685
r232 32 33 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=11.425 $Y=0.43
+ $X2=11.425 $Y2=0.6
r233 30 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.34 $Y=0.345
+ $X2=11.425 $Y2=0.43
r234 30 31 105.364 $w=1.68e-07 $l=1.615e-06 $layer=LI1_cond $X=11.34 $Y=0.345
+ $X2=9.725 $Y2=0.345
r235 28 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.64 $Y=0.43
+ $X2=9.725 $Y2=0.345
r236 28 29 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=9.64 $Y=0.43
+ $X2=9.64 $Y2=1.11
r237 27 50 10.5458 $w=2.95e-07 $l=3.41746e-07 $layer=LI1_cond $X=8.62 $Y=1.195
+ $X2=8.417 $Y2=1.45
r238 26 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.555 $Y=1.195
+ $X2=9.64 $Y2=1.11
r239 26 27 61 $w=1.68e-07 $l=9.35e-07 $layer=LI1_cond $X=9.555 $Y=1.195 $X2=8.62
+ $Y2=1.195
r240 23 51 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=8.38 $Y=1.79
+ $X2=8.38 $Y2=1.45
r241 22 51 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.38 $Y=1.285
+ $X2=8.38 $Y2=1.45
r242 18 20 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=12.705 $Y=1.885
+ $X2=12.705 $Y2=2.46
r243 17 70 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=12.705 $Y=0.74
+ $X2=12.705 $Y2=1.22
r244 14 18 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=12.705 $Y=1.795
+ $X2=12.705 $Y2=1.885
r245 14 71 95.2339 $w=1.8e-07 $l=2.45e-07 $layer=POLY_cond $X=12.705 $Y=1.795
+ $X2=12.705 $Y2=1.55
r246 12 22 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=8.33 $Y=0.9
+ $X2=8.33 $Y2=1.285
r247 7 23 44.3718 $w=2.77e-07 $l=2.90086e-07 $layer=POLY_cond $X=8.305 $Y=2.045
+ $X2=8.38 $Y2=1.79
r248 7 9 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=8.305 $Y=2.045
+ $X2=8.305 $Y2=2.54
r249 2 66 600 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=13.765
+ $Y=1.995 $X2=13.91 $Y2=2.17
r250 1 46 182 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_NDIFF $count=1 $X=13.845
+ $Y=0.9 $X2=13.985 $Y2=1.17
.ends

.subckt PM_SKY130_FD_SC_LS__SDFBBN_2%SET_B 2 3 5 8 11 14 15 17 18 19 22 24 27 32
+ 33 34
c140 34 0 1.96837e-19 $X=12.12 $Y=1.22
c141 33 0 1.11129e-19 $X=12.12 $Y=1.385
c142 27 0 1.46444e-19 $X=8.955 $Y=1.615
c143 18 0 1.44347e-19 $X=12.095 $Y=1.665
r144 33 43 8.72119 $w=3.68e-07 $l=2.8e-07 $layer=LI1_cond $X=12.14 $Y=1.385
+ $X2=12.14 $Y2=1.665
r145 32 35 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=12.12 $Y=1.385
+ $X2=12.12 $Y2=1.55
r146 32 34 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=12.12 $Y=1.385
+ $X2=12.12 $Y2=1.22
r147 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.12
+ $Y=1.385 $X2=12.12 $Y2=1.385
r148 27 30 40.9207 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=8.937 $Y=1.615
+ $X2=8.937 $Y2=1.78
r149 27 29 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=8.937 $Y=1.615
+ $X2=8.937 $Y2=1.45
r150 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.955
+ $Y=1.615 $X2=8.955 $Y2=1.615
r151 24 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=1.665
+ $X2=12.24 $Y2=1.665
r152 22 28 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=9.36 $Y=1.615
+ $X2=8.955 $Y2=1.615
r153 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=1.665
+ $X2=9.36 $Y2=1.665
r154 19 21 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.505 $Y=1.665
+ $X2=9.36 $Y2=1.665
r155 18 24 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=12.095 $Y=1.665
+ $X2=12.24 $Y2=1.665
r156 18 19 3.20544 $w=1.4e-07 $l=2.59e-06 $layer=MET1_cond $X=12.095 $Y=1.665
+ $X2=9.505 $Y2=1.665
r157 15 17 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=12.195 $Y=1.885
+ $X2=12.195 $Y2=2.46
r158 14 34 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=12.185 $Y=0.74
+ $X2=12.185 $Y2=1.22
r159 11 15 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=12.195 $Y=1.795
+ $X2=12.195 $Y2=1.885
r160 11 35 95.2339 $w=1.8e-07 $l=2.45e-07 $layer=POLY_cond $X=12.195 $Y=1.795
+ $X2=12.195 $Y2=1.55
r161 8 29 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=8.935 $Y=0.9
+ $X2=8.935 $Y2=1.45
r162 3 5 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=8.845 $Y=2.045
+ $X2=8.845 $Y2=2.54
r163 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=8.845 $Y=1.955
+ $X2=8.845 $Y2=2.045
r164 2 30 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=8.845 $Y=1.955
+ $X2=8.845 $Y2=1.78
.ends

.subckt PM_SKY130_FD_SC_LS__SDFBBN_2%A_688_98# 1 2 7 9 13 14 15 19 22 23 28 29
+ 30 31 32 35 37 38 40 41 42 46 48 50 55 59 60 61
c181 60 0 1.36467e-19 $X=4.28 $Y=1.505
c182 31 0 1.21918e-19 $X=10.78 $Y=2.085
c183 19 0 9.35685e-20 $X=6.21 $Y=0.835
c184 7 0 4.09367e-20 $X=4.265 $Y=1.765
r185 60 65 48.4693 $w=3.58e-07 $l=3.6e-07 $layer=POLY_cond $X=4.28 $Y=1.552
+ $X2=4.64 $Y2=1.552
r186 60 63 2.01955 $w=3.58e-07 $l=1.5e-08 $layer=POLY_cond $X=4.28 $Y=1.552
+ $X2=4.265 $Y2=1.552
r187 59 62 8.5712 $w=3.78e-07 $l=1.65e-07 $layer=LI1_cond $X=4.255 $Y=1.505
+ $X2=4.255 $Y2=1.67
r188 59 61 8.5712 $w=3.78e-07 $l=1.65e-07 $layer=LI1_cond $X=4.255 $Y=1.505
+ $X2=4.255 $Y2=1.34
r189 59 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.28
+ $Y=1.505 $X2=4.28 $Y2=1.505
r190 55 62 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=4.15 $Y=1.95
+ $X2=4.15 $Y2=1.67
r191 52 61 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.15 $Y=1.17
+ $X2=4.15 $Y2=1.34
r192 51 57 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.675 $Y=2.035
+ $X2=3.55 $Y2=2.035
r193 50 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.065 $Y=2.035
+ $X2=4.15 $Y2=1.95
r194 50 51 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=4.065 $Y=2.035
+ $X2=3.675 $Y2=2.035
r195 46 57 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.55 $Y=2.12
+ $X2=3.55 $Y2=2.035
r196 46 48 32.0379 $w=2.48e-07 $l=6.95e-07 $layer=LI1_cond $X=3.55 $Y=2.12
+ $X2=3.55 $Y2=2.815
r197 42 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.065 $Y=1.085
+ $X2=4.15 $Y2=1.17
r198 42 44 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=4.065 $Y=1.085
+ $X2=3.585 $Y2=1.085
r199 39 40 55.4135 $w=1.85e-07 $l=1.5e-07 $layer=POLY_cond $X=6.227 $Y=2.095
+ $X2=6.227 $Y2=2.245
r200 35 37 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=10.78 $Y=2.465
+ $X2=10.78 $Y2=2.75
r201 33 41 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=10.77 $Y=1.185
+ $X2=10.77 $Y2=1.995
r202 32 35 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=10.78 $Y=2.375
+ $X2=10.78 $Y2=2.465
r203 31 41 36.5962 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=10.78 $Y=2.085
+ $X2=10.78 $Y2=1.995
r204 31 32 112.726 $w=1.8e-07 $l=2.9e-07 $layer=POLY_cond $X=10.78 $Y=2.085
+ $X2=10.78 $Y2=2.375
r205 29 33 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.695 $Y=1.11
+ $X2=10.77 $Y2=1.185
r206 29 30 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=10.695 $Y=1.11
+ $X2=9.985 $Y2=1.11
r207 26 30 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.91 $Y=1.035
+ $X2=9.985 $Y2=1.11
r208 26 28 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=9.91 $Y=1.035
+ $X2=9.91 $Y2=0.685
r209 25 28 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=9.91 $Y=0.255
+ $X2=9.91 $Y2=0.685
r210 24 38 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.285 $Y=0.18
+ $X2=6.21 $Y2=0.18
r211 23 25 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.835 $Y=0.18
+ $X2=9.91 $Y2=0.255
r212 23 24 1820.32 $w=1.5e-07 $l=3.55e-06 $layer=POLY_cond $X=9.835 $Y=0.18
+ $X2=6.285 $Y2=0.18
r213 22 40 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=6.23 $Y=2.64
+ $X2=6.23 $Y2=2.245
r214 19 39 646.085 $w=1.5e-07 $l=1.26e-06 $layer=POLY_cond $X=6.21 $Y=0.835
+ $X2=6.21 $Y2=2.095
r215 16 38 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.21 $Y=0.255
+ $X2=6.21 $Y2=0.18
r216 16 19 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.21 $Y=0.255
+ $X2=6.21 $Y2=0.835
r217 14 38 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.135 $Y=0.18
+ $X2=6.21 $Y2=0.18
r218 14 15 728.128 $w=1.5e-07 $l=1.42e-06 $layer=POLY_cond $X=6.135 $Y=0.18
+ $X2=4.715 $Y2=0.18
r219 11 65 23.1716 $w=1.5e-07 $l=2.12e-07 $layer=POLY_cond $X=4.64 $Y=1.34
+ $X2=4.64 $Y2=1.552
r220 11 13 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.64 $Y=1.34
+ $X2=4.64 $Y2=0.86
r221 10 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.64 $Y=0.255
+ $X2=4.715 $Y2=0.18
r222 10 13 310.223 $w=1.5e-07 $l=6.05e-07 $layer=POLY_cond $X=4.64 $Y=0.255
+ $X2=4.64 $Y2=0.86
r223 7 63 23.1716 $w=1.5e-07 $l=2.13e-07 $layer=POLY_cond $X=4.265 $Y=1.765
+ $X2=4.265 $Y2=1.552
r224 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.265 $Y=1.765
+ $X2=4.265 $Y2=2.4
r225 2 57 400 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=3.445
+ $Y=1.84 $X2=3.59 $Y2=2.115
r226 2 48 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=3.445
+ $Y=1.84 $X2=3.59 $Y2=2.815
r227 1 44 182 $w=1.7e-07 $l=6.63551e-07 $layer=licon1_NDIFF $count=1 $X=3.44
+ $Y=0.49 $X2=3.585 $Y2=1.085
.ends

.subckt PM_SKY130_FD_SC_LS__SDFBBN_2%A_2216_410# 1 2 3 10 12 13 15 17 19 20 24
+ 26 28 31 33 35 36 37 40 42 44 47 54 58 60 64 66 68 71 73 79 83 85 91 93 97
c208 47 0 7.20841e-20 $X=11.67 $Y=0.98
c209 19 0 2.75443e-20 $X=11.67 $Y=2.05
r210 92 97 10.142 $w=3.3e-07 $l=5.8e-08 $layer=POLY_cond $X=14.65 $Y=1.595
+ $X2=14.65 $Y2=1.537
r211 91 94 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=14.65 $Y=1.595
+ $X2=14.65 $Y2=1.76
r212 91 93 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=14.65 $Y=1.595
+ $X2=14.65 $Y2=1.43
r213 91 92 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=14.65
+ $Y=1.595 $X2=14.65 $Y2=1.595
r214 87 88 11.2939 $w=2.48e-07 $l=2.45e-07 $layer=LI1_cond $X=13.31 $Y=2.345
+ $X2=13.31 $Y2=2.59
r215 85 87 5.53173 $w=2.48e-07 $l=1.2e-07 $layer=LI1_cond $X=13.31 $Y=2.225
+ $X2=13.31 $Y2=2.345
r216 81 83 8.52431 $w=3.63e-07 $l=1.65e-07 $layer=LI1_cond $X=12.92 $Y=0.777
+ $X2=13.085 $Y2=0.777
r217 74 95 14.5084 $w=2.99e-07 $l=9e-08 $layer=POLY_cond $X=11.245 $Y=2.215
+ $X2=11.245 $Y2=2.125
r218 73 76 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=11.245 $Y=2.215
+ $X2=11.245 $Y2=2.345
r219 73 74 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.245
+ $Y=2.215 $X2=11.245 $Y2=2.215
r220 71 94 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=14.57 $Y=2.505
+ $X2=14.57 $Y2=1.76
r221 68 89 13.6427 $w=2.52e-07 $l=2.93581e-07 $layer=LI1_cond $X=14.57 $Y=1.005
+ $X2=14.487 $Y2=0.75
r222 68 93 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=14.57 $Y=1.005
+ $X2=14.57 $Y2=1.43
r223 67 88 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.435 $Y=2.59
+ $X2=13.31 $Y2=2.59
r224 66 71 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=14.485 $Y=2.59
+ $X2=14.57 $Y2=2.505
r225 66 67 68.5027 $w=1.68e-07 $l=1.05e-06 $layer=LI1_cond $X=14.485 $Y=2.59
+ $X2=13.435 $Y2=2.59
r226 62 88 3.91831 $w=2.48e-07 $l=8.5e-08 $layer=LI1_cond $X=13.31 $Y=2.675
+ $X2=13.31 $Y2=2.59
r227 62 64 6.45368 $w=2.48e-07 $l=1.4e-07 $layer=LI1_cond $X=13.31 $Y=2.675
+ $X2=13.31 $Y2=2.815
r228 60 89 3.04159 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=14.32 $Y=0.75
+ $X2=14.487 $Y2=0.75
r229 60 83 80.5722 $w=1.68e-07 $l=1.235e-06 $layer=LI1_cond $X=14.32 $Y=0.75
+ $X2=13.085 $Y2=0.75
r230 59 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.135 $Y=2.345
+ $X2=11.97 $Y2=2.345
r231 58 87 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.185 $Y=2.345
+ $X2=13.31 $Y2=2.345
r232 58 59 68.5027 $w=1.68e-07 $l=1.05e-06 $layer=LI1_cond $X=13.185 $Y=2.345
+ $X2=12.135 $Y2=2.345
r233 55 76 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.41 $Y=2.345
+ $X2=11.245 $Y2=2.345
r234 54 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.805 $Y=2.345
+ $X2=11.97 $Y2=2.345
r235 54 55 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=11.805 $Y=2.345
+ $X2=11.41 $Y2=2.345
r236 51 52 14.2163 $w=3.56e-07 $l=1.05e-07 $layer=POLY_cond $X=15.66 $Y=1.557
+ $X2=15.765 $Y2=1.557
r237 50 51 46.7107 $w=3.56e-07 $l=3.45e-07 $layer=POLY_cond $X=15.315 $Y=1.557
+ $X2=15.66 $Y2=1.557
r238 49 50 11.5084 $w=3.56e-07 $l=8.5e-08 $layer=POLY_cond $X=15.23 $Y=1.557
+ $X2=15.315 $Y2=1.557
r239 45 47 61.5319 $w=1.5e-07 $l=1.2e-07 $layer=POLY_cond $X=11.55 $Y=0.98
+ $X2=11.67 $Y2=0.98
r240 42 44 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=16.76 $Y=1.845
+ $X2=16.76 $Y2=2.42
r241 38 40 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=16.72 $Y=1.35
+ $X2=16.72 $Y2=0.79
r242 37 52 13.7431 $w=3.56e-07 $l=1.16189e-07 $layer=POLY_cond $X=15.855
+ $Y=1.497 $X2=15.765 $Y2=1.557
r243 36 42 95.1138 $w=1.79e-07 $l=3.5444e-07 $layer=POLY_cond $X=16.747 $Y=1.497
+ $X2=16.76 $Y2=1.845
r244 36 38 40.9898 $w=1.79e-07 $l=1.59931e-07 $layer=POLY_cond $X=16.747
+ $Y=1.497 $X2=16.72 $Y2=1.35
r245 36 37 160.643 $w=2.95e-07 $l=7.9e-07 $layer=POLY_cond $X=16.645 $Y=1.497
+ $X2=15.855 $Y2=1.497
r246 33 52 23.0368 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=15.765 $Y=1.765
+ $X2=15.765 $Y2=1.557
r247 33 35 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=15.765 $Y=1.765
+ $X2=15.765 $Y2=2.4
r248 29 51 23.0368 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=15.66 $Y=1.35
+ $X2=15.66 $Y2=1.557
r249 29 31 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=15.66 $Y=1.35
+ $X2=15.66 $Y2=0.74
r250 26 50 23.0368 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=15.315 $Y=1.765
+ $X2=15.315 $Y2=1.557
r251 26 28 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=15.315 $Y=1.765
+ $X2=15.315 $Y2=2.4
r252 22 49 23.0368 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=15.23 $Y=1.35
+ $X2=15.23 $Y2=1.557
r253 22 24 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=15.23 $Y=1.35
+ $X2=15.23 $Y2=0.74
r254 21 97 12.8918 $w=2.15e-07 $l=1.65e-07 $layer=POLY_cond $X=14.815 $Y=1.537
+ $X2=14.65 $Y2=1.537
r255 20 49 17.6588 $w=3.56e-07 $l=8.44097e-08 $layer=POLY_cond $X=15.155
+ $Y=1.537 $X2=15.23 $Y2=1.557
r256 20 21 101.481 $w=2.15e-07 $l=3.4e-07 $layer=POLY_cond $X=15.155 $Y=1.537
+ $X2=14.815 $Y2=1.537
r257 18 47 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.67 $Y=1.055
+ $X2=11.67 $Y2=0.98
r258 18 19 510.202 $w=1.5e-07 $l=9.95e-07 $layer=POLY_cond $X=11.67 $Y=1.055
+ $X2=11.67 $Y2=2.05
r259 15 45 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.55 $Y=0.905
+ $X2=11.55 $Y2=0.98
r260 15 17 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=11.55 $Y=0.905
+ $X2=11.55 $Y2=0.62
r261 14 95 18.89 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.41 $Y=2.125
+ $X2=11.245 $Y2=2.125
r262 13 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=11.595 $Y=2.125
+ $X2=11.67 $Y2=2.05
r263 13 14 94.8617 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=11.595 $Y=2.125
+ $X2=11.41 $Y2=2.125
r264 10 74 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=11.17 $Y=2.465
+ $X2=11.245 $Y2=2.215
r265 10 12 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=11.17 $Y=2.465
+ $X2=11.17 $Y2=2.75
r266 3 85 600 $w=1.7e-07 $l=3.31625e-07 $layer=licon1_PDIFF $count=1 $X=13.2
+ $Y=1.96 $X2=13.35 $Y2=2.225
r267 3 64 600 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=13.2
+ $Y=1.96 $X2=13.35 $Y2=2.815
r268 2 79 300 $w=1.7e-07 $l=5.32588e-07 $layer=licon1_PDIFF $count=2 $X=11.825
+ $Y=1.96 $X2=11.97 $Y2=2.425
r269 1 81 182 $w=1.7e-07 $l=4.69814e-07 $layer=licon1_NDIFF $count=1 $X=12.78
+ $Y=0.37 $X2=12.92 $Y2=0.775
.ends

.subckt PM_SKY130_FD_SC_LS__SDFBBN_2%A_1997_82# 1 2 7 9 12 20 23 24 25 26 29 30
+ 32 37 40 44 46 51
c160 40 0 1.85877e-19 $X=10.945 $Y=0.685
c161 25 0 1.62439e-20 $X=10.91 $Y=1.835
r162 51 54 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=13.2 $Y=1.635
+ $X2=13.2 $Y2=1.805
r163 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.2
+ $Y=1.635 $X2=13.2 $Y2=1.635
r164 46 48 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=12.58 $Y=1.805
+ $X2=12.58 $Y2=2.005
r165 44 45 11.3956 $w=1.82e-07 $l=1.7e-07 $layer=LI1_cond $X=11.652 $Y=1.835
+ $X2=11.652 $Y2=2.005
r166 40 42 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=11.025 $Y=0.685
+ $X2=11.025 $Y2=1.025
r167 35 37 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=10.47 $Y=2.185
+ $X2=10.825 $Y2=2.185
r168 33 46 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.665 $Y=1.805
+ $X2=12.58 $Y2=1.805
r169 32 54 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.035 $Y=1.805
+ $X2=13.2 $Y2=1.805
r170 32 33 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=13.035 $Y=1.805
+ $X2=12.665 $Y2=1.805
r171 31 45 1.129 $w=1.7e-07 $l=9.8e-08 $layer=LI1_cond $X=11.75 $Y=2.005
+ $X2=11.652 $Y2=2.005
r172 30 48 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.495 $Y=2.005
+ $X2=12.58 $Y2=2.005
r173 30 31 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=12.495 $Y=2.005
+ $X2=11.75 $Y2=2.005
r174 29 44 5.7679 $w=1.82e-07 $l=9.0802e-08 $layer=LI1_cond $X=11.64 $Y=1.75
+ $X2=11.652 $Y2=1.835
r175 28 29 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=11.64 $Y=1.11
+ $X2=11.64 $Y2=1.75
r176 27 42 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.11 $Y=1.025
+ $X2=11.025 $Y2=1.025
r177 26 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.555 $Y=1.025
+ $X2=11.64 $Y2=1.11
r178 26 27 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=11.555 $Y=1.025
+ $X2=11.11 $Y2=1.025
r179 24 44 1.129 $w=1.7e-07 $l=9.7e-08 $layer=LI1_cond $X=11.555 $Y=1.835
+ $X2=11.652 $Y2=1.835
r180 24 25 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=11.555 $Y=1.835
+ $X2=10.91 $Y2=1.835
r181 23 37 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.825 $Y=2.1
+ $X2=10.825 $Y2=2.185
r182 22 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.825 $Y=1.92
+ $X2=10.91 $Y2=1.835
r183 22 23 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=10.825 $Y=1.92
+ $X2=10.825 $Y2=2.1
r184 20 35 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=10.47 $Y=2.815
+ $X2=10.47 $Y2=2.27
r185 16 40 37.5696 $w=2.48e-07 $l=8.15e-07 $layer=LI1_cond $X=10.125 $Y=0.725
+ $X2=10.94 $Y2=0.725
r186 10 52 38.5562 $w=2.99e-07 $l=1.94808e-07 $layer=POLY_cond $X=13.135 $Y=1.47
+ $X2=13.2 $Y2=1.635
r187 10 12 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=13.135 $Y=1.47
+ $X2=13.135 $Y2=0.74
r188 7 52 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=13.125 $Y=1.885
+ $X2=13.2 $Y2=1.635
r189 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=13.125 $Y=1.885
+ $X2=13.125 $Y2=2.46
r190 2 35 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=10.32
+ $Y=2.12 $X2=10.47 $Y2=2.265
r191 2 20 600 $w=1.7e-07 $l=7.66339e-07 $layer=licon1_PDIFF $count=1 $X=10.32
+ $Y=2.12 $X2=10.47 $Y2=2.815
r192 1 40 91 $w=1.7e-07 $l=1.08885e-06 $layer=licon1_NDIFF $count=2 $X=9.985
+ $Y=0.41 $X2=10.945 $Y2=0.685
r193 1 16 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=9.985
+ $Y=0.41 $X2=10.125 $Y2=0.685
.ends

.subckt PM_SKY130_FD_SC_LS__SDFBBN_2%RESET_B 1 3 6 8
r32 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=14.11
+ $Y=1.67 $X2=14.11 $Y2=1.67
r33 4 11 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=14.2 $Y=1.505
+ $X2=14.11 $Y2=1.67
r34 4 6 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=14.2 $Y=1.505
+ $X2=14.2 $Y2=1.11
r35 1 11 52.2586 $w=2.99e-07 $l=2.62202e-07 $layer=POLY_cond $X=14.135 $Y=1.92
+ $X2=14.11 $Y2=1.67
r36 1 3 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=14.135 $Y=1.92
+ $X2=14.135 $Y2=2.315
.ends

.subckt PM_SKY130_FD_SC_LS__SDFBBN_2%A_3272_94# 1 2 7 9 10 12 13 15 16 18 21 25
+ 31 34 38
c66 25 0 1.7776e-19 $X=16.535 $Y=2.065
c67 7 0 1.00299e-19 $X=17.285 $Y=1.765
r68 38 39 1.69321 $w=4.27e-07 $l=1.5e-08 $layer=POLY_cond $X=17.735 $Y=1.492
+ $X2=17.75 $Y2=1.492
r69 37 38 46.8454 $w=4.27e-07 $l=4.15e-07 $layer=POLY_cond $X=17.32 $Y=1.492
+ $X2=17.735 $Y2=1.492
r70 36 37 3.95082 $w=4.27e-07 $l=3.5e-08 $layer=POLY_cond $X=17.285 $Y=1.492
+ $X2=17.32 $Y2=1.492
r71 32 36 9.59485 $w=4.27e-07 $l=8.5e-08 $layer=POLY_cond $X=17.2 $Y=1.492
+ $X2=17.285 $Y2=1.492
r72 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=17.2
+ $Y=1.385 $X2=17.2 $Y2=1.385
r73 29 34 1.50311 $w=3.3e-07 $l=1.8e-07 $layer=LI1_cond $X=16.7 $Y=1.385
+ $X2=16.52 $Y2=1.385
r74 29 31 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=16.7 $Y=1.385 $X2=17.2
+ $Y2=1.385
r75 25 27 22.7287 $w=3.58e-07 $l=7.1e-07 $layer=LI1_cond $X=16.52 $Y=2.065
+ $X2=16.52 $Y2=2.775
r76 23 34 4.97762 $w=3.45e-07 $l=1.65e-07 $layer=LI1_cond $X=16.52 $Y=1.55
+ $X2=16.52 $Y2=1.385
r77 23 25 16.4863 $w=3.58e-07 $l=5.15e-07 $layer=LI1_cond $X=16.52 $Y=1.55
+ $X2=16.52 $Y2=2.065
r78 19 34 4.97762 $w=3.45e-07 $l=1.72337e-07 $layer=LI1_cond $X=16.505 $Y=1.22
+ $X2=16.52 $Y2=1.385
r79 19 21 20.0804 $w=3.28e-07 $l=5.75e-07 $layer=LI1_cond $X=16.505 $Y=1.22
+ $X2=16.505 $Y2=0.645
r80 16 39 27.4666 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=17.75 $Y=1.22
+ $X2=17.75 $Y2=1.492
r81 16 18 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=17.75 $Y=1.22
+ $X2=17.75 $Y2=0.74
r82 13 38 27.4666 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=17.735 $Y=1.765
+ $X2=17.735 $Y2=1.492
r83 13 15 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=17.735 $Y=1.765
+ $X2=17.735 $Y2=2.4
r84 10 37 27.4666 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=17.32 $Y=1.22
+ $X2=17.32 $Y2=1.492
r85 10 12 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=17.32 $Y=1.22
+ $X2=17.32 $Y2=0.74
r86 7 36 27.4666 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=17.285 $Y=1.765
+ $X2=17.285 $Y2=1.492
r87 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=17.285 $Y=1.765
+ $X2=17.285 $Y2=2.4
r88 2 27 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=16.395
+ $Y=1.92 $X2=16.535 $Y2=2.775
r89 2 25 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=16.395
+ $Y=1.92 $X2=16.535 $Y2=2.065
r90 1 21 91 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_NDIFF $count=2 $X=16.36
+ $Y=0.47 $X2=16.505 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_LS__SDFBBN_2%A_27_464# 1 2 9 12 13 14 17 20
c41 9 0 2.57379e-20 $X=1.065 $Y=2.39
r42 15 17 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=2.02 $Y=2.905
+ $X2=2.02 $Y2=2.465
r43 13 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.855 $Y=2.99
+ $X2=2.02 $Y2=2.905
r44 13 14 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=1.855 $Y=2.99
+ $X2=1.235 $Y2=2.99
r45 12 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.15 $Y=2.905
+ $X2=1.235 $Y2=2.99
r46 11 12 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=1.15 $Y=2.475
+ $X2=1.15 $Y2=2.905
r47 10 20 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.365 $Y=2.39
+ $X2=0.24 $Y2=2.39
r48 9 11 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.065 $Y=2.39
+ $X2=1.15 $Y2=2.475
r49 9 10 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.065 $Y=2.39 $X2=0.365
+ $Y2=2.39
r50 2 17 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=1.87
+ $Y=2.32 $X2=2.02 $Y2=2.465
r51 1 20 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.32 $X2=0.28 $Y2=2.47
.ends

.subckt PM_SKY130_FD_SC_LS__SDFBBN_2%VPWR 1 2 3 4 5 6 7 8 9 10 11 12 39 43 47 49
+ 53 57 61 65 69 73 77 83 87 89 94 95 97 98 100 101 102 104 109 117 122 131 150
+ 154 160 163 166 169 172 175 179 186 188 192
c210 47 0 1.36467e-19 $X=4.04 $Y=2.425
c211 43 0 3.52871e-20 $X=2.58 $Y=2.465
r212 191 192 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=18 $Y=3.33 $X2=18
+ $Y2=3.33
r213 188 189 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=17.04 $Y=3.33
+ $X2=17.04 $Y2=3.33
r214 185 186 9.96101 $w=5.68e-07 $l=1.65e-07 $layer=LI1_cond $X=15.005 $Y=3.13
+ $X2=15.17 $Y2=3.13
r215 183 185 0.167871 $w=5.68e-07 $l=8e-09 $layer=LI1_cond $X=14.997 $Y=3.13
+ $X2=15.005 $Y2=3.13
r216 181 183 7.49123 $w=5.68e-07 $l=3.57e-07 $layer=LI1_cond $X=14.64 $Y=3.13
+ $X2=14.997 $Y2=3.13
r217 181 182 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.64 $Y=3.33
+ $X2=14.64 $Y2=3.33
r218 178 181 4.09185 $w=5.68e-07 $l=1.95e-07 $layer=LI1_cond $X=14.445 $Y=3.13
+ $X2=14.64 $Y2=3.13
r219 178 179 9.96101 $w=5.68e-07 $l=1.65e-07 $layer=LI1_cond $X=14.445 $Y=3.13
+ $X2=14.28 $Y2=3.13
r220 175 176 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r221 172 173 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r222 169 170 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r223 167 170 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r224 166 167 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r225 163 164 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r226 160 161 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r227 158 192 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=17.52 $Y=3.33
+ $X2=18 $Y2=3.33
r228 158 189 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=17.52 $Y=3.33
+ $X2=17.04 $Y2=3.33
r229 157 158 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=17.52 $Y=3.33
+ $X2=17.52 $Y2=3.33
r230 155 188 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=17.225 $Y=3.33
+ $X2=17.06 $Y2=3.33
r231 155 157 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=17.225 $Y=3.33
+ $X2=17.52 $Y2=3.33
r232 154 191 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=17.875 $Y=3.33
+ $X2=18.057 $Y2=3.33
r233 154 157 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=17.875 $Y=3.33
+ $X2=17.52 $Y2=3.33
r234 153 189 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=16.56 $Y=3.33
+ $X2=17.04 $Y2=3.33
r235 152 153 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=16.56 $Y=3.33
+ $X2=16.56 $Y2=3.33
r236 150 188 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=16.895 $Y=3.33
+ $X2=17.06 $Y2=3.33
r237 150 152 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=16.895 $Y=3.33
+ $X2=16.56 $Y2=3.33
r238 149 153 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=15.6 $Y=3.33
+ $X2=16.56 $Y2=3.33
r239 149 182 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=15.6 $Y=3.33
+ $X2=14.64 $Y2=3.33
r240 148 186 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=15.6 $Y=3.33
+ $X2=15.17 $Y2=3.33
r241 148 149 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=15.6 $Y=3.33
+ $X2=15.6 $Y2=3.33
r242 145 182 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.16 $Y=3.33
+ $X2=14.64 $Y2=3.33
r243 144 179 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=14.16 $Y=3.33
+ $X2=14.28 $Y2=3.33
r244 144 145 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=14.16 $Y=3.33
+ $X2=14.16 $Y2=3.33
r245 142 145 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=14.16 $Y2=3.33
r246 141 144 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=12.72 $Y=3.33
+ $X2=14.16 $Y2=3.33
r247 141 142 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r248 138 142 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=12.72 $Y2=3.33
r249 138 176 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=11.28 $Y2=3.33
r250 137 138 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r251 135 175 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.56 $Y=3.33
+ $X2=11.395 $Y2=3.33
r252 135 137 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=11.56 $Y=3.33
+ $X2=12.24 $Y2=3.33
r253 134 176 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=11.28 $Y2=3.33
r254 133 134 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r255 131 175 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.23 $Y=3.33
+ $X2=11.395 $Y2=3.33
r256 131 133 90.6845 $w=1.68e-07 $l=1.39e-06 $layer=LI1_cond $X=11.23 $Y=3.33
+ $X2=9.84 $Y2=3.33
r257 130 134 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=9.84 $Y2=3.33
r258 129 130 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r259 127 172 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.695 $Y=3.33
+ $X2=8.53 $Y2=3.33
r260 127 129 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=8.695 $Y=3.33
+ $X2=9.36 $Y2=3.33
r261 126 173 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=8.4 $Y2=3.33
r262 126 170 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=5.04 $Y2=3.33
r263 125 126 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r264 123 169 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.215 $Y=3.33
+ $X2=5.09 $Y2=3.33
r265 123 125 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.215 $Y=3.33
+ $X2=5.52 $Y2=3.33
r266 122 172 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.365 $Y=3.33
+ $X2=8.53 $Y2=3.33
r267 122 125 185.61 $w=1.68e-07 $l=2.845e-06 $layer=LI1_cond $X=8.365 $Y=3.33
+ $X2=5.52 $Y2=3.33
r268 121 167 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r269 121 164 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=2.64 $Y2=3.33
r270 120 121 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r271 118 163 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.745 $Y=3.33
+ $X2=2.58 $Y2=3.33
r272 118 120 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=2.745 $Y=3.33
+ $X2=3.6 $Y2=3.33
r273 117 166 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.875 $Y=3.33
+ $X2=4.04 $Y2=3.33
r274 117 120 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3.875 $Y=3.33
+ $X2=3.6 $Y2=3.33
r275 116 164 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r276 115 116 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r277 113 116 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r278 113 161 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r279 112 115 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r280 112 113 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r281 110 160 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=0.73 $Y2=3.33
r282 110 112 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=1.2 $Y2=3.33
r283 109 163 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.415 $Y=3.33
+ $X2=2.58 $Y2=3.33
r284 109 115 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.415 $Y=3.33
+ $X2=2.16 $Y2=3.33
r285 107 161 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r286 106 107 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r287 104 160 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.73 $Y2=3.33
r288 104 106 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.24 $Y2=3.33
r289 102 130 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=9.12 $Y=3.33
+ $X2=9.36 $Y2=3.33
r290 102 173 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=9.12 $Y=3.33
+ $X2=8.4 $Y2=3.33
r291 100 148 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=15.825 $Y=3.33
+ $X2=15.6 $Y2=3.33
r292 100 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=15.825 $Y=3.33
+ $X2=15.99 $Y2=3.33
r293 99 152 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=16.155 $Y=3.33
+ $X2=16.56 $Y2=3.33
r294 99 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=16.155 $Y=3.33
+ $X2=15.99 $Y2=3.33
r295 97 137 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=12.305 $Y=3.33
+ $X2=12.24 $Y2=3.33
r296 97 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.305 $Y=3.33
+ $X2=12.47 $Y2=3.33
r297 96 141 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=12.635 $Y=3.33
+ $X2=12.72 $Y2=3.33
r298 96 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.635 $Y=3.33
+ $X2=12.47 $Y2=3.33
r299 94 129 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=9.465 $Y=3.33
+ $X2=9.36 $Y2=3.33
r300 94 95 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.465 $Y=3.33
+ $X2=9.63 $Y2=3.33
r301 93 133 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=9.795 $Y=3.33
+ $X2=9.84 $Y2=3.33
r302 93 95 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.795 $Y=3.33
+ $X2=9.63 $Y2=3.33
r303 89 92 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=18 $Y=1.985 $X2=18
+ $Y2=2.815
r304 87 191 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=18 $Y=3.245
+ $X2=18.057 $Y2=3.33
r305 87 92 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=18 $Y=3.245 $X2=18
+ $Y2=2.815
r306 83 86 26.1919 $w=3.28e-07 $l=7.5e-07 $layer=LI1_cond $X=17.06 $Y=2.045
+ $X2=17.06 $Y2=2.795
r307 81 188 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=17.06 $Y=3.245
+ $X2=17.06 $Y2=3.33
r308 81 86 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=17.06 $Y=3.245
+ $X2=17.06 $Y2=2.795
r309 77 80 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=15.99 $Y=2.115
+ $X2=15.99 $Y2=2.815
r310 75 101 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=15.99 $Y=3.245
+ $X2=15.99 $Y2=3.33
r311 75 80 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=15.99 $Y=3.245
+ $X2=15.99 $Y2=2.815
r312 71 183 3.68532 $w=3.45e-07 $l=2.85e-07 $layer=LI1_cond $X=14.997 $Y=2.845
+ $X2=14.997 $Y2=3.13
r313 71 73 23.2159 $w=3.43e-07 $l=6.95e-07 $layer=LI1_cond $X=14.997 $Y=2.845
+ $X2=14.997 $Y2=2.15
r314 67 98 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.47 $Y=3.245
+ $X2=12.47 $Y2=3.33
r315 67 69 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=12.47 $Y=3.245
+ $X2=12.47 $Y2=2.79
r316 63 175 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.395 $Y=3.245
+ $X2=11.395 $Y2=3.33
r317 63 65 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=11.395 $Y=3.245
+ $X2=11.395 $Y2=2.79
r318 59 95 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.63 $Y=3.245
+ $X2=9.63 $Y2=3.33
r319 59 61 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=9.63 $Y=3.245
+ $X2=9.63 $Y2=2.455
r320 55 172 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.53 $Y=3.245
+ $X2=8.53 $Y2=3.33
r321 55 57 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=8.53 $Y=3.245
+ $X2=8.53 $Y2=2.63
r322 51 169 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.09 $Y=3.245
+ $X2=5.09 $Y2=3.33
r323 51 53 31.8074 $w=2.48e-07 $l=6.9e-07 $layer=LI1_cond $X=5.09 $Y=3.245
+ $X2=5.09 $Y2=2.555
r324 50 166 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.205 $Y=3.33
+ $X2=4.04 $Y2=3.33
r325 49 169 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.965 $Y=3.33
+ $X2=5.09 $Y2=3.33
r326 49 50 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=4.965 $Y=3.33
+ $X2=4.205 $Y2=3.33
r327 45 166 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.04 $Y=3.245
+ $X2=4.04 $Y2=3.33
r328 45 47 28.6365 $w=3.28e-07 $l=8.2e-07 $layer=LI1_cond $X=4.04 $Y=3.245
+ $X2=4.04 $Y2=2.425
r329 41 163 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.58 $Y=3.245
+ $X2=2.58 $Y2=3.33
r330 41 43 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=2.58 $Y=3.245
+ $X2=2.58 $Y2=2.465
r331 37 160 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=3.33
r332 37 39 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=2.81
r333 12 92 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=17.81
+ $Y=1.84 $X2=17.96 $Y2=2.815
r334 12 89 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=17.81
+ $Y=1.84 $X2=17.96 $Y2=1.985
r335 11 86 400 $w=1.7e-07 $l=9.81071e-07 $layer=licon1_PDIFF $count=1 $X=16.835
+ $Y=1.92 $X2=17.06 $Y2=2.795
r336 11 83 400 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_PDIFF $count=1 $X=16.835
+ $Y=1.92 $X2=17.06 $Y2=2.045
r337 10 80 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=15.84
+ $Y=1.84 $X2=15.99 $Y2=2.815
r338 10 77 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=15.84
+ $Y=1.84 $X2=15.99 $Y2=2.115
r339 9 185 600 $w=1.7e-07 $l=1.35542e-06 $layer=licon1_PDIFF $count=1 $X=14.21
+ $Y=1.995 $X2=15.005 $Y2=3.01
r340 9 178 600 $w=1.7e-07 $l=1.12639e-06 $layer=licon1_PDIFF $count=1 $X=14.21
+ $Y=1.995 $X2=14.445 $Y2=3.01
r341 9 73 300 $w=1.7e-07 $l=8.69051e-07 $layer=licon1_PDIFF $count=2 $X=14.21
+ $Y=1.995 $X2=15.005 $Y2=2.15
r342 8 69 600 $w=1.7e-07 $l=9.24608e-07 $layer=licon1_PDIFF $count=1 $X=12.27
+ $Y=1.96 $X2=12.47 $Y2=2.79
r343 7 65 600 $w=1.7e-07 $l=3.16228e-07 $layer=licon1_PDIFF $count=1 $X=11.245
+ $Y=2.54 $X2=11.395 $Y2=2.79
r344 6 61 300 $w=1.7e-07 $l=4.00999e-07 $layer=licon1_PDIFF $count=2 $X=9.485
+ $Y=2.12 $X2=9.63 $Y2=2.455
r345 5 57 600 $w=1.7e-07 $l=5.80172e-07 $layer=licon1_PDIFF $count=1 $X=8.38
+ $Y=2.12 $X2=8.53 $Y2=2.63
r346 4 53 600 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=1 $X=4.905
+ $Y=2.32 $X2=5.05 $Y2=2.555
r347 3 47 300 $w=1.7e-07 $l=6.55725e-07 $layer=licon1_PDIFF $count=2 $X=3.89
+ $Y=1.84 $X2=4.04 $Y2=2.425
r348 2 43 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=2.435
+ $Y=2.32 $X2=2.58 $Y2=2.465
r349 1 39 600 $w=1.7e-07 $l=5.6e-07 $layer=licon1_PDIFF $count=1 $X=0.58 $Y=2.32
+ $X2=0.73 $Y2=2.81
.ends

.subckt PM_SKY130_FD_SC_LS__SDFBBN_2%A_197_119# 1 2 3 4 15 17 19 20 23 24 25 26
+ 28 29 32 33 34 36 37 38 40 41 42 44 45 46 48 49 50 51 56 57 58 60 61 63 64 68
c223 48 0 1.91291e-19 $X=6.03 $Y=0.84
c224 45 0 7.90252e-20 $X=5.945 $Y=0.925
c225 26 0 1.01507e-19 $X=1.69 $Y=1.205
c226 17 0 8.27414e-20 $X=1.57 $Y=2.515
c227 15 0 1.49963e-19 $X=1.53 $Y=2.425
r228 66 68 8.49906 $w=3.53e-07 $l=1.65e-07 $layer=LI1_cond $X=6.505 $Y=2.557
+ $X2=6.67 $Y2=2.557
r229 59 60 89.0535 $w=1.68e-07 $l=1.365e-06 $layer=LI1_cond $X=7.62 $Y=1.015
+ $X2=7.62 $Y2=2.38
r230 57 59 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.535 $Y=0.93
+ $X2=7.62 $Y2=1.015
r231 57 58 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=7.535 $Y=0.93
+ $X2=7.115 $Y2=0.93
r232 54 58 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.95 $Y=0.845
+ $X2=7.115 $Y2=0.93
r233 54 56 1.22229 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=6.95 $Y=0.845
+ $X2=6.95 $Y2=0.81
r234 53 56 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=6.95 $Y=0.435
+ $X2=6.95 $Y2=0.81
r235 51 60 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.535 $Y=2.465
+ $X2=7.62 $Y2=2.38
r236 51 68 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=7.535 $Y=2.465
+ $X2=6.67 $Y2=2.465
r237 49 53 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.785 $Y=0.35
+ $X2=6.95 $Y2=0.435
r238 49 50 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.785 $Y=0.35
+ $X2=6.115 $Y2=0.35
r239 47 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.03 $Y=0.435
+ $X2=6.115 $Y2=0.35
r240 47 48 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=6.03 $Y=0.435
+ $X2=6.03 $Y2=0.84
r241 45 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.945 $Y=0.925
+ $X2=6.03 $Y2=0.84
r242 45 46 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=5.945 $Y=0.925
+ $X2=5.28 $Y2=0.925
r243 44 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.195 $Y=0.84
+ $X2=5.28 $Y2=0.925
r244 43 44 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=5.195 $Y=0.425
+ $X2=5.195 $Y2=0.84
r245 41 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.11 $Y=0.34
+ $X2=5.195 $Y2=0.425
r246 41 42 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=5.11 $Y=0.34
+ $X2=4.52 $Y2=0.34
r247 39 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.435 $Y=0.425
+ $X2=4.52 $Y2=0.34
r248 39 40 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=4.435 $Y=0.425
+ $X2=4.435 $Y2=0.66
r249 37 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.35 $Y=0.745
+ $X2=4.435 $Y2=0.66
r250 37 38 53.1711 $w=1.68e-07 $l=8.15e-07 $layer=LI1_cond $X=4.35 $Y=0.745
+ $X2=3.535 $Y2=0.745
r251 36 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.45 $Y=0.66
+ $X2=3.535 $Y2=0.745
r252 35 36 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=3.45 $Y=0.425
+ $X2=3.45 $Y2=0.66
r253 33 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.365 $Y=0.34
+ $X2=3.45 $Y2=0.425
r254 33 34 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=3.365 $Y=0.34
+ $X2=2.77 $Y2=0.34
r255 31 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.685 $Y=0.425
+ $X2=2.77 $Y2=0.34
r256 31 32 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=2.685 $Y=0.425
+ $X2=2.685 $Y2=1.12
r257 30 64 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.155 $Y=1.205
+ $X2=2.07 $Y2=1.205
r258 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.6 $Y=1.205
+ $X2=2.685 $Y2=1.12
r259 29 30 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=2.6 $Y=1.205
+ $X2=2.155 $Y2=1.205
r260 27 64 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.07 $Y=1.29
+ $X2=2.07 $Y2=1.205
r261 27 28 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.07 $Y=1.29
+ $X2=2.07 $Y2=1.96
r262 25 64 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.985 $Y=1.205
+ $X2=2.07 $Y2=1.205
r263 25 26 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.985 $Y=1.205
+ $X2=1.69 $Y2=1.205
r264 23 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.985 $Y=2.045
+ $X2=2.07 $Y2=1.96
r265 23 24 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.985 $Y=2.045
+ $X2=1.655 $Y2=2.045
r266 21 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.57 $Y=2.13
+ $X2=1.655 $Y2=2.045
r267 21 61 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.57 $Y=2.13
+ $X2=1.57 $Y2=2.3
r268 20 26 6.89401 $w=1.7e-07 $l=1.39155e-07 $layer=LI1_cond $X=1.587 $Y=1.12
+ $X2=1.69 $Y2=1.205
r269 19 63 4.51862 $w=2.05e-07 $l=1.65e-07 $layer=LI1_cond $X=1.587 $Y=0.955
+ $X2=1.587 $Y2=0.79
r270 19 20 8.92683 $w=2.03e-07 $l=1.65e-07 $layer=LI1_cond $X=1.587 $Y=0.955
+ $X2=1.587 $Y2=1.12
r271 15 61 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=1.53 $Y=2.425
+ $X2=1.53 $Y2=2.3
r272 15 17 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=1.53 $Y=2.425
+ $X2=1.53 $Y2=2.515
r273 4 66 600 $w=1.7e-07 $l=2.81069e-07 $layer=licon1_PDIFF $count=1 $X=6.305
+ $Y=2.32 $X2=6.505 $Y2=2.515
r274 3 17 600 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=1.42
+ $Y=2.32 $X2=1.57 $Y2=2.515
r275 2 56 182 $w=1.7e-07 $l=2.8801e-07 $layer=licon1_NDIFF $count=1 $X=6.74
+ $Y=0.625 $X2=6.95 $Y2=0.81
r276 1 63 91 $w=1.7e-07 $l=6.3e-07 $layer=licon1_NDIFF $count=2 $X=0.985
+ $Y=0.595 $X2=1.525 $Y2=0.79
.ends

.subckt PM_SKY130_FD_SC_LS__SDFBBN_2%Q_N 1 2 9 15 19 20 23
r30 20 25 4.72801 $w=3.38e-07 $l=1.15e-07 $layer=LI1_cond $X=15.545 $Y=1.665
+ $X2=15.545 $Y2=1.78
r31 20 23 5.0075 $w=3.38e-07 $l=1.15e-07 $layer=LI1_cond $X=15.545 $Y=1.665
+ $X2=15.545 $Y2=1.55
r32 19 23 16.1832 $w=2.33e-07 $l=3.3e-07 $layer=LI1_cond $X=15.492 $Y=1.22
+ $X2=15.492 $Y2=1.55
r33 15 17 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=15.5 $Y=1.985
+ $X2=15.5 $Y2=2.815
r34 15 25 9.45003 $w=2.48e-07 $l=2.05e-07 $layer=LI1_cond $X=15.5 $Y=1.985
+ $X2=15.5 $Y2=1.78
r35 7 19 6.73378 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=15.445 $Y=1.055
+ $X2=15.445 $Y2=1.22
r36 7 9 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=15.445 $Y=1.055
+ $X2=15.445 $Y2=0.515
r37 2 17 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=15.39
+ $Y=1.84 $X2=15.54 $Y2=2.815
r38 2 15 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=15.39
+ $Y=1.84 $X2=15.54 $Y2=1.985
r39 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=15.305
+ $Y=0.37 $X2=15.445 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__SDFBBN_2%Q 1 2 9 13 14 20 26
c27 26 0 1.00299e-19 $X=17.55 $Y=1.82
r28 17 20 0.371756 $w=3.08e-07 $l=1e-08 $layer=LI1_cond $X=17.55 $Y=1.975
+ $X2=17.55 $Y2=1.985
r29 14 17 0.483283 $w=3.08e-07 $l=1.3e-08 $layer=LI1_cond $X=17.55 $Y=1.962
+ $X2=17.55 $Y2=1.975
r30 14 26 7.61225 $w=3.08e-07 $l=1.42e-07 $layer=LI1_cond $X=17.55 $Y=1.962
+ $X2=17.55 $Y2=1.82
r31 14 23 28.5508 $w=3.08e-07 $l=7.68e-07 $layer=LI1_cond $X=17.55 $Y=2.047
+ $X2=17.55 $Y2=2.815
r32 14 20 2.30489 $w=3.08e-07 $l=6.2e-08 $layer=LI1_cond $X=17.55 $Y=2.047
+ $X2=17.55 $Y2=1.985
r33 13 26 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=17.62 $Y=1.05
+ $X2=17.62 $Y2=1.82
r34 7 13 8.53494 $w=3.33e-07 $l=1.67e-07 $layer=LI1_cond $X=17.537 $Y=0.883
+ $X2=17.537 $Y2=1.05
r35 7 9 12.6597 $w=3.33e-07 $l=3.68e-07 $layer=LI1_cond $X=17.537 $Y=0.883
+ $X2=17.537 $Y2=0.515
r36 2 23 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=17.36
+ $Y=1.84 $X2=17.51 $Y2=2.815
r37 2 20 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=17.36
+ $Y=1.84 $X2=17.51 $Y2=1.985
r38 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=17.395
+ $Y=0.37 $X2=17.535 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__SDFBBN_2%VGND 1 2 3 4 5 6 7 8 9 10 31 33 37 41 45 49
+ 51 55 59 63 67 69 72 73 75 76 78 79 80 89 96 101 119 123 132 135 138 148 152
r191 151 152 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=18 $Y=0 $X2=18
+ $Y2=0
r192 148 149 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=17.04 $Y=0
+ $X2=17.04 $Y2=0
r193 139 143 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=11.76 $Y2=0
r194 138 139 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r195 135 136 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r196 132 133 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r197 129 130 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r198 127 152 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=17.52 $Y=0
+ $X2=18 $Y2=0
r199 127 149 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=17.52 $Y=0
+ $X2=17.04 $Y2=0
r200 126 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=17.52 $Y=0
+ $X2=17.52 $Y2=0
r201 124 148 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=17.2 $Y=0
+ $X2=17.035 $Y2=0
r202 124 126 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=17.2 $Y=0
+ $X2=17.52 $Y2=0
r203 123 151 4.01803 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=17.88 $Y=0
+ $X2=18.06 $Y2=0
r204 123 126 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=17.88 $Y=0
+ $X2=17.52 $Y2=0
r205 122 149 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=16.56 $Y=0
+ $X2=17.04 $Y2=0
r206 121 122 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=16.56 $Y=0
+ $X2=16.56 $Y2=0
r207 119 148 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=16.87 $Y=0
+ $X2=17.035 $Y2=0
r208 119 121 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=16.87 $Y=0
+ $X2=16.56 $Y2=0
r209 118 122 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=15.6 $Y=0
+ $X2=16.56 $Y2=0
r210 117 118 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=15.6 $Y=0
+ $X2=15.6 $Y2=0
r211 115 118 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=14.64 $Y=0
+ $X2=15.6 $Y2=0
r212 114 115 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=14.64 $Y=0
+ $X2=14.64 $Y2=0
r213 112 115 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=14.64 $Y2=0
r214 112 143 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=11.76 $Y2=0
r215 111 114 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=12.24 $Y=0
+ $X2=14.64 $Y2=0
r216 111 112 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r217 109 111 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=12.055 $Y=0
+ $X2=12.24 $Y2=0
r218 107 108 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r219 105 108 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=6 $Y=0 $X2=8.88
+ $Y2=0
r220 105 136 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.52
+ $Y2=0
r221 104 107 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=6 $Y=0 $X2=8.88
+ $Y2=0
r222 104 105 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=6 $Y=0 $X2=6
+ $Y2=0
r223 102 135 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.72 $Y=0
+ $X2=5.585 $Y2=0
r224 102 104 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=5.72 $Y=0 $X2=6
+ $Y2=0
r225 101 138 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.055 $Y=0
+ $X2=9.22 $Y2=0
r226 101 107 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=9.055 $Y=0
+ $X2=8.88 $Y2=0
r227 100 136 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=0
+ $X2=5.52 $Y2=0
r228 100 133 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0
+ $X2=4.08 $Y2=0
r229 99 100 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r230 97 132 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.18 $Y=0
+ $X2=4.055 $Y2=0
r231 97 99 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=4.18 $Y=0 $X2=4.56
+ $Y2=0
r232 96 135 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.45 $Y=0
+ $X2=5.585 $Y2=0
r233 96 99 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=5.45 $Y=0 $X2=4.56
+ $Y2=0
r234 95 133 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r235 94 95 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r236 92 95 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r237 91 94 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r238 91 92 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r239 89 132 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.93 $Y=0
+ $X2=4.055 $Y2=0
r240 89 94 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=3.93 $Y=0 $X2=3.6
+ $Y2=0
r241 88 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r242 87 88 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r243 85 88 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=0.72 $Y=0
+ $X2=2.16 $Y2=0
r244 85 130 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0
+ $X2=0.24 $Y2=0
r245 84 87 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.72 $Y=0 $X2=2.16
+ $Y2=0
r246 84 85 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r247 82 129 4.67962 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=0.47 $Y=0
+ $X2=0.235 $Y2=0
r248 82 84 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.47 $Y=0 $X2=0.72
+ $Y2=0
r249 80 139 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=9.12 $Y=0
+ $X2=9.36 $Y2=0
r250 80 108 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=9.12 $Y=0
+ $X2=8.88 $Y2=0
r251 78 117 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=15.78 $Y=0
+ $X2=15.6 $Y2=0
r252 78 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=15.78 $Y=0
+ $X2=15.945 $Y2=0
r253 77 121 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=16.11 $Y=0
+ $X2=16.56 $Y2=0
r254 77 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=16.11 $Y=0
+ $X2=15.945 $Y2=0
r255 75 114 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=14.825 $Y=0
+ $X2=14.64 $Y2=0
r256 75 76 7.75133 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=14.825 $Y=0
+ $X2=14.967 $Y2=0
r257 74 117 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=15.11 $Y=0
+ $X2=15.6 $Y2=0
r258 74 76 7.75133 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=15.11 $Y=0
+ $X2=14.967 $Y2=0
r259 72 87 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=2.18 $Y=0 $X2=2.16
+ $Y2=0
r260 72 73 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.18 $Y=0 $X2=2.305
+ $Y2=0
r261 71 91 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=2.43 $Y=0 $X2=2.64
+ $Y2=0
r262 71 73 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.43 $Y=0 $X2=2.305
+ $Y2=0
r263 67 151 3.12513 $w=2.5e-07 $l=1.09087e-07 $layer=LI1_cond $X=18.005 $Y=0.085
+ $X2=18.06 $Y2=0
r264 67 69 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=18.005 $Y=0.085
+ $X2=18.005 $Y2=0.515
r265 63 65 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=17.035 $Y=0.515
+ $X2=17.035 $Y2=0.885
r266 61 148 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=17.035 $Y=0.085
+ $X2=17.035 $Y2=0
r267 61 63 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=17.035 $Y=0.085
+ $X2=17.035 $Y2=0.515
r268 57 79 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=15.945 $Y=0.085
+ $X2=15.945 $Y2=0
r269 57 59 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=15.945 $Y=0.085
+ $X2=15.945 $Y2=0.515
r270 53 76 0.432977 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=14.967 $Y=0.085
+ $X2=14.967 $Y2=0
r271 53 55 17.3877 $w=2.83e-07 $l=4.3e-07 $layer=LI1_cond $X=14.967 $Y=0.085
+ $X2=14.967 $Y2=0.515
r272 52 138 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.385 $Y=0
+ $X2=9.22 $Y2=0
r273 51 145 10.6025 $w=3.73e-07 $l=3.45e-07 $layer=LI1_cond $X=11.867 $Y=0
+ $X2=11.867 $Y2=0.345
r274 51 109 5.38787 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=11.867 $Y=0
+ $X2=12.055 $Y2=0
r275 51 143 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r276 51 52 149.727 $w=1.68e-07 $l=2.295e-06 $layer=LI1_cond $X=11.68 $Y=0
+ $X2=9.385 $Y2=0
r277 47 138 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.22 $Y=0.085
+ $X2=9.22 $Y2=0
r278 47 49 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=9.22 $Y=0.085
+ $X2=9.22 $Y2=0.77
r279 43 135 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.585 $Y=0.085
+ $X2=5.585 $Y2=0
r280 43 45 17.9269 $w=2.68e-07 $l=4.2e-07 $layer=LI1_cond $X=5.585 $Y=0.085
+ $X2=5.585 $Y2=0.505
r281 39 132 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.055 $Y=0.085
+ $X2=4.055 $Y2=0
r282 39 41 11.0635 $w=2.48e-07 $l=2.4e-07 $layer=LI1_cond $X=4.055 $Y=0.085
+ $X2=4.055 $Y2=0.325
r283 35 73 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.305 $Y=0.085
+ $X2=2.305 $Y2=0
r284 35 37 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=2.305 $Y=0.085
+ $X2=2.305 $Y2=0.76
r285 31 129 3.08656 $w=3.3e-07 $l=1.14782e-07 $layer=LI1_cond $X=0.305 $Y=0.085
+ $X2=0.235 $Y2=0
r286 31 33 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.305 $Y=0.085
+ $X2=0.305 $Y2=0.765
r287 10 69 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=17.825
+ $Y=0.37 $X2=17.965 $Y2=0.515
r288 9 65 182 $w=1.7e-07 $l=5.21368e-07 $layer=licon1_NDIFF $count=1 $X=16.795
+ $Y=0.47 $X2=17.035 $Y2=0.885
r289 9 63 182 $w=1.7e-07 $l=2.61534e-07 $layer=licon1_NDIFF $count=1 $X=16.795
+ $Y=0.47 $X2=17.035 $Y2=0.515
r290 8 59 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=15.735
+ $Y=0.37 $X2=15.875 $Y2=0.515
r291 7 55 91 $w=1.7e-07 $l=9.12414e-07 $layer=licon1_NDIFF $count=2 $X=14.275
+ $Y=0.9 $X2=15.015 $Y2=0.515
r292 6 145 182 $w=1.7e-07 $l=2.70555e-07 $layer=licon1_NDIFF $count=1 $X=11.625
+ $Y=0.41 $X2=11.865 $Y2=0.345
r293 5 49 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=9.01
+ $Y=0.625 $X2=9.22 $Y2=0.77
r294 4 45 182 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=1 $X=5.39
+ $Y=0.36 $X2=5.545 $Y2=0.505
r295 3 41 182 $w=1.7e-07 $l=2.91033e-07 $layer=licon1_NDIFF $count=1 $X=3.875
+ $Y=0.49 $X2=4.095 $Y2=0.325
r296 2 37 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=2.205
+ $Y=0.595 $X2=2.345 $Y2=0.76
r297 1 33 182 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_NDIFF $count=1 $X=0.16
+ $Y=0.595 $X2=0.305 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LS__SDFBBN_2%A_1473_73# 1 2 7 10 11 19
c40 19 0 8.54043e-20 $X=8.665 $Y=0.77
r41 16 19 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=8.535 $Y=0.77
+ $X2=8.665 $Y2=0.77
r42 11 14 4.33861 $w=4.23e-07 $l=1.6e-07 $layer=LI1_cond $X=7.557 $Y=0.35
+ $X2=7.557 $Y2=0.51
r43 10 16 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.535 $Y=0.605
+ $X2=8.535 $Y2=0.77
r44 9 10 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=8.535 $Y=0.435
+ $X2=8.535 $Y2=0.605
r45 8 11 6.14847 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=7.77 $Y=0.35
+ $X2=7.557 $Y2=0.35
r46 7 9 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.45 $Y=0.35
+ $X2=8.535 $Y2=0.435
r47 7 8 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=8.45 $Y=0.35 $X2=7.77
+ $Y2=0.35
r48 2 19 182 $w=1.7e-07 $l=3.245e-07 $layer=licon1_NDIFF $count=1 $X=8.405
+ $Y=0.625 $X2=8.665 $Y2=0.77
r49 1 14 182 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_NDIFF $count=1 $X=7.365
+ $Y=0.365 $X2=7.555 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_LS__SDFBBN_2%A_2452_74# 1 2 9 15 16
c24 16 0 6.88126e-20 $X=13.265 $Y=0.375
r25 15 16 8.91885 $w=2.38e-07 $l=1.65e-07 $layer=LI1_cond $X=13.43 $Y=0.375
+ $X2=13.265 $Y2=0.375
r26 9 12 4.80185 $w=4.18e-07 $l=1.75e-07 $layer=LI1_cond $X=12.445 $Y=0.34
+ $X2=12.445 $Y2=0.515
r27 8 9 6.07598 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=12.655 $Y=0.34
+ $X2=12.445 $Y2=0.34
r28 8 16 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=12.655 $Y=0.34
+ $X2=13.265 $Y2=0.34
r29 2 15 182 $w=1.7e-07 $l=2.39165e-07 $layer=licon1_NDIFF $count=1 $X=13.21
+ $Y=0.37 $X2=13.43 $Y2=0.41
r30 1 12 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=12.26
+ $Y=0.37 $X2=12.445 $Y2=0.515
.ends

