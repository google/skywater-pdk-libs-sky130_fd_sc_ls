* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__nand4bb_2 A_N B_N C D VGND VNB VPB VPWR Y
X0 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X1 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X2 VPWR B_N a_231_74# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X4 a_886_74# C a_678_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X5 a_373_74# a_27_368# Y VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X6 Y a_27_368# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X7 VPWR a_231_74# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X8 VGND D a_886_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X9 a_27_368# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_678_74# C a_886_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X11 Y a_27_368# a_373_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X12 a_373_74# a_231_74# a_678_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X13 a_678_74# a_231_74# a_373_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X14 a_886_74# D VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X15 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X16 Y a_231_74# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X17 VGND B_N a_231_74# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X18 a_27_368# A_N VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X19 VPWR a_27_368# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
.ends
