* File: sky130_fd_sc_ls__dlrbn_2.spice
* Created: Fri Aug 28 13:18:03 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__dlrbn_2.pex.spice"
.subckt sky130_fd_sc_ls__dlrbn_2  VNB VPB D GATE_N RESET_B VPWR Q Q_N VGND
* 
* VGND	VGND
* Q_N	Q_N
* Q	Q
* VPWR	VPWR
* RESET_B	RESET_B
* GATE_N	GATE_N
* D	D
* VPB	VPB
* VNB	VNB
MM1009 N_VGND_M1009_d N_D_M1009_g N_A_27_112#_M1009_s VNB NSHORT L=0.15 W=0.55
+ AD=0.129591 AS=0.15675 PD=0.997674 PS=1.67 NRD=17.988 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75000.8 A=0.0825 P=1.4 MULT=1
MM1007 N_A_230_74#_M1007_d N_GATE_N_M1007_g N_VGND_M1009_d VNB NSHORT L=0.15
+ W=0.74 AD=0.2109 AS=0.174359 PD=2.05 PS=1.34233 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75000.7 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1019 N_VGND_M1019_d N_A_230_74#_M1019_g N_A_363_74#_M1019_s VNB NSHORT L=0.15
+ W=0.74 AD=0.205591 AS=0.2109 PD=1.3942 PS=2.05 NRD=28.368 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001.7 A=0.111 P=1.78 MULT=1
MM1002 A_592_74# N_A_27_112#_M1002_g N_VGND_M1019_d VNB NSHORT L=0.15 W=0.64
+ AD=0.0768 AS=0.177809 PD=0.88 PS=1.2058 NRD=12.18 NRS=19.68 M=1 R=4.26667
+ SA=75000.9 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1001 N_A_670_74#_M1001_d N_A_230_74#_M1001_g A_592_74# VNB NSHORT L=0.15
+ W=0.64 AD=0.147321 AS=0.0768 PD=1.31623 PS=0.88 NRD=15.936 NRS=12.18 M=1
+ R=4.26667 SA=75001.3 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1010 A_790_74# N_A_363_74#_M1010_g N_A_670_74#_M1001_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.0966792 PD=0.66 PS=0.863774 NRD=18.564 NRS=24.276 M=1
+ R=2.8 SA=75001.9 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1020 N_VGND_M1020_d N_A_838_48#_M1020_g A_790_74# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75002.3
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1025 A_1066_74# N_A_670_74#_M1025_g N_A_838_48#_M1025_s VNB NSHORT L=0.15
+ W=0.74 AD=0.0888 AS=0.2109 PD=0.98 PS=2.05 NRD=10.536 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75002 A=0.111 P=1.78 MULT=1
MM1026 N_VGND_M1026_d N_RESET_B_M1026_g A_1066_74# VNB NSHORT L=0.15 W=0.74
+ AD=0.1628 AS=0.0888 PD=1.18 PS=0.98 NRD=0 NRS=10.536 M=1 R=4.93333 SA=75000.6
+ SB=75001.7 A=0.111 P=1.78 MULT=1
MM1012 N_VGND_M1026_d N_A_838_48#_M1012_g N_Q_M1012_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1628 AS=0.1036 PD=1.18 PS=1.02 NRD=25.944 NRS=0 M=1 R=4.93333 SA=75001.2
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1027 N_VGND_M1027_d N_A_838_48#_M1027_g N_Q_M1012_s VNB NSHORT L=0.15 W=0.74
+ AD=0.133522 AS=0.1036 PD=1.16899 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.6
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1011 N_A_1446_368#_M1011_d N_A_838_48#_M1011_g N_VGND_M1027_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.1824 AS=0.115478 PD=1.85 PS=1.01101 NRD=0 NRS=13.116 M=1
+ R=4.26667 SA=75002.1 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1014 N_VGND_M1014_d N_A_1446_368#_M1014_g N_Q_N_M1014_s VNB NSHORT L=0.15
+ W=0.74 AD=0.2109 AS=0.1184 PD=2.05 PS=1.06 NRD=0 NRS=3.24 M=1 R=4.93333
+ SA=75000.2 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1024 N_VGND_M1024_d N_A_1446_368#_M1024_g N_Q_N_M1014_s VNB NSHORT L=0.15
+ W=0.74 AD=0.2109 AS=0.1184 PD=2.05 PS=1.06 NRD=0 NRS=3.24 M=1 R=4.93333
+ SA=75000.7 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1013 N_VPWR_M1013_d N_D_M1013_g N_A_27_112#_M1013_s VPB PHIGHVT L=0.15 W=0.84
+ AD=0.2226 AS=0.2478 PD=1.37 PS=2.27 NRD=2.3443 NRS=2.3443 M=1 R=5.6 SA=75000.2
+ SB=75000.9 A=0.126 P=1.98 MULT=1
MM1006 N_A_230_74#_M1006_d N_GATE_N_M1006_g N_VPWR_M1013_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.2478 AS=0.2226 PD=2.27 PS=1.37 NRD=2.3443 NRS=56.2829 M=1 R=5.6
+ SA=75000.9 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1022 N_VPWR_M1022_d N_A_230_74#_M1022_g N_A_363_74#_M1022_s VPB PHIGHVT L=0.15
+ W=0.84 AD=0.230498 AS=0.383 PD=1.49739 PS=2.88 NRD=51.4367 NRS=23.443 M=1
+ R=5.6 SA=75000.3 SB=75002.4 A=0.126 P=1.98 MULT=1
MM1016 A_595_392# N_A_27_112#_M1016_g N_VPWR_M1022_d VPB PHIGHVT L=0.15 W=1
+ AD=0.12 AS=0.274402 PD=1.24 PS=1.78261 NRD=12.7853 NRS=19.6803 M=1 R=6.66667
+ SA=75000.8 SB=75002.2 A=0.15 P=2.3 MULT=1
MM1003 N_A_670_74#_M1003_d N_A_363_74#_M1003_g A_595_392# VPB PHIGHVT L=0.15 W=1
+ AD=0.24493 AS=0.12 PD=1.97183 PS=1.24 NRD=2.9353 NRS=12.7853 M=1 R=6.66667
+ SA=75001.2 SB=75001.8 A=0.15 P=2.3 MULT=1
MM1000 A_783_508# N_A_230_74#_M1000_g N_A_670_74#_M1003_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.09975 AS=0.10287 PD=0.895 PS=0.828169 NRD=85.5965 NRS=51.5943 M=1
+ R=2.8 SA=75001.6 SB=75003.4 A=0.063 P=1.14 MULT=1
MM1021 N_VPWR_M1021_d N_A_838_48#_M1021_g A_783_508# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.122182 AS=0.09975 PD=0.951818 PS=0.895 NRD=70.3487 NRS=85.5965 M=1 R=2.8
+ SA=75002.3 SB=75002.8 A=0.063 P=1.14 MULT=1
MM1015 N_A_838_48#_M1015_d N_A_670_74#_M1015_g N_VPWR_M1021_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.1736 AS=0.325818 PD=1.43 PS=2.53818 NRD=3.5066 NRS=34.2977 M=1
+ R=7.46667 SA=75001.3 SB=75002.1 A=0.168 P=2.54 MULT=1
MM1017 N_VPWR_M1017_d N_RESET_B_M1017_g N_A_838_48#_M1015_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.196 AS=0.1736 PD=1.47 PS=1.43 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75001.7 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1004 N_VPWR_M1017_d N_A_838_48#_M1004_g N_Q_M1004_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.196 AS=0.168 PD=1.47 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.2 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1023 N_VPWR_M1023_d N_A_838_48#_M1023_g N_Q_M1004_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.204347 AS=0.168 PD=1.55849 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.7 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1005 N_A_1446_368#_M1005_d N_A_838_48#_M1005_g N_VPWR_M1023_d VPB PHIGHVT
+ L=0.15 W=1 AD=0.295 AS=0.182453 PD=2.59 PS=1.39151 NRD=1.9503 NRS=12.7853 M=1
+ R=6.66667 SA=75003 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1008 N_Q_N_M1008_d N_A_1446_368#_M1008_g N_VPWR_M1008_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1018 N_Q_N_M1008_d N_A_1446_368#_M1018_g N_VPWR_M1018_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75000.2 A=0.168 P=2.54 MULT=1
DX28_noxref VNB VPB NWDIODE A=17.754 P=22.92
c_93 VNB 0 1.25688e-19 $X=0 $Y=0
c_1106 A_595_392# 0 1.09527e-19 $X=2.975 $Y=1.96
*
.include "sky130_fd_sc_ls__dlrbn_2.pxi.spice"
*
.ends
*
*
