* File: sky130_fd_sc_ls__dfrtp_2.pex.spice
* Created: Fri Aug 28 13:14:39 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__DFRTP_2%D 2 4 5 7 10 12 13 14 19 20 23
r35 23 25 40.9207 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=0.402 $Y=1.845
+ $X2=0.402 $Y2=2.01
r36 23 24 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.845 $X2=0.385 $Y2=1.845
r37 19 21 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=0.402 $Y=1.165
+ $X2=0.402 $Y2=1
r38 19 20 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.165 $X2=0.385 $Y2=1.165
r39 14 24 5.91795 $w=3.68e-07 $l=1.9e-07 $layer=LI1_cond $X=0.31 $Y=2.035
+ $X2=0.31 $Y2=1.845
r40 13 24 5.60648 $w=3.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.31 $Y=1.665
+ $X2=0.31 $Y2=1.845
r41 12 13 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.31 $Y=1.295
+ $X2=0.31 $Y2=1.665
r42 12 20 4.04912 $w=3.68e-07 $l=1.3e-07 $layer=LI1_cond $X=0.31 $Y=1.295
+ $X2=0.31 $Y2=1.165
r43 10 21 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=0.51 $Y=0.6 $X2=0.51
+ $Y2=1
r44 5 7 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.495 $Y=2.465
+ $X2=0.495 $Y2=2.75
r45 4 5 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.495 $Y=2.375 $X2=0.495
+ $Y2=2.465
r46 4 25 141.879 $w=1.8e-07 $l=3.65e-07 $layer=POLY_cond $X=0.495 $Y=2.375
+ $X2=0.495 $Y2=2.01
r47 2 23 2.68759 $w=3.65e-07 $l=1.7e-08 $layer=POLY_cond $X=0.402 $Y=1.828
+ $X2=0.402 $Y2=1.845
r48 1 19 2.68759 $w=3.65e-07 $l=1.7e-08 $layer=POLY_cond $X=0.402 $Y=1.182
+ $X2=0.402 $Y2=1.165
r49 1 2 102.129 $w=3.65e-07 $l=6.46e-07 $layer=POLY_cond $X=0.402 $Y=1.182
+ $X2=0.402 $Y2=1.828
.ends

.subckt PM_SKY130_FD_SC_LS__DFRTP_2%CLK 1 3 5 7 8
c45 8 0 1.55106e-19 $X=2.16 $Y=1.665
c46 5 0 2.84391e-19 $X=1.985 $Y=1.435
c47 3 0 1.62267e-19 $X=1.905 $Y=2.45
r48 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.96
+ $Y=1.61 $X2=1.96 $Y2=1.61
r49 8 12 5.6351 $w=4.33e-07 $l=2e-07 $layer=LI1_cond $X=2.16 $Y=1.55 $X2=1.96
+ $Y2=1.55
r50 5 11 40.1136 $w=3.43e-07 $l=1.90788e-07 $layer=POLY_cond $X=1.985 $Y=1.435
+ $X2=1.952 $Y2=1.61
r51 5 7 151.027 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=1.985 $Y=1.435
+ $X2=1.985 $Y2=0.965
r52 1 11 38.7084 $w=3.43e-07 $l=1.87029e-07 $layer=POLY_cond $X=1.905 $Y=1.775
+ $X2=1.952 $Y2=1.61
r53 1 3 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=1.905 $Y=1.775
+ $X2=1.905 $Y2=2.45
.ends

.subckt PM_SKY130_FD_SC_LS__DFRTP_2%A_495_390# 1 2 7 9 11 13 15 17 19 20 21 22
+ 24 27 28 30 33 34 35 38 39 42 45 49 54 60 63
c193 49 0 9.01765e-20 $X=2.832 $Y=0.415
c194 45 0 1.55106e-19 $X=2.967 $Y=1.95
c195 38 0 1.33493e-19 $X=7.12 $Y=2.14
c196 28 0 8.54071e-20 $X=4.305 $Y=0.415
c197 21 0 4.38853e-20 $X=6.355 $Y=1.27
c198 15 0 3.65694e-19 $X=4.04 $Y=0.9
c199 7 0 6.12976e-20 $X=3.41 $Y=1.99
r200 62 63 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=7.12 $Y=1.18
+ $X2=7.37 $Y2=1.18
r201 60 69 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=6.88 $Y=1.18 $X2=6.88
+ $Y2=1.27
r202 59 62 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=6.88 $Y=1.18
+ $X2=7.12 $Y2=1.18
r203 59 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.88
+ $Y=1.18 $X2=6.88 $Y2=1.18
r204 54 56 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=4.39 $Y=0.415
+ $X2=4.39 $Y2=0.7
r205 52 53 6.07947 $w=4.73e-07 $l=8.5e-08 $layer=LI1_cond $X=2.832 $Y=0.72
+ $X2=2.832 $Y2=0.805
r206 49 52 7.68008 $w=4.73e-07 $l=3.05e-07 $layer=LI1_cond $X=2.832 $Y=0.415
+ $X2=2.832 $Y2=0.72
r207 48 65 13.3477 $w=3.25e-07 $l=9e-08 $layer=POLY_cond $X=3.34 $Y=1.82
+ $X2=3.34 $Y2=1.73
r208 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.34
+ $Y=1.82 $X2=3.34 $Y2=1.82
r209 45 47 12.2 $w=3.73e-07 $l=3.73e-07 $layer=LI1_cond $X=2.967 $Y=1.95
+ $X2=3.34 $Y2=1.95
r210 44 45 11.5131 $w=3.73e-07 $l=3.52e-07 $layer=LI1_cond $X=2.615 $Y=1.95
+ $X2=2.967 $Y2=1.95
r211 42 63 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.37 $Y=1.015
+ $X2=7.37 $Y2=1.18
r212 41 42 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=7.37 $Y=0.425
+ $X2=7.37 $Y2=1.015
r213 39 72 25.8214 $w=3.64e-07 $l=1.95e-07 $layer=POLY_cond $X=7.12 $Y=2.182
+ $X2=7.315 $Y2=2.182
r214 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.12
+ $Y=2.14 $X2=7.12 $Y2=2.14
r215 36 62 0.716491 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=7.12 $Y=1.345
+ $X2=7.12 $Y2=1.18
r216 36 38 27.7634 $w=3.28e-07 $l=7.95e-07 $layer=LI1_cond $X=7.12 $Y=1.345
+ $X2=7.12 $Y2=2.14
r217 34 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.285 $Y=0.34
+ $X2=7.37 $Y2=0.425
r218 34 35 104.385 $w=1.68e-07 $l=1.6e-06 $layer=LI1_cond $X=7.285 $Y=0.34
+ $X2=5.685 $Y2=0.34
r219 32 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.6 $Y=0.425
+ $X2=5.685 $Y2=0.34
r220 32 33 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=5.6 $Y=0.425
+ $X2=5.6 $Y2=0.615
r221 31 56 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.475 $Y=0.7
+ $X2=4.39 $Y2=0.7
r222 30 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.515 $Y=0.7
+ $X2=5.6 $Y2=0.615
r223 30 31 67.8503 $w=1.68e-07 $l=1.04e-06 $layer=LI1_cond $X=5.515 $Y=0.7
+ $X2=4.475 $Y2=0.7
r224 29 49 6.83586 $w=1.7e-07 $l=2.38e-07 $layer=LI1_cond $X=3.07 $Y=0.415
+ $X2=2.832 $Y2=0.415
r225 28 54 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.305 $Y=0.415
+ $X2=4.39 $Y2=0.415
r226 28 29 80.5722 $w=1.68e-07 $l=1.235e-06 $layer=LI1_cond $X=4.305 $Y=0.415
+ $X2=3.07 $Y2=0.415
r227 27 45 4.25738 $w=2.05e-07 $l=3.25e-07 $layer=LI1_cond $X=2.967 $Y=1.625
+ $X2=2.967 $Y2=1.95
r228 27 53 44.3636 $w=2.03e-07 $l=8.2e-07 $layer=LI1_cond $X=2.967 $Y=1.625
+ $X2=2.967 $Y2=0.805
r229 22 72 23.572 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=7.315 $Y=2.39
+ $X2=7.315 $Y2=2.182
r230 22 24 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.315 $Y=2.39
+ $X2=7.315 $Y2=2.675
r231 20 69 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.715 $Y=1.27
+ $X2=6.88 $Y2=1.27
r232 20 21 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=6.715 $Y=1.27
+ $X2=6.355 $Y2=1.27
r233 17 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.28 $Y=1.195
+ $X2=6.355 $Y2=1.27
r234 17 19 146.207 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=6.28 $Y=1.195
+ $X2=6.28 $Y2=0.74
r235 13 25 80.845 $w=2.02e-07 $l=3.58295e-07 $layer=POLY_cond $X=4.04 $Y=1.405
+ $X2=3.97 $Y2=1.73
r236 13 15 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=4.04 $Y=1.405
+ $X2=4.04 $Y2=0.9
r237 12 65 20.86 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.505 $Y=1.73
+ $X2=3.34 $Y2=1.73
r238 11 25 9.80621 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=3.825 $Y=1.73
+ $X2=3.97 $Y2=1.73
r239 11 12 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.825 $Y=1.73
+ $X2=3.505 $Y2=1.73
r240 7 48 39.3126 $w=3.25e-07 $l=2.0199e-07 $layer=POLY_cond $X=3.41 $Y=1.99
+ $X2=3.34 $Y2=1.82
r241 7 9 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=3.41 $Y=1.99 $X2=3.41
+ $Y2=2.525
r242 2 44 600 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_PDIFF $count=1 $X=2.475
+ $Y=1.95 $X2=2.615 $Y2=2.11
r243 1 52 182 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_NDIFF $count=1 $X=2.61
+ $Y=0.595 $X2=2.76 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_LS__DFRTP_2%A_839_359# 1 2 7 9 12 16 19 20 23 29 31 32
c87 20 0 1.69473e-19 $X=4.445 $Y=1.04
c88 16 0 3.76464e-20 $X=4.36 $Y=1.96
c89 12 0 1.99579e-19 $X=4.43 $Y=0.9
c90 7 0 1.18794e-19 $X=4.275 $Y=2.21
r91 29 32 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=6.18 $Y=2.02
+ $X2=6.18 $Y2=1.855
r92 25 31 3.70735 $w=2.5e-07 $l=1.21589e-07 $layer=LI1_cond $X=6.1 $Y=1.13
+ $X2=6.02 $Y2=1.042
r93 25 32 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=6.1 $Y=1.13 $X2=6.1
+ $Y2=1.855
r94 21 31 3.70735 $w=2.5e-07 $l=8.7e-08 $layer=LI1_cond $X=6.02 $Y=0.955
+ $X2=6.02 $Y2=1.042
r95 21 23 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=6.02 $Y=0.955
+ $X2=6.02 $Y2=0.86
r96 19 31 2.76166 $w=1.7e-07 $l=1.65997e-07 $layer=LI1_cond $X=5.855 $Y=1.04
+ $X2=6.02 $Y2=1.042
r97 19 20 91.9893 $w=1.68e-07 $l=1.41e-06 $layer=LI1_cond $X=5.855 $Y=1.04
+ $X2=4.445 $Y2=1.04
r98 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.36
+ $Y=1.96 $X2=4.36 $Y2=1.96
r99 14 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.36 $Y=1.125
+ $X2=4.445 $Y2=1.04
r100 14 16 54.4759 $w=1.68e-07 $l=8.35e-07 $layer=LI1_cond $X=4.36 $Y=1.125
+ $X2=4.36 $Y2=1.96
r101 10 17 38.5495 $w=3.2e-07 $l=1.90526e-07 $layer=POLY_cond $X=4.43 $Y=1.795
+ $X2=4.375 $Y2=1.96
r102 10 12 458.926 $w=1.5e-07 $l=8.95e-07 $layer=POLY_cond $X=4.43 $Y=1.795
+ $X2=4.43 $Y2=0.9
r103 7 17 51.3527 $w=3.2e-07 $l=2.95804e-07 $layer=POLY_cond $X=4.275 $Y=2.21
+ $X2=4.375 $Y2=1.96
r104 7 9 101.22 $w=1.5e-07 $l=3.15e-07 $layer=POLY_cond $X=4.275 $Y=2.21
+ $X2=4.275 $Y2=2.525
r105 2 29 300 $w=1.7e-07 $l=3.71786e-07 $layer=licon1_PDIFF $count=2 $X=5.98
+ $Y=1.735 $X2=6.18 $Y2=2.02
r106 1 23 182 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_NDIFF $count=1 $X=5.88
+ $Y=0.37 $X2=6.02 $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_LS__DFRTP_2%RESET_B 4 6 8 11 12 13 17 19 20 22 23 25 28
+ 30 33 35 36 37 38 41 43 46 49 50 53 61
c210 50 0 1.62267e-19 $X=1.12 $Y=1.305
c211 49 0 1.26266e-19 $X=1.12 $Y=1.305
c212 43 0 3.83476e-20 $X=7.92 $Y=2.035
c213 37 0 4.38853e-20 $X=7.775 $Y=2.035
c214 33 0 3.76464e-20 $X=4.88 $Y=1.26
c215 12 0 7.77791e-20 $X=4.715 $Y=0.18
c216 8 0 1.67618e-19 $X=0.962 $Y=2.358
r217 60 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.23
+ $Y=2.11 $X2=8.23 $Y2=2.11
r218 53 55 36.1309 $w=5.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.09 $Y=1.985
+ $X2=1.09 $Y2=2.15
r219 53 54 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.12
+ $Y=1.985 $X2=1.12 $Y2=1.985
r220 50 54 27.9879 $w=2.78e-07 $l=6.8e-07 $layer=LI1_cond $X=1.145 $Y=1.305
+ $X2=1.145 $Y2=1.985
r221 49 51 47.4091 $w=5.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.09 $Y=1.305
+ $X2=1.09 $Y2=1.14
r222 49 50 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.12
+ $Y=1.305 $X2=1.12 $Y2=1.305
r223 46 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=2.035
+ $X2=1.2 $Y2=2.035
r224 44 61 10.0636 $w=3.53e-07 $l=3.1e-07 $layer=LI1_cond $X=7.92 $Y=2.097
+ $X2=8.23 $Y2=2.097
r225 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=2.035
+ $X2=7.92 $Y2=2.035
r226 41 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.12
+ $Y=1.96 $X2=5.12 $Y2=1.96
r227 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=2.035
+ $X2=5.04 $Y2=2.035
r228 38 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.185 $Y=2.035
+ $X2=5.04 $Y2=2.035
r229 37 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.775 $Y=2.035
+ $X2=7.92 $Y2=2.035
r230 37 38 3.20544 $w=1.4e-07 $l=2.59e-06 $layer=MET1_cond $X=7.775 $Y=2.035
+ $X2=5.185 $Y2=2.035
r231 36 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.345 $Y=2.035
+ $X2=1.2 $Y2=2.035
r232 35 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.895 $Y=2.035
+ $X2=5.04 $Y2=2.035
r233 35 36 4.39356 $w=1.4e-07 $l=3.55e-06 $layer=MET1_cond $X=4.895 $Y=2.035
+ $X2=1.345 $Y2=2.035
r234 31 33 46.1489 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.79 $Y=1.26 $X2=4.88
+ $Y2=1.26
r235 26 60 38.6072 $w=2.91e-07 $l=1.69926e-07 $layer=POLY_cond $X=8.24 $Y=1.945
+ $X2=8.23 $Y2=2.11
r236 26 28 681.979 $w=1.5e-07 $l=1.33e-06 $layer=POLY_cond $X=8.24 $Y=1.945
+ $X2=8.24 $Y2=0.615
r237 23 60 57.6553 $w=2.91e-07 $l=2.82489e-07 $layer=POLY_cond $X=8.235 $Y=2.39
+ $X2=8.23 $Y2=2.11
r238 23 25 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=8.235 $Y=2.39
+ $X2=8.235 $Y2=2.675
r239 20 57 49.7565 $w=4.18e-07 $l=3.16228e-07 $layer=POLY_cond $X=4.895 $Y=2.21
+ $X2=5.045 $Y2=1.96
r240 20 22 101.22 $w=1.5e-07 $l=3.15e-07 $layer=POLY_cond $X=4.895 $Y=2.21
+ $X2=4.895 $Y2=2.525
r241 19 57 39.9551 $w=4.18e-07 $l=2.33345e-07 $layer=POLY_cond $X=4.88 $Y=1.795
+ $X2=5.045 $Y2=1.96
r242 18 33 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.88 $Y=1.335
+ $X2=4.88 $Y2=1.26
r243 18 19 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=4.88 $Y=1.335
+ $X2=4.88 $Y2=1.795
r244 15 31 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.79 $Y=1.185
+ $X2=4.79 $Y2=1.26
r245 15 17 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.79 $Y=1.185
+ $X2=4.79 $Y2=0.9
r246 14 17 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=4.79 $Y=0.255
+ $X2=4.79 $Y2=0.9
r247 12 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.715 $Y=0.18
+ $X2=4.79 $Y2=0.255
r248 12 13 1917.74 $w=1.5e-07 $l=3.74e-06 $layer=POLY_cond $X=4.715 $Y=0.18
+ $X2=0.975 $Y2=0.18
r249 11 30 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.945 $Y=2.75
+ $X2=0.945 $Y2=2.465
r250 8 30 35.9967 $w=2.15e-07 $l=1.07e-07 $layer=POLY_cond $X=0.962 $Y=2.358
+ $X2=0.962 $Y2=2.465
r251 8 55 62.0823 $w=2.15e-07 $l=2.08e-07 $layer=POLY_cond $X=0.962 $Y=2.358
+ $X2=0.962 $Y2=2.15
r252 6 53 10.0949 $w=5.3e-07 $l=1e-07 $layer=POLY_cond $X=1.09 $Y=1.885 $X2=1.09
+ $Y2=1.985
r253 5 49 10.0949 $w=5.3e-07 $l=1e-07 $layer=POLY_cond $X=1.09 $Y=1.405 $X2=1.09
+ $Y2=1.305
r254 5 6 48.4555 $w=5.3e-07 $l=4.8e-07 $layer=POLY_cond $X=1.09 $Y=1.405
+ $X2=1.09 $Y2=1.885
r255 4 51 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=0.9 $Y=0.6 $X2=0.9
+ $Y2=1.14
r256 1 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.9 $Y=0.255
+ $X2=0.975 $Y2=0.18
r257 1 4 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=0.9 $Y=0.255 $X2=0.9
+ $Y2=0.6
.ends

.subckt PM_SKY130_FD_SC_LS__DFRTP_2%A_697_463# 1 2 3 12 14 16 18 19 25 28 29 31
+ 36 41 43 44 47
c126 29 0 1.1997e-19 $X=4.785 $Y=1.435
c127 25 0 9.10107e-20 $X=4.615 $Y=2.485
c128 19 0 1.18794e-19 $X=3.935 $Y=2.637
r129 43 44 5.53573 $w=3.13e-07 $l=8.5e-08 $layer=LI1_cond $X=4.092 $Y=2.485
+ $X2=4.092 $Y2=2.4
r130 39 41 5.91385 $w=3.78e-07 $l=1.95e-07 $layer=LI1_cond $X=3.825 $Y=0.86
+ $X2=4.02 $Y2=0.86
r131 34 47 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=4.785 $Y=2.445
+ $X2=4.7 $Y2=2.445
r132 34 36 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=4.785 $Y=2.445
+ $X2=5.12 $Y2=2.445
r133 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.52
+ $Y=1.41 $X2=5.52 $Y2=1.41
r134 29 31 30.2516 $w=2.78e-07 $l=7.35e-07 $layer=LI1_cond $X=4.785 $Y=1.435
+ $X2=5.52 $Y2=1.435
r135 28 47 2.11342 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.7 $Y=2.32 $X2=4.7
+ $Y2=2.445
r136 27 29 7.36005 $w=2.8e-07 $l=1.77482e-07 $layer=LI1_cond $X=4.7 $Y=1.575
+ $X2=4.785 $Y2=1.435
r137 27 28 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=4.7 $Y=1.575
+ $X2=4.7 $Y2=2.32
r138 26 43 4.34843 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=4.25 $Y=2.485
+ $X2=4.092 $Y2=2.485
r139 25 47 4.3182 $w=2.1e-07 $l=1.03078e-07 $layer=LI1_cond $X=4.615 $Y=2.485
+ $X2=4.7 $Y2=2.445
r140 25 26 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=4.615 $Y=2.485
+ $X2=4.25 $Y2=2.485
r141 23 41 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.02 $Y=1.05
+ $X2=4.02 $Y2=0.86
r142 23 44 88.0749 $w=1.68e-07 $l=1.35e-06 $layer=LI1_cond $X=4.02 $Y=1.05
+ $X2=4.02 $Y2=2.4
r143 19 43 5.56099 $w=3.13e-07 $l=1.52e-07 $layer=LI1_cond $X=4.092 $Y=2.637
+ $X2=4.092 $Y2=2.485
r144 19 21 14.0854 $w=2.23e-07 $l=2.75e-07 $layer=LI1_cond $X=3.935 $Y=2.637
+ $X2=3.66 $Y2=2.637
r145 18 32 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=5.73 $Y=1.41
+ $X2=5.52 $Y2=1.41
r146 14 18 64.0286 $w=1.97e-07 $l=2.70647e-07 $layer=POLY_cond $X=5.905 $Y=1.66
+ $X2=5.862 $Y2=1.41
r147 14 16 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.905 $Y=1.66
+ $X2=5.905 $Y2=2.235
r148 10 18 43.2316 $w=1.97e-07 $l=1.9139e-07 $layer=POLY_cond $X=5.805 $Y=1.245
+ $X2=5.862 $Y2=1.41
r149 10 12 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=5.805 $Y=1.245
+ $X2=5.805 $Y2=0.74
r150 3 36 600 $w=1.7e-07 $l=2.22711e-07 $layer=licon1_PDIFF $count=1 $X=4.97
+ $Y=2.315 $X2=5.12 $Y2=2.475
r151 2 21 600 $w=1.7e-07 $l=3.72357e-07 $layer=licon1_PDIFF $count=1 $X=3.485
+ $Y=2.315 $X2=3.66 $Y2=2.61
r152 1 39 182 $w=1.7e-07 $l=2.82489e-07 $layer=licon1_NDIFF $count=1 $X=3.615
+ $Y=0.69 $X2=3.825 $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_LS__DFRTP_2%A_309_390# 1 2 7 9 10 12 14 15 16 17 18 19
+ 21 24 26 31 32 33 36 38 39 43 46 47 50 51 55
c178 55 0 1.67618e-19 $X=1.69 $Y=2.075
c179 51 0 1.26266e-19 $X=1.665 $Y=1.06
c180 50 0 2.55513e-19 $X=2.565 $Y=1.43
c181 32 0 3.77492e-20 $X=7.255 $Y=1.66
c182 24 0 2.30448e-19 $X=3.915 $Y=2.525
c183 17 0 4.65981e-20 $X=3.465 $Y=1.275
c184 10 0 8.54071e-20 $X=2.535 $Y=1.41
c185 7 0 1.98071e-19 $X=2.4 $Y=1.875
r186 59 63 31.482 $w=4.44e-07 $l=2.9e-07 $layer=POLY_cond $X=2.6 $Y=1.537
+ $X2=2.89 $Y2=1.537
r187 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.6
+ $Y=1.61 $X2=2.6 $Y2=1.61
r188 52 55 6.64871 $w=2.58e-07 $l=1.5e-07 $layer=LI1_cond $X=1.54 $Y=2.03
+ $X2=1.69 $Y2=2.03
r189 50 58 9.63385 $w=2.4e-07 $l=1.8e-07 $layer=LI1_cond $X=2.565 $Y=1.43
+ $X2=2.565 $Y2=1.61
r190 49 50 13.4452 $w=2.38e-07 $l=2.8e-07 $layer=LI1_cond $X=2.565 $Y=1.15
+ $X2=2.565 $Y2=1.43
r191 48 51 3.16872 $w=1.8e-07 $l=2.1e-07 $layer=LI1_cond $X=1.875 $Y=1.06
+ $X2=1.665 $Y2=1.06
r192 47 49 9.49129 $w=1.54e-07 $l=1.58745e-07 $layer=LI1_cond $X=2.445 $Y=1.06
+ $X2=2.565 $Y2=1.15
r193 47 48 35.1212 $w=1.78e-07 $l=5.7e-07 $layer=LI1_cond $X=2.445 $Y=1.06
+ $X2=1.875 $Y2=1.06
r194 46 52 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.54 $Y=1.9 $X2=1.54
+ $Y2=2.03
r195 45 51 3.36599 $w=2.95e-07 $l=1.63936e-07 $layer=LI1_cond $X=1.54 $Y=1.15
+ $X2=1.665 $Y2=1.06
r196 45 46 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=1.54 $Y=1.15
+ $X2=1.54 $Y2=1.9
r197 41 51 3.36599 $w=2.95e-07 $l=9e-08 $layer=LI1_cond $X=1.665 $Y=0.97
+ $X2=1.665 $Y2=1.06
r198 41 43 9.4665 $w=4.18e-07 $l=3.45e-07 $layer=LI1_cond $X=1.665 $Y=0.97
+ $X2=1.665 $Y2=0.625
r199 34 36 497.383 $w=1.5e-07 $l=9.7e-07 $layer=POLY_cond $X=7.33 $Y=1.585
+ $X2=7.33 $Y2=0.615
r200 32 34 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.255 $Y=1.66
+ $X2=7.33 $Y2=1.585
r201 32 33 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=7.255 $Y=1.66
+ $X2=6.485 $Y2=1.66
r202 29 39 105.158 $w=1.8e-07 $l=2.65e-07 $layer=POLY_cond $X=6.41 $Y=2.885
+ $X2=6.41 $Y2=3.15
r203 29 31 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.41 $Y=2.885
+ $X2=6.41 $Y2=2.31
r204 28 33 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.41 $Y=1.735
+ $X2=6.485 $Y2=1.66
r205 28 31 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.41 $Y=1.735
+ $X2=6.41 $Y2=2.31
r206 27 38 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.99 $Y=3.15
+ $X2=3.915 $Y2=3.15
r207 26 39 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=6.32 $Y=3.15 $X2=6.41
+ $Y2=3.15
r208 26 27 1194.74 $w=1.5e-07 $l=2.33e-06 $layer=POLY_cond $X=6.32 $Y=3.15
+ $X2=3.99 $Y2=3.15
r209 22 38 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.915 $Y=3.075
+ $X2=3.915 $Y2=3.15
r210 22 24 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=3.915 $Y=3.075
+ $X2=3.915 $Y2=2.525
r211 19 21 96.4 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=3.54 $Y=1.2 $X2=3.54
+ $Y2=0.9
r212 18 63 43.7957 $w=4.44e-07 $l=3.46026e-07 $layer=POLY_cond $X=3.085 $Y=1.275
+ $X2=2.89 $Y2=1.537
r213 17 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.465 $Y=1.275
+ $X2=3.54 $Y2=1.2
r214 17 18 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=3.465 $Y=1.275
+ $X2=3.085 $Y2=1.275
r215 15 38 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.84 $Y=3.15
+ $X2=3.915 $Y2=3.15
r216 15 16 448.67 $w=1.5e-07 $l=8.75e-07 $layer=POLY_cond $X=3.84 $Y=3.15
+ $X2=2.965 $Y2=3.15
r217 14 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.89 $Y=3.075
+ $X2=2.965 $Y2=3.15
r218 13 63 28.433 $w=1.5e-07 $l=3.38e-07 $layer=POLY_cond $X=2.89 $Y=1.875
+ $X2=2.89 $Y2=1.537
r219 13 14 615.319 $w=1.5e-07 $l=1.2e-06 $layer=POLY_cond $X=2.89 $Y=1.875
+ $X2=2.89 $Y2=3.075
r220 10 59 7.05631 $w=4.44e-07 $l=6.5e-08 $layer=POLY_cond $X=2.535 $Y=1.537
+ $X2=2.6 $Y2=1.537
r221 10 60 14.6554 $w=4.44e-07 $l=1.35e-07 $layer=POLY_cond $X=2.535 $Y=1.537
+ $X2=2.4 $Y2=1.537
r222 10 12 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.535 $Y=1.41
+ $X2=2.535 $Y2=0.965
r223 7 60 28.433 $w=1.5e-07 $l=3.38e-07 $layer=POLY_cond $X=2.4 $Y=1.875 $X2=2.4
+ $Y2=1.537
r224 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.4 $Y=1.875 $X2=2.4
+ $Y2=2.45
r225 2 55 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.545
+ $Y=1.95 $X2=1.69 $Y2=2.075
r226 1 43 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=1.565
+ $Y=0.48 $X2=1.71 $Y2=0.625
.ends

.subckt PM_SKY130_FD_SC_LS__DFRTP_2%A_1525_212# 1 2 9 13 14 15 17 18 19 21 27 30
+ 31 32 33 36 38 39 43
c118 39 0 1.33493e-19 $X=7.79 $Y=1.225
c119 36 0 4.37308e-20 $X=9.29 $Y=2.105
c120 21 0 4.77539e-20 $X=8.715 $Y=2.61
c121 13 0 3.83476e-20 $X=7.735 $Y=2.065
r122 39 46 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.79 $Y=1.225
+ $X2=7.79 $Y2=1.39
r123 39 45 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.79 $Y=1.225
+ $X2=7.79 $Y2=1.06
r124 38 41 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=7.79 $Y=1.225 $X2=7.79
+ $Y2=1.305
r125 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.79
+ $Y=1.225 $X2=7.79 $Y2=1.225
r126 35 36 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=9.29 $Y=1.39
+ $X2=9.29 $Y2=2.105
r127 34 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.01 $Y=1.305
+ $X2=8.845 $Y2=1.305
r128 33 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.205 $Y=1.305
+ $X2=9.29 $Y2=1.39
r129 33 34 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=9.205 $Y=1.305
+ $X2=9.01 $Y2=1.305
r130 31 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.205 $Y=2.19
+ $X2=9.29 $Y2=2.105
r131 31 32 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=9.205 $Y=2.19
+ $X2=8.885 $Y2=2.19
r132 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.8 $Y=2.275
+ $X2=8.885 $Y2=2.19
r133 29 30 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=8.8 $Y=2.275
+ $X2=8.8 $Y2=2.445
r134 25 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.845 $Y=1.22
+ $X2=8.845 $Y2=1.305
r135 25 27 21.1281 $w=3.28e-07 $l=6.05e-07 $layer=LI1_cond $X=8.845 $Y=1.22
+ $X2=8.845 $Y2=0.615
r136 21 30 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.715 $Y=2.61
+ $X2=8.8 $Y2=2.445
r137 21 23 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=8.715 $Y=2.61
+ $X2=8.59 $Y2=2.61
r138 20 41 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.955 $Y=1.305
+ $X2=7.79 $Y2=1.305
r139 19 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.68 $Y=1.305
+ $X2=8.845 $Y2=1.305
r140 19 20 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=8.68 $Y=1.305
+ $X2=7.955 $Y2=1.305
r141 18 46 299.968 $w=1.5e-07 $l=5.85e-07 $layer=POLY_cond $X=7.72 $Y=1.975
+ $X2=7.72 $Y2=1.39
r142 15 17 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.735 $Y=2.39
+ $X2=7.735 $Y2=2.675
r143 14 15 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=7.735 $Y=2.3
+ $X2=7.735 $Y2=2.39
r144 13 18 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=7.735 $Y=2.065
+ $X2=7.735 $Y2=1.975
r145 13 14 91.3468 $w=1.8e-07 $l=2.35e-07 $layer=POLY_cond $X=7.735 $Y=2.065
+ $X2=7.735 $Y2=2.3
r146 9 45 228.181 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=7.72 $Y=0.615
+ $X2=7.72 $Y2=1.06
r147 2 23 600 $w=1.7e-07 $l=3.44964e-07 $layer=licon1_PDIFF $count=1 $X=8.31
+ $Y=2.465 $X2=8.59 $Y2=2.61
r148 1 27 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=8.705
+ $Y=0.405 $X2=8.845 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_LS__DFRTP_2%A_1271_74# 1 2 9 12 13 15 16 17 19 20 22 25
+ 27 28 29 31 34 36 37 41 42 43 48 50
c148 41 0 1.53326e-19 $X=7.54 $Y=2.475
c149 17 0 4.77539e-20 $X=9.035 $Y=1.63
c150 12 0 1.36674e-19 $X=8.945 $Y=2.3
r151 54 58 13.0505 $w=2.77e-07 $l=7.5e-08 $layer=POLY_cond $X=8.87 $Y=1.722
+ $X2=8.945 $Y2=1.722
r152 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.87
+ $Y=1.725 $X2=8.87 $Y2=1.725
r153 50 53 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=8.87 $Y=1.645 $X2=8.87
+ $Y2=1.725
r154 46 48 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=6.44 $Y=1.6 $X2=6.6
+ $Y2=1.6
r155 42 50 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.705 $Y=1.645
+ $X2=8.87 $Y2=1.645
r156 42 43 70.4599 $w=1.68e-07 $l=1.08e-06 $layer=LI1_cond $X=8.705 $Y=1.645
+ $X2=7.625 $Y2=1.645
r157 40 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.54 $Y=1.73
+ $X2=7.625 $Y2=1.645
r158 40 41 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=7.54 $Y=1.73
+ $X2=7.54 $Y2=2.475
r159 37 39 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=6.685 $Y=2.64
+ $X2=7.09 $Y2=2.64
r160 36 41 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.455 $Y=2.64
+ $X2=7.54 $Y2=2.475
r161 36 39 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=7.455 $Y=2.64
+ $X2=7.09 $Y2=2.64
r162 32 45 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.525 $Y=0.72
+ $X2=6.44 $Y2=0.72
r163 32 34 19.5915 $w=2.48e-07 $l=4.25e-07 $layer=LI1_cond $X=6.525 $Y=0.72
+ $X2=6.95 $Y2=0.72
r164 31 37 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.6 $Y=2.475
+ $X2=6.685 $Y2=2.64
r165 30 48 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.6 $Y=1.685
+ $X2=6.6 $Y2=1.6
r166 30 31 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=6.6 $Y=1.685
+ $X2=6.6 $Y2=2.475
r167 29 46 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.44 $Y=1.515
+ $X2=6.44 $Y2=1.6
r168 28 45 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.44 $Y=0.845
+ $X2=6.44 $Y2=0.72
r169 28 29 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.44 $Y=0.845
+ $X2=6.44 $Y2=1.515
r170 23 27 18.8402 $w=1.65e-07 $l=9.60469e-08 $layer=POLY_cond $X=9.61 $Y=1.555
+ $X2=9.562 $Y2=1.63
r171 23 25 417.904 $w=1.5e-07 $l=8.15e-07 $layer=POLY_cond $X=9.61 $Y=1.555
+ $X2=9.61 $Y2=0.74
r172 20 22 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=9.53 $Y=1.97
+ $X2=9.53 $Y2=2.465
r173 19 20 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=9.53 $Y=1.88 $X2=9.53
+ $Y2=1.97
r174 18 27 18.8402 $w=1.65e-07 $l=8.95824e-08 $layer=POLY_cond $X=9.53 $Y=1.705
+ $X2=9.562 $Y2=1.63
r175 18 19 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=9.53 $Y=1.705
+ $X2=9.53 $Y2=1.88
r176 17 58 25.7246 $w=2.77e-07 $l=1.29399e-07 $layer=POLY_cond $X=9.035 $Y=1.63
+ $X2=8.945 $Y2=1.722
r177 16 27 6.66866 $w=1.5e-07 $l=1.22e-07 $layer=POLY_cond $X=9.44 $Y=1.63
+ $X2=9.562 $Y2=1.63
r178 16 17 207.67 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=9.44 $Y=1.63
+ $X2=9.035 $Y2=1.63
r179 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=8.945 $Y=2.39
+ $X2=8.945 $Y2=2.675
r180 12 13 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=8.945 $Y=2.3
+ $X2=8.945 $Y2=2.39
r181 11 58 12.8788 $w=1.8e-07 $l=1.68e-07 $layer=POLY_cond $X=8.945 $Y=1.89
+ $X2=8.945 $Y2=1.722
r182 11 12 159.371 $w=1.8e-07 $l=4.1e-07 $layer=POLY_cond $X=8.945 $Y=1.89
+ $X2=8.945 $Y2=2.3
r183 7 54 41.7617 $w=2.77e-07 $l=3.12538e-07 $layer=POLY_cond $X=8.63 $Y=1.555
+ $X2=8.87 $Y2=1.722
r184 7 9 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=8.63 $Y=1.555 $X2=8.63
+ $Y2=0.615
r185 2 39 300 $w=1.7e-07 $l=1.09135e-06 $layer=licon1_PDIFF $count=2 $X=6.485
+ $Y=1.81 $X2=7.09 $Y2=2.64
r186 1 45 182 $w=1.7e-07 $l=3.83732e-07 $layer=licon1_NDIFF $count=1 $X=6.355
+ $Y=0.37 $X2=6.52 $Y2=0.68
r187 1 34 182 $w=1.7e-07 $l=7.33809e-07 $layer=licon1_NDIFF $count=1 $X=6.355
+ $Y=0.37 $X2=6.95 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_LS__DFRTP_2%A_1921_409# 1 2 7 10 11 13 16 18 21 22 24 27
+ 29 30 33 37 41 46 49
c72 49 0 4.37308e-20 $X=10.09 $Y=1.375
c73 33 0 1.36674e-19 $X=9.755 $Y=2.195
r74 47 49 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=10.09 $Y=1.465
+ $X2=10.09 $Y2=1.375
r75 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.09
+ $Y=1.465 $X2=10.09 $Y2=1.465
r76 44 46 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=9.825 $Y=1.465
+ $X2=10.09 $Y2=1.465
r77 42 44 1.22229 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=9.79 $Y=1.465
+ $X2=9.825 $Y2=1.465
r78 39 42 2.13598 $w=2.6e-07 $l=1.65e-07 $layer=LI1_cond $X=9.79 $Y=1.63
+ $X2=9.79 $Y2=1.465
r79 39 41 17.7299 $w=2.58e-07 $l=4e-07 $layer=LI1_cond $X=9.79 $Y=1.63 $X2=9.79
+ $Y2=2.03
r80 35 44 0.716491 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=9.825 $Y=1.3
+ $X2=9.825 $Y2=1.465
r81 35 37 27.4142 $w=3.28e-07 $l=7.85e-07 $layer=LI1_cond $X=9.825 $Y=1.3
+ $X2=9.825 $Y2=0.515
r82 33 41 6.31279 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=9.755 $Y=2.195
+ $X2=9.755 $Y2=2.03
r83 25 30 18.8402 $w=1.65e-07 $l=8.21584e-08 $layer=POLY_cond $X=11.03 $Y=1.3
+ $X2=11.015 $Y2=1.375
r84 25 27 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=11.03 $Y=1.3
+ $X2=11.03 $Y2=0.74
r85 22 24 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=11.015 $Y=1.765
+ $X2=11.015 $Y2=2.4
r86 21 22 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=11.015 $Y=1.675
+ $X2=11.015 $Y2=1.765
r87 20 30 18.8402 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=11.015 $Y=1.45
+ $X2=11.015 $Y2=1.375
r88 20 21 87.4597 $w=1.8e-07 $l=2.25e-07 $layer=POLY_cond $X=11.015 $Y=1.45
+ $X2=11.015 $Y2=1.675
r89 19 29 13.2179 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=10.675 $Y=1.375
+ $X2=10.575 $Y2=1.375
r90 18 30 6.66866 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=10.925 $Y=1.375
+ $X2=11.015 $Y2=1.375
r91 18 19 128.191 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=10.925 $Y=1.375
+ $X2=10.675 $Y2=1.375
r92 14 29 10.9219 $w=1.5e-07 $l=8.66025e-08 $layer=POLY_cond $X=10.6 $Y=1.3
+ $X2=10.575 $Y2=1.375
r93 14 16 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=10.6 $Y=1.3 $X2=10.6
+ $Y2=0.74
r94 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=10.565 $Y=1.765
+ $X2=10.565 $Y2=2.4
r95 10 11 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=10.565 $Y=1.675
+ $X2=10.565 $Y2=1.765
r96 9 29 10.9219 $w=1.8e-07 $l=7.98436e-08 $layer=POLY_cond $X=10.565 $Y=1.45
+ $X2=10.575 $Y2=1.375
r97 9 10 87.4597 $w=1.8e-07 $l=2.25e-07 $layer=POLY_cond $X=10.565 $Y=1.45
+ $X2=10.565 $Y2=1.675
r98 8 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.255 $Y=1.375
+ $X2=10.09 $Y2=1.375
r99 7 29 13.2179 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=10.475 $Y=1.375
+ $X2=10.575 $Y2=1.375
r100 7 8 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=10.475 $Y=1.375
+ $X2=10.255 $Y2=1.375
r101 2 33 300 $w=1.7e-07 $l=2.12132e-07 $layer=licon1_PDIFF $count=2 $X=9.605
+ $Y=2.045 $X2=9.755 $Y2=2.195
r102 1 37 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.685
+ $Y=0.37 $X2=9.825 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__DFRTP_2%VPWR 1 2 3 4 5 6 7 8 9 28 30 34 38 42 44 48
+ 54 58 62 66 68 73 74 75 77 82 87 95 107 111 120 123 126 129 132 135 139
r159 138 139 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r160 135 136 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r161 132 133 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r162 129 130 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r163 127 130 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r164 126 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r165 123 124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r166 120 121 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r167 117 118 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r168 115 139 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=11.28 $Y2=3.33
r169 115 136 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=10.32 $Y2=3.33
r170 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r171 112 135 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.48 $Y=3.33
+ $X2=10.315 $Y2=3.33
r172 112 114 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=10.48 $Y=3.33
+ $X2=10.8 $Y2=3.33
r173 111 138 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=11.155 $Y=3.33
+ $X2=11.337 $Y2=3.33
r174 111 114 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=11.155 $Y=3.33
+ $X2=10.8 $Y2=3.33
r175 110 136 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=10.32 $Y2=3.33
r176 109 110 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r177 107 135 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.15 $Y=3.33
+ $X2=10.315 $Y2=3.33
r178 107 109 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=10.15 $Y=3.33
+ $X2=9.84 $Y2=3.33
r179 106 110 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=9.84 $Y2=3.33
r180 106 133 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=7.92 $Y2=3.33
r181 105 106 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r182 103 132 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.125 $Y=3.33
+ $X2=7.96 $Y2=3.33
r183 103 105 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=8.125 $Y=3.33
+ $X2=8.88 $Y2=3.33
r184 102 133 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r185 101 102 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r186 99 102 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=7.44 $Y2=3.33
r187 98 101 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=6 $Y=3.33
+ $X2=7.44 $Y2=3.33
r188 98 99 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r189 96 129 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.845 $Y=3.33
+ $X2=5.68 $Y2=3.33
r190 96 98 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=5.845 $Y=3.33
+ $X2=6 $Y2=3.33
r191 95 132 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.795 $Y=3.33
+ $X2=7.96 $Y2=3.33
r192 95 101 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=7.795 $Y=3.33
+ $X2=7.44 $Y2=3.33
r193 94 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r194 93 94 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r195 91 94 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=4.08 $Y2=3.33
r196 91 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r197 90 93 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.64 $Y=3.33
+ $X2=4.08 $Y2=3.33
r198 90 91 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r199 88 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.285 $Y=3.33
+ $X2=2.12 $Y2=3.33
r200 88 90 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=2.285 $Y=3.33
+ $X2=2.64 $Y2=3.33
r201 87 126 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.42 $Y=3.33
+ $X2=4.585 $Y2=3.33
r202 87 93 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=4.42 $Y=3.33
+ $X2=4.08 $Y2=3.33
r203 86 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r204 86 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r205 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r206 83 120 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.345 $Y=3.33
+ $X2=1.18 $Y2=3.33
r207 83 85 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.345 $Y=3.33
+ $X2=1.68 $Y2=3.33
r208 82 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.955 $Y=3.33
+ $X2=2.12 $Y2=3.33
r209 82 85 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.955 $Y=3.33
+ $X2=1.68 $Y2=3.33
r210 81 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r211 81 118 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r212 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r213 78 117 4.75569 $w=1.7e-07 $l=2.18e-07 $layer=LI1_cond $X=0.435 $Y=3.33
+ $X2=0.217 $Y2=3.33
r214 78 80 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.435 $Y=3.33
+ $X2=0.72 $Y2=3.33
r215 77 120 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.015 $Y=3.33
+ $X2=1.18 $Y2=3.33
r216 77 80 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.015 $Y=3.33
+ $X2=0.72 $Y2=3.33
r217 75 99 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=5.76 $Y=3.33
+ $X2=6 $Y2=3.33
r218 75 130 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=5.76 $Y=3.33
+ $X2=5.52 $Y2=3.33
r219 73 105 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=9.09 $Y=3.33
+ $X2=8.88 $Y2=3.33
r220 73 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.09 $Y=3.33
+ $X2=9.255 $Y2=3.33
r221 72 109 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=9.42 $Y=3.33
+ $X2=9.84 $Y2=3.33
r222 72 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.42 $Y=3.33
+ $X2=9.255 $Y2=3.33
r223 68 71 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=11.28 $Y=1.985
+ $X2=11.28 $Y2=2.815
r224 66 138 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=11.28 $Y=3.245
+ $X2=11.337 $Y2=3.33
r225 66 71 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=11.28 $Y=3.245
+ $X2=11.28 $Y2=2.815
r226 62 65 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=10.315 $Y=1.985
+ $X2=10.315 $Y2=2.815
r227 60 135 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.315 $Y=3.245
+ $X2=10.315 $Y2=3.33
r228 60 65 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=10.315 $Y=3.245
+ $X2=10.315 $Y2=2.815
r229 56 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.255 $Y=3.245
+ $X2=9.255 $Y2=3.33
r230 56 58 19.9058 $w=3.28e-07 $l=5.7e-07 $layer=LI1_cond $X=9.255 $Y=3.245
+ $X2=9.255 $Y2=2.675
r231 52 132 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.96 $Y=3.245
+ $X2=7.96 $Y2=3.33
r232 52 54 19.9058 $w=3.28e-07 $l=5.7e-07 $layer=LI1_cond $X=7.96 $Y=3.245
+ $X2=7.96 $Y2=2.675
r233 48 51 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=5.68 $Y=1.91
+ $X2=5.68 $Y2=2.59
r234 46 129 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.68 $Y=3.245
+ $X2=5.68 $Y2=3.33
r235 46 51 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=5.68 $Y=3.245
+ $X2=5.68 $Y2=2.59
r236 45 126 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.75 $Y=3.33
+ $X2=4.585 $Y2=3.33
r237 44 129 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.515 $Y=3.33
+ $X2=5.68 $Y2=3.33
r238 44 45 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=5.515 $Y=3.33
+ $X2=4.75 $Y2=3.33
r239 40 126 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.585 $Y=3.245
+ $X2=4.585 $Y2=3.33
r240 40 42 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=4.585 $Y=3.245
+ $X2=4.585 $Y2=2.84
r241 36 123 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.12 $Y=3.245
+ $X2=2.12 $Y2=3.33
r242 36 38 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=2.12 $Y=3.245
+ $X2=2.12 $Y2=2.825
r243 32 120 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.18 $Y=3.245
+ $X2=1.18 $Y2=3.33
r244 32 34 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=1.18 $Y=3.245
+ $X2=1.18 $Y2=2.815
r245 28 117 3.01048 $w=3.3e-07 $l=1.08305e-07 $layer=LI1_cond $X=0.27 $Y=3.245
+ $X2=0.217 $Y2=3.33
r246 28 30 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=0.27 $Y=3.245
+ $X2=0.27 $Y2=2.75
r247 9 71 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=11.09
+ $Y=1.84 $X2=11.24 $Y2=2.815
r248 9 68 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=11.09
+ $Y=1.84 $X2=11.24 $Y2=1.985
r249 8 65 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=10.17
+ $Y=1.84 $X2=10.315 $Y2=2.815
r250 8 62 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=10.17
+ $Y=1.84 $X2=10.315 $Y2=1.985
r251 7 58 600 $w=1.7e-07 $l=3.23381e-07 $layer=licon1_PDIFF $count=1 $X=9.02
+ $Y=2.465 $X2=9.255 $Y2=2.675
r252 6 54 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=7.81
+ $Y=2.465 $X2=7.96 $Y2=2.675
r253 5 51 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=5.535
+ $Y=1.735 $X2=5.68 $Y2=2.59
r254 5 48 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=5.535
+ $Y=1.735 $X2=5.68 $Y2=1.91
r255 4 42 600 $w=1.7e-07 $l=6.31664e-07 $layer=licon1_PDIFF $count=1 $X=4.35
+ $Y=2.315 $X2=4.585 $Y2=2.84
r256 3 38 600 $w=1.7e-07 $l=9.42404e-07 $layer=licon1_PDIFF $count=1 $X=1.98
+ $Y=1.95 $X2=2.12 $Y2=2.825
r257 2 34 600 $w=1.7e-07 $l=3.45868e-07 $layer=licon1_PDIFF $count=1 $X=1.02
+ $Y=2.54 $X2=1.18 $Y2=2.815
r258 1 30 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.54 $X2=0.27 $Y2=2.75
.ends

.subckt PM_SKY130_FD_SC_LS__DFRTP_2%A_30_78# 1 2 3 4 13 17 20 21 23 26 27 30 32
+ 36 39 42 47
c128 42 0 9.78499e-20 $X=3.325 $Y=0.88
c129 39 0 3.37508e-19 $X=3.195 $Y=2.495
c130 30 0 1.40697e-19 $X=3.68 $Y=2.185
c131 26 0 1.73746e-19 $X=3.405 $Y=1.22
r132 45 47 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3.405 $Y=1.305
+ $X2=3.68 $Y2=1.305
r133 42 44 8.79328 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=3.365 $Y=0.88
+ $X2=3.365 $Y2=1.045
r134 39 40 1.37299 $w=3.11e-07 $l=3.5e-08 $layer=LI1_cond $X=3.157 $Y=2.495
+ $X2=3.157 $Y2=2.53
r135 37 39 8.82637 $w=3.11e-07 $l=2.25e-07 $layer=LI1_cond $X=3.157 $Y=2.27
+ $X2=3.157 $Y2=2.495
r136 32 34 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=0.295 $Y=0.6
+ $X2=0.295 $Y2=0.745
r137 29 47 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.68 $Y=1.39
+ $X2=3.68 $Y2=1.305
r138 29 30 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=3.68 $Y=1.39
+ $X2=3.68 $Y2=2.185
r139 28 37 4.27302 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=3.37 $Y=2.27
+ $X2=3.157 $Y2=2.27
r140 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.595 $Y=2.27
+ $X2=3.68 $Y2=2.185
r141 27 28 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=3.595 $Y=2.27
+ $X2=3.37 $Y2=2.27
r142 26 45 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.405 $Y=1.22
+ $X2=3.405 $Y2=1.305
r143 26 44 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.405 $Y=1.22
+ $X2=3.405 $Y2=1.045
r144 23 40 4.27302 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=2.945 $Y=2.53
+ $X2=3.157 $Y2=2.53
r145 23 24 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=2.945 $Y=2.53
+ $X2=2.485 $Y2=2.53
r146 22 36 0.571601 $w=2.3e-07 $l=2.90086e-07 $layer=LI1_cond $X=0.89 $Y=2.445
+ $X2=0.635 $Y2=2.52
r147 21 24 56.3077 $w=2.34e-07 $l=1.1217e-06 $layer=LI1_cond $X=1.405 $Y=2.445
+ $X2=2.485 $Y2=2.53
r148 21 22 25.8047 $w=2.28e-07 $l=5.15e-07 $layer=LI1_cond $X=1.405 $Y=2.445
+ $X2=0.89 $Y2=2.445
r149 20 36 6.1674 $w=1.85e-07 $l=2.40728e-07 $layer=LI1_cond $X=0.75 $Y=2.33
+ $X2=0.635 $Y2=2.52
r150 19 20 97.861 $w=1.68e-07 $l=1.5e-06 $layer=LI1_cond $X=0.75 $Y=0.83
+ $X2=0.75 $Y2=2.33
r151 15 36 6.1674 $w=1.85e-07 $l=1.51987e-07 $layer=LI1_cond $X=0.735 $Y=2.63
+ $X2=0.635 $Y2=2.52
r152 15 17 6.65455 $w=1.98e-07 $l=1.2e-07 $layer=LI1_cond $X=0.735 $Y=2.63
+ $X2=0.735 $Y2=2.75
r153 14 34 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.46 $Y=0.745
+ $X2=0.295 $Y2=0.745
r154 13 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.665 $Y=0.745
+ $X2=0.75 $Y2=0.83
r155 13 14 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=0.665 $Y=0.745
+ $X2=0.46 $Y2=0.745
r156 4 39 600 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_PDIFF $count=1 $X=3.07
+ $Y=2.315 $X2=3.195 $Y2=2.495
r157 3 17 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=0.57
+ $Y=2.54 $X2=0.72 $Y2=2.75
r158 2 42 182 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_NDIFF $count=1 $X=3.18
+ $Y=0.69 $X2=3.325 $Y2=0.88
r159 1 32 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.15
+ $Y=0.39 $X2=0.295 $Y2=0.6
.ends

.subckt PM_SKY130_FD_SC_LS__DFRTP_2%Q 1 2 7 8 9 10 11 12 13
r22 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=10.815 $Y=2.405
+ $X2=10.815 $Y2=2.775
r23 11 12 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=10.815 $Y=1.985
+ $X2=10.815 $Y2=2.405
r24 10 11 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=10.815 $Y=1.665
+ $X2=10.815 $Y2=1.985
r25 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=10.815 $Y=1.295
+ $X2=10.815 $Y2=1.665
r26 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=10.815 $Y=0.925
+ $X2=10.815 $Y2=1.295
r27 7 8 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=10.815 $Y=0.515
+ $X2=10.815 $Y2=0.925
r28 2 13 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=10.64
+ $Y=1.84 $X2=10.79 $Y2=2.815
r29 2 11 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=10.64
+ $Y=1.84 $X2=10.79 $Y2=1.985
r30 1 7 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.675
+ $Y=0.37 $X2=10.815 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__DFRTP_2%VGND 1 2 3 4 5 6 7 24 26 30 34 38 42 44 46
+ 48 50 55 63 71 76 81 87 90 100 103 106 110
c116 110 0 1.99579e-19 $X=11.28 $Y=0
r117 109 110 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r118 106 107 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r119 103 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r120 100 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r121 90 91 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r122 88 91 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r123 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r124 85 110 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=11.28 $Y2=0
r125 85 107 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=10.32 $Y2=0
r126 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=0 $X2=10.8
+ $Y2=0
r127 82 106 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.47 $Y=0
+ $X2=10.345 $Y2=0
r128 82 84 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=10.47 $Y=0 $X2=10.8
+ $Y2=0
r129 81 109 4.01803 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=11.16 $Y=0
+ $X2=11.34 $Y2=0
r130 81 84 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=11.16 $Y=0 $X2=10.8
+ $Y2=0
r131 80 107 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=10.32 $Y2=0
r132 80 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=9.36 $Y2=0
r133 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r134 77 103 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.48 $Y=0
+ $X2=9.355 $Y2=0
r135 77 79 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=9.48 $Y=0 $X2=9.84
+ $Y2=0
r136 76 106 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.22 $Y=0
+ $X2=10.345 $Y2=0
r137 76 79 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=10.22 $Y=0 $X2=9.84
+ $Y2=0
r138 75 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0
+ $X2=9.36 $Y2=0
r139 75 101 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.88 $Y=0
+ $X2=7.92 $Y2=0
r140 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r141 72 100 10.1275 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=8.19 $Y=0 $X2=7.98
+ $Y2=0
r142 72 74 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=8.19 $Y=0 $X2=8.88
+ $Y2=0
r143 71 103 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.23 $Y=0
+ $X2=9.355 $Y2=0
r144 71 74 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=9.23 $Y=0 $X2=8.88
+ $Y2=0
r145 70 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=7.92 $Y2=0
r146 69 70 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r147 67 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r148 66 69 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=5.52 $Y=0 $X2=7.44
+ $Y2=0
r149 66 67 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r150 64 66 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=5.345 $Y=0
+ $X2=5.52 $Y2=0
r151 63 100 10.1275 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=7.77 $Y=0 $X2=7.98
+ $Y2=0
r152 63 69 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=7.77 $Y=0 $X2=7.44
+ $Y2=0
r153 62 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r154 61 62 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r155 59 62 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=4.56 $Y2=0
r156 59 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r157 58 61 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=2.64 $Y=0 $X2=4.56
+ $Y2=0
r158 58 59 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r159 56 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.425 $Y=0 $X2=2.26
+ $Y2=0
r160 56 58 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.425 $Y=0
+ $X2=2.64 $Y2=0
r161 55 97 7.59257 $w=4.23e-07 $l=2.8e-07 $layer=LI1_cond $X=5.132 $Y=0
+ $X2=5.132 $Y2=0.28
r162 55 64 6.14847 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=5.132 $Y=0
+ $X2=5.345 $Y2=0
r163 55 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r164 55 61 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=4.92 $Y=0 $X2=4.56
+ $Y2=0
r165 53 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r166 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r167 50 87 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=1.005 $Y=0 $X2=1.145
+ $Y2=0
r168 50 52 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.005 $Y=0
+ $X2=0.72 $Y2=0
r169 48 70 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=5.76 $Y=0
+ $X2=7.44 $Y2=0
r170 48 67 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=5.76 $Y=0
+ $X2=5.52 $Y2=0
r171 44 109 3.12513 $w=2.5e-07 $l=1.09087e-07 $layer=LI1_cond $X=11.285 $Y=0.085
+ $X2=11.34 $Y2=0
r172 44 46 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=11.285 $Y=0.085
+ $X2=11.285 $Y2=0.515
r173 40 106 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=10.345 $Y=0.085
+ $X2=10.345 $Y2=0
r174 40 42 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=10.345 $Y=0.085
+ $X2=10.345 $Y2=0.515
r175 36 103 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.355 $Y=0.085
+ $X2=9.355 $Y2=0
r176 36 38 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=9.355 $Y=0.085
+ $X2=9.355 $Y2=0.515
r177 32 100 1.60615 $w=4.2e-07 $l=8.5e-08 $layer=LI1_cond $X=7.98 $Y=0.085
+ $X2=7.98 $Y2=0
r178 32 34 12.7592 $w=4.18e-07 $l=4.65e-07 $layer=LI1_cond $X=7.98 $Y=0.085
+ $X2=7.98 $Y2=0.55
r179 28 90 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.26 $Y=0.085
+ $X2=2.26 $Y2=0
r180 28 30 22.0012 $w=3.28e-07 $l=6.3e-07 $layer=LI1_cond $X=2.26 $Y=0.085
+ $X2=2.26 $Y2=0.715
r181 27 87 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=1.285 $Y=0 $X2=1.145
+ $Y2=0
r182 26 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.095 $Y=0 $X2=2.26
+ $Y2=0
r183 26 27 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=2.095 $Y=0
+ $X2=1.285 $Y2=0
r184 22 87 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.145 $Y=0.085
+ $X2=1.145 $Y2=0
r185 22 24 21.1967 $w=2.78e-07 $l=5.15e-07 $layer=LI1_cond $X=1.145 $Y=0.085
+ $X2=1.145 $Y2=0.6
r186 7 46 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=11.105
+ $Y=0.37 $X2=11.245 $Y2=0.515
r187 6 42 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=10.24
+ $Y=0.37 $X2=10.385 $Y2=0.515
r188 5 38 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.255
+ $Y=0.37 $X2=9.395 $Y2=0.515
r189 4 34 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=7.795
+ $Y=0.405 $X2=7.98 $Y2=0.55
r190 3 97 182 $w=1.7e-07 $l=5.2607e-07 $layer=licon1_NDIFF $count=1 $X=4.865
+ $Y=0.69 $X2=5.13 $Y2=0.28
r191 2 30 182 $w=1.7e-07 $l=2.52982e-07 $layer=licon1_NDIFF $count=1 $X=2.06
+ $Y=0.595 $X2=2.26 $Y2=0.715
r192 1 24 182 $w=1.7e-07 $l=2.84341e-07 $layer=licon1_NDIFF $count=1 $X=0.975
+ $Y=0.39 $X2=1.15 $Y2=0.6
.ends

