* File: sky130_fd_sc_ls__nand3_1.pxi.spice
* Created: Wed Sep  2 11:12:05 2020
* 
x_PM_SKY130_FD_SC_LS__NAND3_1%C N_C_c_36_n N_C_c_37_n N_C_M1003_g N_C_c_38_n
+ N_C_M1001_g C C PM_SKY130_FD_SC_LS__NAND3_1%C
x_PM_SKY130_FD_SC_LS__NAND3_1%B N_B_c_59_n N_B_M1000_g N_B_c_60_n N_B_M1004_g B
+ B B PM_SKY130_FD_SC_LS__NAND3_1%B
x_PM_SKY130_FD_SC_LS__NAND3_1%A N_A_c_93_n N_A_M1005_g N_A_c_94_n N_A_M1002_g A
+ PM_SKY130_FD_SC_LS__NAND3_1%A
x_PM_SKY130_FD_SC_LS__NAND3_1%VPWR N_VPWR_M1003_s N_VPWR_M1004_d N_VPWR_c_122_n
+ N_VPWR_c_123_n N_VPWR_c_124_n N_VPWR_c_125_n N_VPWR_c_126_n VPWR
+ N_VPWR_c_127_n N_VPWR_c_121_n PM_SKY130_FD_SC_LS__NAND3_1%VPWR
x_PM_SKY130_FD_SC_LS__NAND3_1%Y N_Y_M1005_d N_Y_M1003_d N_Y_M1002_d N_Y_c_153_n
+ N_Y_c_154_n N_Y_c_150_n N_Y_c_155_n N_Y_c_151_n N_Y_c_152_n N_Y_c_157_n Y Y Y
+ N_Y_c_158_n PM_SKY130_FD_SC_LS__NAND3_1%Y
x_PM_SKY130_FD_SC_LS__NAND3_1%VGND N_VGND_M1001_s N_VGND_c_197_n N_VGND_c_198_n
+ N_VGND_c_199_n VGND N_VGND_c_200_n N_VGND_c_201_n
+ PM_SKY130_FD_SC_LS__NAND3_1%VGND
cc_1 VNB N_C_c_36_n 0.0557536f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.385
cc_2 VNB N_C_c_37_n 0.0231155f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.765
cc_3 VNB N_C_c_38_n 0.0208066f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.22
cc_4 VNB C 0.0311109f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_5 VNB N_B_c_59_n 0.0180991f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.385
cc_6 VNB N_B_c_60_n 0.0394073f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=2.4
cc_7 VNB B 0.00244094f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=0.74
cc_8 VNB N_A_c_93_n 0.0229091f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.385
cc_9 VNB N_A_c_94_n 0.04016f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=2.4
cc_10 VNB A 0.00684394f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=0.74
cc_11 VNB N_VPWR_c_121_n 0.103974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_Y_c_150_n 0.02133f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.385
cc_13 VNB N_Y_c_151_n 0.0320047f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_Y_c_152_n 0.0146427f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_VGND_c_197_n 0.0344107f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.22
cc_16 VNB N_VGND_c_198_n 0.0123263f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_17 VNB N_VGND_c_199_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_18 VNB N_VGND_c_200_n 0.0529515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_VGND_c_201_n 0.18517f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VPB N_C_c_37_n 0.0276786f $X=-0.19 $Y=1.66 $X2=0.655 $Y2=1.765
cc_21 VPB N_B_c_60_n 0.0228813f $X=-0.19 $Y=1.66 $X2=0.655 $Y2=2.4
cc_22 VPB N_A_c_94_n 0.0282492f $X=-0.19 $Y=1.66 $X2=0.655 $Y2=2.4
cc_23 VPB N_VPWR_c_122_n 0.012885f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=0.74
cc_24 VPB N_VPWR_c_123_n 0.0563116f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_25 VPB N_VPWR_c_124_n 0.00976973f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.385
cc_26 VPB N_VPWR_c_125_n 0.0213359f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.365
cc_27 VPB N_VPWR_c_126_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_28 VPB N_VPWR_c_127_n 0.0253045f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_29 VPB N_VPWR_c_121_n 0.0651959f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_30 VPB N_Y_c_153_n 0.00881636f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_31 VPB N_Y_c_154_n 0.00807857f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_32 VPB N_Y_c_155_n 0.0557338f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_33 VPB N_Y_c_151_n 0.00301672f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_34 VPB N_Y_c_157_n 0.0165104f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_35 VPB N_Y_c_158_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_36 N_C_c_38_n N_B_c_59_n 0.0329663f $X=0.7 $Y=1.22 $X2=-0.19 $Y2=-0.245
cc_37 C N_B_c_59_n 0.00239222f $X=0.635 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_38 N_C_c_37_n N_B_c_60_n 0.0545563f $X=0.655 $Y=1.765 $X2=0 $Y2=0
cc_39 N_C_c_38_n B 0.0034981f $X=0.7 $Y=1.22 $X2=0 $Y2=0
cc_40 C B 0.0296912f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_41 N_C_c_36_n N_VPWR_c_123_n 0.00546342f $X=0.565 $Y=1.385 $X2=0 $Y2=0
cc_42 N_C_c_37_n N_VPWR_c_123_n 0.0270742f $X=0.655 $Y=1.765 $X2=0 $Y2=0
cc_43 C N_VPWR_c_123_n 0.0149317f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_44 N_C_c_37_n N_VPWR_c_125_n 0.00320971f $X=0.655 $Y=1.765 $X2=0 $Y2=0
cc_45 N_C_c_37_n N_VPWR_c_121_n 0.00458775f $X=0.655 $Y=1.765 $X2=0 $Y2=0
cc_46 N_C_c_37_n N_Y_c_154_n 0.0113732f $X=0.655 $Y=1.765 $X2=0 $Y2=0
cc_47 C N_Y_c_154_n 0.0191701f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_48 N_C_c_37_n N_Y_c_158_n 0.0207938f $X=0.655 $Y=1.765 $X2=0 $Y2=0
cc_49 N_C_c_36_n N_VGND_c_197_n 0.00199394f $X=0.565 $Y=1.385 $X2=0 $Y2=0
cc_50 N_C_c_38_n N_VGND_c_197_n 0.0151342f $X=0.7 $Y=1.22 $X2=0 $Y2=0
cc_51 C N_VGND_c_197_n 0.0259403f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_52 N_C_c_38_n N_VGND_c_200_n 0.00383152f $X=0.7 $Y=1.22 $X2=0 $Y2=0
cc_53 N_C_c_38_n N_VGND_c_201_n 0.0075725f $X=0.7 $Y=1.22 $X2=0 $Y2=0
cc_54 N_B_c_59_n N_A_c_93_n 0.0246919f $X=1.09 $Y=1.22 $X2=-0.19 $Y2=-0.245
cc_55 B N_A_c_93_n 0.00897929f $X=1.115 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_56 N_B_c_60_n N_A_c_94_n 0.0525007f $X=1.105 $Y=1.765 $X2=0 $Y2=0
cc_57 B N_A_c_94_n 4.06701e-19 $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_58 N_B_c_60_n A 0.00202352f $X=1.105 $Y=1.765 $X2=0 $Y2=0
cc_59 B A 0.0244362f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_60 N_B_c_60_n N_VPWR_c_124_n 0.00899555f $X=1.105 $Y=1.765 $X2=0 $Y2=0
cc_61 N_B_c_60_n N_VPWR_c_125_n 0.00445602f $X=1.105 $Y=1.765 $X2=0 $Y2=0
cc_62 N_B_c_60_n N_VPWR_c_121_n 0.00858056f $X=1.105 $Y=1.765 $X2=0 $Y2=0
cc_63 N_B_c_60_n N_Y_c_153_n 0.0140392f $X=1.105 $Y=1.765 $X2=0 $Y2=0
cc_64 B N_Y_c_153_n 0.0232997f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_65 N_B_c_60_n N_Y_c_154_n 0.00250598f $X=1.105 $Y=1.765 $X2=0 $Y2=0
cc_66 B N_Y_c_154_n 0.00245488f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_67 N_B_c_59_n N_Y_c_150_n 7.56255e-19 $X=1.09 $Y=1.22 $X2=0 $Y2=0
cc_68 B N_Y_c_150_n 0.0172672f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_69 N_B_c_60_n N_Y_c_155_n 9.53135e-19 $X=1.105 $Y=1.765 $X2=0 $Y2=0
cc_70 B N_Y_c_152_n 0.00754251f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_71 N_B_c_60_n N_Y_c_158_n 0.0132766f $X=1.105 $Y=1.765 $X2=0 $Y2=0
cc_72 N_B_c_59_n N_VGND_c_197_n 0.00251629f $X=1.09 $Y=1.22 $X2=0 $Y2=0
cc_73 B N_VGND_c_197_n 0.023155f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_74 N_B_c_59_n N_VGND_c_200_n 0.00304348f $X=1.09 $Y=1.22 $X2=0 $Y2=0
cc_75 B N_VGND_c_200_n 0.00930091f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_76 N_B_c_59_n N_VGND_c_201_n 0.00371612f $X=1.09 $Y=1.22 $X2=0 $Y2=0
cc_77 B N_VGND_c_201_n 0.0106938f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_78 B A_233_74# 0.00988329f $X=1.115 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_79 N_A_c_94_n N_VPWR_c_124_n 0.00868976f $X=1.675 $Y=1.765 $X2=0 $Y2=0
cc_80 N_A_c_94_n N_VPWR_c_127_n 0.00445602f $X=1.675 $Y=1.765 $X2=0 $Y2=0
cc_81 N_A_c_94_n N_VPWR_c_121_n 0.00862449f $X=1.675 $Y=1.765 $X2=0 $Y2=0
cc_82 N_A_c_94_n N_Y_c_153_n 0.0129889f $X=1.675 $Y=1.765 $X2=0 $Y2=0
cc_83 A N_Y_c_153_n 0.0123606f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_84 N_A_c_93_n N_Y_c_150_n 0.00846119f $X=1.66 $Y=1.22 $X2=0 $Y2=0
cc_85 N_A_c_94_n N_Y_c_155_n 0.0144859f $X=1.675 $Y=1.765 $X2=0 $Y2=0
cc_86 N_A_c_93_n N_Y_c_151_n 0.00394268f $X=1.66 $Y=1.22 $X2=0 $Y2=0
cc_87 N_A_c_94_n N_Y_c_151_n 0.0124478f $X=1.675 $Y=1.765 $X2=0 $Y2=0
cc_88 A N_Y_c_151_n 0.0280999f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_89 N_A_c_93_n N_Y_c_152_n 0.00296171f $X=1.66 $Y=1.22 $X2=0 $Y2=0
cc_90 N_A_c_94_n N_Y_c_152_n 0.00101144f $X=1.675 $Y=1.765 $X2=0 $Y2=0
cc_91 A N_Y_c_152_n 0.0138478f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_92 N_A_c_94_n N_Y_c_157_n 0.0049413f $X=1.675 $Y=1.765 $X2=0 $Y2=0
cc_93 A N_Y_c_157_n 0.0151534f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_94 N_A_c_94_n N_Y_c_158_n 9.35896e-19 $X=1.675 $Y=1.765 $X2=0 $Y2=0
cc_95 N_A_c_93_n N_VGND_c_200_n 0.00434272f $X=1.66 $Y=1.22 $X2=0 $Y2=0
cc_96 N_A_c_93_n N_VGND_c_201_n 0.00822158f $X=1.66 $Y=1.22 $X2=0 $Y2=0
cc_97 N_VPWR_M1004_d N_Y_c_153_n 0.0033342f $X=1.18 $Y=1.84 $X2=0 $Y2=0
cc_98 N_VPWR_c_124_n N_Y_c_153_n 0.0248957f $X=1.38 $Y=2.145 $X2=0 $Y2=0
cc_99 N_VPWR_c_123_n N_Y_c_154_n 0.00568224f $X=0.35 $Y=1.985 $X2=0 $Y2=0
cc_100 N_VPWR_c_124_n N_Y_c_155_n 0.0345826f $X=1.38 $Y=2.145 $X2=0 $Y2=0
cc_101 N_VPWR_c_127_n N_Y_c_155_n 0.0230718f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_102 N_VPWR_c_121_n N_Y_c_155_n 0.0190639f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_103 N_VPWR_c_123_n N_Y_c_158_n 0.0846658f $X=0.35 $Y=1.985 $X2=0 $Y2=0
cc_104 N_VPWR_c_124_n N_Y_c_158_n 0.0368642f $X=1.38 $Y=2.145 $X2=0 $Y2=0
cc_105 N_VPWR_c_125_n N_Y_c_158_n 0.0191315f $X=1.215 $Y=3.33 $X2=0 $Y2=0
cc_106 N_VPWR_c_121_n N_Y_c_158_n 0.0155112f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_107 N_Y_c_150_n N_VGND_c_200_n 0.0142249f $X=1.875 $Y=0.515 $X2=0 $Y2=0
cc_108 N_Y_c_150_n N_VGND_c_201_n 0.011867f $X=1.875 $Y=0.515 $X2=0 $Y2=0
cc_109 N_Y_c_152_n N_VGND_c_201_n 0.00749433f $X=2.17 $Y=0.925 $X2=0 $Y2=0
