* File: sky130_fd_sc_ls__o211ai_1.pxi.spice
* Created: Wed Sep  2 11:17:32 2020
* 
x_PM_SKY130_FD_SC_LS__O211AI_1%A1 N_A1_c_46_n N_A1_M1005_g N_A1_M1006_g A1
+ N_A1_c_48_n PM_SKY130_FD_SC_LS__O211AI_1%A1
x_PM_SKY130_FD_SC_LS__O211AI_1%A2 N_A2_c_70_n N_A2_M1000_g N_A2_M1001_g A2 A2 A2
+ A2 A2 PM_SKY130_FD_SC_LS__O211AI_1%A2
x_PM_SKY130_FD_SC_LS__O211AI_1%B1 N_B1_M1002_g N_B1_c_106_n N_B1_M1003_g B1 B1
+ B1 B1 PM_SKY130_FD_SC_LS__O211AI_1%B1
x_PM_SKY130_FD_SC_LS__O211AI_1%C1 N_C1_c_140_n N_C1_M1007_g N_C1_c_141_n
+ N_C1_M1004_g C1 PM_SKY130_FD_SC_LS__O211AI_1%C1
x_PM_SKY130_FD_SC_LS__O211AI_1%VPWR N_VPWR_M1005_s N_VPWR_M1003_d N_VPWR_c_168_n
+ N_VPWR_c_169_n N_VPWR_c_170_n N_VPWR_c_171_n N_VPWR_c_172_n VPWR
+ N_VPWR_c_173_n N_VPWR_c_167_n PM_SKY130_FD_SC_LS__O211AI_1%VPWR
x_PM_SKY130_FD_SC_LS__O211AI_1%Y N_Y_M1007_d N_Y_M1000_d N_Y_M1004_d N_Y_c_200_n
+ N_Y_c_201_n N_Y_c_202_n N_Y_c_203_n N_Y_c_198_n N_Y_c_205_n Y Y N_Y_c_199_n
+ PM_SKY130_FD_SC_LS__O211AI_1%Y
x_PM_SKY130_FD_SC_LS__O211AI_1%A_31_74# N_A_31_74#_M1006_s N_A_31_74#_M1001_d
+ N_A_31_74#_c_239_n N_A_31_74#_c_240_n N_A_31_74#_c_241_n N_A_31_74#_c_242_n
+ PM_SKY130_FD_SC_LS__O211AI_1%A_31_74#
x_PM_SKY130_FD_SC_LS__O211AI_1%VGND N_VGND_M1006_d N_VGND_c_264_n VGND
+ N_VGND_c_265_n N_VGND_c_266_n N_VGND_c_267_n N_VGND_c_268_n
+ PM_SKY130_FD_SC_LS__O211AI_1%VGND
cc_1 VNB N_A1_c_46_n 0.0609482f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_2 VNB N_A1_M1006_g 0.0310333f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=0.74
cc_3 VNB N_A1_c_48_n 0.0050357f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_4 VNB N_A2_c_70_n 0.0305436f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_5 VNB N_A2_M1001_g 0.0224026f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=0.74
cc_6 VNB A2 0.0130937f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_7 VNB A2 4.83307e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_B1_M1002_g 0.024159f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_9 VNB N_B1_c_106_n 0.030671f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=0.74
cc_10 VNB B1 0.00339768f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_11 VNB B1 0.00548062f $X=-0.19 $Y=-0.245 $X2=0.35 $Y2=1.465
cc_12 VNB N_C1_c_140_n 0.0236718f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_13 VNB N_C1_c_141_n 0.0431153f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.3
cc_14 VNB C1 0.00370468f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_VPWR_c_167_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_Y_c_198_n 0.0310722f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_Y_c_199_n 0.0239756f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_31_74#_c_239_n 0.02581f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_31_74#_c_240_n 0.00796953f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_20 VNB N_A_31_74#_c_241_n 0.00898165f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_21 VNB N_A_31_74#_c_242_n 0.00260143f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.665
cc_22 VNB N_VGND_c_264_n 0.00641543f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=0.74
cc_23 VNB N_VGND_c_265_n 0.0197879f $X=-0.19 $Y=-0.245 $X2=0.35 $Y2=1.465
cc_24 VNB N_VGND_c_266_n 0.0547577f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_267_n 0.194045f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_268_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VPB N_A1_c_46_n 0.0262772f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_28 VPB N_A1_c_48_n 0.00974946f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_29 VPB N_A2_c_70_n 0.0261842f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_30 VPB A2 0.00329681f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_31 VPB N_B1_c_106_n 0.0249238f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=0.74
cc_32 VPB N_C1_c_141_n 0.0277275f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=1.3
cc_33 VPB N_VPWR_c_168_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_34 VPB N_VPWR_c_169_n 0.0496032f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_35 VPB N_VPWR_c_170_n 0.00651803f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.665
cc_36 VPB N_VPWR_c_171_n 0.038365f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_37 VPB N_VPWR_c_172_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_38 VPB N_VPWR_c_173_n 0.0246348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_39 VPB N_VPWR_c_167_n 0.0695765f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_40 VPB N_Y_c_200_n 0.00339366f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_41 VPB N_Y_c_201_n 0.00816189f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_42 VPB N_Y_c_202_n 0.00553073f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_43 VPB N_Y_c_203_n 0.0544339f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_44 VPB N_Y_c_198_n 0.00725909f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_45 VPB N_Y_c_205_n 0.0211491f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 N_A1_c_46_n N_A2_c_70_n 0.0741905f $X=0.505 $Y=1.765 $X2=-0.19 $Y2=-0.245
cc_47 N_A1_c_48_n N_A2_c_70_n 2.46571e-19 $X=0.27 $Y=1.465 $X2=-0.19 $Y2=-0.245
cc_48 N_A1_M1006_g N_A2_M1001_g 0.0278145f $X=0.515 $Y=0.74 $X2=0 $Y2=0
cc_49 N_A1_c_46_n A2 0.00304525f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_50 N_A1_c_48_n A2 0.0230252f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_51 N_A1_c_46_n A2 0.00721826f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_52 N_A1_c_48_n A2 0.01146f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_53 N_A1_c_46_n N_VPWR_c_169_n 0.0118646f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_54 N_A1_c_48_n N_VPWR_c_169_n 0.0222392f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_55 N_A1_c_46_n N_VPWR_c_171_n 0.00461464f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_56 N_A1_c_46_n N_VPWR_c_167_n 0.00912251f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_57 N_A1_M1006_g N_A_31_74#_c_239_n 0.00968761f $X=0.515 $Y=0.74 $X2=0 $Y2=0
cc_58 N_A1_M1006_g N_A_31_74#_c_240_n 0.0152543f $X=0.515 $Y=0.74 $X2=0 $Y2=0
cc_59 N_A1_c_46_n N_A_31_74#_c_241_n 0.00265581f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_60 N_A1_M1006_g N_A_31_74#_c_241_n 0.00206782f $X=0.515 $Y=0.74 $X2=0 $Y2=0
cc_61 N_A1_c_48_n N_A_31_74#_c_241_n 0.0260039f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_62 N_A1_M1006_g N_VGND_c_264_n 0.00539757f $X=0.515 $Y=0.74 $X2=0 $Y2=0
cc_63 N_A1_M1006_g N_VGND_c_265_n 0.00434272f $X=0.515 $Y=0.74 $X2=0 $Y2=0
cc_64 N_A1_M1006_g N_VGND_c_267_n 0.00824496f $X=0.515 $Y=0.74 $X2=0 $Y2=0
cc_65 N_A2_M1001_g N_B1_M1002_g 0.0143797f $X=1.015 $Y=0.74 $X2=0 $Y2=0
cc_66 N_A2_c_70_n N_B1_c_106_n 0.0400176f $X=0.925 $Y=1.765 $X2=0 $Y2=0
cc_67 A2 N_B1_c_106_n 4.1782e-19 $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_68 N_A2_c_70_n B1 4.19259e-19 $X=0.925 $Y=1.765 $X2=0 $Y2=0
cc_69 A2 B1 0.0197279f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_70 N_A2_c_70_n N_VPWR_c_171_n 0.00461464f $X=0.925 $Y=1.765 $X2=0 $Y2=0
cc_71 A2 N_VPWR_c_171_n 0.00615262f $X=0.72 $Y=1.665 $X2=0 $Y2=0
cc_72 N_A2_c_70_n N_VPWR_c_167_n 0.00911524f $X=0.925 $Y=1.765 $X2=0 $Y2=0
cc_73 A2 N_VPWR_c_167_n 0.00794958f $X=0.72 $Y=1.665 $X2=0 $Y2=0
cc_74 A2 A_116_368# 0.0112331f $X=0.72 $Y=1.665 $X2=-0.19 $Y2=-0.245
cc_75 N_A2_c_70_n N_Y_c_200_n 0.0127786f $X=0.925 $Y=1.765 $X2=0 $Y2=0
cc_76 N_A2_c_70_n N_Y_c_202_n 0.00236795f $X=0.925 $Y=1.765 $X2=0 $Y2=0
cc_77 A2 N_Y_c_202_n 0.00338979f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_78 A2 N_Y_c_202_n 0.00627449f $X=0.72 $Y=1.665 $X2=0 $Y2=0
cc_79 N_A2_M1001_g N_A_31_74#_c_239_n 9.1183e-19 $X=1.015 $Y=0.74 $X2=0 $Y2=0
cc_80 N_A2_c_70_n N_A_31_74#_c_240_n 0.00127493f $X=0.925 $Y=1.765 $X2=0 $Y2=0
cc_81 N_A2_M1001_g N_A_31_74#_c_240_n 0.0128142f $X=1.015 $Y=0.74 $X2=0 $Y2=0
cc_82 A2 N_A_31_74#_c_240_n 0.041574f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_83 N_A2_M1001_g N_A_31_74#_c_242_n 4.33993e-19 $X=1.015 $Y=0.74 $X2=0 $Y2=0
cc_84 N_A2_M1001_g N_VGND_c_264_n 0.00956268f $X=1.015 $Y=0.74 $X2=0 $Y2=0
cc_85 N_A2_M1001_g N_VGND_c_266_n 0.00383152f $X=1.015 $Y=0.74 $X2=0 $Y2=0
cc_86 N_A2_M1001_g N_VGND_c_267_n 0.00757954f $X=1.015 $Y=0.74 $X2=0 $Y2=0
cc_87 N_B1_M1002_g N_C1_c_140_n 0.0233562f $X=1.48 $Y=0.74 $X2=-0.19 $Y2=-0.245
cc_88 B1 N_C1_c_140_n 0.00938955f $X=1.595 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_89 N_B1_c_106_n N_C1_c_141_n 0.0505679f $X=1.645 $Y=1.765 $X2=0 $Y2=0
cc_90 B1 N_C1_c_141_n 0.00330338f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_91 N_B1_c_106_n C1 2.81336e-19 $X=1.645 $Y=1.765 $X2=0 $Y2=0
cc_92 B1 C1 0.00880658f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_93 B1 C1 0.0192202f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_94 N_B1_c_106_n N_VPWR_c_170_n 0.0182161f $X=1.645 $Y=1.765 $X2=0 $Y2=0
cc_95 N_B1_c_106_n N_VPWR_c_171_n 0.00413917f $X=1.645 $Y=1.765 $X2=0 $Y2=0
cc_96 N_B1_c_106_n N_VPWR_c_167_n 0.00819732f $X=1.645 $Y=1.765 $X2=0 $Y2=0
cc_97 N_B1_c_106_n N_Y_c_200_n 0.0138629f $X=1.645 $Y=1.765 $X2=0 $Y2=0
cc_98 N_B1_c_106_n N_Y_c_201_n 0.0193702f $X=1.645 $Y=1.765 $X2=0 $Y2=0
cc_99 B1 N_Y_c_201_n 0.0252014f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_100 N_B1_c_106_n N_Y_c_202_n 0.00136199f $X=1.645 $Y=1.765 $X2=0 $Y2=0
cc_101 B1 N_Y_c_202_n 0.00421666f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_102 N_B1_c_106_n N_Y_c_203_n 9.66739e-19 $X=1.645 $Y=1.765 $X2=0 $Y2=0
cc_103 B1 N_Y_c_199_n 0.0338432f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_104 B1 N_A_31_74#_c_240_n 0.0016373f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_105 N_B1_M1002_g N_A_31_74#_c_242_n 8.38786e-19 $X=1.48 $Y=0.74 $X2=0 $Y2=0
cc_106 N_B1_M1002_g N_VGND_c_264_n 6.58032e-19 $X=1.48 $Y=0.74 $X2=0 $Y2=0
cc_107 N_B1_M1002_g N_VGND_c_266_n 0.00461464f $X=1.48 $Y=0.74 $X2=0 $Y2=0
cc_108 B1 N_VGND_c_266_n 0.00653424f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_109 N_B1_M1002_g N_VGND_c_267_n 0.00910985f $X=1.48 $Y=0.74 $X2=0 $Y2=0
cc_110 B1 N_VGND_c_267_n 0.00794958f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_111 B1 A_311_74# 0.0161056f $X=1.595 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_112 N_C1_c_141_n N_VPWR_c_170_n 0.00766779f $X=2.145 $Y=1.765 $X2=0 $Y2=0
cc_113 N_C1_c_141_n N_VPWR_c_173_n 0.00445602f $X=2.145 $Y=1.765 $X2=0 $Y2=0
cc_114 N_C1_c_141_n N_VPWR_c_167_n 0.00861477f $X=2.145 $Y=1.765 $X2=0 $Y2=0
cc_115 N_C1_c_141_n N_Y_c_201_n 0.0136234f $X=2.145 $Y=1.765 $X2=0 $Y2=0
cc_116 C1 N_Y_c_201_n 0.0125099f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_117 N_C1_c_141_n N_Y_c_203_n 0.0130597f $X=2.145 $Y=1.765 $X2=0 $Y2=0
cc_118 N_C1_c_140_n N_Y_c_198_n 0.00339074f $X=2.05 $Y=1.22 $X2=0 $Y2=0
cc_119 N_C1_c_141_n N_Y_c_198_n 0.0139137f $X=2.145 $Y=1.765 $X2=0 $Y2=0
cc_120 C1 N_Y_c_198_n 0.0188818f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_121 N_C1_c_141_n N_Y_c_205_n 0.00239008f $X=2.145 $Y=1.765 $X2=0 $Y2=0
cc_122 C1 N_Y_c_205_n 0.00626023f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_123 N_C1_c_140_n N_Y_c_199_n 0.0112973f $X=2.05 $Y=1.22 $X2=0 $Y2=0
cc_124 N_C1_c_141_n N_Y_c_199_n 0.00108361f $X=2.145 $Y=1.765 $X2=0 $Y2=0
cc_125 C1 N_Y_c_199_n 0.0192616f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_126 N_C1_c_140_n N_VGND_c_266_n 0.00377174f $X=2.05 $Y=1.22 $X2=0 $Y2=0
cc_127 N_C1_c_140_n N_VGND_c_267_n 0.00628921f $X=2.05 $Y=1.22 $X2=0 $Y2=0
cc_128 N_VPWR_c_170_n N_Y_c_200_n 0.0485394f $X=1.87 $Y=2.305 $X2=0 $Y2=0
cc_129 N_VPWR_c_171_n N_Y_c_200_n 0.0146357f $X=1.705 $Y=3.33 $X2=0 $Y2=0
cc_130 N_VPWR_c_167_n N_Y_c_200_n 0.0121141f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_131 N_VPWR_M1003_d N_Y_c_201_n 0.00250873f $X=1.72 $Y=1.84 $X2=0 $Y2=0
cc_132 N_VPWR_c_170_n N_Y_c_201_n 0.0202249f $X=1.87 $Y=2.305 $X2=0 $Y2=0
cc_133 N_VPWR_c_170_n N_Y_c_203_n 0.0350101f $X=1.87 $Y=2.305 $X2=0 $Y2=0
cc_134 N_VPWR_c_173_n N_Y_c_203_n 0.0250797f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_135 N_VPWR_c_167_n N_Y_c_203_n 0.0207259f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_136 N_Y_c_202_n N_A_31_74#_c_240_n 0.00821726f $X=1.455 $Y=1.885 $X2=0 $Y2=0
cc_137 N_Y_c_199_n N_VGND_c_266_n 0.0216534f $X=2.682 $Y=0.725 $X2=0 $Y2=0
cc_138 N_Y_c_199_n N_VGND_c_267_n 0.0246737f $X=2.682 $Y=0.725 $X2=0 $Y2=0
cc_139 N_A_31_74#_c_240_n N_VGND_M1006_d 0.00256964f $X=1.145 $Y=1.045 $X2=-0.19
+ $Y2=-0.245
cc_140 N_A_31_74#_c_239_n N_VGND_c_264_n 0.0169251f $X=0.3 $Y=0.515 $X2=0 $Y2=0
cc_141 N_A_31_74#_c_240_n N_VGND_c_264_n 0.0201026f $X=1.145 $Y=1.045 $X2=0
+ $Y2=0
cc_142 N_A_31_74#_c_242_n N_VGND_c_264_n 0.0161397f $X=1.23 $Y=0.515 $X2=0 $Y2=0
cc_143 N_A_31_74#_c_239_n N_VGND_c_265_n 0.0145639f $X=0.3 $Y=0.515 $X2=0 $Y2=0
cc_144 N_A_31_74#_c_242_n N_VGND_c_266_n 0.011066f $X=1.23 $Y=0.515 $X2=0 $Y2=0
cc_145 N_A_31_74#_c_239_n N_VGND_c_267_n 0.0119984f $X=0.3 $Y=0.515 $X2=0 $Y2=0
cc_146 N_A_31_74#_c_242_n N_VGND_c_267_n 0.00915947f $X=1.23 $Y=0.515 $X2=0
+ $Y2=0
