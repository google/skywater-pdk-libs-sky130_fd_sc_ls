* File: sky130_fd_sc_ls__o311a_4.pex.spice
* Created: Wed Sep  2 11:21:27 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__O311A_4%A_83_244# 1 2 3 4 13 15 16 18 19 21 22 24 25
+ 27 28 30 31 33 34 36 37 42 43 44 45 48 50 54 56 58 61 64 65 71 73 77
c189 64 0 1.56729e-19 $X=2.1 $Y=1.385
c190 50 0 9.98244e-21 $X=4.09 $Y=2.035
c191 22 0 4.74979e-20 $X=0.995 $Y=1.22
c192 13 0 4.66086e-20 $X=0.505 $Y=1.765
r193 86 87 46.6828 $w=4.13e-07 $l=4e-07 $layer=POLY_cond $X=1.69 $Y=1.492
+ $X2=2.09 $Y2=1.492
r194 85 86 27.4261 $w=4.13e-07 $l=2.35e-07 $layer=POLY_cond $X=1.455 $Y=1.492
+ $X2=1.69 $Y2=1.492
r195 82 83 4.66828 $w=4.13e-07 $l=4e-08 $layer=POLY_cond $X=0.955 $Y=1.492
+ $X2=0.995 $Y2=1.492
r196 81 82 45.5157 $w=4.13e-07 $l=3.9e-07 $layer=POLY_cond $X=0.565 $Y=1.492
+ $X2=0.955 $Y2=1.492
r197 80 81 7.00242 $w=4.13e-07 $l=6e-08 $layer=POLY_cond $X=0.505 $Y=1.492
+ $X2=0.565 $Y2=1.492
r198 77 79 16.7345 $w=2.26e-07 $l=3.1e-07 $layer=LI1_cond $X=5.615 $Y=2.075
+ $X2=5.925 $Y2=2.075
r199 73 75 5.30124 $w=2.48e-07 $l=1.15e-07 $layer=LI1_cond $X=4.46 $Y=1.1
+ $X2=4.46 $Y2=1.215
r200 67 69 2.44458 $w=3.28e-07 $l=7e-08 $layer=LI1_cond $X=2.82 $Y=2.035
+ $X2=2.82 $Y2=2.105
r201 65 67 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=2.82 $Y=1.805
+ $X2=2.82 $Y2=2.035
r202 64 89 10.5036 $w=4.13e-07 $l=9e-08 $layer=POLY_cond $X=2.1 $Y=1.492
+ $X2=2.19 $Y2=1.492
r203 64 87 1.16707 $w=4.13e-07 $l=1e-08 $layer=POLY_cond $X=2.1 $Y=1.492
+ $X2=2.09 $Y2=1.492
r204 63 64 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.1
+ $Y=1.385 $X2=2.1 $Y2=1.385
r205 61 77 2.4068 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.615 $Y=1.95
+ $X2=5.615 $Y2=2.075
r206 60 61 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=5.615 $Y=1.3
+ $X2=5.615 $Y2=1.95
r207 59 75 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.585 $Y=1.215
+ $X2=4.46 $Y2=1.215
r208 58 60 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.53 $Y=1.215
+ $X2=5.615 $Y2=1.3
r209 58 59 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=5.53 $Y=1.215
+ $X2=4.585 $Y2=1.215
r210 57 71 8.61065 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=4.42 $Y=2.055
+ $X2=4.255 $Y2=2.04
r211 56 77 5.36542 $w=2.26e-07 $l=9.44722e-08 $layer=LI1_cond $X=5.53 $Y=2.055
+ $X2=5.615 $Y2=2.075
r212 56 57 72.4171 $w=1.68e-07 $l=1.11e-06 $layer=LI1_cond $X=5.53 $Y=2.055
+ $X2=4.42 $Y2=2.055
r213 52 71 0.89609 $w=3.3e-07 $l=1e-07 $layer=LI1_cond $X=4.255 $Y=2.14
+ $X2=4.255 $Y2=2.04
r214 52 54 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=4.255 $Y=2.14
+ $X2=4.255 $Y2=2.815
r215 51 67 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.985 $Y=2.035
+ $X2=2.82 $Y2=2.035
r216 50 71 8.61065 $w=1.7e-07 $l=1.67481e-07 $layer=LI1_cond $X=4.09 $Y=2.035
+ $X2=4.255 $Y2=2.04
r217 50 51 72.0909 $w=1.68e-07 $l=1.105e-06 $layer=LI1_cond $X=4.09 $Y=2.035
+ $X2=2.985 $Y2=2.035
r218 46 69 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=2.82 $Y=2.12
+ $X2=2.82 $Y2=2.105
r219 46 48 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=2.82 $Y=2.12
+ $X2=2.82 $Y2=2.815
r220 44 65 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.655 $Y=1.805
+ $X2=2.82 $Y2=1.805
r221 44 45 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=2.655 $Y=1.805
+ $X2=2.265 $Y2=1.805
r222 43 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.18 $Y=1.72
+ $X2=2.265 $Y2=1.805
r223 42 63 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.18 $Y=1.55
+ $X2=2.18 $Y2=1.385
r224 42 43 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.18 $Y=1.55
+ $X2=2.18 $Y2=1.72
r225 40 85 4.08475 $w=4.13e-07 $l=3.5e-08 $layer=POLY_cond $X=1.42 $Y=1.492
+ $X2=1.455 $Y2=1.492
r226 40 83 49.6005 $w=4.13e-07 $l=4.25e-07 $layer=POLY_cond $X=1.42 $Y=1.492
+ $X2=0.995 $Y2=1.492
r227 39 40 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.42
+ $Y=1.385 $X2=1.42 $Y2=1.385
r228 37 63 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.095 $Y=1.385
+ $X2=2.18 $Y2=1.385
r229 37 39 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.095 $Y=1.385
+ $X2=1.42 $Y2=1.385
r230 34 89 26.6457 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=2.19 $Y=1.22
+ $X2=2.19 $Y2=1.492
r231 34 36 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.19 $Y=1.22
+ $X2=2.19 $Y2=0.74
r232 31 87 26.6457 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=2.09 $Y=1.765
+ $X2=2.09 $Y2=1.492
r233 31 33 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.09 $Y=1.765
+ $X2=2.09 $Y2=2.4
r234 28 86 26.6457 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=1.69 $Y=1.22
+ $X2=1.69 $Y2=1.492
r235 28 30 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.69 $Y=1.22
+ $X2=1.69 $Y2=0.74
r236 25 85 26.6457 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=1.455 $Y=1.765
+ $X2=1.455 $Y2=1.492
r237 25 27 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.455 $Y=1.765
+ $X2=1.455 $Y2=2.4
r238 22 83 26.6457 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=0.995 $Y=1.22
+ $X2=0.995 $Y2=1.492
r239 22 24 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.995 $Y=1.22
+ $X2=0.995 $Y2=0.74
r240 19 82 26.6457 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=0.955 $Y=1.765
+ $X2=0.955 $Y2=1.492
r241 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.955 $Y=1.765
+ $X2=0.955 $Y2=2.4
r242 16 81 26.6457 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=0.565 $Y=1.22
+ $X2=0.565 $Y2=1.492
r243 16 18 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.565 $Y=1.22
+ $X2=0.565 $Y2=0.74
r244 13 80 26.6457 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=1.492
r245 13 15 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.4
r246 4 79 600 $w=1.7e-07 $l=2.24499e-07 $layer=licon1_PDIFF $count=1 $X=5.765
+ $Y=1.96 $X2=5.925 $Y2=2.115
r247 3 71 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=4.105
+ $Y=1.96 $X2=4.255 $Y2=2.105
r248 3 54 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=4.105
+ $Y=1.96 $X2=4.255 $Y2=2.815
r249 2 69 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.67
+ $Y=1.96 $X2=2.82 $Y2=2.105
r250 2 48 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=2.67
+ $Y=1.96 $X2=2.82 $Y2=2.815
r251 1 73 182 $w=1.7e-07 $l=8.12588e-07 $layer=licon1_NDIFF $count=1 $X=4.2
+ $Y=0.39 $X2=4.42 $Y2=1.1
.ends

.subckt PM_SKY130_FD_SC_LS__O311A_4%B1 2 3 5 6 10 12 14 15 16 19 21 22 24 26 31
+ 33 38 39 44
c110 24 0 1.03664e-19 $X=4.08 $Y=1.47
c111 3 0 9.98244e-21 $X=2.595 $Y=1.885
r112 38 41 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=5.195 $Y=1.635
+ $X2=5.195 $Y2=1.785
r113 38 40 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.195 $Y=1.635
+ $X2=5.195 $Y2=1.47
r114 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.195
+ $Y=1.635 $X2=5.195 $Y2=1.635
r115 31 39 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=5.04 $Y=1.635
+ $X2=5.195 $Y2=1.635
r116 31 44 6.71605 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=5.04 $Y=1.635
+ $X2=4.925 $Y2=1.635
r117 30 36 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.67 $Y=1.385
+ $X2=2.67 $Y2=1.55
r118 30 33 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.67 $Y=1.385
+ $X2=2.67 $Y2=1.295
r119 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.67
+ $Y=1.385 $X2=2.67 $Y2=1.385
r120 26 44 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=4.165 $Y=1.555
+ $X2=4.925 $Y2=1.555
r121 24 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.08 $Y=1.47
+ $X2=4.165 $Y2=1.555
r122 23 24 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=4.08 $Y=1.265
+ $X2=4.08 $Y2=1.47
r123 22 29 7.35588 $w=3.4e-07 $l=2.89206e-07 $layer=LI1_cond $X=2.91 $Y=1.18
+ $X2=2.707 $Y2=1.385
r124 21 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.995 $Y=1.18
+ $X2=4.08 $Y2=1.265
r125 21 22 70.7861 $w=1.68e-07 $l=1.085e-06 $layer=LI1_cond $X=3.995 $Y=1.18
+ $X2=2.91 $Y2=1.18
r126 19 40 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=5.145 $Y=0.71
+ $X2=5.145 $Y2=1.47
r127 15 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.03 $Y=1.785
+ $X2=5.195 $Y2=1.785
r128 15 16 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=5.03 $Y=1.785
+ $X2=4.62 $Y2=1.785
r129 12 16 26.9307 $w=1.5e-07 $l=1.3784e-07 $layer=POLY_cond $X=4.53 $Y=1.885
+ $X2=4.62 $Y2=1.785
r130 12 14 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=4.53 $Y=1.885
+ $X2=4.53 $Y2=2.46
r131 8 10 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=3.18 $Y=1.22
+ $X2=3.18 $Y2=0.71
r132 7 33 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.835 $Y=1.295
+ $X2=2.67 $Y2=1.295
r133 6 8 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.105 $Y=1.295
+ $X2=3.18 $Y2=1.22
r134 6 7 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=3.105 $Y=1.295
+ $X2=2.835 $Y2=1.295
r135 3 5 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.595 $Y=1.885
+ $X2=2.595 $Y2=2.46
r136 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.595 $Y=1.795
+ $X2=2.595 $Y2=1.885
r137 2 36 95.2339 $w=1.8e-07 $l=2.45e-07 $layer=POLY_cond $X=2.595 $Y=1.795
+ $X2=2.595 $Y2=1.55
.ends

.subckt PM_SKY130_FD_SC_LS__O311A_4%C1 1 3 4 6 8 11 13 14 17 19 21
c73 17 0 1.03664e-19 $X=4.715 $Y=0.71
r74 26 27 9.64 $w=4.75e-07 $l=9.5e-08 $layer=POLY_cond $X=4.03 $Y=1.602
+ $X2=4.125 $Y2=1.602
r75 24 26 37.5453 $w=4.75e-07 $l=3.7e-07 $layer=POLY_cond $X=3.66 $Y=1.602
+ $X2=4.03 $Y2=1.602
r76 21 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.66
+ $Y=1.6 $X2=3.66 $Y2=1.6
r77 15 17 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.715 $Y=1.32
+ $X2=4.715 $Y2=0.71
r78 14 27 32.1576 $w=4.75e-07 $l=2.41607e-07 $layer=POLY_cond $X=4.2 $Y=1.395
+ $X2=4.125 $Y2=1.602
r79 13 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.64 $Y=1.395
+ $X2=4.715 $Y2=1.32
r80 13 14 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=4.64 $Y=1.395
+ $X2=4.2 $Y2=1.395
r81 9 27 30.117 $w=1.5e-07 $l=2.82e-07 $layer=POLY_cond $X=4.125 $Y=1.32
+ $X2=4.125 $Y2=1.602
r82 9 11 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.125 $Y=1.32
+ $X2=4.125 $Y2=0.71
r83 6 26 30.117 $w=1.5e-07 $l=2.83e-07 $layer=POLY_cond $X=4.03 $Y=1.885
+ $X2=4.03 $Y2=1.602
r84 6 8 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=4.03 $Y=1.885
+ $X2=4.03 $Y2=2.46
r85 5 19 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.255 $Y=1.69 $X2=3.165
+ $Y2=1.69
r86 4 24 41.2902 $w=4.75e-07 $l=2.04316e-07 $layer=POLY_cond $X=3.495 $Y=1.69
+ $X2=3.66 $Y2=1.602
r87 4 5 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=3.495 $Y=1.69
+ $X2=3.255 $Y2=1.69
r88 1 19 77.9482 $w=1.8e-07 $l=1.95e-07 $layer=POLY_cond $X=3.165 $Y=1.885
+ $X2=3.165 $Y2=1.69
r89 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.165 $Y=1.885
+ $X2=3.165 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_LS__O311A_4%A3 3 5 7 8 10 13 15 22
c59 15 0 1.46209e-19 $X=6 $Y=1.665
r60 22 23 6.16368 $w=3.91e-07 $l=5e-08 $layer=POLY_cond $X=6.16 $Y=1.652
+ $X2=6.21 $Y2=1.652
r61 20 22 15.4092 $w=3.91e-07 $l=1.25e-07 $layer=POLY_cond $X=6.035 $Y=1.652
+ $X2=6.16 $Y2=1.652
r62 18 20 42.5294 $w=3.91e-07 $l=3.45e-07 $layer=POLY_cond $X=5.69 $Y=1.652
+ $X2=6.035 $Y2=1.652
r63 17 18 1.8491 $w=3.91e-07 $l=1.5e-08 $layer=POLY_cond $X=5.675 $Y=1.652
+ $X2=5.69 $Y2=1.652
r64 15 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.035
+ $Y=1.585 $X2=6.035 $Y2=1.585
r65 11 23 25.3065 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=6.21 $Y=1.42
+ $X2=6.21 $Y2=1.652
r66 11 13 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=6.21 $Y=1.42
+ $X2=6.21 $Y2=0.71
r67 8 22 25.3065 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=6.16 $Y=1.885
+ $X2=6.16 $Y2=1.652
r68 8 10 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.16 $Y=1.885
+ $X2=6.16 $Y2=2.46
r69 5 18 25.3065 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=5.69 $Y=1.885
+ $X2=5.69 $Y2=1.652
r70 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.69 $Y=1.885
+ $X2=5.69 $Y2=2.46
r71 1 17 25.3065 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=5.675 $Y=1.42
+ $X2=5.675 $Y2=1.652
r72 1 3 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=5.675 $Y=1.42
+ $X2=5.675 $Y2=0.71
.ends

.subckt PM_SKY130_FD_SC_LS__O311A_4%A2 2 3 5 8 11 12 14 15 17 18 19 23 24 25 33
+ 37
c79 23 0 2.29863e-19 $X=6.69 $Y=1.385
r80 33 35 31.7105 $w=3.42e-07 $l=2.25e-07 $layer=POLY_cond $X=8.145 $Y=1.35
+ $X2=8.37 $Y2=1.35
r81 32 33 5.63743 $w=3.42e-07 $l=4e-08 $layer=POLY_cond $X=8.105 $Y=1.35
+ $X2=8.145 $Y2=1.35
r82 24 37 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.37 $Y=1.215 $X2=8.37
+ $Y2=1.3
r83 24 25 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=8.37 $Y=1.305
+ $X2=8.37 $Y2=1.665
r84 24 37 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=8.37 $Y=1.305
+ $X2=8.37 $Y2=1.3
r85 24 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.37
+ $Y=1.305 $X2=8.37 $Y2=1.305
r86 23 31 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.69 $Y=1.385
+ $X2=6.69 $Y2=1.55
r87 23 30 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.69 $Y=1.385
+ $X2=6.69 $Y2=1.22
r88 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.69
+ $Y=1.385 $X2=6.69 $Y2=1.385
r89 19 22 5.7933 $w=3.58e-07 $l=2.77263e-07 $layer=LI1_cond $X=6.935 $Y=1.215
+ $X2=6.73 $Y2=1.385
r90 18 24 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.205 $Y=1.215
+ $X2=8.37 $Y2=1.215
r91 18 19 82.8556 $w=1.68e-07 $l=1.27e-06 $layer=LI1_cond $X=8.205 $Y=1.215
+ $X2=6.935 $Y2=1.215
r92 15 33 22.0749 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=8.145 $Y=1.14
+ $X2=8.145 $Y2=1.35
r93 15 17 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=8.145 $Y=1.14
+ $X2=8.145 $Y2=0.71
r94 12 14 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=8.105 $Y=1.885
+ $X2=8.105 $Y2=2.46
r95 11 12 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=8.105 $Y=1.795
+ $X2=8.105 $Y2=1.885
r96 10 32 17.7656 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=8.105 $Y=1.56
+ $X2=8.105 $Y2=1.35
r97 10 11 91.3468 $w=1.8e-07 $l=2.35e-07 $layer=POLY_cond $X=8.105 $Y=1.56
+ $X2=8.105 $Y2=1.795
r98 8 30 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=6.645 $Y=0.71
+ $X2=6.645 $Y2=1.22
r99 3 5 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.615 $Y=1.885
+ $X2=6.615 $Y2=2.46
r100 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.615 $Y=1.795
+ $X2=6.615 $Y2=1.885
r101 2 31 95.2339 $w=1.8e-07 $l=2.45e-07 $layer=POLY_cond $X=6.615 $Y=1.795
+ $X2=6.615 $Y2=1.55
.ends

.subckt PM_SKY130_FD_SC_LS__O311A_4%A1 3 5 7 8 10 13 15 16 24
c58 16 0 8.3654e-20 $X=7.92 $Y=1.665
r59 24 25 8.35467 $w=3.75e-07 $l=6.5e-08 $layer=POLY_cond $X=7.635 $Y=1.677
+ $X2=7.7 $Y2=1.677
r60 22 24 3.21333 $w=3.75e-07 $l=2.5e-08 $layer=POLY_cond $X=7.61 $Y=1.677
+ $X2=7.635 $Y2=1.677
r61 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.61
+ $Y=1.635 $X2=7.61 $Y2=1.635
r62 20 22 54.6267 $w=3.75e-07 $l=4.25e-07 $layer=POLY_cond $X=7.185 $Y=1.677
+ $X2=7.61 $Y2=1.677
r63 19 20 1.928 $w=3.75e-07 $l=1.5e-08 $layer=POLY_cond $X=7.17 $Y=1.677
+ $X2=7.185 $Y2=1.677
r64 16 23 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=7.92 $Y=1.635
+ $X2=7.61 $Y2=1.635
r65 15 23 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=7.44 $Y=1.635
+ $X2=7.61 $Y2=1.635
r66 11 25 24.2915 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.7 $Y=1.47 $X2=7.7
+ $Y2=1.677
r67 11 13 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=7.7 $Y=1.47 $X2=7.7
+ $Y2=0.71
r68 8 24 24.2915 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=7.635 $Y=1.885
+ $X2=7.635 $Y2=1.677
r69 8 10 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=7.635 $Y=1.885
+ $X2=7.635 $Y2=2.46
r70 5 20 24.2915 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=7.185 $Y=1.885
+ $X2=7.185 $Y2=1.677
r71 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=7.185 $Y=1.885
+ $X2=7.185 $Y2=2.46
r72 1 19 24.2915 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.17 $Y=1.47
+ $X2=7.17 $Y2=1.677
r73 1 3 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=7.17 $Y=1.47 $X2=7.17
+ $Y2=0.71
.ends

.subckt PM_SKY130_FD_SC_LS__O311A_4%VPWR 1 2 3 4 5 6 19 21 27 31 35 41 43 44 49
+ 54 55 56 57 58 60 65 78 79 85 88 91
r127 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r128 88 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r129 86 89 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r130 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r131 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r132 78 79 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r133 76 79 0.936549 $w=4.9e-07 $l=3.36e-06 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=8.4 $Y2=3.33
r134 75 78 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=5.04 $Y=3.33
+ $X2=8.4 $Y2=3.33
r135 75 76 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r136 73 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r137 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r138 70 91 13.6095 $w=1.7e-07 $l=3.48e-07 $layer=LI1_cond $X=3.92 $Y=3.33
+ $X2=3.572 $Y2=3.33
r139 70 72 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=3.92 $Y=3.33
+ $X2=4.56 $Y2=3.33
r140 69 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r141 69 89 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.16 $Y2=3.33
r142 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r143 66 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.48 $Y=3.33
+ $X2=2.315 $Y2=3.33
r144 66 68 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=2.48 $Y=3.33
+ $X2=3.12 $Y2=3.33
r145 65 91 13.6095 $w=1.7e-07 $l=3.47e-07 $layer=LI1_cond $X=3.225 $Y=3.33
+ $X2=3.572 $Y2=3.33
r146 65 68 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=3.225 $Y=3.33
+ $X2=3.12 $Y2=3.33
r147 64 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r148 64 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r149 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r150 61 82 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.182 $Y2=3.33
r151 61 63 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.72 $Y2=3.33
r152 60 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.065 $Y=3.33
+ $X2=1.23 $Y2=3.33
r153 60 63 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.065 $Y=3.33
+ $X2=0.72 $Y2=3.33
r154 58 73 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=3.33
+ $X2=4.56 $Y2=3.33
r155 58 92 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=4.32 $Y=3.33
+ $X2=3.6 $Y2=3.33
r156 56 57 8.89604 $w=4.23e-07 $l=1.7e-07 $layer=LI1_cond $X=6.38 $Y=2.255
+ $X2=6.55 $Y2=2.255
r157 54 72 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=4.59 $Y=3.33 $X2=4.56
+ $Y2=3.33
r158 54 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.59 $Y=3.33
+ $X2=4.755 $Y2=3.33
r159 53 75 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=4.92 $Y=3.33
+ $X2=5.04 $Y2=3.33
r160 53 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.92 $Y=3.33
+ $X2=4.755 $Y2=3.33
r161 49 57 23.32 $w=4.23e-07 $l=8.6e-07 $layer=LI1_cond $X=7.41 $Y=2.182
+ $X2=6.55 $Y2=2.182
r162 46 52 4.88517 $w=1.7e-07 $l=1.79374e-07 $layer=LI1_cond $X=4.92 $Y=2.455
+ $X2=4.755 $Y2=2.425
r163 46 56 95.2513 $w=1.68e-07 $l=1.46e-06 $layer=LI1_cond $X=4.92 $Y=2.455
+ $X2=6.38 $Y2=2.455
r164 44 55 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.755 $Y=3.245
+ $X2=4.755 $Y2=3.33
r165 43 52 2.881 $w=3.3e-07 $l=1.15e-07 $layer=LI1_cond $X=4.755 $Y=2.54
+ $X2=4.755 $Y2=2.425
r166 43 44 24.6204 $w=3.28e-07 $l=7.05e-07 $layer=LI1_cond $X=4.755 $Y=2.54
+ $X2=4.755 $Y2=3.245
r167 39 91 2.84707 $w=6.95e-07 $l=8.5e-08 $layer=LI1_cond $X=3.572 $Y=3.245
+ $X2=3.572 $Y2=3.33
r168 39 41 13.5957 $w=6.93e-07 $l=7.9e-07 $layer=LI1_cond $X=3.572 $Y=3.245
+ $X2=3.572 $Y2=2.455
r169 35 38 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=2.315 $Y=2.145
+ $X2=2.315 $Y2=2.825
r170 33 88 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.315 $Y=3.245
+ $X2=2.315 $Y2=3.33
r171 33 38 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=2.315 $Y=3.245
+ $X2=2.315 $Y2=2.825
r172 32 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.395 $Y=3.33
+ $X2=1.23 $Y2=3.33
r173 31 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.15 $Y=3.33
+ $X2=2.315 $Y2=3.33
r174 31 32 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=2.15 $Y=3.33
+ $X2=1.395 $Y2=3.33
r175 27 30 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.23 $Y=2.145
+ $X2=1.23 $Y2=2.825
r176 25 85 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.23 $Y=3.245
+ $X2=1.23 $Y2=3.33
r177 25 30 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=1.23 $Y=3.245
+ $X2=1.23 $Y2=2.825
r178 21 24 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=0.24 $Y=1.985
+ $X2=0.24 $Y2=2.815
r179 19 82 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.182 $Y2=3.33
r180 19 24 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.24 $Y2=2.815
r181 6 49 600 $w=1.7e-07 $l=2.85307e-07 $layer=licon1_PDIFF $count=1 $X=7.26
+ $Y=1.96 $X2=7.41 $Y2=2.18
r182 5 52 300 $w=1.7e-07 $l=5.85214e-07 $layer=licon1_PDIFF $count=2 $X=4.605
+ $Y=1.96 $X2=4.755 $Y2=2.475
r183 4 41 150 $w=1.7e-07 $l=7.73886e-07 $layer=licon1_PDIFF $count=4 $X=3.24
+ $Y=1.96 $X2=3.805 $Y2=2.455
r184 3 38 400 $w=1.7e-07 $l=1.05734e-06 $layer=licon1_PDIFF $count=1 $X=2.165
+ $Y=1.84 $X2=2.315 $Y2=2.825
r185 3 35 400 $w=1.7e-07 $l=3.72525e-07 $layer=licon1_PDIFF $count=1 $X=2.165
+ $Y=1.84 $X2=2.315 $Y2=2.145
r186 2 30 400 $w=1.7e-07 $l=1.08038e-06 $layer=licon1_PDIFF $count=1 $X=1.03
+ $Y=1.84 $X2=1.23 $Y2=2.825
r187 2 27 400 $w=1.7e-07 $l=3.9246e-07 $layer=licon1_PDIFF $count=1 $X=1.03
+ $Y=1.84 $X2=1.23 $Y2=2.145
r188 1 24 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r189 1 21 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_LS__O311A_4%X 1 2 3 4 13 15 16 19 25 27 29 33 39 42 45
+ 48 51
c69 27 0 4.66086e-20 $X=1.565 $Y=1.805
c70 13 0 4.74979e-20 $X=0.615 $Y=1.225
r71 48 51 2.9826 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.24 $Y=1.225 $X2=0.24
+ $Y2=1.31
r72 48 51 1.75372 $w=2.28e-07 $l=3.5e-08 $layer=LI1_cond $X=0.24 $Y=1.345
+ $X2=0.24 $Y2=1.31
r73 45 46 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=0.78 $Y=0.965
+ $X2=0.78 $Y2=1.225
r74 42 44 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=0.73 $Y=1.565
+ $X2=0.73 $Y2=1.805
r75 41 48 6.76434 $w=2.28e-07 $l=1.35e-07 $layer=LI1_cond $X=0.24 $Y=1.48
+ $X2=0.24 $Y2=1.345
r76 37 39 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=1.905 $Y=0.88
+ $X2=1.905 $Y2=0.515
r77 33 35 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=1.73 $Y=1.985
+ $X2=1.73 $Y2=2.815
r78 31 33 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=1.73 $Y=1.89
+ $X2=1.73 $Y2=1.985
r79 30 45 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=0.965
+ $X2=0.78 $Y2=0.965
r80 29 37 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.74 $Y=0.965
+ $X2=1.905 $Y2=0.88
r81 29 30 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=1.74 $Y=0.965
+ $X2=0.945 $Y2=0.965
r82 28 44 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=1.805
+ $X2=0.73 $Y2=1.805
r83 27 31 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.565 $Y=1.805
+ $X2=1.73 $Y2=1.89
r84 27 28 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.565 $Y=1.805
+ $X2=0.895 $Y2=1.805
r85 23 45 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=0.88
+ $X2=0.78 $Y2=0.965
r86 23 25 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=0.78 $Y=0.88
+ $X2=0.78 $Y2=0.515
r87 19 21 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=0.73 $Y=1.985
+ $X2=0.73 $Y2=2.815
r88 17 44 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=1.89
+ $X2=0.73 $Y2=1.805
r89 17 19 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=0.73 $Y=1.89
+ $X2=0.73 $Y2=1.985
r90 16 41 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.355 $Y=1.565
+ $X2=0.24 $Y2=1.48
r91 15 42 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.565 $Y=1.565
+ $X2=0.73 $Y2=1.565
r92 15 16 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=0.565 $Y=1.565
+ $X2=0.355 $Y2=1.565
r93 14 48 4.03528 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=0.355 $Y=1.225
+ $X2=0.24 $Y2=1.225
r94 13 46 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=1.225
+ $X2=0.78 $Y2=1.225
r95 13 14 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.615 $Y=1.225
+ $X2=0.355 $Y2=1.225
r96 4 35 400 $w=1.7e-07 $l=1.07034e-06 $layer=licon1_PDIFF $count=1 $X=1.53
+ $Y=1.84 $X2=1.73 $Y2=2.815
r97 4 33 400 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=1 $X=1.53
+ $Y=1.84 $X2=1.73 $Y2=1.985
r98 3 21 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.84 $X2=0.73 $Y2=2.815
r99 3 19 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.84 $X2=0.73 $Y2=1.985
r100 2 39 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.765
+ $Y=0.37 $X2=1.905 $Y2=0.515
r101 1 25 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.64
+ $Y=0.37 $X2=0.78 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__O311A_4%A_1034_392# 1 2 3 14 18 24 25
r36 23 25 8.52431 $w=3.63e-07 $l=1.65e-07 $layer=LI1_cond $X=6.385 $Y=2.892
+ $X2=6.55 $Y2=2.892
r37 23 24 6.36223 $w=3.63e-07 $l=1.65e-07 $layer=LI1_cond $X=6.385 $Y=2.892
+ $X2=6.22 $Y2=2.892
r38 18 21 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=8.36 $Y=2.135
+ $X2=8.36 $Y2=2.815
r39 16 21 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=8.36 $Y=2.905 $X2=8.36
+ $Y2=2.815
r40 14 16 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.195 $Y=2.99
+ $X2=8.36 $Y2=2.905
r41 14 25 107.321 $w=1.68e-07 $l=1.645e-06 $layer=LI1_cond $X=8.195 $Y=2.99
+ $X2=6.55 $Y2=2.99
r42 12 24 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=5.39 $Y=2.835
+ $X2=6.22 $Y2=2.835
r43 3 21 400 $w=1.7e-07 $l=9.40705e-07 $layer=licon1_PDIFF $count=1 $X=8.18
+ $Y=1.96 $X2=8.36 $Y2=2.815
r44 3 18 400 $w=1.7e-07 $l=2.52785e-07 $layer=licon1_PDIFF $count=1 $X=8.18
+ $Y=1.96 $X2=8.36 $Y2=2.135
r45 2 23 600 $w=1.7e-07 $l=9.16938e-07 $layer=licon1_PDIFF $count=1 $X=6.235
+ $Y=1.96 $X2=6.385 $Y2=2.805
r46 1 12 600 $w=1.7e-07 $l=9.38576e-07 $layer=licon1_PDIFF $count=1 $X=5.17
+ $Y=1.96 $X2=5.39 $Y2=2.795
.ends

.subckt PM_SKY130_FD_SC_LS__O311A_4%A_1338_392# 1 2 7 13
r11 11 13 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=7.9 $Y=2.565 $X2=7.9
+ $Y2=2.135
r12 7 11 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=7.775 $Y=2.65
+ $X2=7.9 $Y2=2.565
r13 7 9 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=7.775 $Y=2.65
+ $X2=6.92 $Y2=2.65
r14 2 13 300 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=2 $X=7.71
+ $Y=1.96 $X2=7.86 $Y2=2.135
r15 1 9 600 $w=1.7e-07 $l=7.96743e-07 $layer=licon1_PDIFF $count=1 $X=6.69
+ $Y=1.96 $X2=6.92 $Y2=2.65
.ends

.subckt PM_SKY130_FD_SC_LS__O311A_4%VGND 1 2 3 4 5 6 19 21 25 29 33 37 41 44 45
+ 46 48 57 64 69 76 77 83 86 89 92
c99 21 0 1.56729e-19 $X=0.35 $Y=0.515
r100 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r101 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r102 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r103 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r104 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r105 77 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=7.92
+ $Y2=0
r106 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r107 74 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.095 $Y=0 $X2=7.93
+ $Y2=0
r108 74 76 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=8.095 $Y=0 $X2=8.4
+ $Y2=0
r109 73 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=7.92
+ $Y2=0
r110 73 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=6.96
+ $Y2=0
r111 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r112 70 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.095 $Y=0 $X2=6.93
+ $Y2=0
r113 70 72 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=7.095 $Y=0 $X2=7.44
+ $Y2=0
r114 69 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.765 $Y=0 $X2=7.93
+ $Y2=0
r115 69 72 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=7.765 $Y=0
+ $X2=7.44 $Y2=0
r116 68 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6.96
+ $Y2=0
r117 68 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r118 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r119 65 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.095 $Y=0 $X2=5.93
+ $Y2=0
r120 65 67 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=6.095 $Y=0
+ $X2=6.48 $Y2=0
r121 64 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.765 $Y=0 $X2=6.93
+ $Y2=0
r122 64 67 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=6.765 $Y=0
+ $X2=6.48 $Y2=0
r123 63 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r124 62 63 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r125 59 62 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=2.64 $Y=0 $X2=5.52
+ $Y2=0
r126 59 60 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r127 57 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.765 $Y=0 $X2=5.93
+ $Y2=0
r128 57 62 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=5.765 $Y=0 $X2=5.52
+ $Y2=0
r129 56 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r130 56 84 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.2
+ $Y2=0
r131 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r132 53 83 10.6558 $w=1.7e-07 $l=2.28e-07 $layer=LI1_cond $X=1.57 $Y=0 $X2=1.342
+ $Y2=0
r133 53 55 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=1.57 $Y=0 $X2=2.16
+ $Y2=0
r134 52 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r135 52 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r136 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r137 49 80 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=0
+ $X2=0.222 $Y2=0
r138 49 51 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=0
+ $X2=0.72 $Y2=0
r139 48 83 10.6558 $w=1.7e-07 $l=2.27e-07 $layer=LI1_cond $X=1.115 $Y=0
+ $X2=1.342 $Y2=0
r140 48 51 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.115 $Y=0
+ $X2=0.72 $Y2=0
r141 46 63 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=4.32 $Y=0 $X2=5.52
+ $Y2=0
r142 46 60 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=4.32 $Y=0
+ $X2=2.64 $Y2=0
r143 44 55 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=2.24 $Y=0 $X2=2.16
+ $Y2=0
r144 44 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.24 $Y=0 $X2=2.405
+ $Y2=0
r145 43 59 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=2.57 $Y=0 $X2=2.64
+ $Y2=0
r146 43 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.57 $Y=0 $X2=2.405
+ $Y2=0
r147 39 92 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.93 $Y=0.085
+ $X2=7.93 $Y2=0
r148 39 41 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=7.93 $Y=0.085
+ $X2=7.93 $Y2=0.535
r149 35 89 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.93 $Y=0.085
+ $X2=6.93 $Y2=0
r150 35 37 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=6.93 $Y=0.085
+ $X2=6.93 $Y2=0.535
r151 31 86 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.93 $Y=0.085
+ $X2=5.93 $Y2=0
r152 31 33 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=5.93 $Y=0.085
+ $X2=5.93 $Y2=0.535
r153 27 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.405 $Y=0.085
+ $X2=2.405 $Y2=0
r154 27 29 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.405 $Y=0.085
+ $X2=2.405 $Y2=0.515
r155 23 83 1.82608 $w=4.55e-07 $l=8.5e-08 $layer=LI1_cond $X=1.342 $Y=0.085
+ $X2=1.342 $Y2=0
r156 23 25 11.3036 $w=4.53e-07 $l=4.3e-07 $layer=LI1_cond $X=1.342 $Y=0.085
+ $X2=1.342 $Y2=0.515
r157 19 80 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.222 $Y2=0
r158 19 21 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.28 $Y2=0.515
r159 6 41 182 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=1 $X=7.775
+ $Y=0.39 $X2=7.93 $Y2=0.535
r160 5 37 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=6.72
+ $Y=0.39 $X2=6.93 $Y2=0.535
r161 4 33 182 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_NDIFF $count=1 $X=5.75
+ $Y=0.39 $X2=5.93 $Y2=0.535
r162 3 29 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.265
+ $Y=0.37 $X2=2.405 $Y2=0.515
r163 2 25 182 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_NDIFF $count=1 $X=1.07
+ $Y=0.37 $X2=1.34 $Y2=0.515
r164 1 21 91 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.35 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__O311A_4%A_564_78# 1 2 3 4 5 18 20 21 23 26 30 32 36
+ 38 40 42 46 48
r83 40 50 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.4 $Y=0.79 $X2=8.4
+ $Y2=0.875
r84 40 42 12.6769 $w=2.48e-07 $l=2.75e-07 $layer=LI1_cond $X=8.4 $Y=0.79 $X2=8.4
+ $Y2=0.515
r85 39 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.595 $Y=0.875
+ $X2=7.43 $Y2=0.875
r86 38 50 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.275 $Y=0.875
+ $X2=8.4 $Y2=0.875
r87 38 39 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=8.275 $Y=0.875
+ $X2=7.595 $Y2=0.875
r88 34 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.43 $Y=0.79 $X2=7.43
+ $Y2=0.875
r89 34 36 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=7.43 $Y=0.79
+ $X2=7.43 $Y2=0.515
r90 33 46 8.61065 $w=1.7e-07 $l=1.86145e-07 $layer=LI1_cond $X=6.595 $Y=0.875
+ $X2=6.43 $Y2=0.92
r91 32 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.265 $Y=0.875
+ $X2=7.43 $Y2=0.875
r92 32 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.265 $Y=0.875
+ $X2=6.595 $Y2=0.875
r93 28 46 0.89609 $w=3.3e-07 $l=1.3e-07 $layer=LI1_cond $X=6.43 $Y=0.79 $X2=6.43
+ $Y2=0.92
r94 28 30 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=6.43 $Y=0.79
+ $X2=6.43 $Y2=0.535
r95 27 45 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.595 $Y=0.875
+ $X2=5.43 $Y2=0.875
r96 26 46 8.61065 $w=1.7e-07 $l=1.86145e-07 $layer=LI1_cond $X=6.265 $Y=0.875
+ $X2=6.43 $Y2=0.92
r97 26 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.265 $Y=0.875
+ $X2=5.595 $Y2=0.875
r98 23 45 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.43 $Y=0.79 $X2=5.43
+ $Y2=0.875
r99 23 25 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=5.43 $Y=0.79
+ $X2=5.43 $Y2=0.535
r100 22 25 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=5.43 $Y=0.425
+ $X2=5.43 $Y2=0.535
r101 20 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.265 $Y=0.34
+ $X2=5.43 $Y2=0.425
r102 20 21 139.289 $w=1.68e-07 $l=2.135e-06 $layer=LI1_cond $X=5.265 $Y=0.34
+ $X2=3.13 $Y2=0.34
r103 16 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.965 $Y=0.425
+ $X2=3.13 $Y2=0.34
r104 16 18 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=2.965 $Y=0.425
+ $X2=2.965 $Y2=0.67
r105 5 50 182 $w=1.7e-07 $l=5.50568e-07 $layer=licon1_NDIFF $count=1 $X=8.22
+ $Y=0.39 $X2=8.36 $Y2=0.875
r106 5 42 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=8.22
+ $Y=0.39 $X2=8.36 $Y2=0.515
r107 4 48 182 $w=1.7e-07 $l=5.70044e-07 $layer=licon1_NDIFF $count=1 $X=7.245
+ $Y=0.39 $X2=7.43 $Y2=0.875
r108 4 36 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=7.245
+ $Y=0.39 $X2=7.43 $Y2=0.515
r109 3 30 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=6.285
+ $Y=0.39 $X2=6.43 $Y2=0.535
r110 2 45 182 $w=1.7e-07 $l=5.80582e-07 $layer=licon1_NDIFF $count=1 $X=5.22
+ $Y=0.39 $X2=5.43 $Y2=0.875
r111 2 25 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=5.22
+ $Y=0.39 $X2=5.43 $Y2=0.535
r112 1 18 182 $w=1.7e-07 $l=3.44964e-07 $layer=licon1_NDIFF $count=1 $X=2.82
+ $Y=0.39 $X2=2.965 $Y2=0.67
.ends

.subckt PM_SKY130_FD_SC_LS__O311A_4%A_651_78# 1 2 9 12 13 14
r20 14 17 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=4.93 $Y=0.68
+ $X2=4.93 $Y2=0.775
r21 12 13 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.91 $Y=0.76
+ $X2=4.075 $Y2=0.76
r22 9 14 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.765 $Y=0.68
+ $X2=4.93 $Y2=0.68
r23 9 13 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.765 $Y=0.68
+ $X2=4.075 $Y2=0.68
r24 2 17 182 $w=1.7e-07 $l=4.49583e-07 $layer=licon1_NDIFF $count=1 $X=4.79
+ $Y=0.39 $X2=4.93 $Y2=0.775
r25 1 12 91 $w=1.7e-07 $l=8.19375e-07 $layer=licon1_NDIFF $count=2 $X=3.255
+ $Y=0.39 $X2=3.91 $Y2=0.76
.ends

