* File: sky130_fd_sc_ls__nor3_1.pxi.spice
* Created: Fri Aug 28 13:38:10 2020
* 
x_PM_SKY130_FD_SC_LS__NOR3_1%A N_A_c_38_n N_A_M1004_g N_A_c_39_n N_A_M1003_g A A
+ PM_SKY130_FD_SC_LS__NOR3_1%A
x_PM_SKY130_FD_SC_LS__NOR3_1%B N_B_c_66_n N_B_M1001_g N_B_M1005_g B
+ PM_SKY130_FD_SC_LS__NOR3_1%B
x_PM_SKY130_FD_SC_LS__NOR3_1%C N_C_M1002_g N_C_c_100_n N_C_M1000_g C N_C_c_101_n
+ PM_SKY130_FD_SC_LS__NOR3_1%C
x_PM_SKY130_FD_SC_LS__NOR3_1%VPWR N_VPWR_M1003_s N_VPWR_c_121_n N_VPWR_c_122_n
+ N_VPWR_c_123_n VPWR N_VPWR_c_124_n N_VPWR_c_120_n
+ PM_SKY130_FD_SC_LS__NOR3_1%VPWR
x_PM_SKY130_FD_SC_LS__NOR3_1%Y N_Y_M1004_d N_Y_M1002_d N_Y_M1000_d N_Y_c_147_n
+ N_Y_c_148_n N_Y_c_149_n N_Y_c_150_n N_Y_c_151_n Y Y Y Y
+ PM_SKY130_FD_SC_LS__NOR3_1%Y
x_PM_SKY130_FD_SC_LS__NOR3_1%VGND N_VGND_M1004_s N_VGND_M1005_d N_VGND_c_195_n
+ N_VGND_c_196_n N_VGND_c_197_n N_VGND_c_198_n N_VGND_c_199_n VGND
+ N_VGND_c_200_n N_VGND_c_201_n N_VGND_c_202_n N_VGND_c_203_n
+ PM_SKY130_FD_SC_LS__NOR3_1%VGND
cc_1 VNB N_A_c_38_n 0.0204394f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.22
cc_2 VNB N_A_c_39_n 0.0626151f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.765
cc_3 VNB A 0.00896353f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_B_c_66_n 0.0305391f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.22
cc_5 VNB N_B_M1005_g 0.0218836f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_6 VNB B 0.00387716f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_7 VNB N_C_M1002_g 0.0310069f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_8 VNB N_C_c_100_n 0.0597531f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_9 VNB N_C_c_101_n 0.00431086f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_10 VNB N_VPWR_c_120_n 0.0840719f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_Y_c_147_n 0.00369654f $X=-0.19 $Y=-0.245 $X2=0.345 $Y2=1.385
cc_12 VNB N_Y_c_148_n 0.00168586f $X=-0.19 $Y=-0.245 $X2=0.232 $Y2=1.295
cc_13 VNB N_Y_c_149_n 0.0160949f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_Y_c_150_n 0.0227723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_Y_c_151_n 0.00398282f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_VGND_c_195_n 0.0120272f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_17 VNB N_VGND_c_196_n 0.0158675f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_VGND_c_197_n 0.0110726f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_19 VNB N_VGND_c_198_n 0.00568581f $X=-0.19 $Y=-0.245 $X2=0.232 $Y2=1.385
cc_20 VNB N_VGND_c_199_n 0.00626527f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_200_n 0.0150599f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_201_n 0.0191515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_202_n 0.138456f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_203_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VPB N_A_c_39_n 0.0248333f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.765
cc_26 VPB A 0.00799838f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_27 VPB N_B_c_66_n 0.022515f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.22
cc_28 VPB B 0.00373582f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_29 VPB N_C_c_100_n 0.0295642f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_30 VPB N_C_c_101_n 0.00740333f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_31 VPB N_VPWR_c_121_n 0.0140744f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_32 VPB N_VPWR_c_122_n 0.0397688f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_33 VPB N_VPWR_c_123_n 0.0063263f $X=-0.19 $Y=1.66 $X2=0.345 $Y2=1.385
cc_34 VPB N_VPWR_c_124_n 0.0397956f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_35 VPB N_VPWR_c_120_n 0.0524524f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_36 VPB N_Y_c_147_n 0.00222773f $X=-0.19 $Y=1.66 $X2=0.345 $Y2=1.385
cc_37 VPB Y 0.0502611f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_38 N_A_c_39_n N_B_c_66_n 0.0843072f $X=0.495 $Y=1.765 $X2=-0.19 $Y2=-0.245
cc_39 N_A_c_38_n N_B_M1005_g 0.0113716f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_40 N_A_c_39_n N_B_M1005_g 0.0034836f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_41 N_A_c_39_n B 4.32665e-19 $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_42 N_A_c_39_n N_VPWR_c_121_n 0.00116809f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_43 A N_VPWR_c_121_n 0.0226331f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_44 N_A_c_39_n N_VPWR_c_122_n 0.00942805f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_45 N_A_c_39_n N_VPWR_c_123_n 0.00222199f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_46 N_A_c_39_n N_VPWR_c_124_n 0.00413917f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_47 N_A_c_39_n N_VPWR_c_120_n 0.00817532f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_48 N_A_c_38_n N_Y_c_147_n 0.00310315f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_49 N_A_c_39_n N_Y_c_147_n 0.0306567f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_50 A N_Y_c_147_n 0.0429724f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_51 N_A_c_38_n N_Y_c_148_n 2.26494e-19 $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_52 N_A_c_38_n N_Y_c_151_n 0.00948239f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_53 N_A_c_38_n N_VGND_c_196_n 0.00707603f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_54 N_A_c_39_n N_VGND_c_197_n 0.00172545f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_55 A N_VGND_c_197_n 0.0221597f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_56 N_A_c_38_n N_VGND_c_198_n 4.67172e-19 $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_57 N_A_c_38_n N_VGND_c_199_n 0.00286134f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_58 N_A_c_39_n N_VGND_c_199_n 9.27443e-19 $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_59 N_A_c_38_n N_VGND_c_200_n 0.00383152f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_60 N_A_c_38_n N_VGND_c_202_n 0.00757637f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_61 N_B_M1005_g N_C_M1002_g 0.0280261f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_62 N_B_c_66_n N_C_c_100_n 0.0695475f $X=0.915 $Y=1.765 $X2=0 $Y2=0
cc_63 B N_C_c_100_n 0.00409357f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_64 N_B_c_66_n N_C_c_101_n 3.30611e-19 $X=0.915 $Y=1.765 $X2=0 $Y2=0
cc_65 B N_C_c_101_n 0.0388906f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_66 N_B_c_66_n N_VPWR_c_122_n 5.45278e-19 $X=0.915 $Y=1.765 $X2=0 $Y2=0
cc_67 N_B_c_66_n N_VPWR_c_123_n 4.70981e-19 $X=0.915 $Y=1.765 $X2=0 $Y2=0
cc_68 N_B_c_66_n N_VPWR_c_124_n 0.00291649f $X=0.915 $Y=1.765 $X2=0 $Y2=0
cc_69 N_B_c_66_n N_VPWR_c_120_n 0.00359917f $X=0.915 $Y=1.765 $X2=0 $Y2=0
cc_70 N_B_c_66_n N_Y_c_147_n 0.00651562f $X=0.915 $Y=1.765 $X2=0 $Y2=0
cc_71 N_B_M1005_g N_Y_c_147_n 0.00356835f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_72 B N_Y_c_147_n 0.0368991f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_73 N_B_M1005_g N_Y_c_148_n 2.26494e-19 $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_74 N_B_c_66_n N_Y_c_149_n 0.00464439f $X=0.915 $Y=1.765 $X2=0 $Y2=0
cc_75 N_B_M1005_g N_Y_c_149_n 0.0157822f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_76 B N_Y_c_149_n 0.0357518f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_77 N_B_M1005_g N_Y_c_150_n 5.9203e-19 $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_78 N_B_c_66_n N_Y_c_151_n 4.44413e-19 $X=0.915 $Y=1.765 $X2=0 $Y2=0
cc_79 N_B_c_66_n Y 0.0441341f $X=0.915 $Y=1.765 $X2=0 $Y2=0
cc_80 B Y 0.0351114f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_81 N_B_M1005_g N_VGND_c_196_n 4.66889e-19 $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_82 N_B_M1005_g N_VGND_c_198_n 0.00803107f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_83 N_B_M1005_g N_VGND_c_200_n 0.00383152f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_84 N_B_M1005_g N_VGND_c_202_n 0.00757637f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_85 N_C_c_100_n N_VPWR_c_124_n 0.00291649f $X=1.425 $Y=1.765 $X2=0 $Y2=0
cc_86 N_C_c_100_n N_VPWR_c_120_n 0.00363572f $X=1.425 $Y=1.765 $X2=0 $Y2=0
cc_87 N_C_M1002_g N_Y_c_149_n 0.0193333f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_88 N_C_c_100_n N_Y_c_149_n 0.00302572f $X=1.425 $Y=1.765 $X2=0 $Y2=0
cc_89 N_C_c_101_n N_Y_c_149_n 0.0276802f $X=1.65 $Y=1.465 $X2=0 $Y2=0
cc_90 N_C_M1002_g N_Y_c_150_n 0.00889319f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_91 N_C_c_100_n Y 0.0396925f $X=1.425 $Y=1.765 $X2=0 $Y2=0
cc_92 N_C_c_101_n Y 0.0265942f $X=1.65 $Y=1.465 $X2=0 $Y2=0
cc_93 N_C_M1002_g N_VGND_c_198_n 0.00503266f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_94 N_C_M1002_g N_VGND_c_201_n 0.00434272f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_95 N_C_M1002_g N_VGND_c_202_n 0.00824429f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_96 N_VPWR_c_121_n N_Y_c_147_n 0.0134237f $X=0.27 $Y=2.115 $X2=0 $Y2=0
cc_97 N_VPWR_c_123_n N_Y_c_147_n 0.0255419f $X=0.27 $Y=2.455 $X2=0 $Y2=0
cc_98 N_VPWR_c_124_n N_Y_c_147_n 0.00421728f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_99 N_VPWR_c_120_n N_Y_c_147_n 0.00350217f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_100 N_VPWR_c_124_n Y 0.048615f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_101 N_VPWR_c_120_n Y 0.0396953f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_102 A_114_368# N_Y_c_147_n 0.00244646f $X=0.57 $Y=1.84 $X2=0.615 $Y2=1.95
cc_103 A_114_368# Y 0.00369906f $X=0.57 $Y=1.84 $X2=1.595 $Y2=2.32
cc_104 A_198_368# Y 0.00259008f $X=0.99 $Y=1.84 $X2=1.595 $Y2=2.32
cc_105 N_Y_c_149_n N_VGND_M1005_d 0.00253871f $X=1.475 $Y=1.005 $X2=0 $Y2=0
cc_106 N_Y_c_148_n N_VGND_c_196_n 0.0130608f $X=0.71 $Y=0.53 $X2=0 $Y2=0
cc_107 N_Y_c_151_n N_VGND_c_197_n 0.0104845f $X=0.71 $Y=0.965 $X2=0 $Y2=0
cc_108 N_Y_c_148_n N_VGND_c_198_n 0.0130983f $X=0.71 $Y=0.53 $X2=0 $Y2=0
cc_109 N_Y_c_149_n N_VGND_c_198_n 0.0215485f $X=1.475 $Y=1.005 $X2=0 $Y2=0
cc_110 N_Y_c_150_n N_VGND_c_198_n 0.0142986f $X=1.64 $Y=0.515 $X2=0 $Y2=0
cc_111 N_Y_c_148_n N_VGND_c_200_n 0.00791198f $X=0.71 $Y=0.53 $X2=0 $Y2=0
cc_112 N_Y_c_150_n N_VGND_c_201_n 0.0145639f $X=1.64 $Y=0.515 $X2=0 $Y2=0
cc_113 N_Y_c_148_n N_VGND_c_202_n 0.00688042f $X=0.71 $Y=0.53 $X2=0 $Y2=0
cc_114 N_Y_c_150_n N_VGND_c_202_n 0.0119984f $X=1.64 $Y=0.515 $X2=0 $Y2=0
