* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__dlxtn_4 D GATE_N VGND VNB VPB VPWR Q
M1000 VPWR a_840_395# Q VPB phighvt w=1.12e+06u l=150000u
+  ad=2.3143e+12p pd=1.737e+07u as=7.56e+11p ps=5.83e+06u
M1001 a_658_79# a_27_115# VGND VNB nshort w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=1.78397e+12p ps=1.439e+07u
M1002 a_591_392# a_27_115# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1003 VGND a_840_395# a_895_123# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1004 VPWR D a_27_115# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=2.478e+11p ps=2.27e+06u
M1005 a_840_395# a_675_392# VPWR VPB phighvt w=840000u l=150000u
+  ad=2.982e+11p pd=2.39e+06u as=0p ps=0u
M1006 VPWR a_675_392# a_840_395# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND a_230_424# a_369_392# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1008 Q a_840_395# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Q a_840_395# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND a_675_392# a_840_395# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1011 VPWR a_230_424# a_369_392# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=2.478e+11p ps=2.27e+06u
M1012 VPWR a_840_395# a_789_508# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1013 a_895_123# a_369_392# a_675_392# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=3.259e+11p ps=2.57e+06u
M1014 VGND D a_27_115# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1015 VPWR a_840_395# Q VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Q a_840_395# VGND VNB nshort w=740000u l=150000u
+  ad=5.143e+11p pd=4.35e+06u as=0p ps=0u
M1017 a_230_424# GATE_N VPWR VPB phighvt w=840000u l=150000u
+  ad=2.478e+11p pd=2.27e+06u as=0p ps=0u
M1018 Q a_840_395# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_789_508# a_230_424# a_675_392# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=3.475e+11p ps=2.84e+06u
M1020 a_230_424# GATE_N VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1021 a_840_395# a_675_392# VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND a_840_395# Q VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VGND a_840_395# Q VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_675_392# a_369_392# a_591_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_675_392# a_230_424# a_658_79# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
