* File: sky130_fd_sc_ls__sdfrtp_1.pxi.spice
* Created: Wed Sep  2 11:27:16 2020
* 
x_PM_SKY130_FD_SC_LS__SDFRTP_1%SCE N_SCE_c_308_n N_SCE_M1033_g N_SCE_c_309_n
+ N_SCE_M1020_g N_SCE_c_310_n N_SCE_c_311_n N_SCE_M1017_g N_SCE_M1024_g
+ N_SCE_c_300_n N_SCE_c_301_n N_SCE_c_302_n N_SCE_c_303_n N_SCE_c_304_n SCE SCE
+ SCE N_SCE_c_305_n N_SCE_c_306_n N_SCE_c_307_n SCE N_SCE_c_315_n
+ PM_SKY130_FD_SC_LS__SDFRTP_1%SCE
x_PM_SKY130_FD_SC_LS__SDFRTP_1%A_27_88# N_A_27_88#_M1033_s N_A_27_88#_M1020_s
+ N_A_27_88#_c_395_n N_A_27_88#_M1005_g N_A_27_88#_M1022_g N_A_27_88#_c_403_n
+ N_A_27_88#_c_396_n N_A_27_88#_c_397_n N_A_27_88#_c_405_n N_A_27_88#_c_398_n
+ N_A_27_88#_c_406_n N_A_27_88#_c_407_n N_A_27_88#_c_399_n N_A_27_88#_c_408_n
+ N_A_27_88#_c_400_n N_A_27_88#_c_401_n N_A_27_88#_c_409_n
+ PM_SKY130_FD_SC_LS__SDFRTP_1%A_27_88#
x_PM_SKY130_FD_SC_LS__SDFRTP_1%D N_D_c_485_n N_D_M1011_g N_D_c_479_n N_D_c_480_n
+ N_D_M1006_g N_D_c_487_n N_D_c_481_n D N_D_c_482_n N_D_c_483_n N_D_c_484_n
+ PM_SKY130_FD_SC_LS__SDFRTP_1%D
x_PM_SKY130_FD_SC_LS__SDFRTP_1%SCD N_SCD_M1026_g N_SCD_M1012_g N_SCD_c_537_n
+ N_SCD_c_541_n SCD SCD N_SCD_c_539_n PM_SKY130_FD_SC_LS__SDFRTP_1%SCD
x_PM_SKY130_FD_SC_LS__SDFRTP_1%CLK N_CLK_c_577_n N_CLK_c_578_n N_CLK_c_579_n
+ N_CLK_M1028_g N_CLK_c_580_n N_CLK_M1027_g N_CLK_c_581_n N_CLK_c_586_n CLK
+ N_CLK_c_583_n N_CLK_c_584_n PM_SKY130_FD_SC_LS__SDFRTP_1%CLK
x_PM_SKY130_FD_SC_LS__SDFRTP_1%A_1034_392# N_A_1034_392#_M1032_d
+ N_A_1034_392#_M1030_d N_A_1034_392#_c_664_n N_A_1034_392#_c_665_n
+ N_A_1034_392#_M1039_g N_A_1034_392#_c_644_n N_A_1034_392#_M1000_g
+ N_A_1034_392#_c_646_n N_A_1034_392#_M1003_g N_A_1034_392#_c_647_n
+ N_A_1034_392#_c_667_n N_A_1034_392#_M1014_g N_A_1034_392#_c_668_n
+ N_A_1034_392#_c_648_n N_A_1034_392#_c_649_n N_A_1034_392#_c_650_n
+ N_A_1034_392#_c_651_n N_A_1034_392#_c_669_n N_A_1034_392#_c_652_n
+ N_A_1034_392#_c_653_n N_A_1034_392#_c_654_n N_A_1034_392#_c_680_p
+ N_A_1034_392#_c_707_p N_A_1034_392#_c_655_n N_A_1034_392#_c_656_n
+ N_A_1034_392#_c_657_n N_A_1034_392#_c_658_n N_A_1034_392#_c_785_p
+ N_A_1034_392#_c_672_n N_A_1034_392#_c_659_n N_A_1034_392#_c_660_n
+ N_A_1034_392#_c_661_n N_A_1034_392#_c_662_n N_A_1034_392#_c_663_n
+ PM_SKY130_FD_SC_LS__SDFRTP_1%A_1034_392#
x_PM_SKY130_FD_SC_LS__SDFRTP_1%A_1367_93# N_A_1367_93#_M1031_d
+ N_A_1367_93#_M1013_d N_A_1367_93#_M1019_g N_A_1367_93#_c_871_n
+ N_A_1367_93#_c_872_n N_A_1367_93#_M1008_g N_A_1367_93#_c_865_n
+ N_A_1367_93#_c_866_n N_A_1367_93#_c_867_n N_A_1367_93#_c_868_n
+ N_A_1367_93#_c_875_n N_A_1367_93#_c_876_n N_A_1367_93#_c_869_n
+ N_A_1367_93#_c_870_n PM_SKY130_FD_SC_LS__SDFRTP_1%A_1367_93#
x_PM_SKY130_FD_SC_LS__SDFRTP_1%RESET_B N_RESET_B_M1037_g N_RESET_B_M1038_g
+ N_RESET_B_c_977_n N_RESET_B_c_978_n N_RESET_B_c_987_n N_RESET_B_c_988_n
+ N_RESET_B_M1007_g N_RESET_B_c_980_n N_RESET_B_c_981_n N_RESET_B_c_982_n
+ N_RESET_B_c_990_n N_RESET_B_M1009_g N_RESET_B_M1036_g N_RESET_B_c_984_n
+ N_RESET_B_c_992_n N_RESET_B_c_993_n N_RESET_B_M1016_g N_RESET_B_c_994_n
+ N_RESET_B_c_985_n N_RESET_B_c_995_n N_RESET_B_c_996_n N_RESET_B_c_997_n
+ N_RESET_B_c_998_n N_RESET_B_c_999_n RESET_B N_RESET_B_c_1001_n
+ N_RESET_B_c_1002_n N_RESET_B_c_1003_n N_RESET_B_c_1004_n
+ PM_SKY130_FD_SC_LS__SDFRTP_1%RESET_B
x_PM_SKY130_FD_SC_LS__SDFRTP_1%A_1234_119# N_A_1234_119#_M1035_d
+ N_A_1234_119#_M1039_d N_A_1234_119#_M1009_d N_A_1234_119#_M1031_g
+ N_A_1234_119#_c_1207_n N_A_1234_119#_c_1216_n N_A_1234_119#_M1013_g
+ N_A_1234_119#_c_1217_n N_A_1234_119#_c_1208_n N_A_1234_119#_c_1209_n
+ N_A_1234_119#_c_1253_n N_A_1234_119#_c_1210_n N_A_1234_119#_c_1211_n
+ N_A_1234_119#_c_1212_n N_A_1234_119#_c_1213_n N_A_1234_119#_c_1214_n
+ N_A_1234_119#_c_1221_n PM_SKY130_FD_SC_LS__SDFRTP_1%A_1234_119#
x_PM_SKY130_FD_SC_LS__SDFRTP_1%A_835_98# N_A_835_98#_M1028_s N_A_835_98#_M1027_s
+ N_A_835_98#_c_1354_n N_A_835_98#_M1030_g N_A_835_98#_c_1342_n
+ N_A_835_98#_M1032_g N_A_835_98#_c_1355_n N_A_835_98#_c_1356_n
+ N_A_835_98#_c_1357_n N_A_835_98#_c_1343_n N_A_835_98#_c_1344_n
+ N_A_835_98#_M1035_g N_A_835_98#_c_1358_n N_A_835_98#_c_1359_n
+ N_A_835_98#_c_1360_n N_A_835_98#_M1029_g N_A_835_98#_c_1361_n
+ N_A_835_98#_c_1362_n N_A_835_98#_c_1363_n N_A_835_98#_M1018_g
+ N_A_835_98#_c_1345_n N_A_835_98#_c_1346_n N_A_835_98#_c_1347_n
+ N_A_835_98#_M1002_g N_A_835_98#_c_1367_n N_A_835_98#_c_1349_n
+ N_A_835_98#_c_1373_n N_A_835_98#_c_1374_n N_A_835_98#_c_1376_n
+ N_A_835_98#_c_1350_n N_A_835_98#_c_1351_n N_A_835_98#_c_1352_n
+ N_A_835_98#_c_1353_n PM_SKY130_FD_SC_LS__SDFRTP_1%A_835_98#
x_PM_SKY130_FD_SC_LS__SDFRTP_1%A_1997_272# N_A_1997_272#_M1021_d
+ N_A_1997_272#_M1016_d N_A_1997_272#_M1001_g N_A_1997_272#_c_1544_n
+ N_A_1997_272#_c_1555_n N_A_1997_272#_c_1556_n N_A_1997_272#_M1034_g
+ N_A_1997_272#_c_1545_n N_A_1997_272#_c_1546_n N_A_1997_272#_c_1547_n
+ N_A_1997_272#_c_1548_n N_A_1997_272#_c_1549_n N_A_1997_272#_c_1550_n
+ N_A_1997_272#_c_1551_n N_A_1997_272#_c_1557_n N_A_1997_272#_c_1552_n
+ N_A_1997_272#_c_1553_n PM_SKY130_FD_SC_LS__SDFRTP_1%A_1997_272#
x_PM_SKY130_FD_SC_LS__SDFRTP_1%A_1745_74# N_A_1745_74#_M1003_d
+ N_A_1745_74#_M1018_d N_A_1745_74#_M1021_g N_A_1745_74#_c_1661_n
+ N_A_1745_74#_c_1672_n N_A_1745_74#_c_1673_n N_A_1745_74#_M1023_g
+ N_A_1745_74#_c_1662_n N_A_1745_74#_c_1663_n N_A_1745_74#_c_1674_n
+ N_A_1745_74#_c_1675_n N_A_1745_74#_M1010_g N_A_1745_74#_M1025_g
+ N_A_1745_74#_c_1676_n N_A_1745_74#_c_1677_n N_A_1745_74#_c_1665_n
+ N_A_1745_74#_c_1666_n N_A_1745_74#_c_1679_n N_A_1745_74#_c_1680_n
+ N_A_1745_74#_c_1681_n N_A_1745_74#_c_1667_n N_A_1745_74#_c_1668_n
+ N_A_1745_74#_c_1669_n N_A_1745_74#_c_1670_n
+ PM_SKY130_FD_SC_LS__SDFRTP_1%A_1745_74#
x_PM_SKY130_FD_SC_LS__SDFRTP_1%A_2399_424# N_A_2399_424#_M1025_d
+ N_A_2399_424#_M1010_d N_A_2399_424#_c_1832_n N_A_2399_424#_M1015_g
+ N_A_2399_424#_M1004_g N_A_2399_424#_c_1828_n N_A_2399_424#_c_1834_n
+ N_A_2399_424#_c_1829_n N_A_2399_424#_c_1854_p N_A_2399_424#_c_1830_n
+ N_A_2399_424#_c_1831_n PM_SKY130_FD_SC_LS__SDFRTP_1%A_2399_424#
x_PM_SKY130_FD_SC_LS__SDFRTP_1%VPWR N_VPWR_M1020_d N_VPWR_M1026_d N_VPWR_M1027_d
+ N_VPWR_M1008_d N_VPWR_M1013_s N_VPWR_M1034_d N_VPWR_M1023_d N_VPWR_M1015_s
+ N_VPWR_c_1875_n N_VPWR_c_1876_n N_VPWR_c_1877_n N_VPWR_c_1878_n
+ N_VPWR_c_1879_n N_VPWR_c_1880_n N_VPWR_c_1881_n N_VPWR_c_1882_n
+ N_VPWR_c_1883_n N_VPWR_c_1884_n N_VPWR_c_1885_n N_VPWR_c_1886_n
+ N_VPWR_c_1887_n N_VPWR_c_1888_n N_VPWR_c_1889_n VPWR N_VPWR_c_1890_n
+ N_VPWR_c_1891_n N_VPWR_c_1892_n N_VPWR_c_1893_n N_VPWR_c_1894_n
+ N_VPWR_c_1874_n N_VPWR_c_1896_n N_VPWR_c_1897_n N_VPWR_c_1898_n
+ N_VPWR_c_1899_n N_VPWR_c_1900_n PM_SKY130_FD_SC_LS__SDFRTP_1%VPWR
x_PM_SKY130_FD_SC_LS__SDFRTP_1%A_300_464# N_A_300_464#_M1006_d
+ N_A_300_464#_M1035_s N_A_300_464#_M1011_d N_A_300_464#_M1038_d
+ N_A_300_464#_M1039_s N_A_300_464#_c_2049_n N_A_300_464#_c_2072_n
+ N_A_300_464#_c_2041_n N_A_300_464#_c_2042_n N_A_300_464#_c_2051_n
+ N_A_300_464#_c_2052_n N_A_300_464#_c_2053_n N_A_300_464#_c_2043_n
+ N_A_300_464#_c_2044_n N_A_300_464#_c_2054_n N_A_300_464#_c_2045_n
+ N_A_300_464#_c_2046_n N_A_300_464#_c_2055_n N_A_300_464#_c_2056_n
+ N_A_300_464#_c_2047_n N_A_300_464#_c_2058_n N_A_300_464#_c_2048_n
+ N_A_300_464#_c_2059_n PM_SKY130_FD_SC_LS__SDFRTP_1%A_300_464#
x_PM_SKY130_FD_SC_LS__SDFRTP_1%Q N_Q_M1004_d N_Q_M1015_d Q Q Q Q Q Q Q Q
+ PM_SKY130_FD_SC_LS__SDFRTP_1%Q
x_PM_SKY130_FD_SC_LS__SDFRTP_1%VGND N_VGND_M1033_d N_VGND_M1037_d N_VGND_M1028_d
+ N_VGND_M1007_d N_VGND_M1001_d N_VGND_M1025_s N_VGND_M1004_s N_VGND_c_2231_n
+ N_VGND_c_2232_n N_VGND_c_2233_n N_VGND_c_2234_n N_VGND_c_2235_n
+ N_VGND_c_2236_n N_VGND_c_2237_n N_VGND_c_2238_n VGND N_VGND_c_2239_n
+ N_VGND_c_2240_n N_VGND_c_2241_n N_VGND_c_2242_n N_VGND_c_2243_n
+ N_VGND_c_2244_n N_VGND_c_2245_n N_VGND_c_2246_n N_VGND_c_2247_n
+ N_VGND_c_2248_n N_VGND_c_2249_n N_VGND_c_2250_n N_VGND_c_2251_n
+ N_VGND_c_2252_n PM_SKY130_FD_SC_LS__SDFRTP_1%VGND
x_PM_SKY130_FD_SC_LS__SDFRTP_1%noxref_24 N_noxref_24_M1005_s N_noxref_24_M1012_d
+ N_noxref_24_c_2364_n N_noxref_24_c_2365_n N_noxref_24_c_2366_n
+ PM_SKY130_FD_SC_LS__SDFRTP_1%noxref_24
cc_1 VNB N_SCE_M1033_g 0.062352f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.65
cc_2 VNB N_SCE_c_300_n 0.0148916f $X=-0.19 $Y=-0.245 $X2=2.625 $Y2=0.9
cc_3 VNB N_SCE_c_301_n 0.0107474f $X=-0.19 $Y=-0.245 $X2=2.625 $Y2=1.05
cc_4 VNB N_SCE_c_302_n 0.0132325f $X=-0.19 $Y=-0.245 $X2=2.345 $Y2=1.575
cc_5 VNB N_SCE_c_303_n 0.0055883f $X=-0.19 $Y=-0.245 $X2=2.51 $Y2=1.425
cc_6 VNB N_SCE_c_304_n 0.0319913f $X=-0.19 $Y=-0.245 $X2=2.51 $Y2=1.425
cc_7 VNB N_SCE_c_305_n 0.0331371f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=1.67
cc_8 VNB N_SCE_c_306_n 0.0119307f $X=-0.19 $Y=-0.245 $X2=2.51 $Y2=1.26
cc_9 VNB N_SCE_c_307_n 0.0110089f $X=-0.19 $Y=-0.245 $X2=1.623 $Y2=1.662
cc_10 VNB N_A_27_88#_c_395_n 0.0192577f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.245
cc_11 VNB N_A_27_88#_c_396_n 0.0282802f $X=-0.19 $Y=-0.245 $X2=2.65 $Y2=0.9
cc_12 VNB N_A_27_88#_c_397_n 0.0187337f $X=-0.19 $Y=-0.245 $X2=2.625 $Y2=0.9
cc_13 VNB N_A_27_88#_c_398_n 0.0167058f $X=-0.19 $Y=-0.245 $X2=2.51 $Y2=1.425
cc_14 VNB N_A_27_88#_c_399_n 0.0130086f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_88#_c_400_n 0.00840348f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.67
cc_16 VNB N_A_27_88#_c_401_n 0.0522403f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.67
cc_17 VNB N_D_c_479_n 0.00442527f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.65
cc_18 VNB N_D_c_480_n 0.0150551f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.245
cc_19 VNB N_D_c_481_n 0.0209259f $X=-0.19 $Y=-0.245 $X2=2.6 $Y2=1.05
cc_20 VNB N_D_c_482_n 0.0321108f $X=-0.19 $Y=-0.245 $X2=2.625 $Y2=0.9
cc_21 VNB N_D_c_483_n 0.00935279f $X=-0.19 $Y=-0.245 $X2=2.625 $Y2=1.05
cc_22 VNB N_D_c_484_n 0.0161524f $X=-0.19 $Y=-0.245 $X2=2.345 $Y2=1.575
cc_23 VNB N_SCD_M1012_g 0.0413981f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_SCD_c_537_n 0.00371437f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.835
cc_25 VNB SCD 0.00356111f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.245
cc_26 VNB N_SCD_c_539_n 0.0155097f $X=-0.19 $Y=-0.245 $X2=2.65 $Y2=0.9
cc_27 VNB N_CLK_c_577_n 0.0269111f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.835
cc_28 VNB N_CLK_c_578_n 0.0142729f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.155
cc_29 VNB N_CLK_c_579_n 0.0155025f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.505
cc_30 VNB N_CLK_c_580_n 0.00413196f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.245
cc_31 VNB N_CLK_c_581_n 0.00963216f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.245
cc_32 VNB CLK 0.00427259f $X=-0.19 $Y=-0.245 $X2=2.6 $Y2=1.26
cc_33 VNB N_CLK_c_583_n 0.0396101f $X=-0.19 $Y=-0.245 $X2=2.65 $Y2=0.615
cc_34 VNB N_CLK_c_584_n 0.0120835f $X=-0.19 $Y=-0.245 $X2=2.625 $Y2=0.9
cc_35 VNB N_A_1034_392#_c_644_n 0.0112522f $X=-0.19 $Y=-0.245 $X2=1.005
+ $Y2=2.245
cc_36 VNB N_A_1034_392#_M1000_g 0.0379064f $X=-0.19 $Y=-0.245 $X2=2.6 $Y2=1.26
cc_37 VNB N_A_1034_392#_c_646_n 0.0161967f $X=-0.19 $Y=-0.245 $X2=2.65 $Y2=0.615
cc_38 VNB N_A_1034_392#_c_647_n 0.00792759f $X=-0.19 $Y=-0.245 $X2=2.345
+ $Y2=1.575
cc_39 VNB N_A_1034_392#_c_648_n 0.00991314f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_1034_392#_c_649_n 6.30651e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_1034_392#_c_650_n 0.0334399f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_1034_392#_c_651_n 0.00321642f $X=-0.19 $Y=-0.245 $X2=0.495
+ $Y2=1.67
cc_43 VNB N_A_1034_392#_c_652_n 0.00171326f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=1.67
cc_44 VNB N_A_1034_392#_c_653_n 0.00375765f $X=-0.19 $Y=-0.245 $X2=2.51 $Y2=1.26
cc_45 VNB N_A_1034_392#_c_654_n 8.10761e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_1034_392#_c_655_n 0.00889307f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_1034_392#_c_656_n 0.00224396f $X=-0.19 $Y=-0.245 $X2=0.96
+ $Y2=1.662
cc_48 VNB N_A_1034_392#_c_657_n 0.00270816f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_1034_392#_c_658_n 0.00419892f $X=-0.19 $Y=-0.245 $X2=1.68
+ $Y2=1.662
cc_50 VNB N_A_1034_392#_c_659_n 4.42537e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_1034_392#_c_660_n 0.0363807f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_1034_392#_c_661_n 0.00354363f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_1034_392#_c_662_n 0.0114218f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_1034_392#_c_663_n 0.0259737f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_1367_93#_M1019_g 0.0317694f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.64
cc_56 VNB N_A_1367_93#_c_865_n 0.00358202f $X=-0.19 $Y=-0.245 $X2=2.65 $Y2=0.615
cc_57 VNB N_A_1367_93#_c_866_n 0.0256217f $X=-0.19 $Y=-0.245 $X2=2.65 $Y2=0.615
cc_58 VNB N_A_1367_93#_c_867_n 0.00667339f $X=-0.19 $Y=-0.245 $X2=2.625 $Y2=1.05
cc_59 VNB N_A_1367_93#_c_868_n 4.38526e-19 $X=-0.19 $Y=-0.245 $X2=2.345
+ $Y2=1.575
cc_60 VNB N_A_1367_93#_c_869_n 0.00364646f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_61 VNB N_A_1367_93#_c_870_n 0.00552017f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_RESET_B_M1037_g 0.0484041f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.65
cc_63 VNB N_RESET_B_c_977_n 0.271956f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.64
cc_64 VNB N_RESET_B_c_978_n 0.012806f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.64
cc_65 VNB N_RESET_B_M1007_g 0.0265319f $X=-0.19 $Y=-0.245 $X2=2.6 $Y2=1.05
cc_66 VNB N_RESET_B_c_980_n 0.0260909f $X=-0.19 $Y=-0.245 $X2=2.6 $Y2=1.26
cc_67 VNB N_RESET_B_c_981_n 0.0069569f $X=-0.19 $Y=-0.245 $X2=2.65 $Y2=0.9
cc_68 VNB N_RESET_B_c_982_n 0.0202613f $X=-0.19 $Y=-0.245 $X2=2.65 $Y2=0.615
cc_69 VNB N_RESET_B_M1036_g 0.0378564f $X=-0.19 $Y=-0.245 $X2=2.51 $Y2=1.425
cc_70 VNB N_RESET_B_c_984_n 0.0109809f $X=-0.19 $Y=-0.245 $X2=2.535 $Y2=1.575
cc_71 VNB N_RESET_B_c_985_n 0.0164222f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=1.67
cc_72 VNB N_A_1234_119#_M1031_g 0.0268916f $X=-0.19 $Y=-0.245 $X2=1.005
+ $Y2=2.245
cc_73 VNB N_A_1234_119#_c_1207_n 0.0175736f $X=-0.19 $Y=-0.245 $X2=1.005
+ $Y2=2.64
cc_74 VNB N_A_1234_119#_c_1208_n 0.00374454f $X=-0.19 $Y=-0.245 $X2=1.795
+ $Y2=1.575
cc_75 VNB N_A_1234_119#_c_1209_n 0.00425843f $X=-0.19 $Y=-0.245 $X2=2.51
+ $Y2=1.425
cc_76 VNB N_A_1234_119#_c_1210_n 4.99311e-19 $X=-0.19 $Y=-0.245 $X2=0.635
+ $Y2=1.58
cc_77 VNB N_A_1234_119#_c_1211_n 0.00215276f $X=-0.19 $Y=-0.245 $X2=1.115
+ $Y2=1.58
cc_78 VNB N_A_1234_119#_c_1212_n 0.00602363f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_1234_119#_c_1213_n 0.0279564f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_1234_119#_c_1214_n 0.00301829f $X=-0.19 $Y=-0.245 $X2=0.495
+ $Y2=1.67
cc_81 VNB N_A_835_98#_c_1342_n 0.0155098f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.835
cc_82 VNB N_A_835_98#_c_1343_n 0.0316816f $X=-0.19 $Y=-0.245 $X2=2.65 $Y2=0.9
cc_83 VNB N_A_835_98#_c_1344_n 0.0159412f $X=-0.19 $Y=-0.245 $X2=2.65 $Y2=0.615
cc_84 VNB N_A_835_98#_c_1345_n 0.0179478f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_835_98#_c_1346_n 0.00460795f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_835_98#_c_1347_n 0.0208108f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.67
cc_87 VNB N_A_835_98#_M1002_g 0.0235073f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=1.67
cc_88 VNB N_A_835_98#_c_1349_n 0.0124432f $X=-0.19 $Y=-0.245 $X2=1.623 $Y2=1.662
cc_89 VNB N_A_835_98#_c_1350_n 0.0012852f $X=-0.19 $Y=-0.245 $X2=1.609 $Y2=1.662
cc_90 VNB N_A_835_98#_c_1351_n 0.00365945f $X=-0.19 $Y=-0.245 $X2=1.795
+ $Y2=1.662
cc_91 VNB N_A_835_98#_c_1352_n 0.00140775f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_835_98#_c_1353_n 0.0546007f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_1997_272#_M1001_g 0.0393068f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.64
cc_94 VNB N_A_1997_272#_c_1544_n 0.0235946f $X=-0.19 $Y=-0.245 $X2=1.005
+ $Y2=2.155
cc_95 VNB N_A_1997_272#_c_1545_n 0.0152817f $X=-0.19 $Y=-0.245 $X2=2.6 $Y2=1.26
cc_96 VNB N_A_1997_272#_c_1546_n 0.0073172f $X=-0.19 $Y=-0.245 $X2=2.625 $Y2=0.9
cc_97 VNB N_A_1997_272#_c_1547_n 0.00658513f $X=-0.19 $Y=-0.245 $X2=2.535
+ $Y2=1.425
cc_98 VNB N_A_1997_272#_c_1548_n 0.00719764f $X=-0.19 $Y=-0.245 $X2=2.51
+ $Y2=1.425
cc_99 VNB N_A_1997_272#_c_1549_n 0.00239418f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_A_1997_272#_c_1550_n 0.00890748f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_A_1997_272#_c_1551_n 0.00132368f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_A_1997_272#_c_1552_n 4.91246e-19 $X=-0.19 $Y=-0.245 $X2=0.495
+ $Y2=1.67
cc_103 VNB N_A_1997_272#_c_1553_n 6.26987e-19 $X=-0.19 $Y=-0.245 $X2=0.96
+ $Y2=1.67
cc_104 VNB N_A_1745_74#_M1021_g 0.0220606f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.64
cc_105 VNB N_A_1745_74#_c_1661_n 0.0178723f $X=-0.19 $Y=-0.245 $X2=1.005
+ $Y2=2.245
cc_106 VNB N_A_1745_74#_c_1662_n 0.0372707f $X=-0.19 $Y=-0.245 $X2=2.65
+ $Y2=0.615
cc_107 VNB N_A_1745_74#_c_1663_n 0.0476514f $X=-0.19 $Y=-0.245 $X2=2.65
+ $Y2=0.615
cc_108 VNB N_A_1745_74#_M1025_g 0.0313727f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_A_1745_74#_c_1665_n 0.0027518f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_A_1745_74#_c_1666_n 0.00220477f $X=-0.19 $Y=-0.245 $X2=0.495
+ $Y2=1.67
cc_111 VNB N_A_1745_74#_c_1667_n 0.00284242f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_A_1745_74#_c_1668_n 0.00104193f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_A_1745_74#_c_1669_n 8.69032e-19 $X=-0.19 $Y=-0.245 $X2=0.96
+ $Y2=1.662
cc_114 VNB N_A_1745_74#_c_1670_n 0.0278597f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_A_2399_424#_M1004_g 0.0281108f $X=-0.19 $Y=-0.245 $X2=1.005
+ $Y2=2.245
cc_116 VNB N_A_2399_424#_c_1828_n 0.0900229f $X=-0.19 $Y=-0.245 $X2=2.6 $Y2=1.05
cc_117 VNB N_A_2399_424#_c_1829_n 0.016101f $X=-0.19 $Y=-0.245 $X2=1.795
+ $Y2=1.575
cc_118 VNB N_A_2399_424#_c_1830_n 8.47259e-19 $X=-0.19 $Y=-0.245 $X2=1.595
+ $Y2=1.58
cc_119 VNB N_A_2399_424#_c_1831_n 0.00458466f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_VPWR_c_1874_n 0.561729f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_A_300_464#_c_2041_n 0.0223051f $X=-0.19 $Y=-0.245 $X2=2.345
+ $Y2=1.575
cc_122 VNB N_A_300_464#_c_2042_n 0.0037881f $X=-0.19 $Y=-0.245 $X2=2.51
+ $Y2=1.425
cc_123 VNB N_A_300_464#_c_2043_n 9.90482e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_A_300_464#_c_2044_n 0.00159941f $X=-0.19 $Y=-0.245 $X2=0.495
+ $Y2=1.67
cc_125 VNB N_A_300_464#_c_2045_n 0.00524388f $X=-0.19 $Y=-0.245 $X2=0.96
+ $Y2=1.67
cc_126 VNB N_A_300_464#_c_2046_n 0.00161435f $X=-0.19 $Y=-0.245 $X2=0.96
+ $Y2=1.67
cc_127 VNB N_A_300_464#_c_2047_n 0.00255764f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_A_300_464#_c_2048_n 0.00434949f $X=-0.19 $Y=-0.245 $X2=0.96
+ $Y2=1.662
cc_129 VNB Q 0.0259999f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.245
cc_130 VNB Q 0.00837931f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.64
cc_131 VNB Q 0.027119f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.64
cc_132 VNB N_VGND_c_2231_n 0.0181638f $X=-0.19 $Y=-0.245 $X2=2.535 $Y2=1.425
cc_133 VNB N_VGND_c_2232_n 0.0123129f $X=-0.19 $Y=-0.245 $X2=2.535 $Y2=1.575
cc_134 VNB N_VGND_c_2233_n 0.012879f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_135 VNB N_VGND_c_2234_n 0.0100142f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_VGND_c_2235_n 0.00854448f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=1.67
cc_137 VNB N_VGND_c_2236_n 0.0169646f $X=-0.19 $Y=-0.245 $X2=2.51 $Y2=1.26
cc_138 VNB N_VGND_c_2237_n 0.021767f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.662
cc_139 VNB N_VGND_c_2238_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_VGND_c_2239_n 0.0177976f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.662
cc_141 VNB N_VGND_c_2240_n 0.0636435f $X=-0.19 $Y=-0.245 $X2=1.694 $Y2=1.662
cc_142 VNB N_VGND_c_2241_n 0.0552549f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_143 VNB N_VGND_c_2242_n 0.0611983f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_144 VNB N_VGND_c_2243_n 0.0297773f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_145 VNB N_VGND_c_2244_n 0.0188435f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_146 VNB N_VGND_c_2245_n 0.0194697f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_147 VNB N_VGND_c_2246_n 0.704864f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_148 VNB N_VGND_c_2247_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_149 VNB N_VGND_c_2248_n 0.0038619f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_150 VNB N_VGND_c_2249_n 0.0140297f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_151 VNB N_VGND_c_2250_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_152 VNB N_VGND_c_2251_n 0.00622769f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_153 VNB N_VGND_c_2252_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_154 VNB N_noxref_24_c_2364_n 0.0131255f $X=-0.19 $Y=-0.245 $X2=0.505
+ $Y2=2.245
cc_155 VNB N_noxref_24_c_2365_n 0.00667823f $X=-0.19 $Y=-0.245 $X2=0.505
+ $Y2=2.64
cc_156 VNB N_noxref_24_c_2366_n 0.00408915f $X=-0.19 $Y=-0.245 $X2=1.005
+ $Y2=2.64
cc_157 VPB N_SCE_c_308_n 0.0195456f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.155
cc_158 VPB N_SCE_c_309_n 0.0273001f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.245
cc_159 VPB N_SCE_c_310_n 0.0184657f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.155
cc_160 VPB N_SCE_c_311_n 0.02161f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.245
cc_161 VPB N_SCE_c_303_n 0.00300633f $X=-0.19 $Y=1.66 $X2=2.51 $Y2=1.425
cc_162 VPB N_SCE_c_305_n 0.0253807f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=1.67
cc_163 VPB N_SCE_c_307_n 0.00455267f $X=-0.19 $Y=1.66 $X2=1.623 $Y2=1.662
cc_164 VPB N_SCE_c_315_n 0.00736556f $X=-0.19 $Y=1.66 $X2=1.795 $Y2=1.662
cc_165 VPB N_A_27_88#_M1022_g 0.0278498f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.245
cc_166 VPB N_A_27_88#_c_403_n 0.061022f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.64
cc_167 VPB N_A_27_88#_c_397_n 0.0161852f $X=-0.19 $Y=1.66 $X2=2.625 $Y2=0.9
cc_168 VPB N_A_27_88#_c_405_n 0.0338402f $X=-0.19 $Y=1.66 $X2=1.795 $Y2=1.575
cc_169 VPB N_A_27_88#_c_406_n 0.00159951f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_170 VPB N_A_27_88#_c_407_n 0.00598053f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_171 VPB N_A_27_88#_c_408_n 0.0129728f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_172 VPB N_A_27_88#_c_409_n 0.0236923f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.67
cc_173 VPB N_D_c_485_n 0.0213045f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.835
cc_174 VPB N_D_c_479_n 0.0247476f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.65
cc_175 VPB N_D_c_487_n 0.0297202f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.155
cc_176 VPB N_SCD_c_537_n 0.0317264f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.835
cc_177 VPB N_SCD_c_541_n 0.0316323f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.155
cc_178 VPB SCD 0.00353385f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.245
cc_179 VPB N_CLK_c_580_n 0.00946347f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.245
cc_180 VPB N_CLK_c_586_n 0.0260162f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.64
cc_181 VPB N_A_1034_392#_c_664_n 0.0159033f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.64
cc_182 VPB N_A_1034_392#_c_665_n 0.020429f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.64
cc_183 VPB N_A_1034_392#_c_644_n 0.0132049f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.245
cc_184 VPB N_A_1034_392#_c_667_n 0.0607238f $X=-0.19 $Y=1.66 $X2=1.795 $Y2=1.575
cc_185 VPB N_A_1034_392#_c_668_n 0.00243629f $X=-0.19 $Y=1.66 $X2=2.51 $Y2=1.425
cc_186 VPB N_A_1034_392#_c_669_n 0.00144735f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.67
cc_187 VPB N_A_1034_392#_c_652_n 0.0019321f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=1.67
cc_188 VPB N_A_1034_392#_c_658_n 0.00116335f $X=-0.19 $Y=1.66 $X2=1.68 $Y2=1.662
cc_189 VPB N_A_1034_392#_c_672_n 0.00218598f $X=-0.19 $Y=1.66 $X2=1.795
+ $Y2=1.662
cc_190 VPB N_A_1034_392#_c_662_n 0.0177172f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_191 VPB N_A_1367_93#_c_871_n 0.0233517f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.245
cc_192 VPB N_A_1367_93#_c_872_n 0.0211965f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.64
cc_193 VPB N_A_1367_93#_c_865_n 0.00197089f $X=-0.19 $Y=1.66 $X2=2.65 $Y2=0.615
cc_194 VPB N_A_1367_93#_c_866_n 0.0231052f $X=-0.19 $Y=1.66 $X2=2.65 $Y2=0.615
cc_195 VPB N_A_1367_93#_c_875_n 0.00178601f $X=-0.19 $Y=1.66 $X2=2.51 $Y2=1.425
cc_196 VPB N_A_1367_93#_c_876_n 0.00224162f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_197 VPB N_A_1367_93#_c_870_n 0.00122099f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_198 VPB N_RESET_B_M1037_g 0.00778474f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.65
cc_199 VPB N_RESET_B_c_987_n 0.0402754f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.835
cc_200 VPB N_RESET_B_c_988_n 0.0302343f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.155
cc_201 VPB N_RESET_B_c_982_n 0.010477f $X=-0.19 $Y=1.66 $X2=2.65 $Y2=0.615
cc_202 VPB N_RESET_B_c_990_n 0.0167021f $X=-0.19 $Y=1.66 $X2=2.625 $Y2=0.9
cc_203 VPB N_RESET_B_c_984_n 0.00936563f $X=-0.19 $Y=1.66 $X2=2.535 $Y2=1.575
cc_204 VPB N_RESET_B_c_992_n 0.0136009f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_205 VPB N_RESET_B_c_993_n 0.0233932f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_206 VPB N_RESET_B_c_994_n 0.0216309f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_207 VPB N_RESET_B_c_995_n 0.0232387f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=1.67
cc_208 VPB N_RESET_B_c_996_n 0.00156846f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.67
cc_209 VPB N_RESET_B_c_997_n 0.0217281f $X=-0.19 $Y=1.66 $X2=2.51 $Y2=1.425
cc_210 VPB N_RESET_B_c_998_n 0.0020849f $X=-0.19 $Y=1.66 $X2=2.51 $Y2=1.26
cc_211 VPB N_RESET_B_c_999_n 0.00628945f $X=-0.19 $Y=1.66 $X2=1.2 $Y2=1.662
cc_212 VPB RESET_B 0.00299651f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_213 VPB N_RESET_B_c_1001_n 0.00803059f $X=-0.19 $Y=1.66 $X2=1.694 $Y2=1.662
cc_214 VPB N_RESET_B_c_1002_n 0.0598827f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_215 VPB N_RESET_B_c_1003_n 0.00324614f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_216 VPB N_RESET_B_c_1004_n 0.0327579f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_217 VPB N_A_1234_119#_c_1207_n 0.0164911f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.64
cc_218 VPB N_A_1234_119#_c_1216_n 0.015497f $X=-0.19 $Y=1.66 $X2=2.6 $Y2=1.26
cc_219 VPB N_A_1234_119#_c_1217_n 5.61498e-19 $X=-0.19 $Y=1.66 $X2=2.65
+ $Y2=0.615
cc_220 VPB N_A_1234_119#_c_1209_n 0.00733755f $X=-0.19 $Y=1.66 $X2=2.51
+ $Y2=1.425
cc_221 VPB N_A_1234_119#_c_1210_n 0.0125171f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_222 VPB N_A_1234_119#_c_1213_n 0.00754174f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_223 VPB N_A_1234_119#_c_1221_n 0.00112616f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=1.67
cc_224 VPB N_A_835_98#_c_1354_n 0.0162237f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.245
cc_225 VPB N_A_835_98#_c_1355_n 0.0722917f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.64
cc_226 VPB N_A_835_98#_c_1356_n 0.0597215f $X=-0.19 $Y=1.66 $X2=2.6 $Y2=1.05
cc_227 VPB N_A_835_98#_c_1357_n 0.0123764f $X=-0.19 $Y=1.66 $X2=2.6 $Y2=1.26
cc_228 VPB N_A_835_98#_c_1358_n 0.00781624f $X=-0.19 $Y=1.66 $X2=2.345 $Y2=1.575
cc_229 VPB N_A_835_98#_c_1359_n 0.0174462f $X=-0.19 $Y=1.66 $X2=1.795 $Y2=1.575
cc_230 VPB N_A_835_98#_c_1360_n 0.0158544f $X=-0.19 $Y=1.66 $X2=2.535 $Y2=1.425
cc_231 VPB N_A_835_98#_c_1361_n 0.187923f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_232 VPB N_A_835_98#_c_1362_n 0.0078517f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_233 VPB N_A_835_98#_c_1363_n 0.0132688f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_234 VPB N_A_835_98#_M1018_g 0.00887153f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_235 VPB N_A_835_98#_c_1345_n 0.0193138f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_236 VPB N_A_835_98#_c_1346_n 0.00438317f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_237 VPB N_A_835_98#_c_1367_n 0.0089865f $X=-0.19 $Y=1.66 $X2=2.51 $Y2=1.425
cc_238 VPB N_A_835_98#_c_1352_n 0.00789082f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_239 VPB N_A_835_98#_c_1353_n 0.0281488f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_240 VPB N_A_1997_272#_c_1544_n 0.0211446f $X=-0.19 $Y=1.66 $X2=1.005
+ $Y2=2.155
cc_241 VPB N_A_1997_272#_c_1555_n 0.0298064f $X=-0.19 $Y=1.66 $X2=1.005
+ $Y2=2.245
cc_242 VPB N_A_1997_272#_c_1556_n 0.0223998f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.64
cc_243 VPB N_A_1997_272#_c_1557_n 0.00909249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_244 VPB N_A_1997_272#_c_1552_n 0.00705302f $X=-0.19 $Y=1.66 $X2=0.495
+ $Y2=1.67
cc_245 VPB N_A_1745_74#_c_1661_n 0.00901615f $X=-0.19 $Y=1.66 $X2=1.005
+ $Y2=2.245
cc_246 VPB N_A_1745_74#_c_1672_n 0.0207522f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.64
cc_247 VPB N_A_1745_74#_c_1673_n 0.0222832f $X=-0.19 $Y=1.66 $X2=2.6 $Y2=1.05
cc_248 VPB N_A_1745_74#_c_1674_n 0.0425889f $X=-0.19 $Y=1.66 $X2=2.625 $Y2=0.9
cc_249 VPB N_A_1745_74#_c_1675_n 0.018388f $X=-0.19 $Y=1.66 $X2=2.345 $Y2=1.575
cc_250 VPB N_A_1745_74#_c_1676_n 0.00552913f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_251 VPB N_A_1745_74#_c_1677_n 0.00178486f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_252 VPB N_A_1745_74#_c_1666_n 0.00223832f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.67
cc_253 VPB N_A_1745_74#_c_1679_n 0.00730775f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=1.67
cc_254 VPB N_A_1745_74#_c_1680_n 0.00277122f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=1.67
cc_255 VPB N_A_1745_74#_c_1681_n 0.00536408f $X=-0.19 $Y=1.66 $X2=2.51 $Y2=1.425
cc_256 VPB N_A_2399_424#_c_1832_n 0.021165f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.245
cc_257 VPB N_A_2399_424#_c_1828_n 0.00855036f $X=-0.19 $Y=1.66 $X2=2.6 $Y2=1.05
cc_258 VPB N_A_2399_424#_c_1834_n 0.0138904f $X=-0.19 $Y=1.66 $X2=2.65 $Y2=0.615
cc_259 VPB N_A_2399_424#_c_1830_n 0.0133083f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.58
cc_260 VPB N_VPWR_c_1875_n 0.00651803f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_261 VPB N_VPWR_c_1876_n 0.00662228f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_262 VPB N_VPWR_c_1877_n 0.00396467f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_263 VPB N_VPWR_c_1878_n 0.0144445f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=1.67
cc_264 VPB N_VPWR_c_1879_n 0.02311f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=1.67
cc_265 VPB N_VPWR_c_1880_n 0.0144685f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_266 VPB N_VPWR_c_1881_n 0.0127921f $X=-0.19 $Y=1.66 $X2=1.2 $Y2=1.662
cc_267 VPB N_VPWR_c_1882_n 0.0158276f $X=-0.19 $Y=1.66 $X2=1.68 $Y2=1.665
cc_268 VPB N_VPWR_c_1883_n 0.0193772f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_269 VPB N_VPWR_c_1884_n 0.0352503f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_270 VPB N_VPWR_c_1885_n 0.00601569f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_271 VPB N_VPWR_c_1886_n 0.0523435f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_272 VPB N_VPWR_c_1887_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_273 VPB N_VPWR_c_1888_n 0.020808f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_274 VPB N_VPWR_c_1889_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_275 VPB N_VPWR_c_1890_n 0.0191515f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_276 VPB N_VPWR_c_1891_n 0.0596953f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_277 VPB N_VPWR_c_1892_n 0.0608368f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_278 VPB N_VPWR_c_1893_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_279 VPB N_VPWR_c_1894_n 0.0181474f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_280 VPB N_VPWR_c_1874_n 0.127177f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_281 VPB N_VPWR_c_1896_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_282 VPB N_VPWR_c_1897_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_283 VPB N_VPWR_c_1898_n 0.00443527f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_284 VPB N_VPWR_c_1899_n 0.00223798f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_285 VPB N_VPWR_c_1900_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_286 VPB N_A_300_464#_c_2049_n 0.00671604f $X=-0.19 $Y=1.66 $X2=2.6 $Y2=1.26
cc_287 VPB N_A_300_464#_c_2042_n 0.00666589f $X=-0.19 $Y=1.66 $X2=2.51 $Y2=1.425
cc_288 VPB N_A_300_464#_c_2051_n 8.30015e-19 $X=-0.19 $Y=1.66 $X2=2.535
+ $Y2=1.575
cc_289 VPB N_A_300_464#_c_2052_n 0.00843413f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_290 VPB N_A_300_464#_c_2053_n 0.00361747f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_291 VPB N_A_300_464#_c_2054_n 0.00289353f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=1.67
cc_292 VPB N_A_300_464#_c_2055_n 0.00709116f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.67
cc_293 VPB N_A_300_464#_c_2056_n 0.00189746f $X=-0.19 $Y=1.66 $X2=2.51 $Y2=1.425
cc_294 VPB N_A_300_464#_c_2047_n 0.00530074f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_295 VPB N_A_300_464#_c_2058_n 0.0025381f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_296 VPB N_A_300_464#_c_2059_n 0.00836287f $X=-0.19 $Y=1.66 $X2=1.694
+ $Y2=1.662
cc_297 VPB Q 0.0544732f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.64
cc_298 N_SCE_c_302_n N_A_27_88#_c_403_n 0.00644926f $X=2.345 $Y=1.575 $X2=0
+ $Y2=0
cc_299 N_SCE_c_303_n N_A_27_88#_c_403_n 0.00212198f $X=2.51 $Y=1.425 $X2=0 $Y2=0
cc_300 N_SCE_c_304_n N_A_27_88#_c_403_n 0.0178777f $X=2.51 $Y=1.425 $X2=0 $Y2=0
cc_301 N_SCE_M1033_g N_A_27_88#_c_396_n 0.00834942f $X=0.495 $Y=0.65 $X2=0 $Y2=0
cc_302 N_SCE_M1033_g N_A_27_88#_c_397_n 0.0131974f $X=0.495 $Y=0.65 $X2=0 $Y2=0
cc_303 N_SCE_c_305_n N_A_27_88#_c_397_n 0.0103131f $X=0.96 $Y=1.67 $X2=0 $Y2=0
cc_304 N_SCE_c_307_n N_A_27_88#_c_397_n 0.0273678f $X=1.623 $Y=1.662 $X2=0 $Y2=0
cc_305 N_SCE_c_309_n N_A_27_88#_c_405_n 0.0130468f $X=0.505 $Y=2.245 $X2=0 $Y2=0
cc_306 N_SCE_c_311_n N_A_27_88#_c_405_n 8.82207e-19 $X=1.005 $Y=2.245 $X2=0
+ $Y2=0
cc_307 N_SCE_M1033_g N_A_27_88#_c_398_n 0.0204376f $X=0.495 $Y=0.65 $X2=0 $Y2=0
cc_308 N_SCE_c_305_n N_A_27_88#_c_398_n 0.0032453f $X=0.96 $Y=1.67 $X2=0 $Y2=0
cc_309 N_SCE_c_307_n N_A_27_88#_c_398_n 0.0382971f $X=1.623 $Y=1.662 $X2=0 $Y2=0
cc_310 N_SCE_c_302_n N_A_27_88#_c_406_n 0.0233402f $X=2.345 $Y=1.575 $X2=0 $Y2=0
cc_311 N_SCE_c_303_n N_A_27_88#_c_407_n 0.0291709f $X=2.51 $Y=1.425 $X2=0 $Y2=0
cc_312 N_SCE_c_304_n N_A_27_88#_c_407_n 3.60884e-19 $X=2.51 $Y=1.425 $X2=0 $Y2=0
cc_313 N_SCE_c_308_n N_A_27_88#_c_408_n 0.00495347f $X=0.505 $Y=2.155 $X2=0
+ $Y2=0
cc_314 N_SCE_c_309_n N_A_27_88#_c_408_n 4.59028e-19 $X=0.505 $Y=2.245 $X2=0
+ $Y2=0
cc_315 N_SCE_M1033_g N_A_27_88#_c_400_n 7.61834e-19 $X=0.495 $Y=0.65 $X2=0 $Y2=0
cc_316 N_SCE_c_307_n N_A_27_88#_c_400_n 0.0212113f $X=1.623 $Y=1.662 $X2=0 $Y2=0
cc_317 N_SCE_M1033_g N_A_27_88#_c_401_n 0.00727818f $X=0.495 $Y=0.65 $X2=0 $Y2=0
cc_318 N_SCE_c_305_n N_A_27_88#_c_401_n 0.00441678f $X=0.96 $Y=1.67 $X2=0 $Y2=0
cc_319 N_SCE_c_307_n N_A_27_88#_c_401_n 0.008287f $X=1.623 $Y=1.662 $X2=0 $Y2=0
cc_320 N_SCE_c_308_n N_A_27_88#_c_409_n 0.00636452f $X=0.505 $Y=2.155 $X2=0
+ $Y2=0
cc_321 N_SCE_c_309_n N_A_27_88#_c_409_n 0.00700767f $X=0.505 $Y=2.245 $X2=0
+ $Y2=0
cc_322 N_SCE_c_310_n N_A_27_88#_c_409_n 0.00899514f $X=1.005 $Y=2.155 $X2=0
+ $Y2=0
cc_323 N_SCE_c_311_n N_A_27_88#_c_409_n 0.007641f $X=1.005 $Y=2.245 $X2=0 $Y2=0
cc_324 N_SCE_c_302_n N_A_27_88#_c_409_n 0.0109158f $X=2.345 $Y=1.575 $X2=0 $Y2=0
cc_325 N_SCE_c_305_n N_A_27_88#_c_409_n 0.00381149f $X=0.96 $Y=1.67 $X2=0 $Y2=0
cc_326 N_SCE_c_307_n N_A_27_88#_c_409_n 0.101415f $X=1.623 $Y=1.662 $X2=0 $Y2=0
cc_327 N_SCE_c_311_n N_D_c_485_n 0.0373647f $X=1.005 $Y=2.245 $X2=-0.19
+ $Y2=-0.245
cc_328 N_SCE_c_310_n N_D_c_479_n 0.0062192f $X=1.005 $Y=2.155 $X2=0 $Y2=0
cc_329 N_SCE_c_307_n N_D_c_479_n 0.00447951f $X=1.623 $Y=1.662 $X2=0 $Y2=0
cc_330 N_SCE_c_315_n N_D_c_479_n 0.00929488f $X=1.795 $Y=1.662 $X2=0 $Y2=0
cc_331 N_SCE_c_303_n N_D_c_480_n 0.00129438f $X=2.51 $Y=1.425 $X2=0 $Y2=0
cc_332 N_SCE_c_304_n N_D_c_480_n 0.00957253f $X=2.51 $Y=1.425 $X2=0 $Y2=0
cc_333 N_SCE_c_310_n N_D_c_487_n 0.0098871f $X=1.005 $Y=2.155 $X2=0 $Y2=0
cc_334 N_SCE_c_307_n N_D_c_487_n 0.00173212f $X=1.623 $Y=1.662 $X2=0 $Y2=0
cc_335 N_SCE_c_302_n N_D_c_481_n 0.00657898f $X=2.345 $Y=1.575 $X2=0 $Y2=0
cc_336 N_SCE_c_305_n N_D_c_481_n 0.00663484f $X=0.96 $Y=1.67 $X2=0 $Y2=0
cc_337 N_SCE_c_307_n N_D_c_481_n 0.00195725f $X=1.623 $Y=1.662 $X2=0 $Y2=0
cc_338 N_SCE_c_315_n N_D_c_481_n 0.0037388f $X=1.795 $Y=1.662 $X2=0 $Y2=0
cc_339 N_SCE_c_301_n N_D_c_482_n 0.00800462f $X=2.625 $Y=1.05 $X2=0 $Y2=0
cc_340 N_SCE_c_302_n N_D_c_482_n 0.00281358f $X=2.345 $Y=1.575 $X2=0 $Y2=0
cc_341 N_SCE_c_304_n N_D_c_482_n 3.01001e-19 $X=2.51 $Y=1.425 $X2=0 $Y2=0
cc_342 N_SCE_c_300_n N_D_c_483_n 2.00624e-19 $X=2.625 $Y=0.9 $X2=0 $Y2=0
cc_343 N_SCE_c_301_n N_D_c_483_n 2.26947e-19 $X=2.625 $Y=1.05 $X2=0 $Y2=0
cc_344 N_SCE_c_306_n N_D_c_483_n 9.5263e-19 $X=2.51 $Y=1.26 $X2=0 $Y2=0
cc_345 N_SCE_c_307_n N_D_c_483_n 0.0338107f $X=1.623 $Y=1.662 $X2=0 $Y2=0
cc_346 N_SCE_c_300_n N_D_c_484_n 0.00692407f $X=2.625 $Y=0.9 $X2=0 $Y2=0
cc_347 N_SCE_c_301_n N_D_c_484_n 5.10539e-19 $X=2.625 $Y=1.05 $X2=0 $Y2=0
cc_348 N_SCE_c_300_n N_SCD_M1012_g 0.0408623f $X=2.625 $Y=0.9 $X2=0 $Y2=0
cc_349 N_SCE_c_303_n N_SCD_M1012_g 0.00402266f $X=2.51 $Y=1.425 $X2=0 $Y2=0
cc_350 N_SCE_c_306_n N_SCD_M1012_g 0.0171335f $X=2.51 $Y=1.26 $X2=0 $Y2=0
cc_351 N_SCE_c_303_n SCD 0.0144929f $X=2.51 $Y=1.425 $X2=0 $Y2=0
cc_352 N_SCE_c_303_n N_SCD_c_539_n 0.002632f $X=2.51 $Y=1.425 $X2=0 $Y2=0
cc_353 N_SCE_c_304_n N_SCD_c_539_n 0.00936322f $X=2.51 $Y=1.425 $X2=0 $Y2=0
cc_354 N_SCE_c_309_n N_VPWR_c_1875_n 0.00657693f $X=0.505 $Y=2.245 $X2=0 $Y2=0
cc_355 N_SCE_c_311_n N_VPWR_c_1875_n 0.0146782f $X=1.005 $Y=2.245 $X2=0 $Y2=0
cc_356 N_SCE_c_309_n N_VPWR_c_1890_n 0.00445602f $X=0.505 $Y=2.245 $X2=0 $Y2=0
cc_357 N_SCE_c_311_n N_VPWR_c_1891_n 0.00413917f $X=1.005 $Y=2.245 $X2=0 $Y2=0
cc_358 N_SCE_c_309_n N_VPWR_c_1874_n 0.00860873f $X=0.505 $Y=2.245 $X2=0 $Y2=0
cc_359 N_SCE_c_311_n N_VPWR_c_1874_n 0.00817532f $X=1.005 $Y=2.245 $X2=0 $Y2=0
cc_360 N_SCE_c_311_n N_A_300_464#_c_2049_n 0.00181955f $X=1.005 $Y=2.245 $X2=0
+ $Y2=0
cc_361 N_SCE_c_301_n N_A_300_464#_c_2041_n 0.00703396f $X=2.625 $Y=1.05 $X2=0
+ $Y2=0
cc_362 N_SCE_c_303_n N_A_300_464#_c_2041_n 0.00943064f $X=2.51 $Y=1.425 $X2=0
+ $Y2=0
cc_363 N_SCE_c_306_n N_A_300_464#_c_2041_n 0.00186472f $X=2.51 $Y=1.26 $X2=0
+ $Y2=0
cc_364 N_SCE_c_300_n N_A_300_464#_c_2048_n 0.00663897f $X=2.625 $Y=0.9 $X2=0
+ $Y2=0
cc_365 N_SCE_c_301_n N_A_300_464#_c_2048_n 0.00472894f $X=2.625 $Y=1.05 $X2=0
+ $Y2=0
cc_366 N_SCE_c_302_n N_A_300_464#_c_2048_n 0.00336351f $X=2.345 $Y=1.575 $X2=0
+ $Y2=0
cc_367 N_SCE_c_303_n N_A_300_464#_c_2048_n 0.0208536f $X=2.51 $Y=1.425 $X2=0
+ $Y2=0
cc_368 N_SCE_c_304_n N_A_300_464#_c_2048_n 0.0013723f $X=2.51 $Y=1.425 $X2=0
+ $Y2=0
cc_369 N_SCE_c_306_n N_A_300_464#_c_2048_n 0.00193022f $X=2.51 $Y=1.26 $X2=0
+ $Y2=0
cc_370 N_SCE_M1033_g N_VGND_c_2231_n 0.0142996f $X=0.495 $Y=0.65 $X2=0 $Y2=0
cc_371 N_SCE_M1033_g N_VGND_c_2239_n 0.00438299f $X=0.495 $Y=0.65 $X2=0 $Y2=0
cc_372 N_SCE_c_300_n N_VGND_c_2240_n 9.15902e-19 $X=2.625 $Y=0.9 $X2=0 $Y2=0
cc_373 N_SCE_M1033_g N_VGND_c_2246_n 0.00439883f $X=0.495 $Y=0.65 $X2=0 $Y2=0
cc_374 N_SCE_c_300_n N_noxref_24_c_2364_n 0.0120947f $X=2.625 $Y=0.9 $X2=0 $Y2=0
cc_375 N_SCE_M1033_g N_noxref_24_c_2365_n 8.90151e-19 $X=0.495 $Y=0.65 $X2=0
+ $Y2=0
cc_376 N_SCE_c_300_n N_noxref_24_c_2366_n 0.001431f $X=2.625 $Y=0.9 $X2=0 $Y2=0
cc_377 N_A_27_88#_c_403_n N_D_c_479_n 0.0190261f $X=2.525 $Y=1.995 $X2=0 $Y2=0
cc_378 N_A_27_88#_c_406_n N_D_c_479_n 0.00102504f $X=2.207 $Y=2.002 $X2=0 $Y2=0
cc_379 N_A_27_88#_c_409_n N_D_c_479_n 0.00492692f $X=2.035 $Y=2.002 $X2=0 $Y2=0
cc_380 N_A_27_88#_c_409_n N_D_c_487_n 0.0190388f $X=2.035 $Y=2.002 $X2=0 $Y2=0
cc_381 N_A_27_88#_c_409_n N_D_c_481_n 7.9327e-19 $X=2.035 $Y=2.002 $X2=0 $Y2=0
cc_382 N_A_27_88#_c_403_n N_D_c_482_n 0.00133757f $X=2.525 $Y=1.995 $X2=0 $Y2=0
cc_383 N_A_27_88#_c_400_n N_D_c_482_n 2.69613e-19 $X=1.21 $Y=1.1 $X2=0 $Y2=0
cc_384 N_A_27_88#_c_401_n N_D_c_482_n 0.0143534f $X=1.21 $Y=1.1 $X2=0 $Y2=0
cc_385 N_A_27_88#_c_395_n N_D_c_483_n 0.00484268f $X=1.485 $Y=0.935 $X2=0 $Y2=0
cc_386 N_A_27_88#_c_400_n N_D_c_483_n 0.0250153f $X=1.21 $Y=1.1 $X2=0 $Y2=0
cc_387 N_A_27_88#_c_401_n N_D_c_483_n 0.0014755f $X=1.21 $Y=1.1 $X2=0 $Y2=0
cc_388 N_A_27_88#_c_395_n N_D_c_484_n 0.0356736f $X=1.485 $Y=0.935 $X2=0 $Y2=0
cc_389 N_A_27_88#_c_403_n N_SCD_c_537_n 0.0132707f $X=2.525 $Y=1.995 $X2=0 $Y2=0
cc_390 N_A_27_88#_c_407_n N_SCD_c_537_n 0.00290511f $X=2.51 $Y=1.995 $X2=0 $Y2=0
cc_391 N_A_27_88#_M1022_g N_SCD_c_541_n 0.0500024f $X=2.6 $Y=2.64 $X2=0 $Y2=0
cc_392 N_A_27_88#_c_403_n SCD 3.43581e-19 $X=2.525 $Y=1.995 $X2=0 $Y2=0
cc_393 N_A_27_88#_c_407_n SCD 0.0207487f $X=2.51 $Y=1.995 $X2=0 $Y2=0
cc_394 N_A_27_88#_c_405_n N_VPWR_c_1875_n 0.0246172f $X=0.28 $Y=2.465 $X2=0
+ $Y2=0
cc_395 N_A_27_88#_c_409_n N_VPWR_c_1875_n 0.0234317f $X=2.035 $Y=2.002 $X2=0
+ $Y2=0
cc_396 N_A_27_88#_M1022_g N_VPWR_c_1876_n 0.00139732f $X=2.6 $Y=2.64 $X2=0 $Y2=0
cc_397 N_A_27_88#_c_405_n N_VPWR_c_1890_n 0.0145938f $X=0.28 $Y=2.465 $X2=0
+ $Y2=0
cc_398 N_A_27_88#_M1022_g N_VPWR_c_1891_n 0.00427501f $X=2.6 $Y=2.64 $X2=0 $Y2=0
cc_399 N_A_27_88#_M1022_g N_VPWR_c_1874_n 0.00443648f $X=2.6 $Y=2.64 $X2=0 $Y2=0
cc_400 N_A_27_88#_c_405_n N_VPWR_c_1874_n 0.0120466f $X=0.28 $Y=2.465 $X2=0
+ $Y2=0
cc_401 N_A_27_88#_c_403_n N_A_300_464#_c_2049_n 0.0037654f $X=2.525 $Y=1.995
+ $X2=0 $Y2=0
cc_402 N_A_27_88#_c_409_n N_A_300_464#_c_2049_n 0.031029f $X=2.035 $Y=2.002
+ $X2=0 $Y2=0
cc_403 N_A_27_88#_M1022_g N_A_300_464#_c_2072_n 0.0081817f $X=2.6 $Y=2.64 $X2=0
+ $Y2=0
cc_404 N_A_27_88#_c_407_n N_A_300_464#_c_2072_n 0.031029f $X=2.51 $Y=1.995 $X2=0
+ $Y2=0
cc_405 N_A_27_88#_M1022_g N_A_300_464#_c_2058_n 0.0103508f $X=2.6 $Y=2.64 $X2=0
+ $Y2=0
cc_406 N_A_27_88#_c_406_n N_A_300_464#_c_2058_n 0.031029f $X=2.207 $Y=2.002
+ $X2=0 $Y2=0
cc_407 N_A_27_88#_c_395_n N_VGND_c_2231_n 0.00578639f $X=1.485 $Y=0.935 $X2=0
+ $Y2=0
cc_408 N_A_27_88#_c_396_n N_VGND_c_2231_n 0.0179429f $X=0.28 $Y=0.65 $X2=0 $Y2=0
cc_409 N_A_27_88#_c_398_n N_VGND_c_2231_n 0.0279517f $X=1.045 $Y=1.157 $X2=0
+ $Y2=0
cc_410 N_A_27_88#_c_396_n N_VGND_c_2239_n 0.00862619f $X=0.28 $Y=0.65 $X2=0
+ $Y2=0
cc_411 N_A_27_88#_c_395_n N_VGND_c_2240_n 9.09582e-19 $X=1.485 $Y=0.935 $X2=0
+ $Y2=0
cc_412 N_A_27_88#_c_396_n N_VGND_c_2246_n 0.00876292f $X=0.28 $Y=0.65 $X2=0
+ $Y2=0
cc_413 N_A_27_88#_c_395_n N_noxref_24_c_2364_n 0.0108727f $X=1.485 $Y=0.935
+ $X2=0 $Y2=0
cc_414 N_A_27_88#_c_395_n N_noxref_24_c_2365_n 0.00859442f $X=1.485 $Y=0.935
+ $X2=0 $Y2=0
cc_415 N_A_27_88#_c_400_n N_noxref_24_c_2365_n 0.0133426f $X=1.21 $Y=1.1 $X2=0
+ $Y2=0
cc_416 N_A_27_88#_c_401_n N_noxref_24_c_2365_n 0.0017694f $X=1.21 $Y=1.1 $X2=0
+ $Y2=0
cc_417 N_D_c_485_n N_VPWR_c_1875_n 0.00237824f $X=1.425 $Y=2.245 $X2=0 $Y2=0
cc_418 N_D_c_485_n N_VPWR_c_1891_n 0.00444483f $X=1.425 $Y=2.245 $X2=0 $Y2=0
cc_419 N_D_c_485_n N_VPWR_c_1874_n 0.00859301f $X=1.425 $Y=2.245 $X2=0 $Y2=0
cc_420 N_D_c_483_n N_A_300_464#_M1006_d 0.00160189f $X=1.935 $Y=1.1 $X2=-0.19
+ $Y2=-0.245
cc_421 N_D_c_485_n N_A_300_464#_c_2049_n 0.0115052f $X=1.425 $Y=2.245 $X2=0
+ $Y2=0
cc_422 N_D_c_487_n N_A_300_464#_c_2049_n 0.00629416f $X=1.425 $Y=2.16 $X2=0
+ $Y2=0
cc_423 N_D_c_482_n N_A_300_464#_c_2048_n 6.08332e-19 $X=1.935 $Y=1.1 $X2=0 $Y2=0
cc_424 N_D_c_483_n N_A_300_464#_c_2048_n 0.0234915f $X=1.935 $Y=1.1 $X2=0 $Y2=0
cc_425 N_D_c_484_n N_A_300_464#_c_2048_n 0.00517774f $X=1.935 $Y=0.935 $X2=0
+ $Y2=0
cc_426 N_D_c_484_n N_VGND_c_2240_n 9.15902e-19 $X=1.935 $Y=0.935 $X2=0 $Y2=0
cc_427 N_D_c_482_n N_noxref_24_c_2364_n 5.66605e-19 $X=1.935 $Y=1.1 $X2=0 $Y2=0
cc_428 N_D_c_483_n N_noxref_24_c_2364_n 0.0128576f $X=1.935 $Y=1.1 $X2=0 $Y2=0
cc_429 N_D_c_484_n N_noxref_24_c_2364_n 0.011902f $X=1.935 $Y=0.935 $X2=0 $Y2=0
cc_430 N_D_c_484_n N_noxref_24_c_2365_n 0.00113655f $X=1.935 $Y=0.935 $X2=0
+ $Y2=0
cc_431 N_D_c_483_n noxref_25 0.00198619f $X=1.935 $Y=1.1 $X2=-0.19 $Y2=-0.245
cc_432 N_SCD_M1012_g N_RESET_B_M1037_g 0.0329664f $X=3.04 $Y=0.615 $X2=0 $Y2=0
cc_433 SCD N_RESET_B_M1037_g 0.00424522f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_434 N_SCD_c_539_n N_RESET_B_M1037_g 0.0255034f $X=3.05 $Y=1.605 $X2=0 $Y2=0
cc_435 N_SCD_c_537_n N_RESET_B_c_988_n 0.0255034f $X=3.05 $Y=2.08 $X2=0 $Y2=0
cc_436 N_SCD_c_541_n N_RESET_B_c_994_n 0.0163311f $X=3.05 $Y=2.245 $X2=0 $Y2=0
cc_437 N_SCD_c_541_n N_VPWR_c_1876_n 0.0091757f $X=3.05 $Y=2.245 $X2=0 $Y2=0
cc_438 N_SCD_c_541_n N_VPWR_c_1891_n 0.00413917f $X=3.05 $Y=2.245 $X2=0 $Y2=0
cc_439 N_SCD_c_541_n N_VPWR_c_1874_n 0.00408796f $X=3.05 $Y=2.245 $X2=0 $Y2=0
cc_440 N_SCD_c_541_n N_A_300_464#_c_2072_n 0.0176382f $X=3.05 $Y=2.245 $X2=0
+ $Y2=0
cc_441 SCD N_A_300_464#_c_2072_n 0.0208238f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_442 N_SCD_M1012_g N_A_300_464#_c_2041_n 0.0123829f $X=3.04 $Y=0.615 $X2=0
+ $Y2=0
cc_443 SCD N_A_300_464#_c_2041_n 0.0149629f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_444 N_SCD_c_539_n N_A_300_464#_c_2041_n 0.00280161f $X=3.05 $Y=1.605 $X2=0
+ $Y2=0
cc_445 N_SCD_M1012_g N_A_300_464#_c_2042_n 0.00207067f $X=3.04 $Y=0.615 $X2=0
+ $Y2=0
cc_446 N_SCD_c_541_n N_A_300_464#_c_2042_n 0.00216808f $X=3.05 $Y=2.245 $X2=0
+ $Y2=0
cc_447 SCD N_A_300_464#_c_2042_n 0.0535746f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_448 N_SCD_c_539_n N_A_300_464#_c_2042_n 7.6448e-19 $X=3.05 $Y=1.605 $X2=0
+ $Y2=0
cc_449 N_SCD_c_541_n N_A_300_464#_c_2052_n 7.16633e-19 $X=3.05 $Y=2.245 $X2=0
+ $Y2=0
cc_450 N_SCD_c_541_n N_A_300_464#_c_2058_n 0.00170376f $X=3.05 $Y=2.245 $X2=0
+ $Y2=0
cc_451 N_SCD_M1012_g N_A_300_464#_c_2048_n 0.00135432f $X=3.04 $Y=0.615 $X2=0
+ $Y2=0
cc_452 N_SCD_M1012_g N_VGND_c_2240_n 9.09315e-19 $X=3.04 $Y=0.615 $X2=0 $Y2=0
cc_453 N_SCD_M1012_g N_noxref_24_c_2364_n 0.00698763f $X=3.04 $Y=0.615 $X2=0
+ $Y2=0
cc_454 N_SCD_M1012_g N_noxref_24_c_2366_n 0.01038f $X=3.04 $Y=0.615 $X2=0 $Y2=0
cc_455 N_CLK_c_586_n N_A_1034_392#_c_668_n 2.76703e-19 $X=4.62 $Y=1.885 $X2=0
+ $Y2=0
cc_456 N_CLK_c_579_n N_A_1034_392#_c_648_n 9.25509e-19 $X=4.595 $Y=1.41 $X2=0
+ $Y2=0
cc_457 N_CLK_c_583_n N_RESET_B_M1037_g 0.0424626f $X=3.95 $Y=1.115 $X2=0 $Y2=0
cc_458 N_CLK_c_584_n N_RESET_B_M1037_g 0.00119114f $X=3.95 $Y=1.115 $X2=0 $Y2=0
cc_459 N_CLK_c_579_n N_RESET_B_c_977_n 0.0100723f $X=4.595 $Y=1.41 $X2=0 $Y2=0
cc_460 N_CLK_c_583_n N_RESET_B_c_977_n 0.00359522f $X=3.95 $Y=1.115 $X2=0 $Y2=0
cc_461 N_CLK_c_584_n N_RESET_B_c_977_n 0.00490098f $X=3.95 $Y=1.115 $X2=0 $Y2=0
cc_462 N_CLK_c_578_n N_RESET_B_c_987_n 0.0213278f $X=4.115 $Y=1.515 $X2=0 $Y2=0
cc_463 N_CLK_c_586_n N_RESET_B_c_987_n 0.00545707f $X=4.62 $Y=1.885 $X2=0 $Y2=0
cc_464 N_CLK_c_584_n N_RESET_B_c_987_n 0.00126249f $X=3.95 $Y=1.115 $X2=0 $Y2=0
cc_465 CLK N_RESET_B_c_995_n 0.00643157f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_466 CLK N_RESET_B_c_996_n 0.00140609f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_467 N_CLK_c_584_n N_RESET_B_c_996_n 0.00301017f $X=3.95 $Y=1.115 $X2=0 $Y2=0
cc_468 N_CLK_c_578_n N_RESET_B_c_1001_n 7.57348e-19 $X=4.115 $Y=1.515 $X2=0
+ $Y2=0
cc_469 N_CLK_c_586_n N_RESET_B_c_1001_n 4.10028e-19 $X=4.62 $Y=1.885 $X2=0 $Y2=0
cc_470 N_CLK_c_584_n N_RESET_B_c_1001_n 0.0294475f $X=3.95 $Y=1.115 $X2=0 $Y2=0
cc_471 CLK N_A_835_98#_M1028_s 0.00369825f $X=3.995 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_472 N_CLK_c_586_n N_A_835_98#_c_1354_n 0.0374504f $X=4.62 $Y=1.885 $X2=0
+ $Y2=0
cc_473 N_CLK_c_579_n N_A_835_98#_c_1342_n 0.0210768f $X=4.595 $Y=1.41 $X2=0
+ $Y2=0
cc_474 N_CLK_c_579_n N_A_835_98#_c_1373_n 0.00608321f $X=4.595 $Y=1.41 $X2=0
+ $Y2=0
cc_475 N_CLK_c_579_n N_A_835_98#_c_1374_n 0.00991602f $X=4.595 $Y=1.41 $X2=0
+ $Y2=0
cc_476 CLK N_A_835_98#_c_1374_n 0.00756644f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_477 N_CLK_c_577_n N_A_835_98#_c_1376_n 3.39015e-19 $X=4.52 $Y=1.515 $X2=0
+ $Y2=0
cc_478 N_CLK_c_579_n N_A_835_98#_c_1376_n 0.00237757f $X=4.595 $Y=1.41 $X2=0
+ $Y2=0
cc_479 CLK N_A_835_98#_c_1376_n 0.00917328f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_480 N_CLK_c_583_n N_A_835_98#_c_1376_n 4.97991e-19 $X=3.95 $Y=1.115 $X2=0
+ $Y2=0
cc_481 N_CLK_c_584_n N_A_835_98#_c_1376_n 0.0149736f $X=3.95 $Y=1.115 $X2=0
+ $Y2=0
cc_482 N_CLK_c_579_n N_A_835_98#_c_1350_n 0.00320422f $X=4.595 $Y=1.41 $X2=0
+ $Y2=0
cc_483 N_CLK_c_581_n N_A_835_98#_c_1350_n 3.3312e-19 $X=4.62 $Y=1.515 $X2=0
+ $Y2=0
cc_484 CLK N_A_835_98#_c_1350_n 0.0151786f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_485 N_CLK_c_584_n N_A_835_98#_c_1350_n 0.00544275f $X=3.95 $Y=1.115 $X2=0
+ $Y2=0
cc_486 N_CLK_c_577_n N_A_835_98#_c_1351_n 7.23018e-19 $X=4.52 $Y=1.515 $X2=0
+ $Y2=0
cc_487 N_CLK_c_579_n N_A_835_98#_c_1351_n 0.00789222f $X=4.595 $Y=1.41 $X2=0
+ $Y2=0
cc_488 CLK N_A_835_98#_c_1351_n 0.0060775f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_489 N_CLK_c_584_n N_A_835_98#_c_1351_n 0.00509028f $X=3.95 $Y=1.115 $X2=0
+ $Y2=0
cc_490 N_CLK_c_577_n N_A_835_98#_c_1352_n 0.00128369f $X=4.52 $Y=1.515 $X2=0
+ $Y2=0
cc_491 N_CLK_c_581_n N_A_835_98#_c_1352_n 0.00595774f $X=4.62 $Y=1.515 $X2=0
+ $Y2=0
cc_492 N_CLK_c_586_n N_A_835_98#_c_1352_n 0.0197097f $X=4.62 $Y=1.885 $X2=0
+ $Y2=0
cc_493 CLK N_A_835_98#_c_1352_n 0.0398499f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_494 N_CLK_c_581_n N_A_835_98#_c_1353_n 0.0261211f $X=4.62 $Y=1.515 $X2=0
+ $Y2=0
cc_495 CLK N_A_835_98#_c_1353_n 2.04525e-19 $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_496 N_CLK_c_586_n N_VPWR_c_1877_n 0.0164315f $X=4.62 $Y=1.885 $X2=0 $Y2=0
cc_497 N_CLK_c_586_n N_VPWR_c_1884_n 0.00302783f $X=4.62 $Y=1.885 $X2=0 $Y2=0
cc_498 N_CLK_c_586_n N_VPWR_c_1874_n 0.00396658f $X=4.62 $Y=1.885 $X2=0 $Y2=0
cc_499 N_CLK_c_583_n N_A_300_464#_c_2041_n 8.58559e-19 $X=3.95 $Y=1.115 $X2=0
+ $Y2=0
cc_500 N_CLK_c_584_n N_A_300_464#_c_2041_n 0.0146802f $X=3.95 $Y=1.115 $X2=0
+ $Y2=0
cc_501 N_CLK_c_583_n N_A_300_464#_c_2042_n 0.0029155f $X=3.95 $Y=1.115 $X2=0
+ $Y2=0
cc_502 N_CLK_c_584_n N_A_300_464#_c_2042_n 0.0428479f $X=3.95 $Y=1.115 $X2=0
+ $Y2=0
cc_503 N_CLK_c_586_n N_A_300_464#_c_2051_n 0.0102356f $X=4.62 $Y=1.885 $X2=0
+ $Y2=0
cc_504 N_CLK_c_586_n N_A_300_464#_c_2052_n 5.41016e-19 $X=4.62 $Y=1.885 $X2=0
+ $Y2=0
cc_505 N_CLK_c_586_n N_A_300_464#_c_2053_n 0.00644616f $X=4.62 $Y=1.885 $X2=0
+ $Y2=0
cc_506 N_CLK_c_586_n N_A_300_464#_c_2059_n 0.00874826f $X=4.62 $Y=1.885 $X2=0
+ $Y2=0
cc_507 N_CLK_c_579_n N_VGND_c_2232_n 0.00165174f $X=4.595 $Y=1.41 $X2=0 $Y2=0
cc_508 N_CLK_c_583_n N_VGND_c_2232_n 4.3252e-19 $X=3.95 $Y=1.115 $X2=0 $Y2=0
cc_509 N_CLK_c_584_n N_VGND_c_2232_n 0.00858263f $X=3.95 $Y=1.115 $X2=0 $Y2=0
cc_510 N_CLK_c_579_n N_VGND_c_2233_n 0.0028517f $X=4.595 $Y=1.41 $X2=0 $Y2=0
cc_511 N_CLK_c_579_n N_VGND_c_2246_n 9.39239e-19 $X=4.595 $Y=1.41 $X2=0 $Y2=0
cc_512 N_A_1034_392#_c_655_n N_A_1367_93#_M1031_d 0.00176461f $X=9.065 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_513 N_A_1034_392#_M1000_g N_A_1367_93#_M1019_g 0.033412f $X=6.525 $Y=0.805
+ $X2=0 $Y2=0
cc_514 N_A_1034_392#_c_650_n N_A_1367_93#_M1019_g 0.00311064f $X=7.05 $Y=0.34
+ $X2=0 $Y2=0
cc_515 N_A_1034_392#_c_653_n N_A_1367_93#_M1019_g 0.00262964f $X=7.135 $Y=0.58
+ $X2=0 $Y2=0
cc_516 N_A_1034_392#_c_680_p N_A_1367_93#_M1019_g 0.0026982f $X=7.22 $Y=0.665
+ $X2=0 $Y2=0
cc_517 N_A_1034_392#_c_662_n N_A_1367_93#_c_871_n 5.85563e-19 $X=6.085 $Y=1.635
+ $X2=0 $Y2=0
cc_518 N_A_1034_392#_c_644_n N_A_1367_93#_c_866_n 0.033412f $X=6.45 $Y=1.635
+ $X2=0 $Y2=0
cc_519 N_A_1034_392#_c_662_n N_A_1367_93#_c_866_n 0.0010868f $X=6.085 $Y=1.635
+ $X2=0 $Y2=0
cc_520 N_A_1034_392#_c_654_n N_A_1367_93#_c_867_n 0.0520186f $X=7.93 $Y=0.665
+ $X2=0 $Y2=0
cc_521 N_A_1034_392#_c_655_n N_A_1367_93#_c_867_n 0.00353238f $X=9.065 $Y=0.34
+ $X2=0 $Y2=0
cc_522 N_A_1034_392#_c_654_n N_A_1367_93#_c_868_n 0.00761753f $X=7.93 $Y=0.665
+ $X2=0 $Y2=0
cc_523 N_A_1034_392#_c_680_p N_A_1367_93#_c_868_n 0.0103944f $X=7.22 $Y=0.665
+ $X2=0 $Y2=0
cc_524 N_A_1034_392#_c_658_n N_A_1367_93#_c_875_n 0.0139231f $X=9.33 $Y=2.125
+ $X2=0 $Y2=0
cc_525 N_A_1034_392#_c_663_n N_A_1367_93#_c_875_n 0.00323506f $X=9.085 $Y=1.105
+ $X2=0 $Y2=0
cc_526 N_A_1034_392#_c_646_n N_A_1367_93#_c_869_n 0.014712f $X=8.65 $Y=1.085
+ $X2=0 $Y2=0
cc_527 N_A_1034_392#_c_647_n N_A_1367_93#_c_869_n 0.00243289f $X=8.725 $Y=1.16
+ $X2=0 $Y2=0
cc_528 N_A_1034_392#_c_655_n N_A_1367_93#_c_869_n 0.0257761f $X=9.065 $Y=0.34
+ $X2=0 $Y2=0
cc_529 N_A_1034_392#_c_657_n N_A_1367_93#_c_869_n 0.0141828f $X=9.15 $Y=0.94
+ $X2=0 $Y2=0
cc_530 N_A_1034_392#_c_660_n N_A_1367_93#_c_869_n 5.79172e-19 $X=9.25 $Y=1.105
+ $X2=0 $Y2=0
cc_531 N_A_1034_392#_c_661_n N_A_1367_93#_c_869_n 0.0131302f $X=9.33 $Y=1.105
+ $X2=0 $Y2=0
cc_532 N_A_1034_392#_c_663_n N_A_1367_93#_c_869_n 0.00313966f $X=9.085 $Y=1.105
+ $X2=0 $Y2=0
cc_533 N_A_1034_392#_c_658_n N_A_1367_93#_c_870_n 0.0197161f $X=9.33 $Y=2.125
+ $X2=0 $Y2=0
cc_534 N_A_1034_392#_c_660_n N_A_1367_93#_c_870_n 2.26254e-19 $X=9.25 $Y=1.105
+ $X2=0 $Y2=0
cc_535 N_A_1034_392#_c_661_n N_A_1367_93#_c_870_n 0.0131446f $X=9.33 $Y=1.105
+ $X2=0 $Y2=0
cc_536 N_A_1034_392#_c_663_n N_A_1367_93#_c_870_n 0.00960948f $X=9.085 $Y=1.105
+ $X2=0 $Y2=0
cc_537 N_A_1034_392#_M1000_g N_RESET_B_c_977_n 0.00882199f $X=6.525 $Y=0.805
+ $X2=0 $Y2=0
cc_538 N_A_1034_392#_c_650_n N_RESET_B_c_977_n 0.0294278f $X=7.05 $Y=0.34 $X2=0
+ $Y2=0
cc_539 N_A_1034_392#_c_651_n N_RESET_B_c_977_n 0.00992957f $X=5.62 $Y=0.34 $X2=0
+ $Y2=0
cc_540 N_A_1034_392#_c_650_n N_RESET_B_M1007_g 0.00466687f $X=7.05 $Y=0.34 $X2=0
+ $Y2=0
cc_541 N_A_1034_392#_c_653_n N_RESET_B_M1007_g 0.00445709f $X=7.135 $Y=0.58
+ $X2=0 $Y2=0
cc_542 N_A_1034_392#_c_654_n N_RESET_B_M1007_g 0.0128143f $X=7.93 $Y=0.665 $X2=0
+ $Y2=0
cc_543 N_A_1034_392#_c_707_p N_RESET_B_M1007_g 0.0035287f $X=8.015 $Y=0.58 $X2=0
+ $Y2=0
cc_544 N_A_1034_392#_c_656_n N_RESET_B_M1007_g 6.46496e-19 $X=8.1 $Y=0.34 $X2=0
+ $Y2=0
cc_545 N_A_1034_392#_c_664_n N_RESET_B_c_995_n 0.00340123f $X=6.135 $Y=2.12
+ $X2=0 $Y2=0
cc_546 N_A_1034_392#_c_644_n N_RESET_B_c_995_n 0.00373244f $X=6.45 $Y=1.635
+ $X2=0 $Y2=0
cc_547 N_A_1034_392#_c_668_n N_RESET_B_c_995_n 0.0144672f $X=5.45 $Y=2.085 $X2=0
+ $Y2=0
cc_548 N_A_1034_392#_c_669_n N_RESET_B_c_995_n 0.017308f $X=5.63 $Y=1.71 $X2=0
+ $Y2=0
cc_549 N_A_1034_392#_c_652_n N_RESET_B_c_995_n 0.0161553f $X=6.085 $Y=1.71 $X2=0
+ $Y2=0
cc_550 N_A_1034_392#_c_662_n N_RESET_B_c_995_n 0.00379596f $X=6.085 $Y=1.635
+ $X2=0 $Y2=0
cc_551 N_A_1034_392#_c_667_n N_RESET_B_c_997_n 0.00642678f $X=9.89 $Y=2.465
+ $X2=0 $Y2=0
cc_552 N_A_1034_392#_c_658_n N_RESET_B_c_997_n 0.0173785f $X=9.33 $Y=2.125 $X2=0
+ $Y2=0
cc_553 N_A_1034_392#_c_672_n N_RESET_B_c_997_n 0.0197423f $X=9.81 $Y=2.215 $X2=0
+ $Y2=0
cc_554 N_A_1034_392#_c_646_n N_A_1234_119#_M1031_g 0.0286306f $X=8.65 $Y=1.085
+ $X2=0 $Y2=0
cc_555 N_A_1034_392#_c_655_n N_A_1234_119#_M1031_g 0.0116373f $X=9.065 $Y=0.34
+ $X2=0 $Y2=0
cc_556 N_A_1034_392#_c_647_n N_A_1234_119#_c_1207_n 0.0152066f $X=8.725 $Y=1.16
+ $X2=0 $Y2=0
cc_557 N_A_1034_392#_c_658_n N_A_1234_119#_c_1207_n 4.45404e-19 $X=9.33 $Y=2.125
+ $X2=0 $Y2=0
cc_558 N_A_1034_392#_c_665_n N_A_1234_119#_c_1217_n 0.00187655f $X=6.135 $Y=2.21
+ $X2=0 $Y2=0
cc_559 N_A_1034_392#_c_644_n N_A_1234_119#_c_1217_n 7.28544e-19 $X=6.45 $Y=1.635
+ $X2=0 $Y2=0
cc_560 N_A_1034_392#_M1000_g N_A_1234_119#_c_1208_n 0.0102762f $X=6.525 $Y=0.805
+ $X2=0 $Y2=0
cc_561 N_A_1034_392#_c_650_n N_A_1234_119#_c_1208_n 0.0118472f $X=7.05 $Y=0.34
+ $X2=0 $Y2=0
cc_562 N_A_1034_392#_c_664_n N_A_1234_119#_c_1209_n 6.14864e-19 $X=6.135 $Y=2.12
+ $X2=0 $Y2=0
cc_563 N_A_1034_392#_c_665_n N_A_1234_119#_c_1209_n 3.40922e-19 $X=6.135 $Y=2.21
+ $X2=0 $Y2=0
cc_564 N_A_1034_392#_M1000_g N_A_1234_119#_c_1209_n 0.00689529f $X=6.525
+ $Y=0.805 $X2=0 $Y2=0
cc_565 N_A_1034_392#_c_644_n N_A_1234_119#_c_1214_n 5.90653e-19 $X=6.45 $Y=1.635
+ $X2=0 $Y2=0
cc_566 N_A_1034_392#_M1000_g N_A_1234_119#_c_1214_n 0.00636651f $X=6.525
+ $Y=0.805 $X2=0 $Y2=0
cc_567 N_A_1034_392#_c_650_n N_A_1234_119#_c_1214_n 0.019863f $X=7.05 $Y=0.34
+ $X2=0 $Y2=0
cc_568 N_A_1034_392#_c_680_p N_A_1234_119#_c_1214_n 0.00486547f $X=7.22 $Y=0.665
+ $X2=0 $Y2=0
cc_569 N_A_1034_392#_c_668_n N_A_835_98#_c_1354_n 0.00260802f $X=5.45 $Y=2.085
+ $X2=0 $Y2=0
cc_570 N_A_1034_392#_c_669_n N_A_835_98#_c_1354_n 6.43092e-19 $X=5.63 $Y=1.71
+ $X2=0 $Y2=0
cc_571 N_A_1034_392#_c_648_n N_A_835_98#_c_1342_n 0.00994075f $X=5.36 $Y=0.78
+ $X2=0 $Y2=0
cc_572 N_A_1034_392#_c_649_n N_A_835_98#_c_1342_n 8.65367e-19 $X=5.54 $Y=1.545
+ $X2=0 $Y2=0
cc_573 N_A_1034_392#_c_659_n N_A_835_98#_c_1342_n 0.00190639f $X=5.422 $Y=1.285
+ $X2=0 $Y2=0
cc_574 N_A_1034_392#_c_664_n N_A_835_98#_c_1355_n 0.0111158f $X=6.135 $Y=2.12
+ $X2=0 $Y2=0
cc_575 N_A_1034_392#_c_665_n N_A_835_98#_c_1355_n 0.0130881f $X=6.135 $Y=2.21
+ $X2=0 $Y2=0
cc_576 N_A_1034_392#_c_668_n N_A_835_98#_c_1355_n 4.97235e-19 $X=5.45 $Y=2.085
+ $X2=0 $Y2=0
cc_577 N_A_1034_392#_c_669_n N_A_835_98#_c_1355_n 0.0104193f $X=5.63 $Y=1.71
+ $X2=0 $Y2=0
cc_578 N_A_1034_392#_c_665_n N_A_835_98#_c_1356_n 0.00899632f $X=6.135 $Y=2.21
+ $X2=0 $Y2=0
cc_579 N_A_1034_392#_c_650_n N_A_835_98#_c_1343_n 0.00139627f $X=7.05 $Y=0.34
+ $X2=0 $Y2=0
cc_580 N_A_1034_392#_c_652_n N_A_835_98#_c_1343_n 0.00441445f $X=6.085 $Y=1.71
+ $X2=0 $Y2=0
cc_581 N_A_1034_392#_c_662_n N_A_835_98#_c_1343_n 0.0160947f $X=6.085 $Y=1.635
+ $X2=0 $Y2=0
cc_582 N_A_1034_392#_M1000_g N_A_835_98#_c_1344_n 0.0223555f $X=6.525 $Y=0.805
+ $X2=0 $Y2=0
cc_583 N_A_1034_392#_c_648_n N_A_835_98#_c_1344_n 0.00472785f $X=5.36 $Y=0.78
+ $X2=0 $Y2=0
cc_584 N_A_1034_392#_c_650_n N_A_835_98#_c_1344_n 0.00330666f $X=7.05 $Y=0.34
+ $X2=0 $Y2=0
cc_585 N_A_1034_392#_c_665_n N_A_835_98#_c_1358_n 0.00151278f $X=6.135 $Y=2.21
+ $X2=0 $Y2=0
cc_586 N_A_1034_392#_c_665_n N_A_835_98#_c_1360_n 0.0132738f $X=6.135 $Y=2.21
+ $X2=0 $Y2=0
cc_587 N_A_1034_392#_c_644_n N_A_835_98#_c_1360_n 0.00109872f $X=6.45 $Y=1.635
+ $X2=0 $Y2=0
cc_588 N_A_1034_392#_c_667_n N_A_835_98#_c_1362_n 0.00644632f $X=9.89 $Y=2.465
+ $X2=0 $Y2=0
cc_589 N_A_1034_392#_c_667_n N_A_835_98#_M1018_g 0.0153501f $X=9.89 $Y=2.465
+ $X2=0 $Y2=0
cc_590 N_A_1034_392#_c_658_n N_A_835_98#_M1018_g 0.00856179f $X=9.33 $Y=2.125
+ $X2=0 $Y2=0
cc_591 N_A_1034_392#_c_667_n N_A_835_98#_c_1345_n 0.00418242f $X=9.89 $Y=2.465
+ $X2=0 $Y2=0
cc_592 N_A_1034_392#_c_658_n N_A_835_98#_c_1345_n 0.0121351f $X=9.33 $Y=2.125
+ $X2=0 $Y2=0
cc_593 N_A_1034_392#_c_672_n N_A_835_98#_c_1345_n 0.00479207f $X=9.81 $Y=2.215
+ $X2=0 $Y2=0
cc_594 N_A_1034_392#_c_660_n N_A_835_98#_c_1346_n 0.019069f $X=9.25 $Y=1.105
+ $X2=0 $Y2=0
cc_595 N_A_1034_392#_c_661_n N_A_835_98#_c_1346_n 0.00163879f $X=9.33 $Y=1.105
+ $X2=0 $Y2=0
cc_596 N_A_1034_392#_c_663_n N_A_835_98#_c_1346_n 0.00141289f $X=9.085 $Y=1.105
+ $X2=0 $Y2=0
cc_597 N_A_1034_392#_c_658_n N_A_835_98#_c_1347_n 0.00153175f $X=9.33 $Y=2.125
+ $X2=0 $Y2=0
cc_598 N_A_1034_392#_c_655_n N_A_835_98#_M1002_g 0.00301232f $X=9.065 $Y=0.34
+ $X2=0 $Y2=0
cc_599 N_A_1034_392#_c_657_n N_A_835_98#_M1002_g 0.00129859f $X=9.15 $Y=0.94
+ $X2=0 $Y2=0
cc_600 N_A_1034_392#_c_660_n N_A_835_98#_M1002_g 0.00125371f $X=9.25 $Y=1.105
+ $X2=0 $Y2=0
cc_601 N_A_1034_392#_c_660_n N_A_835_98#_c_1349_n 0.0194128f $X=9.25 $Y=1.105
+ $X2=0 $Y2=0
cc_602 N_A_1034_392#_c_661_n N_A_835_98#_c_1349_n 3.65519e-19 $X=9.33 $Y=1.105
+ $X2=0 $Y2=0
cc_603 N_A_1034_392#_c_649_n N_A_835_98#_c_1350_n 0.00564461f $X=5.54 $Y=1.545
+ $X2=0 $Y2=0
cc_604 N_A_1034_392#_c_668_n N_A_835_98#_c_1352_n 0.0196012f $X=5.45 $Y=2.085
+ $X2=0 $Y2=0
cc_605 N_A_1034_392#_c_649_n N_A_835_98#_c_1352_n 0.0237013f $X=5.54 $Y=1.545
+ $X2=0 $Y2=0
cc_606 N_A_1034_392#_c_669_n N_A_835_98#_c_1352_n 0.00652762f $X=5.63 $Y=1.71
+ $X2=0 $Y2=0
cc_607 N_A_1034_392#_c_659_n N_A_835_98#_c_1352_n 0.00267749f $X=5.422 $Y=1.285
+ $X2=0 $Y2=0
cc_608 N_A_1034_392#_c_668_n N_A_835_98#_c_1353_n 0.00634613f $X=5.45 $Y=2.085
+ $X2=0 $Y2=0
cc_609 N_A_1034_392#_c_649_n N_A_835_98#_c_1353_n 0.0141907f $X=5.54 $Y=1.545
+ $X2=0 $Y2=0
cc_610 N_A_1034_392#_c_650_n N_A_835_98#_c_1353_n 0.00385788f $X=7.05 $Y=0.34
+ $X2=0 $Y2=0
cc_611 N_A_1034_392#_c_669_n N_A_835_98#_c_1353_n 0.0120447f $X=5.63 $Y=1.71
+ $X2=0 $Y2=0
cc_612 N_A_1034_392#_c_652_n N_A_835_98#_c_1353_n 0.0116804f $X=6.085 $Y=1.71
+ $X2=0 $Y2=0
cc_613 N_A_1034_392#_c_659_n N_A_835_98#_c_1353_n 0.0122529f $X=5.422 $Y=1.285
+ $X2=0 $Y2=0
cc_614 N_A_1034_392#_c_662_n N_A_835_98#_c_1353_n 0.021574f $X=6.085 $Y=1.635
+ $X2=0 $Y2=0
cc_615 N_A_1034_392#_c_667_n N_A_1997_272#_c_1555_n 0.0218756f $X=9.89 $Y=2.465
+ $X2=0 $Y2=0
cc_616 N_A_1034_392#_c_672_n N_A_1997_272#_c_1555_n 2.75032e-19 $X=9.81 $Y=2.215
+ $X2=0 $Y2=0
cc_617 N_A_1034_392#_c_667_n N_A_1997_272#_c_1556_n 0.0293409f $X=9.89 $Y=2.465
+ $X2=0 $Y2=0
cc_618 N_A_1034_392#_c_655_n N_A_1745_74#_M1003_d 0.00630965f $X=9.065 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_619 N_A_1034_392#_c_657_n N_A_1745_74#_M1003_d 0.0113887f $X=9.15 $Y=0.94
+ $X2=-0.19 $Y2=-0.245
cc_620 N_A_1034_392#_c_658_n N_A_1745_74#_M1018_d 0.00749069f $X=9.33 $Y=2.125
+ $X2=0 $Y2=0
cc_621 N_A_1034_392#_c_785_p N_A_1745_74#_M1018_d 0.0039098f $X=9.415 $Y=2.252
+ $X2=0 $Y2=0
cc_622 N_A_1034_392#_c_672_n N_A_1745_74#_M1018_d 0.00176657f $X=9.81 $Y=2.215
+ $X2=0 $Y2=0
cc_623 N_A_1034_392#_c_667_n N_A_1745_74#_c_1677_n 0.0220662f $X=9.89 $Y=2.465
+ $X2=0 $Y2=0
cc_624 N_A_1034_392#_c_785_p N_A_1745_74#_c_1677_n 0.0101735f $X=9.415 $Y=2.252
+ $X2=0 $Y2=0
cc_625 N_A_1034_392#_c_672_n N_A_1745_74#_c_1677_n 0.0386883f $X=9.81 $Y=2.215
+ $X2=0 $Y2=0
cc_626 N_A_1034_392#_c_657_n N_A_1745_74#_c_1665_n 0.00768735f $X=9.15 $Y=0.94
+ $X2=0 $Y2=0
cc_627 N_A_1034_392#_c_660_n N_A_1745_74#_c_1665_n 4.55554e-19 $X=9.25 $Y=1.105
+ $X2=0 $Y2=0
cc_628 N_A_1034_392#_c_661_n N_A_1745_74#_c_1665_n 0.0116456f $X=9.33 $Y=1.105
+ $X2=0 $Y2=0
cc_629 N_A_1034_392#_c_658_n N_A_1745_74#_c_1666_n 0.0375442f $X=9.33 $Y=2.125
+ $X2=0 $Y2=0
cc_630 N_A_1034_392#_c_667_n N_A_1745_74#_c_1679_n 0.00443076f $X=9.89 $Y=2.465
+ $X2=0 $Y2=0
cc_631 N_A_1034_392#_c_672_n N_A_1745_74#_c_1679_n 0.0125258f $X=9.81 $Y=2.215
+ $X2=0 $Y2=0
cc_632 N_A_1034_392#_c_667_n N_A_1745_74#_c_1680_n 9.16255e-19 $X=9.89 $Y=2.465
+ $X2=0 $Y2=0
cc_633 N_A_1034_392#_c_658_n N_A_1745_74#_c_1680_n 0.0141314f $X=9.33 $Y=2.125
+ $X2=0 $Y2=0
cc_634 N_A_1034_392#_c_672_n N_A_1745_74#_c_1680_n 0.0111216f $X=9.81 $Y=2.215
+ $X2=0 $Y2=0
cc_635 N_A_1034_392#_c_667_n N_A_1745_74#_c_1681_n 0.0062593f $X=9.89 $Y=2.465
+ $X2=0 $Y2=0
cc_636 N_A_1034_392#_c_672_n N_A_1745_74#_c_1681_n 0.0202186f $X=9.81 $Y=2.215
+ $X2=0 $Y2=0
cc_637 N_A_1034_392#_c_646_n N_A_1745_74#_c_1667_n 5.77109e-19 $X=8.65 $Y=1.085
+ $X2=0 $Y2=0
cc_638 N_A_1034_392#_c_655_n N_A_1745_74#_c_1667_n 0.00648023f $X=9.065 $Y=0.34
+ $X2=0 $Y2=0
cc_639 N_A_1034_392#_c_657_n N_A_1745_74#_c_1667_n 0.0264512f $X=9.15 $Y=0.94
+ $X2=0 $Y2=0
cc_640 N_A_1034_392#_c_660_n N_A_1745_74#_c_1667_n 2.06488e-19 $X=9.25 $Y=1.105
+ $X2=0 $Y2=0
cc_641 N_A_1034_392#_c_661_n N_A_1745_74#_c_1667_n 7.15367e-19 $X=9.33 $Y=1.105
+ $X2=0 $Y2=0
cc_642 N_A_1034_392#_c_660_n N_A_1745_74#_c_1668_n 6.39686e-19 $X=9.25 $Y=1.105
+ $X2=0 $Y2=0
cc_643 N_A_1034_392#_c_661_n N_A_1745_74#_c_1668_n 0.0144646f $X=9.33 $Y=1.105
+ $X2=0 $Y2=0
cc_644 N_A_1034_392#_c_667_n N_VPWR_c_1886_n 0.00304676f $X=9.89 $Y=2.465 $X2=0
+ $Y2=0
cc_645 N_A_1034_392#_c_665_n N_VPWR_c_1874_n 9.49986e-19 $X=6.135 $Y=2.21 $X2=0
+ $Y2=0
cc_646 N_A_1034_392#_c_667_n N_VPWR_c_1874_n 0.00375875f $X=9.89 $Y=2.465 $X2=0
+ $Y2=0
cc_647 N_A_1034_392#_M1030_d N_A_300_464#_c_2053_n 0.00695361f $X=5.17 $Y=1.96
+ $X2=0 $Y2=0
cc_648 N_A_1034_392#_c_668_n N_A_300_464#_c_2053_n 0.016647f $X=5.45 $Y=2.085
+ $X2=0 $Y2=0
cc_649 N_A_1034_392#_c_669_n N_A_300_464#_c_2053_n 0.0134529f $X=5.63 $Y=1.71
+ $X2=0 $Y2=0
cc_650 N_A_1034_392#_c_652_n N_A_300_464#_c_2053_n 0.0029069f $X=6.085 $Y=1.71
+ $X2=0 $Y2=0
cc_651 N_A_1034_392#_c_648_n N_A_300_464#_c_2043_n 0.0311322f $X=5.36 $Y=0.78
+ $X2=0 $Y2=0
cc_652 N_A_1034_392#_c_650_n N_A_300_464#_c_2043_n 0.013349f $X=7.05 $Y=0.34
+ $X2=0 $Y2=0
cc_653 N_A_1034_392#_M1000_g N_A_300_464#_c_2044_n 3.66002e-19 $X=6.525 $Y=0.805
+ $X2=0 $Y2=0
cc_654 N_A_1034_392#_c_648_n N_A_300_464#_c_2044_n 0.00571418f $X=5.36 $Y=0.78
+ $X2=0 $Y2=0
cc_655 N_A_1034_392#_c_659_n N_A_300_464#_c_2044_n 0.00980399f $X=5.422 $Y=1.285
+ $X2=0 $Y2=0
cc_656 N_A_1034_392#_c_665_n N_A_300_464#_c_2054_n 0.00798244f $X=6.135 $Y=2.21
+ $X2=0 $Y2=0
cc_657 N_A_1034_392#_M1000_g N_A_300_464#_c_2045_n 0.00615688f $X=6.525 $Y=0.805
+ $X2=0 $Y2=0
cc_658 N_A_1034_392#_c_652_n N_A_300_464#_c_2045_n 0.0160606f $X=6.085 $Y=1.71
+ $X2=0 $Y2=0
cc_659 N_A_1034_392#_c_662_n N_A_300_464#_c_2045_n 0.00626971f $X=6.085 $Y=1.635
+ $X2=0 $Y2=0
cc_660 N_A_1034_392#_c_652_n N_A_300_464#_c_2046_n 0.0145081f $X=6.085 $Y=1.71
+ $X2=0 $Y2=0
cc_661 N_A_1034_392#_c_659_n N_A_300_464#_c_2046_n 0.0135231f $X=5.422 $Y=1.285
+ $X2=0 $Y2=0
cc_662 N_A_1034_392#_c_662_n N_A_300_464#_c_2046_n 3.38485e-19 $X=6.085 $Y=1.635
+ $X2=0 $Y2=0
cc_663 N_A_1034_392#_c_664_n N_A_300_464#_c_2055_n 0.00392277f $X=6.135 $Y=2.12
+ $X2=0 $Y2=0
cc_664 N_A_1034_392#_c_665_n N_A_300_464#_c_2055_n 0.00875358f $X=6.135 $Y=2.21
+ $X2=0 $Y2=0
cc_665 N_A_1034_392#_c_644_n N_A_300_464#_c_2055_n 0.00224934f $X=6.45 $Y=1.635
+ $X2=0 $Y2=0
cc_666 N_A_1034_392#_c_652_n N_A_300_464#_c_2055_n 0.00770757f $X=6.085 $Y=1.71
+ $X2=0 $Y2=0
cc_667 N_A_1034_392#_c_662_n N_A_300_464#_c_2055_n 6.46491e-19 $X=6.085 $Y=1.635
+ $X2=0 $Y2=0
cc_668 N_A_1034_392#_c_664_n N_A_300_464#_c_2056_n 0.00121768f $X=6.135 $Y=2.12
+ $X2=0 $Y2=0
cc_669 N_A_1034_392#_c_665_n N_A_300_464#_c_2056_n 0.00154832f $X=6.135 $Y=2.21
+ $X2=0 $Y2=0
cc_670 N_A_1034_392#_c_669_n N_A_300_464#_c_2056_n 0.0116978f $X=5.63 $Y=1.71
+ $X2=0 $Y2=0
cc_671 N_A_1034_392#_c_652_n N_A_300_464#_c_2056_n 0.016874f $X=6.085 $Y=1.71
+ $X2=0 $Y2=0
cc_672 N_A_1034_392#_c_662_n N_A_300_464#_c_2056_n 0.00278662f $X=6.085 $Y=1.635
+ $X2=0 $Y2=0
cc_673 N_A_1034_392#_c_664_n N_A_300_464#_c_2047_n 0.00549102f $X=6.135 $Y=2.12
+ $X2=0 $Y2=0
cc_674 N_A_1034_392#_c_644_n N_A_300_464#_c_2047_n 0.0116747f $X=6.45 $Y=1.635
+ $X2=0 $Y2=0
cc_675 N_A_1034_392#_M1000_g N_A_300_464#_c_2047_n 0.00522785f $X=6.525 $Y=0.805
+ $X2=0 $Y2=0
cc_676 N_A_1034_392#_c_652_n N_A_300_464#_c_2047_n 0.025176f $X=6.085 $Y=1.71
+ $X2=0 $Y2=0
cc_677 N_A_1034_392#_c_662_n N_A_300_464#_c_2047_n 0.00170375f $X=6.085 $Y=1.635
+ $X2=0 $Y2=0
cc_678 N_A_1034_392#_c_654_n N_VGND_M1007_d 0.0170064f $X=7.93 $Y=0.665 $X2=0
+ $Y2=0
cc_679 N_A_1034_392#_c_707_p N_VGND_M1007_d 0.00275919f $X=8.015 $Y=0.58 $X2=0
+ $Y2=0
cc_680 N_A_1034_392#_c_656_n N_VGND_M1007_d 7.93589e-19 $X=8.1 $Y=0.34 $X2=0
+ $Y2=0
cc_681 N_A_1034_392#_c_648_n N_VGND_c_2233_n 0.0189029f $X=5.36 $Y=0.78 $X2=0
+ $Y2=0
cc_682 N_A_1034_392#_c_651_n N_VGND_c_2233_n 0.0144411f $X=5.62 $Y=0.34 $X2=0
+ $Y2=0
cc_683 N_A_1034_392#_c_650_n N_VGND_c_2241_n 0.103356f $X=7.05 $Y=0.34 $X2=0
+ $Y2=0
cc_684 N_A_1034_392#_c_651_n N_VGND_c_2241_n 0.0276098f $X=5.62 $Y=0.34 $X2=0
+ $Y2=0
cc_685 N_A_1034_392#_c_654_n N_VGND_c_2241_n 0.00402072f $X=7.93 $Y=0.665 $X2=0
+ $Y2=0
cc_686 N_A_1034_392#_c_646_n N_VGND_c_2242_n 0.00278271f $X=8.65 $Y=1.085 $X2=0
+ $Y2=0
cc_687 N_A_1034_392#_c_654_n N_VGND_c_2242_n 0.00335833f $X=7.93 $Y=0.665 $X2=0
+ $Y2=0
cc_688 N_A_1034_392#_c_655_n N_VGND_c_2242_n 0.0734255f $X=9.065 $Y=0.34 $X2=0
+ $Y2=0
cc_689 N_A_1034_392#_c_656_n N_VGND_c_2242_n 0.0118998f $X=8.1 $Y=0.34 $X2=0
+ $Y2=0
cc_690 N_A_1034_392#_c_646_n N_VGND_c_2246_n 0.00358525f $X=8.65 $Y=1.085 $X2=0
+ $Y2=0
cc_691 N_A_1034_392#_c_650_n N_VGND_c_2246_n 0.0538367f $X=7.05 $Y=0.34 $X2=0
+ $Y2=0
cc_692 N_A_1034_392#_c_651_n N_VGND_c_2246_n 0.0138923f $X=5.62 $Y=0.34 $X2=0
+ $Y2=0
cc_693 N_A_1034_392#_c_654_n N_VGND_c_2246_n 0.0122484f $X=7.93 $Y=0.665 $X2=0
+ $Y2=0
cc_694 N_A_1034_392#_c_655_n N_VGND_c_2246_n 0.0415191f $X=9.065 $Y=0.34 $X2=0
+ $Y2=0
cc_695 N_A_1034_392#_c_656_n N_VGND_c_2246_n 0.00655543f $X=8.1 $Y=0.34 $X2=0
+ $Y2=0
cc_696 N_A_1034_392#_c_650_n N_VGND_c_2249_n 0.0118008f $X=7.05 $Y=0.34 $X2=0
+ $Y2=0
cc_697 N_A_1034_392#_c_654_n N_VGND_c_2249_n 0.0246013f $X=7.93 $Y=0.665 $X2=0
+ $Y2=0
cc_698 N_A_1034_392#_c_656_n N_VGND_c_2249_n 0.0135793f $X=8.1 $Y=0.34 $X2=0
+ $Y2=0
cc_699 N_A_1034_392#_c_680_p A_1397_119# 0.00349303f $X=7.22 $Y=0.665 $X2=-0.19
+ $Y2=-0.245
cc_700 N_A_1367_93#_M1019_g N_RESET_B_c_977_n 0.00882199f $X=6.91 $Y=0.805 $X2=0
+ $Y2=0
cc_701 N_A_1367_93#_c_868_n N_RESET_B_c_977_n 2.57602e-19 $X=7.325 $Y=1.005
+ $X2=0 $Y2=0
cc_702 N_A_1367_93#_M1019_g N_RESET_B_M1007_g 0.0398707f $X=6.91 $Y=0.805 $X2=0
+ $Y2=0
cc_703 N_A_1367_93#_c_865_n N_RESET_B_M1007_g 0.00127951f $X=7.185 $Y=1.64 $X2=0
+ $Y2=0
cc_704 N_A_1367_93#_c_867_n N_RESET_B_M1007_g 0.00681742f $X=8.27 $Y=1.005 $X2=0
+ $Y2=0
cc_705 N_A_1367_93#_c_868_n N_RESET_B_M1007_g 0.00424625f $X=7.325 $Y=1.005
+ $X2=0 $Y2=0
cc_706 N_A_1367_93#_c_867_n N_RESET_B_c_980_n 0.0117401f $X=8.27 $Y=1.005 $X2=0
+ $Y2=0
cc_707 N_A_1367_93#_c_865_n N_RESET_B_c_981_n 0.00932005f $X=7.185 $Y=1.64 $X2=0
+ $Y2=0
cc_708 N_A_1367_93#_c_866_n N_RESET_B_c_981_n 0.0083853f $X=7.185 $Y=1.64 $X2=0
+ $Y2=0
cc_709 N_A_1367_93#_M1019_g N_RESET_B_c_982_n 0.0024449f $X=6.91 $Y=0.805 $X2=0
+ $Y2=0
cc_710 N_A_1367_93#_c_871_n N_RESET_B_c_982_n 0.00501376f $X=7.06 $Y=2.14 $X2=0
+ $Y2=0
cc_711 N_A_1367_93#_c_865_n N_RESET_B_c_982_n 0.00103605f $X=7.185 $Y=1.64 $X2=0
+ $Y2=0
cc_712 N_A_1367_93#_c_866_n N_RESET_B_c_982_n 0.0173421f $X=7.185 $Y=1.64 $X2=0
+ $Y2=0
cc_713 N_A_1367_93#_c_872_n N_RESET_B_c_990_n 0.01292f $X=7.06 $Y=2.23 $X2=0
+ $Y2=0
cc_714 N_A_1367_93#_c_871_n N_RESET_B_c_995_n 0.0101236f $X=7.06 $Y=2.14 $X2=0
+ $Y2=0
cc_715 N_A_1367_93#_c_865_n N_RESET_B_c_995_n 0.00823427f $X=7.185 $Y=1.64 $X2=0
+ $Y2=0
cc_716 N_A_1367_93#_c_866_n N_RESET_B_c_995_n 0.00318126f $X=7.185 $Y=1.64 $X2=0
+ $Y2=0
cc_717 N_A_1367_93#_M1013_d N_RESET_B_c_997_n 0.00464147f $X=8.77 $Y=1.735 $X2=0
+ $Y2=0
cc_718 N_A_1367_93#_c_876_n N_RESET_B_c_997_n 0.0360053f $X=8.92 $Y=1.88 $X2=0
+ $Y2=0
cc_719 N_A_1367_93#_c_872_n N_RESET_B_c_1002_n 0.00501376f $X=7.06 $Y=2.23 $X2=0
+ $Y2=0
cc_720 N_A_1367_93#_c_867_n N_A_1234_119#_M1031_g 0.01076f $X=8.27 $Y=1.005
+ $X2=0 $Y2=0
cc_721 N_A_1367_93#_c_869_n N_A_1234_119#_M1031_g 0.0114957f $X=8.435 $Y=0.81
+ $X2=0 $Y2=0
cc_722 N_A_1367_93#_c_870_n N_A_1234_119#_M1031_g 9.26224e-19 $X=8.865 $Y=1.715
+ $X2=0 $Y2=0
cc_723 N_A_1367_93#_c_869_n N_A_1234_119#_c_1207_n 0.00716915f $X=8.435 $Y=0.81
+ $X2=0 $Y2=0
cc_724 N_A_1367_93#_c_870_n N_A_1234_119#_c_1207_n 0.0102608f $X=8.865 $Y=1.715
+ $X2=0 $Y2=0
cc_725 N_A_1367_93#_c_875_n N_A_1234_119#_c_1216_n 0.00282141f $X=8.865 $Y=1.855
+ $X2=0 $Y2=0
cc_726 N_A_1367_93#_c_876_n N_A_1234_119#_c_1216_n 0.0109404f $X=8.92 $Y=1.88
+ $X2=0 $Y2=0
cc_727 N_A_1367_93#_c_870_n N_A_1234_119#_c_1216_n 0.00260822f $X=8.865 $Y=1.715
+ $X2=0 $Y2=0
cc_728 N_A_1367_93#_M1019_g N_A_1234_119#_c_1208_n 0.004969f $X=6.91 $Y=0.805
+ $X2=0 $Y2=0
cc_729 N_A_1367_93#_c_868_n N_A_1234_119#_c_1208_n 0.00929856f $X=7.325 $Y=1.005
+ $X2=0 $Y2=0
cc_730 N_A_1367_93#_M1019_g N_A_1234_119#_c_1209_n 0.00772383f $X=6.91 $Y=0.805
+ $X2=0 $Y2=0
cc_731 N_A_1367_93#_c_871_n N_A_1234_119#_c_1209_n 0.00919528f $X=7.06 $Y=2.14
+ $X2=0 $Y2=0
cc_732 N_A_1367_93#_c_872_n N_A_1234_119#_c_1209_n 9.97148e-19 $X=7.06 $Y=2.23
+ $X2=0 $Y2=0
cc_733 N_A_1367_93#_c_865_n N_A_1234_119#_c_1209_n 0.0517809f $X=7.185 $Y=1.64
+ $X2=0 $Y2=0
cc_734 N_A_1367_93#_c_866_n N_A_1234_119#_c_1209_n 0.00937107f $X=7.185 $Y=1.64
+ $X2=0 $Y2=0
cc_735 N_A_1367_93#_c_868_n N_A_1234_119#_c_1209_n 0.00480628f $X=7.325 $Y=1.005
+ $X2=0 $Y2=0
cc_736 N_A_1367_93#_c_872_n N_A_1234_119#_c_1253_n 0.0116684f $X=7.06 $Y=2.23
+ $X2=0 $Y2=0
cc_737 N_A_1367_93#_c_865_n N_A_1234_119#_c_1253_n 0.0034045f $X=7.185 $Y=1.64
+ $X2=0 $Y2=0
cc_738 N_A_1367_93#_c_866_n N_A_1234_119#_c_1253_n 0.00356794f $X=7.185 $Y=1.64
+ $X2=0 $Y2=0
cc_739 N_A_1367_93#_c_871_n N_A_1234_119#_c_1210_n 0.00330246f $X=7.06 $Y=2.14
+ $X2=0 $Y2=0
cc_740 N_A_1367_93#_c_872_n N_A_1234_119#_c_1210_n 0.00151519f $X=7.06 $Y=2.23
+ $X2=0 $Y2=0
cc_741 N_A_1367_93#_c_865_n N_A_1234_119#_c_1210_n 0.0170101f $X=7.185 $Y=1.64
+ $X2=0 $Y2=0
cc_742 N_A_1367_93#_c_866_n N_A_1234_119#_c_1210_n 0.00147646f $X=7.185 $Y=1.64
+ $X2=0 $Y2=0
cc_743 N_A_1367_93#_c_865_n N_A_1234_119#_c_1211_n 0.0270592f $X=7.185 $Y=1.64
+ $X2=0 $Y2=0
cc_744 N_A_1367_93#_c_866_n N_A_1234_119#_c_1211_n 7.33487e-19 $X=7.185 $Y=1.64
+ $X2=0 $Y2=0
cc_745 N_A_1367_93#_c_867_n N_A_1234_119#_c_1211_n 0.0135416f $X=8.27 $Y=1.005
+ $X2=0 $Y2=0
cc_746 N_A_1367_93#_c_867_n N_A_1234_119#_c_1212_n 0.0457531f $X=8.27 $Y=1.005
+ $X2=0 $Y2=0
cc_747 N_A_1367_93#_c_869_n N_A_1234_119#_c_1212_n 0.00357705f $X=8.435 $Y=0.81
+ $X2=0 $Y2=0
cc_748 N_A_1367_93#_c_870_n N_A_1234_119#_c_1212_n 0.0123924f $X=8.865 $Y=1.715
+ $X2=0 $Y2=0
cc_749 N_A_1367_93#_c_867_n N_A_1234_119#_c_1213_n 0.00365093f $X=8.27 $Y=1.005
+ $X2=0 $Y2=0
cc_750 N_A_1367_93#_c_869_n N_A_1234_119#_c_1213_n 4.74815e-19 $X=8.435 $Y=0.81
+ $X2=0 $Y2=0
cc_751 N_A_1367_93#_c_870_n N_A_1234_119#_c_1213_n 0.00153128f $X=8.865 $Y=1.715
+ $X2=0 $Y2=0
cc_752 N_A_1367_93#_M1019_g N_A_1234_119#_c_1214_n 0.00107029f $X=6.91 $Y=0.805
+ $X2=0 $Y2=0
cc_753 N_A_1367_93#_c_872_n N_A_1234_119#_c_1221_n 0.00554019f $X=7.06 $Y=2.23
+ $X2=0 $Y2=0
cc_754 N_A_1367_93#_c_872_n N_A_835_98#_c_1358_n 0.00284772f $X=7.06 $Y=2.23
+ $X2=0 $Y2=0
cc_755 N_A_1367_93#_c_872_n N_A_835_98#_c_1360_n 0.0278287f $X=7.06 $Y=2.23
+ $X2=0 $Y2=0
cc_756 N_A_1367_93#_c_872_n N_A_835_98#_c_1361_n 0.0095327f $X=7.06 $Y=2.23
+ $X2=0 $Y2=0
cc_757 N_A_1367_93#_c_876_n N_A_835_98#_c_1361_n 0.00408637f $X=8.92 $Y=1.88
+ $X2=0 $Y2=0
cc_758 N_A_1367_93#_c_875_n N_A_835_98#_M1018_g 0.0075382f $X=8.865 $Y=1.855
+ $X2=0 $Y2=0
cc_759 N_A_1367_93#_c_870_n N_A_835_98#_M1018_g 4.14175e-19 $X=8.865 $Y=1.715
+ $X2=0 $Y2=0
cc_760 N_A_1367_93#_c_870_n N_A_835_98#_c_1346_n 0.00134852f $X=8.865 $Y=1.715
+ $X2=0 $Y2=0
cc_761 N_A_1367_93#_c_869_n N_A_1745_74#_M1003_d 0.00295216f $X=8.435 $Y=0.81
+ $X2=-0.19 $Y2=-0.245
cc_762 N_A_1367_93#_c_876_n N_A_1745_74#_c_1677_n 0.0117842f $X=8.92 $Y=1.88
+ $X2=0 $Y2=0
cc_763 N_A_1367_93#_c_872_n N_VPWR_c_1878_n 0.00454716f $X=7.06 $Y=2.23 $X2=0
+ $Y2=0
cc_764 N_A_1367_93#_c_875_n N_VPWR_c_1880_n 0.0728f $X=8.865 $Y=1.855 $X2=0
+ $Y2=0
cc_765 N_A_1367_93#_c_869_n N_VPWR_c_1880_n 0.00559467f $X=8.435 $Y=0.81 $X2=0
+ $Y2=0
cc_766 N_A_1367_93#_c_876_n N_VPWR_c_1886_n 0.00629779f $X=8.92 $Y=1.88 $X2=0
+ $Y2=0
cc_767 N_A_1367_93#_c_872_n N_VPWR_c_1874_n 9.43083e-19 $X=7.06 $Y=2.23 $X2=0
+ $Y2=0
cc_768 N_A_1367_93#_c_876_n N_VPWR_c_1874_n 0.00766223f $X=8.92 $Y=1.88 $X2=0
+ $Y2=0
cc_769 N_A_1367_93#_M1019_g N_A_300_464#_c_2047_n 3.24142e-19 $X=6.91 $Y=0.805
+ $X2=0 $Y2=0
cc_770 N_A_1367_93#_c_866_n N_A_300_464#_c_2047_n 2.29181e-19 $X=7.185 $Y=1.64
+ $X2=0 $Y2=0
cc_771 N_A_1367_93#_c_867_n N_VGND_M1007_d 0.00911951f $X=8.27 $Y=1.005 $X2=0
+ $Y2=0
cc_772 N_A_1367_93#_c_868_n A_1397_119# 0.00204263f $X=7.325 $Y=1.005 $X2=-0.19
+ $Y2=-0.245
cc_773 N_RESET_B_c_980_n N_A_1234_119#_M1031_g 0.0052575f $X=7.595 $Y=1.19 $X2=0
+ $Y2=0
cc_774 N_RESET_B_c_997_n N_A_1234_119#_c_1207_n 3.01246e-19 $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_775 N_RESET_B_c_997_n N_A_1234_119#_c_1216_n 0.0082395f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_776 N_RESET_B_c_995_n N_A_1234_119#_c_1217_n 0.00861368f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_777 N_RESET_B_M1007_g N_A_1234_119#_c_1208_n 3.96747e-19 $X=7.3 $Y=0.805
+ $X2=0 $Y2=0
cc_778 N_RESET_B_c_995_n N_A_1234_119#_c_1209_n 0.0240634f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_779 N_RESET_B_c_995_n N_A_1234_119#_c_1253_n 0.0215639f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_780 N_RESET_B_c_982_n N_A_1234_119#_c_1210_n 0.0113497f $X=7.67 $Y=1.815
+ $X2=0 $Y2=0
cc_781 N_RESET_B_c_990_n N_A_1234_119#_c_1210_n 0.0182508f $X=7.685 $Y=2.23
+ $X2=0 $Y2=0
cc_782 N_RESET_B_c_995_n N_A_1234_119#_c_1210_n 0.0273088f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_783 N_RESET_B_c_998_n N_A_1234_119#_c_1210_n 0.01197f $X=8.065 $Y=2.035 $X2=0
+ $Y2=0
cc_784 N_RESET_B_c_999_n N_A_1234_119#_c_1210_n 0.0389238f $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_785 N_RESET_B_c_1002_n N_A_1234_119#_c_1210_n 0.0165391f $X=7.685 $Y=2.022
+ $X2=0 $Y2=0
cc_786 N_RESET_B_c_980_n N_A_1234_119#_c_1211_n 0.00404376f $X=7.595 $Y=1.19
+ $X2=0 $Y2=0
cc_787 N_RESET_B_c_982_n N_A_1234_119#_c_1211_n 0.00501753f $X=7.67 $Y=1.815
+ $X2=0 $Y2=0
cc_788 N_RESET_B_c_980_n N_A_1234_119#_c_1212_n 7.39613e-19 $X=7.595 $Y=1.19
+ $X2=0 $Y2=0
cc_789 N_RESET_B_c_982_n N_A_1234_119#_c_1212_n 0.00710493f $X=7.67 $Y=1.815
+ $X2=0 $Y2=0
cc_790 N_RESET_B_c_995_n N_A_1234_119#_c_1212_n 0.00357593f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_791 N_RESET_B_c_997_n N_A_1234_119#_c_1212_n 0.00581394f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_792 N_RESET_B_c_998_n N_A_1234_119#_c_1212_n 0.00371961f $X=8.065 $Y=2.035
+ $X2=0 $Y2=0
cc_793 N_RESET_B_c_999_n N_A_1234_119#_c_1212_n 0.0172409f $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_794 N_RESET_B_c_1002_n N_A_1234_119#_c_1212_n 0.00735754f $X=7.685 $Y=2.022
+ $X2=0 $Y2=0
cc_795 N_RESET_B_c_980_n N_A_1234_119#_c_1213_n 0.0182615f $X=7.595 $Y=1.19
+ $X2=0 $Y2=0
cc_796 N_RESET_B_c_982_n N_A_1234_119#_c_1213_n 6.54113e-19 $X=7.67 $Y=1.815
+ $X2=0 $Y2=0
cc_797 N_RESET_B_c_997_n N_A_1234_119#_c_1213_n 0.00593186f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_798 N_RESET_B_c_999_n N_A_1234_119#_c_1213_n 6.74459e-19 $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_799 N_RESET_B_c_1002_n N_A_1234_119#_c_1213_n 0.0093828f $X=7.685 $Y=2.022
+ $X2=0 $Y2=0
cc_800 N_RESET_B_c_995_n N_A_835_98#_M1027_s 0.0011277f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_801 N_RESET_B_c_995_n N_A_835_98#_c_1354_n 0.00350083f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_802 N_RESET_B_c_977_n N_A_835_98#_c_1342_n 0.0103973f $X=7.225 $Y=0.18 $X2=0
+ $Y2=0
cc_803 N_RESET_B_c_995_n N_A_835_98#_c_1355_n 0.00218847f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_804 N_RESET_B_c_977_n N_A_835_98#_c_1344_n 0.00882199f $X=7.225 $Y=0.18 $X2=0
+ $Y2=0
cc_805 N_RESET_B_c_995_n N_A_835_98#_c_1360_n 0.0038794f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_806 N_RESET_B_c_990_n N_A_835_98#_c_1361_n 0.00949691f $X=7.685 $Y=2.23 $X2=0
+ $Y2=0
cc_807 N_RESET_B_c_997_n N_A_835_98#_M1018_g 0.0137675f $X=10.655 $Y=2.035 $X2=0
+ $Y2=0
cc_808 N_RESET_B_c_997_n N_A_835_98#_c_1345_n 0.00383889f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_809 N_RESET_B_c_997_n N_A_835_98#_c_1346_n 2.83807e-19 $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_810 N_RESET_B_c_977_n N_A_835_98#_c_1374_n 0.00129274f $X=7.225 $Y=0.18 $X2=0
+ $Y2=0
cc_811 N_RESET_B_c_977_n N_A_835_98#_c_1351_n 0.00782328f $X=7.225 $Y=0.18 $X2=0
+ $Y2=0
cc_812 N_RESET_B_c_987_n N_A_835_98#_c_1352_n 0.00113917f $X=3.93 $Y=1.995 $X2=0
+ $Y2=0
cc_813 N_RESET_B_c_988_n N_A_835_98#_c_1352_n 0.0013004f $X=3.695 $Y=1.995 $X2=0
+ $Y2=0
cc_814 N_RESET_B_c_995_n N_A_835_98#_c_1352_n 0.0467967f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_815 N_RESET_B_c_996_n N_A_835_98#_c_1352_n 0.0028417f $X=4.225 $Y=2.035 $X2=0
+ $Y2=0
cc_816 N_RESET_B_c_1001_n N_A_835_98#_c_1352_n 0.0281446f $X=3.95 $Y=1.995 $X2=0
+ $Y2=0
cc_817 N_RESET_B_c_995_n N_A_835_98#_c_1353_n 0.0016494f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_818 N_RESET_B_M1036_g N_A_1997_272#_M1001_g 0.0312551f $X=10.6 $Y=0.58 $X2=0
+ $Y2=0
cc_819 N_RESET_B_c_984_n N_A_1997_272#_c_1544_n 0.0225363f $X=10.715 $Y=1.82
+ $X2=0 $Y2=0
cc_820 N_RESET_B_c_985_n N_A_1997_272#_c_1544_n 0.00643996f $X=10.715 $Y=1.375
+ $X2=0 $Y2=0
cc_821 N_RESET_B_c_1003_n N_A_1997_272#_c_1544_n 0.00119422f $X=10.805 $Y=1.985
+ $X2=0 $Y2=0
cc_822 N_RESET_B_c_992_n N_A_1997_272#_c_1555_n 0.00511887f $X=10.885 $Y=2.375
+ $X2=0 $Y2=0
cc_823 N_RESET_B_c_997_n N_A_1997_272#_c_1555_n 0.00508273f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_824 N_RESET_B_c_1004_n N_A_1997_272#_c_1555_n 0.0128577f $X=10.885 $Y=1.985
+ $X2=0 $Y2=0
cc_825 N_RESET_B_c_993_n N_A_1997_272#_c_1556_n 0.0138023f $X=10.885 $Y=2.465
+ $X2=0 $Y2=0
cc_826 N_RESET_B_c_984_n N_A_1997_272#_c_1545_n 0.00935059f $X=10.715 $Y=1.82
+ $X2=0 $Y2=0
cc_827 N_RESET_B_c_985_n N_A_1997_272#_c_1545_n 0.0053082f $X=10.715 $Y=1.375
+ $X2=0 $Y2=0
cc_828 RESET_B N_A_1997_272#_c_1545_n 0.00164136f $X=10.715 $Y=1.95 $X2=0 $Y2=0
cc_829 N_RESET_B_c_1003_n N_A_1997_272#_c_1545_n 0.0191591f $X=10.805 $Y=1.985
+ $X2=0 $Y2=0
cc_830 N_RESET_B_c_1004_n N_A_1997_272#_c_1545_n 0.00143438f $X=10.885 $Y=1.985
+ $X2=0 $Y2=0
cc_831 N_RESET_B_M1036_g N_A_1997_272#_c_1546_n 0.00111706f $X=10.6 $Y=0.58
+ $X2=0 $Y2=0
cc_832 N_RESET_B_M1036_g N_A_1997_272#_c_1549_n 7.22053e-19 $X=10.6 $Y=0.58
+ $X2=0 $Y2=0
cc_833 N_RESET_B_c_997_n N_A_1997_272#_c_1551_n 0.0131744f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_834 N_RESET_B_c_993_n N_A_1997_272#_c_1557_n 0.00680136f $X=10.885 $Y=2.465
+ $X2=0 $Y2=0
cc_835 N_RESET_B_c_1003_n N_A_1997_272#_c_1557_n 9.92047e-19 $X=10.805 $Y=1.985
+ $X2=0 $Y2=0
cc_836 N_RESET_B_c_984_n N_A_1997_272#_c_1552_n 0.00366777f $X=10.715 $Y=1.82
+ $X2=0 $Y2=0
cc_837 N_RESET_B_c_993_n N_A_1997_272#_c_1552_n 0.00111437f $X=10.885 $Y=2.465
+ $X2=0 $Y2=0
cc_838 RESET_B N_A_1997_272#_c_1552_n 0.00158814f $X=10.715 $Y=1.95 $X2=0 $Y2=0
cc_839 N_RESET_B_c_1003_n N_A_1997_272#_c_1552_n 0.0232461f $X=10.805 $Y=1.985
+ $X2=0 $Y2=0
cc_840 N_RESET_B_c_1004_n N_A_1997_272#_c_1552_n 0.00858202f $X=10.885 $Y=1.985
+ $X2=0 $Y2=0
cc_841 N_RESET_B_c_997_n N_A_1745_74#_M1018_d 0.00297016f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_842 N_RESET_B_M1036_g N_A_1745_74#_M1021_g 0.0518692f $X=10.6 $Y=0.58 $X2=0
+ $Y2=0
cc_843 N_RESET_B_c_985_n N_A_1745_74#_c_1661_n 0.0117915f $X=10.715 $Y=1.375
+ $X2=0 $Y2=0
cc_844 N_RESET_B_c_1003_n N_A_1745_74#_c_1661_n 3.43698e-19 $X=10.805 $Y=1.985
+ $X2=0 $Y2=0
cc_845 N_RESET_B_c_1004_n N_A_1745_74#_c_1661_n 0.00946465f $X=10.885 $Y=1.985
+ $X2=0 $Y2=0
cc_846 N_RESET_B_c_993_n N_A_1745_74#_c_1672_n 0.00946465f $X=10.885 $Y=2.465
+ $X2=0 $Y2=0
cc_847 N_RESET_B_c_993_n N_A_1745_74#_c_1673_n 0.00921795f $X=10.885 $Y=2.465
+ $X2=0 $Y2=0
cc_848 N_RESET_B_M1036_g N_A_1745_74#_c_1663_n 0.00646231f $X=10.6 $Y=0.58 $X2=0
+ $Y2=0
cc_849 N_RESET_B_c_985_n N_A_1745_74#_c_1663_n 0.0030434f $X=10.715 $Y=1.375
+ $X2=0 $Y2=0
cc_850 N_RESET_B_c_992_n N_A_1745_74#_c_1676_n 0.00946465f $X=10.885 $Y=2.375
+ $X2=0 $Y2=0
cc_851 N_RESET_B_c_997_n N_A_1745_74#_c_1677_n 0.00561127f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_852 N_RESET_B_c_984_n N_A_1745_74#_c_1679_n 6.20198e-19 $X=10.715 $Y=1.82
+ $X2=0 $Y2=0
cc_853 N_RESET_B_c_997_n N_A_1745_74#_c_1679_n 0.0131083f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_854 RESET_B N_A_1745_74#_c_1679_n 2.51275e-19 $X=10.715 $Y=1.95 $X2=0 $Y2=0
cc_855 N_RESET_B_c_1003_n N_A_1745_74#_c_1679_n 0.00608543f $X=10.805 $Y=1.985
+ $X2=0 $Y2=0
cc_856 N_RESET_B_c_997_n N_A_1745_74#_c_1680_n 0.0053742f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_857 N_RESET_B_c_992_n N_A_1745_74#_c_1681_n 0.00159843f $X=10.885 $Y=2.375
+ $X2=0 $Y2=0
cc_858 N_RESET_B_c_993_n N_A_1745_74#_c_1681_n 2.78257e-19 $X=10.885 $Y=2.465
+ $X2=0 $Y2=0
cc_859 N_RESET_B_c_997_n N_A_1745_74#_c_1681_n 0.020931f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_860 RESET_B N_A_1745_74#_c_1681_n 3.29892e-19 $X=10.715 $Y=1.95 $X2=0 $Y2=0
cc_861 N_RESET_B_c_1003_n N_A_1745_74#_c_1681_n 0.00622512f $X=10.805 $Y=1.985
+ $X2=0 $Y2=0
cc_862 N_RESET_B_c_1004_n N_A_1745_74#_c_1681_n 6.08738e-19 $X=10.885 $Y=1.985
+ $X2=0 $Y2=0
cc_863 N_RESET_B_M1036_g N_A_1745_74#_c_1670_n 0.015752f $X=10.6 $Y=0.58 $X2=0
+ $Y2=0
cc_864 N_RESET_B_c_985_n N_A_1745_74#_c_1670_n 0.00357206f $X=10.715 $Y=1.375
+ $X2=0 $Y2=0
cc_865 N_RESET_B_c_995_n N_VPWR_M1027_d 6.6495e-19 $X=7.775 $Y=2.035 $X2=0 $Y2=0
cc_866 N_RESET_B_c_997_n N_VPWR_M1013_s 0.00689173f $X=10.655 $Y=2.035 $X2=0
+ $Y2=0
cc_867 N_RESET_B_c_994_n N_VPWR_c_1876_n 0.00571347f $X=3.56 $Y=2.245 $X2=0
+ $Y2=0
cc_868 N_RESET_B_c_990_n N_VPWR_c_1878_n 0.00404752f $X=7.685 $Y=2.23 $X2=0
+ $Y2=0
cc_869 N_RESET_B_c_995_n N_VPWR_c_1878_n 7.58628e-19 $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_870 N_RESET_B_c_982_n N_VPWR_c_1880_n 0.00146391f $X=7.67 $Y=1.815 $X2=0
+ $Y2=0
cc_871 N_RESET_B_c_990_n N_VPWR_c_1880_n 0.00504716f $X=7.685 $Y=2.23 $X2=0
+ $Y2=0
cc_872 N_RESET_B_c_997_n N_VPWR_c_1880_n 0.0185404f $X=10.655 $Y=2.035 $X2=0
+ $Y2=0
cc_873 N_RESET_B_c_998_n N_VPWR_c_1880_n 5.19261e-19 $X=8.065 $Y=2.035 $X2=0
+ $Y2=0
cc_874 N_RESET_B_c_999_n N_VPWR_c_1880_n 0.0183634f $X=7.92 $Y=2.035 $X2=0 $Y2=0
cc_875 N_RESET_B_c_1002_n N_VPWR_c_1880_n 0.00295171f $X=7.685 $Y=2.022 $X2=0
+ $Y2=0
cc_876 N_RESET_B_c_993_n N_VPWR_c_1881_n 0.00720194f $X=10.885 $Y=2.465 $X2=0
+ $Y2=0
cc_877 N_RESET_B_c_997_n N_VPWR_c_1881_n 0.00652534f $X=10.655 $Y=2.035 $X2=0
+ $Y2=0
cc_878 RESET_B N_VPWR_c_1881_n 6.45709e-19 $X=10.715 $Y=1.95 $X2=0 $Y2=0
cc_879 N_RESET_B_c_1003_n N_VPWR_c_1881_n 0.00292772f $X=10.805 $Y=1.985 $X2=0
+ $Y2=0
cc_880 N_RESET_B_c_1004_n N_VPWR_c_1881_n 6.5955e-19 $X=10.885 $Y=1.985 $X2=0
+ $Y2=0
cc_881 N_RESET_B_c_994_n N_VPWR_c_1884_n 0.00445602f $X=3.56 $Y=2.245 $X2=0
+ $Y2=0
cc_882 N_RESET_B_c_993_n N_VPWR_c_1888_n 0.00445602f $X=10.885 $Y=2.465 $X2=0
+ $Y2=0
cc_883 N_RESET_B_c_990_n N_VPWR_c_1874_n 9.43083e-19 $X=7.685 $Y=2.23 $X2=0
+ $Y2=0
cc_884 N_RESET_B_c_993_n N_VPWR_c_1874_n 0.00896147f $X=10.885 $Y=2.465 $X2=0
+ $Y2=0
cc_885 N_RESET_B_c_994_n N_VPWR_c_1874_n 0.00453497f $X=3.56 $Y=2.245 $X2=0
+ $Y2=0
cc_886 N_RESET_B_c_988_n N_A_300_464#_c_2072_n 8.77027e-19 $X=3.695 $Y=1.995
+ $X2=0 $Y2=0
cc_887 N_RESET_B_M1037_g N_A_300_464#_c_2041_n 0.0137342f $X=3.5 $Y=0.615 $X2=0
+ $Y2=0
cc_888 N_RESET_B_M1037_g N_A_300_464#_c_2042_n 0.0186001f $X=3.5 $Y=0.615 $X2=0
+ $Y2=0
cc_889 N_RESET_B_c_988_n N_A_300_464#_c_2042_n 0.0187601f $X=3.695 $Y=1.995
+ $X2=0 $Y2=0
cc_890 N_RESET_B_c_994_n N_A_300_464#_c_2042_n 0.00445911f $X=3.56 $Y=2.245
+ $X2=0 $Y2=0
cc_891 N_RESET_B_c_996_n N_A_300_464#_c_2042_n 0.00108729f $X=4.225 $Y=2.035
+ $X2=0 $Y2=0
cc_892 N_RESET_B_c_1001_n N_A_300_464#_c_2042_n 0.0243953f $X=3.95 $Y=1.995
+ $X2=0 $Y2=0
cc_893 N_RESET_B_c_995_n N_A_300_464#_c_2051_n 0.00515092f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_894 N_RESET_B_c_987_n N_A_300_464#_c_2052_n 0.00525707f $X=3.93 $Y=1.995
+ $X2=0 $Y2=0
cc_895 N_RESET_B_c_994_n N_A_300_464#_c_2052_n 0.0137348f $X=3.56 $Y=2.245 $X2=0
+ $Y2=0
cc_896 N_RESET_B_c_995_n N_A_300_464#_c_2052_n 0.00101627f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_897 N_RESET_B_c_996_n N_A_300_464#_c_2052_n 0.00440623f $X=4.225 $Y=2.035
+ $X2=0 $Y2=0
cc_898 N_RESET_B_c_1001_n N_A_300_464#_c_2052_n 0.0258218f $X=3.95 $Y=1.995
+ $X2=0 $Y2=0
cc_899 N_RESET_B_c_995_n N_A_300_464#_c_2053_n 0.0138526f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_900 N_RESET_B_c_995_n N_A_300_464#_c_2045_n 0.00360371f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_901 N_RESET_B_c_995_n N_A_300_464#_c_2055_n 0.0179072f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_902 N_RESET_B_c_995_n N_A_300_464#_c_2056_n 0.0167674f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_903 N_RESET_B_c_995_n N_A_300_464#_c_2047_n 0.0094217f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_904 N_RESET_B_c_994_n N_A_300_464#_c_2059_n 0.00511769f $X=3.56 $Y=2.245
+ $X2=0 $Y2=0
cc_905 N_RESET_B_M1037_g N_VGND_c_2232_n 0.00141396f $X=3.5 $Y=0.615 $X2=0 $Y2=0
cc_906 N_RESET_B_c_977_n N_VGND_c_2232_n 0.0208132f $X=7.225 $Y=0.18 $X2=0 $Y2=0
cc_907 N_RESET_B_c_977_n N_VGND_c_2233_n 0.02563f $X=7.225 $Y=0.18 $X2=0 $Y2=0
cc_908 N_RESET_B_M1036_g N_VGND_c_2234_n 0.00390833f $X=10.6 $Y=0.58 $X2=0 $Y2=0
cc_909 N_RESET_B_c_977_n N_VGND_c_2237_n 0.0242452f $X=7.225 $Y=0.18 $X2=0 $Y2=0
cc_910 N_RESET_B_c_978_n N_VGND_c_2240_n 0.0064002f $X=3.575 $Y=0.18 $X2=0 $Y2=0
cc_911 N_RESET_B_c_977_n N_VGND_c_2241_n 0.0512939f $X=7.225 $Y=0.18 $X2=0 $Y2=0
cc_912 N_RESET_B_M1036_g N_VGND_c_2243_n 0.00460063f $X=10.6 $Y=0.58 $X2=0 $Y2=0
cc_913 N_RESET_B_c_977_n N_VGND_c_2246_n 0.0903551f $X=7.225 $Y=0.18 $X2=0 $Y2=0
cc_914 N_RESET_B_c_978_n N_VGND_c_2246_n 0.0113744f $X=3.575 $Y=0.18 $X2=0 $Y2=0
cc_915 N_RESET_B_M1036_g N_VGND_c_2246_n 0.00906826f $X=10.6 $Y=0.58 $X2=0 $Y2=0
cc_916 N_RESET_B_c_977_n N_VGND_c_2249_n 0.00939536f $X=7.225 $Y=0.18 $X2=0
+ $Y2=0
cc_917 N_RESET_B_M1037_g N_noxref_24_c_2366_n 0.00190559f $X=3.5 $Y=0.615 $X2=0
+ $Y2=0
cc_918 N_A_1234_119#_c_1217_n N_A_835_98#_c_1356_n 0.00396944f $X=6.71 $Y=2.555
+ $X2=0 $Y2=0
cc_919 N_A_1234_119#_c_1214_n N_A_835_98#_c_1344_n 0.00566398f $X=6.31 $Y=0.81
+ $X2=0 $Y2=0
cc_920 N_A_1234_119#_c_1217_n N_A_835_98#_c_1360_n 0.00979816f $X=6.71 $Y=2.555
+ $X2=0 $Y2=0
cc_921 N_A_1234_119#_c_1209_n N_A_835_98#_c_1360_n 0.00327177f $X=6.795 $Y=2.32
+ $X2=0 $Y2=0
cc_922 N_A_1234_119#_c_1221_n N_A_835_98#_c_1360_n 0.00504398f $X=6.795 $Y=2.522
+ $X2=0 $Y2=0
cc_923 N_A_1234_119#_c_1216_n N_A_835_98#_c_1361_n 0.0102036f $X=8.695 $Y=1.66
+ $X2=0 $Y2=0
cc_924 N_A_1234_119#_c_1253_n N_A_835_98#_c_1361_n 0.003989f $X=7.495 $Y=2.405
+ $X2=0 $Y2=0
cc_925 N_A_1234_119#_c_1210_n N_A_835_98#_c_1361_n 0.00777265f $X=7.58 $Y=2.32
+ $X2=0 $Y2=0
cc_926 N_A_1234_119#_c_1221_n N_A_835_98#_c_1361_n 0.00119096f $X=6.795 $Y=2.522
+ $X2=0 $Y2=0
cc_927 N_A_1234_119#_c_1216_n N_A_835_98#_c_1362_n 0.00230914f $X=8.695 $Y=1.66
+ $X2=0 $Y2=0
cc_928 N_A_1234_119#_c_1216_n N_A_835_98#_M1018_g 0.00557664f $X=8.695 $Y=1.66
+ $X2=0 $Y2=0
cc_929 N_A_1234_119#_c_1207_n N_A_835_98#_c_1346_n 0.00717177f $X=8.605 $Y=1.52
+ $X2=0 $Y2=0
cc_930 N_A_1234_119#_c_1253_n N_VPWR_M1008_d 0.00772988f $X=7.495 $Y=2.405 $X2=0
+ $Y2=0
cc_931 N_A_1234_119#_c_1210_n N_VPWR_M1008_d 7.78169e-19 $X=7.58 $Y=2.32 $X2=0
+ $Y2=0
cc_932 N_A_1234_119#_c_1253_n N_VPWR_c_1878_n 0.0222224f $X=7.495 $Y=2.405 $X2=0
+ $Y2=0
cc_933 N_A_1234_119#_c_1210_n N_VPWR_c_1878_n 0.00949227f $X=7.58 $Y=2.32 $X2=0
+ $Y2=0
cc_934 N_A_1234_119#_c_1221_n N_VPWR_c_1878_n 0.00341149f $X=6.795 $Y=2.522
+ $X2=0 $Y2=0
cc_935 N_A_1234_119#_c_1210_n N_VPWR_c_1879_n 0.00714098f $X=7.58 $Y=2.32 $X2=0
+ $Y2=0
cc_936 N_A_1234_119#_c_1207_n N_VPWR_c_1880_n 0.00460268f $X=8.605 $Y=1.52 $X2=0
+ $Y2=0
cc_937 N_A_1234_119#_c_1216_n N_VPWR_c_1880_n 0.00728995f $X=8.695 $Y=1.66 $X2=0
+ $Y2=0
cc_938 N_A_1234_119#_c_1210_n N_VPWR_c_1880_n 0.0222061f $X=7.58 $Y=2.32 $X2=0
+ $Y2=0
cc_939 N_A_1234_119#_c_1217_n N_VPWR_c_1892_n 0.00833207f $X=6.71 $Y=2.555 $X2=0
+ $Y2=0
cc_940 N_A_1234_119#_c_1221_n N_VPWR_c_1892_n 0.00291643f $X=6.795 $Y=2.522
+ $X2=0 $Y2=0
cc_941 N_A_1234_119#_c_1216_n N_VPWR_c_1874_n 9.39239e-19 $X=8.695 $Y=1.66 $X2=0
+ $Y2=0
cc_942 N_A_1234_119#_c_1217_n N_VPWR_c_1874_n 0.0118132f $X=6.71 $Y=2.555 $X2=0
+ $Y2=0
cc_943 N_A_1234_119#_c_1253_n N_VPWR_c_1874_n 0.0104334f $X=7.495 $Y=2.405 $X2=0
+ $Y2=0
cc_944 N_A_1234_119#_c_1210_n N_VPWR_c_1874_n 0.0154819f $X=7.58 $Y=2.32 $X2=0
+ $Y2=0
cc_945 N_A_1234_119#_c_1221_n N_VPWR_c_1874_n 0.00457064f $X=6.795 $Y=2.522
+ $X2=0 $Y2=0
cc_946 N_A_1234_119#_c_1214_n N_A_300_464#_c_2044_n 0.0168132f $X=6.31 $Y=0.81
+ $X2=0 $Y2=0
cc_947 N_A_1234_119#_c_1217_n N_A_300_464#_c_2054_n 0.0139482f $X=6.71 $Y=2.555
+ $X2=0 $Y2=0
cc_948 N_A_1234_119#_c_1209_n N_A_300_464#_c_2054_n 0.00242728f $X=6.795 $Y=2.32
+ $X2=0 $Y2=0
cc_949 N_A_1234_119#_c_1221_n N_A_300_464#_c_2054_n 0.00168203f $X=6.795
+ $Y=2.522 $X2=0 $Y2=0
cc_950 N_A_1234_119#_c_1208_n N_A_300_464#_c_2045_n 0.00533227f $X=6.71 $Y=0.945
+ $X2=0 $Y2=0
cc_951 N_A_1234_119#_c_1209_n N_A_300_464#_c_2045_n 0.0135847f $X=6.795 $Y=2.32
+ $X2=0 $Y2=0
cc_952 N_A_1234_119#_c_1214_n N_A_300_464#_c_2045_n 0.0268176f $X=6.31 $Y=0.81
+ $X2=0 $Y2=0
cc_953 N_A_1234_119#_c_1217_n N_A_300_464#_c_2055_n 0.0207396f $X=6.71 $Y=2.555
+ $X2=0 $Y2=0
cc_954 N_A_1234_119#_c_1209_n N_A_300_464#_c_2055_n 0.0135339f $X=6.795 $Y=2.32
+ $X2=0 $Y2=0
cc_955 N_A_1234_119#_c_1209_n N_A_300_464#_c_2047_n 0.0490008f $X=6.795 $Y=2.32
+ $X2=0 $Y2=0
cc_956 N_A_1234_119#_c_1253_n A_1343_461# 6.70978e-19 $X=7.495 $Y=2.405
+ $X2=-0.19 $Y2=-0.245
cc_957 N_A_1234_119#_c_1221_n A_1343_461# 0.00461414f $X=6.795 $Y=2.522
+ $X2=-0.19 $Y2=-0.245
cc_958 N_A_1234_119#_M1031_g N_VGND_c_2242_n 0.00278271f $X=8.22 $Y=0.69 $X2=0
+ $Y2=0
cc_959 N_A_1234_119#_M1031_g N_VGND_c_2246_n 0.00358525f $X=8.22 $Y=0.69 $X2=0
+ $Y2=0
cc_960 N_A_1234_119#_M1031_g N_VGND_c_2249_n 0.00111149f $X=8.22 $Y=0.69 $X2=0
+ $Y2=0
cc_961 N_A_1234_119#_c_1208_n A_1320_119# 0.00177672f $X=6.71 $Y=0.945 $X2=-0.19
+ $Y2=-0.245
cc_962 N_A_835_98#_c_1347_n N_A_1997_272#_M1001_g 0.0100846f $X=9.7 $Y=1.51
+ $X2=0 $Y2=0
cc_963 N_A_835_98#_M1002_g N_A_1997_272#_M1001_g 0.0520068f $X=9.785 $Y=0.58
+ $X2=0 $Y2=0
cc_964 N_A_835_98#_c_1347_n N_A_1997_272#_c_1544_n 0.019486f $X=9.7 $Y=1.51
+ $X2=0 $Y2=0
cc_965 N_A_835_98#_c_1347_n N_A_1997_272#_c_1551_n 6.49074e-19 $X=9.7 $Y=1.51
+ $X2=0 $Y2=0
cc_966 N_A_835_98#_c_1362_n N_A_1745_74#_c_1677_n 0.00244716f $X=9.145 $Y=2.9
+ $X2=0 $Y2=0
cc_967 N_A_835_98#_M1018_g N_A_1745_74#_c_1677_n 0.00467021f $X=9.145 $Y=2.235
+ $X2=0 $Y2=0
cc_968 N_A_835_98#_M1002_g N_A_1745_74#_c_1665_n 0.00653104f $X=9.785 $Y=0.58
+ $X2=0 $Y2=0
cc_969 N_A_835_98#_c_1349_n N_A_1745_74#_c_1665_n 0.00549286f $X=9.785 $Y=1.045
+ $X2=0 $Y2=0
cc_970 N_A_835_98#_c_1345_n N_A_1745_74#_c_1666_n 0.0090777f $X=9.625 $Y=1.585
+ $X2=0 $Y2=0
cc_971 N_A_835_98#_c_1347_n N_A_1745_74#_c_1666_n 0.00911046f $X=9.7 $Y=1.51
+ $X2=0 $Y2=0
cc_972 N_A_835_98#_c_1345_n N_A_1745_74#_c_1679_n 2.60059e-19 $X=9.625 $Y=1.585
+ $X2=0 $Y2=0
cc_973 N_A_835_98#_c_1349_n N_A_1745_74#_c_1679_n 3.58986e-19 $X=9.785 $Y=1.045
+ $X2=0 $Y2=0
cc_974 N_A_835_98#_M1002_g N_A_1745_74#_c_1667_n 0.00822927f $X=9.785 $Y=0.58
+ $X2=0 $Y2=0
cc_975 N_A_835_98#_c_1347_n N_A_1745_74#_c_1668_n 0.00212136f $X=9.7 $Y=1.51
+ $X2=0 $Y2=0
cc_976 N_A_835_98#_c_1349_n N_A_1745_74#_c_1668_n 3.68292e-19 $X=9.785 $Y=1.045
+ $X2=0 $Y2=0
cc_977 N_A_835_98#_c_1347_n N_A_1745_74#_c_1670_n 0.00241471f $X=9.7 $Y=1.51
+ $X2=0 $Y2=0
cc_978 N_A_835_98#_c_1349_n N_A_1745_74#_c_1670_n 0.00651625f $X=9.785 $Y=1.045
+ $X2=0 $Y2=0
cc_979 N_A_835_98#_c_1352_n N_VPWR_M1027_d 0.00264501f $X=4.927 $Y=1.852 $X2=0
+ $Y2=0
cc_980 N_A_835_98#_c_1354_n N_VPWR_c_1877_n 0.00850453f $X=5.095 $Y=1.875 $X2=0
+ $Y2=0
cc_981 N_A_835_98#_c_1355_n N_VPWR_c_1877_n 0.00158412f $X=5.615 $Y=3.075 $X2=0
+ $Y2=0
cc_982 N_A_835_98#_c_1357_n N_VPWR_c_1877_n 0.00232909f $X=5.69 $Y=3.15 $X2=0
+ $Y2=0
cc_983 N_A_835_98#_c_1358_n N_VPWR_c_1878_n 0.00612345f $X=6.64 $Y=2.89 $X2=0
+ $Y2=0
cc_984 N_A_835_98#_c_1361_n N_VPWR_c_1878_n 0.025635f $X=9.055 $Y=3.15 $X2=0
+ $Y2=0
cc_985 N_A_835_98#_c_1361_n N_VPWR_c_1879_n 0.0260958f $X=9.055 $Y=3.15 $X2=0
+ $Y2=0
cc_986 N_A_835_98#_c_1361_n N_VPWR_c_1880_n 0.0170937f $X=9.055 $Y=3.15 $X2=0
+ $Y2=0
cc_987 N_A_835_98#_c_1362_n N_VPWR_c_1880_n 0.00527525f $X=9.145 $Y=2.9 $X2=0
+ $Y2=0
cc_988 N_A_835_98#_c_1361_n N_VPWR_c_1886_n 0.0217861f $X=9.055 $Y=3.15 $X2=0
+ $Y2=0
cc_989 N_A_835_98#_c_1354_n N_VPWR_c_1892_n 0.00303678f $X=5.095 $Y=1.875 $X2=0
+ $Y2=0
cc_990 N_A_835_98#_c_1357_n N_VPWR_c_1892_n 0.0484762f $X=5.69 $Y=3.15 $X2=0
+ $Y2=0
cc_991 N_A_835_98#_c_1354_n N_VPWR_c_1874_n 0.00394737f $X=5.095 $Y=1.875 $X2=0
+ $Y2=0
cc_992 N_A_835_98#_c_1356_n N_VPWR_c_1874_n 0.025222f $X=6.55 $Y=3.15 $X2=0
+ $Y2=0
cc_993 N_A_835_98#_c_1357_n N_VPWR_c_1874_n 0.00688721f $X=5.69 $Y=3.15 $X2=0
+ $Y2=0
cc_994 N_A_835_98#_c_1361_n N_VPWR_c_1874_n 0.0749028f $X=9.055 $Y=3.15 $X2=0
+ $Y2=0
cc_995 N_A_835_98#_c_1367_n N_VPWR_c_1874_n 0.00503906f $X=6.64 $Y=3.15 $X2=0
+ $Y2=0
cc_996 N_A_835_98#_M1027_s N_A_300_464#_c_2051_n 0.00851724f $X=4.275 $Y=1.96
+ $X2=0 $Y2=0
cc_997 N_A_835_98#_c_1352_n N_A_300_464#_c_2051_n 0.017483f $X=4.927 $Y=1.852
+ $X2=0 $Y2=0
cc_998 N_A_835_98#_c_1354_n N_A_300_464#_c_2053_n 0.0151931f $X=5.095 $Y=1.875
+ $X2=0 $Y2=0
cc_999 N_A_835_98#_c_1355_n N_A_300_464#_c_2053_n 0.0148953f $X=5.615 $Y=3.075
+ $X2=0 $Y2=0
cc_1000 N_A_835_98#_c_1356_n N_A_300_464#_c_2053_n 7.24606e-19 $X=6.55 $Y=3.15
+ $X2=0 $Y2=0
cc_1001 N_A_835_98#_c_1352_n N_A_300_464#_c_2053_n 0.0189828f $X=4.927 $Y=1.852
+ $X2=0 $Y2=0
cc_1002 N_A_835_98#_c_1353_n N_A_300_464#_c_2053_n 4.87888e-19 $X=5.115 $Y=1.635
+ $X2=0 $Y2=0
cc_1003 N_A_835_98#_c_1343_n N_A_300_464#_c_2044_n 0.00777044f $X=6.02 $Y=1.225
+ $X2=0 $Y2=0
cc_1004 N_A_835_98#_c_1344_n N_A_300_464#_c_2044_n 0.00423903f $X=6.095 $Y=1.115
+ $X2=0 $Y2=0
cc_1005 N_A_835_98#_c_1355_n N_A_300_464#_c_2054_n 0.00760865f $X=5.615 $Y=3.075
+ $X2=0 $Y2=0
cc_1006 N_A_835_98#_c_1356_n N_A_300_464#_c_2054_n 0.00469098f $X=6.55 $Y=3.15
+ $X2=0 $Y2=0
cc_1007 N_A_835_98#_c_1360_n N_A_300_464#_c_2054_n 4.59946e-19 $X=6.64 $Y=2.8
+ $X2=0 $Y2=0
cc_1008 N_A_835_98#_c_1343_n N_A_300_464#_c_2045_n 0.0119917f $X=6.02 $Y=1.225
+ $X2=0 $Y2=0
cc_1009 N_A_835_98#_c_1343_n N_A_300_464#_c_2046_n 0.00599778f $X=6.02 $Y=1.225
+ $X2=0 $Y2=0
cc_1010 N_A_835_98#_c_1353_n N_A_300_464#_c_2046_n 7.71387e-19 $X=5.115 $Y=1.635
+ $X2=0 $Y2=0
cc_1011 N_A_835_98#_c_1360_n N_A_300_464#_c_2055_n 3.77807e-19 $X=6.64 $Y=2.8
+ $X2=0 $Y2=0
cc_1012 N_A_835_98#_c_1355_n N_A_300_464#_c_2056_n 0.00126396f $X=5.615 $Y=3.075
+ $X2=0 $Y2=0
cc_1013 N_A_835_98#_c_1353_n N_A_300_464#_c_2047_n 0.00425605f $X=5.115 $Y=1.635
+ $X2=0 $Y2=0
cc_1014 N_A_835_98#_c_1374_n N_VGND_M1028_d 0.0075575f $X=4.81 $Y=1.005 $X2=0
+ $Y2=0
cc_1015 N_A_835_98#_c_1350_n N_VGND_M1028_d 0.00430243f $X=4.927 $Y=1.455 $X2=0
+ $Y2=0
cc_1016 N_A_835_98#_c_1351_n N_VGND_c_2232_n 0.0156989f $X=4.45 $Y=0.625 $X2=0
+ $Y2=0
cc_1017 N_A_835_98#_c_1342_n N_VGND_c_2233_n 0.0021556f $X=5.145 $Y=1.41 $X2=0
+ $Y2=0
cc_1018 N_A_835_98#_c_1374_n N_VGND_c_2233_n 0.0250191f $X=4.81 $Y=1.005 $X2=0
+ $Y2=0
cc_1019 N_A_835_98#_c_1351_n N_VGND_c_2233_n 0.0135218f $X=4.45 $Y=0.625 $X2=0
+ $Y2=0
cc_1020 N_A_835_98#_c_1353_n N_VGND_c_2233_n 2.25597e-19 $X=5.115 $Y=1.635 $X2=0
+ $Y2=0
cc_1021 N_A_835_98#_M1002_g N_VGND_c_2234_n 0.0018065f $X=9.785 $Y=0.58 $X2=0
+ $Y2=0
cc_1022 N_A_835_98#_c_1351_n N_VGND_c_2237_n 0.0100041f $X=4.45 $Y=0.625 $X2=0
+ $Y2=0
cc_1023 N_A_835_98#_M1002_g N_VGND_c_2242_n 0.00411612f $X=9.785 $Y=0.58 $X2=0
+ $Y2=0
cc_1024 N_A_835_98#_c_1342_n N_VGND_c_2246_n 9.10391e-19 $X=5.145 $Y=1.41 $X2=0
+ $Y2=0
cc_1025 N_A_835_98#_M1002_g N_VGND_c_2246_n 0.00752295f $X=9.785 $Y=0.58 $X2=0
+ $Y2=0
cc_1026 N_A_835_98#_c_1351_n N_VGND_c_2246_n 0.0112422f $X=4.45 $Y=0.625 $X2=0
+ $Y2=0
cc_1027 N_A_1997_272#_c_1546_n N_A_1745_74#_M1021_g 0.00755075f $X=11.175
+ $Y=0.58 $X2=0 $Y2=0
cc_1028 N_A_1997_272#_c_1549_n N_A_1745_74#_M1021_g 0.00686241f $X=11.34 $Y=0.84
+ $X2=0 $Y2=0
cc_1029 N_A_1997_272#_c_1550_n N_A_1745_74#_M1021_g 3.28981e-19 $X=11.65
+ $Y=1.445 $X2=0 $Y2=0
cc_1030 N_A_1997_272#_c_1547_n N_A_1745_74#_c_1661_n 0.0096742f $X=11.565
+ $Y=1.53 $X2=0 $Y2=0
cc_1031 N_A_1997_272#_c_1552_n N_A_1745_74#_c_1661_n 0.012401f $X=11.127 $Y=2.52
+ $X2=0 $Y2=0
cc_1032 N_A_1997_272#_c_1553_n N_A_1745_74#_c_1661_n 0.00480843f $X=11.225
+ $Y=1.53 $X2=0 $Y2=0
cc_1033 N_A_1997_272#_c_1552_n N_A_1745_74#_c_1672_n 0.00856137f $X=11.127
+ $Y=2.52 $X2=0 $Y2=0
cc_1034 N_A_1997_272#_c_1557_n N_A_1745_74#_c_1673_n 0.00688539f $X=11.11
+ $Y=2.75 $X2=0 $Y2=0
cc_1035 N_A_1997_272#_c_1552_n N_A_1745_74#_c_1673_n 0.00314773f $X=11.127
+ $Y=2.52 $X2=0 $Y2=0
cc_1036 N_A_1997_272#_c_1547_n N_A_1745_74#_c_1662_n 0.00243079f $X=11.565
+ $Y=1.53 $X2=0 $Y2=0
cc_1037 N_A_1997_272#_c_1548_n N_A_1745_74#_c_1662_n 0.00158858f $X=11.565
+ $Y=0.84 $X2=0 $Y2=0
cc_1038 N_A_1997_272#_c_1550_n N_A_1745_74#_c_1662_n 0.0150077f $X=11.65
+ $Y=1.445 $X2=0 $Y2=0
cc_1039 N_A_1997_272#_c_1545_n N_A_1745_74#_c_1663_n 0.00191851f $X=11.14
+ $Y=1.53 $X2=0 $Y2=0
cc_1040 N_A_1997_272#_c_1548_n N_A_1745_74#_c_1663_n 0.00173828f $X=11.565
+ $Y=0.84 $X2=0 $Y2=0
cc_1041 N_A_1997_272#_c_1549_n N_A_1745_74#_c_1663_n 0.00908089f $X=11.34
+ $Y=0.84 $X2=0 $Y2=0
cc_1042 N_A_1997_272#_c_1550_n N_A_1745_74#_c_1663_n 0.00419353f $X=11.65
+ $Y=1.445 $X2=0 $Y2=0
cc_1043 N_A_1997_272#_c_1553_n N_A_1745_74#_c_1663_n 0.00279652f $X=11.225
+ $Y=1.53 $X2=0 $Y2=0
cc_1044 N_A_1997_272#_c_1547_n N_A_1745_74#_c_1674_n 0.00200907f $X=11.565
+ $Y=1.53 $X2=0 $Y2=0
cc_1045 N_A_1997_272#_c_1552_n N_A_1745_74#_c_1674_n 2.62811e-19 $X=11.127
+ $Y=2.52 $X2=0 $Y2=0
cc_1046 N_A_1997_272#_c_1552_n N_A_1745_74#_c_1675_n 4.34489e-19 $X=11.127
+ $Y=2.52 $X2=0 $Y2=0
cc_1047 N_A_1997_272#_c_1546_n N_A_1745_74#_M1025_g 0.00345625f $X=11.175
+ $Y=0.58 $X2=0 $Y2=0
cc_1048 N_A_1997_272#_c_1548_n N_A_1745_74#_M1025_g 0.00399686f $X=11.565
+ $Y=0.84 $X2=0 $Y2=0
cc_1049 N_A_1997_272#_c_1550_n N_A_1745_74#_M1025_g 0.00292154f $X=11.65
+ $Y=1.445 $X2=0 $Y2=0
cc_1050 N_A_1997_272#_c_1547_n N_A_1745_74#_c_1676_n 0.00270233f $X=11.565
+ $Y=1.53 $X2=0 $Y2=0
cc_1051 N_A_1997_272#_c_1552_n N_A_1745_74#_c_1676_n 0.00843513f $X=11.127
+ $Y=2.52 $X2=0 $Y2=0
cc_1052 N_A_1997_272#_c_1556_n N_A_1745_74#_c_1677_n 0.00953641f $X=10.31
+ $Y=2.465 $X2=0 $Y2=0
cc_1053 N_A_1997_272#_M1001_g N_A_1745_74#_c_1666_n 5.63627e-19 $X=10.145
+ $Y=0.58 $X2=0 $Y2=0
cc_1054 N_A_1997_272#_c_1544_n N_A_1745_74#_c_1666_n 0.00475655f $X=10.31
+ $Y=1.84 $X2=0 $Y2=0
cc_1055 N_A_1997_272#_c_1551_n N_A_1745_74#_c_1666_n 0.0105779f $X=10.315
+ $Y=1.525 $X2=0 $Y2=0
cc_1056 N_A_1997_272#_c_1544_n N_A_1745_74#_c_1679_n 0.0112071f $X=10.31 $Y=1.84
+ $X2=0 $Y2=0
cc_1057 N_A_1997_272#_c_1555_n N_A_1745_74#_c_1679_n 0.00484392f $X=10.31
+ $Y=2.375 $X2=0 $Y2=0
cc_1058 N_A_1997_272#_c_1551_n N_A_1745_74#_c_1679_n 0.0232183f $X=10.315
+ $Y=1.525 $X2=0 $Y2=0
cc_1059 N_A_1997_272#_c_1555_n N_A_1745_74#_c_1681_n 0.011498f $X=10.31 $Y=2.375
+ $X2=0 $Y2=0
cc_1060 N_A_1997_272#_c_1556_n N_A_1745_74#_c_1681_n 0.00503711f $X=10.31
+ $Y=2.465 $X2=0 $Y2=0
cc_1061 N_A_1997_272#_M1001_g N_A_1745_74#_c_1667_n 0.00279105f $X=10.145
+ $Y=0.58 $X2=0 $Y2=0
cc_1062 N_A_1997_272#_c_1545_n N_A_1745_74#_c_1669_n 0.00534862f $X=11.14
+ $Y=1.53 $X2=0 $Y2=0
cc_1063 N_A_1997_272#_c_1547_n N_A_1745_74#_c_1669_n 0.0057529f $X=11.565
+ $Y=1.53 $X2=0 $Y2=0
cc_1064 N_A_1997_272#_c_1548_n N_A_1745_74#_c_1669_n 0.00391205f $X=11.565
+ $Y=0.84 $X2=0 $Y2=0
cc_1065 N_A_1997_272#_c_1550_n N_A_1745_74#_c_1669_n 0.0139087f $X=11.65
+ $Y=1.445 $X2=0 $Y2=0
cc_1066 N_A_1997_272#_c_1553_n N_A_1745_74#_c_1669_n 0.0134734f $X=11.225
+ $Y=1.53 $X2=0 $Y2=0
cc_1067 N_A_1997_272#_M1001_g N_A_1745_74#_c_1670_n 0.0145056f $X=10.145 $Y=0.58
+ $X2=0 $Y2=0
cc_1068 N_A_1997_272#_c_1544_n N_A_1745_74#_c_1670_n 0.00481612f $X=10.31
+ $Y=1.84 $X2=0 $Y2=0
cc_1069 N_A_1997_272#_c_1545_n N_A_1745_74#_c_1670_n 0.0525955f $X=11.14 $Y=1.53
+ $X2=0 $Y2=0
cc_1070 N_A_1997_272#_c_1549_n N_A_1745_74#_c_1670_n 0.0263803f $X=11.34 $Y=0.84
+ $X2=0 $Y2=0
cc_1071 N_A_1997_272#_c_1551_n N_A_1745_74#_c_1670_n 0.023139f $X=10.315
+ $Y=1.525 $X2=0 $Y2=0
cc_1072 N_A_1997_272#_c_1547_n N_A_2399_424#_c_1828_n 9.19806e-19 $X=11.565
+ $Y=1.53 $X2=0 $Y2=0
cc_1073 N_A_1997_272#_c_1550_n N_A_2399_424#_c_1828_n 4.60428e-19 $X=11.65
+ $Y=1.445 $X2=0 $Y2=0
cc_1074 N_A_1997_272#_c_1548_n N_A_2399_424#_c_1829_n 0.00457908f $X=11.565
+ $Y=0.84 $X2=0 $Y2=0
cc_1075 N_A_1997_272#_c_1550_n N_A_2399_424#_c_1829_n 0.0171651f $X=11.65
+ $Y=1.445 $X2=0 $Y2=0
cc_1076 N_A_1997_272#_c_1547_n N_A_2399_424#_c_1831_n 0.00962353f $X=11.565
+ $Y=1.53 $X2=0 $Y2=0
cc_1077 N_A_1997_272#_c_1550_n N_A_2399_424#_c_1831_n 0.00719431f $X=11.65
+ $Y=1.445 $X2=0 $Y2=0
cc_1078 N_A_1997_272#_c_1556_n N_VPWR_c_1881_n 0.00624782f $X=10.31 $Y=2.465
+ $X2=0 $Y2=0
cc_1079 N_A_1997_272#_c_1557_n N_VPWR_c_1881_n 0.0299967f $X=11.11 $Y=2.75 $X2=0
+ $Y2=0
cc_1080 N_A_1997_272#_c_1547_n N_VPWR_c_1882_n 0.0110039f $X=11.565 $Y=1.53
+ $X2=0 $Y2=0
cc_1081 N_A_1997_272#_c_1552_n N_VPWR_c_1882_n 0.067513f $X=11.127 $Y=2.52 $X2=0
+ $Y2=0
cc_1082 N_A_1997_272#_c_1556_n N_VPWR_c_1886_n 0.00377777f $X=10.31 $Y=2.465
+ $X2=0 $Y2=0
cc_1083 N_A_1997_272#_c_1557_n N_VPWR_c_1888_n 0.015771f $X=11.11 $Y=2.75 $X2=0
+ $Y2=0
cc_1084 N_A_1997_272#_c_1556_n N_VPWR_c_1874_n 0.00662633f $X=10.31 $Y=2.465
+ $X2=0 $Y2=0
cc_1085 N_A_1997_272#_c_1557_n N_VPWR_c_1874_n 0.0130108f $X=11.11 $Y=2.75 $X2=0
+ $Y2=0
cc_1086 N_A_1997_272#_c_1548_n N_VGND_M1025_s 0.00480139f $X=11.565 $Y=0.84
+ $X2=0 $Y2=0
cc_1087 N_A_1997_272#_M1001_g N_VGND_c_2234_n 0.01204f $X=10.145 $Y=0.58 $X2=0
+ $Y2=0
cc_1088 N_A_1997_272#_c_1546_n N_VGND_c_2234_n 0.0142227f $X=11.175 $Y=0.58
+ $X2=0 $Y2=0
cc_1089 N_A_1997_272#_c_1549_n N_VGND_c_2234_n 0.00176365f $X=11.34 $Y=0.84
+ $X2=0 $Y2=0
cc_1090 N_A_1997_272#_c_1546_n N_VGND_c_2235_n 0.0158614f $X=11.175 $Y=0.58
+ $X2=0 $Y2=0
cc_1091 N_A_1997_272#_c_1548_n N_VGND_c_2235_n 0.0143444f $X=11.565 $Y=0.84
+ $X2=0 $Y2=0
cc_1092 N_A_1997_272#_M1001_g N_VGND_c_2242_n 0.00383152f $X=10.145 $Y=0.58
+ $X2=0 $Y2=0
cc_1093 N_A_1997_272#_c_1546_n N_VGND_c_2243_n 0.0143883f $X=11.175 $Y=0.58
+ $X2=0 $Y2=0
cc_1094 N_A_1997_272#_c_1548_n N_VGND_c_2243_n 0.00329108f $X=11.565 $Y=0.84
+ $X2=0 $Y2=0
cc_1095 N_A_1997_272#_M1001_g N_VGND_c_2246_n 0.0075694f $X=10.145 $Y=0.58 $X2=0
+ $Y2=0
cc_1096 N_A_1997_272#_c_1546_n N_VGND_c_2246_n 0.0119301f $X=11.175 $Y=0.58
+ $X2=0 $Y2=0
cc_1097 N_A_1997_272#_c_1548_n N_VGND_c_2246_n 0.00670825f $X=11.565 $Y=0.84
+ $X2=0 $Y2=0
cc_1098 N_A_1745_74#_c_1662_n N_A_2399_424#_c_1828_n 0.00328297f $X=11.88
+ $Y=1.275 $X2=0 $Y2=0
cc_1099 N_A_1745_74#_c_1674_n N_A_2399_424#_c_1834_n 7.20279e-19 $X=11.83
+ $Y=1.915 $X2=0 $Y2=0
cc_1100 N_A_1745_74#_c_1675_n N_A_2399_424#_c_1834_n 0.0133065f $X=11.92
+ $Y=2.045 $X2=0 $Y2=0
cc_1101 N_A_1745_74#_M1025_g N_A_2399_424#_c_1829_n 0.0137683f $X=11.955
+ $Y=0.645 $X2=0 $Y2=0
cc_1102 N_A_1745_74#_c_1661_n N_A_2399_424#_c_1830_n 0.00247742f $X=11.32
+ $Y=1.84 $X2=0 $Y2=0
cc_1103 N_A_1745_74#_c_1674_n N_A_2399_424#_c_1830_n 0.00929958f $X=11.83
+ $Y=1.915 $X2=0 $Y2=0
cc_1104 N_A_1745_74#_c_1675_n N_A_2399_424#_c_1830_n 0.00208502f $X=11.92
+ $Y=2.045 $X2=0 $Y2=0
cc_1105 N_A_1745_74#_c_1661_n N_A_2399_424#_c_1831_n 0.00108268f $X=11.32
+ $Y=1.84 $X2=0 $Y2=0
cc_1106 N_A_1745_74#_c_1662_n N_A_2399_424#_c_1831_n 5.99943e-19 $X=11.88
+ $Y=1.275 $X2=0 $Y2=0
cc_1107 N_A_1745_74#_c_1677_n N_VPWR_c_1881_n 0.0266532f $X=10.145 $Y=2.715
+ $X2=0 $Y2=0
cc_1108 N_A_1745_74#_c_1681_n N_VPWR_c_1881_n 0.00216548f $X=10.23 $Y=2.55 $X2=0
+ $Y2=0
cc_1109 N_A_1745_74#_c_1672_n N_VPWR_c_1882_n 0.00344007f $X=11.335 $Y=2.375
+ $X2=0 $Y2=0
cc_1110 N_A_1745_74#_c_1673_n N_VPWR_c_1882_n 0.00777412f $X=11.335 $Y=2.465
+ $X2=0 $Y2=0
cc_1111 N_A_1745_74#_c_1674_n N_VPWR_c_1882_n 0.0100207f $X=11.83 $Y=1.915 $X2=0
+ $Y2=0
cc_1112 N_A_1745_74#_c_1675_n N_VPWR_c_1882_n 0.00892462f $X=11.92 $Y=2.045
+ $X2=0 $Y2=0
cc_1113 N_A_1745_74#_c_1675_n N_VPWR_c_1883_n 0.00463887f $X=11.92 $Y=2.045
+ $X2=0 $Y2=0
cc_1114 N_A_1745_74#_c_1677_n N_VPWR_c_1886_n 0.0274952f $X=10.145 $Y=2.715
+ $X2=0 $Y2=0
cc_1115 N_A_1745_74#_c_1673_n N_VPWR_c_1888_n 0.00405947f $X=11.335 $Y=2.465
+ $X2=0 $Y2=0
cc_1116 N_A_1745_74#_c_1675_n N_VPWR_c_1893_n 0.00445602f $X=11.92 $Y=2.045
+ $X2=0 $Y2=0
cc_1117 N_A_1745_74#_c_1673_n N_VPWR_c_1874_n 0.00767502f $X=11.335 $Y=2.465
+ $X2=0 $Y2=0
cc_1118 N_A_1745_74#_c_1675_n N_VPWR_c_1874_n 0.00862869f $X=11.92 $Y=2.045
+ $X2=0 $Y2=0
cc_1119 N_A_1745_74#_c_1677_n N_VPWR_c_1874_n 0.0335089f $X=10.145 $Y=2.715
+ $X2=0 $Y2=0
cc_1120 N_A_1745_74#_c_1677_n A_1993_508# 0.00423971f $X=10.145 $Y=2.715
+ $X2=-0.19 $Y2=-0.245
cc_1121 N_A_1745_74#_c_1667_n N_VGND_c_2234_n 0.0159689f $X=9.57 $Y=0.56 $X2=0
+ $Y2=0
cc_1122 N_A_1745_74#_c_1670_n N_VGND_c_2234_n 0.0191133f $X=11.065 $Y=1.185
+ $X2=0 $Y2=0
cc_1123 N_A_1745_74#_M1021_g N_VGND_c_2235_n 0.00322527f $X=10.96 $Y=0.58 $X2=0
+ $Y2=0
cc_1124 N_A_1745_74#_c_1662_n N_VGND_c_2235_n 0.00195495f $X=11.88 $Y=1.275
+ $X2=0 $Y2=0
cc_1125 N_A_1745_74#_M1025_g N_VGND_c_2235_n 0.00927494f $X=11.955 $Y=0.645
+ $X2=0 $Y2=0
cc_1126 N_A_1745_74#_M1025_g N_VGND_c_2236_n 0.00296233f $X=11.955 $Y=0.645
+ $X2=0 $Y2=0
cc_1127 N_A_1745_74#_c_1667_n N_VGND_c_2242_n 0.0151251f $X=9.57 $Y=0.56 $X2=0
+ $Y2=0
cc_1128 N_A_1745_74#_M1021_g N_VGND_c_2243_n 0.00434272f $X=10.96 $Y=0.58 $X2=0
+ $Y2=0
cc_1129 N_A_1745_74#_M1025_g N_VGND_c_2244_n 0.00383152f $X=11.955 $Y=0.645
+ $X2=0 $Y2=0
cc_1130 N_A_1745_74#_M1021_g N_VGND_c_2246_n 0.00825669f $X=10.96 $Y=0.58 $X2=0
+ $Y2=0
cc_1131 N_A_1745_74#_M1025_g N_VGND_c_2246_n 0.00762539f $X=11.955 $Y=0.645
+ $X2=0 $Y2=0
cc_1132 N_A_1745_74#_c_1667_n N_VGND_c_2246_n 0.0125365f $X=9.57 $Y=0.56 $X2=0
+ $Y2=0
cc_1133 N_A_2399_424#_c_1834_n N_VPWR_c_1882_n 0.0345631f $X=12.145 $Y=2.265
+ $X2=0 $Y2=0
cc_1134 N_A_2399_424#_c_1832_n N_VPWR_c_1883_n 0.0215785f $X=12.93 $Y=1.765
+ $X2=0 $Y2=0
cc_1135 N_A_2399_424#_c_1828_n N_VPWR_c_1883_n 0.00731242f $X=12.84 $Y=1.465
+ $X2=0 $Y2=0
cc_1136 N_A_2399_424#_c_1854_p N_VPWR_c_1883_n 0.0253438f $X=12.745 $Y=1.465
+ $X2=0 $Y2=0
cc_1137 N_A_2399_424#_c_1830_n N_VPWR_c_1883_n 0.0776081f $X=12.145 $Y=2.1 $X2=0
+ $Y2=0
cc_1138 N_A_2399_424#_c_1834_n N_VPWR_c_1893_n 0.0145938f $X=12.145 $Y=2.265
+ $X2=0 $Y2=0
cc_1139 N_A_2399_424#_c_1832_n N_VPWR_c_1894_n 0.00413917f $X=12.93 $Y=1.765
+ $X2=0 $Y2=0
cc_1140 N_A_2399_424#_c_1832_n N_VPWR_c_1874_n 0.00821237f $X=12.93 $Y=1.765
+ $X2=0 $Y2=0
cc_1141 N_A_2399_424#_c_1834_n N_VPWR_c_1874_n 0.0120466f $X=12.145 $Y=2.265
+ $X2=0 $Y2=0
cc_1142 N_A_2399_424#_M1004_g Q 0.00853833f $X=12.945 $Y=0.74 $X2=0 $Y2=0
cc_1143 N_A_2399_424#_M1004_g Q 0.00339956f $X=12.945 $Y=0.74 $X2=0 $Y2=0
cc_1144 N_A_2399_424#_c_1832_n Q 0.00791945f $X=12.93 $Y=1.765 $X2=0 $Y2=0
cc_1145 N_A_2399_424#_M1004_g Q 0.0228636f $X=12.945 $Y=0.74 $X2=0 $Y2=0
cc_1146 N_A_2399_424#_c_1854_p Q 0.0238691f $X=12.745 $Y=1.465 $X2=0 $Y2=0
cc_1147 N_A_2399_424#_c_1829_n N_VGND_c_2235_n 0.00917009f $X=12.17 $Y=0.645
+ $X2=0 $Y2=0
cc_1148 N_A_2399_424#_M1004_g N_VGND_c_2236_n 0.00647412f $X=12.945 $Y=0.74
+ $X2=0 $Y2=0
cc_1149 N_A_2399_424#_c_1828_n N_VGND_c_2236_n 0.00577732f $X=12.84 $Y=1.465
+ $X2=0 $Y2=0
cc_1150 N_A_2399_424#_c_1829_n N_VGND_c_2236_n 0.0504216f $X=12.17 $Y=0.645
+ $X2=0 $Y2=0
cc_1151 N_A_2399_424#_c_1854_p N_VGND_c_2236_n 0.0209147f $X=12.745 $Y=1.465
+ $X2=0 $Y2=0
cc_1152 N_A_2399_424#_c_1829_n N_VGND_c_2244_n 0.011066f $X=12.17 $Y=0.645 $X2=0
+ $Y2=0
cc_1153 N_A_2399_424#_M1004_g N_VGND_c_2245_n 0.00434272f $X=12.945 $Y=0.74
+ $X2=0 $Y2=0
cc_1154 N_A_2399_424#_M1004_g N_VGND_c_2246_n 0.00828941f $X=12.945 $Y=0.74
+ $X2=0 $Y2=0
cc_1155 N_A_2399_424#_c_1829_n N_VGND_c_2246_n 0.00915947f $X=12.17 $Y=0.645
+ $X2=0 $Y2=0
cc_1156 N_VPWR_c_1875_n N_A_300_464#_c_2049_n 0.0195202f $X=0.78 $Y=2.465 $X2=0
+ $Y2=0
cc_1157 N_VPWR_c_1891_n N_A_300_464#_c_2049_n 0.0471516f $X=3.095 $Y=3.33 $X2=0
+ $Y2=0
cc_1158 N_VPWR_c_1874_n N_A_300_464#_c_2049_n 0.0391751f $X=13.2 $Y=3.33 $X2=0
+ $Y2=0
cc_1159 N_VPWR_M1026_d N_A_300_464#_c_2072_n 0.0104311f $X=3.11 $Y=2.32 $X2=0
+ $Y2=0
cc_1160 N_VPWR_c_1876_n N_A_300_464#_c_2072_n 0.0214041f $X=3.26 $Y=2.79 $X2=0
+ $Y2=0
cc_1161 N_VPWR_c_1874_n N_A_300_464#_c_2072_n 0.0190648f $X=13.2 $Y=3.33 $X2=0
+ $Y2=0
cc_1162 N_VPWR_c_1884_n N_A_300_464#_c_2051_n 0.00543175f $X=4.705 $Y=3.33 $X2=0
+ $Y2=0
cc_1163 N_VPWR_c_1874_n N_A_300_464#_c_2051_n 0.0102994f $X=13.2 $Y=3.33 $X2=0
+ $Y2=0
cc_1164 N_VPWR_M1026_d N_A_300_464#_c_2052_n 8.43866e-19 $X=3.11 $Y=2.32 $X2=0
+ $Y2=0
cc_1165 N_VPWR_c_1884_n N_A_300_464#_c_2052_n 0.00409815f $X=4.705 $Y=3.33 $X2=0
+ $Y2=0
cc_1166 N_VPWR_c_1874_n N_A_300_464#_c_2052_n 0.0145667f $X=13.2 $Y=3.33 $X2=0
+ $Y2=0
cc_1167 N_VPWR_M1027_d N_A_300_464#_c_2053_n 0.00387164f $X=4.72 $Y=1.96 $X2=0
+ $Y2=0
cc_1168 N_VPWR_c_1877_n N_A_300_464#_c_2053_n 0.0167709f $X=4.87 $Y=2.835 $X2=0
+ $Y2=0
cc_1169 N_VPWR_c_1884_n N_A_300_464#_c_2053_n 7.54393e-19 $X=4.705 $Y=3.33 $X2=0
+ $Y2=0
cc_1170 N_VPWR_c_1892_n N_A_300_464#_c_2053_n 0.0103722f $X=7.205 $Y=3.33 $X2=0
+ $Y2=0
cc_1171 N_VPWR_c_1874_n N_A_300_464#_c_2053_n 0.0213354f $X=13.2 $Y=3.33 $X2=0
+ $Y2=0
cc_1172 N_VPWR_c_1892_n N_A_300_464#_c_2054_n 0.00535093f $X=7.205 $Y=3.33 $X2=0
+ $Y2=0
cc_1173 N_VPWR_c_1874_n N_A_300_464#_c_2054_n 0.00675054f $X=13.2 $Y=3.33 $X2=0
+ $Y2=0
cc_1174 N_VPWR_c_1876_n N_A_300_464#_c_2058_n 0.00906648f $X=3.26 $Y=2.79 $X2=0
+ $Y2=0
cc_1175 N_VPWR_c_1876_n N_A_300_464#_c_2059_n 0.0176069f $X=3.26 $Y=2.79 $X2=0
+ $Y2=0
cc_1176 N_VPWR_c_1884_n N_A_300_464#_c_2059_n 0.0144865f $X=4.705 $Y=3.33 $X2=0
+ $Y2=0
cc_1177 N_VPWR_c_1874_n N_A_300_464#_c_2059_n 0.012005f $X=13.2 $Y=3.33 $X2=0
+ $Y2=0
cc_1178 N_VPWR_c_1883_n Q 0.0779559f $X=12.705 $Y=1.985 $X2=0 $Y2=0
cc_1179 N_VPWR_c_1894_n Q 0.0112891f $X=13.2 $Y=3.33 $X2=0 $Y2=0
cc_1180 N_VPWR_c_1874_n Q 0.00934413f $X=13.2 $Y=3.33 $X2=0 $Y2=0
cc_1181 N_A_300_464#_c_2072_n A_535_464# 0.00940297f $X=3.445 $Y=2.43 $X2=-0.19
+ $Y2=-0.245
cc_1182 N_A_300_464#_M1006_d N_noxref_24_c_2364_n 0.0106902f $X=1.95 $Y=0.405
+ $X2=0 $Y2=0
cc_1183 N_A_300_464#_c_2041_n N_noxref_24_c_2364_n 0.0126305f $X=3.445 $Y=1.005
+ $X2=0 $Y2=0
cc_1184 N_A_300_464#_c_2048_n N_noxref_24_c_2364_n 0.019982f $X=2.435 $Y=0.68
+ $X2=0 $Y2=0
cc_1185 N_A_300_464#_c_2041_n N_noxref_24_c_2366_n 0.0234737f $X=3.445 $Y=1.005
+ $X2=0 $Y2=0
cc_1186 N_A_300_464#_c_2048_n N_noxref_24_c_2366_n 0.00520956f $X=2.435 $Y=0.68
+ $X2=0 $Y2=0
cc_1187 Q N_VGND_c_2236_n 0.0293763f $X=13.115 $Y=0.47 $X2=0 $Y2=0
cc_1188 Q N_VGND_c_2245_n 0.0145639f $X=13.115 $Y=0.47 $X2=0 $Y2=0
cc_1189 Q N_VGND_c_2246_n 0.0119984f $X=13.115 $Y=0.47 $X2=0 $Y2=0
cc_1190 N_VGND_c_2240_n N_noxref_24_c_2364_n 0.10468f $X=3.59 $Y=0 $X2=0 $Y2=0
cc_1191 N_VGND_c_2246_n N_noxref_24_c_2364_n 0.0610965f $X=13.2 $Y=0 $X2=0 $Y2=0
cc_1192 N_VGND_c_2231_n N_noxref_24_c_2365_n 0.0259562f $X=0.71 $Y=0.65 $X2=0
+ $Y2=0
cc_1193 N_VGND_c_2240_n N_noxref_24_c_2365_n 0.0225398f $X=3.59 $Y=0 $X2=0 $Y2=0
cc_1194 N_VGND_c_2246_n N_noxref_24_c_2365_n 0.0125704f $X=13.2 $Y=0 $X2=0 $Y2=0
cc_1195 N_VGND_c_2232_n N_noxref_24_c_2366_n 0.0118481f $X=3.715 $Y=0.565 $X2=0
+ $Y2=0
cc_1196 N_VGND_c_2240_n N_noxref_24_c_2366_n 0.0243596f $X=3.59 $Y=0 $X2=0 $Y2=0
cc_1197 N_VGND_c_2246_n N_noxref_24_c_2366_n 0.0134194f $X=13.2 $Y=0 $X2=0 $Y2=0
cc_1198 N_noxref_24_c_2364_n noxref_25 0.00198134f $X=3.06 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_1199 N_noxref_24_c_2364_n noxref_26 0.00226367f $X=3.06 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
