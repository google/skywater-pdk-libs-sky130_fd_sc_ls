# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ls__dfsbp_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ls__dfsbp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  12.96000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.475000 0.980000 0.805000 1.990000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.065000 1.820000 12.425000 2.980000 ;
        RECT 12.085000 0.350000 12.425000 1.130000 ;
        RECT 12.255000 1.130000 12.425000 1.820000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.130000 1.820000 10.435000 2.970000 ;
        RECT 10.175000 0.350000 10.435000 1.820000 ;
    END
  END Q_N
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.225000 1.580000 5.635000 2.020000 ;
        RECT 8.285000 1.180000 8.640000 1.780000 ;
      LAYER mcon ;
        RECT 5.435000 1.580000 5.605000 1.750000 ;
        RECT 8.315000 1.580000 8.485000 1.750000 ;
      LAYER met1 ;
        RECT 5.375000 1.550000 5.665000 1.595000 ;
        RECT 5.375000 1.595000 8.545000 1.735000 ;
        RECT 5.375000 1.735000 5.665000 1.780000 ;
        RECT 8.255000 1.550000 8.545000 1.595000 ;
        RECT 8.255000 1.735000 8.545000 1.780000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.315000 1.180000 1.775000 1.550000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 12.960000 0.085000 ;
        RECT  0.545000  0.085000  0.795000 0.810000 ;
        RECT  1.605000  0.085000  1.865000 1.010000 ;
        RECT  3.990000  0.085000  4.240000 0.845000 ;
        RECT  5.340000  0.085000  6.160000 0.680000 ;
        RECT  8.100000  0.085000  8.845000 0.670000 ;
        RECT  9.665000  0.085000  9.995000 0.840000 ;
        RECT 10.605000  0.085000 10.855000 1.130000 ;
        RECT 11.585000  0.085000 11.915000 1.030000 ;
        RECT 12.595000  0.085000 12.845000 1.130000 ;
      LAYER mcon ;
        RECT  0.155000 -0.085000  0.325000 0.085000 ;
        RECT  0.635000 -0.085000  0.805000 0.085000 ;
        RECT  1.115000 -0.085000  1.285000 0.085000 ;
        RECT  1.595000 -0.085000  1.765000 0.085000 ;
        RECT  2.075000 -0.085000  2.245000 0.085000 ;
        RECT  2.555000 -0.085000  2.725000 0.085000 ;
        RECT  3.035000 -0.085000  3.205000 0.085000 ;
        RECT  3.515000 -0.085000  3.685000 0.085000 ;
        RECT  3.995000 -0.085000  4.165000 0.085000 ;
        RECT  4.475000 -0.085000  4.645000 0.085000 ;
        RECT  4.955000 -0.085000  5.125000 0.085000 ;
        RECT  5.435000 -0.085000  5.605000 0.085000 ;
        RECT  5.915000 -0.085000  6.085000 0.085000 ;
        RECT  6.395000 -0.085000  6.565000 0.085000 ;
        RECT  6.875000 -0.085000  7.045000 0.085000 ;
        RECT  7.355000 -0.085000  7.525000 0.085000 ;
        RECT  7.835000 -0.085000  8.005000 0.085000 ;
        RECT  8.315000 -0.085000  8.485000 0.085000 ;
        RECT  8.795000 -0.085000  8.965000 0.085000 ;
        RECT  9.275000 -0.085000  9.445000 0.085000 ;
        RECT  9.755000 -0.085000  9.925000 0.085000 ;
        RECT 10.235000 -0.085000 10.405000 0.085000 ;
        RECT 10.715000 -0.085000 10.885000 0.085000 ;
        RECT 11.195000 -0.085000 11.365000 0.085000 ;
        RECT 11.675000 -0.085000 11.845000 0.085000 ;
        RECT 12.155000 -0.085000 12.325000 0.085000 ;
        RECT 12.635000 -0.085000 12.805000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 12.960000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 3.245000 12.960000 3.415000 ;
        RECT  0.565000 2.530000  0.895000 3.245000 ;
        RECT  1.575000 2.530000  1.905000 3.245000 ;
        RECT  4.020000 2.735000  4.350000 3.245000 ;
        RECT  5.700000 2.530000  6.070000 3.245000 ;
        RECT  8.090000 2.650000  8.260000 3.245000 ;
        RECT  9.630000 2.630000  9.960000 3.245000 ;
        RECT 10.605000 1.820000 10.860000 3.245000 ;
        RECT 11.615000 1.820000 11.865000 3.245000 ;
        RECT 12.595000 1.820000 12.845000 3.245000 ;
      LAYER mcon ;
        RECT  0.155000 3.245000  0.325000 3.415000 ;
        RECT  0.635000 3.245000  0.805000 3.415000 ;
        RECT  1.115000 3.245000  1.285000 3.415000 ;
        RECT  1.595000 3.245000  1.765000 3.415000 ;
        RECT  2.075000 3.245000  2.245000 3.415000 ;
        RECT  2.555000 3.245000  2.725000 3.415000 ;
        RECT  3.035000 3.245000  3.205000 3.415000 ;
        RECT  3.515000 3.245000  3.685000 3.415000 ;
        RECT  3.995000 3.245000  4.165000 3.415000 ;
        RECT  4.475000 3.245000  4.645000 3.415000 ;
        RECT  4.955000 3.245000  5.125000 3.415000 ;
        RECT  5.435000 3.245000  5.605000 3.415000 ;
        RECT  5.915000 3.245000  6.085000 3.415000 ;
        RECT  6.395000 3.245000  6.565000 3.415000 ;
        RECT  6.875000 3.245000  7.045000 3.415000 ;
        RECT  7.355000 3.245000  7.525000 3.415000 ;
        RECT  7.835000 3.245000  8.005000 3.415000 ;
        RECT  8.315000 3.245000  8.485000 3.415000 ;
        RECT  8.795000 3.245000  8.965000 3.415000 ;
        RECT  9.275000 3.245000  9.445000 3.415000 ;
        RECT  9.755000 3.245000  9.925000 3.415000 ;
        RECT 10.235000 3.245000 10.405000 3.415000 ;
        RECT 10.715000 3.245000 10.885000 3.415000 ;
        RECT 11.195000 3.245000 11.365000 3.415000 ;
        RECT 11.675000 3.245000 11.845000 3.415000 ;
        RECT 12.155000 3.245000 12.325000 3.415000 ;
        RECT 12.635000 3.245000 12.805000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 12.960000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.115000 0.350000  0.365000 0.810000 ;
      RECT  0.115000 0.810000  0.285000 2.190000 ;
      RECT  0.115000 2.190000  2.615000 2.230000 ;
      RECT  0.115000 2.230000  1.795000 2.360000 ;
      RECT  0.115000 2.360000  0.365000 2.980000 ;
      RECT  0.975000 0.350000  1.435000 1.010000 ;
      RECT  0.975000 1.010000  1.145000 1.720000 ;
      RECT  0.975000 1.720000  2.275000 1.890000 ;
      RECT  0.975000 1.890000  1.455000 2.020000 ;
      RECT  1.625000 2.060000  2.615000 2.190000 ;
      RECT  1.945000 1.300000  2.275000 1.720000 ;
      RECT  2.045000 0.255000  3.110000 0.425000 ;
      RECT  2.045000 0.425000  2.215000 1.130000 ;
      RECT  2.105000 2.400000  2.275000 2.905000 ;
      RECT  2.105000 2.905000  3.845000 3.075000 ;
      RECT  2.445000 0.595000  2.770000 0.925000 ;
      RECT  2.445000 0.925000  2.615000 2.060000 ;
      RECT  2.445000 2.230000  2.615000 2.295000 ;
      RECT  2.445000 2.295000  2.865000 2.735000 ;
      RECT  2.785000 1.435000  3.115000 2.105000 ;
      RECT  2.940000 0.425000  3.110000 1.435000 ;
      RECT  3.065000 2.295000  3.455000 2.735000 ;
      RECT  3.280000 0.465000  3.530000 0.925000 ;
      RECT  3.285000 0.925000  3.530000 1.095000 ;
      RECT  3.285000 1.095000  4.185000 1.265000 ;
      RECT  3.285000 1.265000  3.455000 2.295000 ;
      RECT  3.625000 1.435000  3.845000 2.395000 ;
      RECT  3.625000 2.395000  4.690000 2.565000 ;
      RECT  3.625000 2.565000  3.845000 2.905000 ;
      RECT  4.015000 1.265000  4.185000 1.515000 ;
      RECT  4.015000 1.515000  5.015000 1.685000 ;
      RECT  4.140000 1.855000  4.470000 2.055000 ;
      RECT  4.140000 2.055000  5.030000 2.225000 ;
      RECT  4.355000 1.015000  4.580000 1.345000 ;
      RECT  4.410000 0.350000  4.880000 1.015000 ;
      RECT  4.520000 2.565000  4.690000 2.905000 ;
      RECT  4.520000 2.905000  5.530000 3.075000 ;
      RECT  4.750000 1.240000  5.915000 1.410000 ;
      RECT  4.750000 1.410000  5.015000 1.515000 ;
      RECT  4.750000 1.685000  5.015000 1.885000 ;
      RECT  4.860000 2.225000  5.030000 2.295000 ;
      RECT  4.860000 2.295000  5.190000 2.735000 ;
      RECT  5.360000 2.190000  6.500000 2.360000 ;
      RECT  5.360000 2.360000  5.530000 2.905000 ;
      RECT  5.585000 1.120000  5.915000 1.240000 ;
      RECT  6.330000 0.280000  7.555000 0.450000 ;
      RECT  6.330000 0.450000  6.500000 1.120000 ;
      RECT  6.330000 1.120000  6.875000 1.450000 ;
      RECT  6.330000 1.450000  6.500000 2.190000 ;
      RECT  6.670000 0.620000  7.215000 0.950000 ;
      RECT  6.780000 1.680000  7.215000 1.850000 ;
      RECT  6.780000 1.850000  7.030000 2.480000 ;
      RECT  6.780000 2.480000  7.920000 2.650000 ;
      RECT  6.780000 2.650000  7.470000 2.980000 ;
      RECT  7.045000 0.950000  7.215000 1.680000 ;
      RECT  7.250000 2.020000  7.580000 2.310000 ;
      RECT  7.385000 0.450000  7.555000 2.020000 ;
      RECT  7.725000 0.840000  9.435000 1.010000 ;
      RECT  7.725000 1.010000  8.055000 1.780000 ;
      RECT  7.750000 1.950000  9.570000 2.120000 ;
      RECT  7.750000 2.120000  8.790000 2.480000 ;
      RECT  8.460000 2.480000  8.790000 2.915000 ;
      RECT  8.900000 1.350000  9.570000 1.950000 ;
      RECT  9.015000 2.290000  9.910000 2.460000 ;
      RECT  9.015000 2.460000  9.345000 2.620000 ;
      RECT  9.105000 0.635000  9.435000 0.840000 ;
      RECT  9.105000 1.010000  9.910000 1.180000 ;
      RECT  9.740000 1.180000  9.910000 2.290000 ;
      RECT 11.085000 0.350000 11.415000 1.300000 ;
      RECT 11.085000 1.300000 12.085000 1.630000 ;
      RECT 11.085000 1.630000 11.415000 2.860000 ;
  END
END sky130_fd_sc_ls__dfsbp_2
