# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ls__dlrbp_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ls__dlrbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.160000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.208500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.435000 1.450000 0.805000 1.780000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.130000 0.350000 6.460000 1.010000 ;
        RECT 6.130000 1.010000 6.670000 1.180000 ;
        RECT 6.200000 2.060000 6.670000 2.980000 ;
        RECT 6.500000 1.180000 6.670000 2.060000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.604200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.710000 0.350000 8.055000 1.040000 ;
        RECT 7.715000 1.820000 8.055000 2.980000 ;
        RECT 7.885000 1.040000 8.055000 1.820000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.425000 1.180000 5.795000 1.550000 ;
    END
  END RESET_B
  PIN GATE
    ANTENNAGATEAREA  0.237000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.975000 1.450000 1.305000 1.780000 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 8.160000 0.085000 ;
        RECT 0.625000  0.085000 0.955000 1.280000 ;
        RECT 2.320000  0.085000 2.650000 0.410000 ;
        RECT 4.240000  0.085000 4.570000 1.060000 ;
        RECT 5.620000  0.085000 5.950000 1.010000 ;
        RECT 7.200000  0.085000 7.530000 0.940000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
        RECT 6.395000 -0.085000 6.565000 0.085000 ;
        RECT 6.875000 -0.085000 7.045000 0.085000 ;
        RECT 7.355000 -0.085000 7.525000 0.085000 ;
        RECT 7.835000 -0.085000 8.005000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.160000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 8.160000 3.415000 ;
        RECT 0.650000 2.730000 0.980000 3.245000 ;
        RECT 2.350000 2.730000 2.685000 3.245000 ;
        RECT 4.405000 2.650000 5.080000 3.245000 ;
        RECT 5.780000 2.060000 6.030000 3.245000 ;
        RECT 7.210000 2.100000 7.540000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
        RECT 6.395000 3.245000 6.565000 3.415000 ;
        RECT 6.875000 3.245000 7.045000 3.415000 ;
        RECT 7.355000 3.245000 7.525000 3.415000 ;
        RECT 7.835000 3.245000 8.005000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 8.160000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.095000 0.690000 0.445000 1.280000 ;
      RECT 0.095000 1.280000 0.265000 1.970000 ;
      RECT 0.095000 1.970000 0.445000 2.390000 ;
      RECT 0.095000 2.390000 2.675000 2.560000 ;
      RECT 0.095000 2.560000 0.445000 2.850000 ;
      RECT 1.185000 0.500000 1.645000 0.580000 ;
      RECT 1.185000 0.580000 2.990000 0.750000 ;
      RECT 1.185000 0.750000 1.645000 1.280000 ;
      RECT 1.185000 1.970000 1.645000 2.220000 ;
      RECT 1.475000 1.280000 1.645000 1.420000 ;
      RECT 1.475000 1.420000 1.875000 1.750000 ;
      RECT 1.475000 1.750000 1.645000 1.970000 ;
      RECT 1.815000 1.940000 2.215000 2.220000 ;
      RECT 1.825000 0.920000 2.215000 1.130000 ;
      RECT 1.825000 1.130000 3.395000 1.250000 ;
      RECT 2.045000 1.250000 3.395000 1.300000 ;
      RECT 2.045000 1.300000 2.215000 1.940000 ;
      RECT 2.505000 1.470000 2.835000 1.800000 ;
      RECT 2.505000 1.800000 2.675000 2.390000 ;
      RECT 2.820000 0.255000 3.905000 0.510000 ;
      RECT 2.820000 0.510000 2.990000 0.580000 ;
      RECT 2.855000 1.970000 3.175000 2.140000 ;
      RECT 2.855000 2.140000 3.025000 2.905000 ;
      RECT 2.855000 2.905000 4.015000 3.075000 ;
      RECT 3.005000 1.300000 3.395000 1.480000 ;
      RECT 3.005000 1.480000 3.175000 1.970000 ;
      RECT 3.190000 0.710000 3.750000 0.960000 ;
      RECT 3.195000 2.405000 3.515000 2.735000 ;
      RECT 3.345000 1.650000 4.915000 1.820000 ;
      RECT 3.345000 1.820000 3.515000 2.405000 ;
      RECT 3.580000 0.960000 3.750000 1.650000 ;
      RECT 3.685000 2.050000 4.015000 2.905000 ;
      RECT 4.225000 1.990000 5.580000 2.320000 ;
      RECT 4.585000 1.350000 4.915000 1.650000 ;
      RECT 4.800000 0.350000 5.255000 1.130000 ;
      RECT 5.085000 1.130000 5.255000 1.720000 ;
      RECT 5.085000 1.720000 6.330000 1.890000 ;
      RECT 5.085000 1.890000 5.580000 1.990000 ;
      RECT 5.250000 2.320000 5.580000 2.980000 ;
      RECT 6.005000 1.350000 6.330000 1.720000 ;
      RECT 6.690000 0.350000 7.020000 0.840000 ;
      RECT 6.840000 0.840000 7.020000 1.320000 ;
      RECT 6.840000 1.320000 7.715000 1.650000 ;
      RECT 6.840000 1.650000 7.010000 2.980000 ;
  END
END sky130_fd_sc_ls__dlrbp_1
