* File: sky130_fd_sc_ls__nor2b_1.pxi.spice
* Created: Wed Sep  2 11:14:20 2020
* 
x_PM_SKY130_FD_SC_LS__NOR2B_1%B_N N_B_N_c_40_n N_B_N_M1003_g N_B_N_c_41_n
+ N_B_N_M1004_g N_B_N_c_42_n B_N PM_SKY130_FD_SC_LS__NOR2B_1%B_N
x_PM_SKY130_FD_SC_LS__NOR2B_1%A N_A_c_67_n N_A_M1002_g N_A_c_68_n N_A_M1005_g A
+ PM_SKY130_FD_SC_LS__NOR2B_1%A
x_PM_SKY130_FD_SC_LS__NOR2B_1%A_27_112# N_A_27_112#_M1004_s N_A_27_112#_M1003_s
+ N_A_27_112#_c_97_n N_A_27_112#_M1000_g N_A_27_112#_M1001_g N_A_27_112#_c_107_n
+ N_A_27_112#_c_102_n N_A_27_112#_c_99_n N_A_27_112#_c_104_n N_A_27_112#_c_105_n
+ N_A_27_112#_c_100_n PM_SKY130_FD_SC_LS__NOR2B_1%A_27_112#
x_PM_SKY130_FD_SC_LS__NOR2B_1%VPWR N_VPWR_M1003_d N_VPWR_c_161_n VPWR
+ N_VPWR_c_162_n N_VPWR_c_163_n N_VPWR_c_160_n N_VPWR_c_165_n
+ PM_SKY130_FD_SC_LS__NOR2B_1%VPWR
x_PM_SKY130_FD_SC_LS__NOR2B_1%Y N_Y_M1005_d N_Y_M1000_d N_Y_c_185_n N_Y_c_186_n
+ N_Y_c_187_n Y Y Y N_Y_c_190_n N_Y_c_188_n Y PM_SKY130_FD_SC_LS__NOR2B_1%Y
x_PM_SKY130_FD_SC_LS__NOR2B_1%VGND N_VGND_M1004_d N_VGND_M1001_d N_VGND_c_216_n
+ N_VGND_c_217_n N_VGND_c_218_n N_VGND_c_219_n N_VGND_c_220_n VGND
+ N_VGND_c_221_n N_VGND_c_222_n PM_SKY130_FD_SC_LS__NOR2B_1%VGND
cc_1 VNB N_B_N_c_40_n 0.0198761f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=1.765
cc_2 VNB N_B_N_c_41_n 0.0233618f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.22
cc_3 VNB N_B_N_c_42_n 0.0628724f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.385
cc_4 VNB B_N 0.017759f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_5 VNB N_A_c_67_n 0.0438471f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=1.765
cc_6 VNB N_A_c_68_n 0.0201157f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.22
cc_7 VNB A 0.00407508f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=1.385
cc_8 VNB N_A_27_112#_c_97_n 0.0348031f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=1.385
cc_9 VNB N_A_27_112#_M1001_g 0.0253088f $X=-0.19 $Y=-0.245 $X2=0.275 $Y2=1.385
cc_10 VNB N_A_27_112#_c_99_n 0.00853715f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_27_112#_c_100_n 0.0111198f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_VPWR_c_160_n 0.103974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_Y_c_185_n 0.00208979f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_14 VNB N_Y_c_186_n 0.012465f $X=-0.19 $Y=-0.245 $X2=0.275 $Y2=1.385
cc_15 VNB N_Y_c_187_n 0.00221952f $X=-0.19 $Y=-0.245 $X2=0.275 $Y2=1.385
cc_16 VNB N_Y_c_188_n 0.0242534f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_VGND_c_216_n 0.0131348f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_18 VNB N_VGND_c_217_n 0.0129133f $X=-0.19 $Y=-0.245 $X2=0.275 $Y2=1.385
cc_19 VNB N_VGND_c_218_n 0.011907f $X=-0.19 $Y=-0.245 $X2=0.275 $Y2=1.385
cc_20 VNB N_VGND_c_219_n 0.0302402f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_220_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_221_n 0.0193208f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_222_n 0.178959f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VPB N_B_N_c_40_n 0.0284988f $X=-0.19 $Y=1.66 $X2=0.705 $Y2=1.765
cc_25 VPB N_A_c_67_n 0.0233735f $X=-0.19 $Y=1.66 $X2=0.705 $Y2=1.765
cc_26 VPB N_A_27_112#_c_97_n 0.0261384f $X=-0.19 $Y=1.66 $X2=0.705 $Y2=1.385
cc_27 VPB N_A_27_112#_c_102_n 0.0349344f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_28 VPB N_A_27_112#_c_99_n 0.00202686f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_29 VPB N_A_27_112#_c_104_n 0.0141291f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_30 VPB N_A_27_112#_c_105_n 0.0101533f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_31 VPB N_A_27_112#_c_100_n 5.62371e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_32 VPB N_VPWR_c_161_n 0.0171513f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=0.835
cc_33 VPB N_VPWR_c_162_n 0.0301039f $X=-0.19 $Y=1.66 $X2=0.275 $Y2=1.385
cc_34 VPB N_VPWR_c_163_n 0.0349999f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_35 VPB N_VPWR_c_160_n 0.081687f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_36 VPB N_VPWR_c_165_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_37 VPB Y 0.0449044f $X=-0.19 $Y=1.66 $X2=0.275 $Y2=1.295
cc_38 VPB N_Y_c_190_n 0.0129713f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_39 VPB N_Y_c_188_n 0.00785541f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_40 N_B_N_c_40_n N_A_c_67_n 0.0348946f $X=0.705 $Y=1.765 $X2=-0.19 $Y2=-0.245
cc_41 N_B_N_c_41_n N_A_c_68_n 0.0094315f $X=0.72 $Y=1.22 $X2=0 $Y2=0
cc_42 N_B_N_c_40_n A 8.64176e-19 $X=0.705 $Y=1.765 $X2=0 $Y2=0
cc_43 N_B_N_c_41_n A 3.04755e-19 $X=0.72 $Y=1.22 $X2=0 $Y2=0
cc_44 N_B_N_c_41_n N_A_27_112#_c_107_n 0.00851666f $X=0.72 $Y=1.22 $X2=0 $Y2=0
cc_45 N_B_N_c_42_n N_A_27_112#_c_107_n 0.00741677f $X=0.615 $Y=1.385 $X2=0 $Y2=0
cc_46 B_N N_A_27_112#_c_107_n 0.0152451f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_47 N_B_N_c_40_n N_A_27_112#_c_102_n 0.0151932f $X=0.705 $Y=1.765 $X2=0 $Y2=0
cc_48 N_B_N_c_40_n N_A_27_112#_c_99_n 0.0142882f $X=0.705 $Y=1.765 $X2=0 $Y2=0
cc_49 N_B_N_c_41_n N_A_27_112#_c_99_n 0.00809053f $X=0.72 $Y=1.22 $X2=0 $Y2=0
cc_50 N_B_N_c_42_n N_A_27_112#_c_99_n 0.0046103f $X=0.615 $Y=1.385 $X2=0 $Y2=0
cc_51 B_N N_A_27_112#_c_99_n 0.026737f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_52 N_B_N_c_40_n N_A_27_112#_c_104_n 0.00128638f $X=0.705 $Y=1.765 $X2=0 $Y2=0
cc_53 N_B_N_c_40_n N_A_27_112#_c_105_n 0.0142951f $X=0.705 $Y=1.765 $X2=0 $Y2=0
cc_54 N_B_N_c_42_n N_A_27_112#_c_105_n 0.00858089f $X=0.615 $Y=1.385 $X2=0 $Y2=0
cc_55 B_N N_A_27_112#_c_105_n 0.0105909f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_56 N_B_N_c_40_n N_VPWR_c_161_n 0.00901804f $X=0.705 $Y=1.765 $X2=0 $Y2=0
cc_57 N_B_N_c_40_n N_VPWR_c_162_n 0.00393873f $X=0.705 $Y=1.765 $X2=0 $Y2=0
cc_58 N_B_N_c_40_n N_VPWR_c_160_n 0.00462577f $X=0.705 $Y=1.765 $X2=0 $Y2=0
cc_59 N_B_N_c_41_n N_VGND_c_216_n 0.00905753f $X=0.72 $Y=1.22 $X2=0 $Y2=0
cc_60 N_B_N_c_41_n N_VGND_c_219_n 0.00360585f $X=0.72 $Y=1.22 $X2=0 $Y2=0
cc_61 N_B_N_c_41_n N_VGND_c_222_n 0.00487769f $X=0.72 $Y=1.22 $X2=0 $Y2=0
cc_62 N_A_c_67_n N_A_27_112#_c_97_n 0.0820914f $X=1.315 $Y=1.765 $X2=0 $Y2=0
cc_63 A N_A_27_112#_c_97_n 2.21841e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_64 N_A_c_68_n N_A_27_112#_M1001_g 0.0219036f $X=1.33 $Y=1.22 $X2=0 $Y2=0
cc_65 A N_A_27_112#_M1001_g 7.63572e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_66 N_A_c_67_n N_A_27_112#_c_102_n 4.75567e-19 $X=1.315 $Y=1.765 $X2=0 $Y2=0
cc_67 N_A_c_67_n N_A_27_112#_c_99_n 0.00323847f $X=1.315 $Y=1.765 $X2=0 $Y2=0
cc_68 N_A_c_68_n N_A_27_112#_c_99_n 6.54906e-19 $X=1.33 $Y=1.22 $X2=0 $Y2=0
cc_69 A N_A_27_112#_c_99_n 0.0199505f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_70 N_A_c_67_n N_A_27_112#_c_104_n 0.0188422f $X=1.315 $Y=1.765 $X2=0 $Y2=0
cc_71 A N_A_27_112#_c_104_n 0.0244703f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_72 N_A_c_67_n N_A_27_112#_c_100_n 0.00565934f $X=1.315 $Y=1.765 $X2=0 $Y2=0
cc_73 A N_A_27_112#_c_100_n 0.0187161f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_74 N_A_c_67_n N_VPWR_c_161_n 0.0216963f $X=1.315 $Y=1.765 $X2=0 $Y2=0
cc_75 N_A_c_67_n N_VPWR_c_163_n 0.00413917f $X=1.315 $Y=1.765 $X2=0 $Y2=0
cc_76 N_A_c_67_n N_VPWR_c_160_n 0.00817532f $X=1.315 $Y=1.765 $X2=0 $Y2=0
cc_77 N_A_c_68_n N_Y_c_185_n 0.00516456f $X=1.33 $Y=1.22 $X2=0 $Y2=0
cc_78 N_A_c_68_n N_Y_c_187_n 0.00443842f $X=1.33 $Y=1.22 $X2=0 $Y2=0
cc_79 N_A_c_67_n N_VGND_c_216_n 0.00139337f $X=1.315 $Y=1.765 $X2=0 $Y2=0
cc_80 N_A_c_68_n N_VGND_c_216_n 0.0139704f $X=1.33 $Y=1.22 $X2=0 $Y2=0
cc_81 A N_VGND_c_216_n 0.0185651f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_82 N_A_c_68_n N_VGND_c_221_n 0.00383152f $X=1.33 $Y=1.22 $X2=0 $Y2=0
cc_83 N_A_c_68_n N_VGND_c_222_n 0.00758292f $X=1.33 $Y=1.22 $X2=0 $Y2=0
cc_84 N_A_27_112#_c_104_n N_VPWR_M1003_d 0.00631766f $X=1.535 $Y=1.805 $X2=-0.19
+ $Y2=-0.245
cc_85 N_A_27_112#_c_97_n N_VPWR_c_161_n 0.00328565f $X=1.735 $Y=1.765 $X2=0
+ $Y2=0
cc_86 N_A_27_112#_c_102_n N_VPWR_c_161_n 0.0339233f $X=0.48 $Y=1.985 $X2=0 $Y2=0
cc_87 N_A_27_112#_c_104_n N_VPWR_c_161_n 0.0219335f $X=1.535 $Y=1.805 $X2=0
+ $Y2=0
cc_88 N_A_27_112#_c_102_n N_VPWR_c_162_n 0.0066794f $X=0.48 $Y=1.985 $X2=0 $Y2=0
cc_89 N_A_27_112#_c_97_n N_VPWR_c_163_n 0.00461464f $X=1.735 $Y=1.765 $X2=0
+ $Y2=0
cc_90 N_A_27_112#_c_97_n N_VPWR_c_160_n 0.00913435f $X=1.735 $Y=1.765 $X2=0
+ $Y2=0
cc_91 N_A_27_112#_c_102_n N_VPWR_c_160_n 0.00997343f $X=0.48 $Y=1.985 $X2=0
+ $Y2=0
cc_92 N_A_27_112#_c_104_n A_278_368# 0.00331953f $X=1.535 $Y=1.805 $X2=-0.19
+ $Y2=-0.245
cc_93 N_A_27_112#_c_100_n A_278_368# 0.00300337f $X=1.81 $Y=1.485 $X2=-0.19
+ $Y2=-0.245
cc_94 N_A_27_112#_M1001_g N_Y_c_185_n 0.0130905f $X=1.835 $Y=0.74 $X2=0 $Y2=0
cc_95 N_A_27_112#_c_97_n N_Y_c_186_n 4.58216e-19 $X=1.735 $Y=1.765 $X2=0 $Y2=0
cc_96 N_A_27_112#_M1001_g N_Y_c_186_n 0.0127588f $X=1.835 $Y=0.74 $X2=0 $Y2=0
cc_97 N_A_27_112#_c_100_n N_Y_c_186_n 0.0138485f $X=1.81 $Y=1.485 $X2=0 $Y2=0
cc_98 N_A_27_112#_c_97_n N_Y_c_187_n 9.00201e-19 $X=1.735 $Y=1.765 $X2=0 $Y2=0
cc_99 N_A_27_112#_M1001_g N_Y_c_187_n 0.00116669f $X=1.835 $Y=0.74 $X2=0 $Y2=0
cc_100 N_A_27_112#_c_100_n N_Y_c_187_n 0.0221208f $X=1.81 $Y=1.485 $X2=0 $Y2=0
cc_101 N_A_27_112#_c_97_n N_Y_c_190_n 0.0161624f $X=1.735 $Y=1.765 $X2=0 $Y2=0
cc_102 N_A_27_112#_c_100_n N_Y_c_190_n 0.0143134f $X=1.81 $Y=1.485 $X2=0 $Y2=0
cc_103 N_A_27_112#_c_97_n N_Y_c_188_n 0.00546429f $X=1.735 $Y=1.765 $X2=0 $Y2=0
cc_104 N_A_27_112#_M1001_g N_Y_c_188_n 0.00539566f $X=1.835 $Y=0.74 $X2=0 $Y2=0
cc_105 N_A_27_112#_c_100_n N_Y_c_188_n 0.031807f $X=1.81 $Y=1.485 $X2=0 $Y2=0
cc_106 N_A_27_112#_M1001_g N_VGND_c_216_n 6.08003e-19 $X=1.835 $Y=0.74 $X2=0
+ $Y2=0
cc_107 N_A_27_112#_c_107_n N_VGND_c_216_n 0.02666f $X=0.61 $Y=0.845 $X2=0 $Y2=0
cc_108 N_A_27_112#_M1001_g N_VGND_c_218_n 0.00521557f $X=1.835 $Y=0.74 $X2=0
+ $Y2=0
cc_109 N_A_27_112#_c_107_n N_VGND_c_219_n 0.00820401f $X=0.61 $Y=0.845 $X2=0
+ $Y2=0
cc_110 N_A_27_112#_M1001_g N_VGND_c_221_n 0.00434272f $X=1.835 $Y=0.74 $X2=0
+ $Y2=0
cc_111 N_A_27_112#_M1001_g N_VGND_c_222_n 0.00824687f $X=1.835 $Y=0.74 $X2=0
+ $Y2=0
cc_112 N_A_27_112#_c_107_n N_VGND_c_222_n 0.0148718f $X=0.61 $Y=0.845 $X2=0
+ $Y2=0
cc_113 N_VPWR_c_161_n Y 0.0262913f $X=1.09 $Y=2.145 $X2=0 $Y2=0
cc_114 N_VPWR_c_163_n Y 0.019544f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_115 N_VPWR_c_160_n Y 0.0161768f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_116 N_Y_c_186_n N_VGND_M1001_d 0.00568412f $X=2.145 $Y=1.065 $X2=0 $Y2=0
cc_117 N_Y_c_185_n N_VGND_c_216_n 0.0350754f $X=1.62 $Y=0.515 $X2=0 $Y2=0
cc_118 N_Y_c_187_n N_VGND_c_216_n 0.00181371f $X=1.785 $Y=1.065 $X2=0 $Y2=0
cc_119 N_Y_c_185_n N_VGND_c_218_n 0.0173103f $X=1.62 $Y=0.515 $X2=0 $Y2=0
cc_120 N_Y_c_186_n N_VGND_c_218_n 0.0220189f $X=2.145 $Y=1.065 $X2=0 $Y2=0
cc_121 N_Y_c_185_n N_VGND_c_221_n 0.0109942f $X=1.62 $Y=0.515 $X2=0 $Y2=0
cc_122 N_Y_c_185_n N_VGND_c_222_n 0.00904371f $X=1.62 $Y=0.515 $X2=0 $Y2=0
