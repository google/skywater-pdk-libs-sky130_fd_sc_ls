* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__dlrtn_2 D GATE_N RESET_B VGND VNB VPB VPWR Q
M1000 VGND RESET_B a_1153_74# VNB nshort w=740000u l=150000u
+  ad=2.30995e+12p pd=1.387e+07u as=1.776e+11p ps=1.96e+06u
M1001 a_232_98# GATE_N VGND VNB nshort w=740000u l=150000u
+  ad=2.257e+11p pd=2.09e+06u as=0p ps=0u
M1002 a_1153_74# a_670_392# a_913_406# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1003 Q a_913_406# VGND VNB nshort w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1004 VGND a_232_98# a_373_82# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.294e+11p ps=2.1e+06u
M1005 a_670_392# a_373_82# a_586_392# VPB phighvt w=1e+06u l=150000u
+  ad=3.371e+11p pd=2.78e+06u as=2.7e+11p ps=2.54e+06u
M1006 Q a_913_406# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=2.7852e+12p ps=1.673e+07u
M1007 VGND a_913_406# Q VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_697_74# a_27_136# VGND VNB nshort w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1009 a_670_392# a_232_98# a_697_74# VNB nshort w=640000u l=150000u
+  ad=1.915e+11p pd=1.93e+06u as=0p ps=0u
M1010 VPWR a_913_406# a_778_504# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=2.898e+11p ps=2.22e+06u
M1011 a_586_392# a_27_136# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR a_913_406# Q VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND D a_27_136# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1014 VPWR D a_27_136# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=2.478e+11p ps=2.27e+06u
M1015 VGND a_913_406# a_870_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.155e+11p ps=1.39e+06u
M1016 VPWR a_232_98# a_373_82# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=2.478e+11p ps=2.27e+06u
M1017 a_913_406# a_670_392# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.472e+11p pd=2.86e+06u as=0p ps=0u
M1018 VPWR RESET_B a_913_406# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_870_74# a_373_82# a_670_392# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_778_504# a_232_98# a_670_392# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_232_98# GATE_N VPWR VPB phighvt w=840000u l=150000u
+  ad=2.478e+11p pd=2.27e+06u as=0p ps=0u
.ends
