* File: sky130_fd_sc_ls__dfsbp_2.pxi.spice
* Created: Wed Sep  2 11:01:35 2020
* 
x_PM_SKY130_FD_SC_LS__DFSBP_2%D N_D_c_278_n N_D_c_283_n N_D_M1027_g N_D_c_284_n
+ N_D_M1017_g D D N_D_c_280_n N_D_c_281_n N_D_c_286_n
+ PM_SKY130_FD_SC_LS__DFSBP_2%D
x_PM_SKY130_FD_SC_LS__DFSBP_2%CLK N_CLK_c_313_n N_CLK_M1031_g N_CLK_c_314_n
+ N_CLK_M1029_g CLK PM_SKY130_FD_SC_LS__DFSBP_2%CLK
x_PM_SKY130_FD_SC_LS__DFSBP_2%A_398_74# N_A_398_74#_M1015_d N_A_398_74#_M1002_d
+ N_A_398_74#_c_346_n N_A_398_74#_c_365_n N_A_398_74#_c_366_n
+ N_A_398_74#_M1003_g N_A_398_74#_c_347_n N_A_398_74#_M1034_g
+ N_A_398_74#_M1018_g N_A_398_74#_c_368_n N_A_398_74#_M1013_g
+ N_A_398_74#_c_349_n N_A_398_74#_c_468_p N_A_398_74#_c_350_n
+ N_A_398_74#_c_351_n N_A_398_74#_c_369_n N_A_398_74#_c_370_n
+ N_A_398_74#_c_352_n N_A_398_74#_c_353_n N_A_398_74#_c_354_n
+ N_A_398_74#_c_374_n N_A_398_74#_c_386_p N_A_398_74#_c_375_n
+ N_A_398_74#_c_376_n N_A_398_74#_c_377_n N_A_398_74#_c_378_n
+ N_A_398_74#_c_379_n N_A_398_74#_c_380_n N_A_398_74#_c_355_n
+ N_A_398_74#_c_356_n N_A_398_74#_c_357_n N_A_398_74#_c_358_n
+ N_A_398_74#_c_359_n N_A_398_74#_c_388_p N_A_398_74#_c_360_n
+ N_A_398_74#_c_361_n N_A_398_74#_c_382_n N_A_398_74#_c_362_n
+ N_A_398_74#_c_363_n PM_SKY130_FD_SC_LS__DFSBP_2%A_398_74#
x_PM_SKY130_FD_SC_LS__DFSBP_2%A_757_401# N_A_757_401#_M1026_s
+ N_A_757_401#_M1005_d N_A_757_401#_c_626_n N_A_757_401#_M1004_g
+ N_A_757_401#_c_621_n N_A_757_401#_M1022_g N_A_757_401#_c_627_n
+ N_A_757_401#_c_622_n N_A_757_401#_c_623_n N_A_757_401#_c_628_n
+ N_A_757_401#_c_629_n N_A_757_401#_c_630_n N_A_757_401#_c_631_n
+ N_A_757_401#_c_624_n N_A_757_401#_c_632_n N_A_757_401#_c_625_n
+ PM_SKY130_FD_SC_LS__DFSBP_2%A_757_401#
x_PM_SKY130_FD_SC_LS__DFSBP_2%A_595_97# N_A_595_97#_M1014_d N_A_595_97#_M1003_d
+ N_A_595_97#_c_731_n N_A_595_97#_c_732_n N_A_595_97#_M1005_g
+ N_A_595_97#_M1026_g N_A_595_97#_c_714_n N_A_595_97#_c_715_n
+ N_A_595_97#_c_734_n N_A_595_97#_M1032_g N_A_595_97#_c_716_n
+ N_A_595_97#_M1008_g N_A_595_97#_c_717_n N_A_595_97#_c_718_n
+ N_A_595_97#_c_719_n N_A_595_97#_c_720_n N_A_595_97#_c_721_n
+ N_A_595_97#_c_722_n N_A_595_97#_c_723_n N_A_595_97#_c_724_n
+ N_A_595_97#_c_738_n N_A_595_97#_c_781_n N_A_595_97#_c_725_n
+ N_A_595_97#_c_726_n N_A_595_97#_c_727_n N_A_595_97#_c_728_n
+ N_A_595_97#_c_729_n N_A_595_97#_c_730_n PM_SKY130_FD_SC_LS__DFSBP_2%A_595_97#
x_PM_SKY130_FD_SC_LS__DFSBP_2%SET_B N_SET_B_M1023_g N_SET_B_c_884_n
+ N_SET_B_c_898_n N_SET_B_M1036_g N_SET_B_c_885_n N_SET_B_M1037_g
+ N_SET_B_c_886_n N_SET_B_c_887_n N_SET_B_c_888_n N_SET_B_c_900_n
+ N_SET_B_M1021_g N_SET_B_c_889_n N_SET_B_c_890_n N_SET_B_c_891_n
+ N_SET_B_c_892_n N_SET_B_c_893_n SET_B N_SET_B_c_895_n N_SET_B_c_896_n
+ PM_SKY130_FD_SC_LS__DFSBP_2%SET_B
x_PM_SKY130_FD_SC_LS__DFSBP_2%A_225_74# N_A_225_74#_M1031_s N_A_225_74#_M1029_s
+ N_A_225_74#_M1015_g N_A_225_74#_c_1009_n N_A_225_74#_M1002_g
+ N_A_225_74#_c_1021_n N_A_225_74#_c_1010_n N_A_225_74#_c_1022_n
+ N_A_225_74#_c_1023_n N_A_225_74#_M1014_g N_A_225_74#_c_1024_n
+ N_A_225_74#_c_1025_n N_A_225_74#_c_1026_n N_A_225_74#_M1012_g
+ N_A_225_74#_c_1027_n N_A_225_74#_M1033_g N_A_225_74#_c_1012_n
+ N_A_225_74#_c_1013_n N_A_225_74#_M1035_g N_A_225_74#_c_1015_n
+ N_A_225_74#_c_1016_n N_A_225_74#_c_1033_n N_A_225_74#_c_1017_n
+ N_A_225_74#_c_1035_n N_A_225_74#_c_1036_n N_A_225_74#_c_1037_n
+ N_A_225_74#_c_1018_n N_A_225_74#_c_1019_n N_A_225_74#_c_1039_n
+ PM_SKY130_FD_SC_LS__DFSBP_2%A_225_74#
x_PM_SKY130_FD_SC_LS__DFSBP_2%A_1501_92# N_A_1501_92#_M1000_d
+ N_A_1501_92#_M1007_s N_A_1501_92#_M1019_g N_A_1501_92#_c_1203_n
+ N_A_1501_92#_c_1204_n N_A_1501_92#_M1010_g N_A_1501_92#_c_1198_n
+ N_A_1501_92#_c_1199_n N_A_1501_92#_c_1235_n N_A_1501_92#_c_1218_n
+ N_A_1501_92#_c_1207_n N_A_1501_92#_c_1200_n N_A_1501_92#_c_1201_n
+ N_A_1501_92#_c_1209_n N_A_1501_92#_c_1202_n
+ PM_SKY130_FD_SC_LS__DFSBP_2%A_1501_92#
x_PM_SKY130_FD_SC_LS__DFSBP_2%A_1339_74# N_A_1339_74#_M1018_d
+ N_A_1339_74#_M1033_d N_A_1339_74#_M1021_d N_A_1339_74#_M1000_g
+ N_A_1339_74#_c_1306_n N_A_1339_74#_c_1307_n N_A_1339_74#_c_1320_n
+ N_A_1339_74#_M1007_g N_A_1339_74#_c_1308_n N_A_1339_74#_c_1321_n
+ N_A_1339_74#_M1024_g N_A_1339_74#_M1009_g N_A_1339_74#_c_1322_n
+ N_A_1339_74#_M1028_g N_A_1339_74#_M1020_g N_A_1339_74#_c_1311_n
+ N_A_1339_74#_c_1312_n N_A_1339_74#_M1006_g N_A_1339_74#_c_1324_n
+ N_A_1339_74#_M1030_g N_A_1339_74#_c_1314_n N_A_1339_74#_c_1336_n
+ N_A_1339_74#_c_1326_n N_A_1339_74#_c_1315_n N_A_1339_74#_c_1327_n
+ N_A_1339_74#_c_1316_n N_A_1339_74#_c_1329_n N_A_1339_74#_c_1330_n
+ N_A_1339_74#_c_1331_n N_A_1339_74#_c_1332_n N_A_1339_74#_c_1333_n
+ N_A_1339_74#_c_1317_n PM_SKY130_FD_SC_LS__DFSBP_2%A_1339_74#
x_PM_SKY130_FD_SC_LS__DFSBP_2%A_2221_74# N_A_2221_74#_M1006_s
+ N_A_2221_74#_M1030_s N_A_2221_74#_c_1506_n N_A_2221_74#_M1016_g
+ N_A_2221_74#_M1001_g N_A_2221_74#_c_1507_n N_A_2221_74#_M1025_g
+ N_A_2221_74#_M1011_g N_A_2221_74#_c_1501_n N_A_2221_74#_c_1502_n
+ N_A_2221_74#_c_1503_n N_A_2221_74#_c_1504_n N_A_2221_74#_c_1505_n
+ PM_SKY130_FD_SC_LS__DFSBP_2%A_2221_74#
x_PM_SKY130_FD_SC_LS__DFSBP_2%A_27_74# N_A_27_74#_M1027_s N_A_27_74#_M1014_s
+ N_A_27_74#_M1017_s N_A_27_74#_M1003_s N_A_27_74#_c_1570_n N_A_27_74#_c_1571_n
+ N_A_27_74#_c_1576_n N_A_27_74#_c_1577_n N_A_27_74#_c_1578_n
+ N_A_27_74#_c_1572_n N_A_27_74#_c_1573_n N_A_27_74#_c_1580_n
+ N_A_27_74#_c_1623_n N_A_27_74#_c_1574_n PM_SKY130_FD_SC_LS__DFSBP_2%A_27_74#
x_PM_SKY130_FD_SC_LS__DFSBP_2%VPWR N_VPWR_M1017_d N_VPWR_M1029_d N_VPWR_M1004_d
+ N_VPWR_M1036_d N_VPWR_M1010_d N_VPWR_M1007_d N_VPWR_M1028_d N_VPWR_M1030_d
+ N_VPWR_M1025_s N_VPWR_c_1641_n N_VPWR_c_1642_n N_VPWR_c_1643_n N_VPWR_c_1644_n
+ N_VPWR_c_1645_n N_VPWR_c_1646_n N_VPWR_c_1647_n N_VPWR_c_1648_n
+ N_VPWR_c_1649_n N_VPWR_c_1650_n N_VPWR_c_1651_n N_VPWR_c_1652_n
+ N_VPWR_c_1653_n N_VPWR_c_1654_n VPWR N_VPWR_c_1655_n N_VPWR_c_1656_n
+ N_VPWR_c_1657_n N_VPWR_c_1658_n N_VPWR_c_1659_n N_VPWR_c_1660_n
+ N_VPWR_c_1661_n N_VPWR_c_1662_n N_VPWR_c_1663_n N_VPWR_c_1664_n
+ N_VPWR_c_1665_n N_VPWR_c_1666_n N_VPWR_c_1667_n N_VPWR_c_1640_n
+ PM_SKY130_FD_SC_LS__DFSBP_2%VPWR
x_PM_SKY130_FD_SC_LS__DFSBP_2%Q_N N_Q_N_M1009_d N_Q_N_M1024_s Q_N Q_N Q_N Q_N
+ Q_N Q_N PM_SKY130_FD_SC_LS__DFSBP_2%Q_N
x_PM_SKY130_FD_SC_LS__DFSBP_2%Q N_Q_M1001_s N_Q_M1016_d N_Q_c_1824_n
+ N_Q_c_1825_n N_Q_c_1821_n Q Q Q PM_SKY130_FD_SC_LS__DFSBP_2%Q
x_PM_SKY130_FD_SC_LS__DFSBP_2%VGND N_VGND_M1027_d N_VGND_M1031_d N_VGND_M1022_d
+ N_VGND_M1023_d N_VGND_M1037_d N_VGND_M1009_s N_VGND_M1020_s N_VGND_M1006_d
+ N_VGND_M1011_d N_VGND_c_1853_n N_VGND_c_1854_n N_VGND_c_1855_n N_VGND_c_1856_n
+ N_VGND_c_1857_n N_VGND_c_1858_n N_VGND_c_1859_n N_VGND_c_1860_n
+ N_VGND_c_1861_n N_VGND_c_1862_n N_VGND_c_1863_n VGND N_VGND_c_1864_n
+ N_VGND_c_1865_n N_VGND_c_1866_n N_VGND_c_1867_n N_VGND_c_1868_n
+ N_VGND_c_1869_n N_VGND_c_1870_n N_VGND_c_1871_n N_VGND_c_1872_n
+ N_VGND_c_1873_n N_VGND_c_1874_n N_VGND_c_1875_n N_VGND_c_1876_n
+ N_VGND_c_1877_n N_VGND_c_1878_n PM_SKY130_FD_SC_LS__DFSBP_2%VGND
cc_1 VNB N_D_c_278_n 0.0447809f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.795
cc_2 VNB N_D_M1027_g 0.0283644f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.58
cc_3 VNB N_D_c_280_n 0.025337f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.145
cc_4 VNB N_D_c_281_n 0.00250659f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.145
cc_5 VNB N_CLK_c_313_n 0.0199636f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.175
cc_6 VNB N_CLK_c_314_n 0.0361334f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.375
cc_7 VNB CLK 0.00845272f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.58
cc_8 VNB N_A_398_74#_c_346_n 0.0152453f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.58
cc_9 VNB N_A_398_74#_c_347_n 0.0218688f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_10 VNB N_A_398_74#_M1034_g 0.0428034f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.145
cc_11 VNB N_A_398_74#_c_349_n 0.00150841f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.295
cc_12 VNB N_A_398_74#_c_350_n 0.0225218f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_398_74#_c_351_n 0.00264685f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_398_74#_c_352_n 0.00184302f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_398_74#_c_353_n 0.0017748f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_398_74#_c_354_n 0.0180595f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_398_74#_c_355_n 0.00252917f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_398_74#_c_356_n 0.00213435f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_398_74#_c_357_n 0.0185305f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_398_74#_c_358_n 0.00189911f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_398_74#_c_359_n 0.00652496f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_398_74#_c_360_n 0.00733674f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_398_74#_c_361_n 0.0309266f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_398_74#_c_362_n 0.00534817f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_398_74#_c_363_n 0.0194713f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_757_401#_c_621_n 0.0184264f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.75
cc_27 VNB N_A_757_401#_c_622_n 0.0584491f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_757_401#_c_623_n 0.00815564f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.145
cc_29 VNB N_A_757_401#_c_624_n 0.018262f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.825
cc_30 VNB N_A_757_401#_c_625_n 0.0154979f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_595_97#_M1026_g 0.0511561f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_595_97#_c_714_n 0.0160274f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.145
cc_33 VNB N_A_595_97#_c_715_n 0.0157366f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.98
cc_34 VNB N_A_595_97#_c_716_n 0.021832f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.99
cc_35 VNB N_A_595_97#_c_717_n 0.00650115f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.295
cc_36 VNB N_A_595_97#_c_718_n 0.00248621f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_595_97#_c_719_n 0.0013452f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_595_97#_c_720_n 0.00289252f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_595_97#_c_721_n 0.0134003f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_595_97#_c_722_n 0.00439152f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_595_97#_c_723_n 0.00427182f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_595_97#_c_724_n 8.90541e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_595_97#_c_725_n 0.00213571f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_595_97#_c_726_n 0.00547595f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_595_97#_c_727_n 0.00856216f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_595_97#_c_728_n 0.00247208f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_595_97#_c_729_n 0.0185631f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_595_97#_c_730_n 0.0380798f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_SET_B_c_884_n 0.0341432f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.98
cc_50 VNB N_SET_B_c_885_n 0.016029f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.465
cc_51 VNB N_SET_B_c_886_n 0.0185076f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_52 VNB N_SET_B_c_887_n 0.00564647f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_53 VNB N_SET_B_c_888_n 0.00734157f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_SET_B_c_889_n 0.0186942f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.98
cc_55 VNB N_SET_B_c_890_n 0.012641f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.825
cc_56 VNB N_SET_B_c_891_n 0.0137927f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.825
cc_57 VNB N_SET_B_c_892_n 0.00275558f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.825
cc_58 VNB N_SET_B_c_893_n 0.00127012f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB SET_B 6.91838e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_SET_B_c_895_n 0.0405859f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_SET_B_c_896_n 0.00406556f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_225_74#_M1015_g 0.0224523f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.465
cc_63 VNB N_A_225_74#_c_1009_n 0.0123708f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.75
cc_64 VNB N_A_225_74#_c_1010_n 0.0289831f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.145
cc_65 VNB N_A_225_74#_M1014_g 0.0210047f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.825
cc_66 VNB N_A_225_74#_c_1012_n 0.00841887f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_225_74#_c_1013_n 8.10901e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_225_74#_M1035_g 0.0446676f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_225_74#_c_1015_n 0.0254751f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_225_74#_c_1016_n 0.0195076f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_225_74#_c_1017_n 0.0104758f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_225_74#_c_1018_n 0.00365457f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_225_74#_c_1019_n 0.0130637f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_1501_92#_M1019_g 0.0323321f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.465
cc_75 VNB N_A_1501_92#_c_1198_n 0.00698987f $X=-0.19 $Y=-0.245 $X2=0.64
+ $Y2=1.145
cc_76 VNB N_A_1501_92#_c_1199_n 0.0327285f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.98
cc_77 VNB N_A_1501_92#_c_1200_n 0.0133421f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_1501_92#_c_1201_n 0.00405333f $X=-0.19 $Y=-0.245 $X2=0.64
+ $Y2=1.665
cc_79 VNB N_A_1501_92#_c_1202_n 0.0100146f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_1339_74#_M1000_g 0.0361264f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_81 VNB N_A_1339_74#_c_1306_n 0.0185463f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_1339_74#_c_1307_n 0.00960128f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_1339_74#_c_1308_n 0.0297435f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.98
cc_84 VNB N_A_1339_74#_M1009_g 0.0259325f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.295
cc_85 VNB N_A_1339_74#_M1020_g 0.0258655f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_1339_74#_c_1311_n 0.0759793f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_1339_74#_c_1312_n 0.0332441f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_1339_74#_M1006_g 0.0364692f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_1339_74#_c_1314_n 0.0109531f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_1339_74#_c_1315_n 0.00581877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_1339_74#_c_1316_n 0.00629293f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_1339_74#_c_1317_n 0.0116128f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_2221_74#_M1001_g 0.0230317f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_94 VNB N_A_2221_74#_M1011_g 0.0260184f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.98
cc_95 VNB N_A_2221_74#_c_1501_n 0.0123246f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.99
cc_96 VNB N_A_2221_74#_c_1502_n 3.56488e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_2221_74#_c_1503_n 0.0072339f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_A_2221_74#_c_1504_n 6.27903e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_A_2221_74#_c_1505_n 0.0736247f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_A_27_74#_c_1570_n 0.0146704f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_A_27_74#_c_1571_n 0.040185f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.145
cc_102 VNB N_A_27_74#_c_1572_n 0.00621313f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.665
cc_103 VNB N_A_27_74#_c_1573_n 0.00791533f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_A_27_74#_c_1574_n 0.00628546f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_VPWR_c_1640_n 0.541827f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB Q_N 0.00397681f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.58
cc_107 VNB N_Q_c_1821_n 0.00141953f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB Q 0.00240191f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.145
cc_109 VNB Q 0.00429087f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.145
cc_110 VNB N_VGND_c_1853_n 0.0077412f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.825
cc_111 VNB N_VGND_c_1854_n 0.0221343f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_1855_n 0.00564229f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_1856_n 0.0119517f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_1857_n 0.0176142f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_VGND_c_1858_n 0.0194608f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_VGND_c_1859_n 0.0112908f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_VGND_c_1860_n 0.010678f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_VGND_c_1861_n 0.0505285f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_VGND_c_1862_n 0.0171743f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_VGND_c_1863_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_VGND_c_1864_n 0.0173909f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_VGND_c_1865_n 0.0558487f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB N_VGND_c_1866_n 0.0245702f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_VGND_c_1867_n 0.0206041f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_1868_n 0.0189349f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_1869_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_VGND_c_1870_n 0.00481148f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_1871_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_1872_n 0.0311101f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_1873_n 0.0239278f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_1874_n 0.0493081f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_VGND_c_1875_n 0.0419048f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_VGND_c_1876_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_VGND_c_1877_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_VGND_c_1878_n 0.720699f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VPB N_D_c_278_n 0.0126976f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.795
cc_137 VPB N_D_c_283_n 0.0313518f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.375
cc_138 VPB N_D_c_284_n 0.0313209f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.465
cc_139 VPB N_D_c_281_n 0.00207792f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.145
cc_140 VPB N_D_c_286_n 0.0244664f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.825
cc_141 VPB N_CLK_c_314_n 0.0230735f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.375
cc_142 VPB N_A_398_74#_c_346_n 0.00815295f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.58
cc_143 VPB N_A_398_74#_c_365_n 0.0405022f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_144 VPB N_A_398_74#_c_366_n 0.0141711f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.465
cc_145 VPB N_A_398_74#_c_347_n 0.016956f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_146 VPB N_A_398_74#_c_368_n 0.0666525f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.825
cc_147 VPB N_A_398_74#_c_369_n 0.022414f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_148 VPB N_A_398_74#_c_370_n 0.00314412f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_149 VPB N_A_398_74#_c_352_n 0.00298749f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_150 VPB N_A_398_74#_c_353_n 0.00605175f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_151 VPB N_A_398_74#_c_354_n 0.0223789f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_152 VPB N_A_398_74#_c_374_n 0.00196411f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_153 VPB N_A_398_74#_c_375_n 0.00401063f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_154 VPB N_A_398_74#_c_376_n 0.0154208f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_155 VPB N_A_398_74#_c_377_n 0.00260501f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_156 VPB N_A_398_74#_c_378_n 0.00197994f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_157 VPB N_A_398_74#_c_379_n 0.00567462f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_158 VPB N_A_398_74#_c_380_n 6.92221e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_159 VPB N_A_398_74#_c_356_n 0.0042866f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_160 VPB N_A_398_74#_c_382_n 0.00176185f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_161 VPB N_A_398_74#_c_362_n 0.00577418f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_162 VPB N_A_757_401#_c_626_n 0.0143184f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.58
cc_163 VPB N_A_757_401#_c_627_n 0.012156f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_164 VPB N_A_757_401#_c_628_n 0.0176706f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=0.98
cc_165 VPB N_A_757_401#_c_629_n 0.00575682f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.825
cc_166 VPB N_A_757_401#_c_630_n 0.00369936f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.145
cc_167 VPB N_A_757_401#_c_631_n 0.0358692f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_168 VPB N_A_757_401#_c_632_n 0.0111833f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_169 VPB N_A_757_401#_c_625_n 0.0114856f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_170 VPB N_A_595_97#_c_731_n 0.0141168f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_171 VPB N_A_595_97#_c_732_n 0.0229683f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.465
cc_172 VPB N_A_595_97#_c_715_n 0.00124104f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=0.98
cc_173 VPB N_A_595_97#_c_734_n 0.0239255f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.825
cc_174 VPB N_A_595_97#_c_720_n 0.0076856f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_175 VPB N_A_595_97#_c_723_n 0.00348451f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_176 VPB N_A_595_97#_c_724_n 0.00251531f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_177 VPB N_A_595_97#_c_738_n 0.00296251f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_178 VPB N_A_595_97#_c_726_n 0.00116107f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_179 VPB N_A_595_97#_c_727_n 0.0227484f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_180 VPB N_SET_B_c_884_n 0.00480279f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.98
cc_181 VPB N_SET_B_c_898_n 0.0696341f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.58
cc_182 VPB N_SET_B_c_888_n 0.0437509f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_183 VPB N_SET_B_c_900_n 0.0266701f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.145
cc_184 VPB N_SET_B_c_891_n 0.0194185f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.825
cc_185 VPB N_SET_B_c_892_n 0.00103414f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.825
cc_186 VPB N_SET_B_c_893_n 0.00776991f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_187 VPB SET_B 0.00113364f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_188 VPB N_SET_B_c_896_n 0.00291878f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_189 VPB N_A_225_74#_c_1009_n 0.0210337f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.75
cc_190 VPB N_A_225_74#_c_1021_n 0.0744152f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_191 VPB N_A_225_74#_c_1022_n 0.0524229f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.145
cc_192 VPB N_A_225_74#_c_1023_n 0.0125859f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=0.98
cc_193 VPB N_A_225_74#_c_1024_n 0.00736242f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.145
cc_194 VPB N_A_225_74#_c_1025_n 0.0131636f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_195 VPB N_A_225_74#_c_1026_n 0.0134614f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.295
cc_196 VPB N_A_225_74#_c_1027_n 0.255448f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_197 VPB N_A_225_74#_M1033_g 0.0103307f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_198 VPB N_A_225_74#_c_1012_n 0.0321991f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_199 VPB N_A_225_74#_c_1013_n 0.0139489f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_200 VPB N_A_225_74#_c_1015_n 5.35904e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_201 VPB N_A_225_74#_c_1016_n 0.011123f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_202 VPB N_A_225_74#_c_1033_n 0.0089864f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_203 VPB N_A_225_74#_c_1017_n 0.00236347f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_204 VPB N_A_225_74#_c_1035_n 0.00592994f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_205 VPB N_A_225_74#_c_1036_n 0.00539283f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_206 VPB N_A_225_74#_c_1037_n 0.00468204f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_207 VPB N_A_225_74#_c_1018_n 5.33031e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_208 VPB N_A_225_74#_c_1039_n 8.57544e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_209 VPB N_A_1501_92#_c_1203_n 0.0304315f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_210 VPB N_A_1501_92#_c_1204_n 0.020379f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_211 VPB N_A_1501_92#_c_1198_n 0.00214188f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.145
cc_212 VPB N_A_1501_92#_c_1199_n 0.0128253f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=0.98
cc_213 VPB N_A_1501_92#_c_1207_n 0.0122039f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.99
cc_214 VPB N_A_1501_92#_c_1201_n 0.00244032f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.665
cc_215 VPB N_A_1501_92#_c_1209_n 0.010941f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_216 VPB N_A_1339_74#_c_1306_n 0.010501f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_217 VPB N_A_1339_74#_c_1307_n 0.00495563f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_218 VPB N_A_1339_74#_c_1320_n 0.0169614f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.145
cc_219 VPB N_A_1339_74#_c_1321_n 0.0171539f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.825
cc_220 VPB N_A_1339_74#_c_1322_n 0.0164743f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.665
cc_221 VPB N_A_1339_74#_c_1312_n 0.0151996f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_222 VPB N_A_1339_74#_c_1324_n 0.017828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_223 VPB N_A_1339_74#_c_1314_n 0.00851496f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_224 VPB N_A_1339_74#_c_1326_n 0.00170136f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_225 VPB N_A_1339_74#_c_1327_n 0.00744422f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_226 VPB N_A_1339_74#_c_1316_n 0.0323112f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_227 VPB N_A_1339_74#_c_1329_n 0.013245f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_228 VPB N_A_1339_74#_c_1330_n 0.00363179f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_229 VPB N_A_1339_74#_c_1331_n 0.00938777f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_230 VPB N_A_1339_74#_c_1332_n 0.00456694f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_231 VPB N_A_1339_74#_c_1333_n 0.00487964f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_232 VPB N_A_1339_74#_c_1317_n 0.00741432f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_233 VPB N_A_2221_74#_c_1506_n 0.016293f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.58
cc_234 VPB N_A_2221_74#_c_1507_n 0.017358f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_235 VPB N_A_2221_74#_c_1502_n 0.0146147f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_236 VPB N_A_2221_74#_c_1505_n 0.0168634f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_237 VPB N_A_27_74#_c_1571_n 0.0250181f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.145
cc_238 VPB N_A_27_74#_c_1576_n 0.0274899f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.825
cc_239 VPB N_A_27_74#_c_1577_n 0.0257471f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.99
cc_240 VPB N_A_27_74#_c_1578_n 0.0138378f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_241 VPB N_A_27_74#_c_1572_n 0.00269752f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.665
cc_242 VPB N_A_27_74#_c_1580_n 0.0109364f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.825
cc_243 VPB N_VPWR_c_1641_n 0.017335f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.825
cc_244 VPB N_VPWR_c_1642_n 0.00646119f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_245 VPB N_VPWR_c_1643_n 0.00579142f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_246 VPB N_VPWR_c_1644_n 0.00912606f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_247 VPB N_VPWR_c_1645_n 0.00811575f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_248 VPB N_VPWR_c_1646_n 0.0222249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_249 VPB N_VPWR_c_1647_n 0.0254075f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_250 VPB N_VPWR_c_1648_n 0.0157883f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_251 VPB N_VPWR_c_1649_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_252 VPB N_VPWR_c_1650_n 0.0644986f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_253 VPB N_VPWR_c_1651_n 0.0559624f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_254 VPB N_VPWR_c_1652_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_255 VPB N_VPWR_c_1653_n 0.0179825f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_256 VPB N_VPWR_c_1654_n 0.00487897f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_257 VPB N_VPWR_c_1655_n 0.0180274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_258 VPB N_VPWR_c_1656_n 0.0215753f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_259 VPB N_VPWR_c_1657_n 0.049432f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_260 VPB N_VPWR_c_1658_n 0.0312072f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_261 VPB N_VPWR_c_1659_n 0.0400196f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_262 VPB N_VPWR_c_1660_n 0.0219379f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_263 VPB N_VPWR_c_1661_n 0.0203698f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_264 VPB N_VPWR_c_1662_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_265 VPB N_VPWR_c_1663_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_266 VPB N_VPWR_c_1664_n 0.00436868f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_267 VPB N_VPWR_c_1665_n 0.00490136f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_268 VPB N_VPWR_c_1666_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_269 VPB N_VPWR_c_1667_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_270 VPB N_VPWR_c_1640_n 0.151502f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_271 VPB Q_N 0.00107477f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.58
cc_272 VPB Q_N 6.77734e-19 $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.75
cc_273 VPB Q_N 0.00238354f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_274 VPB N_Q_c_1824_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.465
cc_275 VPB N_Q_c_1825_n 0.00198321f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_276 VPB N_Q_c_1821_n 0.00104928f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_277 N_D_c_280_n N_CLK_c_313_n 0.00232413f $X=0.64 $Y=1.145 $X2=-0.19
+ $Y2=-0.245
cc_278 N_D_c_278_n N_CLK_c_314_n 0.00972409f $X=0.61 $Y=1.795 $X2=0 $Y2=0
cc_279 N_D_c_278_n N_A_225_74#_c_1017_n 0.00357638f $X=0.61 $Y=1.795 $X2=0 $Y2=0
cc_280 N_D_c_278_n N_A_225_74#_c_1036_n 0.00302188f $X=0.61 $Y=1.795 $X2=0 $Y2=0
cc_281 N_D_c_283_n N_A_225_74#_c_1036_n 9.40485e-19 $X=0.505 $Y=2.375 $X2=0
+ $Y2=0
cc_282 N_D_c_281_n N_A_225_74#_c_1036_n 0.0224944f $X=0.64 $Y=1.145 $X2=0 $Y2=0
cc_283 N_D_M1027_g N_A_225_74#_c_1019_n 0.00616966f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_284 N_D_c_280_n N_A_225_74#_c_1019_n 0.00357638f $X=0.64 $Y=1.145 $X2=0 $Y2=0
cc_285 N_D_c_281_n N_A_225_74#_c_1019_n 0.0556869f $X=0.64 $Y=1.145 $X2=0 $Y2=0
cc_286 N_D_M1027_g N_A_27_74#_c_1570_n 0.00146243f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_287 N_D_M1027_g N_A_27_74#_c_1571_n 0.00600966f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_288 N_D_c_280_n N_A_27_74#_c_1571_n 0.0320429f $X=0.64 $Y=1.145 $X2=0 $Y2=0
cc_289 N_D_c_281_n N_A_27_74#_c_1571_n 0.0697394f $X=0.64 $Y=1.145 $X2=0 $Y2=0
cc_290 N_D_c_283_n N_A_27_74#_c_1576_n 0.00433476f $X=0.505 $Y=2.375 $X2=0 $Y2=0
cc_291 N_D_c_284_n N_A_27_74#_c_1576_n 0.00528173f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_292 N_D_c_283_n N_A_27_74#_c_1577_n 0.0216554f $X=0.505 $Y=2.375 $X2=0 $Y2=0
cc_293 N_D_c_281_n N_A_27_74#_c_1577_n 0.0227191f $X=0.64 $Y=1.145 $X2=0 $Y2=0
cc_294 N_D_c_286_n N_A_27_74#_c_1577_n 0.00140505f $X=0.64 $Y=1.825 $X2=0 $Y2=0
cc_295 N_D_c_284_n N_VPWR_c_1641_n 0.0138303f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_296 N_D_c_284_n N_VPWR_c_1655_n 0.00413917f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_297 N_D_c_284_n N_VPWR_c_1640_n 0.00859049f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_298 N_D_M1027_g N_VGND_c_1853_n 0.0137856f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_299 N_D_c_280_n N_VGND_c_1853_n 0.00175174f $X=0.64 $Y=1.145 $X2=0 $Y2=0
cc_300 N_D_c_281_n N_VGND_c_1853_n 0.0220022f $X=0.64 $Y=1.145 $X2=0 $Y2=0
cc_301 N_D_M1027_g N_VGND_c_1864_n 0.00383152f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_302 N_D_M1027_g N_VGND_c_1878_n 0.00761198f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_303 N_CLK_c_313_n N_A_225_74#_M1015_g 0.0131368f $X=1.485 $Y=1.22 $X2=0 $Y2=0
cc_304 N_CLK_c_314_n N_A_225_74#_M1015_g 0.0210236f $X=1.515 $Y=1.715 $X2=0
+ $Y2=0
cc_305 CLK N_A_225_74#_M1015_g 0.00369616f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_306 N_CLK_c_314_n N_A_225_74#_c_1009_n 0.0477833f $X=1.515 $Y=1.715 $X2=0
+ $Y2=0
cc_307 N_CLK_c_313_n N_A_225_74#_c_1017_n 0.00330079f $X=1.485 $Y=1.22 $X2=0
+ $Y2=0
cc_308 N_CLK_c_314_n N_A_225_74#_c_1017_n 0.0065169f $X=1.515 $Y=1.715 $X2=0
+ $Y2=0
cc_309 CLK N_A_225_74#_c_1017_n 0.0286813f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_310 N_CLK_c_314_n N_A_225_74#_c_1035_n 0.00313913f $X=1.515 $Y=1.715 $X2=0
+ $Y2=0
cc_311 N_CLK_c_314_n N_A_225_74#_c_1037_n 0.00952984f $X=1.515 $Y=1.715 $X2=0
+ $Y2=0
cc_312 N_CLK_c_314_n N_A_225_74#_c_1018_n 0.00111203f $X=1.515 $Y=1.715 $X2=0
+ $Y2=0
cc_313 CLK N_A_225_74#_c_1018_n 0.0203335f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_314 N_CLK_c_313_n N_A_225_74#_c_1019_n 0.00765617f $X=1.485 $Y=1.22 $X2=0
+ $Y2=0
cc_315 N_CLK_c_314_n N_A_225_74#_c_1019_n 0.00114511f $X=1.515 $Y=1.715 $X2=0
+ $Y2=0
cc_316 CLK N_A_225_74#_c_1019_n 0.00762435f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_317 N_CLK_c_314_n N_A_225_74#_c_1039_n 0.00477306f $X=1.515 $Y=1.715 $X2=0
+ $Y2=0
cc_318 CLK N_A_225_74#_c_1039_n 0.0353587f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_319 N_CLK_c_314_n N_A_27_74#_c_1577_n 0.0161052f $X=1.515 $Y=1.715 $X2=0
+ $Y2=0
cc_320 CLK N_A_27_74#_c_1572_n 0.00324184f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_321 N_CLK_c_314_n N_VPWR_c_1641_n 0.0127906f $X=1.515 $Y=1.715 $X2=0 $Y2=0
cc_322 N_CLK_c_314_n N_VPWR_c_1642_n 0.0238569f $X=1.515 $Y=1.715 $X2=0 $Y2=0
cc_323 N_CLK_c_314_n N_VPWR_c_1656_n 0.0048608f $X=1.515 $Y=1.715 $X2=0 $Y2=0
cc_324 N_CLK_c_314_n N_VPWR_c_1640_n 0.00480464f $X=1.515 $Y=1.715 $X2=0 $Y2=0
cc_325 N_CLK_c_313_n N_VGND_c_1853_n 0.00299692f $X=1.485 $Y=1.22 $X2=0 $Y2=0
cc_326 N_CLK_c_313_n N_VGND_c_1854_n 0.00434272f $X=1.485 $Y=1.22 $X2=0 $Y2=0
cc_327 N_CLK_c_313_n N_VGND_c_1855_n 0.00300619f $X=1.485 $Y=1.22 $X2=0 $Y2=0
cc_328 CLK N_VGND_c_1855_n 0.0142803f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_329 N_CLK_c_313_n N_VGND_c_1878_n 0.00825157f $X=1.485 $Y=1.22 $X2=0 $Y2=0
cc_330 N_A_398_74#_c_353_n N_A_757_401#_c_626_n 0.00778145f $X=3.735 $Y=1.6
+ $X2=0 $Y2=0
cc_331 N_A_398_74#_c_374_n N_A_757_401#_c_626_n 0.00832316f $X=3.735 $Y=2.905
+ $X2=0 $Y2=0
cc_332 N_A_398_74#_c_386_p N_A_757_401#_c_626_n 0.00969066f $X=4.52 $Y=2.48
+ $X2=0 $Y2=0
cc_333 N_A_398_74#_c_375_n N_A_757_401#_c_626_n 0.00264629f $X=4.605 $Y=2.905
+ $X2=0 $Y2=0
cc_334 N_A_398_74#_c_388_p N_A_757_401#_c_626_n 0.00204235f $X=3.735 $Y=2.48
+ $X2=0 $Y2=0
cc_335 N_A_398_74#_M1034_g N_A_757_401#_c_621_n 0.0485648f $X=3.58 $Y=0.695
+ $X2=0 $Y2=0
cc_336 N_A_398_74#_c_386_p N_A_757_401#_c_627_n 0.00488545f $X=4.52 $Y=2.48
+ $X2=0 $Y2=0
cc_337 N_A_398_74#_M1034_g N_A_757_401#_c_622_n 0.00296636f $X=3.58 $Y=0.695
+ $X2=0 $Y2=0
cc_338 N_A_398_74#_c_354_n N_A_757_401#_c_623_n 0.00158807f $X=3.735 $Y=1.6
+ $X2=0 $Y2=0
cc_339 N_A_398_74#_c_365_n N_A_757_401#_c_628_n 0.00182462f $X=2.95 $Y=1.94
+ $X2=0 $Y2=0
cc_340 N_A_398_74#_c_353_n N_A_757_401#_c_628_n 0.00938262f $X=3.735 $Y=1.6
+ $X2=0 $Y2=0
cc_341 N_A_398_74#_c_354_n N_A_757_401#_c_628_n 0.00700413f $X=3.735 $Y=1.6
+ $X2=0 $Y2=0
cc_342 N_A_398_74#_c_386_p N_A_757_401#_c_629_n 0.0167319f $X=4.52 $Y=2.48 $X2=0
+ $Y2=0
cc_343 N_A_398_74#_c_353_n N_A_757_401#_c_630_n 0.0182267f $X=3.735 $Y=1.6 $X2=0
+ $Y2=0
cc_344 N_A_398_74#_c_386_p N_A_757_401#_c_630_n 0.0259281f $X=4.52 $Y=2.48 $X2=0
+ $Y2=0
cc_345 N_A_398_74#_c_353_n N_A_757_401#_c_631_n 0.00412226f $X=3.735 $Y=1.6
+ $X2=0 $Y2=0
cc_346 N_A_398_74#_c_386_p N_A_757_401#_c_631_n 0.00190513f $X=4.52 $Y=2.48
+ $X2=0 $Y2=0
cc_347 N_A_398_74#_M1034_g N_A_757_401#_c_624_n 3.1275e-19 $X=3.58 $Y=0.695
+ $X2=0 $Y2=0
cc_348 N_A_398_74#_c_376_n N_A_757_401#_c_632_n 0.0226037f $X=5.36 $Y=2.99 $X2=0
+ $Y2=0
cc_349 N_A_398_74#_c_380_n N_A_757_401#_c_632_n 0.00879771f $X=5.53 $Y=2.275
+ $X2=0 $Y2=0
cc_350 N_A_398_74#_c_353_n N_A_757_401#_c_625_n 0.00214471f $X=3.735 $Y=1.6
+ $X2=0 $Y2=0
cc_351 N_A_398_74#_c_354_n N_A_757_401#_c_625_n 0.00953288f $X=3.735 $Y=1.6
+ $X2=0 $Y2=0
cc_352 N_A_398_74#_c_359_n N_A_595_97#_M1014_d 0.00383506f $X=2.95 $Y=1.435
+ $X2=-0.19 $Y2=-0.245
cc_353 N_A_398_74#_c_375_n N_A_595_97#_c_732_n 0.00705669f $X=4.605 $Y=2.905
+ $X2=0 $Y2=0
cc_354 N_A_398_74#_c_376_n N_A_595_97#_c_732_n 0.00387126f $X=5.36 $Y=2.99 $X2=0
+ $Y2=0
cc_355 N_A_398_74#_c_378_n N_A_595_97#_c_732_n 5.12569e-19 $X=5.445 $Y=2.905
+ $X2=0 $Y2=0
cc_356 N_A_398_74#_c_356_n N_A_595_97#_c_715_n 0.00715673f $X=6.415 $Y=2.19
+ $X2=0 $Y2=0
cc_357 N_A_398_74#_c_378_n N_A_595_97#_c_734_n 0.00397946f $X=5.445 $Y=2.905
+ $X2=0 $Y2=0
cc_358 N_A_398_74#_c_379_n N_A_595_97#_c_734_n 0.0175786f $X=6.33 $Y=2.275 $X2=0
+ $Y2=0
cc_359 N_A_398_74#_c_356_n N_A_595_97#_c_734_n 0.00475761f $X=6.415 $Y=2.19
+ $X2=0 $Y2=0
cc_360 N_A_398_74#_c_355_n N_A_595_97#_c_716_n 0.00482959f $X=6.415 $Y=1.12
+ $X2=0 $Y2=0
cc_361 N_A_398_74#_c_358_n N_A_595_97#_c_716_n 0.00103022f $X=6.5 $Y=0.365 $X2=0
+ $Y2=0
cc_362 N_A_398_74#_c_363_n N_A_595_97#_c_716_n 0.0283274f $X=6.71 $Y=1.12 $X2=0
+ $Y2=0
cc_363 N_A_398_74#_c_360_n N_A_595_97#_c_717_n 0.00505169f $X=6.71 $Y=1.285
+ $X2=0 $Y2=0
cc_364 N_A_398_74#_c_361_n N_A_595_97#_c_717_n 0.0283274f $X=6.71 $Y=1.285 $X2=0
+ $Y2=0
cc_365 N_A_398_74#_M1034_g N_A_595_97#_c_718_n 0.00609952f $X=3.58 $Y=0.695
+ $X2=0 $Y2=0
cc_366 N_A_398_74#_c_359_n N_A_595_97#_c_718_n 0.0344769f $X=2.95 $Y=1.435 $X2=0
+ $Y2=0
cc_367 N_A_398_74#_M1034_g N_A_595_97#_c_719_n 0.00510302f $X=3.58 $Y=0.695
+ $X2=0 $Y2=0
cc_368 N_A_398_74#_c_359_n N_A_595_97#_c_719_n 0.0128205f $X=2.95 $Y=1.435 $X2=0
+ $Y2=0
cc_369 N_A_398_74#_c_365_n N_A_595_97#_c_720_n 0.0080703f $X=2.95 $Y=1.94 $X2=0
+ $Y2=0
cc_370 N_A_398_74#_c_366_n N_A_595_97#_c_720_n 5.4629e-19 $X=3.005 $Y=2.24 $X2=0
+ $Y2=0
cc_371 N_A_398_74#_c_347_n N_A_595_97#_c_720_n 0.0217142f $X=3.505 $Y=1.6 $X2=0
+ $Y2=0
cc_372 N_A_398_74#_M1034_g N_A_595_97#_c_720_n 0.00457084f $X=3.58 $Y=0.695
+ $X2=0 $Y2=0
cc_373 N_A_398_74#_c_352_n N_A_595_97#_c_720_n 0.0490068f $X=2.95 $Y=1.6 $X2=0
+ $Y2=0
cc_374 N_A_398_74#_c_353_n N_A_595_97#_c_720_n 0.0631092f $X=3.735 $Y=1.6 $X2=0
+ $Y2=0
cc_375 N_A_398_74#_c_359_n N_A_595_97#_c_720_n 0.0124678f $X=2.95 $Y=1.435 $X2=0
+ $Y2=0
cc_376 N_A_398_74#_M1034_g N_A_595_97#_c_721_n 0.0143046f $X=3.58 $Y=0.695 $X2=0
+ $Y2=0
cc_377 N_A_398_74#_c_353_n N_A_595_97#_c_721_n 0.0173132f $X=3.735 $Y=1.6 $X2=0
+ $Y2=0
cc_378 N_A_398_74#_c_354_n N_A_595_97#_c_721_n 0.00286357f $X=3.735 $Y=1.6 $X2=0
+ $Y2=0
cc_379 N_A_398_74#_M1034_g N_A_595_97#_c_722_n 0.0015524f $X=3.58 $Y=0.695 $X2=0
+ $Y2=0
cc_380 N_A_398_74#_c_353_n N_A_595_97#_c_722_n 0.00579354f $X=3.735 $Y=1.6 $X2=0
+ $Y2=0
cc_381 N_A_398_74#_c_354_n N_A_595_97#_c_722_n 7.68037e-19 $X=3.735 $Y=1.6 $X2=0
+ $Y2=0
cc_382 N_A_398_74#_c_353_n N_A_595_97#_c_724_n 0.0139492f $X=3.735 $Y=1.6 $X2=0
+ $Y2=0
cc_383 N_A_398_74#_c_354_n N_A_595_97#_c_724_n 0.00180184f $X=3.735 $Y=1.6 $X2=0
+ $Y2=0
cc_384 N_A_398_74#_c_365_n N_A_595_97#_c_738_n 6.08094e-19 $X=2.95 $Y=1.94 $X2=0
+ $Y2=0
cc_385 N_A_398_74#_c_366_n N_A_595_97#_c_738_n 0.00544933f $X=3.005 $Y=2.24
+ $X2=0 $Y2=0
cc_386 N_A_398_74#_c_347_n N_A_595_97#_c_738_n 0.00513144f $X=3.505 $Y=1.6 $X2=0
+ $Y2=0
cc_387 N_A_398_74#_c_369_n N_A_595_97#_c_738_n 0.0242908f $X=3.625 $Y=2.99 $X2=0
+ $Y2=0
cc_388 N_A_398_74#_c_352_n N_A_595_97#_c_738_n 0.00379884f $X=2.95 $Y=1.6 $X2=0
+ $Y2=0
cc_389 N_A_398_74#_c_353_n N_A_595_97#_c_738_n 0.00757356f $X=3.735 $Y=1.6 $X2=0
+ $Y2=0
cc_390 N_A_398_74#_c_374_n N_A_595_97#_c_738_n 0.0129106f $X=3.735 $Y=2.905
+ $X2=0 $Y2=0
cc_391 N_A_398_74#_c_388_p N_A_595_97#_c_738_n 0.0142749f $X=3.735 $Y=2.48 $X2=0
+ $Y2=0
cc_392 N_A_398_74#_M1034_g N_A_595_97#_c_781_n 0.00254046f $X=3.58 $Y=0.695
+ $X2=0 $Y2=0
cc_393 N_A_398_74#_c_347_n N_A_595_97#_c_725_n 0.00220182f $X=3.505 $Y=1.6 $X2=0
+ $Y2=0
cc_394 N_A_398_74#_M1034_g N_A_595_97#_c_725_n 0.00428676f $X=3.58 $Y=0.695
+ $X2=0 $Y2=0
cc_395 N_A_398_74#_c_359_n N_A_595_97#_c_725_n 0.0140647f $X=2.95 $Y=1.435 $X2=0
+ $Y2=0
cc_396 N_A_398_74#_c_360_n N_A_595_97#_c_728_n 0.0126088f $X=6.71 $Y=1.285 $X2=0
+ $Y2=0
cc_397 N_A_398_74#_c_376_n N_SET_B_c_898_n 0.00332799f $X=5.36 $Y=2.99 $X2=0
+ $Y2=0
cc_398 N_A_398_74#_c_378_n N_SET_B_c_898_n 0.0155453f $X=5.445 $Y=2.905 $X2=0
+ $Y2=0
cc_399 N_A_398_74#_c_380_n N_SET_B_c_898_n 0.00836468f $X=5.53 $Y=2.275 $X2=0
+ $Y2=0
cc_400 N_A_398_74#_c_362_n N_SET_B_c_885_n 0.00186884f $X=7.415 $Y=2.02 $X2=0
+ $Y2=0
cc_401 N_A_398_74#_c_368_n N_SET_B_c_891_n 5.88676e-19 $X=7.53 $Y=2.465 $X2=0
+ $Y2=0
cc_402 N_A_398_74#_c_379_n N_SET_B_c_891_n 0.0218509f $X=6.33 $Y=2.275 $X2=0
+ $Y2=0
cc_403 N_A_398_74#_c_356_n N_SET_B_c_891_n 0.0209674f $X=6.415 $Y=2.19 $X2=0
+ $Y2=0
cc_404 N_A_398_74#_c_360_n N_SET_B_c_891_n 0.0165581f $X=6.71 $Y=1.285 $X2=0
+ $Y2=0
cc_405 N_A_398_74#_c_361_n N_SET_B_c_891_n 0.00557641f $X=6.71 $Y=1.285 $X2=0
+ $Y2=0
cc_406 N_A_398_74#_c_382_n N_SET_B_c_891_n 0.00611943f $X=7.415 $Y=2.185 $X2=0
+ $Y2=0
cc_407 N_A_398_74#_c_362_n N_SET_B_c_891_n 0.0189131f $X=7.415 $Y=2.02 $X2=0
+ $Y2=0
cc_408 N_A_398_74#_c_379_n N_SET_B_c_892_n 0.00163184f $X=6.33 $Y=2.275 $X2=0
+ $Y2=0
cc_409 N_A_398_74#_c_380_n N_SET_B_c_892_n 7.6844e-19 $X=5.53 $Y=2.275 $X2=0
+ $Y2=0
cc_410 N_A_398_74#_c_379_n N_SET_B_c_893_n 0.00795886f $X=6.33 $Y=2.275 $X2=0
+ $Y2=0
cc_411 N_A_398_74#_c_380_n N_SET_B_c_893_n 0.0138178f $X=5.53 $Y=2.275 $X2=0
+ $Y2=0
cc_412 N_A_398_74#_c_349_n N_A_225_74#_M1015_g 0.00164183f $X=2.13 $Y=0.515
+ $X2=0 $Y2=0
cc_413 N_A_398_74#_c_351_n N_A_225_74#_M1015_g 0.00266901f $X=2.215 $Y=0.34
+ $X2=0 $Y2=0
cc_414 N_A_398_74#_c_468_p N_A_225_74#_c_1009_n 0.00431056f $X=2.19 $Y=2.665
+ $X2=0 $Y2=0
cc_415 N_A_398_74#_c_370_n N_A_225_74#_c_1009_n 0.00130182f $X=2.275 $Y=2.99
+ $X2=0 $Y2=0
cc_416 N_A_398_74#_c_365_n N_A_225_74#_c_1021_n 0.0237933f $X=2.95 $Y=1.94 $X2=0
+ $Y2=0
cc_417 N_A_398_74#_c_366_n N_A_225_74#_c_1021_n 0.0135716f $X=3.005 $Y=2.24
+ $X2=0 $Y2=0
cc_418 N_A_398_74#_c_468_p N_A_225_74#_c_1021_n 0.00613358f $X=2.19 $Y=2.665
+ $X2=0 $Y2=0
cc_419 N_A_398_74#_c_369_n N_A_225_74#_c_1021_n 0.0104889f $X=3.625 $Y=2.99
+ $X2=0 $Y2=0
cc_420 N_A_398_74#_c_352_n N_A_225_74#_c_1021_n 3.80029e-19 $X=2.95 $Y=1.6 $X2=0
+ $Y2=0
cc_421 N_A_398_74#_c_346_n N_A_225_74#_c_1010_n 0.0105031f $X=2.95 $Y=1.765
+ $X2=0 $Y2=0
cc_422 N_A_398_74#_c_350_n N_A_225_74#_c_1010_n 0.00132303f $X=2.94 $Y=0.34
+ $X2=0 $Y2=0
cc_423 N_A_398_74#_c_352_n N_A_225_74#_c_1010_n 0.00111273f $X=2.95 $Y=1.6 $X2=0
+ $Y2=0
cc_424 N_A_398_74#_c_359_n N_A_225_74#_c_1010_n 0.00549547f $X=2.95 $Y=1.435
+ $X2=0 $Y2=0
cc_425 N_A_398_74#_c_366_n N_A_225_74#_c_1022_n 0.00882199f $X=3.005 $Y=2.24
+ $X2=0 $Y2=0
cc_426 N_A_398_74#_c_369_n N_A_225_74#_c_1022_n 0.0121725f $X=3.625 $Y=2.99
+ $X2=0 $Y2=0
cc_427 N_A_398_74#_M1034_g N_A_225_74#_M1014_g 0.0110915f $X=3.58 $Y=0.695 $X2=0
+ $Y2=0
cc_428 N_A_398_74#_c_349_n N_A_225_74#_M1014_g 0.00397637f $X=2.13 $Y=0.515
+ $X2=0 $Y2=0
cc_429 N_A_398_74#_c_350_n N_A_225_74#_M1014_g 0.0109068f $X=2.94 $Y=0.34 $X2=0
+ $Y2=0
cc_430 N_A_398_74#_c_359_n N_A_225_74#_M1014_g 0.0197485f $X=2.95 $Y=1.435 $X2=0
+ $Y2=0
cc_431 N_A_398_74#_c_366_n N_A_225_74#_c_1024_n 0.00256863f $X=3.005 $Y=2.24
+ $X2=0 $Y2=0
cc_432 N_A_398_74#_c_374_n N_A_225_74#_c_1024_n 0.00287635f $X=3.735 $Y=2.905
+ $X2=0 $Y2=0
cc_433 N_A_398_74#_c_369_n N_A_225_74#_c_1025_n 0.0168575f $X=3.625 $Y=2.99
+ $X2=0 $Y2=0
cc_434 N_A_398_74#_c_365_n N_A_225_74#_c_1026_n 0.00221552f $X=2.95 $Y=1.94
+ $X2=0 $Y2=0
cc_435 N_A_398_74#_c_366_n N_A_225_74#_c_1026_n 0.00734034f $X=3.005 $Y=2.24
+ $X2=0 $Y2=0
cc_436 N_A_398_74#_c_347_n N_A_225_74#_c_1026_n 0.00516549f $X=3.505 $Y=1.6
+ $X2=0 $Y2=0
cc_437 N_A_398_74#_c_353_n N_A_225_74#_c_1026_n 0.00136066f $X=3.735 $Y=1.6
+ $X2=0 $Y2=0
cc_438 N_A_398_74#_c_374_n N_A_225_74#_c_1026_n 0.00288643f $X=3.735 $Y=2.905
+ $X2=0 $Y2=0
cc_439 N_A_398_74#_c_388_p N_A_225_74#_c_1026_n 0.00123961f $X=3.735 $Y=2.48
+ $X2=0 $Y2=0
cc_440 N_A_398_74#_c_368_n N_A_225_74#_c_1027_n 0.00130792f $X=7.53 $Y=2.465
+ $X2=0 $Y2=0
cc_441 N_A_398_74#_c_369_n N_A_225_74#_c_1027_n 0.00654236f $X=3.625 $Y=2.99
+ $X2=0 $Y2=0
cc_442 N_A_398_74#_c_386_p N_A_225_74#_c_1027_n 0.00661182f $X=4.52 $Y=2.48
+ $X2=0 $Y2=0
cc_443 N_A_398_74#_c_376_n N_A_225_74#_c_1027_n 0.0149209f $X=5.36 $Y=2.99 $X2=0
+ $Y2=0
cc_444 N_A_398_74#_c_377_n N_A_225_74#_c_1027_n 0.00419347f $X=4.69 $Y=2.99
+ $X2=0 $Y2=0
cc_445 N_A_398_74#_c_368_n N_A_225_74#_M1033_g 0.0023442f $X=7.53 $Y=2.465 $X2=0
+ $Y2=0
cc_446 N_A_398_74#_c_379_n N_A_225_74#_M1033_g 0.0015933f $X=6.33 $Y=2.275 $X2=0
+ $Y2=0
cc_447 N_A_398_74#_c_356_n N_A_225_74#_M1033_g 0.00241483f $X=6.415 $Y=2.19
+ $X2=0 $Y2=0
cc_448 N_A_398_74#_c_362_n N_A_225_74#_M1033_g 4.18952e-19 $X=7.415 $Y=2.02
+ $X2=0 $Y2=0
cc_449 N_A_398_74#_c_368_n N_A_225_74#_c_1012_n 0.00100919f $X=7.53 $Y=2.465
+ $X2=0 $Y2=0
cc_450 N_A_398_74#_c_356_n N_A_225_74#_c_1013_n 0.00195167f $X=6.415 $Y=2.19
+ $X2=0 $Y2=0
cc_451 N_A_398_74#_c_360_n N_A_225_74#_c_1013_n 0.00122013f $X=6.71 $Y=1.285
+ $X2=0 $Y2=0
cc_452 N_A_398_74#_c_361_n N_A_225_74#_c_1013_n 0.0172549f $X=6.71 $Y=1.285
+ $X2=0 $Y2=0
cc_453 N_A_398_74#_c_362_n N_A_225_74#_c_1013_n 2.64138e-19 $X=7.415 $Y=2.02
+ $X2=0 $Y2=0
cc_454 N_A_398_74#_c_356_n N_A_225_74#_M1035_g 9.168e-19 $X=6.415 $Y=2.19 $X2=0
+ $Y2=0
cc_455 N_A_398_74#_c_357_n N_A_225_74#_M1035_g 0.00565608f $X=7.385 $Y=0.365
+ $X2=0 $Y2=0
cc_456 N_A_398_74#_c_360_n N_A_225_74#_M1035_g 3.65769e-19 $X=6.71 $Y=1.285
+ $X2=0 $Y2=0
cc_457 N_A_398_74#_c_361_n N_A_225_74#_M1035_g 0.0180888f $X=6.71 $Y=1.285 $X2=0
+ $Y2=0
cc_458 N_A_398_74#_c_362_n N_A_225_74#_M1035_g 0.0107513f $X=7.415 $Y=2.02 $X2=0
+ $Y2=0
cc_459 N_A_398_74#_c_363_n N_A_225_74#_M1035_g 0.016767f $X=6.71 $Y=1.12 $X2=0
+ $Y2=0
cc_460 N_A_398_74#_c_346_n N_A_225_74#_c_1015_n 0.019666f $X=2.95 $Y=1.765 $X2=0
+ $Y2=0
cc_461 N_A_398_74#_c_349_n N_A_225_74#_c_1015_n 7.55533e-19 $X=2.13 $Y=0.515
+ $X2=0 $Y2=0
cc_462 N_A_398_74#_c_350_n N_A_225_74#_c_1015_n 9.27593e-19 $X=2.94 $Y=0.34
+ $X2=0 $Y2=0
cc_463 N_A_398_74#_c_352_n N_A_225_74#_c_1015_n 3.80029e-19 $X=2.95 $Y=1.6 $X2=0
+ $Y2=0
cc_464 N_A_398_74#_c_359_n N_A_225_74#_c_1015_n 8.1877e-19 $X=2.95 $Y=1.435
+ $X2=0 $Y2=0
cc_465 N_A_398_74#_c_349_n N_A_225_74#_c_1016_n 0.00106057f $X=2.13 $Y=0.515
+ $X2=0 $Y2=0
cc_466 N_A_398_74#_M1002_d N_A_225_74#_c_1037_n 0.00293855f $X=2.04 $Y=1.79
+ $X2=0 $Y2=0
cc_467 N_A_398_74#_c_349_n N_A_225_74#_c_1018_n 0.0147852f $X=2.13 $Y=0.515
+ $X2=0 $Y2=0
cc_468 N_A_398_74#_c_362_n N_A_1501_92#_M1019_g 0.0209879f $X=7.415 $Y=2.02
+ $X2=0 $Y2=0
cc_469 N_A_398_74#_c_368_n N_A_1501_92#_c_1203_n 0.023087f $X=7.53 $Y=2.465
+ $X2=0 $Y2=0
cc_470 N_A_398_74#_c_382_n N_A_1501_92#_c_1203_n 2.82185e-19 $X=7.415 $Y=2.185
+ $X2=0 $Y2=0
cc_471 N_A_398_74#_c_362_n N_A_1501_92#_c_1203_n 0.00523185f $X=7.415 $Y=2.02
+ $X2=0 $Y2=0
cc_472 N_A_398_74#_c_368_n N_A_1501_92#_c_1204_n 0.0281745f $X=7.53 $Y=2.465
+ $X2=0 $Y2=0
cc_473 N_A_398_74#_c_362_n N_A_1501_92#_c_1198_n 0.0563716f $X=7.415 $Y=2.02
+ $X2=0 $Y2=0
cc_474 N_A_398_74#_c_368_n N_A_1501_92#_c_1199_n 0.00341447f $X=7.53 $Y=2.465
+ $X2=0 $Y2=0
cc_475 N_A_398_74#_c_362_n N_A_1501_92#_c_1199_n 0.00557226f $X=7.415 $Y=2.02
+ $X2=0 $Y2=0
cc_476 N_A_398_74#_c_362_n N_A_1501_92#_c_1218_n 0.013418f $X=7.415 $Y=2.02
+ $X2=0 $Y2=0
cc_477 N_A_398_74#_c_357_n N_A_1339_74#_M1018_d 0.00226519f $X=7.385 $Y=0.365
+ $X2=-0.19 $Y2=-0.245
cc_478 N_A_398_74#_c_357_n N_A_1339_74#_c_1336_n 0.0335956f $X=7.385 $Y=0.365
+ $X2=0 $Y2=0
cc_479 N_A_398_74#_c_360_n N_A_1339_74#_c_1336_n 0.0135629f $X=6.71 $Y=1.285
+ $X2=0 $Y2=0
cc_480 N_A_398_74#_c_361_n N_A_1339_74#_c_1336_n 0.00395514f $X=6.71 $Y=1.285
+ $X2=0 $Y2=0
cc_481 N_A_398_74#_c_362_n N_A_1339_74#_c_1336_n 0.02548f $X=7.415 $Y=2.02 $X2=0
+ $Y2=0
cc_482 N_A_398_74#_c_363_n N_A_1339_74#_c_1336_n 0.00921999f $X=6.71 $Y=1.12
+ $X2=0 $Y2=0
cc_483 N_A_398_74#_c_368_n N_A_1339_74#_c_1326_n 0.00589256f $X=7.53 $Y=2.465
+ $X2=0 $Y2=0
cc_484 N_A_398_74#_c_379_n N_A_1339_74#_c_1326_n 0.00938866f $X=6.33 $Y=2.275
+ $X2=0 $Y2=0
cc_485 N_A_398_74#_c_356_n N_A_1339_74#_c_1326_n 0.0167066f $X=6.415 $Y=2.19
+ $X2=0 $Y2=0
cc_486 N_A_398_74#_c_382_n N_A_1339_74#_c_1326_n 0.0180759f $X=7.415 $Y=2.185
+ $X2=0 $Y2=0
cc_487 N_A_398_74#_c_362_n N_A_1339_74#_c_1326_n 0.00780717f $X=7.415 $Y=2.02
+ $X2=0 $Y2=0
cc_488 N_A_398_74#_c_355_n N_A_1339_74#_c_1315_n 0.00454611f $X=6.415 $Y=1.12
+ $X2=0 $Y2=0
cc_489 N_A_398_74#_c_356_n N_A_1339_74#_c_1315_n 0.0064862f $X=6.415 $Y=2.19
+ $X2=0 $Y2=0
cc_490 N_A_398_74#_c_360_n N_A_1339_74#_c_1315_n 0.0257548f $X=6.71 $Y=1.285
+ $X2=0 $Y2=0
cc_491 N_A_398_74#_c_361_n N_A_1339_74#_c_1315_n 9.90303e-19 $X=6.71 $Y=1.285
+ $X2=0 $Y2=0
cc_492 N_A_398_74#_c_362_n N_A_1339_74#_c_1315_n 0.0517761f $X=7.415 $Y=2.02
+ $X2=0 $Y2=0
cc_493 N_A_398_74#_c_363_n N_A_1339_74#_c_1315_n 0.00131891f $X=6.71 $Y=1.12
+ $X2=0 $Y2=0
cc_494 N_A_398_74#_c_356_n N_A_1339_74#_c_1330_n 0.00802298f $X=6.415 $Y=2.19
+ $X2=0 $Y2=0
cc_495 N_A_398_74#_c_360_n N_A_1339_74#_c_1330_n 0.00416021f $X=6.71 $Y=1.285
+ $X2=0 $Y2=0
cc_496 N_A_398_74#_c_361_n N_A_1339_74#_c_1330_n 3.84168e-19 $X=6.71 $Y=1.285
+ $X2=0 $Y2=0
cc_497 N_A_398_74#_c_362_n N_A_1339_74#_c_1330_n 0.012655f $X=7.415 $Y=2.02
+ $X2=0 $Y2=0
cc_498 N_A_398_74#_c_368_n N_A_1339_74#_c_1331_n 0.0147927f $X=7.53 $Y=2.465
+ $X2=0 $Y2=0
cc_499 N_A_398_74#_c_382_n N_A_1339_74#_c_1331_n 0.0263641f $X=7.415 $Y=2.185
+ $X2=0 $Y2=0
cc_500 N_A_398_74#_c_368_n N_A_1339_74#_c_1332_n 0.0103428f $X=7.53 $Y=2.465
+ $X2=0 $Y2=0
cc_501 N_A_398_74#_c_368_n N_A_1339_74#_c_1333_n 0.00695105f $X=7.53 $Y=2.465
+ $X2=0 $Y2=0
cc_502 N_A_398_74#_c_382_n N_A_1339_74#_c_1333_n 0.0244552f $X=7.415 $Y=2.185
+ $X2=0 $Y2=0
cc_503 N_A_398_74#_c_362_n N_A_1339_74#_c_1333_n 0.00525436f $X=7.415 $Y=2.02
+ $X2=0 $Y2=0
cc_504 N_A_398_74#_M1002_d N_A_27_74#_c_1578_n 0.00599509f $X=2.04 $Y=1.79 $X2=0
+ $Y2=0
cc_505 N_A_398_74#_c_365_n N_A_27_74#_c_1578_n 0.00236432f $X=2.95 $Y=1.94 $X2=0
+ $Y2=0
cc_506 N_A_398_74#_c_366_n N_A_27_74#_c_1578_n 0.00248169f $X=3.005 $Y=2.24
+ $X2=0 $Y2=0
cc_507 N_A_398_74#_c_468_p N_A_27_74#_c_1578_n 0.0389929f $X=2.19 $Y=2.665 $X2=0
+ $Y2=0
cc_508 N_A_398_74#_c_369_n N_A_27_74#_c_1578_n 0.0356935f $X=3.625 $Y=2.99 $X2=0
+ $Y2=0
cc_509 N_A_398_74#_c_352_n N_A_27_74#_c_1578_n 0.0100447f $X=2.95 $Y=1.6 $X2=0
+ $Y2=0
cc_510 N_A_398_74#_c_346_n N_A_27_74#_c_1572_n 0.00362357f $X=2.95 $Y=1.765
+ $X2=0 $Y2=0
cc_511 N_A_398_74#_c_349_n N_A_27_74#_c_1572_n 0.0119039f $X=2.13 $Y=0.515 $X2=0
+ $Y2=0
cc_512 N_A_398_74#_c_352_n N_A_27_74#_c_1572_n 0.0468227f $X=2.95 $Y=1.6 $X2=0
+ $Y2=0
cc_513 N_A_398_74#_c_359_n N_A_27_74#_c_1572_n 0.0228448f $X=2.95 $Y=1.435 $X2=0
+ $Y2=0
cc_514 N_A_398_74#_c_349_n N_A_27_74#_c_1574_n 0.0206338f $X=2.13 $Y=0.515 $X2=0
+ $Y2=0
cc_515 N_A_398_74#_c_350_n N_A_27_74#_c_1574_n 0.0237903f $X=2.94 $Y=0.34 $X2=0
+ $Y2=0
cc_516 N_A_398_74#_c_359_n N_A_27_74#_c_1574_n 0.0119198f $X=2.95 $Y=1.435 $X2=0
+ $Y2=0
cc_517 N_A_398_74#_c_386_p N_VPWR_M1004_d 0.0160077f $X=4.52 $Y=2.48 $X2=0 $Y2=0
cc_518 N_A_398_74#_c_375_n N_VPWR_M1004_d 0.00424497f $X=4.605 $Y=2.905 $X2=0
+ $Y2=0
cc_519 N_A_398_74#_c_378_n N_VPWR_M1036_d 0.00485888f $X=5.445 $Y=2.905 $X2=0
+ $Y2=0
cc_520 N_A_398_74#_c_379_n N_VPWR_M1036_d 0.0160983f $X=6.33 $Y=2.275 $X2=0
+ $Y2=0
cc_521 N_A_398_74#_c_468_p N_VPWR_c_1642_n 0.0243941f $X=2.19 $Y=2.665 $X2=0
+ $Y2=0
cc_522 N_A_398_74#_c_370_n N_VPWR_c_1642_n 0.0128267f $X=2.275 $Y=2.99 $X2=0
+ $Y2=0
cc_523 N_A_398_74#_c_369_n N_VPWR_c_1643_n 0.0147319f $X=3.625 $Y=2.99 $X2=0
+ $Y2=0
cc_524 N_A_398_74#_c_374_n N_VPWR_c_1643_n 0.0129054f $X=3.735 $Y=2.905 $X2=0
+ $Y2=0
cc_525 N_A_398_74#_c_386_p N_VPWR_c_1643_n 0.0259107f $X=4.52 $Y=2.48 $X2=0
+ $Y2=0
cc_526 N_A_398_74#_c_375_n N_VPWR_c_1643_n 0.0134405f $X=4.605 $Y=2.905 $X2=0
+ $Y2=0
cc_527 N_A_398_74#_c_377_n N_VPWR_c_1643_n 0.0150385f $X=4.69 $Y=2.99 $X2=0
+ $Y2=0
cc_528 N_A_398_74#_c_376_n N_VPWR_c_1644_n 0.0151625f $X=5.36 $Y=2.99 $X2=0
+ $Y2=0
cc_529 N_A_398_74#_c_378_n N_VPWR_c_1644_n 0.0293715f $X=5.445 $Y=2.905 $X2=0
+ $Y2=0
cc_530 N_A_398_74#_c_379_n N_VPWR_c_1644_n 0.0299399f $X=6.33 $Y=2.275 $X2=0
+ $Y2=0
cc_531 N_A_398_74#_c_368_n N_VPWR_c_1651_n 0.0032704f $X=7.53 $Y=2.465 $X2=0
+ $Y2=0
cc_532 N_A_398_74#_c_369_n N_VPWR_c_1657_n 0.100928f $X=3.625 $Y=2.99 $X2=0
+ $Y2=0
cc_533 N_A_398_74#_c_370_n N_VPWR_c_1657_n 0.01218f $X=2.275 $Y=2.99 $X2=0 $Y2=0
cc_534 N_A_398_74#_c_376_n N_VPWR_c_1658_n 0.0546768f $X=5.36 $Y=2.99 $X2=0
+ $Y2=0
cc_535 N_A_398_74#_c_377_n N_VPWR_c_1658_n 0.0115893f $X=4.69 $Y=2.99 $X2=0
+ $Y2=0
cc_536 N_A_398_74#_c_368_n N_VPWR_c_1640_n 0.00420718f $X=7.53 $Y=2.465 $X2=0
+ $Y2=0
cc_537 N_A_398_74#_c_369_n N_VPWR_c_1640_n 0.0531785f $X=3.625 $Y=2.99 $X2=0
+ $Y2=0
cc_538 N_A_398_74#_c_370_n N_VPWR_c_1640_n 0.00660793f $X=2.275 $Y=2.99 $X2=0
+ $Y2=0
cc_539 N_A_398_74#_c_386_p N_VPWR_c_1640_n 0.0122674f $X=4.52 $Y=2.48 $X2=0
+ $Y2=0
cc_540 N_A_398_74#_c_376_n N_VPWR_c_1640_n 0.028344f $X=5.36 $Y=2.99 $X2=0 $Y2=0
cc_541 N_A_398_74#_c_377_n N_VPWR_c_1640_n 0.00583135f $X=4.69 $Y=2.99 $X2=0
+ $Y2=0
cc_542 N_A_398_74#_c_353_n A_706_463# 6.51072e-19 $X=3.735 $Y=1.6 $X2=-0.19
+ $Y2=-0.245
cc_543 N_A_398_74#_c_374_n A_706_463# 0.00138456f $X=3.735 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_544 N_A_398_74#_c_388_p A_706_463# 0.00144701f $X=3.735 $Y=2.48 $X2=-0.19
+ $Y2=-0.245
cc_545 N_A_398_74#_c_379_n A_1258_341# 0.00893904f $X=6.33 $Y=2.275 $X2=-0.19
+ $Y2=-0.245
cc_546 N_A_398_74#_c_356_n A_1258_341# 0.00767253f $X=6.415 $Y=2.19 $X2=-0.19
+ $Y2=-0.245
cc_547 N_A_398_74#_c_351_n N_VGND_c_1855_n 0.0110038f $X=2.215 $Y=0.34 $X2=0
+ $Y2=0
cc_548 N_A_398_74#_M1034_g N_VGND_c_1856_n 0.00159069f $X=3.58 $Y=0.695 $X2=0
+ $Y2=0
cc_549 N_A_398_74#_M1034_g N_VGND_c_1865_n 0.00476381f $X=3.58 $Y=0.695 $X2=0
+ $Y2=0
cc_550 N_A_398_74#_c_350_n N_VGND_c_1865_n 0.0588317f $X=2.94 $Y=0.34 $X2=0
+ $Y2=0
cc_551 N_A_398_74#_c_351_n N_VGND_c_1865_n 0.0121867f $X=2.215 $Y=0.34 $X2=0
+ $Y2=0
cc_552 N_A_398_74#_c_358_n N_VGND_c_1873_n 0.0113619f $X=6.5 $Y=0.365 $X2=0
+ $Y2=0
cc_553 N_A_398_74#_c_363_n N_VGND_c_1873_n 3.97182e-19 $X=6.71 $Y=1.12 $X2=0
+ $Y2=0
cc_554 N_A_398_74#_c_357_n N_VGND_c_1874_n 0.0593621f $X=7.385 $Y=0.365 $X2=0
+ $Y2=0
cc_555 N_A_398_74#_c_358_n N_VGND_c_1874_n 0.0105206f $X=6.5 $Y=0.365 $X2=0
+ $Y2=0
cc_556 N_A_398_74#_c_363_n N_VGND_c_1874_n 0.00281891f $X=6.71 $Y=1.12 $X2=0
+ $Y2=0
cc_557 N_A_398_74#_c_357_n N_VGND_c_1875_n 0.0070631f $X=7.385 $Y=0.365 $X2=0
+ $Y2=0
cc_558 N_A_398_74#_c_362_n N_VGND_c_1875_n 0.00572644f $X=7.415 $Y=2.02 $X2=0
+ $Y2=0
cc_559 N_A_398_74#_M1034_g N_VGND_c_1878_n 0.00509887f $X=3.58 $Y=0.695 $X2=0
+ $Y2=0
cc_560 N_A_398_74#_c_350_n N_VGND_c_1878_n 0.0338596f $X=2.94 $Y=0.34 $X2=0
+ $Y2=0
cc_561 N_A_398_74#_c_351_n N_VGND_c_1878_n 0.00660921f $X=2.215 $Y=0.34 $X2=0
+ $Y2=0
cc_562 N_A_398_74#_c_357_n N_VGND_c_1878_n 0.0385992f $X=7.385 $Y=0.365 $X2=0
+ $Y2=0
cc_563 N_A_398_74#_c_358_n N_VGND_c_1878_n 0.00652894f $X=6.5 $Y=0.365 $X2=0
+ $Y2=0
cc_564 N_A_398_74#_c_363_n N_VGND_c_1878_n 0.00358754f $X=6.71 $Y=1.12 $X2=0
+ $Y2=0
cc_565 N_A_398_74#_c_355_n A_1261_74# 0.00221695f $X=6.415 $Y=1.12 $X2=-0.19
+ $Y2=-0.245
cc_566 N_A_398_74#_c_362_n A_1453_118# 0.00353049f $X=7.415 $Y=2.02 $X2=-0.19
+ $Y2=-0.245
cc_567 N_A_757_401#_c_629_n N_A_595_97#_c_731_n 0.00456609f $X=4.86 $Y=2.14
+ $X2=0 $Y2=0
cc_568 N_A_757_401#_c_630_n N_A_595_97#_c_731_n 0.00118759f $X=4.305 $Y=1.99
+ $X2=0 $Y2=0
cc_569 N_A_757_401#_c_631_n N_A_595_97#_c_731_n 0.0152588f $X=4.305 $Y=1.99
+ $X2=0 $Y2=0
cc_570 N_A_757_401#_c_632_n N_A_595_97#_c_731_n 0.00148749f $X=5.025 $Y=2.14
+ $X2=0 $Y2=0
cc_571 N_A_757_401#_c_629_n N_A_595_97#_c_732_n 0.00868233f $X=4.86 $Y=2.14
+ $X2=0 $Y2=0
cc_572 N_A_757_401#_c_630_n N_A_595_97#_c_732_n 2.77028e-19 $X=4.305 $Y=1.99
+ $X2=0 $Y2=0
cc_573 N_A_757_401#_c_632_n N_A_595_97#_c_732_n 0.012978f $X=5.025 $Y=2.14 $X2=0
+ $Y2=0
cc_574 N_A_757_401#_c_622_n N_A_595_97#_M1026_g 0.0201634f $X=4.295 $Y=1.09
+ $X2=0 $Y2=0
cc_575 N_A_757_401#_c_624_n N_A_595_97#_M1026_g 0.0194663f $X=4.715 $Y=0.58
+ $X2=0 $Y2=0
cc_576 N_A_757_401#_c_625_n N_A_595_97#_M1026_g 0.00519936f $X=4.305 $Y=1.825
+ $X2=0 $Y2=0
cc_577 N_A_757_401#_c_621_n N_A_595_97#_c_718_n 0.00117593f $X=3.94 $Y=1.015
+ $X2=0 $Y2=0
cc_578 N_A_757_401#_c_628_n N_A_595_97#_c_720_n 5.46737e-19 $X=3.875 $Y=2.08
+ $X2=0 $Y2=0
cc_579 N_A_757_401#_c_622_n N_A_595_97#_c_721_n 0.00856275f $X=4.295 $Y=1.09
+ $X2=0 $Y2=0
cc_580 N_A_757_401#_c_623_n N_A_595_97#_c_721_n 0.00961364f $X=4.015 $Y=1.09
+ $X2=0 $Y2=0
cc_581 N_A_757_401#_c_624_n N_A_595_97#_c_721_n 0.0137257f $X=4.715 $Y=0.58
+ $X2=0 $Y2=0
cc_582 N_A_757_401#_c_622_n N_A_595_97#_c_722_n 0.00316276f $X=4.295 $Y=1.09
+ $X2=0 $Y2=0
cc_583 N_A_757_401#_c_624_n N_A_595_97#_c_722_n 0.005833f $X=4.715 $Y=0.58 $X2=0
+ $Y2=0
cc_584 N_A_757_401#_c_622_n N_A_595_97#_c_723_n 0.00378094f $X=4.295 $Y=1.09
+ $X2=0 $Y2=0
cc_585 N_A_757_401#_c_629_n N_A_595_97#_c_723_n 0.0119117f $X=4.86 $Y=2.14 $X2=0
+ $Y2=0
cc_586 N_A_757_401#_c_630_n N_A_595_97#_c_723_n 0.0210386f $X=4.305 $Y=1.99
+ $X2=0 $Y2=0
cc_587 N_A_757_401#_c_631_n N_A_595_97#_c_723_n 0.00144642f $X=4.305 $Y=1.99
+ $X2=0 $Y2=0
cc_588 N_A_757_401#_c_624_n N_A_595_97#_c_723_n 0.0239403f $X=4.715 $Y=0.58
+ $X2=0 $Y2=0
cc_589 N_A_757_401#_c_625_n N_A_595_97#_c_723_n 0.0120775f $X=4.305 $Y=1.825
+ $X2=0 $Y2=0
cc_590 N_A_757_401#_c_627_n N_A_595_97#_c_724_n 0.00424988f $X=4.14 $Y=2.08
+ $X2=0 $Y2=0
cc_591 N_A_757_401#_c_630_n N_A_595_97#_c_724_n 0.0037144f $X=4.305 $Y=1.99
+ $X2=0 $Y2=0
cc_592 N_A_757_401#_c_631_n N_A_595_97#_c_724_n 5.49386e-19 $X=4.305 $Y=1.99
+ $X2=0 $Y2=0
cc_593 N_A_757_401#_c_626_n N_A_595_97#_c_738_n 3.77018e-19 $X=3.875 $Y=2.24
+ $X2=0 $Y2=0
cc_594 N_A_757_401#_c_623_n N_A_595_97#_c_781_n 0.00117593f $X=4.015 $Y=1.09
+ $X2=0 $Y2=0
cc_595 N_A_757_401#_c_622_n N_A_595_97#_c_726_n 6.62687e-19 $X=4.295 $Y=1.09
+ $X2=0 $Y2=0
cc_596 N_A_757_401#_c_629_n N_A_595_97#_c_726_n 0.00823228f $X=4.86 $Y=2.14
+ $X2=0 $Y2=0
cc_597 N_A_757_401#_c_630_n N_A_595_97#_c_726_n 0.00148595f $X=4.305 $Y=1.99
+ $X2=0 $Y2=0
cc_598 N_A_757_401#_c_631_n N_A_595_97#_c_726_n 2.79593e-19 $X=4.305 $Y=1.99
+ $X2=0 $Y2=0
cc_599 N_A_757_401#_c_624_n N_A_595_97#_c_726_n 0.017608f $X=4.715 $Y=0.58 $X2=0
+ $Y2=0
cc_600 N_A_757_401#_c_632_n N_A_595_97#_c_726_n 0.0135425f $X=5.025 $Y=2.14
+ $X2=0 $Y2=0
cc_601 N_A_757_401#_c_625_n N_A_595_97#_c_726_n 0.00244526f $X=4.305 $Y=1.825
+ $X2=0 $Y2=0
cc_602 N_A_757_401#_c_629_n N_A_595_97#_c_727_n 6.15625e-19 $X=4.86 $Y=2.14
+ $X2=0 $Y2=0
cc_603 N_A_757_401#_c_631_n N_A_595_97#_c_727_n 0.00379936f $X=4.305 $Y=1.99
+ $X2=0 $Y2=0
cc_604 N_A_757_401#_c_624_n N_A_595_97#_c_727_n 8.22839e-19 $X=4.715 $Y=0.58
+ $X2=0 $Y2=0
cc_605 N_A_757_401#_c_632_n N_A_595_97#_c_727_n 9.65695e-19 $X=5.025 $Y=2.14
+ $X2=0 $Y2=0
cc_606 N_A_757_401#_c_625_n N_A_595_97#_c_727_n 0.0150128f $X=4.305 $Y=1.825
+ $X2=0 $Y2=0
cc_607 N_A_757_401#_c_632_n N_A_595_97#_c_729_n 4.98461e-19 $X=5.025 $Y=2.14
+ $X2=0 $Y2=0
cc_608 N_A_757_401#_c_632_n N_SET_B_c_898_n 0.00678902f $X=5.025 $Y=2.14 $X2=0
+ $Y2=0
cc_609 N_A_757_401#_c_624_n N_SET_B_c_889_n 0.00257545f $X=4.715 $Y=0.58 $X2=0
+ $Y2=0
cc_610 N_A_757_401#_c_626_n N_A_225_74#_c_1024_n 0.0025248f $X=3.875 $Y=2.24
+ $X2=0 $Y2=0
cc_611 N_A_757_401#_c_626_n N_A_225_74#_c_1026_n 0.0239602f $X=3.875 $Y=2.24
+ $X2=0 $Y2=0
cc_612 N_A_757_401#_c_628_n N_A_225_74#_c_1026_n 0.00250032f $X=3.875 $Y=2.08
+ $X2=0 $Y2=0
cc_613 N_A_757_401#_c_626_n N_A_225_74#_c_1027_n 0.00989848f $X=3.875 $Y=2.24
+ $X2=0 $Y2=0
cc_614 N_A_757_401#_c_626_n N_VPWR_c_1643_n 0.00286806f $X=3.875 $Y=2.24 $X2=0
+ $Y2=0
cc_615 N_A_757_401#_c_626_n N_VPWR_c_1640_n 6.59927e-19 $X=3.875 $Y=2.24 $X2=0
+ $Y2=0
cc_616 N_A_757_401#_c_621_n N_VGND_c_1856_n 0.0112772f $X=3.94 $Y=1.015 $X2=0
+ $Y2=0
cc_617 N_A_757_401#_c_622_n N_VGND_c_1856_n 0.00479662f $X=4.295 $Y=1.09 $X2=0
+ $Y2=0
cc_618 N_A_757_401#_c_624_n N_VGND_c_1856_n 0.0411686f $X=4.715 $Y=0.58 $X2=0
+ $Y2=0
cc_619 N_A_757_401#_c_621_n N_VGND_c_1865_n 0.00413255f $X=3.94 $Y=1.015 $X2=0
+ $Y2=0
cc_620 N_A_757_401#_c_624_n N_VGND_c_1872_n 0.0208755f $X=4.715 $Y=0.58 $X2=0
+ $Y2=0
cc_621 N_A_757_401#_c_624_n N_VGND_c_1873_n 0.0120077f $X=4.715 $Y=0.58 $X2=0
+ $Y2=0
cc_622 N_A_757_401#_c_621_n N_VGND_c_1878_n 0.00428305f $X=3.94 $Y=1.015 $X2=0
+ $Y2=0
cc_623 N_A_757_401#_c_624_n N_VGND_c_1878_n 0.0172297f $X=4.715 $Y=0.58 $X2=0
+ $Y2=0
cc_624 N_A_595_97#_M1026_g N_SET_B_c_884_n 0.0317616f $X=4.93 $Y=0.58 $X2=0
+ $Y2=0
cc_625 N_A_595_97#_c_726_n N_SET_B_c_884_n 0.00434007f $X=4.882 $Y=1.325 $X2=0
+ $Y2=0
cc_626 N_A_595_97#_c_727_n N_SET_B_c_884_n 0.0197563f $X=4.85 $Y=1.72 $X2=0
+ $Y2=0
cc_627 N_A_595_97#_c_728_n N_SET_B_c_884_n 7.95332e-19 $X=5.75 $Y=1.285 $X2=0
+ $Y2=0
cc_628 N_A_595_97#_c_729_n N_SET_B_c_884_n 0.0131004f $X=5.585 $Y=1.265 $X2=0
+ $Y2=0
cc_629 N_A_595_97#_c_730_n N_SET_B_c_884_n 0.0208717f $X=5.75 $Y=1.195 $X2=0
+ $Y2=0
cc_630 N_A_595_97#_c_731_n N_SET_B_c_898_n 0.0129088f $X=4.8 $Y=2.15 $X2=0 $Y2=0
cc_631 N_A_595_97#_c_732_n N_SET_B_c_898_n 0.0114098f $X=4.8 $Y=2.24 $X2=0 $Y2=0
cc_632 N_A_595_97#_c_734_n N_SET_B_c_898_n 0.0049383f $X=6.215 $Y=1.63 $X2=0
+ $Y2=0
cc_633 N_A_595_97#_c_729_n N_SET_B_c_898_n 9.56033e-19 $X=5.585 $Y=1.265 $X2=0
+ $Y2=0
cc_634 N_A_595_97#_M1026_g N_SET_B_c_889_n 0.0460006f $X=4.93 $Y=0.58 $X2=0
+ $Y2=0
cc_635 N_A_595_97#_c_729_n N_SET_B_c_890_n 3.91223e-19 $X=5.585 $Y=1.265 $X2=0
+ $Y2=0
cc_636 N_A_595_97#_c_714_n N_SET_B_c_891_n 0.0040413f $X=6.125 $Y=1.195 $X2=0
+ $Y2=0
cc_637 N_A_595_97#_c_734_n N_SET_B_c_891_n 0.0136427f $X=6.215 $Y=1.63 $X2=0
+ $Y2=0
cc_638 N_A_595_97#_c_728_n N_SET_B_c_891_n 0.010821f $X=5.75 $Y=1.285 $X2=0
+ $Y2=0
cc_639 N_A_595_97#_c_730_n N_SET_B_c_891_n 0.00611328f $X=5.75 $Y=1.195 $X2=0
+ $Y2=0
cc_640 N_A_595_97#_c_734_n N_SET_B_c_892_n 0.00154203f $X=6.215 $Y=1.63 $X2=0
+ $Y2=0
cc_641 N_A_595_97#_c_726_n N_SET_B_c_892_n 0.00204547f $X=4.882 $Y=1.325 $X2=0
+ $Y2=0
cc_642 N_A_595_97#_c_729_n N_SET_B_c_892_n 0.00882985f $X=5.585 $Y=1.265 $X2=0
+ $Y2=0
cc_643 N_A_595_97#_c_730_n N_SET_B_c_892_n 0.00215733f $X=5.75 $Y=1.195 $X2=0
+ $Y2=0
cc_644 N_A_595_97#_c_731_n N_SET_B_c_893_n 8.23032e-19 $X=4.8 $Y=2.15 $X2=0
+ $Y2=0
cc_645 N_A_595_97#_c_734_n N_SET_B_c_893_n 0.00727859f $X=6.215 $Y=1.63 $X2=0
+ $Y2=0
cc_646 N_A_595_97#_c_726_n N_SET_B_c_893_n 0.0182485f $X=4.882 $Y=1.325 $X2=0
+ $Y2=0
cc_647 N_A_595_97#_c_727_n N_SET_B_c_893_n 0.0010606f $X=4.85 $Y=1.72 $X2=0
+ $Y2=0
cc_648 N_A_595_97#_c_729_n N_SET_B_c_893_n 0.0282062f $X=5.585 $Y=1.265 $X2=0
+ $Y2=0
cc_649 N_A_595_97#_c_730_n N_SET_B_c_893_n 0.00114191f $X=5.75 $Y=1.195 $X2=0
+ $Y2=0
cc_650 N_A_595_97#_c_738_n N_A_225_74#_c_1021_n 3.09534e-19 $X=3.37 $Y=2.515
+ $X2=0 $Y2=0
cc_651 N_A_595_97#_c_725_n N_A_225_74#_c_1010_n 3.39751e-19 $X=3.407 $Y=1.18
+ $X2=0 $Y2=0
cc_652 N_A_595_97#_c_718_n N_A_225_74#_M1014_g 0.001333f $X=3.365 $Y=0.695 $X2=0
+ $Y2=0
cc_653 N_A_595_97#_c_719_n N_A_225_74#_M1014_g 4.88269e-19 $X=3.407 $Y=1.095
+ $X2=0 $Y2=0
cc_654 N_A_595_97#_c_720_n N_A_225_74#_c_1026_n 0.0036049f $X=3.37 $Y=2.295
+ $X2=0 $Y2=0
cc_655 N_A_595_97#_c_738_n N_A_225_74#_c_1026_n 0.00777105f $X=3.37 $Y=2.515
+ $X2=0 $Y2=0
cc_656 N_A_595_97#_c_732_n N_A_225_74#_c_1027_n 0.00882199f $X=4.8 $Y=2.24 $X2=0
+ $Y2=0
cc_657 N_A_595_97#_c_734_n N_A_225_74#_c_1027_n 0.00907339f $X=6.215 $Y=1.63
+ $X2=0 $Y2=0
cc_658 N_A_595_97#_c_734_n N_A_225_74#_M1033_g 0.0282114f $X=6.215 $Y=1.63 $X2=0
+ $Y2=0
cc_659 N_A_595_97#_c_734_n N_A_225_74#_c_1013_n 0.00736296f $X=6.215 $Y=1.63
+ $X2=0 $Y2=0
cc_660 N_A_595_97#_c_734_n N_A_1339_74#_c_1326_n 8.23374e-19 $X=6.215 $Y=1.63
+ $X2=0 $Y2=0
cc_661 N_A_595_97#_c_734_n N_A_1339_74#_c_1331_n 0.0016275f $X=6.215 $Y=1.63
+ $X2=0 $Y2=0
cc_662 N_A_595_97#_c_720_n N_A_27_74#_c_1578_n 0.00584793f $X=3.37 $Y=2.295
+ $X2=0 $Y2=0
cc_663 N_A_595_97#_c_738_n N_A_27_74#_c_1578_n 0.0312384f $X=3.37 $Y=2.515 $X2=0
+ $Y2=0
cc_664 N_A_595_97#_c_734_n N_VPWR_c_1644_n 0.0127991f $X=6.215 $Y=1.63 $X2=0
+ $Y2=0
cc_665 N_A_595_97#_c_734_n N_VPWR_c_1640_n 9.49986e-19 $X=6.215 $Y=1.63 $X2=0
+ $Y2=0
cc_666 N_A_595_97#_M1026_g N_VGND_c_1856_n 0.00316744f $X=4.93 $Y=0.58 $X2=0
+ $Y2=0
cc_667 N_A_595_97#_c_718_n N_VGND_c_1856_n 0.0121682f $X=3.365 $Y=0.695 $X2=0
+ $Y2=0
cc_668 N_A_595_97#_c_721_n N_VGND_c_1856_n 0.0102353f $X=4.015 $Y=1.18 $X2=0
+ $Y2=0
cc_669 N_A_595_97#_c_723_n N_VGND_c_1856_n 0.00161263f $X=4.75 $Y=1.6 $X2=0
+ $Y2=0
cc_670 N_A_595_97#_c_718_n N_VGND_c_1865_n 0.00747853f $X=3.365 $Y=0.695 $X2=0
+ $Y2=0
cc_671 N_A_595_97#_M1026_g N_VGND_c_1872_n 0.00433139f $X=4.93 $Y=0.58 $X2=0
+ $Y2=0
cc_672 N_A_595_97#_M1026_g N_VGND_c_1873_n 0.00145723f $X=4.93 $Y=0.58 $X2=0
+ $Y2=0
cc_673 N_A_595_97#_c_716_n N_VGND_c_1873_n 0.00739087f $X=6.23 $Y=1.12 $X2=0
+ $Y2=0
cc_674 N_A_595_97#_c_728_n N_VGND_c_1873_n 0.0129342f $X=5.75 $Y=1.285 $X2=0
+ $Y2=0
cc_675 N_A_595_97#_c_729_n N_VGND_c_1873_n 0.0072628f $X=5.585 $Y=1.265 $X2=0
+ $Y2=0
cc_676 N_A_595_97#_c_730_n N_VGND_c_1873_n 0.0129582f $X=5.75 $Y=1.195 $X2=0
+ $Y2=0
cc_677 N_A_595_97#_c_716_n N_VGND_c_1874_n 0.00292261f $X=6.23 $Y=1.12 $X2=0
+ $Y2=0
cc_678 N_A_595_97#_M1026_g N_VGND_c_1878_n 0.00822f $X=4.93 $Y=0.58 $X2=0 $Y2=0
cc_679 N_A_595_97#_c_716_n N_VGND_c_1878_n 0.00872613f $X=6.23 $Y=1.12 $X2=0
+ $Y2=0
cc_680 N_A_595_97#_c_718_n N_VGND_c_1878_n 0.00847688f $X=3.365 $Y=0.695 $X2=0
+ $Y2=0
cc_681 N_SET_B_c_898_n N_A_225_74#_c_1027_n 0.00900792f $X=5.315 $Y=2.24 $X2=0
+ $Y2=0
cc_682 N_SET_B_c_891_n N_A_225_74#_c_1012_n 0.00362468f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_683 N_SET_B_c_891_n N_A_225_74#_c_1013_n 0.00681575f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_684 N_SET_B_c_891_n N_A_225_74#_M1035_g 0.00266496f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_685 N_SET_B_c_885_n N_A_1501_92#_M1019_g 0.0389792f $X=7.97 $Y=1.09 $X2=0
+ $Y2=0
cc_686 N_SET_B_c_895_n N_A_1501_92#_M1019_g 0.00214118f $X=8.475 $Y=1.165 $X2=0
+ $Y2=0
cc_687 N_SET_B_c_888_n N_A_1501_92#_c_1203_n 0.016712f $X=8.4 $Y=2.375 $X2=0
+ $Y2=0
cc_688 N_SET_B_c_900_n N_A_1501_92#_c_1204_n 0.0266936f $X=8.4 $Y=2.465 $X2=0
+ $Y2=0
cc_689 N_SET_B_c_885_n N_A_1501_92#_c_1198_n 0.00272879f $X=7.97 $Y=1.09 $X2=0
+ $Y2=0
cc_690 N_SET_B_c_886_n N_A_1501_92#_c_1198_n 0.00543494f $X=8.31 $Y=1.165 $X2=0
+ $Y2=0
cc_691 N_SET_B_c_887_n N_A_1501_92#_c_1198_n 0.00453006f $X=8.045 $Y=1.165 $X2=0
+ $Y2=0
cc_692 N_SET_B_c_891_n N_A_1501_92#_c_1198_n 0.0259693f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_693 SET_B N_A_1501_92#_c_1198_n 0.00256053f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_694 N_SET_B_c_895_n N_A_1501_92#_c_1198_n 0.00140589f $X=8.475 $Y=1.165 $X2=0
+ $Y2=0
cc_695 N_SET_B_c_896_n N_A_1501_92#_c_1198_n 0.0354924f $X=8.475 $Y=1.345 $X2=0
+ $Y2=0
cc_696 N_SET_B_c_887_n N_A_1501_92#_c_1199_n 0.0104285f $X=8.045 $Y=1.165 $X2=0
+ $Y2=0
cc_697 N_SET_B_c_891_n N_A_1501_92#_c_1199_n 0.01006f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_698 SET_B N_A_1501_92#_c_1199_n 0.00139253f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_699 N_SET_B_c_895_n N_A_1501_92#_c_1199_n 0.0171448f $X=8.475 $Y=1.165 $X2=0
+ $Y2=0
cc_700 N_SET_B_c_896_n N_A_1501_92#_c_1199_n 0.00179807f $X=8.475 $Y=1.345 $X2=0
+ $Y2=0
cc_701 N_SET_B_c_886_n N_A_1501_92#_c_1235_n 0.0175303f $X=8.31 $Y=1.165 $X2=0
+ $Y2=0
cc_702 N_SET_B_c_891_n N_A_1501_92#_c_1235_n 0.00610939f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_703 SET_B N_A_1501_92#_c_1235_n 0.00196951f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_704 N_SET_B_c_896_n N_A_1501_92#_c_1235_n 0.0268551f $X=8.475 $Y=1.345 $X2=0
+ $Y2=0
cc_705 N_SET_B_c_885_n N_A_1501_92#_c_1218_n 0.0115671f $X=7.97 $Y=1.09 $X2=0
+ $Y2=0
cc_706 N_SET_B_c_888_n N_A_1501_92#_c_1209_n 6.87016e-19 $X=8.4 $Y=2.375 $X2=0
+ $Y2=0
cc_707 N_SET_B_c_900_n N_A_1501_92#_c_1209_n 4.63768e-19 $X=8.4 $Y=2.465 $X2=0
+ $Y2=0
cc_708 N_SET_B_c_895_n N_A_1339_74#_M1000_g 0.0217685f $X=8.475 $Y=1.165 $X2=0
+ $Y2=0
cc_709 N_SET_B_c_896_n N_A_1339_74#_M1000_g 0.00107899f $X=8.475 $Y=1.345 $X2=0
+ $Y2=0
cc_710 N_SET_B_c_888_n N_A_1339_74#_c_1307_n 0.00455626f $X=8.4 $Y=2.375 $X2=0
+ $Y2=0
cc_711 N_SET_B_c_896_n N_A_1339_74#_c_1307_n 9.08428e-19 $X=8.475 $Y=1.345 $X2=0
+ $Y2=0
cc_712 N_SET_B_c_891_n N_A_1339_74#_c_1326_n 0.00158223f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_713 N_SET_B_c_891_n N_A_1339_74#_c_1315_n 0.0132819f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_714 N_SET_B_c_888_n N_A_1339_74#_c_1327_n 0.0127871f $X=8.4 $Y=2.375 $X2=0
+ $Y2=0
cc_715 N_SET_B_c_900_n N_A_1339_74#_c_1327_n 0.00636464f $X=8.4 $Y=2.465 $X2=0
+ $Y2=0
cc_716 N_SET_B_c_891_n N_A_1339_74#_c_1327_n 0.00979116f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_717 SET_B N_A_1339_74#_c_1327_n 0.0030363f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_718 N_SET_B_c_896_n N_A_1339_74#_c_1327_n 0.0116201f $X=8.475 $Y=1.345 $X2=0
+ $Y2=0
cc_719 N_SET_B_c_888_n N_A_1339_74#_c_1316_n 0.0170386f $X=8.4 $Y=2.375 $X2=0
+ $Y2=0
cc_720 N_SET_B_c_900_n N_A_1339_74#_c_1316_n 0.00268127f $X=8.4 $Y=2.465 $X2=0
+ $Y2=0
cc_721 SET_B N_A_1339_74#_c_1316_n 0.00218127f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_722 N_SET_B_c_895_n N_A_1339_74#_c_1316_n 0.00125511f $X=8.475 $Y=1.165 $X2=0
+ $Y2=0
cc_723 N_SET_B_c_896_n N_A_1339_74#_c_1316_n 0.0392467f $X=8.475 $Y=1.345 $X2=0
+ $Y2=0
cc_724 N_SET_B_c_900_n N_A_1339_74#_c_1329_n 0.00722925f $X=8.4 $Y=2.465 $X2=0
+ $Y2=0
cc_725 N_SET_B_c_891_n N_A_1339_74#_c_1330_n 0.0177625f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_726 N_SET_B_c_900_n N_A_1339_74#_c_1333_n 4.54623e-19 $X=8.4 $Y=2.465 $X2=0
+ $Y2=0
cc_727 N_SET_B_c_891_n N_A_1339_74#_c_1333_n 0.00223482f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_728 N_SET_B_c_891_n N_VPWR_M1036_d 0.00303119f $X=8.255 $Y=1.665 $X2=0 $Y2=0
cc_729 N_SET_B_c_898_n N_VPWR_c_1644_n 0.00180402f $X=5.315 $Y=2.24 $X2=0 $Y2=0
cc_730 N_SET_B_c_900_n N_VPWR_c_1645_n 0.00478933f $X=8.4 $Y=2.465 $X2=0 $Y2=0
cc_731 N_SET_B_c_900_n N_VPWR_c_1659_n 0.00446404f $X=8.4 $Y=2.465 $X2=0 $Y2=0
cc_732 N_SET_B_c_900_n N_VPWR_c_1640_n 0.00460642f $X=8.4 $Y=2.465 $X2=0 $Y2=0
cc_733 N_SET_B_c_891_n A_1258_341# 0.00256567f $X=8.255 $Y=1.665 $X2=-0.19
+ $Y2=-0.245
cc_734 N_SET_B_c_889_n N_VGND_c_1872_n 0.00383152f $X=5.295 $Y=0.865 $X2=0 $Y2=0
cc_735 N_SET_B_c_889_n N_VGND_c_1873_n 0.0116257f $X=5.295 $Y=0.865 $X2=0 $Y2=0
cc_736 N_SET_B_c_885_n N_VGND_c_1874_n 0.00434252f $X=7.97 $Y=1.09 $X2=0 $Y2=0
cc_737 N_SET_B_c_885_n N_VGND_c_1875_n 0.00536598f $X=7.97 $Y=1.09 $X2=0 $Y2=0
cc_738 N_SET_B_c_885_n N_VGND_c_1878_n 0.00479212f $X=7.97 $Y=1.09 $X2=0 $Y2=0
cc_739 N_SET_B_c_889_n N_VGND_c_1878_n 0.00752325f $X=5.295 $Y=0.865 $X2=0 $Y2=0
cc_740 N_A_225_74#_M1035_g N_A_1501_92#_M1019_g 0.0562485f $X=7.19 $Y=0.8 $X2=0
+ $Y2=0
cc_741 N_A_225_74#_c_1012_n N_A_1501_92#_c_1203_n 3.89004e-19 $X=7.115 $Y=1.735
+ $X2=0 $Y2=0
cc_742 N_A_225_74#_M1035_g N_A_1501_92#_c_1199_n 0.00477807f $X=7.19 $Y=0.8
+ $X2=0 $Y2=0
cc_743 N_A_225_74#_M1035_g N_A_1339_74#_c_1336_n 0.0111291f $X=7.19 $Y=0.8 $X2=0
+ $Y2=0
cc_744 N_A_225_74#_M1033_g N_A_1339_74#_c_1326_n 0.0093209f $X=6.72 $Y=2.46
+ $X2=0 $Y2=0
cc_745 N_A_225_74#_c_1012_n N_A_1339_74#_c_1326_n 0.00229379f $X=7.115 $Y=1.735
+ $X2=0 $Y2=0
cc_746 N_A_225_74#_c_1013_n N_A_1339_74#_c_1326_n 0.00166017f $X=6.81 $Y=1.735
+ $X2=0 $Y2=0
cc_747 N_A_225_74#_c_1012_n N_A_1339_74#_c_1315_n 0.00233299f $X=7.115 $Y=1.735
+ $X2=0 $Y2=0
cc_748 N_A_225_74#_M1035_g N_A_1339_74#_c_1315_n 0.0164602f $X=7.19 $Y=0.8 $X2=0
+ $Y2=0
cc_749 N_A_225_74#_c_1012_n N_A_1339_74#_c_1330_n 0.0144662f $X=7.115 $Y=1.735
+ $X2=0 $Y2=0
cc_750 N_A_225_74#_c_1013_n N_A_1339_74#_c_1330_n 0.00313929f $X=6.81 $Y=1.735
+ $X2=0 $Y2=0
cc_751 N_A_225_74#_c_1027_n N_A_1339_74#_c_1331_n 3.82837e-19 $X=6.63 $Y=3.15
+ $X2=0 $Y2=0
cc_752 N_A_225_74#_M1033_g N_A_1339_74#_c_1331_n 0.0144344f $X=6.72 $Y=2.46
+ $X2=0 $Y2=0
cc_753 N_A_225_74#_c_1012_n N_A_1339_74#_c_1331_n 0.00199255f $X=7.115 $Y=1.735
+ $X2=0 $Y2=0
cc_754 N_A_225_74#_M1029_s N_A_27_74#_c_1577_n 0.0126187f $X=1.145 $Y=1.79 $X2=0
+ $Y2=0
cc_755 N_A_225_74#_c_1035_n N_A_27_74#_c_1577_n 0.0190006f $X=1.305 $Y=1.87
+ $X2=0 $Y2=0
cc_756 N_A_225_74#_c_1036_n N_A_27_74#_c_1577_n 0.0142272f $X=1.145 $Y=1.87
+ $X2=0 $Y2=0
cc_757 N_A_225_74#_c_1037_n N_A_27_74#_c_1577_n 0.0057885f $X=1.945 $Y=1.805
+ $X2=0 $Y2=0
cc_758 N_A_225_74#_c_1009_n N_A_27_74#_c_1578_n 0.0149932f $X=1.965 $Y=1.715
+ $X2=0 $Y2=0
cc_759 N_A_225_74#_c_1021_n N_A_27_74#_c_1578_n 0.025647f $X=2.485 $Y=3.075
+ $X2=0 $Y2=0
cc_760 N_A_225_74#_c_1016_n N_A_27_74#_c_1578_n 0.00492213f $X=2.41 $Y=1.465
+ $X2=0 $Y2=0
cc_761 N_A_225_74#_c_1037_n N_A_27_74#_c_1578_n 0.0278803f $X=1.945 $Y=1.805
+ $X2=0 $Y2=0
cc_762 N_A_225_74#_M1015_g N_A_27_74#_c_1572_n 7.39226e-19 $X=1.915 $Y=0.74
+ $X2=0 $Y2=0
cc_763 N_A_225_74#_c_1009_n N_A_27_74#_c_1572_n 0.00116731f $X=1.965 $Y=1.715
+ $X2=0 $Y2=0
cc_764 N_A_225_74#_c_1021_n N_A_27_74#_c_1572_n 0.00988666f $X=2.485 $Y=3.075
+ $X2=0 $Y2=0
cc_765 N_A_225_74#_c_1010_n N_A_27_74#_c_1572_n 0.00583176f $X=2.825 $Y=1.12
+ $X2=0 $Y2=0
cc_766 N_A_225_74#_M1014_g N_A_27_74#_c_1572_n 0.00236295f $X=2.9 $Y=0.695 $X2=0
+ $Y2=0
cc_767 N_A_225_74#_c_1015_n N_A_27_74#_c_1572_n 0.0188485f $X=2.485 $Y=1.12
+ $X2=0 $Y2=0
cc_768 N_A_225_74#_c_1037_n N_A_27_74#_c_1572_n 0.0135406f $X=1.945 $Y=1.805
+ $X2=0 $Y2=0
cc_769 N_A_225_74#_c_1018_n N_A_27_74#_c_1572_n 0.0302859f $X=2.11 $Y=1.465
+ $X2=0 $Y2=0
cc_770 N_A_225_74#_c_1009_n N_A_27_74#_c_1623_n 0.00185704f $X=1.965 $Y=1.715
+ $X2=0 $Y2=0
cc_771 N_A_225_74#_c_1037_n N_A_27_74#_c_1623_n 0.0112057f $X=1.945 $Y=1.805
+ $X2=0 $Y2=0
cc_772 N_A_225_74#_c_1010_n N_A_27_74#_c_1574_n 0.00610954f $X=2.825 $Y=1.12
+ $X2=0 $Y2=0
cc_773 N_A_225_74#_M1014_g N_A_27_74#_c_1574_n 4.22296e-19 $X=2.9 $Y=0.695 $X2=0
+ $Y2=0
cc_774 N_A_225_74#_c_1015_n N_A_27_74#_c_1574_n 9.83875e-19 $X=2.485 $Y=1.12
+ $X2=0 $Y2=0
cc_775 N_A_225_74#_c_1037_n N_VPWR_M1029_d 0.00196757f $X=1.945 $Y=1.805 $X2=0
+ $Y2=0
cc_776 N_A_225_74#_c_1009_n N_VPWR_c_1642_n 0.00746791f $X=1.965 $Y=1.715 $X2=0
+ $Y2=0
cc_777 N_A_225_74#_c_1021_n N_VPWR_c_1642_n 3.21585e-19 $X=2.485 $Y=3.075 $X2=0
+ $Y2=0
cc_778 N_A_225_74#_c_1023_n N_VPWR_c_1642_n 0.00272925f $X=2.56 $Y=3.15 $X2=0
+ $Y2=0
cc_779 N_A_225_74#_c_1025_n N_VPWR_c_1643_n 7.29299e-19 $X=3.455 $Y=3.075 $X2=0
+ $Y2=0
cc_780 N_A_225_74#_c_1027_n N_VPWR_c_1643_n 0.0250524f $X=6.63 $Y=3.15 $X2=0
+ $Y2=0
cc_781 N_A_225_74#_c_1027_n N_VPWR_c_1644_n 0.0290026f $X=6.63 $Y=3.15 $X2=0
+ $Y2=0
cc_782 N_A_225_74#_M1033_g N_VPWR_c_1644_n 0.0055399f $X=6.72 $Y=2.46 $X2=0
+ $Y2=0
cc_783 N_A_225_74#_c_1027_n N_VPWR_c_1651_n 0.0262434f $X=6.63 $Y=3.15 $X2=0
+ $Y2=0
cc_784 N_A_225_74#_c_1009_n N_VPWR_c_1657_n 0.0048608f $X=1.965 $Y=1.715 $X2=0
+ $Y2=0
cc_785 N_A_225_74#_c_1023_n N_VPWR_c_1657_n 0.0368442f $X=2.56 $Y=3.15 $X2=0
+ $Y2=0
cc_786 N_A_225_74#_c_1027_n N_VPWR_c_1658_n 0.0322942f $X=6.63 $Y=3.15 $X2=0
+ $Y2=0
cc_787 N_A_225_74#_c_1009_n N_VPWR_c_1640_n 0.00480464f $X=1.965 $Y=1.715 $X2=0
+ $Y2=0
cc_788 N_A_225_74#_c_1022_n N_VPWR_c_1640_n 0.0189646f $X=3.365 $Y=3.15 $X2=0
+ $Y2=0
cc_789 N_A_225_74#_c_1023_n N_VPWR_c_1640_n 0.00604517f $X=2.56 $Y=3.15 $X2=0
+ $Y2=0
cc_790 N_A_225_74#_c_1027_n N_VPWR_c_1640_n 0.0880736f $X=6.63 $Y=3.15 $X2=0
+ $Y2=0
cc_791 N_A_225_74#_c_1033_n N_VPWR_c_1640_n 0.00441524f $X=3.455 $Y=3.15 $X2=0
+ $Y2=0
cc_792 N_A_225_74#_c_1019_n N_VGND_c_1853_n 0.0363632f $X=1.27 $Y=0.515 $X2=0
+ $Y2=0
cc_793 N_A_225_74#_c_1019_n N_VGND_c_1854_n 0.0203368f $X=1.27 $Y=0.515 $X2=0
+ $Y2=0
cc_794 N_A_225_74#_M1015_g N_VGND_c_1855_n 0.0115939f $X=1.915 $Y=0.74 $X2=0
+ $Y2=0
cc_795 N_A_225_74#_c_1019_n N_VGND_c_1855_n 0.0268179f $X=1.27 $Y=0.515 $X2=0
+ $Y2=0
cc_796 N_A_225_74#_M1015_g N_VGND_c_1865_n 0.00383152f $X=1.915 $Y=0.74 $X2=0
+ $Y2=0
cc_797 N_A_225_74#_M1014_g N_VGND_c_1865_n 7.53287e-19 $X=2.9 $Y=0.695 $X2=0
+ $Y2=0
cc_798 N_A_225_74#_M1015_g N_VGND_c_1878_n 0.00762539f $X=1.915 $Y=0.74 $X2=0
+ $Y2=0
cc_799 N_A_225_74#_c_1019_n N_VGND_c_1878_n 0.0167889f $X=1.27 $Y=0.515 $X2=0
+ $Y2=0
cc_800 N_A_1501_92#_c_1235_n N_A_1339_74#_M1000_g 0.0152859f $X=9.105 $Y=0.925
+ $X2=0 $Y2=0
cc_801 N_A_1501_92#_c_1201_n N_A_1339_74#_M1000_g 0.00338973f $X=9.825 $Y=2.29
+ $X2=0 $Y2=0
cc_802 N_A_1501_92#_c_1202_n N_A_1339_74#_M1000_g 0.00714524f $X=9.27 $Y=0.8
+ $X2=0 $Y2=0
cc_803 N_A_1501_92#_c_1202_n N_A_1339_74#_c_1306_n 0.00226453f $X=9.27 $Y=0.8
+ $X2=0 $Y2=0
cc_804 N_A_1501_92#_c_1209_n N_A_1339_74#_c_1307_n 9.92746e-19 $X=9.18 $Y=2.375
+ $X2=0 $Y2=0
cc_805 N_A_1501_92#_c_1207_n N_A_1339_74#_c_1320_n 0.0086189f $X=9.74 $Y=2.375
+ $X2=0 $Y2=0
cc_806 N_A_1501_92#_c_1201_n N_A_1339_74#_c_1320_n 0.00483477f $X=9.825 $Y=2.29
+ $X2=0 $Y2=0
cc_807 N_A_1501_92#_c_1209_n N_A_1339_74#_c_1320_n 8.18421e-19 $X=9.18 $Y=2.375
+ $X2=0 $Y2=0
cc_808 N_A_1501_92#_c_1207_n N_A_1339_74#_c_1308_n 0.00364281f $X=9.74 $Y=2.375
+ $X2=0 $Y2=0
cc_809 N_A_1501_92#_c_1201_n N_A_1339_74#_c_1308_n 0.0201283f $X=9.825 $Y=2.29
+ $X2=0 $Y2=0
cc_810 N_A_1501_92#_c_1201_n N_A_1339_74#_c_1321_n 0.00332862f $X=9.825 $Y=2.29
+ $X2=0 $Y2=0
cc_811 N_A_1501_92#_c_1209_n N_A_1339_74#_c_1321_n 0.00371656f $X=9.18 $Y=2.375
+ $X2=0 $Y2=0
cc_812 N_A_1501_92#_c_1200_n N_A_1339_74#_M1009_g 0.00412514f $X=9.74 $Y=1.095
+ $X2=0 $Y2=0
cc_813 N_A_1501_92#_c_1201_n N_A_1339_74#_M1009_g 0.00391208f $X=9.825 $Y=2.29
+ $X2=0 $Y2=0
cc_814 N_A_1501_92#_c_1202_n N_A_1339_74#_M1009_g 0.00398937f $X=9.27 $Y=0.8
+ $X2=0 $Y2=0
cc_815 N_A_1501_92#_c_1201_n N_A_1339_74#_c_1312_n 0.00138342f $X=9.825 $Y=2.29
+ $X2=0 $Y2=0
cc_816 N_A_1501_92#_M1019_g N_A_1339_74#_c_1336_n 3.11108e-19 $X=7.58 $Y=0.8
+ $X2=0 $Y2=0
cc_817 N_A_1501_92#_M1019_g N_A_1339_74#_c_1315_n 6.18383e-19 $X=7.58 $Y=0.8
+ $X2=0 $Y2=0
cc_818 N_A_1501_92#_c_1203_n N_A_1339_74#_c_1327_n 0.0111898f $X=7.95 $Y=2.375
+ $X2=0 $Y2=0
cc_819 N_A_1501_92#_c_1204_n N_A_1339_74#_c_1327_n 0.00528f $X=7.95 $Y=2.465
+ $X2=0 $Y2=0
cc_820 N_A_1501_92#_M1007_s N_A_1339_74#_c_1316_n 0.00624391f $X=9.035 $Y=1.84
+ $X2=0 $Y2=0
cc_821 N_A_1501_92#_c_1235_n N_A_1339_74#_c_1316_n 0.00784261f $X=9.105 $Y=0.925
+ $X2=0 $Y2=0
cc_822 N_A_1501_92#_c_1207_n N_A_1339_74#_c_1316_n 0.0146209f $X=9.74 $Y=2.375
+ $X2=0 $Y2=0
cc_823 N_A_1501_92#_c_1200_n N_A_1339_74#_c_1316_n 0.0107886f $X=9.74 $Y=1.095
+ $X2=0 $Y2=0
cc_824 N_A_1501_92#_c_1201_n N_A_1339_74#_c_1316_n 0.0485702f $X=9.825 $Y=2.29
+ $X2=0 $Y2=0
cc_825 N_A_1501_92#_c_1209_n N_A_1339_74#_c_1316_n 0.0419706f $X=9.18 $Y=2.375
+ $X2=0 $Y2=0
cc_826 N_A_1501_92#_c_1202_n N_A_1339_74#_c_1316_n 0.0286983f $X=9.27 $Y=0.8
+ $X2=0 $Y2=0
cc_827 N_A_1501_92#_c_1204_n N_A_1339_74#_c_1329_n 5.12307e-19 $X=7.95 $Y=2.465
+ $X2=0 $Y2=0
cc_828 N_A_1501_92#_c_1209_n N_A_1339_74#_c_1329_n 0.00954915f $X=9.18 $Y=2.375
+ $X2=0 $Y2=0
cc_829 N_A_1501_92#_c_1204_n N_A_1339_74#_c_1331_n 9.77004e-19 $X=7.95 $Y=2.465
+ $X2=0 $Y2=0
cc_830 N_A_1501_92#_c_1203_n N_A_1339_74#_c_1333_n 0.00628426f $X=7.95 $Y=2.375
+ $X2=0 $Y2=0
cc_831 N_A_1501_92#_c_1204_n N_A_1339_74#_c_1333_n 0.00760762f $X=7.95 $Y=2.465
+ $X2=0 $Y2=0
cc_832 N_A_1501_92#_c_1198_n N_A_1339_74#_c_1333_n 0.0237116f $X=7.89 $Y=1.615
+ $X2=0 $Y2=0
cc_833 N_A_1501_92#_c_1199_n N_A_1339_74#_c_1333_n 8.67582e-19 $X=7.89 $Y=1.615
+ $X2=0 $Y2=0
cc_834 N_A_1501_92#_c_1207_n N_A_1339_74#_c_1317_n 2.15983e-19 $X=9.74 $Y=2.375
+ $X2=0 $Y2=0
cc_835 N_A_1501_92#_c_1200_n N_A_1339_74#_c_1317_n 0.00717173f $X=9.74 $Y=1.095
+ $X2=0 $Y2=0
cc_836 N_A_1501_92#_c_1201_n N_A_1339_74#_c_1317_n 9.58673e-19 $X=9.825 $Y=2.29
+ $X2=0 $Y2=0
cc_837 N_A_1501_92#_c_1207_n N_VPWR_M1007_d 0.00546255f $X=9.74 $Y=2.375 $X2=0
+ $Y2=0
cc_838 N_A_1501_92#_c_1201_n N_VPWR_M1007_d 0.0079206f $X=9.825 $Y=2.29 $X2=0
+ $Y2=0
cc_839 N_A_1501_92#_c_1204_n N_VPWR_c_1645_n 0.00539382f $X=7.95 $Y=2.465 $X2=0
+ $Y2=0
cc_840 N_A_1501_92#_c_1207_n N_VPWR_c_1646_n 0.0221894f $X=9.74 $Y=2.375 $X2=0
+ $Y2=0
cc_841 N_A_1501_92#_c_1204_n N_VPWR_c_1651_n 0.00422316f $X=7.95 $Y=2.465 $X2=0
+ $Y2=0
cc_842 N_A_1501_92#_c_1209_n N_VPWR_c_1659_n 0.00541079f $X=9.18 $Y=2.375 $X2=0
+ $Y2=0
cc_843 N_A_1501_92#_c_1204_n N_VPWR_c_1640_n 0.00453881f $X=7.95 $Y=2.465 $X2=0
+ $Y2=0
cc_844 N_A_1501_92#_c_1209_n N_VPWR_c_1640_n 0.00910369f $X=9.18 $Y=2.375 $X2=0
+ $Y2=0
cc_845 N_A_1501_92#_c_1200_n Q_N 0.00736666f $X=9.74 $Y=1.095 $X2=0 $Y2=0
cc_846 N_A_1501_92#_c_1201_n Q_N 0.0342331f $X=9.825 $Y=2.29 $X2=0 $Y2=0
cc_847 N_A_1501_92#_c_1201_n Q_N 0.00124835f $X=9.825 $Y=2.29 $X2=0 $Y2=0
cc_848 N_A_1501_92#_c_1235_n N_VGND_M1037_d 0.0237418f $X=9.105 $Y=0.925 $X2=0
+ $Y2=0
cc_849 N_A_1501_92#_c_1200_n N_VGND_M1009_s 0.00461825f $X=9.74 $Y=1.095 $X2=0
+ $Y2=0
cc_850 N_A_1501_92#_c_1200_n N_VGND_c_1857_n 0.0213705f $X=9.74 $Y=1.095 $X2=0
+ $Y2=0
cc_851 N_A_1501_92#_c_1202_n N_VGND_c_1857_n 0.0138209f $X=9.27 $Y=0.8 $X2=0
+ $Y2=0
cc_852 N_A_1501_92#_c_1202_n N_VGND_c_1866_n 0.00623106f $X=9.27 $Y=0.8 $X2=0
+ $Y2=0
cc_853 N_A_1501_92#_M1019_g N_VGND_c_1874_n 0.00311027f $X=7.58 $Y=0.8 $X2=0
+ $Y2=0
cc_854 N_A_1501_92#_c_1235_n N_VGND_c_1875_n 0.0586839f $X=9.105 $Y=0.925 $X2=0
+ $Y2=0
cc_855 N_A_1501_92#_M1019_g N_VGND_c_1878_n 0.00321167f $X=7.58 $Y=0.8 $X2=0
+ $Y2=0
cc_856 N_A_1501_92#_c_1235_n N_VGND_c_1878_n 0.0123962f $X=9.105 $Y=0.925 $X2=0
+ $Y2=0
cc_857 N_A_1501_92#_c_1218_n N_VGND_c_1878_n 0.0124246f $X=8.055 $Y=0.925 $X2=0
+ $Y2=0
cc_858 N_A_1501_92#_c_1202_n N_VGND_c_1878_n 0.00984494f $X=9.27 $Y=0.8 $X2=0
+ $Y2=0
cc_859 N_A_1501_92#_c_1218_n A_1531_118# 0.00412701f $X=8.055 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_860 N_A_1339_74#_c_1324_n N_A_2221_74#_c_1506_n 0.0157102f $X=11.475 $Y=1.765
+ $X2=0 $Y2=0
cc_861 N_A_1339_74#_M1006_g N_A_2221_74#_M1001_g 0.0226536f $X=11.465 $Y=0.69
+ $X2=0 $Y2=0
cc_862 N_A_1339_74#_M1020_g N_A_2221_74#_c_1501_n 0.00404932f $X=10.475 $Y=0.74
+ $X2=0 $Y2=0
cc_863 N_A_1339_74#_M1006_g N_A_2221_74#_c_1501_n 0.0189532f $X=11.465 $Y=0.69
+ $X2=0 $Y2=0
cc_864 N_A_1339_74#_c_1322_n N_A_2221_74#_c_1502_n 0.00261093f $X=10.47 $Y=1.765
+ $X2=0 $Y2=0
cc_865 N_A_1339_74#_c_1312_n N_A_2221_74#_c_1502_n 0.00223156f $X=10.56 $Y=1.49
+ $X2=0 $Y2=0
cc_866 N_A_1339_74#_c_1324_n N_A_2221_74#_c_1502_n 0.0137849f $X=11.475 $Y=1.765
+ $X2=0 $Y2=0
cc_867 N_A_1339_74#_c_1314_n N_A_2221_74#_c_1502_n 0.00580251f $X=11.475
+ $Y=1.557 $X2=0 $Y2=0
cc_868 N_A_1339_74#_M1006_g N_A_2221_74#_c_1503_n 0.00696112f $X=11.465 $Y=0.69
+ $X2=0 $Y2=0
cc_869 N_A_1339_74#_c_1314_n N_A_2221_74#_c_1503_n 0.013869f $X=11.475 $Y=1.557
+ $X2=0 $Y2=0
cc_870 N_A_1339_74#_M1020_g N_A_2221_74#_c_1504_n 8.258e-19 $X=10.475 $Y=0.74
+ $X2=0 $Y2=0
cc_871 N_A_1339_74#_c_1311_n N_A_2221_74#_c_1504_n 0.0290202f $X=11.385 $Y=1.49
+ $X2=0 $Y2=0
cc_872 N_A_1339_74#_M1006_g N_A_2221_74#_c_1504_n 0.00110532f $X=11.465 $Y=0.69
+ $X2=0 $Y2=0
cc_873 N_A_1339_74#_c_1314_n N_A_2221_74#_c_1504_n 7.90981e-19 $X=11.475
+ $Y=1.557 $X2=0 $Y2=0
cc_874 N_A_1339_74#_M1006_g N_A_2221_74#_c_1505_n 0.00280567f $X=11.465 $Y=0.69
+ $X2=0 $Y2=0
cc_875 N_A_1339_74#_c_1314_n N_A_2221_74#_c_1505_n 0.0228968f $X=11.475 $Y=1.557
+ $X2=0 $Y2=0
cc_876 N_A_1339_74#_c_1327_n N_VPWR_c_1645_n 0.0147304f $X=8.46 $Y=2.215 $X2=0
+ $Y2=0
cc_877 N_A_1339_74#_c_1329_n N_VPWR_c_1645_n 0.0172613f $X=8.625 $Y=2.75 $X2=0
+ $Y2=0
cc_878 N_A_1339_74#_c_1331_n N_VPWR_c_1645_n 0.00924952f $X=7.47 $Y=2.73 $X2=0
+ $Y2=0
cc_879 N_A_1339_74#_c_1321_n N_VPWR_c_1646_n 0.00902525f $X=10.02 $Y=1.765 $X2=0
+ $Y2=0
cc_880 N_A_1339_74#_c_1322_n N_VPWR_c_1646_n 4.59453e-19 $X=10.47 $Y=1.765 $X2=0
+ $Y2=0
cc_881 N_A_1339_74#_c_1322_n N_VPWR_c_1647_n 0.0081876f $X=10.47 $Y=1.765 $X2=0
+ $Y2=0
cc_882 N_A_1339_74#_c_1311_n N_VPWR_c_1647_n 0.0109752f $X=11.385 $Y=1.49 $X2=0
+ $Y2=0
cc_883 N_A_1339_74#_c_1324_n N_VPWR_c_1647_n 0.00442583f $X=11.475 $Y=1.765
+ $X2=0 $Y2=0
cc_884 N_A_1339_74#_c_1324_n N_VPWR_c_1648_n 0.012094f $X=11.475 $Y=1.765 $X2=0
+ $Y2=0
cc_885 N_A_1339_74#_c_1331_n N_VPWR_c_1651_n 0.0298791f $X=7.47 $Y=2.73 $X2=0
+ $Y2=0
cc_886 N_A_1339_74#_c_1332_n N_VPWR_c_1651_n 0.00628522f $X=7.75 $Y=2.3 $X2=0
+ $Y2=0
cc_887 N_A_1339_74#_c_1321_n N_VPWR_c_1653_n 0.00413917f $X=10.02 $Y=1.765 $X2=0
+ $Y2=0
cc_888 N_A_1339_74#_c_1322_n N_VPWR_c_1653_n 0.00417628f $X=10.47 $Y=1.765 $X2=0
+ $Y2=0
cc_889 N_A_1339_74#_c_1329_n N_VPWR_c_1659_n 0.0103126f $X=8.625 $Y=2.75 $X2=0
+ $Y2=0
cc_890 N_A_1339_74#_c_1324_n N_VPWR_c_1660_n 0.00481995f $X=11.475 $Y=1.765
+ $X2=0 $Y2=0
cc_891 N_A_1339_74#_c_1321_n N_VPWR_c_1640_n 0.00817726f $X=10.02 $Y=1.765 $X2=0
+ $Y2=0
cc_892 N_A_1339_74#_c_1322_n N_VPWR_c_1640_n 0.00770846f $X=10.47 $Y=1.765 $X2=0
+ $Y2=0
cc_893 N_A_1339_74#_c_1324_n N_VPWR_c_1640_n 0.00508379f $X=11.475 $Y=1.765
+ $X2=0 $Y2=0
cc_894 N_A_1339_74#_c_1327_n N_VPWR_c_1640_n 0.0129045f $X=8.46 $Y=2.215 $X2=0
+ $Y2=0
cc_895 N_A_1339_74#_c_1329_n N_VPWR_c_1640_n 0.0115456f $X=8.625 $Y=2.75 $X2=0
+ $Y2=0
cc_896 N_A_1339_74#_c_1331_n N_VPWR_c_1640_n 0.0249947f $X=7.47 $Y=2.73 $X2=0
+ $Y2=0
cc_897 N_A_1339_74#_c_1332_n N_VPWR_c_1640_n 0.011801f $X=7.75 $Y=2.3 $X2=0
+ $Y2=0
cc_898 N_A_1339_74#_c_1332_n A_1521_508# 0.00159274f $X=7.75 $Y=2.3 $X2=-0.19
+ $Y2=-0.245
cc_899 N_A_1339_74#_c_1333_n A_1521_508# 0.00130845f $X=7.92 $Y=2.3 $X2=-0.19
+ $Y2=-0.245
cc_900 N_A_1339_74#_c_1321_n Q_N 4.63609e-19 $X=10.02 $Y=1.765 $X2=0 $Y2=0
cc_901 N_A_1339_74#_M1009_g Q_N 0.00249434f $X=10.045 $Y=0.74 $X2=0 $Y2=0
cc_902 N_A_1339_74#_c_1322_n Q_N 0.00172358f $X=10.47 $Y=1.765 $X2=0 $Y2=0
cc_903 N_A_1339_74#_M1020_g Q_N 0.0170389f $X=10.475 $Y=0.74 $X2=0 $Y2=0
cc_904 N_A_1339_74#_c_1312_n Q_N 0.0334259f $X=10.56 $Y=1.49 $X2=0 $Y2=0
cc_905 N_A_1339_74#_c_1321_n Q_N 4.35663e-19 $X=10.02 $Y=1.765 $X2=0 $Y2=0
cc_906 N_A_1339_74#_c_1322_n Q_N 0.00197146f $X=10.47 $Y=1.765 $X2=0 $Y2=0
cc_907 N_A_1339_74#_c_1312_n Q_N 0.00208351f $X=10.56 $Y=1.49 $X2=0 $Y2=0
cc_908 N_A_1339_74#_c_1322_n Q_N 0.0125507f $X=10.47 $Y=1.765 $X2=0 $Y2=0
cc_909 N_A_1339_74#_M1006_g Q 4.4789e-19 $X=11.465 $Y=0.69 $X2=0 $Y2=0
cc_910 N_A_1339_74#_M1000_g N_VGND_c_1857_n 0.00440494f $X=8.975 $Y=0.8 $X2=0
+ $Y2=0
cc_911 N_A_1339_74#_c_1308_n N_VGND_c_1857_n 6.73898e-19 $X=9.93 $Y=1.49 $X2=0
+ $Y2=0
cc_912 N_A_1339_74#_M1009_g N_VGND_c_1857_n 0.0136519f $X=10.045 $Y=0.74 $X2=0
+ $Y2=0
cc_913 N_A_1339_74#_M1020_g N_VGND_c_1857_n 5.19194e-19 $X=10.475 $Y=0.74 $X2=0
+ $Y2=0
cc_914 N_A_1339_74#_M1020_g N_VGND_c_1858_n 0.00510543f $X=10.475 $Y=0.74 $X2=0
+ $Y2=0
cc_915 N_A_1339_74#_c_1311_n N_VGND_c_1858_n 0.00886118f $X=11.385 $Y=1.49 $X2=0
+ $Y2=0
cc_916 N_A_1339_74#_M1006_g N_VGND_c_1858_n 0.00422013f $X=11.465 $Y=0.69 $X2=0
+ $Y2=0
cc_917 N_A_1339_74#_M1006_g N_VGND_c_1859_n 0.00744279f $X=11.465 $Y=0.69 $X2=0
+ $Y2=0
cc_918 N_A_1339_74#_M1009_g N_VGND_c_1862_n 0.00383152f $X=10.045 $Y=0.74 $X2=0
+ $Y2=0
cc_919 N_A_1339_74#_M1020_g N_VGND_c_1862_n 0.00422942f $X=10.475 $Y=0.74 $X2=0
+ $Y2=0
cc_920 N_A_1339_74#_M1000_g N_VGND_c_1866_n 0.00434252f $X=8.975 $Y=0.8 $X2=0
+ $Y2=0
cc_921 N_A_1339_74#_M1006_g N_VGND_c_1867_n 0.00434272f $X=11.465 $Y=0.69 $X2=0
+ $Y2=0
cc_922 N_A_1339_74#_M1000_g N_VGND_c_1875_n 0.00754579f $X=8.975 $Y=0.8 $X2=0
+ $Y2=0
cc_923 N_A_1339_74#_M1000_g N_VGND_c_1878_n 0.00479212f $X=8.975 $Y=0.8 $X2=0
+ $Y2=0
cc_924 N_A_1339_74#_M1009_g N_VGND_c_1878_n 0.0075754f $X=10.045 $Y=0.74 $X2=0
+ $Y2=0
cc_925 N_A_1339_74#_M1020_g N_VGND_c_1878_n 0.00788596f $X=10.475 $Y=0.74 $X2=0
+ $Y2=0
cc_926 N_A_1339_74#_M1006_g N_VGND_c_1878_n 0.00826311f $X=11.465 $Y=0.69 $X2=0
+ $Y2=0
cc_927 N_A_2221_74#_c_1502_n N_VPWR_c_1647_n 0.0698272f $X=11.25 $Y=1.985 $X2=0
+ $Y2=0
cc_928 N_A_2221_74#_c_1506_n N_VPWR_c_1648_n 0.00911255f $X=12.005 $Y=1.765
+ $X2=0 $Y2=0
cc_929 N_A_2221_74#_c_1502_n N_VPWR_c_1648_n 0.0697922f $X=11.25 $Y=1.985 $X2=0
+ $Y2=0
cc_930 N_A_2221_74#_c_1503_n N_VPWR_c_1648_n 0.0199046f $X=11.94 $Y=1.465 $X2=0
+ $Y2=0
cc_931 N_A_2221_74#_c_1505_n N_VPWR_c_1648_n 0.00205259f $X=12.455 $Y=1.532
+ $X2=0 $Y2=0
cc_932 N_A_2221_74#_c_1507_n N_VPWR_c_1650_n 0.00954146f $X=12.455 $Y=1.765
+ $X2=0 $Y2=0
cc_933 N_A_2221_74#_c_1502_n N_VPWR_c_1660_n 0.0097982f $X=11.25 $Y=1.985 $X2=0
+ $Y2=0
cc_934 N_A_2221_74#_c_1506_n N_VPWR_c_1661_n 0.00445602f $X=12.005 $Y=1.765
+ $X2=0 $Y2=0
cc_935 N_A_2221_74#_c_1507_n N_VPWR_c_1661_n 0.00411612f $X=12.455 $Y=1.765
+ $X2=0 $Y2=0
cc_936 N_A_2221_74#_c_1506_n N_VPWR_c_1640_n 0.00862391f $X=12.005 $Y=1.765
+ $X2=0 $Y2=0
cc_937 N_A_2221_74#_c_1507_n N_VPWR_c_1640_n 0.00751023f $X=12.455 $Y=1.765
+ $X2=0 $Y2=0
cc_938 N_A_2221_74#_c_1502_n N_VPWR_c_1640_n 0.0111907f $X=11.25 $Y=1.985 $X2=0
+ $Y2=0
cc_939 N_A_2221_74#_c_1501_n Q_N 0.00476669f $X=11.25 $Y=0.515 $X2=0 $Y2=0
cc_940 N_A_2221_74#_c_1502_n Q_N 0.00530548f $X=11.25 $Y=1.985 $X2=0 $Y2=0
cc_941 N_A_2221_74#_c_1504_n Q_N 0.00865359f $X=11.25 $Y=1.465 $X2=0 $Y2=0
cc_942 N_A_2221_74#_c_1506_n N_Q_c_1824_n 0.0110945f $X=12.005 $Y=1.765 $X2=0
+ $Y2=0
cc_943 N_A_2221_74#_c_1507_n N_Q_c_1824_n 0.0130738f $X=12.455 $Y=1.765 $X2=0
+ $Y2=0
cc_944 N_A_2221_74#_c_1506_n N_Q_c_1825_n 0.00230932f $X=12.005 $Y=1.765 $X2=0
+ $Y2=0
cc_945 N_A_2221_74#_c_1507_n N_Q_c_1825_n 0.00240464f $X=12.455 $Y=1.765 $X2=0
+ $Y2=0
cc_946 N_A_2221_74#_c_1503_n N_Q_c_1825_n 0.00140951f $X=11.94 $Y=1.465 $X2=0
+ $Y2=0
cc_947 N_A_2221_74#_c_1505_n N_Q_c_1825_n 0.00807114f $X=12.455 $Y=1.532 $X2=0
+ $Y2=0
cc_948 N_A_2221_74#_M1001_g N_Q_c_1821_n 0.0025553f $X=12.035 $Y=0.74 $X2=0
+ $Y2=0
cc_949 N_A_2221_74#_c_1507_n N_Q_c_1821_n 0.0030228f $X=12.455 $Y=1.765 $X2=0
+ $Y2=0
cc_950 N_A_2221_74#_M1011_g N_Q_c_1821_n 0.00866774f $X=12.465 $Y=0.74 $X2=0
+ $Y2=0
cc_951 N_A_2221_74#_c_1503_n N_Q_c_1821_n 0.0249855f $X=11.94 $Y=1.465 $X2=0
+ $Y2=0
cc_952 N_A_2221_74#_c_1505_n N_Q_c_1821_n 0.0358812f $X=12.455 $Y=1.532 $X2=0
+ $Y2=0
cc_953 N_A_2221_74#_M1001_g Q 0.00746865f $X=12.035 $Y=0.74 $X2=0 $Y2=0
cc_954 N_A_2221_74#_M1011_g Q 0.0081896f $X=12.465 $Y=0.74 $X2=0 $Y2=0
cc_955 N_A_2221_74#_M1001_g Q 0.00416712f $X=12.035 $Y=0.74 $X2=0 $Y2=0
cc_956 N_A_2221_74#_M1011_g Q 0.00215589f $X=12.465 $Y=0.74 $X2=0 $Y2=0
cc_957 N_A_2221_74#_c_1501_n Q 0.00238899f $X=11.25 $Y=0.515 $X2=0 $Y2=0
cc_958 N_A_2221_74#_c_1505_n Q 0.00244427f $X=12.455 $Y=1.532 $X2=0 $Y2=0
cc_959 N_A_2221_74#_c_1501_n N_VGND_c_1858_n 0.051504f $X=11.25 $Y=0.515 $X2=0
+ $Y2=0
cc_960 N_A_2221_74#_M1001_g N_VGND_c_1859_n 0.00737997f $X=12.035 $Y=0.74 $X2=0
+ $Y2=0
cc_961 N_A_2221_74#_c_1501_n N_VGND_c_1859_n 0.0270962f $X=11.25 $Y=0.515 $X2=0
+ $Y2=0
cc_962 N_A_2221_74#_c_1503_n N_VGND_c_1859_n 0.019673f $X=11.94 $Y=1.465 $X2=0
+ $Y2=0
cc_963 N_A_2221_74#_c_1505_n N_VGND_c_1859_n 0.00301993f $X=12.455 $Y=1.532
+ $X2=0 $Y2=0
cc_964 N_A_2221_74#_M1011_g N_VGND_c_1861_n 0.00646793f $X=12.465 $Y=0.74 $X2=0
+ $Y2=0
cc_965 N_A_2221_74#_c_1501_n N_VGND_c_1867_n 0.0145639f $X=11.25 $Y=0.515 $X2=0
+ $Y2=0
cc_966 N_A_2221_74#_M1001_g N_VGND_c_1868_n 0.00434272f $X=12.035 $Y=0.74 $X2=0
+ $Y2=0
cc_967 N_A_2221_74#_M1011_g N_VGND_c_1868_n 0.00422942f $X=12.465 $Y=0.74 $X2=0
+ $Y2=0
cc_968 N_A_2221_74#_M1001_g N_VGND_c_1878_n 0.00821312f $X=12.035 $Y=0.74 $X2=0
+ $Y2=0
cc_969 N_A_2221_74#_M1011_g N_VGND_c_1878_n 0.00787255f $X=12.465 $Y=0.74 $X2=0
+ $Y2=0
cc_970 N_A_2221_74#_c_1501_n N_VGND_c_1878_n 0.0119984f $X=11.25 $Y=0.515 $X2=0
+ $Y2=0
cc_971 N_A_27_74#_c_1578_n N_VPWR_M1029_d 0.00134035f $X=2.445 $Y=2.145 $X2=0
+ $Y2=0
cc_972 N_A_27_74#_c_1623_n N_VPWR_M1029_d 0.00532631f $X=1.71 $Y=2.145 $X2=0
+ $Y2=0
cc_973 N_A_27_74#_c_1576_n N_VPWR_c_1641_n 0.0302173f $X=0.28 $Y=2.75 $X2=0
+ $Y2=0
cc_974 N_A_27_74#_c_1577_n N_VPWR_c_1641_n 0.0275301f $X=1.625 $Y=2.275 $X2=0
+ $Y2=0
cc_975 N_A_27_74#_c_1577_n N_VPWR_c_1642_n 0.00106645f $X=1.625 $Y=2.275 $X2=0
+ $Y2=0
cc_976 N_A_27_74#_c_1578_n N_VPWR_c_1642_n 0.00270804f $X=2.445 $Y=2.145 $X2=0
+ $Y2=0
cc_977 N_A_27_74#_c_1623_n N_VPWR_c_1642_n 0.0124964f $X=1.71 $Y=2.145 $X2=0
+ $Y2=0
cc_978 N_A_27_74#_c_1576_n N_VPWR_c_1655_n 0.011066f $X=0.28 $Y=2.75 $X2=0 $Y2=0
cc_979 N_A_27_74#_c_1576_n N_VPWR_c_1640_n 0.00915947f $X=0.28 $Y=2.75 $X2=0
+ $Y2=0
cc_980 N_A_27_74#_c_1570_n N_VGND_c_1853_n 0.0172562f $X=0.28 $Y=0.58 $X2=0
+ $Y2=0
cc_981 N_A_27_74#_c_1570_n N_VGND_c_1864_n 0.0109681f $X=0.28 $Y=0.58 $X2=0
+ $Y2=0
cc_982 N_A_27_74#_c_1570_n N_VGND_c_1878_n 0.00912188f $X=0.28 $Y=0.58 $X2=0
+ $Y2=0
cc_983 N_VPWR_c_1647_n Q_N 0.0870143f $X=10.695 $Y=1.985 $X2=0 $Y2=0
cc_984 N_VPWR_c_1646_n Q_N 0.0131276f $X=9.795 $Y=2.805 $X2=0 $Y2=0
cc_985 N_VPWR_c_1653_n Q_N 0.0128835f $X=10.605 $Y=3.33 $X2=0 $Y2=0
cc_986 N_VPWR_c_1640_n Q_N 0.0109343f $X=12.72 $Y=3.33 $X2=0 $Y2=0
cc_987 N_VPWR_c_1661_n N_Q_c_1824_n 0.0158009f $X=12.595 $Y=3.33 $X2=0 $Y2=0
cc_988 N_VPWR_c_1640_n N_Q_c_1824_n 0.0129424f $X=12.72 $Y=3.33 $X2=0 $Y2=0
cc_989 N_VPWR_c_1648_n N_Q_c_1825_n 0.0783173f $X=11.78 $Y=1.985 $X2=0 $Y2=0
cc_990 N_VPWR_c_1650_n N_Q_c_1825_n 0.0887573f $X=12.68 $Y=1.985 $X2=0 $Y2=0
cc_991 Q_N N_VGND_c_1857_n 0.0182946f $X=10.235 $Y=0.47 $X2=0 $Y2=0
cc_992 Q_N N_VGND_c_1858_n 0.0297335f $X=10.235 $Y=0.47 $X2=0 $Y2=0
cc_993 Q_N N_VGND_c_1862_n 0.0114106f $X=10.235 $Y=0.47 $X2=0 $Y2=0
cc_994 Q_N N_VGND_c_1878_n 0.00936481f $X=10.235 $Y=0.47 $X2=0 $Y2=0
cc_995 Q N_VGND_c_1859_n 0.0263849f $X=12.155 $Y=0.47 $X2=0 $Y2=0
cc_996 Q N_VGND_c_1861_n 0.0308798f $X=12.155 $Y=0.47 $X2=0 $Y2=0
cc_997 Q N_VGND_c_1868_n 0.0149085f $X=12.155 $Y=0.47 $X2=0 $Y2=0
cc_998 Q N_VGND_c_1878_n 0.0122037f $X=12.155 $Y=0.47 $X2=0 $Y2=0
