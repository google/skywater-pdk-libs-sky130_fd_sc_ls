* NGSPICE file created from sky130_fd_sc_ls__o21ba_1.ext - technology: sky130A

.subckt sky130_fd_sc_ls__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
M1000 X a_200_392# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=1.052e+12p ps=8.29e+06u
M1001 VPWR a_281_244# a_200_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=4.2e+11p ps=2.84e+06u
M1002 a_200_392# A2 a_116_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1003 a_200_392# a_281_244# a_27_74# VNB nshort w=640000u l=150000u
+  ad=2.176e+11p pd=1.96e+06u as=3.712e+11p ps=3.72e+06u
M1004 VGND B1_N a_281_244# VNB nshort w=550000u l=150000u
+  ad=5.587e+11p pd=4.44e+06u as=2.75e+11p ps=2.1e+06u
M1005 VPWR B1_N a_281_244# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=3.108e+11p ps=2.42e+06u
M1006 a_116_392# A1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND A1 a_27_74# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_27_74# A2 VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 X a_200_392# VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
.ends

