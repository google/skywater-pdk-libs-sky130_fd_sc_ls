# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ls__sdlclkp_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ls__sdlclkp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.680000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN GATE
    ANTENNAGATEAREA  0.208500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.805000 1.630000 1.285000 2.150000 ;
    END
  END GATE
  PIN GCLK
    ANTENNADIFFAREA  0.632800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.235000 1.820000 7.585000 2.980000 ;
        RECT 7.240000 0.350000 7.585000 1.130000 ;
        RECT 7.415000 1.130000 7.585000 1.820000 ;
    END
  END GCLK
  PIN SCE
    ANTENNAGATEAREA  0.208500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.290000 0.545000 1.960000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.459000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 5.330000 1.355000 5.660000 1.780000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 7.680000 0.085000 ;
        RECT 0.115000  0.085000 0.365000 1.120000 ;
        RECT 1.055000  0.085000 1.385000 0.370000 ;
        RECT 3.750000  0.085000 3.920000 0.710000 ;
        RECT 5.410000  0.085000 5.660000 1.130000 ;
        RECT 6.815000  0.085000 7.065000 1.130000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
        RECT 6.395000 -0.085000 6.565000 0.085000 ;
        RECT 6.875000 -0.085000 7.045000 0.085000 ;
        RECT 7.355000 -0.085000 7.525000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.680000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 7.680000 3.415000 ;
        RECT 0.115000 2.130000 0.445000 3.245000 ;
        RECT 1.515000 2.660000 1.845000 3.245000 ;
        RECT 3.985000 2.440000 4.315000 3.245000 ;
        RECT 5.585000 2.835000 5.990000 3.245000 ;
        RECT 6.695000 2.060000 7.025000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
        RECT 6.395000 3.245000 6.565000 3.415000 ;
        RECT 6.875000 3.245000 7.045000 3.415000 ;
        RECT 7.355000 3.245000 7.525000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 7.680000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.545000 0.540000 2.375000 0.710000 ;
      RECT 0.545000 0.710000 0.885000 1.120000 ;
      RECT 0.715000 1.120000 0.885000 1.290000 ;
      RECT 0.715000 1.290000 1.625000 1.460000 ;
      RECT 0.955000 2.320000 2.860000 2.490000 ;
      RECT 0.955000 2.490000 1.285000 2.980000 ;
      RECT 1.455000 1.460000 1.625000 2.320000 ;
      RECT 1.565000 0.880000 1.895000 0.950000 ;
      RECT 1.565000 0.950000 1.965000 1.120000 ;
      RECT 1.795000 1.120000 1.965000 1.545000 ;
      RECT 1.795000 1.545000 2.900000 1.715000 ;
      RECT 1.795000 1.715000 2.380000 2.150000 ;
      RECT 2.125000 0.350000 2.375000 0.540000 ;
      RECT 2.125000 0.710000 2.375000 0.780000 ;
      RECT 2.135000 1.030000 2.715000 1.200000 ;
      RECT 2.135000 1.200000 2.415000 1.360000 ;
      RECT 2.545000 0.255000 3.580000 0.425000 ;
      RECT 2.545000 0.425000 2.715000 1.030000 ;
      RECT 2.610000 1.885000 2.860000 2.320000 ;
      RECT 2.610000 2.490000 2.860000 2.755000 ;
      RECT 2.625000 1.385000 2.900000 1.545000 ;
      RECT 2.885000 0.595000 3.240000 0.925000 ;
      RECT 3.060000 2.425000 3.390000 2.755000 ;
      RECT 3.070000 0.925000 3.240000 1.220000 ;
      RECT 3.070000 1.220000 4.320000 1.550000 ;
      RECT 3.070000 1.550000 3.390000 2.425000 ;
      RECT 3.410000 0.425000 3.580000 0.880000 ;
      RECT 3.410000 0.880000 4.260000 1.050000 ;
      RECT 3.600000 1.740000 4.820000 2.120000 ;
      RECT 4.090000 0.255000 5.230000 0.425000 ;
      RECT 4.090000 0.425000 4.260000 0.880000 ;
      RECT 4.430000 0.595000 4.680000 1.050000 ;
      RECT 4.490000 1.050000 4.680000 1.740000 ;
      RECT 4.490000 2.120000 4.820000 2.495000 ;
      RECT 4.490000 2.495000 6.000000 2.665000 ;
      RECT 4.490000 2.665000 4.820000 2.900000 ;
      RECT 4.900000 0.425000 5.230000 1.130000 ;
      RECT 4.990000 1.130000 5.160000 1.995000 ;
      RECT 4.990000 1.995000 5.380000 2.325000 ;
      RECT 5.830000 1.220000 6.305000 1.550000 ;
      RECT 5.830000 1.550000 6.000000 2.495000 ;
      RECT 6.165000 0.450000 6.645000 1.050000 ;
      RECT 6.195000 1.720000 6.645000 1.890000 ;
      RECT 6.195000 1.890000 6.525000 2.875000 ;
      RECT 6.475000 1.050000 6.645000 1.300000 ;
      RECT 6.475000 1.300000 7.245000 1.630000 ;
      RECT 6.475000 1.630000 6.645000 1.720000 ;
  END
END sky130_fd_sc_ls__sdlclkp_1
