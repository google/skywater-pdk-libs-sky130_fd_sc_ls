* File: sky130_fd_sc_ls__a21bo_1.pex.spice
* Created: Fri Aug 28 12:50:07 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__A21BO_1%A2 1 2 3 5 9 11 12 16
r32 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=0.405 $X2=0.27 $Y2=0.405
r33 12 16 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=0.27 $Y=0.555
+ $X2=0.27 $Y2=0.405
r34 11 15 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=0.46 $Y=0.405
+ $X2=0.27 $Y2=0.405
r35 9 10 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.535 $Y=1 $X2=0.535
+ $Y2=1.395
r36 6 11 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=0.535 $Y=0.57
+ $X2=0.46 $Y2=0.405
r37 6 9 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=0.535 $Y=0.57
+ $X2=0.535 $Y2=1
r38 3 5 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.52 $Y=1.885
+ $X2=0.52 $Y2=2.46
r39 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.52 $Y=1.795 $X2=0.52
+ $Y2=1.885
r40 1 10 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.52 $Y=1.485 $X2=0.52
+ $Y2=1.395
r41 1 2 120.5 $w=1.8e-07 $l=3.1e-07 $layer=POLY_cond $X=0.52 $Y=1.485 $X2=0.52
+ $Y2=1.795
.ends

.subckt PM_SKY130_FD_SC_LS__A21BO_1%A1 3 5 7 8
c36 5 0 1.15205e-19 $X=1 $Y=1.885
r37 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.985
+ $Y=1.615 $X2=0.985 $Y2=1.615
r38 8 12 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=1.2 $Y=1.615
+ $X2=0.985 $Y2=1.615
r39 5 11 55.8646 $w=2.93e-07 $l=2.77399e-07 $layer=POLY_cond $X=1 $Y=1.885
+ $X2=0.985 $Y2=1.615
r40 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1 $Y=1.885 $X2=1
+ $Y2=2.46
r41 1 11 38.5916 $w=2.93e-07 $l=2.05122e-07 $layer=POLY_cond $X=0.895 $Y=1.45
+ $X2=0.985 $Y2=1.615
r42 1 3 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=0.895 $Y=1.45
+ $X2=0.895 $Y2=1
.ends

.subckt PM_SKY130_FD_SC_LS__A21BO_1%A_272_110# 1 2 7 9 11 12 14 15 17 19 21 22
+ 27 29 34
r66 31 34 8.00764 $w=5.88e-07 $l=3.95e-07 $layer=LI1_cond $X=2.16 $Y=0.645
+ $X2=2.555 $Y2=0.645
r67 25 30 0.0912679 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=2.245 $Y=1.945
+ $X2=2.08 $Y2=1.945
r68 25 27 13.1378 $w=2.48e-07 $l=2.85e-07 $layer=LI1_cond $X=2.245 $Y=1.945
+ $X2=2.53 $Y2=1.945
r69 23 31 8.20854 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=2.16 $Y=0.94
+ $X2=2.16 $Y2=0.645
r70 23 29 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=2.16 $Y=0.94
+ $X2=2.16 $Y2=1.1
r71 22 38 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=2.08 $Y=1.265
+ $X2=2.08 $Y2=1.47
r72 21 29 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.08 $Y=1.265
+ $X2=2.08 $Y2=1.1
r73 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.08
+ $Y=1.265 $X2=2.08 $Y2=1.265
r74 19 30 13.7904 $w=3.3e-07 $l=3.4e-07 $layer=LI1_cond $X=2.08 $Y=1.605
+ $X2=2.08 $Y2=1.945
r75 19 21 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=2.08 $Y=1.605
+ $X2=2.08 $Y2=1.265
r76 16 17 6.66866 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=1.54 $Y=1.47 $X2=1.45
+ $Y2=1.47
r77 15 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.915 $Y=1.47
+ $X2=2.08 $Y2=1.47
r78 15 16 192.287 $w=1.5e-07 $l=3.75e-07 $layer=POLY_cond $X=1.915 $Y=1.47
+ $X2=1.54 $Y2=1.47
r79 12 14 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.45 $Y=1.885
+ $X2=1.45 $Y2=2.46
r80 11 12 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.45 $Y=1.795 $X2=1.45
+ $Y2=1.885
r81 10 17 18.8402 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=1.45 $Y=1.545
+ $X2=1.45 $Y2=1.47
r82 10 11 97.1774 $w=1.8e-07 $l=2.5e-07 $layer=POLY_cond $X=1.45 $Y=1.545
+ $X2=1.45 $Y2=1.795
r83 7 17 18.8402 $w=1.65e-07 $l=8.21584e-08 $layer=POLY_cond $X=1.435 $Y=1.395
+ $X2=1.45 $Y2=1.47
r84 7 9 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.435 $Y=1.395
+ $X2=1.435 $Y2=1
r85 2 27 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=2.405
+ $Y=1.84 $X2=2.53 $Y2=1.985
r86 1 34 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=2.41
+ $Y=0.37 $X2=2.555 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_LS__A21BO_1%B1_N 1 3 6 8
r32 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.68
+ $Y=1.385 $X2=2.68 $Y2=1.385
r33 8 12 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=2.68 $Y=1.295 $X2=2.68
+ $Y2=1.385
r34 4 11 38.9026 $w=2.7e-07 $l=2.05122e-07 $layer=POLY_cond $X=2.77 $Y=1.22
+ $X2=2.68 $Y2=1.385
r35 4 6 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.77 $Y=1.22 $X2=2.77
+ $Y2=0.645
r36 1 11 77.2841 $w=2.7e-07 $l=4.15812e-07 $layer=POLY_cond $X=2.755 $Y=1.765
+ $X2=2.68 $Y2=1.385
r37 1 3 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.755 $Y=1.765
+ $X2=2.755 $Y2=2.26
.ends

.subckt PM_SKY130_FD_SC_LS__A21BO_1%A_194_136# 1 2 9 11 13 16 18 19 22 28 30 33
+ 34 37
c83 34 0 6.82625e-20 $X=1.667 $Y=1.94
c84 33 0 9.10919e-20 $X=3.17 $Y=2.24
c85 11 0 1.9051e-19 $X=3.29 $Y=1.765
r86 37 40 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.25 $Y=1.485
+ $X2=3.25 $Y2=1.65
r87 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.25
+ $Y=1.485 $X2=3.25 $Y2=1.485
r88 33 40 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=3.17 $Y=2.24 $X2=3.17
+ $Y2=1.65
r89 31 35 1.64875 $w=1.7e-07 $l=9.3e-08 $layer=LI1_cond $X=1.76 $Y=2.325
+ $X2=1.667 $Y2=2.325
r90 30 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.085 $Y=2.325
+ $X2=3.17 $Y2=2.24
r91 30 31 86.4438 $w=1.68e-07 $l=1.325e-06 $layer=LI1_cond $X=3.085 $Y=2.325
+ $X2=1.76 $Y2=2.325
r92 26 35 4.81226 $w=1.85e-07 $l=8.5e-08 $layer=LI1_cond $X=1.667 $Y=2.41
+ $X2=1.667 $Y2=2.325
r93 26 28 2.99754 $w=1.83e-07 $l=5e-08 $layer=LI1_cond $X=1.667 $Y=2.41
+ $X2=1.667 $Y2=2.46
r94 23 35 4.81226 $w=1.85e-07 $l=8.5e-08 $layer=LI1_cond $X=1.667 $Y=2.24
+ $X2=1.667 $Y2=2.325
r95 23 25 8.09337 $w=1.83e-07 $l=1.35e-07 $layer=LI1_cond $X=1.667 $Y=2.24
+ $X2=1.667 $Y2=2.105
r96 22 34 5.60801 $w=1.83e-07 $l=9.2e-08 $layer=LI1_cond $X=1.667 $Y=2.032
+ $X2=1.667 $Y2=1.94
r97 22 25 4.37641 $w=1.83e-07 $l=7.3e-08 $layer=LI1_cond $X=1.667 $Y=2.032
+ $X2=1.667 $Y2=2.105
r98 20 34 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=1.66 $Y=1.28
+ $X2=1.66 $Y2=1.94
r99 18 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.575 $Y=1.195
+ $X2=1.66 $Y2=1.28
r100 18 19 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=1.575 $Y=1.195
+ $X2=1.315 $Y2=1.195
r101 14 19 8.10976 $w=1.7e-07 $l=2.23495e-07 $layer=LI1_cond $X=1.13 $Y=1.11
+ $X2=1.315 $Y2=1.195
r102 14 16 9.49987 $w=3.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.13 $Y=1.11
+ $X2=1.13 $Y2=0.805
r103 11 38 57.6553 $w=2.91e-07 $l=2.99333e-07 $layer=POLY_cond $X=3.29 $Y=1.765
+ $X2=3.25 $Y2=1.485
r104 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.29 $Y=1.765
+ $X2=3.29 $Y2=2.4
r105 7 38 38.6072 $w=2.91e-07 $l=1.67481e-07 $layer=POLY_cond $X=3.245 $Y=1.32
+ $X2=3.25 $Y2=1.485
r106 7 9 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.245 $Y=1.32
+ $X2=3.245 $Y2=0.74
r107 2 28 300 $w=1.7e-07 $l=5.70088e-07 $layer=licon1_PDIFF $count=2 $X=1.525
+ $Y=1.96 $X2=1.675 $Y2=2.46
r108 2 25 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.96 $X2=1.675 $Y2=2.105
r109 1 16 91 $w=1.7e-07 $l=2.13542e-07 $layer=licon1_NDIFF $count=2 $X=0.97
+ $Y=0.68 $X2=1.13 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LS__A21BO_1%A_34_392# 1 2 7 9 11 13 15
c30 7 0 4.69421e-20 $X=0.295 $Y=2.12
r31 13 20 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.225 $Y=2.12
+ $X2=1.225 $Y2=2.035
r32 13 15 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=1.225 $Y=2.12
+ $X2=1.225 $Y2=2.815
r33 12 18 5.07788 $w=1.7e-07 $l=1.67481e-07 $layer=LI1_cond $X=0.46 $Y=2.035
+ $X2=0.295 $Y2=2.03
r34 11 20 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.06 $Y=2.035
+ $X2=1.225 $Y2=2.035
r35 11 12 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=1.06 $Y=2.035 $X2=0.46
+ $Y2=2.035
r36 7 18 2.68829 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=0.295 $Y=2.12 $X2=0.295
+ $Y2=2.03
r37 7 9 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=0.295 $Y=2.12
+ $X2=0.295 $Y2=2.815
r38 2 20 400 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=1 $X=1.075
+ $Y=1.96 $X2=1.225 $Y2=2.115
r39 2 15 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=1.075
+ $Y=1.96 $X2=1.225 $Y2=2.815
r40 1 18 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.17
+ $Y=1.96 $X2=0.295 $Y2=2.105
r41 1 9 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.17
+ $Y=1.96 $X2=0.295 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_LS__A21BO_1%VPWR 1 2 11 15 17 19 29 30 33 36
r38 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r39 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r40 30 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r41 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r42 27 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.23 $Y=3.33
+ $X2=3.065 $Y2=3.33
r43 27 29 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.23 $Y=3.33 $X2=3.6
+ $Y2=3.33
r44 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r45 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r46 23 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r47 22 25 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r48 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r49 20 33 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=0.86 $Y=3.33 $X2=0.76
+ $Y2=3.33
r50 20 22 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.86 $Y=3.33 $X2=1.2
+ $Y2=3.33
r51 19 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.9 $Y=3.33
+ $X2=3.065 $Y2=3.33
r52 19 25 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=2.9 $Y=3.33 $X2=2.64
+ $Y2=3.33
r53 17 26 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.64 $Y2=3.33
r54 17 23 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.2 $Y2=3.33
r55 13 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.065 $Y=3.245
+ $X2=3.065 $Y2=3.33
r56 13 15 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=3.065 $Y=3.245
+ $X2=3.065 $Y2=2.745
r57 9 33 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=0.76 $Y=3.245 $X2=0.76
+ $Y2=3.33
r58 9 11 43.8091 $w=1.98e-07 $l=7.9e-07 $layer=LI1_cond $X=0.76 $Y=3.245
+ $X2=0.76 $Y2=2.455
r59 2 15 600 $w=1.7e-07 $l=1.01573e-06 $layer=licon1_PDIFF $count=1 $X=2.83
+ $Y=1.84 $X2=3.065 $Y2=2.745
r60 1 11 300 $w=1.7e-07 $l=5.71577e-07 $layer=licon1_PDIFF $count=2 $X=0.595
+ $Y=1.96 $X2=0.76 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_LS__A21BO_1%X 1 2 9 13 14 15 16 24 33
r25 21 24 0.106379 $w=3.23e-07 $l=3e-09 $layer=LI1_cond $X=3.592 $Y=1.982
+ $X2=3.592 $Y2=1.985
r26 15 16 13.1201 $w=3.23e-07 $l=3.7e-07 $layer=LI1_cond $X=3.592 $Y=2.405
+ $X2=3.592 $Y2=2.775
r27 14 21 0.567357 $w=3.23e-07 $l=1.6e-08 $layer=LI1_cond $X=3.592 $Y=1.966
+ $X2=3.592 $Y2=1.982
r28 14 33 7.78643 $w=3.23e-07 $l=1.46e-07 $layer=LI1_cond $X=3.592 $Y=1.966
+ $X2=3.592 $Y2=1.82
r29 14 15 12.5528 $w=3.23e-07 $l=3.54e-07 $layer=LI1_cond $X=3.592 $Y=2.051
+ $X2=3.592 $Y2=2.405
r30 14 24 2.34035 $w=3.23e-07 $l=6.6e-08 $layer=LI1_cond $X=3.592 $Y=2.051
+ $X2=3.592 $Y2=1.985
r31 13 33 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.67 $Y=1.13 $X2=3.67
+ $Y2=1.82
r32 7 13 10.9702 $w=4.58e-07 $l=2.3e-07 $layer=LI1_cond $X=3.525 $Y=0.9
+ $X2=3.525 $Y2=1.13
r33 7 9 10.0107 $w=4.58e-07 $l=3.85e-07 $layer=LI1_cond $X=3.525 $Y=0.9
+ $X2=3.525 $Y2=0.515
r34 2 16 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=3.365
+ $Y=1.84 $X2=3.515 $Y2=2.815
r35 2 24 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=3.365
+ $Y=1.84 $X2=3.515 $Y2=1.985
r36 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.32
+ $Y=0.37 $X2=3.46 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__A21BO_1%VGND 1 2 3 11 14 18 21 24 25 27 28 29 35 44
+ 45 48
c59 18 0 1.9051e-19 $X=3.005 $Y=0.665
r60 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r61 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r62 42 45 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r63 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r64 39 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.815 $Y=0 $X2=1.65
+ $Y2=0
r65 39 41 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=1.815 $Y=0 $X2=2.64
+ $Y2=0
r66 38 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r67 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r68 35 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.485 $Y=0 $X2=1.65
+ $Y2=0
r69 35 37 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.485 $Y=0 $X2=1.2
+ $Y2=0
r70 33 38 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r71 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r72 29 42 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.64
+ $Y2=0
r73 29 49 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r74 27 41 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=2.9 $Y=0 $X2=2.64
+ $Y2=0
r75 27 28 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=2.9 $Y=0 $X2=3.007
+ $Y2=0
r76 26 44 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=3.115 $Y=0 $X2=3.6
+ $Y2=0
r77 26 28 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=3.115 $Y=0 $X2=3.007
+ $Y2=0
r78 24 32 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.605 $Y=0 $X2=0.24
+ $Y2=0
r79 24 25 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=0 $X2=0.69
+ $Y2=0
r80 23 37 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=0.775 $Y=0 $X2=1.2
+ $Y2=0
r81 23 25 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=0 $X2=0.69
+ $Y2=0
r82 21 22 11.7247 $w=3.85e-07 $l=3.7e-07 $layer=LI1_cond $X=0.32 $Y=1.09
+ $X2=0.69 $Y2=1.09
r83 16 28 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=3.007 $Y=0.085
+ $X2=3.007 $Y2=0
r84 16 18 31.0892 $w=2.13e-07 $l=5.8e-07 $layer=LI1_cond $X=3.007 $Y=0.085
+ $X2=3.007 $Y2=0.665
r85 12 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.65 $Y=0.085
+ $X2=1.65 $Y2=0
r86 12 14 26.1919 $w=3.28e-07 $l=7.5e-07 $layer=LI1_cond $X=1.65 $Y=0.085
+ $X2=1.65 $Y2=0.835
r87 11 22 5.54671 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=0.69 $Y=0.84 $X2=0.69
+ $Y2=1.09
r88 10 25 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=0.085
+ $X2=0.69 $Y2=0
r89 10 11 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=0.69 $Y=0.085
+ $X2=0.69 $Y2=0.84
r90 3 18 182 $w=1.7e-07 $l=3.66367e-07 $layer=licon1_NDIFF $count=1 $X=2.845
+ $Y=0.37 $X2=3.005 $Y2=0.665
r91 2 14 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=1.51
+ $Y=0.68 $X2=1.65 $Y2=0.835
r92 1 21 182 $w=1.7e-07 $l=4.68348e-07 $layer=licon1_NDIFF $count=1 $X=0.195
+ $Y=0.68 $X2=0.32 $Y2=1.09
.ends

