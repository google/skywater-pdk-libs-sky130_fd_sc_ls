* File: sky130_fd_sc_ls__mux4_2.pex.spice
* Created: Wed Sep  2 11:10:59 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__MUX4_2%S0 3 5 6 8 11 13 15 18 19 21 23 24 25 27 30
+ 33 35 39 43 46 47 48 52 54 58 60 67
c163 67 0 9.37441e-20 $X=4.56 $Y=1.22
c164 58 0 1.77444e-19 $X=0.6 $Y=1.385
c165 52 0 4.5023e-20 $X=4.56 $Y=1.385
c166 48 0 2.33726e-19 $X=4.56 $Y=1.195
c167 43 0 1.72582e-19 $X=1.485 $Y=1.195
c168 30 0 1.35612e-19 $X=2.94 $Y=1.615
c169 13 0 2.52602e-19 $X=3.015 $Y=1.885
r170 58 61 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.6 $Y=1.385
+ $X2=0.6 $Y2=1.55
r171 58 60 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.6 $Y=1.385
+ $X2=0.6 $Y2=1.22
r172 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.6
+ $Y=1.385 $X2=0.6 $Y2=1.385
r173 54 59 3.24852 $w=3.38e-07 $l=9e-08 $layer=LI1_cond $X=0.62 $Y=1.295
+ $X2=0.62 $Y2=1.385
r174 54 72 3.60947 $w=3.38e-07 $l=1e-07 $layer=LI1_cond $X=0.62 $Y=1.295
+ $X2=0.62 $Y2=1.195
r175 54 72 4.76605 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=0.805 $Y=1.195
+ $X2=0.62 $Y2=1.195
r176 52 67 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.56 $Y=1.385
+ $X2=4.56 $Y2=1.22
r177 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.56
+ $Y=1.385 $X2=4.56 $Y2=1.385
r178 48 51 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=4.56 $Y=1.195
+ $X2=4.56 $Y2=1.385
r179 46 63 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.68 $Y=1.425
+ $X2=1.68 $Y2=1.26
r180 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.68
+ $Y=1.425 $X2=1.68 $Y2=1.425
r181 43 54 33.6483 $w=2.38e-07 $l=6.8e-07 $layer=LI1_cond $X=1.485 $Y=1.195
+ $X2=0.805 $Y2=1.195
r182 43 45 9.35333 $w=3e-07 $l=3.07083e-07 $layer=LI1_cond $X=1.485 $Y=1.195
+ $X2=1.665 $Y2=1.425
r183 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.64
+ $Y=1.585 $X2=5.64 $Y2=1.585
r184 37 39 13.0183 $w=2.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.61 $Y=1.28
+ $X2=5.61 $Y2=1.585
r185 36 48 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.725 $Y=1.195
+ $X2=4.56 $Y2=1.195
r186 35 37 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=5.475 $Y=1.195
+ $X2=5.61 $Y2=1.28
r187 35 36 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=5.475 $Y=1.195
+ $X2=4.725 $Y2=1.195
r188 34 47 3.05049 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.105 $Y=1.195
+ $X2=2.97 $Y2=1.195
r189 33 48 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.395 $Y=1.195
+ $X2=4.56 $Y2=1.195
r190 33 34 84.1604 $w=1.68e-07 $l=1.29e-06 $layer=LI1_cond $X=4.395 $Y=1.195
+ $X2=3.105 $Y2=1.195
r191 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.94
+ $Y=1.615 $X2=2.94 $Y2=1.615
r192 28 47 3.46198 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.97 $Y=1.28
+ $X2=2.97 $Y2=1.195
r193 28 30 14.2988 $w=2.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.97 $Y=1.28
+ $X2=2.97 $Y2=1.615
r194 27 47 3.46198 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.97 $Y=1.11
+ $X2=2.97 $Y2=1.195
r195 26 27 22.1952 $w=2.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.97 $Y=0.59
+ $X2=2.97 $Y2=1.11
r196 24 26 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=2.835 $Y=0.505
+ $X2=2.97 $Y2=0.59
r197 24 25 76.984 $w=1.68e-07 $l=1.18e-06 $layer=LI1_cond $X=2.835 $Y=0.505
+ $X2=1.655 $Y2=0.505
r198 23 43 5.72868 $w=3e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.57 $Y=1.11
+ $X2=1.485 $Y2=1.195
r199 22 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.57 $Y=0.59
+ $X2=1.655 $Y2=0.505
r200 22 23 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.57 $Y=0.59
+ $X2=1.57 $Y2=1.11
r201 19 40 61.4066 $w=2.86e-07 $l=3.21714e-07 $layer=POLY_cond $X=5.685 $Y=1.885
+ $X2=5.64 $Y2=1.585
r202 19 21 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.685 $Y=1.885
+ $X2=5.685 $Y2=2.46
r203 18 67 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.47 $Y=0.74
+ $X2=4.47 $Y2=1.22
r204 13 31 55.8646 $w=2.93e-07 $l=3.05205e-07 $layer=POLY_cond $X=3.015 $Y=1.885
+ $X2=2.94 $Y2=1.615
r205 13 15 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.015 $Y=1.885
+ $X2=3.015 $Y2=2.46
r206 11 63 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=1.59 $Y=0.74
+ $X2=1.59 $Y2=1.26
r207 6 8 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.645 $Y=1.885
+ $X2=0.645 $Y2=2.46
r208 5 6 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.645 $Y=1.795
+ $X2=0.645 $Y2=1.885
r209 5 61 95.2339 $w=1.8e-07 $l=2.45e-07 $layer=POLY_cond $X=0.645 $Y=1.795
+ $X2=0.645 $Y2=1.55
r210 3 60 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=0.515 $Y=0.79
+ $X2=0.515 $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_LS__MUX4_2%A1 3 5 7 8
c31 8 0 1.14029e-19 $X=1.2 $Y=1.665
r32 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.14
+ $Y=1.615 $X2=1.14 $Y2=1.615
r33 5 11 55.6066 $w=2.97e-07 $l=3.11769e-07 $layer=POLY_cond $X=1.245 $Y=1.885
+ $X2=1.155 $Y2=1.615
r34 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.245 $Y=1.885
+ $X2=1.245 $Y2=2.46
r35 1 11 38.5662 $w=2.97e-07 $l=1.86145e-07 $layer=POLY_cond $X=1.2 $Y=1.45
+ $X2=1.155 $Y2=1.615
r36 1 3 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.2 $Y=1.45 $X2=1.2
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__MUX4_2%A_31_94# 1 2 7 9 12 14 16 19 25 28 31 32 33
+ 34 37 43 48 51 61
c120 48 0 1.66876e-19 $X=2.22 $Y=1.615
c121 33 0 4.5023e-20 $X=4.895 $Y=2.035
c122 14 0 1.11429e-19 $X=4.995 $Y=1.885
c123 7 0 3.08193e-19 $X=2.295 $Y=1.885
r124 63 64 2.37898 $w=4.88e-07 $l=4.5e-08 $layer=LI1_cond $X=0.34 $Y=2.105
+ $X2=0.34 $Y2=2.15
r125 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.1
+ $Y=1.625 $X2=5.1 $Y2=1.625
r126 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.22
+ $Y=1.615 $X2=2.22 $Y2=1.615
r127 44 51 13.8971 $w=3.38e-07 $l=4.1e-07 $layer=LI1_cond $X=5.095 $Y=2.035
+ $X2=5.095 $Y2=1.625
r128 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=2.035
+ $X2=5.04 $Y2=2.035
r129 41 48 17.2866 $w=2.78e-07 $l=4.2e-07 $layer=LI1_cond $X=2.185 $Y=2.035
+ $X2=2.185 $Y2=1.615
r130 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=2.035
+ $X2=2.16 $Y2=2.035
r131 37 63 1.70868 $w=4.88e-07 $l=7e-08 $layer=LI1_cond $X=0.34 $Y=2.035
+ $X2=0.34 $Y2=2.105
r132 37 61 8.23575 $w=4.88e-07 $l=1.15e-07 $layer=LI1_cond $X=0.34 $Y=2.035
+ $X2=0.34 $Y2=1.92
r133 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=2.035
+ $X2=0.24 $Y2=2.035
r134 34 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.305 $Y=2.035
+ $X2=2.16 $Y2=2.035
r135 33 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.895 $Y=2.035
+ $X2=5.04 $Y2=2.035
r136 33 34 3.20544 $w=1.4e-07 $l=2.59e-06 $layer=MET1_cond $X=4.895 $Y=2.035
+ $X2=2.305 $Y2=2.035
r137 32 36 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.385 $Y=2.035
+ $X2=0.24 $Y2=2.035
r138 31 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.015 $Y=2.035
+ $X2=2.16 $Y2=2.035
r139 31 32 2.01732 $w=1.4e-07 $l=1.63e-06 $layer=MET1_cond $X=2.015 $Y=2.035
+ $X2=0.385 $Y2=2.035
r140 30 61 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=0.18 $Y=1.01
+ $X2=0.18 $Y2=1.92
r141 28 30 11.4978 $w=3.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.28 $Y=0.75
+ $X2=0.28 $Y2=1.01
r142 25 64 23.2235 $w=3.28e-07 $l=6.65e-07 $layer=LI1_cond $X=0.42 $Y=2.815
+ $X2=0.42 $Y2=2.15
r143 17 50 38.5916 $w=2.93e-07 $l=1.96074e-07 $layer=POLY_cond $X=5.16 $Y=1.46
+ $X2=5.092 $Y2=1.625
r144 17 19 369.191 $w=1.5e-07 $l=7.2e-07 $layer=POLY_cond $X=5.16 $Y=1.46
+ $X2=5.16 $Y2=0.74
r145 14 50 54.2196 $w=2.93e-07 $l=3.04664e-07 $layer=POLY_cond $X=4.995 $Y=1.885
+ $X2=5.092 $Y2=1.625
r146 14 16 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=4.995 $Y=1.885
+ $X2=4.995 $Y2=2.46
r147 10 47 38.7288 $w=3.45e-07 $l=2.33345e-07 $layer=POLY_cond $X=2.46 $Y=1.45
+ $X2=2.295 $Y2=1.615
r148 10 12 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=2.46 $Y=1.45
+ $X2=2.46 $Y2=0.74
r149 7 47 53.3984 $w=3.45e-07 $l=2.7e-07 $layer=POLY_cond $X=2.295 $Y=1.885
+ $X2=2.295 $Y2=1.615
r150 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.295 $Y=1.885
+ $X2=2.295 $Y2=2.46
r151 2 63 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.275
+ $Y=1.96 $X2=0.42 $Y2=2.105
r152 2 25 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.275
+ $Y=1.96 $X2=0.42 $Y2=2.815
r153 1 28 182 $w=1.7e-07 $l=3.44964e-07 $layer=licon1_NDIFF $count=1 $X=0.155
+ $Y=0.47 $X2=0.3 $Y2=0.75
.ends

.subckt PM_SKY130_FD_SC_LS__MUX4_2%A0 3 5 6 7 9 11
c39 5 0 1.72518e-19 $X=3.48 $Y=1.405
r40 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.48
+ $Y=1.615 $X2=3.48 $Y2=1.615
r41 11 15 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=3.6 $Y=1.615 $X2=3.48
+ $Y2=1.615
r42 7 14 57.5577 $w=2.71e-07 $l=2.91633e-07 $layer=POLY_cond $X=3.435 $Y=1.885
+ $X2=3.48 $Y2=1.615
r43 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.435 $Y=1.885
+ $X2=3.435 $Y2=2.46
r44 6 14 1.68328 $w=3.3e-07 $l=8.75758e-08 $layer=POLY_cond $X=3.48 $Y=1.615
+ $X2=3.48 $Y2=1.615
r45 5 10 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.48 $Y=1.405
+ $X2=3.48 $Y2=1.24
r46 5 6 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=3.48 $Y=1.405 $X2=3.48
+ $Y2=1.615
r47 3 10 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=3.39 $Y=0.74 $X2=3.39
+ $Y2=1.24
.ends

.subckt PM_SKY130_FD_SC_LS__MUX4_2%A3 3 5 7 8
c34 5 0 1.22296e-19 $X=4.125 $Y=1.885
r35 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.02
+ $Y=1.615 $X2=4.02 $Y2=1.615
r36 5 11 56.1368 $w=2.89e-07 $l=3.15214e-07 $layer=POLY_cond $X=4.125 $Y=1.885
+ $X2=4.027 $Y2=1.615
r37 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=4.125 $Y=1.885
+ $X2=4.125 $Y2=2.46
r38 1 11 38.6247 $w=2.89e-07 $l=1.89658e-07 $layer=POLY_cond $X=4.08 $Y=1.45
+ $X2=4.027 $Y2=1.615
r39 1 3 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=4.08 $Y=1.45 $X2=4.08
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__MUX4_2%A2 3 5 6 8 9 10 14 16
r44 14 17 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.18 $Y=1.385
+ $X2=6.18 $Y2=1.55
r45 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.18 $Y=1.385
+ $X2=6.18 $Y2=1.22
r46 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.18
+ $Y=1.385 $X2=6.18 $Y2=1.385
r47 10 15 7.50428 $w=4.28e-07 $l=2.8e-07 $layer=LI1_cond $X=6.13 $Y=1.665
+ $X2=6.13 $Y2=1.385
r48 9 15 2.41209 $w=4.28e-07 $l=9e-08 $layer=LI1_cond $X=6.13 $Y=1.295 $X2=6.13
+ $Y2=1.385
r49 6 8 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.105 $Y=1.885
+ $X2=6.105 $Y2=2.46
r50 5 6 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.105 $Y=1.795 $X2=6.105
+ $Y2=1.885
r51 5 17 95.2339 $w=1.8e-07 $l=2.45e-07 $layer=POLY_cond $X=6.105 $Y=1.795
+ $X2=6.105 $Y2=1.55
r52 3 16 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=6.09 $Y=0.74 $X2=6.09
+ $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_LS__MUX4_2%A_1500_94# 1 2 7 9 10 12 14 19 23 26 27
c54 26 0 1.84046e-19 $X=8.23 $Y=1.615
r55 26 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.23
+ $Y=1.615 $X2=8.23 $Y2=1.615
r56 21 26 6.31733 $w=2.57e-07 $l=1.68953e-07 $layer=LI1_cond $X=8.325 $Y=1.78
+ $X2=8.317 $Y2=1.615
r57 21 23 17.2866 $w=2.48e-07 $l=3.75e-07 $layer=LI1_cond $X=8.325 $Y=1.78
+ $X2=8.325 $Y2=2.155
r58 17 26 6.31733 $w=2.57e-07 $l=1.65e-07 $layer=LI1_cond $X=8.317 $Y=1.45
+ $X2=8.317 $Y2=1.615
r59 17 19 15.2209 $w=2.63e-07 $l=3.5e-07 $layer=LI1_cond $X=8.317 $Y=1.45
+ $X2=8.317 $Y2=1.1
r60 13 27 96.1737 $w=3.3e-07 $l=5.5e-07 $layer=POLY_cond $X=7.68 $Y=1.615
+ $X2=8.23 $Y2=1.615
r61 13 14 5.03009 $w=3.3e-07 $l=1.13049e-07 $layer=POLY_cond $X=7.68 $Y=1.615
+ $X2=7.59 $Y2=1.667
r62 10 14 37.0704 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=7.59 $Y=1.885
+ $X2=7.59 $Y2=1.667
r63 10 12 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=7.59 $Y=1.885
+ $X2=7.59 $Y2=2.46
r64 7 14 37.0704 $w=1.5e-07 $l=2.24375e-07 $layer=POLY_cond $X=7.575 $Y=1.45
+ $X2=7.59 $Y2=1.667
r65 7 9 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=7.575 $Y=1.45 $X2=7.575
+ $Y2=0.97
r66 2 23 600 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_PDIFF $count=1 $X=8.225
+ $Y=1.94 $X2=8.365 $Y2=2.155
r67 1 19 182 $w=1.7e-07 $l=5.70088e-07 $layer=licon1_NDIFF $count=1 $X=8.205
+ $Y=0.6 $X2=8.355 $Y2=1.1
.ends

.subckt PM_SKY130_FD_SC_LS__MUX4_2%S1 4 5 7 8 9 13 14 15 16 18 20
c78 5 0 2.55801e-19 $X=7.14 $Y=1.885
r79 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.065
+ $Y=1.615 $X2=7.065 $Y2=1.615
r80 20 24 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=7.44 $Y=1.615
+ $X2=7.065 $Y2=1.615
r81 16 18 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=8.725 $Y=1.865
+ $X2=8.725 $Y2=2.44
r82 15 16 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=8.725 $Y=1.775
+ $X2=8.725 $Y2=1.865
r83 14 19 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=8.725 $Y=1.405
+ $X2=8.725 $Y2=1.315
r84 14 15 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=8.725 $Y=1.405
+ $X2=8.725 $Y2=1.775
r85 13 19 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=8.71 $Y=0.92
+ $X2=8.71 $Y2=1.315
r86 10 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.71 $Y=0.26
+ $X2=8.71 $Y2=0.92
r87 8 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.635 $Y=0.185
+ $X2=8.71 $Y2=0.26
r88 8 9 764.021 $w=1.5e-07 $l=1.49e-06 $layer=POLY_cond $X=8.635 $Y=0.185
+ $X2=7.145 $Y2=0.185
r89 5 23 55.8646 $w=2.93e-07 $l=3.05205e-07 $layer=POLY_cond $X=7.14 $Y=1.885
+ $X2=7.065 $Y2=1.615
r90 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=7.14 $Y=1.885
+ $X2=7.14 $Y2=2.46
r91 2 23 38.5916 $w=2.93e-07 $l=1.67481e-07 $layer=POLY_cond $X=7.07 $Y=1.45
+ $X2=7.065 $Y2=1.615
r92 2 4 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=7.07 $Y=1.45 $X2=7.07
+ $Y2=0.74
r93 1 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.07 $Y=0.26
+ $X2=7.145 $Y2=0.185
r94 1 4 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=7.07 $Y=0.26 $X2=7.07
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__MUX4_2%A_1429_74# 1 2 7 9 10 12 13 15 16 18 19 22 24
+ 26 29 31 32 38 45
c104 26 0 7.17547e-20 $X=8.96 $Y=2.99
r105 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.22
+ $Y=1.515 $X2=9.22 $Y2=1.515
r106 42 45 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=9.045 $Y=1.515
+ $X2=9.22 $Y2=1.515
r107 38 40 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=7.365 $Y=2.805
+ $X2=7.365 $Y2=2.99
r108 32 35 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=7.285 $Y=0.34
+ $X2=7.285 $Y2=0.515
r109 30 42 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.045 $Y=1.68
+ $X2=9.045 $Y2=1.515
r110 30 31 79.9198 $w=1.68e-07 $l=1.225e-06 $layer=LI1_cond $X=9.045 $Y=1.68
+ $X2=9.045 $Y2=2.905
r111 29 42 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.045 $Y=1.35
+ $X2=9.045 $Y2=1.515
r112 28 29 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=9.045 $Y=0.425
+ $X2=9.045 $Y2=1.35
r113 27 40 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.53 $Y=2.99
+ $X2=7.365 $Y2=2.99
r114 26 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.96 $Y=2.99
+ $X2=9.045 $Y2=2.905
r115 26 27 93.2941 $w=1.68e-07 $l=1.43e-06 $layer=LI1_cond $X=8.96 $Y=2.99
+ $X2=7.53 $Y2=2.99
r116 25 32 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.45 $Y=0.34
+ $X2=7.285 $Y2=0.34
r117 24 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.96 $Y=0.34
+ $X2=9.045 $Y2=0.425
r118 24 25 98.5134 $w=1.68e-07 $l=1.51e-06 $layer=LI1_cond $X=8.96 $Y=0.34
+ $X2=7.45 $Y2=0.34
r119 22 23 4.07324 $w=3.55e-07 $l=3e-08 $layer=POLY_cond $X=10.03 $Y=1.557
+ $X2=10.06 $Y2=1.557
r120 21 22 57.0254 $w=3.55e-07 $l=4.2e-07 $layer=POLY_cond $X=9.61 $Y=1.557
+ $X2=10.03 $Y2=1.557
r121 20 21 1.35775 $w=3.55e-07 $l=1e-08 $layer=POLY_cond $X=9.6 $Y=1.557
+ $X2=9.61 $Y2=1.557
r122 19 46 52.4584 $w=3.3e-07 $l=3e-07 $layer=POLY_cond $X=9.52 $Y=1.515
+ $X2=9.22 $Y2=1.515
r123 19 20 11.1738 $w=3.55e-07 $l=9.87927e-08 $layer=POLY_cond $X=9.52 $Y=1.515
+ $X2=9.6 $Y2=1.557
r124 16 23 22.9692 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=10.06 $Y=1.765
+ $X2=10.06 $Y2=1.557
r125 16 18 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=10.06 $Y=1.765
+ $X2=10.06 $Y2=2.4
r126 13 22 22.9692 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=10.03 $Y=1.35
+ $X2=10.03 $Y2=1.557
r127 13 15 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=10.03 $Y=1.35
+ $X2=10.03 $Y2=0.87
r128 10 21 22.9692 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=9.61 $Y=1.765
+ $X2=9.61 $Y2=1.557
r129 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=9.61 $Y=1.765
+ $X2=9.61 $Y2=2.4
r130 7 20 22.9692 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=9.6 $Y=1.35 $X2=9.6
+ $Y2=1.557
r131 7 9 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=9.6 $Y=1.35 $X2=9.6
+ $Y2=0.87
r132 2 38 600 $w=1.7e-07 $l=9.16938e-07 $layer=licon1_PDIFF $count=1 $X=7.215
+ $Y=1.96 $X2=7.365 $Y2=2.805
r133 1 35 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=7.145
+ $Y=0.37 $X2=7.285 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__MUX4_2%VPWR 1 2 3 4 5 18 24 28 30 34 38 40 45 46 48
+ 49 50 62 69 75 78 82
c98 18 0 6.34146e-20 $X=0.92 $Y=2.115
r99 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r100 78 79 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r101 76 79 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=9.36 $Y2=3.33
r102 75 76 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r103 73 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=10.32 $Y2=3.33
r104 73 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=9.36 $Y2=3.33
r105 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r106 70 78 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.47 $Y=3.33
+ $X2=9.385 $Y2=3.33
r107 70 72 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=9.47 $Y=3.33
+ $X2=9.84 $Y2=3.33
r108 69 81 4.01803 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=10.2 $Y=3.33
+ $X2=10.38 $Y2=3.33
r109 69 72 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=10.2 $Y=3.33
+ $X2=9.84 $Y2=3.33
r110 68 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r111 67 68 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r112 64 67 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.08 $Y=3.33 $X2=6
+ $Y2=3.33
r113 64 65 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r114 62 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.165 $Y=3.33
+ $X2=6.33 $Y2=3.33
r115 62 67 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=6.165 $Y=3.33
+ $X2=6 $Y2=3.33
r116 61 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r117 60 61 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r118 58 61 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=3.6 $Y2=3.33
r119 57 60 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=3.6
+ $Y2=3.33
r120 57 58 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r121 54 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r122 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r123 50 68 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=5.28 $Y=3.33 $X2=6
+ $Y2=3.33
r124 50 65 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=5.28 $Y=3.33
+ $X2=4.08 $Y2=3.33
r125 48 60 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=3.615 $Y=3.33
+ $X2=3.6 $Y2=3.33
r126 48 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.615 $Y=3.33
+ $X2=3.78 $Y2=3.33
r127 47 64 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=3.945 $Y=3.33
+ $X2=4.08 $Y2=3.33
r128 47 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.945 $Y=3.33
+ $X2=3.78 $Y2=3.33
r129 45 53 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=0.755 $Y=3.33
+ $X2=0.72 $Y2=3.33
r130 45 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.755 $Y=3.33
+ $X2=0.92 $Y2=3.33
r131 44 57 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=1.085 $Y=3.33
+ $X2=1.2 $Y2=3.33
r132 44 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.085 $Y=3.33
+ $X2=0.92 $Y2=3.33
r133 40 43 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=10.325 $Y=1.985
+ $X2=10.325 $Y2=2.815
r134 38 81 3.12513 $w=2.5e-07 $l=1.09087e-07 $layer=LI1_cond $X=10.325 $Y=3.245
+ $X2=10.38 $Y2=3.33
r135 38 43 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=10.325 $Y=3.245
+ $X2=10.325 $Y2=2.815
r136 34 37 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=9.385 $Y=2.015
+ $X2=9.385 $Y2=2.795
r137 32 78 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.385 $Y=3.245
+ $X2=9.385 $Y2=3.33
r138 32 37 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=9.385 $Y=3.245
+ $X2=9.385 $Y2=2.795
r139 31 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.495 $Y=3.33
+ $X2=6.33 $Y2=3.33
r140 30 78 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.3 $Y=3.33
+ $X2=9.385 $Y2=3.33
r141 30 31 183 $w=1.68e-07 $l=2.805e-06 $layer=LI1_cond $X=9.3 $Y=3.33 $X2=6.495
+ $Y2=3.33
r142 26 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.33 $Y=3.245
+ $X2=6.33 $Y2=3.33
r143 26 28 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=6.33 $Y=3.245
+ $X2=6.33 $Y2=2.805
r144 22 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.78 $Y=3.245
+ $X2=3.78 $Y2=3.33
r145 22 24 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=3.78 $Y=3.245
+ $X2=3.78 $Y2=2.455
r146 18 21 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=0.92 $Y=2.115
+ $X2=0.92 $Y2=2.815
r147 16 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.92 $Y=3.245
+ $X2=0.92 $Y2=3.33
r148 16 21 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.92 $Y=3.245
+ $X2=0.92 $Y2=2.815
r149 5 43 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=10.135
+ $Y=1.84 $X2=10.285 $Y2=2.815
r150 5 40 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=10.135
+ $Y=1.84 $X2=10.285 $Y2=1.985
r151 4 37 400 $w=1.7e-07 $l=1.10959e-06 $layer=licon1_PDIFF $count=1 $X=8.8
+ $Y=1.94 $X2=9.385 $Y2=2.795
r152 4 34 400 $w=1.7e-07 $l=6.21369e-07 $layer=licon1_PDIFF $count=1 $X=8.8
+ $Y=1.94 $X2=9.385 $Y2=2.015
r153 3 28 600 $w=1.7e-07 $l=9.16938e-07 $layer=licon1_PDIFF $count=1 $X=6.18
+ $Y=1.96 $X2=6.33 $Y2=2.805
r154 2 24 300 $w=1.7e-07 $l=6.15366e-07 $layer=licon1_PDIFF $count=2 $X=3.51
+ $Y=1.96 $X2=3.78 $Y2=2.455
r155 1 21 400 $w=1.7e-07 $l=9.4975e-07 $layer=licon1_PDIFF $count=1 $X=0.72
+ $Y=1.96 $X2=0.92 $Y2=2.815
r156 1 18 400 $w=1.7e-07 $l=2.66458e-07 $layer=licon1_PDIFF $count=1 $X=0.72
+ $Y=1.96 $X2=0.92 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_LS__MUX4_2%A_333_74# 1 2 3 4 13 19 22 23 24 25 26 28 29
+ 31 35 37 38 48
c126 38 0 3.59869e-19 $X=2.97 $Y=1.95
c127 29 0 1.65994e-19 $X=6.73 $Y=1.195
c128 19 0 8.57259e-20 $X=4.115 $Y=2.035
r129 40 42 8.98947 $w=9.48e-07 $l=7e-07 $layer=LI1_cond $X=2.97 $Y=2.115
+ $X2=2.97 $Y2=2.815
r130 37 40 1.02737 $w=9.48e-07 $l=8e-08 $layer=LI1_cond $X=2.97 $Y=2.035
+ $X2=2.97 $Y2=2.115
r131 37 38 11.5385 $w=9.48e-07 $l=8.5e-08 $layer=LI1_cond $X=2.97 $Y=2.035
+ $X2=2.97 $Y2=1.95
r132 33 48 3.77418 $w=2.45e-07 $l=8.5e-08 $layer=LI1_cond $X=6.73 $Y=2.075
+ $X2=6.645 $Y2=2.075
r133 33 35 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=6.73 $Y=2.075
+ $X2=6.9 $Y2=2.075
r134 29 31 69.1551 $w=1.68e-07 $l=1.06e-06 $layer=LI1_cond $X=6.73 $Y=1.195
+ $X2=7.79 $Y2=1.195
r135 28 48 2.68609 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.645 $Y=1.95
+ $X2=6.645 $Y2=2.075
r136 27 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.645 $Y=1.28
+ $X2=6.73 $Y2=1.195
r137 27 28 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.645 $Y=1.28
+ $X2=6.645 $Y2=1.95
r138 26 46 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=5.52 $Y=2.08
+ $X2=5.52 $Y2=2.405
r139 25 48 3.77418 $w=2.45e-07 $l=8.74643e-08 $layer=LI1_cond $X=6.56 $Y=2.08
+ $X2=6.645 $Y2=2.075
r140 25 26 45.8576 $w=2.38e-07 $l=9.55e-07 $layer=LI1_cond $X=6.56 $Y=2.08
+ $X2=5.605 $Y2=2.08
r141 23 46 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.435 $Y=2.405
+ $X2=5.52 $Y2=2.405
r142 23 24 75.0267 $w=1.68e-07 $l=1.15e-06 $layer=LI1_cond $X=5.435 $Y=2.405
+ $X2=4.285 $Y2=2.405
r143 22 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.2 $Y=2.32
+ $X2=4.285 $Y2=2.405
r144 21 22 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=4.2 $Y=2.12 $X2=4.2
+ $Y2=2.32
r145 20 37 11.3727 $w=1.7e-07 $l=4.75e-07 $layer=LI1_cond $X=3.445 $Y=2.035
+ $X2=2.97 $Y2=2.035
r146 19 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.115 $Y=2.035
+ $X2=4.2 $Y2=2.12
r147 19 20 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.115 $Y=2.035
+ $X2=3.445 $Y2=2.035
r148 17 38 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=2.58 $Y=1.09
+ $X2=2.58 $Y2=1.95
r149 13 17 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.495 $Y=0.925
+ $X2=2.58 $Y2=1.09
r150 13 15 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=2.495 $Y=0.925
+ $X2=2.08 $Y2=0.925
r151 4 35 600 $w=1.7e-07 $l=2.19203e-07 $layer=licon1_PDIFF $count=1 $X=6.745
+ $Y=1.96 $X2=6.9 $Y2=2.115
r152 3 42 400 $w=1.7e-07 $l=9.89432e-07 $layer=licon1_PDIFF $count=1 $X=2.37
+ $Y=1.96 $X2=2.66 $Y2=2.815
r153 3 40 400 $w=1.7e-07 $l=3.59235e-07 $layer=licon1_PDIFF $count=1 $X=2.37
+ $Y=1.96 $X2=2.66 $Y2=2.115
r154 2 31 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=7.65
+ $Y=0.6 $X2=7.79 $Y2=1.195
r155 1 15 182 $w=1.7e-07 $l=7.33723e-07 $layer=licon1_NDIFF $count=1 $X=1.665
+ $Y=0.37 $X2=2.08 $Y2=0.925
.ends

.subckt PM_SKY130_FD_SC_LS__MUX4_2%A_909_74# 1 2 3 4 13 17 19 23 25 29 31 33 36
+ 38 42 47 48 50
c130 17 0 9.37441e-20 $X=6.69 $Y=0.855
c131 2 0 1.65994e-19 $X=6.715 $Y=0.37
r132 50 52 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=7.93 $Y=0.68
+ $X2=7.93 $Y2=0.855
r133 48 49 9.75 $w=2.44e-07 $l=1.95e-07 $layer=LI1_cond $X=7.815 $Y=2.455
+ $X2=7.815 $Y2=2.65
r134 38 40 7.07246 $w=5.73e-07 $l=3.4e-07 $layer=LI1_cond $X=4.817 $Y=0.515
+ $X2=4.817 $Y2=0.855
r135 35 36 117.433 $w=1.68e-07 $l=1.8e-06 $layer=LI1_cond $X=8.705 $Y=0.765
+ $X2=8.705 $Y2=2.565
r136 34 50 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.015 $Y=0.68
+ $X2=7.93 $Y2=0.68
r137 33 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.62 $Y=0.68
+ $X2=8.705 $Y2=0.765
r138 33 34 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=8.62 $Y=0.68
+ $X2=8.015 $Y2=0.68
r139 32 49 2.85362 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.98 $Y=2.65
+ $X2=7.815 $Y2=2.65
r140 31 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.62 $Y=2.65
+ $X2=8.705 $Y2=2.565
r141 31 32 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=8.62 $Y=2.65
+ $X2=7.98 $Y2=2.65
r142 27 48 3.99587 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.815 $Y=2.37
+ $X2=7.815 $Y2=2.455
r143 27 29 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=7.815 $Y=2.37
+ $X2=7.815 $Y2=2.115
r144 26 47 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.94 $Y=0.855
+ $X2=6.815 $Y2=0.855
r145 25 52 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.845 $Y=0.855
+ $X2=7.93 $Y2=0.855
r146 25 26 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=7.845 $Y=0.855
+ $X2=6.94 $Y2=0.855
r147 21 47 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.815 $Y=0.77
+ $X2=6.815 $Y2=0.855
r148 21 23 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=6.815 $Y=0.77
+ $X2=6.815 $Y2=0.515
r149 20 42 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.945 $Y=2.455
+ $X2=5.86 $Y2=2.455
r150 19 48 2.85362 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.65 $Y=2.455
+ $X2=7.815 $Y2=2.455
r151 19 20 111.235 $w=1.68e-07 $l=1.705e-06 $layer=LI1_cond $X=7.65 $Y=2.455
+ $X2=5.945 $Y2=2.455
r152 18 40 8.04321 $w=1.7e-07 $l=2.88e-07 $layer=LI1_cond $X=5.105 $Y=0.855
+ $X2=4.817 $Y2=0.855
r153 17 47 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.69 $Y=0.855
+ $X2=6.815 $Y2=0.855
r154 17 18 103.406 $w=1.68e-07 $l=1.585e-06 $layer=LI1_cond $X=6.69 $Y=0.855
+ $X2=5.105 $Y2=0.855
r155 13 42 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=5.86 $Y=2.785
+ $X2=5.86 $Y2=2.455
r156 13 15 20.0525 $w=2.48e-07 $l=4.35e-07 $layer=LI1_cond $X=5.775 $Y=2.785
+ $X2=5.34 $Y2=2.785
r157 4 29 300 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=2 $X=7.665
+ $Y=1.96 $X2=7.815 $Y2=2.115
r158 3 15 600 $w=1.7e-07 $l=9.10041e-07 $layer=licon1_PDIFF $count=1 $X=5.07
+ $Y=1.96 $X2=5.34 $Y2=2.745
r159 2 47 182 $w=1.7e-07 $l=5.50568e-07 $layer=licon1_NDIFF $count=1 $X=6.715
+ $Y=0.37 $X2=6.855 $Y2=0.855
r160 2 23 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=6.715
+ $Y=0.37 $X2=6.855 $Y2=0.515
r161 1 38 91 $w=1.7e-07 $l=3.75566e-07 $layer=licon1_NDIFF $count=2 $X=4.545
+ $Y=0.37 $X2=4.855 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__MUX4_2%X 1 2 7 8 9 10 11 12 13 36
c24 11 0 5.38206e-20 $X=9.755 $Y=1.95
r25 34 36 1.31708 $w=3.48e-07 $l=4e-08 $layer=LI1_cond $X=9.825 $Y=1.995
+ $X2=9.825 $Y2=2.035
r26 12 13 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=9.825 $Y=2.405
+ $X2=9.825 $Y2=2.775
r27 11 34 0.75732 $w=3.48e-07 $l=2.3e-08 $layer=LI1_cond $X=9.825 $Y=1.972
+ $X2=9.825 $Y2=1.995
r28 11 45 5.05604 $w=3.48e-07 $l=1.52e-07 $layer=LI1_cond $X=9.825 $Y=1.972
+ $X2=9.825 $Y2=1.82
r29 11 12 11.4586 $w=3.48e-07 $l=3.48e-07 $layer=LI1_cond $X=9.825 $Y=2.057
+ $X2=9.825 $Y2=2.405
r30 11 36 0.724393 $w=3.48e-07 $l=2.2e-08 $layer=LI1_cond $X=9.825 $Y=2.057
+ $X2=9.825 $Y2=2.035
r31 10 45 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=9.815 $Y=1.665
+ $X2=9.815 $Y2=1.82
r32 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=9.815 $Y=1.295
+ $X2=9.815 $Y2=1.665
r33 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=9.815 $Y=0.925
+ $X2=9.815 $Y2=1.295
r34 8 27 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=9.815 $Y=0.925
+ $X2=9.815 $Y2=0.645
r35 7 27 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=9.815 $Y=0.555
+ $X2=9.815 $Y2=0.645
r36 2 11 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=9.685
+ $Y=1.84 $X2=9.835 $Y2=1.985
r37 2 13 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=9.685
+ $Y=1.84 $X2=9.835 $Y2=2.815
r38 1 27 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.675
+ $Y=0.5 $X2=9.815 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_LS__MUX4_2%VGND 1 2 3 4 5 18 24 28 32 34 36 39 40 42 43
+ 44 50 64 68 74 77 81
r91 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=0 $X2=10.32
+ $Y2=0
r92 77 78 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r93 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r94 72 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0 $X2=10.32
+ $Y2=0
r95 72 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0 $X2=9.36
+ $Y2=0
r96 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r97 69 77 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.47 $Y=0 $X2=9.385
+ $Y2=0
r98 69 71 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=9.47 $Y=0 $X2=9.84
+ $Y2=0
r99 68 80 3.96842 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=10.16 $Y=0 $X2=10.36
+ $Y2=0
r100 68 71 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=10.16 $Y=0 $X2=9.84
+ $Y2=0
r101 67 78 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=6.48 $Y=0
+ $X2=9.36 $Y2=0
r102 66 67 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r103 64 77 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.3 $Y=0 $X2=9.385
+ $Y2=0
r104 64 66 183.979 $w=1.68e-07 $l=2.82e-06 $layer=LI1_cond $X=9.3 $Y=0 $X2=6.48
+ $Y2=0
r105 63 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r106 62 63 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6
+ $Y2=0
r107 60 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r108 59 62 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.08 $Y=0 $X2=6
+ $Y2=0
r109 59 60 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r110 57 74 11.015 $w=1.7e-07 $l=2.4e-07 $layer=LI1_cond $X=3.925 $Y=0 $X2=3.685
+ $Y2=0
r111 57 59 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=3.925 $Y=0
+ $X2=4.08 $Y2=0
r112 56 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r113 55 56 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r114 53 56 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r115 52 55 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r116 52 53 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r117 50 74 11.015 $w=1.7e-07 $l=2.4e-07 $layer=LI1_cond $X=3.445 $Y=0 $X2=3.685
+ $Y2=0
r118 50 55 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=3.445 $Y=0
+ $X2=3.12 $Y2=0
r119 48 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r120 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r121 44 63 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=5.28 $Y=0 $X2=6
+ $Y2=0
r122 44 60 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=5.28 $Y=0 $X2=4.08
+ $Y2=0
r123 42 62 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=6.14 $Y=0 $X2=6
+ $Y2=0
r124 42 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.14 $Y=0 $X2=6.305
+ $Y2=0
r125 41 66 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=6.47 $Y=0 $X2=6.48
+ $Y2=0
r126 41 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.47 $Y=0 $X2=6.305
+ $Y2=0
r127 39 47 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=0.82 $Y=0 $X2=0.72
+ $Y2=0
r128 39 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.82 $Y=0 $X2=0.985
+ $Y2=0
r129 38 52 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=1.15 $Y=0 $X2=1.2
+ $Y2=0
r130 38 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.15 $Y=0 $X2=0.985
+ $Y2=0
r131 34 80 3.17474 $w=2.5e-07 $l=1.16619e-07 $layer=LI1_cond $X=10.285 $Y=0.085
+ $X2=10.36 $Y2=0
r132 34 36 25.8147 $w=2.48e-07 $l=5.6e-07 $layer=LI1_cond $X=10.285 $Y=0.085
+ $X2=10.285 $Y2=0.645
r133 30 77 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.385 $Y=0.085
+ $X2=9.385 $Y2=0
r134 30 32 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=9.385 $Y=0.085
+ $X2=9.385 $Y2=0.675
r135 26 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.305 $Y=0.085
+ $X2=6.305 $Y2=0
r136 26 28 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=6.305 $Y=0.085
+ $X2=6.305 $Y2=0.515
r137 22 74 1.96841 $w=4.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.685 $Y=0.085
+ $X2=3.685 $Y2=0
r138 22 24 10.7149 $w=4.78e-07 $l=4.3e-07 $layer=LI1_cond $X=3.685 $Y=0.085
+ $X2=3.685 $Y2=0.515
r139 18 20 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=0.985 $Y=0.515
+ $X2=0.985 $Y2=0.855
r140 16 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.985 $Y=0.085
+ $X2=0.985 $Y2=0
r141 16 18 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.985 $Y=0.085
+ $X2=0.985 $Y2=0.515
r142 5 36 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.105
+ $Y=0.5 $X2=10.245 $Y2=0.645
r143 4 32 91 $w=1.7e-07 $l=6.36396e-07 $layer=licon1_NDIFF $count=2 $X=8.785
+ $Y=0.6 $X2=9.385 $Y2=0.675
r144 3 28 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=6.165
+ $Y=0.37 $X2=6.305 $Y2=0.515
r145 2 24 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=3.465
+ $Y=0.37 $X2=3.65 $Y2=0.515
r146 1 20 182 $w=1.7e-07 $l=5.55068e-07 $layer=licon1_NDIFF $count=1 $X=0.59
+ $Y=0.47 $X2=0.985 $Y2=0.855
r147 1 18 182 $w=1.7e-07 $l=4.16893e-07 $layer=licon1_NDIFF $count=1 $X=0.59
+ $Y=0.47 $X2=0.985 $Y2=0.515
.ends

