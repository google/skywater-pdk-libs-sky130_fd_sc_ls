* File: sky130_fd_sc_ls__o221ai_2.spice
* Created: Fri Aug 28 13:48:06 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__o221ai_2.pex.spice"
.subckt sky130_fd_sc_ls__o221ai_2  VNB VPB C1 B1 B2 A1 A2 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A2	A2
* A1	A1
* B2	B2
* B1	B1
* C1	C1
* VPB	VPB
* VNB	VNB
MM1015 N_Y_M1015_d N_C1_M1015_g N_A_27_74#_M1015_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1016 N_Y_M1015_d N_C1_M1016_g N_A_27_74#_M1016_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1010 N_A_27_74#_M1010_d N_B1_M1010_g N_A_311_85#_M1010_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75003.6 A=0.111 P=1.78 MULT=1
MM1005 N_A_27_74#_M1010_d N_B2_M1005_g N_A_311_85#_M1005_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75003.1 A=0.111 P=1.78 MULT=1
MM1019 N_A_27_74#_M1019_d N_B2_M1019_g N_A_311_85#_M1005_s VNB NSHORT L=0.15
+ W=0.74 AD=0.14985 AS=0.1036 PD=1.145 PS=1.02 NRD=15.804 NRS=0 M=1 R=4.93333
+ SA=75001.1 SB=75002.7 A=0.111 P=1.78 MULT=1
MM1011 N_A_27_74#_M1019_d N_B1_M1011_g N_A_311_85#_M1011_s VNB NSHORT L=0.15
+ W=0.74 AD=0.14985 AS=0.1036 PD=1.145 PS=1.02 NRD=4.452 NRS=0 M=1 R=4.93333
+ SA=75001.6 SB=75002.1 A=0.111 P=1.78 MULT=1
MM1003 N_VGND_M1003_d N_A1_M1003_g N_A_311_85#_M1011_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1406 AS=0.1036 PD=1.12 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75002.1
+ SB=75001.7 A=0.111 P=1.78 MULT=1
MM1002 N_A_311_85#_M1002_d N_A2_M1002_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.74
+ AD=0.1221 AS=0.1406 PD=1.07 PS=1.12 NRD=6.48 NRS=4.86 M=1 R=4.93333 SA=75002.6
+ SB=75001.2 A=0.111 P=1.78 MULT=1
MM1008 N_A_311_85#_M1002_d N_A2_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1221 AS=0.1258 PD=1.07 PS=1.08 NRD=1.62 NRS=9.72 M=1 R=4.93333 SA=75003.1
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1017 N_VGND_M1008_s N_A1_M1017_g N_A_311_85#_M1017_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1258 AS=0.2146 PD=1.08 PS=2.06 NRD=0 NRS=0 M=1 R=4.93333 SA=75003.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1013 N_Y_M1013_d N_C1_M1013_g N_VPWR_M1013_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75004.9 A=0.168 P=2.54 MULT=1
MM1014 N_Y_M1013_d N_C1_M1014_g N_VPWR_M1014_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.3696 PD=1.42 PS=1.78 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75004.5 A=0.168 P=2.54 MULT=1
MM1000 N_A_376_368#_M1000_d N_B1_M1000_g N_VPWR_M1014_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.1876 AS=0.3696 PD=1.455 PS=1.78 NRD=1.7533 NRS=1.7533 M=1
+ R=7.46667 SA=75001.5 SB=75003.7 A=0.168 P=2.54 MULT=1
MM1007 N_A_376_368#_M1000_d N_B2_M1007_g N_Y_M1007_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.1876 AS=0.1764 PD=1.455 PS=1.435 NRD=7.8997 NRS=4.3931 M=1 R=7.46667
+ SA=75002 SB=75003.2 A=0.168 P=2.54 MULT=1
MM1009 N_A_376_368#_M1009_d N_B2_M1009_g N_Y_M1007_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.196 AS=0.1764 PD=1.47 PS=1.435 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75002.4 SB=75002.7 A=0.168 P=2.54 MULT=1
MM1012 N_A_376_368#_M1009_d N_B1_M1012_g N_VPWR_M1012_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.196 AS=0.224 PD=1.47 PS=1.52 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75002.9 SB=75002.2 A=0.168 P=2.54 MULT=1
MM1006 N_VPWR_M1012_s N_A1_M1006_g N_A_776_368#_M1006_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.224 AS=0.196 PD=1.52 PS=1.47 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75003.5 SB=75001.7 A=0.168 P=2.54 MULT=1
MM1001 N_Y_M1001_d N_A2_M1001_g N_A_776_368#_M1006_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75004 SB=75001.2 A=0.168 P=2.54 MULT=1
MM1004 N_Y_M1001_d N_A2_M1004_g N_A_776_368#_M1004_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75004.4 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1018 N_VPWR_M1018_d N_A1_M1018_g N_A_776_368#_M1004_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.3864 AS=0.168 PD=2.93 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75004.9 SB=75000.3 A=0.168 P=2.54 MULT=1
DX20_noxref VNB VPB NWDIODE A=11.4204 P=16
*
.include "sky130_fd_sc_ls__o221ai_2.pxi.spice"
*
.ends
*
*
