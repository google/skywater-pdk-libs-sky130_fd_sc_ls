* File: sky130_fd_sc_ls__sdfrbp_1.pex.spice
* Created: Fri Aug 28 14:02:22 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__SDFRBP_1%A_27_74# 1 2 9 11 13 16 19 22 23 25 27 32
+ 34
c77 34 0 4.33637e-20 $X=2.5 $Y=1.995
c78 25 0 1.73275e-20 $X=2.365 $Y=2.135
r79 34 37 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=2.53 $Y=1.995
+ $X2=2.53 $Y2=2.135
r80 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.5
+ $Y=1.995 $X2=2.5 $Y2=1.995
r81 31 32 12.4206 $w=9.23e-07 $l=1.65e-07 $layer=LI1_cond $X=0.89 $Y=2.512
+ $X2=1.055 $Y2=2.512
r82 25 37 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.365 $Y=2.135
+ $X2=2.53 $Y2=2.135
r83 25 32 85.4652 $w=1.68e-07 $l=1.31e-06 $layer=LI1_cond $X=2.365 $Y=2.135
+ $X2=1.055 $Y2=2.135
r84 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.23
+ $Y=1.145 $X2=1.23 $Y2=1.145
r85 20 27 0.221902 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=0.365 $Y=1.145
+ $X2=0.24 $Y2=1.145
r86 20 22 30.208 $w=3.28e-07 $l=8.65e-07 $layer=LI1_cond $X=0.365 $Y=1.145
+ $X2=1.23 $Y2=1.145
r87 19 31 9.10054 $w=9.23e-07 $l=6.9e-07 $layer=LI1_cond $X=0.2 $Y=2.512
+ $X2=0.89 $Y2=2.512
r88 18 27 7.38875 $w=2.1e-07 $l=1.83916e-07 $layer=LI1_cond $X=0.2 $Y=1.31
+ $X2=0.24 $Y2=1.145
r89 18 19 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=0.2 $Y=1.31 $X2=0.2
+ $Y2=2.05
r90 14 27 7.38875 $w=2.1e-07 $l=1.65e-07 $layer=LI1_cond $X=0.24 $Y=0.98
+ $X2=0.24 $Y2=1.145
r91 14 16 18.4391 $w=2.48e-07 $l=4e-07 $layer=LI1_cond $X=0.24 $Y=0.98 $X2=0.24
+ $Y2=0.58
r92 11 35 52.2586 $w=2.99e-07 $l=2.57391e-07 $layer=POLY_cond $X=2.485 $Y=2.245
+ $X2=2.5 $Y2=1.995
r93 11 13 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.485 $Y=2.245
+ $X2=2.485 $Y2=2.64
r94 7 23 45.5222 $w=2.7e-07 $l=3.27261e-07 $layer=POLY_cond $X=1.485 $Y=0.98
+ $X2=1.23 $Y2=1.145
r95 7 9 187.16 $w=1.5e-07 $l=3.65e-07 $layer=POLY_cond $X=1.485 $Y=0.98
+ $X2=1.485 $Y2=0.615
r96 2 31 150 $w=1.7e-07 $l=8.24318e-07 $layer=licon1_PDIFF $count=4 $X=0.135
+ $Y=2.32 $X2=0.89 $Y2=2.465
r97 1 16 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRBP_1%SCE 3 6 7 9 11 12 14 19 20 21 22 23 26 27
+ 31 32 33 38 46 49 51 60 62
c97 27 0 3.49301e-19 $X=2.51 $Y=1.425
c98 21 0 1.69076e-19 $X=2.625 $Y=0.9
r99 51 60 2.36399 $w=3.88e-07 $l=8e-08 $layer=LI1_cond $X=1.6 $Y=1.685 $X2=1.68
+ $Y2=1.685
r100 44 46 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.45 $Y=1.715
+ $X2=1.615 $Y2=1.715
r101 44 45 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.45
+ $Y=1.715 $X2=1.45 $Y2=1.715
r102 42 44 58.5785 $w=3.3e-07 $l=3.35e-07 $layer=POLY_cond $X=1.115 $Y=1.715
+ $X2=1.45 $Y2=1.715
r103 38 42 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.025 $Y=1.715
+ $X2=1.115 $Y2=1.715
r104 38 40 44.5896 $w=3.3e-07 $l=2.55e-07 $layer=POLY_cond $X=1.025 $Y=1.715
+ $X2=0.77 $Y2=1.715
r105 33 62 7.07103 $w=3.88e-07 $l=1.13e-07 $layer=LI1_cond $X=1.682 $Y=1.685
+ $X2=1.795 $Y2=1.685
r106 33 60 0.0590996 $w=3.88e-07 $l=2e-09 $layer=LI1_cond $X=1.682 $Y=1.685
+ $X2=1.68 $Y2=1.685
r107 33 51 0.0886495 $w=3.88e-07 $l=3e-09 $layer=LI1_cond $X=1.597 $Y=1.685
+ $X2=1.6 $Y2=1.685
r108 33 45 4.34382 $w=3.88e-07 $l=1.47e-07 $layer=LI1_cond $X=1.597 $Y=1.685
+ $X2=1.45 $Y2=1.685
r109 32 45 7.38745 $w=3.88e-07 $l=2.5e-07 $layer=LI1_cond $X=1.2 $Y=1.685
+ $X2=1.45 $Y2=1.685
r110 31 32 14.1839 $w=3.88e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.685
+ $X2=1.2 $Y2=1.685
r111 31 40 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.77
+ $Y=1.715 $X2=0.77 $Y2=1.715
r112 27 49 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.51 $Y=1.425
+ $X2=2.51 $Y2=1.26
r113 26 29 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=2.56 $Y=1.425
+ $X2=2.56 $Y2=1.575
r114 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.51
+ $Y=1.425 $X2=2.51 $Y2=1.425
r115 23 29 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.395 $Y=1.575
+ $X2=2.56 $Y2=1.575
r116 23 62 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=2.395 $Y=1.575
+ $X2=1.795 $Y2=1.575
r117 22 49 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=2.6 $Y=1.05 $X2=2.6
+ $Y2=1.26
r118 21 22 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=2.625 $Y=0.9
+ $X2=2.625 $Y2=1.05
r119 20 40 34.9723 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=0.57 $Y=1.715
+ $X2=0.77 $Y2=1.715
r120 19 21 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.65 $Y=0.615
+ $X2=2.65 $Y2=0.9
r121 12 14 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.615 $Y=2.245
+ $X2=1.615 $Y2=2.64
r122 11 12 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.615 $Y=2.155
+ $X2=1.615 $Y2=2.245
r123 10 46 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.615 $Y=1.88
+ $X2=1.615 $Y2=1.715
r124 10 11 106.895 $w=1.8e-07 $l=2.75e-07 $layer=POLY_cond $X=1.615 $Y=1.88
+ $X2=1.615 $Y2=2.155
r125 7 9 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.115 $Y=2.245
+ $X2=1.115 $Y2=2.64
r126 6 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.115 $Y=2.155
+ $X2=1.115 $Y2=2.245
r127 5 42 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.115 $Y=1.88
+ $X2=1.115 $Y2=1.715
r128 5 6 106.895 $w=1.8e-07 $l=2.75e-07 $layer=POLY_cond $X=1.115 $Y=1.88
+ $X2=1.115 $Y2=2.155
r129 1 20 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=0.495 $Y=1.55
+ $X2=0.57 $Y2=1.715
r130 1 3 497.383 $w=1.5e-07 $l=9.7e-07 $layer=POLY_cond $X=0.495 $Y=1.55
+ $X2=0.495 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRBP_1%D 3 6 7 9 10 13 14
c46 14 0 3.42316e-19 $X=1.935 $Y=1.145
c47 7 0 4.33637e-20 $X=2.035 $Y=2.245
r48 13 16 40.8147 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=1.947 $Y=1.145
+ $X2=1.947 $Y2=1.31
r49 13 15 46.504 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=1.947 $Y=1.145
+ $X2=1.947 $Y2=0.98
r50 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.935
+ $Y=1.145 $X2=1.935 $Y2=1.145
r51 10 14 6.1 $w=4.98e-07 $l=2.55e-07 $layer=LI1_cond $X=1.68 $Y=1.06 $X2=1.935
+ $Y2=1.06
r52 7 9 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.035 $Y=2.245
+ $X2=2.035 $Y2=2.64
r53 6 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.035 $Y=2.155 $X2=2.035
+ $Y2=2.245
r54 6 16 328.46 $w=1.8e-07 $l=8.45e-07 $layer=POLY_cond $X=2.035 $Y=2.155
+ $X2=2.035 $Y2=1.31
r55 3 15 187.16 $w=1.5e-07 $l=3.65e-07 $layer=POLY_cond $X=1.97 $Y=0.615
+ $X2=1.97 $Y2=0.98
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRBP_1%SCD 3 6 10 11 12 13 17
c42 12 0 1.58733e-19 $X=3.12 $Y=1.665
c43 11 0 7.60406e-20 $X=3.05 $Y=2.245
c44 6 0 1.93733e-19 $X=3.04 $Y=0.615
r45 12 13 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.1 $Y=1.605 $X2=3.1
+ $Y2=2.035
r46 12 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.05
+ $Y=1.605 $X2=3.05 $Y2=1.605
r47 10 17 83.0591 $w=3.3e-07 $l=4.75e-07 $layer=POLY_cond $X=3.05 $Y=2.08
+ $X2=3.05 $Y2=1.605
r48 10 11 38.3209 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.05 $Y=2.08
+ $X2=3.05 $Y2=2.245
r49 9 17 38.0424 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.05 $Y=1.44
+ $X2=3.05 $Y2=1.605
r50 6 9 423.032 $w=1.5e-07 $l=8.25e-07 $layer=POLY_cond $X=3.04 $Y=0.615
+ $X2=3.04 $Y2=1.44
r51 3 11 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.035 $Y=2.64
+ $X2=3.035 $Y2=2.245
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRBP_1%CLK 1 2 3 5 7 10 12 13 14 18 19 23
c61 23 0 3.88236e-19 $X=4.08 $Y=1.295
c62 13 0 1.4151e-19 $X=4.62 $Y=1.885
r63 21 23 0.542222 $w=4.5e-07 $l=2e-08 $layer=LI1_cond $X=4.06 $Y=1.405 $X2=4.08
+ $Y2=1.405
r64 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.95
+ $Y=1.115 $X2=3.95 $Y2=1.115
r65 14 21 4.60977 $w=2.73e-07 $l=1.1e-07 $layer=LI1_cond $X=3.922 $Y=1.295
+ $X2=3.922 $Y2=1.405
r66 14 19 7.54326 $w=2.73e-07 $l=1.8e-07 $layer=LI1_cond $X=3.922 $Y=1.295
+ $X2=3.922 $Y2=1.115
r67 14 23 0.867556 $w=4.5e-07 $l=3.2e-08 $layer=LI1_cond $X=4.112 $Y=1.405
+ $X2=4.08 $Y2=1.405
r68 11 18 51.5841 $w=3.3e-07 $l=2.95e-07 $layer=POLY_cond $X=3.95 $Y=1.41
+ $X2=3.95 $Y2=1.115
r69 10 13 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=4.645 $Y=2.46
+ $X2=4.645 $Y2=1.885
r70 7 13 37.4512 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=4.62 $Y=1.785 $X2=4.62
+ $Y2=1.885
r71 6 12 23.6879 $w=1.75e-07 $l=1.05e-07 $layer=POLY_cond $X=4.62 $Y=1.62
+ $X2=4.62 $Y2=1.515
r72 6 7 54.7102 $w=2e-07 $l=1.65e-07 $layer=POLY_cond $X=4.62 $Y=1.62 $X2=4.62
+ $Y2=1.785
r73 3 12 23.6879 $w=1.75e-07 $l=1.16833e-07 $layer=POLY_cond $X=4.595 $Y=1.41
+ $X2=4.62 $Y2=1.515
r74 3 5 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=4.595 $Y=1.41
+ $X2=4.595 $Y2=0.965
r75 2 11 28.6974 $w=2.1e-07 $l=2.11069e-07 $layer=POLY_cond $X=4.115 $Y=1.515
+ $X2=3.95 $Y2=1.41
r76 1 12 2.7459 $w=2.1e-07 $l=1e-07 $layer=POLY_cond $X=4.52 $Y=1.515 $X2=4.62
+ $Y2=1.515
r77 1 2 127.894 $w=2.1e-07 $l=4.05e-07 $layer=POLY_cond $X=4.52 $Y=1.515
+ $X2=4.115 $Y2=1.515
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRBP_1%A_1034_392# 1 2 8 9 11 12 16 18 20 21 22 23
+ 25 26 33 35 36 37 38 40 44 45 46 48 49 50 52 54 57 61 68 69 73 75
c217 69 0 1.6856e-19 $X=9.27 $Y=1.07
c218 68 0 1.89827e-19 $X=9.27 $Y=1.07
c219 46 0 1.61901e-19 $X=7.22 $Y=0.665
c220 9 0 1.58245e-19 $X=6.135 $Y=2.21
r221 69 81 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=9.27 $Y=1.07 $X2=9.27
+ $Y2=1.16
r222 68 69 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.27
+ $Y=1.07 $X2=9.27 $Y2=1.07
r223 65 68 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=8.91 $Y=0.99
+ $X2=9.27 $Y2=0.99
r224 60 61 9.72653 $w=4.03e-07 $l=2.15e-07 $layer=LI1_cond $X=5.422 $Y=1.07
+ $X2=5.422 $Y2=1.285
r225 57 58 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.67
+ $Y=2.065 $X2=9.67 $Y2=2.065
r226 55 73 0.201461 $w=2.5e-07 $l=1.15e-07 $layer=LI1_cond $X=9.63 $Y=1.575
+ $X2=9.63 $Y2=1.46
r227 55 57 22.5879 $w=2.48e-07 $l=4.9e-07 $layer=LI1_cond $X=9.63 $Y=1.575
+ $X2=9.63 $Y2=2.065
r228 54 73 18.0382 $w=2.28e-07 $l=3.6e-07 $layer=LI1_cond $X=9.27 $Y=1.46
+ $X2=9.63 $Y2=1.46
r229 54 68 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=9.27 $Y=1.345
+ $X2=9.27 $Y2=1.075
r230 52 65 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.91 $Y=0.905
+ $X2=8.91 $Y2=0.99
r231 51 52 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=8.91 $Y=0.425
+ $X2=8.91 $Y2=0.905
r232 49 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.825 $Y=0.34
+ $X2=8.91 $Y2=0.425
r233 49 50 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=8.825 $Y=0.34
+ $X2=8.1 $Y2=0.34
r234 47 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.015 $Y=0.425
+ $X2=8.1 $Y2=0.34
r235 47 48 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=8.015 $Y=0.425
+ $X2=8.015 $Y2=0.58
r236 45 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.93 $Y=0.665
+ $X2=8.015 $Y2=0.58
r237 45 46 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=7.93 $Y=0.665
+ $X2=7.22 $Y2=0.665
r238 44 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.135 $Y=0.58
+ $X2=7.22 $Y2=0.665
r239 43 44 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=7.135 $Y=0.425
+ $X2=7.135 $Y2=0.58
r240 41 78 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.085 $Y=1.71
+ $X2=6.085 $Y2=1.875
r241 41 75 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=6.085 $Y=1.71
+ $X2=6.085 $Y2=1.635
r242 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.085
+ $Y=1.71 $X2=6.085 $Y2=1.71
r243 38 40 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=5.63 $Y=1.71
+ $X2=6.085 $Y2=1.71
r244 36 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.05 $Y=0.34
+ $X2=7.135 $Y2=0.425
r245 36 37 93.2941 $w=1.68e-07 $l=1.43e-06 $layer=LI1_cond $X=7.05 $Y=0.34
+ $X2=5.62 $Y2=0.34
r246 35 38 10.1667 $w=1.78e-07 $l=1.65e-07 $layer=LI1_cond $X=5.54 $Y=1.545
+ $X2=5.54 $Y2=1.71
r247 35 61 16.0202 $w=1.78e-07 $l=2.6e-07 $layer=LI1_cond $X=5.54 $Y=1.545
+ $X2=5.54 $Y2=1.285
r248 33 60 8.25206 $w=4.03e-07 $l=2.9e-07 $layer=LI1_cond $X=5.417 $Y=0.78
+ $X2=5.417 $Y2=1.07
r249 30 37 8.41448 $w=1.7e-07 $l=2.41793e-07 $layer=LI1_cond $X=5.417 $Y=0.425
+ $X2=5.62 $Y2=0.34
r250 30 33 10.1017 $w=4.03e-07 $l=3.55e-07 $layer=LI1_cond $X=5.417 $Y=0.425
+ $X2=5.417 $Y2=0.78
r251 26 38 23.1061 $w=1.78e-07 $l=3.75e-07 $layer=LI1_cond $X=5.54 $Y=2.085
+ $X2=5.54 $Y2=1.71
r252 26 28 5.76222 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=5.45 $Y=2.085
+ $X2=5.32 $Y2=2.085
r253 23 58 60.889 $w=3.02e-07 $l=3.46215e-07 $layer=POLY_cond $X=9.77 $Y=2.37
+ $X2=9.682 $Y2=2.065
r254 23 25 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=9.77 $Y=2.37
+ $X2=9.77 $Y2=2.655
r255 21 81 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.105 $Y=1.16
+ $X2=9.27 $Y2=1.16
r256 21 22 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=9.105 $Y=1.16
+ $X2=8.735 $Y2=1.16
r257 18 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.66 $Y=1.085
+ $X2=8.735 $Y2=1.16
r258 18 20 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=8.66 $Y=1.085
+ $X2=8.66 $Y2=0.69
r259 14 16 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=6.525 $Y=1.545
+ $X2=6.525 $Y2=0.805
r260 13 75 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.25 $Y=1.635
+ $X2=6.085 $Y2=1.635
r261 12 14 27.2212 $w=1.8e-07 $l=1.21861e-07 $layer=POLY_cond $X=6.45 $Y=1.635
+ $X2=6.525 $Y2=1.545
r262 12 13 77.7419 $w=1.8e-07 $l=2e-07 $layer=POLY_cond $X=6.45 $Y=1.635
+ $X2=6.25 $Y2=1.635
r263 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.135 $Y=2.21
+ $X2=6.135 $Y2=2.495
r264 8 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.135 $Y=2.12 $X2=6.135
+ $Y2=2.21
r265 8 78 95.2339 $w=1.8e-07 $l=2.45e-07 $layer=POLY_cond $X=6.135 $Y=2.12
+ $X2=6.135 $Y2=1.875
r266 2 28 600 $w=1.7e-07 $l=2.33238e-07 $layer=licon1_PDIFF $count=1 $X=5.17
+ $Y=1.96 $X2=5.32 $Y2=2.13
r267 1 33 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=5.22
+ $Y=0.595 $X2=5.36 $Y2=0.78
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRBP_1%A_1367_93# 1 2 9 13 17 18 21 23 24 26 32 33
c111 33 0 1.6856e-19 $X=8.57 $Y=0.842
c112 24 0 4.08738e-20 $X=8.81 $Y=1.415
c113 9 0 1.43931e-19 $X=6.91 $Y=0.805
r114 39 41 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=6.91 $Y=1.64
+ $X2=6.945 $Y2=1.64
r115 31 33 3.0204 $w=4.93e-07 $l=1.25e-07 $layer=LI1_cond $X=8.445 $Y=0.842
+ $X2=8.57 $Y2=0.842
r116 31 32 9.72819 $w=4.93e-07 $l=1.75e-07 $layer=LI1_cond $X=8.445 $Y=0.842
+ $X2=8.27 $Y2=0.842
r117 26 28 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=8.81 $Y=1.88
+ $X2=8.81 $Y2=2.59
r118 24 35 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=8.81 $Y=1.33
+ $X2=8.57 $Y2=1.33
r119 24 26 21.4354 $w=2.48e-07 $l=4.65e-07 $layer=LI1_cond $X=8.81 $Y=1.415
+ $X2=8.81 $Y2=1.88
r120 23 35 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.57 $Y=1.245
+ $X2=8.57 $Y2=1.33
r121 22 33 7.09362 $w=1.7e-07 $l=2.48e-07 $layer=LI1_cond $X=8.57 $Y=1.09
+ $X2=8.57 $Y2=0.842
r122 22 23 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=8.57 $Y=1.09
+ $X2=8.57 $Y2=1.245
r123 21 32 65.5668 $w=1.68e-07 $l=1.005e-06 $layer=LI1_cond $X=7.265 $Y=1.005
+ $X2=8.27 $Y2=1.005
r124 18 41 34.9723 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=7.145 $Y=1.64
+ $X2=6.945 $Y2=1.64
r125 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.145
+ $Y=1.64 $X2=7.145 $Y2=1.64
r126 15 21 7.07814 $w=1.7e-07 $l=1.56844e-07 $layer=LI1_cond $X=7.145 $Y=1.09
+ $X2=7.265 $Y2=1.005
r127 15 17 26.4102 $w=2.38e-07 $l=5.5e-07 $layer=LI1_cond $X=7.145 $Y=1.09
+ $X2=7.145 $Y2=1.64
r128 11 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.945 $Y=1.805
+ $X2=6.945 $Y2=1.64
r129 11 13 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.945 $Y=1.805
+ $X2=6.945 $Y2=2.495
r130 7 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.91 $Y=1.475
+ $X2=6.91 $Y2=1.64
r131 7 9 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=6.91 $Y=1.475
+ $X2=6.91 $Y2=0.805
r132 2 28 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=8.62
+ $Y=1.735 $X2=8.77 $Y2=2.59
r133 2 26 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=8.62
+ $Y=1.735 $X2=8.77 $Y2=1.88
r134 1 31 182 $w=1.7e-07 $l=5.0951e-07 $layer=licon1_NDIFF $count=1 $X=8.295
+ $Y=0.37 $X2=8.445 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRBP_1%RESET_B 4 7 8 9 10 11 15 16 18 20 23 27 34
+ 37 41 43 44 45 46 47 48 56 60 62 65 67 68 69
c249 68 0 1.5378e-19 $X=10.9 $Y=1.845
c250 67 0 2.44776e-20 $X=10.9 $Y=1.845
c251 60 0 1.4151e-19 $X=3.95 $Y=1.995
c252 44 0 8.18376e-20 $X=10.81 $Y=2.37
c253 41 0 6.47027e-20 $X=10.81 $Y=1.335
c254 34 0 9.37604e-20 $X=3.56 $Y=2.245
c255 15 0 1.75393e-19 $X=7.3 $Y=0.805
c256 10 0 1.98276e-19 $X=3.93 $Y=1.995
r257 68 77 5.91795 $w=3.68e-07 $l=1.9e-07 $layer=LI1_cond $X=10.88 $Y=1.845
+ $X2=10.88 $Y2=2.035
r258 67 70 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.9 $Y=1.845
+ $X2=10.9 $Y2=2.01
r259 67 69 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.9 $Y=1.845
+ $X2=10.9 $Y2=1.68
r260 67 68 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.9
+ $Y=1.845 $X2=10.9 $Y2=1.845
r261 64 65 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.86
+ $Y=1.96 $X2=7.86 $Y2=1.96
r262 62 64 39.5449 $w=3.23e-07 $l=2.65e-07 $layer=POLY_cond $X=7.595 $Y=2.002
+ $X2=7.86 $Y2=2.002
r263 59 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.95
+ $Y=1.995 $X2=3.95 $Y2=1.995
r264 56 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=2.035
+ $X2=10.8 $Y2=2.035
r265 54 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=2.035
+ $X2=7.92 $Y2=2.035
r266 50 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=2.035
+ $X2=4.08 $Y2=2.035
r267 48 54 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.065 $Y=2.035
+ $X2=7.92 $Y2=2.035
r268 47 56 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=10.655 $Y=2.035
+ $X2=10.8 $Y2=2.035
r269 47 48 3.20544 $w=1.4e-07 $l=2.59e-06 $layer=MET1_cond $X=10.655 $Y=2.035
+ $X2=8.065 $Y2=2.035
r270 46 50 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.225 $Y=2.035
+ $X2=4.08 $Y2=2.035
r271 45 54 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.775 $Y=2.035
+ $X2=7.92 $Y2=2.035
r272 45 46 4.39356 $w=1.4e-07 $l=3.55e-06 $layer=MET1_cond $X=7.775 $Y=2.035
+ $X2=4.225 $Y2=2.035
r273 43 44 47.3682 $w=2.1e-07 $l=1.5e-07 $layer=POLY_cond $X=10.81 $Y=2.22
+ $X2=10.81 $Y2=2.37
r274 43 70 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=10.84 $Y=2.22
+ $X2=10.84 $Y2=2.01
r275 39 41 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=10.545 $Y=1.335
+ $X2=10.81 $Y2=1.335
r276 35 37 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=7.3 $Y=1.19
+ $X2=7.595 $Y2=1.19
r277 28 41 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.81 $Y=1.41
+ $X2=10.81 $Y2=1.335
r278 28 69 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=10.81 $Y=1.41
+ $X2=10.81 $Y2=1.68
r279 27 44 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=10.795 $Y=2.655
+ $X2=10.795 $Y2=2.37
r280 21 39 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.545 $Y=1.26
+ $X2=10.545 $Y2=1.335
r281 21 23 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=10.545 $Y=1.26
+ $X2=10.545 $Y2=0.58
r282 20 62 20.7134 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.595 $Y=1.795
+ $X2=7.595 $Y2=2.002
r283 19 37 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.595 $Y=1.265
+ $X2=7.595 $Y2=1.19
r284 19 20 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=7.595 $Y=1.265
+ $X2=7.595 $Y2=1.795
r285 16 62 29.8452 $w=3.23e-07 $l=2.91314e-07 $layer=POLY_cond $X=7.395 $Y=2.21
+ $X2=7.595 $Y2=2.002
r286 16 18 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.395 $Y=2.21
+ $X2=7.395 $Y2=2.495
r287 13 35 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.3 $Y=1.115
+ $X2=7.3 $Y2=1.19
r288 13 15 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=7.3 $Y=1.115
+ $X2=7.3 $Y2=0.805
r289 12 15 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=7.3 $Y=0.255
+ $X2=7.3 $Y2=0.805
r290 11 34 67.3007 $w=2.7e-07 $l=2.5e-07 $layer=POLY_cond $X=3.56 $Y=1.995
+ $X2=3.56 $Y2=2.245
r291 11 33 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.56 $Y=1.995
+ $X2=3.56 $Y2=1.83
r292 10 59 2.92121 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=3.93 $Y=1.995
+ $X2=3.95 $Y2=1.995
r293 10 11 41.0924 $w=3.3e-07 $l=2.35e-07 $layer=POLY_cond $X=3.93 $Y=1.995
+ $X2=3.695 $Y2=1.995
r294 8 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.225 $Y=0.18
+ $X2=7.3 $Y2=0.255
r295 8 9 1871.6 $w=1.5e-07 $l=3.65e-06 $layer=POLY_cond $X=7.225 $Y=0.18
+ $X2=3.575 $Y2=0.18
r296 7 34 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.605 $Y=2.64
+ $X2=3.605 $Y2=2.245
r297 4 33 623.011 $w=1.5e-07 $l=1.215e-06 $layer=POLY_cond $X=3.5 $Y=0.615
+ $X2=3.5 $Y2=1.83
r298 1 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.5 $Y=0.255
+ $X2=3.575 $Y2=0.18
r299 1 4 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=3.5 $Y=0.255 $X2=3.5
+ $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRBP_1%A_1234_119# 1 2 3 12 14 16 17 21 24 26 27
+ 30 33 35 39 43 44 46 47 50
c138 43 0 7.56682e-20 $X=6.77 $Y=2.075
c139 35 0 2.13861e-20 $X=8.15 $Y=1.41
c140 24 0 1.75393e-19 $X=6.77 $Y=1.985
c141 21 0 1.51844e-20 $X=6.685 $Y=0.945
c142 17 0 1.58245e-19 $X=6.685 $Y=2.555
r143 50 51 59.3371 $w=2.64e-07 $l=3.25e-07 $layer=POLY_cond $X=8.22 $Y=1.452
+ $X2=8.545 $Y2=1.452
r144 46 47 10.0337 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=7.6 $Y=2.53 $X2=7.6
+ $Y2=2.32
r145 39 41 4.78707 $w=3.23e-07 $l=1.35e-07 $layer=LI1_cond $X=6.307 $Y=0.81
+ $X2=6.307 $Y2=0.945
r146 36 50 12.7803 $w=2.64e-07 $l=7e-08 $layer=POLY_cond $X=8.15 $Y=1.452
+ $X2=8.22 $Y2=1.452
r147 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.15
+ $Y=1.41 $X2=8.15 $Y2=1.41
r148 33 35 22.0379 $w=2.83e-07 $l=5.45e-07 $layer=LI1_cond $X=7.605 $Y=1.402
+ $X2=8.15 $Y2=1.402
r149 31 44 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=7.52 $Y=2.165 $X2=7.52
+ $Y2=2.075
r150 31 47 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=7.52 $Y=2.165
+ $X2=7.52 $Y2=2.32
r151 30 44 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=7.52 $Y=1.985 $X2=7.52
+ $Y2=2.075
r152 29 33 7.39867 $w=2.85e-07 $l=1.80566e-07 $layer=LI1_cond $X=7.52 $Y=1.545
+ $X2=7.605 $Y2=1.402
r153 29 30 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=7.52 $Y=1.545
+ $X2=7.52 $Y2=1.985
r154 28 43 1.13756 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=6.855 $Y=2.075
+ $X2=6.77 $Y2=2.075
r155 27 44 1.13756 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=7.435 $Y=2.075
+ $X2=7.52 $Y2=2.075
r156 27 28 35.7374 $w=1.78e-07 $l=5.8e-07 $layer=LI1_cond $X=7.435 $Y=2.075
+ $X2=6.855 $Y2=2.075
r157 25 43 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=6.77 $Y=2.165 $X2=6.77
+ $Y2=2.075
r158 25 26 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=6.77 $Y=2.165
+ $X2=6.77 $Y2=2.385
r159 24 43 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=6.77 $Y=1.985 $X2=6.77
+ $Y2=2.075
r160 23 24 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=6.77 $Y=1.03
+ $X2=6.77 $Y2=1.985
r161 22 41 4.53325 $w=1.7e-07 $l=1.63e-07 $layer=LI1_cond $X=6.47 $Y=0.945
+ $X2=6.307 $Y2=0.945
r162 21 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.685 $Y=0.945
+ $X2=6.77 $Y2=1.03
r163 21 22 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=6.685 $Y=0.945
+ $X2=6.47 $Y2=0.945
r164 17 26 7.85115 $w=3.4e-07 $l=2.08207e-07 $layer=LI1_cond $X=6.685 $Y=2.555
+ $X2=6.77 $Y2=2.385
r165 17 19 11.016 $w=3.38e-07 $l=3.25e-07 $layer=LI1_cond $X=6.685 $Y=2.555
+ $X2=6.36 $Y2=2.555
r166 14 51 15.9823 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=8.545 $Y=1.66
+ $X2=8.545 $Y2=1.452
r167 14 16 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=8.545 $Y=1.66
+ $X2=8.545 $Y2=2.235
r168 10 50 15.9823 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=8.22 $Y=1.245
+ $X2=8.22 $Y2=1.452
r169 10 12 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=8.22 $Y=1.245
+ $X2=8.22 $Y2=0.69
r170 3 46 600 $w=1.7e-07 $l=3.11087e-07 $layer=licon1_PDIFF $count=1 $X=7.47
+ $Y=2.285 $X2=7.62 $Y2=2.53
r171 2 19 600 $w=1.7e-07 $l=3.36749e-07 $layer=licon1_PDIFF $count=1 $X=6.21
+ $Y=2.285 $X2=6.36 $Y2=2.555
r172 1 39 182 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=1 $X=6.17
+ $Y=0.595 $X2=6.31 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRBP_1%A_835_98# 1 2 7 9 10 12 14 15 16 17 19 21
+ 24 26 28 29 33 34 35 38 40 41 44 46 50 53
c179 53 0 1.8996e-19 $X=5.115 $Y=1.635
c180 50 0 9.37604e-20 $X=4.93 $Y=1.852
c181 38 0 1.87652e-19 $X=9.755 $Y=0.58
c182 35 0 6.22599e-20 $X=9.07 $Y=1.585
c183 34 0 2.17443e-21 $X=9.68 $Y=1.585
c184 24 0 7.56682e-20 $X=6.585 $Y=2.495
c185 19 0 1.51844e-20 $X=6.095 $Y=1.115
c186 7 0 1.94423e-19 $X=5.095 $Y=1.875
r187 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.115
+ $Y=1.635 $X2=5.115 $Y2=1.635
r188 50 52 5.09481 $w=4.43e-07 $l=2.95354e-07 $layer=LI1_cond $X=4.93 $Y=1.852
+ $X2=5.115 $Y2=1.635
r189 49 50 14.0451 $w=4.43e-07 $l=5.1e-07 $layer=LI1_cond $X=4.42 $Y=1.852
+ $X2=4.93 $Y2=1.852
r190 46 47 9.03704 $w=3.51e-07 $l=2.6e-07 $layer=LI1_cond $X=4.335 $Y=0.665
+ $X2=4.335 $Y2=0.925
r191 44 50 4.57747 $w=2.3e-07 $l=3.97e-07 $layer=LI1_cond $X=4.93 $Y=1.455
+ $X2=4.93 $Y2=1.852
r192 43 44 22.2973 $w=2.28e-07 $l=4.45e-07 $layer=LI1_cond $X=4.93 $Y=1.01
+ $X2=4.93 $Y2=1.455
r193 42 47 4.99104 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=4.535 $Y=0.925
+ $X2=4.335 $Y2=0.925
r194 41 43 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=4.815 $Y=0.925
+ $X2=4.93 $Y2=1.01
r195 41 42 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=4.815 $Y=0.925
+ $X2=4.535 $Y2=0.925
r196 36 38 476.872 $w=1.5e-07 $l=9.3e-07 $layer=POLY_cond $X=9.755 $Y=1.51
+ $X2=9.755 $Y2=0.58
r197 34 36 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.68 $Y=1.585
+ $X2=9.755 $Y2=1.51
r198 34 35 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=9.68 $Y=1.585
+ $X2=9.07 $Y2=1.585
r199 31 33 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=8.995 $Y=2.81
+ $X2=8.995 $Y2=2.235
r200 30 35 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.995 $Y=1.66
+ $X2=9.07 $Y2=1.585
r201 30 33 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=8.995 $Y=1.66
+ $X2=8.995 $Y2=2.235
r202 28 31 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=8.995 $Y=2.9
+ $X2=8.995 $Y2=2.81
r203 28 29 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=8.995 $Y=2.9
+ $X2=8.995 $Y2=3.075
r204 27 40 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.66 $Y=3.15
+ $X2=6.585 $Y2=3.15
r205 26 29 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=8.905 $Y=3.15
+ $X2=8.995 $Y2=3.075
r206 26 27 1151.16 $w=1.5e-07 $l=2.245e-06 $layer=POLY_cond $X=8.905 $Y=3.15
+ $X2=6.66 $Y2=3.15
r207 22 40 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.585 $Y=3.075
+ $X2=6.585 $Y2=3.15
r208 22 24 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.585 $Y=3.075
+ $X2=6.585 $Y2=2.495
r209 19 21 99.6133 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=6.095 $Y=1.115
+ $X2=6.095 $Y2=0.805
r210 18 53 37.7859 $w=5.23e-07 $l=5.69122e-07 $layer=POLY_cond $X=5.71 $Y=1.225
+ $X2=5.33 $Y2=1.635
r211 17 19 28.2037 $w=2.2e-07 $l=1.42653e-07 $layer=POLY_cond $X=6.02 $Y=1.225
+ $X2=6.095 $Y2=1.115
r212 17 18 90.4236 $w=2.2e-07 $l=3.1e-07 $layer=POLY_cond $X=6.02 $Y=1.225
+ $X2=5.71 $Y2=1.225
r213 15 40 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.51 $Y=3.15
+ $X2=6.585 $Y2=3.15
r214 15 16 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=6.51 $Y=3.15
+ $X2=5.69 $Y2=3.15
r215 14 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.615 $Y=3.075
+ $X2=5.69 $Y2=3.15
r216 13 53 46.2206 $w=2.61e-07 $l=3.86814e-07 $layer=POLY_cond $X=5.615 $Y=1.875
+ $X2=5.33 $Y2=1.635
r217 13 14 615.319 $w=1.5e-07 $l=1.2e-06 $layer=POLY_cond $X=5.615 $Y=1.875
+ $X2=5.615 $Y2=3.075
r218 10 18 44.3687 $w=5.23e-07 $l=6.50961e-07 $layer=POLY_cond $X=5.145 $Y=1.41
+ $X2=5.71 $Y2=1.225
r219 10 12 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=5.145 $Y=1.41
+ $X2=5.145 $Y2=0.965
r220 7 53 46.2206 $w=2.61e-07 $l=3.37639e-07 $layer=POLY_cond $X=5.095 $Y=1.875
+ $X2=5.33 $Y2=1.635
r221 7 9 187.98 $w=1.5e-07 $l=5.85e-07 $layer=POLY_cond $X=5.095 $Y=1.875
+ $X2=5.095 $Y2=2.46
r222 2 49 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=4.275
+ $Y=1.96 $X2=4.42 $Y2=2.085
r223 1 46 182 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_NDIFF $count=1 $X=4.175
+ $Y=0.49 $X2=4.32 $Y2=0.665
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRBP_1%A_2008_48# 1 2 9 11 12 13 15 18 21 22 25 28
+ 29 31 32 34 35 37
c136 29 0 1.60243e-20 $X=11.675 $Y=0.665
c137 21 0 2.44776e-20 $X=10.855 $Y=2.405
c138 18 0 6.47027e-20 $X=10.36 $Y=1.815
r139 37 39 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=11.12 $Y=0.55
+ $X2=11.12 $Y2=0.665
r140 33 34 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=11.76 $Y=0.75
+ $X2=11.76 $Y2=1.63
r141 31 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.675 $Y=1.715
+ $X2=11.76 $Y2=1.63
r142 31 32 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=11.675 $Y=1.715
+ $X2=11.405 $Y2=1.715
r143 30 39 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.285 $Y=0.665
+ $X2=11.12 $Y2=0.665
r144 29 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.675 $Y=0.665
+ $X2=11.76 $Y2=0.75
r145 29 30 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=11.675 $Y=0.665
+ $X2=11.285 $Y2=0.665
r146 28 35 3.70735 $w=2.5e-07 $l=2.28583e-07 $layer=LI1_cond $X=11.32 $Y=2.32
+ $X2=11.13 $Y2=2.405
r147 27 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.32 $Y=1.8
+ $X2=11.405 $Y2=1.715
r148 27 28 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=11.32 $Y=1.8
+ $X2=11.32 $Y2=2.32
r149 23 35 3.70735 $w=2.5e-07 $l=1.46458e-07 $layer=LI1_cond $X=11.02 $Y=2.49
+ $X2=11.13 $Y2=2.405
r150 23 25 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=11.02 $Y=2.49
+ $X2=11.02 $Y2=2.655
r151 21 35 2.76166 $w=1.7e-07 $l=2.75e-07 $layer=LI1_cond $X=10.855 $Y=2.405
+ $X2=11.13 $Y2=2.405
r152 21 22 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=10.855 $Y=2.405
+ $X2=10.525 $Y2=2.405
r153 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.36
+ $Y=1.815 $X2=10.36 $Y2=1.815
r154 16 22 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=10.395 $Y=2.32
+ $X2=10.525 $Y2=2.405
r155 16 18 22.384 $w=2.58e-07 $l=5.05e-07 $layer=LI1_cond $X=10.395 $Y=2.32
+ $X2=10.395 $Y2=1.815
r156 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=10.16 $Y=2.37
+ $X2=10.16 $Y2=2.655
r157 12 13 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=10.16 $Y=2.28
+ $X2=10.16 $Y2=2.37
r158 11 19 34.2225 $w=3.69e-07 $l=2.17612e-07 $layer=POLY_cond $X=10.16 $Y=1.98
+ $X2=10.282 $Y2=1.815
r159 11 12 116.613 $w=1.8e-07 $l=3e-07 $layer=POLY_cond $X=10.16 $Y=1.98
+ $X2=10.16 $Y2=2.28
r160 7 19 58.6339 $w=3.69e-07 $l=3.89654e-07 $layer=POLY_cond $X=10.115 $Y=1.5
+ $X2=10.282 $Y2=1.815
r161 7 9 471.745 $w=1.5e-07 $l=9.2e-07 $layer=POLY_cond $X=10.115 $Y=1.5
+ $X2=10.115 $Y2=0.58
r162 2 25 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=10.87
+ $Y=2.445 $X2=11.02 $Y2=2.655
r163 1 37 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=10.98
+ $Y=0.37 $X2=11.12 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRBP_1%A_1747_74# 1 2 7 9 10 11 12 14 16 17 19 20
+ 22 23 24 26 27 29 32 40 42 45 47 51 52 56 58 59 61
c180 58 0 8.18376e-20 $X=10.01 $Y=2.425
c181 10 0 1.78926e-19 $X=11.26 $Y=1.02
c182 7 0 1.60243e-20 $X=10.905 $Y=0.87
r183 68 69 4.6235 $w=4.17e-07 $l=4e-08 $layer=POLY_cond $X=11.925 $Y=1.5
+ $X2=11.965 $Y2=1.5
r184 64 65 15.0154 $w=2.6e-07 $l=3.2e-07 $layer=LI1_cond $X=9.69 $Y=1.175
+ $X2=10.01 $Y2=1.175
r185 59 65 4.30428 $w=4.3e-07 $l=1.05119e-07 $layer=LI1_cond $X=10.095 $Y=1.22
+ $X2=10.01 $Y2=1.175
r186 59 61 31.2232 $w=4.28e-07 $l=1.165e-06 $layer=LI1_cond $X=10.095 $Y=1.22
+ $X2=11.26 $Y2=1.22
r187 57 65 3.22376 $w=1.7e-07 $l=2.6e-07 $layer=LI1_cond $X=10.01 $Y=1.435
+ $X2=10.01 $Y2=1.175
r188 57 58 64.5882 $w=1.68e-07 $l=9.9e-07 $layer=LI1_cond $X=10.01 $Y=1.435
+ $X2=10.01 $Y2=2.425
r189 56 64 3.22376 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=9.69 $Y=1.005
+ $X2=9.69 $Y2=1.175
r190 55 56 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=9.69 $Y=0.735
+ $X2=9.69 $Y2=1.005
r191 52 54 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=9.325 $Y=2.59
+ $X2=9.545 $Y2=2.59
r192 51 58 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.925 $Y=2.59
+ $X2=10.01 $Y2=2.425
r193 51 54 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=9.925 $Y=2.59
+ $X2=9.545 $Y2=2.59
r194 47 55 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.605 $Y=0.57
+ $X2=9.69 $Y2=0.735
r195 47 49 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=9.605 $Y=0.57
+ $X2=9.37 $Y2=0.57
r196 43 52 7.17723 $w=3.3e-07 $l=2.13014e-07 $layer=LI1_cond $X=9.215 $Y=2.425
+ $X2=9.325 $Y2=2.59
r197 43 45 26.4538 $w=2.18e-07 $l=5.05e-07 $layer=LI1_cond $X=9.215 $Y=2.425
+ $X2=9.215 $Y2=1.92
r198 38 40 53.8404 $w=1.5e-07 $l=1.05e-07 $layer=POLY_cond $X=11.245 $Y=2.295
+ $X2=11.35 $Y2=2.295
r199 30 42 34.7346 $w=1.65e-07 $l=1.72337e-07 $layer=POLY_cond $X=12.93 $Y=1.355
+ $X2=12.915 $Y2=1.52
r200 30 32 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=12.93 $Y=1.355
+ $X2=12.93 $Y2=0.645
r201 27 29 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=12.915 $Y=2.045
+ $X2=12.915 $Y2=2.54
r202 26 27 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=12.915 $Y=1.955
+ $X2=12.915 $Y2=2.045
r203 25 42 34.7346 $w=1.65e-07 $l=1.65e-07 $layer=POLY_cond $X=12.915 $Y=1.685
+ $X2=12.915 $Y2=1.52
r204 25 26 104.952 $w=1.8e-07 $l=2.7e-07 $layer=POLY_cond $X=12.915 $Y=1.685
+ $X2=12.915 $Y2=1.955
r205 24 69 10.9026 $w=4.17e-07 $l=8.44097e-08 $layer=POLY_cond $X=12.04 $Y=1.52
+ $X2=11.965 $Y2=1.5
r206 23 42 3.90195 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=12.825 $Y=1.52
+ $X2=12.915 $Y2=1.52
r207 23 24 137.266 $w=3.3e-07 $l=7.85e-07 $layer=POLY_cond $X=12.825 $Y=1.52
+ $X2=12.04 $Y2=1.52
r208 20 69 26.8826 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=11.965 $Y=1.235
+ $X2=11.965 $Y2=1.5
r209 20 22 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=11.965 $Y=1.235
+ $X2=11.965 $Y2=0.74
r210 17 68 26.8826 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=11.925 $Y=1.765
+ $X2=11.925 $Y2=1.5
r211 17 19 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=11.925 $Y=1.765
+ $X2=11.925 $Y2=2.4
r212 16 40 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.35 $Y=2.22
+ $X2=11.35 $Y2=2.295
r213 15 68 66.4628 $w=4.17e-07 $l=5.75e-07 $layer=POLY_cond $X=11.35 $Y=1.5
+ $X2=11.925 $Y2=1.5
r214 15 16 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=11.35 $Y=1.685
+ $X2=11.35 $Y2=2.22
r215 12 38 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.245 $Y=2.37
+ $X2=11.245 $Y2=2.295
r216 12 14 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=11.245 $Y=2.37
+ $X2=11.245 $Y2=2.655
r217 11 15 10.4029 $w=4.17e-07 $l=3.06716e-07 $layer=POLY_cond $X=11.26 $Y=1.235
+ $X2=11.35 $Y2=1.5
r218 11 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.26
+ $Y=1.27 $X2=11.26 $Y2=1.27
r219 10 34 182.032 $w=1.5e-07 $l=3.55e-07 $layer=POLY_cond $X=11.26 $Y=0.945
+ $X2=10.905 $Y2=0.945
r220 10 11 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=11.26 $Y=1.02
+ $X2=11.26 $Y2=1.235
r221 7 34 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.905 $Y=0.87
+ $X2=10.905 $Y2=0.945
r222 7 9 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=10.905 $Y=0.87
+ $X2=10.905 $Y2=0.58
r223 2 54 600 $w=1.7e-07 $l=1.06637e-06 $layer=licon1_PDIFF $count=1 $X=9.07
+ $Y=1.735 $X2=9.545 $Y2=2.59
r224 2 45 300 $w=1.7e-07 $l=2.48948e-07 $layer=licon1_PDIFF $count=2 $X=9.07
+ $Y=1.735 $X2=9.22 $Y2=1.92
r225 1 49 182 $w=1.7e-07 $l=7.28166e-07 $layer=licon1_NDIFF $count=1 $X=8.735
+ $Y=0.37 $X2=9.37 $Y2=0.57
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRBP_1%A_2513_424# 1 2 9 11 13 16 20 24 27
r50 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.38
+ $Y=1.465 $X2=13.38 $Y2=1.465
r51 22 27 0.820356 $w=3.3e-07 $l=1.43e-07 $layer=LI1_cond $X=12.855 $Y=1.465
+ $X2=12.712 $Y2=1.465
r52 22 24 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=12.855 $Y=1.465
+ $X2=13.38 $Y2=1.465
r53 18 27 5.82594 $w=2.85e-07 $l=1.65e-07 $layer=LI1_cond $X=12.712 $Y=1.63
+ $X2=12.712 $Y2=1.465
r54 18 20 25.6772 $w=2.83e-07 $l=6.35e-07 $layer=LI1_cond $X=12.712 $Y=1.63
+ $X2=12.712 $Y2=2.265
r55 14 27 5.82594 $w=2.85e-07 $l=1.65e-07 $layer=LI1_cond $X=12.712 $Y=1.3
+ $X2=12.712 $Y2=1.465
r56 14 16 26.486 $w=2.83e-07 $l=6.55e-07 $layer=LI1_cond $X=12.712 $Y=1.3
+ $X2=12.712 $Y2=0.645
r57 11 25 61.4066 $w=2.86e-07 $l=3.26343e-07 $layer=POLY_cond $X=13.435 $Y=1.765
+ $X2=13.38 $Y2=1.465
r58 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=13.435 $Y=1.765
+ $X2=13.435 $Y2=2.4
r59 7 25 38.6549 $w=2.86e-07 $l=1.83916e-07 $layer=POLY_cond $X=13.42 $Y=1.3
+ $X2=13.38 $Y2=1.465
r60 7 9 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=13.42 $Y=1.3 $X2=13.42
+ $Y2=0.74
r61 2 20 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=12.565
+ $Y=2.12 $X2=12.69 $Y2=2.265
r62 1 16 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=12.59
+ $Y=0.37 $X2=12.715 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRBP_1%VPWR 1 2 3 4 5 6 7 8 27 31 35 39 43 49 52
+ 55 59 64 65 67 68 70 71 73 75 84 101 105 110 115 122 123 126 129 132 135 138
c186 2 0 1.19423e-19 $X=3.11 $Y=2.32
r187 138 139 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=3.33
+ $X2=13.2 $Y2=3.33
r188 135 136 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r189 132 133 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r190 129 130 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r191 126 127 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r192 123 139 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=3.33
+ $X2=13.2 $Y2=3.33
r193 122 123 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=3.33
+ $X2=13.68 $Y2=3.33
r194 120 138 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=13.325 $Y=3.33
+ $X2=13.185 $Y2=3.33
r195 120 122 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=13.325 $Y=3.33
+ $X2=13.68 $Y2=3.33
r196 119 139 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=13.2 $Y2=3.33
r197 119 136 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=11.76 $Y2=3.33
r198 118 119 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r199 116 135 10.508 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=11.815 $Y=3.33
+ $X2=11.592 $Y2=3.33
r200 116 118 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=11.815 $Y=3.33
+ $X2=12.72 $Y2=3.33
r201 115 138 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=13.045 $Y=3.33
+ $X2=13.185 $Y2=3.33
r202 115 118 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=13.045 $Y=3.33
+ $X2=12.72 $Y2=3.33
r203 114 136 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=11.76 $Y2=3.33
r204 114 133 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=10.32 $Y2=3.33
r205 113 114 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r206 111 132 8.88104 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=10.65 $Y=3.33
+ $X2=10.477 $Y2=3.33
r207 111 113 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=10.65 $Y=3.33
+ $X2=11.28 $Y2=3.33
r208 110 135 10.508 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=11.37 $Y=3.33
+ $X2=11.592 $Y2=3.33
r209 110 113 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=11.37 $Y=3.33
+ $X2=11.28 $Y2=3.33
r210 109 133 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=10.32 $Y2=3.33
r211 109 130 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=8.4 $Y2=3.33
r212 108 109 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r213 106 129 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.485 $Y=3.33
+ $X2=8.36 $Y2=3.33
r214 106 108 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=8.485 $Y=3.33
+ $X2=8.88 $Y2=3.33
r215 105 132 8.88104 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=10.305 $Y=3.33
+ $X2=10.477 $Y2=3.33
r216 105 108 92.9679 $w=1.68e-07 $l=1.425e-06 $layer=LI1_cond $X=10.305 $Y=3.33
+ $X2=8.88 $Y2=3.33
r217 104 130 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r218 103 104 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r219 101 129 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.235 $Y=3.33
+ $X2=8.36 $Y2=3.33
r220 101 103 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=8.235 $Y=3.33
+ $X2=7.92 $Y2=3.33
r221 96 99 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=5.04 $Y=3.33
+ $X2=6.96 $Y2=3.33
r222 96 97 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r223 94 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r224 93 94 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r225 91 94 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r226 91 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r227 90 93 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.6 $Y=3.33 $X2=4.56
+ $Y2=3.33
r228 90 91 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r229 88 126 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.425 $Y=3.33
+ $X2=3.26 $Y2=3.33
r230 88 90 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.425 $Y=3.33
+ $X2=3.6 $Y2=3.33
r231 87 127 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=3.12 $Y2=3.33
r232 86 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r233 84 126 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.095 $Y=3.33
+ $X2=3.26 $Y2=3.33
r234 84 86 92.3155 $w=1.68e-07 $l=1.415e-06 $layer=LI1_cond $X=3.095 $Y=3.33
+ $X2=1.68 $Y2=3.33
r235 83 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r236 82 83 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r237 79 83 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r238 78 82 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=3.33 $X2=1.2
+ $Y2=3.33
r239 78 79 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r240 75 104 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.92 $Y2=3.33
r241 75 97 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=5.04 $Y2=3.33
r242 75 99 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r243 73 74 5.78802 $w=4.43e-07 $l=1.2e-07 $layer=LI1_cond $X=11.592 $Y=2.815
+ $X2=11.592 $Y2=2.695
r244 70 99 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=7.025 $Y=3.33
+ $X2=6.96 $Y2=3.33
r245 70 71 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=7.025 $Y=3.33
+ $X2=7.145 $Y2=3.33
r246 69 103 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=7.265 $Y=3.33
+ $X2=7.92 $Y2=3.33
r247 69 71 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=7.265 $Y=3.33
+ $X2=7.145 $Y2=3.33
r248 67 93 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=4.705 $Y=3.33
+ $X2=4.56 $Y2=3.33
r249 67 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.705 $Y=3.33
+ $X2=4.87 $Y2=3.33
r250 66 96 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=5.035 $Y=3.33
+ $X2=5.04 $Y2=3.33
r251 66 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.035 $Y=3.33
+ $X2=4.87 $Y2=3.33
r252 64 82 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=1.225 $Y=3.33
+ $X2=1.2 $Y2=3.33
r253 64 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.225 $Y=3.33
+ $X2=1.39 $Y2=3.33
r254 63 86 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=1.555 $Y=3.33
+ $X2=1.68 $Y2=3.33
r255 63 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.555 $Y=3.33
+ $X2=1.39 $Y2=3.33
r256 59 62 17.0809 $w=2.78e-07 $l=4.15e-07 $layer=LI1_cond $X=13.185 $Y=1.985
+ $X2=13.185 $Y2=2.4
r257 57 138 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=13.185 $Y=3.245
+ $X2=13.185 $Y2=3.33
r258 57 62 34.7791 $w=2.78e-07 $l=8.45e-07 $layer=LI1_cond $X=13.185 $Y=3.245
+ $X2=13.185 $Y2=2.4
r259 55 74 28.0595 $w=2.28e-07 $l=5.6e-07 $layer=LI1_cond $X=11.7 $Y=2.135
+ $X2=11.7 $Y2=2.695
r260 52 135 1.76584 $w=4.45e-07 $l=8.5e-08 $layer=LI1_cond $X=11.592 $Y=3.245
+ $X2=11.592 $Y2=3.33
r261 51 73 2.64155 $w=4.43e-07 $l=1.02e-07 $layer=LI1_cond $X=11.592 $Y=2.917
+ $X2=11.592 $Y2=2.815
r262 51 52 8.49441 $w=4.43e-07 $l=3.28e-07 $layer=LI1_cond $X=11.592 $Y=2.917
+ $X2=11.592 $Y2=3.245
r263 47 132 1.03204 $w=3.45e-07 $l=8.5e-08 $layer=LI1_cond $X=10.477 $Y=3.245
+ $X2=10.477 $Y2=3.33
r264 47 49 14.0297 $w=3.43e-07 $l=4.2e-07 $layer=LI1_cond $X=10.477 $Y=3.245
+ $X2=10.477 $Y2=2.825
r265 43 46 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=8.36 $Y=1.88
+ $X2=8.36 $Y2=2.59
r266 41 129 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.36 $Y=3.245
+ $X2=8.36 $Y2=3.33
r267 41 46 30.194 $w=2.48e-07 $l=6.55e-07 $layer=LI1_cond $X=8.36 $Y=3.245
+ $X2=8.36 $Y2=2.59
r268 37 71 0.135687 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=7.145 $Y=3.245
+ $X2=7.145 $Y2=3.33
r269 37 39 31.9323 $w=2.38e-07 $l=6.65e-07 $layer=LI1_cond $X=7.145 $Y=3.245
+ $X2=7.145 $Y2=2.58
r270 33 68 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.87 $Y=3.245
+ $X2=4.87 $Y2=3.33
r271 33 35 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=4.87 $Y=3.245
+ $X2=4.87 $Y2=2.835
r272 29 126 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.26 $Y=3.245
+ $X2=3.26 $Y2=3.33
r273 29 31 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.26 $Y=3.245
+ $X2=3.26 $Y2=2.815
r274 25 65 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.39 $Y=3.245
+ $X2=1.39 $Y2=3.33
r275 25 27 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=1.39 $Y=3.245
+ $X2=1.39 $Y2=2.475
r276 8 62 300 $w=1.7e-07 $l=3.60832e-07 $layer=licon1_PDIFF $count=2 $X=12.99
+ $Y=2.12 $X2=13.175 $Y2=2.4
r277 8 59 600 $w=1.7e-07 $l=2.79464e-07 $layer=licon1_PDIFF $count=1 $X=12.99
+ $Y=2.12 $X2=13.21 $Y2=1.985
r278 7 73 600 $w=1.7e-07 $l=4.65242e-07 $layer=licon1_PDIFF $count=1 $X=11.32
+ $Y=2.445 $X2=11.535 $Y2=2.815
r279 7 55 300 $w=1.7e-07 $l=5.06828e-07 $layer=licon1_PDIFF $count=2 $X=11.32
+ $Y=2.445 $X2=11.695 $Y2=2.135
r280 6 49 600 $w=1.7e-07 $l=4.85386e-07 $layer=licon1_PDIFF $count=1 $X=10.235
+ $Y=2.445 $X2=10.475 $Y2=2.825
r281 5 46 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=8.185
+ $Y=1.735 $X2=8.32 $Y2=2.59
r282 5 43 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=8.185
+ $Y=1.735 $X2=8.32 $Y2=1.88
r283 4 39 600 $w=1.7e-07 $l=3.62319e-07 $layer=licon1_PDIFF $count=1 $X=7.02
+ $Y=2.285 $X2=7.17 $Y2=2.58
r284 3 35 600 $w=1.7e-07 $l=9.47035e-07 $layer=licon1_PDIFF $count=1 $X=4.72
+ $Y=1.96 $X2=4.87 $Y2=2.835
r285 2 31 600 $w=1.7e-07 $l=5.65044e-07 $layer=licon1_PDIFF $count=1 $X=3.11
+ $Y=2.32 $X2=3.26 $Y2=2.815
r286 1 27 300 $w=1.7e-07 $l=2.66458e-07 $layer=licon1_PDIFF $count=2 $X=1.19
+ $Y=2.32 $X2=1.39 $Y2=2.475
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRBP_1%A_409_81# 1 2 3 4 5 16 18 20 23 26 27 28 32
+ 35 37 38 39 40 41 43 45 50 54 57
c172 57 0 7.60406e-20 $X=3.83 $Y=2.475
c173 38 0 1.43931e-19 $X=6.345 $Y=1.285
c174 26 0 1.94423e-19 $X=4.555 $Y=2.52
c175 23 0 1.19423e-19 $X=3.53 $Y=2.33
r176 55 57 15.1867 $w=2.41e-07 $l=3e-07 $layer=LI1_cond $X=3.53 $Y=2.475
+ $X2=3.83 $Y2=2.475
r177 50 52 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=2.435 $Y=0.68
+ $X2=2.435 $Y2=1.005
r178 45 47 0.520034 $w=4.58e-07 $l=2e-08 $layer=LI1_cond $X=2.325 $Y=2.475
+ $X2=2.325 $Y2=2.495
r179 42 43 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=6.43 $Y=1.37
+ $X2=6.43 $Y2=2.045
r180 40 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.345 $Y=2.13
+ $X2=6.43 $Y2=2.045
r181 40 41 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=6.345 $Y=2.13
+ $X2=6.075 $Y2=2.13
r182 38 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.345 $Y=1.285
+ $X2=6.43 $Y2=1.37
r183 38 39 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=6.345 $Y=1.285
+ $X2=5.975 $Y2=1.285
r184 37 60 3.21189 $w=2.5e-07 $l=1.7e-07 $layer=LI1_cond $X=5.95 $Y=2.385
+ $X2=5.95 $Y2=2.555
r185 36 41 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.95 $Y=2.215
+ $X2=6.075 $Y2=2.13
r186 36 37 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=5.95 $Y=2.215
+ $X2=5.95 $Y2=2.385
r187 35 39 6.81835 $w=1.7e-07 $l=1.23386e-07 $layer=LI1_cond $X=5.887 $Y=1.2
+ $X2=5.975 $Y2=1.285
r188 35 58 12.9922 $w=1.73e-07 $l=2.05e-07 $layer=LI1_cond $X=5.887 $Y=1.2
+ $X2=5.887 $Y2=0.995
r189 30 58 5.54545 $w=1.78e-07 $l=9e-08 $layer=LI1_cond $X=5.885 $Y=0.905
+ $X2=5.885 $Y2=0.995
r190 30 32 5.85354 $w=1.78e-07 $l=9.5e-08 $layer=LI1_cond $X=5.885 $Y=0.905
+ $X2=5.885 $Y2=0.81
r191 28 60 3.74091 $w=1.95e-07 $l=1.57321e-07 $layer=LI1_cond $X=5.825 $Y=2.482
+ $X2=5.95 $Y2=2.555
r192 28 29 67.1142 $w=1.93e-07 $l=1.18e-06 $layer=LI1_cond $X=5.825 $Y=2.482
+ $X2=4.645 $Y2=2.482
r193 27 57 21.6506 $w=2.41e-07 $l=4.41928e-07 $layer=LI1_cond $X=4.25 $Y=2.52
+ $X2=3.83 $Y2=2.475
r194 26 29 5.46269 $w=2.01e-07 $l=1.07331e-07 $layer=LI1_cond $X=4.555 $Y=2.52
+ $X2=4.645 $Y2=2.482
r195 26 27 16.9136 $w=1.98e-07 $l=3.05e-07 $layer=LI1_cond $X=4.555 $Y=2.52
+ $X2=4.25 $Y2=2.52
r196 23 55 2.78154 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=3.53 $Y=2.33
+ $X2=3.53 $Y2=2.475
r197 22 23 80.8984 $w=1.68e-07 $l=1.24e-06 $layer=LI1_cond $X=3.53 $Y=1.09
+ $X2=3.53 $Y2=2.33
r198 20 55 5.37722 $w=2.41e-07 $l=8.5e-08 $layer=LI1_cond $X=3.445 $Y=2.475
+ $X2=3.53 $Y2=2.475
r199 20 54 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=3.445 $Y=2.475
+ $X2=2.945 $Y2=2.475
r200 19 52 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.6 $Y=1.005
+ $X2=2.435 $Y2=1.005
r201 18 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.445 $Y=1.005
+ $X2=3.53 $Y2=1.09
r202 18 19 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=3.445 $Y=1.005
+ $X2=2.6 $Y2=1.005
r203 17 47 5.34566 $w=2.1e-07 $l=2.3e-07 $layer=LI1_cond $X=2.555 $Y=2.495
+ $X2=2.325 $Y2=2.495
r204 16 54 5.98033 $w=2.08e-07 $l=1.05e-07 $layer=LI1_cond $X=2.84 $Y=2.495
+ $X2=2.945 $Y2=2.495
r205 16 17 15.0519 $w=2.08e-07 $l=2.85e-07 $layer=LI1_cond $X=2.84 $Y=2.495
+ $X2=2.555 $Y2=2.495
r206 5 60 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=5.765
+ $Y=2.285 $X2=5.91 $Y2=2.495
r207 4 57 300 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=2 $X=3.68
+ $Y=2.32 $X2=3.83 $Y2=2.475
r208 3 45 300 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=2 $X=2.11
+ $Y=2.32 $X2=2.26 $Y2=2.475
r209 2 32 182 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_NDIFF $count=1 $X=5.755
+ $Y=0.595 $X2=5.88 $Y2=0.81
r210 1 50 182 $w=1.7e-07 $l=5.09264e-07 $layer=licon1_NDIFF $count=1 $X=2.045
+ $Y=0.405 $X2=2.435 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRBP_1%Q_N 1 2 7 8 9 10 11 12 13
r21 13 40 1.3969 $w=3.28e-07 $l=4e-08 $layer=LI1_cond $X=12.18 $Y=2.775
+ $X2=12.18 $Y2=2.815
r22 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=12.18 $Y=2.405
+ $X2=12.18 $Y2=2.775
r23 12 34 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=12.18 $Y=2.405
+ $X2=12.18 $Y2=2.055
r24 11 34 0.69845 $w=3.28e-07 $l=2e-08 $layer=LI1_cond $X=12.18 $Y=2.035
+ $X2=12.18 $Y2=2.055
r25 10 11 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=12.18 $Y=1.665
+ $X2=12.18 $Y2=2.035
r26 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=12.18 $Y=1.295
+ $X2=12.18 $Y2=1.665
r27 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=12.18 $Y=0.925
+ $X2=12.18 $Y2=1.295
r28 7 8 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=12.18 $Y=0.515
+ $X2=12.18 $Y2=0.925
r29 2 40 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=12
+ $Y=1.84 $X2=12.15 $Y2=2.815
r30 2 34 400 $w=1.7e-07 $l=2.80134e-07 $layer=licon1_PDIFF $count=1 $X=12
+ $Y=1.84 $X2=12.15 $Y2=2.055
r31 1 7 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=12.04
+ $Y=0.37 $X2=12.18 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRBP_1%Q 1 2 9 10 11 12 13 28 32 43
r20 41 43 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=13.75 $Y=1.13
+ $X2=13.75 $Y2=1.82
r21 29 32 1.02897 $w=2.78e-07 $l=2.5e-08 $layer=LI1_cond $X=13.695 $Y=1.96
+ $X2=13.695 $Y2=1.985
r22 21 28 0.726197 $w=3.63e-07 $l=2.3e-08 $layer=LI1_cond $X=13.652 $Y=0.948
+ $X2=13.652 $Y2=0.925
r23 12 13 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=13.695 $Y=2.405
+ $X2=13.695 $Y2=2.775
r24 11 29 0.205793 $w=2.78e-07 $l=5e-09 $layer=LI1_cond $X=13.695 $Y=1.955
+ $X2=13.695 $Y2=1.96
r25 11 43 7.32213 $w=2.78e-07 $l=1.35e-07 $layer=LI1_cond $X=13.695 $Y=1.955
+ $X2=13.695 $Y2=1.82
r26 11 12 15.0229 $w=2.78e-07 $l=3.65e-07 $layer=LI1_cond $X=13.695 $Y=2.04
+ $X2=13.695 $Y2=2.405
r27 11 32 2.26373 $w=2.78e-07 $l=5.5e-08 $layer=LI1_cond $X=13.695 $Y=2.04
+ $X2=13.695 $Y2=1.985
r28 10 41 8.08227 $w=3.63e-07 $l=1.51e-07 $layer=LI1_cond $X=13.652 $Y=0.979
+ $X2=13.652 $Y2=1.13
r29 10 21 0.978787 $w=3.63e-07 $l=3.1e-08 $layer=LI1_cond $X=13.652 $Y=0.979
+ $X2=13.652 $Y2=0.948
r30 10 28 0.978787 $w=3.63e-07 $l=3.1e-08 $layer=LI1_cond $X=13.652 $Y=0.894
+ $X2=13.652 $Y2=0.925
r31 9 10 11.9665 $w=3.63e-07 $l=3.79e-07 $layer=LI1_cond $X=13.652 $Y=0.515
+ $X2=13.652 $Y2=0.894
r32 2 13 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=13.51
+ $Y=1.84 $X2=13.66 $Y2=2.815
r33 2 32 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=13.51
+ $Y=1.84 $X2=13.66 $Y2=1.985
r34 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=13.495
+ $Y=0.37 $X2=13.635 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRBP_1%VGND 1 2 3 4 5 6 7 24 28 32 36 38 42 45 46
+ 47 49 54 63 67 75 82 83 86 89 93 99 103 109
c138 83 0 6.07903e-20 $X=13.68 $Y=0
c139 28 0 1.58089e-19 $X=3.715 $Y=0.565
r140 109 110 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.2 $Y=0
+ $X2=13.2 $Y2=0
r141 104 110 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=13.2 $Y2=0
r142 103 106 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=11.675 $Y=0
+ $X2=11.675 $Y2=0.325
r143 103 104 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r144 99 100 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r145 93 96 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=7.595 $Y=0
+ $X2=7.595 $Y2=0.325
r146 93 94 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r147 89 90 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r148 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r149 83 110 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=0
+ $X2=13.2 $Y2=0
r150 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=0
+ $X2=13.68 $Y2=0
r151 80 109 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.29 $Y=0
+ $X2=13.205 $Y2=0
r152 80 82 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=13.29 $Y=0
+ $X2=13.68 $Y2=0
r153 79 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=11.76 $Y2=0
r154 79 100 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=10.32 $Y2=0
r155 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r156 76 99 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.495 $Y=0
+ $X2=10.33 $Y2=0
r157 76 78 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=10.495 $Y=0
+ $X2=11.28 $Y2=0
r158 75 103 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.51 $Y=0
+ $X2=11.675 $Y2=0
r159 75 78 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=11.51 $Y=0
+ $X2=11.28 $Y2=0
r160 74 100 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=10.32 $Y2=0
r161 73 74 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=9.84 $Y=0
+ $X2=9.84 $Y2=0
r162 71 74 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=7.92 $Y=0
+ $X2=9.84 $Y2=0
r163 71 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=7.44
+ $Y2=0
r164 70 73 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=7.92 $Y=0 $X2=9.84
+ $Y2=0
r165 70 71 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r166 68 93 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.76 $Y=0 $X2=7.595
+ $Y2=0
r167 68 70 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=7.76 $Y=0 $X2=7.92
+ $Y2=0
r168 67 99 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.165 $Y=0
+ $X2=10.33 $Y2=0
r169 67 73 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=10.165 $Y=0
+ $X2=9.84 $Y2=0
r170 65 66 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r171 63 93 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.43 $Y=0 $X2=7.595
+ $Y2=0
r172 63 65 155.925 $w=1.68e-07 $l=2.39e-06 $layer=LI1_cond $X=7.43 $Y=0 $X2=5.04
+ $Y2=0
r173 62 66 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r174 62 90 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=3.6
+ $Y2=0
r175 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r176 59 89 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=3.88 $Y=0 $X2=3.735
+ $Y2=0
r177 59 61 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.88 $Y=0 $X2=4.56
+ $Y2=0
r178 58 90 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=3.6
+ $Y2=0
r179 58 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r180 57 58 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r181 55 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=0.71
+ $Y2=0
r182 55 57 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=1.2
+ $Y2=0
r183 54 89 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=3.59 $Y=0 $X2=3.735
+ $Y2=0
r184 54 57 155.925 $w=1.68e-07 $l=2.39e-06 $layer=LI1_cond $X=3.59 $Y=0 $X2=1.2
+ $Y2=0
r185 52 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r186 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r187 49 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.71
+ $Y2=0
r188 49 51 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0
+ $X2=0.24 $Y2=0
r189 47 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r190 47 66 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6.96 $Y=0
+ $X2=5.04 $Y2=0
r191 45 61 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=4.705 $Y=0
+ $X2=4.56 $Y2=0
r192 45 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.705 $Y=0 $X2=4.87
+ $Y2=0
r193 44 65 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=5.035 $Y=0 $X2=5.04
+ $Y2=0
r194 44 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.035 $Y=0 $X2=4.87
+ $Y2=0
r195 40 109 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.205 $Y=0.085
+ $X2=13.205 $Y2=0
r196 40 42 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=13.205 $Y=0.085
+ $X2=13.205 $Y2=0.515
r197 39 103 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.84 $Y=0
+ $X2=11.675 $Y2=0
r198 38 109 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.12 $Y=0
+ $X2=13.205 $Y2=0
r199 38 39 83.508 $w=1.68e-07 $l=1.28e-06 $layer=LI1_cond $X=13.12 $Y=0
+ $X2=11.84 $Y2=0
r200 34 99 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.33 $Y=0.085
+ $X2=10.33 $Y2=0
r201 34 36 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=10.33 $Y=0.085
+ $X2=10.33 $Y2=0.58
r202 30 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.87 $Y=0.085
+ $X2=4.87 $Y2=0
r203 30 32 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=4.87 $Y=0.085
+ $X2=4.87 $Y2=0.585
r204 26 89 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.735 $Y=0.085
+ $X2=3.735 $Y2=0
r205 26 28 19.0749 $w=2.88e-07 $l=4.8e-07 $layer=LI1_cond $X=3.735 $Y=0.085
+ $X2=3.735 $Y2=0.565
r206 22 86 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0
r207 22 24 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0.58
r208 7 42 91 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_NDIFF $count=2 $X=13.005
+ $Y=0.37 $X2=13.205 $Y2=0.515
r209 6 106 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=11.535
+ $Y=0.18 $X2=11.675 $Y2=0.325
r210 5 36 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=10.19
+ $Y=0.37 $X2=10.33 $Y2=0.58
r211 4 96 182 $w=1.7e-07 $l=3.63731e-07 $layer=licon1_NDIFF $count=1 $X=7.375
+ $Y=0.595 $X2=7.595 $Y2=0.325
r212 3 32 182 $w=1.7e-07 $l=2.04939e-07 $layer=licon1_NDIFF $count=1 $X=4.67
+ $Y=0.595 $X2=4.87 $Y2=0.585
r213 2 28 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=3.575
+ $Y=0.405 $X2=3.715 $Y2=0.565
r214 1 24 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRBP_1%noxref_25 1 2 9 11 12 13
r33 13 16 7.40856 $w=3.48e-07 $l=2.25e-07 $layer=LI1_cond $X=3.235 $Y=0.34
+ $X2=3.235 $Y2=0.565
r34 11 13 4.974 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=3.06 $Y=0.34 $X2=3.235
+ $Y2=0.34
r35 11 12 111.235 $w=1.68e-07 $l=1.705e-06 $layer=LI1_cond $X=3.06 $Y=0.34
+ $X2=1.355 $Y2=0.34
r36 7 12 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.23 $Y=0.425
+ $X2=1.355 $Y2=0.34
r37 7 9 8.98906 $w=2.48e-07 $l=1.95e-07 $layer=LI1_cond $X=1.23 $Y=0.425
+ $X2=1.23 $Y2=0.62
r38 2 16 182 $w=1.7e-07 $l=2.22711e-07 $layer=licon1_NDIFF $count=1 $X=3.115
+ $Y=0.405 $X2=3.265 $Y2=0.565
r39 1 9 182 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_NDIFF $count=1 $X=1.125
+ $Y=0.405 $X2=1.27 $Y2=0.62
.ends

