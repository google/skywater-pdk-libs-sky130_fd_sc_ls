* File: sky130_fd_sc_ls__o2111ai_4.spice
* Created: Wed Sep  2 11:17:04 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__o2111ai_4.pex.spice"
.subckt sky130_fd_sc_ls__o2111ai_4  VNB VPB D1 C1 B1 A1 A2 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A2	A2
* A1	A1
* B1	B1
* C1	C1
* D1	D1
* VPB	VPB
* VNB	VNB
MM1008 N_A_27_74#_M1008_d N_D1_M1008_g N_Y_M1008_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.1295 PD=2.05 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75000.2
+ SB=75003.3 A=0.111 P=1.78 MULT=1
MM1010 N_A_27_74#_M1010_d N_D1_M1010_g N_Y_M1008_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.7
+ SB=75002.8 A=0.111 P=1.78 MULT=1
MM1024 N_A_27_74#_M1010_d N_D1_M1024_g N_Y_M1024_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75002.4 A=0.111 P=1.78 MULT=1
MM1030 N_A_27_74#_M1030_d N_D1_M1030_g N_Y_M1024_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.6
+ SB=75001.9 A=0.111 P=1.78 MULT=1
MM1006 N_A_27_74#_M1030_d N_C1_M1006_g N_A_472_74#_M1006_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002
+ SB=75001.5 A=0.111 P=1.78 MULT=1
MM1018 N_A_27_74#_M1018_d N_C1_M1018_g N_A_472_74#_M1006_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75002.4 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1022 N_A_27_74#_M1018_d N_C1_M1022_g N_A_472_74#_M1022_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75002.9 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1033 N_A_27_74#_M1033_d N_C1_M1033_g N_A_472_74#_M1022_s VNB NSHORT L=0.15
+ W=0.74 AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75003.3 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1007 N_A_472_74#_M1007_d N_B1_M1007_g N_A_841_74#_M1007_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75005.2 A=0.111 P=1.78 MULT=1
MM1012 N_A_472_74#_M1007_d N_B1_M1012_g N_A_841_74#_M1012_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75004.8 A=0.111 P=1.78 MULT=1
MM1021 N_A_472_74#_M1021_d N_B1_M1021_g N_A_841_74#_M1012_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.1 SB=75004.4 A=0.111 P=1.78 MULT=1
MM1027 N_A_472_74#_M1021_d N_B1_M1027_g N_A_841_74#_M1027_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75001.5 SB=75003.9 A=0.111 P=1.78 MULT=1
MM1002 N_A_841_74#_M1027_s N_A1_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1295 AS=0.1295 PD=1.09 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75002
+ SB=75003.4 A=0.111 P=1.78 MULT=1
MM1005 N_A_841_74#_M1005_d N_A1_M1005_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.5
+ SB=75002.9 A=0.111 P=1.78 MULT=1
MM1009 N_A_841_74#_M1005_d N_A1_M1009_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.9
+ SB=75002.5 A=0.111 P=1.78 MULT=1
MM1017 N_A_841_74#_M1017_d N_A1_M1017_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75003.4
+ SB=75002.1 A=0.111 P=1.78 MULT=1
MM1001 N_A_841_74#_M1017_d N_A2_M1001_g N_VGND_M1001_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75003.8
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1013 N_A_841_74#_M1013_d N_A2_M1013_g N_VGND_M1001_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1332 AS=0.1295 PD=1.1 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75004.3
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1015 N_A_841_74#_M1013_d N_A2_M1015_g N_VGND_M1015_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1332 AS=0.1036 PD=1.1 PS=1.02 NRD=12.972 NRS=0 M=1 R=4.93333 SA=75004.8
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1025 N_A_841_74#_M1025_d N_A2_M1025_g N_VGND_M1015_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75005.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1028 N_VPWR_M1028_d N_D1_M1028_g N_Y_M1028_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.224 AS=1.176 PD=1.52 PS=4.34 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75001 SB=75003.1 A=0.168 P=2.54 MULT=1
MM1032 N_VPWR_M1028_d N_D1_M1032_g N_Y_M1032_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.224 AS=0.168 PD=1.52 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75001.5 SB=75002.5 A=0.168 P=2.54 MULT=1
MM1003 N_VPWR_M1003_d N_C1_M1003_g N_Y_M1032_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.4032 AS=0.168 PD=1.84 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002 SB=75002.1 A=0.168 P=2.54 MULT=1
MM1004 N_VPWR_M1003_d N_C1_M1004_g N_Y_M1004_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.4032 AS=0.168 PD=1.84 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.8 SB=75001.2 A=0.168 P=2.54 MULT=1
MM1014 N_VPWR_M1014_d N_B1_M1014_g N_Y_M1004_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.224 AS=0.168 PD=1.52 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75003.3 SB=75000.8 A=0.168 P=2.54 MULT=1
MM1019 N_VPWR_M1014_d N_B1_M1019_g N_Y_M1019_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.224 AS=0.3304 PD=1.52 PS=2.83 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75003.8 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1000 N_A_954_368#_M1000_d N_A1_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.15
+ W=1.12 AD=1.5848 AS=0.1764 PD=5.07 PS=1.435 NRD=2.6201 NRS=4.3931 M=1
+ R=7.46667 SA=75001.3 SB=75003.5 A=0.168 P=2.54 MULT=1
MM1016 N_A_954_368#_M1016_d N_A1_M1016_g N_VPWR_M1000_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.1764 PD=1.42 PS=1.435 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.8 SB=75003.1 A=0.168 P=2.54 MULT=1
MM1023 N_A_954_368#_M1016_d N_A1_M1023_g N_VPWR_M1023_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.3 SB=75002.6 A=0.168 P=2.54 MULT=1
MM1026 N_A_954_368#_M1026_d N_A1_M1026_g N_VPWR_M1023_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.1764 AS=0.168 PD=1.435 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.7 SB=75002.2 A=0.168 P=2.54 MULT=1
MM1011 N_A_954_368#_M1026_d N_A2_M1011_g N_Y_M1011_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.1764 AS=0.1876 PD=1.435 PS=1.455 NRD=4.3931 NRS=7.8997 M=1 R=7.46667
+ SA=75003.2 SB=75001.7 A=0.168 P=2.54 MULT=1
MM1020 N_A_954_368#_M1020_d N_A2_M1020_g N_Y_M1011_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.196 AS=0.1876 PD=1.47 PS=1.455 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75003.7 SB=75001.2 A=0.168 P=2.54 MULT=1
MM1029 N_A_954_368#_M1020_d N_A2_M1029_g N_Y_M1029_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.196 AS=0.196 PD=1.47 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75004.2 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1031 N_A_954_368#_M1031_d N_A2_M1031_g N_Y_M1029_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.196 PD=2.83 PS=1.47 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75004.7 SB=75000.2 A=0.168 P=2.54 MULT=1
DX34_noxref VNB VPB NWDIODE A=19.4556 P=24.64
*
.include "sky130_fd_sc_ls__o2111ai_4.pxi.spice"
*
.ends
*
*
