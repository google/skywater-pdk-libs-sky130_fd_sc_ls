* File: sky130_fd_sc_ls__nand2b_1.pxi.spice
* Created: Wed Sep  2 11:11:43 2020
* 
x_PM_SKY130_FD_SC_LS__NAND2B_1%A_N N_A_N_M1002_g N_A_N_c_45_n N_A_N_M1003_g A_N
+ A_N N_A_N_c_44_n PM_SKY130_FD_SC_LS__NAND2B_1%A_N
x_PM_SKY130_FD_SC_LS__NAND2B_1%B N_B_c_74_n N_B_M1001_g N_B_M1000_g B N_B_c_76_n
+ PM_SKY130_FD_SC_LS__NAND2B_1%B
x_PM_SKY130_FD_SC_LS__NAND2B_1%A_27_112# N_A_27_112#_M1002_s N_A_27_112#_M1003_s
+ N_A_27_112#_M1005_g N_A_27_112#_c_110_n N_A_27_112#_M1004_g
+ N_A_27_112#_c_111_n N_A_27_112#_c_112_n N_A_27_112#_c_113_n
+ N_A_27_112#_c_125_n N_A_27_112#_c_117_n N_A_27_112#_c_118_n
+ N_A_27_112#_c_114_n N_A_27_112#_c_115_n PM_SKY130_FD_SC_LS__NAND2B_1%A_27_112#
x_PM_SKY130_FD_SC_LS__NAND2B_1%VPWR N_VPWR_M1003_d N_VPWR_M1004_d N_VPWR_c_179_n
+ N_VPWR_c_180_n N_VPWR_c_181_n N_VPWR_c_182_n VPWR N_VPWR_c_183_n
+ N_VPWR_c_178_n N_VPWR_c_185_n PM_SKY130_FD_SC_LS__NAND2B_1%VPWR
x_PM_SKY130_FD_SC_LS__NAND2B_1%Y N_Y_M1005_d N_Y_M1001_d N_Y_c_210_n N_Y_c_207_n
+ N_Y_c_208_n N_Y_c_209_n Y Y N_Y_c_214_n PM_SKY130_FD_SC_LS__NAND2B_1%Y
x_PM_SKY130_FD_SC_LS__NAND2B_1%VGND N_VGND_M1002_d N_VGND_c_241_n VGND
+ N_VGND_c_242_n N_VGND_c_243_n N_VGND_c_244_n N_VGND_c_245_n
+ PM_SKY130_FD_SC_LS__NAND2B_1%VGND
cc_1 VNB N_A_N_M1002_g 0.031967f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.835
cc_2 VNB A_N 0.0177819f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_3 VNB N_A_N_c_44_n 0.0658387f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.532
cc_4 VNB N_B_c_74_n 0.0271918f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.3
cc_5 VNB N_B_M1000_g 0.0274125f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.26
cc_6 VNB N_B_c_76_n 0.00182951f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.532
cc_7 VNB N_A_27_112#_M1005_g 0.0248499f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_8 VNB N_A_27_112#_c_110_n 0.0344014f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_27_112#_c_111_n 0.0188303f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.465
cc_10 VNB N_A_27_112#_c_112_n 0.0153597f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.54
cc_11 VNB N_A_27_112#_c_113_n 0.00869634f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.54
cc_12 VNB N_A_27_112#_c_114_n 0.00981133f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_112#_c_115_n 0.00161243f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_VPWR_c_178_n 0.103974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_Y_c_207_n 0.027835f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_Y_c_208_n 0.0250664f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.532
cc_17 VNB N_Y_c_209_n 0.0158601f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.465
cc_18 VNB N_VGND_c_241_n 0.0155608f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.26
cc_19 VNB N_VGND_c_242_n 0.0182319f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_243_n 0.0364261f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.54
cc_21 VNB N_VGND_c_244_n 0.175015f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_245_n 0.0126977f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.54
cc_23 VPB N_A_N_c_45_n 0.0222398f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_24 VPB A_N 0.0113319f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_25 VPB N_A_N_c_44_n 0.00793031f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.532
cc_26 VPB N_B_c_74_n 0.0286805f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.3
cc_27 VPB N_B_c_76_n 0.0029888f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.532
cc_28 VPB N_A_27_112#_c_110_n 0.0247857f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_29 VPB N_A_27_112#_c_117_n 0.00136663f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_30 VPB N_A_27_112#_c_118_n 0.0333833f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_31 VPB N_VPWR_c_179_n 0.0194035f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_32 VPB N_VPWR_c_180_n 0.0221346f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.54
cc_33 VPB N_VPWR_c_181_n 0.0221383f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.54
cc_34 VPB N_VPWR_c_182_n 0.00623744f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.54
cc_35 VPB N_VPWR_c_183_n 0.0126445f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_36 VPB N_VPWR_c_178_n 0.0738319f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_37 VPB N_VPWR_c_185_n 0.0264241f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_38 VPB N_Y_c_210_n 0.0169104f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.26
cc_39 VPB N_Y_c_208_n 0.0314126f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.532
cc_40 VPB Y 0.00319648f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.465
cc_41 N_A_N_c_45_n N_B_c_74_n 0.0205137f $X=0.505 $Y=1.765 $X2=-0.19 $Y2=-0.245
cc_42 A_N N_B_c_74_n 0.0026624f $X=0.635 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_43 N_A_N_c_44_n N_B_c_74_n 0.0177315f $X=0.505 $Y=1.532 $X2=-0.19 $Y2=-0.245
cc_44 N_A_N_M1002_g N_B_M1000_g 0.00900688f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_45 A_N N_B_M1000_g 0.00113012f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_46 N_A_N_c_44_n N_B_M1000_g 0.00121331f $X=0.505 $Y=1.532 $X2=0 $Y2=0
cc_47 A_N N_B_c_76_n 0.0350659f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_48 N_A_N_c_44_n N_B_c_76_n 5.61835e-19 $X=0.505 $Y=1.532 $X2=0 $Y2=0
cc_49 N_A_N_M1002_g N_A_27_112#_c_111_n 0.0020078f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_50 N_A_N_M1002_g N_A_27_112#_c_112_n 0.015445f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_51 A_N N_A_27_112#_c_112_n 0.0348645f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_52 N_A_N_c_44_n N_A_27_112#_c_112_n 0.00556316f $X=0.505 $Y=1.532 $X2=0 $Y2=0
cc_53 A_N N_A_27_112#_c_113_n 0.0226786f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_54 N_A_N_c_44_n N_A_27_112#_c_113_n 0.00613776f $X=0.505 $Y=1.532 $X2=0 $Y2=0
cc_55 N_A_N_c_45_n N_A_27_112#_c_125_n 0.0128974f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_56 A_N N_A_27_112#_c_125_n 0.0283317f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_57 N_A_N_c_44_n N_A_27_112#_c_125_n 8.10409e-19 $X=0.505 $Y=1.532 $X2=0 $Y2=0
cc_58 N_A_N_c_45_n N_A_27_112#_c_118_n 0.00957412f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_59 A_N N_A_27_112#_c_118_n 0.0267404f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_60 N_A_N_c_44_n N_A_27_112#_c_118_n 0.0015638f $X=0.505 $Y=1.532 $X2=0 $Y2=0
cc_61 N_A_N_c_45_n N_VPWR_c_179_n 0.00737625f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_62 N_A_N_c_45_n N_VPWR_c_178_n 0.00462577f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_63 N_A_N_c_45_n N_VPWR_c_185_n 0.00393873f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_64 N_A_N_M1002_g N_VGND_c_241_n 0.010935f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_65 N_A_N_M1002_g N_VGND_c_242_n 0.003901f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_66 N_A_N_M1002_g N_VGND_c_244_n 0.00425985f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_67 N_B_M1000_g N_A_27_112#_M1005_g 0.0373434f $X=1.27 $Y=0.74 $X2=0 $Y2=0
cc_68 N_B_c_74_n N_A_27_112#_c_110_n 0.0717248f $X=1.175 $Y=1.765 $X2=0 $Y2=0
cc_69 N_B_c_76_n N_A_27_112#_c_110_n 6.73156e-19 $X=1.18 $Y=1.515 $X2=0 $Y2=0
cc_70 N_B_c_74_n N_A_27_112#_c_112_n 0.00118672f $X=1.175 $Y=1.765 $X2=0 $Y2=0
cc_71 N_B_M1000_g N_A_27_112#_c_112_n 0.0156214f $X=1.27 $Y=0.74 $X2=0 $Y2=0
cc_72 N_B_c_76_n N_A_27_112#_c_112_n 0.0202397f $X=1.18 $Y=1.515 $X2=0 $Y2=0
cc_73 N_B_c_74_n N_A_27_112#_c_125_n 0.012472f $X=1.175 $Y=1.765 $X2=0 $Y2=0
cc_74 N_B_c_76_n N_A_27_112#_c_125_n 0.0210863f $X=1.18 $Y=1.515 $X2=0 $Y2=0
cc_75 N_B_c_74_n N_A_27_112#_c_117_n 0.00349194f $X=1.175 $Y=1.765 $X2=0 $Y2=0
cc_76 N_B_c_74_n N_A_27_112#_c_118_n 7.20757e-19 $X=1.175 $Y=1.765 $X2=0 $Y2=0
cc_77 N_B_c_74_n N_A_27_112#_c_114_n 0.00330428f $X=1.175 $Y=1.765 $X2=0 $Y2=0
cc_78 N_B_c_76_n N_A_27_112#_c_114_n 0.0341497f $X=1.18 $Y=1.515 $X2=0 $Y2=0
cc_79 N_B_M1000_g N_A_27_112#_c_115_n 0.00330428f $X=1.27 $Y=0.74 $X2=0 $Y2=0
cc_80 N_B_c_74_n N_VPWR_c_179_n 0.00711266f $X=1.175 $Y=1.765 $X2=0 $Y2=0
cc_81 N_B_c_74_n N_VPWR_c_180_n 6.06947e-19 $X=1.175 $Y=1.765 $X2=0 $Y2=0
cc_82 N_B_c_74_n N_VPWR_c_181_n 0.00291513f $X=1.175 $Y=1.765 $X2=0 $Y2=0
cc_83 N_B_c_74_n N_VPWR_c_178_n 0.00364726f $X=1.175 $Y=1.765 $X2=0 $Y2=0
cc_84 N_B_c_74_n Y 0.014114f $X=1.175 $Y=1.765 $X2=0 $Y2=0
cc_85 N_B_c_74_n N_Y_c_214_n 0.00587989f $X=1.175 $Y=1.765 $X2=0 $Y2=0
cc_86 N_B_M1000_g N_VGND_c_241_n 0.0172792f $X=1.27 $Y=0.74 $X2=0 $Y2=0
cc_87 N_B_M1000_g N_VGND_c_243_n 0.00383152f $X=1.27 $Y=0.74 $X2=0 $Y2=0
cc_88 N_B_M1000_g N_VGND_c_244_n 0.0075725f $X=1.27 $Y=0.74 $X2=0 $Y2=0
cc_89 N_A_27_112#_c_125_n N_VPWR_M1003_d 0.0187431f $X=1.515 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_90 N_A_27_112#_c_125_n N_VPWR_c_179_n 0.0213973f $X=1.515 $Y=2.035 $X2=0
+ $Y2=0
cc_91 N_A_27_112#_c_118_n N_VPWR_c_179_n 0.0271251f $X=0.28 $Y=2.115 $X2=0 $Y2=0
cc_92 N_A_27_112#_c_110_n N_VPWR_c_180_n 0.00833347f $X=1.675 $Y=1.765 $X2=0
+ $Y2=0
cc_93 N_A_27_112#_c_110_n N_VPWR_c_181_n 0.00413917f $X=1.675 $Y=1.765 $X2=0
+ $Y2=0
cc_94 N_A_27_112#_c_110_n N_VPWR_c_178_n 0.00818241f $X=1.675 $Y=1.765 $X2=0
+ $Y2=0
cc_95 N_A_27_112#_c_118_n N_VPWR_c_178_n 0.00997343f $X=0.28 $Y=2.115 $X2=0
+ $Y2=0
cc_96 N_A_27_112#_c_118_n N_VPWR_c_185_n 0.0066794f $X=0.28 $Y=2.115 $X2=0 $Y2=0
cc_97 N_A_27_112#_c_125_n N_Y_M1001_d 0.00930652f $X=1.515 $Y=2.035 $X2=0 $Y2=0
cc_98 N_A_27_112#_c_117_n N_Y_M1001_d 0.00135982f $X=1.6 $Y=1.95 $X2=0 $Y2=0
cc_99 N_A_27_112#_c_110_n N_Y_c_210_n 0.0181072f $X=1.675 $Y=1.765 $X2=0 $Y2=0
cc_100 N_A_27_112#_c_125_n N_Y_c_210_n 0.00643277f $X=1.515 $Y=2.035 $X2=0 $Y2=0
cc_101 N_A_27_112#_c_114_n N_Y_c_210_n 0.00488923f $X=1.75 $Y=1.465 $X2=0 $Y2=0
cc_102 N_A_27_112#_M1005_g N_Y_c_207_n 0.0221957f $X=1.66 $Y=0.74 $X2=0 $Y2=0
cc_103 N_A_27_112#_M1005_g N_Y_c_208_n 0.00292854f $X=1.66 $Y=0.74 $X2=0 $Y2=0
cc_104 N_A_27_112#_c_110_n N_Y_c_208_n 0.0210207f $X=1.675 $Y=1.765 $X2=0 $Y2=0
cc_105 N_A_27_112#_c_125_n N_Y_c_208_n 0.00712937f $X=1.515 $Y=2.035 $X2=0 $Y2=0
cc_106 N_A_27_112#_c_117_n N_Y_c_208_n 0.0120524f $X=1.6 $Y=1.95 $X2=0 $Y2=0
cc_107 N_A_27_112#_c_114_n N_Y_c_208_n 0.0251716f $X=1.75 $Y=1.465 $X2=0 $Y2=0
cc_108 N_A_27_112#_c_115_n N_Y_c_208_n 0.00637596f $X=1.715 $Y=1.3 $X2=0 $Y2=0
cc_109 N_A_27_112#_c_110_n N_Y_c_209_n 4.59055e-19 $X=1.675 $Y=1.765 $X2=0 $Y2=0
cc_110 N_A_27_112#_c_112_n N_Y_c_209_n 0.0142393f $X=1.515 $Y=1.045 $X2=0 $Y2=0
cc_111 N_A_27_112#_c_114_n N_Y_c_209_n 0.0049152f $X=1.75 $Y=1.465 $X2=0 $Y2=0
cc_112 N_A_27_112#_c_110_n Y 0.00283699f $X=1.675 $Y=1.765 $X2=0 $Y2=0
cc_113 N_A_27_112#_c_125_n N_Y_c_214_n 0.0307866f $X=1.515 $Y=2.035 $X2=0 $Y2=0
cc_114 N_A_27_112#_c_112_n N_VGND_M1002_d 0.00761754f $X=1.515 $Y=1.045
+ $X2=-0.19 $Y2=-0.245
cc_115 N_A_27_112#_M1005_g N_VGND_c_241_n 0.00188096f $X=1.66 $Y=0.74 $X2=0
+ $Y2=0
cc_116 N_A_27_112#_c_111_n N_VGND_c_241_n 0.0112176f $X=0.28 $Y=0.835 $X2=0
+ $Y2=0
cc_117 N_A_27_112#_c_112_n N_VGND_c_241_n 0.0447655f $X=1.515 $Y=1.045 $X2=0
+ $Y2=0
cc_118 N_A_27_112#_c_111_n N_VGND_c_242_n 0.00651231f $X=0.28 $Y=0.835 $X2=0
+ $Y2=0
cc_119 N_A_27_112#_M1005_g N_VGND_c_243_n 0.00461464f $X=1.66 $Y=0.74 $X2=0
+ $Y2=0
cc_120 N_A_27_112#_M1005_g N_VGND_c_244_n 0.00913279f $X=1.66 $Y=0.74 $X2=0
+ $Y2=0
cc_121 N_A_27_112#_c_111_n N_VGND_c_244_n 0.00849993f $X=0.28 $Y=0.835 $X2=0
+ $Y2=0
cc_122 N_A_27_112#_c_112_n A_269_74# 0.00485986f $X=1.515 $Y=1.045 $X2=-0.19
+ $Y2=-0.245
cc_123 N_VPWR_M1004_d N_Y_c_210_n 0.0109667f $X=1.75 $Y=1.84 $X2=0 $Y2=0
cc_124 N_VPWR_c_180_n N_Y_c_210_n 0.0206146f $X=1.9 $Y=2.815 $X2=0 $Y2=0
cc_125 N_VPWR_c_179_n Y 0.021048f $X=0.82 $Y=2.455 $X2=0 $Y2=0
cc_126 N_VPWR_c_180_n Y 0.0132475f $X=1.9 $Y=2.815 $X2=0 $Y2=0
cc_127 N_VPWR_c_181_n Y 0.0209023f $X=1.735 $Y=3.33 $X2=0 $Y2=0
cc_128 N_VPWR_c_178_n Y 0.0169394f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_129 N_Y_c_207_n N_VGND_c_241_n 0.0128668f $X=1.94 $Y=0.515 $X2=0 $Y2=0
cc_130 N_Y_c_207_n N_VGND_c_243_n 0.0177591f $X=1.94 $Y=0.515 $X2=0 $Y2=0
cc_131 N_Y_c_207_n N_VGND_c_244_n 0.0146995f $X=1.94 $Y=0.515 $X2=0 $Y2=0
