* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__bufinv_8 A VGND VNB VPB VPWR Y
M1000 Y a_183_48# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=1.4896e+12p pd=1.162e+07u as=2.184e+12p ps=1.734e+07u
M1001 Y a_183_48# VGND VNB nshort w=740000u l=150000u
+  ad=8.954e+11p pd=8.34e+06u as=1.5392e+12p ps=1.304e+07u
M1002 VPWR a_183_48# Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VGND a_183_48# Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_183_48# a_27_368# VGND VNB nshort w=740000u l=150000u
+  ad=4.292e+11p pd=4.12e+06u as=0p ps=0u
M1005 VGND a_183_48# Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y a_183_48# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR a_183_48# Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_183_48# a_27_368# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y a_183_48# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 Y a_183_48# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND a_183_48# Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND a_27_368# a_183_48# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR A a_27_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.304e+11p ps=2.83e+06u
M1014 a_183_48# a_27_368# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=6.664e+11p pd=5.67e+06u as=0p ps=0u
M1015 Y a_183_48# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR a_183_48# Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 Y a_183_48# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR a_27_368# a_183_48# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR a_183_48# Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND a_183_48# Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND A a_27_368# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1022 Y a_183_48# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_183_48# a_27_368# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
