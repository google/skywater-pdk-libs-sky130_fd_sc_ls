* File: sky130_fd_sc_ls__a32oi_1.pxi.spice
* Created: Fri Aug 28 13:00:35 2020
* 
x_PM_SKY130_FD_SC_LS__A32OI_1%B2 N_B2_c_46_n N_B2_M1006_g N_B2_c_47_n
+ N_B2_M1002_g B2 PM_SKY130_FD_SC_LS__A32OI_1%B2
x_PM_SKY130_FD_SC_LS__A32OI_1%B1 N_B1_c_67_n N_B1_M1008_g N_B1_c_68_n
+ N_B1_M1004_g B1 PM_SKY130_FD_SC_LS__A32OI_1%B1
x_PM_SKY130_FD_SC_LS__A32OI_1%A1 N_A1_c_95_n N_A1_M1009_g N_A1_c_96_n
+ N_A1_M1005_g A1 PM_SKY130_FD_SC_LS__A32OI_1%A1
x_PM_SKY130_FD_SC_LS__A32OI_1%A2 N_A2_c_124_n N_A2_M1007_g N_A2_c_125_n
+ N_A2_M1001_g A2 A2 A2 PM_SKY130_FD_SC_LS__A32OI_1%A2
x_PM_SKY130_FD_SC_LS__A32OI_1%A3 N_A3_c_159_n N_A3_M1000_g N_A3_c_160_n
+ N_A3_M1003_g A3 PM_SKY130_FD_SC_LS__A32OI_1%A3
x_PM_SKY130_FD_SC_LS__A32OI_1%A_27_368# N_A_27_368#_M1006_s N_A_27_368#_M1004_d
+ N_A_27_368#_M1001_d N_A_27_368#_c_183_n N_A_27_368#_c_184_n
+ N_A_27_368#_c_185_n N_A_27_368#_c_195_n N_A_27_368#_c_196_n
+ N_A_27_368#_c_197_n N_A_27_368#_c_186_n N_A_27_368#_c_187_n
+ N_A_27_368#_c_202_n PM_SKY130_FD_SC_LS__A32OI_1%A_27_368#
x_PM_SKY130_FD_SC_LS__A32OI_1%Y N_Y_M1008_d N_Y_M1006_d N_Y_c_232_n N_Y_c_246_n
+ N_Y_c_233_n N_Y_c_234_n N_Y_c_236_n Y N_Y_c_238_n
+ PM_SKY130_FD_SC_LS__A32OI_1%Y
x_PM_SKY130_FD_SC_LS__A32OI_1%VPWR N_VPWR_M1009_d N_VPWR_M1003_d N_VPWR_c_281_n
+ N_VPWR_c_282_n VPWR N_VPWR_c_283_n N_VPWR_c_284_n N_VPWR_c_285_n
+ N_VPWR_c_280_n PM_SKY130_FD_SC_LS__A32OI_1%VPWR
x_PM_SKY130_FD_SC_LS__A32OI_1%VGND N_VGND_M1002_s N_VGND_M1000_d N_VGND_c_320_n
+ N_VGND_c_321_n N_VGND_c_322_n N_VGND_c_323_n VGND N_VGND_c_324_n
+ N_VGND_c_325_n PM_SKY130_FD_SC_LS__A32OI_1%VGND
cc_1 VNB N_B2_c_46_n 0.0677571f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_2 VNB N_B2_c_47_n 0.0199632f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.22
cc_3 VNB B2 0.00806923f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_B1_c_67_n 0.0229989f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_5 VNB N_B1_c_68_n 0.048622f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.22
cc_6 VNB B1 0.00758946f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_7 VNB N_A1_c_95_n 0.0498088f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_8 VNB N_A1_c_96_n 0.0231454f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.22
cc_9 VNB A1 0.00429394f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_10 VNB N_A2_c_124_n 0.0174586f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_11 VNB N_A2_c_125_n 0.0380544f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.22
cc_12 VNB A2 0.00819917f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_13 VNB N_A3_c_159_n 0.0223315f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_14 VNB N_A3_c_160_n 0.0445355f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.22
cc_15 VNB A3 0.0219295f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_16 VNB N_Y_c_232_n 0.0100996f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_Y_c_233_n 0.00159849f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_Y_c_234_n 0.00778594f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.385
cc_19 VNB N_VPWR_c_280_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_320_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_21 VNB N_VGND_c_321_n 0.0377474f $X=-0.19 $Y=-0.245 $X2=0.355 $Y2=1.385
cc_22 VNB N_VGND_c_322_n 0.0128247f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.385
cc_23 VNB N_VGND_c_323_n 0.0344702f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_324_n 0.0649785f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_325_n 0.215051f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VPB N_B2_c_46_n 0.0293876f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_27 VPB N_B1_c_68_n 0.0226345f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.22
cc_28 VPB N_A1_c_95_n 0.0253782f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_29 VPB N_A2_c_125_n 0.0250856f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.22
cc_30 VPB N_A3_c_160_n 0.0281228f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.22
cc_31 VPB N_A_27_368#_c_183_n 0.0436022f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=1.295
cc_32 VPB N_A_27_368#_c_184_n 0.00667982f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_33 VPB N_A_27_368#_c_185_n 0.00983167f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_34 VPB N_A_27_368#_c_186_n 0.0102405f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_35 VPB N_A_27_368#_c_187_n 0.00243101f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_36 VPB N_Y_c_232_n 0.00132726f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_37 VPB N_Y_c_236_n 0.00462141f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_38 VPB Y 0.0101401f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_39 VPB N_Y_c_238_n 0.00893879f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_40 VPB N_VPWR_c_281_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_41 VPB N_VPWR_c_282_n 0.0564565f $X=-0.19 $Y=1.66 $X2=0.355 $Y2=1.385
cc_42 VPB N_VPWR_c_283_n 0.0425054f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=1.385
cc_43 VPB N_VPWR_c_284_n 0.0183219f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_44 VPB N_VPWR_c_285_n 0.018879f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_45 VPB N_VPWR_c_280_n 0.0590517f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 N_B2_c_47_n N_B1_c_67_n 0.0321121f $X=0.52 $Y=1.22 $X2=-0.19 $Y2=-0.245
cc_47 N_B2_c_46_n N_B1_c_68_n 0.0666062f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_48 N_B2_c_46_n N_A_27_368#_c_183_n 0.0163614f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_49 B2 N_A_27_368#_c_183_n 0.0197435f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_50 N_B2_c_46_n N_A_27_368#_c_184_n 0.011054f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_51 N_B2_c_46_n N_A_27_368#_c_185_n 0.00262441f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_52 N_B2_c_47_n N_Y_c_232_n 0.00939717f $X=0.52 $Y=1.22 $X2=0 $Y2=0
cc_53 B2 N_Y_c_232_n 0.0279669f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_54 N_B2_c_47_n N_Y_c_233_n 0.00269193f $X=0.52 $Y=1.22 $X2=0 $Y2=0
cc_55 N_B2_c_46_n N_Y_c_236_n 0.00380161f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_56 N_B2_c_46_n N_VPWR_c_283_n 0.00278257f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_57 N_B2_c_46_n N_VPWR_c_280_n 0.0035783f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_58 N_B2_c_46_n N_VGND_c_321_n 0.00217022f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_59 N_B2_c_47_n N_VGND_c_321_n 0.00533858f $X=0.52 $Y=1.22 $X2=0 $Y2=0
cc_60 B2 N_VGND_c_321_n 0.0263177f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_61 N_B2_c_47_n N_VGND_c_324_n 0.00460063f $X=0.52 $Y=1.22 $X2=0 $Y2=0
cc_62 N_B2_c_47_n N_VGND_c_325_n 0.00910551f $X=0.52 $Y=1.22 $X2=0 $Y2=0
cc_63 N_B1_c_68_n N_A1_c_95_n 0.049683f $X=1.005 $Y=1.765 $X2=-0.19 $Y2=-0.245
cc_64 B1 N_A1_c_95_n 0.0020937f $X=1.115 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_65 N_B1_c_68_n A1 3.96911e-19 $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_66 B1 A1 0.0253469f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_67 N_B1_c_68_n N_A_27_368#_c_183_n 7.61749e-19 $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_68 N_B1_c_68_n N_A_27_368#_c_184_n 0.014165f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_69 N_B1_c_67_n N_Y_c_232_n 0.00474996f $X=0.91 $Y=1.22 $X2=0 $Y2=0
cc_70 N_B1_c_68_n N_Y_c_232_n 0.00378083f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_71 B1 N_Y_c_232_n 0.0279522f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_72 N_B1_c_68_n N_Y_c_246_n 0.0123778f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_73 N_B1_c_67_n N_Y_c_234_n 0.0228512f $X=0.91 $Y=1.22 $X2=0 $Y2=0
cc_74 N_B1_c_68_n N_Y_c_234_n 0.00194662f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_75 B1 N_Y_c_234_n 0.0284419f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_76 N_B1_c_68_n N_Y_c_236_n 0.00750061f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_77 N_B1_c_68_n Y 6.16746e-19 $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_78 N_B1_c_68_n N_Y_c_238_n 0.0147928f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_79 B1 N_Y_c_238_n 0.0268776f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_80 N_B1_c_68_n N_VPWR_c_283_n 0.00278271f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_81 N_B1_c_68_n N_VPWR_c_285_n 2.50377e-19 $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_82 N_B1_c_68_n N_VPWR_c_280_n 0.00355672f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_83 N_B1_c_67_n N_VGND_c_324_n 0.00291649f $X=0.91 $Y=1.22 $X2=0 $Y2=0
cc_84 N_B1_c_67_n N_VGND_c_325_n 0.0036383f $X=0.91 $Y=1.22 $X2=0 $Y2=0
cc_85 N_A1_c_96_n N_A2_c_124_n 0.033517f $X=1.88 $Y=1.22 $X2=-0.19 $Y2=-0.245
cc_86 A1 N_A2_c_124_n 3.10488e-19 $X=1.595 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_87 N_A1_c_95_n N_A2_c_125_n 0.0522235f $X=1.615 $Y=1.765 $X2=0 $Y2=0
cc_88 N_A1_c_96_n A2 0.0118388f $X=1.88 $Y=1.22 $X2=0 $Y2=0
cc_89 A1 A2 0.0277288f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_90 N_A1_c_95_n N_A_27_368#_c_184_n 0.00180441f $X=1.615 $Y=1.765 $X2=0 $Y2=0
cc_91 N_A1_c_95_n N_A_27_368#_c_195_n 0.00530604f $X=1.615 $Y=1.765 $X2=0 $Y2=0
cc_92 N_A1_c_95_n N_A_27_368#_c_196_n 0.00711821f $X=1.615 $Y=1.765 $X2=0 $Y2=0
cc_93 N_A1_c_95_n N_A_27_368#_c_197_n 0.0141783f $X=1.615 $Y=1.765 $X2=0 $Y2=0
cc_94 N_A1_c_95_n N_Y_c_246_n 7.14972e-19 $X=1.615 $Y=1.765 $X2=0 $Y2=0
cc_95 N_A1_c_95_n N_Y_c_234_n 0.00179345f $X=1.615 $Y=1.765 $X2=0 $Y2=0
cc_96 N_A1_c_96_n N_Y_c_234_n 0.00905028f $X=1.88 $Y=1.22 $X2=0 $Y2=0
cc_97 A1 N_Y_c_234_n 0.0237588f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_98 N_A1_c_95_n Y 0.0246832f $X=1.615 $Y=1.765 $X2=0 $Y2=0
cc_99 N_A1_c_95_n N_Y_c_238_n 0.00582717f $X=1.615 $Y=1.765 $X2=0 $Y2=0
cc_100 A1 N_Y_c_238_n 0.0257356f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_101 N_A1_c_95_n N_VPWR_c_283_n 0.00415318f $X=1.615 $Y=1.765 $X2=0 $Y2=0
cc_102 N_A1_c_95_n N_VPWR_c_285_n 0.00797106f $X=1.615 $Y=1.765 $X2=0 $Y2=0
cc_103 N_A1_c_95_n N_VPWR_c_280_n 0.00415839f $X=1.615 $Y=1.765 $X2=0 $Y2=0
cc_104 N_A1_c_96_n N_VGND_c_324_n 0.00433162f $X=1.88 $Y=1.22 $X2=0 $Y2=0
cc_105 N_A1_c_96_n N_VGND_c_325_n 0.00822327f $X=1.88 $Y=1.22 $X2=0 $Y2=0
cc_106 N_A2_c_124_n N_A3_c_159_n 0.0241574f $X=2.27 $Y=1.22 $X2=-0.19 $Y2=-0.245
cc_107 A2 N_A3_c_159_n 0.00950494f $X=2.075 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_108 N_A2_c_125_n N_A3_c_160_n 0.0391014f $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_109 A2 N_A3_c_160_n 4.18785e-19 $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_110 N_A2_c_125_n A3 0.00121116f $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_111 A2 A3 0.0223908f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_112 N_A2_c_125_n N_A_27_368#_c_197_n 0.0143515f $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_113 N_A2_c_125_n N_A_27_368#_c_186_n 0.0121655f $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_114 A2 N_A_27_368#_c_186_n 0.0035826f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_115 N_A2_c_125_n N_A_27_368#_c_187_n 2.71519e-19 $X=2.405 $Y=1.765 $X2=0
+ $Y2=0
cc_116 N_A2_c_125_n N_A_27_368#_c_202_n 5.73569e-19 $X=2.405 $Y=1.765 $X2=0
+ $Y2=0
cc_117 N_A2_c_124_n N_Y_c_234_n 9.06958e-19 $X=2.27 $Y=1.22 $X2=0 $Y2=0
cc_118 A2 N_Y_c_234_n 0.0401943f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_119 N_A2_c_125_n Y 0.00697427f $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_120 A2 Y 0.0202848f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_121 N_A2_c_125_n N_VPWR_c_284_n 0.00415318f $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_122 N_A2_c_125_n N_VPWR_c_285_n 0.00811382f $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_123 N_A2_c_125_n N_VPWR_c_280_n 0.00414564f $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_124 N_A2_c_124_n N_VGND_c_323_n 0.00141413f $X=2.27 $Y=1.22 $X2=0 $Y2=0
cc_125 A2 N_VGND_c_323_n 0.025354f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_126 N_A2_c_124_n N_VGND_c_324_n 0.00303293f $X=2.27 $Y=1.22 $X2=0 $Y2=0
cc_127 A2 N_VGND_c_324_n 0.0132057f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_128 N_A2_c_124_n N_VGND_c_325_n 0.00372643f $X=2.27 $Y=1.22 $X2=0 $Y2=0
cc_129 A2 N_VGND_c_325_n 0.0159188f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_130 A2 A_391_74# 0.00780801f $X=2.075 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_131 A2 A_469_74# 0.0100426f $X=2.075 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_132 N_A3_c_160_n N_A_27_368#_c_186_n 0.0066684f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_133 A3 N_A_27_368#_c_186_n 0.00167971f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_134 N_A3_c_160_n N_A_27_368#_c_187_n 0.00584689f $X=2.855 $Y=1.765 $X2=0
+ $Y2=0
cc_135 N_A3_c_160_n N_A_27_368#_c_202_n 0.00183357f $X=2.855 $Y=1.765 $X2=0
+ $Y2=0
cc_136 N_A3_c_160_n N_VPWR_c_282_n 0.0109613f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_137 A3 N_VPWR_c_282_n 0.014999f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_138 N_A3_c_160_n N_VPWR_c_284_n 0.00445602f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_139 N_A3_c_160_n N_VPWR_c_285_n 4.26569e-19 $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_140 N_A3_c_160_n N_VPWR_c_280_n 0.00861168f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_141 N_A3_c_159_n N_VGND_c_323_n 0.0159756f $X=2.84 $Y=1.22 $X2=0 $Y2=0
cc_142 N_A3_c_160_n N_VGND_c_323_n 0.00111834f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_143 A3 N_VGND_c_323_n 0.0259407f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_144 N_A3_c_159_n N_VGND_c_324_n 0.00383152f $X=2.84 $Y=1.22 $X2=0 $Y2=0
cc_145 N_A3_c_159_n N_VGND_c_325_n 0.00758792f $X=2.84 $Y=1.22 $X2=0 $Y2=0
cc_146 N_A_27_368#_c_184_n N_Y_M1006_d 0.00250873f $X=1.115 $Y=2.99 $X2=0 $Y2=0
cc_147 N_A_27_368#_c_184_n N_Y_c_246_n 0.018923f $X=1.115 $Y=2.99 $X2=0 $Y2=0
cc_148 N_A_27_368#_c_183_n N_Y_c_236_n 0.0035248f $X=0.28 $Y=1.985 $X2=0 $Y2=0
cc_149 N_A_27_368#_c_195_n Y 0.00733332f $X=1.28 $Y=2.49 $X2=0 $Y2=0
cc_150 N_A_27_368#_c_197_n Y 0.0483435f $X=2.465 $Y=2.405 $X2=0 $Y2=0
cc_151 N_A_27_368#_c_186_n Y 0.0121588f $X=2.63 $Y=1.985 $X2=0 $Y2=0
cc_152 N_A_27_368#_M1004_d N_Y_c_238_n 0.00424779f $X=1.08 $Y=1.84 $X2=0 $Y2=0
cc_153 N_A_27_368#_c_195_n N_Y_c_238_n 0.0240481f $X=1.28 $Y=2.49 $X2=0 $Y2=0
cc_154 N_A_27_368#_c_197_n N_Y_c_238_n 0.00295908f $X=2.465 $Y=2.405 $X2=0 $Y2=0
cc_155 N_A_27_368#_c_197_n N_VPWR_M1009_d 0.0137245f $X=2.465 $Y=2.405 $X2=-0.19
+ $Y2=1.66
cc_156 N_A_27_368#_c_186_n N_VPWR_c_282_n 0.0335221f $X=2.63 $Y=1.985 $X2=0
+ $Y2=0
cc_157 N_A_27_368#_c_187_n N_VPWR_c_282_n 0.0324512f $X=2.63 $Y=2.815 $X2=0
+ $Y2=0
cc_158 N_A_27_368#_c_202_n N_VPWR_c_282_n 0.0121024f $X=2.63 $Y=2.405 $X2=0
+ $Y2=0
cc_159 N_A_27_368#_c_184_n N_VPWR_c_283_n 0.0659319f $X=1.115 $Y=2.99 $X2=0
+ $Y2=0
cc_160 N_A_27_368#_c_185_n N_VPWR_c_283_n 0.0235712f $X=0.445 $Y=2.99 $X2=0
+ $Y2=0
cc_161 N_A_27_368#_c_187_n N_VPWR_c_284_n 0.0123628f $X=2.63 $Y=2.815 $X2=0
+ $Y2=0
cc_162 N_A_27_368#_c_184_n N_VPWR_c_285_n 0.0119072f $X=1.115 $Y=2.99 $X2=0
+ $Y2=0
cc_163 N_A_27_368#_c_196_n N_VPWR_c_285_n 0.0158719f $X=1.28 $Y=2.815 $X2=0
+ $Y2=0
cc_164 N_A_27_368#_c_197_n N_VPWR_c_285_n 0.043859f $X=2.465 $Y=2.405 $X2=0
+ $Y2=0
cc_165 N_A_27_368#_c_187_n N_VPWR_c_285_n 0.0141508f $X=2.63 $Y=2.815 $X2=0
+ $Y2=0
cc_166 N_A_27_368#_c_184_n N_VPWR_c_280_n 0.0367158f $X=1.115 $Y=2.99 $X2=0
+ $Y2=0
cc_167 N_A_27_368#_c_185_n N_VPWR_c_280_n 0.0127563f $X=0.445 $Y=2.99 $X2=0
+ $Y2=0
cc_168 N_A_27_368#_c_197_n N_VPWR_c_280_n 0.0124275f $X=2.465 $Y=2.405 $X2=0
+ $Y2=0
cc_169 N_A_27_368#_c_187_n N_VPWR_c_280_n 0.0101999f $X=2.63 $Y=2.815 $X2=0
+ $Y2=0
cc_170 N_A_27_368#_c_202_n N_VPWR_c_280_n 0.00181649f $X=2.63 $Y=2.405 $X2=0
+ $Y2=0
cc_171 Y N_VPWR_M1009_d 0.0125184f $X=2.075 $Y=1.95 $X2=-0.19 $Y2=-0.245
cc_172 N_Y_c_233_n N_VGND_c_321_n 0.0284176f $X=0.785 $Y=0.68 $X2=0 $Y2=0
cc_173 N_Y_c_233_n N_VGND_c_324_n 0.00758556f $X=0.785 $Y=0.68 $X2=0 $Y2=0
cc_174 N_Y_c_234_n N_VGND_c_324_n 0.0457898f $X=1.665 $Y=0.495 $X2=0 $Y2=0
cc_175 N_Y_c_233_n N_VGND_c_325_n 0.00627867f $X=0.785 $Y=0.68 $X2=0 $Y2=0
cc_176 N_Y_c_234_n N_VGND_c_325_n 0.037678f $X=1.665 $Y=0.495 $X2=0 $Y2=0
