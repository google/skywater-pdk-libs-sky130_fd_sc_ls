* File: sky130_fd_sc_ls__decaphe_6.pex.spice
* Created: Fri Aug 28 13:12:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__DECAPHE_6%VGND 1 7 8 9 12 15 26 29
r17 28 29 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r18 26 28 0.245473 $w=9.94e-07 $l=2e-08 $layer=LI1_cond $X=2.62 $Y=0.497
+ $X2=2.64 $Y2=0.497
r19 22 23 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r20 20 22 3.66319 $w=1.532e-06 $l=4.6e-07 $layer=LI1_cond $X=0.26 $Y=0.757
+ $X2=0.72 $Y2=0.757
r21 18 23 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r22 17 20 0.159269 $w=1.532e-06 $l=2e-08 $layer=LI1_cond $X=0.24 $Y=0.757
+ $X2=0.26 $Y2=0.757
r23 17 18 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r24 13 22 1.55287 $w=1.532e-06 $l=1.95e-07 $layer=LI1_cond $X=0.915 $Y=0.757
+ $X2=0.72 $Y2=0.757
r25 12 15 25.2123 $w=1.82e-06 $l=1.18579e-06 $layer=POLY_cond $X=0.915 $Y=1.515
+ $X2=1.44 $Y2=2.467
r26 12 13 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.915
+ $Y=1.515 $X2=0.915 $Y2=1.515
r27 9 29 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.44 $Y=0 $X2=2.64
+ $Y2=0
r28 9 23 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=0.72
+ $Y2=0
r29 8 13 2.95945 $w=1.532e-06 $l=3.88844e-07 $layer=LI1_cond $X=1.195 $Y=0.497
+ $X2=0.915 $Y2=0.757
r30 7 26 4.9262 $w=1.165e-06 $l=4.42e-07 $layer=LI1_cond $X=2.178 $Y=0.497
+ $X2=2.62 $Y2=0.497
r31 7 8 10.2941 $w=1.163e-06 $l=9.83e-07 $layer=LI1_cond $X=2.178 $Y=0.497
+ $X2=1.195 $Y2=0.497
r32 1 26 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=2.485
+ $Y=0.235 $X2=2.62 $Y2=0.38
r33 1 20 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=2.485
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LS__DECAPHE_6%VPWR 1 9 10 15 17 29 37
r17 29 32 0.13762 $w=1.773e-06 $l=2e-08 $layer=LI1_cond $X=2.62 $Y=2.332
+ $X2=2.64 $Y2=2.332
r18 22 37 0.00529514 $w=2.88e-06 $l=1.22e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.44 $Y2=3.208
r19 22 32 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r20 21 24 0.13762 $w=1.773e-06 $l=2e-08 $layer=LI1_cond $X=0.24 $Y=2.332
+ $X2=0.26 $Y2=2.332
r21 21 22 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r22 18 29 2.16751 $w=1.773e-06 $l=3.15e-07 $layer=LI1_cond $X=2.305 $Y=2.332
+ $X2=2.62 $Y2=2.332
r23 17 18 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.305
+ $Y=1.335 $X2=2.305 $Y2=1.335
r24 14 18 4.67908 $w=1.773e-06 $l=6.8e-07 $layer=LI1_cond $X=1.625 $Y=2.332
+ $X2=2.305 $Y2=2.332
r25 14 24 9.39256 $w=1.773e-06 $l=1.365e-06 $layer=LI1_cond $X=1.625 $Y=2.332
+ $X2=0.26 $Y2=2.332
r26 13 17 24.0843 $w=1.395e-06 $l=6.8e-07 $layer=POLY_cond $X=1.625 $Y=0.802
+ $X2=2.305 $Y2=0.802
r27 13 15 9.23771 $w=1.395e-06 $l=1.65e-07 $layer=POLY_cond $X=1.625 $Y=0.802
+ $X2=1.46 $Y2=0.802
r28 13 14 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.625
+ $Y=1.335 $X2=1.625 $Y2=1.335
r29 10 37 4.34028e-05 $w=2.88e-06 $l=1e-09 $layer=MET1_cond $X=1.44 $Y=3.207
+ $X2=1.44 $Y2=3.208
r30 9 15 0.931401 $w=1.035e-06 $l=2e-08 $layer=POLY_cond $X=1.44 $Y=0.622
+ $X2=1.46 $Y2=0.622
r31 1 29 400 $w=1.7e-07 $l=1.17556e-06 $layer=licon1_PDIFF $count=1 $X=2.485
+ $Y=1.84 $X2=2.62 $Y2=2.95
r32 1 29 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.485
+ $Y=1.84 $X2=2.62 $Y2=1.985
r33 1 24 400 $w=1.7e-07 $l=1.17083e-06 $layer=licon1_PDIFF $count=1 $X=2.485
+ $Y=1.84 $X2=0.26 $Y2=2.95
r34 1 24 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=2.485
+ $Y=1.84 $X2=0.26 $Y2=1.985
.ends

