* File: sky130_fd_sc_ls__o21ba_1.pex.spice
* Created: Wed Sep  2 11:18:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__O21BA_1%A1 2 5 6 8 9 10 14 16
r29 14 16 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.395 $Y=1.295
+ $X2=0.395 $Y2=1.13
r30 9 10 10.033 $w=4.23e-07 $l=3.7e-07 $layer=LI1_cond $X=0.337 $Y=1.295
+ $X2=0.337 $Y2=1.665
r31 9 14 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.385
+ $Y=1.295 $X2=0.385 $Y2=1.295
r32 6 8 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.505 $Y=1.885
+ $X2=0.505 $Y2=2.46
r33 5 16 141.387 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=0.495 $Y=0.69
+ $X2=0.495 $Y2=1.13
r34 2 6 43.3633 $w=2.89e-07 $l=3.10161e-07 $layer=POLY_cond $X=0.395 $Y=1.625
+ $X2=0.505 $Y2=1.885
r35 1 14 1.64869 $w=3.5e-07 $l=1e-08 $layer=POLY_cond $X=0.395 $Y=1.305
+ $X2=0.395 $Y2=1.295
r36 1 2 52.7581 $w=3.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.395 $Y=1.305
+ $X2=0.395 $Y2=1.625
.ends

.subckt PM_SKY130_FD_SC_LS__O21BA_1%A2 1 3 6 8 9 10 11 15
r39 10 11 9.21977 $w=4.78e-07 $l=3.7e-07 $layer=LI1_cond $X=1.075 $Y=1.295
+ $X2=1.075 $Y2=1.665
r40 10 15 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1 $Y=1.295
+ $X2=1 $Y2=1.295
r41 9 15 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1 $Y=1.635 $X2=1
+ $Y2=1.295
r42 8 15 42.4377 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1 $Y=1.13 $X2=1
+ $Y2=1.295
r43 6 8 141.387 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=1.065 $Y=0.69
+ $X2=1.065 $Y2=1.13
r44 1 9 43.19 $w=2.79e-07 $l=2.85044e-07 $layer=POLY_cond $X=0.925 $Y=1.885
+ $X2=1 $Y2=1.635
r45 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.925 $Y=1.885
+ $X2=0.925 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_LS__O21BA_1%A_281_244# 1 2 8 9 11 14 18 20 22 23 26 28
+ 30 34 37
r61 31 34 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.22 $Y=0.845
+ $X2=2.555 $Y2=0.845
r62 26 28 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=2.305 $Y=1.985
+ $X2=2.52 $Y2=1.985
r63 24 31 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.22 $Y=1.01
+ $X2=2.22 $Y2=0.845
r64 24 30 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=2.22 $Y=1.01
+ $X2=2.22 $Y2=1.22
r65 23 37 29.847 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.14 $Y=1.385
+ $X2=1.975 $Y2=1.385
r66 22 30 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.14 $Y=1.385
+ $X2=2.14 $Y2=1.22
r67 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.14
+ $Y=1.385 $X2=2.14 $Y2=1.385
r68 20 26 6.81649 $w=3.3e-07 $l=2.33345e-07 $layer=LI1_cond $X=2.14 $Y=1.82
+ $X2=2.305 $Y2=1.985
r69 20 22 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=2.14 $Y=1.82
+ $X2=2.14 $Y2=1.385
r70 17 18 2.30962 $w=2.9e-07 $l=9e-08 $layer=POLY_cond $X=1.585 $Y=1.365
+ $X2=1.495 $Y2=1.365
r71 17 37 80.672 $w=2.9e-07 $l=3.9e-07 $layer=POLY_cond $X=1.585 $Y=1.365
+ $X2=1.975 $Y2=1.365
r72 12 18 31.696 $w=1.65e-07 $l=1.52315e-07 $layer=POLY_cond $X=1.51 $Y=1.22
+ $X2=1.495 $Y2=1.365
r73 12 14 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.51 $Y=1.22
+ $X2=1.51 $Y2=0.69
r74 9 11 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.495 $Y=1.885
+ $X2=1.495 $Y2=2.46
r75 8 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.495 $Y=1.795 $X2=1.495
+ $Y2=1.885
r76 7 18 31.696 $w=1.65e-07 $l=1.45e-07 $layer=POLY_cond $X=1.495 $Y=1.51
+ $X2=1.495 $Y2=1.365
r77 7 8 110.782 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=1.495 $Y=1.51
+ $X2=1.495 $Y2=1.795
r78 2 28 600 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_PDIFF $count=1 $X=2.305
+ $Y=1.84 $X2=2.52 $Y2=1.985
r79 1 34 182 $w=1.7e-07 $l=4.81871e-07 $layer=licon1_NDIFF $count=1 $X=2.195
+ $Y=0.56 $X2=2.555 $Y2=0.845
.ends

.subckt PM_SKY130_FD_SC_LS__O21BA_1%B1_N 1 3 4 6 7
c31 1 0 9.60317e-20 $X=2.75 $Y=1.765
r32 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.68
+ $Y=1.385 $X2=2.68 $Y2=1.385
r33 7 11 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=2.68 $Y=1.295 $X2=2.68
+ $Y2=1.385
r34 4 10 38.9026 $w=2.7e-07 $l=2.05122e-07 $layer=POLY_cond $X=2.77 $Y=1.22
+ $X2=2.68 $Y2=1.385
r35 4 6 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=2.77 $Y=1.22 $X2=2.77
+ $Y2=0.835
r36 1 10 77.2841 $w=2.7e-07 $l=4.13521e-07 $layer=POLY_cond $X=2.75 $Y=1.765
+ $X2=2.68 $Y2=1.385
r37 1 3 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.75 $Y=1.765 $X2=2.75
+ $Y2=2.26
.ends

.subckt PM_SKY130_FD_SC_LS__O21BA_1%A_200_392# 1 2 7 9 12 18 21 22 25 27 31 32
+ 36
r80 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.25
+ $Y=1.485 $X2=3.25 $Y2=1.485
r81 33 36 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=3.14 $Y=1.485
+ $X2=3.25 $Y2=1.485
r82 30 31 7.80118 $w=5.18e-07 $l=8.5e-08 $layer=LI1_cond $X=1.7 $Y=2.23
+ $X2=1.785 $Y2=2.23
r83 27 30 11.0407 $w=5.18e-07 $l=4.8e-07 $layer=LI1_cond $X=1.22 $Y=2.23 $X2=1.7
+ $Y2=2.23
r84 24 33 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.14 $Y=1.65
+ $X2=3.14 $Y2=1.485
r85 24 25 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.14 $Y=1.65
+ $X2=3.14 $Y2=2.32
r86 22 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.055 $Y=2.405
+ $X2=3.14 $Y2=2.32
r87 22 31 82.8556 $w=1.68e-07 $l=1.27e-06 $layer=LI1_cond $X=3.055 $Y=2.405
+ $X2=1.785 $Y2=2.405
r88 21 30 7.40362 $w=1.7e-07 $l=2.6e-07 $layer=LI1_cond $X=1.7 $Y=1.97 $X2=1.7
+ $Y2=2.23
r89 21 32 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=1.7 $Y=1.97 $X2=1.7
+ $Y2=1.03
r90 16 32 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.78 $Y=0.865
+ $X2=1.78 $Y2=1.03
r91 16 18 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=1.78 $Y=0.865
+ $X2=1.78 $Y2=0.515
r92 10 37 38.561 $w=2.98e-07 $l=2.03101e-07 $layer=POLY_cond $X=3.34 $Y=1.32
+ $X2=3.255 $Y2=1.485
r93 10 12 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.34 $Y=1.32
+ $X2=3.34 $Y2=0.74
r94 7 37 57.1617 $w=2.98e-07 $l=3.1749e-07 $layer=POLY_cond $X=3.335 $Y=1.765
+ $X2=3.255 $Y2=1.485
r95 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.335 $Y=1.765
+ $X2=3.335 $Y2=2.4
r96 2 27 300 $w=1.7e-07 $l=6.15244e-07 $layer=licon1_PDIFF $count=2 $X=1 $Y=1.96
+ $X2=1.22 $Y2=2.475
r97 2 27 600 $w=1.7e-07 $l=2.94788e-07 $layer=licon1_PDIFF $count=1 $X=1 $Y=1.96
+ $X2=1.22 $Y2=2.135
r98 1 18 91 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_NDIFF $count=2 $X=1.585
+ $Y=0.37 $X2=1.78 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__O21BA_1%VPWR 1 2 3 10 12 18 22 24 26 31 38 39 45 48
r45 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r46 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r47 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r48 39 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r49 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r50 36 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.225 $Y=3.33
+ $X2=3.06 $Y2=3.33
r51 36 38 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=3.225 $Y=3.33
+ $X2=3.6 $Y2=3.33
r52 35 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r53 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r54 32 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.885 $Y=3.33
+ $X2=1.72 $Y2=3.33
r55 32 34 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=1.885 $Y=3.33
+ $X2=2.64 $Y2=3.33
r56 31 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.895 $Y=3.33
+ $X2=3.06 $Y2=3.33
r57 31 34 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.895 $Y=3.33
+ $X2=2.64 $Y2=3.33
r58 30 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r59 30 43 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.24 $Y2=3.33
r60 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r61 27 42 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.222 $Y2=3.33
r62 27 29 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=1.2 $Y2=3.33
r63 26 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.555 $Y=3.33
+ $X2=1.72 $Y2=3.33
r64 26 29 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=1.555 $Y=3.33
+ $X2=1.2 $Y2=3.33
r65 24 35 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.64 $Y2=3.33
r66 24 46 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r67 20 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.06 $Y=3.245
+ $X2=3.06 $Y2=3.33
r68 20 22 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=3.06 $Y=3.245
+ $X2=3.06 $Y2=2.78
r69 16 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.72 $Y=3.245
+ $X2=1.72 $Y2=3.33
r70 16 18 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=1.72 $Y=3.245
+ $X2=1.72 $Y2=2.78
r71 12 15 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.28 $Y=2.135
+ $X2=0.28 $Y2=2.815
r72 10 42 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.222 $Y2=3.33
r73 10 15 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.28 $Y2=2.815
r74 3 22 600 $w=1.7e-07 $l=1.05095e-06 $layer=licon1_PDIFF $count=1 $X=2.825
+ $Y=1.84 $X2=3.06 $Y2=2.78
r75 2 18 600 $w=1.7e-07 $l=8.91852e-07 $layer=licon1_PDIFF $count=1 $X=1.57
+ $Y=1.96 $X2=1.72 $Y2=2.78
r76 1 15 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.28 $Y2=2.815
r77 1 12 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.28 $Y2=2.135
.ends

.subckt PM_SKY130_FD_SC_LS__O21BA_1%X 1 2 9 13 14 15 16 23 32
c26 14 0 9.60317e-20 $X=3.515 $Y=1.95
r27 21 23 1.12043 $w=3.58e-07 $l=3.5e-08 $layer=LI1_cond $X=3.575 $Y=2 $X2=3.575
+ $Y2=2.035
r28 15 16 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=3.575 $Y=2.405
+ $X2=3.575 $Y2=2.775
r29 14 21 0.800308 $w=3.58e-07 $l=2.5e-08 $layer=LI1_cond $X=3.575 $Y=1.975
+ $X2=3.575 $Y2=2
r30 14 32 8.1909 $w=3.58e-07 $l=1.55e-07 $layer=LI1_cond $X=3.575 $Y=1.975
+ $X2=3.575 $Y2=1.82
r31 14 15 11.0442 $w=3.58e-07 $l=3.45e-07 $layer=LI1_cond $X=3.575 $Y=2.06
+ $X2=3.575 $Y2=2.405
r32 14 23 0.800308 $w=3.58e-07 $l=2.5e-08 $layer=LI1_cond $X=3.575 $Y=2.06
+ $X2=3.575 $Y2=2.035
r33 13 32 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.67 $Y=1.13 $X2=3.67
+ $Y2=1.82
r34 7 13 9.06106 $w=3.63e-07 $l=1.82e-07 $layer=LI1_cond $X=3.572 $Y=0.948
+ $X2=3.572 $Y2=1.13
r35 7 9 13.6714 $w=3.63e-07 $l=4.33e-07 $layer=LI1_cond $X=3.572 $Y=0.948
+ $X2=3.572 $Y2=0.515
r36 2 14 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=3.41
+ $Y=1.84 $X2=3.56 $Y2=1.985
r37 2 16 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=3.41
+ $Y=1.84 $X2=3.56 $Y2=2.815
r38 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.415
+ $Y=0.37 $X2=3.555 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__O21BA_1%A_27_74# 1 2 9 11 12 15
r27 13 15 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.28 $Y=0.79
+ $X2=1.28 $Y2=0.515
r28 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.115 $Y=0.875
+ $X2=1.28 $Y2=0.79
r29 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.115 $Y=0.875
+ $X2=0.445 $Y2=0.875
r30 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=0.79
+ $X2=0.445 $Y2=0.875
r31 7 9 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=0.28 $Y=0.79 $X2=0.28
+ $Y2=0.515
r32 2 15 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.14
+ $Y=0.37 $X2=1.28 $Y2=0.515
r33 1 9 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__O21BA_1%VGND 1 2 9 13 15 17 22 32 33 36 39
r40 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r41 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r42 33 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r43 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r44 30 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.22 $Y=0 $X2=3.055
+ $Y2=0
r45 30 32 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=3.22 $Y=0 $X2=3.6
+ $Y2=0
r46 29 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r47 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r48 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r49 25 28 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r50 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r51 23 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=0.78
+ $Y2=0
r52 23 25 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=1.2
+ $Y2=0
r53 22 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.89 $Y=0 $X2=3.055
+ $Y2=0
r54 22 28 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.89 $Y=0 $X2=2.64
+ $Y2=0
r55 20 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r56 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r57 17 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.78
+ $Y2=0
r58 17 19 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.24
+ $Y2=0
r59 15 29 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.64
+ $Y2=0
r60 15 26 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.2
+ $Y2=0
r61 11 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.055 $Y=0.085
+ $X2=3.055 $Y2=0
r62 11 13 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=3.055 $Y=0.085
+ $X2=3.055 $Y2=0.495
r63 7 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=0.085 $X2=0.78
+ $Y2=0
r64 7 9 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=0.78 $Y=0.085 $X2=0.78
+ $Y2=0.525
r65 2 13 91 $w=1.7e-07 $l=3.10805e-07 $layer=licon1_NDIFF $count=2 $X=2.845
+ $Y=0.56 $X2=3.125 $Y2=0.495
r66 1 9 182 $w=1.7e-07 $l=2.76857e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.78 $Y2=0.525
.ends

