* File: sky130_fd_sc_ls__inv_1.pxi.spice
* Created: Fri Aug 28 13:28:04 2020
* 
x_PM_SKY130_FD_SC_LS__INV_1%A N_A_c_25_n N_A_M1000_g N_A_M1001_g N_A_c_22_n
+ N_A_c_23_n A N_A_c_24_n PM_SKY130_FD_SC_LS__INV_1%A
x_PM_SKY130_FD_SC_LS__INV_1%VPWR N_VPWR_M1000_s N_VPWR_c_43_n VPWR N_VPWR_c_44_n
+ N_VPWR_c_45_n N_VPWR_c_42_n N_VPWR_c_47_n PM_SKY130_FD_SC_LS__INV_1%VPWR
x_PM_SKY130_FD_SC_LS__INV_1%Y N_Y_M1001_d N_Y_M1000_d Y Y Y Y Y Y Y
+ PM_SKY130_FD_SC_LS__INV_1%Y
x_PM_SKY130_FD_SC_LS__INV_1%VGND N_VGND_M1001_s N_VGND_c_68_n VGND N_VGND_c_69_n
+ N_VGND_c_70_n N_VGND_c_71_n N_VGND_c_72_n PM_SKY130_FD_SC_LS__INV_1%VGND
cc_1 VNB N_A_M1001_g 0.0324221f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=0.74
cc_2 VNB N_A_c_22_n 0.0799619f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=1.465
cc_3 VNB N_A_c_23_n 0.019289f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.532
cc_4 VNB N_A_c_24_n 0.0156043f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.465
cc_5 VNB N_VPWR_c_42_n 0.0641695f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB Y 0.054464f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_VGND_c_68_n 0.0443804f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=0.74
cc_8 VNB N_VGND_c_69_n 0.017577f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_9 VNB N_VGND_c_70_n 0.0194697f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_VGND_c_71_n 0.129238f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_VGND_c_72_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VPB N_A_c_25_n 0.0220613f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.765
cc_13 VPB N_A_c_23_n 0.00849648f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.532
cc_14 VPB N_A_c_24_n 0.0227034f $X=-0.19 $Y=1.66 $X2=0.65 $Y2=1.465
cc_15 VPB N_VPWR_c_43_n 0.0517561f $X=-0.19 $Y=1.66 $X2=0.935 $Y2=0.74
cc_16 VPB N_VPWR_c_44_n 0.017577f $X=-0.19 $Y=1.66 $X2=0.65 $Y2=1.465
cc_17 VPB N_VPWR_c_45_n 0.0194697f $X=-0.19 $Y=1.66 $X2=0.65 $Y2=1.54
cc_18 VPB N_VPWR_c_42_n 0.0647565f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_19 VPB N_VPWR_c_47_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_20 VPB Y 0.0535665f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_21 N_A_c_25_n N_VPWR_c_43_n 0.0249269f $X=0.925 $Y=1.765 $X2=0 $Y2=0
cc_22 N_A_c_22_n N_VPWR_c_43_n 0.00176665f $X=0.835 $Y=1.465 $X2=0 $Y2=0
cc_23 N_A_c_24_n N_VPWR_c_43_n 0.0283244f $X=0.65 $Y=1.465 $X2=0 $Y2=0
cc_24 N_A_c_25_n N_VPWR_c_45_n 0.00445602f $X=0.925 $Y=1.765 $X2=0 $Y2=0
cc_25 N_A_c_25_n N_VPWR_c_42_n 0.00865246f $X=0.925 $Y=1.765 $X2=0 $Y2=0
cc_26 N_A_c_25_n Y 0.0207035f $X=0.925 $Y=1.765 $X2=0 $Y2=0
cc_27 N_A_M1001_g Y 0.0212856f $X=0.935 $Y=0.74 $X2=0 $Y2=0
cc_28 N_A_c_23_n Y 0.0169685f $X=0.925 $Y=1.532 $X2=0 $Y2=0
cc_29 N_A_c_24_n Y 0.0388343f $X=0.65 $Y=1.465 $X2=0 $Y2=0
cc_30 N_A_M1001_g N_VGND_c_68_n 0.0198727f $X=0.935 $Y=0.74 $X2=0 $Y2=0
cc_31 N_A_c_22_n N_VGND_c_68_n 0.00764098f $X=0.835 $Y=1.465 $X2=0 $Y2=0
cc_32 N_A_c_24_n N_VGND_c_68_n 0.0283907f $X=0.65 $Y=1.465 $X2=0 $Y2=0
cc_33 N_A_M1001_g N_VGND_c_70_n 0.00434272f $X=0.935 $Y=0.74 $X2=0 $Y2=0
cc_34 N_A_M1001_g N_VGND_c_71_n 0.00828751f $X=0.935 $Y=0.74 $X2=0 $Y2=0
cc_35 N_VPWR_c_43_n Y 0.0394385f $X=0.65 $Y=2.115 $X2=0 $Y2=0
cc_36 N_VPWR_c_45_n Y 0.0145938f $X=1.2 $Y=3.33 $X2=0 $Y2=0
cc_37 N_VPWR_c_42_n Y 0.0120466f $X=1.2 $Y=3.33 $X2=0 $Y2=0
cc_38 Y N_VGND_c_68_n 0.0308485f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_39 Y N_VGND_c_70_n 0.0145639f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_40 Y N_VGND_c_71_n 0.0119984f $X=1.115 $Y=0.47 $X2=0 $Y2=0
