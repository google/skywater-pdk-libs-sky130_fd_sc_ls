* File: sky130_fd_sc_ls__sdfxtp_2.spice
* Created: Fri Aug 28 14:05:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__sdfxtp_2.pex.spice"
.subckt sky130_fd_sc_ls__sdfxtp_2  VNB VPB SCE D SCD CLK VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* CLK	CLK
* SCD	SCD
* D	D
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1030 N_VGND_M1030_d N_SCE_M1030_g N_A_27_74#_M1030_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0735 AS=0.1386 PD=0.77 PS=1.5 NRD=19.992 NRS=7.14 M=1 R=2.8 SA=75000.3
+ SB=75002.8 A=0.063 P=1.14 MULT=1
MM1014 A_223_74# N_A_27_74#_M1014_g N_VGND_M1030_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0735 PD=0.66 PS=0.77 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.8
+ SB=75002.3 A=0.063 P=1.14 MULT=1
MM1015 N_A_300_453#_M1015_d N_D_M1015_g A_223_74# VNB NSHORT L=0.15 W=0.42
+ AD=0.11655 AS=0.0504 PD=0.975 PS=0.66 NRD=38.568 NRS=18.564 M=1 R=2.8
+ SA=75001.1 SB=75001.9 A=0.063 P=1.14 MULT=1
MM1012 A_442_74# N_SCE_M1012_g N_A_300_453#_M1015_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.11655 PD=0.66 PS=0.975 NRD=18.564 NRS=39.996 M=1 R=2.8
+ SA=75001.8 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1000 N_VGND_M1000_d N_SCD_M1000_g A_442_74# VNB NSHORT L=0.15 W=0.42
+ AD=0.0968897 AS=0.0504 PD=0.84 PS=0.66 NRD=32.856 NRS=18.564 M=1 R=2.8
+ SA=75002.2 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1029 N_A_634_74#_M1029_d N_CLK_M1029_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.17071 PD=2.05 PS=1.48 NRD=0 NRS=4.044 M=1 R=4.93333 SA=75001.7
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1028 N_A_846_74#_M1028_d N_A_634_74#_M1028_g N_VGND_M1028_s VNB NSHORT L=0.15
+ W=0.74 AD=0.2109 AS=0.2627 PD=2.05 PS=2.19 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75000.3 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1033 N_A_1044_100#_M1033_d N_A_634_74#_M1033_g N_A_300_453#_M1033_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.15225 AS=0.1197 PD=1.145 PS=1.41 NRD=71.424 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75004.4 A=0.063 P=1.14 MULT=1
MM1002 A_1219_100# N_A_846_74#_M1002_g N_A_1044_100#_M1033_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0882 AS=0.15225 PD=0.84 PS=1.145 NRD=44.28 NRS=55.704 M=1 R=2.8
+ SA=75001.1 SB=75003.5 A=0.063 P=1.14 MULT=1
MM1008 N_VGND_M1008_d N_A_1287_320#_M1008_g A_1219_100# VNB NSHORT L=0.15 W=0.42
+ AD=0.195473 AS=0.0882 PD=1.25567 PS=0.84 NRD=117.252 NRS=44.28 M=1 R=2.8
+ SA=75001.7 SB=75002.9 A=0.063 P=1.14 MULT=1
MM1003 N_A_1287_320#_M1003_d N_A_1044_100#_M1003_g N_VGND_M1008_d VNB NSHORT
+ L=0.15 W=0.55 AD=0.18975 AS=0.255977 PD=1.24 PS=1.64433 NRD=0 NRS=90.54 M=1
+ R=3.66667 SA=75002.1 SB=75002.1 A=0.0825 P=1.4 MULT=1
MM1010 N_A_1592_424#_M1010_d N_A_846_74#_M1010_g N_A_1287_320#_M1003_d VNB
+ NSHORT L=0.15 W=0.55 AD=0.10674 AS=0.18975 PD=1.03196 PS=1.24 NRD=0 NRS=89.448
+ M=1 R=3.66667 SA=75003 SB=75001.3 A=0.0825 P=1.4 MULT=1
MM1020 A_1787_74# N_A_634_74#_M1020_g N_A_1592_424#_M1010_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.0815103 PD=0.66 PS=0.788041 NRD=18.564 NRS=22.848 M=1
+ R=2.8 SA=75003.3 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1021 N_VGND_M1021_d N_A_1829_398#_M1021_g A_1787_74# VNB NSHORT L=0.15 W=0.42
+ AD=0.0821897 AS=0.0504 PD=0.78931 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8
+ SA=75003.7 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1016 N_A_1829_398#_M1016_d N_A_1592_424#_M1016_g N_VGND_M1021_d VNB NSHORT
+ L=0.15 W=0.74 AD=0.2109 AS=0.14481 PD=2.05 PS=1.39069 NRD=0 NRS=11.34 M=1
+ R=4.93333 SA=75002.5 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1001 N_VGND_M1001_d N_A_1829_398#_M1001_g N_Q_M1001_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2627 AS=0.12025 PD=2.19 PS=1.065 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.3
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1023 N_VGND_M1023_d N_A_1829_398#_M1023_g N_Q_M1001_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2294 AS=0.12025 PD=2.1 PS=1.065 NRD=4.044 NRS=7.296 M=1 R=4.93333
+ SA=75000.8 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1024 N_VPWR_M1024_d N_SCE_M1024_g N_A_27_74#_M1024_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.112 AS=0.1888 PD=0.99 PS=1.87 NRD=18.4589 NRS=3.0732 M=1 R=4.26667
+ SA=75000.2 SB=75003 A=0.096 P=1.58 MULT=1
MM1022 A_216_453# N_SCE_M1022_g N_VPWR_M1024_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0864 AS=0.112 PD=0.91 PS=0.99 NRD=24.625 NRS=3.0732 M=1 R=4.26667
+ SA=75000.7 SB=75002.5 A=0.096 P=1.58 MULT=1
MM1013 N_A_300_453#_M1013_d N_D_M1013_g A_216_453# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1744 AS=0.0864 PD=1.185 PS=0.91 NRD=40.0107 NRS=24.625 M=1 R=4.26667
+ SA=75001.1 SB=75002.1 A=0.096 P=1.58 MULT=1
MM1006 A_439_453# N_A_27_74#_M1006_g N_A_300_453#_M1013_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0864 AS=0.1744 PD=0.91 PS=1.185 NRD=24.625 NRS=41.5473 M=1
+ R=4.26667 SA=75001.8 SB=75001.4 A=0.096 P=1.58 MULT=1
MM1017 N_VPWR_M1017_d N_SCD_M1017_g A_439_453# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.209136 AS=0.0864 PD=1.34545 PS=0.91 NRD=49.25 NRS=24.625 M=1 R=4.26667
+ SA=75002.3 SB=75001 A=0.096 P=1.58 MULT=1
MM1004 N_A_634_74#_M1004_d N_CLK_M1004_g N_VPWR_M1017_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.3304 AS=0.365989 PD=2.83 PS=2.35455 NRD=1.7533 NRS=28.1316 M=1
+ R=7.46667 SA=75001.8 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1027 N_A_846_74#_M1027_d N_A_634_74#_M1027_g N_VPWR_M1027_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.3304 AS=0.6426 PD=2.83 PS=3.56 NRD=1.7533 NRS=29.8849 M=1
+ R=7.46667 SA=75000.4 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1026 N_A_1044_100#_M1026_d N_A_846_74#_M1026_g N_A_300_453#_M1026_s VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.063 AS=0.1239 PD=0.72 PS=1.43 NRD=4.6886 NRS=4.6886
+ M=1 R=2.8 SA=75000.2 SB=75004.4 A=0.063 P=1.14 MULT=1
MM1031 A_1210_508# N_A_634_74#_M1031_g N_A_1044_100#_M1026_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.084 AS=0.063 PD=0.82 PS=0.72 NRD=68.0044 NRS=4.6886 M=1 R=2.8
+ SA=75000.7 SB=75004 A=0.063 P=1.14 MULT=1
MM1005 N_VPWR_M1005_d N_A_1287_320#_M1005_g A_1210_508# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.084 PD=0.913333 PS=0.82 NRD=4.6886 NRS=68.0044 M=1 R=2.8
+ SA=75001.2 SB=75003.4 A=0.063 P=1.14 MULT=1
MM1007 N_A_1287_320#_M1007_d N_A_1044_100#_M1007_g N_VPWR_M1005_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.2226 AS=0.2226 PD=1.37 PS=1.82667 NRD=2.3443 NRS=56.2829
+ M=1 R=5.6 SA=75001 SB=75002 A=0.126 P=1.98 MULT=1
MM1025 N_A_1592_424#_M1025_d N_A_634_74#_M1025_g N_A_1287_320#_M1007_d VPB
+ PHIGHVT L=0.15 W=0.84 AD=0.1962 AS=0.2226 PD=1.66667 PS=1.37 NRD=2.3443
+ NRS=56.2829 M=1 R=5.6 SA=75001.7 SB=75001.3 A=0.126 P=1.98 MULT=1
MM1011 A_1704_496# N_A_846_74#_M1011_g N_A_1592_424#_M1025_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1344 AS=0.0981 PD=1.06 PS=0.833333 NRD=124.287 NRS=56.2829 M=1
+ R=2.8 SA=75002.9 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1032 N_VPWR_M1032_d N_A_1829_398#_M1032_g A_1704_496# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.126207 AS=0.1344 PD=0.976056 PS=1.06 NRD=4.6886 NRS=124.287 M=1
+ R=2.8 SA=75003.7 SB=75001 A=0.063 P=1.14 MULT=1
MM1018 N_A_1829_398#_M1018_d N_A_1592_424#_M1018_g N_VPWR_M1032_d VPB PHIGHVT
+ L=0.15 W=1 AD=0.295 AS=0.300493 PD=2.59 PS=2.32394 NRD=1.9503 NRS=1.9503 M=1
+ R=6.66667 SA=75002 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1009 N_Q_M1009_d N_A_1829_398#_M1009_g N_VPWR_M1009_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1019 N_Q_M1009_d N_A_1829_398#_M1019_g N_VPWR_M1019_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75000.2 A=0.168 P=2.54 MULT=1
DX34_noxref VNB VPB NWDIODE A=23.0268 P=28.48
c_127 VNB 0 1.87953e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_ls__sdfxtp_2.pxi.spice"
*
.ends
*
*
