* File: sky130_fd_sc_ls__sdlclkp_1.spice
* Created: Fri Aug 28 14:06:13 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__sdlclkp_1.pex.spice"
.subckt sky130_fd_sc_ls__sdlclkp_1  VNB VPB SCE GATE CLK VPWR GCLK VGND
* 
* VGND	VGND
* GCLK	GCLK
* VPWR	VPWR
* CLK	CLK
* GATE	GATE
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1009 N_A_114_112#_M1009_d N_SCE_M1009_g N_VGND_M1009_s VNB NSHORT L=0.15
+ W=0.55 AD=0.077 AS=0.15675 PD=0.83 PS=1.67 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75001.2 A=0.0825 P=1.4 MULT=1
MM1008 N_VGND_M1008_d N_GATE_M1008_g N_A_114_112#_M1009_d VNB NSHORT L=0.15
+ W=0.55 AD=0.161184 AS=0.077 PD=1.20233 PS=0.83 NRD=51.936 NRS=0 M=1 R=3.66667
+ SA=75000.6 SB=75000.8 A=0.0825 P=1.4 MULT=1
MM1000 N_A_318_74#_M1000_d N_A_288_48#_M1000_g N_VGND_M1008_d VNB NSHORT L=0.15
+ W=0.74 AD=0.2109 AS=0.216866 PD=2.05 PS=1.61767 NRD=0 NRS=38.604 M=1 R=4.93333
+ SA=75001 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1015 N_A_566_74#_M1015_d N_A_288_48#_M1015_g N_A_114_112#_M1015_s VNB NSHORT
+ L=0.15 W=0.55 AD=0.10467 AS=0.29425 PD=1.02629 PS=2.17 NRD=0 NRS=54.54 M=1
+ R=3.66667 SA=75000.5 SB=75001.4 A=0.0825 P=1.4 MULT=1
MM1012 A_667_80# N_A_318_74#_M1012_g N_A_566_74#_M1015_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.0799299 PD=0.63 PS=0.783711 NRD=14.28 NRS=22.848 M=1
+ R=2.8 SA=75001 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1013 N_VGND_M1013_d N_A_709_54#_M1013_g A_667_80# VNB NSHORT L=0.15 W=0.42
+ AD=0.109562 AS=0.0441 PD=0.919655 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.3
+ SB=75000.9 A=0.063 P=1.14 MULT=1
MM1007 N_A_709_54#_M1007_d N_A_566_74#_M1007_g N_VGND_M1013_d VNB NSHORT L=0.15
+ W=0.74 AD=0.2072 AS=0.193038 PD=2.04 PS=1.62034 NRD=0 NRS=40.536 M=1 R=4.93333
+ SA=75001.2 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1002 N_VGND_M1002_d N_CLK_M1002_g N_A_288_48#_M1002_s VNB NSHORT L=0.15 W=0.74
+ AD=0.124942 AS=0.2072 PD=1.14217 PS=2.04 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.9 A=0.111 P=1.78 MULT=1
MM1003 A_1166_94# N_CLK_M1003_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.64
+ AD=0.0672 AS=0.108058 PD=0.85 PS=0.987826 NRD=9.372 NRS=8.436 M=1 R=4.26667
+ SA=75000.7 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1005 N_A_1238_94#_M1005_d N_A_709_54#_M1005_g A_1166_94# VNB NSHORT L=0.15
+ W=0.64 AD=0.1824 AS=0.0672 PD=1.85 PS=0.85 NRD=0 NRS=9.372 M=1 R=4.26667
+ SA=75001 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1018 N_GCLK_M1018_d N_A_1238_94#_M1018_g N_VGND_M1018_s VNB NSHORT L=0.15
+ W=0.74 AD=0.2072 AS=0.2664 PD=2.04 PS=2.2 NRD=0 NRS=12.156 M=1 R=4.93333
+ SA=75000.3 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1014 A_116_424# N_SCE_M1014_g N_VPWR_M1014_s VPB PHIGHVT L=0.15 W=0.84
+ AD=0.1008 AS=0.2478 PD=1.08 PS=2.27 NRD=15.2281 NRS=2.3443 M=1 R=5.6
+ SA=75000.2 SB=75000.6 A=0.126 P=1.98 MULT=1
MM1019 N_A_114_112#_M1019_d N_GATE_M1019_g A_116_424# VPB PHIGHVT L=0.15 W=0.84
+ AD=0.2478 AS=0.1008 PD=2.27 PS=1.08 NRD=2.3443 NRS=15.2281 M=1 R=5.6
+ SA=75000.6 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1004 N_A_318_74#_M1004_d N_A_288_48#_M1004_g N_VPWR_M1004_s VPB PHIGHVT L=0.15
+ W=0.84 AD=0.2478 AS=0.4033 PD=2.27 PS=3.02 NRD=2.3443 NRS=99.682 M=1 R=5.6
+ SA=75000.3 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1006 N_A_566_74#_M1006_d N_A_318_74#_M1006_g N_A_114_112#_M1006_s VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.207317 AS=0.2478 PD=1.82667 PS=2.27 NRD=2.3443 NRS=2.3443
+ M=1 R=5.6 SA=75000.2 SB=75000.7 A=0.126 P=1.98 MULT=1
MM1020 A_722_492# N_A_288_48#_M1020_g N_A_566_74#_M1006_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0504 AS=0.103658 PD=0.66 PS=0.913333 NRD=30.4759 NRS=44.5417 M=1
+ R=2.8 SA=75000.6 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1001 N_VPWR_M1001_d N_A_709_54#_M1001_g A_722_492# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0912545 AS=0.0504 PD=0.804545 PS=0.66 NRD=4.6886 NRS=30.4759 M=1 R=2.8
+ SA=75000.9 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1016 N_A_709_54#_M1016_d N_A_566_74#_M1016_g N_VPWR_M1001_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.3304 AS=0.243345 PD=2.83 PS=2.14545 NRD=1.7533 NRS=11.426 M=1
+ R=7.46667 SA=75000.7 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1021 N_VPWR_M1021_d N_CLK_M1021_g N_A_288_48#_M1021_s VPB PHIGHVT L=0.15
+ W=0.84 AD=0.281825 AS=0.2478 PD=1.675 PS=2.27 NRD=65.7783 NRS=2.3443 M=1 R=5.6
+ SA=75000.2 SB=75002 A=0.126 P=1.98 MULT=1
MM1010 N_A_1238_94#_M1010_d N_CLK_M1010_g N_VPWR_M1021_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.126 AS=0.281825 PD=1.14 PS=1.675 NRD=2.3443 NRS=65.7783 M=1 R=5.6
+ SA=75000.9 SB=75001.3 A=0.126 P=1.98 MULT=1
MM1017 N_VPWR_M1017_d N_A_709_54#_M1017_g N_A_1238_94#_M1010_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.1596 AS=0.126 PD=1.26429 PS=1.14 NRD=14.0658 NRS=2.3443 M=1
+ R=5.6 SA=75001.4 SB=75000.8 A=0.126 P=1.98 MULT=1
MM1011 N_GCLK_M1011_d N_A_1238_94#_M1011_g N_VPWR_M1017_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.4256 AS=0.2128 PD=3 PS=1.68571 NRD=16.7056 NRS=2.6201 M=1
+ R=7.46667 SA=75001.4 SB=75000.3 A=0.168 P=2.54 MULT=1
DX22_noxref VNB VPB NWDIODE A=15.0772 P=20
*
.include "sky130_fd_sc_ls__sdlclkp_1.pxi.spice"
*
.ends
*
*
