* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__dlrtp_4 D GATE RESET_B VGND VNB VPB VPWR Q
X0 Q a_797_48# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X1 a_797_48# a_640_74# a_938_74# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X2 VPWR a_640_74# a_797_48# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X3 a_562_392# a_240_394# a_640_74# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 VGND a_27_126# a_559_74# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X5 a_364_120# a_240_394# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X6 a_27_126# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X7 a_747_508# a_797_48# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 VPWR a_797_48# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X9 a_797_48# a_640_74# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X10 VGND a_797_48# Q VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X11 a_938_74# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X12 VGND RESET_B a_938_74# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X13 VPWR RESET_B a_797_48# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X14 a_27_126# D VGND VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X15 Q a_797_48# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X16 VPWR a_27_126# a_562_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X17 VGND GATE a_240_394# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X18 VPWR a_797_48# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X19 VGND a_797_48# Q VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X20 a_364_120# a_240_394# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X21 Q a_797_48# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X22 a_559_74# a_364_120# a_640_74# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X23 Q a_797_48# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X24 a_640_74# a_240_394# a_755_74# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X25 a_797_48# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X26 a_938_74# a_640_74# a_797_48# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X27 a_755_74# a_797_48# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X28 VPWR GATE a_240_394# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X29 a_640_74# a_364_120# a_747_508# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
.ends
