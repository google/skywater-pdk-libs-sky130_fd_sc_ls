* File: sky130_fd_sc_ls__mux2i_2.pex.spice
* Created: Wed Sep  2 11:10:39 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__MUX2I_2%A0 1 3 4 6 7 9 10 12 13 14 22
c52 7 0 3.78814e-19 $X=1.005 $Y=1.765
c53 4 0 1.51809e-19 $X=0.515 $Y=1.765
r54 22 23 1.62472 $w=4.45e-07 $l=1.5e-08 $layer=POLY_cond $X=1.005 $Y=1.492
+ $X2=1.02 $Y2=1.492
r55 20 22 8.1236 $w=4.45e-07 $l=7.5e-08 $layer=POLY_cond $X=0.93 $Y=1.492
+ $X2=1.005 $Y2=1.492
r56 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.93
+ $Y=1.385 $X2=0.93 $Y2=1.385
r57 18 20 44.9506 $w=4.45e-07 $l=4.15e-07 $layer=POLY_cond $X=0.515 $Y=1.492
+ $X2=0.93 $Y2=1.492
r58 17 18 1.62472 $w=4.45e-07 $l=1.5e-08 $layer=POLY_cond $X=0.5 $Y=1.492
+ $X2=0.515 $Y2=1.492
r59 14 21 8.40972 $w=3.68e-07 $l=2.7e-07 $layer=LI1_cond $X=1.2 $Y=1.365
+ $X2=0.93 $Y2=1.365
r60 13 21 6.54089 $w=3.68e-07 $l=2.1e-07 $layer=LI1_cond $X=0.72 $Y=1.365
+ $X2=0.93 $Y2=1.365
r61 10 23 28.4889 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=1.02 $Y=1.22
+ $X2=1.02 $Y2=1.492
r62 10 12 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.02 $Y=1.22 $X2=1.02
+ $Y2=0.74
r63 7 22 28.4889 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=1.005 $Y=1.765
+ $X2=1.005 $Y2=1.492
r64 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.005 $Y=1.765
+ $X2=1.005 $Y2=2.4
r65 4 18 28.4889 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=0.515 $Y=1.765
+ $X2=0.515 $Y2=1.492
r66 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.515 $Y=1.765
+ $X2=0.515 $Y2=2.4
r67 1 17 28.4889 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=0.5 $Y=1.22 $X2=0.5
+ $Y2=1.492
r68 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.5 $Y=1.22 $X2=0.5
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__MUX2I_2%A1 3 5 7 8 10 12 15 17 18 19 20 26 29
c63 20 0 2.4396e-19 $X=3.12 $Y=1.665
r64 29 30 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.38
+ $Y=1.515 $X2=2.38 $Y2=1.515
r65 26 27 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.7
+ $Y=1.515 $X2=1.7 $Y2=1.515
r66 19 20 16.034 $w=3.43e-07 $l=4.8e-07 $layer=LI1_cond $X=2.64 $Y=1.602
+ $X2=3.12 $Y2=1.602
r67 19 30 8.68508 $w=3.43e-07 $l=2.6e-07 $layer=LI1_cond $X=2.64 $Y=1.602
+ $X2=2.38 $Y2=1.602
r68 18 30 7.34891 $w=3.43e-07 $l=2.2e-07 $layer=LI1_cond $X=2.16 $Y=1.602
+ $X2=2.38 $Y2=1.602
r69 18 27 15.3659 $w=3.43e-07 $l=4.6e-07 $layer=LI1_cond $X=2.16 $Y=1.602
+ $X2=1.7 $Y2=1.602
r70 17 27 0.668083 $w=3.43e-07 $l=2e-08 $layer=LI1_cond $X=1.68 $Y=1.602 $X2=1.7
+ $Y2=1.602
r71 13 29 37.0704 $w=1.5e-07 $l=2.14369e-07 $layer=POLY_cond $X=2.47 $Y=1.35
+ $X2=2.455 $Y2=1.557
r72 13 15 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.47 $Y=1.35
+ $X2=2.47 $Y2=0.74
r73 10 29 37.0704 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.455 $Y=1.765
+ $X2=2.455 $Y2=1.557
r74 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.455 $Y=1.765
+ $X2=2.455 $Y2=2.4
r75 9 26 5.03009 $w=3.3e-07 $l=1.08995e-07 $layer=POLY_cond $X=1.715 $Y=1.515
+ $X2=1.625 $Y2=1.557
r76 8 29 5.03009 $w=3.3e-07 $l=1.08995e-07 $layer=POLY_cond $X=2.365 $Y=1.515
+ $X2=2.455 $Y2=1.557
r77 8 9 113.66 $w=3.3e-07 $l=6.5e-07 $layer=POLY_cond $X=2.365 $Y=1.515
+ $X2=1.715 $Y2=1.515
r78 5 26 37.0704 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.625 $Y=1.765
+ $X2=1.625 $Y2=1.557
r79 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.625 $Y=1.765
+ $X2=1.625 $Y2=2.4
r80 1 26 37.0704 $w=1.5e-07 $l=2.14369e-07 $layer=POLY_cond $X=1.61 $Y=1.35
+ $X2=1.625 $Y2=1.557
r81 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.61 $Y=1.35 $X2=1.61
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__MUX2I_2%S 1 3 4 6 7 9 10 12 13 15 16 18 19 23 26 27
+ 28 37 48 50
c94 4 0 5.75093e-20 $X=3.615 $Y=1.765
r95 37 38 1.928 $w=3.75e-07 $l=1.5e-08 $layer=POLY_cond $X=4.065 $Y=1.557
+ $X2=4.08 $Y2=1.557
r96 35 37 4.49867 $w=3.75e-07 $l=3.5e-08 $layer=POLY_cond $X=4.03 $Y=1.557
+ $X2=4.065 $Y2=1.557
r97 35 36 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.03
+ $Y=1.515 $X2=4.03 $Y2=1.515
r98 33 35 53.3413 $w=3.75e-07 $l=4.15e-07 $layer=POLY_cond $X=3.615 $Y=1.557
+ $X2=4.03 $Y2=1.557
r99 32 33 1.928 $w=3.75e-07 $l=1.5e-08 $layer=POLY_cond $X=3.6 $Y=1.557
+ $X2=3.615 $Y2=1.557
r100 28 50 8.99479 $w=5.78e-07 $l=1.15e-07 $layer=LI1_cond $X=4.56 $Y=1.72
+ $X2=4.675 $Y2=1.72
r101 28 48 5.37376 $w=5.78e-07 $l=2.1e-07 $layer=LI1_cond $X=4.56 $Y=1.72
+ $X2=4.35 $Y2=1.72
r102 27 48 7.58926 $w=4.08e-07 $l=2.7e-07 $layer=LI1_cond $X=4.08 $Y=1.635
+ $X2=4.35 $Y2=1.635
r103 27 36 1.40542 $w=4.08e-07 $l=5e-08 $layer=LI1_cond $X=4.08 $Y=1.635
+ $X2=4.03 $Y2=1.635
r104 26 36 12.0866 $w=4.08e-07 $l=4.3e-07 $layer=LI1_cond $X=3.6 $Y=1.635
+ $X2=4.03 $Y2=1.635
r105 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.645
+ $Y=1.515 $X2=5.645 $Y2=1.515
r106 21 23 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=5.645 $Y=1.84
+ $X2=5.645 $Y2=1.515
r107 19 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.48 $Y=1.925
+ $X2=5.645 $Y2=1.84
r108 19 50 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=5.48 $Y=1.925
+ $X2=4.675 $Y2=1.925
r109 16 24 38.532 $w=3.11e-07 $l=2.06325e-07 $layer=POLY_cond $X=5.745 $Y=1.35
+ $X2=5.652 $Y2=1.515
r110 16 18 141.387 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=5.745 $Y=1.35
+ $X2=5.745 $Y2=0.91
r111 13 24 51.7056 $w=3.11e-07 $l=2.88531e-07 $layer=POLY_cond $X=5.735 $Y=1.765
+ $X2=5.652 $Y2=1.515
r112 13 15 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.735 $Y=1.765
+ $X2=5.735 $Y2=2.34
r113 10 38 24.2915 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.08 $Y=1.35
+ $X2=4.08 $Y2=1.557
r114 10 12 157.453 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=4.08 $Y=1.35
+ $X2=4.08 $Y2=0.86
r115 7 37 24.2915 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=4.065 $Y=1.765
+ $X2=4.065 $Y2=1.557
r116 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.065 $Y=1.765
+ $X2=4.065 $Y2=2.4
r117 4 33 24.2915 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.615 $Y=1.765
+ $X2=3.615 $Y2=1.557
r118 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.615 $Y=1.765
+ $X2=3.615 $Y2=2.4
r119 1 32 24.2915 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.6 $Y=1.35 $X2=3.6
+ $Y2=1.557
r120 1 3 157.453 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=3.6 $Y=1.35 $X2=3.6
+ $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_LS__MUX2I_2%A_922_72# 1 2 7 9 10 12 13 15 16 18 21 24 25
+ 28 34 36 37 41
c77 13 0 6.86239e-20 $X=5.15 $Y=1.765
r78 41 42 1.88281 $w=3.84e-07 $l=1.5e-08 $layer=POLY_cond $X=5.15 $Y=1.552
+ $X2=5.165 $Y2=1.552
r79 38 39 1.88281 $w=3.84e-07 $l=1.5e-08 $layer=POLY_cond $X=4.685 $Y=1.552
+ $X2=4.7 $Y2=1.552
r80 36 37 5.902 $w=3.53e-07 $l=8.5e-08 $layer=LI1_cond $X=5.972 $Y=2.265
+ $X2=5.972 $Y2=2.18
r81 32 34 3.55013 $w=2.62e-07 $l=1.28662e-07 $layer=LI1_cond $X=6.065 $Y=1.18
+ $X2=5.972 $Y2=1.095
r82 32 37 65.2406 $w=1.68e-07 $l=1e-06 $layer=LI1_cond $X=6.065 $Y=1.18
+ $X2=6.065 $Y2=2.18
r83 26 34 3.55013 $w=2.62e-07 $l=8.5e-08 $layer=LI1_cond $X=5.972 $Y=1.01
+ $X2=5.972 $Y2=1.095
r84 26 28 8.92738 $w=3.53e-07 $l=2.75e-07 $layer=LI1_cond $X=5.972 $Y=1.01
+ $X2=5.972 $Y2=0.735
r85 24 34 2.9446 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=5.795 $Y=1.095
+ $X2=5.972 $Y2=1.095
r86 24 25 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=5.795 $Y=1.095
+ $X2=5.24 $Y2=1.095
r87 22 41 9.41406 $w=3.84e-07 $l=7.5e-08 $layer=POLY_cond $X=5.075 $Y=1.552
+ $X2=5.15 $Y2=1.552
r88 22 39 47.0703 $w=3.84e-07 $l=3.75e-07 $layer=POLY_cond $X=5.075 $Y=1.552
+ $X2=4.7 $Y2=1.552
r89 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.075
+ $Y=1.505 $X2=5.075 $Y2=1.505
r90 19 25 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.075 $Y=1.18
+ $X2=5.24 $Y2=1.095
r91 19 21 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=5.075 $Y=1.18
+ $X2=5.075 $Y2=1.505
r92 16 42 24.8669 $w=1.5e-07 $l=2.12e-07 $layer=POLY_cond $X=5.165 $Y=1.34
+ $X2=5.165 $Y2=1.552
r93 16 18 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.165 $Y=1.34
+ $X2=5.165 $Y2=0.86
r94 13 41 24.8669 $w=1.5e-07 $l=2.13e-07 $layer=POLY_cond $X=5.15 $Y=1.765
+ $X2=5.15 $Y2=1.552
r95 13 15 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.15 $Y=1.765
+ $X2=5.15 $Y2=2.4
r96 10 39 24.8669 $w=1.5e-07 $l=2.13e-07 $layer=POLY_cond $X=4.7 $Y=1.765
+ $X2=4.7 $Y2=1.552
r97 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.7 $Y=1.765
+ $X2=4.7 $Y2=2.4
r98 7 38 24.8669 $w=1.5e-07 $l=2.12e-07 $layer=POLY_cond $X=4.685 $Y=1.34
+ $X2=4.685 $Y2=1.552
r99 7 9 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.685 $Y=1.34 $X2=4.685
+ $Y2=0.86
r100 2 36 300 $w=1.7e-07 $l=4.94343e-07 $layer=licon1_PDIFF $count=2 $X=5.81
+ $Y=1.84 $X2=5.96 $Y2=2.265
r101 1 28 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.82
+ $Y=0.59 $X2=5.96 $Y2=0.735
.ends

.subckt PM_SKY130_FD_SC_LS__MUX2I_2%Y 1 2 3 4 5 6 22 29 31 32 35 36 41 42 43 57
+ 58 62
c68 58 0 1.51809e-19 $X=0.265 $Y=1.82
c69 41 0 1.92364e-19 $X=0.155 $Y=1.95
c70 31 0 4.77058e-20 $X=2.58 $Y=0.34
r71 57 59 1.44055 $w=3.58e-07 $l=4.5e-08 $layer=LI1_cond $X=0.265 $Y=1.985
+ $X2=0.265 $Y2=2.03
r72 57 58 8.51103 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=0.265 $Y=1.985
+ $X2=0.265 $Y2=1.82
r73 48 62 2.56098 $w=3.58e-07 $l=8e-08 $layer=LI1_cond $X=0.265 $Y=2.115
+ $X2=0.265 $Y2=2.035
r74 42 43 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=0.265 $Y=2.405
+ $X2=0.265 $Y2=2.775
r75 41 62 0.0960369 $w=3.58e-07 $l=3e-09 $layer=LI1_cond $X=0.265 $Y=2.032
+ $X2=0.265 $Y2=2.035
r76 41 59 0.0640246 $w=3.58e-07 $l=2e-09 $layer=LI1_cond $X=0.265 $Y=2.032
+ $X2=0.265 $Y2=2.03
r77 41 42 9.21954 $w=3.58e-07 $l=2.88e-07 $layer=LI1_cond $X=0.265 $Y=2.117
+ $X2=0.265 $Y2=2.405
r78 41 48 0.0640246 $w=3.58e-07 $l=2e-09 $layer=LI1_cond $X=0.265 $Y=2.117
+ $X2=0.265 $Y2=2.115
r79 36 39 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=2.745 $Y=0.34
+ $X2=2.745 $Y2=0.495
r80 35 58 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=0.17 $Y=1.01
+ $X2=0.17 $Y2=1.82
r81 32 34 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=0.45 $Y=0.34
+ $X2=1.315 $Y2=0.34
r82 31 36 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.58 $Y=0.34
+ $X2=2.745 $Y2=0.34
r83 31 34 82.5294 $w=1.68e-07 $l=1.265e-06 $layer=LI1_cond $X=2.58 $Y=0.34
+ $X2=1.315 $Y2=0.34
r84 27 29 89.0535 $w=1.68e-07 $l=1.365e-06 $layer=LI1_cond $X=1.315 $Y=2.03
+ $X2=2.68 $Y2=2.03
r85 25 59 5.14255 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=0.445 $Y=2.03
+ $X2=0.265 $Y2=2.03
r86 25 27 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=0.445 $Y=2.03
+ $X2=1.315 $Y2=2.03
r87 20 35 9.06106 $w=3.63e-07 $l=1.82e-07 $layer=LI1_cond $X=0.267 $Y=0.828
+ $X2=0.267 $Y2=1.01
r88 20 22 9.88259 $w=3.63e-07 $l=3.13e-07 $layer=LI1_cond $X=0.267 $Y=0.828
+ $X2=0.267 $Y2=0.515
r89 19 32 8.06639 $w=1.7e-07 $l=2.21459e-07 $layer=LI1_cond $X=0.267 $Y=0.425
+ $X2=0.45 $Y2=0.34
r90 19 22 2.84164 $w=3.63e-07 $l=9e-08 $layer=LI1_cond $X=0.267 $Y=0.425
+ $X2=0.267 $Y2=0.515
r91 6 29 600 $w=1.7e-07 $l=2.54165e-07 $layer=licon1_PDIFF $count=1 $X=2.53
+ $Y=1.84 $X2=2.68 $Y2=2.03
r92 5 27 600 $w=1.7e-07 $l=3.1603e-07 $layer=licon1_PDIFF $count=1 $X=1.08
+ $Y=1.84 $X2=1.315 $Y2=2.03
r93 4 57 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
r94 4 43 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r95 3 39 182 $w=1.7e-07 $l=2.54951e-07 $layer=licon1_NDIFF $count=1 $X=2.545
+ $Y=0.37 $X2=2.745 $Y2=0.495
r96 2 34 182 $w=1.7e-07 $l=2.34521e-07 $layer=licon1_NDIFF $count=1 $X=1.095
+ $Y=0.37 $X2=1.315 $Y2=0.34
r97 1 22 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.14
+ $Y=0.37 $X2=0.285 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__MUX2I_2%A_118_368# 1 2 13 16 17 18
c36 13 0 3.09973e-20 $X=3.84 $Y=2.175
r37 17 18 8.63679 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=3.015 $Y=2.232
+ $X2=3.185 $Y2=2.232
r38 13 18 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=3.84 $Y=2.175
+ $X2=3.185 $Y2=2.175
r39 10 16 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=2.37
+ $X2=0.78 $Y2=2.37
r40 10 17 135.048 $w=1.68e-07 $l=2.07e-06 $layer=LI1_cond $X=0.945 $Y=2.37
+ $X2=3.015 $Y2=2.37
r41 2 13 600 $w=1.7e-07 $l=4.03082e-07 $layer=licon1_PDIFF $count=1 $X=3.69
+ $Y=1.84 $X2=3.84 $Y2=2.175
r42 1 16 300 $w=1.7e-07 $l=6.17738e-07 $layer=licon1_PDIFF $count=2 $X=0.59
+ $Y=1.84 $X2=0.78 $Y2=2.37
.ends

.subckt PM_SKY130_FD_SC_LS__MUX2I_2%A_340_368# 1 2 9 11 14 15 16 21
c44 11 0 6.86239e-20 $X=4.76 $Y=2.595
r45 21 23 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=4.925 $Y=2.265
+ $X2=4.925 $Y2=2.595
r46 16 18 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=3.44 $Y=2.595
+ $X2=3.44 $Y2=2.71
r47 14 15 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.23 $Y=2.79
+ $X2=2.395 $Y2=2.79
r48 12 16 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.525 $Y=2.595
+ $X2=3.44 $Y2=2.595
r49 11 23 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.76 $Y=2.595
+ $X2=4.925 $Y2=2.595
r50 11 12 80.5722 $w=1.68e-07 $l=1.235e-06 $layer=LI1_cond $X=4.76 $Y=2.595
+ $X2=3.525 $Y2=2.595
r51 9 18 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.355 $Y=2.71
+ $X2=3.44 $Y2=2.71
r52 9 15 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.355 $Y=2.71
+ $X2=2.395 $Y2=2.71
r53 2 21 300 $w=1.7e-07 $l=4.94343e-07 $layer=licon1_PDIFF $count=2 $X=4.775
+ $Y=1.84 $X2=4.925 $Y2=2.265
r54 1 14 300 $w=1.7e-07 $l=1.18575e-06 $layer=licon1_PDIFF $count=2 $X=1.7
+ $Y=1.84 $X2=2.23 $Y2=2.79
.ends

.subckt PM_SKY130_FD_SC_LS__MUX2I_2%VPWR 1 2 3 12 16 21 22 24 25 26 28 41 42 45
c66 45 0 3.09973e-20 $X=3.27 $Y=3.05
r67 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r68 39 42 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33 $X2=6
+ $Y2=3.33
r69 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r70 36 39 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r71 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r72 33 35 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=3.47 $Y=3.33
+ $X2=4.08 $Y2=3.33
r73 30 31 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r74 28 33 5.70203 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=3.272 $Y=3.33
+ $X2=3.47 $Y2=3.33
r75 28 45 8.16922 $w=3.93e-07 $l=2.8e-07 $layer=LI1_cond $X=3.272 $Y=3.33
+ $X2=3.272 $Y2=3.05
r76 28 30 184.957 $w=1.68e-07 $l=2.835e-06 $layer=LI1_cond $X=3.075 $Y=3.33
+ $X2=0.24 $Y2=3.33
r77 26 36 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r78 26 31 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=0.24 $Y2=3.33
r79 26 28 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r80 24 38 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=5.26 $Y=3.33
+ $X2=5.04 $Y2=3.33
r81 24 25 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.26 $Y=3.33
+ $X2=5.425 $Y2=3.33
r82 23 41 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=5.59 $Y=3.33 $X2=6
+ $Y2=3.33
r83 23 25 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.59 $Y=3.33
+ $X2=5.425 $Y2=3.33
r84 21 35 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=4.21 $Y=3.33
+ $X2=4.08 $Y2=3.33
r85 21 22 8.88104 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=4.21 $Y=3.33
+ $X2=4.382 $Y2=3.33
r86 20 38 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=4.555 $Y=3.33
+ $X2=5.04 $Y2=3.33
r87 20 22 8.88104 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=4.555 $Y=3.33
+ $X2=4.382 $Y2=3.33
r88 16 19 19.2074 $w=3.28e-07 $l=5.5e-07 $layer=LI1_cond $X=5.425 $Y=2.265
+ $X2=5.425 $Y2=2.815
r89 14 25 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.425 $Y=3.245
+ $X2=5.425 $Y2=3.33
r90 14 19 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=5.425 $Y=3.245
+ $X2=5.425 $Y2=2.815
r91 10 22 1.03204 $w=3.45e-07 $l=8.5e-08 $layer=LI1_cond $X=4.382 $Y=3.245
+ $X2=4.382 $Y2=3.33
r92 10 12 8.35104 $w=3.43e-07 $l=2.5e-07 $layer=LI1_cond $X=4.382 $Y=3.245
+ $X2=4.382 $Y2=2.995
r93 3 19 600 $w=1.7e-07 $l=1.07034e-06 $layer=licon1_PDIFF $count=1 $X=5.225
+ $Y=1.84 $X2=5.425 $Y2=2.815
r94 3 16 600 $w=1.7e-07 $l=5.15388e-07 $layer=licon1_PDIFF $count=1 $X=5.225
+ $Y=1.84 $X2=5.425 $Y2=2.265
r95 2 12 600 $w=1.7e-07 $l=1.26934e-06 $layer=licon1_PDIFF $count=1 $X=4.14
+ $Y=1.84 $X2=4.38 $Y2=2.995
r96 1 45 600 $w=1.7e-07 $l=1.29455e-06 $layer=licon1_PDIFF $count=1 $X=3.095
+ $Y=1.84 $X2=3.27 $Y2=3.05
.ends

.subckt PM_SKY130_FD_SC_LS__MUX2I_2%A_115_74# 1 2 7 9 13 18 22 27 28
r63 27 28 9.33524 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=4.925 $Y=0.665
+ $X2=4.735 $Y2=0.665
r64 22 24 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=3.165 $Y=0.745
+ $X2=3.165 $Y2=0.835
r65 18 20 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=2.325 $Y=0.68
+ $X2=2.325 $Y2=0.835
r66 13 16 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=0.805 $Y=0.68
+ $X2=0.805 $Y2=0.8
r67 12 22 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.25 $Y=0.745
+ $X2=3.165 $Y2=0.745
r68 12 28 96.8824 $w=1.68e-07 $l=1.485e-06 $layer=LI1_cond $X=3.25 $Y=0.745
+ $X2=4.735 $Y2=0.745
r69 10 20 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.41 $Y=0.835
+ $X2=2.325 $Y2=0.835
r70 9 24 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.08 $Y=0.835
+ $X2=3.165 $Y2=0.835
r71 9 10 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.08 $Y=0.835
+ $X2=2.41 $Y2=0.835
r72 8 13 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.97 $Y=0.68
+ $X2=0.805 $Y2=0.68
r73 7 18 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.24 $Y=0.68
+ $X2=2.325 $Y2=0.68
r74 7 8 82.8556 $w=1.68e-07 $l=1.27e-06 $layer=LI1_cond $X=2.24 $Y=0.68 $X2=0.97
+ $Y2=0.68
r75 2 27 182 $w=1.7e-07 $l=2.43926e-07 $layer=licon1_NDIFF $count=1 $X=4.76
+ $Y=0.49 $X2=4.925 $Y2=0.665
r76 1 16 182 $w=1.7e-07 $l=5.32729e-07 $layer=licon1_NDIFF $count=1 $X=0.575
+ $Y=0.37 $X2=0.805 $Y2=0.8
.ends

.subckt PM_SKY130_FD_SC_LS__MUX2I_2%A_337_74# 1 2 10 15 16
c30 16 0 7.88763e-20 $X=3.65 $Y=1.13
r31 15 16 9.80174 $w=2.58e-07 $l=1.9e-07 $layer=LI1_cond $X=3.84 $Y=1.13
+ $X2=3.65 $Y2=1.13
r32 10 12 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=1.905 $Y=1.02
+ $X2=1.905 $Y2=1.175
r33 8 12 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.07 $Y=1.175
+ $X2=1.905 $Y2=1.175
r34 8 16 103.08 $w=1.68e-07 $l=1.58e-06 $layer=LI1_cond $X=2.07 $Y=1.175
+ $X2=3.65 $Y2=1.175
r35 2 15 182 $w=1.7e-07 $l=6.72458e-07 $layer=licon1_NDIFF $count=1 $X=3.675
+ $Y=0.49 $X2=3.84 $Y2=1.085
r36 1 10 182 $w=1.7e-07 $l=7.51997e-07 $layer=licon1_NDIFF $count=1 $X=1.685
+ $Y=0.37 $X2=1.905 $Y2=1.02
.ends

.subckt PM_SKY130_FD_SC_LS__MUX2I_2%VGND 1 2 3 12 16 20 23 24 26 27 28 40 46 47
+ 50
c64 12 0 3.11705e-20 $X=3.305 $Y=0.325
r65 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r66 47 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.52
+ $Y2=0
r67 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r68 44 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.615 $Y=0 $X2=5.45
+ $Y2=0
r69 44 46 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=5.615 $Y=0 $X2=6
+ $Y2=0
r70 43 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r71 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r72 40 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.285 $Y=0 $X2=5.45
+ $Y2=0
r73 40 42 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=5.285 $Y=0 $X2=5.04
+ $Y2=0
r74 39 43 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=5.04
+ $Y2=0
r75 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r76 31 35 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=3.12
+ $Y2=0
r77 31 32 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r78 28 39 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r79 28 32 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=3.12 $Y=0 $X2=0.24
+ $Y2=0
r80 28 35 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r81 26 38 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=4.21 $Y=0 $X2=4.08
+ $Y2=0
r82 26 27 8.88104 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=4.21 $Y=0 $X2=4.382
+ $Y2=0
r83 25 42 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=4.555 $Y=0 $X2=5.04
+ $Y2=0
r84 25 27 8.88104 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=4.555 $Y=0 $X2=4.382
+ $Y2=0
r85 23 35 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=3.14 $Y=0 $X2=3.12
+ $Y2=0
r86 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.14 $Y=0 $X2=3.305
+ $Y2=0
r87 22 38 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=3.47 $Y=0 $X2=4.08
+ $Y2=0
r88 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.47 $Y=0 $X2=3.305
+ $Y2=0
r89 18 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.45 $Y=0.085
+ $X2=5.45 $Y2=0
r90 18 20 19.9058 $w=3.28e-07 $l=5.7e-07 $layer=LI1_cond $X=5.45 $Y=0.085
+ $X2=5.45 $Y2=0.655
r91 14 27 1.03204 $w=3.45e-07 $l=8.5e-08 $layer=LI1_cond $X=4.382 $Y=0.085
+ $X2=4.382 $Y2=0
r92 14 16 8.01699 $w=3.43e-07 $l=2.4e-07 $layer=LI1_cond $X=4.382 $Y=0.085
+ $X2=4.382 $Y2=0.325
r93 10 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.305 $Y=0.085
+ $X2=3.305 $Y2=0
r94 10 12 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=3.305 $Y=0.085
+ $X2=3.305 $Y2=0.325
r95 3 20 182 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_NDIFF $count=1 $X=5.24
+ $Y=0.49 $X2=5.45 $Y2=0.655
r96 2 16 182 $w=1.7e-07 $l=2.96226e-07 $layer=licon1_NDIFF $count=1 $X=4.155
+ $Y=0.49 $X2=4.38 $Y2=0.325
r97 1 12 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=3.16
+ $Y=0.18 $X2=3.305 $Y2=0.325
.ends

