* File: sky130_fd_sc_ls__dlrtp_4.pex.spice
* Created: Wed Sep  2 11:04:11 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__DLRTP_4%D 3 5 7 8 12
c26 5 0 1.89325e-19 $X=0.505 $Y=1.895
r27 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.615 $X2=0.385 $Y2=1.615
r28 8 12 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=0.24 $Y=1.615
+ $X2=0.385 $Y2=1.615
r29 5 11 55.6741 $w=3.24e-07 $l=3.25331e-07 $layer=POLY_cond $X=0.505 $Y=1.895
+ $X2=0.407 $Y2=1.615
r30 5 7 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.505 $Y=1.895
+ $X2=0.505 $Y2=2.39
r31 1 11 38.5661 $w=3.24e-07 $l=2.04316e-07 $layer=POLY_cond $X=0.495 $Y=1.45
+ $X2=0.407 $Y2=1.615
r32 1 3 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=0.495 $Y=1.45
+ $X2=0.495 $Y2=0.905
.ends

.subckt PM_SKY130_FD_SC_LS__DLRTP_4%GATE 1 3 6 8
c33 6 0 3.6533e-19 $X=1.19 $Y=0.81
r34 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.165
+ $Y=1.615 $X2=1.165 $Y2=1.615
r35 4 11 38.6072 $w=2.91e-07 $l=1.77059e-07 $layer=POLY_cond $X=1.19 $Y=1.45
+ $X2=1.165 $Y2=1.615
r36 4 6 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=1.19 $Y=1.45 $X2=1.19
+ $Y2=0.81
r37 1 11 57.6553 $w=2.91e-07 $l=2.99333e-07 $layer=POLY_cond $X=1.125 $Y=1.895
+ $X2=1.165 $Y2=1.615
r38 1 3 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.125 $Y=1.895
+ $X2=1.125 $Y2=2.39
.ends

.subckt PM_SKY130_FD_SC_LS__DLRTP_4%A_240_394# 1 2 7 9 10 12 13 15 16 17 20 22
+ 23 24 29 31 32 35 36 37 41 48 52 53 54
c149 53 0 1.30138e-19 $X=3.985 $Y=1.39
c150 37 0 5.47968e-20 $X=3.005 $Y=0.34
c151 32 0 1.82632e-19 $X=2.835 $Y=0.855
c152 24 0 1.89325e-19 $X=1.46 $Y=2.075
c153 17 0 1.84143e-19 $X=3.215 $Y=1.765
c154 13 0 1.78764e-19 $X=3.125 $Y=1.885
r155 52 54 8.48463 $w=2.98e-07 $l=1.65e-07 $layer=LI1_cond $X=4 $Y=1.39 $X2=4
+ $Y2=1.225
r156 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.985
+ $Y=1.39 $X2=3.985 $Y2=1.39
r157 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.735
+ $Y=1.615 $X2=1.735 $Y2=1.615
r158 45 48 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=1.545 $Y=1.615
+ $X2=1.735 $Y2=1.615
r159 43 44 13.9266 $w=3.88e-07 $l=3.45e-07 $layer=LI1_cond $X=1.435 $Y=0.855
+ $X2=1.435 $Y2=1.2
r160 41 43 7.97845 $w=3.88e-07 $l=2.7e-07 $layer=LI1_cond $X=1.435 $Y=0.585
+ $X2=1.435 $Y2=0.855
r161 38 54 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=3.935 $Y=0.425
+ $X2=3.935 $Y2=1.225
r162 36 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.85 $Y=0.34
+ $X2=3.935 $Y2=0.425
r163 36 37 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=3.85 $Y=0.34
+ $X2=3.005 $Y2=0.34
r164 34 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.92 $Y=0.425
+ $X2=3.005 $Y2=0.34
r165 34 35 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.92 $Y=0.425
+ $X2=2.92 $Y2=0.77
r166 33 43 5.6248 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=1.63 $Y=0.855
+ $X2=1.435 $Y2=0.855
r167 32 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.835 $Y=0.855
+ $X2=2.92 $Y2=0.77
r168 32 33 78.615 $w=1.68e-07 $l=1.205e-06 $layer=LI1_cond $X=2.835 $Y=0.855
+ $X2=1.63 $Y2=0.855
r169 30 45 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.545 $Y=1.78
+ $X2=1.545 $Y2=1.615
r170 30 31 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.545 $Y=1.78
+ $X2=1.545 $Y2=1.95
r171 29 45 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.545 $Y=1.45
+ $X2=1.545 $Y2=1.615
r172 29 44 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.545 $Y=1.45
+ $X2=1.545 $Y2=1.2
r173 24 31 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.46 $Y=2.075
+ $X2=1.545 $Y2=1.95
r174 24 26 3.91831 $w=2.48e-07 $l=8.5e-08 $layer=LI1_cond $X=1.46 $Y=2.075
+ $X2=1.375 $Y2=2.075
r175 22 49 63.8244 $w=3.3e-07 $l=3.65e-07 $layer=POLY_cond $X=2.1 $Y=1.615
+ $X2=1.735 $Y2=1.615
r176 22 23 5.03009 $w=3.3e-07 $l=1.13049e-07 $layer=POLY_cond $X=2.1 $Y=1.615
+ $X2=2.19 $Y2=1.667
r177 18 53 38.7956 $w=3.51e-07 $l=2.56562e-07 $layer=POLY_cond $X=3.7 $Y=1.225
+ $X2=3.887 $Y2=1.39
r178 18 20 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=3.7 $Y=1.225
+ $X2=3.7 $Y2=0.58
r179 16 53 51.4957 $w=3.51e-07 $l=4.88748e-07 $layer=POLY_cond $X=3.625 $Y=1.765
+ $X2=3.887 $Y2=1.39
r180 16 17 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=3.625 $Y=1.765
+ $X2=3.215 $Y2=1.765
r181 13 17 26.9307 $w=1.5e-07 $l=1.58745e-07 $layer=POLY_cond $X=3.125 $Y=1.885
+ $X2=3.215 $Y2=1.765
r182 13 15 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.125 $Y=1.885
+ $X2=3.125 $Y2=2.46
r183 10 23 37.0704 $w=1.5e-07 $l=2.24375e-07 $layer=POLY_cond $X=2.205 $Y=1.45
+ $X2=2.19 $Y2=1.667
r184 10 12 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.205 $Y=1.45
+ $X2=2.205 $Y2=0.97
r185 7 23 37.0704 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=2.19 $Y=1.885
+ $X2=2.19 $Y2=1.667
r186 7 9 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.19 $Y=1.885
+ $X2=2.19 $Y2=2.38
r187 2 26 600 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=1.2
+ $Y=1.97 $X2=1.375 $Y2=2.115
r188 1 41 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.265
+ $Y=0.44 $X2=1.405 $Y2=0.585
.ends

.subckt PM_SKY130_FD_SC_LS__DLRTP_4%A_27_126# 1 2 9 11 13 16 18 19 21 22 25 27
+ 30
c89 30 0 1.08744e-19 $X=2.66 $Y=1.635
c90 25 0 1.25148e-19 $X=2.58 $Y=2.37
c91 11 0 1.75896e-19 $X=2.735 $Y=1.885
c92 9 0 1.68329e-19 $X=2.72 $Y=0.69
r93 30 33 8.51388 $w=2.88e-07 $l=1.65e-07 $layer=LI1_cond $X=2.64 $Y=1.635
+ $X2=2.64 $Y2=1.8
r94 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.66
+ $Y=1.635 $X2=2.66 $Y2=1.635
r95 27 28 6.86755 $w=6.04e-07 $l=3.4e-07 $layer=LI1_cond $X=0.485 $Y=2.115
+ $X2=0.485 $Y2=2.455
r96 25 33 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=2.58 $Y=2.37
+ $X2=2.58 $Y2=1.8
r97 23 28 8.35964 $w=1.7e-07 $l=3.7e-07 $layer=LI1_cond $X=0.855 $Y=2.455
+ $X2=0.485 $Y2=2.455
r98 22 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.495 $Y=2.455
+ $X2=2.58 $Y2=2.37
r99 22 23 106.995 $w=1.68e-07 $l=1.64e-06 $layer=LI1_cond $X=2.495 $Y=2.455
+ $X2=0.855 $Y2=2.455
r100 21 27 10.3858 $w=6.04e-07 $l=3.5812e-07 $layer=LI1_cond $X=0.77 $Y=1.95
+ $X2=0.485 $Y2=2.115
r101 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.77 $Y=1.28
+ $X2=0.77 $Y2=1.95
r102 18 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.685 $Y=1.195
+ $X2=0.77 $Y2=1.28
r103 18 19 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=0.685 $Y=1.195
+ $X2=0.445 $Y2=1.195
r104 14 19 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=1.11
+ $X2=0.445 $Y2=1.195
r105 14 16 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=0.28 $Y=1.11
+ $X2=0.28 $Y2=0.905
r106 11 31 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=2.735 $Y=1.885
+ $X2=2.66 $Y2=1.635
r107 11 13 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.735 $Y=1.885
+ $X2=2.735 $Y2=2.46
r108 7 31 38.5562 $w=2.99e-07 $l=1.92678e-07 $layer=POLY_cond $X=2.72 $Y=1.47
+ $X2=2.66 $Y2=1.635
r109 7 9 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=2.72 $Y=1.47 $X2=2.72
+ $Y2=0.69
r110 2 27 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.97 $X2=0.28 $Y2=2.115
r111 1 16 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.63 $X2=0.28 $Y2=0.905
.ends

.subckt PM_SKY130_FD_SC_LS__DLRTP_4%A_364_120# 1 2 9 10 12 14 15 16 18 20 21 22
+ 25 35 39 45 48
c106 35 0 1.75896e-19 $X=2.155 $Y=2.11
c107 25 0 1.30138e-19 $X=3.82 $Y=2.215
c108 16 0 1.82698e-19 $X=2.24 $Y=1.195
r109 45 48 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.2 $Y=1.285
+ $X2=3.2 $Y2=1.12
r110 44 46 8.58894 $w=3.83e-07 $l=1.65e-07 $layer=LI1_cond $X=3.147 $Y=1.285
+ $X2=3.147 $Y2=1.45
r111 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.2
+ $Y=1.285 $X2=3.2 $Y2=1.285
r112 37 39 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=2.93 $Y=2.055
+ $X2=3.04 $Y2=2.055
r113 33 35 11.7071 $w=1.78e-07 $l=1.9e-07 $layer=LI1_cond $X=1.965 $Y=2.11
+ $X2=2.155 $Y2=2.11
r114 29 31 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.975 $Y=1.195
+ $X2=2.155 $Y2=1.195
r115 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.82
+ $Y=2.215 $X2=3.82 $Y2=2.215
r116 23 25 24.0965 $w=3.28e-07 $l=6.9e-07 $layer=LI1_cond $X=3.82 $Y=2.905
+ $X2=3.82 $Y2=2.215
r117 21 23 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.655 $Y=2.99
+ $X2=3.82 $Y2=2.905
r118 21 22 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=3.655 $Y=2.99
+ $X2=3.015 $Y2=2.99
r119 20 39 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.04 $Y=1.97
+ $X2=3.04 $Y2=2.055
r120 20 46 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=3.04 $Y=1.97
+ $X2=3.04 $Y2=1.45
r121 18 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.93 $Y=2.905
+ $X2=3.015 $Y2=2.99
r122 17 37 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.93 $Y=2.14
+ $X2=2.93 $Y2=2.055
r123 17 18 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=2.93 $Y=2.14
+ $X2=2.93 $Y2=2.905
r124 16 31 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.24 $Y=1.195
+ $X2=2.155 $Y2=1.195
r125 15 44 2.69402 $w=3.83e-07 $l=9e-08 $layer=LI1_cond $X=3.147 $Y=1.195
+ $X2=3.147 $Y2=1.285
r126 15 16 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=2.955 $Y=1.195
+ $X2=2.24 $Y2=1.195
r127 14 35 1.06262 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=2.155 $Y=2.02
+ $X2=2.155 $Y2=2.11
r128 13 31 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.155 $Y=1.28
+ $X2=2.155 $Y2=1.195
r129 13 14 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=2.155 $Y=1.28
+ $X2=2.155 $Y2=2.02
r130 10 26 50.1894 $w=3.66e-07 $l=3.02903e-07 $layer=POLY_cond $X=3.66 $Y=2.465
+ $X2=3.777 $Y2=2.215
r131 10 12 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.66 $Y=2.465
+ $X2=3.66 $Y2=2.75
r132 9 48 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.125 $Y=0.69
+ $X2=3.125 $Y2=1.12
r133 2 33 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.82
+ $Y=1.96 $X2=1.965 $Y2=2.11
r134 1 29 182 $w=1.7e-07 $l=6.68019e-07 $layer=licon1_NDIFF $count=1 $X=1.82
+ $Y=0.6 $X2=1.975 $Y2=1.195
.ends

.subckt PM_SKY130_FD_SC_LS__DLRTP_4%A_797_48# 1 2 3 10 12 13 14 15 17 19 20 22
+ 25 27 29 32 34 36 39 41 43 46 48 54 58 59 63 72 81 84 85 86 87 97
c192 48 0 1.13625e-19 $X=5.11 $Y=2.272
c193 14 0 7.47035e-20 $X=4.135 $Y=0.94
r194 94 95 27.0642 $w=3.74e-07 $l=2.1e-07 $layer=POLY_cond $X=7.985 $Y=1.532
+ $X2=8.195 $Y2=1.532
r195 93 94 28.3529 $w=3.74e-07 $l=2.2e-07 $layer=POLY_cond $X=7.765 $Y=1.532
+ $X2=7.985 $Y2=1.532
r196 92 93 36.0856 $w=3.74e-07 $l=2.8e-07 $layer=POLY_cond $X=7.485 $Y=1.532
+ $X2=7.765 $Y2=1.532
r197 89 90 38.6631 $w=3.74e-07 $l=3e-07 $layer=POLY_cond $X=7.035 $Y=1.532
+ $X2=7.335 $Y2=1.532
r198 86 87 8.63679 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=6.765 $Y=1.545
+ $X2=6.935 $Y2=1.545
r199 81 83 10.2135 $w=1.78e-07 $l=1.65e-07 $layer=LI1_cond $X=5.27 $Y=0.785
+ $X2=5.27 $Y2=0.95
r200 73 97 9.66578 $w=3.74e-07 $l=7.5e-08 $layer=POLY_cond $X=8.43 $Y=1.532
+ $X2=8.505 $Y2=1.532
r201 73 95 30.2861 $w=3.74e-07 $l=2.35e-07 $layer=POLY_cond $X=8.43 $Y=1.532
+ $X2=8.195 $Y2=1.532
r202 72 73 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.43
+ $Y=1.465 $X2=8.43 $Y2=1.465
r203 70 92 9.66578 $w=3.74e-07 $l=7.5e-08 $layer=POLY_cond $X=7.41 $Y=1.532
+ $X2=7.485 $Y2=1.532
r204 70 90 9.66578 $w=3.74e-07 $l=7.5e-08 $layer=POLY_cond $X=7.41 $Y=1.532
+ $X2=7.335 $Y2=1.532
r205 69 72 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=7.41 $Y=1.465
+ $X2=8.43 $Y2=1.465
r206 69 87 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=7.41 $Y=1.465
+ $X2=6.935 $Y2=1.465
r207 69 70 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.41
+ $Y=1.465 $X2=7.41 $Y2=1.465
r208 66 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.44 $Y=1.705
+ $X2=6.275 $Y2=1.705
r209 66 86 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=6.44 $Y=1.705
+ $X2=6.765 $Y2=1.705
r210 61 85 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.275 $Y=1.79
+ $X2=6.275 $Y2=1.705
r211 61 63 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=6.275 $Y=1.79
+ $X2=6.275 $Y2=1.985
r212 60 84 2.11342 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.44 $Y=1.705
+ $X2=5.315 $Y2=1.705
r213 59 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.11 $Y=1.705
+ $X2=6.275 $Y2=1.705
r214 59 60 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.11 $Y=1.705
+ $X2=5.44 $Y2=1.705
r215 58 76 4.60977 $w=2.48e-07 $l=1e-07 $layer=LI1_cond $X=5.315 $Y=1.965
+ $X2=5.315 $Y2=2.065
r216 55 84 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=5.315 $Y=1.79
+ $X2=5.315 $Y2=1.705
r217 55 58 8.0671 $w=2.48e-07 $l=1.75e-07 $layer=LI1_cond $X=5.315 $Y=1.79
+ $X2=5.315 $Y2=1.965
r218 54 84 4.3182 $w=2.1e-07 $l=1.03078e-07 $layer=LI1_cond $X=5.275 $Y=1.62
+ $X2=5.315 $Y2=1.705
r219 54 83 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.275 $Y=1.62
+ $X2=5.275 $Y2=0.95
r220 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.36
+ $Y=2.215 $X2=4.36 $Y2=2.215
r221 48 78 9.18462 $w=3.28e-07 $l=2.63e-07 $layer=LI1_cond $X=5.275 $Y=2.272
+ $X2=5.275 $Y2=2.535
r222 48 76 7.93363 $w=3.28e-07 $l=2.07e-07 $layer=LI1_cond $X=5.275 $Y=2.272
+ $X2=5.275 $Y2=2.065
r223 48 50 20.8273 $w=4.13e-07 $l=7.5e-07 $layer=LI1_cond $X=5.11 $Y=2.272
+ $X2=4.36 $Y2=2.272
r224 44 97 15.4652 $w=3.74e-07 $l=2.85769e-07 $layer=POLY_cond $X=8.625 $Y=1.3
+ $X2=8.505 $Y2=1.532
r225 44 46 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=8.625 $Y=1.3
+ $X2=8.625 $Y2=0.74
r226 41 97 24.2268 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=8.505 $Y=1.765
+ $X2=8.505 $Y2=1.532
r227 41 43 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.505 $Y=1.765
+ $X2=8.505 $Y2=2.4
r228 37 95 24.2268 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=8.195 $Y=1.3
+ $X2=8.195 $Y2=1.532
r229 37 39 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=8.195 $Y=1.3
+ $X2=8.195 $Y2=0.74
r230 34 94 24.2268 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=7.985 $Y=1.765
+ $X2=7.985 $Y2=1.532
r231 34 36 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.985 $Y=1.765
+ $X2=7.985 $Y2=2.4
r232 30 93 24.2268 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=7.765 $Y=1.3
+ $X2=7.765 $Y2=1.532
r233 30 32 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=7.765 $Y=1.3
+ $X2=7.765 $Y2=0.74
r234 27 92 24.2268 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=7.485 $Y=1.765
+ $X2=7.485 $Y2=1.532
r235 27 29 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.485 $Y=1.765
+ $X2=7.485 $Y2=2.4
r236 23 90 24.2268 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=7.335 $Y=1.3
+ $X2=7.335 $Y2=1.532
r237 23 25 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=7.335 $Y=1.3
+ $X2=7.335 $Y2=0.74
r238 20 89 24.2268 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=7.035 $Y=1.765
+ $X2=7.035 $Y2=1.532
r239 20 22 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.035 $Y=1.765
+ $X2=7.035 $Y2=2.4
r240 19 51 38.5562 $w=2.99e-07 $l=1.98997e-07 $layer=POLY_cond $X=4.435 $Y=2.05
+ $X2=4.36 $Y2=2.215
r241 18 19 530.713 $w=1.5e-07 $l=1.035e-06 $layer=POLY_cond $X=4.435 $Y=1.015
+ $X2=4.435 $Y2=2.05
r242 15 51 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=4.285 $Y=2.465
+ $X2=4.36 $Y2=2.215
r243 15 17 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.285 $Y=2.465
+ $X2=4.285 $Y2=2.75
r244 13 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.36 $Y=0.94
+ $X2=4.435 $Y2=1.015
r245 13 14 115.372 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=4.36 $Y=0.94
+ $X2=4.135 $Y2=0.94
r246 10 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.06 $Y=0.865
+ $X2=4.135 $Y2=0.94
r247 10 12 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.06 $Y=0.865
+ $X2=4.06 $Y2=0.58
r248 3 63 300 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=2 $X=6.075
+ $Y=1.84 $X2=6.275 $Y2=1.985
r249 2 78 600 $w=1.7e-07 $l=7.66339e-07 $layer=licon1_PDIFF $count=1 $X=5.125
+ $Y=1.84 $X2=5.275 $Y2=2.535
r250 2 58 600 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_PDIFF $count=1 $X=5.125
+ $Y=1.84 $X2=5.275 $Y2=1.965
r251 1 81 182 $w=1.7e-07 $l=4.79922e-07 $layer=licon1_NDIFF $count=1 $X=5.125
+ $Y=0.37 $X2=5.265 $Y2=0.785
.ends

.subckt PM_SKY130_FD_SC_LS__DLRTP_4%A_640_74# 1 2 9 11 13 14 18 21 22 24 25 27
+ 34 35 36 39 43 44
c110 44 0 4.97491e-20 $X=3.325 $Y=2.405
c111 36 0 1.78764e-19 $X=3.68 $Y=1.81
c112 34 0 7.47035e-20 $X=3.595 $Y=1.725
c113 27 0 1.68329e-19 $X=3.51 $Y=0.76
c114 22 0 1.13625e-19 $X=5.5 $Y=1.765
r115 46 48 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=3.38 $Y=1.81
+ $X2=3.595 $Y2=1.81
r116 43 44 8.55689 $w=2.78e-07 $l=1.65e-07 $layer=LI1_cond $X=3.325 $Y=2.57
+ $X2=3.325 $Y2=2.405
r117 40 49 11.7243 $w=3.7e-07 $l=9e-08 $layer=POLY_cond $X=4.93 $Y=1.515
+ $X2=4.93 $Y2=1.425
r118 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.885
+ $Y=1.515 $X2=4.885 $Y2=1.515
r119 37 39 8.0671 $w=2.98e-07 $l=2.1e-07 $layer=LI1_cond $X=4.87 $Y=1.725
+ $X2=4.87 $Y2=1.515
r120 36 48 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.68 $Y=1.81
+ $X2=3.595 $Y2=1.81
r121 35 37 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=4.72 $Y=1.81
+ $X2=4.87 $Y2=1.725
r122 35 36 67.8503 $w=1.68e-07 $l=1.04e-06 $layer=LI1_cond $X=4.72 $Y=1.81
+ $X2=3.68 $Y2=1.81
r123 34 48 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.595 $Y=1.725
+ $X2=3.595 $Y2=1.81
r124 33 34 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=3.595 $Y=0.925
+ $X2=3.595 $Y2=1.725
r125 31 46 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.38 $Y=1.895
+ $X2=3.38 $Y2=1.81
r126 31 44 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=3.38 $Y=1.895
+ $X2=3.38 $Y2=2.405
r127 27 33 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.51 $Y=0.76
+ $X2=3.595 $Y2=0.925
r128 27 29 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=3.51 $Y=0.76
+ $X2=3.37 $Y2=0.76
r129 25 26 89.6095 $w=1.8e-07 $l=2.25e-07 $layer=POLY_cond $X=5.5 $Y=1.425
+ $X2=5.5 $Y2=1.2
r130 22 24 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=5.5 $Y=1.765
+ $X2=5.5 $Y2=2.26
r131 21 22 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.5 $Y=1.675 $X2=5.5
+ $Y2=1.765
r132 20 25 29.1532 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=5.5 $Y=1.5 $X2=5.5
+ $Y2=1.425
r133 20 21 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=5.5 $Y=1.5 $X2=5.5
+ $Y2=1.675
r134 18 26 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=5.485 $Y=0.69
+ $X2=5.485 $Y2=1.2
r135 15 49 23.9667 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=5.14 $Y=1.425
+ $X2=4.93 $Y2=1.425
r136 14 25 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=5.41 $Y=1.425 $X2=5.5
+ $Y2=1.425
r137 14 15 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=5.41 $Y=1.425
+ $X2=5.14 $Y2=1.425
r138 11 40 50.1287 $w=3.7e-07 $l=3.04138e-07 $layer=POLY_cond $X=5.05 $Y=1.765
+ $X2=4.93 $Y2=1.515
r139 11 13 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=5.05 $Y=1.765
+ $X2=5.05 $Y2=2.26
r140 7 49 27.3315 $w=3.7e-07 $l=1.52971e-07 $layer=POLY_cond $X=5.05 $Y=1.35
+ $X2=4.93 $Y2=1.425
r141 7 9 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.05 $Y=1.35 $X2=5.05
+ $Y2=0.69
r142 2 43 600 $w=1.7e-07 $l=6.80882e-07 $layer=licon1_PDIFF $count=1 $X=3.2
+ $Y=1.96 $X2=3.35 $Y2=2.57
r143 1 29 182 $w=1.7e-07 $l=4.67333e-07 $layer=licon1_NDIFF $count=1 $X=3.2
+ $Y=0.37 $X2=3.37 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_LS__DLRTP_4%RESET_B 1 3 5 6 8 9 11 13 14 16 17 18 28
c64 28 0 3.8972e-20 $X=6.5 $Y=1.285
r65 26 28 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=6.39 $Y=1.285
+ $X2=6.5 $Y2=1.285
r66 26 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.39
+ $Y=1.285 $X2=6.39 $Y2=1.285
r67 24 26 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=6.345 $Y=1.285
+ $X2=6.39 $Y2=1.285
r68 23 24 60.3271 $w=3.3e-07 $l=3.45e-07 $layer=POLY_cond $X=6 $Y=1.285
+ $X2=6.345 $Y2=1.285
r69 21 23 14.8632 $w=3.3e-07 $l=8.5e-08 $layer=POLY_cond $X=5.915 $Y=1.285 $X2=6
+ $Y2=1.285
r70 18 27 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=6.48 $Y=1.285 $X2=6.39
+ $Y2=1.285
r71 17 27 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=6 $Y=1.285 $X2=6.39
+ $Y2=1.285
r72 14 16 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=6.5 $Y=1.765 $X2=6.5
+ $Y2=2.26
r73 13 14 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.5 $Y=1.675 $X2=6.5
+ $Y2=1.765
r74 12 28 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.5 $Y=1.45 $X2=6.5
+ $Y2=1.285
r75 12 13 87.4597 $w=1.8e-07 $l=2.25e-07 $layer=POLY_cond $X=6.5 $Y=1.45 $X2=6.5
+ $Y2=1.675
r76 9 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.345 $Y=1.12
+ $X2=6.345 $Y2=1.285
r77 9 11 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=6.345 $Y=1.12
+ $X2=6.345 $Y2=0.69
r78 6 8 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=6 $Y=1.765 $X2=6
+ $Y2=2.26
r79 5 6 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6 $Y=1.675 $X2=6
+ $Y2=1.765
r80 4 23 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6 $Y=1.45 $X2=6
+ $Y2=1.285
r81 4 5 87.4597 $w=1.8e-07 $l=2.25e-07 $layer=POLY_cond $X=6 $Y=1.45 $X2=6
+ $Y2=1.675
r82 1 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.915 $Y=1.12
+ $X2=5.915 $Y2=1.285
r83 1 3 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=5.915 $Y=1.12
+ $X2=5.915 $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_LS__DLRTP_4%VPWR 1 2 3 4 5 6 7 26 30 34 38 42 48 50 52
+ 55 56 58 59 61 62 63 65 73 88 93 96 99 103
r113 102 103 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r114 96 97 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r115 93 94 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r116 91 103 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=8.88 $Y2=3.33
r117 90 91 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r118 88 102 4.58274 $w=1.7e-07 $l=2.62e-07 $layer=LI1_cond $X=8.595 $Y=3.33
+ $X2=8.857 $Y2=3.33
r119 88 90 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=8.595 $Y=3.33
+ $X2=8.4 $Y2=3.33
r120 87 91 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=8.4 $Y2=3.33
r121 86 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r122 84 87 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=7.44 $Y2=3.33
r123 83 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r124 81 84 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6.48 $Y2=3.33
r125 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r126 78 99 12.0744 $w=1.7e-07 $l=2.8e-07 $layer=LI1_cond $X=4.905 $Y=3.33
+ $X2=4.625 $Y2=3.33
r127 78 80 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=4.905 $Y=3.33
+ $X2=5.52 $Y2=3.33
r128 77 97 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=2.64 $Y2=3.33
r129 76 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r130 74 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.665 $Y=3.33
+ $X2=2.5 $Y2=3.33
r131 74 76 92.3155 $w=1.68e-07 $l=1.415e-06 $layer=LI1_cond $X=2.665 $Y=3.33
+ $X2=4.08 $Y2=3.33
r132 73 99 12.0744 $w=1.7e-07 $l=2.8e-07 $layer=LI1_cond $X=4.345 $Y=3.33
+ $X2=4.625 $Y2=3.33
r133 73 76 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=4.345 $Y=3.33
+ $X2=4.08 $Y2=3.33
r134 72 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r135 71 72 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r136 69 72 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r137 69 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r138 68 71 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r139 68 69 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r140 66 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.98 $Y=3.33
+ $X2=0.815 $Y2=3.33
r141 66 68 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.98 $Y=3.33
+ $X2=1.2 $Y2=3.33
r142 65 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.335 $Y=3.33
+ $X2=2.5 $Y2=3.33
r143 65 71 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.335 $Y=3.33
+ $X2=2.16 $Y2=3.33
r144 63 81 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r145 63 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r146 63 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r147 61 86 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=7.595 $Y=3.33
+ $X2=7.44 $Y2=3.33
r148 61 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.595 $Y=3.33
+ $X2=7.76 $Y2=3.33
r149 60 90 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=7.925 $Y=3.33
+ $X2=8.4 $Y2=3.33
r150 60 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.925 $Y=3.33
+ $X2=7.76 $Y2=3.33
r151 58 83 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=6.645 $Y=3.33
+ $X2=6.48 $Y2=3.33
r152 58 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.645 $Y=3.33
+ $X2=6.81 $Y2=3.33
r153 57 86 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=6.975 $Y=3.33
+ $X2=7.44 $Y2=3.33
r154 57 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.975 $Y=3.33
+ $X2=6.81 $Y2=3.33
r155 55 80 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=5.61 $Y=3.33 $X2=5.52
+ $Y2=3.33
r156 55 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.61 $Y=3.33
+ $X2=5.775 $Y2=3.33
r157 54 83 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=5.94 $Y=3.33
+ $X2=6.48 $Y2=3.33
r158 54 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.94 $Y=3.33
+ $X2=5.775 $Y2=3.33
r159 50 102 3.18343 $w=3.3e-07 $l=1.32868e-07 $layer=LI1_cond $X=8.76 $Y=3.245
+ $X2=8.857 $Y2=3.33
r160 50 52 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=8.76 $Y=3.245
+ $X2=8.76 $Y2=2.225
r161 46 62 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.76 $Y=3.245
+ $X2=7.76 $Y2=3.33
r162 46 48 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=7.76 $Y=3.245
+ $X2=7.76 $Y2=2.225
r163 42 45 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=6.81 $Y=2.045
+ $X2=6.81 $Y2=2.815
r164 40 59 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.81 $Y=3.245
+ $X2=6.81 $Y2=3.33
r165 40 45 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=6.81 $Y=3.245
+ $X2=6.81 $Y2=2.815
r166 36 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.775 $Y=3.245
+ $X2=5.775 $Y2=3.33
r167 36 38 41.034 $w=3.28e-07 $l=1.175e-06 $layer=LI1_cond $X=5.775 $Y=3.245
+ $X2=5.775 $Y2=2.07
r168 32 99 2.35715 $w=5.6e-07 $l=8.5e-08 $layer=LI1_cond $X=4.625 $Y=3.245
+ $X2=4.625 $Y2=3.33
r169 32 34 9.18417 $w=5.58e-07 $l=4.3e-07 $layer=LI1_cond $X=4.625 $Y=3.245
+ $X2=4.625 $Y2=2.815
r170 28 96 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.5 $Y=3.245 $X2=2.5
+ $Y2=3.33
r171 28 30 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=2.5 $Y=3.245
+ $X2=2.5 $Y2=2.805
r172 24 93 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=3.245
+ $X2=0.815 $Y2=3.33
r173 24 26 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.815 $Y=3.245
+ $X2=0.815 $Y2=2.875
r174 7 52 300 $w=1.7e-07 $l=4.66396e-07 $layer=licon1_PDIFF $count=2 $X=8.58
+ $Y=1.84 $X2=8.76 $Y2=2.225
r175 6 48 300 $w=1.7e-07 $l=4.74579e-07 $layer=licon1_PDIFF $count=2 $X=7.56
+ $Y=1.84 $X2=7.76 $Y2=2.225
r176 5 45 600 $w=1.7e-07 $l=1.08616e-06 $layer=licon1_PDIFF $count=1 $X=6.575
+ $Y=1.84 $X2=6.81 $Y2=2.815
r177 5 42 300 $w=1.7e-07 $l=3.21559e-07 $layer=licon1_PDIFF $count=2 $X=6.575
+ $Y=1.84 $X2=6.81 $Y2=2.045
r178 4 38 300 $w=1.7e-07 $l=3.14484e-07 $layer=licon1_PDIFF $count=2 $X=5.575
+ $Y=1.84 $X2=5.775 $Y2=2.07
r179 3 34 600 $w=1.7e-07 $l=3.85357e-07 $layer=licon1_PDIFF $count=1 $X=4.36
+ $Y=2.54 $X2=4.625 $Y2=2.815
r180 2 30 600 $w=1.7e-07 $l=9.55301e-07 $layer=licon1_PDIFF $count=1 $X=2.265
+ $Y=1.96 $X2=2.5 $Y2=2.805
r181 1 26 600 $w=1.7e-07 $l=1.01573e-06 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.97 $X2=0.815 $Y2=2.875
.ends

.subckt PM_SKY130_FD_SC_LS__DLRTP_4%Q 1 2 3 4 15 19 21 23 24 25 29 35 37 39 43
+ 45 48 49
r77 48 49 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=8.88 $Y=1.295
+ $X2=8.88 $Y2=1.665
r78 47 49 6.76434 $w=2.28e-07 $l=1.35e-07 $layer=LI1_cond $X=8.88 $Y=1.8
+ $X2=8.88 $Y2=1.665
r79 46 48 8.26753 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=8.88 $Y=1.13
+ $X2=8.88 $Y2=1.295
r80 40 45 4.08801 $w=2.5e-07 $l=9.5e-08 $layer=LI1_cond $X=8.505 $Y=1.005
+ $X2=8.41 $Y2=1.005
r81 39 46 6.8319 $w=2.5e-07 $l=1.73205e-07 $layer=LI1_cond $X=8.765 $Y=1.005
+ $X2=8.88 $Y2=1.13
r82 39 40 11.9854 $w=2.48e-07 $l=2.6e-07 $layer=LI1_cond $X=8.765 $Y=1.005
+ $X2=8.505 $Y2=1.005
r83 38 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.425 $Y=1.885
+ $X2=8.26 $Y2=1.885
r84 37 47 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=8.765 $Y=1.885
+ $X2=8.88 $Y2=1.8
r85 37 38 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=8.765 $Y=1.885
+ $X2=8.425 $Y2=1.885
r86 33 45 2.34704 $w=1.9e-07 $l=1.25e-07 $layer=LI1_cond $X=8.41 $Y=0.88
+ $X2=8.41 $Y2=1.005
r87 33 35 20.4306 $w=1.88e-07 $l=3.5e-07 $layer=LI1_cond $X=8.41 $Y=0.88
+ $X2=8.41 $Y2=0.53
r88 29 31 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=8.26 $Y=1.985
+ $X2=8.26 $Y2=2.815
r89 27 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.26 $Y=1.97 $X2=8.26
+ $Y2=1.885
r90 27 29 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=8.26 $Y=1.97
+ $X2=8.26 $Y2=1.985
r91 26 42 3.47681 $w=2.5e-07 $l=1.3e-07 $layer=LI1_cond $X=7.645 $Y=1.005
+ $X2=7.515 $Y2=1.005
r92 25 45 4.08801 $w=2.5e-07 $l=9.5e-08 $layer=LI1_cond $X=8.315 $Y=1.005
+ $X2=8.41 $Y2=1.005
r93 25 26 30.8855 $w=2.48e-07 $l=6.7e-07 $layer=LI1_cond $X=8.315 $Y=1.005
+ $X2=7.645 $Y2=1.005
r94 23 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.095 $Y=1.885
+ $X2=8.26 $Y2=1.885
r95 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.095 $Y=1.885
+ $X2=7.425 $Y2=1.885
r96 19 42 3.34309 $w=2.6e-07 $l=1.25e-07 $layer=LI1_cond $X=7.515 $Y=0.88
+ $X2=7.515 $Y2=1.005
r97 19 21 15.5137 $w=2.58e-07 $l=3.5e-07 $layer=LI1_cond $X=7.515 $Y=0.88
+ $X2=7.515 $Y2=0.53
r98 15 17 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=7.3 $Y=1.985 $X2=7.3
+ $Y2=2.815
r99 13 24 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=7.3 $Y=1.97
+ $X2=7.425 $Y2=1.885
r100 13 15 0.691466 $w=2.48e-07 $l=1.5e-08 $layer=LI1_cond $X=7.3 $Y=1.97
+ $X2=7.3 $Y2=1.985
r101 4 31 400 $w=1.7e-07 $l=1.07034e-06 $layer=licon1_PDIFF $count=1 $X=8.06
+ $Y=1.84 $X2=8.26 $Y2=2.815
r102 4 29 400 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=1 $X=8.06
+ $Y=1.84 $X2=8.26 $Y2=1.985
r103 3 17 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=7.11
+ $Y=1.84 $X2=7.26 $Y2=2.815
r104 3 15 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=7.11
+ $Y=1.84 $X2=7.26 $Y2=1.985
r105 2 45 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=8.27
+ $Y=0.37 $X2=8.41 $Y2=0.965
r106 2 35 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=8.27
+ $Y=0.37 $X2=8.41 $Y2=0.53
r107 1 42 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=7.41
+ $Y=0.37 $X2=7.55 $Y2=0.965
r108 1 21 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=7.41
+ $Y=0.37 $X2=7.55 $Y2=0.53
.ends

.subckt PM_SKY130_FD_SC_LS__DLRTP_4%VGND 1 2 3 4 5 6 7 26 30 34 38 40 44 48 50
+ 52 55 56 57 59 71 75 80 86 89 92 95 98 102
c122 44 0 3.8972e-20 $X=7.12 $Y=0.53
r123 101 102 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r124 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r125 95 96 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r126 93 96 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.96
+ $Y2=0
r127 92 93 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6 $Y2=0
r128 89 90 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r129 86 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r130 84 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=8.88
+ $Y2=0
r131 84 99 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=7.92
+ $Y2=0
r132 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r133 81 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.145 $Y=0 $X2=7.98
+ $Y2=0
r134 81 83 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=8.145 $Y=0 $X2=8.4
+ $Y2=0
r135 80 101 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=8.675 $Y=0
+ $X2=8.897 $Y2=0
r136 80 83 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=8.675 $Y=0 $X2=8.4
+ $Y2=0
r137 79 99 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=7.92
+ $Y2=0
r138 79 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=6.96
+ $Y2=0
r139 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r140 76 95 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=7.215 $Y=0 $X2=7.085
+ $Y2=0
r141 76 78 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=7.215 $Y=0
+ $X2=7.44 $Y2=0
r142 75 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.815 $Y=0 $X2=7.98
+ $Y2=0
r143 75 78 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=7.815 $Y=0
+ $X2=7.44 $Y2=0
r144 71 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.965 $Y=0 $X2=6.13
+ $Y2=0
r145 71 73 91.6631 $w=1.68e-07 $l=1.405e-06 $layer=LI1_cond $X=5.965 $Y=0
+ $X2=4.56 $Y2=0
r146 70 90 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.08 $Y=0
+ $X2=2.64 $Y2=0
r147 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r148 67 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.665 $Y=0 $X2=2.5
+ $Y2=0
r149 67 69 92.3155 $w=1.68e-07 $l=1.415e-06 $layer=LI1_cond $X=2.665 $Y=0
+ $X2=4.08 $Y2=0
r150 66 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r151 65 66 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r152 63 66 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r153 63 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r154 62 65 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r155 62 63 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r156 60 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.01 $Y=0 $X2=0.845
+ $Y2=0
r157 60 62 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.01 $Y=0 $X2=1.2
+ $Y2=0
r158 59 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.335 $Y=0 $X2=2.5
+ $Y2=0
r159 59 65 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.335 $Y=0
+ $X2=2.16 $Y2=0
r160 57 93 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.56 $Y=0 $X2=6
+ $Y2=0
r161 57 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r162 57 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r163 55 69 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=4.19 $Y=0 $X2=4.08
+ $Y2=0
r164 55 56 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.19 $Y=0 $X2=4.315
+ $Y2=0
r165 54 73 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=4.44 $Y=0 $X2=4.56
+ $Y2=0
r166 54 56 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.44 $Y=0 $X2=4.315
+ $Y2=0
r167 50 101 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=8.84 $Y=0.085
+ $X2=8.897 $Y2=0
r168 50 52 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=8.84 $Y=0.085
+ $X2=8.84 $Y2=0.53
r169 46 98 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.98 $Y=0.085
+ $X2=7.98 $Y2=0
r170 46 48 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=7.98 $Y=0.085
+ $X2=7.98 $Y2=0.53
r171 42 95 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=7.085 $Y=0.085
+ $X2=7.085 $Y2=0
r172 42 44 19.7245 $w=2.58e-07 $l=4.45e-07 $layer=LI1_cond $X=7.085 $Y=0.085
+ $X2=7.085 $Y2=0.53
r173 41 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.295 $Y=0 $X2=6.13
+ $Y2=0
r174 40 95 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.955 $Y=0 $X2=7.085
+ $Y2=0
r175 40 41 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=6.955 $Y=0
+ $X2=6.295 $Y2=0
r176 36 92 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.13 $Y=0.085
+ $X2=6.13 $Y2=0
r177 36 38 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=6.13 $Y=0.085
+ $X2=6.13 $Y2=0.515
r178 32 56 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.315 $Y=0.085
+ $X2=4.315 $Y2=0
r179 32 34 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=4.315 $Y=0.085
+ $X2=4.315 $Y2=0.58
r180 28 89 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.5 $Y=0.085 $X2=2.5
+ $Y2=0
r181 28 30 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.5 $Y=0.085
+ $X2=2.5 $Y2=0.515
r182 24 86 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.845 $Y=0.085
+ $X2=0.845 $Y2=0
r183 24 26 24.0965 $w=3.28e-07 $l=6.9e-07 $layer=LI1_cond $X=0.845 $Y=0.085
+ $X2=0.845 $Y2=0.775
r184 7 52 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=8.7
+ $Y=0.37 $X2=8.84 $Y2=0.53
r185 6 48 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=7.84
+ $Y=0.37 $X2=7.98 $Y2=0.53
r186 5 44 91 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=2 $X=6.975
+ $Y=0.37 $X2=7.12 $Y2=0.53
r187 4 38 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=5.99
+ $Y=0.37 $X2=6.13 $Y2=0.515
r188 3 34 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.135
+ $Y=0.37 $X2=4.275 $Y2=0.58
r189 2 30 182 $w=1.7e-07 $l=2.59037e-07 $layer=licon1_NDIFF $count=1 $X=2.28
+ $Y=0.6 $X2=2.5 $Y2=0.515
r190 1 26 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.63 $X2=0.845 $Y2=0.775
.ends

.subckt PM_SKY130_FD_SC_LS__DLRTP_4%A_938_74# 1 2 3 12 14 15 17 19 20 22 24
r47 22 29 2.91016 $w=2.6e-07 $l=9e-08 $layer=LI1_cond $X=6.595 $Y=0.77 $X2=6.595
+ $Y2=0.86
r48 22 24 11.5244 $w=2.58e-07 $l=2.6e-07 $layer=LI1_cond $X=6.595 $Y=0.77
+ $X2=6.595 $Y2=0.51
r49 21 27 4.10122 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=5.785 $Y=0.86
+ $X2=5.66 $Y2=0.86
r50 20 29 4.20357 $w=1.8e-07 $l=1.3e-07 $layer=LI1_cond $X=6.465 $Y=0.86
+ $X2=6.595 $Y2=0.86
r51 20 21 41.899 $w=1.78e-07 $l=6.8e-07 $layer=LI1_cond $X=6.465 $Y=0.86
+ $X2=5.785 $Y2=0.86
r52 17 27 2.95288 $w=2.5e-07 $l=9e-08 $layer=LI1_cond $X=5.66 $Y=0.77 $X2=5.66
+ $Y2=0.86
r53 17 19 12.6769 $w=2.48e-07 $l=2.75e-07 $layer=LI1_cond $X=5.66 $Y=0.77
+ $X2=5.66 $Y2=0.495
r54 16 19 2.0744 $w=2.48e-07 $l=4.5e-08 $layer=LI1_cond $X=5.66 $Y=0.45 $X2=5.66
+ $Y2=0.495
r55 14 16 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.535 $Y=0.365
+ $X2=5.66 $Y2=0.45
r56 14 15 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=5.535 $Y=0.365
+ $X2=5 $Y2=0.365
r57 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.835 $Y=0.45
+ $X2=5 $Y2=0.365
r58 10 12 2.26996 $w=3.28e-07 $l=6.5e-08 $layer=LI1_cond $X=4.835 $Y=0.45
+ $X2=4.835 $Y2=0.515
r59 3 29 182 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_NDIFF $count=1 $X=6.42
+ $Y=0.37 $X2=6.56 $Y2=0.86
r60 3 24 182 $w=1.7e-07 $l=1.9799e-07 $layer=licon1_NDIFF $count=1 $X=6.42
+ $Y=0.37 $X2=6.56 $Y2=0.51
r61 2 27 182 $w=1.7e-07 $l=5.50568e-07 $layer=licon1_NDIFF $count=1 $X=5.56
+ $Y=0.37 $X2=5.7 $Y2=0.855
r62 2 19 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=5.56
+ $Y=0.37 $X2=5.7 $Y2=0.495
r63 1 12 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=4.69
+ $Y=0.37 $X2=4.835 $Y2=0.515
.ends

