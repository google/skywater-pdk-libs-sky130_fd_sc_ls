* File: sky130_fd_sc_ls__a2111o_2.pxi.spice
* Created: Wed Sep  2 10:46:40 2020
* 
x_PM_SKY130_FD_SC_LS__A2111O_2%A_91_244# N_A_91_244#_M1013_s N_A_91_244#_M1004_d
+ N_A_91_244#_M1008_d N_A_91_244#_M1002_s N_A_91_244#_c_94_n N_A_91_244#_M1009_g
+ N_A_91_244#_c_81_n N_A_91_244#_M1005_g N_A_91_244#_c_82_n N_A_91_244#_M1006_g
+ N_A_91_244#_c_95_n N_A_91_244#_M1010_g N_A_91_244#_c_83_n N_A_91_244#_c_84_n
+ N_A_91_244#_c_85_n N_A_91_244#_c_97_n N_A_91_244#_c_98_n N_A_91_244#_c_99_n
+ N_A_91_244#_c_100_n N_A_91_244#_c_86_n N_A_91_244#_c_87_n N_A_91_244#_c_88_n
+ N_A_91_244#_c_89_n N_A_91_244#_c_90_n N_A_91_244#_c_91_n N_A_91_244#_c_92_n
+ N_A_91_244#_c_93_n PM_SKY130_FD_SC_LS__A2111O_2%A_91_244#
x_PM_SKY130_FD_SC_LS__A2111O_2%D1 N_D1_c_192_n N_D1_M1002_g N_D1_M1013_g D1 D1
+ PM_SKY130_FD_SC_LS__A2111O_2%D1
x_PM_SKY130_FD_SC_LS__A2111O_2%C1 N_C1_c_224_n N_C1_M1003_g N_C1_M1004_g C1 C1
+ C1 C1 N_C1_c_226_n PM_SKY130_FD_SC_LS__A2111O_2%C1
x_PM_SKY130_FD_SC_LS__A2111O_2%B1 N_B1_M1012_g N_B1_c_257_n N_B1_M1001_g B1
+ N_B1_c_258_n PM_SKY130_FD_SC_LS__A2111O_2%B1
x_PM_SKY130_FD_SC_LS__A2111O_2%A2 N_A2_c_287_n N_A2_M1011_g N_A2_M1007_g A2 A2
+ PM_SKY130_FD_SC_LS__A2111O_2%A2
x_PM_SKY130_FD_SC_LS__A2111O_2%A1 N_A1_M1008_g N_A1_c_322_n N_A1_M1000_g
+ N_A1_c_319_n A1 N_A1_c_320_n N_A1_c_321_n PM_SKY130_FD_SC_LS__A2111O_2%A1
x_PM_SKY130_FD_SC_LS__A2111O_2%VPWR N_VPWR_M1009_s N_VPWR_M1010_s N_VPWR_M1011_d
+ N_VPWR_c_349_n N_VPWR_c_350_n N_VPWR_c_351_n N_VPWR_c_352_n N_VPWR_c_353_n
+ N_VPWR_c_354_n VPWR N_VPWR_c_355_n N_VPWR_c_356_n N_VPWR_c_348_n
+ N_VPWR_c_358_n PM_SKY130_FD_SC_LS__A2111O_2%VPWR
x_PM_SKY130_FD_SC_LS__A2111O_2%X N_X_M1005_s N_X_M1009_d N_X_c_401_n X X X X X
+ PM_SKY130_FD_SC_LS__A2111O_2%X
x_PM_SKY130_FD_SC_LS__A2111O_2%A_630_368# N_A_630_368#_M1001_d
+ N_A_630_368#_M1000_d N_A_630_368#_c_425_n N_A_630_368#_c_422_n
+ N_A_630_368#_c_432_n N_A_630_368#_c_423_n N_A_630_368#_c_424_n
+ PM_SKY130_FD_SC_LS__A2111O_2%A_630_368#
x_PM_SKY130_FD_SC_LS__A2111O_2%VGND N_VGND_M1005_d N_VGND_M1006_d N_VGND_M1013_d
+ N_VGND_M1012_d N_VGND_c_448_n N_VGND_c_449_n N_VGND_c_450_n N_VGND_c_451_n
+ N_VGND_c_452_n N_VGND_c_453_n N_VGND_c_454_n VGND N_VGND_c_455_n
+ N_VGND_c_456_n N_VGND_c_457_n N_VGND_c_458_n N_VGND_c_459_n N_VGND_c_460_n
+ PM_SKY130_FD_SC_LS__A2111O_2%VGND
cc_1 VNB N_A_91_244#_c_81_n 0.021272f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=1.22
cc_2 VNB N_A_91_244#_c_82_n 0.0189136f $X=-0.19 $Y=-0.245 $X2=0.99 $Y2=1.22
cc_3 VNB N_A_91_244#_c_83_n 0.0144821f $X=-0.19 $Y=-0.245 $X2=1.275 $Y2=1.55
cc_4 VNB N_A_91_244#_c_84_n 0.00164528f $X=-0.19 $Y=-0.245 $X2=1.275 $Y2=1.95
cc_5 VNB N_A_91_244#_c_85_n 0.0247935f $X=-0.19 $Y=-0.245 $X2=1.78 $Y2=1.095
cc_6 VNB N_A_91_244#_c_86_n 0.0159334f $X=-0.19 $Y=-0.245 $X2=1.945 $Y2=0.515
cc_7 VNB N_A_91_244#_c_87_n 0.00754392f $X=-0.19 $Y=-0.245 $X2=2.76 $Y2=1.095
cc_8 VNB N_A_91_244#_c_88_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=2.845 $Y2=0.515
cc_9 VNB N_A_91_244#_c_89_n 0.0208031f $X=-0.19 $Y=-0.245 $X2=4.19 $Y2=1.095
cc_10 VNB N_A_91_244#_c_90_n 0.0281813f $X=-0.19 $Y=-0.245 $X2=4.355 $Y2=0.515
cc_11 VNB N_A_91_244#_c_91_n 0.00237125f $X=-0.19 $Y=-0.245 $X2=1.905 $Y2=1.095
cc_12 VNB N_A_91_244#_c_92_n 0.0086793f $X=-0.19 $Y=-0.245 $X2=2.885 $Y2=1.095
cc_13 VNB N_A_91_244#_c_93_n 0.0954235f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.492
cc_14 VNB N_D1_c_192_n 0.0257447f $X=-0.19 $Y=-0.245 $X2=1.82 $Y2=0.37
cc_15 VNB N_D1_M1013_g 0.0327351f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB D1 0.00943624f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_C1_c_224_n 0.0262092f $X=-0.19 $Y=-0.245 $X2=1.82 $Y2=0.37
cc_18 VNB N_C1_M1004_g 0.0238646f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_C1_c_226_n 0.00167125f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=0.74
cc_20 VNB N_B1_M1012_g 0.0272326f $X=-0.19 $Y=-0.245 $X2=4.215 $Y2=0.37
cc_21 VNB N_B1_c_257_n 0.0262417f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_B1_c_258_n 0.00166777f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A2_c_287_n 0.021813f $X=-0.19 $Y=-0.245 $X2=1.82 $Y2=0.37
cc_24 VNB N_A2_M1007_g 0.0254699f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB A2 0.00423229f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A1_M1008_g 0.0321165f $X=-0.19 $Y=-0.245 $X2=4.215 $Y2=0.37
cc_27 VNB N_A1_c_319_n 0.00982321f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A1_c_320_n 0.0439496f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.765
cc_29 VNB N_A1_c_321_n 0.00813406f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.4
cc_30 VNB N_VPWR_c_348_n 0.203486f $X=-0.19 $Y=-0.245 $X2=2.845 $Y2=0.515
cc_31 VNB N_X_c_401_n 0.00350677f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB X 8.01576e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_448_n 0.0141006f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.765
cc_34 VNB N_VGND_c_449_n 0.0502297f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.4
cc_35 VNB N_VGND_c_450_n 0.016021f $X=-0.19 $Y=-0.245 $X2=0.99 $Y2=1.22
cc_36 VNB N_VGND_c_451_n 0.00333244f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=2.4
cc_37 VNB N_VGND_c_452_n 0.00790127f $X=-0.19 $Y=-0.245 $X2=1.78 $Y2=1.095
cc_38 VNB N_VGND_c_453_n 0.0245715f $X=-0.19 $Y=-0.245 $X2=1.36 $Y2=2.035
cc_39 VNB N_VGND_c_454_n 0.00677473f $X=-0.19 $Y=-0.245 $X2=1.92 $Y2=2.12
cc_40 VNB N_VGND_c_455_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_456_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=2.845 $Y2=0.515
cc_42 VNB N_VGND_c_457_n 0.0334725f $X=-0.19 $Y=-0.245 $X2=4.355 $Y2=0.515
cc_43 VNB N_VGND_c_458_n 0.302009f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_459_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=1.92 $Y2=2.115
cc_45 VNB N_VGND_c_460_n 0.0103896f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.492
cc_46 VPB N_A_91_244#_c_94_n 0.0174317f $X=-0.19 $Y=1.66 $X2=0.545 $Y2=1.765
cc_47 VPB N_A_91_244#_c_95_n 0.0172125f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=1.765
cc_48 VPB N_A_91_244#_c_84_n 0.00889688f $X=-0.19 $Y=1.66 $X2=1.275 $Y2=1.95
cc_49 VPB N_A_91_244#_c_97_n 0.0241081f $X=-0.19 $Y=1.66 $X2=1.755 $Y2=2.035
cc_50 VPB N_A_91_244#_c_98_n 2.25523e-19 $X=-0.19 $Y=1.66 $X2=1.36 $Y2=2.035
cc_51 VPB N_A_91_244#_c_99_n 6.27129e-19 $X=-0.19 $Y=1.66 $X2=1.92 $Y2=2.12
cc_52 VPB N_A_91_244#_c_100_n 0.0139581f $X=-0.19 $Y=1.66 $X2=1.92 $Y2=2.815
cc_53 VPB N_A_91_244#_c_93_n 0.017011f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=1.492
cc_54 VPB N_D1_c_192_n 0.0306614f $X=-0.19 $Y=1.66 $X2=1.82 $Y2=0.37
cc_55 VPB D1 0.00917945f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_C1_c_224_n 0.0265214f $X=-0.19 $Y=1.66 $X2=1.82 $Y2=0.37
cc_57 VPB N_C1_c_226_n 0.00205145f $X=-0.19 $Y=1.66 $X2=0.56 $Y2=0.74
cc_58 VPB N_B1_c_257_n 0.0286834f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_B1_c_258_n 0.00278595f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_A2_c_287_n 0.0273391f $X=-0.19 $Y=1.66 $X2=1.82 $Y2=0.37
cc_61 VPB A2 0.00493565f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_A1_c_322_n 0.0216608f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_A1_c_319_n 0.00628072f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_A1_c_320_n 0.0145157f $X=-0.19 $Y=1.66 $X2=0.545 $Y2=1.765
cc_65 VPB N_A1_c_321_n 0.0117196f $X=-0.19 $Y=1.66 $X2=0.545 $Y2=2.4
cc_66 VPB N_VPWR_c_349_n 0.011928f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_350_n 0.0647053f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_351_n 0.0151005f $X=-0.19 $Y=1.66 $X2=0.56 $Y2=0.74
cc_69 VPB N_VPWR_c_352_n 0.00695663f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=1.765
cc_70 VPB N_VPWR_c_353_n 0.0650664f $X=-0.19 $Y=1.66 $X2=1.275 $Y2=1.55
cc_71 VPB N_VPWR_c_354_n 0.00691066f $X=-0.19 $Y=1.66 $X2=1.275 $Y2=1.95
cc_72 VPB N_VPWR_c_355_n 0.0184862f $X=-0.19 $Y=1.66 $X2=1.755 $Y2=2.035
cc_73 VPB N_VPWR_c_356_n 0.0236066f $X=-0.19 $Y=1.66 $X2=2.885 $Y2=0.515
cc_74 VPB N_VPWR_c_348_n 0.105208f $X=-0.19 $Y=1.66 $X2=2.845 $Y2=0.515
cc_75 VPB N_VPWR_c_358_n 0.00614127f $X=-0.19 $Y=1.66 $X2=4.355 $Y2=0.515
cc_76 VPB X 0.00357774f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_A_630_368#_c_422_n 0.00327016f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_A_630_368#_c_423_n 0.00743317f $X=-0.19 $Y=1.66 $X2=0.545 $Y2=1.765
cc_79 VPB N_A_630_368#_c_424_n 0.0360166f $X=-0.19 $Y=1.66 $X2=0.545 $Y2=2.4
cc_80 N_A_91_244#_c_84_n N_D1_c_192_n 6.74178e-19 $X=1.275 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_81 N_A_91_244#_c_99_n N_D1_c_192_n 0.00332314f $X=1.92 $Y=2.12 $X2=-0.19
+ $Y2=-0.245
cc_82 N_A_91_244#_c_100_n N_D1_c_192_n 0.0124227f $X=1.92 $Y=2.815 $X2=-0.19
+ $Y2=-0.245
cc_83 N_A_91_244#_c_87_n N_D1_c_192_n 0.00130632f $X=2.76 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_84 N_A_91_244#_c_91_n N_D1_c_192_n 0.00291196f $X=1.905 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_85 N_A_91_244#_c_93_n N_D1_c_192_n 0.0033277f $X=0.995 $Y=1.492 $X2=-0.19
+ $Y2=-0.245
cc_86 N_A_91_244#_c_86_n N_D1_M1013_g 0.00159319f $X=1.945 $Y=0.515 $X2=0 $Y2=0
cc_87 N_A_91_244#_c_87_n N_D1_M1013_g 0.0140963f $X=2.76 $Y=1.095 $X2=0 $Y2=0
cc_88 N_A_91_244#_c_83_n D1 0.0146967f $X=1.275 $Y=1.55 $X2=0 $Y2=0
cc_89 N_A_91_244#_c_84_n D1 0.0169762f $X=1.275 $Y=1.95 $X2=0 $Y2=0
cc_90 N_A_91_244#_c_85_n D1 0.0173741f $X=1.78 $Y=1.095 $X2=0 $Y2=0
cc_91 N_A_91_244#_c_97_n D1 0.0153495f $X=1.755 $Y=2.035 $X2=0 $Y2=0
cc_92 N_A_91_244#_c_99_n D1 0.0265363f $X=1.92 $Y=2.12 $X2=0 $Y2=0
cc_93 N_A_91_244#_c_87_n D1 0.0183652f $X=2.76 $Y=1.095 $X2=0 $Y2=0
cc_94 N_A_91_244#_c_91_n D1 0.0220075f $X=1.905 $Y=1.095 $X2=0 $Y2=0
cc_95 N_A_91_244#_c_93_n D1 9.56934e-19 $X=0.995 $Y=1.492 $X2=0 $Y2=0
cc_96 N_A_91_244#_c_100_n N_C1_c_224_n 0.00123511f $X=1.92 $Y=2.815 $X2=-0.19
+ $Y2=-0.245
cc_97 N_A_91_244#_c_87_n N_C1_c_224_n 0.0011446f $X=2.76 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_98 N_A_91_244#_c_87_n N_C1_M1004_g 0.0132453f $X=2.76 $Y=1.095 $X2=0 $Y2=0
cc_99 N_A_91_244#_c_88_n N_C1_M1004_g 3.97481e-19 $X=2.845 $Y=0.515 $X2=0 $Y2=0
cc_100 N_A_91_244#_c_87_n N_C1_c_226_n 0.0244947f $X=2.76 $Y=1.095 $X2=0 $Y2=0
cc_101 N_A_91_244#_c_92_n N_C1_c_226_n 0.00124816f $X=2.885 $Y=1.095 $X2=0 $Y2=0
cc_102 N_A_91_244#_c_88_n N_B1_M1012_g 0.00979642f $X=2.845 $Y=0.515 $X2=0 $Y2=0
cc_103 N_A_91_244#_c_89_n N_B1_M1012_g 0.0123033f $X=4.19 $Y=1.095 $X2=0 $Y2=0
cc_104 N_A_91_244#_c_92_n N_B1_M1012_g 0.00154264f $X=2.885 $Y=1.095 $X2=0 $Y2=0
cc_105 N_A_91_244#_c_89_n N_B1_c_257_n 0.00126003f $X=4.19 $Y=1.095 $X2=0 $Y2=0
cc_106 N_A_91_244#_c_89_n N_B1_c_258_n 0.0229301f $X=4.19 $Y=1.095 $X2=0 $Y2=0
cc_107 N_A_91_244#_c_92_n N_B1_c_258_n 0.00196319f $X=2.885 $Y=1.095 $X2=0 $Y2=0
cc_108 N_A_91_244#_c_89_n N_A2_c_287_n 0.00465926f $X=4.19 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_109 N_A_91_244#_c_88_n N_A2_M1007_g 9.95982e-19 $X=2.845 $Y=0.515 $X2=0 $Y2=0
cc_110 N_A_91_244#_c_89_n N_A2_M1007_g 0.0149964f $X=4.19 $Y=1.095 $X2=0 $Y2=0
cc_111 N_A_91_244#_c_90_n N_A2_M1007_g 0.00218322f $X=4.355 $Y=0.515 $X2=0 $Y2=0
cc_112 N_A_91_244#_c_89_n A2 0.0544915f $X=4.19 $Y=1.095 $X2=0 $Y2=0
cc_113 N_A_91_244#_c_89_n N_A1_M1008_g 0.0135439f $X=4.19 $Y=1.095 $X2=0 $Y2=0
cc_114 N_A_91_244#_c_90_n N_A1_M1008_g 0.0125612f $X=4.355 $Y=0.515 $X2=0 $Y2=0
cc_115 N_A_91_244#_c_89_n N_A1_c_319_n 0.00676585f $X=4.19 $Y=1.095 $X2=0 $Y2=0
cc_116 N_A_91_244#_c_89_n N_A1_c_320_n 0.00121887f $X=4.19 $Y=1.095 $X2=0 $Y2=0
cc_117 N_A_91_244#_c_89_n N_A1_c_321_n 0.0132907f $X=4.19 $Y=1.095 $X2=0 $Y2=0
cc_118 N_A_91_244#_c_84_n N_VPWR_M1010_s 0.0021071f $X=1.275 $Y=1.95 $X2=0 $Y2=0
cc_119 N_A_91_244#_c_98_n N_VPWR_M1010_s 0.00504875f $X=1.36 $Y=2.035 $X2=0
+ $Y2=0
cc_120 N_A_91_244#_c_94_n N_VPWR_c_350_n 0.008783f $X=0.545 $Y=1.765 $X2=0 $Y2=0
cc_121 N_A_91_244#_c_94_n N_VPWR_c_351_n 5.61406e-19 $X=0.545 $Y=1.765 $X2=0
+ $Y2=0
cc_122 N_A_91_244#_c_95_n N_VPWR_c_351_n 0.012555f $X=0.995 $Y=1.765 $X2=0 $Y2=0
cc_123 N_A_91_244#_c_97_n N_VPWR_c_351_n 0.00198924f $X=1.755 $Y=2.035 $X2=0
+ $Y2=0
cc_124 N_A_91_244#_c_98_n N_VPWR_c_351_n 0.0152886f $X=1.36 $Y=2.035 $X2=0 $Y2=0
cc_125 N_A_91_244#_c_100_n N_VPWR_c_351_n 0.0335663f $X=1.92 $Y=2.815 $X2=0
+ $Y2=0
cc_126 N_A_91_244#_c_100_n N_VPWR_c_353_n 0.0145938f $X=1.92 $Y=2.815 $X2=0
+ $Y2=0
cc_127 N_A_91_244#_c_94_n N_VPWR_c_355_n 0.00445602f $X=0.545 $Y=1.765 $X2=0
+ $Y2=0
cc_128 N_A_91_244#_c_95_n N_VPWR_c_355_n 0.00413917f $X=0.995 $Y=1.765 $X2=0
+ $Y2=0
cc_129 N_A_91_244#_c_94_n N_VPWR_c_348_n 0.00861209f $X=0.545 $Y=1.765 $X2=0
+ $Y2=0
cc_130 N_A_91_244#_c_95_n N_VPWR_c_348_n 0.00817726f $X=0.995 $Y=1.765 $X2=0
+ $Y2=0
cc_131 N_A_91_244#_c_100_n N_VPWR_c_348_n 0.0120466f $X=1.92 $Y=2.815 $X2=0
+ $Y2=0
cc_132 N_A_91_244#_c_81_n N_X_c_401_n 0.00267578f $X=0.56 $Y=1.22 $X2=0 $Y2=0
cc_133 N_A_91_244#_c_82_n N_X_c_401_n 0.00139568f $X=0.99 $Y=1.22 $X2=0 $Y2=0
cc_134 N_A_91_244#_c_83_n N_X_c_401_n 0.0319992f $X=1.275 $Y=1.55 $X2=0 $Y2=0
cc_135 N_A_91_244#_c_93_n N_X_c_401_n 0.0251153f $X=0.995 $Y=1.492 $X2=0 $Y2=0
cc_136 N_A_91_244#_c_94_n X 0.0162357f $X=0.545 $Y=1.765 $X2=0 $Y2=0
cc_137 N_A_91_244#_c_95_n X 0.00857619f $X=0.995 $Y=1.765 $X2=0 $Y2=0
cc_138 N_A_91_244#_c_84_n X 0.0191743f $X=1.275 $Y=1.95 $X2=0 $Y2=0
cc_139 N_A_91_244#_c_98_n X 0.00870628f $X=1.36 $Y=2.035 $X2=0 $Y2=0
cc_140 N_A_91_244#_c_93_n X 0.0201749f $X=0.995 $Y=1.492 $X2=0 $Y2=0
cc_141 N_A_91_244#_c_83_n N_VGND_M1006_d 0.00288214f $X=1.275 $Y=1.55 $X2=0
+ $Y2=0
cc_142 N_A_91_244#_c_87_n N_VGND_M1013_d 0.00218982f $X=2.76 $Y=1.095 $X2=0
+ $Y2=0
cc_143 N_A_91_244#_c_89_n N_VGND_M1012_d 0.0059981f $X=4.19 $Y=1.095 $X2=0 $Y2=0
cc_144 N_A_91_244#_c_81_n N_VGND_c_449_n 0.0159149f $X=0.56 $Y=1.22 $X2=0 $Y2=0
cc_145 N_A_91_244#_c_82_n N_VGND_c_449_n 5.58177e-19 $X=0.99 $Y=1.22 $X2=0 $Y2=0
cc_146 N_A_91_244#_c_93_n N_VGND_c_449_n 0.00155918f $X=0.995 $Y=1.492 $X2=0
+ $Y2=0
cc_147 N_A_91_244#_c_81_n N_VGND_c_450_n 4.71636e-19 $X=0.56 $Y=1.22 $X2=0 $Y2=0
cc_148 N_A_91_244#_c_82_n N_VGND_c_450_n 0.0128397f $X=0.99 $Y=1.22 $X2=0 $Y2=0
cc_149 N_A_91_244#_c_83_n N_VGND_c_450_n 0.020572f $X=1.275 $Y=1.55 $X2=0 $Y2=0
cc_150 N_A_91_244#_c_85_n N_VGND_c_450_n 7.22336e-19 $X=1.78 $Y=1.095 $X2=0
+ $Y2=0
cc_151 N_A_91_244#_c_86_n N_VGND_c_450_n 0.0217548f $X=1.945 $Y=0.515 $X2=0
+ $Y2=0
cc_152 N_A_91_244#_c_93_n N_VGND_c_450_n 0.00147793f $X=0.995 $Y=1.492 $X2=0
+ $Y2=0
cc_153 N_A_91_244#_c_86_n N_VGND_c_451_n 0.0186004f $X=1.945 $Y=0.515 $X2=0
+ $Y2=0
cc_154 N_A_91_244#_c_87_n N_VGND_c_451_n 0.020332f $X=2.76 $Y=1.095 $X2=0 $Y2=0
cc_155 N_A_91_244#_c_88_n N_VGND_c_451_n 0.0186004f $X=2.845 $Y=0.515 $X2=0
+ $Y2=0
cc_156 N_A_91_244#_c_88_n N_VGND_c_452_n 0.018474f $X=2.845 $Y=0.515 $X2=0 $Y2=0
cc_157 N_A_91_244#_c_89_n N_VGND_c_452_n 0.0389277f $X=4.19 $Y=1.095 $X2=0 $Y2=0
cc_158 N_A_91_244#_c_90_n N_VGND_c_452_n 0.01706f $X=4.355 $Y=0.515 $X2=0 $Y2=0
cc_159 N_A_91_244#_c_86_n N_VGND_c_453_n 0.011066f $X=1.945 $Y=0.515 $X2=0 $Y2=0
cc_160 N_A_91_244#_c_81_n N_VGND_c_455_n 0.00383152f $X=0.56 $Y=1.22 $X2=0 $Y2=0
cc_161 N_A_91_244#_c_82_n N_VGND_c_455_n 0.00383152f $X=0.99 $Y=1.22 $X2=0 $Y2=0
cc_162 N_A_91_244#_c_88_n N_VGND_c_456_n 0.0109942f $X=2.845 $Y=0.515 $X2=0
+ $Y2=0
cc_163 N_A_91_244#_c_90_n N_VGND_c_457_n 0.0145639f $X=4.355 $Y=0.515 $X2=0
+ $Y2=0
cc_164 N_A_91_244#_c_81_n N_VGND_c_458_n 0.0075754f $X=0.56 $Y=1.22 $X2=0 $Y2=0
cc_165 N_A_91_244#_c_82_n N_VGND_c_458_n 0.0075754f $X=0.99 $Y=1.22 $X2=0 $Y2=0
cc_166 N_A_91_244#_c_86_n N_VGND_c_458_n 0.00915947f $X=1.945 $Y=0.515 $X2=0
+ $Y2=0
cc_167 N_A_91_244#_c_88_n N_VGND_c_458_n 0.00904371f $X=2.845 $Y=0.515 $X2=0
+ $Y2=0
cc_168 N_A_91_244#_c_90_n N_VGND_c_458_n 0.0119984f $X=4.355 $Y=0.515 $X2=0
+ $Y2=0
cc_169 N_A_91_244#_c_89_n A_771_74# 0.00366293f $X=4.19 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_170 N_D1_c_192_n N_C1_c_224_n 0.0933439f $X=2.145 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_171 D1 N_C1_c_224_n 0.00255274f $X=2.075 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_172 N_D1_M1013_g N_C1_M1004_g 0.0281796f $X=2.16 $Y=0.74 $X2=0 $Y2=0
cc_173 N_D1_c_192_n N_C1_c_226_n 0.00456229f $X=2.145 $Y=1.765 $X2=0 $Y2=0
cc_174 D1 N_C1_c_226_n 0.036282f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_175 N_D1_c_192_n N_VPWR_c_351_n 0.00383557f $X=2.145 $Y=1.765 $X2=0 $Y2=0
cc_176 N_D1_c_192_n N_VPWR_c_353_n 0.00445602f $X=2.145 $Y=1.765 $X2=0 $Y2=0
cc_177 N_D1_c_192_n N_VPWR_c_348_n 0.00862666f $X=2.145 $Y=1.765 $X2=0 $Y2=0
cc_178 N_D1_M1013_g N_VGND_c_451_n 0.0140324f $X=2.16 $Y=0.74 $X2=0 $Y2=0
cc_179 N_D1_M1013_g N_VGND_c_453_n 0.00383152f $X=2.16 $Y=0.74 $X2=0 $Y2=0
cc_180 N_D1_M1013_g N_VGND_c_458_n 0.00762539f $X=2.16 $Y=0.74 $X2=0 $Y2=0
cc_181 N_C1_M1004_g N_B1_M1012_g 0.0195038f $X=2.63 $Y=0.74 $X2=0 $Y2=0
cc_182 N_C1_c_224_n N_B1_c_257_n 0.0587037f $X=2.535 $Y=1.765 $X2=0 $Y2=0
cc_183 N_C1_c_226_n N_B1_c_257_n 0.0137282f $X=2.61 $Y=1.515 $X2=0 $Y2=0
cc_184 N_C1_c_224_n N_B1_c_258_n 0.00127792f $X=2.535 $Y=1.765 $X2=0 $Y2=0
cc_185 N_C1_c_226_n N_B1_c_258_n 0.0277337f $X=2.61 $Y=1.515 $X2=0 $Y2=0
cc_186 N_C1_c_224_n N_VPWR_c_353_n 0.00303293f $X=2.535 $Y=1.765 $X2=0 $Y2=0
cc_187 N_C1_c_226_n N_VPWR_c_353_n 0.00909385f $X=2.61 $Y=1.515 $X2=0 $Y2=0
cc_188 N_C1_c_224_n N_VPWR_c_348_n 0.00372419f $X=2.535 $Y=1.765 $X2=0 $Y2=0
cc_189 N_C1_c_226_n N_VPWR_c_348_n 0.0106888f $X=2.61 $Y=1.515 $X2=0 $Y2=0
cc_190 N_C1_c_226_n A_522_368# 0.0141247f $X=2.61 $Y=1.515 $X2=-0.19 $Y2=-0.245
cc_191 N_C1_c_226_n N_A_630_368#_c_425_n 0.00784442f $X=2.61 $Y=1.515 $X2=0
+ $Y2=0
cc_192 N_C1_c_224_n N_A_630_368#_c_422_n 0.00107752f $X=2.535 $Y=1.765 $X2=0
+ $Y2=0
cc_193 N_C1_c_226_n N_A_630_368#_c_422_n 0.0338558f $X=2.61 $Y=1.515 $X2=0 $Y2=0
cc_194 N_C1_M1004_g N_VGND_c_451_n 0.0110514f $X=2.63 $Y=0.74 $X2=0 $Y2=0
cc_195 N_C1_M1004_g N_VGND_c_456_n 0.00383152f $X=2.63 $Y=0.74 $X2=0 $Y2=0
cc_196 N_C1_M1004_g N_VGND_c_458_n 0.00757637f $X=2.63 $Y=0.74 $X2=0 $Y2=0
cc_197 N_B1_c_257_n N_A2_c_287_n 0.0450961f $X=3.075 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_198 N_B1_c_258_n N_A2_c_287_n 7.1218e-19 $X=3.15 $Y=1.515 $X2=-0.19
+ $Y2=-0.245
cc_199 N_B1_M1012_g N_A2_M1007_g 0.0187776f $X=3.06 $Y=0.74 $X2=0 $Y2=0
cc_200 N_B1_c_257_n A2 0.00230997f $X=3.075 $Y=1.765 $X2=0 $Y2=0
cc_201 N_B1_c_258_n A2 0.0366314f $X=3.15 $Y=1.515 $X2=0 $Y2=0
cc_202 N_B1_c_257_n N_VPWR_c_352_n 6.63234e-19 $X=3.075 $Y=1.765 $X2=0 $Y2=0
cc_203 N_B1_c_257_n N_VPWR_c_353_n 0.00445602f $X=3.075 $Y=1.765 $X2=0 $Y2=0
cc_204 N_B1_c_257_n N_VPWR_c_348_n 0.00860014f $X=3.075 $Y=1.765 $X2=0 $Y2=0
cc_205 N_B1_c_257_n N_A_630_368#_c_425_n 0.00339629f $X=3.075 $Y=1.765 $X2=0
+ $Y2=0
cc_206 N_B1_c_258_n N_A_630_368#_c_425_n 0.0131798f $X=3.15 $Y=1.515 $X2=0 $Y2=0
cc_207 N_B1_c_257_n N_A_630_368#_c_422_n 0.0128839f $X=3.075 $Y=1.765 $X2=0
+ $Y2=0
cc_208 N_B1_M1012_g N_VGND_c_451_n 5.17244e-19 $X=3.06 $Y=0.74 $X2=0 $Y2=0
cc_209 N_B1_M1012_g N_VGND_c_452_n 0.00589272f $X=3.06 $Y=0.74 $X2=0 $Y2=0
cc_210 N_B1_M1012_g N_VGND_c_456_n 0.00434272f $X=3.06 $Y=0.74 $X2=0 $Y2=0
cc_211 N_B1_M1012_g N_VGND_c_458_n 0.0082236f $X=3.06 $Y=0.74 $X2=0 $Y2=0
cc_212 N_A2_M1007_g N_A1_M1008_g 0.0442642f $X=3.78 $Y=0.74 $X2=0 $Y2=0
cc_213 N_A2_c_287_n N_A1_c_322_n 0.0264386f $X=3.615 $Y=1.765 $X2=0 $Y2=0
cc_214 A2 N_A1_c_322_n 0.00205152f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_215 N_A2_c_287_n N_A1_c_319_n 0.0470099f $X=3.615 $Y=1.765 $X2=0 $Y2=0
cc_216 A2 N_A1_c_319_n 0.0166734f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_217 A2 N_A1_c_321_n 0.0346459f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_218 N_A2_c_287_n N_VPWR_c_352_n 0.010989f $X=3.615 $Y=1.765 $X2=0 $Y2=0
cc_219 N_A2_c_287_n N_VPWR_c_353_n 0.00413917f $X=3.615 $Y=1.765 $X2=0 $Y2=0
cc_220 N_A2_c_287_n N_VPWR_c_348_n 0.00818558f $X=3.615 $Y=1.765 $X2=0 $Y2=0
cc_221 N_A2_c_287_n N_A_630_368#_c_422_n 0.00507867f $X=3.615 $Y=1.765 $X2=0
+ $Y2=0
cc_222 N_A2_c_287_n N_A_630_368#_c_432_n 0.0164172f $X=3.615 $Y=1.765 $X2=0
+ $Y2=0
cc_223 A2 N_A_630_368#_c_432_n 0.0477758f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_224 N_A2_c_287_n N_A_630_368#_c_424_n 8.54227e-19 $X=3.615 $Y=1.765 $X2=0
+ $Y2=0
cc_225 N_A2_M1007_g N_VGND_c_452_n 0.0215908f $X=3.78 $Y=0.74 $X2=0 $Y2=0
cc_226 N_A2_M1007_g N_VGND_c_457_n 0.00383152f $X=3.78 $Y=0.74 $X2=0 $Y2=0
cc_227 N_A2_M1007_g N_VGND_c_458_n 0.0075694f $X=3.78 $Y=0.74 $X2=0 $Y2=0
cc_228 N_A1_c_322_n N_VPWR_c_352_n 0.00734374f $X=4.155 $Y=1.765 $X2=0 $Y2=0
cc_229 N_A1_c_322_n N_VPWR_c_356_n 0.00445602f $X=4.155 $Y=1.765 $X2=0 $Y2=0
cc_230 N_A1_c_322_n N_VPWR_c_348_n 0.00861623f $X=4.155 $Y=1.765 $X2=0 $Y2=0
cc_231 N_A1_c_322_n N_A_630_368#_c_432_n 0.0129877f $X=4.155 $Y=1.765 $X2=0
+ $Y2=0
cc_232 N_A1_c_322_n N_A_630_368#_c_423_n 9.1767e-19 $X=4.155 $Y=1.765 $X2=0
+ $Y2=0
cc_233 N_A1_c_320_n N_A_630_368#_c_423_n 0.0050009f $X=4.53 $Y=1.515 $X2=0 $Y2=0
cc_234 N_A1_c_321_n N_A_630_368#_c_423_n 0.0159673f $X=4.53 $Y=1.515 $X2=0 $Y2=0
cc_235 N_A1_c_322_n N_A_630_368#_c_424_n 0.0103816f $X=4.155 $Y=1.765 $X2=0
+ $Y2=0
cc_236 N_A1_M1008_g N_VGND_c_452_n 0.00189477f $X=4.14 $Y=0.74 $X2=0 $Y2=0
cc_237 N_A1_M1008_g N_VGND_c_457_n 0.00434272f $X=4.14 $Y=0.74 $X2=0 $Y2=0
cc_238 N_A1_M1008_g N_VGND_c_458_n 0.00824773f $X=4.14 $Y=0.74 $X2=0 $Y2=0
cc_239 N_VPWR_c_350_n X 0.0763579f $X=0.32 $Y=1.985 $X2=0 $Y2=0
cc_240 N_VPWR_c_351_n X 0.0472744f $X=1.22 $Y=2.455 $X2=0 $Y2=0
cc_241 N_VPWR_c_355_n X 0.0112472f $X=1.055 $Y=3.33 $X2=0 $Y2=0
cc_242 N_VPWR_c_348_n X 0.00927661f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_243 N_VPWR_c_352_n N_A_630_368#_c_422_n 0.0271521f $X=3.86 $Y=2.455 $X2=0
+ $Y2=0
cc_244 N_VPWR_c_353_n N_A_630_368#_c_422_n 0.0163786f $X=3.675 $Y=3.33 $X2=0
+ $Y2=0
cc_245 N_VPWR_c_348_n N_A_630_368#_c_422_n 0.0135239f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_246 N_VPWR_M1011_d N_A_630_368#_c_432_n 0.0059417f $X=3.69 $Y=1.84 $X2=0
+ $Y2=0
cc_247 N_VPWR_c_352_n N_A_630_368#_c_432_n 0.0234793f $X=3.86 $Y=2.455 $X2=0
+ $Y2=0
cc_248 N_VPWR_c_352_n N_A_630_368#_c_424_n 0.0266947f $X=3.86 $Y=2.455 $X2=0
+ $Y2=0
cc_249 N_VPWR_c_356_n N_A_630_368#_c_424_n 0.0145938f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_250 N_VPWR_c_348_n N_A_630_368#_c_424_n 0.0120466f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_251 N_X_c_401_n N_VGND_c_449_n 0.0293294f $X=0.775 $Y=0.515 $X2=0 $Y2=0
cc_252 N_X_c_401_n N_VGND_c_450_n 0.0182488f $X=0.775 $Y=0.515 $X2=0 $Y2=0
cc_253 N_X_c_401_n N_VGND_c_455_n 0.00749631f $X=0.775 $Y=0.515 $X2=0 $Y2=0
cc_254 N_X_c_401_n N_VGND_c_458_n 0.0062048f $X=0.775 $Y=0.515 $X2=0 $Y2=0
