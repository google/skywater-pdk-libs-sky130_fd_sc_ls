* File: sky130_fd_sc_ls__o21ba_2.pex.spice
* Created: Fri Aug 28 13:46:00 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__O21BA_2%B1_N 3 5 7 8 12
c27 5 0 1.07789e-19 $X=0.505 $Y=1.765
c28 3 0 5.63373e-20 $X=0.485 $Y=0.645
r29 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.29
+ $Y=1.465 $X2=0.29 $Y2=1.465
r30 8 12 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=0.29 $Y=1.665 $X2=0.29
+ $Y2=1.465
r31 5 11 56.2063 $w=3.85e-07 $l=3.65377e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.36 $Y2=1.465
r32 5 7 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.26
r33 1 11 39.305 $w=3.85e-07 $l=2.18746e-07 $layer=POLY_cond $X=0.485 $Y=1.3
+ $X2=0.36 $Y2=1.465
r34 1 3 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.485 $Y=1.3
+ $X2=0.485 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_LS__O21BA_2%A_177_48# 1 2 9 11 13 16 18 20 21 25 31 33
+ 38 41 42 47
c101 38 0 1.92475e-19 $X=2.465 $Y=1.095
r102 46 47 14.8933 $w=3.56e-07 $l=1.1e-07 $layer=POLY_cond $X=1.39 $Y=1.532
+ $X2=1.5 $Y2=1.532
r103 45 46 46.0337 $w=3.56e-07 $l=3.4e-07 $layer=POLY_cond $X=1.05 $Y=1.532
+ $X2=1.39 $Y2=1.532
r104 44 45 12.1854 $w=3.56e-07 $l=9e-08 $layer=POLY_cond $X=0.96 $Y=1.532
+ $X2=1.05 $Y2=1.532
r105 41 43 12.7457 $w=3.93e-07 $l=4.25e-07 $layer=LI1_cond $X=2.577 $Y=1.985
+ $X2=2.577 $Y2=2.41
r106 41 42 8.6272 $w=3.93e-07 $l=1.65e-07 $layer=LI1_cond $X=2.577 $Y=1.985
+ $X2=2.577 $Y2=1.82
r107 36 47 2.0309 $w=3.56e-07 $l=1.5e-08 $layer=POLY_cond $X=1.515 $Y=1.532
+ $X2=1.5 $Y2=1.532
r108 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.515
+ $Y=1.465 $X2=1.515 $Y2=1.465
r109 33 35 17.702 $w=2.55e-07 $l=3.7e-07 $layer=LI1_cond $X=1.515 $Y=1.095
+ $X2=1.515 $Y2=1.465
r110 31 43 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=2.61 $Y=2.695
+ $X2=2.61 $Y2=2.41
r111 27 38 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.465 $Y=1.18
+ $X2=2.465 $Y2=1.095
r112 27 42 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=2.465 $Y=1.18
+ $X2=2.465 $Y2=1.82
r113 23 38 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=2.105 $Y=1.095
+ $X2=2.465 $Y2=1.095
r114 23 25 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=2.105 $Y=1.01
+ $X2=2.105 $Y2=0.515
r115 22 33 3.11056 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.68 $Y=1.095
+ $X2=1.515 $Y2=1.095
r116 21 23 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=1.98 $Y=1.095
+ $X2=2.105 $Y2=1.095
r117 21 22 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.98 $Y=1.095
+ $X2=1.68 $Y2=1.095
r118 18 47 23.0368 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=1.5 $Y=1.765
+ $X2=1.5 $Y2=1.532
r119 18 20 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.5 $Y=1.765
+ $X2=1.5 $Y2=2.4
r120 14 46 23.0368 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=1.39 $Y=1.3
+ $X2=1.39 $Y2=1.532
r121 14 16 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.39 $Y=1.3
+ $X2=1.39 $Y2=0.74
r122 11 45 23.0368 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=1.05 $Y=1.765
+ $X2=1.05 $Y2=1.532
r123 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.05 $Y=1.765
+ $X2=1.05 $Y2=2.4
r124 7 44 23.0368 $w=1.5e-07 $l=1.87e-07 $layer=POLY_cond $X=0.96 $Y=1.345
+ $X2=0.96 $Y2=1.532
r125 7 9 310.223 $w=1.5e-07 $l=6.05e-07 $layer=POLY_cond $X=0.96 $Y=1.345
+ $X2=0.96 $Y2=0.74
r126 2 41 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.46
+ $Y=1.84 $X2=2.61 $Y2=1.985
r127 2 31 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=2.46
+ $Y=1.84 $X2=2.61 $Y2=2.695
r128 1 25 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=2.01
+ $Y=0.37 $X2=2.145 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__O21BA_2%A_27_74# 1 2 9 11 13 14 15 18 20 21 23 24 28
+ 32
c87 15 0 1.92475e-19 $X=2.285 $Y=1.35
c88 9 0 2.05372e-19 $X=2.36 $Y=0.74
r89 32 33 4.70956 $w=5.44e-07 $l=2.1e-07 $layer=LI1_cond $X=0.455 $Y=2.115
+ $X2=0.455 $Y2=2.325
r90 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.055
+ $Y=1.515 $X2=2.055 $Y2=1.515
r91 26 28 26.11 $w=3.18e-07 $l=7.25e-07 $layer=LI1_cond $X=2.05 $Y=2.24 $X2=2.05
+ $Y2=1.515
r92 25 33 7.68949 $w=1.7e-07 $l=3.4e-07 $layer=LI1_cond $X=0.795 $Y=2.325
+ $X2=0.455 $Y2=2.325
r93 24 26 7.68211 $w=1.7e-07 $l=1.9799e-07 $layer=LI1_cond $X=1.89 $Y=2.325
+ $X2=2.05 $Y2=2.24
r94 24 25 71.4385 $w=1.68e-07 $l=1.095e-06 $layer=LI1_cond $X=1.89 $Y=2.325
+ $X2=0.795 $Y2=2.325
r95 23 32 9.98939 $w=5.44e-07 $l=3.27261e-07 $layer=LI1_cond $X=0.71 $Y=1.95
+ $X2=0.455 $Y2=2.115
r96 22 23 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=0.71 $Y=1.13
+ $X2=0.71 $Y2=1.95
r97 20 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.625 $Y=1.045
+ $X2=0.71 $Y2=1.13
r98 20 21 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.625 $Y=1.045
+ $X2=0.355 $Y2=1.045
r99 16 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.23 $Y=0.96
+ $X2=0.355 $Y2=1.045
r100 16 18 14.5208 $w=2.48e-07 $l=3.15e-07 $layer=LI1_cond $X=0.23 $Y=0.96
+ $X2=0.23 $Y2=0.645
r101 14 29 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=2.285 $Y=1.515
+ $X2=2.055 $Y2=1.515
r102 14 15 5.03009 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.285 $Y=1.515
+ $X2=2.285 $Y2=1.35
r103 11 15 37.0704 $w=1.5e-07 $l=4.62304e-07 $layer=POLY_cond $X=2.385 $Y=1.765
+ $X2=2.285 $Y2=1.35
r104 11 13 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.385 $Y=1.765
+ $X2=2.385 $Y2=2.34
r105 7 15 37.0704 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.36 $Y=1.35
+ $X2=2.285 $Y2=1.35
r106 7 9 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.36 $Y=1.35 $X2=2.36
+ $Y2=0.74
r107 2 32 300 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.115
r108 1 18 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.27 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_LS__O21BA_2%A2 1 3 4 6 7
c32 7 0 1.75261e-19 $X=3.12 $Y=1.295
c33 1 0 2.53695e-20 $X=2.79 $Y=1.22
r34 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.88
+ $Y=1.385 $X2=2.88 $Y2=1.385
r35 7 11 7.47531 $w=3.68e-07 $l=2.4e-07 $layer=LI1_cond $X=3.12 $Y=1.365
+ $X2=2.88 $Y2=1.365
r36 4 10 77.2841 $w=2.7e-07 $l=4.01871e-07 $layer=POLY_cond $X=2.835 $Y=1.765
+ $X2=2.88 $Y2=1.385
r37 4 6 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.835 $Y=1.765
+ $X2=2.835 $Y2=2.34
r38 1 10 38.9026 $w=2.7e-07 $l=2.05122e-07 $layer=POLY_cond $X=2.79 $Y=1.22
+ $X2=2.88 $Y2=1.385
r39 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.79 $Y=1.22 $X2=2.79
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__O21BA_2%A1 1 3 4 6 7
c22 7 0 2.53695e-20 $X=3.6 $Y=1.295
r23 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.57
+ $Y=1.385 $X2=3.57 $Y2=1.385
r24 7 11 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=3.57 $Y=1.295 $X2=3.57
+ $Y2=1.385
r25 4 10 38.7084 $w=3.43e-07 $l=2.22486e-07 $layer=POLY_cond $X=3.36 $Y=1.22
+ $X2=3.495 $Y2=1.385
r26 4 6 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.36 $Y=1.22 $X2=3.36
+ $Y2=0.74
r27 1 10 68.9212 $w=3.43e-07 $l=4.48776e-07 $layer=POLY_cond $X=3.345 $Y=1.765
+ $X2=3.495 $Y2=1.385
r28 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.345 $Y=1.765
+ $X2=3.345 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_LS__O21BA_2%VPWR 1 2 3 14 16 18 22 24 29 35 38 48
r44 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r45 41 44 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r46 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r47 38 41 10.9789 $w=6.68e-07 $l=6.15e-07 $layer=LI1_cond $X=1.9 $Y=2.715
+ $X2=1.9 $Y2=3.33
r48 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r49 33 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r50 33 44 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.16 $Y2=3.33
r51 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r52 30 41 9.03384 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=2.235 $Y=3.33
+ $X2=1.9 $Y2=3.33
r53 30 32 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=2.235 $Y=3.33
+ $X2=3.12 $Y2=3.33
r54 29 47 4.76062 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=3.405 $Y=3.33
+ $X2=3.622 $Y2=3.33
r55 29 32 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=3.405 $Y=3.33
+ $X2=3.12 $Y2=3.33
r56 28 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r57 28 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r58 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r59 25 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.98 $Y=3.33
+ $X2=0.815 $Y2=3.33
r60 25 27 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.98 $Y=3.33 $X2=1.2
+ $Y2=3.33
r61 24 41 9.03384 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=1.565 $Y=3.33
+ $X2=1.9 $Y2=3.33
r62 24 27 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.565 $Y=3.33
+ $X2=1.2 $Y2=3.33
r63 22 44 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.16 $Y2=3.33
r64 22 42 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r65 18 21 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=3.57 $Y=1.985
+ $X2=3.57 $Y2=2.695
r66 16 47 3.00555 $w=3.3e-07 $l=1.07912e-07 $layer=LI1_cond $X=3.57 $Y=3.245
+ $X2=3.622 $Y2=3.33
r67 16 21 19.2074 $w=3.28e-07 $l=5.5e-07 $layer=LI1_cond $X=3.57 $Y=3.245
+ $X2=3.57 $Y2=2.695
r68 12 35 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=3.245
+ $X2=0.815 $Y2=3.33
r69 12 14 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=0.815 $Y=3.245
+ $X2=0.815 $Y2=2.745
r70 3 21 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=3.42
+ $Y=1.84 $X2=3.57 $Y2=2.695
r71 3 18 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=3.42
+ $Y=1.84 $X2=3.57 $Y2=1.985
r72 2 38 300 $w=1.7e-07 $l=1.09487e-06 $layer=licon1_PDIFF $count=2 $X=1.575
+ $Y=1.84 $X2=2.07 $Y2=2.715
r73 1 14 600 $w=1.7e-07 $l=1.01573e-06 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.84 $X2=0.815 $Y2=2.745
.ends

.subckt PM_SKY130_FD_SC_LS__O21BA_2%X 1 2 8 12 14 15 26
c35 15 0 5.63373e-20 $X=1.115 $Y=0.84
c36 12 0 1.07789e-19 $X=1.275 $Y=1.985
r37 19 26 1.3969 $w=3.28e-07 $l=4e-08 $layer=LI1_cond $X=1.175 $Y=0.965
+ $X2=1.175 $Y2=0.925
r38 15 28 7.69388 $w=3.28e-07 $l=1.43e-07 $layer=LI1_cond $X=1.175 $Y=0.987
+ $X2=1.175 $Y2=1.13
r39 15 19 0.768295 $w=3.28e-07 $l=2.2e-08 $layer=LI1_cond $X=1.175 $Y=0.987
+ $X2=1.175 $Y2=0.965
r40 15 26 0.803218 $w=3.28e-07 $l=2.3e-08 $layer=LI1_cond $X=1.175 $Y=0.902
+ $X2=1.175 $Y2=0.925
r41 14 15 13.515 $w=3.28e-07 $l=3.87e-07 $layer=LI1_cond $X=1.175 $Y=0.515
+ $X2=1.175 $Y2=0.902
r42 9 12 8.29759 $w=2.48e-07 $l=1.8e-07 $layer=LI1_cond $X=1.095 $Y=1.945
+ $X2=1.275 $Y2=1.945
r43 8 9 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.095 $Y=1.82
+ $X2=1.095 $Y2=1.945
r44 8 28 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.095 $Y=1.82
+ $X2=1.095 $Y2=1.13
r45 2 12 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.125
+ $Y=1.84 $X2=1.275 $Y2=1.985
r46 1 14 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.035
+ $Y=0.37 $X2=1.175 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__O21BA_2%VGND 1 2 3 12 16 20 23 24 25 31 35 42 43 46
+ 49
r56 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r57 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r58 43 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r59 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r60 40 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.24 $Y=0 $X2=3.075
+ $Y2=0
r61 40 42 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=3.24 $Y=0 $X2=3.6
+ $Y2=0
r62 39 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r63 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r64 36 46 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.77 $Y=0 $X2=1.645
+ $Y2=0
r65 36 38 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=1.77 $Y=0 $X2=2.64
+ $Y2=0
r66 35 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.91 $Y=0 $X2=3.075
+ $Y2=0
r67 35 38 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=2.91 $Y=0 $X2=2.64
+ $Y2=0
r68 34 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r69 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r70 31 46 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.52 $Y=0 $X2=1.645
+ $Y2=0
r71 31 33 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.52 $Y=0 $X2=1.2
+ $Y2=0
r72 29 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r73 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r74 25 39 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.64
+ $Y2=0
r75 25 47 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r76 23 28 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.535 $Y=0 $X2=0.24
+ $Y2=0
r77 23 24 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.535 $Y=0 $X2=0.66
+ $Y2=0
r78 22 33 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=0.785 $Y=0 $X2=1.2
+ $Y2=0
r79 22 24 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.785 $Y=0 $X2=0.66
+ $Y2=0
r80 18 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.075 $Y=0.085
+ $X2=3.075 $Y2=0
r81 18 20 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=3.075 $Y=0.085
+ $X2=3.075 $Y2=0.335
r82 14 46 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.645 $Y=0.085
+ $X2=1.645 $Y2=0
r83 14 16 25.5842 $w=2.48e-07 $l=5.55e-07 $layer=LI1_cond $X=1.645 $Y=0.085
+ $X2=1.645 $Y2=0.64
r84 10 24 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.66 $Y=0.085
+ $X2=0.66 $Y2=0
r85 10 12 24.2013 $w=2.48e-07 $l=5.25e-07 $layer=LI1_cond $X=0.66 $Y=0.085
+ $X2=0.66 $Y2=0.61
r86 3 20 182 $w=1.7e-07 $l=2.26826e-07 $layer=licon1_NDIFF $count=1 $X=2.865
+ $Y=0.37 $X2=3.075 $Y2=0.335
r87 2 16 182 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_NDIFF $count=1 $X=1.465
+ $Y=0.37 $X2=1.605 $Y2=0.64
r88 1 12 182 $w=1.7e-07 $l=3.01993e-07 $layer=licon1_NDIFF $count=1 $X=0.56
+ $Y=0.37 $X2=0.7 $Y2=0.61
.ends

.subckt PM_SKY130_FD_SC_LS__O21BA_2%A_487_74# 1 2 7 10 15
c28 7 0 3.01108e-20 $X=3.41 $Y=0.755
r29 15 17 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=3.575 $Y=0.515
+ $X2=3.575 $Y2=0.755
r30 10 12 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=2.575 $Y=0.595
+ $X2=2.575 $Y2=0.755
r31 8 12 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.74 $Y=0.755
+ $X2=2.575 $Y2=0.755
r32 7 17 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.41 $Y=0.755
+ $X2=3.575 $Y2=0.755
r33 7 8 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.41 $Y=0.755 $X2=2.74
+ $Y2=0.755
r34 2 15 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.435
+ $Y=0.37 $X2=3.575 $Y2=0.515
r35 1 10 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=2.435
+ $Y=0.37 $X2=2.575 $Y2=0.595
.ends

