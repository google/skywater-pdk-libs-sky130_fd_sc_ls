* File: sky130_fd_sc_ls__dfstp_4.pex.spice
* Created: Wed Sep  2 11:01:56 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__DFSTP_4%D 2 4 7 9 11 12 13 17 18 21
c35 18 0 1.4091e-19 $X=0.64 $Y=1.145
r36 21 23 39.7991 $w=3.9e-07 $l=1.65e-07 $layer=POLY_cond $X=0.61 $Y=1.825
+ $X2=0.61 $Y2=1.99
r37 21 22 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.64
+ $Y=1.825 $X2=0.64 $Y2=1.825
r38 17 19 45.456 $w=3.9e-07 $l=1.65e-07 $layer=POLY_cond $X=0.61 $Y=1.145
+ $X2=0.61 $Y2=0.98
r39 17 18 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.64
+ $Y=1.145 $X2=0.64 $Y2=1.145
r40 13 22 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=0.64 $Y=1.665
+ $X2=0.64 $Y2=1.825
r41 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.64 $Y=1.295
+ $X2=0.64 $Y2=1.665
r42 12 18 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=0.64 $Y=1.295
+ $X2=0.64 $Y2=1.145
r43 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.505 $Y=2.445
+ $X2=0.505 $Y2=2.73
r44 7 19 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=0.495 $Y=0.58 $X2=0.495
+ $Y2=0.98
r45 4 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.505 $Y=2.355 $X2=0.505
+ $Y2=2.445
r46 4 23 141.879 $w=1.8e-07 $l=3.65e-07 $layer=POLY_cond $X=0.505 $Y=2.355
+ $X2=0.505 $Y2=1.99
r47 2 21 4.27811 $w=3.9e-07 $l=3e-08 $layer=POLY_cond $X=0.61 $Y=1.795 $X2=0.61
+ $Y2=1.825
r48 1 17 4.27811 $w=3.9e-07 $l=3e-08 $layer=POLY_cond $X=0.61 $Y=1.175 $X2=0.61
+ $Y2=1.145
r49 1 2 88.4142 $w=3.9e-07 $l=6.2e-07 $layer=POLY_cond $X=0.61 $Y=1.175 $X2=0.61
+ $Y2=1.795
.ends

.subckt PM_SKY130_FD_SC_LS__DFSTP_4%CLK 1 3 4 6 7
c32 4 0 2.37719e-19 $X=1.515 $Y=1.765
r33 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.465
+ $Y=1.385 $X2=1.465 $Y2=1.385
r34 7 11 6.69663 $w=3.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.68 $Y=1.365
+ $X2=1.465 $Y2=1.365
r35 4 10 77.2841 $w=2.7e-07 $l=4.04228e-07 $layer=POLY_cond $X=1.515 $Y=1.765
+ $X2=1.465 $Y2=1.385
r36 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.515 $Y=1.765
+ $X2=1.515 $Y2=2.4
r37 1 10 38.9026 $w=2.7e-07 $l=1.74714e-07 $layer=POLY_cond $X=1.485 $Y=1.22
+ $X2=1.465 $Y2=1.385
r38 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.485 $Y=1.22 $X2=1.485
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__DFSTP_4%A_398_74# 1 2 7 9 10 14 18 19 21 24 28 30 31
+ 32 33 36 43 44 47 48 51 52 53 55 56 57 61 62 63 66 67 69 70 71 74 76 84
c261 70 0 8.24247e-20 $X=6.53 $Y=1.285
c262 69 0 2.80241e-20 $X=6.53 $Y=1.285
c263 67 0 1.99261e-20 $X=3.71 $Y=2.25
c264 57 0 1.62371e-19 $X=5.51 $Y=2.18
r265 74 76 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.21 $Y=2.185
+ $X2=7.21 $Y2=2.02
r266 74 75 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.21
+ $Y=2.185 $X2=7.21 $Y2=2.185
r267 70 84 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.53 $Y=1.285
+ $X2=6.53 $Y2=1.12
r268 69 72 8.60763 $w=3.88e-07 $l=1.65e-07 $layer=LI1_cond $X=6.5 $Y=1.285
+ $X2=6.5 $Y2=1.45
r269 69 71 8.60763 $w=3.88e-07 $l=1.65e-07 $layer=LI1_cond $X=6.5 $Y=1.285
+ $X2=6.5 $Y2=1.12
r270 69 70 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.53
+ $Y=1.285 $X2=6.53 $Y2=1.285
r271 64 76 104.059 $w=1.68e-07 $l=1.595e-06 $layer=LI1_cond $X=7.29 $Y=0.425
+ $X2=7.29 $Y2=2.02
r272 62 64 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.205 $Y=0.34
+ $X2=7.29 $Y2=0.425
r273 62 63 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=7.205 $Y=0.34
+ $X2=6.475 $Y2=0.34
r274 61 72 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=6.39 $Y=2.095
+ $X2=6.39 $Y2=1.45
r275 58 63 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.39 $Y=0.425
+ $X2=6.475 $Y2=0.34
r276 58 71 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=6.39 $Y=0.425
+ $X2=6.39 $Y2=1.12
r277 56 61 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.305 $Y=2.18
+ $X2=6.39 $Y2=2.095
r278 56 57 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=6.305 $Y=2.18
+ $X2=5.51 $Y2=2.18
r279 54 57 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.425 $Y=2.265
+ $X2=5.51 $Y2=2.18
r280 54 55 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=5.425 $Y=2.265
+ $X2=5.425 $Y2=2.905
r281 52 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.34 $Y=2.99
+ $X2=5.425 $Y2=2.905
r282 52 53 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=5.34 $Y=2.99
+ $X2=4.685 $Y2=2.99
r283 51 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.6 $Y=2.905
+ $X2=4.685 $Y2=2.99
r284 50 51 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=4.6 $Y=2.335
+ $X2=4.6 $Y2=2.905
r285 49 67 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.795 $Y=2.25
+ $X2=3.71 $Y2=2.25
r286 48 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.515 $Y=2.25
+ $X2=4.6 $Y2=2.335
r287 48 49 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=4.515 $Y=2.25
+ $X2=3.795 $Y2=2.25
r288 46 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.71 $Y=2.335
+ $X2=3.71 $Y2=2.25
r289 46 47 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=3.71 $Y=2.335
+ $X2=3.71 $Y2=2.905
r290 44 80 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=3.71 $Y=1.635
+ $X2=3.585 $Y2=1.635
r291 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.71
+ $Y=1.635 $X2=3.71 $Y2=1.635
r292 41 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.71 $Y=2.165
+ $X2=3.71 $Y2=2.25
r293 41 43 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.71 $Y=2.165
+ $X2=3.71 $Y2=1.635
r294 39 66 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=3.03 $Y=0.425
+ $X2=3.03 $Y2=1.455
r295 37 79 2.3474 $w=3.08e-07 $l=1.5e-08 $layer=POLY_cond $X=2.95 $Y=1.62
+ $X2=2.95 $Y2=1.635
r296 36 66 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.95 $Y=1.62
+ $X2=2.95 $Y2=1.455
r297 36 37 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.95
+ $Y=1.62 $X2=2.95 $Y2=1.62
r298 32 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.625 $Y=2.99
+ $X2=3.71 $Y2=2.905
r299 32 33 88.0749 $w=1.68e-07 $l=1.35e-06 $layer=LI1_cond $X=3.625 $Y=2.99
+ $X2=2.275 $Y2=2.99
r300 30 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.945 $Y=0.34
+ $X2=3.03 $Y2=0.425
r301 30 31 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=2.945 $Y=0.34
+ $X2=2.215 $Y2=0.34
r302 26 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.19 $Y=2.905
+ $X2=2.275 $Y2=2.99
r303 26 28 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.19 $Y=2.905
+ $X2=2.19 $Y2=2.575
r304 22 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.13 $Y=0.425
+ $X2=2.215 $Y2=0.34
r305 22 24 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=2.13 $Y=0.425
+ $X2=2.13 $Y2=0.515
r306 19 75 55.8714 $w=3.2e-07 $l=3.24037e-07 $layer=POLY_cond $X=7.325 $Y=2.465
+ $X2=7.23 $Y2=2.185
r307 19 21 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.325 $Y=2.465
+ $X2=7.325 $Y2=2.75
r308 18 84 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=6.595 $Y=0.69
+ $X2=6.595 $Y2=1.12
r309 12 80 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.585 $Y=1.47
+ $X2=3.585 $Y2=1.635
r310 12 14 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=3.585 $Y=1.47
+ $X2=3.585 $Y2=0.58
r311 11 79 1.15097 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.115 $Y=1.635
+ $X2=2.95 $Y2=1.635
r312 10 80 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=3.51 $Y=1.635
+ $X2=3.585 $Y2=1.635
r313 10 11 69.0702 $w=3.3e-07 $l=3.95e-07 $layer=POLY_cond $X=3.51 $Y=1.635
+ $X2=3.115 $Y2=1.635
r314 7 79 107.39 $w=3.08e-07 $l=6.31902e-07 $layer=POLY_cond $X=3.005 $Y=2.24
+ $X2=2.95 $Y2=1.635
r315 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.005 $Y=2.24
+ $X2=3.005 $Y2=2.525
r316 2 28 600 $w=1.7e-07 $l=8.0652e-07 $layer=licon1_PDIFF $count=1 $X=2.04
+ $Y=1.84 $X2=2.19 $Y2=2.575
r317 1 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.99
+ $Y=0.37 $X2=2.13 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__DFSTP_4%A_767_402# 1 2 7 9 10 12 13 14 16 17 23 25
+ 32 35
c86 35 0 1.30099e-19 $X=4.395 $Y=0.975
c87 17 0 1.30611e-19 $X=4.855 $Y=1.867
c88 7 0 1.18613e-19 $X=3.925 $Y=2.24
r89 29 32 3.79782 $w=4.38e-07 $l=1.45e-07 $layer=LI1_cond $X=4.94 $Y=2.515
+ $X2=5.085 $Y2=2.515
r90 26 38 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.395 $Y=1.065
+ $X2=4.395 $Y2=1.23
r91 26 35 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.395 $Y=1.065
+ $X2=4.395 $Y2=0.975
r92 25 28 14.8027 $w=3.75e-07 $l=4.55e-07 $layer=LI1_cond $X=4.395 $Y=0.925
+ $X2=4.85 $Y2=0.925
r93 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.395
+ $Y=1.065 $X2=4.395 $Y2=1.065
r94 23 29 6.36164 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=4.94 $Y=2.295
+ $X2=4.94 $Y2=2.515
r95 22 23 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=4.94 $Y=1.995 $X2=4.94
+ $Y2=2.295
r96 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.28
+ $Y=1.865 $X2=4.28 $Y2=1.865
r97 17 22 7.17723 $w=2.55e-07 $l=1.65118e-07 $layer=LI1_cond $X=4.855 $Y=1.867
+ $X2=4.94 $Y2=1.995
r98 17 19 25.9865 $w=2.53e-07 $l=5.75e-07 $layer=LI1_cond $X=4.855 $Y=1.867
+ $X2=4.28 $Y2=1.867
r99 16 20 39.305 $w=3.85e-07 $l=2.33345e-07 $layer=POLY_cond $X=4.305 $Y=1.7
+ $X2=4.14 $Y2=1.865
r100 16 38 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=4.305 $Y=1.7 $X2=4.305
+ $Y2=1.23
r101 13 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.23 $Y=0.975
+ $X2=4.395 $Y2=0.975
r102 13 14 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=4.23 $Y=0.975
+ $X2=4.05 $Y2=0.975
r103 10 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.975 $Y=0.9
+ $X2=4.05 $Y2=0.975
r104 10 12 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.975 $Y=0.9
+ $X2=3.975 $Y2=0.58
r105 7 20 65.5959 $w=3.85e-07 $l=4.70372e-07 $layer=POLY_cond $X=3.925 $Y=2.24
+ $X2=4.14 $Y2=1.865
r106 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.925 $Y=2.24
+ $X2=3.925 $Y2=2.525
r107 2 32 600 $w=1.7e-07 $l=2.64575e-07 $layer=licon1_PDIFF $count=1 $X=4.935
+ $Y=2.315 $X2=5.085 $Y2=2.515
r108 1 28 182 $w=1.7e-07 $l=2.70416e-07 $layer=licon1_NDIFF $count=1 $X=4.67
+ $Y=0.59 $X2=4.85 $Y2=0.785
.ends

.subckt PM_SKY130_FD_SC_LS__DFSTP_4%A_612_74# 1 2 8 9 11 12 14 15 17 20 24 28 30
+ 32 35 36 38 39 44 49 58
c137 44 0 2.27104e-19 $X=4.935 $Y=1.285
c138 35 0 1.18613e-19 $X=3.28 $Y=2.515
c139 9 0 2.33614e-20 $X=4.86 $Y=2.24
c140 8 0 1.3901e-19 $X=4.86 $Y=2.15
r141 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.97
+ $Y=1.365 $X2=5.97 $Y2=1.365
r142 49 52 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=5.97 $Y=1.285 $X2=5.97
+ $Y2=1.365
r143 45 58 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.935 $Y=1.285
+ $X2=5.1 $Y2=1.285
r144 45 55 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.935 $Y=1.285
+ $X2=4.86 $Y2=1.285
r145 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.935
+ $Y=1.285 $X2=4.935 $Y2=1.285
r146 39 41 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=4.05 $Y=1.215
+ $X2=4.05 $Y2=1.485
r147 35 36 10.3362 $w=3.38e-07 $l=2.2e-07 $layer=LI1_cond $X=3.285 $Y=2.515
+ $X2=3.285 $Y2=2.295
r148 33 44 3.11056 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=5.025 $Y=1.285
+ $X2=4.897 $Y2=1.285
r149 32 49 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.805 $Y=1.285
+ $X2=5.97 $Y2=1.285
r150 32 33 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=5.805 $Y=1.285
+ $X2=5.025 $Y2=1.285
r151 31 41 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.135 $Y=1.485
+ $X2=4.05 $Y2=1.485
r152 30 44 9.03877 $w=2.53e-07 $l=2e-07 $layer=LI1_cond $X=4.897 $Y=1.485
+ $X2=4.897 $Y2=1.285
r153 30 31 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=4.77 $Y=1.485
+ $X2=4.135 $Y2=1.485
r154 29 38 2.11342 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.535 $Y=1.215
+ $X2=3.41 $Y2=1.215
r155 28 39 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.965 $Y=1.215
+ $X2=4.05 $Y2=1.215
r156 28 29 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=3.965 $Y=1.215
+ $X2=3.535 $Y2=1.215
r157 26 38 4.3182 $w=2.1e-07 $l=1.03078e-07 $layer=LI1_cond $X=3.37 $Y=1.3
+ $X2=3.41 $Y2=1.215
r158 26 36 64.9144 $w=1.68e-07 $l=9.95e-07 $layer=LI1_cond $X=3.37 $Y=1.3
+ $X2=3.37 $Y2=2.295
r159 22 38 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.41 $Y=1.13 $X2=3.41
+ $Y2=1.215
r160 22 24 25.3537 $w=2.48e-07 $l=5.5e-07 $layer=LI1_cond $X=3.41 $Y=1.13
+ $X2=3.41 $Y2=0.58
r161 18 53 38.6443 $w=2.87e-07 $l=2.0106e-07 $layer=POLY_cond $X=6.05 $Y=1.2
+ $X2=5.97 $Y2=1.365
r162 18 20 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=6.05 $Y=1.2
+ $X2=6.05 $Y2=0.69
r163 15 53 60.4771 $w=2.87e-07 $l=3.21325e-07 $layer=POLY_cond $X=6.025 $Y=1.66
+ $X2=5.97 $Y2=1.365
r164 15 17 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.025 $Y=1.66
+ $X2=6.025 $Y2=2.235
r165 12 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.1 $Y=1.12
+ $X2=5.1 $Y2=1.285
r166 12 14 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=5.1 $Y=1.12 $X2=5.1
+ $Y2=0.8
r167 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.86 $Y=2.24 $X2=4.86
+ $Y2=2.525
r168 8 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=4.86 $Y=2.15 $X2=4.86
+ $Y2=2.24
r169 7 55 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.86 $Y=1.45
+ $X2=4.86 $Y2=1.285
r170 7 8 272.097 $w=1.8e-07 $l=7e-07 $layer=POLY_cond $X=4.86 $Y=1.45 $X2=4.86
+ $Y2=2.15
r171 2 35 600 $w=1.7e-07 $l=2.82843e-07 $layer=licon1_PDIFF $count=1 $X=3.08
+ $Y=2.315 $X2=3.28 $Y2=2.515
r172 1 24 182 $w=1.7e-07 $l=4.01497e-07 $layer=licon1_NDIFF $count=1 $X=3.06
+ $Y=0.37 $X2=3.37 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_LS__DFSTP_4%SET_B 2 3 5 8 10 12 13 14 16 17 19 20 21 22
+ 27 33 34 39
c137 39 0 1.13172e-19 $X=8.35 $Y=1.345
c138 22 0 9.70053e-20 $X=5.665 $Y=1.665
c139 21 0 2.34318e-20 $X=8.255 $Y=1.665
c140 16 0 6.99491e-20 $X=8.195 $Y=2.375
c141 2 0 1.30611e-19 $X=5.31 $Y=2.15
r142 39 46 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=8.35 $Y=1.345
+ $X2=8.35 $Y2=1.665
r143 32 34 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=5.36 $Y=1.825
+ $X2=5.49 $Y2=1.825
r144 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.36
+ $Y=1.825 $X2=5.36 $Y2=1.825
r145 29 32 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=5.31 $Y=1.825
+ $X2=5.36 $Y2=1.825
r146 27 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=1.665
+ $X2=8.4 $Y2=1.665
r147 24 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=1.665
+ $X2=5.52 $Y2=1.665
r148 22 24 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.665 $Y=1.665
+ $X2=5.52 $Y2=1.665
r149 21 27 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.255 $Y=1.665
+ $X2=8.4 $Y2=1.665
r150 21 22 3.20544 $w=1.4e-07 $l=2.59e-06 $layer=MET1_cond $X=8.255 $Y=1.665
+ $X2=5.665 $Y2=1.665
r151 17 19 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=8.195 $Y=2.465
+ $X2=8.195 $Y2=2.75
r152 16 17 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=8.195 $Y=2.375
+ $X2=8.195 $Y2=2.465
r153 16 20 204.073 $w=1.8e-07 $l=5.25e-07 $layer=POLY_cond $X=8.195 $Y=2.375
+ $X2=8.195 $Y2=1.85
r154 14 20 45.5979 $w=4.1e-07 $l=2.05e-07 $layer=POLY_cond $X=8.31 $Y=1.645
+ $X2=8.31 $Y2=1.85
r155 13 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.35
+ $Y=1.345 $X2=8.35 $Y2=1.345
r156 13 14 35.2683 $w=4.1e-07 $l=2.6e-07 $layer=POLY_cond $X=8.31 $Y=1.385
+ $X2=8.31 $Y2=1.645
r157 10 13 86.4346 $w=2.37e-07 $l=6.27495e-07 $layer=POLY_cond $X=7.885 $Y=0.935
+ $X2=8.31 $Y2=1.385
r158 10 12 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.885 $Y=0.935
+ $X2=7.885 $Y2=0.65
r159 6 34 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.49 $Y=1.66
+ $X2=5.49 $Y2=1.825
r160 6 8 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=5.49 $Y=1.66 $X2=5.49
+ $Y2=0.8
r161 3 5 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=5.31 $Y=2.24 $X2=5.31
+ $Y2=2.525
r162 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.31 $Y=2.15 $X2=5.31
+ $Y2=2.24
r163 1 29 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.31 $Y=1.99
+ $X2=5.31 $Y2=1.825
r164 1 2 62.1936 $w=1.8e-07 $l=1.6e-07 $layer=POLY_cond $X=5.31 $Y=1.99 $X2=5.31
+ $Y2=2.15
.ends

.subckt PM_SKY130_FD_SC_LS__DFSTP_4%A_225_74# 1 2 9 11 13 15 16 18 19 22 24 25
+ 26 28 29 34 35 36 39 43 46 47 49 50 54 58 65
c179 35 0 2.80241e-20 $X=7.03 $Y=1.735
c180 26 0 1.22525e-19 $X=3.505 $Y=2.81
r181 64 65 8.48848 $w=3.48e-07 $l=1.65e-07 $layer=LI1_cond $X=1.29 $Y=1.895
+ $X2=1.455 $Y2=1.895
r182 61 64 7.5732 $w=3.48e-07 $l=2.3e-07 $layer=LI1_cond $X=1.06 $Y=1.895
+ $X2=1.29 $Y2=1.895
r183 58 60 17.8607 $w=4.58e-07 $l=4.95e-07 $layer=LI1_cond $X=1.205 $Y=0.515
+ $X2=1.205 $Y2=1.01
r184 54 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.11
+ $Y=1.515 $X2=2.11 $Y2=1.515
r185 52 54 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=2.11 $Y=1.72
+ $X2=2.11 $Y2=1.515
r186 50 52 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.945 $Y=1.805
+ $X2=2.11 $Y2=1.72
r187 50 65 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=1.945 $Y=1.805
+ $X2=1.455 $Y2=1.805
r188 49 61 4.974 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=1.06 $Y=1.72 $X2=1.06
+ $Y2=1.895
r189 49 60 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=1.06 $Y=1.72
+ $X2=1.06 $Y2=1.01
r190 46 55 52.4584 $w=3.3e-07 $l=3e-07 $layer=POLY_cond $X=2.41 $Y=1.515
+ $X2=2.11 $Y2=1.515
r191 43 46 192.287 $w=1.5e-07 $l=3.75e-07 $layer=POLY_cond $X=2.485 $Y=1.14
+ $X2=2.485 $Y2=1.515
r192 42 55 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=2.055 $Y=1.515
+ $X2=2.11 $Y2=1.515
r193 37 39 517.894 $w=1.5e-07 $l=1.01e-06 $layer=POLY_cond $X=7.105 $Y=1.66
+ $X2=7.105 $Y2=0.65
r194 35 37 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.03 $Y=1.735
+ $X2=7.105 $Y2=1.66
r195 35 36 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=7.03 $Y=1.735
+ $X2=6.62 $Y2=1.735
r196 32 34 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.53 $Y=3.035
+ $X2=6.53 $Y2=2.46
r197 31 36 26.9307 $w=1.5e-07 $l=1.89737e-07 $layer=POLY_cond $X=6.53 $Y=1.885
+ $X2=6.62 $Y2=1.735
r198 31 34 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.53 $Y=1.885
+ $X2=6.53 $Y2=2.46
r199 30 47 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.595 $Y=3.15
+ $X2=3.505 $Y2=3.15
r200 29 32 26.9307 $w=1.5e-07 $l=1.53542e-07 $layer=POLY_cond $X=6.44 $Y=3.15
+ $X2=6.53 $Y2=3.035
r201 29 30 1458.82 $w=1.5e-07 $l=2.845e-06 $layer=POLY_cond $X=6.44 $Y=3.15
+ $X2=3.595 $Y2=3.15
r202 26 28 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.505 $Y=2.81
+ $X2=3.505 $Y2=2.525
r203 25 47 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=3.505 $Y=3.075
+ $X2=3.505 $Y2=3.15
r204 24 26 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.505 $Y=2.9
+ $X2=3.505 $Y2=2.81
r205 24 25 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=3.505 $Y=2.9
+ $X2=3.505 $Y2=3.075
r206 20 22 248.691 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=2.985 $Y=1.065
+ $X2=2.985 $Y2=0.58
r207 18 47 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.415 $Y=3.15
+ $X2=3.505 $Y2=3.15
r208 18 19 438.415 $w=1.5e-07 $l=8.55e-07 $layer=POLY_cond $X=3.415 $Y=3.15
+ $X2=2.56 $Y2=3.15
r209 17 43 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.56 $Y=1.14
+ $X2=2.485 $Y2=1.14
r210 16 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.91 $Y=1.14
+ $X2=2.985 $Y2=1.065
r211 16 17 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=2.91 $Y=1.14
+ $X2=2.56 $Y2=1.14
r212 15 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.485 $Y=3.075
+ $X2=2.56 $Y2=3.15
r213 14 46 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.485 $Y=1.68
+ $X2=2.485 $Y2=1.515
r214 14 15 715.309 $w=1.5e-07 $l=1.395e-06 $layer=POLY_cond $X=2.485 $Y=1.68
+ $X2=2.485 $Y2=3.075
r215 11 42 61.9504 $w=2.07e-07 $l=2.58844e-07 $layer=POLY_cond $X=1.965 $Y=1.765
+ $X2=1.947 $Y2=1.515
r216 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.965 $Y=1.765
+ $X2=1.965 $Y2=2.4
r217 7 42 42.1581 $w=2.07e-07 $l=1.80291e-07 $layer=POLY_cond $X=1.915 $Y=1.35
+ $X2=1.947 $Y2=1.515
r218 7 9 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.915 $Y=1.35
+ $X2=1.915 $Y2=0.74
r219 2 64 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.145
+ $Y=1.84 $X2=1.29 $Y2=1.985
r220 1 58 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=1.125
+ $Y=0.37 $X2=1.27 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__DFSTP_4%A_1484_62# 1 2 9 12 13 15 18 21 22 25 29 31
+ 32 37
c90 37 0 1.90022e-19 $X=7.745 $Y=1.49
c91 12 0 7.64129e-20 $X=7.745 $Y=2.375
c92 9 0 1.13172e-19 $X=7.495 $Y=0.65
r93 31 32 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=9.395 $Y=2.815
+ $X2=9.395 $Y2=2.65
r94 27 29 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=9.365 $Y=1.01
+ $X2=9.285 $Y2=0.925
r95 27 32 106.995 $w=1.68e-07 $l=1.64e-06 $layer=LI1_cond $X=9.365 $Y=1.01
+ $X2=9.365 $Y2=2.65
r96 23 29 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.285 $Y=0.84
+ $X2=9.285 $Y2=0.925
r97 23 25 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=9.285 $Y=0.84
+ $X2=9.285 $Y2=0.65
r98 21 29 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.12 $Y=0.925
+ $X2=9.285 $Y2=0.925
r99 21 22 81.2246 $w=1.68e-07 $l=1.245e-06 $layer=LI1_cond $X=9.12 $Y=0.925
+ $X2=7.875 $Y2=0.925
r100 19 37 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=7.71 $Y=1.49
+ $X2=7.745 $Y2=1.49
r101 19 34 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=7.71 $Y=1.49
+ $X2=7.495 $Y2=1.49
r102 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.71
+ $Y=1.49 $X2=7.71 $Y2=1.49
r103 16 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.71 $Y=1.01
+ $X2=7.875 $Y2=0.925
r104 16 18 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=7.71 $Y=1.01
+ $X2=7.71 $Y2=1.49
r105 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.745 $Y=2.465
+ $X2=7.745 $Y2=2.75
r106 12 13 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=7.745 $Y=2.375
+ $X2=7.745 $Y2=2.465
r107 11 37 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.745 $Y=1.655
+ $X2=7.745 $Y2=1.49
r108 11 12 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=7.745 $Y=1.655
+ $X2=7.745 $Y2=2.375
r109 7 34 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.495 $Y=1.325
+ $X2=7.495 $Y2=1.49
r110 7 9 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=7.495 $Y=1.325
+ $X2=7.495 $Y2=0.65
r111 2 31 600 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=9.245
+ $Y=2.54 $X2=9.395 $Y2=2.815
r112 1 25 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=9.145
+ $Y=0.44 $X2=9.285 $Y2=0.65
.ends

.subckt PM_SKY130_FD_SC_LS__DFSTP_4%A_1321_392# 1 2 3 11 14 16 18 19 23 25 27 28
+ 30 32 38 40 41 42 43 47 49 53 54 65 69 71 75
c166 71 0 6.99491e-20 $X=7.63 $Y=2.395
c167 69 0 5.89928e-20 $X=6.95 $Y=1.705
c168 43 0 1.90022e-19 $X=8.255 $Y=2.395
c169 28 0 2.87198e-21 $X=10.52 $Y=1.69
c170 23 0 2.91921e-19 $X=10.13 $Y=0.74
r171 71 73 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=7.63 $Y=2.395
+ $X2=7.63 $Y2=2.565
r172 67 69 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=6.755 $Y=1.705
+ $X2=6.95 $Y2=1.705
r173 63 65 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=6.81 $Y=0.76
+ $X2=6.95 $Y2=0.76
r174 59 61 8.78706 $w=4.79e-07 $l=3.45e-07 $layer=LI1_cond $X=6.755 $Y=2.73
+ $X2=7.1 $Y2=2.73
r175 57 58 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=8.945
+ $Y=2.215 $X2=8.945 $Y2=2.215
r176 53 57 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=8.945 $Y=1.535
+ $X2=8.945 $Y2=2.215
r177 53 54 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=8.945
+ $Y=1.535 $X2=8.945 $Y2=1.535
r178 51 57 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=8.945 $Y=2.31
+ $X2=8.945 $Y2=2.215
r179 50 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.585 $Y=2.395
+ $X2=8.42 $Y2=2.395
r180 49 51 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.78 $Y=2.395
+ $X2=8.945 $Y2=2.31
r181 49 50 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=8.78 $Y=2.395
+ $X2=8.585 $Y2=2.395
r182 45 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.42 $Y=2.48
+ $X2=8.42 $Y2=2.395
r183 45 47 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=8.42 $Y=2.48
+ $X2=8.42 $Y2=2.75
r184 44 71 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.715 $Y=2.395
+ $X2=7.63 $Y2=2.395
r185 43 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.255 $Y=2.395
+ $X2=8.42 $Y2=2.395
r186 43 44 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=8.255 $Y=2.395
+ $X2=7.715 $Y2=2.395
r187 42 61 9.57821 $w=4.79e-07 $l=2.33345e-07 $layer=LI1_cond $X=7.265 $Y=2.565
+ $X2=7.1 $Y2=2.73
r188 41 73 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.545 $Y=2.565
+ $X2=7.63 $Y2=2.565
r189 41 42 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=7.545 $Y=2.565
+ $X2=7.265 $Y2=2.565
r190 40 69 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.95 $Y=1.62
+ $X2=6.95 $Y2=1.705
r191 39 65 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.95 $Y=0.925
+ $X2=6.95 $Y2=0.76
r192 39 40 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=6.95 $Y=0.925
+ $X2=6.95 $Y2=1.62
r193 36 59 6.88815 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=6.755 $Y=2.48
+ $X2=6.755 $Y2=2.73
r194 36 38 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=6.755 $Y=2.48
+ $X2=6.755 $Y2=2.135
r195 35 67 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.755 $Y=1.79
+ $X2=6.755 $Y2=1.705
r196 35 38 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=6.755 $Y=1.79
+ $X2=6.755 $Y2=2.135
r197 30 32 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=10.595 $Y=1.765
+ $X2=10.595 $Y2=2.26
r198 29 34 3.61756 $w=1.5e-07 $l=8.3e-08 $layer=POLY_cond $X=10.22 $Y=1.69
+ $X2=10.137 $Y2=1.69
r199 28 30 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.52 $Y=1.69
+ $X2=10.595 $Y2=1.765
r200 28 29 153.83 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=10.52 $Y=1.69
+ $X2=10.22 $Y2=1.69
r201 25 34 23.3226 $w=1.55e-07 $l=7.88987e-08 $layer=POLY_cond $X=10.145
+ $Y=1.765 $X2=10.137 $Y2=1.69
r202 25 27 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=10.145 $Y=1.765
+ $X2=10.145 $Y2=2.26
r203 21 23 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=10.13 $Y=1.37
+ $X2=10.13 $Y2=0.74
r204 20 54 8.93404 $w=2.45e-07 $l=2.4e-07 $layer=POLY_cond $X=9.26 $Y=1.492
+ $X2=9.02 $Y2=1.492
r205 19 34 61.5716 $w=1.55e-07 $l=1.98e-07 $layer=POLY_cond $X=10.137 $Y=1.492
+ $X2=10.137 $Y2=1.69
r206 19 21 37.9381 $w=1.55e-07 $l=1.25451e-07 $layer=POLY_cond $X=10.137
+ $Y=1.492 $X2=10.13 $Y2=1.37
r207 19 20 201.552 $w=2.45e-07 $l=7.95e-07 $layer=POLY_cond $X=10.055 $Y=1.492
+ $X2=9.26 $Y2=1.492
r208 16 58 49.8219 $w=4.01e-07 $l=3.16228e-07 $layer=POLY_cond $X=9.17 $Y=2.465
+ $X2=9.02 $Y2=2.215
r209 16 18 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=9.17 $Y=2.465
+ $X2=9.17 $Y2=2.75
r210 12 54 16.4793 $w=3.15e-07 $l=1.44859e-07 $layer=POLY_cond $X=9.07 $Y=1.37
+ $X2=9.02 $Y2=1.492
r211 12 14 369.191 $w=1.5e-07 $l=7.2e-07 $layer=POLY_cond $X=9.07 $Y=1.37
+ $X2=9.07 $Y2=0.65
r212 11 58 8.97868 $w=4.8e-07 $l=7.5e-08 $layer=POLY_cond $X=9.02 $Y=2.14
+ $X2=9.02 $Y2=2.215
r213 10 54 16.4793 $w=3.15e-07 $l=1.23e-07 $layer=POLY_cond $X=9.02 $Y=1.615
+ $X2=9.02 $Y2=1.492
r214 10 11 58.5188 $w=4.8e-07 $l=5.25e-07 $layer=POLY_cond $X=9.02 $Y=1.615
+ $X2=9.02 $Y2=2.14
r215 3 47 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=8.27
+ $Y=2.54 $X2=8.42 $Y2=2.75
r216 2 61 300 $w=1.7e-07 $l=1.07436e-06 $layer=licon1_PDIFF $count=2 $X=6.605
+ $Y=1.96 $X2=7.1 $Y2=2.815
r217 2 38 300 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=2 $X=6.605
+ $Y=1.96 $X2=6.755 $Y2=2.135
r218 1 63 182 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_NDIFF $count=1 $X=6.67
+ $Y=0.37 $X2=6.81 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_LS__DFSTP_4%A_1940_74# 1 2 7 9 10 11 12 14 15 17 18 20
+ 21 23 24 26 27 29 31 33 36 38 39 42 49 52
r114 58 59 10.5507 $w=4.34e-07 $l=9.5e-08 $layer=POLY_cond $X=11.92 $Y=1.495
+ $X2=12.015 $Y2=1.495
r115 53 54 6.10829 $w=4.34e-07 $l=5.5e-08 $layer=POLY_cond $X=11.06 $Y=1.495
+ $X2=11.115 $Y2=1.495
r116 50 58 9.99539 $w=4.34e-07 $l=9e-08 $layer=POLY_cond $X=11.83 $Y=1.495
+ $X2=11.92 $Y2=1.495
r117 50 56 29.4309 $w=4.34e-07 $l=2.65e-07 $layer=POLY_cond $X=11.83 $Y=1.495
+ $X2=11.565 $Y2=1.495
r118 49 50 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=11.83
+ $Y=1.485 $X2=11.83 $Y2=1.485
r119 47 56 46.0899 $w=4.34e-07 $l=4.15e-07 $layer=POLY_cond $X=11.15 $Y=1.495
+ $X2=11.565 $Y2=1.495
r120 47 54 3.8871 $w=4.34e-07 $l=3.5e-08 $layer=POLY_cond $X=11.15 $Y=1.495
+ $X2=11.115 $Y2=1.495
r121 46 49 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=11.15 $Y=1.485
+ $X2=11.83 $Y2=1.485
r122 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.15
+ $Y=1.485 $X2=11.15 $Y2=1.485
r123 44 52 6.46576 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=10.535 $Y=1.485
+ $X2=10.37 $Y2=1.485
r124 44 46 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=10.535 $Y=1.485
+ $X2=11.15 $Y2=1.485
r125 40 52 0.364692 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=10.37 $Y=1.65
+ $X2=10.37 $Y2=1.485
r126 40 42 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=10.37 $Y=1.65
+ $X2=10.37 $Y2=1.985
r127 38 52 6.46576 $w=2.5e-07 $l=2.0106e-07 $layer=LI1_cond $X=10.205 $Y=1.405
+ $X2=10.37 $Y2=1.485
r128 38 39 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=10.205 $Y=1.405
+ $X2=10.01 $Y2=1.405
r129 34 39 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.845 $Y=1.32
+ $X2=10.01 $Y2=1.405
r130 34 36 28.1126 $w=3.28e-07 $l=8.05e-07 $layer=LI1_cond $X=9.845 $Y=1.32
+ $X2=9.845 $Y2=0.515
r131 31 61 27.8684 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=12.465 $Y=1.765
+ $X2=12.465 $Y2=1.495
r132 31 33 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=12.465 $Y=1.765
+ $X2=12.465 $Y2=2.4
r133 27 61 7.77419 $w=4.34e-07 $l=7e-08 $layer=POLY_cond $X=12.395 $Y=1.495
+ $X2=12.465 $Y2=1.495
r134 27 59 42.2028 $w=4.34e-07 $l=3.8e-07 $layer=POLY_cond $X=12.395 $Y=1.495
+ $X2=12.015 $Y2=1.495
r135 27 29 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=12.395 $Y=1.32
+ $X2=12.395 $Y2=0.74
r136 24 59 27.8684 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=12.015 $Y=1.765
+ $X2=12.015 $Y2=1.495
r137 24 26 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=12.015 $Y=1.765
+ $X2=12.015 $Y2=2.4
r138 21 58 27.8684 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=11.92 $Y=1.225
+ $X2=11.92 $Y2=1.495
r139 21 23 155.847 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=11.92 $Y=1.225
+ $X2=11.92 $Y2=0.74
r140 18 56 27.8684 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=11.565 $Y=1.765
+ $X2=11.565 $Y2=1.495
r141 18 20 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=11.565 $Y=1.765
+ $X2=11.565 $Y2=2.4
r142 15 54 27.8684 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=11.115 $Y=1.765
+ $X2=11.115 $Y2=1.495
r143 15 17 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=11.115 $Y=1.765
+ $X2=11.115 $Y2=2.4
r144 12 53 27.8684 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=11.06 $Y=1.225
+ $X2=11.06 $Y2=1.495
r145 12 14 155.847 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=11.06 $Y=1.225
+ $X2=11.06 $Y2=0.74
r146 10 53 30.3131 $w=4.34e-07 $l=2.29456e-07 $layer=POLY_cond $X=10.985 $Y=1.3
+ $X2=11.06 $Y2=1.495
r147 10 11 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=10.985 $Y=1.3
+ $X2=10.705 $Y2=1.3
r148 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.63 $Y=1.225
+ $X2=10.705 $Y2=1.3
r149 7 9 155.847 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=10.63 $Y=1.225
+ $X2=10.63 $Y2=0.74
r150 2 42 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=10.22
+ $Y=1.84 $X2=10.37 $Y2=1.985
r151 1 36 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=9.7
+ $Y=0.37 $X2=9.845 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__DFSTP_4%A_27_74# 1 2 3 4 15 18 21 23 25 28 29 30 31
+ 38
c69 25 0 1.22525e-19 $X=2.445 $Y=2.155
r70 35 38 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=2.53 $Y=0.76 $X2=2.69
+ $Y2=0.76
r71 31 33 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.71 $Y=2.155
+ $X2=1.71 $Y2=2.325
r72 27 35 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.53 $Y=0.925
+ $X2=2.53 $Y2=0.76
r73 27 28 74.7005 $w=1.68e-07 $l=1.145e-06 $layer=LI1_cond $X=2.53 $Y=0.925
+ $X2=2.53 $Y2=2.07
r74 26 31 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.795 $Y=2.155
+ $X2=1.71 $Y2=2.155
r75 25 42 11.3196 $w=3.88e-07 $l=4.68615e-07 $layer=LI1_cond $X=2.445 $Y=2.155
+ $X2=2.695 $Y2=2.515
r76 25 28 6.58872 $w=3.88e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.445 $Y=2.155
+ $X2=2.53 $Y2=2.07
r77 25 26 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=2.445 $Y=2.155
+ $X2=1.795 $Y2=2.155
r78 24 30 2.11342 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.365 $Y=2.325
+ $X2=0.24 $Y2=2.325
r79 23 33 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.625 $Y=2.325
+ $X2=1.71 $Y2=2.325
r80 23 24 82.2032 $w=1.68e-07 $l=1.26e-06 $layer=LI1_cond $X=1.625 $Y=2.325
+ $X2=0.365 $Y2=2.325
r81 19 30 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.24 $Y=2.41 $X2=0.24
+ $Y2=2.325
r82 19 21 14.7513 $w=2.48e-07 $l=3.2e-07 $layer=LI1_cond $X=0.24 $Y=2.41
+ $X2=0.24 $Y2=2.73
r83 18 30 4.3182 $w=2.1e-07 $l=1.03078e-07 $layer=LI1_cond $X=0.2 $Y=2.24
+ $X2=0.24 $Y2=2.325
r84 18 29 93.2941 $w=1.68e-07 $l=1.43e-06 $layer=LI1_cond $X=0.2 $Y=2.24 $X2=0.2
+ $Y2=0.81
r85 13 29 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=0.24 $Y=0.685
+ $X2=0.24 $Y2=0.81
r86 13 15 4.84026 $w=2.48e-07 $l=1.05e-07 $layer=LI1_cond $X=0.24 $Y=0.685
+ $X2=0.24 $Y2=0.58
r87 4 42 600 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=1 $X=2.635
+ $Y=2.315 $X2=2.78 $Y2=2.515
r88 3 21 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.52 $X2=0.28 $Y2=2.73
r89 2 38 182 $w=1.7e-07 $l=4.56782e-07 $layer=licon1_NDIFF $count=1 $X=2.545
+ $Y=0.37 $X2=2.69 $Y2=0.76
r90 1 15 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_LS__DFSTP_4%VPWR 1 2 3 4 5 6 7 8 9 10 33 37 40 43 47 51
+ 55 57 61 67 69 71 76 79 80 81 83 88 93 105 109 114 119 124 130 133 136 139 142
+ 145 148 151 155
r175 154 155 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r176 151 152 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r177 148 149 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r178 146 149 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=10.8 $Y2=3.33
r179 145 146 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r180 142 143 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r181 139 140 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r182 136 137 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r183 133 134 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r184 130 131 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r185 128 155 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=12.72 $Y2=3.33
r186 128 152 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=11.76 $Y2=3.33
r187 127 128 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r188 125 151 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.955 $Y=3.33
+ $X2=11.79 $Y2=3.33
r189 125 127 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=11.955 $Y=3.33
+ $X2=12.24 $Y2=3.33
r190 124 154 4.76062 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=12.525 $Y=3.33
+ $X2=12.742 $Y2=3.33
r191 124 127 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=12.525 $Y=3.33
+ $X2=12.24 $Y2=3.33
r192 123 152 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=11.76 $Y2=3.33
r193 123 149 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=10.8 $Y2=3.33
r194 122 123 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r195 120 148 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=11.005 $Y=3.33
+ $X2=10.865 $Y2=3.33
r196 120 122 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=11.005 $Y=3.33
+ $X2=11.28 $Y2=3.33
r197 119 151 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.625 $Y=3.33
+ $X2=11.79 $Y2=3.33
r198 119 122 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=11.625 $Y=3.33
+ $X2=11.28 $Y2=3.33
r199 118 146 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=9.84 $Y2=3.33
r200 118 143 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=8.88 $Y2=3.33
r201 117 118 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r202 115 142 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.03 $Y=3.33
+ $X2=8.905 $Y2=3.33
r203 115 117 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=9.03 $Y=3.33
+ $X2=9.36 $Y2=3.33
r204 114 145 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.755 $Y=3.33
+ $X2=9.88 $Y2=3.33
r205 114 117 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=9.755 $Y=3.33
+ $X2=9.36 $Y2=3.33
r206 113 143 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=8.88 $Y2=3.33
r207 113 140 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=7.92 $Y2=3.33
r208 112 113 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r209 110 139 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.055 $Y=3.33
+ $X2=7.97 $Y2=3.33
r210 110 112 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=8.055 $Y=3.33
+ $X2=8.4 $Y2=3.33
r211 109 142 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.78 $Y=3.33
+ $X2=8.905 $Y2=3.33
r212 109 112 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=8.78 $Y=3.33
+ $X2=8.4 $Y2=3.33
r213 107 108 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r214 105 139 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.885 $Y=3.33
+ $X2=7.97 $Y2=3.33
r215 105 107 122.979 $w=1.68e-07 $l=1.885e-06 $layer=LI1_cond $X=7.885 $Y=3.33
+ $X2=6 $Y2=3.33
r216 104 108 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6 $Y2=3.33
r217 104 137 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=4.08 $Y2=3.33
r218 103 104 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r219 101 136 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.155 $Y=3.33
+ $X2=4.07 $Y2=3.33
r220 101 103 89.0535 $w=1.68e-07 $l=1.365e-06 $layer=LI1_cond $X=4.155 $Y=3.33
+ $X2=5.52 $Y2=3.33
r221 100 137 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r222 99 100 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r223 97 100 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.6 $Y2=3.33
r224 97 134 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r225 96 99 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=3.6 $Y2=3.33
r226 96 97 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r227 94 133 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.905 $Y=3.33
+ $X2=1.74 $Y2=3.33
r228 94 96 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.905 $Y=3.33
+ $X2=2.16 $Y2=3.33
r229 93 136 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.985 $Y=3.33
+ $X2=4.07 $Y2=3.33
r230 93 99 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=3.985 $Y=3.33
+ $X2=3.6 $Y2=3.33
r231 92 134 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r232 92 131 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r233 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r234 89 130 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=0.73 $Y2=3.33
r235 89 91 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=1.2 $Y2=3.33
r236 88 133 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.575 $Y=3.33
+ $X2=1.74 $Y2=3.33
r237 88 91 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.575 $Y=3.33
+ $X2=1.2 $Y2=3.33
r238 86 131 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r239 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r240 83 130 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.73 $Y2=3.33
r241 83 85 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.24 $Y2=3.33
r242 81 140 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=7.92 $Y2=3.33
r243 81 108 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6 $Y2=3.33
r244 79 103 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=5.68 $Y=3.33
+ $X2=5.52 $Y2=3.33
r245 79 80 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.68 $Y=3.33
+ $X2=5.81 $Y2=3.33
r246 78 107 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=5.94 $Y=3.33 $X2=6
+ $Y2=3.33
r247 78 80 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.94 $Y=3.33
+ $X2=5.81 $Y2=3.33
r248 73 76 4.37928 $w=2.48e-07 $l=9.5e-08 $layer=LI1_cond $X=4.07 $Y=2.63
+ $X2=4.165 $Y2=2.63
r249 69 154 3.00555 $w=3.3e-07 $l=1.07912e-07 $layer=LI1_cond $X=12.69 $Y=3.245
+ $X2=12.742 $Y2=3.33
r250 69 71 29.3349 $w=3.28e-07 $l=8.4e-07 $layer=LI1_cond $X=12.69 $Y=3.245
+ $X2=12.69 $Y2=2.405
r251 65 151 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.79 $Y=3.245
+ $X2=11.79 $Y2=3.33
r252 65 67 31.7795 $w=3.28e-07 $l=9.1e-07 $layer=LI1_cond $X=11.79 $Y=3.245
+ $X2=11.79 $Y2=2.335
r253 61 64 34.1617 $w=2.78e-07 $l=8.3e-07 $layer=LI1_cond $X=10.865 $Y=1.985
+ $X2=10.865 $Y2=2.815
r254 59 148 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=10.865 $Y=3.245
+ $X2=10.865 $Y2=3.33
r255 59 64 17.6982 $w=2.78e-07 $l=4.3e-07 $layer=LI1_cond $X=10.865 $Y=3.245
+ $X2=10.865 $Y2=2.815
r256 58 145 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.005 $Y=3.33
+ $X2=9.88 $Y2=3.33
r257 57 148 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=10.725 $Y=3.33
+ $X2=10.865 $Y2=3.33
r258 57 58 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=10.725 $Y=3.33
+ $X2=10.005 $Y2=3.33
r259 53 145 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.88 $Y=3.245
+ $X2=9.88 $Y2=3.33
r260 53 55 58.0831 $w=2.48e-07 $l=1.26e-06 $layer=LI1_cond $X=9.88 $Y=3.245
+ $X2=9.88 $Y2=1.985
r261 49 142 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.905 $Y=3.245
+ $X2=8.905 $Y2=3.33
r262 49 51 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=8.905 $Y=3.245
+ $X2=8.905 $Y2=2.815
r263 45 139 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.97 $Y=3.245
+ $X2=7.97 $Y2=3.33
r264 45 47 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=7.97 $Y=3.245
+ $X2=7.97 $Y2=2.815
r265 41 80 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=5.81 $Y=3.245
+ $X2=5.81 $Y2=3.33
r266 41 43 28.5895 $w=2.58e-07 $l=6.45e-07 $layer=LI1_cond $X=5.81 $Y=3.245
+ $X2=5.81 $Y2=2.6
r267 40 136 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.07 $Y=3.245
+ $X2=4.07 $Y2=3.33
r268 39 73 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.07 $Y=2.755
+ $X2=4.07 $Y2=2.63
r269 39 40 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=4.07 $Y=2.755
+ $X2=4.07 $Y2=3.245
r270 35 133 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.74 $Y=3.245
+ $X2=1.74 $Y2=3.33
r271 35 37 17.6359 $w=3.28e-07 $l=5.05e-07 $layer=LI1_cond $X=1.74 $Y=3.245
+ $X2=1.74 $Y2=2.74
r272 31 130 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=3.33
r273 31 33 17.9851 $w=3.28e-07 $l=5.15e-07 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=2.73
r274 10 71 300 $w=1.7e-07 $l=6.3559e-07 $layer=licon1_PDIFF $count=2 $X=12.54
+ $Y=1.84 $X2=12.69 $Y2=2.405
r275 9 67 300 $w=1.7e-07 $l=5.65044e-07 $layer=licon1_PDIFF $count=2 $X=11.64
+ $Y=1.84 $X2=11.79 $Y2=2.335
r276 8 64 600 $w=1.7e-07 $l=1.07941e-06 $layer=licon1_PDIFF $count=1 $X=10.67
+ $Y=1.84 $X2=10.89 $Y2=2.815
r277 8 61 300 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_PDIFF $count=2 $X=10.67
+ $Y=1.84 $X2=10.89 $Y2=1.985
r278 7 55 300 $w=1.7e-07 $l=1.99687e-07 $layer=licon1_PDIFF $count=2 $X=9.79
+ $Y=1.84 $X2=9.92 $Y2=1.985
r279 6 51 600 $w=1.7e-07 $l=3.33729e-07 $layer=licon1_PDIFF $count=1 $X=8.815
+ $Y=2.54 $X2=8.945 $Y2=2.815
r280 5 47 600 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=7.82
+ $Y=2.54 $X2=7.97 $Y2=2.815
r281 4 43 600 $w=1.7e-07 $l=5.07888e-07 $layer=licon1_PDIFF $count=1 $X=5.385
+ $Y=2.315 $X2=5.77 $Y2=2.6
r282 3 76 600 $w=1.7e-07 $l=3.47851e-07 $layer=licon1_PDIFF $count=1 $X=4
+ $Y=2.315 $X2=4.165 $Y2=2.59
r283 2 37 600 $w=1.7e-07 $l=9.72111e-07 $layer=licon1_PDIFF $count=1 $X=1.59
+ $Y=1.84 $X2=1.74 $Y2=2.74
r284 1 33 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=2.52 $X2=0.73 $Y2=2.73
.ends

.subckt PM_SKY130_FD_SC_LS__DFSTP_4%Q 1 2 3 4 15 17 18 19 21 27 31 33 37 39 40
+ 41 52
c73 18 0 1.09343e-19 $X=11.01 $Y=1.065
c74 15 0 1.85451e-19 $X=10.845 $Y=0.515
r75 51 52 4.56667 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=12.24 $Y=1.985
+ $X2=12.125 $Y2=1.985
r76 41 51 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=12.72 $Y=1.985
+ $X2=12.24 $Y2=1.985
r77 41 45 2.85155 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=12.72 $Y=1.985
+ $X2=12.72 $Y2=1.82
r78 40 45 7.76646 $w=2.28e-07 $l=1.55e-07 $layer=LI1_cond $X=12.72 $Y=1.665
+ $X2=12.72 $Y2=1.82
r79 39 40 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=12.72 $Y=1.295
+ $X2=12.72 $Y2=1.665
r80 38 39 7.2654 $w=2.28e-07 $l=1.45e-07 $layer=LI1_cond $X=12.72 $Y=1.15
+ $X2=12.72 $Y2=1.295
r81 34 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.345 $Y=1.065
+ $X2=12.18 $Y2=1.065
r82 33 38 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=12.605 $Y=1.065
+ $X2=12.72 $Y2=1.15
r83 33 34 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=12.605 $Y=1.065
+ $X2=12.345 $Y2=1.065
r84 29 51 2.85155 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=12.24 $Y=2.15
+ $X2=12.24 $Y2=1.985
r85 29 31 11.775 $w=2.28e-07 $l=2.35e-07 $layer=LI1_cond $X=12.24 $Y=2.15
+ $X2=12.24 $Y2=2.385
r86 25 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.18 $Y=0.98
+ $X2=12.18 $Y2=1.065
r87 25 27 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=12.18 $Y=0.98
+ $X2=12.18 $Y2=0.515
r88 24 36 3.54079 $w=2.6e-07 $l=1.4e-07 $layer=LI1_cond $X=11.455 $Y=1.95
+ $X2=11.315 $Y2=1.95
r89 24 52 29.6976 $w=2.58e-07 $l=6.7e-07 $layer=LI1_cond $X=11.455 $Y=1.95
+ $X2=12.125 $Y2=1.95
r90 19 36 3.28787 $w=2.8e-07 $l=1.3e-07 $layer=LI1_cond $X=11.315 $Y=2.08
+ $X2=11.315 $Y2=1.95
r91 19 21 12.5534 $w=2.78e-07 $l=3.05e-07 $layer=LI1_cond $X=11.315 $Y=2.08
+ $X2=11.315 $Y2=2.385
r92 17 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.015 $Y=1.065
+ $X2=12.18 $Y2=1.065
r93 17 18 65.5668 $w=1.68e-07 $l=1.005e-06 $layer=LI1_cond $X=12.015 $Y=1.065
+ $X2=11.01 $Y2=1.065
r94 13 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=10.845 $Y=0.98
+ $X2=11.01 $Y2=1.065
r95 13 15 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=10.845 $Y=0.98
+ $X2=10.845 $Y2=0.515
r96 4 51 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=12.09
+ $Y=1.84 $X2=12.24 $Y2=1.985
r97 4 31 300 $w=1.7e-07 $l=6.15447e-07 $layer=licon1_PDIFF $count=2 $X=12.09
+ $Y=1.84 $X2=12.24 $Y2=2.385
r98 3 36 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=11.19
+ $Y=1.84 $X2=11.34 $Y2=1.985
r99 3 21 300 $w=1.7e-07 $l=6.15447e-07 $layer=licon1_PDIFF $count=2 $X=11.19
+ $Y=1.84 $X2=11.34 $Y2=2.385
r100 2 27 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=11.995
+ $Y=0.37 $X2=12.18 $Y2=0.515
r101 1 15 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.705
+ $Y=0.37 $X2=10.845 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__DFSTP_4%VGND 1 2 3 4 5 6 7 8 27 29 33 37 41 45 49 51
+ 53 56 57 58 60 65 84 89 94 100 103 106 110 119 121 124 130
c144 33 0 9.68091e-20 $X=1.7 $Y=0.495
r145 129 130 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r146 125 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=11.28 $Y2=0
r147 124 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r148 124 125 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r149 121 122 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r150 117 119 9.64943 $w=7.53e-07 $l=7e-08 $layer=LI1_cond $X=8.88 $Y=0.292
+ $X2=8.95 $Y2=0.292
r151 117 118 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r152 115 117 1.505 $w=7.53e-07 $l=9.5e-08 $layer=LI1_cond $X=8.785 $Y=0.292
+ $X2=8.88 $Y2=0.292
r153 113 118 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0
+ $X2=8.88 $Y2=0
r154 112 115 6.09921 $w=7.53e-07 $l=3.85e-07 $layer=LI1_cond $X=8.4 $Y=0.292
+ $X2=8.785 $Y2=0.292
r155 112 113 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r156 109 112 4.75263 $w=7.53e-07 $l=3e-07 $layer=LI1_cond $X=8.1 $Y=0.292
+ $X2=8.4 $Y2=0.292
r157 109 110 11.1544 $w=7.53e-07 $l=1.65e-07 $layer=LI1_cond $X=8.1 $Y=0.292
+ $X2=7.935 $Y2=0.292
r158 106 107 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r159 103 104 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0
+ $X2=1.68 $Y2=0
r160 101 104 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0
+ $X2=1.68 $Y2=0
r161 100 101 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0
+ $X2=0.72 $Y2=0
r162 98 130 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=12.72 $Y2=0
r163 98 125 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=11.76 $Y2=0
r164 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r165 95 124 13.2917 $w=1.7e-07 $l=3.33e-07 $layer=LI1_cond $X=11.845 $Y=0
+ $X2=11.512 $Y2=0
r166 95 97 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=11.845 $Y=0
+ $X2=12.24 $Y2=0
r167 94 129 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=12.515 $Y=0
+ $X2=12.737 $Y2=0
r168 94 97 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=12.515 $Y=0
+ $X2=12.24 $Y2=0
r169 93 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=11.28 $Y2=0
r170 93 122 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=10.32 $Y2=0
r171 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=0 $X2=10.8
+ $Y2=0
r172 90 121 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.51 $Y=0
+ $X2=10.345 $Y2=0
r173 90 92 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=10.51 $Y=0 $X2=10.8
+ $Y2=0
r174 89 124 13.2917 $w=1.7e-07 $l=3.32e-07 $layer=LI1_cond $X=11.18 $Y=0
+ $X2=11.512 $Y2=0
r175 89 92 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=11.18 $Y=0 $X2=10.8
+ $Y2=0
r176 88 122 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=10.32 $Y2=0
r177 88 118 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=8.88 $Y2=0
r178 87 119 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=9.84 $Y=0 $X2=8.95
+ $Y2=0
r179 87 88 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r180 84 121 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.18 $Y=0
+ $X2=10.345 $Y2=0
r181 84 87 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=10.18 $Y=0 $X2=9.84
+ $Y2=0
r182 83 113 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.4
+ $Y2=0
r183 82 110 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=7.92 $Y=0
+ $X2=7.935 $Y2=0
r184 82 83 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r185 79 82 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=6 $Y=0 $X2=7.92
+ $Y2=0
r186 79 80 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6
+ $Y2=0
r187 76 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r188 75 76 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r189 73 76 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.52
+ $Y2=0
r190 73 107 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0
+ $X2=4.08 $Y2=0
r191 72 75 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.56 $Y=0 $X2=5.52
+ $Y2=0
r192 72 73 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r193 70 106 9.73034 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=4.42 $Y=0
+ $X2=4.222 $Y2=0
r194 70 72 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=4.42 $Y=0 $X2=4.56
+ $Y2=0
r195 69 107 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=4.08 $Y2=0
r196 69 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=1.68 $Y2=0
r197 68 69 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r198 66 103 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.865 $Y=0
+ $X2=1.74 $Y2=0
r199 66 68 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.865 $Y=0 $X2=2.16
+ $Y2=0
r200 65 106 9.73034 $w=1.7e-07 $l=1.97e-07 $layer=LI1_cond $X=4.025 $Y=0
+ $X2=4.222 $Y2=0
r201 65 68 121.674 $w=1.68e-07 $l=1.865e-06 $layer=LI1_cond $X=4.025 $Y=0
+ $X2=2.16 $Y2=0
r202 63 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0
+ $X2=0.72 $Y2=0
r203 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r204 60 100 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.545 $Y=0
+ $X2=0.67 $Y2=0
r205 60 62 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0
+ $X2=0.24 $Y2=0
r206 58 83 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=6.48 $Y=0
+ $X2=7.92 $Y2=0
r207 58 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r208 57 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.835 $Y=0 $X2=6
+ $Y2=0
r209 56 75 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=5.67 $Y=0 $X2=5.52
+ $Y2=0
r210 56 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.67 $Y=0 $X2=5.835
+ $Y2=0
r211 51 129 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=12.68 $Y=0.085
+ $X2=12.737 $Y2=0
r212 51 53 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=12.68 $Y=0.085
+ $X2=12.68 $Y2=0.645
r213 47 124 2.7522 $w=6.65e-07 $l=8.5e-08 $layer=LI1_cond $X=11.512 $Y=0.085
+ $X2=11.512 $Y2=0
r214 47 49 9.89238 $w=6.63e-07 $l=5.5e-07 $layer=LI1_cond $X=11.512 $Y=0.085
+ $X2=11.512 $Y2=0.635
r215 43 121 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.345 $Y=0.085
+ $X2=10.345 $Y2=0
r216 43 45 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=10.345 $Y=0.085
+ $X2=10.345 $Y2=0.515
r217 39 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.835 $Y=0.085
+ $X2=5.835 $Y2=0
r218 39 41 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=5.835 $Y=0.085
+ $X2=5.835 $Y2=0.515
r219 35 106 1.43204 $w=3.95e-07 $l=8.5e-08 $layer=LI1_cond $X=4.222 $Y=0.085
+ $X2=4.222 $Y2=0
r220 35 37 12.5456 $w=3.93e-07 $l=4.3e-07 $layer=LI1_cond $X=4.222 $Y=0.085
+ $X2=4.222 $Y2=0.515
r221 31 103 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.74 $Y=0.085
+ $X2=1.74 $Y2=0
r222 31 33 18.9001 $w=2.48e-07 $l=4.1e-07 $layer=LI1_cond $X=1.74 $Y=0.085
+ $X2=1.74 $Y2=0.495
r223 30 100 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.795 $Y=0
+ $X2=0.67 $Y2=0
r224 29 103 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.615 $Y=0
+ $X2=1.74 $Y2=0
r225 29 30 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=1.615 $Y=0
+ $X2=0.795 $Y2=0
r226 25 100 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.67 $Y=0.085
+ $X2=0.67 $Y2=0
r227 25 27 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=0.67 $Y=0.085
+ $X2=0.67 $Y2=0.58
r228 8 53 182 $w=1.7e-07 $l=3.65205e-07 $layer=licon1_NDIFF $count=1 $X=12.47
+ $Y=0.37 $X2=12.68 $Y2=0.645
r229 7 49 91 $w=1.7e-07 $l=6.89891e-07 $layer=licon1_NDIFF $count=2 $X=11.135
+ $Y=0.37 $X2=11.705 $Y2=0.635
r230 6 45 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.205
+ $Y=0.37 $X2=10.345 $Y2=0.515
r231 5 115 121.333 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_NDIFF $count=1
+ $X=7.96 $Y=0.44 $X2=8.785 $Y2=0.585
r232 5 109 121.333 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1
+ $X=7.96 $Y=0.44 $X2=8.1 $Y2=0.585
r233 4 41 91 $w=1.7e-07 $l=3.05205e-07 $layer=licon1_NDIFF $count=2 $X=5.565
+ $Y=0.59 $X2=5.835 $Y2=0.515
r234 3 37 182 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_NDIFF $count=1 $X=4.05
+ $Y=0.37 $X2=4.22 $Y2=0.515
r235 2 33 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.56
+ $Y=0.37 $X2=1.7 $Y2=0.495
r236 1 27 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.58
.ends

