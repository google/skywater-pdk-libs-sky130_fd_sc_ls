* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__or4b_1 A B C D_N VGND VNB VPB VPWR X
M1000 VGND C a_228_74# VNB nshort w=550000u l=150000u
+  ad=7.8175e+11p pd=6.35e+06u as=6.6275e+11p ps=4.61e+06u
M1001 a_356_368# a_27_74# a_228_74# VPB phighvt w=1e+06u l=150000u
+  ad=2.7e+11p pd=2.54e+06u as=2.95e+11p ps=2.59e+06u
M1002 VPWR A a_524_368# VPB phighvt w=1e+06u l=150000u
+  ad=8.712e+11p pd=5.69e+06u as=3.9e+11p ps=2.78e+06u
M1003 a_524_368# B a_440_368# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1004 X a_228_74# VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1005 X a_228_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=0p ps=0u
M1006 VPWR D_N a_27_74# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=2.478e+11p ps=2.27e+06u
M1007 a_228_74# B VGND VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND D_N a_27_74# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1009 a_440_368# C a_356_368# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_228_74# a_27_74# VGND VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND A a_228_74# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
