* File: sky130_fd_sc_ls__nor4b_1.pex.spice
* Created: Fri Aug 28 13:40:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__NOR4B_1%D_N 2 3 5 8 10 13
c40 13 0 1.706e-19 $X=0.61 $Y=1.275
r41 13 16 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.61 $Y=1.275
+ $X2=0.61 $Y2=1.44
r42 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.61 $Y=1.275
+ $X2=0.61 $Y2=1.11
r43 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.61
+ $Y=1.275 $X2=0.61 $Y2=1.275
r44 10 14 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=0.72 $Y=1.275
+ $X2=0.61 $Y2=1.275
r45 8 15 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.67 $Y=0.645
+ $X2=0.67 $Y2=1.11
r46 3 5 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.655 $Y=1.765
+ $X2=0.655 $Y2=2.26
r47 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.655 $Y=1.675 $X2=0.655
+ $Y2=1.765
r48 2 16 91.3468 $w=1.8e-07 $l=2.35e-07 $layer=POLY_cond $X=0.655 $Y=1.675
+ $X2=0.655 $Y2=1.44
.ends

.subckt PM_SKY130_FD_SC_LS__NOR4B_1%A 1 3 6 8 12
c34 12 0 1.02415e-19 $X=1.15 $Y=1.515
r35 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.15
+ $Y=1.515 $X2=1.15 $Y2=1.515
r36 8 12 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.15 $Y=1.665
+ $X2=1.15 $Y2=1.515
r37 4 11 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=1.24 $Y=1.35
+ $X2=1.15 $Y2=1.515
r38 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.24 $Y=1.35 $X2=1.24
+ $Y2=0.74
r39 1 11 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=1.225 $Y=1.765
+ $X2=1.15 $Y2=1.515
r40 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.225 $Y=1.765
+ $X2=1.225 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__NOR4B_1%B 1 3 6 8 12
r31 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.69
+ $Y=1.515 $X2=1.69 $Y2=1.515
r32 8 12 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.69 $Y=1.665
+ $X2=1.69 $Y2=1.515
r33 4 11 38.5562 $w=2.99e-07 $l=1.74714e-07 $layer=POLY_cond $X=1.67 $Y=1.35
+ $X2=1.69 $Y2=1.515
r34 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.67 $Y=1.35 $X2=1.67
+ $Y2=0.74
r35 1 11 52.2586 $w=2.99e-07 $l=2.7157e-07 $layer=POLY_cond $X=1.645 $Y=1.765
+ $X2=1.69 $Y2=1.515
r36 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.645 $Y=1.765
+ $X2=1.645 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__NOR4B_1%C 1 3 6 8 12
r32 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.23
+ $Y=1.515 $X2=2.23 $Y2=1.515
r33 8 12 4.93904 $w=3.48e-07 $l=1.5e-07 $layer=LI1_cond $X=2.22 $Y=1.665
+ $X2=2.22 $Y2=1.515
r34 4 11 38.5562 $w=2.99e-07 $l=1.74714e-07 $layer=POLY_cond $X=2.25 $Y=1.35
+ $X2=2.23 $Y2=1.515
r35 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.25 $Y=1.35 $X2=2.25
+ $Y2=0.74
r36 1 11 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=2.155 $Y=1.765
+ $X2=2.23 $Y2=1.515
r37 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.155 $Y=1.765
+ $X2=2.155 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__NOR4B_1%A_57_368# 1 2 9 11 13 18 21 25 28 29 30 34
r70 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.77
+ $Y=1.515 $X2=2.77 $Y2=1.515
r71 31 34 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=2.65 $Y=1.515
+ $X2=2.77 $Y2=1.515
r72 28 30 1.22049 $w=4.88e-07 $l=5e-08 $layer=LI1_cond $X=0.35 $Y=1.985 $X2=0.35
+ $Y2=2.035
r73 28 29 9.45624 $w=4.88e-07 $l=1.65e-07 $layer=LI1_cond $X=0.35 $Y=1.985
+ $X2=0.35 $Y2=1.82
r74 22 25 5.37222 $w=5.88e-07 $l=2.65e-07 $layer=LI1_cond $X=0.19 $Y=0.645
+ $X2=0.455 $Y2=0.645
r75 20 31 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.65 $Y=1.68
+ $X2=2.65 $Y2=1.515
r76 20 21 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=2.65 $Y=1.68 $X2=2.65
+ $Y2=1.95
r77 19 30 7.03003 $w=1.7e-07 $l=2.45e-07 $layer=LI1_cond $X=0.595 $Y=2.035
+ $X2=0.35 $Y2=2.035
r78 18 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.565 $Y=2.035
+ $X2=2.65 $Y2=1.95
r79 18 19 128.524 $w=1.68e-07 $l=1.97e-06 $layer=LI1_cond $X=2.565 $Y=2.035
+ $X2=0.595 $Y2=2.035
r80 14 22 8.20854 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=0.19 $Y=0.94
+ $X2=0.19 $Y2=0.645
r81 14 29 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=0.19 $Y=0.94
+ $X2=0.19 $Y2=1.82
r82 11 35 52.2586 $w=2.99e-07 $l=2.7157e-07 $layer=POLY_cond $X=2.725 $Y=1.765
+ $X2=2.77 $Y2=1.515
r83 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.725 $Y=1.765
+ $X2=2.725 $Y2=2.4
r84 7 35 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=2.68 $Y=1.35
+ $X2=2.77 $Y2=1.515
r85 7 9 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.68 $Y=1.35 $X2=2.68
+ $Y2=0.74
r86 2 28 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.285
+ $Y=1.84 $X2=0.43 $Y2=1.985
r87 1 25 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=0.31
+ $Y=0.37 $X2=0.455 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_LS__NOR4B_1%VPWR 1 6 9 10 11 21 22
r26 21 22 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r27 18 21 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=3.12 $Y2=3.33
r28 18 19 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r29 15 19 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r30 14 15 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r31 11 22 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=3.12 $Y2=3.33
r32 11 19 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r33 9 14 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=0.835 $Y=3.33
+ $X2=0.72 $Y2=3.33
r34 9 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.835 $Y=3.33 $X2=1
+ $Y2=3.33
r35 8 18 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=1.165 $Y=3.33 $X2=1.2
+ $Y2=3.33
r36 8 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.165 $Y=3.33 $X2=1
+ $Y2=3.33
r37 4 10 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1 $Y=3.245 $X2=1
+ $Y2=3.33
r38 4 6 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=1 $Y=3.245 $X2=1
+ $Y2=2.455
r39 1 6 300 $w=1.7e-07 $l=7.3775e-07 $layer=licon1_PDIFF $count=2 $X=0.73
+ $Y=1.84 $X2=1 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_LS__NOR4B_1%Y 1 2 3 12 14 15 18 20 24 25 26 27 43
c59 15 0 6.81849e-20 $X=1.62 $Y=1.095
r60 26 27 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.09 $Y=2.405
+ $X2=3.09 $Y2=2.775
r61 25 43 7.82243 $w=3.68e-07 $l=1.42e-07 $layer=LI1_cond $X=3.09 $Y=1.992
+ $X2=3.09 $Y2=1.85
r62 25 26 10.2163 $w=3.68e-07 $l=3.28e-07 $layer=LI1_cond $X=3.09 $Y=2.077
+ $X2=3.09 $Y2=2.405
r63 22 43 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.19 $Y=1.18
+ $X2=3.19 $Y2=1.85
r64 21 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.63 $Y=1.095
+ $X2=2.465 $Y2=1.095
r65 20 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.105 $Y=1.095
+ $X2=3.19 $Y2=1.18
r66 20 21 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=3.105 $Y=1.095
+ $X2=2.63 $Y2=1.095
r67 16 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.465 $Y=1.01
+ $X2=2.465 $Y2=1.095
r68 16 18 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=2.465 $Y=1.01
+ $X2=2.465 $Y2=0.515
r69 14 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.3 $Y=1.095
+ $X2=2.465 $Y2=1.095
r70 14 15 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.3 $Y=1.095
+ $X2=1.62 $Y2=1.095
r71 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.455 $Y=1.01
+ $X2=1.62 $Y2=1.095
r72 10 12 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=1.455 $Y=1.01
+ $X2=1.455 $Y2=0.515
r73 3 25 400 $w=1.7e-07 $l=3.46627e-07 $layer=licon1_PDIFF $count=1 $X=2.8
+ $Y=1.84 $X2=3.07 $Y2=2.015
r74 3 27 400 $w=1.7e-07 $l=1.10176e-06 $layer=licon1_PDIFF $count=1 $X=2.8
+ $Y=1.84 $X2=3.07 $Y2=2.815
r75 2 18 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.325
+ $Y=0.37 $X2=2.465 $Y2=0.515
r76 1 12 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.315
+ $Y=0.37 $X2=1.455 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__NOR4B_1%VGND 1 2 3 12 16 18 20 23 24 26 27 28 37 43
r43 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r44 40 43 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r45 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r46 37 42 4.53027 $w=1.7e-07 $l=2.8e-07 $layer=LI1_cond $X=2.8 $Y=0 $X2=3.08
+ $Y2=0
r47 37 39 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=2.8 $Y=0 $X2=2.64
+ $Y2=0
r48 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r49 28 40 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r50 28 32 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r51 28 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r52 26 35 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=1.79 $Y=0 $X2=1.68
+ $Y2=0
r53 26 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.79 $Y=0 $X2=1.955
+ $Y2=0
r54 25 39 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.12 $Y=0 $X2=2.64
+ $Y2=0
r55 25 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.12 $Y=0 $X2=1.955
+ $Y2=0
r56 23 31 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=0.79 $Y=0 $X2=0.72
+ $Y2=0
r57 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.79 $Y=0 $X2=0.955
+ $Y2=0
r58 22 35 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.12 $Y=0 $X2=1.68
+ $Y2=0
r59 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.12 $Y=0 $X2=0.955
+ $Y2=0
r60 18 42 3.23591 $w=3.3e-07 $l=1.51658e-07 $layer=LI1_cond $X=2.965 $Y=0.085
+ $X2=3.08 $Y2=0
r61 18 20 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=2.965 $Y=0.085
+ $X2=2.965 $Y2=0.595
r62 14 27 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.955 $Y=0.085
+ $X2=1.955 $Y2=0
r63 14 16 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=1.955 $Y=0.085
+ $X2=1.955 $Y2=0.595
r64 10 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.955 $Y=0.085
+ $X2=0.955 $Y2=0
r65 10 12 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=0.955 $Y=0.085
+ $X2=0.955 $Y2=0.645
r66 3 20 182 $w=1.7e-07 $l=3.1285e-07 $layer=licon1_NDIFF $count=1 $X=2.755
+ $Y=0.37 $X2=2.965 $Y2=0.595
r67 2 16 182 $w=1.7e-07 $l=3.1285e-07 $layer=licon1_NDIFF $count=1 $X=1.745
+ $Y=0.37 $X2=1.955 $Y2=0.595
r68 1 12 182 $w=1.7e-07 $l=3.65205e-07 $layer=licon1_NDIFF $count=1 $X=0.745
+ $Y=0.37 $X2=0.955 $Y2=0.645
.ends

