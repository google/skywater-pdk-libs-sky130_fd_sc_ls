* NGSPICE file created from sky130_fd_sc_ls__sdfrtp_2.ext - technology: sky130A

.subckt sky130_fd_sc_ls__sdfrtp_2 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
M1000 a_1320_119# a_1034_392# a_1234_119# VNB nshort w=420000u l=150000u
+  ad=9.87e+10p pd=1.31e+06u as=1.176e+11p ps=1.4e+06u
M1001 a_1234_119# RESET_B VPWR VPB phighvt w=420000u l=150000u
+  ad=2.499e+11p pd=2.87e+06u as=3.0042e+12p ps=2.284e+07u
M1002 a_2078_74# a_835_98# a_1824_74# VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=5.504e+11p ps=3.72e+06u
M1003 VGND a_2082_446# a_2078_74# VNB nshort w=420000u l=150000u
+  ad=2.07625e+12p pd=1.687e+07u as=0p ps=0u
M1004 a_390_81# D a_340_464# VPB phighvt w=640000u l=150000u
+  ad=4.983e+11p pd=5.16e+06u as=1.728e+11p ps=1.82e+06u
M1005 a_312_81# a_27_74# a_225_81# VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=2.499e+11p ps=2.87e+06u
M1006 a_390_81# D a_312_81# VNB nshort w=420000u l=150000u
+  ad=3.738e+11p pd=3.46e+06u as=0p ps=0u
M1007 a_2082_446# a_1824_74# a_2242_74# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=8.82e+10p ps=1.26e+06u
M1008 a_1332_457# a_835_98# a_1234_119# VPB phighvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1009 VGND RESET_B a_1397_119# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1010 a_2492_392# a_1824_74# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.95e+11p pd=2.59e+06u as=0p ps=0u
M1011 a_225_81# SCD a_545_81# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1012 Q a_2492_392# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=0p ps=0u
M1013 a_2082_446# RESET_B VPWR VPB phighvt w=420000u l=150000u
+  ad=1.26e+11p pd=1.44e+06u as=0p ps=0u
M1014 a_2242_74# RESET_B VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_1367_93# a_1234_119# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=4.9755e+11p pd=3.13e+06u as=0p ps=0u
M1016 a_1824_74# a_1034_392# a_1367_93# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.627e+11p ps=2.19e+06u
M1017 a_512_464# a_27_74# a_390_81# VPB phighvt w=640000u l=150000u
+  ad=2.56e+11p pd=2.08e+06u as=0p ps=0u
M1018 a_1824_74# a_835_98# a_1367_93# VPB phighvt w=1e+06u l=150000u
+  ad=4.4725e+11p pd=3.66e+06u as=0p ps=0u
M1019 a_1397_119# a_1367_93# a_1320_119# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR a_2492_392# Q VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_2492_392# a_1824_74# VGND VNB nshort w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=0p ps=0u
M1022 VPWR SCE a_27_74# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.888e+11p ps=1.87e+06u
M1023 VGND a_2492_392# Q VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.072e+11p ps=2.04e+06u
M1024 VPWR a_1824_74# a_2082_446# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_340_464# SCE VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_545_81# SCE a_390_81# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VPWR SCD a_512_464# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VPWR CLK a_835_98# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.95e+11p ps=2.59e+06u
M1029 VGND CLK a_835_98# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.619e+11p ps=2.38e+06u
M1030 a_1034_392# a_835_98# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.95e+11p pd=2.59e+06u as=0p ps=0u
M1031 VGND SCE a_27_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1032 a_1034_392# a_835_98# VGND VNB nshort w=740000u l=150000u
+  ad=1.961e+11p pd=2.01e+06u as=0p ps=0u
M1033 VPWR a_1367_93# a_1332_457# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_1234_119# a_835_98# a_390_81# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_1367_93# a_1234_119# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 VGND RESET_B a_225_81# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_2037_508# a_1034_392# a_1824_74# VPB phighvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1038 VPWR a_2082_446# a_2037_508# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_390_81# RESET_B VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1040 a_1234_119# a_1034_392# a_390_81# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1041 Q a_2492_392# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

