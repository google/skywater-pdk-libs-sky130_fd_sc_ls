* File: sky130_fd_sc_ls__o41a_4.spice
* Created: Fri Aug 28 13:55:55 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__o41a_4.pex.spice"
.subckt sky130_fd_sc_ls__o41a_4  VNB VPB B1 A4 A3 A1 A2 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A2	A2
* A1	A1
* A3	A3
* A4	A4
* B1	B1
* VPB	VPB
* VNB	VNB
MM1006 N_X_M1006_d N_A_110_48#_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.2627 PD=1.02 PS=2.19 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75000.3
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1012 N_X_M1006_d N_A_110_48#_M1012_g N_VGND_M1012_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.7
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1016 N_X_M1016_d N_A_110_48#_M1016_g N_VGND_M1012_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.2
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1024 N_X_M1016_d N_A_110_48#_M1024_g N_VGND_M1024_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1003 N_A_523_124#_M1003_d N_B1_M1003_g N_A_110_48#_M1003_s VNB NSHORT L=0.15
+ W=0.64 AD=0.1824 AS=0.0896 PD=1.85 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75004.5 A=0.096 P=1.58 MULT=1
MM1011 N_A_523_124#_M1011_d N_B1_M1011_g N_A_110_48#_M1003_s VNB NSHORT L=0.15
+ W=0.64 AD=0.1184 AS=0.0896 PD=1.01 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75004 A=0.096 P=1.58 MULT=1
MM1002 N_A_523_124#_M1011_d N_A3_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.64
+ AD=0.1184 AS=0.19135 PD=1.01 PS=1.26 NRD=16.872 NRS=60 M=1 R=4.26667
+ SA=75001.2 SB=75003.5 A=0.096 P=1.58 MULT=1
MM1001 N_A_523_124#_M1001_d N_A4_M1001_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.19135 PD=0.92 PS=1.26 NRD=0 NRS=0 M=1 R=4.26667 SA=75001.9
+ SB=75002.9 A=0.096 P=1.58 MULT=1
MM1026 N_A_523_124#_M1001_d N_A4_M1026_g N_VGND_M1026_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75002.3
+ SB=75002.4 A=0.096 P=1.58 MULT=1
MM1013 N_A_523_124#_M1013_d N_A3_M1013_g N_VGND_M1026_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0928 AS=0.0896 PD=0.93 PS=0.92 NRD=0.936 NRS=0 M=1 R=4.26667 SA=75002.7
+ SB=75002 A=0.096 P=1.58 MULT=1
MM1005 N_A_523_124#_M1013_d N_A2_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0928 AS=0.0896 PD=0.93 PS=0.92 NRD=0.936 NRS=0 M=1 R=4.26667 SA=75003.2
+ SB=75001.6 A=0.096 P=1.58 MULT=1
MM1007 N_A_523_124#_M1007_d N_A1_M1007_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75003.6
+ SB=75001.1 A=0.096 P=1.58 MULT=1
MM1009 N_A_523_124#_M1007_d N_A1_M1009_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.113125 PD=0.92 PS=1.005 NRD=0 NRS=0 M=1 R=4.26667 SA=75004
+ SB=75000.7 A=0.096 P=1.58 MULT=1
MM1020 N_A_523_124#_M1020_d N_A2_M1020_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.64
+ AD=0.1824 AS=0.113125 PD=1.85 PS=1.005 NRD=0 NRS=13.116 M=1 R=4.26667
+ SA=75004.5 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1000 N_X_M1000_d N_A_110_48#_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75002.3 A=0.168 P=2.54 MULT=1
MM1004 N_X_M1000_d N_A_110_48#_M1004_g N_VPWR_M1004_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75001.9 A=0.168 P=2.54 MULT=1
MM1014 N_X_M1014_d N_A_110_48#_M1014_g N_VPWR_M1004_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75001.4 A=0.168 P=2.54 MULT=1
MM1021 N_X_M1014_d N_A_110_48#_M1021_g N_VPWR_M1021_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.228743 PD=1.42 PS=1.72 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.6 SB=75001 A=0.168 P=2.54 MULT=1
MM1010 N_A_110_48#_M1010_d N_B1_M1010_g N_VPWR_M1021_s VPB PHIGHVT L=0.15 W=0.84
+ AD=0.126 AS=0.171557 PD=1.14 PS=1.29 NRD=2.3443 NRS=22.261 M=1 R=5.6
+ SA=75002.1 SB=75000.7 A=0.126 P=1.98 MULT=1
MM1018 N_A_110_48#_M1010_d N_B1_M1018_g N_VPWR_M1018_s VPB PHIGHVT L=0.15 W=0.84
+ AD=0.126 AS=0.2478 PD=1.14 PS=2.27 NRD=2.3443 NRS=2.3443 M=1 R=5.6 SA=75002.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1015 N_A_762_368#_M1015_d N_A3_M1015_g N_A_851_368#_M1015_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75003.5 A=0.168 P=2.54 MULT=1
MM1022 N_A_851_368#_M1015_s N_A4_M1022_g N_A_110_48#_M1022_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.1736 PD=1.42 PS=1.43 NRD=1.7533 NRS=2.6201 M=1 R=7.46667
+ SA=75000.7 SB=75003.1 A=0.168 P=2.54 MULT=1
MM1025 N_A_851_368#_M1025_d N_A4_M1025_g N_A_110_48#_M1022_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.1736 PD=1.42 PS=1.43 NRD=1.7533 NRS=2.6201 M=1 R=7.46667
+ SA=75001.1 SB=75002.6 A=0.168 P=2.54 MULT=1
MM1019 N_A_762_368#_M1019_d N_A3_M1019_g N_A_851_368#_M1025_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.6 SB=75002.2 A=0.168 P=2.54 MULT=1
MM1017 N_A_762_368#_M1019_d N_A2_M1017_g N_A_1213_368#_M1017_s VPB PHIGHVT
+ L=0.15 W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1
+ R=7.46667 SA=75002 SB=75001.7 A=0.168 P=2.54 MULT=1
MM1008 N_A_1213_368#_M1017_s N_A1_M1008_g N_VPWR_M1008_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.1904 PD=1.42 PS=1.46 NRD=1.7533 NRS=5.2599 M=1 R=7.46667
+ SA=75002.5 SB=75001.3 A=0.168 P=2.54 MULT=1
MM1027 N_A_1213_368#_M1027_d N_A1_M1027_g N_VPWR_M1008_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.196 AS=0.1904 PD=1.47 PS=1.46 NRD=10.5395 NRS=5.2599 M=1 R=7.46667
+ SA=75003 SB=75000.8 A=0.168 P=2.54 MULT=1
MM1023 N_A_762_368#_M1023_d N_A2_M1023_g N_A_1213_368#_M1027_d VPB PHIGHVT
+ L=0.15 W=1.12 AD=0.3864 AS=0.196 PD=2.93 PS=1.47 NRD=10.5395 NRS=1.7533 M=1
+ R=7.46667 SA=75003.5 SB=75000.3 A=0.168 P=2.54 MULT=1
DX28_noxref VNB VPB NWDIODE A=15.8844 P=20.8
*
.include "sky130_fd_sc_ls__o41a_4.pxi.spice"
*
.ends
*
*
