* File: sky130_fd_sc_ls__dfbbn_1.pxi.spice
* Created: Wed Sep  2 11:00:23 2020
* 
x_PM_SKY130_FD_SC_LS__DFBBN_1%CLK_N N_CLK_N_M1033_g N_CLK_N_c_276_n
+ N_CLK_N_M1030_g CLK_N N_CLK_N_c_277_n PM_SKY130_FD_SC_LS__DFBBN_1%CLK_N
x_PM_SKY130_FD_SC_LS__DFBBN_1%D N_D_M1013_g N_D_c_307_n N_D_c_311_n N_D_M1037_g
+ D D N_D_c_309_n PM_SKY130_FD_SC_LS__DFBBN_1%D
x_PM_SKY130_FD_SC_LS__DFBBN_1%A_474_405# N_A_474_405#_M1016_d
+ N_A_474_405#_M1019_s N_A_474_405#_M1027_d N_A_474_405#_M1011_g
+ N_A_474_405#_c_355_n N_A_474_405#_M1015_g N_A_474_405#_M1021_g
+ N_A_474_405#_c_351_n N_A_474_405#_M1017_g N_A_474_405#_c_357_n
+ N_A_474_405#_c_358_n N_A_474_405#_c_359_n N_A_474_405#_c_360_n
+ N_A_474_405#_c_352_n N_A_474_405#_c_353_n N_A_474_405#_c_423_p
+ N_A_474_405#_c_362_n N_A_474_405#_c_363_n N_A_474_405#_c_364_n
+ N_A_474_405#_c_365_n N_A_474_405#_c_366_n N_A_474_405#_c_367_n
+ PM_SKY130_FD_SC_LS__DFBBN_1%A_474_405#
x_PM_SKY130_FD_SC_LS__DFBBN_1%A_200_74# N_A_200_74#_M1034_d N_A_200_74#_M1031_d
+ N_A_200_74#_c_534_n N_A_200_74#_M1035_g N_A_200_74#_M1004_g
+ N_A_200_74#_c_519_n N_A_200_74#_M1003_g N_A_200_74#_c_520_n
+ N_A_200_74#_M1018_g N_A_200_74#_c_536_n N_A_200_74#_c_521_n
+ N_A_200_74#_c_537_n N_A_200_74#_c_538_n N_A_200_74#_c_539_n
+ N_A_200_74#_c_540_n N_A_200_74#_c_554_n N_A_200_74#_c_522_n
+ N_A_200_74#_c_541_n N_A_200_74#_c_523_n N_A_200_74#_c_524_n
+ N_A_200_74#_c_525_n N_A_200_74#_c_543_n N_A_200_74#_c_526_n
+ N_A_200_74#_c_527_n N_A_200_74#_c_545_n N_A_200_74#_c_528_n
+ N_A_200_74#_c_558_n N_A_200_74#_c_529_n N_A_200_74#_c_530_n
+ N_A_200_74#_c_531_n N_A_200_74#_c_532_n N_A_200_74#_c_533_n
+ PM_SKY130_FD_SC_LS__DFBBN_1%A_200_74#
x_PM_SKY130_FD_SC_LS__DFBBN_1%A_595_119# N_A_595_119#_M1001_d
+ N_A_595_119#_M1035_d N_A_595_119#_c_740_n N_A_595_119#_c_741_n
+ N_A_595_119#_c_749_n N_A_595_119#_M1019_g N_A_595_119#_M1016_g
+ N_A_595_119#_c_743_n N_A_595_119#_c_762_n N_A_595_119#_c_769_n
+ N_A_595_119#_c_750_n N_A_595_119#_c_744_n N_A_595_119#_c_745_n
+ N_A_595_119#_c_746_n N_A_595_119#_c_747_n
+ PM_SKY130_FD_SC_LS__DFBBN_1%A_595_119#
x_PM_SKY130_FD_SC_LS__DFBBN_1%A_978_357# N_A_978_357#_M1008_s
+ N_A_978_357#_M1005_s N_A_978_357#_c_848_n N_A_978_357#_M1020_g
+ N_A_978_357#_M1026_g N_A_978_357#_M1032_g N_A_978_357#_c_850_n
+ N_A_978_357#_c_866_n N_A_978_357#_M1039_g N_A_978_357#_c_851_n
+ N_A_978_357#_c_852_n N_A_978_357#_c_853_n N_A_978_357#_c_854_n
+ N_A_978_357#_c_855_n N_A_978_357#_c_912_p N_A_978_357#_c_941_p
+ N_A_978_357#_c_856_n N_A_978_357#_c_857_n N_A_978_357#_c_858_n
+ N_A_978_357#_c_859_n N_A_978_357#_c_860_n N_A_978_357#_c_868_n
+ N_A_978_357#_c_869_n N_A_978_357#_c_861_n N_A_978_357#_c_938_p
+ N_A_978_357#_c_862_n N_A_978_357#_c_863_n
+ PM_SKY130_FD_SC_LS__DFBBN_1%A_978_357#
x_PM_SKY130_FD_SC_LS__DFBBN_1%SET_B N_SET_B_c_1027_n N_SET_B_M1027_g
+ N_SET_B_M1022_g N_SET_B_c_1029_n N_SET_B_c_1030_n N_SET_B_c_1035_n
+ N_SET_B_M1007_g N_SET_B_M1014_g N_SET_B_c_1036_n N_SET_B_c_1051_n SET_B
+ N_SET_B_c_1037_n N_SET_B_c_1032_n PM_SKY130_FD_SC_LS__DFBBN_1%SET_B
x_PM_SKY130_FD_SC_LS__DFBBN_1%A_27_74# N_A_27_74#_M1033_s N_A_27_74#_M1030_s
+ N_A_27_74#_M1034_g N_A_27_74#_c_1158_n N_A_27_74#_M1031_g N_A_27_74#_c_1159_n
+ N_A_27_74#_c_1160_n N_A_27_74#_M1001_g N_A_27_74#_c_1162_n N_A_27_74#_c_1175_n
+ N_A_27_74#_c_1176_n N_A_27_74#_c_1177_n N_A_27_74#_c_1178_n
+ N_A_27_74#_c_1179_n N_A_27_74#_M1036_g N_A_27_74#_M1024_g N_A_27_74#_c_1164_n
+ N_A_27_74#_c_1165_n N_A_27_74#_c_1180_n N_A_27_74#_c_1181_n
+ N_A_27_74#_c_1182_n N_A_27_74#_M1012_g N_A_27_74#_c_1166_n N_A_27_74#_c_1183_n
+ N_A_27_74#_c_1167_n N_A_27_74#_c_1185_n N_A_27_74#_c_1186_n
+ N_A_27_74#_c_1168_n N_A_27_74#_c_1169_n N_A_27_74#_c_1170_n
+ N_A_27_74#_c_1200_n N_A_27_74#_c_1171_n N_A_27_74#_c_1172_n
+ N_A_27_74#_c_1173_n PM_SKY130_FD_SC_LS__DFBBN_1%A_27_74#
x_PM_SKY130_FD_SC_LS__DFBBN_1%A_1534_446# N_A_1534_446#_M1032_d
+ N_A_1534_446#_M1007_s N_A_1534_446#_M1028_d N_A_1534_446#_c_1354_n
+ N_A_1534_446#_M1010_g N_A_1534_446#_M1038_g N_A_1534_446#_c_1356_n
+ N_A_1534_446#_M1023_g N_A_1534_446#_M1025_g N_A_1534_446#_c_1344_n
+ N_A_1534_446#_c_1345_n N_A_1534_446#_c_1346_n N_A_1534_446#_c_1347_n
+ N_A_1534_446#_c_1359_n N_A_1534_446#_M1002_g N_A_1534_446#_c_1348_n
+ N_A_1534_446#_M1000_g N_A_1534_446#_c_1349_n N_A_1534_446#_c_1350_n
+ N_A_1534_446#_c_1360_n N_A_1534_446#_c_1361_n N_A_1534_446#_c_1362_n
+ N_A_1534_446#_c_1481_p N_A_1534_446#_c_1363_n N_A_1534_446#_c_1351_n
+ N_A_1534_446#_c_1364_n N_A_1534_446#_c_1365_n N_A_1534_446#_c_1366_n
+ N_A_1534_446#_c_1367_n N_A_1534_446#_c_1368_n N_A_1534_446#_c_1369_n
+ N_A_1534_446#_c_1352_n N_A_1534_446#_c_1353_n
+ PM_SKY130_FD_SC_LS__DFBBN_1%A_1534_446#
x_PM_SKY130_FD_SC_LS__DFBBN_1%A_1349_114# N_A_1349_114#_M1024_d
+ N_A_1349_114#_M1003_d N_A_1349_114#_M1029_g N_A_1349_114#_c_1554_n
+ N_A_1349_114#_M1028_g N_A_1349_114#_c_1555_n N_A_1349_114#_c_1559_n
+ N_A_1349_114#_c_1560_n N_A_1349_114#_c_1561_n N_A_1349_114#_c_1556_n
+ N_A_1349_114#_c_1563_n N_A_1349_114#_c_1564_n N_A_1349_114#_c_1633_n
+ N_A_1349_114#_c_1565_n N_A_1349_114#_c_1637_n N_A_1349_114#_c_1566_n
+ N_A_1349_114#_c_1567_n N_A_1349_114#_c_1557_n N_A_1349_114#_c_1569_n
+ N_A_1349_114#_c_1570_n N_A_1349_114#_c_1571_n
+ PM_SKY130_FD_SC_LS__DFBBN_1%A_1349_114#
x_PM_SKY130_FD_SC_LS__DFBBN_1%RESET_B N_RESET_B_c_1703_n N_RESET_B_M1005_g
+ N_RESET_B_M1008_g RESET_B N_RESET_B_c_1705_n
+ PM_SKY130_FD_SC_LS__DFBBN_1%RESET_B
x_PM_SKY130_FD_SC_LS__DFBBN_1%A_2412_410# N_A_2412_410#_M1000_s
+ N_A_2412_410#_M1002_s N_A_2412_410#_c_1741_n N_A_2412_410#_M1006_g
+ N_A_2412_410#_M1009_g N_A_2412_410#_c_1736_n N_A_2412_410#_c_1737_n
+ N_A_2412_410#_c_1738_n N_A_2412_410#_c_1739_n N_A_2412_410#_c_1740_n
+ PM_SKY130_FD_SC_LS__DFBBN_1%A_2412_410#
x_PM_SKY130_FD_SC_LS__DFBBN_1%VPWR N_VPWR_M1030_d N_VPWR_M1037_d N_VPWR_M1020_d
+ N_VPWR_M1017_s N_VPWR_M1010_d N_VPWR_M1007_d N_VPWR_M1005_d N_VPWR_M1002_d
+ N_VPWR_c_1793_n N_VPWR_c_1794_n N_VPWR_c_1795_n N_VPWR_c_1796_n
+ N_VPWR_c_1797_n N_VPWR_c_1798_n N_VPWR_c_1799_n N_VPWR_c_1800_n
+ N_VPWR_c_1801_n N_VPWR_c_1802_n VPWR N_VPWR_c_1803_n N_VPWR_c_1804_n
+ N_VPWR_c_1805_n N_VPWR_c_1806_n N_VPWR_c_1807_n N_VPWR_c_1808_n
+ N_VPWR_c_1809_n N_VPWR_c_1792_n N_VPWR_c_1811_n N_VPWR_c_1812_n
+ N_VPWR_c_1813_n N_VPWR_c_1814_n N_VPWR_c_1815_n N_VPWR_c_1816_n
+ PM_SKY130_FD_SC_LS__DFBBN_1%VPWR
x_PM_SKY130_FD_SC_LS__DFBBN_1%A_311_119# N_A_311_119#_M1013_s
+ N_A_311_119#_M1004_d N_A_311_119#_M1037_s N_A_311_119#_M1036_d
+ N_A_311_119#_c_1968_n N_A_311_119#_c_1952_n N_A_311_119#_c_1953_n
+ N_A_311_119#_c_1954_n N_A_311_119#_c_1955_n N_A_311_119#_c_1962_n
+ N_A_311_119#_c_1956_n N_A_311_119#_c_1963_n N_A_311_119#_c_1964_n
+ N_A_311_119#_c_1957_n N_A_311_119#_c_1958_n N_A_311_119#_c_1966_n
+ N_A_311_119#_c_1959_n N_A_311_119#_c_1960_n N_A_311_119#_c_1961_n
+ PM_SKY130_FD_SC_LS__DFBBN_1%A_311_119#
x_PM_SKY130_FD_SC_LS__DFBBN_1%Q_N N_Q_N_M1025_d N_Q_N_M1023_d N_Q_N_c_2081_n
+ N_Q_N_c_2082_n Q_N Q_N Q_N Q_N N_Q_N_c_2083_n PM_SKY130_FD_SC_LS__DFBBN_1%Q_N
x_PM_SKY130_FD_SC_LS__DFBBN_1%Q N_Q_M1009_d N_Q_M1006_d Q Q Q Q Q Q Q
+ PM_SKY130_FD_SC_LS__DFBBN_1%Q
x_PM_SKY130_FD_SC_LS__DFBBN_1%VGND N_VGND_M1033_d N_VGND_M1013_d N_VGND_M1022_d
+ N_VGND_M1038_d N_VGND_M1008_d N_VGND_M1000_d N_VGND_c_2133_n N_VGND_c_2134_n
+ N_VGND_c_2135_n N_VGND_c_2136_n N_VGND_c_2137_n N_VGND_c_2138_n VGND
+ N_VGND_c_2139_n N_VGND_c_2140_n N_VGND_c_2141_n N_VGND_c_2142_n
+ N_VGND_c_2143_n N_VGND_c_2144_n N_VGND_c_2145_n N_VGND_c_2146_n
+ N_VGND_c_2147_n N_VGND_c_2148_n N_VGND_c_2149_n N_VGND_c_2150_n
+ N_VGND_c_2151_n N_VGND_c_2152_n PM_SKY130_FD_SC_LS__DFBBN_1%VGND
x_PM_SKY130_FD_SC_LS__DFBBN_1%A_867_119# N_A_867_119#_M1016_s
+ N_A_867_119#_M1026_d N_A_867_119#_c_2265_n N_A_867_119#_c_2266_n
+ N_A_867_119#_c_2267_n N_A_867_119#_c_2268_n
+ PM_SKY130_FD_SC_LS__DFBBN_1%A_867_119#
x_PM_SKY130_FD_SC_LS__DFBBN_1%A_1818_76# N_A_1818_76#_M1014_d
+ N_A_1818_76#_M1029_d N_A_1818_76#_c_2301_n N_A_1818_76#_c_2297_n
+ N_A_1818_76#_c_2298_n PM_SKY130_FD_SC_LS__DFBBN_1%A_1818_76#
cc_1 VNB N_CLK_N_M1033_g 0.0292041f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_CLK_N_c_276_n 0.0461135f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.765
cc_3 VNB N_CLK_N_c_277_n 0.016346f $X=-0.19 $Y=-0.245 $X2=0.33 $Y2=1.465
cc_4 VNB N_D_M1013_g 0.0216814f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_5 VNB N_D_c_307_n 0.00955404f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_6 VNB D 0.00815265f $X=-0.19 $Y=-0.245 $X2=0.33 $Y2=1.465
cc_7 VNB N_D_c_309_n 0.0419609f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_474_405#_M1011_g 0.0386017f $X=-0.19 $Y=-0.245 $X2=0.33 $Y2=1.465
cc_9 VNB N_A_474_405#_M1021_g 0.0371582f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_474_405#_c_351_n 0.00822764f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_474_405#_c_352_n 0.001941f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_474_405#_c_353_n 0.00390787f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_200_74#_c_519_n 0.00800468f $X=-0.19 $Y=-0.245 $X2=0.31 $Y2=1.465
cc_14 VNB N_A_200_74#_c_520_n 0.0207162f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_200_74#_c_521_n 0.0109425f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_200_74#_c_522_n 0.00448218f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_200_74#_c_523_n 0.00350452f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_200_74#_c_524_n 0.00156732f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_200_74#_c_525_n 0.0113538f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_200_74#_c_526_n 0.00999574f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_200_74#_c_527_n 0.00789892f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_200_74#_c_528_n 0.0410328f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_200_74#_c_529_n 0.0020871f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_200_74#_c_530_n 0.0334343f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_200_74#_c_531_n 0.00271411f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_200_74#_c_532_n 0.0161806f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_200_74#_c_533_n 0.0432725f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_595_119#_c_740_n 0.0253592f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_29 VNB N_A_595_119#_c_741_n 0.00607878f $X=-0.19 $Y=-0.245 $X2=0.375
+ $Y2=1.465
cc_30 VNB N_A_595_119#_M1016_g 0.0255867f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_595_119#_c_743_n 0.012552f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_595_119#_c_744_n 0.00722226f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_595_119#_c_745_n 0.00105081f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_595_119#_c_746_n 0.00780945f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_595_119#_c_747_n 0.0276674f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_978_357#_c_848_n 0.0279397f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_37 VNB N_A_978_357#_M1026_g 0.0200752f $X=-0.19 $Y=-0.245 $X2=0.33 $Y2=1.465
cc_38 VNB N_A_978_357#_c_850_n 0.00600683f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_978_357#_c_851_n 0.0147484f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_978_357#_c_852_n 0.00469357f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_978_357#_c_853_n 0.044764f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_978_357#_c_854_n 0.00290409f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_978_357#_c_855_n 0.00330882f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_978_357#_c_856_n 0.00430743f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_978_357#_c_857_n 0.0320602f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_978_357#_c_858_n 9.45324e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_978_357#_c_859_n 0.0128172f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_978_357#_c_860_n 0.00393056f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_978_357#_c_861_n 4.53958e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_978_357#_c_862_n 0.0026653f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_978_357#_c_863_n 0.0144593f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_SET_B_c_1027_n 0.00645524f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.3
cc_53 VNB N_SET_B_M1022_g 0.0344333f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_54 VNB N_SET_B_c_1029_n 0.0354185f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_55 VNB N_SET_B_c_1030_n 0.00426394f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_SET_B_M1014_g 0.0183433f $X=-0.19 $Y=-0.245 $X2=0.31 $Y2=1.665
cc_57 VNB N_SET_B_c_1032_n 0.00175833f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_27_74#_M1034_g 0.0194417f $X=-0.19 $Y=-0.245 $X2=0.375 $Y2=1.465
cc_59 VNB N_A_27_74#_c_1158_n 0.0366106f $X=-0.19 $Y=-0.245 $X2=0.33 $Y2=1.465
cc_60 VNB N_A_27_74#_c_1159_n 0.131917f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_27_74#_c_1160_n 0.0113774f $X=-0.19 $Y=-0.245 $X2=0.31 $Y2=1.665
cc_62 VNB N_A_27_74#_M1001_g 0.047777f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_27_74#_c_1162_n 0.274447f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_27_74#_M1024_g 0.0303562f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_27_74#_c_1164_n 0.0403591f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_27_74#_c_1165_n 0.0092319f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_27_74#_c_1166_n 0.00749069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_27_74#_c_1167_n 0.0182231f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_27_74#_c_1168_n 0.0247745f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_27_74#_c_1169_n 0.00333636f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_27_74#_c_1170_n 0.00916851f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_27_74#_c_1171_n 0.00330574f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_27_74#_c_1172_n 7.77832e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_27_74#_c_1173_n 0.00267069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_1534_446#_M1038_g 0.0407631f $X=-0.19 $Y=-0.245 $X2=0.31 $Y2=1.665
cc_76 VNB N_A_1534_446#_M1025_g 0.0235282f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_1534_446#_c_1344_n 0.0485932f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_1534_446#_c_1345_n 0.0256101f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_1534_446#_c_1346_n 0.0152755f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_1534_446#_c_1347_n 0.0014249f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_1534_446#_c_1348_n 0.0197433f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_1534_446#_c_1349_n 0.028512f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_1534_446#_c_1350_n 0.00915926f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_1534_446#_c_1351_n 0.0136932f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_1534_446#_c_1352_n 0.00592654f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_1534_446#_c_1353_n 0.00271654f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_1349_114#_M1029_g 0.0297354f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_1349_114#_c_1554_n 0.0240305f $X=-0.19 $Y=-0.245 $X2=0.33
+ $Y2=1.465
cc_89 VNB N_A_1349_114#_c_1555_n 0.00203818f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_1349_114#_c_1556_n 0.00622688f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_1349_114#_c_1557_n 0.00214252f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_RESET_B_c_1703_n 0.0300381f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.3
cc_93 VNB N_RESET_B_M1008_g 0.0240606f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_94 VNB N_RESET_B_c_1705_n 0.00190844f $X=-0.19 $Y=-0.245 $X2=0.33 $Y2=1.465
cc_95 VNB N_A_2412_410#_M1009_g 0.0261447f $X=-0.19 $Y=-0.245 $X2=0.33 $Y2=1.465
cc_96 VNB N_A_2412_410#_c_1736_n 0.0616339f $X=-0.19 $Y=-0.245 $X2=0.31
+ $Y2=1.665
cc_97 VNB N_A_2412_410#_c_1737_n 0.0132214f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_A_2412_410#_c_1738_n 0.00107535f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_A_2412_410#_c_1739_n 0.00316228f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_A_2412_410#_c_1740_n 4.95953e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_VPWR_c_1792_n 0.561729f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_A_311_119#_c_1952_n 0.00190227f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_A_311_119#_c_1953_n 0.00165852f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_A_311_119#_c_1954_n 0.00763927f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_A_311_119#_c_1955_n 0.00381808f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_A_311_119#_c_1956_n 0.00475828f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_A_311_119#_c_1957_n 0.00554809f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_A_311_119#_c_1958_n 0.00226481f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_A_311_119#_c_1959_n 0.0127551f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_A_311_119#_c_1960_n 0.0115642f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_A_311_119#_c_1961_n 0.0114046f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_Q_N_c_2081_n 0.00882806f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_Q_N_c_2082_n 0.00164555f $X=-0.19 $Y=-0.245 $X2=0.31 $Y2=1.465
cc_114 VNB N_Q_N_c_2083_n 0.00232427f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB Q 0.0550644f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_116 VNB N_VGND_c_2133_n 0.00222691f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_VGND_c_2134_n 0.00951027f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_VGND_c_2135_n 0.00588277f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_VGND_c_2136_n 0.010469f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_VGND_c_2137_n 0.0159801f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_VGND_c_2138_n 0.00938486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_VGND_c_2139_n 0.0173909f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB N_VGND_c_2140_n 0.0308837f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_VGND_c_2141_n 0.0788352f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_2142_n 0.0629314f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_2143_n 0.0530939f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_VGND_c_2144_n 0.0334456f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_2145_n 0.0189533f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_2146_n 0.679646f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_2147_n 0.00501873f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_2148_n 0.00486067f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_VGND_c_2149_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_VGND_c_2150_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_VGND_c_2151_n 0.00631189f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_VGND_c_2152_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_A_867_119#_c_2265_n 0.00536288f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_A_867_119#_c_2266_n 0.016861f $X=-0.19 $Y=-0.245 $X2=0.33 $Y2=1.465
cc_138 VNB N_A_867_119#_c_2267_n 0.00260666f $X=-0.19 $Y=-0.245 $X2=0.33
+ $Y2=1.465
cc_139 VNB N_A_867_119#_c_2268_n 0.00281812f $X=-0.19 $Y=-0.245 $X2=0.31
+ $Y2=1.665
cc_140 VNB N_A_1818_76#_c_2297_n 0.00162264f $X=-0.19 $Y=-0.245 $X2=0.33
+ $Y2=1.465
cc_141 VNB N_A_1818_76#_c_2298_n 0.0108274f $X=-0.19 $Y=-0.245 $X2=0.31
+ $Y2=1.465
cc_142 VPB N_CLK_N_c_276_n 0.028884f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.765
cc_143 VPB N_CLK_N_c_277_n 0.00727431f $X=-0.19 $Y=1.66 $X2=0.33 $Y2=1.465
cc_144 VPB N_D_c_307_n 0.0390947f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_145 VPB N_D_c_311_n 0.022836f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_146 VPB N_A_474_405#_M1011_g 0.0200101f $X=-0.19 $Y=1.66 $X2=0.33 $Y2=1.465
cc_147 VPB N_A_474_405#_c_355_n 0.0497235f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_148 VPB N_A_474_405#_c_351_n 0.0511255f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_149 VPB N_A_474_405#_c_357_n 0.00180125f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_150 VPB N_A_474_405#_c_358_n 0.0223541f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_151 VPB N_A_474_405#_c_359_n 0.00131809f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_152 VPB N_A_474_405#_c_360_n 0.00509739f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_153 VPB N_A_474_405#_c_353_n 0.004099f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_154 VPB N_A_474_405#_c_362_n 0.0077751f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_155 VPB N_A_474_405#_c_363_n 0.00775337f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_156 VPB N_A_474_405#_c_364_n 0.00127831f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_157 VPB N_A_474_405#_c_365_n 0.00559253f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_158 VPB N_A_474_405#_c_366_n 0.00211414f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_159 VPB N_A_474_405#_c_367_n 4.51177e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_160 VPB N_A_200_74#_c_534_n 0.050545f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_161 VPB N_A_200_74#_c_519_n 0.0434238f $X=-0.19 $Y=1.66 $X2=0.31 $Y2=1.465
cc_162 VPB N_A_200_74#_c_536_n 0.01055f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_163 VPB N_A_200_74#_c_537_n 0.013262f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_164 VPB N_A_200_74#_c_538_n 0.00401663f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_165 VPB N_A_200_74#_c_539_n 0.00579154f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_166 VPB N_A_200_74#_c_540_n 0.0197982f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_167 VPB N_A_200_74#_c_541_n 0.00425894f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_168 VPB N_A_200_74#_c_524_n 0.00329882f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_169 VPB N_A_200_74#_c_543_n 0.00824568f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_170 VPB N_A_200_74#_c_526_n 0.00300768f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_171 VPB N_A_200_74#_c_545_n 2.50324e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_172 VPB N_A_595_119#_c_741_n 0.0153521f $X=-0.19 $Y=1.66 $X2=0.375 $Y2=1.465
cc_173 VPB N_A_595_119#_c_749_n 0.0223393f $X=-0.19 $Y=1.66 $X2=0.33 $Y2=1.465
cc_174 VPB N_A_595_119#_c_750_n 0.00552766f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_175 VPB N_A_595_119#_c_746_n 0.00925066f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_176 VPB N_A_595_119#_c_747_n 0.0137598f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_177 VPB N_A_978_357#_c_848_n 0.0489003f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_178 VPB N_A_978_357#_c_850_n 0.00819504f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_179 VPB N_A_978_357#_c_866_n 0.0232824f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_180 VPB N_A_978_357#_c_859_n 0.0061671f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_181 VPB N_A_978_357#_c_868_n 0.00377786f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_182 VPB N_A_978_357#_c_869_n 0.0019404f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_183 VPB N_A_978_357#_c_861_n 0.00225867f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_184 VPB N_SET_B_c_1027_n 0.0626085f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.3
cc_185 VPB N_SET_B_c_1030_n 0.0072325f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_186 VPB N_SET_B_c_1035_n 0.023649f $X=-0.19 $Y=1.66 $X2=0.375 $Y2=1.465
cc_187 VPB N_SET_B_c_1036_n 0.0402022f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_188 VPB N_SET_B_c_1037_n 0.00567459f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_189 VPB N_SET_B_c_1032_n 0.00578177f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_190 VPB N_A_27_74#_c_1158_n 0.0258152f $X=-0.19 $Y=1.66 $X2=0.33 $Y2=1.465
cc_191 VPB N_A_27_74#_c_1175_n 0.0382587f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_192 VPB N_A_27_74#_c_1176_n 0.00713209f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_193 VPB N_A_27_74#_c_1177_n 0.00649329f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_194 VPB N_A_27_74#_c_1178_n 0.0150721f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_195 VPB N_A_27_74#_c_1179_n 0.0219944f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_196 VPB N_A_27_74#_c_1180_n 0.00604086f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_197 VPB N_A_27_74#_c_1181_n 0.0300633f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_198 VPB N_A_27_74#_c_1182_n 0.0220152f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_199 VPB N_A_27_74#_c_1183_n 0.0135635f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_200 VPB N_A_27_74#_c_1167_n 0.00818693f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_201 VPB N_A_27_74#_c_1185_n 0.00805193f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_202 VPB N_A_27_74#_c_1186_n 0.0357063f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_203 VPB N_A_27_74#_c_1172_n 0.00276102f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_204 VPB N_A_1534_446#_c_1354_n 0.016653f $X=-0.19 $Y=1.66 $X2=0.375 $Y2=1.465
cc_205 VPB N_A_1534_446#_M1038_g 0.0251872f $X=-0.19 $Y=1.66 $X2=0.31 $Y2=1.665
cc_206 VPB N_A_1534_446#_c_1356_n 0.0206419f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_207 VPB N_A_1534_446#_c_1345_n 0.00774128f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_208 VPB N_A_1534_446#_c_1347_n 0.00790101f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_209 VPB N_A_1534_446#_c_1359_n 0.0181732f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_210 VPB N_A_1534_446#_c_1360_n 0.0269403f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_211 VPB N_A_1534_446#_c_1361_n 0.00314814f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_212 VPB N_A_1534_446#_c_1362_n 0.0773091f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_213 VPB N_A_1534_446#_c_1363_n 0.0168669f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_214 VPB N_A_1534_446#_c_1364_n 0.00164807f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_215 VPB N_A_1534_446#_c_1365_n 0.00302121f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_216 VPB N_A_1534_446#_c_1366_n 0.012225f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_217 VPB N_A_1534_446#_c_1367_n 0.0013767f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_218 VPB N_A_1534_446#_c_1368_n 0.0057012f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_219 VPB N_A_1534_446#_c_1369_n 0.00598454f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_220 VPB N_A_1349_114#_c_1554_n 0.0406877f $X=-0.19 $Y=1.66 $X2=0.33 $Y2=1.465
cc_221 VPB N_A_1349_114#_c_1559_n 0.00336771f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_222 VPB N_A_1349_114#_c_1560_n 0.0111543f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_223 VPB N_A_1349_114#_c_1561_n 0.00123654f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_224 VPB N_A_1349_114#_c_1556_n 0.00159665f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_225 VPB N_A_1349_114#_c_1563_n 0.00633533f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_226 VPB N_A_1349_114#_c_1564_n 3.23201e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_227 VPB N_A_1349_114#_c_1565_n 0.00181786f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_228 VPB N_A_1349_114#_c_1566_n 0.00795334f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_229 VPB N_A_1349_114#_c_1567_n 0.00377263f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_230 VPB N_A_1349_114#_c_1557_n 0.00227416f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_231 VPB N_A_1349_114#_c_1569_n 0.00209164f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_232 VPB N_A_1349_114#_c_1570_n 0.00228549f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_233 VPB N_A_1349_114#_c_1571_n 0.00124141f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_234 VPB N_RESET_B_c_1703_n 0.0305223f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.3
cc_235 VPB N_RESET_B_c_1705_n 0.00326259f $X=-0.19 $Y=1.66 $X2=0.33 $Y2=1.465
cc_236 VPB N_A_2412_410#_c_1741_n 0.0209332f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_237 VPB N_A_2412_410#_c_1736_n 0.00925563f $X=-0.19 $Y=1.66 $X2=0.31
+ $Y2=1.665
cc_238 VPB N_A_2412_410#_c_1738_n 0.00742978f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_239 VPB N_VPWR_c_1793_n 0.00770537f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_240 VPB N_VPWR_c_1794_n 0.00830745f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_241 VPB N_VPWR_c_1795_n 0.00339119f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_242 VPB N_VPWR_c_1796_n 0.00912283f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_243 VPB N_VPWR_c_1797_n 0.0230104f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_244 VPB N_VPWR_c_1798_n 0.0150833f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_245 VPB N_VPWR_c_1799_n 0.0366962f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_246 VPB N_VPWR_c_1800_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_247 VPB N_VPWR_c_1801_n 0.0185253f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_248 VPB N_VPWR_c_1802_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_249 VPB N_VPWR_c_1803_n 0.0197879f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_250 VPB N_VPWR_c_1804_n 0.0637933f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_251 VPB N_VPWR_c_1805_n 0.0448784f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_252 VPB N_VPWR_c_1806_n 0.0196646f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_253 VPB N_VPWR_c_1807_n 0.0477054f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_254 VPB N_VPWR_c_1808_n 0.0329211f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_255 VPB N_VPWR_c_1809_n 0.0197489f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_256 VPB N_VPWR_c_1792_n 0.186632f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_257 VPB N_VPWR_c_1811_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_258 VPB N_VPWR_c_1812_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_259 VPB N_VPWR_c_1813_n 0.0151559f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_260 VPB N_VPWR_c_1814_n 0.0139421f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_261 VPB N_VPWR_c_1815_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_262 VPB N_VPWR_c_1816_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_263 VPB N_A_311_119#_c_1962_n 0.0102675f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_264 VPB N_A_311_119#_c_1963_n 0.0126293f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_265 VPB N_A_311_119#_c_1964_n 0.00421304f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_266 VPB N_A_311_119#_c_1957_n 0.00994381f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_267 VPB N_A_311_119#_c_1966_n 0.00148905f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_268 VPB N_A_311_119#_c_1959_n 0.0148724f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_269 VPB Q_N 0.0037781f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_270 VPB Q_N 0.0154766f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_271 VPB N_Q_N_c_2083_n 0.00191248f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_272 VPB Q 0.0543585f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_273 N_CLK_N_c_276_n N_A_200_74#_c_536_n 6.23973e-19 $X=0.495 $Y=1.765 $X2=0
+ $Y2=0
cc_274 N_CLK_N_c_276_n N_A_27_74#_c_1158_n 0.0473574f $X=0.495 $Y=1.765 $X2=0
+ $Y2=0
cc_275 N_CLK_N_c_277_n N_A_27_74#_c_1158_n 2.76539e-19 $X=0.33 $Y=1.465 $X2=0
+ $Y2=0
cc_276 N_CLK_N_M1033_g N_A_27_74#_c_1160_n 0.0271107f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_277 N_CLK_N_c_276_n N_A_27_74#_c_1185_n 0.0016558f $X=0.495 $Y=1.765 $X2=0
+ $Y2=0
cc_278 N_CLK_N_c_277_n N_A_27_74#_c_1185_n 0.0249655f $X=0.33 $Y=1.465 $X2=0
+ $Y2=0
cc_279 N_CLK_N_c_276_n N_A_27_74#_c_1186_n 0.0104891f $X=0.495 $Y=1.765 $X2=0
+ $Y2=0
cc_280 N_CLK_N_M1033_g N_A_27_74#_c_1168_n 0.00159319f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_281 N_CLK_N_M1033_g N_A_27_74#_c_1169_n 0.0145993f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_282 N_CLK_N_c_276_n N_A_27_74#_c_1169_n 9.73098e-19 $X=0.495 $Y=1.765 $X2=0
+ $Y2=0
cc_283 N_CLK_N_c_277_n N_A_27_74#_c_1169_n 0.00971403f $X=0.33 $Y=1.465 $X2=0
+ $Y2=0
cc_284 N_CLK_N_c_276_n N_A_27_74#_c_1170_n 0.00158295f $X=0.495 $Y=1.765 $X2=0
+ $Y2=0
cc_285 N_CLK_N_c_277_n N_A_27_74#_c_1170_n 0.0209549f $X=0.33 $Y=1.465 $X2=0
+ $Y2=0
cc_286 N_CLK_N_c_276_n N_A_27_74#_c_1200_n 0.0139266f $X=0.495 $Y=1.765 $X2=0
+ $Y2=0
cc_287 N_CLK_N_c_277_n N_A_27_74#_c_1200_n 0.00433199f $X=0.33 $Y=1.465 $X2=0
+ $Y2=0
cc_288 N_CLK_N_M1033_g N_A_27_74#_c_1171_n 0.00383463f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_289 N_CLK_N_c_276_n N_A_27_74#_c_1172_n 0.00487653f $X=0.495 $Y=1.765 $X2=0
+ $Y2=0
cc_290 N_CLK_N_c_277_n N_A_27_74#_c_1172_n 0.0113335f $X=0.33 $Y=1.465 $X2=0
+ $Y2=0
cc_291 N_CLK_N_c_276_n N_A_27_74#_c_1173_n 0.00233952f $X=0.495 $Y=1.765 $X2=0
+ $Y2=0
cc_292 N_CLK_N_c_277_n N_A_27_74#_c_1173_n 0.0267562f $X=0.33 $Y=1.465 $X2=0
+ $Y2=0
cc_293 N_CLK_N_c_276_n N_VPWR_c_1793_n 0.00486623f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_294 N_CLK_N_c_276_n N_VPWR_c_1803_n 0.00445602f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_295 N_CLK_N_c_276_n N_VPWR_c_1792_n 0.00861134f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_296 N_CLK_N_M1033_g N_VGND_c_2133_n 0.0125189f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_297 N_CLK_N_M1033_g N_VGND_c_2139_n 0.00383152f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_298 N_CLK_N_M1033_g N_VGND_c_2146_n 0.00761198f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_299 N_D_M1013_g N_A_474_405#_M1011_g 0.0157832f $X=1.915 $Y=0.805 $X2=0 $Y2=0
cc_300 N_D_c_307_n N_A_474_405#_M1011_g 0.0174461f $X=2.01 $Y=2.35 $X2=0 $Y2=0
cc_301 D N_A_474_405#_M1011_g 0.013583f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_302 N_D_c_309_n N_A_474_405#_M1011_g 0.0213648f $X=2.09 $Y=1.345 $X2=0 $Y2=0
cc_303 N_D_c_307_n N_A_474_405#_c_355_n 0.0156185f $X=2.01 $Y=2.35 $X2=0 $Y2=0
cc_304 N_D_c_311_n N_A_474_405#_c_355_n 0.0114171f $X=2.01 $Y=2.44 $X2=0 $Y2=0
cc_305 N_D_c_311_n N_A_474_405#_c_357_n 2.49669e-19 $X=2.01 $Y=2.44 $X2=0 $Y2=0
cc_306 N_D_c_307_n N_A_474_405#_c_365_n 4.06248e-19 $X=2.01 $Y=2.35 $X2=0 $Y2=0
cc_307 N_D_c_311_n N_A_200_74#_c_536_n 0.00308482f $X=2.01 $Y=2.44 $X2=0 $Y2=0
cc_308 N_D_M1013_g N_A_200_74#_c_521_n 0.00280927f $X=1.915 $Y=0.805 $X2=0 $Y2=0
cc_309 N_D_c_311_n N_A_200_74#_c_537_n 0.0102153f $X=2.01 $Y=2.44 $X2=0 $Y2=0
cc_310 N_D_c_307_n N_A_200_74#_c_539_n 0.0120338f $X=2.01 $Y=2.35 $X2=0 $Y2=0
cc_311 N_D_c_311_n N_A_200_74#_c_539_n 0.0159117f $X=2.01 $Y=2.44 $X2=0 $Y2=0
cc_312 D N_A_200_74#_c_540_n 0.0471758f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_313 N_D_c_309_n N_A_200_74#_c_540_n 0.00290311f $X=2.09 $Y=1.345 $X2=0 $Y2=0
cc_314 N_D_c_307_n N_A_200_74#_c_554_n 0.00803175f $X=2.01 $Y=2.35 $X2=0 $Y2=0
cc_315 D N_A_200_74#_c_554_n 0.0133696f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_316 N_D_c_309_n N_A_200_74#_c_554_n 5.80967e-19 $X=2.09 $Y=1.345 $X2=0 $Y2=0
cc_317 D N_A_200_74#_c_522_n 0.00391807f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_318 D N_A_200_74#_c_558_n 0.00187865f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_319 D N_A_200_74#_c_531_n 0.0155335f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_320 N_D_c_309_n N_A_27_74#_c_1158_n 0.00190331f $X=2.09 $Y=1.345 $X2=0 $Y2=0
cc_321 N_D_M1013_g N_A_27_74#_c_1159_n 0.00999521f $X=1.915 $Y=0.805 $X2=0 $Y2=0
cc_322 D N_A_27_74#_M1001_g 0.00260483f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_323 N_D_c_311_n N_VPWR_c_1794_n 0.00177809f $X=2.01 $Y=2.44 $X2=0 $Y2=0
cc_324 N_D_c_311_n N_VPWR_c_1799_n 9.62598e-19 $X=2.01 $Y=2.44 $X2=0 $Y2=0
cc_325 N_D_M1013_g N_A_311_119#_c_1968_n 0.0100459f $X=1.915 $Y=0.805 $X2=0
+ $Y2=0
cc_326 D N_A_311_119#_c_1968_n 0.056469f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_327 N_D_c_309_n N_A_311_119#_c_1968_n 0.00624979f $X=2.09 $Y=1.345 $X2=0
+ $Y2=0
cc_328 N_D_M1013_g N_A_311_119#_c_1952_n 8.06126e-19 $X=1.915 $Y=0.805 $X2=0
+ $Y2=0
cc_329 N_D_M1013_g N_A_311_119#_c_1958_n 0.00774165f $X=1.915 $Y=0.805 $X2=0
+ $Y2=0
cc_330 N_D_c_311_n N_A_311_119#_c_1966_n 0.0065017f $X=2.01 $Y=2.44 $X2=0 $Y2=0
cc_331 N_D_M1013_g N_A_311_119#_c_1959_n 0.0122916f $X=1.915 $Y=0.805 $X2=0
+ $Y2=0
cc_332 N_D_c_307_n N_A_311_119#_c_1959_n 0.0207136f $X=2.01 $Y=2.35 $X2=0 $Y2=0
cc_333 D N_A_311_119#_c_1959_n 0.0262098f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_334 N_D_M1013_g N_VGND_c_2134_n 0.00252054f $X=1.915 $Y=0.805 $X2=0 $Y2=0
cc_335 N_D_M1013_g N_VGND_c_2146_n 9.39239e-19 $X=1.915 $Y=0.805 $X2=0 $Y2=0
cc_336 N_A_474_405#_c_355_n N_A_200_74#_c_534_n 0.051967f $X=2.61 $Y=2.44 $X2=0
+ $Y2=0
cc_337 N_A_474_405#_c_357_n N_A_200_74#_c_534_n 0.00692726f $X=2.72 $Y=2.905
+ $X2=0 $Y2=0
cc_338 N_A_474_405#_c_358_n N_A_200_74#_c_534_n 0.0125015f $X=4.2 $Y=2.99 $X2=0
+ $Y2=0
cc_339 N_A_474_405#_c_365_n N_A_200_74#_c_534_n 0.00217001f $X=2.72 $Y=2.19
+ $X2=0 $Y2=0
cc_340 N_A_474_405#_M1021_g N_A_200_74#_c_519_n 8.87914e-19 $X=6.195 $Y=0.87
+ $X2=0 $Y2=0
cc_341 N_A_474_405#_c_351_n N_A_200_74#_c_519_n 0.0792398f $X=6.41 $Y=2.045
+ $X2=0 $Y2=0
cc_342 N_A_474_405#_c_363_n N_A_200_74#_c_519_n 5.57726e-19 $X=6.12 $Y=2.405
+ $X2=0 $Y2=0
cc_343 N_A_474_405#_c_364_n N_A_200_74#_c_519_n 0.00308463f $X=6.285 $Y=1.795
+ $X2=0 $Y2=0
cc_344 N_A_474_405#_M1011_g N_A_200_74#_c_539_n 0.00296524f $X=2.54 $Y=0.805
+ $X2=0 $Y2=0
cc_345 N_A_474_405#_c_355_n N_A_200_74#_c_539_n 0.00225238f $X=2.61 $Y=2.44
+ $X2=0 $Y2=0
cc_346 N_A_474_405#_c_357_n N_A_200_74#_c_539_n 0.00512815f $X=2.72 $Y=2.905
+ $X2=0 $Y2=0
cc_347 N_A_474_405#_c_365_n N_A_200_74#_c_539_n 0.0192184f $X=2.72 $Y=2.19 $X2=0
+ $Y2=0
cc_348 N_A_474_405#_M1011_g N_A_200_74#_c_540_n 0.0109769f $X=2.54 $Y=0.805
+ $X2=0 $Y2=0
cc_349 N_A_474_405#_c_355_n N_A_200_74#_c_540_n 0.00432778f $X=2.61 $Y=2.44
+ $X2=0 $Y2=0
cc_350 N_A_474_405#_c_365_n N_A_200_74#_c_540_n 0.0325651f $X=2.72 $Y=2.19 $X2=0
+ $Y2=0
cc_351 N_A_474_405#_M1011_g N_A_200_74#_c_522_n 0.00178535f $X=2.54 $Y=0.805
+ $X2=0 $Y2=0
cc_352 N_A_474_405#_M1011_g N_A_200_74#_c_541_n 0.00498597f $X=2.54 $Y=0.805
+ $X2=0 $Y2=0
cc_353 N_A_474_405#_c_355_n N_A_200_74#_c_541_n 3.0079e-19 $X=2.61 $Y=2.44 $X2=0
+ $Y2=0
cc_354 N_A_474_405#_c_358_n N_A_200_74#_c_541_n 0.00330156f $X=4.2 $Y=2.99 $X2=0
+ $Y2=0
cc_355 N_A_474_405#_c_365_n N_A_200_74#_c_541_n 0.0262565f $X=2.72 $Y=2.19 $X2=0
+ $Y2=0
cc_356 N_A_474_405#_M1021_g N_A_200_74#_c_523_n 0.00260546f $X=6.195 $Y=0.87
+ $X2=0 $Y2=0
cc_357 N_A_474_405#_M1021_g N_A_200_74#_c_524_n 0.00127909f $X=6.195 $Y=0.87
+ $X2=0 $Y2=0
cc_358 N_A_474_405#_c_351_n N_A_200_74#_c_524_n 0.00127078f $X=6.41 $Y=2.045
+ $X2=0 $Y2=0
cc_359 N_A_474_405#_c_364_n N_A_200_74#_c_524_n 0.0137339f $X=6.285 $Y=1.795
+ $X2=0 $Y2=0
cc_360 N_A_474_405#_M1021_g N_A_200_74#_c_528_n 0.00706397f $X=6.195 $Y=0.87
+ $X2=0 $Y2=0
cc_361 N_A_474_405#_c_351_n N_A_200_74#_c_528_n 3.56533e-19 $X=6.41 $Y=2.045
+ $X2=0 $Y2=0
cc_362 N_A_474_405#_c_352_n N_A_200_74#_c_528_n 0.0141949f $X=4.73 $Y=1.165
+ $X2=0 $Y2=0
cc_363 N_A_474_405#_c_353_n N_A_200_74#_c_528_n 0.0246337f $X=4.73 $Y=2.305
+ $X2=0 $Y2=0
cc_364 N_A_474_405#_c_364_n N_A_200_74#_c_528_n 0.00188756f $X=6.285 $Y=1.795
+ $X2=0 $Y2=0
cc_365 N_A_474_405#_M1011_g N_A_200_74#_c_531_n 6.10356e-19 $X=2.54 $Y=0.805
+ $X2=0 $Y2=0
cc_366 N_A_474_405#_c_358_n N_A_595_119#_M1035_d 0.00254113f $X=4.2 $Y=2.99
+ $X2=0 $Y2=0
cc_367 N_A_474_405#_c_353_n N_A_595_119#_c_741_n 0.00757396f $X=4.73 $Y=2.305
+ $X2=0 $Y2=0
cc_368 N_A_474_405#_c_358_n N_A_595_119#_c_749_n 0.00559477f $X=4.2 $Y=2.99
+ $X2=0 $Y2=0
cc_369 N_A_474_405#_c_360_n N_A_595_119#_c_749_n 0.00759862f $X=4.365 $Y=2.905
+ $X2=0 $Y2=0
cc_370 N_A_474_405#_c_353_n N_A_595_119#_c_749_n 0.00817868f $X=4.73 $Y=2.305
+ $X2=0 $Y2=0
cc_371 N_A_474_405#_c_366_n N_A_595_119#_c_749_n 0.0134914f $X=4.815 $Y=2.397
+ $X2=0 $Y2=0
cc_372 N_A_474_405#_c_352_n N_A_595_119#_M1016_g 0.00833041f $X=4.73 $Y=1.165
+ $X2=0 $Y2=0
cc_373 N_A_474_405#_c_353_n N_A_595_119#_M1016_g 0.00448696f $X=4.73 $Y=2.305
+ $X2=0 $Y2=0
cc_374 N_A_474_405#_c_353_n N_A_595_119#_c_743_n 0.00646074f $X=4.73 $Y=2.305
+ $X2=0 $Y2=0
cc_375 N_A_474_405#_c_357_n N_A_595_119#_c_762_n 0.00862753f $X=2.72 $Y=2.905
+ $X2=0 $Y2=0
cc_376 N_A_474_405#_c_358_n N_A_595_119#_c_762_n 0.0258603f $X=4.2 $Y=2.99 $X2=0
+ $Y2=0
cc_377 N_A_474_405#_c_357_n N_A_595_119#_c_750_n 0.00561291f $X=2.72 $Y=2.905
+ $X2=0 $Y2=0
cc_378 N_A_474_405#_M1011_g N_A_595_119#_c_745_n 2.98275e-19 $X=2.54 $Y=0.805
+ $X2=0 $Y2=0
cc_379 N_A_474_405#_c_358_n N_A_978_357#_c_848_n 4.73984e-19 $X=4.2 $Y=2.99
+ $X2=0 $Y2=0
cc_380 N_A_474_405#_c_360_n N_A_978_357#_c_848_n 0.00151152f $X=4.365 $Y=2.905
+ $X2=0 $Y2=0
cc_381 N_A_474_405#_c_352_n N_A_978_357#_c_848_n 0.00378209f $X=4.73 $Y=1.165
+ $X2=0 $Y2=0
cc_382 N_A_474_405#_c_353_n N_A_978_357#_c_848_n 0.010802f $X=4.73 $Y=2.305
+ $X2=0 $Y2=0
cc_383 N_A_474_405#_c_423_p N_A_978_357#_c_848_n 0.017662f $X=5.57 $Y=2.405
+ $X2=0 $Y2=0
cc_384 N_A_474_405#_c_366_n N_A_978_357#_c_848_n 4.04324e-19 $X=4.815 $Y=2.397
+ $X2=0 $Y2=0
cc_385 N_A_474_405#_c_352_n N_A_978_357#_M1026_g 0.00781472f $X=4.73 $Y=1.165
+ $X2=0 $Y2=0
cc_386 N_A_474_405#_c_353_n N_A_978_357#_M1026_g 0.00250793f $X=4.73 $Y=2.305
+ $X2=0 $Y2=0
cc_387 N_A_474_405#_M1021_g N_A_978_357#_c_851_n 0.0131218f $X=6.195 $Y=0.87
+ $X2=0 $Y2=0
cc_388 N_A_474_405#_c_351_n N_A_978_357#_c_851_n 0.00667283f $X=6.41 $Y=2.045
+ $X2=0 $Y2=0
cc_389 N_A_474_405#_c_364_n N_A_978_357#_c_851_n 0.0239932f $X=6.285 $Y=1.795
+ $X2=0 $Y2=0
cc_390 N_A_474_405#_M1021_g N_A_978_357#_c_852_n 0.00762346f $X=6.195 $Y=0.87
+ $X2=0 $Y2=0
cc_391 N_A_474_405#_M1021_g N_A_978_357#_c_854_n 3.98045e-19 $X=6.195 $Y=0.87
+ $X2=0 $Y2=0
cc_392 N_A_474_405#_c_352_n N_A_978_357#_c_861_n 0.0106525f $X=4.73 $Y=1.165
+ $X2=0 $Y2=0
cc_393 N_A_474_405#_c_353_n N_A_978_357#_c_861_n 0.0243026f $X=4.73 $Y=2.305
+ $X2=0 $Y2=0
cc_394 N_A_474_405#_c_423_p N_A_978_357#_c_861_n 0.00615851f $X=5.57 $Y=2.405
+ $X2=0 $Y2=0
cc_395 N_A_474_405#_c_351_n N_SET_B_c_1027_n 0.017588f $X=6.41 $Y=2.045
+ $X2=-0.19 $Y2=-0.245
cc_396 N_A_474_405#_c_423_p N_SET_B_c_1027_n 0.0105328f $X=5.57 $Y=2.405
+ $X2=-0.19 $Y2=-0.245
cc_397 N_A_474_405#_c_362_n N_SET_B_c_1027_n 0.00545193f $X=5.655 $Y=2.815
+ $X2=-0.19 $Y2=-0.245
cc_398 N_A_474_405#_c_363_n N_SET_B_c_1027_n 4.6316e-19 $X=6.12 $Y=2.405
+ $X2=-0.19 $Y2=-0.245
cc_399 N_A_474_405#_c_364_n N_SET_B_c_1027_n 0.00415719f $X=6.285 $Y=1.795
+ $X2=-0.19 $Y2=-0.245
cc_400 N_A_474_405#_c_367_n N_SET_B_c_1027_n 0.00361799f $X=5.655 $Y=2.405
+ $X2=-0.19 $Y2=-0.245
cc_401 N_A_474_405#_M1021_g N_SET_B_M1022_g 0.0322389f $X=6.195 $Y=0.87 $X2=0
+ $Y2=0
cc_402 N_A_474_405#_c_352_n N_SET_B_M1022_g 5.41739e-19 $X=4.73 $Y=1.165 $X2=0
+ $Y2=0
cc_403 N_A_474_405#_c_351_n N_SET_B_c_1036_n 0.0033232f $X=6.41 $Y=2.045 $X2=0
+ $Y2=0
cc_404 N_A_474_405#_c_363_n N_SET_B_c_1036_n 0.0124917f $X=6.12 $Y=2.405 $X2=0
+ $Y2=0
cc_405 N_A_474_405#_c_364_n N_SET_B_c_1036_n 0.026357f $X=6.285 $Y=1.795 $X2=0
+ $Y2=0
cc_406 N_A_474_405#_c_367_n N_SET_B_c_1036_n 0.00435015f $X=5.655 $Y=2.405 $X2=0
+ $Y2=0
cc_407 N_A_474_405#_M1027_d N_SET_B_c_1051_n 0.00121073f $X=5.505 $Y=2.12 $X2=0
+ $Y2=0
cc_408 N_A_474_405#_c_353_n N_SET_B_c_1051_n 0.00473289f $X=4.73 $Y=2.305 $X2=0
+ $Y2=0
cc_409 N_A_474_405#_c_423_p N_SET_B_c_1051_n 0.00339938f $X=5.57 $Y=2.405 $X2=0
+ $Y2=0
cc_410 N_A_474_405#_c_364_n N_SET_B_c_1051_n 0.00140895f $X=6.285 $Y=1.795 $X2=0
+ $Y2=0
cc_411 N_A_474_405#_c_367_n N_SET_B_c_1051_n 0.00151694f $X=5.655 $Y=2.405 $X2=0
+ $Y2=0
cc_412 N_A_474_405#_M1027_d N_SET_B_c_1037_n 6.75624e-19 $X=5.505 $Y=2.12 $X2=0
+ $Y2=0
cc_413 N_A_474_405#_c_351_n N_SET_B_c_1037_n 0.00156685f $X=6.41 $Y=2.045 $X2=0
+ $Y2=0
cc_414 N_A_474_405#_c_353_n N_SET_B_c_1037_n 0.0108049f $X=4.73 $Y=2.305 $X2=0
+ $Y2=0
cc_415 N_A_474_405#_c_423_p N_SET_B_c_1037_n 0.00574959f $X=5.57 $Y=2.405 $X2=0
+ $Y2=0
cc_416 N_A_474_405#_c_363_n N_SET_B_c_1037_n 6.76383e-19 $X=6.12 $Y=2.405 $X2=0
+ $Y2=0
cc_417 N_A_474_405#_c_364_n N_SET_B_c_1037_n 0.0190661f $X=6.285 $Y=1.795 $X2=0
+ $Y2=0
cc_418 N_A_474_405#_c_367_n N_SET_B_c_1037_n 0.00940548f $X=5.655 $Y=2.405 $X2=0
+ $Y2=0
cc_419 N_A_474_405#_M1011_g N_A_27_74#_c_1159_n 0.00997995f $X=2.54 $Y=0.805
+ $X2=0 $Y2=0
cc_420 N_A_474_405#_M1011_g N_A_27_74#_M1001_g 0.0820849f $X=2.54 $Y=0.805 $X2=0
+ $Y2=0
cc_421 N_A_474_405#_M1021_g N_A_27_74#_c_1162_n 0.0103107f $X=6.195 $Y=0.87
+ $X2=0 $Y2=0
cc_422 N_A_474_405#_c_358_n N_A_27_74#_c_1179_n 0.0135343f $X=4.2 $Y=2.99 $X2=0
+ $Y2=0
cc_423 N_A_474_405#_c_360_n N_A_27_74#_c_1179_n 0.00442678f $X=4.365 $Y=2.905
+ $X2=0 $Y2=0
cc_424 N_A_474_405#_M1021_g N_A_27_74#_M1024_g 0.0270157f $X=6.195 $Y=0.87 $X2=0
+ $Y2=0
cc_425 N_A_474_405#_c_351_n N_A_1349_114#_c_1569_n 0.00274738f $X=6.41 $Y=2.045
+ $X2=0 $Y2=0
cc_426 N_A_474_405#_c_363_n N_A_1349_114#_c_1569_n 0.00689203f $X=6.12 $Y=2.405
+ $X2=0 $Y2=0
cc_427 N_A_474_405#_c_364_n N_A_1349_114#_c_1569_n 0.00834957f $X=6.285 $Y=1.795
+ $X2=0 $Y2=0
cc_428 N_A_474_405#_c_423_p N_VPWR_M1020_d 0.00527285f $X=5.57 $Y=2.405 $X2=0
+ $Y2=0
cc_429 N_A_474_405#_c_363_n N_VPWR_M1017_s 0.00417768f $X=6.12 $Y=2.405 $X2=0
+ $Y2=0
cc_430 N_A_474_405#_c_364_n N_VPWR_M1017_s 0.00382512f $X=6.285 $Y=1.795 $X2=0
+ $Y2=0
cc_431 N_A_474_405#_c_355_n N_VPWR_c_1794_n 0.00455817f $X=2.61 $Y=2.44 $X2=0
+ $Y2=0
cc_432 N_A_474_405#_c_357_n N_VPWR_c_1794_n 0.0266437f $X=2.72 $Y=2.905 $X2=0
+ $Y2=0
cc_433 N_A_474_405#_c_359_n N_VPWR_c_1794_n 0.0135904f $X=2.805 $Y=2.99 $X2=0
+ $Y2=0
cc_434 N_A_474_405#_c_365_n N_VPWR_c_1794_n 0.00776258f $X=2.72 $Y=2.19 $X2=0
+ $Y2=0
cc_435 N_A_474_405#_c_358_n N_VPWR_c_1795_n 0.00551498f $X=4.2 $Y=2.99 $X2=0
+ $Y2=0
cc_436 N_A_474_405#_c_360_n N_VPWR_c_1795_n 0.00747936f $X=4.365 $Y=2.905 $X2=0
+ $Y2=0
cc_437 N_A_474_405#_c_423_p N_VPWR_c_1795_n 0.0168032f $X=5.57 $Y=2.405 $X2=0
+ $Y2=0
cc_438 N_A_474_405#_c_362_n N_VPWR_c_1795_n 0.0214859f $X=5.655 $Y=2.815 $X2=0
+ $Y2=0
cc_439 N_A_474_405#_c_351_n N_VPWR_c_1796_n 0.0106984f $X=6.41 $Y=2.045 $X2=0
+ $Y2=0
cc_440 N_A_474_405#_c_362_n N_VPWR_c_1796_n 0.0232837f $X=5.655 $Y=2.815 $X2=0
+ $Y2=0
cc_441 N_A_474_405#_c_363_n N_VPWR_c_1796_n 0.0222325f $X=6.12 $Y=2.405 $X2=0
+ $Y2=0
cc_442 N_A_474_405#_c_362_n N_VPWR_c_1801_n 0.0110419f $X=5.655 $Y=2.815 $X2=0
+ $Y2=0
cc_443 N_A_474_405#_c_355_n N_VPWR_c_1804_n 0.00404572f $X=2.61 $Y=2.44 $X2=0
+ $Y2=0
cc_444 N_A_474_405#_c_358_n N_VPWR_c_1804_n 0.113144f $X=4.2 $Y=2.99 $X2=0 $Y2=0
cc_445 N_A_474_405#_c_359_n N_VPWR_c_1804_n 0.0122392f $X=2.805 $Y=2.99 $X2=0
+ $Y2=0
cc_446 N_A_474_405#_c_351_n N_VPWR_c_1805_n 0.00413917f $X=6.41 $Y=2.045 $X2=0
+ $Y2=0
cc_447 N_A_474_405#_c_355_n N_VPWR_c_1792_n 0.00358569f $X=2.61 $Y=2.44 $X2=0
+ $Y2=0
cc_448 N_A_474_405#_c_351_n N_VPWR_c_1792_n 0.0051762f $X=6.41 $Y=2.045 $X2=0
+ $Y2=0
cc_449 N_A_474_405#_c_358_n N_VPWR_c_1792_n 0.065152f $X=4.2 $Y=2.99 $X2=0 $Y2=0
cc_450 N_A_474_405#_c_359_n N_VPWR_c_1792_n 0.00661913f $X=2.805 $Y=2.99 $X2=0
+ $Y2=0
cc_451 N_A_474_405#_c_423_p N_VPWR_c_1792_n 0.00697113f $X=5.57 $Y=2.405 $X2=0
+ $Y2=0
cc_452 N_A_474_405#_c_362_n N_VPWR_c_1792_n 0.00915013f $X=5.655 $Y=2.815 $X2=0
+ $Y2=0
cc_453 N_A_474_405#_c_363_n N_VPWR_c_1792_n 0.0112609f $X=6.12 $Y=2.405 $X2=0
+ $Y2=0
cc_454 N_A_474_405#_c_366_n N_VPWR_c_1792_n 0.0157857f $X=4.815 $Y=2.397 $X2=0
+ $Y2=0
cc_455 N_A_474_405#_c_358_n N_A_311_119#_M1036_d 0.00556203f $X=4.2 $Y=2.99
+ $X2=0 $Y2=0
cc_456 N_A_474_405#_M1011_g N_A_311_119#_c_1968_n 0.00932917f $X=2.54 $Y=0.805
+ $X2=0 $Y2=0
cc_457 N_A_474_405#_M1011_g N_A_311_119#_c_1952_n 0.00804248f $X=2.54 $Y=0.805
+ $X2=0 $Y2=0
cc_458 N_A_474_405#_c_358_n N_A_311_119#_c_1962_n 0.0189745f $X=4.2 $Y=2.99
+ $X2=0 $Y2=0
cc_459 N_A_474_405#_c_360_n N_A_311_119#_c_1962_n 0.0178267f $X=4.365 $Y=2.905
+ $X2=0 $Y2=0
cc_460 N_A_474_405#_c_353_n N_A_311_119#_c_1962_n 0.00455445f $X=4.73 $Y=2.305
+ $X2=0 $Y2=0
cc_461 N_A_474_405#_c_366_n N_A_311_119#_c_1962_n 0.0141437f $X=4.815 $Y=2.397
+ $X2=0 $Y2=0
cc_462 N_A_474_405#_M1019_s N_A_311_119#_c_1963_n 0.0025523f $X=4.235 $Y=2.12
+ $X2=0 $Y2=0
cc_463 N_A_474_405#_c_353_n N_A_311_119#_c_1963_n 0.012934f $X=4.73 $Y=2.305
+ $X2=0 $Y2=0
cc_464 N_A_474_405#_c_366_n N_A_311_119#_c_1963_n 0.0202522f $X=4.815 $Y=2.397
+ $X2=0 $Y2=0
cc_465 N_A_474_405#_c_353_n N_A_311_119#_c_1957_n 0.0559469f $X=4.73 $Y=2.305
+ $X2=0 $Y2=0
cc_466 N_A_474_405#_M1011_g N_A_311_119#_c_1958_n 8.52988e-19 $X=2.54 $Y=0.805
+ $X2=0 $Y2=0
cc_467 N_A_474_405#_c_352_n N_A_311_119#_c_1961_n 0.0140524f $X=4.73 $Y=1.165
+ $X2=0 $Y2=0
cc_468 N_A_474_405#_c_357_n A_537_503# 0.00435802f $X=2.72 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_469 N_A_474_405#_c_358_n A_537_503# 0.00351031f $X=4.2 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_470 N_A_474_405#_c_353_n A_933_424# 0.00239212f $X=4.73 $Y=2.305 $X2=-0.19
+ $Y2=-0.245
cc_471 N_A_474_405#_c_423_p A_933_424# 0.00186433f $X=5.57 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_472 N_A_474_405#_c_366_n A_933_424# 0.00232236f $X=4.815 $Y=2.397 $X2=-0.19
+ $Y2=-0.245
cc_473 N_A_474_405#_M1011_g N_VGND_c_2134_n 0.00177627f $X=2.54 $Y=0.805 $X2=0
+ $Y2=0
cc_474 N_A_474_405#_M1021_g N_VGND_c_2135_n 0.00898422f $X=6.195 $Y=0.87 $X2=0
+ $Y2=0
cc_475 N_A_474_405#_M1011_g N_VGND_c_2146_n 7.22543e-19 $X=2.54 $Y=0.805 $X2=0
+ $Y2=0
cc_476 N_A_474_405#_M1021_g N_VGND_c_2146_n 7.88961e-19 $X=6.195 $Y=0.87 $X2=0
+ $Y2=0
cc_477 N_A_474_405#_c_352_n N_A_867_119#_c_2266_n 0.0189518f $X=4.73 $Y=1.165
+ $X2=0 $Y2=0
cc_478 N_A_474_405#_M1021_g N_A_867_119#_c_2268_n 2.31893e-19 $X=6.195 $Y=0.87
+ $X2=0 $Y2=0
cc_479 N_A_200_74#_c_528_n N_A_595_119#_M1016_g 0.00360788f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_480 N_A_200_74#_c_534_n N_A_595_119#_c_762_n 0.00312608f $X=3.03 $Y=2.44
+ $X2=0 $Y2=0
cc_481 N_A_200_74#_c_541_n N_A_595_119#_c_762_n 0.00809752f $X=3.075 $Y=2.19
+ $X2=0 $Y2=0
cc_482 N_A_200_74#_c_528_n N_A_595_119#_c_769_n 0.00566444f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_483 N_A_200_74#_c_530_n N_A_595_119#_c_769_n 0.00258703f $X=3.35 $Y=1.29
+ $X2=0 $Y2=0
cc_484 N_A_200_74#_c_531_n N_A_595_119#_c_769_n 0.010638f $X=3.35 $Y=1.29 $X2=0
+ $Y2=0
cc_485 N_A_200_74#_c_532_n N_A_595_119#_c_769_n 0.00975616f $X=3.35 $Y=1.125
+ $X2=0 $Y2=0
cc_486 N_A_200_74#_c_534_n N_A_595_119#_c_750_n 0.00308573f $X=3.03 $Y=2.44
+ $X2=0 $Y2=0
cc_487 N_A_200_74#_c_541_n N_A_595_119#_c_750_n 0.0375973f $X=3.075 $Y=2.19
+ $X2=0 $Y2=0
cc_488 N_A_200_74#_c_545_n N_A_595_119#_c_750_n 0.00486726f $X=3.107 $Y=1.77
+ $X2=0 $Y2=0
cc_489 N_A_200_74#_c_528_n N_A_595_119#_c_744_n 0.0170584f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_490 N_A_200_74#_c_558_n N_A_595_119#_c_744_n 3.53962e-19 $X=3.265 $Y=1.295
+ $X2=0 $Y2=0
cc_491 N_A_200_74#_c_530_n N_A_595_119#_c_744_n 0.00564507f $X=3.35 $Y=1.29
+ $X2=0 $Y2=0
cc_492 N_A_200_74#_c_531_n N_A_595_119#_c_744_n 0.0192812f $X=3.35 $Y=1.29 $X2=0
+ $Y2=0
cc_493 N_A_200_74#_c_532_n N_A_595_119#_c_744_n 0.00542458f $X=3.35 $Y=1.125
+ $X2=0 $Y2=0
cc_494 N_A_200_74#_c_558_n N_A_595_119#_c_745_n 0.00201621f $X=3.265 $Y=1.295
+ $X2=0 $Y2=0
cc_495 N_A_200_74#_c_530_n N_A_595_119#_c_745_n 0.00145122f $X=3.35 $Y=1.29
+ $X2=0 $Y2=0
cc_496 N_A_200_74#_c_531_n N_A_595_119#_c_745_n 0.0187186f $X=3.35 $Y=1.29 $X2=0
+ $Y2=0
cc_497 N_A_200_74#_c_532_n N_A_595_119#_c_745_n 0.00905142f $X=3.35 $Y=1.125
+ $X2=0 $Y2=0
cc_498 N_A_200_74#_c_522_n N_A_595_119#_c_746_n 0.0130684f $X=3.107 $Y=1.685
+ $X2=0 $Y2=0
cc_499 N_A_200_74#_c_545_n N_A_595_119#_c_746_n 0.0093116f $X=3.107 $Y=1.77
+ $X2=0 $Y2=0
cc_500 N_A_200_74#_c_528_n N_A_595_119#_c_746_n 0.0194182f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_501 N_A_200_74#_c_530_n N_A_595_119#_c_746_n 0.00147136f $X=3.35 $Y=1.29
+ $X2=0 $Y2=0
cc_502 N_A_200_74#_c_531_n N_A_595_119#_c_746_n 0.00918903f $X=3.35 $Y=1.29
+ $X2=0 $Y2=0
cc_503 N_A_200_74#_c_522_n N_A_595_119#_c_747_n 9.08222e-19 $X=3.107 $Y=1.685
+ $X2=0 $Y2=0
cc_504 N_A_200_74#_c_528_n N_A_595_119#_c_747_n 0.00815023f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_505 N_A_200_74#_c_530_n N_A_595_119#_c_747_n 0.00239727f $X=3.35 $Y=1.29
+ $X2=0 $Y2=0
cc_506 N_A_200_74#_c_528_n N_A_978_357#_c_848_n 0.00428585f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_507 N_A_200_74#_c_528_n N_A_978_357#_M1026_g 0.00705248f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_508 N_A_200_74#_c_523_n N_A_978_357#_c_851_n 0.0120591f $X=6.892 $Y=1.56
+ $X2=0 $Y2=0
cc_509 N_A_200_74#_c_528_n N_A_978_357#_c_851_n 0.045746f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_510 N_A_200_74#_c_529_n N_A_978_357#_c_851_n 2.99413e-19 $X=6.96 $Y=1.295
+ $X2=0 $Y2=0
cc_511 N_A_200_74#_c_523_n N_A_978_357#_c_852_n 0.00817666f $X=6.892 $Y=1.56
+ $X2=0 $Y2=0
cc_512 N_A_200_74#_c_528_n N_A_978_357#_c_852_n 0.0161182f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_513 N_A_200_74#_c_529_n N_A_978_357#_c_852_n 2.5995e-19 $X=6.96 $Y=1.295
+ $X2=0 $Y2=0
cc_514 N_A_200_74#_c_520_n N_A_978_357#_c_853_n 0.00449896f $X=7.98 $Y=1.23
+ $X2=0 $Y2=0
cc_515 N_A_200_74#_c_523_n N_A_978_357#_c_853_n 2.41257e-19 $X=6.892 $Y=1.56
+ $X2=0 $Y2=0
cc_516 N_A_200_74#_c_520_n N_A_978_357#_c_855_n 8.23715e-19 $X=7.98 $Y=1.23
+ $X2=0 $Y2=0
cc_517 N_A_200_74#_c_528_n N_A_978_357#_c_861_n 0.0168823f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_518 N_A_200_74#_c_528_n N_SET_B_M1022_g 0.00712937f $X=6.815 $Y=1.295 $X2=0
+ $Y2=0
cc_519 N_A_200_74#_c_519_n N_SET_B_c_1036_n 0.00935922f $X=6.8 $Y=2.045 $X2=0
+ $Y2=0
cc_520 N_A_200_74#_c_524_n N_SET_B_c_1036_n 0.0103776f $X=6.875 $Y=1.765 $X2=0
+ $Y2=0
cc_521 N_A_200_74#_c_525_n N_SET_B_c_1036_n 0.00541798f $X=7.775 $Y=1.395 $X2=0
+ $Y2=0
cc_522 N_A_200_74#_c_529_n N_SET_B_c_1036_n 0.0122618f $X=6.96 $Y=1.295 $X2=0
+ $Y2=0
cc_523 N_A_200_74#_c_528_n N_SET_B_c_1051_n 0.0113058f $X=6.815 $Y=1.295 $X2=0
+ $Y2=0
cc_524 N_A_200_74#_c_528_n N_SET_B_c_1037_n 0.00178987f $X=6.815 $Y=1.295 $X2=0
+ $Y2=0
cc_525 N_A_200_74#_c_521_n N_A_27_74#_M1034_g 0.00206053f $X=1.14 $Y=0.515 $X2=0
+ $Y2=0
cc_526 N_A_200_74#_c_526_n N_A_27_74#_M1034_g 0.00235546f $X=1.21 $Y=1.82 $X2=0
+ $Y2=0
cc_527 N_A_200_74#_c_536_n N_A_27_74#_c_1158_n 0.0111628f $X=1.17 $Y=2.815 $X2=0
+ $Y2=0
cc_528 N_A_200_74#_c_538_n N_A_27_74#_c_1158_n 0.00456398f $X=1.415 $Y=2.99
+ $X2=0 $Y2=0
cc_529 N_A_200_74#_c_543_n N_A_27_74#_c_1158_n 0.00608516f $X=1.17 $Y=1.985
+ $X2=0 $Y2=0
cc_530 N_A_200_74#_c_526_n N_A_27_74#_c_1158_n 0.00835618f $X=1.21 $Y=1.82 $X2=0
+ $Y2=0
cc_531 N_A_200_74#_c_527_n N_A_27_74#_c_1158_n 0.00266468f $X=1.235 $Y=1.13
+ $X2=0 $Y2=0
cc_532 N_A_200_74#_c_521_n N_A_27_74#_c_1159_n 0.00766647f $X=1.14 $Y=0.515
+ $X2=0 $Y2=0
cc_533 N_A_200_74#_c_522_n N_A_27_74#_M1001_g 0.00420477f $X=3.107 $Y=1.685
+ $X2=0 $Y2=0
cc_534 N_A_200_74#_c_530_n N_A_27_74#_M1001_g 0.0213331f $X=3.35 $Y=1.29 $X2=0
+ $Y2=0
cc_535 N_A_200_74#_c_531_n N_A_27_74#_M1001_g 0.00378881f $X=3.35 $Y=1.29 $X2=0
+ $Y2=0
cc_536 N_A_200_74#_c_532_n N_A_27_74#_M1001_g 0.0126333f $X=3.35 $Y=1.125 $X2=0
+ $Y2=0
cc_537 N_A_200_74#_c_532_n N_A_27_74#_c_1162_n 0.00882199f $X=3.35 $Y=1.125
+ $X2=0 $Y2=0
cc_538 N_A_200_74#_c_522_n N_A_27_74#_c_1175_n 0.00537991f $X=3.107 $Y=1.685
+ $X2=0 $Y2=0
cc_539 N_A_200_74#_c_545_n N_A_27_74#_c_1175_n 0.00745509f $X=3.107 $Y=1.77
+ $X2=0 $Y2=0
cc_540 N_A_200_74#_c_530_n N_A_27_74#_c_1175_n 0.0217028f $X=3.35 $Y=1.29 $X2=0
+ $Y2=0
cc_541 N_A_200_74#_c_531_n N_A_27_74#_c_1175_n 0.00215493f $X=3.35 $Y=1.29 $X2=0
+ $Y2=0
cc_542 N_A_200_74#_c_534_n N_A_27_74#_c_1176_n 0.0213211f $X=3.03 $Y=2.44 $X2=0
+ $Y2=0
cc_543 N_A_200_74#_c_540_n N_A_27_74#_c_1176_n 0.0109949f $X=2.975 $Y=1.77 $X2=0
+ $Y2=0
cc_544 N_A_200_74#_c_534_n N_A_27_74#_c_1177_n 0.0204984f $X=3.03 $Y=2.44 $X2=0
+ $Y2=0
cc_545 N_A_200_74#_c_541_n N_A_27_74#_c_1177_n 3.83539e-19 $X=3.075 $Y=2.19
+ $X2=0 $Y2=0
cc_546 N_A_200_74#_c_534_n N_A_27_74#_c_1179_n 0.0124302f $X=3.03 $Y=2.44 $X2=0
+ $Y2=0
cc_547 N_A_200_74#_c_523_n N_A_27_74#_M1024_g 0.00117954f $X=6.892 $Y=1.56 $X2=0
+ $Y2=0
cc_548 N_A_200_74#_c_520_n N_A_27_74#_c_1164_n 5.75074e-19 $X=7.98 $Y=1.23 $X2=0
+ $Y2=0
cc_549 N_A_200_74#_c_523_n N_A_27_74#_c_1164_n 0.0132432f $X=6.892 $Y=1.56 $X2=0
+ $Y2=0
cc_550 N_A_200_74#_c_525_n N_A_27_74#_c_1164_n 0.0139078f $X=7.775 $Y=1.395
+ $X2=0 $Y2=0
cc_551 N_A_200_74#_c_533_n N_A_27_74#_c_1164_n 0.0213941f $X=7.98 $Y=1.395 $X2=0
+ $Y2=0
cc_552 N_A_200_74#_c_519_n N_A_27_74#_c_1165_n 0.0167975f $X=6.8 $Y=2.045 $X2=0
+ $Y2=0
cc_553 N_A_200_74#_c_523_n N_A_27_74#_c_1165_n 0.00177344f $X=6.892 $Y=1.56
+ $X2=0 $Y2=0
cc_554 N_A_200_74#_c_528_n N_A_27_74#_c_1165_n 0.00661136f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_555 N_A_200_74#_c_525_n N_A_27_74#_c_1180_n 2.0305e-19 $X=7.775 $Y=1.395
+ $X2=0 $Y2=0
cc_556 N_A_200_74#_c_519_n N_A_27_74#_c_1181_n 0.0116454f $X=6.8 $Y=2.045 $X2=0
+ $Y2=0
cc_557 N_A_200_74#_c_519_n N_A_27_74#_c_1182_n 0.0140197f $X=6.8 $Y=2.045 $X2=0
+ $Y2=0
cc_558 N_A_200_74#_c_541_n N_A_27_74#_c_1183_n 0.00111738f $X=3.075 $Y=2.19
+ $X2=0 $Y2=0
cc_559 N_A_200_74#_c_545_n N_A_27_74#_c_1183_n 2.83685e-19 $X=3.107 $Y=1.77
+ $X2=0 $Y2=0
cc_560 N_A_200_74#_c_519_n N_A_27_74#_c_1167_n 0.0205564f $X=6.8 $Y=2.045 $X2=0
+ $Y2=0
cc_561 N_A_200_74#_c_524_n N_A_27_74#_c_1167_n 0.00514147f $X=6.875 $Y=1.765
+ $X2=0 $Y2=0
cc_562 N_A_200_74#_c_525_n N_A_27_74#_c_1167_n 0.0118811f $X=7.775 $Y=1.395
+ $X2=0 $Y2=0
cc_563 N_A_200_74#_c_536_n N_A_27_74#_c_1186_n 0.00477469f $X=1.17 $Y=2.815
+ $X2=0 $Y2=0
cc_564 N_A_200_74#_c_527_n N_A_27_74#_c_1169_n 0.0014153f $X=1.235 $Y=1.13 $X2=0
+ $Y2=0
cc_565 N_A_200_74#_c_526_n N_A_27_74#_c_1171_n 0.0048959f $X=1.21 $Y=1.82 $X2=0
+ $Y2=0
cc_566 N_A_200_74#_c_543_n N_A_27_74#_c_1172_n 0.00575748f $X=1.17 $Y=1.985
+ $X2=0 $Y2=0
cc_567 N_A_200_74#_c_526_n N_A_27_74#_c_1172_n 0.00571013f $X=1.21 $Y=1.82 $X2=0
+ $Y2=0
cc_568 N_A_200_74#_c_543_n N_A_27_74#_c_1173_n 0.00528781f $X=1.17 $Y=1.985
+ $X2=0 $Y2=0
cc_569 N_A_200_74#_c_526_n N_A_27_74#_c_1173_n 0.0251869f $X=1.21 $Y=1.82 $X2=0
+ $Y2=0
cc_570 N_A_200_74#_c_527_n N_A_27_74#_c_1173_n 0.00160233f $X=1.235 $Y=1.13
+ $X2=0 $Y2=0
cc_571 N_A_200_74#_c_520_n N_A_1534_446#_M1038_g 0.0491204f $X=7.98 $Y=1.23
+ $X2=0 $Y2=0
cc_572 N_A_200_74#_c_533_n N_A_1534_446#_c_1362_n 0.00629065f $X=7.98 $Y=1.395
+ $X2=0 $Y2=0
cc_573 N_A_200_74#_c_520_n N_A_1349_114#_c_1555_n 0.0216797f $X=7.98 $Y=1.23
+ $X2=0 $Y2=0
cc_574 N_A_200_74#_c_523_n N_A_1349_114#_c_1555_n 0.0236508f $X=6.892 $Y=1.56
+ $X2=0 $Y2=0
cc_575 N_A_200_74#_c_525_n N_A_1349_114#_c_1555_n 0.0641468f $X=7.775 $Y=1.395
+ $X2=0 $Y2=0
cc_576 N_A_200_74#_c_528_n N_A_1349_114#_c_1555_n 6.67233e-19 $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_577 N_A_200_74#_c_529_n N_A_1349_114#_c_1555_n 0.00293315f $X=6.96 $Y=1.295
+ $X2=0 $Y2=0
cc_578 N_A_200_74#_c_533_n N_A_1349_114#_c_1555_n 0.00161335f $X=7.98 $Y=1.395
+ $X2=0 $Y2=0
cc_579 N_A_200_74#_c_519_n N_A_1349_114#_c_1559_n 0.0127063f $X=6.8 $Y=2.045
+ $X2=0 $Y2=0
cc_580 N_A_200_74#_c_525_n N_A_1349_114#_c_1560_n 0.033189f $X=7.775 $Y=1.395
+ $X2=0 $Y2=0
cc_581 N_A_200_74#_c_533_n N_A_1349_114#_c_1560_n 0.0076278f $X=7.98 $Y=1.395
+ $X2=0 $Y2=0
cc_582 N_A_200_74#_c_519_n N_A_1349_114#_c_1561_n 5.92995e-19 $X=6.8 $Y=2.045
+ $X2=0 $Y2=0
cc_583 N_A_200_74#_c_524_n N_A_1349_114#_c_1561_n 0.015142f $X=6.875 $Y=1.765
+ $X2=0 $Y2=0
cc_584 N_A_200_74#_c_525_n N_A_1349_114#_c_1561_n 0.0132387f $X=7.775 $Y=1.395
+ $X2=0 $Y2=0
cc_585 N_A_200_74#_c_520_n N_A_1349_114#_c_1556_n 0.00868176f $X=7.98 $Y=1.23
+ $X2=0 $Y2=0
cc_586 N_A_200_74#_c_525_n N_A_1349_114#_c_1556_n 0.0289805f $X=7.775 $Y=1.395
+ $X2=0 $Y2=0
cc_587 N_A_200_74#_c_533_n N_A_1349_114#_c_1556_n 0.00735633f $X=7.98 $Y=1.395
+ $X2=0 $Y2=0
cc_588 N_A_200_74#_c_519_n N_A_1349_114#_c_1569_n 0.00573263f $X=6.8 $Y=2.045
+ $X2=0 $Y2=0
cc_589 N_A_200_74#_c_524_n N_A_1349_114#_c_1569_n 0.0150341f $X=6.875 $Y=1.765
+ $X2=0 $Y2=0
cc_590 N_A_200_74#_c_525_n N_A_1349_114#_c_1569_n 0.00347259f $X=7.775 $Y=1.395
+ $X2=0 $Y2=0
cc_591 N_A_200_74#_c_519_n N_A_1349_114#_c_1570_n 0.00227216f $X=6.8 $Y=2.045
+ $X2=0 $Y2=0
cc_592 N_A_200_74#_c_524_n N_A_1349_114#_c_1570_n 0.0023592f $X=6.875 $Y=1.765
+ $X2=0 $Y2=0
cc_593 N_A_200_74#_c_536_n N_VPWR_c_1793_n 0.0407093f $X=1.17 $Y=2.815 $X2=0
+ $Y2=0
cc_594 N_A_200_74#_c_538_n N_VPWR_c_1793_n 0.0119328f $X=1.415 $Y=2.99 $X2=0
+ $Y2=0
cc_595 N_A_200_74#_c_537_n N_VPWR_c_1794_n 0.0128702f $X=1.955 $Y=2.99 $X2=0
+ $Y2=0
cc_596 N_A_200_74#_c_540_n N_VPWR_c_1794_n 0.00224848f $X=2.975 $Y=1.77 $X2=0
+ $Y2=0
cc_597 N_A_200_74#_c_519_n N_VPWR_c_1796_n 0.00144618f $X=6.8 $Y=2.045 $X2=0
+ $Y2=0
cc_598 N_A_200_74#_c_537_n N_VPWR_c_1799_n 0.0469143f $X=1.955 $Y=2.99 $X2=0
+ $Y2=0
cc_599 N_A_200_74#_c_538_n N_VPWR_c_1799_n 0.0293026f $X=1.415 $Y=2.99 $X2=0
+ $Y2=0
cc_600 N_A_200_74#_c_534_n N_VPWR_c_1804_n 9.44495e-19 $X=3.03 $Y=2.44 $X2=0
+ $Y2=0
cc_601 N_A_200_74#_c_519_n N_VPWR_c_1805_n 0.00445602f $X=6.8 $Y=2.045 $X2=0
+ $Y2=0
cc_602 N_A_200_74#_c_519_n N_VPWR_c_1792_n 0.00858696f $X=6.8 $Y=2.045 $X2=0
+ $Y2=0
cc_603 N_A_200_74#_c_537_n N_VPWR_c_1792_n 0.026904f $X=1.955 $Y=2.99 $X2=0
+ $Y2=0
cc_604 N_A_200_74#_c_538_n N_VPWR_c_1792_n 0.0158659f $X=1.415 $Y=2.99 $X2=0
+ $Y2=0
cc_605 N_A_200_74#_c_537_n N_A_311_119#_M1037_s 0.00659884f $X=1.955 $Y=2.99
+ $X2=0 $Y2=0
cc_606 N_A_200_74#_c_528_n N_A_311_119#_c_1954_n 0.00551684f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_607 N_A_200_74#_c_528_n N_A_311_119#_c_1955_n 8.77327e-19 $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_608 N_A_200_74#_c_532_n N_A_311_119#_c_1955_n 0.00635523f $X=3.35 $Y=1.125
+ $X2=0 $Y2=0
cc_609 N_A_200_74#_c_532_n N_A_311_119#_c_1956_n 0.0044168f $X=3.35 $Y=1.125
+ $X2=0 $Y2=0
cc_610 N_A_200_74#_c_528_n N_A_311_119#_c_1963_n 0.00532224f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_611 N_A_200_74#_c_528_n N_A_311_119#_c_1964_n 5.75848e-19 $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_612 N_A_200_74#_c_528_n N_A_311_119#_c_1957_n 0.0131302f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_613 N_A_200_74#_c_521_n N_A_311_119#_c_1958_n 0.0570871f $X=1.14 $Y=0.515
+ $X2=0 $Y2=0
cc_614 N_A_200_74#_c_537_n N_A_311_119#_c_1966_n 0.0149535f $X=1.955 $Y=2.99
+ $X2=0 $Y2=0
cc_615 N_A_200_74#_c_539_n N_A_311_119#_c_1966_n 0.0234566f $X=2.04 $Y=2.905
+ $X2=0 $Y2=0
cc_616 N_A_200_74#_c_543_n N_A_311_119#_c_1966_n 0.0570871f $X=1.17 $Y=1.985
+ $X2=0 $Y2=0
cc_617 N_A_200_74#_c_539_n N_A_311_119#_c_1959_n 0.0347359f $X=2.04 $Y=2.905
+ $X2=0 $Y2=0
cc_618 N_A_200_74#_c_554_n N_A_311_119#_c_1959_n 0.0120098f $X=2.125 $Y=1.77
+ $X2=0 $Y2=0
cc_619 N_A_200_74#_c_527_n N_A_311_119#_c_1959_n 0.0570871f $X=1.235 $Y=1.13
+ $X2=0 $Y2=0
cc_620 N_A_200_74#_c_532_n N_A_311_119#_c_1960_n 0.00150382f $X=3.35 $Y=1.125
+ $X2=0 $Y2=0
cc_621 N_A_200_74#_c_528_n N_A_311_119#_c_1961_n 0.0150322f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_622 N_A_200_74#_c_521_n N_VGND_c_2133_n 0.0165395f $X=1.14 $Y=0.515 $X2=0
+ $Y2=0
cc_623 N_A_200_74#_c_521_n N_VGND_c_2134_n 0.00758914f $X=1.14 $Y=0.515 $X2=0
+ $Y2=0
cc_624 N_A_200_74#_c_528_n N_VGND_c_2135_n 0.00908153f $X=6.815 $Y=1.295 $X2=0
+ $Y2=0
cc_625 N_A_200_74#_c_521_n N_VGND_c_2140_n 0.0159616f $X=1.14 $Y=0.515 $X2=0
+ $Y2=0
cc_626 N_A_200_74#_c_521_n N_VGND_c_2146_n 0.0117867f $X=1.14 $Y=0.515 $X2=0
+ $Y2=0
cc_627 N_A_200_74#_c_528_n N_A_867_119#_c_2265_n 0.00677876f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_628 N_A_200_74#_c_528_n N_A_867_119#_c_2268_n 0.00908153f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_629 N_A_595_119#_c_741_n N_A_978_357#_c_848_n 0.0246055f $X=4.59 $Y=1.955
+ $X2=0 $Y2=0
cc_630 N_A_595_119#_c_749_n N_A_978_357#_c_848_n 0.0528753f $X=4.59 $Y=2.045
+ $X2=0 $Y2=0
cc_631 N_A_595_119#_M1016_g N_A_978_357#_c_848_n 0.0132724f $X=4.695 $Y=0.87
+ $X2=0 $Y2=0
cc_632 N_A_595_119#_M1016_g N_A_978_357#_M1026_g 0.0211547f $X=4.695 $Y=0.87
+ $X2=0 $Y2=0
cc_633 N_A_595_119#_M1016_g N_A_978_357#_c_861_n 2.53172e-19 $X=4.695 $Y=0.87
+ $X2=0 $Y2=0
cc_634 N_A_595_119#_c_745_n N_A_27_74#_M1001_g 0.00526053f $X=3.115 $Y=0.775
+ $X2=0 $Y2=0
cc_635 N_A_595_119#_c_746_n N_A_27_74#_M1001_g 3.07252e-19 $X=3.72 $Y=1.595
+ $X2=0 $Y2=0
cc_636 N_A_595_119#_M1016_g N_A_27_74#_c_1162_n 0.00897756f $X=4.695 $Y=0.87
+ $X2=0 $Y2=0
cc_637 N_A_595_119#_c_750_n N_A_27_74#_c_1175_n 0.00217111f $X=3.495 $Y=2.565
+ $X2=0 $Y2=0
cc_638 N_A_595_119#_c_746_n N_A_27_74#_c_1175_n 0.00872687f $X=3.72 $Y=1.595
+ $X2=0 $Y2=0
cc_639 N_A_595_119#_c_747_n N_A_27_74#_c_1175_n 0.00390887f $X=3.975 $Y=1.47
+ $X2=0 $Y2=0
cc_640 N_A_595_119#_c_750_n N_A_27_74#_c_1177_n 0.00262194f $X=3.495 $Y=2.565
+ $X2=0 $Y2=0
cc_641 N_A_595_119#_c_746_n N_A_27_74#_c_1177_n 0.00121509f $X=3.72 $Y=1.595
+ $X2=0 $Y2=0
cc_642 N_A_595_119#_c_750_n N_A_27_74#_c_1178_n 0.00614852f $X=3.495 $Y=2.565
+ $X2=0 $Y2=0
cc_643 N_A_595_119#_c_762_n N_A_27_74#_c_1179_n 0.00442313f $X=3.41 $Y=2.65
+ $X2=0 $Y2=0
cc_644 N_A_595_119#_c_750_n N_A_27_74#_c_1179_n 0.00492794f $X=3.495 $Y=2.565
+ $X2=0 $Y2=0
cc_645 N_A_595_119#_c_750_n N_A_27_74#_c_1183_n 0.0094144f $X=3.495 $Y=2.565
+ $X2=0 $Y2=0
cc_646 N_A_595_119#_c_749_n N_VPWR_c_1795_n 0.00125011f $X=4.59 $Y=2.045 $X2=0
+ $Y2=0
cc_647 N_A_595_119#_c_749_n N_VPWR_c_1804_n 0.0044313f $X=4.59 $Y=2.045 $X2=0
+ $Y2=0
cc_648 N_A_595_119#_c_749_n N_VPWR_c_1792_n 0.0045818f $X=4.59 $Y=2.045 $X2=0
+ $Y2=0
cc_649 N_A_595_119#_c_769_n N_A_311_119#_M1004_d 0.00979049f $X=3.635 $Y=0.87
+ $X2=0 $Y2=0
cc_650 N_A_595_119#_c_744_n N_A_311_119#_M1004_d 0.00185193f $X=3.72 $Y=1.395
+ $X2=0 $Y2=0
cc_651 N_A_595_119#_c_745_n N_A_311_119#_c_1968_n 0.00837589f $X=3.115 $Y=0.775
+ $X2=0 $Y2=0
cc_652 N_A_595_119#_c_745_n N_A_311_119#_c_1952_n 0.0159264f $X=3.115 $Y=0.775
+ $X2=0 $Y2=0
cc_653 N_A_595_119#_M1016_g N_A_311_119#_c_1954_n 5.72873e-19 $X=4.695 $Y=0.87
+ $X2=0 $Y2=0
cc_654 N_A_595_119#_c_769_n N_A_311_119#_c_1955_n 0.026311f $X=3.635 $Y=0.87
+ $X2=0 $Y2=0
cc_655 N_A_595_119#_c_749_n N_A_311_119#_c_1962_n 0.00186774f $X=4.59 $Y=2.045
+ $X2=0 $Y2=0
cc_656 N_A_595_119#_c_762_n N_A_311_119#_c_1962_n 0.0133863f $X=3.41 $Y=2.65
+ $X2=0 $Y2=0
cc_657 N_A_595_119#_c_750_n N_A_311_119#_c_1962_n 0.0313882f $X=3.495 $Y=2.565
+ $X2=0 $Y2=0
cc_658 N_A_595_119#_M1016_g N_A_311_119#_c_1956_n 0.00145038f $X=4.695 $Y=0.87
+ $X2=0 $Y2=0
cc_659 N_A_595_119#_c_769_n N_A_311_119#_c_1956_n 0.0135471f $X=3.635 $Y=0.87
+ $X2=0 $Y2=0
cc_660 N_A_595_119#_c_744_n N_A_311_119#_c_1956_n 0.00286902f $X=3.72 $Y=1.395
+ $X2=0 $Y2=0
cc_661 N_A_595_119#_c_740_n N_A_311_119#_c_1963_n 0.00431129f $X=4.5 $Y=1.47
+ $X2=0 $Y2=0
cc_662 N_A_595_119#_c_749_n N_A_311_119#_c_1963_n 0.00401235f $X=4.59 $Y=2.045
+ $X2=0 $Y2=0
cc_663 N_A_595_119#_c_746_n N_A_311_119#_c_1963_n 0.0106373f $X=3.72 $Y=1.595
+ $X2=0 $Y2=0
cc_664 N_A_595_119#_c_747_n N_A_311_119#_c_1963_n 9.61154e-19 $X=3.975 $Y=1.47
+ $X2=0 $Y2=0
cc_665 N_A_595_119#_c_750_n N_A_311_119#_c_1964_n 0.0136812f $X=3.495 $Y=2.565
+ $X2=0 $Y2=0
cc_666 N_A_595_119#_c_746_n N_A_311_119#_c_1964_n 0.022168f $X=3.72 $Y=1.595
+ $X2=0 $Y2=0
cc_667 N_A_595_119#_c_747_n N_A_311_119#_c_1964_n 0.00125273f $X=3.975 $Y=1.47
+ $X2=0 $Y2=0
cc_668 N_A_595_119#_c_740_n N_A_311_119#_c_1957_n 0.0134603f $X=4.5 $Y=1.47
+ $X2=0 $Y2=0
cc_669 N_A_595_119#_c_741_n N_A_311_119#_c_1957_n 0.00721254f $X=4.59 $Y=1.955
+ $X2=0 $Y2=0
cc_670 N_A_595_119#_M1016_g N_A_311_119#_c_1957_n 0.00397984f $X=4.695 $Y=0.87
+ $X2=0 $Y2=0
cc_671 N_A_595_119#_c_744_n N_A_311_119#_c_1957_n 0.00632424f $X=3.72 $Y=1.395
+ $X2=0 $Y2=0
cc_672 N_A_595_119#_c_746_n N_A_311_119#_c_1957_n 0.0312801f $X=3.72 $Y=1.595
+ $X2=0 $Y2=0
cc_673 N_A_595_119#_c_747_n N_A_311_119#_c_1957_n 0.00130314f $X=3.975 $Y=1.47
+ $X2=0 $Y2=0
cc_674 N_A_595_119#_c_769_n N_A_311_119#_c_1960_n 0.0057043f $X=3.635 $Y=0.87
+ $X2=0 $Y2=0
cc_675 N_A_595_119#_c_745_n N_A_311_119#_c_1960_n 0.0198509f $X=3.115 $Y=0.775
+ $X2=0 $Y2=0
cc_676 N_A_595_119#_c_740_n N_A_311_119#_c_1961_n 6.95961e-19 $X=4.5 $Y=1.47
+ $X2=0 $Y2=0
cc_677 N_A_595_119#_M1016_g N_A_311_119#_c_1961_n 0.00341236f $X=4.695 $Y=0.87
+ $X2=0 $Y2=0
cc_678 N_A_595_119#_c_744_n N_A_311_119#_c_1961_n 0.0137783f $X=3.72 $Y=1.395
+ $X2=0 $Y2=0
cc_679 N_A_595_119#_c_746_n N_A_311_119#_c_1961_n 0.00657374f $X=3.72 $Y=1.595
+ $X2=0 $Y2=0
cc_680 N_A_595_119#_c_747_n N_A_311_119#_c_1961_n 0.00654668f $X=3.975 $Y=1.47
+ $X2=0 $Y2=0
cc_681 N_A_595_119#_c_740_n N_A_867_119#_c_2265_n 0.00351951f $X=4.5 $Y=1.47
+ $X2=0 $Y2=0
cc_682 N_A_595_119#_M1016_g N_A_867_119#_c_2265_n 0.00948034f $X=4.695 $Y=0.87
+ $X2=0 $Y2=0
cc_683 N_A_595_119#_M1016_g N_A_867_119#_c_2266_n 0.00159671f $X=4.695 $Y=0.87
+ $X2=0 $Y2=0
cc_684 N_A_978_357#_c_848_n N_SET_B_c_1027_n 0.0451902f $X=4.98 $Y=2.045
+ $X2=-0.19 $Y2=-0.245
cc_685 N_A_978_357#_c_851_n N_SET_B_c_1027_n 0.0078907f $X=6.315 $Y=1.42
+ $X2=-0.19 $Y2=-0.245
cc_686 N_A_978_357#_c_861_n N_SET_B_c_1027_n 2.24557e-19 $X=5.125 $Y=1.42
+ $X2=-0.19 $Y2=-0.245
cc_687 N_A_978_357#_c_848_n N_SET_B_M1022_g 0.0121481f $X=4.98 $Y=2.045 $X2=0
+ $Y2=0
cc_688 N_A_978_357#_M1026_g N_SET_B_M1022_g 0.0217173f $X=5.195 $Y=0.87 $X2=0
+ $Y2=0
cc_689 N_A_978_357#_c_851_n N_SET_B_M1022_g 0.0122073f $X=6.315 $Y=1.42 $X2=0
+ $Y2=0
cc_690 N_A_978_357#_c_861_n N_SET_B_M1022_g 8.00353e-19 $X=5.125 $Y=1.42 $X2=0
+ $Y2=0
cc_691 N_A_978_357#_c_850_n N_SET_B_c_1029_n 7.28982e-19 $X=9.51 $Y=1.795 $X2=0
+ $Y2=0
cc_692 N_A_978_357#_c_912_p N_SET_B_c_1029_n 0.00528688f $X=9.3 $Y=1.02 $X2=0
+ $Y2=0
cc_693 N_A_978_357#_c_856_n N_SET_B_c_1029_n 5.89036e-19 $X=9.465 $Y=1.395 $X2=0
+ $Y2=0
cc_694 N_A_978_357#_c_857_n N_SET_B_c_1029_n 0.00828265f $X=9.465 $Y=1.395 $X2=0
+ $Y2=0
cc_695 N_A_978_357#_c_850_n N_SET_B_c_1030_n 0.00343482f $X=9.51 $Y=1.795 $X2=0
+ $Y2=0
cc_696 N_A_978_357#_c_866_n N_SET_B_c_1035_n 0.0301124f $X=9.51 $Y=1.885 $X2=0
+ $Y2=0
cc_697 N_A_978_357#_c_855_n N_SET_B_M1014_g 0.00329169f $X=8.46 $Y=0.935 $X2=0
+ $Y2=0
cc_698 N_A_978_357#_c_912_p N_SET_B_M1014_g 0.0159922f $X=9.3 $Y=1.02 $X2=0
+ $Y2=0
cc_699 N_A_978_357#_c_856_n N_SET_B_M1014_g 0.00354892f $X=9.465 $Y=1.395 $X2=0
+ $Y2=0
cc_700 N_A_978_357#_c_857_n N_SET_B_M1014_g 0.0106664f $X=9.465 $Y=1.395 $X2=0
+ $Y2=0
cc_701 N_A_978_357#_c_863_n N_SET_B_M1014_g 0.0276447f $X=9.465 $Y=1.23 $X2=0
+ $Y2=0
cc_702 N_A_978_357#_c_851_n N_SET_B_c_1036_n 0.0122852f $X=6.315 $Y=1.42 $X2=0
+ $Y2=0
cc_703 N_A_978_357#_c_848_n N_SET_B_c_1051_n 0.00120119f $X=4.98 $Y=2.045 $X2=0
+ $Y2=0
cc_704 N_A_978_357#_c_851_n N_SET_B_c_1051_n 0.00196094f $X=6.315 $Y=1.42 $X2=0
+ $Y2=0
cc_705 N_A_978_357#_c_848_n N_SET_B_c_1037_n 0.00322407f $X=4.98 $Y=2.045 $X2=0
+ $Y2=0
cc_706 N_A_978_357#_c_851_n N_SET_B_c_1037_n 0.0279177f $X=6.315 $Y=1.42 $X2=0
+ $Y2=0
cc_707 N_A_978_357#_c_850_n N_SET_B_c_1032_n 0.00625952f $X=9.51 $Y=1.795 $X2=0
+ $Y2=0
cc_708 N_A_978_357#_c_866_n N_SET_B_c_1032_n 0.00171243f $X=9.51 $Y=1.885 $X2=0
+ $Y2=0
cc_709 N_A_978_357#_c_912_p N_SET_B_c_1032_n 0.023413f $X=9.3 $Y=1.02 $X2=0
+ $Y2=0
cc_710 N_A_978_357#_c_856_n N_SET_B_c_1032_n 0.0162366f $X=9.465 $Y=1.395 $X2=0
+ $Y2=0
cc_711 N_A_978_357#_c_857_n N_SET_B_c_1032_n 0.00100533f $X=9.465 $Y=1.395 $X2=0
+ $Y2=0
cc_712 N_A_978_357#_M1026_g N_A_27_74#_c_1162_n 0.00882199f $X=5.195 $Y=0.87
+ $X2=0 $Y2=0
cc_713 N_A_978_357#_c_853_n N_A_27_74#_c_1162_n 4.42178e-19 $X=8.375 $Y=0.425
+ $X2=0 $Y2=0
cc_714 N_A_978_357#_c_854_n N_A_27_74#_c_1162_n 0.00404452f $X=6.485 $Y=0.425
+ $X2=0 $Y2=0
cc_715 N_A_978_357#_c_852_n N_A_27_74#_M1024_g 0.0114165f $X=6.4 $Y=1.335 $X2=0
+ $Y2=0
cc_716 N_A_978_357#_c_853_n N_A_27_74#_M1024_g 0.0169314f $X=8.375 $Y=0.425
+ $X2=0 $Y2=0
cc_717 N_A_978_357#_c_858_n N_A_1534_446#_M1032_d 0.00741937f $X=10.345 $Y=1.02
+ $X2=-0.19 $Y2=-0.245
cc_718 N_A_978_357#_c_938_p N_A_1534_446#_M1032_d 5.75378e-19 $X=9.465 $Y=1.02
+ $X2=-0.19 $Y2=-0.245
cc_719 N_A_978_357#_c_853_n N_A_1534_446#_M1038_g 0.00372402f $X=8.375 $Y=0.425
+ $X2=0 $Y2=0
cc_720 N_A_978_357#_c_855_n N_A_1534_446#_M1038_g 0.0105501f $X=8.46 $Y=0.935
+ $X2=0 $Y2=0
cc_721 N_A_978_357#_c_941_p N_A_1534_446#_M1038_g 0.00726228f $X=8.545 $Y=1.02
+ $X2=0 $Y2=0
cc_722 N_A_978_357#_c_866_n N_A_1534_446#_c_1363_n 0.0143867f $X=9.51 $Y=1.885
+ $X2=0 $Y2=0
cc_723 N_A_978_357#_M1008_s N_A_1534_446#_c_1351_n 0.0022485f $X=10.595 $Y=0.745
+ $X2=0 $Y2=0
cc_724 N_A_978_357#_c_857_n N_A_1534_446#_c_1351_n 3.26243e-19 $X=9.465 $Y=1.395
+ $X2=0 $Y2=0
cc_725 N_A_978_357#_c_858_n N_A_1534_446#_c_1351_n 0.0428702f $X=10.345 $Y=1.02
+ $X2=0 $Y2=0
cc_726 N_A_978_357#_c_860_n N_A_1534_446#_c_1351_n 0.0231179f $X=10.725 $Y=1.02
+ $X2=0 $Y2=0
cc_727 N_A_978_357#_c_938_p N_A_1534_446#_c_1351_n 0.00613989f $X=9.465 $Y=1.02
+ $X2=0 $Y2=0
cc_728 N_A_978_357#_c_862_n N_A_1534_446#_c_1351_n 0.0143583f $X=10.43 $Y=1.02
+ $X2=0 $Y2=0
cc_729 N_A_978_357#_c_863_n N_A_1534_446#_c_1351_n 0.00239488f $X=9.465 $Y=1.23
+ $X2=0 $Y2=0
cc_730 N_A_978_357#_c_866_n N_A_1534_446#_c_1364_n 4.98568e-19 $X=9.51 $Y=1.885
+ $X2=0 $Y2=0
cc_731 N_A_978_357#_c_866_n N_A_1534_446#_c_1365_n 8.11517e-19 $X=9.51 $Y=1.885
+ $X2=0 $Y2=0
cc_732 N_A_978_357#_M1005_s N_A_1534_446#_c_1366_n 0.0117332f $X=10.555 $Y=1.84
+ $X2=0 $Y2=0
cc_733 N_A_978_357#_c_868_n N_A_1534_446#_c_1366_n 0.014265f $X=10.515 $Y=2.035
+ $X2=0 $Y2=0
cc_734 N_A_978_357#_c_869_n N_A_1534_446#_c_1366_n 0.0201544f $X=10.685 $Y=2.035
+ $X2=0 $Y2=0
cc_735 N_A_978_357#_c_869_n N_A_1534_446#_c_1367_n 0.00713628f $X=10.685
+ $Y=2.035 $X2=0 $Y2=0
cc_736 N_A_978_357#_c_866_n N_A_1534_446#_c_1369_n 7.46086e-19 $X=9.51 $Y=1.885
+ $X2=0 $Y2=0
cc_737 N_A_978_357#_c_860_n N_A_1534_446#_c_1353_n 0.00799877f $X=10.725 $Y=1.02
+ $X2=0 $Y2=0
cc_738 N_A_978_357#_c_856_n N_A_1349_114#_M1029_g 0.00458614f $X=9.465 $Y=1.395
+ $X2=0 $Y2=0
cc_739 N_A_978_357#_c_857_n N_A_1349_114#_M1029_g 0.0207024f $X=9.465 $Y=1.395
+ $X2=0 $Y2=0
cc_740 N_A_978_357#_c_858_n N_A_1349_114#_M1029_g 0.0135044f $X=10.345 $Y=1.02
+ $X2=0 $Y2=0
cc_741 N_A_978_357#_c_859_n N_A_1349_114#_M1029_g 0.00822808f $X=10.43 $Y=1.95
+ $X2=0 $Y2=0
cc_742 N_A_978_357#_c_863_n N_A_1349_114#_M1029_g 0.0225065f $X=9.465 $Y=1.23
+ $X2=0 $Y2=0
cc_743 N_A_978_357#_c_850_n N_A_1349_114#_c_1554_n 0.0179326f $X=9.51 $Y=1.795
+ $X2=0 $Y2=0
cc_744 N_A_978_357#_c_866_n N_A_1349_114#_c_1554_n 0.0561339f $X=9.51 $Y=1.885
+ $X2=0 $Y2=0
cc_745 N_A_978_357#_c_858_n N_A_1349_114#_c_1554_n 9.39932e-19 $X=10.345 $Y=1.02
+ $X2=0 $Y2=0
cc_746 N_A_978_357#_c_859_n N_A_1349_114#_c_1554_n 0.0040159f $X=10.43 $Y=1.95
+ $X2=0 $Y2=0
cc_747 N_A_978_357#_c_868_n N_A_1349_114#_c_1554_n 8.9204e-19 $X=10.515 $Y=2.035
+ $X2=0 $Y2=0
cc_748 N_A_978_357#_c_852_n N_A_1349_114#_c_1555_n 0.02006f $X=6.4 $Y=1.335
+ $X2=0 $Y2=0
cc_749 N_A_978_357#_c_853_n N_A_1349_114#_c_1555_n 0.108619f $X=8.375 $Y=0.425
+ $X2=0 $Y2=0
cc_750 N_A_978_357#_c_855_n N_A_1349_114#_c_1555_n 0.020128f $X=8.46 $Y=0.935
+ $X2=0 $Y2=0
cc_751 N_A_978_357#_c_941_p N_A_1349_114#_c_1555_n 0.00655524f $X=8.545 $Y=1.02
+ $X2=0 $Y2=0
cc_752 N_A_978_357#_c_941_p N_A_1349_114#_c_1556_n 0.00743036f $X=8.545 $Y=1.02
+ $X2=0 $Y2=0
cc_753 N_A_978_357#_c_912_p N_A_1349_114#_c_1563_n 4.73677e-19 $X=9.3 $Y=1.02
+ $X2=0 $Y2=0
cc_754 N_A_978_357#_c_941_p N_A_1349_114#_c_1563_n 0.00452026f $X=8.545 $Y=1.02
+ $X2=0 $Y2=0
cc_755 N_A_978_357#_c_866_n N_A_1349_114#_c_1566_n 0.0143059f $X=9.51 $Y=1.885
+ $X2=0 $Y2=0
cc_756 N_A_978_357#_c_856_n N_A_1349_114#_c_1566_n 0.0091331f $X=9.465 $Y=1.395
+ $X2=0 $Y2=0
cc_757 N_A_978_357#_c_857_n N_A_1349_114#_c_1566_n 2.83373e-19 $X=9.465 $Y=1.395
+ $X2=0 $Y2=0
cc_758 N_A_978_357#_c_868_n N_A_1349_114#_c_1566_n 0.0149789f $X=10.515 $Y=2.035
+ $X2=0 $Y2=0
cc_759 N_A_978_357#_c_856_n N_A_1349_114#_c_1567_n 0.0045977f $X=9.465 $Y=1.395
+ $X2=0 $Y2=0
cc_760 N_A_978_357#_c_857_n N_A_1349_114#_c_1567_n 6.67297e-19 $X=9.465 $Y=1.395
+ $X2=0 $Y2=0
cc_761 N_A_978_357#_c_850_n N_A_1349_114#_c_1557_n 0.00213562f $X=9.51 $Y=1.795
+ $X2=0 $Y2=0
cc_762 N_A_978_357#_c_866_n N_A_1349_114#_c_1557_n 0.00135582f $X=9.51 $Y=1.885
+ $X2=0 $Y2=0
cc_763 N_A_978_357#_c_856_n N_A_1349_114#_c_1557_n 0.00887229f $X=9.465 $Y=1.395
+ $X2=0 $Y2=0
cc_764 N_A_978_357#_c_857_n N_A_1349_114#_c_1557_n 4.87607e-19 $X=9.465 $Y=1.395
+ $X2=0 $Y2=0
cc_765 N_A_978_357#_c_858_n N_A_1349_114#_c_1557_n 0.0143654f $X=10.345 $Y=1.02
+ $X2=0 $Y2=0
cc_766 N_A_978_357#_c_859_n N_A_1349_114#_c_1557_n 0.0397228f $X=10.43 $Y=1.95
+ $X2=0 $Y2=0
cc_767 N_A_978_357#_c_859_n N_RESET_B_c_1703_n 0.00678516f $X=10.43 $Y=1.95
+ $X2=-0.19 $Y2=-0.245
cc_768 N_A_978_357#_c_860_n N_RESET_B_c_1703_n 0.00101541f $X=10.725 $Y=1.02
+ $X2=-0.19 $Y2=-0.245
cc_769 N_A_978_357#_c_869_n N_RESET_B_c_1703_n 0.00340176f $X=10.685 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_770 N_A_978_357#_c_859_n N_RESET_B_M1008_g 0.00606104f $X=10.43 $Y=1.95 $X2=0
+ $Y2=0
cc_771 N_A_978_357#_c_860_n N_RESET_B_M1008_g 0.00307743f $X=10.725 $Y=1.02
+ $X2=0 $Y2=0
cc_772 N_A_978_357#_c_859_n N_RESET_B_c_1705_n 0.0327297f $X=10.43 $Y=1.95 $X2=0
+ $Y2=0
cc_773 N_A_978_357#_c_860_n N_RESET_B_c_1705_n 0.00997949f $X=10.725 $Y=1.02
+ $X2=0 $Y2=0
cc_774 N_A_978_357#_c_869_n N_RESET_B_c_1705_n 0.0109102f $X=10.685 $Y=2.035
+ $X2=0 $Y2=0
cc_775 N_A_978_357#_c_848_n N_VPWR_c_1795_n 0.00908874f $X=4.98 $Y=2.045 $X2=0
+ $Y2=0
cc_776 N_A_978_357#_c_848_n N_VPWR_c_1804_n 0.00413917f $X=4.98 $Y=2.045 $X2=0
+ $Y2=0
cc_777 N_A_978_357#_c_866_n N_VPWR_c_1807_n 0.00314375f $X=9.51 $Y=1.885 $X2=0
+ $Y2=0
cc_778 N_A_978_357#_c_848_n N_VPWR_c_1792_n 0.00414018f $X=4.98 $Y=2.045 $X2=0
+ $Y2=0
cc_779 N_A_978_357#_c_866_n N_VPWR_c_1792_n 0.00390476f $X=9.51 $Y=1.885 $X2=0
+ $Y2=0
cc_780 N_A_978_357#_c_866_n N_VPWR_c_1814_n 0.00330333f $X=9.51 $Y=1.885 $X2=0
+ $Y2=0
cc_781 N_A_978_357#_c_855_n N_VGND_M1038_d 0.00296211f $X=8.46 $Y=0.935 $X2=0
+ $Y2=0
cc_782 N_A_978_357#_c_912_p N_VGND_M1038_d 0.01748f $X=9.3 $Y=1.02 $X2=0 $Y2=0
cc_783 N_A_978_357#_c_941_p N_VGND_M1038_d 8.96084e-19 $X=8.545 $Y=1.02 $X2=0
+ $Y2=0
cc_784 N_A_978_357#_c_851_n N_VGND_c_2135_n 0.0112717f $X=6.315 $Y=1.42 $X2=0
+ $Y2=0
cc_785 N_A_978_357#_c_852_n N_VGND_c_2135_n 0.022822f $X=6.4 $Y=1.335 $X2=0
+ $Y2=0
cc_786 N_A_978_357#_c_854_n N_VGND_c_2135_n 0.014852f $X=6.485 $Y=0.425 $X2=0
+ $Y2=0
cc_787 N_A_978_357#_c_853_n N_VGND_c_2136_n 0.0141848f $X=8.375 $Y=0.425 $X2=0
+ $Y2=0
cc_788 N_A_978_357#_c_855_n N_VGND_c_2136_n 0.0187368f $X=8.46 $Y=0.935 $X2=0
+ $Y2=0
cc_789 N_A_978_357#_c_912_p N_VGND_c_2136_n 0.0135869f $X=9.3 $Y=1.02 $X2=0
+ $Y2=0
cc_790 N_A_978_357#_c_853_n N_VGND_c_2142_n 0.08689f $X=8.375 $Y=0.425 $X2=0
+ $Y2=0
cc_791 N_A_978_357#_c_854_n N_VGND_c_2142_n 0.00789578f $X=6.485 $Y=0.425 $X2=0
+ $Y2=0
cc_792 N_A_978_357#_c_863_n N_VGND_c_2143_n 0.00390708f $X=9.465 $Y=1.23 $X2=0
+ $Y2=0
cc_793 N_A_978_357#_c_853_n N_VGND_c_2146_n 0.0724187f $X=8.375 $Y=0.425 $X2=0
+ $Y2=0
cc_794 N_A_978_357#_c_854_n N_VGND_c_2146_n 0.00563471f $X=6.485 $Y=0.425 $X2=0
+ $Y2=0
cc_795 N_A_978_357#_c_863_n N_VGND_c_2146_n 0.00542671f $X=9.465 $Y=1.23 $X2=0
+ $Y2=0
cc_796 N_A_978_357#_M1026_g N_A_867_119#_c_2265_n 7.14713e-19 $X=5.195 $Y=0.87
+ $X2=0 $Y2=0
cc_797 N_A_978_357#_M1026_g N_A_867_119#_c_2266_n 0.00333342f $X=5.195 $Y=0.87
+ $X2=0 $Y2=0
cc_798 N_A_978_357#_M1026_g N_A_867_119#_c_2268_n 0.00432227f $X=5.195 $Y=0.87
+ $X2=0 $Y2=0
cc_799 N_A_978_357#_c_851_n N_A_867_119#_c_2268_n 0.0112717f $X=6.315 $Y=1.42
+ $X2=0 $Y2=0
cc_800 N_A_978_357#_c_852_n A_1254_119# 0.0103426f $X=6.4 $Y=1.335 $X2=-0.19
+ $Y2=-0.245
cc_801 N_A_978_357#_c_912_p N_A_1818_76#_M1014_d 0.00741543f $X=9.3 $Y=1.02
+ $X2=-0.19 $Y2=-0.245
cc_802 N_A_978_357#_c_858_n N_A_1818_76#_M1029_d 0.0117491f $X=10.345 $Y=1.02
+ $X2=0 $Y2=0
cc_803 N_A_978_357#_c_912_p N_A_1818_76#_c_2301_n 0.0139095f $X=9.3 $Y=1.02
+ $X2=0 $Y2=0
cc_804 N_A_978_357#_c_938_p N_A_1818_76#_c_2301_n 0.0011409f $X=9.465 $Y=1.02
+ $X2=0 $Y2=0
cc_805 N_A_978_357#_c_938_p N_A_1818_76#_c_2298_n 0.00383022f $X=9.465 $Y=1.02
+ $X2=0 $Y2=0
cc_806 N_A_978_357#_c_863_n N_A_1818_76#_c_2298_n 0.0101322f $X=9.465 $Y=1.23
+ $X2=0 $Y2=0
cc_807 N_SET_B_M1022_g N_A_27_74#_c_1162_n 0.0103062f $X=5.695 $Y=0.87 $X2=0
+ $Y2=0
cc_808 N_SET_B_c_1036_n N_A_27_74#_c_1165_n 0.00122312f $X=8.735 $Y=2.035 $X2=0
+ $Y2=0
cc_809 N_SET_B_c_1036_n N_A_27_74#_c_1181_n 0.00254121f $X=8.735 $Y=2.035 $X2=0
+ $Y2=0
cc_810 N_SET_B_c_1036_n N_A_1534_446#_M1007_s 0.00787608f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_811 SET_B N_A_1534_446#_M1007_s 8.97845e-19 $X=8.795 $Y=1.95 $X2=0 $Y2=0
cc_812 N_SET_B_c_1032_n N_A_1534_446#_M1007_s 9.5208e-19 $X=8.895 $Y=1.415 $X2=0
+ $Y2=0
cc_813 N_SET_B_c_1029_n N_A_1534_446#_M1038_g 0.0140919f $X=8.89 $Y=1.58 $X2=0
+ $Y2=0
cc_814 N_SET_B_c_1030_n N_A_1534_446#_M1038_g 0.0095843f $X=8.89 $Y=1.795 $X2=0
+ $Y2=0
cc_815 N_SET_B_c_1035_n N_A_1534_446#_M1038_g 0.0150812f $X=8.89 $Y=1.885 $X2=0
+ $Y2=0
cc_816 N_SET_B_M1014_g N_A_1534_446#_M1038_g 0.0128657f $X=9.015 $Y=0.75 $X2=0
+ $Y2=0
cc_817 N_SET_B_c_1036_n N_A_1534_446#_M1038_g 0.00213512f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_818 N_SET_B_c_1032_n N_A_1534_446#_M1038_g 0.00351656f $X=8.895 $Y=1.415
+ $X2=0 $Y2=0
cc_819 N_SET_B_c_1035_n N_A_1534_446#_c_1361_n 0.00416794f $X=8.89 $Y=1.885
+ $X2=0 $Y2=0
cc_820 N_SET_B_c_1036_n N_A_1534_446#_c_1361_n 0.0215507f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_821 N_SET_B_c_1036_n N_A_1534_446#_c_1362_n 0.00925849f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_822 N_SET_B_c_1035_n N_A_1534_446#_c_1363_n 0.00834036f $X=8.89 $Y=1.885
+ $X2=0 $Y2=0
cc_823 N_SET_B_c_1036_n N_A_1534_446#_c_1368_n 0.00557042f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_824 N_SET_B_c_1035_n N_A_1534_446#_c_1369_n 0.00451111f $X=8.89 $Y=1.885
+ $X2=0 $Y2=0
cc_825 N_SET_B_c_1036_n N_A_1534_446#_c_1369_n 3.27896e-19 $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_826 N_SET_B_c_1036_n N_A_1349_114#_c_1560_n 0.0280202f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_827 N_SET_B_c_1032_n N_A_1349_114#_c_1556_n 0.015133f $X=8.895 $Y=1.415 $X2=0
+ $Y2=0
cc_828 N_SET_B_c_1030_n N_A_1349_114#_c_1563_n 5.53942e-19 $X=8.89 $Y=1.795
+ $X2=0 $Y2=0
cc_829 N_SET_B_c_1036_n N_A_1349_114#_c_1563_n 0.00830114f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_830 N_SET_B_c_1032_n N_A_1349_114#_c_1563_n 0.0150352f $X=8.895 $Y=1.415
+ $X2=0 $Y2=0
cc_831 N_SET_B_c_1035_n N_A_1349_114#_c_1564_n 0.00216378f $X=8.89 $Y=1.885
+ $X2=0 $Y2=0
cc_832 N_SET_B_c_1036_n N_A_1349_114#_c_1564_n 0.0177878f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_833 SET_B N_A_1349_114#_c_1564_n 0.00149807f $X=8.795 $Y=1.95 $X2=0 $Y2=0
cc_834 N_SET_B_c_1032_n N_A_1349_114#_c_1564_n 0.0155323f $X=8.895 $Y=1.415
+ $X2=0 $Y2=0
cc_835 N_SET_B_c_1035_n N_A_1349_114#_c_1633_n 0.0120642f $X=8.89 $Y=1.885 $X2=0
+ $Y2=0
cc_836 N_SET_B_c_1036_n N_A_1349_114#_c_1633_n 0.00762662f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_837 SET_B N_A_1349_114#_c_1633_n 0.00758836f $X=8.795 $Y=1.95 $X2=0 $Y2=0
cc_838 N_SET_B_c_1032_n N_A_1349_114#_c_1633_n 0.0159409f $X=8.895 $Y=1.415
+ $X2=0 $Y2=0
cc_839 N_SET_B_c_1035_n N_A_1349_114#_c_1637_n 0.00172002f $X=8.89 $Y=1.885
+ $X2=0 $Y2=0
cc_840 SET_B N_A_1349_114#_c_1637_n 0.00100326f $X=8.795 $Y=1.95 $X2=0 $Y2=0
cc_841 N_SET_B_c_1035_n N_A_1349_114#_c_1567_n 6.14829e-19 $X=8.89 $Y=1.885
+ $X2=0 $Y2=0
cc_842 SET_B N_A_1349_114#_c_1567_n 0.00127852f $X=8.795 $Y=1.95 $X2=0 $Y2=0
cc_843 N_SET_B_c_1032_n N_A_1349_114#_c_1567_n 0.0131771f $X=8.895 $Y=1.415
+ $X2=0 $Y2=0
cc_844 N_SET_B_c_1036_n N_A_1349_114#_c_1569_n 0.0337565f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_845 N_SET_B_c_1036_n N_A_1349_114#_c_1570_n 0.0129511f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_846 N_SET_B_c_1036_n N_A_1349_114#_c_1571_n 0.00501285f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_847 SET_B N_VPWR_M1007_d 7.45817e-19 $X=8.795 $Y=1.95 $X2=0 $Y2=0
cc_848 N_SET_B_c_1032_n N_VPWR_M1007_d 0.00184442f $X=8.895 $Y=1.415 $X2=0 $Y2=0
cc_849 N_SET_B_c_1027_n N_VPWR_c_1795_n 0.00782017f $X=5.43 $Y=2.045 $X2=0 $Y2=0
cc_850 N_SET_B_c_1027_n N_VPWR_c_1796_n 0.00226109f $X=5.43 $Y=2.045 $X2=0 $Y2=0
cc_851 N_SET_B_c_1036_n N_VPWR_c_1796_n 0.00112478f $X=8.735 $Y=2.035 $X2=0
+ $Y2=0
cc_852 N_SET_B_c_1027_n N_VPWR_c_1801_n 0.00413917f $X=5.43 $Y=2.045 $X2=0 $Y2=0
cc_853 N_SET_B_c_1035_n N_VPWR_c_1806_n 0.00361132f $X=8.89 $Y=1.885 $X2=0 $Y2=0
cc_854 N_SET_B_c_1027_n N_VPWR_c_1792_n 0.00419307f $X=5.43 $Y=2.045 $X2=0 $Y2=0
cc_855 N_SET_B_c_1035_n N_VPWR_c_1792_n 0.00565696f $X=8.89 $Y=1.885 $X2=0 $Y2=0
cc_856 N_SET_B_c_1035_n N_VPWR_c_1813_n 0.00280081f $X=8.89 $Y=1.885 $X2=0 $Y2=0
cc_857 N_SET_B_c_1035_n N_VPWR_c_1814_n 0.00326445f $X=8.89 $Y=1.885 $X2=0 $Y2=0
cc_858 N_SET_B_M1022_g N_VGND_c_2135_n 0.00339793f $X=5.695 $Y=0.87 $X2=0 $Y2=0
cc_859 N_SET_B_M1014_g N_VGND_c_2136_n 0.00301762f $X=9.015 $Y=0.75 $X2=0 $Y2=0
cc_860 N_SET_B_M1014_g N_VGND_c_2143_n 0.00540881f $X=9.015 $Y=0.75 $X2=0 $Y2=0
cc_861 N_SET_B_M1022_g N_VGND_c_2146_n 7.85159e-19 $X=5.695 $Y=0.87 $X2=0 $Y2=0
cc_862 N_SET_B_M1014_g N_VGND_c_2146_n 0.00542671f $X=9.015 $Y=0.75 $X2=0 $Y2=0
cc_863 N_SET_B_M1022_g N_A_867_119#_c_2268_n 0.00901521f $X=5.695 $Y=0.87 $X2=0
+ $Y2=0
cc_864 N_SET_B_M1014_g N_A_1818_76#_c_2301_n 0.00407202f $X=9.015 $Y=0.75 $X2=0
+ $Y2=0
cc_865 N_SET_B_M1014_g N_A_1818_76#_c_2297_n 0.00343135f $X=9.015 $Y=0.75 $X2=0
+ $Y2=0
cc_866 N_A_27_74#_c_1182_n N_A_1534_446#_c_1354_n 0.0275254f $X=7.34 $Y=2.465
+ $X2=0 $Y2=0
cc_867 N_A_27_74#_c_1181_n N_A_1534_446#_c_1361_n 9.55001e-19 $X=7.34 $Y=2.375
+ $X2=0 $Y2=0
cc_868 N_A_27_74#_c_1181_n N_A_1534_446#_c_1362_n 0.0169874f $X=7.34 $Y=2.375
+ $X2=0 $Y2=0
cc_869 N_A_27_74#_M1024_g N_A_1349_114#_c_1555_n 0.00450135f $X=6.67 $Y=0.845
+ $X2=0 $Y2=0
cc_870 N_A_27_74#_c_1164_n N_A_1349_114#_c_1555_n 0.00454853f $X=7.25 $Y=1.27
+ $X2=0 $Y2=0
cc_871 N_A_27_74#_c_1182_n N_A_1349_114#_c_1559_n 0.0264716f $X=7.34 $Y=2.465
+ $X2=0 $Y2=0
cc_872 N_A_27_74#_c_1180_n N_A_1349_114#_c_1560_n 0.00251451f $X=7.34 $Y=1.89
+ $X2=0 $Y2=0
cc_873 N_A_27_74#_c_1181_n N_A_1349_114#_c_1560_n 3.87155e-19 $X=7.34 $Y=2.375
+ $X2=0 $Y2=0
cc_874 N_A_27_74#_c_1180_n N_A_1349_114#_c_1561_n 0.00174329f $X=7.34 $Y=1.89
+ $X2=0 $Y2=0
cc_875 N_A_27_74#_c_1167_n N_A_1349_114#_c_1561_n 0.00489714f $X=7.34 $Y=1.8
+ $X2=0 $Y2=0
cc_876 N_A_27_74#_c_1167_n N_A_1349_114#_c_1556_n 0.00358739f $X=7.34 $Y=1.8
+ $X2=0 $Y2=0
cc_877 N_A_27_74#_c_1181_n N_A_1349_114#_c_1569_n 0.0113548f $X=7.34 $Y=2.375
+ $X2=0 $Y2=0
cc_878 N_A_27_74#_c_1181_n N_A_1349_114#_c_1570_n 0.00822465f $X=7.34 $Y=2.375
+ $X2=0 $Y2=0
cc_879 N_A_27_74#_c_1200_n N_VPWR_M1030_d 0.00454793f $X=0.665 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_880 N_A_27_74#_c_1172_n N_VPWR_M1030_d 0.0015936f $X=0.75 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_881 N_A_27_74#_c_1158_n N_VPWR_c_1793_n 0.00334369f $X=0.945 $Y=1.765 $X2=0
+ $Y2=0
cc_882 N_A_27_74#_c_1186_n N_VPWR_c_1793_n 0.0449718f $X=0.27 $Y=2.815 $X2=0
+ $Y2=0
cc_883 N_A_27_74#_c_1200_n N_VPWR_c_1793_n 0.0145152f $X=0.665 $Y=2.035 $X2=0
+ $Y2=0
cc_884 N_A_27_74#_c_1158_n N_VPWR_c_1799_n 0.0044313f $X=0.945 $Y=1.765 $X2=0
+ $Y2=0
cc_885 N_A_27_74#_c_1186_n N_VPWR_c_1803_n 0.0145938f $X=0.27 $Y=2.815 $X2=0
+ $Y2=0
cc_886 N_A_27_74#_c_1179_n N_VPWR_c_1804_n 9.44495e-19 $X=3.54 $Y=2.44 $X2=0
+ $Y2=0
cc_887 N_A_27_74#_c_1182_n N_VPWR_c_1805_n 0.00292646f $X=7.34 $Y=2.465 $X2=0
+ $Y2=0
cc_888 N_A_27_74#_c_1158_n N_VPWR_c_1792_n 0.00858246f $X=0.945 $Y=1.765 $X2=0
+ $Y2=0
cc_889 N_A_27_74#_c_1182_n N_VPWR_c_1792_n 0.00396444f $X=7.34 $Y=2.465 $X2=0
+ $Y2=0
cc_890 N_A_27_74#_c_1186_n N_VPWR_c_1792_n 0.0120466f $X=0.27 $Y=2.815 $X2=0
+ $Y2=0
cc_891 N_A_27_74#_c_1159_n N_A_311_119#_c_1968_n 0.00187443f $X=2.825 $Y=0.18
+ $X2=0 $Y2=0
cc_892 N_A_27_74#_M1001_g N_A_311_119#_c_1968_n 0.0025009f $X=2.9 $Y=0.805 $X2=0
+ $Y2=0
cc_893 N_A_27_74#_M1001_g N_A_311_119#_c_1952_n 0.00592273f $X=2.9 $Y=0.805
+ $X2=0 $Y2=0
cc_894 N_A_27_74#_c_1159_n N_A_311_119#_c_1953_n 0.00466053f $X=2.825 $Y=0.18
+ $X2=0 $Y2=0
cc_895 N_A_27_74#_c_1162_n N_A_311_119#_c_1954_n 0.00420304f $X=6.595 $Y=0.18
+ $X2=0 $Y2=0
cc_896 N_A_27_74#_M1001_g N_A_311_119#_c_1955_n 0.00141636f $X=2.9 $Y=0.805
+ $X2=0 $Y2=0
cc_897 N_A_27_74#_c_1178_n N_A_311_119#_c_1962_n 0.0064597f $X=3.54 $Y=2.35
+ $X2=0 $Y2=0
cc_898 N_A_27_74#_c_1179_n N_A_311_119#_c_1962_n 0.00591631f $X=3.54 $Y=2.44
+ $X2=0 $Y2=0
cc_899 N_A_27_74#_c_1177_n N_A_311_119#_c_1964_n 0.00371933f $X=3.54 $Y=2.055
+ $X2=0 $Y2=0
cc_900 N_A_27_74#_M1034_g N_A_311_119#_c_1958_n 0.00135176f $X=0.925 $Y=0.74
+ $X2=0 $Y2=0
cc_901 N_A_27_74#_c_1159_n N_A_311_119#_c_1958_n 0.00517374f $X=2.825 $Y=0.18
+ $X2=0 $Y2=0
cc_902 N_A_27_74#_c_1158_n N_A_311_119#_c_1959_n 0.00175436f $X=0.945 $Y=1.765
+ $X2=0 $Y2=0
cc_903 N_A_27_74#_M1001_g N_A_311_119#_c_1960_n 0.0146966f $X=2.9 $Y=0.805 $X2=0
+ $Y2=0
cc_904 N_A_27_74#_c_1162_n N_A_311_119#_c_1960_n 0.0191582f $X=6.595 $Y=0.18
+ $X2=0 $Y2=0
cc_905 N_A_27_74#_c_1169_n N_VGND_M1033_d 0.00210254f $X=0.665 $Y=1.045
+ $X2=-0.19 $Y2=-0.245
cc_906 N_A_27_74#_M1034_g N_VGND_c_2133_n 0.0115341f $X=0.925 $Y=0.74 $X2=0
+ $Y2=0
cc_907 N_A_27_74#_c_1160_n N_VGND_c_2133_n 0.0075099f $X=1 $Y=0.18 $X2=0 $Y2=0
cc_908 N_A_27_74#_c_1168_n N_VGND_c_2133_n 0.0164982f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_909 N_A_27_74#_c_1169_n N_VGND_c_2133_n 0.0158226f $X=0.665 $Y=1.045 $X2=0
+ $Y2=0
cc_910 N_A_27_74#_c_1173_n N_VGND_c_2133_n 0.00102653f $X=0.96 $Y=1.465 $X2=0
+ $Y2=0
cc_911 N_A_27_74#_c_1159_n N_VGND_c_2134_n 0.0272601f $X=2.825 $Y=0.18 $X2=0
+ $Y2=0
cc_912 N_A_27_74#_M1001_g N_VGND_c_2134_n 8.03294e-19 $X=2.9 $Y=0.805 $X2=0
+ $Y2=0
cc_913 N_A_27_74#_c_1162_n N_VGND_c_2135_n 0.0256899f $X=6.595 $Y=0.18 $X2=0
+ $Y2=0
cc_914 N_A_27_74#_M1024_g N_VGND_c_2135_n 0.003017f $X=6.67 $Y=0.845 $X2=0 $Y2=0
cc_915 N_A_27_74#_c_1168_n N_VGND_c_2139_n 0.011066f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_916 N_A_27_74#_c_1160_n N_VGND_c_2140_n 0.0339223f $X=1 $Y=0.18 $X2=0 $Y2=0
cc_917 N_A_27_74#_c_1159_n N_VGND_c_2141_n 0.0774212f $X=2.825 $Y=0.18 $X2=0
+ $Y2=0
cc_918 N_A_27_74#_c_1162_n N_VGND_c_2142_n 0.016002f $X=6.595 $Y=0.18 $X2=0
+ $Y2=0
cc_919 N_A_27_74#_c_1159_n N_VGND_c_2146_n 0.0441429f $X=2.825 $Y=0.18 $X2=0
+ $Y2=0
cc_920 N_A_27_74#_c_1160_n N_VGND_c_2146_n 0.00749832f $X=1 $Y=0.18 $X2=0 $Y2=0
cc_921 N_A_27_74#_c_1162_n N_VGND_c_2146_n 0.0930344f $X=6.595 $Y=0.18 $X2=0
+ $Y2=0
cc_922 N_A_27_74#_c_1166_n N_VGND_c_2146_n 0.00370846f $X=2.9 $Y=0.18 $X2=0
+ $Y2=0
cc_923 N_A_27_74#_c_1168_n N_VGND_c_2146_n 0.00915947f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_924 N_A_27_74#_c_1162_n N_A_867_119#_c_2266_n 0.0188768f $X=6.595 $Y=0.18
+ $X2=0 $Y2=0
cc_925 N_A_27_74#_c_1162_n N_A_867_119#_c_2267_n 0.00766706f $X=6.595 $Y=0.18
+ $X2=0 $Y2=0
cc_926 N_A_1534_446#_c_1351_n N_A_1349_114#_M1029_g 0.0104522f $X=11.215 $Y=0.68
+ $X2=0 $Y2=0
cc_927 N_A_1534_446#_c_1363_n N_A_1349_114#_c_1554_n 0.0128716f $X=9.99 $Y=2.715
+ $X2=0 $Y2=0
cc_928 N_A_1534_446#_c_1364_n N_A_1349_114#_c_1554_n 0.00369207f $X=10.155
+ $Y=2.46 $X2=0 $Y2=0
cc_929 N_A_1534_446#_c_1365_n N_A_1349_114#_c_1554_n 0.00291953f $X=10.155
+ $Y=2.63 $X2=0 $Y2=0
cc_930 N_A_1534_446#_M1038_g N_A_1349_114#_c_1555_n 0.00231064f $X=8.37 $Y=0.91
+ $X2=0 $Y2=0
cc_931 N_A_1534_446#_c_1354_n N_A_1349_114#_c_1559_n 0.00234284f $X=7.76
+ $Y=2.465 $X2=0 $Y2=0
cc_932 N_A_1534_446#_c_1361_n N_A_1349_114#_c_1560_n 0.00898403f $X=8.055
+ $Y=2.215 $X2=0 $Y2=0
cc_933 N_A_1534_446#_c_1362_n N_A_1349_114#_c_1560_n 0.00578365f $X=8.055
+ $Y=2.215 $X2=0 $Y2=0
cc_934 N_A_1534_446#_M1038_g N_A_1349_114#_c_1556_n 0.0115778f $X=8.37 $Y=0.91
+ $X2=0 $Y2=0
cc_935 N_A_1534_446#_M1038_g N_A_1349_114#_c_1563_n 0.0146162f $X=8.37 $Y=0.91
+ $X2=0 $Y2=0
cc_936 N_A_1534_446#_c_1361_n N_A_1349_114#_c_1563_n 8.46766e-19 $X=8.055
+ $Y=2.215 $X2=0 $Y2=0
cc_937 N_A_1534_446#_c_1362_n N_A_1349_114#_c_1563_n 0.0027583f $X=8.055
+ $Y=2.215 $X2=0 $Y2=0
cc_938 N_A_1534_446#_M1007_s N_A_1349_114#_c_1564_n 0.00320628f $X=8.52 $Y=1.96
+ $X2=0 $Y2=0
cc_939 N_A_1534_446#_M1038_g N_A_1349_114#_c_1564_n 0.00598373f $X=8.37 $Y=0.91
+ $X2=0 $Y2=0
cc_940 N_A_1534_446#_c_1361_n N_A_1349_114#_c_1564_n 0.0153418f $X=8.055
+ $Y=2.215 $X2=0 $Y2=0
cc_941 N_A_1534_446#_c_1362_n N_A_1349_114#_c_1564_n 0.00646651f $X=8.055
+ $Y=2.215 $X2=0 $Y2=0
cc_942 N_A_1534_446#_M1007_s N_A_1349_114#_c_1633_n 0.00464867f $X=8.52 $Y=1.96
+ $X2=0 $Y2=0
cc_943 N_A_1534_446#_c_1363_n N_A_1349_114#_c_1633_n 0.0117636f $X=9.99 $Y=2.715
+ $X2=0 $Y2=0
cc_944 N_A_1534_446#_c_1369_n N_A_1349_114#_c_1633_n 0.0398435f $X=8.83 $Y=2.805
+ $X2=0 $Y2=0
cc_945 N_A_1534_446#_M1007_s N_A_1349_114#_c_1565_n 4.32645e-19 $X=8.52 $Y=1.96
+ $X2=0 $Y2=0
cc_946 N_A_1534_446#_c_1361_n N_A_1349_114#_c_1565_n 0.0142611f $X=8.055
+ $Y=2.215 $X2=0 $Y2=0
cc_947 N_A_1534_446#_c_1362_n N_A_1349_114#_c_1565_n 0.00397568f $X=8.055
+ $Y=2.215 $X2=0 $Y2=0
cc_948 N_A_1534_446#_c_1368_n N_A_1349_114#_c_1565_n 0.0139859f $X=8.5 $Y=2.805
+ $X2=0 $Y2=0
cc_949 N_A_1534_446#_M1028_d N_A_1349_114#_c_1566_n 0.00283783f $X=10.005
+ $Y=1.96 $X2=0 $Y2=0
cc_950 N_A_1534_446#_c_1363_n N_A_1349_114#_c_1566_n 0.0135034f $X=9.99 $Y=2.715
+ $X2=0 $Y2=0
cc_951 N_A_1534_446#_c_1364_n N_A_1349_114#_c_1566_n 0.0110004f $X=10.155
+ $Y=2.46 $X2=0 $Y2=0
cc_952 N_A_1534_446#_c_1362_n N_A_1349_114#_c_1569_n 0.00100073f $X=8.055
+ $Y=2.215 $X2=0 $Y2=0
cc_953 N_A_1534_446#_c_1361_n N_A_1349_114#_c_1570_n 0.0174474f $X=8.055
+ $Y=2.215 $X2=0 $Y2=0
cc_954 N_A_1534_446#_c_1362_n N_A_1349_114#_c_1570_n 8.48859e-19 $X=8.055
+ $Y=2.215 $X2=0 $Y2=0
cc_955 N_A_1534_446#_c_1361_n N_A_1349_114#_c_1571_n 0.0118206f $X=8.055
+ $Y=2.215 $X2=0 $Y2=0
cc_956 N_A_1534_446#_c_1362_n N_A_1349_114#_c_1571_n 0.00293763f $X=8.055
+ $Y=2.215 $X2=0 $Y2=0
cc_957 N_A_1534_446#_c_1356_n N_RESET_B_c_1703_n 0.0247424f $X=11.435 $Y=1.765
+ $X2=-0.19 $Y2=-0.245
cc_958 N_A_1534_446#_c_1345_n N_RESET_B_c_1703_n 0.00394665f $X=11.585 $Y=1.477
+ $X2=-0.19 $Y2=-0.245
cc_959 N_A_1534_446#_c_1365_n N_RESET_B_c_1703_n 0.00386334f $X=10.155 $Y=2.63
+ $X2=-0.19 $Y2=-0.245
cc_960 N_A_1534_446#_c_1366_n N_RESET_B_c_1703_n 0.0182209f $X=11.215 $Y=2.375
+ $X2=-0.19 $Y2=-0.245
cc_961 N_A_1534_446#_c_1367_n N_RESET_B_c_1703_n 0.00848787f $X=11.3 $Y=2.29
+ $X2=-0.19 $Y2=-0.245
cc_962 N_A_1534_446#_c_1352_n N_RESET_B_c_1703_n 0.00614026f $X=11.42 $Y=1.485
+ $X2=-0.19 $Y2=-0.245
cc_963 N_A_1534_446#_M1025_g N_RESET_B_M1008_g 0.0144563f $X=11.505 $Y=0.795
+ $X2=0 $Y2=0
cc_964 N_A_1534_446#_c_1345_n N_RESET_B_M1008_g 0.0174418f $X=11.585 $Y=1.477
+ $X2=0 $Y2=0
cc_965 N_A_1534_446#_c_1351_n N_RESET_B_M1008_g 0.013621f $X=11.215 $Y=0.68
+ $X2=0 $Y2=0
cc_966 N_A_1534_446#_c_1353_n N_RESET_B_M1008_g 0.00614026f $X=11.4 $Y=1.32
+ $X2=0 $Y2=0
cc_967 N_A_1534_446#_c_1345_n N_RESET_B_c_1705_n 6.28354e-19 $X=11.585 $Y=1.477
+ $X2=0 $Y2=0
cc_968 N_A_1534_446#_c_1351_n N_RESET_B_c_1705_n 0.00326943f $X=11.215 $Y=0.68
+ $X2=0 $Y2=0
cc_969 N_A_1534_446#_c_1366_n N_RESET_B_c_1705_n 0.00461406f $X=11.215 $Y=2.375
+ $X2=0 $Y2=0
cc_970 N_A_1534_446#_c_1352_n N_RESET_B_c_1705_n 0.0302494f $X=11.42 $Y=1.485
+ $X2=0 $Y2=0
cc_971 N_A_1534_446#_c_1359_n N_A_2412_410#_c_1741_n 0.0130881f $X=12.42
+ $Y=1.975 $X2=0 $Y2=0
cc_972 N_A_1534_446#_c_1360_n N_A_2412_410#_c_1741_n 0.00227172f $X=12.42 $Y=1.9
+ $X2=0 $Y2=0
cc_973 N_A_1534_446#_c_1346_n N_A_2412_410#_M1009_g 0.00197661f $X=12.19 $Y=1.32
+ $X2=0 $Y2=0
cc_974 N_A_1534_446#_c_1348_n N_A_2412_410#_M1009_g 0.016648f $X=12.465 $Y=0.865
+ $X2=0 $Y2=0
cc_975 N_A_1534_446#_c_1346_n N_A_2412_410#_c_1736_n 0.018228f $X=12.19 $Y=1.32
+ $X2=0 $Y2=0
cc_976 N_A_1534_446#_c_1349_n N_A_2412_410#_c_1736_n 0.00217096f $X=12.465
+ $Y=0.94 $X2=0 $Y2=0
cc_977 N_A_1534_446#_c_1350_n N_A_2412_410#_c_1736_n 0.00217986f $X=12.19
+ $Y=1.477 $X2=0 $Y2=0
cc_978 N_A_1534_446#_c_1360_n N_A_2412_410#_c_1736_n 2.79387e-19 $X=12.42 $Y=1.9
+ $X2=0 $Y2=0
cc_979 N_A_1534_446#_M1025_g N_A_2412_410#_c_1737_n 0.00269951f $X=11.505
+ $Y=0.795 $X2=0 $Y2=0
cc_980 N_A_1534_446#_c_1346_n N_A_2412_410#_c_1737_n 0.00692844f $X=12.19
+ $Y=1.32 $X2=0 $Y2=0
cc_981 N_A_1534_446#_c_1348_n N_A_2412_410#_c_1737_n 0.00313626f $X=12.465
+ $Y=0.865 $X2=0 $Y2=0
cc_982 N_A_1534_446#_c_1349_n N_A_2412_410#_c_1737_n 0.0152083f $X=12.465
+ $Y=0.94 $X2=0 $Y2=0
cc_983 N_A_1534_446#_c_1356_n N_A_2412_410#_c_1738_n 0.00151996f $X=11.435
+ $Y=1.765 $X2=0 $Y2=0
cc_984 N_A_1534_446#_c_1344_n N_A_2412_410#_c_1738_n 7.12587e-19 $X=12.115
+ $Y=1.477 $X2=0 $Y2=0
cc_985 N_A_1534_446#_c_1347_n N_A_2412_410#_c_1738_n 0.00535887f $X=12.19
+ $Y=1.825 $X2=0 $Y2=0
cc_986 N_A_1534_446#_c_1359_n N_A_2412_410#_c_1738_n 0.0144691f $X=12.42
+ $Y=1.975 $X2=0 $Y2=0
cc_987 N_A_1534_446#_c_1350_n N_A_2412_410#_c_1738_n 0.00124729f $X=12.19
+ $Y=1.477 $X2=0 $Y2=0
cc_988 N_A_1534_446#_c_1360_n N_A_2412_410#_c_1738_n 0.0141075f $X=12.42 $Y=1.9
+ $X2=0 $Y2=0
cc_989 N_A_1534_446#_c_1349_n N_A_2412_410#_c_1739_n 0.00601101f $X=12.465
+ $Y=0.94 $X2=0 $Y2=0
cc_990 N_A_1534_446#_c_1360_n N_A_2412_410#_c_1739_n 0.00591326f $X=12.42 $Y=1.9
+ $X2=0 $Y2=0
cc_991 N_A_1534_446#_c_1344_n N_A_2412_410#_c_1740_n 0.00411413f $X=12.115
+ $Y=1.477 $X2=0 $Y2=0
cc_992 N_A_1534_446#_c_1346_n N_A_2412_410#_c_1740_n 0.00204812f $X=12.19
+ $Y=1.32 $X2=0 $Y2=0
cc_993 N_A_1534_446#_c_1350_n N_A_2412_410#_c_1740_n 0.00650752f $X=12.19
+ $Y=1.477 $X2=0 $Y2=0
cc_994 N_A_1534_446#_c_1361_n N_VPWR_M1010_d 0.00285892f $X=8.055 $Y=2.215 $X2=0
+ $Y2=0
cc_995 N_A_1534_446#_c_1481_p N_VPWR_M1010_d 0.00654299f $X=8.22 $Y=2.715 $X2=0
+ $Y2=0
cc_996 N_A_1534_446#_c_1368_n N_VPWR_M1010_d 7.35761e-19 $X=8.5 $Y=2.805 $X2=0
+ $Y2=0
cc_997 N_A_1534_446#_c_1363_n N_VPWR_M1007_d 0.00840813f $X=9.99 $Y=2.715 $X2=0
+ $Y2=0
cc_998 N_A_1534_446#_c_1366_n N_VPWR_M1005_d 0.00945087f $X=11.215 $Y=2.375
+ $X2=0 $Y2=0
cc_999 N_A_1534_446#_c_1367_n N_VPWR_M1005_d 0.0053787f $X=11.3 $Y=2.29 $X2=0
+ $Y2=0
cc_1000 N_A_1534_446#_c_1356_n N_VPWR_c_1797_n 0.0114397f $X=11.435 $Y=1.765
+ $X2=0 $Y2=0
cc_1001 N_A_1534_446#_c_1366_n N_VPWR_c_1797_n 0.0227964f $X=11.215 $Y=2.375
+ $X2=0 $Y2=0
cc_1002 N_A_1534_446#_c_1359_n N_VPWR_c_1798_n 0.0102733f $X=12.42 $Y=1.975
+ $X2=0 $Y2=0
cc_1003 N_A_1534_446#_c_1360_n N_VPWR_c_1798_n 0.001526f $X=12.42 $Y=1.9 $X2=0
+ $Y2=0
cc_1004 N_A_1534_446#_c_1354_n N_VPWR_c_1805_n 0.00461464f $X=7.76 $Y=2.465
+ $X2=0 $Y2=0
cc_1005 N_A_1534_446#_c_1481_p N_VPWR_c_1805_n 3.46167e-19 $X=8.22 $Y=2.715
+ $X2=0 $Y2=0
cc_1006 N_A_1534_446#_c_1363_n N_VPWR_c_1806_n 0.00283195f $X=9.99 $Y=2.715
+ $X2=0 $Y2=0
cc_1007 N_A_1534_446#_c_1368_n N_VPWR_c_1806_n 0.00532338f $X=8.5 $Y=2.805 $X2=0
+ $Y2=0
cc_1008 N_A_1534_446#_c_1369_n N_VPWR_c_1806_n 0.013942f $X=8.83 $Y=2.805 $X2=0
+ $Y2=0
cc_1009 N_A_1534_446#_c_1363_n N_VPWR_c_1807_n 0.0256793f $X=9.99 $Y=2.715 $X2=0
+ $Y2=0
cc_1010 N_A_1534_446#_c_1356_n N_VPWR_c_1808_n 0.00413917f $X=11.435 $Y=1.765
+ $X2=0 $Y2=0
cc_1011 N_A_1534_446#_c_1359_n N_VPWR_c_1808_n 0.00513952f $X=12.42 $Y=1.975
+ $X2=0 $Y2=0
cc_1012 N_A_1534_446#_c_1354_n N_VPWR_c_1792_n 0.00913671f $X=7.76 $Y=2.465
+ $X2=0 $Y2=0
cc_1013 N_A_1534_446#_c_1356_n N_VPWR_c_1792_n 0.00822528f $X=11.435 $Y=1.765
+ $X2=0 $Y2=0
cc_1014 N_A_1534_446#_c_1359_n N_VPWR_c_1792_n 0.00523671f $X=12.42 $Y=1.975
+ $X2=0 $Y2=0
cc_1015 N_A_1534_446#_c_1362_n N_VPWR_c_1792_n 6.39414e-19 $X=8.055 $Y=2.215
+ $X2=0 $Y2=0
cc_1016 N_A_1534_446#_c_1481_p N_VPWR_c_1792_n 0.00248878f $X=8.22 $Y=2.715
+ $X2=0 $Y2=0
cc_1017 N_A_1534_446#_c_1363_n N_VPWR_c_1792_n 0.0350508f $X=9.99 $Y=2.715 $X2=0
+ $Y2=0
cc_1018 N_A_1534_446#_c_1368_n N_VPWR_c_1792_n 0.00743467f $X=8.5 $Y=2.805 $X2=0
+ $Y2=0
cc_1019 N_A_1534_446#_c_1369_n N_VPWR_c_1792_n 0.0118463f $X=8.83 $Y=2.805 $X2=0
+ $Y2=0
cc_1020 N_A_1534_446#_c_1354_n N_VPWR_c_1813_n 0.00483717f $X=7.76 $Y=2.465
+ $X2=0 $Y2=0
cc_1021 N_A_1534_446#_c_1362_n N_VPWR_c_1813_n 0.00108791f $X=8.055 $Y=2.215
+ $X2=0 $Y2=0
cc_1022 N_A_1534_446#_c_1481_p N_VPWR_c_1813_n 0.0254526f $X=8.22 $Y=2.715 $X2=0
+ $Y2=0
cc_1023 N_A_1534_446#_c_1368_n N_VPWR_c_1813_n 0.00362066f $X=8.5 $Y=2.805 $X2=0
+ $Y2=0
cc_1024 N_A_1534_446#_c_1369_n N_VPWR_c_1813_n 6.13558e-19 $X=8.83 $Y=2.805
+ $X2=0 $Y2=0
cc_1025 N_A_1534_446#_c_1363_n N_VPWR_c_1814_n 0.0244485f $X=9.99 $Y=2.715 $X2=0
+ $Y2=0
cc_1026 N_A_1534_446#_c_1369_n N_VPWR_c_1814_n 6.21521e-19 $X=8.83 $Y=2.805
+ $X2=0 $Y2=0
cc_1027 N_A_1534_446#_c_1363_n A_1917_392# 0.0052232f $X=9.99 $Y=2.715 $X2=-0.19
+ $Y2=-0.245
cc_1028 N_A_1534_446#_M1025_g N_Q_N_c_2081_n 0.0126598f $X=11.505 $Y=0.795 $X2=0
+ $Y2=0
cc_1029 N_A_1534_446#_c_1349_n N_Q_N_c_2081_n 9.53622e-19 $X=12.465 $Y=0.94
+ $X2=0 $Y2=0
cc_1030 N_A_1534_446#_M1025_g N_Q_N_c_2082_n 0.00219593f $X=11.505 $Y=0.795
+ $X2=0 $Y2=0
cc_1031 N_A_1534_446#_c_1344_n N_Q_N_c_2082_n 0.00254586f $X=12.115 $Y=1.477
+ $X2=0 $Y2=0
cc_1032 N_A_1534_446#_c_1346_n N_Q_N_c_2082_n 9.53622e-19 $X=12.19 $Y=1.32 $X2=0
+ $Y2=0
cc_1033 N_A_1534_446#_c_1352_n N_Q_N_c_2082_n 0.00203513f $X=11.42 $Y=1.485
+ $X2=0 $Y2=0
cc_1034 N_A_1534_446#_c_1356_n Q_N 0.00895694f $X=11.435 $Y=1.765 $X2=0 $Y2=0
cc_1035 N_A_1534_446#_c_1344_n Q_N 0.00531561f $X=12.115 $Y=1.477 $X2=0 $Y2=0
cc_1036 N_A_1534_446#_c_1359_n Q_N 0.00232011f $X=12.42 $Y=1.975 $X2=0 $Y2=0
cc_1037 N_A_1534_446#_c_1360_n Q_N 7.24024e-19 $X=12.42 $Y=1.9 $X2=0 $Y2=0
cc_1038 N_A_1534_446#_c_1367_n Q_N 0.0320405f $X=11.3 $Y=2.29 $X2=0 $Y2=0
cc_1039 N_A_1534_446#_c_1352_n Q_N 6.77959e-19 $X=11.42 $Y=1.485 $X2=0 $Y2=0
cc_1040 N_A_1534_446#_c_1359_n Q_N 0.00127059f $X=12.42 $Y=1.975 $X2=0 $Y2=0
cc_1041 N_A_1534_446#_c_1366_n Q_N 0.0129043f $X=11.215 $Y=2.375 $X2=0 $Y2=0
cc_1042 N_A_1534_446#_M1025_g N_Q_N_c_2083_n 0.00120695f $X=11.505 $Y=0.795
+ $X2=0 $Y2=0
cc_1043 N_A_1534_446#_c_1344_n N_Q_N_c_2083_n 0.0218962f $X=12.115 $Y=1.477
+ $X2=0 $Y2=0
cc_1044 N_A_1534_446#_c_1345_n N_Q_N_c_2083_n 0.00126172f $X=11.585 $Y=1.477
+ $X2=0 $Y2=0
cc_1045 N_A_1534_446#_c_1347_n N_Q_N_c_2083_n 7.24024e-19 $X=12.19 $Y=1.825
+ $X2=0 $Y2=0
cc_1046 N_A_1534_446#_c_1367_n N_Q_N_c_2083_n 0.00477417f $X=11.3 $Y=2.29 $X2=0
+ $Y2=0
cc_1047 N_A_1534_446#_c_1352_n N_Q_N_c_2083_n 0.023841f $X=11.42 $Y=1.485 $X2=0
+ $Y2=0
cc_1048 N_A_1534_446#_c_1353_n N_Q_N_c_2083_n 0.00523611f $X=11.4 $Y=1.32 $X2=0
+ $Y2=0
cc_1049 N_A_1534_446#_c_1348_n Q 8.51067e-19 $X=12.465 $Y=0.865 $X2=0 $Y2=0
cc_1050 N_A_1534_446#_c_1351_n N_VGND_M1008_d 0.0100046f $X=11.215 $Y=0.68 $X2=0
+ $Y2=0
cc_1051 N_A_1534_446#_c_1353_n N_VGND_M1008_d 0.00783804f $X=11.4 $Y=1.32 $X2=0
+ $Y2=0
cc_1052 N_A_1534_446#_M1038_g N_VGND_c_2136_n 5.6876e-19 $X=8.37 $Y=0.91 $X2=0
+ $Y2=0
cc_1053 N_A_1534_446#_M1025_g N_VGND_c_2137_n 0.00513051f $X=11.505 $Y=0.795
+ $X2=0 $Y2=0
cc_1054 N_A_1534_446#_c_1351_n N_VGND_c_2137_n 0.025628f $X=11.215 $Y=0.68 $X2=0
+ $Y2=0
cc_1055 N_A_1534_446#_c_1348_n N_VGND_c_2138_n 0.00549585f $X=12.465 $Y=0.865
+ $X2=0 $Y2=0
cc_1056 N_A_1534_446#_M1038_g N_VGND_c_2142_n 3.43662e-19 $X=8.37 $Y=0.91 $X2=0
+ $Y2=0
cc_1057 N_A_1534_446#_c_1351_n N_VGND_c_2143_n 0.0138172f $X=11.215 $Y=0.68
+ $X2=0 $Y2=0
cc_1058 N_A_1534_446#_M1025_g N_VGND_c_2144_n 0.00514022f $X=11.505 $Y=0.795
+ $X2=0 $Y2=0
cc_1059 N_A_1534_446#_c_1348_n N_VGND_c_2144_n 0.00461464f $X=12.465 $Y=0.865
+ $X2=0 $Y2=0
cc_1060 N_A_1534_446#_M1025_g N_VGND_c_2146_n 0.00528353f $X=11.505 $Y=0.795
+ $X2=0 $Y2=0
cc_1061 N_A_1534_446#_c_1348_n N_VGND_c_2146_n 0.00913666f $X=12.465 $Y=0.865
+ $X2=0 $Y2=0
cc_1062 N_A_1534_446#_c_1349_n N_VGND_c_2146_n 6.2279e-19 $X=12.465 $Y=0.94
+ $X2=0 $Y2=0
cc_1063 N_A_1534_446#_c_1351_n N_VGND_c_2146_n 0.0239625f $X=11.215 $Y=0.68
+ $X2=0 $Y2=0
cc_1064 N_A_1534_446#_c_1351_n N_A_1818_76#_M1029_d 0.00713159f $X=11.215
+ $Y=0.68 $X2=0 $Y2=0
cc_1065 N_A_1534_446#_M1032_d N_A_1818_76#_c_2298_n 0.00219516f $X=9.52 $Y=0.38
+ $X2=0 $Y2=0
cc_1066 N_A_1534_446#_c_1351_n N_A_1818_76#_c_2298_n 0.0466631f $X=11.215
+ $Y=0.68 $X2=0 $Y2=0
cc_1067 N_A_1349_114#_M1029_g N_RESET_B_c_1703_n 6.81196e-19 $X=9.915 $Y=0.75
+ $X2=-0.19 $Y2=-0.245
cc_1068 N_A_1349_114#_c_1554_n N_RESET_B_c_1703_n 0.00498165f $X=9.93 $Y=1.885
+ $X2=-0.19 $Y2=-0.245
cc_1069 N_A_1349_114#_c_1633_n N_VPWR_M1007_d 0.0126897f $X=9.23 $Y=2.375 $X2=0
+ $Y2=0
cc_1070 N_A_1349_114#_c_1637_n N_VPWR_M1007_d 0.00261352f $X=9.315 $Y=2.29 $X2=0
+ $Y2=0
cc_1071 N_A_1349_114#_c_1567_n N_VPWR_M1007_d 0.00154587f $X=9.4 $Y=2.035 $X2=0
+ $Y2=0
cc_1072 N_A_1349_114#_c_1559_n N_VPWR_c_1796_n 0.0101939f $X=7.025 $Y=2.815
+ $X2=0 $Y2=0
cc_1073 N_A_1349_114#_c_1559_n N_VPWR_c_1805_n 0.0241881f $X=7.025 $Y=2.815
+ $X2=0 $Y2=0
cc_1074 N_A_1349_114#_c_1554_n N_VPWR_c_1807_n 0.00361118f $X=9.93 $Y=1.885
+ $X2=0 $Y2=0
cc_1075 N_A_1349_114#_c_1554_n N_VPWR_c_1792_n 0.0056474f $X=9.93 $Y=1.885 $X2=0
+ $Y2=0
cc_1076 N_A_1349_114#_c_1559_n N_VPWR_c_1792_n 0.0196379f $X=7.025 $Y=2.815
+ $X2=0 $Y2=0
cc_1077 N_A_1349_114#_c_1559_n N_VPWR_c_1813_n 3.72769e-19 $X=7.025 $Y=2.815
+ $X2=0 $Y2=0
cc_1078 N_A_1349_114#_c_1566_n A_1917_392# 0.00284769f $X=9.84 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_1079 N_A_1349_114#_M1029_g N_VGND_c_2143_n 0.00390708f $X=9.915 $Y=0.75 $X2=0
+ $Y2=0
cc_1080 N_A_1349_114#_M1029_g N_VGND_c_2146_n 0.00542671f $X=9.915 $Y=0.75 $X2=0
+ $Y2=0
cc_1081 N_A_1349_114#_c_1555_n A_1611_140# 0.0026403f $X=8.035 $Y=0.845
+ $X2=-0.19 $Y2=-0.245
cc_1082 N_A_1349_114#_c_1556_n A_1611_140# 9.34402e-19 $X=8.12 $Y=1.73 $X2=-0.19
+ $Y2=-0.245
cc_1083 N_A_1349_114#_M1029_g N_A_1818_76#_c_2298_n 0.0108598f $X=9.915 $Y=0.75
+ $X2=0 $Y2=0
cc_1084 N_RESET_B_c_1703_n N_VPWR_c_1807_n 0.00314304f $X=10.91 $Y=1.765 $X2=0
+ $Y2=0
cc_1085 N_RESET_B_c_1703_n N_VPWR_c_1792_n 0.00411481f $X=10.91 $Y=1.765 $X2=0
+ $Y2=0
cc_1086 N_RESET_B_M1008_g N_VGND_c_2143_n 5.97925e-19 $X=10.94 $Y=0.955 $X2=0
+ $Y2=0
cc_1087 N_A_2412_410#_c_1741_n N_VPWR_c_1798_n 0.008384f $X=12.945 $Y=1.765
+ $X2=0 $Y2=0
cc_1088 N_A_2412_410#_c_1736_n N_VPWR_c_1798_n 0.00557956f $X=12.855 $Y=1.42
+ $X2=0 $Y2=0
cc_1089 N_A_2412_410#_c_1738_n N_VPWR_c_1798_n 0.0733497f $X=12.195 $Y=2.195
+ $X2=0 $Y2=0
cc_1090 N_A_2412_410#_c_1739_n N_VPWR_c_1798_n 0.016421f $X=12.67 $Y=1.42 $X2=0
+ $Y2=0
cc_1091 N_A_2412_410#_c_1738_n N_VPWR_c_1808_n 0.00858826f $X=12.195 $Y=2.195
+ $X2=0 $Y2=0
cc_1092 N_A_2412_410#_c_1741_n N_VPWR_c_1809_n 0.00445602f $X=12.945 $Y=1.765
+ $X2=0 $Y2=0
cc_1093 N_A_2412_410#_c_1741_n N_VPWR_c_1792_n 0.00865852f $X=12.945 $Y=1.765
+ $X2=0 $Y2=0
cc_1094 N_A_2412_410#_c_1738_n N_VPWR_c_1792_n 0.00874971f $X=12.195 $Y=2.195
+ $X2=0 $Y2=0
cc_1095 N_A_2412_410#_c_1737_n N_Q_N_c_2081_n 0.0657174f $X=12.25 $Y=0.58 $X2=0
+ $Y2=0
cc_1096 N_A_2412_410#_c_1738_n N_Q_N_c_2083_n 0.0999722f $X=12.195 $Y=2.195
+ $X2=0 $Y2=0
cc_1097 N_A_2412_410#_c_1740_n N_Q_N_c_2083_n 0.0240258f $X=12.235 $Y=1.42 $X2=0
+ $Y2=0
cc_1098 N_A_2412_410#_c_1741_n Q 0.0161159f $X=12.945 $Y=1.765 $X2=0 $Y2=0
cc_1099 N_A_2412_410#_M1009_g Q 0.0190895f $X=12.96 $Y=0.74 $X2=0 $Y2=0
cc_1100 N_A_2412_410#_c_1736_n Q 0.0203238f $X=12.855 $Y=1.42 $X2=0 $Y2=0
cc_1101 N_A_2412_410#_c_1737_n Q 0.0118818f $X=12.25 $Y=0.58 $X2=0 $Y2=0
cc_1102 N_A_2412_410#_c_1738_n Q 0.00657635f $X=12.195 $Y=2.195 $X2=0 $Y2=0
cc_1103 N_A_2412_410#_c_1739_n Q 0.026211f $X=12.67 $Y=1.42 $X2=0 $Y2=0
cc_1104 N_A_2412_410#_M1009_g N_VGND_c_2138_n 0.00330721f $X=12.96 $Y=0.74 $X2=0
+ $Y2=0
cc_1105 N_A_2412_410#_c_1736_n N_VGND_c_2138_n 0.0048385f $X=12.855 $Y=1.42
+ $X2=0 $Y2=0
cc_1106 N_A_2412_410#_c_1737_n N_VGND_c_2138_n 0.00252997f $X=12.25 $Y=0.58
+ $X2=0 $Y2=0
cc_1107 N_A_2412_410#_c_1739_n N_VGND_c_2138_n 0.00977708f $X=12.67 $Y=1.42
+ $X2=0 $Y2=0
cc_1108 N_A_2412_410#_c_1737_n N_VGND_c_2144_n 0.011066f $X=12.25 $Y=0.58 $X2=0
+ $Y2=0
cc_1109 N_A_2412_410#_M1009_g N_VGND_c_2145_n 0.00428607f $X=12.96 $Y=0.74 $X2=0
+ $Y2=0
cc_1110 N_A_2412_410#_M1009_g N_VGND_c_2146_n 0.00806216f $X=12.96 $Y=0.74 $X2=0
+ $Y2=0
cc_1111 N_A_2412_410#_c_1737_n N_VGND_c_2146_n 0.00915947f $X=12.25 $Y=0.58
+ $X2=0 $Y2=0
cc_1112 N_VPWR_c_1797_n Q_N 0.0241146f $X=11.21 $Y=2.805 $X2=0 $Y2=0
cc_1113 N_VPWR_c_1798_n Q_N 0.00227754f $X=12.72 $Y=1.985 $X2=0 $Y2=0
cc_1114 N_VPWR_c_1808_n Q_N 0.0155281f $X=12.555 $Y=3.33 $X2=0 $Y2=0
cc_1115 N_VPWR_c_1792_n Q_N 0.0128528f $X=13.2 $Y=3.33 $X2=0 $Y2=0
cc_1116 N_VPWR_c_1798_n Q 0.0779264f $X=12.72 $Y=1.985 $X2=0 $Y2=0
cc_1117 N_VPWR_c_1809_n Q 0.0148169f $X=13.2 $Y=3.33 $X2=0 $Y2=0
cc_1118 N_VPWR_c_1792_n Q 0.0122313f $X=13.2 $Y=3.33 $X2=0 $Y2=0
cc_1119 N_A_311_119#_c_1968_n N_VGND_M1013_d 0.00783807f $X=2.58 $Y=0.925 $X2=0
+ $Y2=0
cc_1120 N_A_311_119#_c_1968_n N_VGND_c_2134_n 0.0287269f $X=2.58 $Y=0.925 $X2=0
+ $Y2=0
cc_1121 N_A_311_119#_c_1952_n N_VGND_c_2134_n 0.0155564f $X=2.665 $Y=0.84 $X2=0
+ $Y2=0
cc_1122 N_A_311_119#_c_1953_n N_VGND_c_2134_n 0.0151473f $X=2.75 $Y=0.34 $X2=0
+ $Y2=0
cc_1123 N_A_311_119#_c_1958_n N_VGND_c_2134_n 0.00409119f $X=1.7 $Y=0.79 $X2=0
+ $Y2=0
cc_1124 N_A_311_119#_c_1958_n N_VGND_c_2140_n 0.00626553f $X=1.7 $Y=0.79 $X2=0
+ $Y2=0
cc_1125 N_A_311_119#_c_1953_n N_VGND_c_2141_n 0.0115893f $X=2.75 $Y=0.34 $X2=0
+ $Y2=0
cc_1126 N_A_311_119#_c_1954_n N_VGND_c_2141_n 0.0115893f $X=3.975 $Y=0.435 $X2=0
+ $Y2=0
cc_1127 N_A_311_119#_c_1960_n N_VGND_c_2141_n 0.0801396f $X=3.46 $Y=0.435 $X2=0
+ $Y2=0
cc_1128 N_A_311_119#_c_1968_n N_VGND_c_2146_n 0.0111714f $X=2.58 $Y=0.925 $X2=0
+ $Y2=0
cc_1129 N_A_311_119#_c_1953_n N_VGND_c_2146_n 0.00583135f $X=2.75 $Y=0.34 $X2=0
+ $Y2=0
cc_1130 N_A_311_119#_c_1954_n N_VGND_c_2146_n 0.00583135f $X=3.975 $Y=0.435
+ $X2=0 $Y2=0
cc_1131 N_A_311_119#_c_1958_n N_VGND_c_2146_n 0.00761936f $X=1.7 $Y=0.79 $X2=0
+ $Y2=0
cc_1132 N_A_311_119#_c_1960_n N_VGND_c_2146_n 0.0413441f $X=3.46 $Y=0.435 $X2=0
+ $Y2=0
cc_1133 N_A_311_119#_c_1968_n A_523_119# 0.00260391f $X=2.58 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_1134 N_A_311_119#_c_1952_n A_523_119# 0.00211902f $X=2.665 $Y=0.84 $X2=-0.19
+ $Y2=-0.245
cc_1135 N_A_311_119#_c_1961_n N_A_867_119#_M1016_s 0.00382131f $X=4.39 $Y=1.08
+ $X2=-0.19 $Y2=-0.245
cc_1136 N_A_311_119#_c_1954_n N_A_867_119#_c_2265_n 0.0167755f $X=3.975 $Y=0.435
+ $X2=0 $Y2=0
cc_1137 N_A_311_119#_c_1956_n N_A_867_119#_c_2265_n 0.0166121f $X=4.06 $Y=0.995
+ $X2=0 $Y2=0
cc_1138 N_A_311_119#_c_1961_n N_A_867_119#_c_2265_n 0.0121158f $X=4.39 $Y=1.08
+ $X2=0 $Y2=0
cc_1139 N_A_311_119#_c_1954_n N_A_867_119#_c_2267_n 0.0159286f $X=3.975 $Y=0.435
+ $X2=0 $Y2=0
cc_1140 N_Q_N_c_2081_n N_VGND_c_2137_n 0.00159581f $X=11.72 $Y=0.57 $X2=0 $Y2=0
cc_1141 N_Q_N_c_2081_n N_VGND_c_2144_n 0.0133729f $X=11.72 $Y=0.57 $X2=0 $Y2=0
cc_1142 N_Q_N_c_2081_n N_VGND_c_2146_n 0.0131093f $X=11.72 $Y=0.57 $X2=0 $Y2=0
cc_1143 Q N_VGND_c_2138_n 0.0176449f $X=13.115 $Y=0.47 $X2=0 $Y2=0
cc_1144 Q N_VGND_c_2145_n 0.0147721f $X=13.115 $Y=0.47 $X2=0 $Y2=0
cc_1145 Q N_VGND_c_2146_n 0.0121589f $X=13.115 $Y=0.47 $X2=0 $Y2=0
cc_1146 N_VGND_c_2135_n N_A_867_119#_c_2266_n 0.0150385f $X=5.98 $Y=0.87 $X2=0
+ $Y2=0
cc_1147 N_VGND_c_2141_n N_A_867_119#_c_2266_n 0.0655844f $X=5.815 $Y=0 $X2=0
+ $Y2=0
cc_1148 N_VGND_c_2146_n N_A_867_119#_c_2266_n 0.0338323f $X=13.2 $Y=0 $X2=0
+ $Y2=0
cc_1149 N_VGND_c_2141_n N_A_867_119#_c_2267_n 0.0222128f $X=5.815 $Y=0 $X2=0
+ $Y2=0
cc_1150 N_VGND_c_2146_n N_A_867_119#_c_2267_n 0.0112618f $X=13.2 $Y=0 $X2=0
+ $Y2=0
cc_1151 N_VGND_c_2135_n N_A_867_119#_c_2268_n 0.030044f $X=5.98 $Y=0.87 $X2=0
+ $Y2=0
cc_1152 N_VGND_c_2146_n N_A_1818_76#_M1029_d 0.00252807f $X=13.2 $Y=0 $X2=0
+ $Y2=0
cc_1153 N_VGND_c_2136_n N_A_1818_76#_c_2297_n 0.0113368f $X=8.8 $Y=0.56 $X2=0
+ $Y2=0
cc_1154 N_VGND_c_2143_n N_A_1818_76#_c_2297_n 0.0174569f $X=11.055 $Y=0 $X2=0
+ $Y2=0
cc_1155 N_VGND_c_2146_n N_A_1818_76#_c_2297_n 0.00963343f $X=13.2 $Y=0 $X2=0
+ $Y2=0
cc_1156 N_VGND_c_2143_n N_A_1818_76#_c_2298_n 0.0661462f $X=11.055 $Y=0 $X2=0
+ $Y2=0
cc_1157 N_VGND_c_2146_n N_A_1818_76#_c_2298_n 0.039116f $X=13.2 $Y=0 $X2=0 $Y2=0
