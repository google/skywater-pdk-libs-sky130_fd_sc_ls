* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
M1000 Y B1 a_159_74# VNB nshort w=740000u l=150000u
+  ad=2.886e+11p pd=2.26e+06u as=1.554e+11p ps=1.9e+06u
M1001 a_159_74# B2 VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=3.922e+11p ps=4.02e+06u
M1002 VPWR A1 a_71_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=4.368e+11p pd=3.02e+06u as=9.856e+11p ps=8.48e+06u
M1003 a_339_74# A1 Y VNB nshort w=740000u l=150000u
+  ad=2.886e+11p pd=2.26e+06u as=0p ps=0u
M1004 Y B2 a_71_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=0p ps=0u
M1005 a_71_368# A2 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND A2 a_339_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_71_368# B1 Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
