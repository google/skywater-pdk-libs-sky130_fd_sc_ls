* File: sky130_fd_sc_ls__buf_4.pex.spice
* Created: Fri Aug 28 13:07:13 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__BUF_4%A_86_260# 1 2 8 9 11 14 16 18 20 23 25 27 30
+ 32 34 37 39 40 47 49 50 51 52 58 61 62
c119 51 0 1.88724e-19 $X=2.285 $Y=1.045
r120 67 68 37.5985 $w=3.91e-07 $l=3.05e-07 $layer=POLY_cond $X=1.565 $Y=1.532
+ $X2=1.87 $Y2=1.532
r121 66 67 17.8747 $w=3.91e-07 $l=1.45e-07 $layer=POLY_cond $X=1.42 $Y=1.532
+ $X2=1.565 $Y2=1.532
r122 63 64 3.08184 $w=3.91e-07 $l=2.5e-08 $layer=POLY_cond $X=0.97 $Y=1.532
+ $X2=0.995 $Y2=1.532
r123 60 62 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=3.16 $Y=1.13
+ $X2=3.08 $Y2=1.045
r124 60 61 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=3.16 $Y=1.13
+ $X2=3.16 $Y2=1.95
r125 56 62 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.08 $Y=0.96
+ $X2=3.08 $Y2=1.045
r126 56 58 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=3.08 $Y=0.96
+ $X2=3.08 $Y2=0.515
r127 52 61 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.075 $Y=2.075
+ $X2=3.16 $Y2=1.95
r128 52 54 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=3.075 $Y=2.075
+ $X2=2.63 $Y2=2.075
r129 50 62 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.915 $Y=1.045
+ $X2=3.08 $Y2=1.045
r130 50 51 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=2.915 $Y=1.045
+ $X2=2.285 $Y2=1.045
r131 48 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.2 $Y=1.13
+ $X2=2.285 $Y2=1.045
r132 48 49 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.2 $Y=1.13 $X2=2.2
+ $Y2=1.3
r133 47 70 11.0946 $w=3.91e-07 $l=9e-08 $layer=POLY_cond $X=1.905 $Y=1.532
+ $X2=1.995 $Y2=1.532
r134 47 68 4.31458 $w=3.91e-07 $l=3.5e-08 $layer=POLY_cond $X=1.905 $Y=1.532
+ $X2=1.87 $Y2=1.532
r135 46 47 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.905
+ $Y=1.465 $X2=1.905 $Y2=1.465
r136 43 66 24.0384 $w=3.91e-07 $l=1.95e-07 $layer=POLY_cond $X=1.225 $Y=1.532
+ $X2=1.42 $Y2=1.532
r137 43 64 28.3529 $w=3.91e-07 $l=2.3e-07 $layer=POLY_cond $X=1.225 $Y=1.532
+ $X2=0.995 $Y2=1.532
r138 42 46 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.225 $Y=1.465
+ $X2=1.905 $Y2=1.465
r139 42 43 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.225
+ $Y=1.465 $X2=1.225 $Y2=1.465
r140 40 49 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.115 $Y=1.465
+ $X2=2.2 $Y2=1.3
r141 40 46 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=2.115 $Y=1.465
+ $X2=1.905 $Y2=1.465
r142 35 70 25.3065 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=1.995 $Y=1.3
+ $X2=1.995 $Y2=1.532
r143 35 37 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.995 $Y=1.3
+ $X2=1.995 $Y2=0.74
r144 32 68 25.3065 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=1.87 $Y=1.765
+ $X2=1.87 $Y2=1.532
r145 32 34 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.87 $Y=1.765
+ $X2=1.87 $Y2=2.4
r146 28 67 25.3065 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=1.565 $Y=1.3
+ $X2=1.565 $Y2=1.532
r147 28 30 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.565 $Y=1.3
+ $X2=1.565 $Y2=0.74
r148 25 66 25.3065 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=1.42 $Y=1.765
+ $X2=1.42 $Y2=1.532
r149 25 27 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.42 $Y=1.765
+ $X2=1.42 $Y2=2.4
r150 21 64 25.3065 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=0.995 $Y=1.3
+ $X2=0.995 $Y2=1.532
r151 21 23 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.995 $Y=1.3
+ $X2=0.995 $Y2=0.74
r152 18 63 25.3065 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=0.97 $Y=1.765
+ $X2=0.97 $Y2=1.532
r153 18 20 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.97 $Y=1.765
+ $X2=0.97 $Y2=2.4
r154 17 39 6.66866 $w=1.5e-07 $l=1.05e-07 $layer=POLY_cond $X=0.64 $Y=1.375
+ $X2=0.535 $Y2=1.375
r155 16 63 30.1682 $w=3.91e-07 $l=1.96924e-07 $layer=POLY_cond $X=0.88 $Y=1.375
+ $X2=0.97 $Y2=1.532
r156 16 17 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=0.88 $Y=1.375
+ $X2=0.64 $Y2=1.375
r157 12 39 18.8402 $w=1.65e-07 $l=8.87412e-08 $layer=POLY_cond $X=0.565 $Y=1.3
+ $X2=0.535 $Y2=1.375
r158 12 14 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.565 $Y=1.3
+ $X2=0.565 $Y2=0.74
r159 9 11 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.52 $Y=1.765
+ $X2=0.52 $Y2=2.4
r160 8 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.52 $Y=1.675 $X2=0.52
+ $Y2=1.765
r161 7 39 18.8402 $w=1.65e-07 $l=8.21584e-08 $layer=POLY_cond $X=0.52 $Y=1.45
+ $X2=0.535 $Y2=1.375
r162 7 8 87.4597 $w=1.8e-07 $l=2.25e-07 $layer=POLY_cond $X=0.52 $Y=1.45
+ $X2=0.52 $Y2=1.675
r163 2 54 600 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=2.48
+ $Y=1.84 $X2=2.63 $Y2=2.115
r164 1 58 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.94
+ $Y=0.37 $X2=3.08 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__BUF_4%A 1 3 4 6 9 11 16 17
r39 17 18 1.58553 $w=3.04e-07 $l=1e-08 $layer=POLY_cond $X=2.855 $Y=1.557
+ $X2=2.865 $Y2=1.557
r40 15 17 18.2336 $w=3.04e-07 $l=1.15e-07 $layer=POLY_cond $X=2.74 $Y=1.557
+ $X2=2.855 $Y2=1.557
r41 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.74
+ $Y=1.515 $X2=2.74 $Y2=1.515
r42 13 15 53.1151 $w=3.04e-07 $l=3.35e-07 $layer=POLY_cond $X=2.405 $Y=1.557
+ $X2=2.74 $Y2=1.557
r43 11 16 4.54912 $w=3.78e-07 $l=1.5e-07 $layer=LI1_cond $X=2.715 $Y=1.665
+ $X2=2.715 $Y2=1.515
r44 7 18 19.2802 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.865 $Y=1.35
+ $X2=2.865 $Y2=1.557
r45 7 9 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.865 $Y=1.35
+ $X2=2.865 $Y2=0.74
r46 4 17 19.2802 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.855 $Y=1.765
+ $X2=2.855 $Y2=1.557
r47 4 6 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.855 $Y=1.765
+ $X2=2.855 $Y2=2.26
r48 1 13 19.2802 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.405 $Y=1.765
+ $X2=2.405 $Y2=1.557
r49 1 3 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.405 $Y=1.765
+ $X2=2.405 $Y2=2.26
.ends

.subckt PM_SKY130_FD_SC_LS__BUF_4%VPWR 1 2 3 4 13 15 21 25 29 31 33 35 40 45 54
+ 57 61
r54 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r55 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r56 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r57 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r58 49 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r59 49 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r60 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r61 46 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.26 $Y=3.33
+ $X2=2.095 $Y2=3.33
r62 46 48 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=2.26 $Y=3.33
+ $X2=2.64 $Y2=3.33
r63 45 60 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=2.915 $Y=3.33
+ $X2=3.137 $Y2=3.33
r64 45 48 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.915 $Y=3.33
+ $X2=2.64 $Y2=3.33
r65 41 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.36 $Y=3.33
+ $X2=1.195 $Y2=3.33
r66 41 43 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.36 $Y=3.33 $X2=1.68
+ $Y2=3.33
r67 40 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.93 $Y=3.33
+ $X2=2.095 $Y2=3.33
r68 40 43 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.93 $Y=3.33
+ $X2=1.68 $Y2=3.33
r69 39 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r70 39 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r71 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r72 36 51 4.70058 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=0.46 $Y=3.33 $X2=0.23
+ $Y2=3.33
r73 36 38 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.46 $Y=3.33
+ $X2=0.72 $Y2=3.33
r74 35 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.03 $Y=3.33
+ $X2=1.195 $Y2=3.33
r75 35 38 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1.03 $Y=3.33
+ $X2=0.72 $Y2=3.33
r76 33 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r77 33 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r78 33 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r79 29 60 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=3.08 $Y=3.245
+ $X2=3.137 $Y2=3.33
r80 29 31 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=3.08 $Y=3.245
+ $X2=3.08 $Y2=2.535
r81 25 28 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=2.095 $Y=1.985
+ $X2=2.095 $Y2=2.815
r82 23 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.095 $Y=3.245
+ $X2=2.095 $Y2=3.33
r83 23 28 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.095 $Y=3.245
+ $X2=2.095 $Y2=2.815
r84 19 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.195 $Y=3.245
+ $X2=1.195 $Y2=3.33
r85 19 21 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=1.195 $Y=3.245
+ $X2=1.195 $Y2=2.225
r86 15 18 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=0.295 $Y=1.985
+ $X2=0.295 $Y2=2.815
r87 13 51 3.0656 $w=3.3e-07 $l=1.12916e-07 $layer=LI1_cond $X=0.295 $Y=3.245
+ $X2=0.23 $Y2=3.33
r88 13 18 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.295 $Y=3.245
+ $X2=0.295 $Y2=2.815
r89 4 31 600 $w=1.7e-07 $l=7.66339e-07 $layer=licon1_PDIFF $count=1 $X=2.93
+ $Y=1.84 $X2=3.08 $Y2=2.535
r90 3 28 600 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.945
+ $Y=1.84 $X2=2.095 $Y2=2.815
r91 3 25 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=1.945
+ $Y=1.84 $X2=2.095 $Y2=1.985
r92 2 21 300 $w=1.7e-07 $l=4.53845e-07 $layer=licon1_PDIFF $count=2 $X=1.045
+ $Y=1.84 $X2=1.195 $Y2=2.225
r93 1 18 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.15
+ $Y=1.84 $X2=0.295 $Y2=2.815
r94 1 15 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.15
+ $Y=1.84 $X2=0.295 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_LS__BUF_4%X 1 2 3 4 15 17 18 21 25 27 31 37 39 40
r65 40 42 11.4662 $w=2.66e-07 $l=2.5e-07 $layer=LI1_cond $X=0.775 $Y=1.295
+ $X2=0.775 $Y2=1.045
r66 35 37 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=1.78 $Y=0.96
+ $X2=1.78 $Y2=0.515
r67 31 33 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=1.645 $Y=1.985
+ $X2=1.645 $Y2=2.815
r68 29 31 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=1.645 $Y=1.97
+ $X2=1.645 $Y2=1.985
r69 28 42 3.35683 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=0.945 $Y=1.045
+ $X2=0.775 $Y2=1.045
r70 27 35 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.615 $Y=1.045
+ $X2=1.78 $Y2=0.96
r71 27 28 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.615 $Y=1.045
+ $X2=0.945 $Y2=1.045
r72 26 39 1.44715 $w=1.7e-07 $l=8.8e-08 $layer=LI1_cond $X=0.835 $Y=1.885
+ $X2=0.747 $Y2=1.885
r73 25 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.56 $Y=1.885
+ $X2=1.645 $Y2=1.97
r74 25 26 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=1.56 $Y=1.885
+ $X2=0.835 $Y2=1.885
r75 21 23 52.6026 $w=1.73e-07 $l=8.3e-07 $layer=LI1_cond $X=0.747 $Y=1.985
+ $X2=0.747 $Y2=2.815
r76 19 39 5.04255 $w=1.75e-07 $l=8.5e-08 $layer=LI1_cond $X=0.747 $Y=1.97
+ $X2=0.747 $Y2=1.885
r77 19 21 0.950649 $w=1.73e-07 $l=1.5e-08 $layer=LI1_cond $X=0.747 $Y=1.97
+ $X2=0.747 $Y2=1.985
r78 18 39 5.04255 $w=1.75e-07 $l=8.5e-08 $layer=LI1_cond $X=0.747 $Y=1.8
+ $X2=0.747 $Y2=1.885
r79 17 40 6.70265 $w=2.66e-07 $l=1.28238e-07 $layer=LI1_cond $X=0.747 $Y=1.41
+ $X2=0.775 $Y2=1.295
r80 17 18 24.7169 $w=1.73e-07 $l=3.9e-07 $layer=LI1_cond $X=0.747 $Y=1.41
+ $X2=0.747 $Y2=1.8
r81 13 42 3.63684 $w=3.3e-07 $l=8.74643e-08 $layer=LI1_cond $X=0.78 $Y=0.96
+ $X2=0.775 $Y2=1.045
r82 13 15 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=0.78 $Y=0.96
+ $X2=0.78 $Y2=0.515
r83 4 33 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.495
+ $Y=1.84 $X2=1.645 $Y2=2.815
r84 4 31 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.495
+ $Y=1.84 $X2=1.645 $Y2=1.985
r85 3 23 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.84 $X2=0.745 $Y2=2.815
r86 3 21 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.84 $X2=0.745 $Y2=1.985
r87 2 37 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.64
+ $Y=0.37 $X2=1.78 $Y2=0.515
r88 1 15 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.64
+ $Y=0.37 $X2=0.78 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__BUF_4%VGND 1 2 3 10 12 16 18 20 22 29 30 36 40
r42 41 43 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r43 40 45 9.77747 $w=6.28e-07 $l=5.15e-07 $layer=LI1_cond $X=2.43 $Y=0 $X2=2.43
+ $Y2=0.515
r44 40 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r45 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r46 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r47 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r48 30 43 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r49 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r50 27 40 8.63246 $w=1.7e-07 $l=3.15e-07 $layer=LI1_cond $X=2.745 $Y=0 $X2=2.43
+ $Y2=0
r51 27 29 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=2.745 $Y=0 $X2=3.12
+ $Y2=0
r52 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r53 26 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r54 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r55 23 33 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.222
+ $Y2=0
r56 23 25 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.72
+ $Y2=0
r57 22 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.115 $Y=0 $X2=1.28
+ $Y2=0
r58 22 25 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.115 $Y=0 $X2=0.72
+ $Y2=0
r59 20 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r60 20 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r61 19 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.445 $Y=0 $X2=1.28
+ $Y2=0
r62 18 40 8.63246 $w=1.7e-07 $l=3.15e-07 $layer=LI1_cond $X=2.115 $Y=0 $X2=2.43
+ $Y2=0
r63 18 19 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.115 $Y=0 $X2=1.445
+ $Y2=0
r64 14 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.28 $Y=0.085
+ $X2=1.28 $Y2=0
r65 14 16 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=1.28 $Y=0.085
+ $X2=1.28 $Y2=0.57
r66 10 33 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.222 $Y2=0
r67 10 12 20.7789 $w=3.28e-07 $l=5.95e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.28 $Y2=0.68
r68 3 45 182 $w=1.7e-07 $l=4.2638e-07 $layer=licon1_NDIFF $count=1 $X=2.07
+ $Y=0.37 $X2=2.43 $Y2=0.515
r69 2 16 182 $w=1.7e-07 $l=2.93428e-07 $layer=licon1_NDIFF $count=1 $X=1.07
+ $Y=0.37 $X2=1.28 $Y2=0.57
r70 1 12 182 $w=1.7e-07 $l=3.75566e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.68
.ends

