* File: sky130_fd_sc_ls__sdlclkp_2.pxi.spice
* Created: Fri Aug 28 14:06:23 2020
* 
x_PM_SKY130_FD_SC_LS__SDLCLKP_2%SCE N_SCE_c_169_n N_SCE_M1011_g N_SCE_c_174_n
+ N_SCE_M1021_g SCE N_SCE_c_171_n N_SCE_c_172_n
+ PM_SKY130_FD_SC_LS__SDLCLKP_2%SCE
x_PM_SKY130_FD_SC_LS__SDLCLKP_2%GATE N_GATE_c_201_n N_GATE_M1000_g
+ N_GATE_M1009_g GATE N_GATE_c_203_n PM_SKY130_FD_SC_LS__SDLCLKP_2%GATE
x_PM_SKY130_FD_SC_LS__SDLCLKP_2%A_318_74# N_A_318_74#_M1002_d
+ N_A_318_74#_M1003_d N_A_318_74#_c_246_n N_A_318_74#_M1017_g
+ N_A_318_74#_M1019_g N_A_318_74#_c_240_n N_A_318_74#_c_241_n
+ N_A_318_74#_c_242_n N_A_318_74#_c_243_n N_A_318_74#_c_244_n
+ N_A_318_74#_c_245_n PM_SKY130_FD_SC_LS__SDLCLKP_2%A_318_74#
x_PM_SKY130_FD_SC_LS__SDLCLKP_2%A_288_48# N_A_288_48#_M1023_s
+ N_A_288_48#_M1013_s N_A_288_48#_c_323_n N_A_288_48#_M1002_g
+ N_A_288_48#_c_324_n N_A_288_48#_c_325_n N_A_288_48#_c_326_n
+ N_A_288_48#_c_343_n N_A_288_48#_c_344_n N_A_288_48#_c_345_n
+ N_A_288_48#_M1003_g N_A_288_48#_c_347_n N_A_288_48#_c_348_n
+ N_A_288_48#_c_327_n N_A_288_48#_c_328_n N_A_288_48#_c_329_n
+ N_A_288_48#_M1022_g N_A_288_48#_c_349_n N_A_288_48#_c_350_n
+ N_A_288_48#_c_351_n N_A_288_48#_M1004_g N_A_288_48#_c_330_n
+ N_A_288_48#_c_331_n N_A_288_48#_c_332_n N_A_288_48#_c_333_n
+ N_A_288_48#_c_334_n N_A_288_48#_c_335_n N_A_288_48#_c_393_p
+ N_A_288_48#_c_336_n N_A_288_48#_c_337_n N_A_288_48#_c_338_n
+ N_A_288_48#_c_339_n N_A_288_48#_c_340_n N_A_288_48#_c_352_n
+ N_A_288_48#_c_341_n PM_SKY130_FD_SC_LS__SDLCLKP_2%A_288_48#
x_PM_SKY130_FD_SC_LS__SDLCLKP_2%A_706_317# N_A_706_317#_M1001_d
+ N_A_706_317#_M1008_d N_A_706_317#_M1020_g N_A_706_317#_c_502_n
+ N_A_706_317#_c_503_n N_A_706_317#_M1012_g N_A_706_317#_M1007_g
+ N_A_706_317#_c_493_n N_A_706_317#_M1010_g N_A_706_317#_c_505_n
+ N_A_706_317#_c_506_n N_A_706_317#_c_507_n N_A_706_317#_c_494_n
+ N_A_706_317#_c_495_n N_A_706_317#_c_509_n N_A_706_317#_c_496_n
+ N_A_706_317#_c_497_n N_A_706_317#_c_498_n N_A_706_317#_c_499_n
+ N_A_706_317#_c_512_n N_A_706_317#_c_513_n N_A_706_317#_c_500_n
+ N_A_706_317#_c_501_n PM_SKY130_FD_SC_LS__SDLCLKP_2%A_706_317#
x_PM_SKY130_FD_SC_LS__SDLCLKP_2%A_580_74# N_A_580_74#_M1022_d
+ N_A_580_74#_M1017_d N_A_580_74#_c_626_n N_A_580_74#_M1008_g
+ N_A_580_74#_c_627_n N_A_580_74#_M1001_g N_A_580_74#_c_636_n
+ N_A_580_74#_c_628_n N_A_580_74#_c_629_n N_A_580_74#_c_633_n
+ N_A_580_74#_c_630_n N_A_580_74#_c_648_n N_A_580_74#_c_631_n
+ PM_SKY130_FD_SC_LS__SDLCLKP_2%A_580_74#
x_PM_SKY130_FD_SC_LS__SDLCLKP_2%CLK N_CLK_c_715_n N_CLK_M1013_g N_CLK_c_710_n
+ N_CLK_M1023_g N_CLK_c_711_n N_CLK_c_712_n N_CLK_c_718_n N_CLK_M1018_g
+ N_CLK_c_713_n N_CLK_M1015_g CLK PM_SKY130_FD_SC_LS__SDLCLKP_2%CLK
x_PM_SKY130_FD_SC_LS__SDLCLKP_2%A_1195_374# N_A_1195_374#_M1007_d
+ N_A_1195_374#_M1018_d N_A_1195_374#_c_775_n N_A_1195_374#_M1006_g
+ N_A_1195_374#_M1005_g N_A_1195_374#_c_776_n N_A_1195_374#_M1014_g
+ N_A_1195_374#_M1016_g N_A_1195_374#_c_777_n N_A_1195_374#_c_768_n
+ N_A_1195_374#_c_778_n N_A_1195_374#_c_779_n N_A_1195_374#_c_769_n
+ N_A_1195_374#_c_770_n N_A_1195_374#_c_771_n N_A_1195_374#_c_772_n
+ N_A_1195_374#_c_773_n N_A_1195_374#_c_774_n
+ PM_SKY130_FD_SC_LS__SDLCLKP_2%A_1195_374#
x_PM_SKY130_FD_SC_LS__SDLCLKP_2%VPWR N_VPWR_M1021_s N_VPWR_M1003_s
+ N_VPWR_M1012_d N_VPWR_M1013_d N_VPWR_M1010_d N_VPWR_M1014_s N_VPWR_c_854_n
+ N_VPWR_c_855_n N_VPWR_c_856_n N_VPWR_c_857_n N_VPWR_c_858_n N_VPWR_c_859_n
+ N_VPWR_c_860_n N_VPWR_c_861_n N_VPWR_c_862_n N_VPWR_c_863_n VPWR
+ N_VPWR_c_864_n N_VPWR_c_865_n N_VPWR_c_866_n N_VPWR_c_867_n N_VPWR_c_868_n
+ N_VPWR_c_869_n N_VPWR_c_870_n N_VPWR_c_853_n
+ PM_SKY130_FD_SC_LS__SDLCLKP_2%VPWR
x_PM_SKY130_FD_SC_LS__SDLCLKP_2%A_114_112# N_A_114_112#_M1011_d
+ N_A_114_112#_M1022_s N_A_114_112#_M1000_d N_A_114_112#_M1017_s
+ N_A_114_112#_c_948_n N_A_114_112#_c_963_n N_A_114_112#_c_949_n
+ N_A_114_112#_c_950_n N_A_114_112#_c_951_n N_A_114_112#_c_954_n
+ N_A_114_112#_c_952_n N_A_114_112#_c_956_n N_A_114_112#_c_957_n
+ N_A_114_112#_c_958_n N_A_114_112#_c_959_n N_A_114_112#_c_953_n
+ PM_SKY130_FD_SC_LS__SDLCLKP_2%A_114_112#
x_PM_SKY130_FD_SC_LS__SDLCLKP_2%GCLK N_GCLK_M1005_d N_GCLK_M1006_d
+ N_GCLK_c_1047_n N_GCLK_c_1048_n GCLK GCLK GCLK GCLK N_GCLK_c_1049_n
+ PM_SKY130_FD_SC_LS__SDLCLKP_2%GCLK
x_PM_SKY130_FD_SC_LS__SDLCLKP_2%VGND N_VGND_M1011_s N_VGND_M1009_d
+ N_VGND_M1020_d N_VGND_M1023_d N_VGND_M1005_s N_VGND_M1016_s N_VGND_c_1084_n
+ N_VGND_c_1085_n N_VGND_c_1086_n N_VGND_c_1087_n N_VGND_c_1088_n
+ N_VGND_c_1089_n N_VGND_c_1090_n N_VGND_c_1091_n N_VGND_c_1092_n
+ N_VGND_c_1093_n N_VGND_c_1094_n VGND N_VGND_c_1095_n N_VGND_c_1096_n
+ N_VGND_c_1097_n N_VGND_c_1098_n N_VGND_c_1099_n N_VGND_c_1100_n
+ PM_SKY130_FD_SC_LS__SDLCLKP_2%VGND
cc_1 VNB N_SCE_c_169_n 0.0160819f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1.778
cc_2 VNB N_SCE_M1011_g 0.0259574f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.835
cc_3 VNB N_SCE_c_171_n 0.0228767f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.455
cc_4 VNB N_SCE_c_172_n 0.0150846f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.455
cc_5 VNB N_GATE_c_201_n 0.00752214f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1.472
cc_6 VNB N_GATE_M1009_g 0.0410235f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_GATE_c_203_n 0.0039698f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1.455
cc_8 VNB N_A_318_74#_M1019_g 0.0290535f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1.455
cc_9 VNB N_A_318_74#_c_240_n 0.00409123f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1.29
cc_10 VNB N_A_318_74#_c_241_n 0.00340601f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.625
cc_11 VNB N_A_318_74#_c_242_n 0.00392562f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_318_74#_c_243_n 0.00407793f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_318_74#_c_244_n 0.0039819f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_318_74#_c_245_n 0.060829f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_288_48#_c_323_n 0.0222943f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.045
cc_16 VNB N_A_288_48#_c_324_n 0.0196979f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_17 VNB N_A_288_48#_c_325_n 0.00949141f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_288_48#_c_326_n 0.0229124f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.455
cc_19 VNB N_A_288_48#_c_327_n 0.0286287f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_288_48#_c_328_n 0.0570075f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_288_48#_c_329_n 0.018287f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_288_48#_c_330_n 0.0017689f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_288_48#_c_331_n 0.00620923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_288_48#_c_332_n 0.0054008f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_288_48#_c_333_n 4.56848e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_288_48#_c_334_n 0.0083234f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_288_48#_c_335_n 0.00200416f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_288_48#_c_336_n 0.0157841f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_288_48#_c_337_n 0.00232637f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_288_48#_c_338_n 0.00425067f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_288_48#_c_339_n 0.0103992f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_288_48#_c_340_n 0.001685f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_288_48#_c_341_n 0.00972167f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_706_317#_M1020_g 0.0516566f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.54
cc_35 VNB N_A_706_317#_M1007_g 0.0244504f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_706_317#_c_493_n 0.0418962f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_706_317#_c_494_n 0.00340445f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_706_317#_c_495_n 0.00882689f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_706_317#_c_496_n 3.62031e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_706_317#_c_497_n 6.10912e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_706_317#_c_498_n 0.0137603f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_706_317#_c_499_n 0.00147549f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_706_317#_c_500_n 0.00121771f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_706_317#_c_501_n 0.00835532f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_580_74#_c_626_n 0.029437f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.045
cc_46 VNB N_A_580_74#_c_627_n 0.019747f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_47 VNB N_A_580_74#_c_628_n 0.00278951f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_580_74#_c_629_n 0.018075f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_580_74#_c_630_n 0.0022609f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_580_74#_c_631_n 0.00177044f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_CLK_c_710_n 0.0198677f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.835
cc_52 VNB N_CLK_c_711_n 0.0548824f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.045
cc_53 VNB N_CLK_c_712_n 0.00279639f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.54
cc_54 VNB N_CLK_c_713_n 0.0169383f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1.455
cc_55 VNB CLK 0.00687956f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1.29
cc_56 VNB N_A_1195_374#_M1005_g 0.0224327f $X=-0.19 $Y=-0.245 $X2=0.402
+ $Y2=1.455
cc_57 VNB N_A_1195_374#_M1016_g 0.0266863f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.625
cc_58 VNB N_A_1195_374#_c_768_n 0.00882336f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_1195_374#_c_769_n 0.012386f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_1195_374#_c_770_n 0.0024413f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_1195_374#_c_771_n 5.02584e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_1195_374#_c_772_n 0.00651904f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_1195_374#_c_773_n 0.00347217f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_1195_374#_c_774_n 0.0808246f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VPWR_c_853_n 0.342803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_114_112#_c_948_n 0.011371f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.455
cc_67 VNB N_A_114_112#_c_949_n 0.00956352f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_114_112#_c_950_n 0.00325069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_114_112#_c_951_n 0.0148174f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.625
cc_70 VNB N_A_114_112#_c_952_n 0.00557558f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_114_112#_c_953_n 0.00641776f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_GCLK_c_1047_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.54
cc_73 VNB N_GCLK_c_1048_n 0.00448002f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.455
cc_74 VNB N_GCLK_c_1049_n 0.0030223f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1084_n 0.010678f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.625
cc_76 VNB N_VGND_c_1085_n 0.0503665f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1086_n 0.00858671f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1087_n 0.006053f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1088_n 0.0133405f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1089_n 0.010359f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1090_n 0.050871f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1091_n 0.0621246f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1092_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1093_n 0.0364191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1094_n 0.00615884f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1095_n 0.0191861f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1096_n 0.0291972f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1097_n 0.0193312f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1098_n 0.017485f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1099_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_VGND_c_1100_n 0.469354f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VPB N_SCE_c_169_n 0.0381764f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=1.778
cc_93 VPB N_SCE_c_174_n 0.0189667f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.045
cc_94 VPB N_SCE_c_172_n 0.0123922f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.455
cc_95 VPB N_GATE_c_201_n 0.0518772f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=1.472
cc_96 VPB N_GATE_c_203_n 0.00506155f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=1.455
cc_97 VPB N_A_318_74#_c_246_n 0.0182613f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.045
cc_98 VPB N_A_318_74#_c_241_n 0.00494693f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.625
cc_99 VPB N_A_318_74#_c_243_n 0.00747384f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 VPB N_A_318_74#_c_244_n 0.00290184f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB N_A_318_74#_c_245_n 0.026766f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_102 VPB N_A_288_48#_c_326_n 9.91146e-19 $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.455
cc_103 VPB N_A_288_48#_c_343_n 0.00878351f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.455
cc_104 VPB N_A_288_48#_c_344_n 0.0202251f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=1.29
cc_105 VPB N_A_288_48#_c_345_n 0.00748337f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.625
cc_106 VPB N_A_288_48#_M1003_g 0.0102221f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.625
cc_107 VPB N_A_288_48#_c_347_n 0.111588f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_A_288_48#_c_348_n 0.0139988f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_109 VPB N_A_288_48#_c_349_n 0.00720327f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_110 VPB N_A_288_48#_c_350_n 0.0214052f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_A_288_48#_c_351_n 0.0191972f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_A_288_48#_c_352_n 0.00725076f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_A_288_48#_c_341_n 0.00292333f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_A_706_317#_c_502_n 0.0117206f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=1.455
cc_115 VPB N_A_706_317#_c_503_n 0.0232286f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.455
cc_116 VPB N_A_706_317#_c_493_n 0.0264042f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_A_706_317#_c_505_n 0.00527081f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_A_706_317#_c_506_n 0.00413045f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_A_706_317#_c_507_n 0.0176004f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_A_706_317#_c_495_n 0.00383352f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_A_706_317#_c_509_n 0.0134329f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_A_706_317#_c_496_n 0.0022385f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_A_706_317#_c_499_n 0.00876761f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_A_706_317#_c_512_n 0.00602039f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_A_706_317#_c_513_n 5.34456e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 VPB N_A_706_317#_c_501_n 0.0340855f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_127 VPB N_A_580_74#_c_626_n 0.0342743f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.045
cc_128 VPB N_A_580_74#_c_633_n 0.00122423f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_129 VPB N_A_580_74#_c_630_n 0.00732221f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_A_580_74#_c_631_n 0.00137316f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_CLK_c_715_n 0.0180833f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=1.472
cc_132 VPB N_CLK_c_711_n 0.00730728f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.045
cc_133 VPB N_CLK_c_712_n 0.00549609f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.54
cc_134 VPB N_CLK_c_718_n 0.0237763f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.54
cc_135 VPB N_A_1195_374#_c_775_n 0.0165013f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.045
cc_136 VPB N_A_1195_374#_c_776_n 0.0174144f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.455
cc_137 VPB N_A_1195_374#_c_777_n 0.00338422f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_A_1195_374#_c_778_n 0.00387888f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_A_1195_374#_c_779_n 0.00275202f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_140 VPB N_A_1195_374#_c_771_n 0.00236962f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_141 VPB N_A_1195_374#_c_774_n 0.0170011f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_142 VPB N_VPWR_c_854_n 0.0116916f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.625
cc_143 VPB N_VPWR_c_855_n 0.0427764f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_144 VPB N_VPWR_c_856_n 0.0163243f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_145 VPB N_VPWR_c_857_n 0.0173524f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_146 VPB N_VPWR_c_858_n 0.0250916f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_147 VPB N_VPWR_c_859_n 0.0130642f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_148 VPB N_VPWR_c_860_n 0.0124065f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_149 VPB N_VPWR_c_861_n 0.064296f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_150 VPB N_VPWR_c_862_n 0.0254743f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_151 VPB N_VPWR_c_863_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_152 VPB N_VPWR_c_864_n 0.0306291f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_153 VPB N_VPWR_c_865_n 0.0663018f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_154 VPB N_VPWR_c_866_n 0.0376907f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_155 VPB N_VPWR_c_867_n 0.0194542f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_156 VPB N_VPWR_c_868_n 0.00626979f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_157 VPB N_VPWR_c_869_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_158 VPB N_VPWR_c_870_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_159 VPB N_VPWR_c_853_n 0.135857f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_160 VPB N_A_114_112#_c_954_n 0.0105766f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_161 VPB N_A_114_112#_c_952_n 0.00853783f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_162 VPB N_A_114_112#_c_956_n 0.0132669f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_163 VPB N_A_114_112#_c_957_n 0.00689851f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_164 VPB N_A_114_112#_c_958_n 0.00890932f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_165 VPB N_A_114_112#_c_959_n 8.47548e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_166 VPB GCLK 0.00194876f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.455
cc_167 VPB GCLK 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_168 VPB N_GCLK_c_1049_n 0.00122468f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_169 N_SCE_c_169_n N_GATE_c_201_n 0.0256071f $X=0.402 $Y=1.778 $X2=-0.19
+ $Y2=-0.245
cc_170 N_SCE_c_174_n N_GATE_c_201_n 0.0523461f $X=0.495 $Y=2.045 $X2=-0.19
+ $Y2=-0.245
cc_171 N_SCE_c_172_n N_GATE_c_201_n 0.00108715f $X=0.385 $Y=1.455 $X2=-0.19
+ $Y2=-0.245
cc_172 N_SCE_M1011_g N_GATE_M1009_g 0.020509f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_173 N_SCE_c_171_n N_GATE_M1009_g 0.0168557f $X=0.385 $Y=1.455 $X2=0 $Y2=0
cc_174 N_SCE_c_172_n N_GATE_M1009_g 0.00149764f $X=0.385 $Y=1.455 $X2=0 $Y2=0
cc_175 N_SCE_c_169_n N_GATE_c_203_n 0.00177127f $X=0.402 $Y=1.778 $X2=0 $Y2=0
cc_176 N_SCE_c_174_n N_GATE_c_203_n 0.00182484f $X=0.495 $Y=2.045 $X2=0 $Y2=0
cc_177 N_SCE_c_172_n N_GATE_c_203_n 0.0194621f $X=0.385 $Y=1.455 $X2=0 $Y2=0
cc_178 N_SCE_c_169_n N_VPWR_c_855_n 0.00483851f $X=0.402 $Y=1.778 $X2=0 $Y2=0
cc_179 N_SCE_c_174_n N_VPWR_c_855_n 0.0215138f $X=0.495 $Y=2.045 $X2=0 $Y2=0
cc_180 N_SCE_c_172_n N_VPWR_c_855_n 0.0246573f $X=0.385 $Y=1.455 $X2=0 $Y2=0
cc_181 N_SCE_c_174_n N_VPWR_c_864_n 0.00413917f $X=0.495 $Y=2.045 $X2=0 $Y2=0
cc_182 N_SCE_c_174_n N_VPWR_c_853_n 0.00817239f $X=0.495 $Y=2.045 $X2=0 $Y2=0
cc_183 N_SCE_M1011_g N_A_114_112#_c_948_n 0.00819024f $X=0.495 $Y=0.835 $X2=0
+ $Y2=0
cc_184 N_SCE_c_171_n N_A_114_112#_c_948_n 0.00147346f $X=0.385 $Y=1.455 $X2=0
+ $Y2=0
cc_185 N_SCE_c_172_n N_A_114_112#_c_948_n 0.00895228f $X=0.385 $Y=1.455 $X2=0
+ $Y2=0
cc_186 N_SCE_M1011_g N_A_114_112#_c_963_n 0.00257503f $X=0.495 $Y=0.835 $X2=0
+ $Y2=0
cc_187 N_SCE_M1011_g N_A_114_112#_c_950_n 0.00333944f $X=0.495 $Y=0.835 $X2=0
+ $Y2=0
cc_188 N_SCE_c_174_n N_A_114_112#_c_958_n 0.00184503f $X=0.495 $Y=2.045 $X2=0
+ $Y2=0
cc_189 N_SCE_M1011_g N_VGND_c_1085_n 0.00819878f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_190 N_SCE_c_171_n N_VGND_c_1085_n 0.00386581f $X=0.385 $Y=1.455 $X2=0 $Y2=0
cc_191 N_SCE_c_172_n N_VGND_c_1085_n 0.0216167f $X=0.385 $Y=1.455 $X2=0 $Y2=0
cc_192 N_SCE_M1011_g N_VGND_c_1095_n 0.00432822f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_193 N_SCE_M1011_g N_VGND_c_1100_n 0.00487769f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_194 N_GATE_M1009_g N_A_318_74#_c_242_n 5.25064e-19 $X=0.925 $Y=0.835 $X2=0
+ $Y2=0
cc_195 N_GATE_M1009_g N_A_288_48#_c_323_n 0.024928f $X=0.925 $Y=0.835 $X2=0
+ $Y2=0
cc_196 N_GATE_c_201_n N_VPWR_c_855_n 0.003245f $X=0.885 $Y=2.045 $X2=0 $Y2=0
cc_197 N_GATE_c_201_n N_VPWR_c_856_n 0.0033262f $X=0.885 $Y=2.045 $X2=0 $Y2=0
cc_198 N_GATE_c_201_n N_VPWR_c_864_n 0.00445602f $X=0.885 $Y=2.045 $X2=0 $Y2=0
cc_199 N_GATE_c_201_n N_VPWR_c_853_n 0.00862666f $X=0.885 $Y=2.045 $X2=0 $Y2=0
cc_200 N_GATE_c_203_n N_A_114_112#_M1000_d 0.00255236f $X=0.96 $Y=1.795 $X2=0
+ $Y2=0
cc_201 N_GATE_c_201_n N_A_114_112#_c_948_n 4.06408e-19 $X=0.885 $Y=2.045 $X2=0
+ $Y2=0
cc_202 N_GATE_M1009_g N_A_114_112#_c_948_n 0.0100761f $X=0.925 $Y=0.835 $X2=0
+ $Y2=0
cc_203 N_GATE_c_203_n N_A_114_112#_c_948_n 0.00615564f $X=0.96 $Y=1.795 $X2=0
+ $Y2=0
cc_204 N_GATE_M1009_g N_A_114_112#_c_963_n 0.00513644f $X=0.925 $Y=0.835 $X2=0
+ $Y2=0
cc_205 N_GATE_M1009_g N_A_114_112#_c_949_n 0.00867681f $X=0.925 $Y=0.835 $X2=0
+ $Y2=0
cc_206 N_GATE_M1009_g N_A_114_112#_c_950_n 0.00231761f $X=0.925 $Y=0.835 $X2=0
+ $Y2=0
cc_207 N_GATE_c_201_n N_A_114_112#_c_951_n 8.19427e-19 $X=0.885 $Y=2.045 $X2=0
+ $Y2=0
cc_208 N_GATE_M1009_g N_A_114_112#_c_951_n 0.00909975f $X=0.925 $Y=0.835 $X2=0
+ $Y2=0
cc_209 N_GATE_c_203_n N_A_114_112#_c_951_n 0.025014f $X=0.96 $Y=1.795 $X2=0
+ $Y2=0
cc_210 N_GATE_c_203_n N_A_114_112#_c_954_n 0.00194498f $X=0.96 $Y=1.795 $X2=0
+ $Y2=0
cc_211 N_GATE_c_201_n N_A_114_112#_c_952_n 0.00495471f $X=0.885 $Y=2.045 $X2=0
+ $Y2=0
cc_212 N_GATE_M1009_g N_A_114_112#_c_952_n 0.00596863f $X=0.925 $Y=0.835 $X2=0
+ $Y2=0
cc_213 N_GATE_c_203_n N_A_114_112#_c_952_n 0.0426646f $X=0.96 $Y=1.795 $X2=0
+ $Y2=0
cc_214 N_GATE_c_201_n N_A_114_112#_c_958_n 0.0124987f $X=0.885 $Y=2.045 $X2=0
+ $Y2=0
cc_215 N_GATE_c_203_n N_A_114_112#_c_958_n 0.0240594f $X=0.96 $Y=1.795 $X2=0
+ $Y2=0
cc_216 N_GATE_M1009_g N_VGND_c_1095_n 0.0034063f $X=0.925 $Y=0.835 $X2=0 $Y2=0
cc_217 N_GATE_M1009_g N_VGND_c_1100_n 0.00487769f $X=0.925 $Y=0.835 $X2=0 $Y2=0
cc_218 N_A_318_74#_c_240_n N_A_288_48#_c_323_n 0.00317258f $X=1.895 $Y=1.545
+ $X2=0 $Y2=0
cc_219 N_A_318_74#_c_242_n N_A_288_48#_c_323_n 0.00411406f $X=1.895 $Y=0.965
+ $X2=0 $Y2=0
cc_220 N_A_318_74#_c_240_n N_A_288_48#_c_324_n 0.00469377f $X=1.895 $Y=1.545
+ $X2=0 $Y2=0
cc_221 N_A_318_74#_c_242_n N_A_288_48#_c_324_n 0.00535989f $X=1.895 $Y=0.965
+ $X2=0 $Y2=0
cc_222 N_A_318_74#_c_243_n N_A_288_48#_c_324_n 2.27576e-19 $X=2.34 $Y=1.847
+ $X2=0 $Y2=0
cc_223 N_A_318_74#_c_240_n N_A_288_48#_c_326_n 0.0120541f $X=1.895 $Y=1.545
+ $X2=0 $Y2=0
cc_224 N_A_318_74#_c_243_n N_A_288_48#_c_326_n 0.00984101f $X=2.34 $Y=1.847
+ $X2=0 $Y2=0
cc_225 N_A_318_74#_c_244_n N_A_288_48#_c_326_n 8.85889e-19 $X=2.855 $Y=1.55
+ $X2=0 $Y2=0
cc_226 N_A_318_74#_c_245_n N_A_288_48#_c_326_n 0.00541276f $X=2.94 $Y=1.507
+ $X2=0 $Y2=0
cc_227 N_A_318_74#_c_243_n N_A_288_48#_c_345_n 0.00530675f $X=2.34 $Y=1.847
+ $X2=0 $Y2=0
cc_228 N_A_318_74#_c_243_n N_A_288_48#_M1003_g 0.0149207f $X=2.34 $Y=1.847 $X2=0
+ $Y2=0
cc_229 N_A_318_74#_c_246_n N_A_288_48#_c_347_n 0.0103572f $X=2.94 $Y=1.82 $X2=0
+ $Y2=0
cc_230 N_A_318_74#_c_241_n N_A_288_48#_c_327_n 0.00115318f $X=2.69 $Y=1.63 $X2=0
+ $Y2=0
cc_231 N_A_318_74#_c_244_n N_A_288_48#_c_327_n 0.00135102f $X=2.855 $Y=1.55
+ $X2=0 $Y2=0
cc_232 N_A_318_74#_c_245_n N_A_288_48#_c_327_n 0.0116193f $X=2.94 $Y=1.507 $X2=0
+ $Y2=0
cc_233 N_A_318_74#_c_240_n N_A_288_48#_c_328_n 0.00644266f $X=1.895 $Y=1.545
+ $X2=0 $Y2=0
cc_234 N_A_318_74#_c_242_n N_A_288_48#_c_328_n 6.5359e-19 $X=1.895 $Y=0.965
+ $X2=0 $Y2=0
cc_235 N_A_318_74#_c_243_n N_A_288_48#_c_328_n 0.00740977f $X=2.34 $Y=1.847
+ $X2=0 $Y2=0
cc_236 N_A_318_74#_c_245_n N_A_288_48#_c_328_n 0.00214647f $X=2.94 $Y=1.507
+ $X2=0 $Y2=0
cc_237 N_A_318_74#_M1019_g N_A_288_48#_c_329_n 0.0202664f $X=3.35 $Y=0.615 $X2=0
+ $Y2=0
cc_238 N_A_318_74#_c_246_n N_A_288_48#_c_349_n 0.00467581f $X=2.94 $Y=1.82 $X2=0
+ $Y2=0
cc_239 N_A_318_74#_c_246_n N_A_288_48#_c_351_n 0.0106814f $X=2.94 $Y=1.82 $X2=0
+ $Y2=0
cc_240 N_A_318_74#_c_242_n N_A_288_48#_c_330_n 0.00502799f $X=1.895 $Y=0.965
+ $X2=0 $Y2=0
cc_241 N_A_318_74#_M1019_g N_A_288_48#_c_331_n 0.0119709f $X=3.35 $Y=0.615 $X2=0
+ $Y2=0
cc_242 N_A_318_74#_M1019_g N_A_288_48#_c_333_n 0.00550364f $X=3.35 $Y=0.615
+ $X2=0 $Y2=0
cc_243 N_A_318_74#_M1019_g N_A_288_48#_c_335_n 0.00115488f $X=3.35 $Y=0.615
+ $X2=0 $Y2=0
cc_244 N_A_318_74#_M1019_g N_A_288_48#_c_339_n 3.86166e-19 $X=3.35 $Y=0.615
+ $X2=0 $Y2=0
cc_245 N_A_318_74#_c_240_n N_A_288_48#_c_339_n 0.023335f $X=1.895 $Y=1.545 $X2=0
+ $Y2=0
cc_246 N_A_318_74#_c_241_n N_A_288_48#_c_339_n 0.0104963f $X=2.69 $Y=1.63 $X2=0
+ $Y2=0
cc_247 N_A_318_74#_c_242_n N_A_288_48#_c_339_n 0.00160791f $X=1.895 $Y=0.965
+ $X2=0 $Y2=0
cc_248 N_A_318_74#_c_243_n N_A_288_48#_c_339_n 0.0247748f $X=2.34 $Y=1.847 $X2=0
+ $Y2=0
cc_249 N_A_318_74#_c_244_n N_A_288_48#_c_339_n 0.00190778f $X=2.855 $Y=1.55
+ $X2=0 $Y2=0
cc_250 N_A_318_74#_c_245_n N_A_288_48#_c_339_n 9.77176e-19 $X=2.94 $Y=1.507
+ $X2=0 $Y2=0
cc_251 N_A_318_74#_M1019_g N_A_706_317#_M1020_g 0.0547363f $X=3.35 $Y=0.615
+ $X2=0 $Y2=0
cc_252 N_A_318_74#_c_245_n N_A_706_317#_M1020_g 0.00691964f $X=2.94 $Y=1.507
+ $X2=0 $Y2=0
cc_253 N_A_318_74#_c_246_n N_A_706_317#_c_501_n 0.00146761f $X=2.94 $Y=1.82
+ $X2=0 $Y2=0
cc_254 N_A_318_74#_c_245_n N_A_706_317#_c_501_n 0.00871293f $X=2.94 $Y=1.507
+ $X2=0 $Y2=0
cc_255 N_A_318_74#_M1019_g N_A_580_74#_c_636_n 0.00840926f $X=3.35 $Y=0.615
+ $X2=0 $Y2=0
cc_256 N_A_318_74#_c_244_n N_A_580_74#_c_636_n 0.00316115f $X=2.855 $Y=1.55
+ $X2=0 $Y2=0
cc_257 N_A_318_74#_c_245_n N_A_580_74#_c_636_n 0.00539885f $X=2.94 $Y=1.507
+ $X2=0 $Y2=0
cc_258 N_A_318_74#_M1019_g N_A_580_74#_c_628_n 0.00883344f $X=3.35 $Y=0.615
+ $X2=0 $Y2=0
cc_259 N_A_318_74#_c_245_n N_A_580_74#_c_628_n 0.00508821f $X=2.94 $Y=1.507
+ $X2=0 $Y2=0
cc_260 N_A_318_74#_c_245_n N_A_580_74#_c_629_n 0.00543726f $X=2.94 $Y=1.507
+ $X2=0 $Y2=0
cc_261 N_A_318_74#_c_246_n N_A_580_74#_c_633_n 0.00644362f $X=2.94 $Y=1.82 $X2=0
+ $Y2=0
cc_262 N_A_318_74#_c_244_n N_A_580_74#_c_633_n 4.94403e-19 $X=2.855 $Y=1.55
+ $X2=0 $Y2=0
cc_263 N_A_318_74#_c_245_n N_A_580_74#_c_633_n 0.00410958f $X=2.94 $Y=1.507
+ $X2=0 $Y2=0
cc_264 N_A_318_74#_c_246_n N_A_580_74#_c_630_n 0.00723476f $X=2.94 $Y=1.82 $X2=0
+ $Y2=0
cc_265 N_A_318_74#_c_244_n N_A_580_74#_c_630_n 0.0213899f $X=2.855 $Y=1.55 $X2=0
+ $Y2=0
cc_266 N_A_318_74#_c_245_n N_A_580_74#_c_630_n 0.0135532f $X=2.94 $Y=1.507 $X2=0
+ $Y2=0
cc_267 N_A_318_74#_c_244_n N_A_580_74#_c_648_n 0.00239474f $X=2.855 $Y=1.55
+ $X2=0 $Y2=0
cc_268 N_A_318_74#_c_245_n N_A_580_74#_c_648_n 0.0116105f $X=2.94 $Y=1.507 $X2=0
+ $Y2=0
cc_269 N_A_318_74#_c_243_n N_VPWR_M1003_s 0.00331237f $X=2.34 $Y=1.847 $X2=0
+ $Y2=0
cc_270 N_A_318_74#_c_246_n N_VPWR_c_853_n 9.39239e-19 $X=2.94 $Y=1.82 $X2=0
+ $Y2=0
cc_271 N_A_318_74#_c_242_n N_A_114_112#_c_948_n 0.00245013f $X=1.895 $Y=0.965
+ $X2=0 $Y2=0
cc_272 N_A_318_74#_c_242_n N_A_114_112#_c_963_n 0.00161039f $X=1.895 $Y=0.965
+ $X2=0 $Y2=0
cc_273 N_A_318_74#_M1002_d N_A_114_112#_c_949_n 0.00669515f $X=1.59 $Y=0.37
+ $X2=0 $Y2=0
cc_274 N_A_318_74#_c_242_n N_A_114_112#_c_949_n 0.0261275f $X=1.895 $Y=0.965
+ $X2=0 $Y2=0
cc_275 N_A_318_74#_c_240_n N_A_114_112#_c_951_n 0.0131979f $X=1.895 $Y=1.545
+ $X2=0 $Y2=0
cc_276 N_A_318_74#_c_242_n N_A_114_112#_c_951_n 0.00393441f $X=1.895 $Y=0.965
+ $X2=0 $Y2=0
cc_277 N_A_318_74#_c_240_n N_A_114_112#_c_952_n 0.0116322f $X=1.895 $Y=1.545
+ $X2=0 $Y2=0
cc_278 N_A_318_74#_c_243_n N_A_114_112#_c_952_n 0.0492499f $X=2.34 $Y=1.847
+ $X2=0 $Y2=0
cc_279 N_A_318_74#_M1003_d N_A_114_112#_c_956_n 0.00594176f $X=2.025 $Y=1.84
+ $X2=0 $Y2=0
cc_280 N_A_318_74#_c_246_n N_A_114_112#_c_956_n 0.00453229f $X=2.94 $Y=1.82
+ $X2=0 $Y2=0
cc_281 N_A_318_74#_c_241_n N_A_114_112#_c_956_n 0.00650951f $X=2.69 $Y=1.63
+ $X2=0 $Y2=0
cc_282 N_A_318_74#_c_243_n N_A_114_112#_c_956_n 0.0326456f $X=2.34 $Y=1.847
+ $X2=0 $Y2=0
cc_283 N_A_318_74#_c_246_n N_A_114_112#_c_957_n 0.00406223f $X=2.94 $Y=1.82
+ $X2=0 $Y2=0
cc_284 N_A_318_74#_c_241_n N_A_114_112#_c_957_n 0.01174f $X=2.69 $Y=1.63 $X2=0
+ $Y2=0
cc_285 N_A_318_74#_c_243_n N_A_114_112#_c_957_n 0.0193405f $X=2.34 $Y=1.847
+ $X2=0 $Y2=0
cc_286 N_A_318_74#_c_244_n N_A_114_112#_c_957_n 0.00915244f $X=2.855 $Y=1.55
+ $X2=0 $Y2=0
cc_287 N_A_318_74#_c_245_n N_A_114_112#_c_957_n 8.54792e-19 $X=2.94 $Y=1.507
+ $X2=0 $Y2=0
cc_288 N_A_318_74#_M1019_g N_VGND_c_1091_n 9.15902e-19 $X=3.35 $Y=0.615 $X2=0
+ $Y2=0
cc_289 N_A_288_48#_c_336_n N_A_706_317#_M1001_d 0.00253411f $X=4.995 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_290 N_A_288_48#_c_331_n N_A_706_317#_M1020_g 0.00371294f $X=3.53 $Y=0.34
+ $X2=0 $Y2=0
cc_291 N_A_288_48#_c_333_n N_A_706_317#_M1020_g 0.00954024f $X=3.615 $Y=0.905
+ $X2=0 $Y2=0
cc_292 N_A_288_48#_c_334_n N_A_706_317#_M1020_g 0.0112741f $X=4.21 $Y=0.99 $X2=0
+ $Y2=0
cc_293 N_A_288_48#_c_335_n N_A_706_317#_M1020_g 0.00209968f $X=3.7 $Y=0.99 $X2=0
+ $Y2=0
cc_294 N_A_288_48#_c_393_p N_A_706_317#_M1020_g 0.00167035f $X=4.295 $Y=0.905
+ $X2=0 $Y2=0
cc_295 N_A_288_48#_c_349_n N_A_706_317#_c_503_n 0.00322812f $X=3.465 $Y=2.84
+ $X2=0 $Y2=0
cc_296 N_A_288_48#_c_351_n N_A_706_317#_c_503_n 0.0316012f $X=3.465 $Y=2.75
+ $X2=0 $Y2=0
cc_297 N_A_288_48#_c_352_n N_A_706_317#_c_506_n 0.0104522f $X=5.145 $Y=1.885
+ $X2=0 $Y2=0
cc_298 N_A_288_48#_c_336_n N_A_706_317#_c_494_n 0.0206246f $X=4.995 $Y=0.34
+ $X2=0 $Y2=0
cc_299 N_A_288_48#_c_338_n N_A_706_317#_c_494_n 0.0307524f $X=5.195 $Y=0.515
+ $X2=0 $Y2=0
cc_300 N_A_288_48#_c_341_n N_A_706_317#_c_495_n 0.0307524f $X=5.152 $Y=1.72
+ $X2=0 $Y2=0
cc_301 N_A_288_48#_M1013_s N_A_706_317#_c_509_n 0.0120995f $X=5.01 $Y=1.74 $X2=0
+ $Y2=0
cc_302 N_A_288_48#_c_352_n N_A_706_317#_c_509_n 0.0203663f $X=5.145 $Y=1.885
+ $X2=0 $Y2=0
cc_303 N_A_288_48#_c_352_n N_A_706_317#_c_496_n 0.00931677f $X=5.145 $Y=1.885
+ $X2=0 $Y2=0
cc_304 N_A_288_48#_c_341_n N_A_706_317#_c_496_n 9.85866e-19 $X=5.152 $Y=1.72
+ $X2=0 $Y2=0
cc_305 N_A_288_48#_c_341_n N_A_706_317#_c_497_n 0.00218999f $X=5.152 $Y=1.72
+ $X2=0 $Y2=0
cc_306 N_A_288_48#_c_351_n N_A_706_317#_c_499_n 2.08922e-19 $X=3.465 $Y=2.75
+ $X2=0 $Y2=0
cc_307 N_A_288_48#_c_352_n N_A_706_317#_c_512_n 0.0149884f $X=5.145 $Y=1.885
+ $X2=0 $Y2=0
cc_308 N_A_288_48#_c_340_n N_A_706_317#_c_500_n 0.0307524f $X=5.177 $Y=1.01
+ $X2=0 $Y2=0
cc_309 N_A_288_48#_c_351_n N_A_706_317#_c_501_n 6.78356e-19 $X=3.465 $Y=2.75
+ $X2=0 $Y2=0
cc_310 N_A_288_48#_c_331_n N_A_580_74#_M1022_d 0.00281472f $X=3.53 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_311 N_A_288_48#_c_334_n N_A_580_74#_c_626_n 0.00123256f $X=4.21 $Y=0.99 $X2=0
+ $Y2=0
cc_312 N_A_288_48#_c_352_n N_A_580_74#_c_626_n 4.31891e-19 $X=5.145 $Y=1.885
+ $X2=0 $Y2=0
cc_313 N_A_288_48#_c_341_n N_A_580_74#_c_626_n 6.29272e-19 $X=5.152 $Y=1.72
+ $X2=0 $Y2=0
cc_314 N_A_288_48#_c_333_n N_A_580_74#_c_627_n 2.03258e-19 $X=3.615 $Y=0.905
+ $X2=0 $Y2=0
cc_315 N_A_288_48#_c_334_n N_A_580_74#_c_627_n 0.00554025f $X=4.21 $Y=0.99 $X2=0
+ $Y2=0
cc_316 N_A_288_48#_c_393_p N_A_580_74#_c_627_n 0.0128024f $X=4.295 $Y=0.905
+ $X2=0 $Y2=0
cc_317 N_A_288_48#_c_336_n N_A_580_74#_c_627_n 0.011853f $X=4.995 $Y=0.34 $X2=0
+ $Y2=0
cc_318 N_A_288_48#_c_337_n N_A_580_74#_c_627_n 0.00273646f $X=4.38 $Y=0.34 $X2=0
+ $Y2=0
cc_319 N_A_288_48#_c_338_n N_A_580_74#_c_627_n 0.00468553f $X=5.195 $Y=0.515
+ $X2=0 $Y2=0
cc_320 N_A_288_48#_c_329_n N_A_580_74#_c_636_n 0.00294277f $X=2.825 $Y=0.995
+ $X2=0 $Y2=0
cc_321 N_A_288_48#_c_331_n N_A_580_74#_c_636_n 0.0254752f $X=3.53 $Y=0.34 $X2=0
+ $Y2=0
cc_322 N_A_288_48#_c_333_n N_A_580_74#_c_636_n 0.0191208f $X=3.615 $Y=0.905
+ $X2=0 $Y2=0
cc_323 N_A_288_48#_c_329_n N_A_580_74#_c_628_n 0.0024498f $X=2.825 $Y=0.995
+ $X2=0 $Y2=0
cc_324 N_A_288_48#_c_330_n N_A_580_74#_c_628_n 0.0051404f $X=2.63 $Y=1.03 $X2=0
+ $Y2=0
cc_325 N_A_288_48#_c_333_n N_A_580_74#_c_628_n 0.00421956f $X=3.615 $Y=0.905
+ $X2=0 $Y2=0
cc_326 N_A_288_48#_c_335_n N_A_580_74#_c_628_n 0.0137149f $X=3.7 $Y=0.99 $X2=0
+ $Y2=0
cc_327 N_A_288_48#_c_339_n N_A_580_74#_c_628_n 0.00638342f $X=2.315 $Y=1.195
+ $X2=0 $Y2=0
cc_328 N_A_288_48#_c_334_n N_A_580_74#_c_629_n 0.0332831f $X=4.21 $Y=0.99 $X2=0
+ $Y2=0
cc_329 N_A_288_48#_c_335_n N_A_580_74#_c_629_n 0.0140682f $X=3.7 $Y=0.99 $X2=0
+ $Y2=0
cc_330 N_A_288_48#_c_347_n N_A_580_74#_c_633_n 0.00487059f $X=3.375 $Y=3.15
+ $X2=0 $Y2=0
cc_331 N_A_288_48#_c_351_n N_A_580_74#_c_630_n 0.00461193f $X=3.465 $Y=2.75
+ $X2=0 $Y2=0
cc_332 N_A_288_48#_c_334_n N_A_580_74#_c_631_n 0.0162324f $X=4.21 $Y=0.99 $X2=0
+ $Y2=0
cc_333 N_A_288_48#_c_352_n N_CLK_c_715_n 0.00685155f $X=5.145 $Y=1.885 $X2=-0.19
+ $Y2=-0.245
cc_334 N_A_288_48#_c_336_n N_CLK_c_710_n 0.00462641f $X=4.995 $Y=0.34 $X2=0
+ $Y2=0
cc_335 N_A_288_48#_c_338_n N_CLK_c_710_n 0.00451642f $X=5.195 $Y=0.515 $X2=0
+ $Y2=0
cc_336 N_A_288_48#_c_340_n N_CLK_c_710_n 0.00219347f $X=5.177 $Y=1.01 $X2=0
+ $Y2=0
cc_337 N_A_288_48#_c_341_n N_CLK_c_710_n 0.00401029f $X=5.152 $Y=1.72 $X2=0
+ $Y2=0
cc_338 N_A_288_48#_c_352_n N_CLK_c_711_n 7.12948e-19 $X=5.145 $Y=1.885 $X2=0
+ $Y2=0
cc_339 N_A_288_48#_c_341_n N_CLK_c_711_n 0.0123032f $X=5.152 $Y=1.72 $X2=0 $Y2=0
cc_340 N_A_288_48#_c_352_n N_CLK_c_718_n 9.78534e-19 $X=5.145 $Y=1.885 $X2=0
+ $Y2=0
cc_341 N_A_288_48#_c_340_n CLK 0.00186086f $X=5.177 $Y=1.01 $X2=0 $Y2=0
cc_342 N_A_288_48#_c_341_n CLK 0.0277686f $X=5.152 $Y=1.72 $X2=0 $Y2=0
cc_343 N_A_288_48#_c_343_n N_VPWR_c_856_n 0.0197695f $X=1.95 $Y=2.845 $X2=0
+ $Y2=0
cc_344 N_A_288_48#_M1003_g N_VPWR_c_856_n 0.00395406f $X=1.95 $Y=2.26 $X2=0
+ $Y2=0
cc_345 N_A_288_48#_c_349_n N_VPWR_c_857_n 0.0105483f $X=3.465 $Y=2.84 $X2=0
+ $Y2=0
cc_346 N_A_288_48#_c_348_n N_VPWR_c_865_n 0.0550819f $X=2.04 $Y=3.15 $X2=0 $Y2=0
cc_347 N_A_288_48#_c_347_n N_VPWR_c_853_n 0.0536609f $X=3.375 $Y=3.15 $X2=0
+ $Y2=0
cc_348 N_A_288_48#_c_348_n N_VPWR_c_853_n 0.0079125f $X=2.04 $Y=3.15 $X2=0 $Y2=0
cc_349 N_A_288_48#_c_330_n N_A_114_112#_M1022_s 0.0122448f $X=2.63 $Y=1.03 $X2=0
+ $Y2=0
cc_350 N_A_288_48#_c_332_n N_A_114_112#_M1022_s 6.86248e-19 $X=2.715 $Y=0.34
+ $X2=0 $Y2=0
cc_351 N_A_288_48#_c_323_n N_A_114_112#_c_948_n 0.00112866f $X=1.515 $Y=1.21
+ $X2=0 $Y2=0
cc_352 N_A_288_48#_c_323_n N_A_114_112#_c_963_n 0.00100301f $X=1.515 $Y=1.21
+ $X2=0 $Y2=0
cc_353 N_A_288_48#_c_323_n N_A_114_112#_c_949_n 0.0150312f $X=1.515 $Y=1.21
+ $X2=0 $Y2=0
cc_354 N_A_288_48#_c_328_n N_A_114_112#_c_949_n 0.00224989f $X=2.48 $Y=1.07
+ $X2=0 $Y2=0
cc_355 N_A_288_48#_c_324_n N_A_114_112#_c_951_n 0.00461745f $X=1.86 $Y=1.285
+ $X2=0 $Y2=0
cc_356 N_A_288_48#_c_325_n N_A_114_112#_c_951_n 0.011085f $X=1.59 $Y=1.285 $X2=0
+ $Y2=0
cc_357 N_A_288_48#_c_326_n N_A_114_112#_c_951_n 2.05828e-19 $X=1.95 $Y=1.675
+ $X2=0 $Y2=0
cc_358 N_A_288_48#_c_326_n N_A_114_112#_c_952_n 0.00231661f $X=1.95 $Y=1.675
+ $X2=0 $Y2=0
cc_359 N_A_288_48#_M1003_g N_A_114_112#_c_952_n 0.00774134f $X=1.95 $Y=2.26
+ $X2=0 $Y2=0
cc_360 N_A_288_48#_M1003_g N_A_114_112#_c_956_n 0.0226838f $X=1.95 $Y=2.26 $X2=0
+ $Y2=0
cc_361 N_A_288_48#_c_347_n N_A_114_112#_c_956_n 0.0144075f $X=3.375 $Y=3.15
+ $X2=0 $Y2=0
cc_362 N_A_288_48#_M1003_g N_A_114_112#_c_957_n 0.0038542f $X=1.95 $Y=2.26 $X2=0
+ $Y2=0
cc_363 N_A_288_48#_M1003_g N_A_114_112#_c_958_n 0.00415884f $X=1.95 $Y=2.26
+ $X2=0 $Y2=0
cc_364 N_A_288_48#_c_323_n N_A_114_112#_c_953_n 0.00504475f $X=1.515 $Y=1.21
+ $X2=0 $Y2=0
cc_365 N_A_288_48#_c_328_n N_A_114_112#_c_953_n 0.00493278f $X=2.48 $Y=1.07
+ $X2=0 $Y2=0
cc_366 N_A_288_48#_c_329_n N_A_114_112#_c_953_n 8.15455e-19 $X=2.825 $Y=0.995
+ $X2=0 $Y2=0
cc_367 N_A_288_48#_c_330_n N_A_114_112#_c_953_n 0.0212796f $X=2.63 $Y=1.03 $X2=0
+ $Y2=0
cc_368 N_A_288_48#_c_332_n N_A_114_112#_c_953_n 0.00632876f $X=2.715 $Y=0.34
+ $X2=0 $Y2=0
cc_369 N_A_288_48#_c_339_n N_A_114_112#_c_953_n 0.0108433f $X=2.315 $Y=1.195
+ $X2=0 $Y2=0
cc_370 N_A_288_48#_c_334_n N_VGND_M1020_d 0.00676444f $X=4.21 $Y=0.99 $X2=0
+ $Y2=0
cc_371 N_A_288_48#_c_393_p N_VGND_M1020_d 0.00511615f $X=4.295 $Y=0.905 $X2=0
+ $Y2=0
cc_372 N_A_288_48#_c_331_n N_VGND_c_1086_n 0.0128817f $X=3.53 $Y=0.34 $X2=0
+ $Y2=0
cc_373 N_A_288_48#_c_334_n N_VGND_c_1086_n 0.013847f $X=4.21 $Y=0.99 $X2=0 $Y2=0
cc_374 N_A_288_48#_c_393_p N_VGND_c_1086_n 0.0224799f $X=4.295 $Y=0.905 $X2=0
+ $Y2=0
cc_375 N_A_288_48#_c_337_n N_VGND_c_1086_n 0.0142952f $X=4.38 $Y=0.34 $X2=0
+ $Y2=0
cc_376 N_A_288_48#_c_336_n N_VGND_c_1087_n 0.011924f $X=4.995 $Y=0.34 $X2=0
+ $Y2=0
cc_377 N_A_288_48#_c_323_n N_VGND_c_1091_n 0.00315544f $X=1.515 $Y=1.21 $X2=0
+ $Y2=0
cc_378 N_A_288_48#_c_329_n N_VGND_c_1091_n 0.00278271f $X=2.825 $Y=0.995 $X2=0
+ $Y2=0
cc_379 N_A_288_48#_c_331_n N_VGND_c_1091_n 0.0641927f $X=3.53 $Y=0.34 $X2=0
+ $Y2=0
cc_380 N_A_288_48#_c_332_n N_VGND_c_1091_n 0.0121867f $X=2.715 $Y=0.34 $X2=0
+ $Y2=0
cc_381 N_A_288_48#_c_336_n N_VGND_c_1093_n 0.0656368f $X=4.995 $Y=0.34 $X2=0
+ $Y2=0
cc_382 N_A_288_48#_c_337_n N_VGND_c_1093_n 0.0121867f $X=4.38 $Y=0.34 $X2=0
+ $Y2=0
cc_383 N_A_288_48#_c_323_n N_VGND_c_1098_n 0.00542971f $X=1.515 $Y=1.21 $X2=0
+ $Y2=0
cc_384 N_A_288_48#_c_323_n N_VGND_c_1100_n 0.00400711f $X=1.515 $Y=1.21 $X2=0
+ $Y2=0
cc_385 N_A_288_48#_c_329_n N_VGND_c_1100_n 0.00363426f $X=2.825 $Y=0.995 $X2=0
+ $Y2=0
cc_386 N_A_288_48#_c_331_n N_VGND_c_1100_n 0.0365608f $X=3.53 $Y=0.34 $X2=0
+ $Y2=0
cc_387 N_A_288_48#_c_332_n N_VGND_c_1100_n 0.00660921f $X=2.715 $Y=0.34 $X2=0
+ $Y2=0
cc_388 N_A_288_48#_c_336_n N_VGND_c_1100_n 0.0371906f $X=4.995 $Y=0.34 $X2=0
+ $Y2=0
cc_389 N_A_288_48#_c_337_n N_VGND_c_1100_n 0.00660921f $X=4.38 $Y=0.34 $X2=0
+ $Y2=0
cc_390 N_A_288_48#_c_331_n A_685_81# 0.00179331f $X=3.53 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_391 N_A_288_48#_c_333_n A_685_81# 0.00376627f $X=3.615 $Y=0.905 $X2=-0.19
+ $Y2=-0.245
cc_392 N_A_706_317#_M1020_g N_A_580_74#_c_626_n 0.012245f $X=3.74 $Y=0.615 $X2=0
+ $Y2=0
cc_393 N_A_706_317#_c_503_n N_A_580_74#_c_626_n 0.00826835f $X=3.855 $Y=2.18
+ $X2=0 $Y2=0
cc_394 N_A_706_317#_c_505_n N_A_580_74#_c_626_n 0.0136209f $X=4.44 $Y=1.84 $X2=0
+ $Y2=0
cc_395 N_A_706_317#_c_506_n N_A_580_74#_c_626_n 0.00501909f $X=4.632 $Y=2.22
+ $X2=0 $Y2=0
cc_396 N_A_706_317#_c_507_n N_A_580_74#_c_626_n 0.00658247f $X=4.605 $Y=2.755
+ $X2=0 $Y2=0
cc_397 N_A_706_317#_c_495_n N_A_580_74#_c_626_n 0.00412716f $X=4.74 $Y=1.755
+ $X2=0 $Y2=0
cc_398 N_A_706_317#_c_499_n N_A_580_74#_c_626_n 9.64431e-19 $X=3.695 $Y=1.75
+ $X2=0 $Y2=0
cc_399 N_A_706_317#_c_512_n N_A_580_74#_c_626_n 0.0020637f $X=4.632 $Y=1.84
+ $X2=0 $Y2=0
cc_400 N_A_706_317#_c_513_n N_A_580_74#_c_626_n 0.00175527f $X=4.632 $Y=2.305
+ $X2=0 $Y2=0
cc_401 N_A_706_317#_c_501_n N_A_580_74#_c_626_n 0.0187668f $X=3.855 $Y=1.75
+ $X2=0 $Y2=0
cc_402 N_A_706_317#_M1020_g N_A_580_74#_c_627_n 0.0154325f $X=3.74 $Y=0.615
+ $X2=0 $Y2=0
cc_403 N_A_706_317#_c_495_n N_A_580_74#_c_627_n 0.0118613f $X=4.74 $Y=1.755
+ $X2=0 $Y2=0
cc_404 N_A_706_317#_M1020_g N_A_580_74#_c_636_n 2.25119e-19 $X=3.74 $Y=0.615
+ $X2=0 $Y2=0
cc_405 N_A_706_317#_M1020_g N_A_580_74#_c_628_n 0.00116521f $X=3.74 $Y=0.615
+ $X2=0 $Y2=0
cc_406 N_A_706_317#_M1020_g N_A_580_74#_c_629_n 0.0107958f $X=3.74 $Y=0.615
+ $X2=0 $Y2=0
cc_407 N_A_706_317#_c_505_n N_A_580_74#_c_629_n 0.0134189f $X=4.44 $Y=1.84 $X2=0
+ $Y2=0
cc_408 N_A_706_317#_c_499_n N_A_580_74#_c_629_n 0.0242682f $X=3.695 $Y=1.75
+ $X2=0 $Y2=0
cc_409 N_A_706_317#_c_501_n N_A_580_74#_c_629_n 0.00367849f $X=3.855 $Y=1.75
+ $X2=0 $Y2=0
cc_410 N_A_706_317#_M1020_g N_A_580_74#_c_630_n 0.00310402f $X=3.74 $Y=0.615
+ $X2=0 $Y2=0
cc_411 N_A_706_317#_c_502_n N_A_580_74#_c_630_n 0.00530736f $X=3.855 $Y=2.09
+ $X2=0 $Y2=0
cc_412 N_A_706_317#_c_499_n N_A_580_74#_c_630_n 0.0255945f $X=3.695 $Y=1.75
+ $X2=0 $Y2=0
cc_413 N_A_706_317#_c_501_n N_A_580_74#_c_630_n 0.00260244f $X=3.855 $Y=1.75
+ $X2=0 $Y2=0
cc_414 N_A_706_317#_M1020_g N_A_580_74#_c_631_n 0.00113382f $X=3.74 $Y=0.615
+ $X2=0 $Y2=0
cc_415 N_A_706_317#_c_505_n N_A_580_74#_c_631_n 0.0209593f $X=4.44 $Y=1.84 $X2=0
+ $Y2=0
cc_416 N_A_706_317#_c_495_n N_A_580_74#_c_631_n 0.0255154f $X=4.74 $Y=1.755
+ $X2=0 $Y2=0
cc_417 N_A_706_317#_c_512_n N_A_580_74#_c_631_n 0.00366862f $X=4.632 $Y=1.84
+ $X2=0 $Y2=0
cc_418 N_A_706_317#_c_506_n N_CLK_c_715_n 0.00430514f $X=4.632 $Y=2.22 $X2=-0.19
+ $Y2=-0.245
cc_419 N_A_706_317#_c_507_n N_CLK_c_715_n 0.00881328f $X=4.605 $Y=2.755
+ $X2=-0.19 $Y2=-0.245
cc_420 N_A_706_317#_c_495_n N_CLK_c_715_n 8.01335e-19 $X=4.74 $Y=1.755 $X2=-0.19
+ $Y2=-0.245
cc_421 N_A_706_317#_c_509_n N_CLK_c_715_n 0.0194685f $X=5.835 $Y=2.305 $X2=-0.19
+ $Y2=-0.245
cc_422 N_A_706_317#_c_496_n N_CLK_c_715_n 0.00249924f $X=5.92 $Y=2.22 $X2=-0.19
+ $Y2=-0.245
cc_423 N_A_706_317#_c_494_n N_CLK_c_710_n 5.87969e-19 $X=4.635 $Y=0.835 $X2=0
+ $Y2=0
cc_424 N_A_706_317#_c_493_n N_CLK_c_711_n 0.042261f $X=6.565 $Y=1.795 $X2=0
+ $Y2=0
cc_425 N_A_706_317#_c_509_n N_CLK_c_711_n 0.00383202f $X=5.835 $Y=2.305 $X2=0
+ $Y2=0
cc_426 N_A_706_317#_c_497_n N_CLK_c_711_n 0.0171337f $X=6.005 $Y=1.465 $X2=0
+ $Y2=0
cc_427 N_A_706_317#_c_493_n N_CLK_c_712_n 0.00331227f $X=6.565 $Y=1.795 $X2=0
+ $Y2=0
cc_428 N_A_706_317#_c_496_n N_CLK_c_712_n 0.0026549f $X=5.92 $Y=2.22 $X2=0 $Y2=0
cc_429 N_A_706_317#_c_497_n N_CLK_c_712_n 0.0030238f $X=6.005 $Y=1.465 $X2=0
+ $Y2=0
cc_430 N_A_706_317#_c_493_n N_CLK_c_718_n 0.0126008f $X=6.565 $Y=1.795 $X2=0
+ $Y2=0
cc_431 N_A_706_317#_c_509_n N_CLK_c_718_n 0.0136085f $X=5.835 $Y=2.305 $X2=0
+ $Y2=0
cc_432 N_A_706_317#_c_496_n N_CLK_c_718_n 0.0179856f $X=5.92 $Y=2.22 $X2=0 $Y2=0
cc_433 N_A_706_317#_M1007_g N_CLK_c_713_n 0.042261f $X=6.275 $Y=0.74 $X2=0 $Y2=0
cc_434 N_A_706_317#_M1007_g CLK 2.78077e-19 $X=6.275 $Y=0.74 $X2=0 $Y2=0
cc_435 N_A_706_317#_c_509_n CLK 0.0072603f $X=5.835 $Y=2.305 $X2=0 $Y2=0
cc_436 N_A_706_317#_c_497_n CLK 0.0199911f $X=6.005 $Y=1.465 $X2=0 $Y2=0
cc_437 N_A_706_317#_c_493_n N_A_1195_374#_c_775_n 0.0238261f $X=6.565 $Y=1.795
+ $X2=0 $Y2=0
cc_438 N_A_706_317#_c_493_n N_A_1195_374#_c_777_n 0.0116766f $X=6.565 $Y=1.795
+ $X2=0 $Y2=0
cc_439 N_A_706_317#_M1007_g N_A_1195_374#_c_768_n 0.0115865f $X=6.275 $Y=0.74
+ $X2=0 $Y2=0
cc_440 N_A_706_317#_c_493_n N_A_1195_374#_c_778_n 0.0142722f $X=6.565 $Y=1.795
+ $X2=0 $Y2=0
cc_441 N_A_706_317#_c_498_n N_A_1195_374#_c_778_n 0.00175142f $X=6.365 $Y=1.465
+ $X2=0 $Y2=0
cc_442 N_A_706_317#_c_493_n N_A_1195_374#_c_779_n 0.00894315f $X=6.565 $Y=1.795
+ $X2=0 $Y2=0
cc_443 N_A_706_317#_c_496_n N_A_1195_374#_c_779_n 0.0103613f $X=5.92 $Y=2.22
+ $X2=0 $Y2=0
cc_444 N_A_706_317#_c_498_n N_A_1195_374#_c_779_n 0.0278654f $X=6.365 $Y=1.465
+ $X2=0 $Y2=0
cc_445 N_A_706_317#_M1007_g N_A_1195_374#_c_770_n 0.0038748f $X=6.275 $Y=0.74
+ $X2=0 $Y2=0
cc_446 N_A_706_317#_c_493_n N_A_1195_374#_c_770_n 0.00861575f $X=6.565 $Y=1.795
+ $X2=0 $Y2=0
cc_447 N_A_706_317#_c_498_n N_A_1195_374#_c_770_n 0.0171756f $X=6.365 $Y=1.465
+ $X2=0 $Y2=0
cc_448 N_A_706_317#_c_493_n N_A_1195_374#_c_772_n 0.00606655f $X=6.565 $Y=1.795
+ $X2=0 $Y2=0
cc_449 N_A_706_317#_c_498_n N_A_1195_374#_c_772_n 0.0164832f $X=6.365 $Y=1.465
+ $X2=0 $Y2=0
cc_450 N_A_706_317#_M1007_g N_A_1195_374#_c_773_n 0.00399952f $X=6.275 $Y=0.74
+ $X2=0 $Y2=0
cc_451 N_A_706_317#_c_493_n N_A_1195_374#_c_774_n 0.0209041f $X=6.565 $Y=1.795
+ $X2=0 $Y2=0
cc_452 N_A_706_317#_c_498_n N_A_1195_374#_c_774_n 3.30771e-19 $X=6.365 $Y=1.465
+ $X2=0 $Y2=0
cc_453 N_A_706_317#_c_505_n N_VPWR_M1012_d 0.00267141f $X=4.44 $Y=1.84 $X2=0
+ $Y2=0
cc_454 N_A_706_317#_c_509_n N_VPWR_M1013_d 0.00809063f $X=5.835 $Y=2.305 $X2=0
+ $Y2=0
cc_455 N_A_706_317#_c_503_n N_VPWR_c_857_n 0.0116652f $X=3.855 $Y=2.18 $X2=0
+ $Y2=0
cc_456 N_A_706_317#_c_505_n N_VPWR_c_857_n 0.0202669f $X=4.44 $Y=1.84 $X2=0
+ $Y2=0
cc_457 N_A_706_317#_c_506_n N_VPWR_c_857_n 0.00844596f $X=4.632 $Y=2.22 $X2=0
+ $Y2=0
cc_458 N_A_706_317#_c_507_n N_VPWR_c_857_n 0.0359497f $X=4.605 $Y=2.755 $X2=0
+ $Y2=0
cc_459 N_A_706_317#_c_513_n N_VPWR_c_857_n 0.0121024f $X=4.632 $Y=2.305 $X2=0
+ $Y2=0
cc_460 N_A_706_317#_c_493_n N_VPWR_c_858_n 5.74698e-19 $X=6.565 $Y=1.795 $X2=0
+ $Y2=0
cc_461 N_A_706_317#_c_509_n N_VPWR_c_858_n 0.0215947f $X=5.835 $Y=2.305 $X2=0
+ $Y2=0
cc_462 N_A_706_317#_c_493_n N_VPWR_c_859_n 0.0103799f $X=6.565 $Y=1.795 $X2=0
+ $Y2=0
cc_463 N_A_706_317#_c_493_n N_VPWR_c_862_n 0.00500894f $X=6.565 $Y=1.795 $X2=0
+ $Y2=0
cc_464 N_A_706_317#_c_503_n N_VPWR_c_865_n 0.00399858f $X=3.855 $Y=2.18 $X2=0
+ $Y2=0
cc_465 N_A_706_317#_c_507_n N_VPWR_c_866_n 0.0137199f $X=4.605 $Y=2.755 $X2=0
+ $Y2=0
cc_466 N_A_706_317#_c_503_n N_VPWR_c_853_n 0.0046122f $X=3.855 $Y=2.18 $X2=0
+ $Y2=0
cc_467 N_A_706_317#_c_493_n N_VPWR_c_853_n 0.00517496f $X=6.565 $Y=1.795 $X2=0
+ $Y2=0
cc_468 N_A_706_317#_c_507_n N_VPWR_c_853_n 0.0136092f $X=4.605 $Y=2.755 $X2=0
+ $Y2=0
cc_469 N_A_706_317#_c_493_n GCLK 0.00100924f $X=6.565 $Y=1.795 $X2=0 $Y2=0
cc_470 N_A_706_317#_M1020_g N_VGND_c_1086_n 0.0012897f $X=3.74 $Y=0.615 $X2=0
+ $Y2=0
cc_471 N_A_706_317#_M1007_g N_VGND_c_1087_n 0.00234521f $X=6.275 $Y=0.74 $X2=0
+ $Y2=0
cc_472 N_A_706_317#_c_497_n N_VGND_c_1087_n 0.00115537f $X=6.005 $Y=1.465 $X2=0
+ $Y2=0
cc_473 N_A_706_317#_M1007_g N_VGND_c_1088_n 0.00356081f $X=6.275 $Y=0.74 $X2=0
+ $Y2=0
cc_474 N_A_706_317#_M1020_g N_VGND_c_1091_n 0.00444804f $X=3.74 $Y=0.615 $X2=0
+ $Y2=0
cc_475 N_A_706_317#_M1007_g N_VGND_c_1096_n 0.00434272f $X=6.275 $Y=0.74 $X2=0
+ $Y2=0
cc_476 N_A_706_317#_M1020_g N_VGND_c_1100_n 0.00409911f $X=3.74 $Y=0.615 $X2=0
+ $Y2=0
cc_477 N_A_706_317#_M1007_g N_VGND_c_1100_n 0.00825669f $X=6.275 $Y=0.74 $X2=0
+ $Y2=0
cc_478 N_A_580_74#_c_626_n N_VPWR_c_857_n 0.00819892f $X=4.38 $Y=1.705 $X2=0
+ $Y2=0
cc_479 N_A_580_74#_c_630_n N_VPWR_c_857_n 0.0115204f $X=3.18 $Y=2.235 $X2=0
+ $Y2=0
cc_480 N_A_580_74#_c_633_n N_VPWR_c_865_n 0.00632793f $X=3.165 $Y=2.465 $X2=0
+ $Y2=0
cc_481 N_A_580_74#_c_626_n N_VPWR_c_866_n 0.00520623f $X=4.38 $Y=1.705 $X2=0
+ $Y2=0
cc_482 N_A_580_74#_c_626_n N_VPWR_c_853_n 0.00526787f $X=4.38 $Y=1.705 $X2=0
+ $Y2=0
cc_483 N_A_580_74#_c_633_n N_VPWR_c_853_n 0.0093378f $X=3.165 $Y=2.465 $X2=0
+ $Y2=0
cc_484 N_A_580_74#_c_633_n N_A_114_112#_c_956_n 0.0263549f $X=3.165 $Y=2.465
+ $X2=0 $Y2=0
cc_485 N_A_580_74#_c_633_n N_A_114_112#_c_957_n 0.00570278f $X=3.165 $Y=2.465
+ $X2=0 $Y2=0
cc_486 N_A_580_74#_c_630_n N_A_114_112#_c_957_n 0.0141982f $X=3.18 $Y=2.235
+ $X2=0 $Y2=0
cc_487 N_A_580_74#_c_627_n N_VGND_c_1086_n 0.00126464f $X=4.42 $Y=1.255 $X2=0
+ $Y2=0
cc_488 N_A_580_74#_c_627_n N_VGND_c_1093_n 9.34772e-19 $X=4.42 $Y=1.255 $X2=0
+ $Y2=0
cc_489 N_CLK_c_718_n N_A_1195_374#_c_777_n 0.0090769f $X=5.9 $Y=1.795 $X2=0
+ $Y2=0
cc_490 N_CLK_c_713_n N_A_1195_374#_c_768_n 0.0016642f $X=5.915 $Y=1.22 $X2=0
+ $Y2=0
cc_491 N_CLK_c_718_n N_A_1195_374#_c_779_n 7.38302e-19 $X=5.9 $Y=1.795 $X2=0
+ $Y2=0
cc_492 N_CLK_c_713_n N_A_1195_374#_c_770_n 7.31697e-19 $X=5.915 $Y=1.22 $X2=0
+ $Y2=0
cc_493 N_CLK_c_715_n N_VPWR_c_858_n 0.00420207f $X=5.37 $Y=1.665 $X2=0 $Y2=0
cc_494 N_CLK_c_718_n N_VPWR_c_858_n 0.00990608f $X=5.9 $Y=1.795 $X2=0 $Y2=0
cc_495 N_CLK_c_718_n N_VPWR_c_862_n 0.00461214f $X=5.9 $Y=1.795 $X2=0 $Y2=0
cc_496 N_CLK_c_715_n N_VPWR_c_866_n 0.00355139f $X=5.37 $Y=1.665 $X2=0 $Y2=0
cc_497 N_CLK_c_715_n N_VPWR_c_853_n 0.0043622f $X=5.37 $Y=1.665 $X2=0 $Y2=0
cc_498 N_CLK_c_718_n N_VPWR_c_853_n 0.00469196f $X=5.9 $Y=1.795 $X2=0 $Y2=0
cc_499 N_CLK_c_710_n N_VGND_c_1087_n 0.00475792f $X=5.41 $Y=1.22 $X2=0 $Y2=0
cc_500 N_CLK_c_711_n N_VGND_c_1087_n 0.00429275f $X=5.9 $Y=1.55 $X2=0 $Y2=0
cc_501 N_CLK_c_713_n N_VGND_c_1087_n 0.0147865f $X=5.915 $Y=1.22 $X2=0 $Y2=0
cc_502 CLK N_VGND_c_1087_n 0.0111858f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_503 N_CLK_c_710_n N_VGND_c_1093_n 0.00430908f $X=5.41 $Y=1.22 $X2=0 $Y2=0
cc_504 N_CLK_c_713_n N_VGND_c_1096_n 0.00398535f $X=5.915 $Y=1.22 $X2=0 $Y2=0
cc_505 N_CLK_c_710_n N_VGND_c_1100_n 0.00821159f $X=5.41 $Y=1.22 $X2=0 $Y2=0
cc_506 N_CLK_c_713_n N_VGND_c_1100_n 0.00786935f $X=5.915 $Y=1.22 $X2=0 $Y2=0
cc_507 N_A_1195_374#_c_778_n N_VPWR_M1010_d 0.00526636f $X=6.87 $Y=1.885 $X2=0
+ $Y2=0
cc_508 N_A_1195_374#_c_777_n N_VPWR_c_858_n 0.0152579f $X=6.34 $Y=2.015 $X2=0
+ $Y2=0
cc_509 N_A_1195_374#_c_775_n N_VPWR_c_859_n 0.00985112f $X=7.15 $Y=1.765 $X2=0
+ $Y2=0
cc_510 N_A_1195_374#_c_777_n N_VPWR_c_859_n 0.0504392f $X=6.34 $Y=2.015 $X2=0
+ $Y2=0
cc_511 N_A_1195_374#_c_778_n N_VPWR_c_859_n 0.0262435f $X=6.87 $Y=1.885 $X2=0
+ $Y2=0
cc_512 N_A_1195_374#_c_774_n N_VPWR_c_859_n 5.22182e-19 $X=7.6 $Y=1.532 $X2=0
+ $Y2=0
cc_513 N_A_1195_374#_c_776_n N_VPWR_c_861_n 0.00963415f $X=7.6 $Y=1.765 $X2=0
+ $Y2=0
cc_514 N_A_1195_374#_c_774_n N_VPWR_c_861_n 3.5215e-19 $X=7.6 $Y=1.532 $X2=0
+ $Y2=0
cc_515 N_A_1195_374#_c_777_n N_VPWR_c_862_n 0.0106883f $X=6.34 $Y=2.015 $X2=0
+ $Y2=0
cc_516 N_A_1195_374#_c_775_n N_VPWR_c_867_n 0.00445602f $X=7.15 $Y=1.765 $X2=0
+ $Y2=0
cc_517 N_A_1195_374#_c_776_n N_VPWR_c_867_n 0.00417277f $X=7.6 $Y=1.765 $X2=0
+ $Y2=0
cc_518 N_A_1195_374#_c_775_n N_VPWR_c_853_n 0.00861719f $X=7.15 $Y=1.765 $X2=0
+ $Y2=0
cc_519 N_A_1195_374#_c_776_n N_VPWR_c_853_n 0.00769535f $X=7.6 $Y=1.765 $X2=0
+ $Y2=0
cc_520 N_A_1195_374#_c_777_n N_VPWR_c_853_n 0.0114226f $X=6.34 $Y=2.015 $X2=0
+ $Y2=0
cc_521 N_A_1195_374#_M1005_g N_GCLK_c_1047_n 0.00969649f $X=7.245 $Y=0.74 $X2=0
+ $Y2=0
cc_522 N_A_1195_374#_M1016_g N_GCLK_c_1047_n 0.00788704f $X=7.675 $Y=0.74 $X2=0
+ $Y2=0
cc_523 N_A_1195_374#_c_768_n N_GCLK_c_1047_n 0.00490352f $X=6.49 $Y=0.515 $X2=0
+ $Y2=0
cc_524 N_A_1195_374#_c_769_n N_GCLK_c_1047_n 0.0103299f $X=6.87 $Y=1.045 $X2=0
+ $Y2=0
cc_525 N_A_1195_374#_M1005_g N_GCLK_c_1048_n 0.00351919f $X=7.245 $Y=0.74 $X2=0
+ $Y2=0
cc_526 N_A_1195_374#_M1016_g N_GCLK_c_1048_n 0.00327512f $X=7.675 $Y=0.74 $X2=0
+ $Y2=0
cc_527 N_A_1195_374#_c_775_n GCLK 0.00241662f $X=7.15 $Y=1.765 $X2=0 $Y2=0
cc_528 N_A_1195_374#_c_776_n GCLK 0.00233168f $X=7.6 $Y=1.765 $X2=0 $Y2=0
cc_529 N_A_1195_374#_c_778_n GCLK 0.00660441f $X=6.87 $Y=1.885 $X2=0 $Y2=0
cc_530 N_A_1195_374#_c_772_n GCLK 9.53215e-19 $X=7.06 $Y=1.465 $X2=0 $Y2=0
cc_531 N_A_1195_374#_c_774_n GCLK 0.00816244f $X=7.6 $Y=1.532 $X2=0 $Y2=0
cc_532 N_A_1195_374#_c_775_n GCLK 0.0119614f $X=7.15 $Y=1.765 $X2=0 $Y2=0
cc_533 N_A_1195_374#_c_776_n GCLK 0.0128557f $X=7.6 $Y=1.765 $X2=0 $Y2=0
cc_534 N_A_1195_374#_c_775_n N_GCLK_c_1049_n 4.20792e-19 $X=7.15 $Y=1.765 $X2=0
+ $Y2=0
cc_535 N_A_1195_374#_M1005_g N_GCLK_c_1049_n 0.00154761f $X=7.245 $Y=0.74 $X2=0
+ $Y2=0
cc_536 N_A_1195_374#_c_776_n N_GCLK_c_1049_n 0.00259359f $X=7.6 $Y=1.765 $X2=0
+ $Y2=0
cc_537 N_A_1195_374#_M1016_g N_GCLK_c_1049_n 0.00413752f $X=7.675 $Y=0.74 $X2=0
+ $Y2=0
cc_538 N_A_1195_374#_c_778_n N_GCLK_c_1049_n 9.86685e-19 $X=6.87 $Y=1.885 $X2=0
+ $Y2=0
cc_539 N_A_1195_374#_c_771_n N_GCLK_c_1049_n 0.00762026f $X=6.955 $Y=1.8 $X2=0
+ $Y2=0
cc_540 N_A_1195_374#_c_772_n N_GCLK_c_1049_n 0.0237053f $X=7.06 $Y=1.465 $X2=0
+ $Y2=0
cc_541 N_A_1195_374#_c_773_n N_GCLK_c_1049_n 0.00759747f $X=7.047 $Y=1.3 $X2=0
+ $Y2=0
cc_542 N_A_1195_374#_c_774_n N_GCLK_c_1049_n 0.0358033f $X=7.6 $Y=1.532 $X2=0
+ $Y2=0
cc_543 N_A_1195_374#_c_769_n N_VGND_M1005_s 0.00432991f $X=6.87 $Y=1.045 $X2=0
+ $Y2=0
cc_544 N_A_1195_374#_c_768_n N_VGND_c_1087_n 0.0202037f $X=6.49 $Y=0.515 $X2=0
+ $Y2=0
cc_545 N_A_1195_374#_c_770_n N_VGND_c_1087_n 0.001765f $X=6.655 $Y=1.045 $X2=0
+ $Y2=0
cc_546 N_A_1195_374#_M1005_g N_VGND_c_1088_n 0.00545557f $X=7.245 $Y=0.74 $X2=0
+ $Y2=0
cc_547 N_A_1195_374#_c_768_n N_VGND_c_1088_n 0.0309452f $X=6.49 $Y=0.515 $X2=0
+ $Y2=0
cc_548 N_A_1195_374#_c_769_n N_VGND_c_1088_n 0.0154159f $X=6.87 $Y=1.045 $X2=0
+ $Y2=0
cc_549 N_A_1195_374#_c_772_n N_VGND_c_1088_n 0.00258618f $X=7.06 $Y=1.465 $X2=0
+ $Y2=0
cc_550 N_A_1195_374#_c_774_n N_VGND_c_1088_n 0.00104582f $X=7.6 $Y=1.532 $X2=0
+ $Y2=0
cc_551 N_A_1195_374#_M1016_g N_VGND_c_1090_n 0.00647412f $X=7.675 $Y=0.74 $X2=0
+ $Y2=0
cc_552 N_A_1195_374#_c_768_n N_VGND_c_1096_n 0.0145639f $X=6.49 $Y=0.515 $X2=0
+ $Y2=0
cc_553 N_A_1195_374#_M1005_g N_VGND_c_1097_n 0.00434272f $X=7.245 $Y=0.74 $X2=0
+ $Y2=0
cc_554 N_A_1195_374#_M1016_g N_VGND_c_1097_n 0.00434272f $X=7.675 $Y=0.74 $X2=0
+ $Y2=0
cc_555 N_A_1195_374#_M1005_g N_VGND_c_1100_n 0.00825283f $X=7.245 $Y=0.74 $X2=0
+ $Y2=0
cc_556 N_A_1195_374#_M1016_g N_VGND_c_1100_n 0.00823907f $X=7.675 $Y=0.74 $X2=0
+ $Y2=0
cc_557 N_A_1195_374#_c_768_n N_VGND_c_1100_n 0.0119984f $X=6.49 $Y=0.515 $X2=0
+ $Y2=0
cc_558 N_VPWR_c_853_n N_A_114_112#_c_954_n 0.00670752f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_559 N_VPWR_M1003_s N_A_114_112#_c_952_n 0.00799893f $X=1.515 $Y=1.84 $X2=0
+ $Y2=0
cc_560 N_VPWR_M1003_s N_A_114_112#_c_956_n 0.00880783f $X=1.515 $Y=1.84 $X2=0
+ $Y2=0
cc_561 N_VPWR_c_856_n N_A_114_112#_c_956_n 0.0138115f $X=1.65 $Y=2.825 $X2=0
+ $Y2=0
cc_562 N_VPWR_c_865_n N_A_114_112#_c_956_n 0.00575553f $X=3.99 $Y=3.33 $X2=0
+ $Y2=0
cc_563 N_VPWR_c_853_n N_A_114_112#_c_956_n 0.0297748f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_564 N_VPWR_c_855_n N_A_114_112#_c_958_n 0.020489f $X=0.27 $Y=2.295 $X2=0
+ $Y2=0
cc_565 N_VPWR_c_856_n N_A_114_112#_c_958_n 0.0229788f $X=1.65 $Y=2.825 $X2=0
+ $Y2=0
cc_566 N_VPWR_c_864_n N_A_114_112#_c_958_n 0.0145621f $X=1.485 $Y=3.33 $X2=0
+ $Y2=0
cc_567 N_VPWR_c_853_n N_A_114_112#_c_958_n 0.0120343f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_568 N_VPWR_M1003_s N_A_114_112#_c_959_n 0.00252977f $X=1.515 $Y=1.84 $X2=0
+ $Y2=0
cc_569 N_VPWR_c_856_n N_A_114_112#_c_959_n 0.0136075f $X=1.65 $Y=2.825 $X2=0
+ $Y2=0
cc_570 N_VPWR_c_853_n N_A_114_112#_c_959_n 0.00116919f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_571 N_VPWR_c_861_n GCLK 0.0866997f $X=7.825 $Y=1.985 $X2=0 $Y2=0
cc_572 N_VPWR_c_859_n GCLK 0.0326636f $X=6.875 $Y=2.305 $X2=0 $Y2=0
cc_573 N_VPWR_c_867_n GCLK 0.0155928f $X=7.74 $Y=3.33 $X2=0 $Y2=0
cc_574 N_VPWR_c_853_n GCLK 0.0127818f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_575 N_A_114_112#_c_949_n N_VGND_M1009_d 0.00932283f $X=2.125 $Y=0.625 $X2=0
+ $Y2=0
cc_576 N_A_114_112#_c_948_n N_VGND_c_1085_n 0.00658627f $X=0.717 $Y=0.948 $X2=0
+ $Y2=0
cc_577 N_A_114_112#_c_950_n N_VGND_c_1085_n 0.00756924f $X=0.89 $Y=0.625 $X2=0
+ $Y2=0
cc_578 N_A_114_112#_c_949_n N_VGND_c_1091_n 0.0151441f $X=2.125 $Y=0.625 $X2=0
+ $Y2=0
cc_579 N_A_114_112#_c_953_n N_VGND_c_1091_n 0.0105752f $X=2.29 $Y=0.53 $X2=0
+ $Y2=0
cc_580 N_A_114_112#_c_949_n N_VGND_c_1095_n 0.00350553f $X=2.125 $Y=0.625 $X2=0
+ $Y2=0
cc_581 N_A_114_112#_c_950_n N_VGND_c_1095_n 0.00842441f $X=0.89 $Y=0.625 $X2=0
+ $Y2=0
cc_582 N_A_114_112#_c_949_n N_VGND_c_1098_n 0.0242087f $X=2.125 $Y=0.625 $X2=0
+ $Y2=0
cc_583 N_A_114_112#_c_949_n N_VGND_c_1100_n 0.0288276f $X=2.125 $Y=0.625 $X2=0
+ $Y2=0
cc_584 N_A_114_112#_c_950_n N_VGND_c_1100_n 0.0111078f $X=0.89 $Y=0.625 $X2=0
+ $Y2=0
cc_585 N_A_114_112#_c_953_n N_VGND_c_1100_n 0.00897192f $X=2.29 $Y=0.53 $X2=0
+ $Y2=0
cc_586 N_GCLK_c_1047_n N_VGND_c_1088_n 0.0164982f $X=7.46 $Y=0.515 $X2=0 $Y2=0
cc_587 N_GCLK_c_1047_n N_VGND_c_1090_n 0.0293763f $X=7.46 $Y=0.515 $X2=0 $Y2=0
cc_588 N_GCLK_c_1047_n N_VGND_c_1097_n 0.0144922f $X=7.46 $Y=0.515 $X2=0 $Y2=0
cc_589 N_GCLK_c_1047_n N_VGND_c_1100_n 0.0118826f $X=7.46 $Y=0.515 $X2=0 $Y2=0
