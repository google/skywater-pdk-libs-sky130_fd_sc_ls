* File: sky130_fd_sc_ls__a221oi_4.spice
* Created: Fri Aug 28 12:53:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__a221oi_4.pex.spice"
.subckt sky130_fd_sc_ls__a221oi_4  VNB VPB C1 A2 A1 B1 B2 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* B2	B2
* B1	B1
* A1	A1
* A2	A2
* C1	C1
* VPB	VPB
* VNB	VNB
MM1014 N_VGND_M1014_d N_C1_M1014_g N_Y_M1014_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1961 PD=1.02 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.5 A=0.111 P=1.78 MULT=1
MM1024 N_VGND_M1014_d N_C1_M1024_g N_Y_M1024_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1028 N_VGND_M1028_d N_C1_M1028_g N_Y_M1024_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1039 N_VGND_M1028_d N_C1_M1039_g N_Y_M1039_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1961 PD=1.02 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1002 N_VGND_M1002_d N_A2_M1002_g N_A_534_74#_M1002_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1961 PD=1.02 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75003.2 A=0.111 P=1.78 MULT=1
MM1006 N_VGND_M1002_d N_A2_M1006_g N_A_534_74#_M1006_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75002.8 A=0.111 P=1.78 MULT=1
MM1019 N_VGND_M1019_d N_A2_M1019_g N_A_534_74#_M1006_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75002.3 A=0.111 P=1.78 MULT=1
MM1021 N_VGND_M1019_d N_A2_M1021_g N_A_534_74#_M1021_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75001.9 A=0.111 P=1.78 MULT=1
MM1009 N_A_534_74#_M1021_s N_A1_M1009_g N_Y_M1009_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.9
+ SB=75001.5 A=0.111 P=1.78 MULT=1
MM1026 N_A_534_74#_M1026_d N_A1_M1026_g N_Y_M1009_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.3
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1033 N_A_534_74#_M1026_d N_A1_M1033_g N_Y_M1033_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.8
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1034 N_A_534_74#_M1034_d N_A1_M1034_g N_Y_M1033_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1961 AS=0.1036 PD=2.01 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75003.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1008 N_A_1326_74#_M1008_d N_B1_M1008_g N_Y_M1008_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1961 AS=0.1036 PD=2.01 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75003.2 A=0.111 P=1.78 MULT=1
MM1010 N_A_1326_74#_M1010_d N_B1_M1010_g N_Y_M1008_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75002.8 A=0.111 P=1.78 MULT=1
MM1029 N_A_1326_74#_M1010_d N_B1_M1029_g N_Y_M1029_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75002.3 A=0.111 P=1.78 MULT=1
MM1037 N_A_1326_74#_M1037_d N_B1_M1037_g N_Y_M1029_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75001.9 A=0.111 P=1.78 MULT=1
MM1004 N_A_1326_74#_M1037_d N_B2_M1004_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.9
+ SB=75001.5 A=0.111 P=1.78 MULT=1
MM1007 N_A_1326_74#_M1007_d N_B2_M1007_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.3
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1022 N_A_1326_74#_M1007_d N_B2_M1022_g N_VGND_M1022_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.8
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1025 N_A_1326_74#_M1025_d N_B2_M1025_g N_VGND_M1022_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1961 AS=0.1036 PD=2.01 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75003.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1000 N_A_114_368#_M1000_d N_C1_M1000_g N_Y_M1000_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.308 PD=1.42 PS=2.79 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75001.5 A=0.168 P=2.54 MULT=1
MM1011 N_A_114_368#_M1000_d N_C1_M1011_g N_Y_M1011_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.6 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1035 N_A_114_368#_M1035_d N_C1_M1035_g N_Y_M1011_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75000.6 A=0.168 P=2.54 MULT=1
MM1036 N_A_114_368#_M1035_d N_C1_M1036_g N_Y_M1036_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.308 PD=1.42 PS=2.79 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.5 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1003 N_A_531_368#_M1003_d N_A2_M1003_g N_VPWR_M1003_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.308 AS=0.168 PD=2.79 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75007.2 A=0.168 P=2.54 MULT=1
MM1017 N_A_531_368#_M1017_d N_A2_M1017_g N_VPWR_M1003_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.6 SB=75006.7 A=0.168 P=2.54 MULT=1
MM1031 N_A_531_368#_M1017_d N_A2_M1031_g N_VPWR_M1031_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75006.3 A=0.168 P=2.54 MULT=1
MM1038 N_A_531_368#_M1038_d N_A2_M1038_g N_VPWR_M1031_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.5 SB=75005.8 A=0.168 P=2.54 MULT=1
MM1005 N_A_531_368#_M1038_d N_A1_M1005_g N_VPWR_M1005_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002 SB=75005.4 A=0.168 P=2.54 MULT=1
MM1015 N_A_531_368#_M1015_d N_A1_M1015_g N_VPWR_M1005_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.4 SB=75004.9 A=0.168 P=2.54 MULT=1
MM1018 N_A_531_368#_M1015_d N_A1_M1018_g N_VPWR_M1018_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.2968 PD=1.42 PS=1.65 NRD=1.7533 NRS=21.9852 M=1 R=7.46667
+ SA=75002.9 SB=75004.5 A=0.168 P=2.54 MULT=1
MM1030 N_A_531_368#_M1030_d N_A1_M1030_g N_VPWR_M1018_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.2968 PD=1.42 PS=1.65 NRD=1.7533 NRS=21.9852 M=1 R=7.46667
+ SA=75003.6 SB=75003.8 A=0.168 P=2.54 MULT=1
MM1001 N_A_531_368#_M1030_d N_B1_M1001_g N_A_114_368#_M1001_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75004 SB=75003.3 A=0.168 P=2.54 MULT=1
MM1016 N_A_531_368#_M1016_d N_B1_M1016_g N_A_114_368#_M1001_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75004.5 SB=75002.9 A=0.168 P=2.54 MULT=1
MM1027 N_A_531_368#_M1016_d N_B1_M1027_g N_A_114_368#_M1027_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75004.9 SB=75002.4 A=0.168 P=2.54 MULT=1
MM1032 N_A_531_368#_M1032_d N_B1_M1032_g N_A_114_368#_M1027_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75005.4 SB=75002 A=0.168 P=2.54 MULT=1
MM1012 N_A_114_368#_M1012_d N_B2_M1012_g N_A_531_368#_M1032_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75005.8 SB=75001.5 A=0.168 P=2.54 MULT=1
MM1013 N_A_114_368#_M1012_d N_B2_M1013_g N_A_531_368#_M1013_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75006.3 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1020 N_A_114_368#_M1020_d N_B2_M1020_g N_A_531_368#_M1013_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75006.7 SB=75000.6 A=0.168 P=2.54 MULT=1
MM1023 N_A_114_368#_M1020_d N_B2_M1023_g N_A_531_368#_M1023_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.308 PD=1.42 PS=2.79 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75007.2 SB=75000.2 A=0.168 P=2.54 MULT=1
DX40_noxref VNB VPB NWDIODE A=20.3484 P=25.6
*
.include "sky130_fd_sc_ls__a221oi_4.pxi.spice"
*
.ends
*
*
