* File: sky130_fd_sc_ls__o211ai_4.pxi.spice
* Created: Wed Sep  2 11:17:46 2020
* 
x_PM_SKY130_FD_SC_LS__O211AI_4%A1 N_A1_M1010_g N_A1_c_133_n N_A1_M1007_g
+ N_A1_c_134_n N_A1_M1009_g N_A1_M1017_g N_A1_c_135_n N_A1_M1013_g N_A1_M1022_g
+ N_A1_c_136_n N_A1_M1023_g N_A1_M1024_g A1 A1 A1 A1 N_A1_c_132_n
+ PM_SKY130_FD_SC_LS__O211AI_4%A1
x_PM_SKY130_FD_SC_LS__O211AI_4%A2 N_A2_M1002_g N_A2_c_220_n N_A2_M1004_g
+ N_A2_M1005_g N_A2_c_221_n N_A2_M1011_g N_A2_M1008_g N_A2_c_222_n N_A2_M1016_g
+ N_A2_M1014_g N_A2_c_223_n N_A2_M1025_g A2 A2 A2 A2 A2 N_A2_c_219_n
+ PM_SKY130_FD_SC_LS__O211AI_4%A2
x_PM_SKY130_FD_SC_LS__O211AI_4%B1 N_B1_c_305_n N_B1_M1006_g N_B1_c_306_n
+ N_B1_c_307_n N_B1_c_308_n N_B1_M1012_g N_B1_c_313_n N_B1_M1001_g N_B1_M1019_g
+ N_B1_c_314_n N_B1_M1021_g N_B1_M1020_g B1 B1 B1 N_B1_c_312_n
+ PM_SKY130_FD_SC_LS__O211AI_4%B1
x_PM_SKY130_FD_SC_LS__O211AI_4%C1 N_C1_c_386_n N_C1_M1003_g N_C1_c_387_n
+ N_C1_M1026_g N_C1_M1000_g N_C1_M1015_g N_C1_c_379_n N_C1_c_380_n N_C1_M1018_g
+ N_C1_c_382_n N_C1_M1027_g N_C1_c_384_n C1 C1 C1
+ PM_SKY130_FD_SC_LS__O211AI_4%C1
x_PM_SKY130_FD_SC_LS__O211AI_4%A_30_368# N_A_30_368#_M1007_d N_A_30_368#_M1009_d
+ N_A_30_368#_M1023_d N_A_30_368#_M1011_d N_A_30_368#_M1025_d
+ N_A_30_368#_c_450_n N_A_30_368#_c_451_n N_A_30_368#_c_462_n
+ N_A_30_368#_c_452_n N_A_30_368#_c_470_n N_A_30_368#_c_474_n
+ N_A_30_368#_c_475_n N_A_30_368#_c_453_n N_A_30_368#_c_454_n
+ N_A_30_368#_c_485_n N_A_30_368#_c_455_n N_A_30_368#_c_456_n
+ N_A_30_368#_c_478_n N_A_30_368#_c_457_n PM_SKY130_FD_SC_LS__O211AI_4%A_30_368#
x_PM_SKY130_FD_SC_LS__O211AI_4%VPWR N_VPWR_M1007_s N_VPWR_M1013_s N_VPWR_M1001_d
+ N_VPWR_M1021_d N_VPWR_M1026_d N_VPWR_c_525_n N_VPWR_c_526_n N_VPWR_c_527_n
+ N_VPWR_c_528_n N_VPWR_c_529_n N_VPWR_c_530_n N_VPWR_c_531_n VPWR
+ N_VPWR_c_532_n N_VPWR_c_533_n N_VPWR_c_534_n N_VPWR_c_524_n N_VPWR_c_536_n
+ N_VPWR_c_537_n N_VPWR_c_538_n N_VPWR_c_539_n N_VPWR_c_540_n
+ PM_SKY130_FD_SC_LS__O211AI_4%VPWR
x_PM_SKY130_FD_SC_LS__O211AI_4%Y N_Y_M1000_d N_Y_M1018_d N_Y_M1004_s N_Y_M1016_s
+ N_Y_M1001_s N_Y_M1003_s N_Y_c_626_n N_Y_c_620_n N_Y_c_621_n N_Y_c_645_n
+ N_Y_c_622_n N_Y_c_623_n N_Y_c_705_p N_Y_c_616_n N_Y_c_617_n N_Y_c_710_p
+ N_Y_c_632_n N_Y_c_637_n N_Y_c_648_n N_Y_c_665_n N_Y_c_669_n Y Y Y Y
+ N_Y_c_619_n PM_SKY130_FD_SC_LS__O211AI_4%Y
x_PM_SKY130_FD_SC_LS__O211AI_4%A_27_74# N_A_27_74#_M1010_d N_A_27_74#_M1017_d
+ N_A_27_74#_M1024_d N_A_27_74#_M1005_s N_A_27_74#_M1014_s N_A_27_74#_M1012_s
+ N_A_27_74#_M1020_s N_A_27_74#_c_713_n N_A_27_74#_c_714_n N_A_27_74#_c_715_n
+ N_A_27_74#_c_716_n N_A_27_74#_c_717_n N_A_27_74#_c_718_n N_A_27_74#_c_719_n
+ N_A_27_74#_c_720_n N_A_27_74#_c_721_n N_A_27_74#_c_722_n N_A_27_74#_c_723_n
+ N_A_27_74#_c_724_n N_A_27_74#_c_725_n N_A_27_74#_c_726_n N_A_27_74#_c_727_n
+ N_A_27_74#_c_728_n N_A_27_74#_c_729_n N_A_27_74#_c_730_n
+ PM_SKY130_FD_SC_LS__O211AI_4%A_27_74#
x_PM_SKY130_FD_SC_LS__O211AI_4%VGND N_VGND_M1010_s N_VGND_M1022_s N_VGND_M1002_d
+ N_VGND_M1008_d N_VGND_c_824_n N_VGND_c_825_n N_VGND_c_826_n N_VGND_c_827_n
+ N_VGND_c_828_n N_VGND_c_829_n VGND N_VGND_c_830_n N_VGND_c_831_n
+ N_VGND_c_832_n N_VGND_c_833_n N_VGND_c_834_n N_VGND_c_835_n N_VGND_c_836_n
+ N_VGND_c_837_n PM_SKY130_FD_SC_LS__O211AI_4%VGND
x_PM_SKY130_FD_SC_LS__O211AI_4%A_834_74# N_A_834_74#_M1006_d N_A_834_74#_M1019_d
+ N_A_834_74#_M1000_s N_A_834_74#_M1015_s N_A_834_74#_M1027_s
+ N_A_834_74#_c_918_n N_A_834_74#_c_919_n N_A_834_74#_c_920_n
+ N_A_834_74#_c_939_n N_A_834_74#_c_921_n N_A_834_74#_c_922_n
+ N_A_834_74#_c_923_n N_A_834_74#_c_924_n N_A_834_74#_c_925_n
+ N_A_834_74#_c_926_n PM_SKY130_FD_SC_LS__O211AI_4%A_834_74#
cc_1 VNB N_A1_M1010_g 0.0336211f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_A1_M1017_g 0.0234895f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_3 VNB N_A1_M1022_g 0.0240453f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=0.74
cc_4 VNB N_A1_M1024_g 0.0239939f $X=-0.19 $Y=-0.245 $X2=1.925 $Y2=0.74
cc_5 VNB A1 0.0166475f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_6 VNB N_A1_c_132_n 0.0775151f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=1.557
cc_7 VNB N_A2_M1002_g 0.0229971f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_8 VNB N_A2_M1005_g 0.0224899f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=2.4
cc_9 VNB N_A2_M1008_g 0.0227896f $X=-0.19 $Y=-0.245 $X2=1.42 $Y2=2.4
cc_10 VNB N_A2_M1014_g 0.0234714f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=2.4
cc_11 VNB A2 0.012529f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A2_c_219_n 0.0718879f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.565
cc_13 VNB N_B1_c_305_n 0.0145385f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.35
cc_14 VNB N_B1_c_306_n 0.0155482f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_B1_c_307_n 0.0091019f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.765
cc_16 VNB N_B1_c_308_n 0.0138218f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=2.4
cc_17 VNB N_B1_M1019_g 0.0222131f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_B1_M1020_g 0.030436f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB B1 0.00651754f $X=-0.19 $Y=-0.245 $X2=1.925 $Y2=1.35
cc_20 VNB N_B1_c_312_n 0.0560168f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.557
cc_21 VNB N_C1_M1000_g 0.0265174f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=2.4
cc_22 VNB N_C1_M1015_g 0.0191198f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_23 VNB N_C1_c_379_n 0.0148877f $X=-0.19 $Y=-0.245 $X2=1.42 $Y2=1.765
cc_24 VNB N_C1_c_380_n 0.0681419f $X=-0.19 $Y=-0.245 $X2=1.42 $Y2=2.4
cc_25 VNB N_C1_M1018_g 0.0190737f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=0.74
cc_26 VNB N_C1_c_382_n 0.0296235f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_C1_M1027_g 0.0264634f $X=-0.19 $Y=-0.245 $X2=1.925 $Y2=1.35
cc_28 VNB N_C1_c_384_n 0.0071842f $X=-0.19 $Y=-0.245 $X2=1.925 $Y2=0.74
cc_29 VNB C1 0.00184575f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_30 VNB N_VPWR_c_524_n 0.342803f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.565
cc_31 VNB N_Y_c_616_n 0.00674473f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.557
cc_32 VNB N_Y_c_617_n 0.00138193f $X=-0.19 $Y=-0.245 $X2=1.42 $Y2=1.557
cc_33 VNB Y 0.0125004f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=1.565
cc_34 VNB N_Y_c_619_n 0.00520142f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_27_74#_c_713_n 0.0277086f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=2.4
cc_36 VNB N_A_27_74#_c_714_n 0.00317099f $X=-0.19 $Y=-0.245 $X2=1.925 $Y2=0.74
cc_37 VNB N_A_27_74#_c_715_n 0.0104987f $X=-0.19 $Y=-0.245 $X2=1.925 $Y2=0.74
cc_38 VNB N_A_27_74#_c_716_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_39 VNB N_A_27_74#_c_717_n 0.00568769f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_40 VNB N_A_27_74#_c_718_n 0.00178908f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_27_74#_c_719_n 0.00324651f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.557
cc_42 VNB N_A_27_74#_c_720_n 0.00178908f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=1.557
cc_43 VNB N_A_27_74#_c_721_n 0.00322912f $X=-0.19 $Y=-0.245 $X2=1.42 $Y2=1.557
cc_44 VNB N_A_27_74#_c_722_n 0.0017926f $X=-0.19 $Y=-0.245 $X2=1.605 $Y2=1.515
cc_45 VNB N_A_27_74#_c_723_n 0.00846513f $X=-0.19 $Y=-0.245 $X2=1.925 $Y2=1.557
cc_46 VNB N_A_27_74#_c_724_n 0.0108245f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_27_74#_c_725_n 0.00381977f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_27_74#_c_726_n 0.00178779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_27_74#_c_727_n 0.00159638f $X=-0.19 $Y=-0.245 $X2=1.605 $Y2=1.565
cc_50 VNB N_A_27_74#_c_728_n 0.00127131f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=1.565
cc_51 VNB N_A_27_74#_c_729_n 0.00143651f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_27_74#_c_730_n 0.00123317f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_824_n 0.00578139f $X=-0.19 $Y=-0.245 $X2=1.42 $Y2=1.765
cc_54 VNB N_VGND_c_825_n 0.00485164f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=0.74
cc_55 VNB N_VGND_c_826_n 0.00250542f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=2.4
cc_56 VNB N_VGND_c_827_n 0.00323505f $X=-0.19 $Y=-0.245 $X2=1.925 $Y2=0.74
cc_57 VNB N_VGND_c_828_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_58 VNB N_VGND_c_829_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_59 VNB N_VGND_c_830_n 0.0191515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_831_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.557
cc_61 VNB N_VGND_c_832_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=1.42 $Y2=1.557
cc_62 VNB N_VGND_c_833_n 0.108808f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.565
cc_63 VNB N_VGND_c_834_n 0.442219f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_835_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_836_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_837_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_834_74#_c_918_n 0.0142521f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=0.74
cc_68 VNB N_A_834_74#_c_919_n 0.00962178f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=2.4
cc_69 VNB N_A_834_74#_c_920_n 0.00375941f $X=-0.19 $Y=-0.245 $X2=1.925 $Y2=0.74
cc_70 VNB N_A_834_74#_c_921_n 0.0138519f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_71 VNB N_A_834_74#_c_922_n 0.0328968f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_834_74#_c_923_n 0.0044358f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.515
cc_73 VNB N_A_834_74#_c_924_n 0.00123647f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.515
cc_74 VNB N_A_834_74#_c_925_n 0.00316884f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=1.557
cc_75 VNB N_A_834_74#_c_926_n 0.0023816f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.557
cc_76 VPB N_A1_c_133_n 0.0208611f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.765
cc_77 VPB N_A1_c_134_n 0.0155127f $X=-0.19 $Y=1.66 $X2=0.97 $Y2=1.765
cc_78 VPB N_A1_c_135_n 0.0155127f $X=-0.19 $Y=1.66 $X2=1.42 $Y2=1.765
cc_79 VPB N_A1_c_136_n 0.0156829f $X=-0.19 $Y=1.66 $X2=1.87 $Y2=1.765
cc_80 VPB A1 0.0168757f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.58
cc_81 VPB N_A1_c_132_n 0.0494113f $X=-0.19 $Y=1.66 $X2=1.87 $Y2=1.557
cc_82 VPB N_A2_c_220_n 0.0151599f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.765
cc_83 VPB N_A2_c_221_n 0.014664f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=0.74
cc_84 VPB N_A2_c_222_n 0.0150436f $X=-0.19 $Y=1.66 $X2=1.425 $Y2=0.74
cc_85 VPB N_A2_c_223_n 0.0188637f $X=-0.19 $Y=1.66 $X2=1.925 $Y2=0.74
cc_86 VPB A2 0.0181712f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_A2_c_219_n 0.0495874f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.565
cc_88 VPB N_B1_c_313_n 0.0195047f $X=-0.19 $Y=1.66 $X2=0.97 $Y2=2.4
cc_89 VPB N_B1_c_314_n 0.0161716f $X=-0.19 $Y=1.66 $X2=1.42 $Y2=2.4
cc_90 VPB B1 0.0101401f $X=-0.19 $Y=1.66 $X2=1.925 $Y2=1.35
cc_91 VPB N_B1_c_312_n 0.03291f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.557
cc_92 VPB N_C1_c_386_n 0.0162998f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.35
cc_93 VPB N_C1_c_387_n 0.0179643f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB N_C1_c_380_n 0.0354584f $X=-0.19 $Y=1.66 $X2=1.42 $Y2=2.4
cc_95 VPB C1 0.0104769f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_96 VPB N_A_30_368#_c_450_n 0.00723723f $X=-0.19 $Y=1.66 $X2=1.42 $Y2=2.4
cc_97 VPB N_A_30_368#_c_451_n 0.035396f $X=-0.19 $Y=1.66 $X2=1.425 $Y2=1.35
cc_98 VPB N_A_30_368#_c_452_n 0.00257348f $X=-0.19 $Y=1.66 $X2=1.87 $Y2=2.4
cc_99 VPB N_A_30_368#_c_453_n 0.0028338f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.58
cc_100 VPB N_A_30_368#_c_454_n 0.0022931f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB N_A_30_368#_c_455_n 0.00737055f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.557
cc_102 VPB N_A_30_368#_c_456_n 0.00563431f $X=-0.19 $Y=1.66 $X2=0.97 $Y2=1.557
cc_103 VPB N_A_30_368#_c_457_n 0.00171072f $X=-0.19 $Y=1.66 $X2=1.925 $Y2=1.557
cc_104 VPB N_VPWR_c_525_n 0.00799266f $X=-0.19 $Y=1.66 $X2=1.425 $Y2=0.74
cc_105 VPB N_VPWR_c_526_n 0.00769929f $X=-0.19 $Y=1.66 $X2=1.87 $Y2=2.4
cc_106 VPB N_VPWR_c_527_n 0.0121832f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB N_VPWR_c_528_n 0.0183788f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_108 VPB N_VPWR_c_529_n 0.00537359f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_109 VPB N_VPWR_c_530_n 0.0186948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_110 VPB N_VPWR_c_531_n 0.0285549f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.515
cc_111 VPB N_VPWR_c_532_n 0.0206041f $X=-0.19 $Y=1.66 $X2=1.42 $Y2=1.557
cc_112 VPB N_VPWR_c_533_n 0.0640488f $X=-0.19 $Y=1.66 $X2=1.87 $Y2=1.557
cc_113 VPB N_VPWR_c_534_n 0.0266338f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_VPWR_c_524_n 0.109013f $X=-0.19 $Y=1.66 $X2=1.2 $Y2=1.565
cc_115 VPB N_VPWR_c_536_n 0.0238275f $X=-0.19 $Y=1.66 $X2=1.68 $Y2=1.565
cc_116 VPB N_VPWR_c_537_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_538_n 0.00608948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_539_n 0.00615051f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_540_n 0.0163237f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_Y_c_620_n 0.0136413f $X=-0.19 $Y=1.66 $X2=1.925 $Y2=1.35
cc_121 VPB N_Y_c_621_n 0.00326487f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_122 VPB N_Y_c_622_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_Y_c_623_n 0.00501938f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.557
cc_124 VPB Y 0.0458711f $X=-0.19 $Y=1.66 $X2=1.68 $Y2=1.565
cc_125 VPB Y 0.061961f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 N_A1_M1024_g N_A2_M1002_g 0.0169515f $X=1.925 $Y=0.74 $X2=0 $Y2=0
cc_127 N_A1_c_136_n N_A2_c_220_n 0.0241875f $X=1.87 $Y=1.765 $X2=0 $Y2=0
cc_128 A1 A2 0.0284975f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_129 N_A1_c_132_n A2 0.00468941f $X=1.87 $Y=1.557 $X2=0 $Y2=0
cc_130 A1 N_A2_c_219_n 2.85015e-19 $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_131 N_A1_c_132_n N_A2_c_219_n 0.0198415f $X=1.87 $Y=1.557 $X2=0 $Y2=0
cc_132 N_A1_c_133_n N_A_30_368#_c_450_n 4.27055e-19 $X=0.52 $Y=1.765 $X2=0 $Y2=0
cc_133 A1 N_A_30_368#_c_450_n 0.026501f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_134 N_A1_c_133_n N_A_30_368#_c_451_n 0.0104891f $X=0.52 $Y=1.765 $X2=0 $Y2=0
cc_135 N_A1_c_134_n N_A_30_368#_c_451_n 6.45594e-19 $X=0.97 $Y=1.765 $X2=0 $Y2=0
cc_136 N_A1_c_133_n N_A_30_368#_c_462_n 0.0120074f $X=0.52 $Y=1.765 $X2=0 $Y2=0
cc_137 N_A1_c_134_n N_A_30_368#_c_462_n 0.0120074f $X=0.97 $Y=1.765 $X2=0 $Y2=0
cc_138 A1 N_A_30_368#_c_462_n 0.0393875f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_139 N_A1_c_132_n N_A_30_368#_c_462_n 0.00131353f $X=1.87 $Y=1.557 $X2=0 $Y2=0
cc_140 N_A1_c_133_n N_A_30_368#_c_452_n 6.45594e-19 $X=0.52 $Y=1.765 $X2=0 $Y2=0
cc_141 N_A1_c_134_n N_A_30_368#_c_452_n 0.0103431f $X=0.97 $Y=1.765 $X2=0 $Y2=0
cc_142 N_A1_c_135_n N_A_30_368#_c_452_n 0.0103431f $X=1.42 $Y=1.765 $X2=0 $Y2=0
cc_143 N_A1_c_136_n N_A_30_368#_c_452_n 6.45594e-19 $X=1.87 $Y=1.765 $X2=0 $Y2=0
cc_144 N_A1_c_135_n N_A_30_368#_c_470_n 0.0120074f $X=1.42 $Y=1.765 $X2=0 $Y2=0
cc_145 N_A1_c_136_n N_A_30_368#_c_470_n 0.0160999f $X=1.87 $Y=1.765 $X2=0 $Y2=0
cc_146 A1 N_A_30_368#_c_470_n 0.0295713f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_147 N_A1_c_132_n N_A_30_368#_c_470_n 0.00131353f $X=1.87 $Y=1.557 $X2=0 $Y2=0
cc_148 N_A1_c_136_n N_A_30_368#_c_474_n 9.50925e-19 $X=1.87 $Y=1.765 $X2=0 $Y2=0
cc_149 N_A1_c_135_n N_A_30_368#_c_475_n 6.22492e-19 $X=1.42 $Y=1.765 $X2=0 $Y2=0
cc_150 N_A1_c_136_n N_A_30_368#_c_475_n 0.00919154f $X=1.87 $Y=1.765 $X2=0 $Y2=0
cc_151 N_A1_c_136_n N_A_30_368#_c_454_n 0.00340501f $X=1.87 $Y=1.765 $X2=0 $Y2=0
cc_152 N_A1_c_134_n N_A_30_368#_c_478_n 4.27055e-19 $X=0.97 $Y=1.765 $X2=0 $Y2=0
cc_153 N_A1_c_135_n N_A_30_368#_c_478_n 4.27055e-19 $X=1.42 $Y=1.765 $X2=0 $Y2=0
cc_154 A1 N_A_30_368#_c_478_n 0.0237598f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_155 N_A1_c_132_n N_A_30_368#_c_478_n 0.00144162f $X=1.87 $Y=1.557 $X2=0 $Y2=0
cc_156 N_A1_c_133_n N_VPWR_c_525_n 0.00486623f $X=0.52 $Y=1.765 $X2=0 $Y2=0
cc_157 N_A1_c_134_n N_VPWR_c_525_n 0.00486623f $X=0.97 $Y=1.765 $X2=0 $Y2=0
cc_158 N_A1_c_135_n N_VPWR_c_526_n 0.00486623f $X=1.42 $Y=1.765 $X2=0 $Y2=0
cc_159 N_A1_c_136_n N_VPWR_c_526_n 0.00331651f $X=1.87 $Y=1.765 $X2=0 $Y2=0
cc_160 N_A1_c_134_n N_VPWR_c_532_n 0.00445602f $X=0.97 $Y=1.765 $X2=0 $Y2=0
cc_161 N_A1_c_135_n N_VPWR_c_532_n 0.00445602f $X=1.42 $Y=1.765 $X2=0 $Y2=0
cc_162 N_A1_c_136_n N_VPWR_c_533_n 0.0044313f $X=1.87 $Y=1.765 $X2=0 $Y2=0
cc_163 N_A1_c_133_n N_VPWR_c_524_n 0.00861133f $X=0.52 $Y=1.765 $X2=0 $Y2=0
cc_164 N_A1_c_134_n N_VPWR_c_524_n 0.00857589f $X=0.97 $Y=1.765 $X2=0 $Y2=0
cc_165 N_A1_c_135_n N_VPWR_c_524_n 0.00857589f $X=1.42 $Y=1.765 $X2=0 $Y2=0
cc_166 N_A1_c_136_n N_VPWR_c_524_n 0.00853875f $X=1.87 $Y=1.765 $X2=0 $Y2=0
cc_167 N_A1_c_133_n N_VPWR_c_536_n 0.00445602f $X=0.52 $Y=1.765 $X2=0 $Y2=0
cc_168 N_A1_M1010_g N_A_27_74#_c_713_n 0.0101077f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_169 N_A1_M1017_g N_A_27_74#_c_713_n 9.62944e-19 $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_170 N_A1_M1010_g N_A_27_74#_c_714_n 0.0115433f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_171 N_A1_M1017_g N_A_27_74#_c_714_n 0.0134851f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_172 A1 N_A_27_74#_c_714_n 0.0510636f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_173 N_A1_c_132_n N_A_27_74#_c_714_n 0.00381149f $X=1.87 $Y=1.557 $X2=0 $Y2=0
cc_174 N_A1_M1010_g N_A_27_74#_c_715_n 0.00214722f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_175 A1 N_A_27_74#_c_715_n 0.0286342f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_176 N_A1_M1017_g N_A_27_74#_c_716_n 3.97481e-19 $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_177 N_A1_M1022_g N_A_27_74#_c_716_n 0.00913563f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_178 N_A1_M1024_g N_A_27_74#_c_716_n 9.66583e-19 $X=1.925 $Y=0.74 $X2=0 $Y2=0
cc_179 N_A1_M1022_g N_A_27_74#_c_717_n 0.0115433f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_180 N_A1_M1024_g N_A_27_74#_c_717_n 0.0179212f $X=1.925 $Y=0.74 $X2=0 $Y2=0
cc_181 A1 N_A_27_74#_c_717_n 0.0317172f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_182 N_A1_c_132_n N_A_27_74#_c_717_n 0.00381149f $X=1.87 $Y=1.557 $X2=0 $Y2=0
cc_183 N_A1_M1024_g N_A_27_74#_c_718_n 3.92313e-19 $X=1.925 $Y=0.74 $X2=0 $Y2=0
cc_184 N_A1_M1022_g N_A_27_74#_c_726_n 0.00157732f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_185 A1 N_A_27_74#_c_726_n 0.0213626f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_186 N_A1_c_132_n N_A_27_74#_c_726_n 0.00232957f $X=1.87 $Y=1.557 $X2=0 $Y2=0
cc_187 N_A1_M1010_g N_VGND_c_824_n 0.00571035f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_188 N_A1_M1017_g N_VGND_c_824_n 0.0104623f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_189 N_A1_M1022_g N_VGND_c_824_n 5.17822e-19 $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_190 N_A1_M1022_g N_VGND_c_825_n 0.00423899f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_191 N_A1_M1024_g N_VGND_c_825_n 0.0103415f $X=1.925 $Y=0.74 $X2=0 $Y2=0
cc_192 N_A1_M1024_g N_VGND_c_826_n 4.71636e-19 $X=1.925 $Y=0.74 $X2=0 $Y2=0
cc_193 N_A1_M1010_g N_VGND_c_830_n 0.00434272f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_194 N_A1_M1017_g N_VGND_c_831_n 0.00383152f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_195 N_A1_M1022_g N_VGND_c_831_n 0.00434272f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_196 N_A1_M1024_g N_VGND_c_832_n 0.00383152f $X=1.925 $Y=0.74 $X2=0 $Y2=0
cc_197 N_A1_M1010_g N_VGND_c_834_n 0.00824376f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_198 N_A1_M1017_g N_VGND_c_834_n 0.0075754f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_199 N_A1_M1022_g N_VGND_c_834_n 0.00820718f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_200 N_A1_M1024_g N_VGND_c_834_n 0.00757637f $X=1.925 $Y=0.74 $X2=0 $Y2=0
cc_201 N_A2_M1014_g N_B1_c_305_n 0.0192395f $X=3.665 $Y=0.74 $X2=-0.19
+ $Y2=-0.245
cc_202 A2 N_B1_c_307_n 0.00563789f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_203 A2 B1 0.0305598f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_204 N_A2_c_219_n B1 0.00111184f $X=3.665 $Y=1.557 $X2=0 $Y2=0
cc_205 N_A2_M1014_g N_B1_c_312_n 3.10152e-19 $X=3.665 $Y=0.74 $X2=0 $Y2=0
cc_206 A2 N_B1_c_312_n 0.00204508f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_207 N_A2_c_219_n N_B1_c_312_n 0.00371778f $X=3.665 $Y=1.557 $X2=0 $Y2=0
cc_208 A2 N_A_30_368#_c_474_n 0.0180181f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_209 N_A2_c_220_n N_A_30_368#_c_453_n 0.0137488f $X=2.37 $Y=1.765 $X2=0 $Y2=0
cc_210 N_A2_c_221_n N_A_30_368#_c_453_n 0.0128349f $X=2.82 $Y=1.765 $X2=0 $Y2=0
cc_211 N_A2_c_222_n N_A_30_368#_c_485_n 0.00769091f $X=3.27 $Y=1.765 $X2=0 $Y2=0
cc_212 N_A2_c_223_n N_A_30_368#_c_485_n 5.87446e-19 $X=3.77 $Y=1.765 $X2=0 $Y2=0
cc_213 N_A2_c_222_n N_A_30_368#_c_455_n 0.0111147f $X=3.27 $Y=1.765 $X2=0 $Y2=0
cc_214 N_A2_c_223_n N_A_30_368#_c_455_n 0.0152643f $X=3.77 $Y=1.765 $X2=0 $Y2=0
cc_215 N_A2_c_222_n N_A_30_368#_c_457_n 0.00175197f $X=3.27 $Y=1.765 $X2=0 $Y2=0
cc_216 N_A2_c_223_n N_VPWR_c_527_n 0.00189254f $X=3.77 $Y=1.765 $X2=0 $Y2=0
cc_217 N_A2_c_220_n N_VPWR_c_533_n 0.00278271f $X=2.37 $Y=1.765 $X2=0 $Y2=0
cc_218 N_A2_c_221_n N_VPWR_c_533_n 0.00278271f $X=2.82 $Y=1.765 $X2=0 $Y2=0
cc_219 N_A2_c_222_n N_VPWR_c_533_n 0.00278257f $X=3.27 $Y=1.765 $X2=0 $Y2=0
cc_220 N_A2_c_223_n N_VPWR_c_533_n 0.00278271f $X=3.77 $Y=1.765 $X2=0 $Y2=0
cc_221 N_A2_c_220_n N_VPWR_c_524_n 0.00354337f $X=2.37 $Y=1.765 $X2=0 $Y2=0
cc_222 N_A2_c_221_n N_VPWR_c_524_n 0.00353823f $X=2.82 $Y=1.765 $X2=0 $Y2=0
cc_223 N_A2_c_222_n N_VPWR_c_524_n 0.00354283f $X=3.27 $Y=1.765 $X2=0 $Y2=0
cc_224 N_A2_c_223_n N_VPWR_c_524_n 0.00359085f $X=3.77 $Y=1.765 $X2=0 $Y2=0
cc_225 N_A2_c_221_n N_Y_c_626_n 0.0120074f $X=2.82 $Y=1.765 $X2=0 $Y2=0
cc_226 N_A2_c_222_n N_Y_c_626_n 0.0151589f $X=3.27 $Y=1.765 $X2=0 $Y2=0
cc_227 A2 N_Y_c_626_n 0.0420324f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_228 N_A2_c_219_n N_Y_c_626_n 0.00146022f $X=3.665 $Y=1.557 $X2=0 $Y2=0
cc_229 N_A2_c_223_n N_Y_c_620_n 0.0139279f $X=3.77 $Y=1.765 $X2=0 $Y2=0
cc_230 A2 N_Y_c_620_n 0.0356307f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_231 N_A2_c_220_n N_Y_c_632_n 0.00869368f $X=2.37 $Y=1.765 $X2=0 $Y2=0
cc_232 N_A2_c_221_n N_Y_c_632_n 0.00904709f $X=2.82 $Y=1.765 $X2=0 $Y2=0
cc_233 N_A2_c_222_n N_Y_c_632_n 4.45174e-19 $X=3.27 $Y=1.765 $X2=0 $Y2=0
cc_234 A2 N_Y_c_632_n 0.0237597f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_235 N_A2_c_219_n N_Y_c_632_n 0.0016057f $X=3.665 $Y=1.557 $X2=0 $Y2=0
cc_236 N_A2_c_223_n N_Y_c_637_n 0.01303f $X=3.77 $Y=1.765 $X2=0 $Y2=0
cc_237 A2 N_Y_c_637_n 0.0254779f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_238 N_A2_c_219_n N_Y_c_637_n 0.00186492f $X=3.665 $Y=1.557 $X2=0 $Y2=0
cc_239 A2 N_A_27_74#_c_717_n 7.722e-19 $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_240 N_A2_M1002_g N_A_27_74#_c_718_n 3.92313e-19 $X=2.355 $Y=0.74 $X2=0 $Y2=0
cc_241 N_A2_M1002_g N_A_27_74#_c_719_n 0.013073f $X=2.355 $Y=0.74 $X2=0 $Y2=0
cc_242 N_A2_M1005_g N_A_27_74#_c_719_n 0.0130918f $X=2.785 $Y=0.74 $X2=0 $Y2=0
cc_243 A2 N_A_27_74#_c_719_n 0.0519686f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_244 N_A2_c_219_n N_A_27_74#_c_719_n 0.00230191f $X=3.665 $Y=1.557 $X2=0 $Y2=0
cc_245 N_A2_M1005_g N_A_27_74#_c_720_n 3.92313e-19 $X=2.785 $Y=0.74 $X2=0 $Y2=0
cc_246 N_A2_M1008_g N_A_27_74#_c_720_n 3.92313e-19 $X=3.215 $Y=0.74 $X2=0 $Y2=0
cc_247 N_A2_M1008_g N_A_27_74#_c_721_n 0.0132118f $X=3.215 $Y=0.74 $X2=0 $Y2=0
cc_248 N_A2_M1014_g N_A_27_74#_c_721_n 0.0136953f $X=3.665 $Y=0.74 $X2=0 $Y2=0
cc_249 A2 N_A_27_74#_c_721_n 0.0534599f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_250 N_A2_c_219_n N_A_27_74#_c_721_n 0.0032112f $X=3.665 $Y=1.557 $X2=0 $Y2=0
cc_251 N_A2_M1014_g N_A_27_74#_c_722_n 3.97896e-19 $X=3.665 $Y=0.74 $X2=0 $Y2=0
cc_252 A2 N_A_27_74#_c_723_n 0.0189979f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_253 A2 N_A_27_74#_c_727_n 0.0153286f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_254 A2 N_A_27_74#_c_728_n 0.0146029f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_255 N_A2_c_219_n N_A_27_74#_c_728_n 0.00238948f $X=3.665 $Y=1.557 $X2=0 $Y2=0
cc_256 A2 N_A_27_74#_c_729_n 0.0153284f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_257 N_A2_c_219_n N_A_27_74#_c_729_n 3.07687e-19 $X=3.665 $Y=1.557 $X2=0 $Y2=0
cc_258 N_A2_M1002_g N_VGND_c_825_n 4.71636e-19 $X=2.355 $Y=0.74 $X2=0 $Y2=0
cc_259 N_A2_M1002_g N_VGND_c_826_n 0.0103289f $X=2.355 $Y=0.74 $X2=0 $Y2=0
cc_260 N_A2_M1005_g N_VGND_c_826_n 0.0103289f $X=2.785 $Y=0.74 $X2=0 $Y2=0
cc_261 N_A2_M1008_g N_VGND_c_826_n 4.71636e-19 $X=3.215 $Y=0.74 $X2=0 $Y2=0
cc_262 N_A2_M1005_g N_VGND_c_827_n 4.71636e-19 $X=2.785 $Y=0.74 $X2=0 $Y2=0
cc_263 N_A2_M1008_g N_VGND_c_827_n 0.0104789f $X=3.215 $Y=0.74 $X2=0 $Y2=0
cc_264 N_A2_M1014_g N_VGND_c_827_n 0.00910824f $X=3.665 $Y=0.74 $X2=0 $Y2=0
cc_265 N_A2_M1005_g N_VGND_c_828_n 0.00383152f $X=2.785 $Y=0.74 $X2=0 $Y2=0
cc_266 N_A2_M1008_g N_VGND_c_828_n 0.00383152f $X=3.215 $Y=0.74 $X2=0 $Y2=0
cc_267 N_A2_M1002_g N_VGND_c_832_n 0.00383152f $X=2.355 $Y=0.74 $X2=0 $Y2=0
cc_268 N_A2_M1014_g N_VGND_c_833_n 0.00444681f $X=3.665 $Y=0.74 $X2=0 $Y2=0
cc_269 N_A2_M1002_g N_VGND_c_834_n 0.00757637f $X=2.355 $Y=0.74 $X2=0 $Y2=0
cc_270 N_A2_M1005_g N_VGND_c_834_n 0.0075754f $X=2.785 $Y=0.74 $X2=0 $Y2=0
cc_271 N_A2_M1008_g N_VGND_c_834_n 0.0075754f $X=3.215 $Y=0.74 $X2=0 $Y2=0
cc_272 N_A2_M1014_g N_VGND_c_834_n 0.00877616f $X=3.665 $Y=0.74 $X2=0 $Y2=0
cc_273 N_A2_M1014_g N_A_834_74#_c_923_n 3.65259e-19 $X=3.665 $Y=0.74 $X2=0 $Y2=0
cc_274 N_B1_c_314_n N_C1_c_386_n 0.028874f $X=5.37 $Y=1.765 $X2=-0.19 $Y2=-0.245
cc_275 B1 N_C1_c_380_n 0.00397058f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_276 N_B1_c_312_n N_C1_c_380_n 0.0148278f $X=5.37 $Y=1.475 $X2=0 $Y2=0
cc_277 B1 C1 0.029855f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_278 N_B1_c_312_n C1 3.61244e-19 $X=5.37 $Y=1.475 $X2=0 $Y2=0
cc_279 N_B1_c_313_n N_A_30_368#_c_455_n 5.94256e-19 $X=4.83 $Y=1.765 $X2=0 $Y2=0
cc_280 N_B1_c_313_n N_A_30_368#_c_456_n 0.00115567f $X=4.83 $Y=1.765 $X2=0 $Y2=0
cc_281 N_B1_c_313_n N_VPWR_c_527_n 0.0128703f $X=4.83 $Y=1.765 $X2=0 $Y2=0
cc_282 N_B1_c_314_n N_VPWR_c_527_n 4.83094e-19 $X=5.37 $Y=1.765 $X2=0 $Y2=0
cc_283 N_B1_c_313_n N_VPWR_c_528_n 0.00413917f $X=4.83 $Y=1.765 $X2=0 $Y2=0
cc_284 N_B1_c_314_n N_VPWR_c_528_n 0.00444681f $X=5.37 $Y=1.765 $X2=0 $Y2=0
cc_285 N_B1_c_313_n N_VPWR_c_529_n 4.73566e-19 $X=4.83 $Y=1.765 $X2=0 $Y2=0
cc_286 N_B1_c_314_n N_VPWR_c_529_n 0.0104404f $X=5.37 $Y=1.765 $X2=0 $Y2=0
cc_287 N_B1_c_313_n N_VPWR_c_524_n 0.00818526f $X=4.83 $Y=1.765 $X2=0 $Y2=0
cc_288 N_B1_c_314_n N_VPWR_c_524_n 0.00878515f $X=5.37 $Y=1.765 $X2=0 $Y2=0
cc_289 N_B1_c_306_n N_Y_c_620_n 0.00626133f $X=4.45 $Y=1.26 $X2=0 $Y2=0
cc_290 N_B1_c_313_n N_Y_c_620_n 0.0172731f $X=4.83 $Y=1.765 $X2=0 $Y2=0
cc_291 B1 N_Y_c_620_n 0.0351028f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_292 N_B1_c_312_n N_Y_c_620_n 0.00148857f $X=5.37 $Y=1.475 $X2=0 $Y2=0
cc_293 N_B1_c_313_n N_Y_c_621_n 0.00507697f $X=4.83 $Y=1.765 $X2=0 $Y2=0
cc_294 N_B1_c_314_n N_Y_c_645_n 0.0131978f $X=5.37 $Y=1.765 $X2=0 $Y2=0
cc_295 B1 N_Y_c_645_n 0.0250576f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_296 N_B1_c_314_n N_Y_c_622_n 4.54343e-19 $X=5.37 $Y=1.765 $X2=0 $Y2=0
cc_297 B1 N_Y_c_648_n 0.0267474f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_298 N_B1_c_312_n N_Y_c_648_n 0.00188247f $X=5.37 $Y=1.475 $X2=0 $Y2=0
cc_299 N_B1_c_305_n N_A_27_74#_c_722_n 3.92031e-19 $X=4.095 $Y=1.185 $X2=0 $Y2=0
cc_300 N_B1_c_305_n N_A_27_74#_c_723_n 0.014886f $X=4.095 $Y=1.185 $X2=0 $Y2=0
cc_301 N_B1_c_306_n N_A_27_74#_c_723_n 0.00449289f $X=4.45 $Y=1.26 $X2=0 $Y2=0
cc_302 N_B1_c_308_n N_A_27_74#_c_723_n 0.014287f $X=4.525 $Y=1.185 $X2=0 $Y2=0
cc_303 B1 N_A_27_74#_c_723_n 0.0762823f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_304 N_B1_c_312_n N_A_27_74#_c_723_n 0.00243496f $X=5.37 $Y=1.475 $X2=0 $Y2=0
cc_305 N_B1_M1019_g N_A_27_74#_c_724_n 0.00822358f $X=4.955 $Y=0.74 $X2=0 $Y2=0
cc_306 N_B1_M1020_g N_A_27_74#_c_724_n 0.0122724f $X=5.385 $Y=0.74 $X2=0 $Y2=0
cc_307 B1 N_A_27_74#_c_724_n 0.0176085f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_308 N_B1_c_312_n N_A_27_74#_c_724_n 0.00224206f $X=5.37 $Y=1.475 $X2=0 $Y2=0
cc_309 N_B1_M1019_g N_A_27_74#_c_725_n 5.58807e-19 $X=4.955 $Y=0.74 $X2=0 $Y2=0
cc_310 N_B1_M1020_g N_A_27_74#_c_725_n 0.00723951f $X=5.385 $Y=0.74 $X2=0 $Y2=0
cc_311 N_B1_M1019_g N_A_27_74#_c_730_n 0.00507129f $X=4.955 $Y=0.74 $X2=0 $Y2=0
cc_312 N_B1_M1020_g N_A_27_74#_c_730_n 5.06799e-19 $X=5.385 $Y=0.74 $X2=0 $Y2=0
cc_313 N_B1_c_305_n N_VGND_c_827_n 5.0386e-19 $X=4.095 $Y=1.185 $X2=0 $Y2=0
cc_314 N_B1_c_305_n N_VGND_c_833_n 0.00430932f $X=4.095 $Y=1.185 $X2=0 $Y2=0
cc_315 N_B1_c_308_n N_VGND_c_833_n 0.00278271f $X=4.525 $Y=1.185 $X2=0 $Y2=0
cc_316 N_B1_M1019_g N_VGND_c_833_n 0.00278271f $X=4.955 $Y=0.74 $X2=0 $Y2=0
cc_317 N_B1_M1020_g N_VGND_c_833_n 0.00278271f $X=5.385 $Y=0.74 $X2=0 $Y2=0
cc_318 N_B1_c_305_n N_VGND_c_834_n 0.00442002f $X=4.095 $Y=1.185 $X2=0 $Y2=0
cc_319 N_B1_c_308_n N_VGND_c_834_n 0.00353428f $X=4.525 $Y=1.185 $X2=0 $Y2=0
cc_320 N_B1_M1019_g N_VGND_c_834_n 0.00353428f $X=4.955 $Y=0.74 $X2=0 $Y2=0
cc_321 N_B1_M1020_g N_VGND_c_834_n 0.00358427f $X=5.385 $Y=0.74 $X2=0 $Y2=0
cc_322 N_B1_M1020_g N_A_834_74#_c_918_n 0.0125531f $X=5.385 $Y=0.74 $X2=0 $Y2=0
cc_323 N_B1_M1020_g N_A_834_74#_c_919_n 0.00573384f $X=5.385 $Y=0.74 $X2=0 $Y2=0
cc_324 N_B1_c_305_n N_A_834_74#_c_923_n 0.00660507f $X=4.095 $Y=1.185 $X2=0
+ $Y2=0
cc_325 N_B1_c_308_n N_A_834_74#_c_923_n 0.0143701f $X=4.525 $Y=1.185 $X2=0 $Y2=0
cc_326 N_B1_M1019_g N_A_834_74#_c_923_n 0.015701f $X=4.955 $Y=0.74 $X2=0 $Y2=0
cc_327 N_C1_c_386_n N_VPWR_c_529_n 0.00558426f $X=5.88 $Y=1.765 $X2=0 $Y2=0
cc_328 N_C1_c_386_n N_VPWR_c_530_n 0.00445602f $X=5.88 $Y=1.765 $X2=0 $Y2=0
cc_329 N_C1_c_387_n N_VPWR_c_530_n 0.00445602f $X=6.33 $Y=1.765 $X2=0 $Y2=0
cc_330 N_C1_c_387_n N_VPWR_c_531_n 0.00399808f $X=6.33 $Y=1.765 $X2=0 $Y2=0
cc_331 N_C1_c_386_n N_VPWR_c_524_n 0.00857513f $X=5.88 $Y=1.765 $X2=0 $Y2=0
cc_332 N_C1_c_387_n N_VPWR_c_524_n 0.00861719f $X=6.33 $Y=1.765 $X2=0 $Y2=0
cc_333 N_C1_c_386_n N_Y_c_645_n 0.0141391f $X=5.88 $Y=1.765 $X2=0 $Y2=0
cc_334 C1 N_Y_c_645_n 0.00507353f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_335 N_C1_c_386_n N_Y_c_622_n 0.010238f $X=5.88 $Y=1.765 $X2=0 $Y2=0
cc_336 N_C1_c_387_n N_Y_c_622_n 0.0144423f $X=6.33 $Y=1.765 $X2=0 $Y2=0
cc_337 N_C1_c_387_n N_Y_c_623_n 0.0139279f $X=6.33 $Y=1.765 $X2=0 $Y2=0
cc_338 N_C1_c_379_n N_Y_c_623_n 0.00966332f $X=7.16 $Y=1.425 $X2=0 $Y2=0
cc_339 N_C1_c_380_n N_Y_c_623_n 0.00240711f $X=6.88 $Y=1.425 $X2=0 $Y2=0
cc_340 C1 N_Y_c_623_n 0.0611122f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_341 N_C1_M1015_g N_Y_c_616_n 0.0109453f $X=6.805 $Y=0.79 $X2=0 $Y2=0
cc_342 N_C1_c_379_n N_Y_c_616_n 0.00190909f $X=7.16 $Y=1.425 $X2=0 $Y2=0
cc_343 N_C1_M1018_g N_Y_c_616_n 0.0149475f $X=7.235 $Y=0.79 $X2=0 $Y2=0
cc_344 C1 N_Y_c_616_n 0.030047f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_345 N_C1_M1000_g N_Y_c_617_n 4.99029e-19 $X=6.375 $Y=0.79 $X2=0 $Y2=0
cc_346 N_C1_c_380_n N_Y_c_617_n 0.00231547f $X=6.88 $Y=1.425 $X2=0 $Y2=0
cc_347 C1 N_Y_c_617_n 0.0144276f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_348 N_C1_c_386_n N_Y_c_665_n 4.27055e-19 $X=5.88 $Y=1.765 $X2=0 $Y2=0
cc_349 N_C1_c_387_n N_Y_c_665_n 4.27055e-19 $X=6.33 $Y=1.765 $X2=0 $Y2=0
cc_350 N_C1_c_380_n N_Y_c_665_n 0.00145364f $X=6.88 $Y=1.425 $X2=0 $Y2=0
cc_351 C1 N_Y_c_665_n 0.0237598f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_352 N_C1_M1027_g N_Y_c_669_n 5.05504e-19 $X=7.665 $Y=0.79 $X2=0 $Y2=0
cc_353 N_C1_c_382_n Y 0.0102519f $X=7.59 $Y=1.425 $X2=0 $Y2=0
cc_354 N_C1_c_380_n N_Y_c_619_n 8.68505e-19 $X=6.88 $Y=1.425 $X2=0 $Y2=0
cc_355 N_C1_M1018_g N_Y_c_619_n 0.00407735f $X=7.235 $Y=0.79 $X2=0 $Y2=0
cc_356 N_C1_c_382_n N_Y_c_619_n 0.0176888f $X=7.59 $Y=1.425 $X2=0 $Y2=0
cc_357 N_C1_M1027_g N_Y_c_619_n 0.00412955f $X=7.665 $Y=0.79 $X2=0 $Y2=0
cc_358 C1 N_Y_c_619_n 0.0250193f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_359 N_C1_M1000_g N_A_27_74#_c_724_n 3.9607e-19 $X=6.375 $Y=0.79 $X2=0 $Y2=0
cc_360 N_C1_M1000_g N_A_27_74#_c_725_n 8.49936e-19 $X=6.375 $Y=0.79 $X2=0 $Y2=0
cc_361 N_C1_M1000_g N_VGND_c_833_n 8.94875e-19 $X=6.375 $Y=0.79 $X2=0 $Y2=0
cc_362 N_C1_M1015_g N_VGND_c_833_n 8.94875e-19 $X=6.805 $Y=0.79 $X2=0 $Y2=0
cc_363 N_C1_M1018_g N_VGND_c_833_n 8.94875e-19 $X=7.235 $Y=0.79 $X2=0 $Y2=0
cc_364 N_C1_M1027_g N_VGND_c_833_n 8.94875e-19 $X=7.665 $Y=0.79 $X2=0 $Y2=0
cc_365 N_C1_M1000_g N_A_834_74#_c_919_n 0.0109245f $X=6.375 $Y=0.79 $X2=0 $Y2=0
cc_366 N_C1_M1015_g N_A_834_74#_c_919_n 7.18637e-19 $X=6.805 $Y=0.79 $X2=0 $Y2=0
cc_367 N_C1_c_380_n N_A_834_74#_c_919_n 0.00727567f $X=6.88 $Y=1.425 $X2=0 $Y2=0
cc_368 C1 N_A_834_74#_c_919_n 0.0280641f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_369 N_C1_M1000_g N_A_834_74#_c_920_n 0.0104623f $X=6.375 $Y=0.79 $X2=0 $Y2=0
cc_370 N_C1_M1015_g N_A_834_74#_c_920_n 0.00831767f $X=6.805 $Y=0.79 $X2=0 $Y2=0
cc_371 N_C1_M1000_g N_A_834_74#_c_939_n 5.7278e-19 $X=6.375 $Y=0.79 $X2=0 $Y2=0
cc_372 N_C1_M1015_g N_A_834_74#_c_939_n 0.00628142f $X=6.805 $Y=0.79 $X2=0 $Y2=0
cc_373 N_C1_M1018_g N_A_834_74#_c_939_n 0.00628142f $X=7.235 $Y=0.79 $X2=0 $Y2=0
cc_374 N_C1_M1027_g N_A_834_74#_c_939_n 5.7278e-19 $X=7.665 $Y=0.79 $X2=0 $Y2=0
cc_375 N_C1_M1018_g N_A_834_74#_c_921_n 0.00831767f $X=7.235 $Y=0.79 $X2=0 $Y2=0
cc_376 N_C1_M1027_g N_A_834_74#_c_921_n 0.013752f $X=7.665 $Y=0.79 $X2=0 $Y2=0
cc_377 N_C1_M1018_g N_A_834_74#_c_922_n 7.09577e-19 $X=7.235 $Y=0.79 $X2=0 $Y2=0
cc_378 N_C1_M1027_g N_A_834_74#_c_922_n 0.0108615f $X=7.665 $Y=0.79 $X2=0 $Y2=0
cc_379 N_C1_M1000_g N_A_834_74#_c_925_n 0.00379107f $X=6.375 $Y=0.79 $X2=0 $Y2=0
cc_380 N_C1_M1015_g N_A_834_74#_c_926_n 0.00229636f $X=6.805 $Y=0.79 $X2=0 $Y2=0
cc_381 N_C1_M1018_g N_A_834_74#_c_926_n 0.00229636f $X=7.235 $Y=0.79 $X2=0 $Y2=0
cc_382 N_A_30_368#_c_462_n N_VPWR_M1007_s 0.00408911f $X=1.03 $Y=2.035 $X2=-0.19
+ $Y2=1.66
cc_383 N_A_30_368#_c_470_n N_VPWR_M1013_s 0.00408911f $X=1.93 $Y=2.035 $X2=0
+ $Y2=0
cc_384 N_A_30_368#_c_451_n N_VPWR_c_525_n 0.0449718f $X=0.295 $Y=2.815 $X2=0
+ $Y2=0
cc_385 N_A_30_368#_c_462_n N_VPWR_c_525_n 0.0136682f $X=1.03 $Y=2.035 $X2=0
+ $Y2=0
cc_386 N_A_30_368#_c_452_n N_VPWR_c_525_n 0.0449718f $X=1.195 $Y=2.815 $X2=0
+ $Y2=0
cc_387 N_A_30_368#_c_452_n N_VPWR_c_526_n 0.0449718f $X=1.195 $Y=2.815 $X2=0
+ $Y2=0
cc_388 N_A_30_368#_c_470_n N_VPWR_c_526_n 0.0136682f $X=1.93 $Y=2.035 $X2=0
+ $Y2=0
cc_389 N_A_30_368#_c_475_n N_VPWR_c_526_n 0.0400262f $X=2.095 $Y=2.815 $X2=0
+ $Y2=0
cc_390 N_A_30_368#_c_454_n N_VPWR_c_526_n 0.0119328f $X=2.26 $Y=2.99 $X2=0 $Y2=0
cc_391 N_A_30_368#_c_455_n N_VPWR_c_527_n 0.0121618f $X=3.88 $Y=2.99 $X2=0 $Y2=0
cc_392 N_A_30_368#_c_456_n N_VPWR_c_527_n 0.041429f $X=4.045 $Y=2.375 $X2=0
+ $Y2=0
cc_393 N_A_30_368#_c_452_n N_VPWR_c_532_n 0.014552f $X=1.195 $Y=2.815 $X2=0
+ $Y2=0
cc_394 N_A_30_368#_c_453_n N_VPWR_c_533_n 0.0441612f $X=2.96 $Y=2.99 $X2=0 $Y2=0
cc_395 N_A_30_368#_c_454_n N_VPWR_c_533_n 0.0236039f $X=2.26 $Y=2.99 $X2=0 $Y2=0
cc_396 N_A_30_368#_c_455_n N_VPWR_c_533_n 0.0659319f $X=3.88 $Y=2.99 $X2=0 $Y2=0
cc_397 N_A_30_368#_c_457_n N_VPWR_c_533_n 0.017869f $X=3.085 $Y=2.99 $X2=0 $Y2=0
cc_398 N_A_30_368#_c_451_n N_VPWR_c_524_n 0.0120466f $X=0.295 $Y=2.815 $X2=0
+ $Y2=0
cc_399 N_A_30_368#_c_452_n N_VPWR_c_524_n 0.0119791f $X=1.195 $Y=2.815 $X2=0
+ $Y2=0
cc_400 N_A_30_368#_c_453_n N_VPWR_c_524_n 0.0249452f $X=2.96 $Y=2.99 $X2=0 $Y2=0
cc_401 N_A_30_368#_c_454_n N_VPWR_c_524_n 0.012761f $X=2.26 $Y=2.99 $X2=0 $Y2=0
cc_402 N_A_30_368#_c_455_n N_VPWR_c_524_n 0.0367158f $X=3.88 $Y=2.99 $X2=0 $Y2=0
cc_403 N_A_30_368#_c_457_n N_VPWR_c_524_n 0.00965079f $X=3.085 $Y=2.99 $X2=0
+ $Y2=0
cc_404 N_A_30_368#_c_451_n N_VPWR_c_536_n 0.0145938f $X=0.295 $Y=2.815 $X2=0
+ $Y2=0
cc_405 N_A_30_368#_c_453_n N_Y_M1004_s 0.00197722f $X=2.96 $Y=2.99 $X2=0 $Y2=0
cc_406 N_A_30_368#_c_455_n N_Y_M1016_s 0.00250873f $X=3.88 $Y=2.99 $X2=0 $Y2=0
cc_407 N_A_30_368#_M1011_d N_Y_c_626_n 0.00381296f $X=2.895 $Y=1.84 $X2=0 $Y2=0
cc_408 N_A_30_368#_c_485_n N_Y_c_626_n 0.0154248f $X=3.045 $Y=2.455 $X2=0 $Y2=0
cc_409 N_A_30_368#_M1025_d N_Y_c_620_n 0.00751585f $X=3.845 $Y=1.84 $X2=0 $Y2=0
cc_410 N_A_30_368#_c_456_n N_Y_c_620_n 0.025036f $X=4.045 $Y=2.375 $X2=0 $Y2=0
cc_411 N_A_30_368#_c_453_n N_Y_c_632_n 0.0160777f $X=2.96 $Y=2.99 $X2=0 $Y2=0
cc_412 N_A_30_368#_c_485_n N_Y_c_632_n 0.0298377f $X=3.045 $Y=2.455 $X2=0 $Y2=0
cc_413 N_A_30_368#_c_455_n N_Y_c_637_n 0.018923f $X=3.88 $Y=2.99 $X2=0 $Y2=0
cc_414 N_VPWR_M1001_d N_Y_c_620_n 0.00566769f $X=4.46 $Y=1.84 $X2=0 $Y2=0
cc_415 N_VPWR_c_527_n N_Y_c_620_n 0.0219924f $X=4.605 $Y=2.375 $X2=0 $Y2=0
cc_416 N_VPWR_c_527_n N_Y_c_621_n 0.0266809f $X=4.605 $Y=2.375 $X2=0 $Y2=0
cc_417 N_VPWR_c_528_n N_Y_c_621_n 0.0146357f $X=5.44 $Y=3.33 $X2=0 $Y2=0
cc_418 N_VPWR_c_529_n N_Y_c_621_n 0.0266809f $X=5.605 $Y=2.375 $X2=0 $Y2=0
cc_419 N_VPWR_c_524_n N_Y_c_621_n 0.0121141f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_420 N_VPWR_M1021_d N_Y_c_645_n 0.00834387f $X=5.445 $Y=1.84 $X2=0 $Y2=0
cc_421 N_VPWR_c_529_n N_Y_c_645_n 0.0202768f $X=5.605 $Y=2.375 $X2=0 $Y2=0
cc_422 N_VPWR_c_529_n N_Y_c_622_n 0.0266809f $X=5.605 $Y=2.375 $X2=0 $Y2=0
cc_423 N_VPWR_c_530_n N_Y_c_622_n 0.014552f $X=6.44 $Y=3.33 $X2=0 $Y2=0
cc_424 N_VPWR_c_531_n N_Y_c_622_n 0.0267725f $X=7.125 $Y=2.455 $X2=0 $Y2=0
cc_425 N_VPWR_c_524_n N_Y_c_622_n 0.0119791f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_426 N_VPWR_M1026_d N_Y_c_623_n 0.023281f $X=6.405 $Y=1.84 $X2=0 $Y2=0
cc_427 N_VPWR_c_531_n N_Y_c_623_n 0.0673425f $X=7.125 $Y=2.455 $X2=0 $Y2=0
cc_428 N_VPWR_c_531_n Y 0.0410158f $X=7.125 $Y=2.455 $X2=0 $Y2=0
cc_429 N_VPWR_c_534_n Y 0.0159573f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_430 N_VPWR_c_524_n Y 0.0170149f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_431 N_Y_c_616_n N_A_834_74#_M1015_s 0.00176461f $X=7.365 $Y=1.095 $X2=0 $Y2=0
cc_432 N_Y_c_617_n N_A_834_74#_c_919_n 0.00697079f $X=6.675 $Y=1.095 $X2=0 $Y2=0
cc_433 N_Y_M1000_d N_A_834_74#_c_920_n 0.00176461f $X=6.45 $Y=0.42 $X2=0 $Y2=0
cc_434 N_Y_c_705_p N_A_834_74#_c_920_n 0.0124895f $X=6.59 $Y=0.885 $X2=0 $Y2=0
cc_435 N_Y_c_616_n N_A_834_74#_c_920_n 0.0030313f $X=7.365 $Y=1.095 $X2=0 $Y2=0
cc_436 N_Y_c_616_n N_A_834_74#_c_939_n 0.0168694f $X=7.365 $Y=1.095 $X2=0 $Y2=0
cc_437 N_Y_M1018_d N_A_834_74#_c_921_n 0.00176461f $X=7.31 $Y=0.42 $X2=0 $Y2=0
cc_438 N_Y_c_616_n N_A_834_74#_c_921_n 0.0030313f $X=7.365 $Y=1.095 $X2=0 $Y2=0
cc_439 N_Y_c_710_p N_A_834_74#_c_921_n 0.0126348f $X=7.45 $Y=0.885 $X2=0 $Y2=0
cc_440 N_Y_c_669_n N_A_834_74#_c_922_n 0.00729487f $X=7.455 $Y=1.095 $X2=0 $Y2=0
cc_441 Y N_A_834_74#_c_922_n 0.0172112f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_442 N_A_27_74#_c_714_n N_VGND_M1010_s 0.00250873f $X=1.125 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_443 N_A_27_74#_c_717_n N_VGND_M1022_s 0.00250873f $X=2.055 $Y=1.095 $X2=0
+ $Y2=0
cc_444 N_A_27_74#_c_719_n N_VGND_M1002_d 0.00176461f $X=2.915 $Y=1.095 $X2=0
+ $Y2=0
cc_445 N_A_27_74#_c_721_n N_VGND_M1008_d 0.00197722f $X=3.795 $Y=1.095 $X2=0
+ $Y2=0
cc_446 N_A_27_74#_c_713_n N_VGND_c_824_n 0.0191765f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_447 N_A_27_74#_c_714_n N_VGND_c_824_n 0.0210288f $X=1.125 $Y=1.095 $X2=0
+ $Y2=0
cc_448 N_A_27_74#_c_716_n N_VGND_c_824_n 0.0182902f $X=1.21 $Y=0.515 $X2=0 $Y2=0
cc_449 N_A_27_74#_c_716_n N_VGND_c_825_n 0.0184106f $X=1.21 $Y=0.515 $X2=0 $Y2=0
cc_450 N_A_27_74#_c_717_n N_VGND_c_825_n 0.0210288f $X=2.055 $Y=1.095 $X2=0
+ $Y2=0
cc_451 N_A_27_74#_c_718_n N_VGND_c_825_n 0.0182488f $X=2.14 $Y=0.515 $X2=0 $Y2=0
cc_452 N_A_27_74#_c_718_n N_VGND_c_826_n 0.0182488f $X=2.14 $Y=0.515 $X2=0 $Y2=0
cc_453 N_A_27_74#_c_719_n N_VGND_c_826_n 0.0171619f $X=2.915 $Y=1.095 $X2=0
+ $Y2=0
cc_454 N_A_27_74#_c_720_n N_VGND_c_826_n 0.0182488f $X=3 $Y=0.515 $X2=0 $Y2=0
cc_455 N_A_27_74#_c_720_n N_VGND_c_827_n 0.0182488f $X=3 $Y=0.515 $X2=0 $Y2=0
cc_456 N_A_27_74#_c_721_n N_VGND_c_827_n 0.0172656f $X=3.795 $Y=1.095 $X2=0
+ $Y2=0
cc_457 N_A_27_74#_c_722_n N_VGND_c_827_n 0.0161219f $X=3.88 $Y=0.515 $X2=0 $Y2=0
cc_458 N_A_27_74#_c_720_n N_VGND_c_828_n 0.00749631f $X=3 $Y=0.515 $X2=0 $Y2=0
cc_459 N_A_27_74#_c_713_n N_VGND_c_830_n 0.0145639f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_460 N_A_27_74#_c_716_n N_VGND_c_831_n 0.0109942f $X=1.21 $Y=0.515 $X2=0 $Y2=0
cc_461 N_A_27_74#_c_718_n N_VGND_c_832_n 0.00749631f $X=2.14 $Y=0.515 $X2=0
+ $Y2=0
cc_462 N_A_27_74#_c_722_n N_VGND_c_833_n 0.00749631f $X=3.88 $Y=0.515 $X2=0
+ $Y2=0
cc_463 N_A_27_74#_c_713_n N_VGND_c_834_n 0.0119984f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_464 N_A_27_74#_c_716_n N_VGND_c_834_n 0.00904371f $X=1.21 $Y=0.515 $X2=0
+ $Y2=0
cc_465 N_A_27_74#_c_718_n N_VGND_c_834_n 0.0062048f $X=2.14 $Y=0.515 $X2=0 $Y2=0
cc_466 N_A_27_74#_c_720_n N_VGND_c_834_n 0.0062048f $X=3 $Y=0.515 $X2=0 $Y2=0
cc_467 N_A_27_74#_c_722_n N_VGND_c_834_n 0.0062048f $X=3.88 $Y=0.515 $X2=0 $Y2=0
cc_468 N_A_27_74#_c_723_n N_VGND_c_834_n 0.00699877f $X=4.725 $Y=1 $X2=0 $Y2=0
cc_469 N_A_27_74#_c_723_n N_A_834_74#_M1006_d 0.0017828f $X=4.725 $Y=1 $X2=-0.19
+ $Y2=-0.245
cc_470 N_A_27_74#_c_724_n N_A_834_74#_M1019_d 0.00176891f $X=5.435 $Y=1.095
+ $X2=0 $Y2=0
cc_471 N_A_27_74#_M1020_s N_A_834_74#_c_918_n 0.00273752f $X=5.46 $Y=0.37 $X2=0
+ $Y2=0
cc_472 N_A_27_74#_c_724_n N_A_834_74#_c_918_n 0.0030313f $X=5.435 $Y=1.095 $X2=0
+ $Y2=0
cc_473 N_A_27_74#_c_725_n N_A_834_74#_c_918_n 0.0203278f $X=5.6 $Y=0.86 $X2=0
+ $Y2=0
cc_474 N_A_27_74#_c_724_n N_A_834_74#_c_919_n 0.0121616f $X=5.435 $Y=1.095 $X2=0
+ $Y2=0
cc_475 N_A_27_74#_c_725_n N_A_834_74#_c_919_n 0.027945f $X=5.6 $Y=0.86 $X2=0
+ $Y2=0
cc_476 N_A_27_74#_M1012_s N_A_834_74#_c_923_n 0.0018154f $X=4.6 $Y=0.37 $X2=0
+ $Y2=0
cc_477 N_A_27_74#_c_722_n N_A_834_74#_c_923_n 0.0127168f $X=3.88 $Y=0.515 $X2=0
+ $Y2=0
cc_478 N_A_27_74#_c_723_n N_A_834_74#_c_923_n 0.0411655f $X=4.725 $Y=1 $X2=0
+ $Y2=0
cc_479 N_A_27_74#_c_724_n N_A_834_74#_c_923_n 0.00491975f $X=5.435 $Y=1.095
+ $X2=0 $Y2=0
cc_480 N_A_27_74#_c_724_n N_A_834_74#_c_924_n 0.0132789f $X=5.435 $Y=1.095 $X2=0
+ $Y2=0
cc_481 N_VGND_c_833_n N_A_834_74#_c_920_n 0.0340834f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_482 N_VGND_c_834_n N_A_834_74#_c_920_n 0.0199188f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_483 N_VGND_c_833_n N_A_834_74#_c_921_n 0.05774f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_484 N_VGND_c_834_n N_A_834_74#_c_921_n 0.0327484f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_485 N_VGND_c_827_n N_A_834_74#_c_923_n 0.00285145f $X=3.43 $Y=0.635 $X2=0
+ $Y2=0
cc_486 N_VGND_c_833_n N_A_834_74#_c_923_n 0.122339f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_487 N_VGND_c_834_n N_A_834_74#_c_923_n 0.0682449f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_488 N_VGND_c_833_n N_A_834_74#_c_925_n 0.0236566f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_489 N_VGND_c_834_n N_A_834_74#_c_925_n 0.0128296f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_490 N_VGND_c_833_n N_A_834_74#_c_926_n 0.023391f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_491 N_VGND_c_834_n N_A_834_74#_c_926_n 0.0127797f $X=7.92 $Y=0 $X2=0 $Y2=0
