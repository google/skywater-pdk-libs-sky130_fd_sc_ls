* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
X0 VPWR A1 a_531_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X1 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X2 a_534_74# A1 Y VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X3 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X4 Y C1 a_114_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X5 a_114_368# B2 a_531_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X6 a_1326_74# B1 Y VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X7 Y B1 a_1326_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X8 a_1326_74# B1 Y VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X9 a_531_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X10 a_531_368# B2 a_114_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X11 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X12 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X13 a_1326_74# B2 VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X14 Y C1 a_114_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X15 VGND B2 a_1326_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X16 a_531_368# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X17 a_531_368# B1 a_114_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X18 a_531_368# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X19 VPWR A1 a_531_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X20 a_531_368# B1 a_114_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X21 Y B1 a_1326_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X22 a_1326_74# B2 VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X23 a_114_368# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X24 a_534_74# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X25 Y A1 a_534_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X26 VGND A2 a_534_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X27 a_114_368# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X28 a_531_368# B2 a_114_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X29 a_114_368# B2 a_531_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X30 VPWR A2 a_531_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X31 VGND B2 a_1326_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X32 a_114_368# B1 a_531_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X33 Y A1 a_534_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X34 a_531_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X35 a_534_74# A1 Y VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X36 VPWR A2 a_531_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X37 a_114_368# B1 a_531_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X38 a_534_74# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X39 VGND A2 a_534_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
.ends
