* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__dlxbn_1 D GATE_N VGND VNB VPB VPWR Q Q_N
X0 a_575_79# a_232_82# a_653_79# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X1 VPWR a_1347_424# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X2 VPWR GATE_N a_232_82# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X3 a_571_392# a_343_80# a_653_79# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 a_653_79# a_343_80# a_852_123# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_653_79# a_232_82# a_805_392# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 a_343_80# a_232_82# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X7 VPWR a_27_120# a_571_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 a_343_80# a_232_82# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X9 a_805_392# a_863_294# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X10 VGND GATE_N a_232_82# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X11 Q a_863_294# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X12 VGND a_27_120# a_575_79# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X13 VPWR a_653_79# a_863_294# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X14 a_852_123# a_863_294# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 Q a_863_294# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X16 a_27_120# D VGND VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X17 VGND a_1347_424# Q_N VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X18 VGND a_653_79# a_863_294# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X19 VGND a_863_294# a_1347_424# VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X20 VPWR a_863_294# a_1347_424# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X21 a_27_120# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
.ends
