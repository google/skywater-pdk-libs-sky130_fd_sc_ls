* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
X0 X a_91_48# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X1 a_968_391# A2 a_91_48# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 X a_91_48# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X3 VPWR C1 a_91_48# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X4 VPWR a_91_48# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X5 VPWR B1 a_91_48# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X6 a_510_125# B1 a_597_125# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X7 a_91_48# A2 a_968_391# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 a_91_48# C1 a_597_125# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X9 a_510_125# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X10 VGND a_91_48# X VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X11 a_597_125# B1 a_510_125# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X12 X a_91_48# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X13 VPWR a_91_48# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X14 a_597_125# C1 a_91_48# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X15 a_91_48# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X16 VGND A1 a_510_125# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X17 VGND A2 a_510_125# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X18 a_91_48# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X19 VGND a_91_48# X VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X20 a_968_391# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X21 X a_91_48# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X22 a_510_125# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X23 VPWR A1 a_968_391# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends
