# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_ls__sdfsbp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_ls__sdfsbp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  17.76000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.385000 0.440000 1.795000 1.230000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 16.865000 1.820000 17.225000 2.980000 ;
        RECT 16.885000 0.350000 17.225000 1.130000 ;
        RECT 17.055000 1.130000 17.225000 1.820000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.558000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 14.850000 0.350000 15.235000 1.410000 ;
        RECT 14.850000 1.410000 15.105000 2.980000 ;
    END
  END Q_N
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.805000 0.950000 3.205000 1.620000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 1.400000 2.295000 1.570000 ;
        RECT 0.425000 1.570000 1.085000 1.800000 ;
        RECT 1.965000 0.900000 2.295000 1.400000 ;
    END
  END SCE
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT  7.775000 1.550000  8.065000 1.595000 ;
        RECT  7.775000 1.595000 13.345000 1.735000 ;
        RECT  7.775000 1.735000  8.065000 1.780000 ;
        RECT 13.055000 1.550000 13.345000 1.595000 ;
        RECT 13.055000 1.735000 13.345000 1.780000 ;
    END
  END SET_B
  PIN VNB
    PORT
      LAYER pwell ;
        RECT 0.000000 0.000000 17.760000 0.245000 ;
    END
  END VNB
  PIN VPB
    PORT
      LAYER nwell ;
        RECT -0.190000 1.660000 17.950000 3.520000 ;
    END
  END VPB
  PIN CLK
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.715000 1.180000 4.195000 1.550000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 17.760000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 17.760000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 17.760000 0.085000 ;
      RECT  0.000000  3.245000 17.760000 3.415000 ;
      RECT  0.085000  0.350000  0.445000 0.900000 ;
      RECT  0.085000  0.900000  1.145000 1.230000 ;
      RECT  0.085000  1.230000  0.255000 1.970000 ;
      RECT  0.085000  1.970000  2.105000 2.140000 ;
      RECT  0.085000  2.140000  0.465000 2.980000 ;
      RECT  0.615000  0.085000  1.020000 0.680000 ;
      RECT  0.635000  2.310000  0.965000 3.245000 ;
      RECT  1.505000  2.310000  3.885000 2.480000 ;
      RECT  1.505000  2.480000  1.955000 2.980000 ;
      RECT  1.775000  1.810000  2.105000 1.970000 ;
      RECT  1.965000  0.400000  2.350000 0.560000 ;
      RECT  1.965000  0.560000  2.635000 0.730000 ;
      RECT  2.465000  0.730000  2.635000 2.310000 ;
      RECT  2.495000  2.650000  2.845000 3.245000 ;
      RECT  2.840000  0.085000  3.170000 0.780000 ;
      RECT  3.075000  1.790000  4.720000 1.960000 ;
      RECT  3.075000  1.960000  3.545000 2.140000 ;
      RECT  3.375000  0.340000  3.650000 1.010000 ;
      RECT  3.375000  1.010000  3.545000 1.790000 ;
      RECT  3.525000  2.650000  4.220000 3.245000 ;
      RECT  3.715000  2.130000  5.370000 2.300000 ;
      RECT  3.715000  2.300000  3.885000 2.310000 ;
      RECT  3.830000  0.085000  4.160000 1.010000 ;
      RECT  4.330000  0.255000  5.560000 0.425000 ;
      RECT  4.330000  0.425000  4.660000 1.010000 ;
      RECT  4.390000  1.350000  4.720000 1.790000 ;
      RECT  4.390000  2.470000  4.720000 2.905000 ;
      RECT  4.390000  2.905000  6.240000 3.075000 ;
      RECT  4.890000  0.595000  5.220000 0.845000 ;
      RECT  4.890000  0.845000  5.060000 2.130000 ;
      RECT  4.890000  2.300000  5.370000 2.735000 ;
      RECT  5.230000  1.290000  5.560000 1.960000 ;
      RECT  5.390000  0.425000  5.560000 1.290000 ;
      RECT  5.540000  2.295000  5.900000 2.735000 ;
      RECT  5.730000  0.470000  6.645000 0.800000 ;
      RECT  5.730000  0.800000  5.900000 2.295000 ;
      RECT  6.070000  0.970000  6.305000 2.165000 ;
      RECT  6.070000  2.165000  7.325000 2.335000 ;
      RECT  6.070000  2.335000  6.240000 2.905000 ;
      RECT  6.410000  2.505000  6.985000 3.245000 ;
      RECT  6.475000  0.800000  6.645000 1.395000 ;
      RECT  6.475000  1.395000  7.665000 1.565000 ;
      RECT  6.635000  1.735000  7.665000 1.995000 ;
      RECT  6.815000  0.085000  7.150000 0.700000 ;
      RECT  6.815000  0.870000  7.710000 1.040000 ;
      RECT  6.815000  1.040000  7.145000 1.225000 ;
      RECT  7.155000  2.335000  7.325000 2.905000 ;
      RECT  7.155000  2.905000  8.165000 3.075000 ;
      RECT  7.355000  1.210000  8.050000 1.380000 ;
      RECT  7.355000  1.380000  7.665000 1.395000 ;
      RECT  7.380000  0.350000  7.710000 0.870000 ;
      RECT  7.495000  1.995000  7.665000 2.295000 ;
      RECT  7.495000  2.295000  7.825000 2.735000 ;
      RECT  7.835000  1.550000  8.225000 1.880000 ;
      RECT  7.880000  0.900000  8.860000 1.175000 ;
      RECT  7.880000  1.175000  8.050000 1.210000 ;
      RECT  7.995000  2.050000  8.565000 2.220000 ;
      RECT  7.995000  2.220000  8.165000 2.905000 ;
      RECT  8.200000  0.085000  8.530000 0.680000 ;
      RECT  8.335000  2.390000  8.665000 3.245000 ;
      RECT  8.395000  1.345000 11.390000 1.515000 ;
      RECT  8.395000  1.515000  8.565000 2.050000 ;
      RECT  8.735000  1.685000  9.065000 1.700000 ;
      RECT  8.735000  1.700000 12.050000 1.870000 ;
      RECT  8.735000  1.870000  9.065000 1.960000 ;
      RECT  8.925000  2.130000 10.125000 2.300000 ;
      RECT  8.925000  2.300000  9.255000 2.980000 ;
      RECT  9.030000  0.350000  9.280000 1.005000 ;
      RECT  9.030000  1.005000 10.210000 1.175000 ;
      RECT  9.425000  2.470000  9.675000 3.245000 ;
      RECT  9.450000  0.085000  9.780000 0.835000 ;
      RECT  9.875000  2.100000 10.125000 2.130000 ;
      RECT  9.875000  2.300000 10.125000 2.905000 ;
      RECT  9.875000  2.905000 11.105000 3.075000 ;
      RECT  9.960000  0.255000 11.210000 0.425000 ;
      RECT  9.960000  0.425000 10.210000 1.005000 ;
      RECT 10.325000  2.040000 12.390000 2.140000 ;
      RECT 10.325000  2.140000 13.975000 2.210000 ;
      RECT 10.325000  2.210000 10.575000 2.700000 ;
      RECT 10.380000  0.595000 10.710000 0.860000 ;
      RECT 10.380000  0.860000 11.550000 1.030000 ;
      RECT 10.380000  1.200000 11.390000 1.345000 ;
      RECT 10.380000  1.515000 11.390000 1.530000 ;
      RECT 10.775000  2.380000 11.105000 2.905000 ;
      RECT 10.880000  0.425000 11.210000 0.690000 ;
      RECT 11.365000  2.385000 11.620000 2.885000 ;
      RECT 11.365000  2.885000 12.740000 3.055000 ;
      RECT 11.380000  0.400000 12.390000 0.730000 ;
      RECT 11.380000  0.730000 11.550000 0.860000 ;
      RECT 11.720000  0.900000 12.050000 1.700000 ;
      RECT 11.820000  2.210000 13.975000 2.310000 ;
      RECT 11.820000  2.310000 12.220000 2.715000 ;
      RECT 12.220000  0.730000 12.390000 2.040000 ;
      RECT 12.410000  2.520000 12.740000 2.885000 ;
      RECT 12.565000  0.960000 14.315000 1.130000 ;
      RECT 12.565000  1.130000 12.895000 1.960000 ;
      RECT 12.940000  2.520000 13.110000 3.245000 ;
      RECT 13.085000  1.300000 13.435000 1.970000 ;
      RECT 13.260000  0.085000 13.590000 0.790000 ;
      RECT 13.310000  2.310000 13.640000 2.980000 ;
      RECT 13.645000  1.300000 13.975000 2.140000 ;
      RECT 13.770000  0.350000 14.100000 0.960000 ;
      RECT 13.870000  2.480000 14.315000 2.910000 ;
      RECT 14.145000  1.130000 14.315000 2.480000 ;
      RECT 14.350000  0.085000 14.680000 0.790000 ;
      RECT 14.485000  1.820000 14.655000 3.245000 ;
      RECT 15.305000  1.820000 15.635000 3.245000 ;
      RECT 15.405000  0.085000 15.655000 1.130000 ;
      RECT 15.865000  0.450000 16.220000 1.300000 ;
      RECT 15.865000  1.300000 16.885000 1.630000 ;
      RECT 15.865000  1.630000 16.195000 2.860000 ;
      RECT 16.415000  1.820000 16.665000 3.245000 ;
      RECT 16.455000  0.085000 16.705000 1.130000 ;
      RECT 17.395000  0.085000 17.645000 1.130000 ;
      RECT 17.395000  1.820000 17.645000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  1.580000  8.005000 1.750000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  1.580000 13.285000 1.750000 ;
      RECT 13.115000  3.245000 13.285000 3.415000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.245000 13.765000 3.415000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000  3.245000 14.245000 3.415000 ;
      RECT 14.555000 -0.085000 14.725000 0.085000 ;
      RECT 14.555000  3.245000 14.725000 3.415000 ;
      RECT 15.035000 -0.085000 15.205000 0.085000 ;
      RECT 15.035000  3.245000 15.205000 3.415000 ;
      RECT 15.515000 -0.085000 15.685000 0.085000 ;
      RECT 15.515000  3.245000 15.685000 3.415000 ;
      RECT 15.995000 -0.085000 16.165000 0.085000 ;
      RECT 15.995000  3.245000 16.165000 3.415000 ;
      RECT 16.475000 -0.085000 16.645000 0.085000 ;
      RECT 16.475000  3.245000 16.645000 3.415000 ;
      RECT 16.955000 -0.085000 17.125000 0.085000 ;
      RECT 16.955000  3.245000 17.125000 3.415000 ;
      RECT 17.435000 -0.085000 17.605000 0.085000 ;
      RECT 17.435000  3.245000 17.605000 3.415000 ;
  END
END sky130_fd_sc_ls__sdfsbp_2
END LIBRARY
