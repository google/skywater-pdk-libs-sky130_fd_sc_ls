* File: sky130_fd_sc_ls__nor3b_2.pex.spice
* Created: Wed Sep  2 11:15:10 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__NOR3B_2%C_N 3 5 7 8
c31 5 0 2.87358e-19 $X=0.5 $Y=1.885
r32 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.59
+ $Y=1.615 $X2=0.59 $Y2=1.615
r33 8 12 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=0.72 $Y=1.615
+ $X2=0.59 $Y2=1.615
r34 5 11 55.1302 $w=3.05e-07 $l=3.08286e-07 $layer=POLY_cond $X=0.5 $Y=1.885
+ $X2=0.582 $Y2=1.615
r35 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.5 $Y=1.885 $X2=0.5
+ $Y2=2.46
r36 1 11 38.5368 $w=3.05e-07 $l=2.01879e-07 $layer=POLY_cond $X=0.5 $Y=1.45
+ $X2=0.582 $Y2=1.615
r37 1 3 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=0.5 $Y=1.45 $X2=0.5
+ $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_LS__NOR3B_2%A_27_392# 1 2 7 9 10 12 13 15 17 18 20 23 27
+ 29 33 35 36 37 46
c82 37 0 1.05511e-19 $X=1.17 $Y=1.195
c83 18 0 1.8273e-19 $X=1.95 $Y=1.765
c84 13 0 1.49881e-19 $X=1.515 $Y=1.22
c85 10 0 1.81847e-19 $X=1.5 $Y=1.765
r86 45 46 2.01955 $w=3.58e-07 $l=1.5e-08 $layer=POLY_cond $X=1.5 $Y=1.492
+ $X2=1.515 $Y2=1.492
r87 41 45 44.4302 $w=3.58e-07 $l=3.3e-07 $layer=POLY_cond $X=1.17 $Y=1.492
+ $X2=1.5 $Y2=1.492
r88 41 43 13.4637 $w=3.58e-07 $l=1e-07 $layer=POLY_cond $X=1.17 $Y=1.492
+ $X2=1.07 $Y2=1.492
r89 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.17
+ $Y=1.385 $X2=1.17 $Y2=1.385
r90 37 40 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=1.17 $Y=1.195
+ $X2=1.17 $Y2=1.385
r91 34 35 3.01551 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.45 $Y=1.195
+ $X2=0.267 $Y2=1.195
r92 33 37 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.005 $Y=1.195
+ $X2=1.17 $Y2=1.195
r93 33 34 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=1.005 $Y=1.195
+ $X2=0.45 $Y2=1.195
r94 29 31 29.3349 $w=2.73e-07 $l=7e-07 $layer=LI1_cond $X=0.222 $Y=2.115
+ $X2=0.222 $Y2=2.815
r95 27 36 7.41084 $w=2.73e-07 $l=1.37e-07 $layer=LI1_cond $X=0.222 $Y=2.087
+ $X2=0.222 $Y2=1.95
r96 27 29 1.1734 $w=2.73e-07 $l=2.8e-08 $layer=LI1_cond $X=0.222 $Y=2.087
+ $X2=0.222 $Y2=2.115
r97 25 35 3.49088 $w=2.67e-07 $l=1.32868e-07 $layer=LI1_cond $X=0.17 $Y=1.28
+ $X2=0.267 $Y2=1.195
r98 25 36 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.17 $Y=1.28
+ $X2=0.17 $Y2=1.95
r99 21 35 3.49088 $w=2.67e-07 $l=8.5e-08 $layer=LI1_cond $X=0.267 $Y=1.11
+ $X2=0.267 $Y2=1.195
r100 21 23 18.7864 $w=3.63e-07 $l=5.95e-07 $layer=LI1_cond $X=0.267 $Y=1.11
+ $X2=0.267 $Y2=0.515
r101 18 20 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.95 $Y=1.765
+ $X2=1.95 $Y2=2.4
r102 17 18 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.95 $Y=1.675
+ $X2=1.95 $Y2=1.765
r103 16 46 58.567 $w=3.58e-07 $l=4.35e-07 $layer=POLY_cond $X=1.95 $Y=1.492
+ $X2=1.515 $Y2=1.492
r104 16 17 56.3629 $w=1.8e-07 $l=1.45e-07 $layer=POLY_cond $X=1.95 $Y=1.53
+ $X2=1.95 $Y2=1.675
r105 13 46 23.1716 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=1.515 $Y=1.22
+ $X2=1.515 $Y2=1.492
r106 13 15 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.515 $Y=1.22
+ $X2=1.515 $Y2=0.74
r107 10 45 23.1716 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=1.5 $Y=1.765
+ $X2=1.5 $Y2=1.492
r108 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.5 $Y=1.765
+ $X2=1.5 $Y2=2.4
r109 7 43 23.1716 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=1.07 $Y=1.22
+ $X2=1.07 $Y2=1.492
r110 7 9 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.07 $Y=1.22 $X2=1.07
+ $Y2=0.74
r111 2 31 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.275 $Y2=2.815
r112 2 29 400 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.275 $Y2=2.115
r113 1 23 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.14
+ $Y=0.37 $X2=0.285 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__NOR3B_2%B 3 5 7 10 12 14 15 17 19
c52 15 0 5.79615e-20 $X=3.12 $Y=1.665
c53 12 0 5.27684e-20 $X=2.85 $Y=1.765
r54 27 28 4.46296 $w=3.78e-07 $l=3.5e-08 $layer=POLY_cond $X=2.815 $Y=1.557
+ $X2=2.85 $Y2=1.557
r55 25 27 5.7381 $w=3.78e-07 $l=4.5e-08 $layer=POLY_cond $X=2.77 $Y=1.557
+ $X2=2.815 $Y2=1.557
r56 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.77
+ $Y=1.515 $X2=2.77 $Y2=1.515
r57 23 25 47.1799 $w=3.78e-07 $l=3.7e-07 $layer=POLY_cond $X=2.4 $Y=1.557
+ $X2=2.77 $Y2=1.557
r58 22 23 1.9127 $w=3.78e-07 $l=1.5e-08 $layer=POLY_cond $X=2.385 $Y=1.557
+ $X2=2.4 $Y2=1.557
r59 20 26 9.11234 $w=4.28e-07 $l=3.4e-07 $layer=LI1_cond $X=3.11 $Y=1.565
+ $X2=2.77 $Y2=1.565
r60 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.11
+ $Y=1.515 $X2=3.11 $Y2=1.515
r61 17 28 12.3802 $w=3.78e-07 $l=1.08995e-07 $layer=POLY_cond $X=2.94 $Y=1.515
+ $X2=2.85 $Y2=1.557
r62 17 19 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=2.94 $Y=1.515
+ $X2=3.11 $Y2=1.515
r63 15 20 0.26801 $w=4.28e-07 $l=1e-08 $layer=LI1_cond $X=3.12 $Y=1.565 $X2=3.11
+ $Y2=1.565
r64 12 28 24.4846 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.85 $Y=1.765
+ $X2=2.85 $Y2=1.557
r65 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.85 $Y=1.765
+ $X2=2.85 $Y2=2.4
r66 8 27 24.4846 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.815 $Y=1.35
+ $X2=2.815 $Y2=1.557
r67 8 10 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.815 $Y=1.35
+ $X2=2.815 $Y2=0.74
r68 5 23 24.4846 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.4 $Y=1.765 $X2=2.4
+ $Y2=1.557
r69 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.4 $Y=1.765 $X2=2.4
+ $Y2=2.4
r70 1 22 24.4846 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.385 $Y=1.35
+ $X2=2.385 $Y2=1.557
r71 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.385 $Y=1.35
+ $X2=2.385 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__NOR3B_2%A 3 5 7 10 12 14 15 16 17 26
c46 17 0 5.27684e-20 $X=4.56 $Y=1.665
c47 10 0 1.81748e-19 $X=4.285 $Y=0.74
c48 5 0 5.79615e-20 $X=3.85 $Y=1.765
r49 26 27 1.93834 $w=3.73e-07 $l=1.5e-08 $layer=POLY_cond $X=4.285 $Y=1.557
+ $X2=4.3 $Y2=1.557
r50 24 26 11.63 $w=3.73e-07 $l=9e-08 $layer=POLY_cond $X=4.195 $Y=1.557
+ $X2=4.285 $Y2=1.557
r51 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.195
+ $Y=1.515 $X2=4.195 $Y2=1.515
r52 22 24 44.5818 $w=3.73e-07 $l=3.45e-07 $layer=POLY_cond $X=3.85 $Y=1.557
+ $X2=4.195 $Y2=1.557
r53 21 22 5.81501 $w=3.73e-07 $l=4.5e-08 $layer=POLY_cond $X=3.805 $Y=1.557
+ $X2=3.85 $Y2=1.557
r54 17 25 9.78236 $w=4.28e-07 $l=3.65e-07 $layer=LI1_cond $X=4.56 $Y=1.565
+ $X2=4.195 $Y2=1.565
r55 16 25 3.08211 $w=4.28e-07 $l=1.15e-07 $layer=LI1_cond $X=4.08 $Y=1.565
+ $X2=4.195 $Y2=1.565
r56 15 16 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=3.6 $Y=1.565
+ $X2=4.08 $Y2=1.565
r57 12 27 24.162 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=4.3 $Y=1.765 $X2=4.3
+ $Y2=1.557
r58 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.3 $Y=1.765
+ $X2=4.3 $Y2=2.4
r59 8 26 24.162 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.285 $Y=1.35
+ $X2=4.285 $Y2=1.557
r60 8 10 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.285 $Y=1.35
+ $X2=4.285 $Y2=0.74
r61 5 22 24.162 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.85 $Y=1.765
+ $X2=3.85 $Y2=1.557
r62 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.85 $Y=1.765
+ $X2=3.85 $Y2=2.4
r63 1 21 24.162 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.805 $Y=1.35
+ $X2=3.805 $Y2=1.557
r64 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.805 $Y=1.35
+ $X2=3.805 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__NOR3B_2%VPWR 1 2 3 12 18 20 22 26 28 33 41 47 50 54
r55 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r56 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r57 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r58 45 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r59 45 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r60 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r61 42 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.79 $Y=3.33
+ $X2=3.625 $Y2=3.33
r62 42 44 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=3.79 $Y=3.33
+ $X2=4.08 $Y2=3.33
r63 41 53 4.14492 $w=1.7e-07 $l=1.87e-07 $layer=LI1_cond $X=4.425 $Y=3.33
+ $X2=4.612 $Y2=3.33
r64 41 44 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=4.425 $Y=3.33
+ $X2=4.08 $Y2=3.33
r65 40 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r66 39 40 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r67 37 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r68 36 39 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=3.12 $Y2=3.33
r69 36 37 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r70 34 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.89 $Y=3.33
+ $X2=0.725 $Y2=3.33
r71 34 36 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.89 $Y=3.33 $X2=1.2
+ $Y2=3.33
r72 33 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.46 $Y=3.33
+ $X2=3.625 $Y2=3.33
r73 33 39 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=3.46 $Y=3.33
+ $X2=3.12 $Y2=3.33
r74 31 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r75 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r76 28 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.56 $Y=3.33
+ $X2=0.725 $Y2=3.33
r77 28 30 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.56 $Y=3.33 $X2=0.24
+ $Y2=3.33
r78 26 40 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=3.12 $Y2=3.33
r79 26 37 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=2.4 $Y=3.33 $X2=1.2
+ $Y2=3.33
r80 22 25 30.4419 $w=2.63e-07 $l=7e-07 $layer=LI1_cond $X=4.557 $Y=2.115
+ $X2=4.557 $Y2=2.815
r81 20 53 3.10315 $w=2.65e-07 $l=1.09087e-07 $layer=LI1_cond $X=4.557 $Y=3.245
+ $X2=4.612 $Y2=3.33
r82 20 25 18.7 $w=2.63e-07 $l=4.3e-07 $layer=LI1_cond $X=4.557 $Y=3.245
+ $X2=4.557 $Y2=2.815
r83 16 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.625 $Y=3.245
+ $X2=3.625 $Y2=3.33
r84 16 18 29.6841 $w=3.28e-07 $l=8.5e-07 $layer=LI1_cond $X=3.625 $Y=3.245
+ $X2=3.625 $Y2=2.395
r85 12 15 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=0.725 $Y=2.115
+ $X2=0.725 $Y2=2.815
r86 10 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.725 $Y=3.245
+ $X2=0.725 $Y2=3.33
r87 10 15 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.725 $Y=3.245
+ $X2=0.725 $Y2=2.815
r88 3 25 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=4.375
+ $Y=1.84 $X2=4.525 $Y2=2.815
r89 3 22 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=4.375
+ $Y=1.84 $X2=4.525 $Y2=2.115
r90 2 18 300 $w=1.7e-07 $l=6.21068e-07 $layer=licon1_PDIFF $count=2 $X=3.485
+ $Y=1.84 $X2=3.625 $Y2=2.395
r91 1 15 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=0.575
+ $Y=1.96 $X2=0.725 $Y2=2.815
r92 1 12 400 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=1 $X=0.575
+ $Y=1.96 $X2=0.725 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_LS__NOR3B_2%A_227_368# 1 2 3 12 16 17 20 24 28 30
r44 26 28 19.2074 $w=2.68e-07 $l=4.5e-07 $layer=LI1_cond $X=3.105 $Y=2.905
+ $X2=3.105 $Y2=2.455
r45 25 30 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.29 $Y=2.99 $X2=2.15
+ $Y2=2.99
r46 24 26 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=2.97 $Y=2.99
+ $X2=3.105 $Y2=2.905
r47 24 25 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.97 $Y=2.99
+ $X2=2.29 $Y2=2.99
r48 20 23 34.1617 $w=2.78e-07 $l=8.3e-07 $layer=LI1_cond $X=2.15 $Y=1.985
+ $X2=2.15 $Y2=2.815
r49 18 30 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.15 $Y=2.905
+ $X2=2.15 $Y2=2.99
r50 18 23 3.70428 $w=2.78e-07 $l=9e-08 $layer=LI1_cond $X=2.15 $Y=2.905 $X2=2.15
+ $Y2=2.815
r51 16 30 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.01 $Y=2.99 $X2=2.15
+ $Y2=2.99
r52 16 17 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=2.01 $Y=2.99
+ $X2=1.44 $Y2=2.99
r53 12 15 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=1.275 $Y=1.985
+ $X2=1.275 $Y2=2.815
r54 10 17 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.275 $Y=2.905
+ $X2=1.44 $Y2=2.99
r55 10 15 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=1.275 $Y=2.905
+ $X2=1.275 $Y2=2.815
r56 3 28 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=2.925
+ $Y=1.84 $X2=3.075 $Y2=2.455
r57 2 23 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.025
+ $Y=1.84 $X2=2.175 $Y2=2.815
r58 2 20 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.025
+ $Y=1.84 $X2=2.175 $Y2=1.985
r59 1 15 400 $w=1.7e-07 $l=1.04265e-06 $layer=licon1_PDIFF $count=1 $X=1.135
+ $Y=1.84 $X2=1.275 $Y2=2.815
r60 1 12 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.135
+ $Y=1.84 $X2=1.275 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_LS__NOR3B_2%Y 1 2 3 4 15 19 23 25 29 31 33 34 35 38
c61 25 0 1.81748e-19 $X=3.925 $Y=1.045
c62 15 0 1.49881e-19 $X=1.285 $Y=0.515
r63 38 45 4.30525 $w=3.6e-07 $l=8.9861e-08 $layer=LI1_cond $X=1.81 $Y=0.95
+ $X2=1.725 $Y2=0.94
r64 35 38 11.2043 $w=3.58e-07 $l=3.5e-07 $layer=LI1_cond $X=2.16 $Y=0.95
+ $X2=1.81 $Y2=0.95
r65 34 45 2.31646 $w=2.37e-07 $l=4.5e-08 $layer=LI1_cond $X=1.68 $Y=0.94
+ $X2=1.725 $Y2=0.94
r66 31 35 11.0442 $w=3.58e-07 $l=3.45e-07 $layer=LI1_cond $X=2.505 $Y=0.95
+ $X2=2.16 $Y2=0.95
r67 31 33 3.88469 $w=2.65e-07 $l=9.5e-08 $layer=LI1_cond $X=2.505 $Y=0.95
+ $X2=2.6 $Y2=0.95
r68 27 29 19.7245 $w=2.58e-07 $l=4.45e-07 $layer=LI1_cond $X=4.055 $Y=0.96
+ $X2=4.055 $Y2=0.515
r69 26 33 3.88469 $w=2.65e-07 $l=1.3435e-07 $layer=LI1_cond $X=2.695 $Y=1.045
+ $X2=2.6 $Y2=0.95
r70 25 27 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=3.925 $Y=1.045
+ $X2=4.055 $Y2=0.96
r71 25 26 80.246 $w=1.68e-07 $l=1.23e-06 $layer=LI1_cond $X=3.925 $Y=1.045
+ $X2=2.695 $Y2=1.045
r72 21 33 2.5638 $w=1.9e-07 $l=1.8e-07 $layer=LI1_cond $X=2.6 $Y=0.77 $X2=2.6
+ $Y2=0.95
r73 21 23 14.8852 $w=1.88e-07 $l=2.55e-07 $layer=LI1_cond $X=2.6 $Y=0.77 $X2=2.6
+ $Y2=0.515
r74 17 45 2.684 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.725 $Y=1.13 $X2=1.725
+ $Y2=0.94
r75 17 19 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=1.725 $Y=1.13
+ $X2=1.725 $Y2=1.985
r76 13 34 21.7747 $w=2.37e-07 $l=4.23e-07 $layer=LI1_cond $X=1.257 $Y=0.94
+ $X2=1.68 $Y2=0.94
r77 13 15 10.6863 $w=2.73e-07 $l=2.55e-07 $layer=LI1_cond $X=1.257 $Y=0.77
+ $X2=1.257 $Y2=0.515
r78 4 19 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=1.575
+ $Y=1.84 $X2=1.725 $Y2=1.985
r79 3 29 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.88
+ $Y=0.37 $X2=4.02 $Y2=0.515
r80 2 33 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=2.46
+ $Y=0.37 $X2=2.6 $Y2=0.965
r81 2 23 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.46
+ $Y=0.37 $X2=2.6 $Y2=0.515
r82 1 13 182 $w=1.7e-07 $l=5.50568e-07 $layer=licon1_NDIFF $count=1 $X=1.145
+ $Y=0.37 $X2=1.285 $Y2=0.855
r83 1 15 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1.145
+ $Y=0.37 $X2=1.285 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__NOR3B_2%A_495_368# 1 2 9 11 13 16
c27 16 0 1.8273e-19 $X=2.625 $Y=2.035
r28 11 18 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.115 $Y=2.12
+ $X2=4.115 $Y2=2.035
r29 11 13 14.7513 $w=2.48e-07 $l=3.2e-07 $layer=LI1_cond $X=4.115 $Y=2.12
+ $X2=4.115 $Y2=2.44
r30 10 16 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.79 $Y=2.035
+ $X2=2.625 $Y2=2.035
r31 9 18 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.99 $Y=2.035
+ $X2=4.115 $Y2=2.035
r32 9 10 78.2888 $w=1.68e-07 $l=1.2e-06 $layer=LI1_cond $X=3.99 $Y=2.035
+ $X2=2.79 $Y2=2.035
r33 2 18 600 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=3.925
+ $Y=1.84 $X2=4.075 $Y2=2.035
r34 2 13 300 $w=1.7e-07 $l=6.7082e-07 $layer=licon1_PDIFF $count=2 $X=3.925
+ $Y=1.84 $X2=4.075 $Y2=2.44
r35 1 16 300 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=2 $X=2.475
+ $Y=1.84 $X2=2.625 $Y2=2.035
.ends

.subckt PM_SKY130_FD_SC_LS__NOR3B_2%VGND 1 2 3 4 15 17 19 21 23 38 44 49 55 58
+ 62 65
r65 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r66 60 62 11.8599 $w=8.53e-07 $l=1.55e-07 $layer=LI1_cond $X=3.6 $Y=0.342
+ $X2=3.755 $Y2=0.342
r67 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r68 57 60 0.14269 $w=8.53e-07 $l=1e-08 $layer=LI1_cond $X=3.59 $Y=0.342 $X2=3.6
+ $Y2=0.342
r69 57 58 19.9932 $w=8.53e-07 $l=7.25e-07 $layer=LI1_cond $X=3.59 $Y=0.342
+ $X2=2.865 $Y2=0.342
r70 54 55 10.7086 $w=6.83e-07 $l=1.65e-07 $layer=LI1_cond $X=2.17 $Y=0.257
+ $X2=2.335 $Y2=0.257
r71 51 54 0.17461 $w=6.83e-07 $l=1e-08 $layer=LI1_cond $X=2.16 $Y=0.257 $X2=2.17
+ $Y2=0.257
r72 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r73 48 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r74 47 51 8.38128 $w=6.83e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=0.257
+ $X2=2.16 $Y2=0.257
r75 47 49 9.83558 $w=6.83e-07 $l=1.15e-07 $layer=LI1_cond $X=1.68 $Y=0.257
+ $X2=1.565 $Y2=0.257
r76 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r77 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r78 42 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r79 42 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r80 41 62 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=4.08 $Y=0 $X2=3.755
+ $Y2=0
r81 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r82 38 64 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=4.355 $Y=0 $X2=4.577
+ $Y2=0
r83 38 41 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.355 $Y=0 $X2=4.08
+ $Y2=0
r84 37 61 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r85 36 58 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.64 $Y=0 $X2=2.865
+ $Y2=0
r86 36 55 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.64 $Y=0 $X2=2.335
+ $Y2=0
r87 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r88 32 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r89 32 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r90 31 49 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=1.565
+ $Y2=0
r91 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r92 29 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.95 $Y=0 $X2=0.785
+ $Y2=0
r93 29 31 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.95 $Y=0 $X2=1.2
+ $Y2=0
r94 26 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r95 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r96 23 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.62 $Y=0 $X2=0.785
+ $Y2=0
r97 23 25 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=0.62 $Y=0 $X2=0.24
+ $Y2=0
r98 21 37 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=2.64
+ $Y2=0
r99 21 52 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=2.16
+ $Y2=0
r100 17 64 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=4.52 $Y=0.085
+ $X2=4.577 $Y2=0
r101 17 19 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=4.52 $Y=0.085
+ $X2=4.52 $Y2=0.515
r102 13 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.785 $Y=0.085
+ $X2=0.785 $Y2=0
r103 13 15 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.785 $Y=0.085
+ $X2=0.785 $Y2=0.515
r104 4 19 91 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=2 $X=4.36
+ $Y=0.37 $X2=4.52 $Y2=0.515
r105 3 57 91 $w=1.7e-07 $l=8.09012e-07 $layer=licon1_NDIFF $count=2 $X=2.89
+ $Y=0.37 $X2=3.59 $Y2=0.605
r106 2 54 91 $w=1.7e-07 $l=6.4846e-07 $layer=licon1_NDIFF $count=2 $X=1.59
+ $Y=0.37 $X2=2.17 $Y2=0.515
r107 1 15 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=0.575
+ $Y=0.37 $X2=0.785 $Y2=0.515
.ends

