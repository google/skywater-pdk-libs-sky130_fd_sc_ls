* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__or3b_1 A B C_N VGND VNB VPB VPWR X
X0 VGND B a_239_74# VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X1 a_239_74# A VGND VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X2 VPWR C_N a_124_424# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X3 a_239_74# a_124_424# a_368_391# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 a_452_391# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_239_74# a_124_424# VGND VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X6 VGND C_N a_124_424# VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X7 VGND a_239_74# X VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X8 a_368_391# B a_452_391# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 VPWR a_239_74# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
.ends
