* File: sky130_fd_sc_ls__einvn_2.pxi.spice
* Created: Wed Sep  2 11:06:43 2020
* 
x_PM_SKY130_FD_SC_LS__EINVN_2%A_115_464# N_A_115_464#_M1009_d
+ N_A_115_464#_M1006_d N_A_115_464#_c_68_n N_A_115_464#_M1001_g
+ N_A_115_464#_c_70_n N_A_115_464#_M1004_g N_A_115_464#_c_72_n
+ N_A_115_464#_c_78_n N_A_115_464#_c_73_n N_A_115_464#_c_74_n
+ N_A_115_464#_c_75_n N_A_115_464#_c_76_n N_A_115_464#_c_77_n
+ PM_SKY130_FD_SC_LS__EINVN_2%A_115_464#
x_PM_SKY130_FD_SC_LS__EINVN_2%TE_B N_TE_B_c_129_n N_TE_B_c_134_n N_TE_B_M1006_g
+ N_TE_B_M1009_g N_TE_B_c_136_n N_TE_B_c_137_n N_TE_B_c_138_n N_TE_B_M1000_g
+ N_TE_B_c_139_n N_TE_B_c_140_n N_TE_B_M1007_g N_TE_B_c_141_n TE_B TE_B
+ N_TE_B_c_131_n N_TE_B_c_132_n PM_SKY130_FD_SC_LS__EINVN_2%TE_B
x_PM_SKY130_FD_SC_LS__EINVN_2%A N_A_c_194_n N_A_M1002_g N_A_c_195_n N_A_c_202_n
+ N_A_M1003_g N_A_c_196_n N_A_c_197_n N_A_M1008_g N_A_c_198_n N_A_M1005_g
+ N_A_c_199_n A A PM_SKY130_FD_SC_LS__EINVN_2%A
x_PM_SKY130_FD_SC_LS__EINVN_2%VPWR N_VPWR_M1006_s N_VPWR_M1000_s N_VPWR_c_245_n
+ N_VPWR_c_246_n N_VPWR_c_247_n VPWR N_VPWR_c_248_n N_VPWR_c_249_n
+ N_VPWR_c_244_n N_VPWR_c_251_n PM_SKY130_FD_SC_LS__EINVN_2%VPWR
x_PM_SKY130_FD_SC_LS__EINVN_2%A_227_368# N_A_227_368#_M1000_d
+ N_A_227_368#_M1007_d N_A_227_368#_M1005_s N_A_227_368#_c_283_n
+ N_A_227_368#_c_284_n N_A_227_368#_c_285_n N_A_227_368#_c_286_n
+ N_A_227_368#_c_304_n N_A_227_368#_c_287_n N_A_227_368#_c_288_n
+ N_A_227_368#_c_289_n PM_SKY130_FD_SC_LS__EINVN_2%A_227_368#
x_PM_SKY130_FD_SC_LS__EINVN_2%Z N_Z_M1002_s N_Z_M1003_d Z Z Z Z Z
+ PM_SKY130_FD_SC_LS__EINVN_2%Z
x_PM_SKY130_FD_SC_LS__EINVN_2%VGND N_VGND_M1009_s N_VGND_M1001_d N_VGND_c_360_n
+ N_VGND_c_361_n N_VGND_c_362_n VGND N_VGND_c_363_n N_VGND_c_364_n
+ N_VGND_c_365_n N_VGND_c_366_n PM_SKY130_FD_SC_LS__EINVN_2%VGND
x_PM_SKY130_FD_SC_LS__EINVN_2%A_231_74# N_A_231_74#_M1001_s N_A_231_74#_M1004_s
+ N_A_231_74#_M1008_d N_A_231_74#_c_397_n N_A_231_74#_c_398_n
+ N_A_231_74#_c_399_n N_A_231_74#_c_400_n N_A_231_74#_c_401_n
+ PM_SKY130_FD_SC_LS__EINVN_2%A_231_74#
cc_1 VNB N_A_115_464#_c_68_n 0.0175732f $X=-0.19 $Y=-0.245 $X2=1.44 $Y2=1.395
cc_2 VNB N_A_115_464#_M1001_g 0.0270981f $X=-0.19 $Y=-0.245 $X2=1.515 $Y2=0.74
cc_3 VNB N_A_115_464#_c_70_n 0.0227696f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=1.395
cc_4 VNB N_A_115_464#_M1004_g 0.021718f $X=-0.19 $Y=-0.245 $X2=1.945 $Y2=0.74
cc_5 VNB N_A_115_464#_c_72_n 0.0052192f $X=-0.19 $Y=-0.245 $X2=1.515 $Y2=1.395
cc_6 VNB N_A_115_464#_c_73_n 0.0111828f $X=-0.19 $Y=-0.245 $X2=0.805 $Y2=1.32
cc_7 VNB N_A_115_464#_c_74_n 0.0121801f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=0.58
cc_8 VNB N_A_115_464#_c_75_n 7.13956e-19 $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=2.3
cc_9 VNB N_A_115_464#_c_76_n 0.0095065f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.485
cc_10 VNB N_A_115_464#_c_77_n 0.0497031f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.395
cc_11 VNB N_TE_B_c_129_n 0.0305908f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=2.32
cc_12 VNB N_TE_B_M1009_g 0.0431726f $X=-0.19 $Y=-0.245 $X2=1.515 $Y2=1.32
cc_13 VNB N_TE_B_c_131_n 0.0227507f $X=-0.19 $Y=-0.245 $X2=0.805 $Y2=2.3
cc_14 VNB N_TE_B_c_132_n 0.0261838f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=0.58
cc_15 VNB N_A_c_194_n 0.0172813f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=0.37
cc_16 VNB N_A_c_195_n 0.0200758f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_c_196_n 0.0135987f $X=-0.19 $Y=-0.245 $X2=1.515 $Y2=1.32
cc_18 VNB N_A_c_197_n 0.020506f $X=-0.19 $Y=-0.245 $X2=1.515 $Y2=0.74
cc_19 VNB N_A_c_198_n 0.0678081f $X=-0.19 $Y=-0.245 $X2=1.59 $Y2=1.395
cc_20 VNB N_A_c_199_n 0.00694111f $X=-0.19 $Y=-0.245 $X2=1.945 $Y2=0.74
cc_21 VNB A 0.02299f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VPWR_c_244_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=0.58
cc_23 VNB Z 5.654e-19 $X=-0.19 $Y=-0.245 $X2=1.44 $Y2=1.395
cc_24 VNB Z 0.00184709f $X=-0.19 $Y=-0.245 $X2=1.16 $Y2=1.395
cc_25 VNB N_VGND_c_360_n 0.0111565f $X=-0.19 $Y=-0.245 $X2=1.44 $Y2=1.395
cc_26 VNB N_VGND_c_361_n 0.0310923f $X=-0.19 $Y=-0.245 $X2=1.515 $Y2=1.32
cc_27 VNB N_VGND_c_362_n 0.00396467f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=1.395
cc_28 VNB N_VGND_c_363_n 0.0329878f $X=-0.19 $Y=-0.245 $X2=1.945 $Y2=0.74
cc_29 VNB N_VGND_c_364_n 0.0398307f $X=-0.19 $Y=-0.245 $X2=0.805 $Y2=2.3
cc_30 VNB N_VGND_c_365_n 0.21764f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=0.58
cc_31 VNB N_VGND_c_366_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_231_74#_c_397_n 0.00810194f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_231_74#_c_398_n 0.00866729f $X=-0.19 $Y=-0.245 $X2=1.59 $Y2=1.395
cc_34 VNB N_A_231_74#_c_399_n 0.00413418f $X=-0.19 $Y=-0.245 $X2=1.945 $Y2=1.32
cc_35 VNB N_A_231_74#_c_400_n 0.0016059f $X=-0.19 $Y=-0.245 $X2=1.945 $Y2=0.74
cc_36 VNB N_A_231_74#_c_401_n 0.015961f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=2.465
cc_37 VPB N_A_115_464#_c_78_n 0.0138241f $X=-0.19 $Y=1.66 $X2=0.725 $Y2=2.465
cc_38 VPB N_A_115_464#_c_75_n 0.0139784f $X=-0.19 $Y=1.66 $X2=0.725 $Y2=2.3
cc_39 VPB N_TE_B_c_129_n 0.0262002f $X=-0.19 $Y=1.66 $X2=0.575 $Y2=2.32
cc_40 VPB N_TE_B_c_134_n 0.0333098f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_41 VPB N_TE_B_M1006_g 0.0117187f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_42 VPB N_TE_B_c_136_n 0.0626593f $X=-0.19 $Y=1.66 $X2=1.515 $Y2=0.74
cc_43 VPB N_TE_B_c_137_n 0.0135918f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_44 VPB N_TE_B_c_138_n 0.0162831f $X=-0.19 $Y=1.66 $X2=1.87 $Y2=1.395
cc_45 VPB N_TE_B_c_139_n 0.0297299f $X=-0.19 $Y=1.66 $X2=1.945 $Y2=0.74
cc_46 VPB N_TE_B_c_140_n 0.0132138f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB N_TE_B_c_141_n 0.00749069f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 VPB N_TE_B_c_132_n 0.0223278f $X=-0.19 $Y=1.66 $X2=0.725 $Y2=0.58
cc_49 VPB N_A_c_195_n 0.00111912f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_A_c_202_n 0.0214236f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_51 VPB N_A_c_198_n 0.0283056f $X=-0.19 $Y=1.66 $X2=1.59 $Y2=1.395
cc_52 VPB N_VPWR_c_245_n 0.0104926f $X=-0.19 $Y=1.66 $X2=1.44 $Y2=1.395
cc_53 VPB N_VPWR_c_246_n 0.0392161f $X=-0.19 $Y=1.66 $X2=1.515 $Y2=1.32
cc_54 VPB N_VPWR_c_247_n 0.00260181f $X=-0.19 $Y=1.66 $X2=1.87 $Y2=1.395
cc_55 VPB N_VPWR_c_248_n 0.0332027f $X=-0.19 $Y=1.66 $X2=1.945 $Y2=0.74
cc_56 VPB N_VPWR_c_249_n 0.0386269f $X=-0.19 $Y=1.66 $X2=0.805 $Y2=2.3
cc_57 VPB N_VPWR_c_244_n 0.053591f $X=-0.19 $Y=1.66 $X2=0.725 $Y2=0.58
cc_58 VPB N_VPWR_c_251_n 0.00345125f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_A_227_368#_c_283_n 0.00455758f $X=-0.19 $Y=1.66 $X2=1.515 $Y2=0.74
cc_60 VPB N_A_227_368#_c_284_n 0.0106744f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_A_227_368#_c_285_n 0.0036265f $X=-0.19 $Y=1.66 $X2=1.59 $Y2=1.395
cc_62 VPB N_A_227_368#_c_286_n 0.00593179f $X=-0.19 $Y=1.66 $X2=1.945 $Y2=0.74
cc_63 VPB N_A_227_368#_c_287_n 0.0121971f $X=-0.19 $Y=1.66 $X2=0.725 $Y2=2.465
cc_64 VPB N_A_227_368#_c_288_n 0.00181992f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_A_227_368#_c_289_n 0.0427462f $X=-0.19 $Y=1.66 $X2=0.805 $Y2=0.81
cc_66 VPB Z 0.00153198f $X=-0.19 $Y=1.66 $X2=1.16 $Y2=1.395
cc_67 VPB Z 2.84451e-19 $X=-0.19 $Y=1.66 $X2=1.515 $Y2=0.74
cc_68 N_A_115_464#_c_75_n N_TE_B_c_129_n 0.0155887f $X=0.725 $Y=2.3 $X2=0 $Y2=0
cc_69 N_A_115_464#_c_76_n N_TE_B_c_129_n 0.00223631f $X=0.995 $Y=1.485 $X2=0
+ $Y2=0
cc_70 N_A_115_464#_c_77_n N_TE_B_c_129_n 0.0170189f $X=0.995 $Y=1.395 $X2=0
+ $Y2=0
cc_71 N_A_115_464#_c_78_n N_TE_B_c_134_n 5.4497e-19 $X=0.725 $Y=2.465 $X2=0
+ $Y2=0
cc_72 N_A_115_464#_c_78_n N_TE_B_M1006_g 0.00896514f $X=0.725 $Y=2.465 $X2=0
+ $Y2=0
cc_73 N_A_115_464#_c_75_n N_TE_B_M1006_g 0.00189951f $X=0.725 $Y=2.3 $X2=0 $Y2=0
cc_74 N_A_115_464#_c_73_n N_TE_B_M1009_g 0.0157368f $X=0.805 $Y=1.32 $X2=0 $Y2=0
cc_75 N_A_115_464#_c_74_n N_TE_B_M1009_g 0.00786676f $X=0.725 $Y=0.58 $X2=0
+ $Y2=0
cc_76 N_A_115_464#_c_78_n N_TE_B_c_136_n 0.00558258f $X=0.725 $Y=2.465 $X2=0
+ $Y2=0
cc_77 N_A_115_464#_c_68_n N_TE_B_c_138_n 0.00943731f $X=1.44 $Y=1.395 $X2=0
+ $Y2=0
cc_78 N_A_115_464#_c_75_n N_TE_B_c_138_n 0.00285535f $X=0.725 $Y=2.3 $X2=0 $Y2=0
cc_79 N_A_115_464#_c_70_n N_TE_B_c_140_n 0.00889072f $X=1.87 $Y=1.395 $X2=0
+ $Y2=0
cc_80 N_A_115_464#_c_73_n N_TE_B_c_132_n 0.0152878f $X=0.805 $Y=1.32 $X2=0 $Y2=0
cc_81 N_A_115_464#_c_75_n N_TE_B_c_132_n 0.0367453f $X=0.725 $Y=2.3 $X2=0 $Y2=0
cc_82 N_A_115_464#_c_76_n N_TE_B_c_132_n 0.0271789f $X=0.995 $Y=1.485 $X2=0
+ $Y2=0
cc_83 N_A_115_464#_c_77_n N_TE_B_c_132_n 3.17368e-19 $X=0.995 $Y=1.395 $X2=0
+ $Y2=0
cc_84 N_A_115_464#_M1004_g N_A_c_194_n 0.0104506f $X=1.945 $Y=0.74 $X2=-0.19
+ $Y2=-0.245
cc_85 N_A_115_464#_c_70_n N_A_c_195_n 0.00490479f $X=1.87 $Y=1.395 $X2=0 $Y2=0
cc_86 N_A_115_464#_c_70_n N_A_c_199_n 0.0104506f $X=1.87 $Y=1.395 $X2=0 $Y2=0
cc_87 N_A_115_464#_c_78_n N_VPWR_c_246_n 0.0456209f $X=0.725 $Y=2.465 $X2=0
+ $Y2=0
cc_88 N_A_115_464#_c_78_n N_VPWR_c_248_n 0.0145841f $X=0.725 $Y=2.465 $X2=0
+ $Y2=0
cc_89 N_A_115_464#_c_78_n N_VPWR_c_244_n 0.0107612f $X=0.725 $Y=2.465 $X2=0
+ $Y2=0
cc_90 N_A_115_464#_c_68_n N_A_227_368#_c_283_n 0.00507112f $X=1.44 $Y=1.395
+ $X2=0 $Y2=0
cc_91 N_A_115_464#_c_75_n N_A_227_368#_c_283_n 0.0117904f $X=0.725 $Y=2.3 $X2=0
+ $Y2=0
cc_92 N_A_115_464#_c_76_n N_A_227_368#_c_283_n 0.003795f $X=0.995 $Y=1.485 $X2=0
+ $Y2=0
cc_93 N_A_115_464#_c_77_n N_A_227_368#_c_283_n 0.0010483f $X=0.995 $Y=1.395
+ $X2=0 $Y2=0
cc_94 N_A_115_464#_c_75_n N_A_227_368#_c_284_n 0.0659097f $X=0.725 $Y=2.3 $X2=0
+ $Y2=0
cc_95 N_A_115_464#_c_68_n N_A_227_368#_c_285_n 0.00116956f $X=1.44 $Y=1.395
+ $X2=0 $Y2=0
cc_96 N_A_115_464#_c_70_n N_A_227_368#_c_285_n 5.4934e-19 $X=1.87 $Y=1.395 $X2=0
+ $Y2=0
cc_97 N_A_115_464#_c_72_n N_A_227_368#_c_285_n 0.00690164f $X=1.515 $Y=1.395
+ $X2=0 $Y2=0
cc_98 N_A_115_464#_M1004_g Z 0.00127446f $X=1.945 $Y=0.74 $X2=0 $Y2=0
cc_99 N_A_115_464#_c_74_n N_VGND_c_361_n 0.0179429f $X=0.725 $Y=0.58 $X2=0 $Y2=0
cc_100 N_A_115_464#_M1001_g N_VGND_c_362_n 0.012411f $X=1.515 $Y=0.74 $X2=0
+ $Y2=0
cc_101 N_A_115_464#_M1004_g N_VGND_c_362_n 0.00950277f $X=1.945 $Y=0.74 $X2=0
+ $Y2=0
cc_102 N_A_115_464#_M1001_g N_VGND_c_363_n 0.00383152f $X=1.515 $Y=0.74 $X2=0
+ $Y2=0
cc_103 N_A_115_464#_c_74_n N_VGND_c_363_n 0.0143708f $X=0.725 $Y=0.58 $X2=0
+ $Y2=0
cc_104 N_A_115_464#_M1004_g N_VGND_c_364_n 0.00383152f $X=1.945 $Y=0.74 $X2=0
+ $Y2=0
cc_105 N_A_115_464#_M1001_g N_VGND_c_365_n 0.00762539f $X=1.515 $Y=0.74 $X2=0
+ $Y2=0
cc_106 N_A_115_464#_M1004_g N_VGND_c_365_n 0.00757637f $X=1.945 $Y=0.74 $X2=0
+ $Y2=0
cc_107 N_A_115_464#_c_74_n N_VGND_c_365_n 0.011923f $X=0.725 $Y=0.58 $X2=0 $Y2=0
cc_108 N_A_115_464#_M1001_g N_A_231_74#_c_397_n 0.00159319f $X=1.515 $Y=0.74
+ $X2=0 $Y2=0
cc_109 N_A_115_464#_c_74_n N_A_231_74#_c_397_n 0.039239f $X=0.725 $Y=0.58 $X2=0
+ $Y2=0
cc_110 N_A_115_464#_c_68_n N_A_231_74#_c_398_n 0.00129671f $X=1.44 $Y=1.395
+ $X2=0 $Y2=0
cc_111 N_A_115_464#_M1001_g N_A_231_74#_c_398_n 0.0142221f $X=1.515 $Y=0.74
+ $X2=0 $Y2=0
cc_112 N_A_115_464#_c_70_n N_A_231_74#_c_398_n 0.00240153f $X=1.87 $Y=1.395
+ $X2=0 $Y2=0
cc_113 N_A_115_464#_M1004_g N_A_231_74#_c_398_n 0.0138457f $X=1.945 $Y=0.74
+ $X2=0 $Y2=0
cc_114 N_A_115_464#_c_73_n N_A_231_74#_c_399_n 0.0111139f $X=0.805 $Y=1.32 $X2=0
+ $Y2=0
cc_115 N_A_115_464#_c_76_n N_A_231_74#_c_399_n 0.00210833f $X=0.995 $Y=1.485
+ $X2=0 $Y2=0
cc_116 N_A_115_464#_c_77_n N_A_231_74#_c_399_n 0.00660264f $X=0.995 $Y=1.395
+ $X2=0 $Y2=0
cc_117 N_TE_B_c_139_n N_A_c_202_n 0.00255103f $X=1.88 $Y=3.11 $X2=0 $Y2=0
cc_118 N_TE_B_c_140_n N_A_c_202_n 0.0104511f $X=1.955 $Y=3.035 $X2=0 $Y2=0
cc_119 N_TE_B_c_134_n N_VPWR_c_246_n 0.00108702f $X=0.5 $Y=2.245 $X2=0 $Y2=0
cc_120 N_TE_B_M1006_g N_VPWR_c_246_n 0.0052938f $X=0.5 $Y=2.64 $X2=0 $Y2=0
cc_121 N_TE_B_c_137_n N_VPWR_c_246_n 0.00624174f $X=0.575 $Y=3.11 $X2=0 $Y2=0
cc_122 N_TE_B_c_132_n N_VPWR_c_246_n 0.0212001f $X=0.385 $Y=1.285 $X2=0 $Y2=0
cc_123 N_TE_B_c_138_n N_VPWR_c_247_n 0.00217316f $X=1.505 $Y=3.035 $X2=0 $Y2=0
cc_124 N_TE_B_c_139_n N_VPWR_c_247_n 0.0181091f $X=1.88 $Y=3.11 $X2=0 $Y2=0
cc_125 N_TE_B_c_140_n N_VPWR_c_247_n 0.00373405f $X=1.955 $Y=3.035 $X2=0 $Y2=0
cc_126 N_TE_B_c_137_n N_VPWR_c_248_n 0.0320947f $X=0.575 $Y=3.11 $X2=0 $Y2=0
cc_127 N_TE_B_c_139_n N_VPWR_c_249_n 0.00784922f $X=1.88 $Y=3.11 $X2=0 $Y2=0
cc_128 N_TE_B_c_136_n N_VPWR_c_244_n 0.0288728f $X=1.43 $Y=3.11 $X2=0 $Y2=0
cc_129 N_TE_B_c_137_n N_VPWR_c_244_n 0.0108306f $X=0.575 $Y=3.11 $X2=0 $Y2=0
cc_130 N_TE_B_c_139_n N_VPWR_c_244_n 0.0144853f $X=1.88 $Y=3.11 $X2=0 $Y2=0
cc_131 N_TE_B_c_141_n N_VPWR_c_244_n 0.00904465f $X=1.505 $Y=3.11 $X2=0 $Y2=0
cc_132 N_TE_B_M1006_g N_A_227_368#_c_284_n 0.00119572f $X=0.5 $Y=2.64 $X2=0
+ $Y2=0
cc_133 N_TE_B_c_136_n N_A_227_368#_c_284_n 0.00558669f $X=1.43 $Y=3.11 $X2=0
+ $Y2=0
cc_134 N_TE_B_c_138_n N_A_227_368#_c_284_n 0.0014444f $X=1.505 $Y=3.035 $X2=0
+ $Y2=0
cc_135 N_TE_B_c_138_n N_A_227_368#_c_285_n 0.0138982f $X=1.505 $Y=3.035 $X2=0
+ $Y2=0
cc_136 N_TE_B_c_140_n N_A_227_368#_c_285_n 0.0124129f $X=1.955 $Y=3.035 $X2=0
+ $Y2=0
cc_137 N_TE_B_c_140_n N_A_227_368#_c_286_n 7.02482e-19 $X=1.955 $Y=3.035 $X2=0
+ $Y2=0
cc_138 N_TE_B_c_138_n N_A_227_368#_c_304_n 6.71925e-19 $X=1.505 $Y=3.035 $X2=0
+ $Y2=0
cc_139 N_TE_B_c_140_n N_A_227_368#_c_304_n 0.0111451f $X=1.955 $Y=3.035 $X2=0
+ $Y2=0
cc_140 N_TE_B_c_139_n N_A_227_368#_c_288_n 0.00181967f $X=1.88 $Y=3.11 $X2=0
+ $Y2=0
cc_141 N_TE_B_c_140_n N_A_227_368#_c_288_n 0.0022238f $X=1.955 $Y=3.035 $X2=0
+ $Y2=0
cc_142 N_TE_B_c_140_n Z 5.12494e-19 $X=1.955 $Y=3.035 $X2=0 $Y2=0
cc_143 N_TE_B_c_140_n Z 2.69789e-19 $X=1.955 $Y=3.035 $X2=0 $Y2=0
cc_144 N_TE_B_M1009_g N_VGND_c_361_n 0.00589946f $X=0.51 $Y=0.58 $X2=0 $Y2=0
cc_145 N_TE_B_c_131_n N_VGND_c_361_n 0.00115809f $X=0.385 $Y=1.285 $X2=0 $Y2=0
cc_146 N_TE_B_c_132_n N_VGND_c_361_n 0.0145115f $X=0.385 $Y=1.285 $X2=0 $Y2=0
cc_147 N_TE_B_M1009_g N_VGND_c_363_n 0.00434272f $X=0.51 $Y=0.58 $X2=0 $Y2=0
cc_148 N_TE_B_M1009_g N_VGND_c_365_n 0.00828991f $X=0.51 $Y=0.58 $X2=0 $Y2=0
cc_149 N_TE_B_M1009_g N_A_231_74#_c_397_n 9.23906e-19 $X=0.51 $Y=0.58 $X2=0
+ $Y2=0
cc_150 N_TE_B_c_138_n N_A_231_74#_c_398_n 3.80991e-19 $X=1.505 $Y=3.035 $X2=0
+ $Y2=0
cc_151 N_TE_B_c_140_n N_A_231_74#_c_398_n 5.78606e-19 $X=1.955 $Y=3.035 $X2=0
+ $Y2=0
cc_152 N_A_c_202_n N_VPWR_c_249_n 0.00278271f $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_153 N_A_c_198_n N_VPWR_c_249_n 0.00278271f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_154 N_A_c_202_n N_VPWR_c_244_n 0.0035377f $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_155 N_A_c_198_n N_VPWR_c_244_n 0.00357317f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_156 N_A_c_202_n N_A_227_368#_c_287_n 0.0127806f $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_157 N_A_c_198_n N_A_227_368#_c_287_n 0.0137046f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_158 N_A_c_198_n N_A_227_368#_c_289_n 0.00351248f $X=2.855 $Y=1.765 $X2=0
+ $Y2=0
cc_159 A N_A_227_368#_c_289_n 0.0175067f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_160 N_A_c_194_n Z 0.00549559f $X=2.375 $Y=1.22 $X2=0 $Y2=0
cc_161 N_A_c_197_n Z 0.00558139f $X=2.81 $Y=1.22 $X2=0 $Y2=0
cc_162 A Z 0.0443015f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_163 N_A_c_194_n Z 0.00212163f $X=2.375 $Y=1.22 $X2=0 $Y2=0
cc_164 N_A_c_195_n Z 0.0138409f $X=2.405 $Y=1.675 $X2=0 $Y2=0
cc_165 N_A_c_202_n Z 0.00529818f $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_166 N_A_c_196_n Z 0.0115492f $X=2.735 $Y=1.295 $X2=0 $Y2=0
cc_167 N_A_c_197_n Z 0.00179582f $X=2.81 $Y=1.22 $X2=0 $Y2=0
cc_168 N_A_c_198_n Z 0.0150869f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_169 N_A_c_199_n Z 0.00290588f $X=2.397 $Y=1.295 $X2=0 $Y2=0
cc_170 N_A_c_202_n Z 0.00179807f $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_171 N_A_c_198_n Z 0.00387064f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_172 N_A_c_202_n Z 0.00723184f $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_173 N_A_c_198_n Z 0.00764814f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_174 N_A_c_194_n N_VGND_c_362_n 6.35276e-19 $X=2.375 $Y=1.22 $X2=0 $Y2=0
cc_175 N_A_c_194_n N_VGND_c_364_n 0.00291649f $X=2.375 $Y=1.22 $X2=0 $Y2=0
cc_176 N_A_c_197_n N_VGND_c_364_n 0.00291649f $X=2.81 $Y=1.22 $X2=0 $Y2=0
cc_177 N_A_c_194_n N_VGND_c_365_n 0.00359269f $X=2.375 $Y=1.22 $X2=0 $Y2=0
cc_178 N_A_c_197_n N_VGND_c_365_n 0.00363003f $X=2.81 $Y=1.22 $X2=0 $Y2=0
cc_179 A N_VGND_c_365_n 0.00283239f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_180 A N_A_231_74#_M1008_d 0.00476174f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_181 N_A_c_194_n N_A_231_74#_c_398_n 3.43633e-19 $X=2.375 $Y=1.22 $X2=0 $Y2=0
cc_182 N_A_c_194_n N_A_231_74#_c_401_n 0.0142515f $X=2.375 $Y=1.22 $X2=0 $Y2=0
cc_183 N_A_c_196_n N_A_231_74#_c_401_n 3.11327e-19 $X=2.735 $Y=1.295 $X2=0 $Y2=0
cc_184 N_A_c_197_n N_A_231_74#_c_401_n 0.0145459f $X=2.81 $Y=1.22 $X2=0 $Y2=0
cc_185 N_A_c_198_n N_A_231_74#_c_401_n 8.45143e-19 $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_186 A N_A_231_74#_c_401_n 0.017603f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_187 N_VPWR_c_247_n N_A_227_368#_c_284_n 0.0280319f $X=1.73 $Y=2.325 $X2=0
+ $Y2=0
cc_188 N_VPWR_c_248_n N_A_227_368#_c_284_n 0.012618f $X=1.58 $Y=3.33 $X2=0 $Y2=0
cc_189 N_VPWR_c_244_n N_A_227_368#_c_284_n 0.00931741f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_190 N_VPWR_M1000_s N_A_227_368#_c_285_n 0.00222494f $X=1.58 $Y=1.84 $X2=0
+ $Y2=0
cc_191 N_VPWR_c_247_n N_A_227_368#_c_285_n 0.0144005f $X=1.73 $Y=2.325 $X2=0
+ $Y2=0
cc_192 N_VPWR_c_247_n N_A_227_368#_c_304_n 0.0490769f $X=1.73 $Y=2.325 $X2=0
+ $Y2=0
cc_193 N_VPWR_c_249_n N_A_227_368#_c_287_n 0.062301f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_194 N_VPWR_c_244_n N_A_227_368#_c_287_n 0.0347031f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_195 N_VPWR_c_247_n N_A_227_368#_c_288_n 0.0120205f $X=1.73 $Y=2.325 $X2=0
+ $Y2=0
cc_196 N_VPWR_c_249_n N_A_227_368#_c_288_n 0.0199669f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_197 N_VPWR_c_244_n N_A_227_368#_c_288_n 0.0107485f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_198 N_A_227_368#_c_287_n N_Z_M1003_d 0.00197722f $X=2.965 $Y=2.99 $X2=0 $Y2=0
cc_199 N_A_227_368#_c_286_n Z 0.00725716f $X=2.155 $Y=1.99 $X2=0 $Y2=0
cc_200 N_A_227_368#_c_289_n Z 0.0350665f $X=3.08 $Y=1.985 $X2=0 $Y2=0
cc_201 N_A_227_368#_c_287_n Z 0.0160777f $X=2.965 $Y=2.99 $X2=0 $Y2=0
cc_202 N_A_227_368#_c_283_n N_A_231_74#_c_398_n 4.64785e-19 $X=1.257 $Y=1.99
+ $X2=0 $Y2=0
cc_203 N_A_227_368#_c_285_n N_A_231_74#_c_398_n 0.0155334f $X=2.015 $Y=1.905
+ $X2=0 $Y2=0
cc_204 N_A_227_368#_c_286_n N_A_231_74#_c_398_n 0.00791107f $X=2.155 $Y=1.99
+ $X2=0 $Y2=0
cc_205 N_A_227_368#_c_283_n N_A_231_74#_c_399_n 0.0079427f $X=1.257 $Y=1.99
+ $X2=0 $Y2=0
cc_206 Z N_A_231_74#_c_398_n 0.00625076f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_207 Z N_A_231_74#_c_398_n 0.00142622f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_208 N_Z_M1002_s N_A_231_74#_c_401_n 0.00174803f $X=2.45 $Y=0.37 $X2=0 $Y2=0
cc_209 Z N_A_231_74#_c_401_n 0.0168802f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_210 N_VGND_c_362_n N_A_231_74#_c_397_n 0.0164982f $X=1.73 $Y=0.61 $X2=0 $Y2=0
cc_211 N_VGND_c_363_n N_A_231_74#_c_397_n 0.011066f $X=1.565 $Y=0 $X2=0 $Y2=0
cc_212 N_VGND_c_365_n N_A_231_74#_c_397_n 0.00915947f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_213 N_VGND_M1001_d N_A_231_74#_c_398_n 0.00184993f $X=1.59 $Y=0.37 $X2=0
+ $Y2=0
cc_214 N_VGND_c_362_n N_A_231_74#_c_398_n 0.0156953f $X=1.73 $Y=0.61 $X2=0 $Y2=0
cc_215 N_VGND_c_362_n N_A_231_74#_c_400_n 0.00985092f $X=1.73 $Y=0.61 $X2=0
+ $Y2=0
cc_216 N_VGND_c_364_n N_A_231_74#_c_400_n 0.00758556f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_217 N_VGND_c_365_n N_A_231_74#_c_400_n 0.00627867f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_218 N_VGND_c_364_n N_A_231_74#_c_401_n 0.038742f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_219 N_VGND_c_365_n N_A_231_74#_c_401_n 0.0327013f $X=3.12 $Y=0 $X2=0 $Y2=0
