* NGSPICE file created from sky130_fd_sc_ls__o2bb2ai_4.ext - technology: sky130A

.subckt sky130_fd_sc_ls__o2bb2ai_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
M1000 a_114_368# A1_N VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=1.344e+12p pd=1.136e+07u as=2.9904e+12p ps=2.55e+07u
M1001 Y B2 a_1215_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=1.344e+12p pd=1.136e+07u as=1.6464e+12p ps=1.414e+07u
M1002 a_857_74# B1 VGND VNB nshort w=740000u l=150000u
+  ad=1.4578e+12p pd=1.43e+07u as=1.3986e+12p ps=1.266e+07u
M1003 a_27_74# A2_N a_114_368# VNB nshort w=740000u l=150000u
+  ad=1.1211e+12p pd=1.043e+07u as=4.477e+11p ps=4.17e+06u
M1004 a_857_74# a_114_368# Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=4.144e+11p ps=4.08e+06u
M1005 VPWR A2_N a_114_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR a_114_368# Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_27_74# A1_N VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND B1 a_857_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_1215_368# B1 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR A1_N a_114_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND B1 a_857_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_114_368# A2_N a_27_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_1215_368# B2 Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Y a_114_368# a_857_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y a_114_368# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Y a_114_368# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR B1 a_1215_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_114_368# A2_N VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR a_114_368# Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 Y B2 a_1215_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_114_368# A2_N a_27_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_857_74# a_114_368# Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_857_74# B2 VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_1215_368# B1 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPWR A2_N a_114_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VGND B2 a_857_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_1215_368# B2 Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 Y a_114_368# a_857_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_114_368# A1_N VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VPWR A1_N a_114_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VGND A1_N a_27_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_27_74# A1_N VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VGND A1_N a_27_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_857_74# B1 VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_857_74# B2 VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_114_368# A2_N VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_27_74# A2_N a_114_368# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 VPWR B1 a_1215_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 VGND B2 a_857_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

