# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_ls__sdfrtp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  13.44000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 0.810000 2.100000 1.265000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.995000 0.350000 13.325000 1.130000 ;
        RECT 13.070000 1.130000 13.325000 2.980000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.411000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT  3.935000 1.920000  4.225000 1.965000 ;
        RECT  3.935000 1.965000 10.945000 2.105000 ;
        RECT  3.935000 2.105000  4.225000 2.150000 ;
        RECT  7.775000 1.920000  8.065000 1.965000 ;
        RECT  7.775000 2.105000  8.065000 2.150000 ;
        RECT 10.655000 1.920000 10.945000 1.965000 ;
        RECT 10.655000 2.105000 10.945000 2.150000 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.945000 1.440000 3.275000 2.150000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.455000 1.490000 2.725000 1.660000 ;
        RECT 0.455000 1.660000 1.795000 1.835000 ;
        RECT 2.345000 1.260000 2.725000 1.490000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.785000 0.920000 4.195000 1.260000 ;
        RECT 3.785000 1.260000 4.640000 1.650000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 13.440000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 13.440000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 13.440000 0.085000 ;
      RECT  0.000000  3.245000 13.440000 3.415000 ;
      RECT  0.115000  0.420000  0.365000 1.050000 ;
      RECT  0.115000  1.050000  1.375000 1.265000 ;
      RECT  0.115000  1.265000  0.285000 2.005000 ;
      RECT  0.115000  2.005000  2.705000 2.175000 ;
      RECT  0.115000  2.175000  0.445000 2.980000 ;
      RECT  0.545000  0.085000  0.875000 0.880000 ;
      RECT  0.615000  2.345000  0.945000 3.245000 ;
      RECT  1.045000  0.935000  1.375000 1.050000 ;
      RECT  1.105000  0.255000  3.410000 0.425000 ;
      RECT  1.105000  0.425000  1.435000 0.640000 ;
      RECT  1.485000  2.345000  3.785000 2.385000 ;
      RECT  1.485000  2.385000  4.230000 2.400000 ;
      RECT  1.485000  2.400000  4.250000 2.420000 ;
      RECT  1.485000  2.420000  6.075000 2.515000 ;
      RECT  1.485000  2.515000  2.555000 2.980000 ;
      RECT  2.035000  1.830000  2.705000 2.005000 ;
      RECT  2.270000  0.595000  2.600000 0.920000 ;
      RECT  2.270000  0.920000  3.615000 1.090000 ;
      RECT  3.060000  0.425000  3.410000 0.750000 ;
      RECT  3.095000  2.685000  3.425000 3.245000 ;
      RECT  3.445000  1.090000  3.615000 2.330000 ;
      RECT  3.445000  2.330000  3.785000 2.345000 ;
      RECT  3.590000  0.085000  3.880000 0.750000 ;
      RECT  3.665000  2.515000  6.075000 2.580000 ;
      RECT  3.665000  2.580000  4.645000 2.585000 ;
      RECT  3.665000  2.585000  4.630000 2.590000 ;
      RECT  3.665000  2.590000  4.610000 2.600000 ;
      RECT  3.665000  2.600000  4.580000 2.620000 ;
      RECT  3.665000  2.620000  3.995000 2.980000 ;
      RECT  3.785000  1.830000  4.165000 2.160000 ;
      RECT  3.920000  2.160000  4.165000 2.190000 ;
      RECT  4.135000  0.500000  4.535000 0.750000 ;
      RECT  4.335000  1.820000  4.980000 2.195000 ;
      RECT  4.335000  2.195000  4.505000 2.250000 ;
      RECT  4.365000  0.750000  4.535000 0.920000 ;
      RECT  4.365000  0.920000  5.045000 1.090000 ;
      RECT  4.555000  2.415000  6.075000 2.420000 ;
      RECT  4.570000  2.410000  6.075000 2.415000 ;
      RECT  4.590000  2.400000  6.075000 2.410000 ;
      RECT  4.615000  2.385000  6.075000 2.400000 ;
      RECT  4.705000  0.085000  5.035000 0.750000 ;
      RECT  4.705000  2.750000  5.035000 3.245000 ;
      RECT  4.810000  1.090000  5.045000 1.455000 ;
      RECT  4.810000  1.455000  5.280000 1.775000 ;
      RECT  4.810000  1.775000  4.980000 1.820000 ;
      RECT  5.155000  1.955000  5.630000 2.215000 ;
      RECT  5.215000  0.255000  7.220000 0.425000 ;
      RECT  5.215000  0.425000  5.620000 1.070000 ;
      RECT  5.215000  1.070000  5.630000 1.285000 ;
      RECT  5.450000  1.285000  5.630000 1.545000 ;
      RECT  5.450000  1.545000  6.200000 1.875000 ;
      RECT  5.450000  1.875000  5.630000 1.955000 ;
      RECT  5.795000  0.595000  5.975000 0.995000 ;
      RECT  5.800000  0.995000  5.975000 1.200000 ;
      RECT  5.800000  1.200000  6.540000 1.370000 ;
      RECT  5.825000  2.045000  6.540000 2.215000 ;
      RECT  5.825000  2.215000  6.075000 2.385000 ;
      RECT  5.825000  2.580000  6.075000 2.725000 ;
      RECT  6.145000  0.595000  6.470000 0.860000 ;
      RECT  6.145000  0.860000  6.880000 1.030000 ;
      RECT  6.250000  2.385000  8.075000 2.490000 ;
      RECT  6.250000  2.490000  6.880000 2.725000 ;
      RECT  6.370000  1.370000  6.540000 2.045000 ;
      RECT  6.710000  1.030000  6.880000 2.320000 ;
      RECT  6.710000  2.320000  8.075000 2.385000 ;
      RECT  7.050000  0.425000  7.220000 0.580000 ;
      RECT  7.050000  0.580000  8.100000 0.750000 ;
      RECT  7.050000  0.920000  8.895000 1.090000 ;
      RECT  7.050000  1.090000  7.325000 1.805000 ;
      RECT  7.205000  2.660000  7.540000 3.245000 ;
      RECT  7.430000  0.085000  7.760000 0.410000 ;
      RECT  7.495000  1.260000  8.315000 1.575000 ;
      RECT  7.495000  1.575000  7.665000 2.320000 ;
      RECT  7.745000  2.490000  8.075000 2.745000 ;
      RECT  7.835000  1.815000  8.165000 2.150000 ;
      RECT  7.930000  0.255000  9.235000 0.425000 ;
      RECT  7.930000  0.425000  8.100000 0.580000 ;
      RECT  8.270000  0.595000  8.655000 0.920000 ;
      RECT  8.385000  1.745000  8.555000 3.245000 ;
      RECT  8.725000  1.090000  8.895000 1.715000 ;
      RECT  8.725000  1.715000  9.005000 2.755000 ;
      RECT  9.065000  0.425000  9.235000 0.940000 ;
      RECT  9.065000  0.940000  9.415000 1.270000 ;
      RECT  9.245000  1.270000  9.415000 2.125000 ;
      RECT  9.245000  2.125000  9.975000 2.380000 ;
      RECT  9.290000  2.550000 10.315000 2.880000 ;
      RECT  9.405000  0.350000  9.755000 0.770000 ;
      RECT  9.585000  0.770000  9.755000 1.095000 ;
      RECT  9.585000  1.095000 11.395000 1.265000 ;
      RECT  9.585000  1.265000  9.755000 1.785000 ;
      RECT  9.585000  1.785000 10.315000 1.955000 ;
      RECT  9.985000  1.435000 10.315000 1.445000 ;
      RECT  9.985000  1.445000 11.735000 1.615000 ;
      RECT 10.145000  1.955000 10.315000 2.550000 ;
      RECT 10.195000  0.085000 10.525000 0.810000 ;
      RECT 10.485000  2.520000 10.735000 3.245000 ;
      RECT 10.640000  1.820000 10.970000 2.150000 ;
      RECT 10.945000  2.520000 11.310000 2.980000 ;
      RECT 11.010000  0.350000 11.340000 0.755000 ;
      RECT 11.010000  0.755000 11.735000 0.925000 ;
      RECT 11.065000  1.265000 11.395000 1.275000 ;
      RECT 11.140000  1.615000 11.310000 2.520000 ;
      RECT 11.480000  2.100000 11.810000 3.245000 ;
      RECT 11.565000  0.925000 11.735000 1.445000 ;
      RECT 11.570000  0.085000 11.905000 0.585000 ;
      RECT 11.980000  2.100000 12.310000 2.980000 ;
      RECT 12.085000  0.350000 12.335000 1.300000 ;
      RECT 12.085000  1.300000 12.870000 1.630000 ;
      RECT 12.085000  1.630000 12.310000 2.100000 ;
      RECT 12.540000  1.820000 12.870000 3.245000 ;
      RECT 12.565000  0.085000 12.815000 1.130000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  1.950000  4.165000 2.120000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  1.950000  8.005000 2.120000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  1.950000 10.885000 2.120000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.245000 13.285000 3.415000 ;
  END
END sky130_fd_sc_ls__sdfrtp_1
END LIBRARY
