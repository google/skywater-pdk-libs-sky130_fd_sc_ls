* File: sky130_fd_sc_ls__a311oi_1.pex.spice
* Created: Fri Aug 28 12:57:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__A311OI_1%A3 1 3 6 8 9 10 11
c27 1 0 4.6169e-20 $X=0.705 $Y=1.765
r28 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.33
+ $Y=1.385 $X2=0.33 $Y2=1.385
r29 11 16 8.72119 $w=3.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.31 $Y=1.665
+ $X2=0.31 $Y2=1.385
r30 10 16 2.80324 $w=3.68e-07 $l=9e-08 $layer=LI1_cond $X=0.31 $Y=1.295 $X2=0.31
+ $Y2=1.385
r31 8 15 49.8355 $w=3.3e-07 $l=2.85e-07 $layer=POLY_cond $X=0.615 $Y=1.385
+ $X2=0.33 $Y2=1.385
r32 8 9 66.2869 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.705 $Y=1.385
+ $X2=0.705 $Y2=1.22
r33 6 9 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.72 $Y=0.74 $X2=0.72
+ $Y2=1.22
r34 1 8 149.859 $w=1.8e-07 $l=3.8e-07 $layer=POLY_cond $X=0.705 $Y=1.765
+ $X2=0.705 $Y2=1.385
r35 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.705 $Y=1.765
+ $X2=0.705 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__A311OI_1%A2 3 5 7 8 12
c32 12 0 4.6169e-20 $X=1.17 $Y=1.515
r33 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.17
+ $Y=1.515 $X2=1.17 $Y2=1.515
r34 8 12 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.17 $Y=1.665
+ $X2=1.17 $Y2=1.515
r35 5 11 52.2586 $w=2.99e-07 $l=2.57391e-07 $layer=POLY_cond $X=1.155 $Y=1.765
+ $X2=1.17 $Y2=1.515
r36 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.155 $Y=1.765
+ $X2=1.155 $Y2=2.4
r37 1 11 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=1.08 $Y=1.35
+ $X2=1.17 $Y2=1.515
r38 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.08 $Y=1.35 $X2=1.08
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__A311OI_1%A1 3 5 7 8 12
r29 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.71
+ $Y=1.515 $X2=1.71 $Y2=1.515
r30 8 12 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.71 $Y=1.665
+ $X2=1.71 $Y2=1.515
r31 5 11 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=1.785 $Y=1.765
+ $X2=1.71 $Y2=1.515
r32 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.785 $Y=1.765
+ $X2=1.785 $Y2=2.4
r33 1 11 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=1.62 $Y=1.35
+ $X2=1.71 $Y2=1.515
r34 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.62 $Y=1.35 $X2=1.62
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__A311OI_1%B1 3 5 7 8 9
c30 5 0 1.56668e-19 $X=2.235 $Y=1.765
r31 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.25
+ $Y=1.515 $X2=2.25 $Y2=1.515
r32 9 14 10.4524 $w=4.28e-07 $l=3.9e-07 $layer=LI1_cond $X=2.64 $Y=1.565
+ $X2=2.25 $Y2=1.565
r33 8 14 2.41209 $w=4.28e-07 $l=9e-08 $layer=LI1_cond $X=2.16 $Y=1.565 $X2=2.25
+ $Y2=1.565
r34 5 13 52.2586 $w=2.99e-07 $l=2.57391e-07 $layer=POLY_cond $X=2.235 $Y=1.765
+ $X2=2.25 $Y2=1.515
r35 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.235 $Y=1.765
+ $X2=2.235 $Y2=2.4
r36 1 13 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=2.16 $Y=1.35
+ $X2=2.25 $Y2=1.515
r37 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.16 $Y=1.35 $X2=2.16
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__A311OI_1%C1 3 5 7 9 10 13 14
c30 14 0 1.56668e-19 $X=3.09 $Y=1.515
r31 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.09
+ $Y=1.515 $X2=3.09 $Y2=1.515
r32 10 14 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=3.09 $Y=1.665
+ $X2=3.09 $Y2=1.515
r33 8 13 49.8355 $w=3.3e-07 $l=2.85e-07 $layer=POLY_cond $X=2.805 $Y=1.515
+ $X2=3.09 $Y2=1.515
r34 8 9 5.03009 $w=3.3e-07 $l=1.08995e-07 $layer=POLY_cond $X=2.805 $Y=1.515
+ $X2=2.715 $Y2=1.557
r35 5 9 37.0704 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.715 $Y=1.765
+ $X2=2.715 $Y2=1.557
r36 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.715 $Y=1.765
+ $X2=2.715 $Y2=2.4
r37 1 9 37.0704 $w=1.5e-07 $l=2.14369e-07 $layer=POLY_cond $X=2.7 $Y=1.35
+ $X2=2.715 $Y2=1.557
r38 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.7 $Y=1.35 $X2=2.7
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__A311OI_1%VPWR 1 2 9 13 16 17 19 20 21 34 35
r35 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r36 31 34 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.68 $Y=3.33
+ $X2=3.12 $Y2=3.33
r37 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r38 25 29 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r39 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r40 21 35 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=3.12 $Y2=3.33
r41 21 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r42 21 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r43 19 28 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=1.265 $Y=3.33
+ $X2=1.2 $Y2=3.33
r44 19 20 9.97069 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=1.265 $Y=3.33
+ $X2=1.47 $Y2=3.33
r45 18 31 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=1.675 $Y=3.33
+ $X2=1.68 $Y2=3.33
r46 18 20 9.97069 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=1.675 $Y=3.33
+ $X2=1.47 $Y2=3.33
r47 16 24 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=0.315 $Y=3.33
+ $X2=0.24 $Y2=3.33
r48 16 17 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.315 $Y=3.33
+ $X2=0.44 $Y2=3.33
r49 15 28 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=1.2 $Y2=3.33
r50 15 17 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.44 $Y2=3.33
r51 11 20 1.53834 $w=4.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.47 $Y=3.245
+ $X2=1.47 $Y2=3.33
r52 11 13 13.6326 $w=4.08e-07 $l=4.85e-07 $layer=LI1_cond $X=1.47 $Y=3.245
+ $X2=1.47 $Y2=2.76
r53 7 17 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.44 $Y=3.245
+ $X2=0.44 $Y2=3.33
r54 7 9 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=0.44 $Y=3.245 $X2=0.44
+ $Y2=2.455
r55 2 13 600 $w=1.7e-07 $l=1.03305e-06 $layer=licon1_PDIFF $count=1 $X=1.23
+ $Y=1.84 $X2=1.47 $Y2=2.76
r56 1 9 300 $w=1.7e-07 $l=6.74611e-07 $layer=licon1_PDIFF $count=2 $X=0.355
+ $Y=1.84 $X2=0.48 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_LS__A311OI_1%A_156_368# 1 2 9 14 16
r27 10 14 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.095 $Y=2.375
+ $X2=0.93 $Y2=2.375
r28 9 16 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.845 $Y=2.375
+ $X2=2.01 $Y2=2.375
r29 9 10 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=1.845 $Y=2.375
+ $X2=1.095 $Y2=2.375
r30 2 16 300 $w=1.7e-07 $l=6.40625e-07 $layer=licon1_PDIFF $count=2 $X=1.86
+ $Y=1.84 $X2=2.01 $Y2=2.41
r31 1 14 300 $w=1.7e-07 $l=6.40625e-07 $layer=licon1_PDIFF $count=2 $X=0.78
+ $Y=1.84 $X2=0.93 $Y2=2.41
.ends

.subckt PM_SKY130_FD_SC_LS__A311OI_1%Y 1 2 3 11 13 14 15 16 20 22 24 28 30 37 45
r69 44 45 11.9052 $w=8.28e-07 $l=1.85e-07 $layer=LI1_cond $X=1.855 $Y=0.765
+ $X2=2.04 $Y2=0.765
r70 30 44 2.52185 $w=8.28e-07 $l=1.75e-07 $layer=LI1_cond $X=1.68 $Y=0.765
+ $X2=1.855 $Y2=0.765
r71 28 30 6.91708 $w=8.28e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=0.765
+ $X2=1.68 $Y2=0.765
r72 28 37 10.8964 $w=8.28e-07 $l=1.15e-07 $layer=LI1_cond $X=1.2 $Y=0.765
+ $X2=1.085 $Y2=0.765
r73 22 27 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.94 $Y=2.12 $X2=2.94
+ $Y2=2.035
r74 22 24 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=2.94 $Y=2.12
+ $X2=2.94 $Y2=2.815
r75 18 20 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=2.915 $Y=1.01
+ $X2=2.915 $Y2=0.515
r76 16 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.75 $Y=1.095
+ $X2=2.915 $Y2=1.01
r77 16 45 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=2.75 $Y=1.095
+ $X2=2.04 $Y2=1.095
r78 14 27 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.775 $Y=2.035
+ $X2=2.94 $Y2=2.035
r79 14 15 126.567 $w=1.68e-07 $l=1.94e-06 $layer=LI1_cond $X=2.775 $Y=2.035
+ $X2=0.835 $Y2=2.035
r80 13 37 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.835 $Y=1.095
+ $X2=1.085 $Y2=1.095
r81 11 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.75 $Y=1.95
+ $X2=0.835 $Y2=2.035
r82 10 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.75 $Y=1.18
+ $X2=0.835 $Y2=1.095
r83 10 11 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=0.75 $Y=1.18
+ $X2=0.75 $Y2=1.95
r84 3 27 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=2.79
+ $Y=1.84 $X2=2.94 $Y2=2.115
r85 3 24 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.79
+ $Y=1.84 $X2=2.94 $Y2=2.815
r86 2 20 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.775
+ $Y=0.37 $X2=2.915 $Y2=0.515
r87 1 44 91 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=2 $X=1.695
+ $Y=0.37 $X2=1.855 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__A311OI_1%VGND 1 2 9 13 16 17 19 20 21 34 35
r34 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r35 32 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r36 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r37 28 31 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.72 $Y=0 $X2=2.16
+ $Y2=0
r38 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r39 25 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r40 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r41 21 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r42 21 29 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r43 19 31 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=2.21 $Y=0 $X2=2.16
+ $Y2=0
r44 19 20 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=2.21 $Y=0 $X2=2.395
+ $Y2=0
r45 18 34 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=2.58 $Y=0 $X2=3.12
+ $Y2=0
r46 18 20 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=2.58 $Y=0 $X2=2.395
+ $Y2=0
r47 16 24 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=0.34 $Y=0 $X2=0.24
+ $Y2=0
r48 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.34 $Y=0 $X2=0.505
+ $Y2=0
r49 15 28 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=0.67 $Y=0 $X2=0.72
+ $Y2=0
r50 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.67 $Y=0 $X2=0.505
+ $Y2=0
r51 11 20 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.395 $Y=0.085
+ $X2=2.395 $Y2=0
r52 11 13 18.3768 $w=3.68e-07 $l=5.9e-07 $layer=LI1_cond $X=2.395 $Y=0.085
+ $X2=2.395 $Y2=0.675
r53 7 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.505 $Y=0.085
+ $X2=0.505 $Y2=0
r54 7 9 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=0.505 $Y=0.085
+ $X2=0.505 $Y2=0.675
r55 2 13 182 $w=1.7e-07 $l=3.76597e-07 $layer=licon1_NDIFF $count=1 $X=2.235
+ $Y=0.37 $X2=2.395 $Y2=0.675
r56 1 9 182 $w=1.7e-07 $l=3.62146e-07 $layer=licon1_NDIFF $count=1 $X=0.38
+ $Y=0.37 $X2=0.505 $Y2=0.675
.ends

