* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
X0 a_472_388# a_200_74# a_412_140# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X1 VGND A_N a_200_74# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X2 X a_472_388# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X3 VPWR a_27_74# a_472_388# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 a_685_140# C a_882_137# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X5 a_412_140# a_200_74# a_472_388# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X6 a_472_388# a_200_74# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 a_412_140# a_27_74# a_685_140# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X8 VPWR a_200_74# a_472_388# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 VGND D a_882_137# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X10 VPWR a_472_388# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X11 a_882_137# D VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X12 a_472_388# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 VPWR a_472_388# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X14 VPWR A_N a_200_74# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 VGND a_472_388# X VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X16 a_685_140# a_27_74# a_412_140# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X17 VGND a_472_388# X VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X18 a_27_74# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 a_27_74# B_N VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X20 X a_472_388# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X21 X a_472_388# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X22 a_472_388# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X23 X a_472_388# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X24 a_882_137# C a_685_140# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X25 a_472_388# a_27_74# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X26 VPWR C a_472_388# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X27 VPWR D a_472_388# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends
