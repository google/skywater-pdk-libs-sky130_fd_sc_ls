* File: sky130_fd_sc_ls__and4_2.pex.spice
* Created: Fri Aug 28 13:05:09 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__AND4_2%A 2 3 5 8 10 11 12 16
c32 11 0 1.05466e-19 $X=0.505 $Y=1.3
r33 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.28
+ $Y=1.465 $X2=0.28 $Y2=1.465
r34 12 16 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=0.28 $Y=1.665 $X2=0.28
+ $Y2=1.465
r35 10 15 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=0.505 $Y=1.465
+ $X2=0.28 $Y2=1.465
r36 10 11 3.90195 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.465
+ $X2=0.505 $Y2=1.3
r37 6 11 34.7346 $w=1.65e-07 $l=1.35e-07 $layer=POLY_cond $X=0.64 $Y=1.3
+ $X2=0.505 $Y2=1.3
r38 6 8 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.64 $Y=1.3 $X2=0.64
+ $Y2=0.74
r39 3 5 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.595 $Y=1.885
+ $X2=0.595 $Y2=2.46
r40 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.595 $Y=1.795 $X2=0.595
+ $Y2=1.885
r41 1 11 34.7346 $w=1.65e-07 $l=3.7229e-07 $layer=POLY_cond $X=0.595 $Y=1.63
+ $X2=0.505 $Y2=1.3
r42 1 2 64.1371 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.595 $Y=1.63
+ $X2=0.595 $Y2=1.795
.ends

.subckt PM_SKY130_FD_SC_LS__AND4_2%B 3 5 6 8 9 10 11 16 18
c42 9 0 1.05466e-19 $X=1.2 $Y=0.555
r43 16 19 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.12 $Y=1.385
+ $X2=1.12 $Y2=1.55
r44 16 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.12 $Y=1.385
+ $X2=1.12 $Y2=1.22
r45 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.12
+ $Y=1.385 $X2=1.12 $Y2=1.385
r46 11 17 2.88111 $w=3.58e-07 $l=9e-08 $layer=LI1_cond $X=1.135 $Y=1.295
+ $X2=1.135 $Y2=1.385
r47 10 11 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=1.135 $Y=0.925
+ $X2=1.135 $Y2=1.295
r48 9 10 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=1.135 $Y=0.555
+ $X2=1.135 $Y2=0.925
r49 6 8 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.045 $Y=1.885
+ $X2=1.045 $Y2=2.46
r50 5 6 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.045 $Y=1.795 $X2=1.045
+ $Y2=1.885
r51 5 19 95.2339 $w=1.8e-07 $l=2.45e-07 $layer=POLY_cond $X=1.045 $Y=1.795
+ $X2=1.045 $Y2=1.55
r52 3 18 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.03 $Y=0.74 $X2=1.03
+ $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_LS__AND4_2%C 3 5 6 8 9 10 11 16 18
c39 18 0 1.05261e-19 $X=1.69 $Y=1.22
r40 16 19 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.69 $Y=1.385
+ $X2=1.69 $Y2=1.55
r41 16 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.69 $Y=1.385
+ $X2=1.69 $Y2=1.22
r42 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.69
+ $Y=1.385 $X2=1.69 $Y2=1.385
r43 11 17 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=1.69 $Y=1.295 $X2=1.69
+ $Y2=1.385
r44 10 11 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.69 $Y=0.925
+ $X2=1.69 $Y2=1.295
r45 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.69 $Y=0.555
+ $X2=1.69 $Y2=0.925
r46 6 8 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.705 $Y=1.885
+ $X2=1.705 $Y2=2.46
r47 5 6 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.705 $Y=1.795 $X2=1.705
+ $Y2=1.885
r48 5 19 95.2339 $w=1.8e-07 $l=2.45e-07 $layer=POLY_cond $X=1.705 $Y=1.795
+ $X2=1.705 $Y2=1.55
r49 3 18 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.6 $Y=0.74 $X2=1.6
+ $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_LS__AND4_2%D 3 6 9 10 11 14 15 16
c41 15 0 1.05261e-19 $X=2.26 $Y=1.385
r42 14 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.26 $Y=1.385
+ $X2=2.26 $Y2=1.55
r43 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.26 $Y=1.385
+ $X2=2.26 $Y2=1.22
r44 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.26
+ $Y=1.385 $X2=2.26 $Y2=1.385
r45 11 15 3.11471 $w=3.68e-07 $l=1e-07 $layer=LI1_cond $X=2.16 $Y=1.365 $X2=2.26
+ $Y2=1.365
r46 9 10 41.3838 $w=1.65e-07 $l=9.5e-08 $layer=POLY_cond $X=2.162 $Y=1.79
+ $X2=2.162 $Y2=1.885
r47 9 17 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=2.17 $Y=1.79 $X2=2.17
+ $Y2=1.55
r48 6 16 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.17 $Y=0.74 $X2=2.17
+ $Y2=1.22
r49 3 10 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.155 $Y=2.46
+ $X2=2.155 $Y2=1.885
.ends

.subckt PM_SKY130_FD_SC_LS__AND4_2%A_56_74# 1 2 3 12 14 16 19 21 23 24 31 34 37
+ 41 46 49 51 55 56 60 62 63
r114 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.57
+ $Y=1.465 $X2=3.57 $Y2=1.465
r115 53 55 29.8588 $w=3.28e-07 $l=8.55e-07 $layer=LI1_cond $X=3.57 $Y=2.32
+ $X2=3.57 $Y2=1.465
r116 52 63 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.095 $Y=2.405
+ $X2=1.93 $Y2=2.405
r117 51 53 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.405 $Y=2.405
+ $X2=3.57 $Y2=2.32
r118 51 52 85.4652 $w=1.68e-07 $l=1.31e-06 $layer=LI1_cond $X=3.405 $Y=2.405
+ $X2=2.095 $Y2=2.405
r119 47 63 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.93 $Y=2.49
+ $X2=1.93 $Y2=2.405
r120 47 49 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=1.93 $Y=2.49
+ $X2=1.93 $Y2=2.815
r121 44 63 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.93 $Y=2.32
+ $X2=1.93 $Y2=2.405
r122 44 46 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=1.93 $Y=2.32
+ $X2=1.93 $Y2=2.105
r123 43 46 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=1.93 $Y=1.89
+ $X2=1.93 $Y2=2.105
r124 42 62 3.05049 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=0.985 $Y=1.805
+ $X2=0.8 $Y2=1.805
r125 41 43 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.765 $Y=1.805
+ $X2=1.93 $Y2=1.89
r126 41 42 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=1.765 $Y=1.805
+ $X2=0.985 $Y2=1.805
r127 37 39 22.1144 $w=3.68e-07 $l=7.1e-07 $layer=LI1_cond $X=0.8 $Y=2.105
+ $X2=0.8 $Y2=2.815
r128 35 62 3.46198 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.8 $Y=1.89 $X2=0.8
+ $Y2=1.805
r129 35 37 6.69663 $w=3.68e-07 $l=2.15e-07 $layer=LI1_cond $X=0.8 $Y=1.89
+ $X2=0.8 $Y2=2.105
r130 34 62 3.46198 $w=2.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=0.7 $Y=1.72
+ $X2=0.8 $Y2=1.805
r131 33 60 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.7 $Y=1.13 $X2=0.7
+ $Y2=1.045
r132 33 34 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=0.7 $Y=1.13 $X2=0.7
+ $Y2=1.72
r133 29 60 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.425 $Y=1.045
+ $X2=0.7 $Y2=1.045
r134 29 31 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=0.425 $Y=0.96
+ $X2=0.425 $Y2=0.515
r135 27 28 6.78005 $w=3.91e-07 $l=5.5e-08 $layer=POLY_cond $X=3.17 $Y=1.532
+ $X2=3.225 $Y2=1.532
r136 26 27 48.6931 $w=3.91e-07 $l=3.95e-07 $layer=POLY_cond $X=2.775 $Y=1.532
+ $X2=3.17 $Y2=1.532
r137 25 26 4.31458 $w=3.91e-07 $l=3.5e-08 $layer=POLY_cond $X=2.74 $Y=1.532
+ $X2=2.775 $Y2=1.532
r138 24 56 44.5896 $w=3.3e-07 $l=2.55e-07 $layer=POLY_cond $X=3.315 $Y=1.465
+ $X2=3.57 $Y2=1.465
r139 24 28 12.4078 $w=3.91e-07 $l=1.1887e-07 $layer=POLY_cond $X=3.315 $Y=1.465
+ $X2=3.225 $Y2=1.532
r140 21 28 25.3065 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=3.225 $Y=1.765
+ $X2=3.225 $Y2=1.532
r141 21 23 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.225 $Y=1.765
+ $X2=3.225 $Y2=2.4
r142 17 27 25.3065 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=3.17 $Y=1.3
+ $X2=3.17 $Y2=1.532
r143 17 19 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.17 $Y=1.3
+ $X2=3.17 $Y2=0.74
r144 14 26 25.3065 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=2.775 $Y=1.765
+ $X2=2.775 $Y2=1.532
r145 14 16 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.775 $Y=1.765
+ $X2=2.775 $Y2=2.4
r146 10 25 25.3065 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=2.74 $Y=1.3
+ $X2=2.74 $Y2=1.532
r147 10 12 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.74 $Y=1.3
+ $X2=2.74 $Y2=0.74
r148 3 49 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=1.78
+ $Y=1.96 $X2=1.93 $Y2=2.815
r149 3 46 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.78
+ $Y=1.96 $X2=1.93 $Y2=2.105
r150 2 39 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=0.67
+ $Y=1.96 $X2=0.82 $Y2=2.815
r151 2 37 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=0.67
+ $Y=1.96 $X2=0.82 $Y2=2.105
r152 1 31 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.28
+ $Y=0.37 $X2=0.425 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__AND4_2%VPWR 1 2 3 4 13 15 21 25 27 29 32 33 35 36 37
+ 46 55
r50 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r51 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r52 49 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r53 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r54 46 54 4.96106 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=3.37 $Y=3.33
+ $X2=3.605 $Y2=3.33
r55 46 48 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.37 $Y=3.33
+ $X2=3.12 $Y2=3.33
r56 45 49 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r57 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r58 42 52 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.24 $Y2=3.33
r59 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r60 39 51 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.222 $Y2=3.33
r61 39 41 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=1.2 $Y2=3.33
r62 37 45 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.16 $Y2=3.33
r63 37 42 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.2 $Y2=3.33
r64 35 44 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=2.3 $Y=3.33 $X2=2.16
+ $Y2=3.33
r65 35 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.3 $Y=3.33
+ $X2=2.465 $Y2=3.33
r66 34 48 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=2.63 $Y=3.33
+ $X2=3.12 $Y2=3.33
r67 34 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.63 $Y=3.33
+ $X2=2.465 $Y2=3.33
r68 32 41 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=1.215 $Y=3.33
+ $X2=1.2 $Y2=3.33
r69 32 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.215 $Y=3.33
+ $X2=1.38 $Y2=3.33
r70 31 44 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=1.545 $Y=3.33
+ $X2=2.16 $Y2=3.33
r71 31 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.545 $Y=3.33
+ $X2=1.38 $Y2=3.33
r72 27 54 3.01886 $w=3.55e-07 $l=1.1025e-07 $layer=LI1_cond $X=3.547 $Y=3.245
+ $X2=3.605 $Y2=3.33
r73 27 29 14.6084 $w=3.53e-07 $l=4.5e-07 $layer=LI1_cond $X=3.547 $Y=3.245
+ $X2=3.547 $Y2=2.795
r74 23 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.465 $Y=3.245
+ $X2=2.465 $Y2=3.33
r75 23 25 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=2.465 $Y=3.245
+ $X2=2.465 $Y2=2.795
r76 19 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.38 $Y=3.245
+ $X2=1.38 $Y2=3.33
r77 19 21 36.6686 $w=3.28e-07 $l=1.05e-06 $layer=LI1_cond $X=1.38 $Y=3.245
+ $X2=1.38 $Y2=2.195
r78 15 18 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=0.28 $Y=2.115 $X2=0.28
+ $Y2=2.815
r79 13 51 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.222 $Y2=3.33
r80 13 18 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.28 $Y2=2.815
r81 4 29 600 $w=1.7e-07 $l=1.07051e-06 $layer=licon1_PDIFF $count=1 $X=3.3
+ $Y=1.84 $X2=3.545 $Y2=2.795
r82 3 25 600 $w=1.7e-07 $l=9.45225e-07 $layer=licon1_PDIFF $count=1 $X=2.23
+ $Y=1.96 $X2=2.465 $Y2=2.795
r83 2 21 300 $w=1.7e-07 $l=3.58748e-07 $layer=licon1_PDIFF $count=2 $X=1.12
+ $Y=1.96 $X2=1.38 $Y2=2.195
r84 1 18 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.28 $Y2=2.815
r85 1 15 400 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.28 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_LS__AND4_2%X 1 2 7 8 9 10 26
r21 10 21 1.44055 $w=3.98e-07 $l=5e-08 $layer=LI1_cond $X=3.035 $Y=2.035
+ $X2=3.035 $Y2=1.985
r22 9 21 9.21954 $w=3.98e-07 $l=3.2e-07 $layer=LI1_cond $X=3.035 $Y=1.665
+ $X2=3.035 $Y2=1.985
r23 8 9 10.6601 $w=3.98e-07 $l=3.7e-07 $layer=LI1_cond $X=3.035 $Y=1.295
+ $X2=3.035 $Y2=1.665
r24 8 30 4.75383 $w=3.98e-07 $l=1.65e-07 $layer=LI1_cond $X=3.035 $Y=1.295
+ $X2=3.035 $Y2=1.13
r25 7 30 5.45223 $w=4.43e-07 $l=2.05e-07 $layer=LI1_cond $X=3.012 $Y=0.925
+ $X2=3.012 $Y2=1.13
r26 7 26 0.388464 $w=4.43e-07 $l=1.5e-08 $layer=LI1_cond $X=3.012 $Y=0.925
+ $X2=3.012 $Y2=0.91
r27 2 21 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.85
+ $Y=1.84 $X2=3 $Y2=1.985
r28 1 26 182 $w=1.7e-07 $l=6.0597e-07 $layer=licon1_NDIFF $count=1 $X=2.815
+ $Y=0.37 $X2=2.955 $Y2=0.91
.ends

.subckt PM_SKY130_FD_SC_LS__AND4_2%VGND 1 2 9 11 12 15 18 19 21 23 32 38
r42 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r43 35 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r44 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r45 32 37 5.51088 $w=1.7e-07 $l=3.1e-07 $layer=LI1_cond $X=3.22 $Y=0 $X2=3.53
+ $Y2=0
r46 32 34 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=3.22 $Y=0 $X2=3.12
+ $Y2=0
r47 31 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r48 30 31 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r49 26 30 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=2.16
+ $Y2=0
r50 26 27 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r51 23 31 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.16
+ $Y2=0
r52 23 27 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=1.92 $Y=0 $X2=0.24
+ $Y2=0
r53 21 22 4.31883 $w=4.33e-07 $l=8.5e-08 $layer=LI1_cond $X=3.437 $Y=0.515
+ $X2=3.437 $Y2=0.6
r54 18 30 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=2.265 $Y=0 $X2=2.16
+ $Y2=0
r55 18 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.265 $Y=0 $X2=2.43
+ $Y2=0
r56 17 34 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=2.595 $Y=0 $X2=3.12
+ $Y2=0
r57 17 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.595 $Y=0 $X2=2.43
+ $Y2=0
r58 15 22 14.5208 $w=2.48e-07 $l=3.15e-07 $layer=LI1_cond $X=3.53 $Y=0.915
+ $X2=3.53 $Y2=0.6
r59 12 21 3.49707 $w=4.33e-07 $l=1.32e-07 $layer=LI1_cond $X=3.437 $Y=0.383
+ $X2=3.437 $Y2=0.515
r60 11 37 3.16431 $w=4.35e-07 $l=1.28662e-07 $layer=LI1_cond $X=3.437 $Y=0.085
+ $X2=3.53 $Y2=0
r61 11 12 7.8949 $w=4.33e-07 $l=2.98e-07 $layer=LI1_cond $X=3.437 $Y=0.085
+ $X2=3.437 $Y2=0.383
r62 7 19 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.43 $Y=0.085 $X2=2.43
+ $Y2=0
r63 7 9 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=2.43 $Y=0.085 $X2=2.43
+ $Y2=0.495
r64 2 21 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.245
+ $Y=0.37 $X2=3.385 $Y2=0.515
r65 2 15 182 $w=1.7e-07 $l=6.56163e-07 $layer=licon1_NDIFF $count=1 $X=3.245
+ $Y=0.37 $X2=3.49 $Y2=0.915
r66 1 9 91 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=2 $X=2.245
+ $Y=0.37 $X2=2.43 $Y2=0.495
.ends

