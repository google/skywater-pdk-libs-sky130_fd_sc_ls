# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ls__mux2_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ls__mux2_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.640000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A0
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.640000 1.450000 7.075000 1.780000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.325000 1.450000 8.175000 1.780000 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  0.738000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 1.350000 0.835000 1.780000 ;
        RECT 0.665000 1.780000 0.835000 2.050000 ;
        RECT 0.665000 2.050000 1.675000 2.155000 ;
        RECT 0.665000 2.155000 3.165000 2.220000 ;
        RECT 1.505000 2.220000 3.165000 2.325000 ;
        RECT 2.995000 1.435000 3.745000 1.765000 ;
        RECT 2.995000 1.765000 3.165000 2.155000 ;
    END
  END S
  PIN X
    ANTENNADIFFAREA  1.576550 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.370000 2.755000 1.710000 ;
        RECT 1.085000 1.710000 2.770000 1.880000 ;
        RECT 1.310000 0.370000 1.640000 1.370000 ;
        RECT 2.330000 0.370000 2.755000 1.370000 ;
        RECT 2.440000 1.880000 2.770000 1.985000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 8.640000 0.085000 ;
        RECT 0.770000  0.085000 1.100000 1.150000 ;
        RECT 1.810000  0.085000 2.140000 1.070000 ;
        RECT 2.925000  0.085000 3.255000 1.255000 ;
        RECT 4.020000  0.085000 4.490000 0.905000 ;
        RECT 5.170000  0.085000 5.575000 0.585000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
        RECT 6.395000 -0.085000 6.565000 0.085000 ;
        RECT 6.875000 -0.085000 7.045000 0.085000 ;
        RECT 7.355000 -0.085000 7.525000 0.085000 ;
        RECT 7.835000 -0.085000 8.005000 0.085000 ;
        RECT 8.315000 -0.085000 8.485000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.640000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 8.640000 3.415000 ;
        RECT 0.650000 2.730000 0.995000 3.245000 ;
        RECT 1.820000 2.835000 2.150000 3.245000 ;
        RECT 3.060000 2.835000 3.390000 3.245000 ;
        RECT 4.130000 2.775000 4.460000 3.245000 ;
        RECT 5.200000 2.775000 5.450000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
        RECT 6.395000 3.245000 6.565000 3.415000 ;
        RECT 6.875000 3.245000 7.045000 3.415000 ;
        RECT 7.355000 3.245000 7.525000 3.415000 ;
        RECT 7.835000 3.245000 8.005000 3.415000 ;
        RECT 8.315000 3.245000 8.485000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 8.640000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085000 0.470000 0.600000 1.150000 ;
      RECT 0.085000 1.150000 0.255000 1.950000 ;
      RECT 0.085000 1.950000 0.445000 2.390000 ;
      RECT 0.085000 2.390000 1.335000 2.495000 ;
      RECT 0.085000 2.495000 3.505000 2.560000 ;
      RECT 0.085000 2.560000 0.445000 2.860000 ;
      RECT 1.165000 2.560000 3.505000 2.665000 ;
      RECT 3.335000 1.935000 4.085000 2.105000 ;
      RECT 3.335000 2.105000 3.505000 2.495000 ;
      RECT 3.520000 0.575000 3.850000 1.095000 ;
      RECT 3.520000 1.095000 5.325000 1.110000 ;
      RECT 3.520000 1.110000 8.020000 1.265000 ;
      RECT 3.675000 2.275000 3.925000 2.435000 ;
      RECT 3.675000 2.435000 5.790000 2.605000 ;
      RECT 3.675000 2.605000 3.925000 2.975000 ;
      RECT 3.915000 1.435000 4.985000 1.765000 ;
      RECT 3.915000 1.765000 4.085000 1.935000 ;
      RECT 4.660000 0.575000 4.990000 0.755000 ;
      RECT 4.660000 0.755000 5.665000 0.770000 ;
      RECT 4.660000 0.770000 7.090000 0.925000 ;
      RECT 4.665000 1.935000 5.140000 2.095000 ;
      RECT 4.665000 2.095000 6.130000 2.265000 ;
      RECT 5.155000 1.265000 8.020000 1.280000 ;
      RECT 5.385000 1.450000 6.470000 1.780000 ;
      RECT 5.495000 0.925000 7.090000 0.940000 ;
      RECT 5.620000 2.605000 5.790000 2.710000 ;
      RECT 5.620000 2.710000 7.115000 2.980000 ;
      RECT 5.835000 0.255000 8.525000 0.425000 ;
      RECT 5.835000 0.425000 6.590000 0.600000 ;
      RECT 5.960000 2.265000 6.130000 2.370000 ;
      RECT 5.960000 2.370000 8.025000 2.540000 ;
      RECT 6.300000 1.780000 6.470000 1.950000 ;
      RECT 6.300000 1.950000 8.525000 2.200000 ;
      RECT 6.760000 0.595000 7.090000 0.770000 ;
      RECT 7.260000 0.425000 7.590000 0.940000 ;
      RECT 7.695000 2.540000 8.025000 2.980000 ;
      RECT 7.770000 0.595000 8.020000 1.110000 ;
      RECT 8.190000 0.425000 8.525000 1.030000 ;
      RECT 8.195000 2.200000 8.525000 2.980000 ;
      RECT 8.355000 1.030000 8.525000 1.950000 ;
  END
END sky130_fd_sc_ls__mux2_4
