* NGSPICE file created from sky130_fd_sc_ls__xnor3_4.ext - technology: sky130A

.subckt sky130_fd_sc_ls__xnor3_4 A B C VGND VNB VPB VPWR X
M1000 a_75_227# A VGND VNB nshort w=640000u l=150000u
+  ad=5.611e+11p pd=4.74e+06u as=2.35215e+12p ps=1.359e+07u
M1001 X a_1057_74# VGND VNB nshort w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=0p ps=0u
M1002 a_324_373# B a_27_373# VNB nshort w=640000u l=150000u
+  ad=3.84e+11p pd=3.76e+06u as=4.635e+11p ps=4.06e+06u
M1003 a_27_373# a_386_23# a_321_77# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=3.739e+11p ps=3.78e+06u
M1004 a_75_227# a_386_23# a_324_373# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_324_373# C a_1057_74# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=2.592e+11p ps=2.09e+06u
M1006 VGND a_1057_74# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_27_373# a_386_23# a_324_373# VPB phighvt w=640000u l=150000u
+  ad=4.87e+11p pd=4.47e+06u as=6.528e+11p ps=5.05e+06u
M1008 X a_1057_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=6.72e+11p pd=5.68e+06u as=2.41e+12p ps=1.554e+07u
M1009 VGND a_1057_74# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_75_227# A VPWR VPB phighvt w=1e+06u l=150000u
+  ad=7.6215e+11p pd=5.69e+06u as=0p ps=0u
M1011 VPWR a_75_227# a_27_373# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND a_75_227# a_27_373# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND C a_1024_300# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1014 VPWR B a_386_23# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.304e+11p ps=2.83e+06u
M1015 a_321_77# B a_27_373# VPB phighvt w=640000u l=150000u
+  ad=5.312e+11p pd=4.67e+06u as=0p ps=0u
M1016 VPWR a_1057_74# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_75_227# a_386_23# a_321_77# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR C a_1024_300# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.888e+11p ps=1.87e+06u
M1019 VPWR a_1057_74# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_321_77# C a_1057_74# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=4.557e+11p ps=3.04e+06u
M1021 VGND B a_386_23# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1022 a_324_373# B a_75_227# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 X a_1057_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_321_77# B a_75_227# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_1057_74# a_1024_300# a_324_373# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_1057_74# a_1024_300# a_321_77# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 X a_1057_74# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

