* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_ls__nand4_2 A B C D VGND VNB VPB VPWR Y
*.PININFO A:I B:I C:I D:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMP0 Y A VPB phighvt m=2 w=1.12 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPB phighvt m=2 w=1.12 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 Y D VPB phighvt m=2 w=1.12 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPB phighvt m=2 w=1.12 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VNB nshort m=2 w=0.74 l=0.15 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
MMN1 sndA B VNB nshort m=2 w=0.74 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C VNB nshort m=2 w=0.74 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VNB nshort m=2 w=0.74 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_sc_ls__nand4_2
