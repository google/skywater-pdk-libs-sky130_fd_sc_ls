* File: sky130_fd_sc_ls__sdfbbn_1.spice
* Created: Wed Sep  2 11:26:31 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__sdfbbn_1.pex.spice"
.subckt sky130_fd_sc_ls__sdfbbn_1  VNB VPB SCD D SCE CLK_N SET_B RESET_B VPWR
+ Q_N Q VGND
* 
* VGND	VGND
* Q	Q
* Q_N	Q_N
* VPWR	VPWR
* RESET_B	RESET_B
* SET_B	SET_B
* CLK_N	CLK_N
* SCE	SCE
* D	D
* SCD	SCD
* VPB	VPB
* VNB	VNB
MM1004 A_119_119# N_SCD_M1004_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.4 A=0.063 P=1.14 MULT=1
MM1030 N_A_197_119#_M1030_d N_SCE_M1030_g A_119_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.0819 AS=0.0504 PD=0.81 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.6
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1000 A_305_119# N_D_M1000_g N_A_197_119#_M1030_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0819 PD=0.66 PS=0.81 NRD=18.564 NRS=31.428 M=1 R=2.8 SA=75001.1
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1031 N_VGND_M1031_d N_A_353_93#_M1031_g A_305_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.1449 AS=0.0504 PD=1.11 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.5
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1017 N_A_353_93#_M1017_d N_SCE_M1017_g N_VGND_M1031_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.1449 PD=1.41 PS=1.11 NRD=0 NRS=117.132 M=1 R=2.8 SA=75002.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1013 N_VGND_M1013_d N_CLK_N_M1013_g N_A_662_82#_M1013_s VNB NSHORT L=0.15
+ W=0.74 AD=0.19615 AS=0.2109 PD=1.41 PS=2.05 NRD=34.056 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.9 A=0.111 P=1.78 MULT=1
MM1014 N_A_867_82#_M1014_d N_A_662_82#_M1014_g N_VGND_M1013_d VNB NSHORT L=0.15
+ W=0.74 AD=0.3219 AS=0.19615 PD=2.35 PS=1.41 NRD=12.156 NRS=34.056 M=1
+ R=4.93333 SA=75000.8 SB=75000.4 A=0.111 P=1.78 MULT=1
MM1019 A_1151_119# N_A_977_243#_M1019_g N_VGND_M1019_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1015 N_A_1159_497#_M1015_d N_A_662_82#_M1015_g A_1151_119# VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1001 N_A_197_119#_M1001_d N_A_867_82#_M1001_g N_A_1159_497#_M1015_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.1491 AS=0.0588 PD=1.55 PS=0.7 NRD=21.42 NRS=0 M=1 R=2.8
+ SA=75001 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1005 N_A_977_243#_M1005_d N_A_1159_497#_M1005_g N_A_1434_78#_M1005_s VNB
+ NSHORT L=0.15 W=0.55 AD=0.1045 AS=0.2602 PD=0.93 PS=2.24 NRD=4.908 NRS=91.212
+ M=1 R=3.66667 SA=75000.3 SB=75004.9 A=0.0825 P=1.4 MULT=1
MM1045 N_A_1434_78#_M1045_d N_A_1579_258#_M1045_g N_A_977_243#_M1005_d VNB
+ NSHORT L=0.15 W=0.55 AD=0.125125 AS=0.1045 PD=1.005 PS=0.93 NRD=15.264 NRS=0
+ M=1 R=3.66667 SA=75000.8 SB=75004.4 A=0.0825 P=1.4 MULT=1
MM1021 N_VGND_M1021_d N_SET_B_M1021_g N_A_1434_78#_M1045_d VNB NSHORT L=0.15
+ W=0.55 AD=0.11275 AS=0.125125 PD=0.96 PS=1.005 NRD=0 NRS=22.908 M=1 R=3.66667
+ SA=75001.4 SB=75003.7 A=0.0825 P=1.4 MULT=1
MM1044 A_1876_119# N_A_977_243#_M1044_g N_VGND_M1021_d VNB NSHORT L=0.15 W=0.55
+ AD=0.066 AS=0.11275 PD=0.79 PS=0.96 NRD=14.172 NRS=28.356 M=1 R=3.66667
+ SA=75002 SB=75003.2 A=0.0825 P=1.4 MULT=1
MM1022 N_A_1954_119#_M1022_d N_A_662_82#_M1022_g A_1876_119# VNB NSHORT L=0.15
+ W=0.55 AD=0.272562 AS=0.066 PD=1.64433 PS=0.79 NRD=0 NRS=14.172 M=1 R=3.66667
+ SA=75002.4 SB=75002.8 A=0.0825 P=1.4 MULT=1
MM1040 A_2164_119# N_A_867_82#_M1040_g N_A_1954_119#_M1022_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0819 AS=0.208138 PD=0.81 PS=1.25567 NRD=39.996 NRS=32.856 M=1
+ R=2.8 SA=75003.4 SB=75002.4 A=0.063 P=1.14 MULT=1
MM1009 N_VGND_M1009_d N_A_2133_410#_M1009_g A_2164_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.128218 AS=0.0819 PD=0.99931 PS=0.81 NRD=71.508 NRS=39.996 M=1 R=2.8
+ SA=75004 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1010 N_A_2392_74#_M1010_d N_SET_B_M1010_g N_VGND_M1009_d VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.225907 PD=1.02 PS=1.76069 NRD=0 NRS=40.584 M=1 R=4.93333
+ SA=75002.7 SB=75001.2 A=0.111 P=1.78 MULT=1
MM1036 N_A_2133_410#_M1036_d N_A_1579_258#_M1036_g N_A_2392_74#_M1010_d VNB
+ NSHORT L=0.15 W=0.74 AD=0.1406 AS=0.1036 PD=1.12 PS=1.02 NRD=16.212 NRS=0 M=1
+ R=4.93333 SA=75003.1 SB=75000.8 A=0.111 P=1.78 MULT=1
MM1028 N_A_2392_74#_M1028_d N_A_1954_119#_M1028_g N_A_2133_410#_M1036_d VNB
+ NSHORT L=0.15 W=0.74 AD=0.2875 AS=0.1406 PD=2.33 PS=1.12 NRD=13.776 NRS=0 M=1
+ R=4.93333 SA=75003.7 SB=75000.3 A=0.111 P=1.78 MULT=1
MM1002 N_VGND_M1002_d N_RESET_B_M1002_g N_A_1579_258#_M1002_s VNB NSHORT L=0.15
+ W=0.42 AD=0.132372 AS=0.1197 PD=0.970345 PS=1.41 NRD=74.328 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001 A=0.063 P=1.14 MULT=1
MM1007 N_Q_N_M1007_d N_A_2133_410#_M1007_g N_VGND_M1002_d VNB NSHORT L=0.15
+ W=0.74 AD=0.2109 AS=0.233228 PD=2.05 PS=1.70966 NRD=0 NRS=5.664 M=1 R=4.93333
+ SA=75000.7 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1018 N_VGND_M1018_d N_A_2133_410#_M1018_g N_A_3078_384#_M1018_s VNB NSHORT
+ L=0.15 W=0.55 AD=0.107506 AS=0.15675 PD=0.937984 PS=1.67 NRD=17.988 NRS=0 M=1
+ R=3.66667 SA=75000.2 SB=75000.7 A=0.0825 P=1.4 MULT=1
MM1034 N_Q_M1034_d N_A_3078_384#_M1034_g N_VGND_M1018_d VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.144644 PD=2.05 PS=1.26202 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1025 N_VPWR_M1025_d N_SCD_M1025_g N_A_27_464#_M1025_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1056 AS=0.1888 PD=0.97 PS=1.87 NRD=3.0732 NRS=3.0732 M=1 R=4.26667
+ SA=75000.2 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1046 A_212_464# N_SCE_M1046_g N_VPWR_M1025_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0864 AS=0.1056 PD=0.91 PS=0.97 NRD=24.625 NRS=12.2928 M=1 R=4.26667
+ SA=75000.7 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1037 N_A_197_119#_M1037_d N_D_M1037_g A_212_464# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.096 AS=0.0864 PD=0.94 PS=0.91 NRD=3.0732 NRS=24.625 M=1 R=4.26667
+ SA=75001.1 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1003 N_A_27_464#_M1003_d N_A_353_93#_M1003_g N_A_197_119#_M1037_d VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.1856 AS=0.096 PD=1.86 PS=0.94 NRD=3.0732 NRS=3.0732 M=1
+ R=4.26667 SA=75001.6 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1016 N_A_353_93#_M1016_d N_SCE_M1016_g N_VPWR_M1016_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1888 AS=0.1888 PD=1.87 PS=1.87 NRD=3.0732 NRS=3.0732 M=1 R=4.26667
+ SA=75000.2 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1026 N_VPWR_M1026_d N_CLK_N_M1026_g N_A_662_82#_M1026_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1038 N_A_867_82#_M1038_d N_A_662_82#_M1038_g N_VPWR_M1026_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1023 A_1081_497# N_A_977_243#_M1023_g N_VPWR_M1023_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0504 AS=0.1239 PD=0.66 PS=1.43 NRD=30.4759 NRS=4.6886 M=1 R=2.8
+ SA=75000.2 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1006 N_A_1159_497#_M1006_d N_A_867_82#_M1006_g A_1081_497# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0897849 AS=0.0504 PD=0.812264 PS=0.66 NRD=46.886 NRS=30.4759 M=1
+ R=2.8 SA=75000.6 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1041 N_A_197_119#_M1041_d N_A_662_82#_M1041_g N_A_1159_497#_M1006_d VPB
+ PHIGHVT L=0.15 W=0.64 AD=0.2208 AS=0.136815 PD=1.97 PS=1.23774 NRD=18.4589
+ NRS=3.0732 M=1 R=4.26667 SA=75000.8 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1042 A_1528_424# N_A_1159_497#_M1042_g N_A_977_243#_M1042_s VPB PHIGHVT L=0.15
+ W=0.84 AD=0.1134 AS=0.3906 PD=1.11 PS=2.61 NRD=18.7544 NRS=3.5066 M=1 R=5.6
+ SA=75000.4 SB=75001.1 A=0.126 P=1.98 MULT=1
MM1033 N_VPWR_M1033_d N_A_1579_258#_M1033_g A_1528_424# VPB PHIGHVT L=0.15
+ W=0.84 AD=0.126 AS=0.1134 PD=1.14 PS=1.11 NRD=2.3443 NRS=18.7544 M=1 R=5.6
+ SA=75000.8 SB=75000.7 A=0.126 P=1.98 MULT=1
MM1043 N_A_977_243#_M1043_d N_SET_B_M1043_g N_VPWR_M1033_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.2436 AS=0.126 PD=2.26 PS=1.14 NRD=2.3443 NRS=2.3443 M=1 R=5.6
+ SA=75001.3 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1011 A_1903_424# N_A_977_243#_M1011_g N_VPWR_M1011_s VPB PHIGHVT L=0.15 W=0.84
+ AD=0.1008 AS=0.2478 PD=1.08 PS=2.27 NRD=15.2281 NRS=2.3443 M=1 R=5.6
+ SA=75000.2 SB=75001.1 A=0.126 P=1.98 MULT=1
MM1029 N_A_1954_119#_M1029_d N_A_867_82#_M1029_g A_1903_424# VPB PHIGHVT L=0.15
+ W=0.84 AD=0.1904 AS=0.1008 PD=1.63333 PS=1.08 NRD=2.3443 NRS=15.2281 M=1 R=5.6
+ SA=75000.6 SB=75000.7 A=0.126 P=1.98 MULT=1
MM1035 A_2088_508# N_A_662_82#_M1035_g N_A_1954_119#_M1029_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0504 AS=0.0952 PD=0.66 PS=0.816667 NRD=30.4759 NRS=44.5417 M=1
+ R=2.8 SA=75001.1 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1008 N_VPWR_M1008_d N_A_2133_410#_M1008_g A_2088_508# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.22775 AS=0.0504 PD=2.07 PS=0.66 NRD=228.54 NRS=30.4759 M=1 R=2.8
+ SA=75001.5 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1039 N_VPWR_M1039_d N_SET_B_M1039_g N_A_2133_410#_M1039_s VPB PHIGHVT L=0.15
+ W=1 AD=0.269075 AS=0.295 PD=1.705 PS=2.59 NRD=42.158 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75001.3 A=0.15 P=2.3 MULT=1
MM1032 A_2509_392# N_A_1579_258#_M1032_g N_VPWR_M1039_d VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.269075 PD=1.27 PS=1.705 NRD=15.7403 NRS=42.158 M=1 R=6.66667
+ SA=75000.8 SB=75000.6 A=0.15 P=2.3 MULT=1
MM1020 N_A_2133_410#_M1020_d N_A_1954_119#_M1020_g A_2509_392# VPB PHIGHVT
+ L=0.15 W=1 AD=0.295 AS=0.135 PD=2.59 PS=1.27 NRD=1.9503 NRS=15.7403 M=1
+ R=6.66667 SA=75001.3 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1027 N_VPWR_M1027_d N_RESET_B_M1027_g N_A_1579_258#_M1027_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.199855 AS=0.3625 PD=1.29455 PS=3.71 NRD=3.0732 NRS=157.403 M=1
+ R=4.26667 SA=75000.2 SB=75001 A=0.096 P=1.58 MULT=1
MM1047 N_Q_N_M1047_d N_A_2133_410#_M1047_g N_VPWR_M1027_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.3304 AS=0.349745 PD=2.83 PS=2.26545 NRD=1.7533 NRS=1.7533 M=1
+ R=7.46667 SA=75000.7 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1024 N_VPWR_M1024_d N_A_2133_410#_M1024_g N_A_3078_384#_M1024_s VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.174 AS=0.2478 PD=1.29 PS=2.27 NRD=22.655 NRS=2.3443 M=1
+ R=5.6 SA=75000.2 SB=75000.8 A=0.126 P=1.98 MULT=1
MM1012 N_Q_M1012_d N_A_3078_384#_M1012_g N_VPWR_M1024_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.3304 AS=0.232 PD=2.83 PS=1.72 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.6 SB=75000.2 A=0.168 P=2.54 MULT=1
DX48_noxref VNB VPB NWDIODE A=32.1616 P=38.3
c_196 VNB 0 1.86341e-19 $X=0 $Y=0
c_2466 A_212_464# 0 1.00461e-19 $X=1.06 $Y=2.32
*
.include "sky130_fd_sc_ls__sdfbbn_1.pxi.spice"
*
.ends
*
*
