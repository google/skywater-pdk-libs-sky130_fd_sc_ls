* NGSPICE file created from sky130_fd_sc_ls__a221oi_2.ext - technology: sky130A

.subckt sky130_fd_sc_ls__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
M1000 a_294_368# B1 a_29_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=1.3776e+12p pd=1.142e+07u as=1.288e+12p ps=1.126e+07u
M1001 VGND B2 a_293_74# VNB nshort w=740000u l=150000u
+  ad=7.696e+11p pd=6.52e+06u as=4.44e+11p ps=4.16e+06u
M1002 a_29_368# B1 a_294_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_293_74# B1 Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=8.362e+11p ps=8.18e+06u
M1004 a_294_368# A1 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=9.52e+11p ps=8.42e+06u
M1005 a_675_74# A2 VGND VNB nshort w=740000u l=150000u
+  ad=7.03e+11p pd=4.86e+06u as=0p ps=0u
M1006 Y A1 a_675_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND A2 a_675_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_293_74# B2 VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR A2 a_294_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_294_368# A2 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_29_368# B2 a_294_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_675_74# A1 Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR A1 a_294_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Y B1 a_293_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y C1 VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Y C1 a_29_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=0p ps=0u
M1017 a_29_368# C1 Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_294_368# B2 a_29_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND C1 Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

