* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__dlrtn_4 D GATE_N RESET_B VGND VNB VPB VPWR Q
X0 VPWR RESET_B a_888_406# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X1 VGND GATE_N a_232_98# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X2 VPWR a_888_406# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X3 a_888_406# a_639_392# a_1035_74# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X4 a_666_74# a_232_98# a_639_392# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X5 a_1035_74# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X6 VPWR GATE_N a_232_98# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X7 VGND RESET_B a_1035_74# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X8 a_348_392# a_232_98# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X9 a_348_392# a_232_98# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X10 a_27_136# D VGND VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X11 VPWR a_639_392# a_888_406# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X12 a_839_74# a_888_406# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 VGND a_888_406# Q VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X14 Q a_888_406# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X15 a_888_406# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X16 VGND a_888_406# Q VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X17 Q a_888_406# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X18 VPWR a_27_136# a_561_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 VGND a_27_136# a_666_74# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X20 a_639_392# a_348_392# a_839_74# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X21 a_639_392# a_232_98# a_747_504# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X22 VPWR a_888_406# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X23 Q a_888_406# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X24 Q a_888_406# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X25 a_888_406# a_639_392# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X26 a_27_136# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X27 a_747_504# a_888_406# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X28 a_561_392# a_348_392# a_639_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X29 a_1035_74# a_639_392# a_888_406# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
.ends
