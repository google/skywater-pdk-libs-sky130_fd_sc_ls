* File: sky130_fd_sc_ls__edfxtp_1.pex.spice
* Created: Fri Aug 28 13:23:13 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__EDFXTP_1%D 2 3 5 8 12 13 18 19 21 23
c46 19 0 6.23793e-20 $X=0.52 $Y=1.145
c47 2 0 1.15294e-19 $X=0.495 $Y=2.375
r48 21 23 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.52 $Y=1.825
+ $X2=0.52 $Y2=1.99
r49 21 22 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.52
+ $Y=1.825 $X2=0.52 $Y2=1.825
r50 18 21 118.906 $w=3.3e-07 $l=6.8e-07 $layer=POLY_cond $X=0.52 $Y=1.145
+ $X2=0.52 $Y2=1.825
r51 18 19 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.52
+ $Y=1.145 $X2=0.52 $Y2=1.145
r52 13 22 4.85239 $w=3.78e-07 $l=1.6e-07 $layer=LI1_cond $X=0.615 $Y=1.665
+ $X2=0.615 $Y2=1.825
r53 12 13 11.2212 $w=3.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.615 $Y=1.295
+ $X2=0.615 $Y2=1.665
r54 12 19 4.54912 $w=3.78e-07 $l=1.5e-07 $layer=LI1_cond $X=0.615 $Y=1.295
+ $X2=0.615 $Y2=1.145
r55 11 18 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.52 $Y=0.98
+ $X2=0.52 $Y2=1.145
r56 8 11 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=0.58 $Y=0.58 $X2=0.58
+ $Y2=0.98
r57 3 5 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.495 $Y=2.465
+ $X2=0.495 $Y2=2.75
r58 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.495 $Y=2.375 $X2=0.495
+ $Y2=2.465
r59 2 23 149.653 $w=1.8e-07 $l=3.85e-07 $layer=POLY_cond $X=0.495 $Y=2.375
+ $X2=0.495 $Y2=1.99
.ends

.subckt PM_SKY130_FD_SC_LS__EDFXTP_1%A_159_446# 1 2 7 9 11 14 16 19 23 24 25 26
+ 27 28 31 35 37 39 41 50
c127 50 0 1.98585e-19 $X=2.38 $Y=1.55
c128 41 0 1.9156e-19 $X=2.22 $Y=1.55
c129 39 0 1.34182e-19 $X=1.79 $Y=1.695
c130 28 0 1.15294e-19 $X=1.305 $Y=1.695
c131 25 0 1.9799e-19 $X=1.57 $Y=0.855
c132 16 0 6.23793e-20 $X=0.885 $Y=2.347
r133 42 50 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=2.22 $Y=1.55
+ $X2=2.38 $Y2=1.55
r134 41 44 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=2.22 $Y=1.55
+ $X2=2.22 $Y2=1.695
r135 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.22
+ $Y=1.55 $X2=2.22 $Y2=1.55
r136 38 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.875 $Y=1.695
+ $X2=1.79 $Y2=1.695
r137 37 44 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.055 $Y=1.695
+ $X2=2.22 $Y2=1.695
r138 37 38 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.055 $Y=1.695
+ $X2=1.875 $Y2=1.695
r139 33 39 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.79 $Y=1.78
+ $X2=1.79 $Y2=1.695
r140 33 35 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=1.79 $Y=1.78
+ $X2=1.79 $Y2=2.495
r141 29 31 5.76222 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=1.695 $Y=0.77
+ $X2=1.695 $Y2=0.645
r142 27 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.705 $Y=1.695
+ $X2=1.79 $Y2=1.695
r143 27 28 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=1.705 $Y=1.695
+ $X2=1.305 $Y2=1.695
r144 25 29 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.57 $Y=0.855
+ $X2=1.695 $Y2=0.77
r145 25 26 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.57 $Y=0.855
+ $X2=1.305 $Y2=0.855
r146 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.14
+ $Y=1.505 $X2=1.14 $Y2=1.505
r147 21 28 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.14 $Y=1.61
+ $X2=1.305 $Y2=1.695
r148 21 23 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=1.14 $Y=1.61
+ $X2=1.14 $Y2=1.505
r149 20 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.14 $Y=0.94
+ $X2=1.305 $Y2=0.855
r150 20 23 19.7312 $w=3.28e-07 $l=5.65e-07 $layer=LI1_cond $X=1.14 $Y=0.94
+ $X2=1.14 $Y2=1.505
r151 18 24 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.14 $Y=1.845
+ $X2=1.14 $Y2=1.505
r152 18 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.14 $Y=1.845
+ $X2=1.14 $Y2=2.01
r153 16 17 40.5765 $w=1.96e-07 $l=1.65e-07 $layer=POLY_cond $X=0.885 $Y=2.347
+ $X2=1.05 $Y2=2.347
r154 12 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.38 $Y=1.385
+ $X2=2.38 $Y2=1.55
r155 12 14 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=2.38 $Y=1.385
+ $X2=2.38 $Y2=0.645
r156 11 17 9.11062 $w=1.5e-07 $l=1.17e-07 $layer=POLY_cond $X=1.05 $Y=2.23
+ $X2=1.05 $Y2=2.347
r157 11 19 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=1.05 $Y=2.23
+ $X2=1.05 $Y2=2.01
r158 7 16 9.11062 $w=1.5e-07 $l=1.18e-07 $layer=POLY_cond $X=0.885 $Y=2.465
+ $X2=0.885 $Y2=2.347
r159 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.885 $Y=2.465
+ $X2=0.885 $Y2=2.75
r160 2 35 600 $w=1.7e-07 $l=3.80657e-07 $layer=licon1_PDIFF $count=1 $X=1.645
+ $Y=2.18 $X2=1.79 $Y2=2.495
r161 1 31 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.595
+ $Y=0.435 $X2=1.735 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_LS__EDFXTP_1%DE 3 5 6 10 11 13 14 16 17 18 19 21 22 26
+ 29 31
c89 31 0 3.25741e-19 $X=1.68 $Y=1.44
c90 26 0 1.98585e-19 $X=1.68 $Y=1.295
c91 10 0 3.01092e-20 $X=1.74 $Y=1.955
r92 29 31 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.68 $Y=1.275
+ $X2=1.68 $Y2=1.44
r93 26 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.68
+ $Y=1.275 $X2=1.68 $Y2=1.275
r94 23 25 141.011 $w=1.5e-07 $l=2.75e-07 $layer=POLY_cond $X=1.74 $Y=2.03
+ $X2=2.015 $Y2=2.03
r95 19 21 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.695 $Y=2.105
+ $X2=2.695 $Y2=2.39
r96 18 25 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.09 $Y=2.03
+ $X2=2.015 $Y2=2.03
r97 17 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.62 $Y=2.03
+ $X2=2.695 $Y2=2.105
r98 17 18 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.62 $Y=2.03
+ $X2=2.09 $Y2=2.03
r99 14 25 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.015 $Y=2.105
+ $X2=2.015 $Y2=2.03
r100 14 16 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.015 $Y=2.105
+ $X2=2.015 $Y2=2.5
r101 11 22 13.5877 $w=2.4e-07 $l=2.14243e-07 $layer=POLY_cond $X=1.95 $Y=0.95
+ $X2=1.77 $Y2=1.025
r102 11 13 98.0067 $w=1.5e-07 $l=3.05e-07 $layer=POLY_cond $X=1.95 $Y=0.95
+ $X2=1.95 $Y2=0.645
r103 10 23 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.74 $Y=1.955
+ $X2=1.74 $Y2=2.03
r104 10 31 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=1.74 $Y=1.955
+ $X2=1.74 $Y2=1.44
r105 7 22 13.5877 $w=2.4e-07 $l=1.21861e-07 $layer=POLY_cond $X=1.68 $Y=1.1
+ $X2=1.77 $Y2=1.025
r106 7 29 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=1.68 $Y=1.1
+ $X2=1.68 $Y2=1.275
r107 5 22 12.1617 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=1.515 $Y=1.025
+ $X2=1.77 $Y2=1.025
r108 5 6 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=1.515 $Y=1.025 $X2=1.045
+ $Y2=1.025
r109 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.97 $Y=0.95
+ $X2=1.045 $Y2=1.025
r110 1 3 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=0.97 $Y=0.95 $X2=0.97
+ $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_LS__EDFXTP_1%A_533_61# 1 2 9 12 13 15 16 18 19 20 21 23
+ 25 26 33 36 40 43 44 45 51 52 55 56 65
c201 44 0 2.65373e-20 $X=11.615 $Y=1.665
r202 55 58 76.7264 $w=5.1e-07 $l=5.05e-07 $layer=POLY_cond $X=2.92 $Y=1.21
+ $X2=2.92 $Y2=1.715
r203 55 57 46.8261 $w=5.1e-07 $l=1.65e-07 $layer=POLY_cond $X=2.92 $Y=1.21
+ $X2=2.92 $Y2=1.045
r204 55 56 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.83
+ $Y=1.21 $X2=2.83 $Y2=1.21
r205 52 65 6.51792 $w=2.38e-07 $l=1.15e-07 $layer=LI1_cond $X=11.765 $Y=1.665
+ $X2=11.765 $Y2=1.55
r206 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=1.665
+ $X2=11.76 $Y2=1.665
r207 48 56 13.983 $w=3.73e-07 $l=4.55e-07 $layer=LI1_cond $X=2.742 $Y=1.665
+ $X2=2.742 $Y2=1.21
r208 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=1.665
+ $X2=2.64 $Y2=1.665
r209 45 47 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.785 $Y=1.665
+ $X2=2.64 $Y2=1.665
r210 44 51 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=11.615 $Y=1.665
+ $X2=11.76 $Y2=1.665
r211 44 45 10.9282 $w=1.4e-07 $l=8.83e-06 $layer=MET1_cond $X=11.615 $Y=1.665
+ $X2=2.785 $Y2=1.665
r212 42 65 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=11.76 $Y=0.81
+ $X2=11.76 $Y2=1.55
r213 40 42 10.9338 $w=3.53e-07 $l=2.4e-07 $layer=LI1_cond $X=11.667 $Y=0.57
+ $X2=11.667 $Y2=0.81
r214 36 43 4.2255 $w=2.85e-07 $l=1.32605e-07 $layer=LI1_cond $X=11.765 $Y=2.095
+ $X2=11.72 $Y2=2.207
r215 35 52 0.240092 $w=2.38e-07 $l=5e-09 $layer=LI1_cond $X=11.765 $Y=1.67
+ $X2=11.765 $Y2=1.665
r216 35 36 20.4078 $w=2.38e-07 $l=4.25e-07 $layer=LI1_cond $X=11.765 $Y=1.67
+ $X2=11.765 $Y2=2.095
r217 31 43 4.2255 $w=2.85e-07 $l=1.13e-07 $layer=LI1_cond $X=11.72 $Y=2.32
+ $X2=11.72 $Y2=2.207
r218 31 33 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=11.72 $Y=2.32
+ $X2=11.72 $Y2=2.435
r219 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.83
+ $Y=2.185 $X2=10.83 $Y2=2.185
r220 26 43 2.20607 $w=2.25e-07 $l=1.65e-07 $layer=LI1_cond $X=11.555 $Y=2.207
+ $X2=11.72 $Y2=2.207
r221 26 28 37.1343 $w=2.23e-07 $l=7.25e-07 $layer=LI1_cond $X=11.555 $Y=2.207
+ $X2=10.83 $Y2=2.207
r222 25 29 38.5562 $w=2.99e-07 $l=1.92678e-07 $layer=POLY_cond $X=10.89 $Y=2.02
+ $X2=10.83 $Y2=2.185
r223 24 25 515.33 $w=1.5e-07 $l=1.005e-06 $layer=POLY_cond $X=10.89 $Y=1.015
+ $X2=10.89 $Y2=2.02
r224 21 29 52.2586 $w=2.99e-07 $l=2.7157e-07 $layer=POLY_cond $X=10.785 $Y=2.435
+ $X2=10.83 $Y2=2.185
r225 21 23 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=10.785 $Y=2.435
+ $X2=10.785 $Y2=2.72
r226 19 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.815 $Y=0.94
+ $X2=10.89 $Y2=1.015
r227 19 20 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=10.815 $Y=0.94
+ $X2=10.375 $Y2=0.94
r228 16 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.3 $Y=0.865
+ $X2=10.375 $Y2=0.94
r229 16 18 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=10.3 $Y=0.865
+ $X2=10.3 $Y2=0.58
r230 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.085 $Y=2.105
+ $X2=3.085 $Y2=2.39
r231 12 13 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.085 $Y=2.015
+ $X2=3.085 $Y2=2.105
r232 12 58 116.613 $w=1.8e-07 $l=3e-07 $layer=POLY_cond $X=3.085 $Y=2.015
+ $X2=3.085 $Y2=1.715
r233 9 57 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.74 $Y=0.645 $X2=2.74
+ $Y2=1.045
r234 2 33 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=11.57
+ $Y=2.29 $X2=11.72 $Y2=2.435
r235 1 40 182 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=1 $X=11.48
+ $Y=0.37 $X2=11.62 $Y2=0.57
.ends

.subckt PM_SKY130_FD_SC_LS__EDFXTP_1%CLK 3 4 6 8 9 11 14 16
c43 14 0 1.4577e-19 $X=3.615 $Y=1.385
r44 14 17 14.2284 $w=3.65e-07 $l=9e-08 $layer=POLY_cond $X=3.632 $Y=1.385
+ $X2=3.632 $Y2=1.475
r45 14 16 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=3.632 $Y=1.385
+ $X2=3.632 $Y2=1.22
r46 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.615
+ $Y=1.385 $X2=3.615 $Y2=1.385
r47 11 15 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=3.615 $Y=1.295
+ $X2=3.615 $Y2=1.385
r48 6 9 83.7788 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=4.06 $Y=1.685 $X2=4.06
+ $Y2=1.475
r49 6 8 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.06 $Y=1.685
+ $X2=4.06 $Y2=2.32
r50 5 17 23.6381 $w=1.5e-07 $l=1.83e-07 $layer=POLY_cond $X=3.815 $Y=1.475
+ $X2=3.632 $Y2=1.475
r51 4 9 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.97 $Y=1.475 $X2=4.06
+ $Y2=1.475
r52 4 5 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=3.97 $Y=1.475
+ $X2=3.815 $Y2=1.475
r53 3 16 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.74 $Y=0.74 $X2=3.74
+ $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_LS__EDFXTP_1%A_958_74# 1 2 7 9 10 12 15 17 18 20 23 25
+ 26 27 32 33 36 37 40 41 42 44 45 46 47 49 50 53 56 59 61 64 65 69 76
c223 69 0 2.65373e-20 $X=10.44 $Y=1.42
c224 56 0 2.80716e-20 $X=6.67 $Y=1.145
c225 53 0 1.6161e-19 $X=6.085 $Y=2.135
c226 40 0 1.62788e-19 $X=7.675 $Y=0.935
c227 10 0 1.96074e-19 $X=6.67 $Y=0.98
r228 69 80 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.44 $Y=1.42
+ $X2=10.44 $Y2=1.585
r229 68 69 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.44
+ $Y=1.42 $X2=10.44 $Y2=1.42
r230 65 68 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=10.44 $Y=1.29
+ $X2=10.44 $Y2=1.42
r231 64 76 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.36 $Y=1.385
+ $X2=9.36 $Y2=1.22
r232 63 64 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.36
+ $Y=1.385 $X2=9.36 $Y2=1.385
r233 61 63 4.29259 $w=2.7e-07 $l=9.5e-08 $layer=LI1_cond $X=9.285 $Y=1.29
+ $X2=9.285 $Y2=1.385
r234 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.67
+ $Y=1.145 $X2=6.67 $Y2=1.145
r235 53 72 46.6452 $w=3.1e-07 $l=3e-07 $layer=POLY_cond $X=6.085 $Y=2.217
+ $X2=6.385 $Y2=2.217
r236 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.085
+ $Y=2.135 $X2=6.085 $Y2=2.135
r237 50 52 5.47436 $w=3.9e-07 $l=1.75e-07 $layer=LI1_cond $X=5.91 $Y=2.06
+ $X2=6.085 $Y2=2.06
r238 48 61 3.44395 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=9.46 $Y=1.29
+ $X2=9.285 $Y2=1.29
r239 47 65 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.275 $Y=1.29
+ $X2=10.44 $Y2=1.29
r240 47 48 53.1711 $w=1.68e-07 $l=8.15e-07 $layer=LI1_cond $X=10.275 $Y=1.29
+ $X2=9.46 $Y2=1.29
r241 45 61 12.2 $w=2.7e-07 $l=3.46627e-07 $layer=LI1_cond $X=9.11 $Y=1.02
+ $X2=9.285 $Y2=1.29
r242 45 46 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.11 $Y=1.02
+ $X2=8.44 $Y2=1.02
r243 44 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.355 $Y=0.935
+ $X2=8.44 $Y2=1.02
r244 43 44 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=8.355 $Y=0.425
+ $X2=8.355 $Y2=0.935
r245 41 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.27 $Y=0.34
+ $X2=8.355 $Y2=0.425
r246 41 42 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=8.27 $Y=0.34
+ $X2=7.76 $Y2=0.34
r247 39 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.675 $Y=0.425
+ $X2=7.76 $Y2=0.34
r248 39 40 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=7.675 $Y=0.425
+ $X2=7.675 $Y2=0.935
r249 37 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.59 $Y=1.02
+ $X2=7.675 $Y2=0.935
r250 37 59 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=7.59 $Y=1.02
+ $X2=6.96 $Y2=1.02
r251 36 59 6.09592 $w=3.73e-07 $l=8.5e-08 $layer=LI1_cond $X=6.875 $Y=1.122
+ $X2=6.96 $Y2=1.122
r252 36 55 6.30002 $w=3.73e-07 $l=2.05e-07 $layer=LI1_cond $X=6.875 $Y=1.122
+ $X2=6.67 $Y2=1.122
r253 35 36 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=6.875 $Y=0.425
+ $X2=6.875 $Y2=0.935
r254 34 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.995 $Y=0.34
+ $X2=5.91 $Y2=0.34
r255 33 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.79 $Y=0.34
+ $X2=6.875 $Y2=0.425
r256 33 34 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=6.79 $Y=0.34
+ $X2=5.995 $Y2=0.34
r257 32 50 5.6248 $w=1.7e-07 $l=2.4e-07 $layer=LI1_cond $X=5.91 $Y=1.82 $X2=5.91
+ $Y2=2.06
r258 31 49 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.91 $Y=0.425
+ $X2=5.91 $Y2=0.34
r259 31 32 91.0107 $w=1.68e-07 $l=1.395e-06 $layer=LI1_cond $X=5.91 $Y=0.425
+ $X2=5.91 $Y2=1.82
r260 27 50 3.08808 $w=3.9e-07 $l=1.18427e-07 $layer=LI1_cond $X=5.825 $Y=1.98
+ $X2=5.91 $Y2=2.06
r261 27 29 6.84263 $w=3.18e-07 $l=1.9e-07 $layer=LI1_cond $X=5.825 $Y=1.98
+ $X2=5.635 $Y2=1.98
r262 25 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.825 $Y=0.34
+ $X2=5.91 $Y2=0.34
r263 25 26 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=5.825 $Y=0.34
+ $X2=5.095 $Y2=0.34
r264 21 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.93 $Y=0.425
+ $X2=5.095 $Y2=0.34
r265 21 23 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=4.93 $Y=0.425
+ $X2=4.93 $Y2=0.515
r266 18 20 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=10.365 $Y=2.435
+ $X2=10.365 $Y2=2.72
r267 17 18 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=10.365 $Y=2.345
+ $X2=10.365 $Y2=2.435
r268 17 80 295.419 $w=1.8e-07 $l=7.6e-07 $layer=POLY_cond $X=10.365 $Y=2.345
+ $X2=10.365 $Y2=1.585
r269 15 76 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=9.4 $Y=0.74 $X2=9.4
+ $Y2=1.22
r270 10 56 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.67 $Y=0.98
+ $X2=6.67 $Y2=1.145
r271 10 12 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.67 $Y=0.98
+ $X2=6.67 $Y2=0.66
r272 7 72 19.7411 $w=1.5e-07 $l=2.48e-07 $layer=POLY_cond $X=6.385 $Y=2.465
+ $X2=6.385 $Y2=2.217
r273 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.385 $Y=2.465
+ $X2=6.385 $Y2=2.75
r274 2 29 600 $w=1.7e-07 $l=2.43721e-07 $layer=licon1_PDIFF $count=1 $X=5.485
+ $Y=1.84 $X2=5.635 $Y2=2.02
r275 1 23 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.79
+ $Y=0.37 $X2=4.93 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__EDFXTP_1%A_763_74# 1 2 11 13 15 17 20 22 23 25 26 28
+ 29 31 34 40 43 44 48 49 51 54 55 57 63 68
c186 57 0 1.6161e-19 $X=6.875 $Y=2.165
c187 49 0 5.61815e-20 $X=4.735 $Y=1.635
r188 63 64 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.9
+ $Y=1.635 $X2=9.9 $Y2=1.635
r189 60 63 11.399 $w=1.78e-07 $l=1.85e-07 $layer=LI1_cond $X=9.715 $Y=1.635
+ $X2=9.9 $Y2=1.635
r190 57 58 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.875
+ $Y=2.165 $X2=6.875 $Y2=2.165
r191 53 60 1.06262 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=9.715 $Y=1.725
+ $X2=9.715 $Y2=1.635
r192 53 54 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=9.715 $Y=1.725
+ $X2=9.715 $Y2=2.41
r193 52 57 14.482 $w=2.78e-07 $l=4.10244e-07 $layer=LI1_cond $X=7.115 $Y=2.495
+ $X2=6.935 $Y2=2.165
r194 51 54 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.63 $Y=2.495
+ $X2=9.715 $Y2=2.41
r195 51 52 164.08 $w=1.68e-07 $l=2.515e-06 $layer=LI1_cond $X=9.63 $Y=2.495
+ $X2=7.115 $Y2=2.495
r196 49 68 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=4.735 $Y=1.635
+ $X2=4.735 $Y2=1.655
r197 49 67 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.735 $Y=1.635
+ $X2=4.735 $Y2=1.47
r198 48 49 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.735
+ $Y=1.635 $X2=4.735 $Y2=1.635
r199 46 48 8.03336 $w=6.68e-07 $l=4.5e-07 $layer=LI1_cond $X=4.285 $Y=1.805
+ $X2=4.735 $Y2=1.805
r200 44 46 2.94557 $w=6.68e-07 $l=1.65e-07 $layer=LI1_cond $X=4.12 $Y=1.805
+ $X2=4.285 $Y2=1.805
r201 43 44 10.5816 $w=6.7e-07 $l=3.751e-07 $layer=LI1_cond $X=4.035 $Y=1.47
+ $X2=4.12 $Y2=1.805
r202 43 55 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=4.035 $Y=1.47
+ $X2=4.035 $Y2=1.01
r203 38 55 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.955 $Y=0.845
+ $X2=3.955 $Y2=1.01
r204 38 40 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=3.955 $Y=0.845
+ $X2=3.955 $Y2=0.515
r205 36 37 87.2331 $w=1.63e-07 $l=2.95e-07 $layer=POLY_cond $X=5.41 $Y=1.672
+ $X2=5.705 $Y2=1.672
r206 32 64 38.5562 $w=2.99e-07 $l=1.69926e-07 $layer=POLY_cond $X=9.91 $Y=1.47
+ $X2=9.9 $Y2=1.635
r207 32 34 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=9.91 $Y=1.47
+ $X2=9.91 $Y2=0.58
r208 29 64 52.2586 $w=2.99e-07 $l=2.82843e-07 $layer=POLY_cond $X=9.83 $Y=1.885
+ $X2=9.9 $Y2=1.635
r209 29 31 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=9.83 $Y=1.885
+ $X2=9.83 $Y2=2.46
r210 26 58 59.9436 $w=3.04e-07 $l=3.13209e-07 $layer=POLY_cond $X=6.835 $Y=2.465
+ $X2=6.862 $Y2=2.165
r211 26 28 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.835 $Y=2.465
+ $X2=6.835 $Y2=2.75
r212 25 58 38.539 $w=3.04e-07 $l=2.09893e-07 $layer=POLY_cond $X=6.76 $Y=2
+ $X2=6.862 $Y2=2.165
r213 24 25 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=6.76 $Y=1.73
+ $X2=6.76 $Y2=2
r214 23 37 22.5683 $w=1.63e-07 $l=8.30662e-08 $layer=POLY_cond $X=5.78 $Y=1.655
+ $X2=5.705 $Y2=1.672
r215 22 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.685 $Y=1.655
+ $X2=6.76 $Y2=1.73
r216 22 23 464.053 $w=1.5e-07 $l=9.05e-07 $layer=POLY_cond $X=6.685 $Y=1.655
+ $X2=5.78 $Y2=1.655
r217 18 37 4.81329 $w=1.5e-07 $l=9.2e-08 $layer=POLY_cond $X=5.705 $Y=1.58
+ $X2=5.705 $Y2=1.672
r218 18 20 471.745 $w=1.5e-07 $l=9.2e-07 $layer=POLY_cond $X=5.705 $Y=1.58
+ $X2=5.705 $Y2=0.66
r219 15 36 4.81329 $w=1.5e-07 $l=9.3e-08 $layer=POLY_cond $X=5.41 $Y=1.765
+ $X2=5.41 $Y2=1.672
r220 15 17 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.41 $Y=1.765
+ $X2=5.41 $Y2=2.4
r221 14 68 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.9 $Y=1.655
+ $X2=4.735 $Y2=1.655
r222 13 36 27.0038 $w=1.63e-07 $l=9.81326e-08 $layer=POLY_cond $X=5.32 $Y=1.655
+ $X2=5.41 $Y2=1.672
r223 13 14 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=5.32 $Y=1.655
+ $X2=4.9 $Y2=1.655
r224 11 67 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=4.715 $Y=0.74
+ $X2=4.715 $Y2=1.47
r225 2 46 600 $w=1.7e-07 $l=2.43721e-07 $layer=licon1_PDIFF $count=1 $X=4.135
+ $Y=1.76 $X2=4.285 $Y2=1.94
r226 1 40 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.815
+ $Y=0.37 $X2=3.955 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__EDFXTP_1%A_1409_64# 1 2 9 12 13 15 17 18 20 23 25 26
+ 27 31 33 38 39 41 48 56
c104 48 0 2.74064e-19 $X=7.46 $Y=1.367
c105 12 0 1.96559e-19 $X=7.34 $Y=2.375
r106 49 50 18.6009 $w=2.23e-07 $l=3.4e-07 $layer=LI1_cond $X=8.015 $Y=1.44
+ $X2=8.355 $Y2=1.44
r107 46 56 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=7.295 $Y=1.365
+ $X2=7.34 $Y2=1.365
r108 46 53 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=7.295 $Y=1.365
+ $X2=7.12 $Y2=1.365
r109 45 48 9.98442 $w=1.83e-07 $l=1.65e-07 $layer=LI1_cond $X=7.295 $Y=1.367
+ $X2=7.46 $Y2=1.367
r110 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.295
+ $Y=1.365 $X2=7.295 $Y2=1.365
r111 41 42 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.775
+ $Y=1.44 $X2=8.775 $Y2=1.44
r112 39 50 4.43115 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.44 $Y=1.44
+ $X2=8.355 $Y2=1.44
r113 39 41 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=8.44 $Y=1.44
+ $X2=8.775 $Y2=1.44
r114 37 50 2.32876 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.355 $Y=1.605
+ $X2=8.355 $Y2=1.44
r115 37 38 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=8.355 $Y=1.605
+ $X2=8.355 $Y2=2.07
r116 33 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.27 $Y=2.155
+ $X2=8.355 $Y2=2.07
r117 33 35 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=8.27 $Y=2.155
+ $X2=8.11 $Y2=2.155
r118 29 49 2.32876 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.015 $Y=1.275
+ $X2=8.015 $Y2=1.44
r119 29 31 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=8.015 $Y=1.275
+ $X2=8.015 $Y2=0.85
r120 27 49 5.36928 $w=2.23e-07 $l=1.18427e-07 $layer=LI1_cond $X=7.93 $Y=1.36
+ $X2=8.015 $Y2=1.44
r121 27 48 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=7.93 $Y=1.36
+ $X2=7.46 $Y2=1.36
r122 25 42 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=8.805 $Y=1.44
+ $X2=8.775 $Y2=1.44
r123 25 26 3.90195 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=8.805 $Y=1.44
+ $X2=8.895 $Y2=1.44
r124 21 26 34.7346 $w=1.65e-07 $l=1.72337e-07 $layer=POLY_cond $X=8.91 $Y=1.275
+ $X2=8.895 $Y2=1.44
r125 21 23 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=8.91 $Y=1.275
+ $X2=8.91 $Y2=0.74
r126 18 20 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=8.895 $Y=1.885
+ $X2=8.895 $Y2=2.46
r127 17 18 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=8.895 $Y=1.795
+ $X2=8.895 $Y2=1.885
r128 16 26 34.7346 $w=1.65e-07 $l=1.65e-07 $layer=POLY_cond $X=8.895 $Y=1.605
+ $X2=8.895 $Y2=1.44
r129 16 17 73.8548 $w=1.8e-07 $l=1.9e-07 $layer=POLY_cond $X=8.895 $Y=1.605
+ $X2=8.895 $Y2=1.795
r130 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.34 $Y=2.465
+ $X2=7.34 $Y2=2.75
r131 12 13 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=7.34 $Y=2.375
+ $X2=7.34 $Y2=2.465
r132 11 56 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.34 $Y=1.53
+ $X2=7.34 $Y2=1.365
r133 11 12 328.46 $w=1.8e-07 $l=8.45e-07 $layer=POLY_cond $X=7.34 $Y=1.53
+ $X2=7.34 $Y2=2.375
r134 7 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.12 $Y=1.2
+ $X2=7.12 $Y2=1.365
r135 7 9 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=7.12 $Y=1.2 $X2=7.12
+ $Y2=0.66
r136 2 35 600 $w=1.7e-07 $l=2.04939e-07 $layer=licon1_PDIFF $count=1 $X=7.96
+ $Y=2.025 $X2=8.11 $Y2=2.155
r137 1 31 182 $w=1.7e-07 $l=4.64758e-07 $layer=licon1_NDIFF $count=1 $X=7.875
+ $Y=0.45 $X2=8.015 $Y2=0.85
.ends

.subckt PM_SKY130_FD_SC_LS__EDFXTP_1%A_1156_90# 1 2 9 11 13 15 16 22 27 28 31 33
c93 9 0 2.85555e-19 $X=7.8 $Y=0.77
r94 31 33 9.38152 $w=2.13e-07 $l=1.65e-07 $layer=LI1_cond $X=7.865 $Y=1.722
+ $X2=7.7 $Y2=1.722
r95 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.865
+ $Y=1.7 $X2=7.865 $Y2=1.7
r96 27 28 10.5918 $w=3.58e-07 $l=2.3e-07 $layer=LI1_cond $X=6.595 $Y=2.75
+ $X2=6.595 $Y2=2.52
r97 23 25 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=6.25 $Y=1.715
+ $X2=6.5 $Y2=1.715
r98 22 25 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=6.585 $Y=1.715
+ $X2=6.5 $Y2=1.715
r99 22 33 72.7433 $w=1.68e-07 $l=1.115e-06 $layer=LI1_cond $X=6.585 $Y=1.715
+ $X2=7.7 $Y2=1.715
r100 19 25 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.5 $Y=1.8 $X2=6.5
+ $Y2=1.715
r101 19 28 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=6.5 $Y=1.8 $X2=6.5
+ $Y2=2.52
r102 16 18 3.94706 $w=1.7e-07 $l=5.5e-08 $layer=LI1_cond $X=6.335 $Y=0.68
+ $X2=6.39 $Y2=0.68
r103 15 23 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.25 $Y=1.63
+ $X2=6.25 $Y2=1.715
r104 14 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.25 $Y=0.765
+ $X2=6.335 $Y2=0.68
r105 14 15 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=6.25 $Y=0.765
+ $X2=6.25 $Y2=1.63
r106 11 32 52.2586 $w=2.99e-07 $l=2.59808e-07 $layer=POLY_cond $X=7.885 $Y=1.95
+ $X2=7.865 $Y2=1.7
r107 11 13 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=7.885 $Y=1.95
+ $X2=7.885 $Y2=2.445
r108 7 32 38.5562 $w=2.99e-07 $l=1.94808e-07 $layer=POLY_cond $X=7.8 $Y=1.535
+ $X2=7.865 $Y2=1.7
r109 7 9 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=7.8 $Y=1.535 $X2=7.8
+ $Y2=0.77
r110 2 27 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=6.46
+ $Y=2.54 $X2=6.61 $Y2=2.75
r111 1 18 182 $w=1.7e-07 $l=7.15821e-07 $layer=licon1_NDIFF $count=1 $X=5.78
+ $Y=0.45 $X2=6.39 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_LS__EDFXTP_1%A_1895_74# 1 2 9 12 13 15 16 18 20 22 23 25
+ 26 29 31 32 35 39 40 42 45 46 49
c137 32 0 1.36277e-19 $X=9.78 $Y=0.92
r138 52 53 27.9638 $w=4.1e-07 $l=7.5e-08 $layer=POLY_cond $X=11.38 $Y=1.26
+ $X2=11.38 $Y2=1.335
r139 46 52 12.2083 $w=4.1e-07 $l=9e-08 $layer=POLY_cond $X=11.38 $Y=1.17
+ $X2=11.38 $Y2=1.26
r140 46 51 45.9078 $w=4.1e-07 $l=1.65e-07 $layer=POLY_cond $X=11.38 $Y=1.17
+ $X2=11.38 $Y2=1.005
r141 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.34
+ $Y=1.17 $X2=11.34 $Y2=1.17
r142 43 49 3.70735 $w=2.5e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.945 $Y=1.17
+ $X2=10.86 $Y2=1.085
r143 43 45 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=10.945 $Y=1.17
+ $X2=11.34 $Y2=1.17
r144 41 49 2.76166 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=10.86 $Y=1.335
+ $X2=10.86 $Y2=1.085
r145 41 42 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=10.86 $Y=1.335
+ $X2=10.86 $Y2=1.755
r146 40 48 16.9994 $w=2.36e-07 $l=3.49929e-07 $layer=LI1_cond $X=10.405 $Y=1.84
+ $X2=10.095 $Y2=1.925
r147 39 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.775 $Y=1.84
+ $X2=10.86 $Y2=1.755
r148 39 40 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=10.775 $Y=1.84
+ $X2=10.405 $Y2=1.84
r149 35 37 33.6513 $w=2.48e-07 $l=7.3e-07 $layer=LI1_cond $X=10.095 $Y=2.105
+ $X2=10.095 $Y2=2.835
r150 33 48 0.361987 $w=2.5e-07 $l=1.7e-07 $layer=LI1_cond $X=10.095 $Y=2.095
+ $X2=10.095 $Y2=1.925
r151 33 35 0.460977 $w=2.48e-07 $l=1e-08 $layer=LI1_cond $X=10.095 $Y=2.095
+ $X2=10.095 $Y2=2.105
r152 31 49 3.70735 $w=2.5e-07 $l=2.03101e-07 $layer=LI1_cond $X=10.775 $Y=0.92
+ $X2=10.86 $Y2=1.085
r153 31 32 64.9144 $w=1.68e-07 $l=9.95e-07 $layer=LI1_cond $X=10.775 $Y=0.92
+ $X2=9.78 $Y2=0.92
r154 27 32 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.615 $Y=0.835
+ $X2=9.78 $Y2=0.92
r155 27 29 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=9.615 $Y=0.835
+ $X2=9.615 $Y2=0.515
r156 23 25 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=12.465 $Y=1.765
+ $X2=12.465 $Y2=2.4
r157 22 23 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=12.465 $Y=1.675
+ $X2=12.465 $Y2=1.765
r158 21 26 18.8402 $w=1.65e-07 $l=8.7892e-08 $layer=POLY_cond $X=12.465 $Y=1.335
+ $X2=12.437 $Y2=1.26
r159 21 22 132.161 $w=1.8e-07 $l=3.4e-07 $layer=POLY_cond $X=12.465 $Y=1.335
+ $X2=12.465 $Y2=1.675
r160 18 26 18.8402 $w=1.65e-07 $l=9.3675e-08 $layer=POLY_cond $X=12.395 $Y=1.185
+ $X2=12.437 $Y2=1.26
r161 18 20 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=12.395 $Y=1.185
+ $X2=12.395 $Y2=0.74
r162 17 52 26.4667 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=11.585 $Y=1.26
+ $X2=11.38 $Y2=1.26
r163 16 26 6.66866 $w=1.5e-07 $l=1.17e-07 $layer=POLY_cond $X=12.32 $Y=1.26
+ $X2=12.437 $Y2=1.26
r164 16 17 376.883 $w=1.5e-07 $l=7.35e-07 $layer=POLY_cond $X=12.32 $Y=1.26
+ $X2=11.585 $Y2=1.26
r165 13 15 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=11.495 $Y=2.215
+ $X2=11.495 $Y2=2.61
r166 12 13 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=11.495 $Y=2.125
+ $X2=11.495 $Y2=2.215
r167 12 53 307.081 $w=1.8e-07 $l=7.9e-07 $layer=POLY_cond $X=11.495 $Y=2.125
+ $X2=11.495 $Y2=1.335
r168 9 51 217.926 $w=1.5e-07 $l=4.25e-07 $layer=POLY_cond $X=11.405 $Y=0.58
+ $X2=11.405 $Y2=1.005
r169 2 37 600 $w=1.7e-07 $l=9.47035e-07 $layer=licon1_PDIFF $count=1 $X=9.905
+ $Y=1.96 $X2=10.055 $Y2=2.835
r170 2 35 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=9.905
+ $Y=1.96 $X2=10.055 $Y2=2.105
r171 1 29 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.475
+ $Y=0.37 $X2=9.615 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__EDFXTP_1%A_27_508# 1 2 3 4 5 6 20 23 25 28 29 30 32
+ 33 34 36 37 40 41 43 45 46 49 54 56 60 64
c178 64 0 1.4577e-19 $X=3.31 $Y=2.39
c179 43 0 5.61815e-20 $X=5.49 $Y=0.7
c180 34 0 3.01092e-20 $X=2.215 $Y=2.035
r181 64 65 0.189441 $w=3.22e-07 $l=5e-09 $layer=LI1_cond $X=3.287 $Y=2.39
+ $X2=3.287 $Y2=2.395
r182 58 60 5.98039 $w=4.58e-07 $l=2.3e-07 $layer=LI1_cond $X=2.955 $Y=0.645
+ $X2=3.185 $Y2=0.645
r183 51 54 4.96245 $w=4.68e-07 $l=1.95e-07 $layer=LI1_cond $X=0.17 $Y=0.575
+ $X2=0.365 $Y2=0.575
r184 47 49 2.76586 $w=2.48e-07 $l=6e-08 $layer=LI1_cond $X=6.12 $Y=2.69 $X2=6.12
+ $Y2=2.75
r185 46 70 20.8849 $w=2.44e-07 $l=4.53211e-07 $layer=LI1_cond $X=5.61 $Y=2.605
+ $X2=5.215 $Y2=2.48
r186 45 47 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.995 $Y=2.605
+ $X2=6.12 $Y2=2.69
r187 45 46 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=5.995 $Y=2.605
+ $X2=5.61 $Y2=2.605
r188 41 66 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=5.49 $Y=1.565
+ $X2=5.215 $Y2=1.565
r189 41 43 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=5.49 $Y=1.48
+ $X2=5.49 $Y2=0.7
r190 40 70 2.85362 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=5.215 $Y=2.31
+ $X2=5.215 $Y2=2.48
r191 39 66 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.215 $Y=1.65
+ $X2=5.215 $Y2=1.565
r192 39 40 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=5.215 $Y=1.65
+ $X2=5.215 $Y2=2.31
r193 38 65 4.47834 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=3.475 $Y=2.395
+ $X2=3.287 $Y2=2.395
r194 37 70 5.3849 $w=2.44e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.13 $Y=2.395
+ $X2=5.215 $Y2=2.48
r195 37 38 107.973 $w=1.68e-07 $l=1.655e-06 $layer=LI1_cond $X=5.13 $Y=2.395
+ $X2=3.475 $Y2=2.395
r196 35 60 6.6364 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=3.185 $Y=0.875
+ $X2=3.185 $Y2=0.645
r197 35 36 70.1337 $w=1.68e-07 $l=1.075e-06 $layer=LI1_cond $X=3.185 $Y=0.875
+ $X2=3.185 $Y2=1.95
r198 33 64 13.4503 $w=3.22e-07 $l=4.38646e-07 $layer=LI1_cond $X=3.1 $Y=2.035
+ $X2=3.287 $Y2=2.39
r199 33 36 5.92483 $w=3.22e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.1 $Y=2.035
+ $X2=3.185 $Y2=1.95
r200 33 34 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=3.1 $Y=2.035
+ $X2=2.215 $Y2=2.035
r201 31 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.13 $Y=2.12
+ $X2=2.215 $Y2=2.035
r202 31 32 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=2.13 $Y=2.12
+ $X2=2.13 $Y2=2.905
r203 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.045 $Y=2.99
+ $X2=2.13 $Y2=2.905
r204 29 30 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=2.045 $Y=2.99
+ $X2=1.535 $Y2=2.99
r205 28 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.45 $Y=2.905
+ $X2=1.535 $Y2=2.99
r206 27 28 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=1.45 $Y=2.35
+ $X2=1.45 $Y2=2.905
r207 26 56 2.90867 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=0.435 $Y=2.265
+ $X2=0.26 $Y2=2.265
r208 25 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.365 $Y=2.265
+ $X2=1.45 $Y2=2.35
r209 25 26 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=1.365 $Y=2.265
+ $X2=0.435 $Y2=2.265
r210 21 56 3.58051 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=2.35
+ $X2=0.26 $Y2=2.265
r211 21 23 13.1708 $w=3.48e-07 $l=4e-07 $layer=LI1_cond $X=0.26 $Y=2.35 $X2=0.26
+ $Y2=2.75
r212 20 56 3.58051 $w=2.6e-07 $l=1.25499e-07 $layer=LI1_cond $X=0.17 $Y=2.18
+ $X2=0.26 $Y2=2.265
r213 19 51 6.76998 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=0.17 $Y=0.81
+ $X2=0.17 $Y2=0.575
r214 19 20 89.3797 $w=1.68e-07 $l=1.37e-06 $layer=LI1_cond $X=0.17 $Y=0.81
+ $X2=0.17 $Y2=2.18
r215 6 49 600 $w=1.7e-07 $l=2.67208e-07 $layer=licon1_PDIFF $count=1 $X=6.03
+ $Y=2.54 $X2=6.16 $Y2=2.75
r216 5 64 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=3.16
+ $Y=2.18 $X2=3.31 $Y2=2.39
r217 4 23 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.54 $X2=0.27 $Y2=2.75
r218 3 43 182 $w=1.7e-07 $l=3.14245e-07 $layer=licon1_NDIFF $count=1 $X=5.345
+ $Y=0.45 $X2=5.49 $Y2=0.7
r219 2 58 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.815
+ $Y=0.435 $X2=2.955 $Y2=0.645
r220 1 54 182 $w=1.7e-07 $l=2.67862e-07 $layer=licon1_NDIFF $count=1 $X=0.22
+ $Y=0.37 $X2=0.365 $Y2=0.575
.ends

.subckt PM_SKY130_FD_SC_LS__EDFXTP_1%VPWR 1 2 3 4 5 6 7 8 27 31 35 39 43 47 51
+ 53 55 60 61 63 64 66 67 69 70 71 89 93 102 109 115 118 121 125
r135 124 125 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r136 121 122 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r137 118 119 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r138 115 116 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r139 113 125 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=12.72 $Y2=3.33
r140 113 122 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=11.28 $Y2=3.33
r141 112 113 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r142 110 121 11.8214 $w=1.7e-07 $l=2.7e-07 $layer=LI1_cond $X=11.385 $Y=3.33
+ $X2=11.115 $Y2=3.33
r143 110 112 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=11.385 $Y=3.33
+ $X2=12.24 $Y2=3.33
r144 109 124 4.02656 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=12.605 $Y=3.33
+ $X2=12.782 $Y2=3.33
r145 109 112 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=12.605 $Y=3.33
+ $X2=12.24 $Y2=3.33
r146 108 122 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=11.28 $Y2=3.33
r147 107 108 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r148 105 108 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=10.8 $Y2=3.33
r149 104 107 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=8.88 $Y=3.33
+ $X2=10.8 $Y2=3.33
r150 104 105 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r151 102 121 11.8214 $w=1.7e-07 $l=2.7e-07 $layer=LI1_cond $X=10.845 $Y=3.33
+ $X2=11.115 $Y2=3.33
r152 102 107 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=10.845 $Y=3.33
+ $X2=10.8 $Y2=3.33
r153 101 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=8.88 $Y2=3.33
r154 101 119 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=7.44 $Y2=3.33
r155 100 101 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r156 98 118 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.74 $Y=3.33
+ $X2=7.575 $Y2=3.33
r157 98 100 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=7.74 $Y=3.33
+ $X2=8.4 $Y2=3.33
r158 97 116 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=5.04 $Y2=3.33
r159 96 97 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r160 94 115 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.27 $Y=3.33
+ $X2=5.145 $Y2=3.33
r161 94 96 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=5.27 $Y=3.33
+ $X2=5.52 $Y2=3.33
r162 93 118 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.41 $Y=3.33
+ $X2=7.575 $Y2=3.33
r163 93 96 123.305 $w=1.68e-07 $l=1.89e-06 $layer=LI1_cond $X=7.41 $Y=3.33
+ $X2=5.52 $Y2=3.33
r164 92 116 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r165 91 92 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r166 89 115 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.02 $Y=3.33
+ $X2=5.145 $Y2=3.33
r167 89 91 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=5.02 $Y=3.33
+ $X2=4.08 $Y2=3.33
r168 88 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r169 87 88 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r170 85 88 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r171 84 87 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.64 $Y=3.33 $X2=3.6
+ $Y2=3.33
r172 84 85 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r173 82 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r174 81 82 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r175 79 82 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r176 78 81 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r177 78 79 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r178 75 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r179 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r180 71 119 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=7.44 $Y2=3.33
r181 71 97 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=5.52 $Y2=3.33
r182 69 100 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=8.505 $Y=3.33
+ $X2=8.4 $Y2=3.33
r183 69 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.505 $Y=3.33
+ $X2=8.67 $Y2=3.33
r184 68 104 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=8.835 $Y=3.33
+ $X2=8.88 $Y2=3.33
r185 68 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.835 $Y=3.33
+ $X2=8.67 $Y2=3.33
r186 66 87 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=3.67 $Y=3.33 $X2=3.6
+ $Y2=3.33
r187 66 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.67 $Y=3.33
+ $X2=3.835 $Y2=3.33
r188 65 91 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=4 $Y=3.33 $X2=4.08
+ $Y2=3.33
r189 65 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4 $Y=3.33 $X2=3.835
+ $Y2=3.33
r190 63 81 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.385 $Y=3.33
+ $X2=2.16 $Y2=3.33
r191 63 64 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.385 $Y=3.33
+ $X2=2.51 $Y2=3.33
r192 62 84 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=2.635 $Y=3.33
+ $X2=2.64 $Y2=3.33
r193 62 64 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.635 $Y=3.33
+ $X2=2.51 $Y2=3.33
r194 60 74 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=0.72 $Y2=3.33
r195 60 61 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=1.07 $Y2=3.33
r196 59 78 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=1.195 $Y=3.33
+ $X2=1.2 $Y2=3.33
r197 59 61 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.195 $Y=3.33
+ $X2=1.07 $Y2=3.33
r198 55 58 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=12.73 $Y=1.985
+ $X2=12.73 $Y2=2.815
r199 53 124 3.1166 $w=2.5e-07 $l=1.07912e-07 $layer=LI1_cond $X=12.73 $Y=3.245
+ $X2=12.782 $Y2=3.33
r200 53 58 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=12.73 $Y=3.245
+ $X2=12.73 $Y2=2.815
r201 49 121 2.26835 $w=5.4e-07 $l=8.5e-08 $layer=LI1_cond $X=11.115 $Y=3.245
+ $X2=11.115 $Y2=3.33
r202 49 51 12.293 $w=5.38e-07 $l=5.55e-07 $layer=LI1_cond $X=11.115 $Y=3.245
+ $X2=11.115 $Y2=2.69
r203 45 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.67 $Y=3.245
+ $X2=8.67 $Y2=3.33
r204 45 47 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=8.67 $Y=3.245
+ $X2=8.67 $Y2=2.835
r205 41 118 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.575 $Y=3.245
+ $X2=7.575 $Y2=3.33
r206 41 43 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=7.575 $Y=3.245
+ $X2=7.575 $Y2=2.835
r207 37 115 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.145 $Y=3.245
+ $X2=5.145 $Y2=3.33
r208 37 39 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=5.145 $Y=3.245
+ $X2=5.145 $Y2=2.815
r209 33 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.835 $Y=3.245
+ $X2=3.835 $Y2=3.33
r210 33 35 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=3.835 $Y=3.245
+ $X2=3.835 $Y2=2.735
r211 29 64 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.51 $Y=3.245
+ $X2=2.51 $Y2=3.33
r212 29 31 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=2.51 $Y=3.245
+ $X2=2.51 $Y2=2.455
r213 25 61 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.07 $Y=3.245
+ $X2=1.07 $Y2=3.33
r214 25 27 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=1.07 $Y=3.245
+ $X2=1.07 $Y2=2.75
r215 8 58 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=12.54
+ $Y=1.84 $X2=12.69 $Y2=2.815
r216 8 55 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=12.54
+ $Y=1.84 $X2=12.69 $Y2=1.985
r217 7 51 600 $w=1.7e-07 $l=3.58887e-07 $layer=licon1_PDIFF $count=1 $X=10.86
+ $Y=2.51 $X2=11.14 $Y2=2.69
r218 6 47 600 $w=1.7e-07 $l=9.44722e-07 $layer=licon1_PDIFF $count=1 $X=8.525
+ $Y=1.96 $X2=8.67 $Y2=2.835
r219 5 43 600 $w=1.7e-07 $l=3.66367e-07 $layer=licon1_PDIFF $count=1 $X=7.415
+ $Y=2.54 $X2=7.575 $Y2=2.835
r220 4 39 600 $w=1.7e-07 $l=1.03562e-06 $layer=licon1_PDIFF $count=1 $X=5.06
+ $Y=1.84 $X2=5.185 $Y2=2.815
r221 3 35 600 $w=1.7e-07 $l=1.03797e-06 $layer=licon1_PDIFF $count=1 $X=3.705
+ $Y=1.76 $X2=3.835 $Y2=2.735
r222 2 31 600 $w=1.7e-07 $l=4.98899e-07 $layer=licon1_PDIFF $count=1 $X=2.09
+ $Y=2.18 $X2=2.47 $Y2=2.455
r223 1 27 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=0.96
+ $Y=2.54 $X2=1.11 $Y2=2.75
.ends

.subckt PM_SKY130_FD_SC_LS__EDFXTP_1%Q 1 2 9 13 14 15 16 17 35 37
r30 23 37 1.74613 $w=3.28e-07 $l=5e-08 $layer=LI1_cond $X=12.24 $Y=1.715
+ $X2=12.24 $Y2=1.665
r31 16 17 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=12.24 $Y=2.405
+ $X2=12.24 $Y2=2.775
r32 15 16 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=12.24 $Y=1.985
+ $X2=12.24 $Y2=2.405
r33 14 37 0.628605 $w=3.28e-07 $l=1.8e-08 $layer=LI1_cond $X=12.24 $Y=1.647
+ $X2=12.24 $Y2=1.665
r34 14 35 3.8025 $w=3.28e-07 $l=9.7e-08 $layer=LI1_cond $X=12.24 $Y=1.647
+ $X2=12.24 $Y2=1.55
r35 14 15 8.8354 $w=3.28e-07 $l=2.53e-07 $layer=LI1_cond $X=12.24 $Y=1.732
+ $X2=12.24 $Y2=1.985
r36 14 23 0.593683 $w=3.28e-07 $l=1.7e-08 $layer=LI1_cond $X=12.24 $Y=1.732
+ $X2=12.24 $Y2=1.715
r37 13 35 17.9269 $w=2.68e-07 $l=4.2e-07 $layer=LI1_cond $X=12.21 $Y=1.13
+ $X2=12.21 $Y2=1.55
r38 7 13 6.17723 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=12.18 $Y=0.965
+ $X2=12.18 $Y2=1.13
r39 7 9 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=12.18 $Y=0.965
+ $X2=12.18 $Y2=0.515
r40 2 17 400 $w=1.7e-07 $l=1.03562e-06 $layer=licon1_PDIFF $count=1 $X=12.115
+ $Y=1.84 $X2=12.24 $Y2=2.815
r41 2 15 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=12.115
+ $Y=1.84 $X2=12.24 $Y2=1.985
r42 1 9 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=12.035
+ $Y=0.37 $X2=12.18 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__EDFXTP_1%VGND 1 2 3 4 5 6 7 8 27 31 35 39 43 47 49
+ 51 54 55 57 58 60 61 62 64 69 78 99 105 108 111 116 122 125
c148 43 0 1.96074e-19 $X=7.335 $Y=0.595
c149 1 0 1.9799e-19 $X=1.045 $Y=0.37
r150 124 125 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r151 120 122 8.97006 $w=7.48e-07 $l=3e-08 $layer=LI1_cond $X=11.28 $Y=0.29
+ $X2=11.31 $Y2=0.29
r152 120 121 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r153 118 120 1.43529 $w=7.48e-07 $l=9e-08 $layer=LI1_cond $X=11.19 $Y=0.29
+ $X2=11.28 $Y2=0.29
r154 115 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=11.28 $Y2=0
r155 114 118 6.21961 $w=7.48e-07 $l=3.9e-07 $layer=LI1_cond $X=10.8 $Y=0.29
+ $X2=11.19 $Y2=0.29
r156 114 116 15.6681 $w=7.48e-07 $l=4.5e-07 $layer=LI1_cond $X=10.8 $Y=0.29
+ $X2=10.35 $Y2=0.29
r157 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=0
+ $X2=10.8 $Y2=0
r158 111 112 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r159 108 109 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r160 105 106 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r161 103 125 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=12.72 $Y2=0
r162 103 121 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=11.28 $Y2=0
r163 102 122 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=12.24 $Y=0
+ $X2=11.31 $Y2=0
r164 102 103 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r165 99 124 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=12.515 $Y=0
+ $X2=12.737 $Y2=0
r166 99 102 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=12.515 $Y=0
+ $X2=12.24 $Y2=0
r167 98 115 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=10.8 $Y2=0
r168 97 116 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=10.32 $Y=0 $X2=10.35
+ $Y2=0
r169 97 98 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r170 95 98 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=8.88 $Y=0
+ $X2=10.32 $Y2=0
r171 94 97 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=8.88 $Y=0
+ $X2=10.32 $Y2=0
r172 94 95 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r173 91 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=8.88
+ $Y2=0
r174 90 91 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r175 88 91 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=8.4
+ $Y2=0
r176 87 90 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=7.44 $Y=0 $X2=8.4
+ $Y2=0
r177 87 88 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r178 85 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r179 84 85 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r180 82 111 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.585 $Y=0
+ $X2=4.46 $Y2=0
r181 82 84 154.947 $w=1.68e-07 $l=2.375e-06 $layer=LI1_cond $X=4.585 $Y=0
+ $X2=6.96 $Y2=0
r182 81 112 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0
+ $X2=4.56 $Y2=0
r183 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r184 78 111 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.335 $Y=0
+ $X2=4.46 $Y2=0
r185 78 80 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=4.335 $Y=0
+ $X2=4.08 $Y2=0
r186 77 81 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r187 77 109 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0
+ $X2=2.16 $Y2=0
r188 76 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r189 74 108 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.33 $Y=0
+ $X2=2.165 $Y2=0
r190 74 76 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=2.33 $Y=0 $X2=3.12
+ $Y2=0
r191 73 109 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0
+ $X2=2.16 $Y2=0
r192 73 106 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r193 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r194 70 105 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.35 $Y=0
+ $X2=1.185 $Y2=0
r195 70 72 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.35 $Y=0 $X2=1.68
+ $Y2=0
r196 69 108 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2 $Y=0 $X2=2.165
+ $Y2=0
r197 69 72 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2 $Y=0 $X2=1.68
+ $Y2=0
r198 67 106 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r199 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r200 64 105 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.02 $Y=0
+ $X2=1.185 $Y2=0
r201 64 66 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.02 $Y=0 $X2=0.72
+ $Y2=0
r202 62 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6.96
+ $Y2=0
r203 62 112 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6.48 $Y=0
+ $X2=4.56 $Y2=0
r204 60 90 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=8.61 $Y=0 $X2=8.4
+ $Y2=0
r205 60 61 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.61 $Y=0 $X2=8.735
+ $Y2=0
r206 59 94 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=8.86 $Y=0 $X2=8.88
+ $Y2=0
r207 59 61 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.86 $Y=0 $X2=8.735
+ $Y2=0
r208 57 84 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=7.17 $Y=0 $X2=6.96
+ $Y2=0
r209 57 58 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.17 $Y=0 $X2=7.295
+ $Y2=0
r210 56 87 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=7.42 $Y=0 $X2=7.44
+ $Y2=0
r211 56 58 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.42 $Y=0 $X2=7.295
+ $Y2=0
r212 54 76 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=3.44 $Y=0 $X2=3.12
+ $Y2=0
r213 54 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.44 $Y=0 $X2=3.525
+ $Y2=0
r214 53 80 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=3.61 $Y=0 $X2=4.08
+ $Y2=0
r215 53 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.61 $Y=0 $X2=3.525
+ $Y2=0
r216 49 124 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=12.68 $Y=0.085
+ $X2=12.737 $Y2=0
r217 49 51 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=12.68 $Y=0.085
+ $X2=12.68 $Y2=0.515
r218 45 61 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.735 $Y=0.085
+ $X2=8.735 $Y2=0
r219 45 47 21.6659 $w=2.48e-07 $l=4.7e-07 $layer=LI1_cond $X=8.735 $Y=0.085
+ $X2=8.735 $Y2=0.555
r220 41 58 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.295 $Y=0.085
+ $X2=7.295 $Y2=0
r221 41 43 23.5098 $w=2.48e-07 $l=5.1e-07 $layer=LI1_cond $X=7.295 $Y=0.085
+ $X2=7.295 $Y2=0.595
r222 37 111 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.46 $Y=0.085
+ $X2=4.46 $Y2=0
r223 37 39 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=4.46 $Y=0.085
+ $X2=4.46 $Y2=0.515
r224 33 55 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.525 $Y=0.085
+ $X2=3.525 $Y2=0
r225 33 35 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=3.525 $Y=0.085
+ $X2=3.525 $Y2=0.505
r226 29 108 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.165 $Y=0.085
+ $X2=2.165 $Y2=0
r227 29 31 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=2.165 $Y=0.085
+ $X2=2.165 $Y2=0.645
r228 25 105 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=0.085
+ $X2=1.185 $Y2=0
r229 25 27 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=1.185 $Y=0.085
+ $X2=1.185 $Y2=0.515
r230 8 51 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=12.47
+ $Y=0.37 $X2=12.68 $Y2=0.515
r231 7 118 91 $w=1.7e-07 $l=8.77596e-07 $layer=licon1_NDIFF $count=2 $X=10.375
+ $Y=0.37 $X2=11.19 $Y2=0.5
r232 6 47 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=8.55
+ $Y=0.37 $X2=8.695 $Y2=0.555
r233 5 43 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=7.195
+ $Y=0.45 $X2=7.335 $Y2=0.595
r234 4 39 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.36
+ $Y=0.37 $X2=4.5 $Y2=0.515
r235 3 35 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=3.38
+ $Y=0.37 $X2=3.525 $Y2=0.505
r236 2 31 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.025
+ $Y=0.435 $X2=2.165 $Y2=0.645
r237 1 27 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1.045
+ $Y=0.37 $X2=1.185 $Y2=0.515
.ends

