* File: sky130_fd_sc_ls__nor4_4.pxi.spice
* Created: Wed Sep  2 11:15:36 2020
* 
x_PM_SKY130_FD_SC_LS__NOR4_4%D N_D_M1002_g N_D_c_105_n N_D_M1000_g N_D_c_106_n
+ N_D_M1012_g N_D_c_107_n N_D_M1013_g N_D_M1020_g N_D_c_108_n N_D_M1018_g D D D
+ N_D_c_109_n N_D_c_104_n PM_SKY130_FD_SC_LS__NOR4_4%D
x_PM_SKY130_FD_SC_LS__NOR4_4%C N_C_M1008_g N_C_c_169_n N_C_M1005_g N_C_c_170_n
+ N_C_M1011_g N_C_c_171_n N_C_M1016_g N_C_M1022_g N_C_c_172_n N_C_M1021_g C C C
+ N_C_c_167_n N_C_c_168_n PM_SKY130_FD_SC_LS__NOR4_4%C
x_PM_SKY130_FD_SC_LS__NOR4_4%B N_B_M1007_g N_B_M1015_g N_B_c_240_n N_B_M1003_g
+ N_B_c_241_n N_B_M1004_g N_B_c_242_n N_B_M1006_g N_B_c_243_n N_B_M1023_g B B B
+ B B B N_B_c_239_n PM_SKY130_FD_SC_LS__NOR4_4%B
x_PM_SKY130_FD_SC_LS__NOR4_4%A N_A_c_320_n N_A_M1001_g N_A_c_312_n N_A_M1010_g
+ N_A_c_321_n N_A_M1009_g N_A_c_322_n N_A_M1014_g N_A_M1017_g N_A_c_323_n
+ N_A_M1019_g N_A_c_315_n A A N_A_c_317_n N_A_c_318_n N_A_c_319_n
+ PM_SKY130_FD_SC_LS__NOR4_4%A
x_PM_SKY130_FD_SC_LS__NOR4_4%A_27_368# N_A_27_368#_M1000_d N_A_27_368#_M1012_d
+ N_A_27_368#_M1018_d N_A_27_368#_M1011_s N_A_27_368#_M1021_s
+ N_A_27_368#_c_386_n N_A_27_368#_c_387_n N_A_27_368#_c_388_n
+ N_A_27_368#_c_395_n N_A_27_368#_c_389_n N_A_27_368#_c_390_n
+ N_A_27_368#_c_400_n N_A_27_368#_c_405_n N_A_27_368#_c_437_p
+ N_A_27_368#_c_409_n N_A_27_368#_c_391_n N_A_27_368#_c_413_n
+ N_A_27_368#_c_392_n PM_SKY130_FD_SC_LS__NOR4_4%A_27_368#
x_PM_SKY130_FD_SC_LS__NOR4_4%Y N_Y_M1002_s N_Y_M1008_s N_Y_M1007_d N_Y_M1010_d
+ N_Y_M1000_s N_Y_M1013_s N_Y_c_453_n N_Y_c_466_n N_Y_c_464_n N_Y_c_468_n
+ N_Y_c_454_n N_Y_c_455_n N_Y_c_456_n N_Y_c_457_n N_Y_c_458_n N_Y_c_477_n
+ N_Y_c_482_n N_Y_c_459_n N_Y_c_460_n N_Y_c_461_n N_Y_c_462_n Y
+ PM_SKY130_FD_SC_LS__NOR4_4%Y
x_PM_SKY130_FD_SC_LS__NOR4_4%A_496_368# N_A_496_368#_M1005_d
+ N_A_496_368#_M1016_d N_A_496_368#_M1003_d N_A_496_368#_M1006_d
+ N_A_496_368#_c_565_n N_A_496_368#_c_559_n N_A_496_368#_c_560_n
+ N_A_496_368#_c_572_n N_A_496_368#_c_561_n N_A_496_368#_c_579_n
+ N_A_496_368#_c_562_n N_A_496_368#_c_585_n N_A_496_368#_c_563_n
+ N_A_496_368#_c_564_n PM_SKY130_FD_SC_LS__NOR4_4%A_496_368#
x_PM_SKY130_FD_SC_LS__NOR4_4%A_879_368# N_A_879_368#_M1003_s
+ N_A_879_368#_M1004_s N_A_879_368#_M1023_s N_A_879_368#_M1009_d
+ N_A_879_368#_M1019_d N_A_879_368#_c_625_n N_A_879_368#_c_626_n
+ N_A_879_368#_c_634_n N_A_879_368#_c_680_n N_A_879_368#_c_638_n
+ N_A_879_368#_c_627_n N_A_879_368#_c_643_n N_A_879_368#_c_628_n
+ N_A_879_368#_c_657_n N_A_879_368#_c_629_n N_A_879_368#_c_630_n
+ N_A_879_368#_c_644_n N_A_879_368#_c_646_n N_A_879_368#_c_668_n
+ PM_SKY130_FD_SC_LS__NOR4_4%A_879_368#
x_PM_SKY130_FD_SC_LS__NOR4_4%VPWR N_VPWR_M1001_s N_VPWR_M1014_s N_VPWR_c_699_n
+ N_VPWR_c_700_n N_VPWR_c_701_n N_VPWR_c_702_n VPWR N_VPWR_c_703_n
+ N_VPWR_c_704_n N_VPWR_c_698_n N_VPWR_c_706_n PM_SKY130_FD_SC_LS__NOR4_4%VPWR
x_PM_SKY130_FD_SC_LS__NOR4_4%VGND N_VGND_M1002_d N_VGND_M1020_d N_VGND_M1022_d
+ N_VGND_M1015_s N_VGND_M1017_s N_VGND_c_778_n N_VGND_c_779_n N_VGND_c_780_n
+ N_VGND_c_781_n N_VGND_c_782_n N_VGND_c_783_n N_VGND_c_784_n N_VGND_c_785_n
+ N_VGND_c_786_n N_VGND_c_787_n N_VGND_c_788_n N_VGND_c_789_n VGND
+ N_VGND_c_790_n N_VGND_c_791_n N_VGND_c_792_n N_VGND_c_793_n N_VGND_c_794_n
+ PM_SKY130_FD_SC_LS__NOR4_4%VGND
cc_1 VNB N_D_M1002_g 0.0350087f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=0.74
cc_2 VNB N_D_M1020_g 0.033152f $X=-0.19 $Y=-0.245 $X2=1.86 $Y2=0.74
cc_3 VNB N_D_c_104_n 0.091975f $X=-0.19 $Y=-0.245 $X2=1.86 $Y2=1.557
cc_4 VNB N_C_M1008_g 0.0340976f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=0.74
cc_5 VNB N_C_M1022_g 0.033152f $X=-0.19 $Y=-0.245 $X2=1.86 $Y2=0.74
cc_6 VNB N_C_c_167_n 0.0012292f $X=-0.19 $Y=-0.245 $X2=1.71 $Y2=1.515
cc_7 VNB N_C_c_168_n 0.0890911f $X=-0.19 $Y=-0.245 $X2=1.86 $Y2=1.557
cc_8 VNB N_B_M1007_g 0.0244877f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=0.74
cc_9 VNB N_B_M1015_g 0.0306733f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=2.4
cc_10 VNB B 0.00861277f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_B_c_239_n 0.120702f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_c_312_n 0.0242527f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_M1010_g 0.0318428f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.765
cc_14 VNB N_A_M1017_g 0.0293697f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=1.765
cc_15 VNB N_A_c_315_n 0.011577f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_16 VNB A 0.0325254f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.515
cc_17 VNB N_A_c_317_n 0.0949378f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.565
cc_18 VNB N_A_c_318_n 0.00425479f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.565
cc_19 VNB N_A_c_319_n 0.00386031f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_Y_c_453_n 0.00746863f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=2.4
cc_21 VNB N_Y_c_454_n 0.00675823f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.515
cc_22 VNB N_Y_c_455_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=1.71 $Y2=1.515
cc_23 VNB N_Y_c_456_n 0.0203308f $X=-0.19 $Y=-0.245 $X2=1.86 $Y2=1.557
cc_24 VNB N_Y_c_457_n 0.00374454f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.565
cc_25 VNB N_Y_c_458_n 0.0197472f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_Y_c_459_n 0.00683417f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_Y_c_460_n 0.0201517f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_Y_c_461_n 0.00230427f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_Y_c_462_n 0.00874911f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB Y 0.0240186f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VPWR_c_698_n 0.362705f $X=-0.19 $Y=-0.245 $X2=1.71 $Y2=1.557
cc_32 VNB N_VGND_c_778_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=1.86 $Y2=0.74
cc_33 VNB N_VGND_c_779_n 0.0316455f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=1.765
cc_34 VNB N_VGND_c_780_n 0.00641221f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_35 VNB N_VGND_c_781_n 0.00571437f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_782_n 0.02962f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.557
cc_37 VNB N_VGND_c_783_n 0.028454f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.557
cc_38 VNB N_VGND_c_784_n 0.0344702f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.557
cc_39 VNB N_VGND_c_785_n 0.0389478f $X=-0.19 $Y=-0.245 $X2=1.71 $Y2=1.515
cc_40 VNB N_VGND_c_786_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=1.71 $Y2=1.515
cc_41 VNB N_VGND_c_787_n 0.0110534f $X=-0.19 $Y=-0.245 $X2=1.86 $Y2=1.557
cc_42 VNB N_VGND_c_788_n 0.0252293f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=1.557
cc_43 VNB N_VGND_c_789_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.565
cc_44 VNB N_VGND_c_790_n 0.0376264f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_791_n 0.455329f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_792_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_793_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_794_n 0.0126522f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VPB N_D_c_105_n 0.0170346f $X=-0.19 $Y=1.66 $X2=0.555 $Y2=1.765
cc_50 VPB N_D_c_106_n 0.0146623f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.765
cc_51 VPB N_D_c_107_n 0.0150427f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=1.765
cc_52 VPB N_D_c_108_n 0.0152896f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=1.765
cc_53 VPB N_D_c_109_n 0.00893755f $X=-0.19 $Y=1.66 $X2=1.71 $Y2=1.515
cc_54 VPB N_D_c_104_n 0.0493687f $X=-0.19 $Y=1.66 $X2=1.86 $Y2=1.557
cc_55 VPB N_C_c_169_n 0.0154934f $X=-0.19 $Y=1.66 $X2=0.555 $Y2=1.765
cc_56 VPB N_C_c_170_n 0.014659f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.765
cc_57 VPB N_C_c_171_n 0.0146598f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=1.765
cc_58 VPB N_C_c_172_n 0.0185749f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=1.765
cc_59 VPB N_C_c_167_n 0.00839727f $X=-0.19 $Y=1.66 $X2=1.71 $Y2=1.515
cc_60 VPB N_C_c_168_n 0.0479246f $X=-0.19 $Y=1.66 $X2=1.86 $Y2=1.557
cc_61 VPB N_B_c_240_n 0.0186627f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.4
cc_62 VPB N_B_c_241_n 0.0148184f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=2.4
cc_63 VPB N_B_c_242_n 0.0148184f $X=-0.19 $Y=1.66 $X2=1.86 $Y2=0.74
cc_64 VPB N_B_c_243_n 0.0154583f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=1.765
cc_65 VPB B 0.0255745f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_B_c_239_n 0.0642716f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_A_c_320_n 0.0165692f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.35
cc_68 VPB N_A_c_321_n 0.0163482f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.4
cc_69 VPB N_A_c_322_n 0.0163482f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=2.4
cc_70 VPB N_A_c_323_n 0.0214854f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=2.4
cc_71 VPB N_A_c_315_n 0.00635608f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.58
cc_72 VPB N_A_c_317_n 0.0235052f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.565
cc_73 VPB N_A_27_368#_c_386_n 0.0237653f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=1.765
cc_74 VPB N_A_27_368#_c_387_n 0.0028338f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=2.4
cc_75 VPB N_A_27_368#_c_388_n 0.0101535f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_76 VPB N_A_27_368#_c_389_n 0.005135f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_A_27_368#_c_390_n 0.00328567f $X=-0.19 $Y=1.66 $X2=0.555 $Y2=1.557
cc_78 VPB N_A_27_368#_c_391_n 0.00171072f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 VPB N_A_27_368#_c_392_n 0.00726038f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 VPB N_Y_c_464_n 0.00707089f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_81 VPB Y 0.0129762f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 VPB N_A_496_368#_c_559_n 0.00213603f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 VPB N_A_496_368#_c_560_n 0.0021839f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=1.765
cc_84 VPB N_A_496_368#_c_561_n 0.0170892f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.58
cc_85 VPB N_A_496_368#_c_562_n 0.00446234f $X=-0.19 $Y=1.66 $X2=0.69 $Y2=1.557
cc_86 VPB N_A_496_368#_c_563_n 0.0021839f $X=-0.19 $Y=1.66 $X2=1.71 $Y2=1.515
cc_87 VPB N_A_496_368#_c_564_n 0.0021839f $X=-0.19 $Y=1.66 $X2=1.71 $Y2=1.515
cc_88 VPB N_A_879_368#_c_625_n 0.00164284f $X=-0.19 $Y=1.66 $X2=1.86 $Y2=0.74
cc_89 VPB N_A_879_368#_c_626_n 0.00558825f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=1.765
cc_90 VPB N_A_879_368#_c_627_n 0.00234561f $X=-0.19 $Y=1.66 $X2=0.69 $Y2=1.515
cc_91 VPB N_A_879_368#_c_628_n 0.00257348f $X=-0.19 $Y=1.66 $X2=1.71 $Y2=1.515
cc_92 VPB N_A_879_368#_c_629_n 0.0154085f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_A_879_368#_c_630_n 0.035396f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_699_n 0.00895818f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.4
cc_95 VPB N_VPWR_c_700_n 0.00900305f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=2.4
cc_96 VPB N_VPWR_c_701_n 0.15727f $X=-0.19 $Y=1.66 $X2=1.86 $Y2=0.74
cc_97 VPB N_VPWR_c_702_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_703_n 0.0186948f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.557
cc_99 VPB N_VPWR_c_704_n 0.0191515f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=1.557
cc_100 VPB N_VPWR_c_698_n 0.0936461f $X=-0.19 $Y=1.66 $X2=1.71 $Y2=1.557
cc_101 VPB N_VPWR_c_706_n 0.00632158f $X=-0.19 $Y=1.66 $X2=1.86 $Y2=1.557
cc_102 N_D_M1020_g N_C_M1008_g 0.0181303f $X=1.86 $Y=0.74 $X2=0 $Y2=0
cc_103 N_D_c_108_n N_C_c_169_n 0.00956654f $X=1.955 $Y=1.765 $X2=0 $Y2=0
cc_104 N_D_c_109_n N_C_c_167_n 0.0135483f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_105 N_D_c_104_n N_C_c_167_n 0.00149052f $X=1.86 $Y=1.557 $X2=0 $Y2=0
cc_106 N_D_c_109_n N_C_c_168_n 0.00156928f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_107 N_D_c_104_n N_C_c_168_n 0.031193f $X=1.86 $Y=1.557 $X2=0 $Y2=0
cc_108 N_D_c_105_n N_A_27_368#_c_387_n 0.0149468f $X=0.555 $Y=1.765 $X2=0 $Y2=0
cc_109 N_D_c_106_n N_A_27_368#_c_387_n 0.0128349f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_110 N_D_c_107_n N_A_27_368#_c_395_n 0.0074736f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_111 N_D_c_108_n N_A_27_368#_c_395_n 8.53333e-19 $X=1.955 $Y=1.765 $X2=0 $Y2=0
cc_112 N_D_c_107_n N_A_27_368#_c_389_n 0.0111147f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_113 N_D_c_108_n N_A_27_368#_c_389_n 0.0127772f $X=1.955 $Y=1.765 $X2=0 $Y2=0
cc_114 N_D_c_108_n N_A_27_368#_c_390_n 0.00336699f $X=1.955 $Y=1.765 $X2=0 $Y2=0
cc_115 N_D_c_108_n N_A_27_368#_c_400_n 0.00544145f $X=1.955 $Y=1.765 $X2=0 $Y2=0
cc_116 N_D_c_107_n N_A_27_368#_c_391_n 0.00175197f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_117 N_D_c_105_n N_Y_c_466_n 0.01477f $X=0.555 $Y=1.765 $X2=0 $Y2=0
cc_118 N_D_c_109_n N_Y_c_466_n 0.0065328f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_119 N_D_c_106_n N_Y_c_468_n 0.0120074f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_120 N_D_c_107_n N_Y_c_468_n 0.0151589f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_121 N_D_c_109_n N_Y_c_468_n 0.0420325f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_122 N_D_c_104_n N_Y_c_468_n 0.00132059f $X=1.86 $Y=1.557 $X2=0 $Y2=0
cc_123 N_D_M1002_g N_Y_c_457_n 0.0162717f $X=0.54 $Y=0.74 $X2=0 $Y2=0
cc_124 N_D_c_109_n N_Y_c_457_n 0.113145f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_125 N_D_M1002_g N_Y_c_458_n 0.00423262f $X=0.54 $Y=0.74 $X2=0 $Y2=0
cc_126 N_D_M1020_g N_Y_c_458_n 0.00160267f $X=1.86 $Y=0.74 $X2=0 $Y2=0
cc_127 N_D_c_104_n N_Y_c_458_n 0.0242986f $X=1.86 $Y=1.557 $X2=0 $Y2=0
cc_128 N_D_c_105_n N_Y_c_477_n 0.0130624f $X=0.555 $Y=1.765 $X2=0 $Y2=0
cc_129 N_D_c_106_n N_Y_c_477_n 0.00904709f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_130 N_D_c_107_n N_Y_c_477_n 4.45174e-19 $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_131 N_D_c_109_n N_Y_c_477_n 0.0237598f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_132 N_D_c_104_n N_Y_c_477_n 0.00144939f $X=1.86 $Y=1.557 $X2=0 $Y2=0
cc_133 N_D_c_108_n N_Y_c_482_n 0.00965096f $X=1.955 $Y=1.765 $X2=0 $Y2=0
cc_134 N_D_c_109_n N_Y_c_482_n 0.0240818f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_135 N_D_c_104_n N_Y_c_482_n 0.00167671f $X=1.86 $Y=1.557 $X2=0 $Y2=0
cc_136 N_D_M1020_g N_Y_c_459_n 0.0159009f $X=1.86 $Y=0.74 $X2=0 $Y2=0
cc_137 N_D_c_104_n N_Y_c_459_n 0.0037027f $X=1.86 $Y=1.557 $X2=0 $Y2=0
cc_138 N_D_M1020_g N_Y_c_460_n 6.34175e-19 $X=1.86 $Y=0.74 $X2=0 $Y2=0
cc_139 N_D_M1002_g Y 0.0176245f $X=0.54 $Y=0.74 $X2=0 $Y2=0
cc_140 N_D_c_105_n Y 0.00661889f $X=0.555 $Y=1.765 $X2=0 $Y2=0
cc_141 N_D_c_109_n Y 0.0349192f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_142 N_D_c_105_n N_VPWR_c_701_n 0.00278271f $X=0.555 $Y=1.765 $X2=0 $Y2=0
cc_143 N_D_c_106_n N_VPWR_c_701_n 0.00278271f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_144 N_D_c_107_n N_VPWR_c_701_n 0.00278257f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_145 N_D_c_108_n N_VPWR_c_701_n 0.00278271f $X=1.955 $Y=1.765 $X2=0 $Y2=0
cc_146 N_D_c_105_n N_VPWR_c_698_n 0.00357472f $X=0.555 $Y=1.765 $X2=0 $Y2=0
cc_147 N_D_c_106_n N_VPWR_c_698_n 0.00353823f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_148 N_D_c_107_n N_VPWR_c_698_n 0.00354283f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_149 N_D_c_108_n N_VPWR_c_698_n 0.00354368f $X=1.955 $Y=1.765 $X2=0 $Y2=0
cc_150 N_D_M1002_g N_VGND_c_779_n 0.00744799f $X=0.54 $Y=0.74 $X2=0 $Y2=0
cc_151 N_D_M1020_g N_VGND_c_780_n 0.0136269f $X=1.86 $Y=0.74 $X2=0 $Y2=0
cc_152 N_D_M1002_g N_VGND_c_790_n 0.00461464f $X=0.54 $Y=0.74 $X2=0 $Y2=0
cc_153 N_D_M1020_g N_VGND_c_790_n 0.00383152f $X=1.86 $Y=0.74 $X2=0 $Y2=0
cc_154 N_D_M1002_g N_VGND_c_791_n 0.00916349f $X=0.54 $Y=0.74 $X2=0 $Y2=0
cc_155 N_D_M1020_g N_VGND_c_791_n 0.00762539f $X=1.86 $Y=0.74 $X2=0 $Y2=0
cc_156 N_C_M1022_g N_B_M1007_g 0.0176979f $X=3.71 $Y=0.74 $X2=0 $Y2=0
cc_157 N_C_c_172_n B 2.76411e-19 $X=3.755 $Y=1.765 $X2=0 $Y2=0
cc_158 N_C_c_167_n B 0.0364929f $X=3.62 $Y=1.515 $X2=0 $Y2=0
cc_159 N_C_c_168_n B 0.00398976f $X=3.71 $Y=1.557 $X2=0 $Y2=0
cc_160 N_C_c_167_n N_B_c_239_n 3.01993e-19 $X=3.62 $Y=1.515 $X2=0 $Y2=0
cc_161 N_C_c_168_n N_B_c_239_n 0.0241886f $X=3.71 $Y=1.557 $X2=0 $Y2=0
cc_162 N_C_c_169_n N_A_27_368#_c_389_n 0.00124692f $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_163 N_C_c_169_n N_A_27_368#_c_390_n 0.00262483f $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_164 N_C_c_169_n N_A_27_368#_c_400_n 0.00544145f $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_165 N_C_c_169_n N_A_27_368#_c_405_n 0.0158616f $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_166 N_C_c_170_n N_A_27_368#_c_405_n 0.0126342f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_167 N_C_c_167_n N_A_27_368#_c_405_n 0.0356825f $X=3.62 $Y=1.515 $X2=0 $Y2=0
cc_168 N_C_c_168_n N_A_27_368#_c_405_n 0.00131847f $X=3.71 $Y=1.557 $X2=0 $Y2=0
cc_169 N_C_c_171_n N_A_27_368#_c_409_n 0.0126853f $X=3.305 $Y=1.765 $X2=0 $Y2=0
cc_170 N_C_c_172_n N_A_27_368#_c_409_n 0.0138931f $X=3.755 $Y=1.765 $X2=0 $Y2=0
cc_171 N_C_c_167_n N_A_27_368#_c_409_n 0.0400603f $X=3.62 $Y=1.515 $X2=0 $Y2=0
cc_172 N_C_c_168_n N_A_27_368#_c_409_n 0.00131212f $X=3.71 $Y=1.557 $X2=0 $Y2=0
cc_173 N_C_c_167_n N_A_27_368#_c_413_n 0.0179213f $X=3.62 $Y=1.515 $X2=0 $Y2=0
cc_174 N_C_c_168_n N_A_27_368#_c_413_n 0.00127084f $X=3.71 $Y=1.557 $X2=0 $Y2=0
cc_175 N_C_c_172_n N_A_27_368#_c_392_n 0.0063565f $X=3.755 $Y=1.765 $X2=0 $Y2=0
cc_176 N_C_M1022_g N_Y_c_454_n 0.0142504f $X=3.71 $Y=0.74 $X2=0 $Y2=0
cc_177 N_C_c_168_n N_Y_c_454_n 0.00198898f $X=3.71 $Y=1.557 $X2=0 $Y2=0
cc_178 N_C_M1022_g N_Y_c_455_n 4.81487e-19 $X=3.71 $Y=0.74 $X2=0 $Y2=0
cc_179 N_C_M1008_g N_Y_c_459_n 0.0133774f $X=2.36 $Y=0.74 $X2=0 $Y2=0
cc_180 N_C_M1008_g N_Y_c_460_n 0.0138796f $X=2.36 $Y=0.74 $X2=0 $Y2=0
cc_181 N_C_M1022_g N_Y_c_460_n 0.00160267f $X=3.71 $Y=0.74 $X2=0 $Y2=0
cc_182 N_C_c_167_n N_Y_c_460_n 0.113128f $X=3.62 $Y=1.515 $X2=0 $Y2=0
cc_183 N_C_c_168_n N_Y_c_460_n 0.0249971f $X=3.71 $Y=1.557 $X2=0 $Y2=0
cc_184 N_C_c_169_n N_A_496_368#_c_565_n 0.0070569f $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_185 N_C_c_170_n N_A_496_368#_c_565_n 0.00804424f $X=2.855 $Y=1.765 $X2=0
+ $Y2=0
cc_186 N_C_c_171_n N_A_496_368#_c_565_n 5.5529e-19 $X=3.305 $Y=1.765 $X2=0 $Y2=0
cc_187 N_C_c_170_n N_A_496_368#_c_559_n 0.0108414f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_188 N_C_c_171_n N_A_496_368#_c_559_n 0.0108414f $X=3.305 $Y=1.765 $X2=0 $Y2=0
cc_189 N_C_c_169_n N_A_496_368#_c_560_n 0.00323911f $X=2.405 $Y=1.765 $X2=0
+ $Y2=0
cc_190 N_C_c_170_n N_A_496_368#_c_560_n 0.00175197f $X=2.855 $Y=1.765 $X2=0
+ $Y2=0
cc_191 N_C_c_170_n N_A_496_368#_c_572_n 5.5529e-19 $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_192 N_C_c_171_n N_A_496_368#_c_572_n 0.00804424f $X=3.305 $Y=1.765 $X2=0
+ $Y2=0
cc_193 N_C_c_172_n N_A_496_368#_c_572_n 0.0127937f $X=3.755 $Y=1.765 $X2=0 $Y2=0
cc_194 N_C_c_172_n N_A_496_368#_c_561_n 0.012762f $X=3.755 $Y=1.765 $X2=0 $Y2=0
cc_195 N_C_c_171_n N_A_496_368#_c_563_n 0.00175197f $X=3.305 $Y=1.765 $X2=0
+ $Y2=0
cc_196 N_C_c_172_n N_A_496_368#_c_563_n 0.00175197f $X=3.755 $Y=1.765 $X2=0
+ $Y2=0
cc_197 N_C_c_169_n N_VPWR_c_701_n 0.0044313f $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_198 N_C_c_170_n N_VPWR_c_701_n 0.00278257f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_199 N_C_c_171_n N_VPWR_c_701_n 0.00278257f $X=3.305 $Y=1.765 $X2=0 $Y2=0
cc_200 N_C_c_172_n N_VPWR_c_701_n 0.00278257f $X=3.755 $Y=1.765 $X2=0 $Y2=0
cc_201 N_C_c_169_n N_VPWR_c_698_n 0.00854206f $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_202 N_C_c_170_n N_VPWR_c_698_n 0.00353822f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_203 N_C_c_171_n N_VPWR_c_698_n 0.00353822f $X=3.305 $Y=1.765 $X2=0 $Y2=0
cc_204 N_C_c_172_n N_VPWR_c_698_n 0.00358623f $X=3.755 $Y=1.765 $X2=0 $Y2=0
cc_205 N_C_M1008_g N_VGND_c_780_n 0.00572988f $X=2.36 $Y=0.74 $X2=0 $Y2=0
cc_206 N_C_M1022_g N_VGND_c_781_n 0.0136269f $X=3.71 $Y=0.74 $X2=0 $Y2=0
cc_207 N_C_M1008_g N_VGND_c_785_n 0.00433162f $X=2.36 $Y=0.74 $X2=0 $Y2=0
cc_208 N_C_M1022_g N_VGND_c_785_n 0.00383152f $X=3.71 $Y=0.74 $X2=0 $Y2=0
cc_209 N_C_M1008_g N_VGND_c_791_n 0.00822119f $X=2.36 $Y=0.74 $X2=0 $Y2=0
cc_210 N_C_M1022_g N_VGND_c_791_n 0.00762539f $X=3.71 $Y=0.74 $X2=0 $Y2=0
cc_211 N_B_c_243_n N_A_c_320_n 0.00916697f $X=6.135 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_212 B N_A_c_320_n 0.00171095f $X=6.395 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_213 B N_A_c_315_n 0.0139806f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_214 N_B_c_239_n N_A_c_315_n 0.0135756f $X=6 $Y=1.515 $X2=0 $Y2=0
cc_215 B N_A_c_317_n 0.00157292f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_216 B N_A_c_319_n 0.0112317f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_217 B N_A_27_368#_c_392_n 0.0159469f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_218 N_B_M1007_g N_Y_c_454_n 0.0114826f $X=4.21 $Y=0.74 $X2=0 $Y2=0
cc_219 B N_Y_c_454_n 0.022854f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_220 N_B_M1007_g N_Y_c_455_n 0.00856181f $X=4.21 $Y=0.74 $X2=0 $Y2=0
cc_221 N_B_M1015_g N_Y_c_455_n 0.0132207f $X=4.64 $Y=0.74 $X2=0 $Y2=0
cc_222 N_B_M1015_g N_Y_c_456_n 0.0134377f $X=4.64 $Y=0.74 $X2=0 $Y2=0
cc_223 B N_Y_c_456_n 0.127864f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_224 N_B_c_239_n N_Y_c_456_n 0.0350022f $X=6 $Y=1.515 $X2=0 $Y2=0
cc_225 N_B_M1007_g N_Y_c_461_n 0.00257802f $X=4.21 $Y=0.74 $X2=0 $Y2=0
cc_226 N_B_M1015_g N_Y_c_461_n 0.00393109f $X=4.64 $Y=0.74 $X2=0 $Y2=0
cc_227 B N_Y_c_461_n 0.0281223f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_228 N_B_c_239_n N_Y_c_461_n 0.00232957f $X=6 $Y=1.515 $X2=0 $Y2=0
cc_229 N_B_c_240_n N_A_496_368#_c_561_n 0.012762f $X=4.765 $Y=1.765 $X2=0 $Y2=0
cc_230 N_B_c_240_n N_A_496_368#_c_579_n 0.0125645f $X=4.765 $Y=1.765 $X2=0 $Y2=0
cc_231 N_B_c_241_n N_A_496_368#_c_579_n 0.00801409f $X=5.215 $Y=1.765 $X2=0
+ $Y2=0
cc_232 N_B_c_242_n N_A_496_368#_c_579_n 5.57313e-19 $X=5.685 $Y=1.765 $X2=0
+ $Y2=0
cc_233 N_B_c_241_n N_A_496_368#_c_562_n 0.0109552f $X=5.215 $Y=1.765 $X2=0 $Y2=0
cc_234 N_B_c_242_n N_A_496_368#_c_562_n 0.0127071f $X=5.685 $Y=1.765 $X2=0 $Y2=0
cc_235 N_B_c_243_n N_A_496_368#_c_562_n 0.00399942f $X=6.135 $Y=1.765 $X2=0
+ $Y2=0
cc_236 N_B_c_241_n N_A_496_368#_c_585_n 5.57313e-19 $X=5.215 $Y=1.765 $X2=0
+ $Y2=0
cc_237 N_B_c_242_n N_A_496_368#_c_585_n 0.00801409f $X=5.685 $Y=1.765 $X2=0
+ $Y2=0
cc_238 N_B_c_243_n N_A_496_368#_c_585_n 0.00655294f $X=6.135 $Y=1.765 $X2=0
+ $Y2=0
cc_239 N_B_c_240_n N_A_496_368#_c_564_n 0.00175197f $X=4.765 $Y=1.765 $X2=0
+ $Y2=0
cc_240 N_B_c_241_n N_A_496_368#_c_564_n 0.00175197f $X=5.215 $Y=1.765 $X2=0
+ $Y2=0
cc_241 B N_A_879_368#_c_625_n 0.0221345f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_242 N_B_c_239_n N_A_879_368#_c_625_n 0.00153044f $X=6 $Y=1.515 $X2=0 $Y2=0
cc_243 N_B_c_240_n N_A_879_368#_c_626_n 0.00805015f $X=4.765 $Y=1.765 $X2=0
+ $Y2=0
cc_244 N_B_c_240_n N_A_879_368#_c_634_n 0.012691f $X=4.765 $Y=1.765 $X2=0 $Y2=0
cc_245 N_B_c_241_n N_A_879_368#_c_634_n 0.012691f $X=5.215 $Y=1.765 $X2=0 $Y2=0
cc_246 B N_A_879_368#_c_634_n 0.046814f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_247 N_B_c_239_n N_A_879_368#_c_634_n 0.00151204f $X=6 $Y=1.515 $X2=0 $Y2=0
cc_248 N_B_c_242_n N_A_879_368#_c_638_n 0.012691f $X=5.685 $Y=1.765 $X2=0 $Y2=0
cc_249 N_B_c_243_n N_A_879_368#_c_638_n 0.012691f $X=6.135 $Y=1.765 $X2=0 $Y2=0
cc_250 B N_A_879_368#_c_638_n 0.0456931f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_251 N_B_c_239_n N_A_879_368#_c_638_n 0.00132059f $X=6 $Y=1.515 $X2=0 $Y2=0
cc_252 N_B_c_243_n N_A_879_368#_c_627_n 2.45464e-19 $X=6.135 $Y=1.765 $X2=0
+ $Y2=0
cc_253 B N_A_879_368#_c_643_n 0.00507353f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_254 B N_A_879_368#_c_644_n 0.018819f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_255 N_B_c_239_n N_A_879_368#_c_644_n 0.00132101f $X=6 $Y=1.515 $X2=0 $Y2=0
cc_256 B N_A_879_368#_c_646_n 0.0206231f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_257 N_B_c_240_n N_VPWR_c_701_n 0.00278257f $X=4.765 $Y=1.765 $X2=0 $Y2=0
cc_258 N_B_c_241_n N_VPWR_c_701_n 0.00278257f $X=5.215 $Y=1.765 $X2=0 $Y2=0
cc_259 N_B_c_242_n N_VPWR_c_701_n 0.00278257f $X=5.685 $Y=1.765 $X2=0 $Y2=0
cc_260 N_B_c_243_n N_VPWR_c_701_n 0.0044313f $X=6.135 $Y=1.765 $X2=0 $Y2=0
cc_261 N_B_c_240_n N_VPWR_c_698_n 0.00358623f $X=4.765 $Y=1.765 $X2=0 $Y2=0
cc_262 N_B_c_241_n N_VPWR_c_698_n 0.00354011f $X=5.215 $Y=1.765 $X2=0 $Y2=0
cc_263 N_B_c_242_n N_VPWR_c_698_n 0.00354011f $X=5.685 $Y=1.765 $X2=0 $Y2=0
cc_264 N_B_c_243_n N_VPWR_c_698_n 0.00854206f $X=6.135 $Y=1.765 $X2=0 $Y2=0
cc_265 N_B_M1007_g N_VGND_c_781_n 0.00432719f $X=4.21 $Y=0.74 $X2=0 $Y2=0
cc_266 N_B_M1015_g N_VGND_c_783_n 0.00510848f $X=4.64 $Y=0.74 $X2=0 $Y2=0
cc_267 N_B_M1007_g N_VGND_c_791_n 0.00820772f $X=4.21 $Y=0.74 $X2=0 $Y2=0
cc_268 N_B_M1015_g N_VGND_c_791_n 0.00825037f $X=4.64 $Y=0.74 $X2=0 $Y2=0
cc_269 N_B_M1007_g N_VGND_c_793_n 0.00434272f $X=4.21 $Y=0.74 $X2=0 $Y2=0
cc_270 N_B_M1015_g N_VGND_c_793_n 0.00434272f $X=4.64 $Y=0.74 $X2=0 $Y2=0
cc_271 N_A_M1010_g N_Y_c_456_n 0.0146105f $X=7.12 $Y=0.74 $X2=0 $Y2=0
cc_272 N_A_c_315_n N_Y_c_456_n 0.0136138f $X=6.585 $Y=1.555 $X2=0 $Y2=0
cc_273 N_A_c_319_n N_Y_c_456_n 0.014057f $X=7.805 $Y=1.405 $X2=0 $Y2=0
cc_274 N_A_M1010_g N_Y_c_462_n 9.31832e-19 $X=7.12 $Y=0.74 $X2=0 $Y2=0
cc_275 N_A_M1017_g N_Y_c_462_n 0.00330748f $X=7.98 $Y=0.74 $X2=0 $Y2=0
cc_276 N_A_c_317_n N_Y_c_462_n 0.0123903f $X=7.98 $Y=1.532 $X2=0 $Y2=0
cc_277 N_A_c_318_n N_Y_c_462_n 0.00433553f $X=8.03 $Y=1.405 $X2=0 $Y2=0
cc_278 N_A_c_319_n N_Y_c_462_n 0.0406673f $X=7.805 $Y=1.405 $X2=0 $Y2=0
cc_279 N_A_c_320_n N_A_496_368#_c_562_n 3.13933e-19 $X=6.585 $Y=1.765 $X2=0
+ $Y2=0
cc_280 N_A_c_320_n N_A_879_368#_c_627_n 0.0104684f $X=6.585 $Y=1.765 $X2=0 $Y2=0
cc_281 N_A_c_321_n N_A_879_368#_c_627_n 6.64834e-19 $X=7.135 $Y=1.765 $X2=0
+ $Y2=0
cc_282 N_A_c_320_n N_A_879_368#_c_643_n 0.0143301f $X=6.585 $Y=1.765 $X2=0 $Y2=0
cc_283 N_A_c_312_n N_A_879_368#_c_643_n 0.00952485f $X=7.045 $Y=1.555 $X2=0
+ $Y2=0
cc_284 N_A_c_321_n N_A_879_368#_c_643_n 0.0132722f $X=7.135 $Y=1.765 $X2=0 $Y2=0
cc_285 N_A_c_319_n N_A_879_368#_c_643_n 0.00612933f $X=7.805 $Y=1.405 $X2=0
+ $Y2=0
cc_286 N_A_c_320_n N_A_879_368#_c_628_n 6.63528e-19 $X=6.585 $Y=1.765 $X2=0
+ $Y2=0
cc_287 N_A_c_321_n N_A_879_368#_c_628_n 0.0105688f $X=7.135 $Y=1.765 $X2=0 $Y2=0
cc_288 N_A_c_322_n N_A_879_368#_c_628_n 0.0105688f $X=7.585 $Y=1.765 $X2=0 $Y2=0
cc_289 N_A_c_323_n N_A_879_368#_c_628_n 6.63528e-19 $X=8.135 $Y=1.765 $X2=0
+ $Y2=0
cc_290 N_A_c_322_n N_A_879_368#_c_657_n 0.0132722f $X=7.585 $Y=1.765 $X2=0 $Y2=0
cc_291 N_A_c_323_n N_A_879_368#_c_657_n 0.0132722f $X=8.135 $Y=1.765 $X2=0 $Y2=0
cc_292 N_A_c_317_n N_A_879_368#_c_657_n 0.00798721f $X=7.98 $Y=1.532 $X2=0 $Y2=0
cc_293 N_A_c_319_n N_A_879_368#_c_657_n 0.0275323f $X=7.805 $Y=1.405 $X2=0 $Y2=0
cc_294 N_A_c_322_n N_A_879_368#_c_629_n 5.90388e-19 $X=7.585 $Y=1.765 $X2=0
+ $Y2=0
cc_295 N_A_c_323_n N_A_879_368#_c_629_n 0.00336601f $X=8.135 $Y=1.765 $X2=0
+ $Y2=0
cc_296 A N_A_879_368#_c_629_n 0.0265584f $X=8.315 $Y=1.21 $X2=0 $Y2=0
cc_297 N_A_c_317_n N_A_879_368#_c_629_n 3.97113e-19 $X=7.98 $Y=1.532 $X2=0 $Y2=0
cc_298 N_A_c_322_n N_A_879_368#_c_630_n 6.63528e-19 $X=7.585 $Y=1.765 $X2=0
+ $Y2=0
cc_299 N_A_c_323_n N_A_879_368#_c_630_n 0.0114814f $X=8.135 $Y=1.765 $X2=0 $Y2=0
cc_300 N_A_c_320_n N_A_879_368#_c_646_n 4.27055e-19 $X=6.585 $Y=1.765 $X2=0
+ $Y2=0
cc_301 N_A_c_321_n N_A_879_368#_c_668_n 5.11086e-19 $X=7.135 $Y=1.765 $X2=0
+ $Y2=0
cc_302 N_A_c_322_n N_A_879_368#_c_668_n 5.11086e-19 $X=7.585 $Y=1.765 $X2=0
+ $Y2=0
cc_303 N_A_c_317_n N_A_879_368#_c_668_n 0.00561879f $X=7.98 $Y=1.532 $X2=0 $Y2=0
cc_304 N_A_c_319_n N_A_879_368#_c_668_n 0.0134236f $X=7.805 $Y=1.405 $X2=0 $Y2=0
cc_305 N_A_c_320_n N_VPWR_c_699_n 0.00610756f $X=6.585 $Y=1.765 $X2=0 $Y2=0
cc_306 N_A_c_321_n N_VPWR_c_699_n 0.00598632f $X=7.135 $Y=1.765 $X2=0 $Y2=0
cc_307 N_A_c_322_n N_VPWR_c_700_n 0.00598632f $X=7.585 $Y=1.765 $X2=0 $Y2=0
cc_308 N_A_c_323_n N_VPWR_c_700_n 0.00737447f $X=8.135 $Y=1.765 $X2=0 $Y2=0
cc_309 N_A_c_320_n N_VPWR_c_701_n 0.00445602f $X=6.585 $Y=1.765 $X2=0 $Y2=0
cc_310 N_A_c_321_n N_VPWR_c_703_n 0.00445602f $X=7.135 $Y=1.765 $X2=0 $Y2=0
cc_311 N_A_c_322_n N_VPWR_c_703_n 0.00445602f $X=7.585 $Y=1.765 $X2=0 $Y2=0
cc_312 N_A_c_323_n N_VPWR_c_704_n 0.00445602f $X=8.135 $Y=1.765 $X2=0 $Y2=0
cc_313 N_A_c_320_n N_VPWR_c_698_n 0.00857881f $X=6.585 $Y=1.765 $X2=0 $Y2=0
cc_314 N_A_c_321_n N_VPWR_c_698_n 0.00857797f $X=7.135 $Y=1.765 $X2=0 $Y2=0
cc_315 N_A_c_322_n N_VPWR_c_698_n 0.00857797f $X=7.585 $Y=1.765 $X2=0 $Y2=0
cc_316 N_A_c_323_n N_VPWR_c_698_n 0.00861291f $X=8.135 $Y=1.765 $X2=0 $Y2=0
cc_317 N_A_M1017_g N_VGND_c_784_n 0.0151922f $X=7.98 $Y=0.74 $X2=0 $Y2=0
cc_318 A N_VGND_c_784_n 0.026357f $X=8.315 $Y=1.21 $X2=0 $Y2=0
cc_319 N_A_c_317_n N_VGND_c_784_n 5.99646e-19 $X=7.98 $Y=1.532 $X2=0 $Y2=0
cc_320 N_A_M1010_g N_VGND_c_788_n 0.00383152f $X=7.12 $Y=0.74 $X2=0 $Y2=0
cc_321 N_A_M1017_g N_VGND_c_788_n 0.00383152f $X=7.98 $Y=0.74 $X2=0 $Y2=0
cc_322 N_A_M1010_g N_VGND_c_791_n 0.00755866f $X=7.12 $Y=0.74 $X2=0 $Y2=0
cc_323 N_A_M1017_g N_VGND_c_791_n 0.00760481f $X=7.98 $Y=0.74 $X2=0 $Y2=0
cc_324 N_A_M1010_g N_VGND_c_794_n 0.0148268f $X=7.12 $Y=0.74 $X2=0 $Y2=0
cc_325 N_A_27_368#_c_387_n N_Y_M1000_s 0.00197722f $X=1.145 $Y=2.99 $X2=0 $Y2=0
cc_326 N_A_27_368#_c_389_n N_Y_M1013_s 0.00250873f $X=2.095 $Y=2.99 $X2=0 $Y2=0
cc_327 N_A_27_368#_M1000_d N_Y_c_466_n 0.00326865f $X=0.135 $Y=1.84 $X2=0 $Y2=0
cc_328 N_A_27_368#_c_386_n N_Y_c_466_n 0.00549591f $X=0.28 $Y=2.455 $X2=0 $Y2=0
cc_329 N_A_27_368#_M1000_d N_Y_c_464_n 0.00397608f $X=0.135 $Y=1.84 $X2=0 $Y2=0
cc_330 N_A_27_368#_c_386_n N_Y_c_464_n 0.0206806f $X=0.28 $Y=2.455 $X2=0 $Y2=0
cc_331 N_A_27_368#_M1012_d N_Y_c_468_n 0.00384138f $X=1.08 $Y=1.84 $X2=0 $Y2=0
cc_332 N_A_27_368#_c_395_n N_Y_c_468_n 0.0154248f $X=1.23 $Y=2.455 $X2=0 $Y2=0
cc_333 N_A_27_368#_c_387_n N_Y_c_477_n 0.0160777f $X=1.145 $Y=2.99 $X2=0 $Y2=0
cc_334 N_A_27_368#_c_395_n N_Y_c_477_n 0.0298377f $X=1.23 $Y=2.455 $X2=0 $Y2=0
cc_335 N_A_27_368#_c_389_n N_Y_c_482_n 0.018923f $X=2.095 $Y=2.99 $X2=0 $Y2=0
cc_336 N_A_27_368#_c_390_n N_Y_c_482_n 0.013092f $X=2.18 $Y=2.12 $X2=0 $Y2=0
cc_337 N_A_27_368#_c_400_n N_Y_c_482_n 0.039994f $X=2.18 $Y=2.4 $X2=0 $Y2=0
cc_338 N_A_27_368#_c_390_n N_Y_c_459_n 0.00568183f $X=2.18 $Y=2.12 $X2=0 $Y2=0
cc_339 N_A_27_368#_M1000_d Y 0.00227207f $X=0.135 $Y=1.84 $X2=0 $Y2=0
cc_340 N_A_27_368#_c_405_n N_A_496_368#_M1005_d 0.00359365f $X=2.97 $Y=2.035
+ $X2=-0.19 $Y2=1.66
cc_341 N_A_27_368#_c_409_n N_A_496_368#_M1016_d 0.00359365f $X=3.895 $Y=2.035
+ $X2=0 $Y2=0
cc_342 N_A_27_368#_c_400_n N_A_496_368#_c_565_n 0.039994f $X=2.18 $Y=2.4 $X2=0
+ $Y2=0
cc_343 N_A_27_368#_c_405_n N_A_496_368#_c_565_n 0.0171813f $X=2.97 $Y=2.035
+ $X2=0 $Y2=0
cc_344 N_A_27_368#_M1011_s N_A_496_368#_c_559_n 0.00197722f $X=2.93 $Y=1.84
+ $X2=0 $Y2=0
cc_345 N_A_27_368#_c_437_p N_A_496_368#_c_559_n 0.014157f $X=3.08 $Y=2.57 $X2=0
+ $Y2=0
cc_346 N_A_27_368#_c_389_n N_A_496_368#_c_560_n 0.0132987f $X=2.095 $Y=2.99
+ $X2=0 $Y2=0
cc_347 N_A_27_368#_c_409_n N_A_496_368#_c_572_n 0.0171813f $X=3.895 $Y=2.035
+ $X2=0 $Y2=0
cc_348 N_A_27_368#_c_392_n N_A_496_368#_c_572_n 0.0298377f $X=3.98 $Y=2.115
+ $X2=0 $Y2=0
cc_349 N_A_27_368#_M1021_s N_A_496_368#_c_561_n 0.00312144f $X=3.83 $Y=1.84
+ $X2=0 $Y2=0
cc_350 N_A_27_368#_c_392_n N_A_496_368#_c_561_n 0.018931f $X=3.98 $Y=2.115 $X2=0
+ $Y2=0
cc_351 N_A_27_368#_c_392_n N_A_879_368#_c_625_n 0.0128665f $X=3.98 $Y=2.115
+ $X2=0 $Y2=0
cc_352 N_A_27_368#_c_392_n N_A_879_368#_c_626_n 0.039691f $X=3.98 $Y=2.115 $X2=0
+ $Y2=0
cc_353 N_A_27_368#_c_387_n N_VPWR_c_701_n 0.0441612f $X=1.145 $Y=2.99 $X2=0
+ $Y2=0
cc_354 N_A_27_368#_c_388_n N_VPWR_c_701_n 0.0236566f $X=0.445 $Y=2.99 $X2=0
+ $Y2=0
cc_355 N_A_27_368#_c_389_n N_VPWR_c_701_n 0.0563945f $X=2.095 $Y=2.99 $X2=0
+ $Y2=0
cc_356 N_A_27_368#_c_391_n N_VPWR_c_701_n 0.017869f $X=1.27 $Y=2.99 $X2=0 $Y2=0
cc_357 N_A_27_368#_c_387_n N_VPWR_c_698_n 0.0249452f $X=1.145 $Y=2.99 $X2=0
+ $Y2=0
cc_358 N_A_27_368#_c_388_n N_VPWR_c_698_n 0.0128296f $X=0.445 $Y=2.99 $X2=0
+ $Y2=0
cc_359 N_A_27_368#_c_389_n N_VPWR_c_698_n 0.0316233f $X=2.095 $Y=2.99 $X2=0
+ $Y2=0
cc_360 N_A_27_368#_c_391_n N_VPWR_c_698_n 0.00965079f $X=1.27 $Y=2.99 $X2=0
+ $Y2=0
cc_361 N_Y_c_453_n N_VGND_M1002_d 0.00326483f $X=0.355 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_362 N_Y_c_457_n N_VGND_M1002_d 5.5277e-19 $X=0.615 $Y=0.765 $X2=-0.19
+ $Y2=-0.245
cc_363 N_Y_c_459_n N_VGND_M1020_d 0.00250873f $X=2.41 $Y=0.765 $X2=0 $Y2=0
cc_364 N_Y_c_454_n N_VGND_M1022_d 0.00250873f $X=4.26 $Y=1.095 $X2=0 $Y2=0
cc_365 N_Y_c_456_n N_VGND_M1015_s 0.0398609f $X=7.24 $Y=1.045 $X2=0 $Y2=0
cc_366 N_Y_c_453_n N_VGND_c_779_n 0.0207726f $X=0.355 $Y=1.095 $X2=0 $Y2=0
cc_367 N_Y_c_457_n N_VGND_c_779_n 0.00427553f $X=0.615 $Y=0.765 $X2=0 $Y2=0
cc_368 N_Y_c_458_n N_VGND_c_779_n 0.0232074f $X=1.74 $Y=0.765 $X2=0 $Y2=0
cc_369 N_Y_c_458_n N_VGND_c_780_n 0.0192747f $X=1.74 $Y=0.765 $X2=0 $Y2=0
cc_370 N_Y_c_459_n N_VGND_c_780_n 0.0209867f $X=2.41 $Y=0.765 $X2=0 $Y2=0
cc_371 N_Y_c_460_n N_VGND_c_780_n 0.0213507f $X=3.59 $Y=0.765 $X2=0 $Y2=0
cc_372 N_Y_c_454_n N_VGND_c_781_n 0.0209867f $X=4.26 $Y=1.095 $X2=0 $Y2=0
cc_373 N_Y_c_455_n N_VGND_c_781_n 0.0191765f $X=4.425 $Y=0.515 $X2=0 $Y2=0
cc_374 N_Y_c_460_n N_VGND_c_781_n 0.0192747f $X=3.59 $Y=0.765 $X2=0 $Y2=0
cc_375 N_Y_c_455_n N_VGND_c_783_n 0.0174363f $X=4.425 $Y=0.515 $X2=0 $Y2=0
cc_376 N_Y_c_456_n N_VGND_c_783_n 0.181264f $X=7.24 $Y=1.045 $X2=0 $Y2=0
cc_377 N_Y_c_462_n N_VGND_c_784_n 0.0265927f $X=7.335 $Y=0.965 $X2=0 $Y2=0
cc_378 N_Y_c_460_n N_VGND_c_785_n 0.0523677f $X=3.59 $Y=0.765 $X2=0 $Y2=0
cc_379 N_Y_c_462_n N_VGND_c_788_n 0.0288054f $X=7.335 $Y=0.965 $X2=0 $Y2=0
cc_380 N_Y_c_458_n N_VGND_c_790_n 0.0499979f $X=1.74 $Y=0.765 $X2=0 $Y2=0
cc_381 N_Y_c_455_n N_VGND_c_791_n 0.0118826f $X=4.425 $Y=0.515 $X2=0 $Y2=0
cc_382 N_Y_c_458_n N_VGND_c_791_n 0.041525f $X=1.74 $Y=0.765 $X2=0 $Y2=0
cc_383 N_Y_c_460_n N_VGND_c_791_n 0.0434345f $X=3.59 $Y=0.765 $X2=0 $Y2=0
cc_384 N_Y_c_462_n N_VGND_c_791_n 0.02303f $X=7.335 $Y=0.965 $X2=0 $Y2=0
cc_385 N_Y_c_455_n N_VGND_c_793_n 0.0144922f $X=4.425 $Y=0.515 $X2=0 $Y2=0
cc_386 N_Y_c_462_n N_VGND_c_794_n 0.0203431f $X=7.335 $Y=0.965 $X2=0 $Y2=0
cc_387 N_A_496_368#_c_561_n N_A_879_368#_M1003_s 0.00312144f $X=4.825 $Y=2.99
+ $X2=-0.19 $Y2=1.66
cc_388 N_A_496_368#_c_562_n N_A_879_368#_M1004_s 0.00218982f $X=5.745 $Y=2.99
+ $X2=0 $Y2=0
cc_389 N_A_496_368#_c_561_n N_A_879_368#_c_626_n 0.018931f $X=4.825 $Y=2.99
+ $X2=0 $Y2=0
cc_390 N_A_496_368#_c_579_n N_A_879_368#_c_626_n 0.0291672f $X=4.99 $Y=2.385
+ $X2=0 $Y2=0
cc_391 N_A_496_368#_M1003_d N_A_879_368#_c_634_n 0.00364166f $X=4.84 $Y=1.84
+ $X2=0 $Y2=0
cc_392 N_A_496_368#_c_579_n N_A_879_368#_c_634_n 0.0164557f $X=4.99 $Y=2.385
+ $X2=0 $Y2=0
cc_393 N_A_496_368#_c_562_n N_A_879_368#_c_680_n 0.0156793f $X=5.745 $Y=2.99
+ $X2=0 $Y2=0
cc_394 N_A_496_368#_M1006_d N_A_879_368#_c_638_n 0.00364166f $X=5.76 $Y=1.84
+ $X2=0 $Y2=0
cc_395 N_A_496_368#_c_585_n N_A_879_368#_c_638_n 0.0164557f $X=5.91 $Y=2.385
+ $X2=0 $Y2=0
cc_396 N_A_496_368#_c_562_n N_A_879_368#_c_627_n 0.00375634f $X=5.745 $Y=2.99
+ $X2=0 $Y2=0
cc_397 N_A_496_368#_c_562_n N_VPWR_c_699_n 0.00294239f $X=5.745 $Y=2.99 $X2=0
+ $Y2=0
cc_398 N_A_496_368#_c_559_n N_VPWR_c_701_n 0.03588f $X=3.365 $Y=2.99 $X2=0 $Y2=0
cc_399 N_A_496_368#_c_560_n N_VPWR_c_701_n 0.0235512f $X=2.795 $Y=2.99 $X2=0
+ $Y2=0
cc_400 N_A_496_368#_c_561_n N_VPWR_c_701_n 0.0719543f $X=4.825 $Y=2.99 $X2=0
+ $Y2=0
cc_401 N_A_496_368#_c_562_n N_VPWR_c_701_n 0.0607196f $X=5.745 $Y=2.99 $X2=0
+ $Y2=0
cc_402 N_A_496_368#_c_563_n N_VPWR_c_701_n 0.0235512f $X=3.53 $Y=2.99 $X2=0
+ $Y2=0
cc_403 N_A_496_368#_c_564_n N_VPWR_c_701_n 0.0235512f $X=4.99 $Y=2.99 $X2=0
+ $Y2=0
cc_404 N_A_496_368#_c_559_n N_VPWR_c_698_n 0.0201952f $X=3.365 $Y=2.99 $X2=0
+ $Y2=0
cc_405 N_A_496_368#_c_560_n N_VPWR_c_698_n 0.0126924f $X=2.795 $Y=2.99 $X2=0
+ $Y2=0
cc_406 N_A_496_368#_c_561_n N_VPWR_c_698_n 0.04125f $X=4.825 $Y=2.99 $X2=0 $Y2=0
cc_407 N_A_496_368#_c_562_n N_VPWR_c_698_n 0.0336395f $X=5.745 $Y=2.99 $X2=0
+ $Y2=0
cc_408 N_A_496_368#_c_563_n N_VPWR_c_698_n 0.0126924f $X=3.53 $Y=2.99 $X2=0
+ $Y2=0
cc_409 N_A_496_368#_c_564_n N_VPWR_c_698_n 0.0126924f $X=4.99 $Y=2.99 $X2=0
+ $Y2=0
cc_410 N_A_879_368#_c_643_n N_VPWR_M1001_s 0.00715624f $X=7.195 $Y=2.035
+ $X2=-0.19 $Y2=1.66
cc_411 N_A_879_368#_c_657_n N_VPWR_M1014_s 0.00671265f $X=8.195 $Y=2.035 $X2=0
+ $Y2=0
cc_412 N_A_879_368#_c_627_n N_VPWR_c_699_n 0.0258971f $X=6.36 $Y=2.445 $X2=0
+ $Y2=0
cc_413 N_A_879_368#_c_643_n N_VPWR_c_699_n 0.0232685f $X=7.195 $Y=2.035 $X2=0
+ $Y2=0
cc_414 N_A_879_368#_c_628_n N_VPWR_c_699_n 0.0266809f $X=7.36 $Y=2.815 $X2=0
+ $Y2=0
cc_415 N_A_879_368#_c_628_n N_VPWR_c_700_n 0.0266809f $X=7.36 $Y=2.815 $X2=0
+ $Y2=0
cc_416 N_A_879_368#_c_657_n N_VPWR_c_700_n 0.0232685f $X=8.195 $Y=2.035 $X2=0
+ $Y2=0
cc_417 N_A_879_368#_c_630_n N_VPWR_c_700_n 0.0266809f $X=8.36 $Y=2.815 $X2=0
+ $Y2=0
cc_418 N_A_879_368#_c_627_n N_VPWR_c_701_n 0.0119166f $X=6.36 $Y=2.445 $X2=0
+ $Y2=0
cc_419 N_A_879_368#_c_628_n N_VPWR_c_703_n 0.014552f $X=7.36 $Y=2.815 $X2=0
+ $Y2=0
cc_420 N_A_879_368#_c_630_n N_VPWR_c_704_n 0.0145938f $X=8.36 $Y=2.815 $X2=0
+ $Y2=0
cc_421 N_A_879_368#_c_627_n N_VPWR_c_698_n 0.00983061f $X=6.36 $Y=2.445 $X2=0
+ $Y2=0
cc_422 N_A_879_368#_c_628_n N_VPWR_c_698_n 0.0119791f $X=7.36 $Y=2.815 $X2=0
+ $Y2=0
cc_423 N_A_879_368#_c_630_n N_VPWR_c_698_n 0.0120466f $X=8.36 $Y=2.815 $X2=0
+ $Y2=0
