* File: sky130_fd_sc_ls__nor2b_2.pxi.spice
* Created: Wed Sep  2 11:14:27 2020
* 
x_PM_SKY130_FD_SC_LS__NOR2B_2%B_N N_B_N_c_63_n N_B_N_M1008_g N_B_N_M1002_g B_N
+ N_B_N_c_62_n PM_SKY130_FD_SC_LS__NOR2B_2%B_N
x_PM_SKY130_FD_SC_LS__NOR2B_2%A_27_392# N_A_27_392#_M1002_s N_A_27_392#_M1008_s
+ N_A_27_392#_c_94_n N_A_27_392#_M1001_g N_A_27_392#_c_102_n N_A_27_392#_M1006_g
+ N_A_27_392#_c_95_n N_A_27_392#_M1004_g N_A_27_392#_c_103_n N_A_27_392#_M1009_g
+ N_A_27_392#_c_96_n N_A_27_392#_c_97_n N_A_27_392#_c_98_n N_A_27_392#_c_99_n
+ N_A_27_392#_c_100_n N_A_27_392#_c_101_n PM_SKY130_FD_SC_LS__NOR2B_2%A_27_392#
x_PM_SKY130_FD_SC_LS__NOR2B_2%A N_A_M1005_g N_A_c_177_n N_A_M1000_g N_A_M1007_g
+ N_A_c_178_n N_A_M1003_g A A N_A_c_176_n PM_SKY130_FD_SC_LS__NOR2B_2%A
x_PM_SKY130_FD_SC_LS__NOR2B_2%VPWR N_VPWR_M1008_d N_VPWR_M1000_d N_VPWR_c_225_n
+ N_VPWR_c_226_n VPWR N_VPWR_c_227_n N_VPWR_c_228_n N_VPWR_c_229_n
+ N_VPWR_c_224_n N_VPWR_c_231_n N_VPWR_c_232_n PM_SKY130_FD_SC_LS__NOR2B_2%VPWR
x_PM_SKY130_FD_SC_LS__NOR2B_2%A_228_368# N_A_228_368#_M1006_s
+ N_A_228_368#_M1009_s N_A_228_368#_M1003_s N_A_228_368#_c_266_n
+ N_A_228_368#_c_267_n N_A_228_368#_c_268_n N_A_228_368#_c_282_n
+ N_A_228_368#_c_283_n N_A_228_368#_c_290_n N_A_228_368#_c_269_n
+ N_A_228_368#_c_270_n PM_SKY130_FD_SC_LS__NOR2B_2%A_228_368#
x_PM_SKY130_FD_SC_LS__NOR2B_2%Y N_Y_M1001_d N_Y_M1005_d N_Y_M1006_d N_Y_c_315_n
+ N_Y_c_316_n N_Y_c_317_n N_Y_c_318_n N_Y_c_319_n N_Y_c_320_n N_Y_c_321_n Y
+ N_Y_c_322_n PM_SKY130_FD_SC_LS__NOR2B_2%Y
x_PM_SKY130_FD_SC_LS__NOR2B_2%VGND N_VGND_M1002_d N_VGND_M1004_s N_VGND_M1007_s
+ N_VGND_c_369_n N_VGND_c_370_n N_VGND_c_371_n N_VGND_c_372_n VGND
+ N_VGND_c_373_n N_VGND_c_374_n N_VGND_c_375_n N_VGND_c_376_n N_VGND_c_377_n
+ N_VGND_c_378_n PM_SKY130_FD_SC_LS__NOR2B_2%VGND
cc_1 VNB N_B_N_M1002_g 0.0367247f $X=-0.19 $Y=-0.245 $X2=0.83 $Y2=0.79
cc_2 VNB B_N 0.00207353f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_3 VNB N_B_N_c_62_n 0.0284009f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=1.635
cc_4 VNB N_A_27_392#_c_94_n 0.018486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_5 VNB N_A_27_392#_c_95_n 0.016567f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=1.635
cc_6 VNB N_A_27_392#_c_96_n 0.0432843f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_27_392#_c_97_n 0.0192881f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_27_392#_c_98_n 0.0121892f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_27_392#_c_99_n 0.0145497f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_27_392#_c_100_n 0.00587637f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_27_392#_c_101_n 0.0823364f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_M1005_g 0.023477f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.46
cc_13 VNB N_A_M1007_g 0.0269184f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.677
cc_14 VNB A 0.00224035f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_c_176_n 0.0444267f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_VPWR_c_224_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_Y_c_315_n 0.00280126f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=1.635
cc_18 VNB N_Y_c_316_n 5.19053e-19 $X=-0.19 $Y=-0.245 $X2=0.83 $Y2=1.677
cc_19 VNB N_Y_c_317_n 0.00135442f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_Y_c_318_n 0.00392956f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_Y_c_319_n 0.00252696f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_Y_c_320_n 0.00292043f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_Y_c_321_n 0.00186002f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_Y_c_322_n 0.0212378f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_369_n 0.0127511f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=1.635
cc_26 VNB N_VGND_c_370_n 0.00277973f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_371_n 0.0120457f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_372_n 0.0279043f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_373_n 0.0292002f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_374_n 0.0185368f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_375_n 0.0167762f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_376_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_377_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_378_n 0.210833f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VPB N_B_N_c_63_n 0.021205f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=1.885
cc_36 VPB B_N 0.00249009f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_37 VPB N_B_N_c_62_n 0.031283f $X=-0.19 $Y=1.66 $X2=0.695 $Y2=1.635
cc_38 VPB N_A_27_392#_c_102_n 0.0176597f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=1.677
cc_39 VPB N_A_27_392#_c_103_n 0.0148823f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_40 VPB N_A_27_392#_c_97_n 0.0558724f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_41 VPB N_A_27_392#_c_101_n 0.0161002f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_42 VPB N_A_c_177_n 0.0152418f $X=-0.19 $Y=1.66 $X2=0.83 $Y2=0.79
cc_43 VPB N_A_c_178_n 0.0199141f $X=-0.19 $Y=1.66 $X2=0.695 $Y2=1.635
cc_44 VPB A 0.00637702f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_45 VPB N_A_c_176_n 0.02384f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_225_n 0.0155045f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_226_n 0.00538737f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_227_n 0.0178682f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_228_n 0.0407833f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_229_n 0.0178682f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_224_n 0.0730651f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_231_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_232_n 0.00460249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_A_228_368#_c_266_n 0.0131449f $X=-0.19 $Y=1.66 $X2=0.695 $Y2=1.635
cc_55 VPB N_A_228_368#_c_267_n 0.00431993f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_A_228_368#_c_268_n 0.00431456f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_A_228_368#_c_269_n 0.015978f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_A_228_368#_c_270_n 0.0341208f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_Y_c_317_n 0.00320608f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 N_B_N_M1002_g N_A_27_392#_c_94_n 0.0171333f $X=0.83 $Y=0.79 $X2=0 $Y2=0
cc_61 N_B_N_c_62_n N_A_27_392#_c_102_n 9.02862e-19 $X=0.695 $Y=1.635 $X2=0 $Y2=0
cc_62 N_B_N_M1002_g N_A_27_392#_c_96_n 0.0106849f $X=0.83 $Y=0.79 $X2=0 $Y2=0
cc_63 N_B_N_c_63_n N_A_27_392#_c_97_n 0.00706891f $X=0.5 $Y=1.885 $X2=0 $Y2=0
cc_64 N_B_N_M1002_g N_A_27_392#_c_97_n 0.00477364f $X=0.83 $Y=0.79 $X2=0 $Y2=0
cc_65 B_N N_A_27_392#_c_97_n 0.025547f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_66 N_B_N_c_62_n N_A_27_392#_c_97_n 0.0129015f $X=0.695 $Y=1.635 $X2=0 $Y2=0
cc_67 N_B_N_M1002_g N_A_27_392#_c_98_n 0.0118985f $X=0.83 $Y=0.79 $X2=0 $Y2=0
cc_68 B_N N_A_27_392#_c_98_n 0.00563709f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_69 N_B_N_M1002_g N_A_27_392#_c_99_n 0.00476166f $X=0.83 $Y=0.79 $X2=0 $Y2=0
cc_70 B_N N_A_27_392#_c_99_n 0.0209889f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_71 N_B_N_c_62_n N_A_27_392#_c_99_n 0.0075801f $X=0.695 $Y=1.635 $X2=0 $Y2=0
cc_72 N_B_N_M1002_g N_A_27_392#_c_100_n 0.00158684f $X=0.83 $Y=0.79 $X2=0 $Y2=0
cc_73 B_N N_A_27_392#_c_100_n 0.00397231f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_74 N_B_N_M1002_g N_A_27_392#_c_101_n 0.0191582f $X=0.83 $Y=0.79 $X2=0 $Y2=0
cc_75 B_N N_A_27_392#_c_101_n 0.00153638f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_76 N_B_N_c_62_n N_A_27_392#_c_101_n 0.00681533f $X=0.695 $Y=1.635 $X2=0 $Y2=0
cc_77 N_B_N_c_63_n N_VPWR_c_225_n 0.0185298f $X=0.5 $Y=1.885 $X2=0 $Y2=0
cc_78 B_N N_VPWR_c_225_n 0.0220821f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_79 N_B_N_c_62_n N_VPWR_c_225_n 0.00301557f $X=0.695 $Y=1.635 $X2=0 $Y2=0
cc_80 N_B_N_c_63_n N_VPWR_c_227_n 0.00413917f $X=0.5 $Y=1.885 $X2=0 $Y2=0
cc_81 N_B_N_c_63_n N_VPWR_c_224_n 0.00821204f $X=0.5 $Y=1.885 $X2=0 $Y2=0
cc_82 N_B_N_c_63_n N_A_228_368#_c_266_n 0.0020061f $X=0.5 $Y=1.885 $X2=0 $Y2=0
cc_83 N_B_N_c_62_n N_A_228_368#_c_266_n 0.00168698f $X=0.695 $Y=1.635 $X2=0
+ $Y2=0
cc_84 N_B_N_c_63_n N_A_228_368#_c_268_n 5.94256e-19 $X=0.5 $Y=1.885 $X2=0 $Y2=0
cc_85 N_B_N_M1002_g N_VGND_c_369_n 0.0080577f $X=0.83 $Y=0.79 $X2=0 $Y2=0
cc_86 N_B_N_M1002_g N_VGND_c_373_n 0.00485498f $X=0.83 $Y=0.79 $X2=0 $Y2=0
cc_87 N_B_N_M1002_g N_VGND_c_378_n 0.00514438f $X=0.83 $Y=0.79 $X2=0 $Y2=0
cc_88 N_A_27_392#_c_95_n N_A_M1005_g 0.0239839f $X=1.915 $Y=1.22 $X2=0 $Y2=0
cc_89 N_A_27_392#_c_101_n N_A_M1005_g 0.0263421f $X=1.915 $Y=1.492 $X2=0 $Y2=0
cc_90 N_A_27_392#_c_103_n N_A_c_177_n 0.00893213f $X=1.96 $Y=1.765 $X2=0 $Y2=0
cc_91 N_A_27_392#_c_101_n A 0.0106625f $X=1.915 $Y=1.492 $X2=0 $Y2=0
cc_92 N_A_27_392#_c_101_n N_A_c_176_n 0.00401348f $X=1.915 $Y=1.492 $X2=0 $Y2=0
cc_93 N_A_27_392#_c_102_n N_VPWR_c_225_n 0.00256389f $X=1.51 $Y=1.765 $X2=0
+ $Y2=0
cc_94 N_A_27_392#_c_97_n N_VPWR_c_225_n 0.0677511f $X=0.275 $Y=2.105 $X2=0 $Y2=0
cc_95 N_A_27_392#_c_98_n N_VPWR_c_225_n 8.30447e-19 $X=1.145 $Y=1.215 $X2=0
+ $Y2=0
cc_96 N_A_27_392#_c_97_n N_VPWR_c_227_n 0.011066f $X=0.275 $Y=2.105 $X2=0 $Y2=0
cc_97 N_A_27_392#_c_102_n N_VPWR_c_228_n 0.00278257f $X=1.51 $Y=1.765 $X2=0
+ $Y2=0
cc_98 N_A_27_392#_c_103_n N_VPWR_c_228_n 0.00278257f $X=1.96 $Y=1.765 $X2=0
+ $Y2=0
cc_99 N_A_27_392#_c_102_n N_VPWR_c_224_n 0.00358623f $X=1.51 $Y=1.765 $X2=0
+ $Y2=0
cc_100 N_A_27_392#_c_103_n N_VPWR_c_224_n 0.00353905f $X=1.96 $Y=1.765 $X2=0
+ $Y2=0
cc_101 N_A_27_392#_c_97_n N_VPWR_c_224_n 0.00915947f $X=0.275 $Y=2.105 $X2=0
+ $Y2=0
cc_102 N_A_27_392#_c_102_n N_A_228_368#_c_266_n 0.01381f $X=1.51 $Y=1.765 $X2=0
+ $Y2=0
cc_103 N_A_27_392#_c_103_n N_A_228_368#_c_266_n 7.07518e-19 $X=1.96 $Y=1.765
+ $X2=0 $Y2=0
cc_104 N_A_27_392#_c_98_n N_A_228_368#_c_266_n 9.32104e-19 $X=1.145 $Y=1.215
+ $X2=0 $Y2=0
cc_105 N_A_27_392#_c_100_n N_A_228_368#_c_266_n 0.0183877f $X=1.31 $Y=1.215
+ $X2=0 $Y2=0
cc_106 N_A_27_392#_c_101_n N_A_228_368#_c_266_n 0.00408351f $X=1.915 $Y=1.492
+ $X2=0 $Y2=0
cc_107 N_A_27_392#_c_102_n N_A_228_368#_c_267_n 0.0108414f $X=1.51 $Y=1.765
+ $X2=0 $Y2=0
cc_108 N_A_27_392#_c_103_n N_A_228_368#_c_267_n 0.0125587f $X=1.96 $Y=1.765
+ $X2=0 $Y2=0
cc_109 N_A_27_392#_c_102_n N_A_228_368#_c_268_n 0.00262934f $X=1.51 $Y=1.765
+ $X2=0 $Y2=0
cc_110 N_A_27_392#_c_103_n N_A_228_368#_c_282_n 0.00245972f $X=1.96 $Y=1.765
+ $X2=0 $Y2=0
cc_111 N_A_27_392#_c_102_n N_A_228_368#_c_283_n 6.22492e-19 $X=1.51 $Y=1.765
+ $X2=0 $Y2=0
cc_112 N_A_27_392#_c_103_n N_A_228_368#_c_283_n 0.00931603f $X=1.96 $Y=1.765
+ $X2=0 $Y2=0
cc_113 N_A_27_392#_c_94_n N_Y_c_315_n 0.00505604f $X=1.435 $Y=1.22 $X2=0 $Y2=0
cc_114 N_A_27_392#_c_94_n N_Y_c_316_n 0.00778619f $X=1.435 $Y=1.22 $X2=0 $Y2=0
cc_115 N_A_27_392#_c_100_n N_Y_c_316_n 0.00421645f $X=1.31 $Y=1.215 $X2=0 $Y2=0
cc_116 N_A_27_392#_c_101_n N_Y_c_316_n 0.00181131f $X=1.915 $Y=1.492 $X2=0 $Y2=0
cc_117 N_A_27_392#_c_94_n N_Y_c_317_n 2.53709e-19 $X=1.435 $Y=1.22 $X2=0 $Y2=0
cc_118 N_A_27_392#_c_102_n N_Y_c_317_n 0.00514255f $X=1.51 $Y=1.765 $X2=0 $Y2=0
cc_119 N_A_27_392#_c_95_n N_Y_c_317_n 0.00100575f $X=1.915 $Y=1.22 $X2=0 $Y2=0
cc_120 N_A_27_392#_c_103_n N_Y_c_317_n 0.00706473f $X=1.96 $Y=1.765 $X2=0 $Y2=0
cc_121 N_A_27_392#_c_100_n N_Y_c_317_n 0.0265536f $X=1.31 $Y=1.215 $X2=0 $Y2=0
cc_122 N_A_27_392#_c_101_n N_Y_c_317_n 0.0312076f $X=1.915 $Y=1.492 $X2=0 $Y2=0
cc_123 N_A_27_392#_c_95_n N_Y_c_318_n 0.0199327f $X=1.915 $Y=1.22 $X2=0 $Y2=0
cc_124 N_A_27_392#_c_101_n N_Y_c_318_n 0.0028271f $X=1.915 $Y=1.492 $X2=0 $Y2=0
cc_125 N_A_27_392#_c_94_n N_VGND_c_369_n 0.00714781f $X=1.435 $Y=1.22 $X2=0
+ $Y2=0
cc_126 N_A_27_392#_c_96_n N_VGND_c_369_n 0.036192f $X=0.615 $Y=0.615 $X2=0 $Y2=0
cc_127 N_A_27_392#_c_98_n N_VGND_c_369_n 0.0131477f $X=1.145 $Y=1.215 $X2=0
+ $Y2=0
cc_128 N_A_27_392#_c_100_n N_VGND_c_369_n 0.0143981f $X=1.31 $Y=1.215 $X2=0
+ $Y2=0
cc_129 N_A_27_392#_c_101_n N_VGND_c_369_n 0.00102906f $X=1.915 $Y=1.492 $X2=0
+ $Y2=0
cc_130 N_A_27_392#_c_94_n N_VGND_c_370_n 4.45911e-19 $X=1.435 $Y=1.22 $X2=0
+ $Y2=0
cc_131 N_A_27_392#_c_95_n N_VGND_c_370_n 0.00825039f $X=1.915 $Y=1.22 $X2=0
+ $Y2=0
cc_132 N_A_27_392#_c_96_n N_VGND_c_373_n 0.0211421f $X=0.615 $Y=0.615 $X2=0
+ $Y2=0
cc_133 N_A_27_392#_c_94_n N_VGND_c_374_n 0.00434272f $X=1.435 $Y=1.22 $X2=0
+ $Y2=0
cc_134 N_A_27_392#_c_95_n N_VGND_c_374_n 0.00444681f $X=1.915 $Y=1.22 $X2=0
+ $Y2=0
cc_135 N_A_27_392#_c_94_n N_VGND_c_378_n 0.00825538f $X=1.435 $Y=1.22 $X2=0
+ $Y2=0
cc_136 N_A_27_392#_c_95_n N_VGND_c_378_n 0.00877997f $X=1.915 $Y=1.22 $X2=0
+ $Y2=0
cc_137 N_A_27_392#_c_96_n N_VGND_c_378_n 0.0231103f $X=0.615 $Y=0.615 $X2=0
+ $Y2=0
cc_138 N_A_c_177_n N_VPWR_c_226_n 0.00356844f $X=2.41 $Y=1.765 $X2=0 $Y2=0
cc_139 N_A_c_178_n N_VPWR_c_226_n 0.0135832f $X=2.86 $Y=1.765 $X2=0 $Y2=0
cc_140 N_A_c_177_n N_VPWR_c_228_n 0.0044313f $X=2.41 $Y=1.765 $X2=0 $Y2=0
cc_141 N_A_c_178_n N_VPWR_c_229_n 0.00413917f $X=2.86 $Y=1.765 $X2=0 $Y2=0
cc_142 N_A_c_177_n N_VPWR_c_224_n 0.00853445f $X=2.41 $Y=1.765 $X2=0 $Y2=0
cc_143 N_A_c_178_n N_VPWR_c_224_n 0.00821204f $X=2.86 $Y=1.765 $X2=0 $Y2=0
cc_144 N_A_c_177_n N_A_228_368#_c_267_n 0.0032261f $X=2.41 $Y=1.765 $X2=0 $Y2=0
cc_145 N_A_c_177_n N_A_228_368#_c_282_n 4.27055e-19 $X=2.41 $Y=1.765 $X2=0 $Y2=0
cc_146 A N_A_228_368#_c_282_n 0.0221462f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_147 N_A_c_177_n N_A_228_368#_c_283_n 0.0095181f $X=2.41 $Y=1.765 $X2=0 $Y2=0
cc_148 N_A_c_178_n N_A_228_368#_c_283_n 4.50629e-19 $X=2.86 $Y=1.765 $X2=0 $Y2=0
cc_149 N_A_c_177_n N_A_228_368#_c_290_n 0.0120074f $X=2.41 $Y=1.765 $X2=0 $Y2=0
cc_150 N_A_c_178_n N_A_228_368#_c_290_n 0.0171961f $X=2.86 $Y=1.765 $X2=0 $Y2=0
cc_151 A N_A_228_368#_c_290_n 0.0282713f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_152 N_A_c_176_n N_A_228_368#_c_290_n 0.00125848f $X=2.845 $Y=1.557 $X2=0
+ $Y2=0
cc_153 N_A_c_178_n N_A_228_368#_c_269_n 0.00314968f $X=2.86 $Y=1.765 $X2=0 $Y2=0
cc_154 N_A_c_178_n N_A_228_368#_c_270_n 0.00526798f $X=2.86 $Y=1.765 $X2=0 $Y2=0
cc_155 N_A_M1005_g N_Y_c_317_n 5.38267e-19 $X=2.365 $Y=0.74 $X2=0 $Y2=0
cc_156 A N_Y_c_317_n 0.0268883f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_157 N_A_M1005_g N_Y_c_318_n 0.0147681f $X=2.365 $Y=0.74 $X2=0 $Y2=0
cc_158 A N_Y_c_318_n 0.0356018f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_159 N_A_M1005_g N_Y_c_319_n 4.49298e-19 $X=2.365 $Y=0.74 $X2=0 $Y2=0
cc_160 N_A_M1007_g N_Y_c_319_n 4.7485e-19 $X=2.845 $Y=0.74 $X2=0 $Y2=0
cc_161 N_A_M1007_g N_Y_c_320_n 0.0188046f $X=2.845 $Y=0.74 $X2=0 $Y2=0
cc_162 A N_Y_c_320_n 7.29585e-19 $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_163 N_A_c_176_n N_Y_c_320_n 9.98122e-19 $X=2.845 $Y=1.557 $X2=0 $Y2=0
cc_164 A N_Y_c_321_n 0.0214748f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_165 N_A_c_176_n N_Y_c_321_n 0.00349435f $X=2.845 $Y=1.557 $X2=0 $Y2=0
cc_166 N_A_M1007_g N_Y_c_322_n 0.00964993f $X=2.845 $Y=0.74 $X2=0 $Y2=0
cc_167 A N_Y_c_322_n 0.00361538f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_168 N_A_M1005_g N_VGND_c_370_n 0.00982302f $X=2.365 $Y=0.74 $X2=0 $Y2=0
cc_169 N_A_M1007_g N_VGND_c_370_n 4.5319e-19 $X=2.845 $Y=0.74 $X2=0 $Y2=0
cc_170 N_A_M1005_g N_VGND_c_372_n 4.40885e-19 $X=2.365 $Y=0.74 $X2=0 $Y2=0
cc_171 N_A_M1007_g N_VGND_c_372_n 0.0111523f $X=2.845 $Y=0.74 $X2=0 $Y2=0
cc_172 N_A_M1005_g N_VGND_c_375_n 0.00383152f $X=2.365 $Y=0.74 $X2=0 $Y2=0
cc_173 N_A_M1007_g N_VGND_c_375_n 0.00444681f $X=2.845 $Y=0.74 $X2=0 $Y2=0
cc_174 N_A_M1005_g N_VGND_c_378_n 0.00758019f $X=2.365 $Y=0.74 $X2=0 $Y2=0
cc_175 N_A_M1007_g N_VGND_c_378_n 0.00877997f $X=2.845 $Y=0.74 $X2=0 $Y2=0
cc_176 N_VPWR_c_225_n N_A_228_368#_c_266_n 0.0630028f $X=0.725 $Y=2.135 $X2=0
+ $Y2=0
cc_177 N_VPWR_c_226_n N_A_228_368#_c_267_n 0.012272f $X=2.635 $Y=2.455 $X2=0
+ $Y2=0
cc_178 N_VPWR_c_228_n N_A_228_368#_c_267_n 0.0594312f $X=2.55 $Y=3.33 $X2=0
+ $Y2=0
cc_179 N_VPWR_c_224_n N_A_228_368#_c_267_n 0.0328875f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_180 N_VPWR_c_225_n N_A_228_368#_c_268_n 0.0121617f $X=0.725 $Y=2.135 $X2=0
+ $Y2=0
cc_181 N_VPWR_c_228_n N_A_228_368#_c_268_n 0.0236039f $X=2.55 $Y=3.33 $X2=0
+ $Y2=0
cc_182 N_VPWR_c_224_n N_A_228_368#_c_268_n 0.012761f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_183 N_VPWR_c_226_n N_A_228_368#_c_283_n 0.0412035f $X=2.635 $Y=2.455 $X2=0
+ $Y2=0
cc_184 N_VPWR_M1000_d N_A_228_368#_c_290_n 0.00384138f $X=2.485 $Y=1.84 $X2=0
+ $Y2=0
cc_185 N_VPWR_c_226_n N_A_228_368#_c_290_n 0.0154248f $X=2.635 $Y=2.455 $X2=0
+ $Y2=0
cc_186 N_VPWR_c_226_n N_A_228_368#_c_270_n 0.0453479f $X=2.635 $Y=2.455 $X2=0
+ $Y2=0
cc_187 N_VPWR_c_229_n N_A_228_368#_c_270_n 0.011066f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_188 N_VPWR_c_224_n N_A_228_368#_c_270_n 0.00915947f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_189 N_A_228_368#_c_267_n N_Y_M1006_d 0.00218242f $X=2.02 $Y=2.99 $X2=0 $Y2=0
cc_190 N_A_228_368#_c_266_n N_Y_c_317_n 0.0609301f $X=1.285 $Y=1.985 $X2=0 $Y2=0
cc_191 N_A_228_368#_c_267_n N_Y_c_317_n 0.0131675f $X=2.02 $Y=2.99 $X2=0 $Y2=0
cc_192 N_A_228_368#_c_282_n N_Y_c_317_n 0.0117998f $X=2.185 $Y=2.12 $X2=0 $Y2=0
cc_193 N_A_228_368#_c_283_n N_Y_c_317_n 0.0401125f $X=2.185 $Y=2.815 $X2=0 $Y2=0
cc_194 N_A_228_368#_c_269_n N_Y_c_322_n 0.0111281f $X=3.125 $Y=2.12 $X2=0 $Y2=0
cc_195 N_Y_c_318_n N_VGND_M1004_s 0.001993f $X=2.495 $Y=1.07 $X2=0 $Y2=0
cc_196 N_Y_c_320_n N_VGND_M1007_s 5.90379e-19 $X=3.005 $Y=1.095 $X2=0 $Y2=0
cc_197 N_Y_c_322_n N_VGND_M1007_s 0.0033108f $X=3.12 $Y=1.095 $X2=0 $Y2=0
cc_198 N_Y_c_315_n N_VGND_c_369_n 0.0174504f $X=1.65 $Y=0.515 $X2=0 $Y2=0
cc_199 N_Y_c_315_n N_VGND_c_370_n 0.0173003f $X=1.65 $Y=0.515 $X2=0 $Y2=0
cc_200 N_Y_c_318_n N_VGND_c_370_n 0.0174872f $X=2.495 $Y=1.07 $X2=0 $Y2=0
cc_201 N_Y_c_319_n N_VGND_c_370_n 0.0164981f $X=2.58 $Y=0.515 $X2=0 $Y2=0
cc_202 N_Y_c_319_n N_VGND_c_372_n 0.0191439f $X=2.58 $Y=0.515 $X2=0 $Y2=0
cc_203 N_Y_c_320_n N_VGND_c_372_n 0.00254062f $X=3.005 $Y=1.095 $X2=0 $Y2=0
cc_204 N_Y_c_322_n N_VGND_c_372_n 0.0198092f $X=3.12 $Y=1.095 $X2=0 $Y2=0
cc_205 N_Y_c_315_n N_VGND_c_374_n 0.0145091f $X=1.65 $Y=0.515 $X2=0 $Y2=0
cc_206 N_Y_c_319_n N_VGND_c_375_n 0.011066f $X=2.58 $Y=0.515 $X2=0 $Y2=0
cc_207 N_Y_c_315_n N_VGND_c_378_n 0.0119768f $X=1.65 $Y=0.515 $X2=0 $Y2=0
cc_208 N_Y_c_319_n N_VGND_c_378_n 0.00915947f $X=2.58 $Y=0.515 $X2=0 $Y2=0
