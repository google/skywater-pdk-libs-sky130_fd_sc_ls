* File: sky130_fd_sc_ls__sedfxbp_2.spice
* Created: Wed Sep  2 11:29:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__sedfxbp_2.pex.spice"
.subckt sky130_fd_sc_ls__sedfxbp_2  VNB VPB D DE SCD SCE CLK VPWR Q Q_N VGND
* 
* VGND	VGND
* Q_N	Q_N
* Q	Q
* VPWR	VPWR
* CLK	CLK
* SCE	SCE
* SCD	SCD
* DE	DE
* D	D
* VPB	VPB
* VNB	VNB
MM1047 A_141_74# N_D_M1047_g N_A_32_74#_M1047_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.1659 PD=0.66 PS=1.63 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.3
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1042 N_VGND_M1042_d N_DE_M1042_g A_141_74# VNB NSHORT L=0.15 W=0.42 AD=0.1197
+ AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.7 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1028 N_VGND_M1028_d N_DE_M1028_g N_A_183_290#_M1028_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0735 AS=0.1197 PD=0.77 PS=1.41 NRD=19.992 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1024 A_527_113# N_A_183_290#_M1024_g N_VGND_M1028_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0735 PD=0.66 PS=0.77 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.7
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1006 N_A_32_74#_M1006_d N_A_575_87#_M1006_g A_527_113# VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.0504 PD=0.7 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8
+ SA=75001.1 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1010 N_A_691_113#_M1010_d N_A_661_87#_M1010_g N_A_32_74#_M1006_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.1491 AS=0.0588 PD=1.55 PS=0.7 NRD=19.992 NRS=0 M=1 R=2.8
+ SA=75001.5 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1039 N_VGND_M1039_d N_SCE_M1039_g N_A_661_87#_M1039_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0819 AS=0.1197 PD=0.81 PS=1.41 NRD=19.992 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1021 A_1091_125# N_SCD_M1021_g N_VGND_M1039_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0819 PD=0.66 PS=0.81 NRD=18.564 NRS=11.424 M=1 R=2.8 SA=75000.7
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1036 N_A_691_113#_M1036_d N_SCE_M1036_g A_1091_125# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1035 N_A_1374_368#_M1035_d N_CLK_M1035_g N_VGND_M1035_s VNB NSHORT L=0.15
+ W=0.74 AD=0.2109 AS=0.2627 PD=2.05 PS=2.19 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75000.3 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1003 N_A_1586_74#_M1003_d N_A_1374_368#_M1003_g N_VGND_M1003_s VNB NSHORT
+ L=0.15 W=0.74 AD=0.2109 AS=0.2109 PD=2.05 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1037 N_A_1784_97#_M1037_d N_A_1374_368#_M1037_g N_A_691_113#_M1037_s VNB
+ NSHORT L=0.15 W=0.42 AD=0.1113 AS=0.1197 PD=0.95 PS=1.41 NRD=71.424 NRS=0 M=1
+ R=2.8 SA=75000.2 SB=75002.3 A=0.063 P=1.14 MULT=1
MM1040 A_1920_97# N_A_1586_74#_M1040_g N_A_1784_97#_M1037_d VNB NSHORT L=0.15
+ W=0.42 AD=0.09765 AS=0.1113 PD=0.885 PS=0.95 NRD=50.712 NRS=0 M=1 R=2.8
+ SA=75000.9 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1034 N_VGND_M1034_d N_A_2013_71#_M1034_g A_1920_97# VNB NSHORT L=0.15 W=0.42
+ AD=0.136292 AS=0.09765 PD=0.990566 PS=0.885 NRD=24.276 NRS=50.712 M=1 R=2.8
+ SA=75001.5 SB=75001 A=0.063 P=1.14 MULT=1
MM1023 N_A_2013_71#_M1023_d N_A_1784_97#_M1023_g N_VGND_M1034_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.1824 AS=0.207683 PD=1.85 PS=1.50943 NRD=0 NRS=46.872 M=1
+ R=4.26667 SA=75001.6 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1009 A_2417_74# N_A_2013_71#_M1009_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0672 AS=0.1824 PD=0.85 PS=1.85 NRD=9.372 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75001.9 A=0.096 P=1.58 MULT=1
MM1011 N_A_2489_74#_M1011_d N_A_1586_74#_M1011_g A_2417_74# VNB NSHORT L=0.15
+ W=0.64 AD=0.129147 AS=0.0672 PD=1.20755 PS=0.85 NRD=0 NRS=9.372 M=1 R=4.26667
+ SA=75000.6 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1013 A_2591_74# N_A_1374_368#_M1013_g N_A_2489_74#_M1011_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.0847528 PD=0.66 PS=0.792453 NRD=18.564 NRS=23.568 M=1
+ R=2.8 SA=75001.1 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1026 N_VGND_M1026_d N_A_575_87#_M1026_g A_2591_74# VNB NSHORT L=0.15 W=0.42
+ AD=0.199681 AS=0.0504 PD=1.28534 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.5
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1014 N_A_575_87#_M1014_d N_A_2489_74#_M1014_g N_VGND_M1026_d VNB NSHORT L=0.15
+ W=0.74 AD=0.2109 AS=0.351819 PD=2.05 PS=2.26466 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1032 N_Q_M1032_d N_A_2489_74#_M1032_g N_VGND_M1032_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.5 A=0.111 P=1.78 MULT=1
MM1043 N_Q_M1032_d N_A_2489_74#_M1043_g N_VGND_M1043_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1027 N_Q_N_M1027_d N_A_575_87#_M1027_g N_VGND_M1043_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1041 N_Q_N_M1027_d N_A_575_87#_M1041_g N_VGND_M1041_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1004 A_132_464# N_D_M1004_g N_A_32_74#_M1004_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0864 AS=0.1888 PD=0.91 PS=1.87 NRD=24.625 NRS=3.0732 M=1 R=4.26667
+ SA=75000.2 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1029 N_VPWR_M1029_d N_A_183_290#_M1029_g A_132_464# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1888 AS=0.0864 PD=1.87 PS=0.91 NRD=3.0732 NRS=24.625 M=1 R=4.26667
+ SA=75000.6 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1017 N_VPWR_M1017_d N_DE_M1017_g N_A_183_290#_M1017_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1696 AS=0.1888 PD=1.17 PS=1.87 NRD=73.8553 NRS=3.0732 M=1
+ R=4.26667 SA=75000.2 SB=75001.7 A=0.096 P=1.58 MULT=1
MM1044 A_578_462# N_DE_M1044_g N_VPWR_M1017_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0768 AS=0.1696 PD=0.88 PS=1.17 NRD=19.9955 NRS=3.0732 M=1 R=4.26667
+ SA=75000.9 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1018 N_A_32_74#_M1018_d N_A_575_87#_M1018_g A_578_462# VPB PHIGHVT L=0.15
+ W=0.64 AD=0.096 AS=0.0768 PD=0.94 PS=0.88 NRD=3.0732 NRS=19.9955 M=1 R=4.26667
+ SA=75001.3 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1033 N_A_691_113#_M1033_d N_SCE_M1033_g N_A_32_74#_M1018_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1888 AS=0.096 PD=1.87 PS=0.94 NRD=3.0732 NRS=3.0732 M=1 R=4.26667
+ SA=75001.7 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1045 N_VPWR_M1045_d N_SCE_M1045_g N_A_661_87#_M1045_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1728 AS=0.1952 PD=1.18 PS=1.89 NRD=73.8553 NRS=6.1464 M=1
+ R=4.26667 SA=75000.2 SB=75001.3 A=0.096 P=1.58 MULT=1
MM1012 A_1088_453# N_SCD_M1012_g N_VPWR_M1045_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0864 AS=0.1728 PD=0.91 PS=1.18 NRD=24.625 NRS=6.1464 M=1 R=4.26667
+ SA=75000.9 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1000 N_A_691_113#_M1000_d N_A_661_87#_M1000_g A_1088_453# VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1888 AS=0.0864 PD=1.87 PS=0.91 NRD=3.0732 NRS=24.625 M=1 R=4.26667
+ SA=75001.3 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1007 N_A_1374_368#_M1007_d N_CLK_M1007_g N_VPWR_M1007_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.3304 AS=0.3304 PD=2.83 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1001 N_A_1586_74#_M1001_d N_A_1374_368#_M1001_g N_VPWR_M1001_s VPB PHIGHVT
+ L=0.15 W=1.12 AD=0.3304 AS=0.3304 PD=2.83 PS=2.83 NRD=1.7533 NRS=1.7533 M=1
+ R=7.46667 SA=75000.2 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1008 N_A_1784_97#_M1008_d N_A_1586_74#_M1008_g N_A_691_113#_M1008_s VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.063 AS=0.1239 PD=0.72 PS=1.43 NRD=4.6886 NRS=4.6886
+ M=1 R=2.8 SA=75000.2 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1019 A_1944_508# N_A_1374_368#_M1019_g N_A_1784_97#_M1008_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0756 AS=0.063 PD=0.78 PS=0.72 NRD=58.6272 NRS=4.6886 M=1 R=2.8
+ SA=75000.7 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1002 N_VPWR_M1002_d N_A_2013_71#_M1002_g A_1944_508# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0999833 AS=0.0756 PD=0.91 PS=0.78 NRD=9.3772 NRS=58.6272 M=1 R=2.8
+ SA=75001.2 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1030 N_A_2013_71#_M1030_d N_A_1784_97#_M1030_g N_VPWR_M1002_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.2478 AS=0.199967 PD=2.27 PS=1.82 NRD=2.3443 NRS=23.443 M=1
+ R=5.6 SA=75000.7 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1046 A_2374_392# N_A_2013_71#_M1046_g N_VPWR_M1046_s VPB PHIGHVT L=0.15 W=1
+ AD=0.4025 AS=0.4032 PD=1.805 PS=2.92 NRD=68.4378 NRS=19.6803 M=1 R=6.66667
+ SA=75000.3 SB=75001.9 A=0.15 P=2.3 MULT=1
MM1015 N_A_2489_74#_M1015_d N_A_1374_368#_M1015_g A_2374_392# VPB PHIGHVT L=0.15
+ W=1 AD=0.234366 AS=0.4025 PD=1.9507 PS=1.805 NRD=1.9503 NRS=68.4378 M=1
+ R=6.66667 SA=75001.3 SB=75000.9 A=0.15 P=2.3 MULT=1
MM1025 A_2672_508# N_A_1586_74#_M1025_g N_A_2489_74#_M1015_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0567 AS=0.0984338 PD=0.69 PS=0.819296 NRD=37.5088 NRS=44.5417 M=1
+ R=2.8 SA=75001.8 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1022 N_VPWR_M1022_d N_A_575_87#_M1022_g A_2672_508# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.114736 AS=0.0567 PD=0.916364 PS=0.69 NRD=53.9386 NRS=37.5088 M=1 R=2.8
+ SA=75002.2 SB=75000.9 A=0.063 P=1.14 MULT=1
MM1020 N_A_575_87#_M1020_d N_A_2489_74#_M1020_g N_VPWR_M1022_d VPB PHIGHVT
+ L=0.15 W=1.12 AD=0.3304 AS=0.305964 PD=2.83 PS=2.44364 NRD=1.7533 NRS=29.0181
+ M=1 R=7.46667 SA=75001.2 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1005 N_Q_M1005_d N_A_2489_74#_M1005_g N_VPWR_M1005_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1016 N_Q_M1005_d N_A_2489_74#_M1016_g N_VPWR_M1016_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1031 N_Q_N_M1031_d N_A_575_87#_M1031_g N_VPWR_M1016_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1038 N_Q_N_M1031_d N_A_575_87#_M1038_g N_VPWR_M1038_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.6 SB=75000.2 A=0.168 P=2.54 MULT=1
DX48_noxref VNB VPB NWDIODE A=32.8476 P=39.04
c_182 VNB 0 1.45871e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_ls__sedfxbp_2.pxi.spice"
*
.ends
*
*
