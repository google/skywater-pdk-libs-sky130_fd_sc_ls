* File: sky130_fd_sc_ls__and3b_2.pex.spice
* Created: Wed Sep  2 10:55:11 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__AND3B_2%A_N 2 5 7 9 10 13 14
r31 13 15 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.395 $Y=1.425
+ $X2=0.395 $Y2=1.26
r32 13 14 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.385
+ $Y=1.425 $X2=0.385 $Y2=1.425
r33 10 14 2.58853 $w=6.68e-07 $l=1.45e-07 $layer=LI1_cond $X=0.24 $Y=1.595
+ $X2=0.385 $Y2=1.595
r34 7 9 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.505 $Y=2.045
+ $X2=0.505 $Y2=2.54
r35 5 15 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=0.495 $Y=0.715
+ $X2=0.495 $Y2=1.26
r36 2 7 50.6449 $w=2.76e-07 $l=3.40588e-07 $layer=POLY_cond $X=0.395 $Y=1.755
+ $X2=0.505 $Y2=2.045
r37 1 13 1.64869 $w=3.5e-07 $l=1e-08 $layer=POLY_cond $X=0.395 $Y=1.435
+ $X2=0.395 $Y2=1.425
r38 1 2 52.7581 $w=3.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.395 $Y=1.435
+ $X2=0.395 $Y2=1.755
.ends

.subckt PM_SKY130_FD_SC_LS__AND3B_2%A_27_88# 1 2 7 9 11 12 14 15 18 22 23 24 29
+ 30 32 34 35
c67 9 0 1.29196e-19 $X=1.79 $Y=1.765
r68 32 35 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.985 $Y=2.1
+ $X2=0.985 $Y2=1.855
r69 29 30 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.065
+ $Y=1.35 $X2=1.065 $Y2=1.35
r70 27 35 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.065 $Y=1.69
+ $X2=1.065 $Y2=1.855
r71 27 29 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=1.065 $Y=1.69
+ $X2=1.065 $Y2=1.35
r72 26 29 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=1.065 $Y=1.09
+ $X2=1.065 $Y2=1.35
r73 25 34 4.64039 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=0.4 $Y=2.185
+ $X2=0.257 $Y2=2.185
r74 24 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.9 $Y=2.185
+ $X2=0.985 $Y2=2.1
r75 24 25 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=0.9 $Y=2.185 $X2=0.4
+ $Y2=2.185
r76 22 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.9 $Y=1.005
+ $X2=1.065 $Y2=1.09
r77 22 23 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=0.9 $Y=1.005
+ $X2=0.375 $Y2=1.005
r78 16 23 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.245 $Y=0.92
+ $X2=0.375 $Y2=1.005
r79 16 18 9.08657 $w=2.58e-07 $l=2.05e-07 $layer=LI1_cond $X=0.245 $Y=0.92
+ $X2=0.245 $Y2=0.715
r80 12 15 43.6107 $w=1.5e-07 $l=2.97405e-07 $layer=POLY_cond $X=1.805 $Y=1.185
+ $X2=1.79 $Y2=1.475
r81 12 14 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.805 $Y=1.185
+ $X2=1.805 $Y2=0.74
r82 9 15 43.6107 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=1.79 $Y=1.765
+ $X2=1.79 $Y2=1.475
r83 9 11 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.79 $Y=1.765
+ $X2=1.79 $Y2=2.34
r84 8 30 8.21848 $w=3.3e-07 $l=4.7e-08 $layer=POLY_cond $X=1.065 $Y=1.397
+ $X2=1.065 $Y2=1.35
r85 7 15 7.81274 $w=4.25e-07 $l=1.22963e-07 $layer=POLY_cond $X=1.7 $Y=1.397
+ $X2=1.79 $Y2=1.475
r86 7 8 61.5041 $w=4.25e-07 $l=4.7e-07 $layer=POLY_cond $X=1.7 $Y=1.397 $X2=1.23
+ $Y2=1.397
r87 2 34 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.12 $X2=0.28 $Y2=2.265
r88 1 18 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.44 $X2=0.28 $Y2=0.715
.ends

.subckt PM_SKY130_FD_SC_LS__AND3B_2%B 1 3 4 6 7 8 9 10
c36 7 0 1.29196e-19 $X=2.16 $Y=0.555
r37 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.285
+ $Y=1.385 $X2=2.285 $Y2=1.385
r38 10 17 7.96751 $w=4.03e-07 $l=2.8e-07 $layer=LI1_cond $X=2.247 $Y=1.665
+ $X2=2.247 $Y2=1.385
r39 9 17 2.56098 $w=4.03e-07 $l=9e-08 $layer=LI1_cond $X=2.247 $Y=1.295
+ $X2=2.247 $Y2=1.385
r40 8 9 10.5285 $w=4.03e-07 $l=3.7e-07 $layer=LI1_cond $X=2.247 $Y=0.925
+ $X2=2.247 $Y2=1.295
r41 7 8 10.5285 $w=4.03e-07 $l=3.7e-07 $layer=LI1_cond $X=2.247 $Y=0.555
+ $X2=2.247 $Y2=0.925
r42 4 16 77.2841 $w=2.7e-07 $l=4.15812e-07 $layer=POLY_cond $X=2.36 $Y=1.765
+ $X2=2.285 $Y2=1.385
r43 4 6 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.36 $Y=1.765
+ $X2=2.36 $Y2=2.34
r44 1 16 38.9026 $w=2.7e-07 $l=2.05122e-07 $layer=POLY_cond $X=2.195 $Y=1.22
+ $X2=2.285 $Y2=1.385
r45 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.195 $Y=1.22 $X2=2.195
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__AND3B_2%C 3 5 7 8
c33 8 0 1.28931e-19 $X=3.12 $Y=1.665
r34 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.855
+ $Y=1.515 $X2=2.855 $Y2=1.515
r35 8 12 7.10226 $w=4.28e-07 $l=2.65e-07 $layer=LI1_cond $X=3.12 $Y=1.565
+ $X2=2.855 $Y2=1.565
r36 5 11 52.2586 $w=2.99e-07 $l=2.7157e-07 $layer=POLY_cond $X=2.81 $Y=1.765
+ $X2=2.855 $Y2=1.515
r37 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.81 $Y=1.765
+ $X2=2.81 $Y2=2.34
r38 1 11 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=2.765 $Y=1.35
+ $X2=2.855 $Y2=1.515
r39 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.765 $Y=1.35
+ $X2=2.765 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__AND3B_2%A_284_368# 1 2 3 12 14 16 19 21 23 26 30 32
+ 36 38 41 43 46 49 56
c100 14 0 1.28931e-19 $X=3.35 $Y=1.765
r101 55 56 6.34211 $w=3.8e-07 $l=5e-08 $layer=POLY_cond $X=3.765 $Y=1.532
+ $X2=3.815 $Y2=1.532
r102 54 55 52.6395 $w=3.8e-07 $l=4.15e-07 $layer=POLY_cond $X=3.35 $Y=1.532
+ $X2=3.765 $Y2=1.532
r103 53 54 1.90263 $w=3.8e-07 $l=1.5e-08 $layer=POLY_cond $X=3.335 $Y=1.532
+ $X2=3.35 $Y2=1.532
r104 50 56 29.8079 $w=3.8e-07 $l=2.35e-07 $layer=POLY_cond $X=4.05 $Y=1.532
+ $X2=3.815 $Y2=1.532
r105 49 52 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.05 $Y=1.465
+ $X2=4.05 $Y2=1.63
r106 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.05
+ $Y=1.465 $X2=4.05 $Y2=1.465
r107 46 47 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=2.585 $Y=2.035
+ $X2=2.585 $Y2=2.325
r108 41 52 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=4.13 $Y=2.24
+ $X2=4.13 $Y2=1.63
r109 39 47 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.75 $Y=2.325
+ $X2=2.585 $Y2=2.325
r110 38 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.045 $Y=2.325
+ $X2=4.13 $Y2=2.24
r111 38 39 84.4866 $w=1.68e-07 $l=1.295e-06 $layer=LI1_cond $X=4.045 $Y=2.325
+ $X2=2.75 $Y2=2.325
r112 34 47 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=2.585 $Y=2.41
+ $X2=2.585 $Y2=2.325
r113 34 36 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=2.585 $Y=2.41
+ $X2=2.585 $Y2=2.715
r114 33 43 3.95098 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=1.755 $Y=2.035
+ $X2=1.577 $Y2=2.035
r115 32 46 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.42 $Y=2.035
+ $X2=2.585 $Y2=2.035
r116 32 33 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=2.42 $Y=2.035
+ $X2=1.755 $Y2=2.035
r117 28 43 2.79095 $w=3.42e-07 $l=9.0802e-08 $layer=LI1_cond $X=1.565 $Y=2.12
+ $X2=1.577 $Y2=2.035
r118 28 30 20.0804 $w=3.28e-07 $l=5.75e-07 $layer=LI1_cond $X=1.565 $Y=2.12
+ $X2=1.565 $Y2=2.695
r119 24 43 2.79095 $w=3.42e-07 $l=8.5e-08 $layer=LI1_cond $X=1.577 $Y=1.95
+ $X2=1.577 $Y2=2.035
r120 24 26 46.5847 $w=3.53e-07 $l=1.435e-06 $layer=LI1_cond $X=1.577 $Y=1.95
+ $X2=1.577 $Y2=0.515
r121 21 56 24.6126 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=3.815 $Y=1.765
+ $X2=3.815 $Y2=1.532
r122 21 23 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.815 $Y=1.765
+ $X2=3.815 $Y2=2.4
r123 17 55 24.6126 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=3.765 $Y=1.3
+ $X2=3.765 $Y2=1.532
r124 17 19 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.765 $Y=1.3
+ $X2=3.765 $Y2=0.74
r125 14 54 24.6126 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=3.35 $Y=1.765
+ $X2=3.35 $Y2=1.532
r126 14 16 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.35 $Y=1.765
+ $X2=3.35 $Y2=2.4
r127 10 53 24.6126 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=3.335 $Y=1.3
+ $X2=3.335 $Y2=1.532
r128 10 12 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.335 $Y=1.3
+ $X2=3.335 $Y2=0.74
r129 3 46 400 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=2.435
+ $Y=1.84 $X2=2.585 $Y2=2.035
r130 3 36 400 $w=1.7e-07 $l=9.47035e-07 $layer=licon1_PDIFF $count=1 $X=2.435
+ $Y=1.84 $X2=2.585 $Y2=2.715
r131 2 43 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.42
+ $Y=1.84 $X2=1.565 $Y2=1.985
r132 2 30 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.42
+ $Y=1.84 $X2=1.565 $Y2=2.695
r133 1 26 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=1.445
+ $Y=0.37 $X2=1.59 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__AND3B_2%VPWR 1 2 3 4 15 19 23 25 27 30 31 32 34 43
+ 47 53 56 60
r54 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r55 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r56 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r57 51 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r58 51 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r59 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r60 48 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.29 $Y=3.33
+ $X2=3.125 $Y2=3.33
r61 48 50 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=3.29 $Y=3.33 $X2=3.6
+ $Y2=3.33
r62 47 59 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=3.875 $Y=3.33
+ $X2=4.097 $Y2=3.33
r63 47 50 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3.875 $Y=3.33
+ $X2=3.6 $Y2=3.33
r64 46 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r65 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r66 43 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.96 $Y=3.33
+ $X2=3.125 $Y2=3.33
r67 43 45 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2.96 $Y=3.33 $X2=2.64
+ $Y2=3.33
r68 42 54 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r69 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r70 39 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.9 $Y=3.33
+ $X2=0.735 $Y2=3.33
r71 39 41 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=0.9 $Y=3.33 $X2=1.68
+ $Y2=3.33
r72 37 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r73 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r74 34 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.57 $Y=3.33
+ $X2=0.735 $Y2=3.33
r75 34 36 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.57 $Y=3.33
+ $X2=0.24 $Y2=3.33
r76 32 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r77 32 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r78 30 41 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=1.9 $Y=3.33 $X2=1.68
+ $Y2=3.33
r79 30 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.9 $Y=3.33
+ $X2=2.065 $Y2=3.33
r80 29 45 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=2.23 $Y=3.33
+ $X2=2.64 $Y2=3.33
r81 29 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.23 $Y=3.33
+ $X2=2.065 $Y2=3.33
r82 25 59 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=4.04 $Y=3.245
+ $X2=4.097 $Y2=3.33
r83 25 27 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=4.04 $Y=3.245
+ $X2=4.04 $Y2=2.715
r84 21 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.125 $Y=3.245
+ $X2=3.125 $Y2=3.33
r85 21 23 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=3.125 $Y=3.245
+ $X2=3.125 $Y2=2.715
r86 17 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.065 $Y=3.245
+ $X2=2.065 $Y2=3.33
r87 17 19 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=2.065 $Y=3.245
+ $X2=2.065 $Y2=2.375
r88 13 53 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.735 $Y=3.245
+ $X2=0.735 $Y2=3.33
r89 13 15 22.3504 $w=3.28e-07 $l=6.4e-07 $layer=LI1_cond $X=0.735 $Y=3.245
+ $X2=0.735 $Y2=2.605
r90 4 27 600 $w=1.7e-07 $l=9.47035e-07 $layer=licon1_PDIFF $count=1 $X=3.89
+ $Y=1.84 $X2=4.04 $Y2=2.715
r91 3 23 600 $w=1.7e-07 $l=9.87737e-07 $layer=licon1_PDIFF $count=1 $X=2.885
+ $Y=1.84 $X2=3.125 $Y2=2.715
r92 2 19 300 $w=1.7e-07 $l=6.27077e-07 $layer=licon1_PDIFF $count=2 $X=1.865
+ $Y=1.84 $X2=2.065 $Y2=2.375
r93 1 15 600 $w=1.7e-07 $l=5.57136e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=2.12 $X2=0.735 $Y2=2.605
.ends

.subckt PM_SKY130_FD_SC_LS__AND3B_2%X 1 2 9 12 13 14 15 28
r30 21 28 1.3969 $w=3.28e-07 $l=4e-08 $layer=LI1_cond $X=3.55 $Y=0.965 $X2=3.55
+ $Y2=0.925
r31 14 15 13.9805 $w=3.03e-07 $l=3.7e-07 $layer=LI1_cond $X=3.562 $Y=1.295
+ $X2=3.562 $Y2=1.665
r32 14 35 6.23453 $w=3.03e-07 $l=1.65e-07 $layer=LI1_cond $X=3.562 $Y=1.295
+ $X2=3.562 $Y2=1.13
r33 13 35 5.07898 $w=3.28e-07 $l=1.43e-07 $layer=LI1_cond $X=3.55 $Y=0.987
+ $X2=3.55 $Y2=1.13
r34 13 21 0.768295 $w=3.28e-07 $l=2.2e-08 $layer=LI1_cond $X=3.55 $Y=0.987
+ $X2=3.55 $Y2=0.965
r35 13 28 0.803218 $w=3.28e-07 $l=2.3e-08 $layer=LI1_cond $X=3.55 $Y=0.902
+ $X2=3.55 $Y2=0.925
r36 12 13 13.515 $w=3.28e-07 $l=3.87e-07 $layer=LI1_cond $X=3.55 $Y=0.515
+ $X2=3.55 $Y2=0.902
r37 10 15 5.85668 $w=3.03e-07 $l=1.55e-07 $layer=LI1_cond $X=3.562 $Y=1.82
+ $X2=3.562 $Y2=1.665
r38 9 10 5.69504 $w=3.43e-07 $l=1.65e-07 $layer=LI1_cond $X=3.582 $Y=1.985
+ $X2=3.582 $Y2=1.82
r39 2 9 600 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=1 $X=3.425
+ $Y=1.84 $X2=3.58 $Y2=1.985
r40 1 12 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.41
+ $Y=0.37 $X2=3.55 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__AND3B_2%VGND 1 2 3 12 16 18 20 23 24 25 27 39 44 48
r46 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r47 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r48 42 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r49 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r50 39 47 3.94362 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=3.895 $Y=0 $X2=4.107
+ $Y2=0
r51 39 41 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.895 $Y=0 $X2=3.6
+ $Y2=0
r52 38 42 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r53 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r54 35 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r55 34 37 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r56 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r57 32 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=0.71
+ $Y2=0
r58 32 34 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=1.2
+ $Y2=0
r59 30 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r60 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r61 27 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.71
+ $Y2=0
r62 27 29 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.24
+ $Y2=0
r63 25 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r64 25 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.2
+ $Y2=0
r65 23 37 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.815 $Y=0 $X2=2.64
+ $Y2=0
r66 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.815 $Y=0 $X2=2.98
+ $Y2=0
r67 22 41 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=3.145 $Y=0 $X2=3.6
+ $Y2=0
r68 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.145 $Y=0 $X2=2.98
+ $Y2=0
r69 18 47 3.19954 $w=2.5e-07 $l=1.22327e-07 $layer=LI1_cond $X=4.02 $Y=0.085
+ $X2=4.107 $Y2=0
r70 18 20 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=4.02 $Y=0.085
+ $X2=4.02 $Y2=0.515
r71 14 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.98 $Y=0.085
+ $X2=2.98 $Y2=0
r72 14 16 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.98 $Y=0.085
+ $X2=2.98 $Y2=0.515
r73 10 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0
r74 10 12 18.6835 $w=3.28e-07 $l=5.35e-07 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0.62
r75 3 20 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.84
+ $Y=0.37 $X2=3.98 $Y2=0.515
r76 2 16 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.84
+ $Y=0.37 $X2=2.98 $Y2=0.515
r77 1 12 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=0.57 $Y=0.44
+ $X2=0.71 $Y2=0.62
.ends

