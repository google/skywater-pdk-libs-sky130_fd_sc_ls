* File: sky130_fd_sc_ls__xnor3_2.pxi.spice
* Created: Wed Sep  2 11:30:39 2020
* 
x_PM_SKY130_FD_SC_LS__XNOR3_2%A_83_247# N_A_83_247#_M1007_d N_A_83_247#_M1000_d
+ N_A_83_247#_M1011_d N_A_83_247#_M1012_d N_A_83_247#_c_175_n
+ N_A_83_247#_M1008_g N_A_83_247#_M1009_g N_A_83_247#_c_177_n
+ N_A_83_247#_c_178_n N_A_83_247#_c_179_n N_A_83_247#_c_198_p
+ N_A_83_247#_c_259_p N_A_83_247#_c_193_p N_A_83_247#_c_199_p
+ N_A_83_247#_c_185_n N_A_83_247#_c_180_n N_A_83_247#_c_186_n
+ N_A_83_247#_c_187_n N_A_83_247#_c_181_n N_A_83_247#_c_182_n
+ N_A_83_247#_c_188_n PM_SKY130_FD_SC_LS__XNOR3_2%A_83_247#
x_PM_SKY130_FD_SC_LS__XNOR3_2%A N_A_M1007_g N_A_c_304_n N_A_M1011_g A
+ N_A_c_305_n PM_SKY130_FD_SC_LS__XNOR3_2%A
x_PM_SKY130_FD_SC_LS__XNOR3_2%A_397_21# N_A_397_21#_M1014_s N_A_397_21#_M1020_s
+ N_A_397_21#_M1002_g N_A_397_21#_c_346_n N_A_397_21#_c_347_n
+ N_A_397_21#_c_357_n N_A_397_21#_M1004_g N_A_397_21#_c_348_n
+ N_A_397_21#_c_349_n N_A_397_21#_M1000_g N_A_397_21#_c_351_n
+ N_A_397_21#_M1012_g N_A_397_21#_c_359_n N_A_397_21#_c_352_n
+ N_A_397_21#_c_353_n N_A_397_21#_c_371_n N_A_397_21#_c_360_n
+ N_A_397_21#_c_354_n N_A_397_21#_c_355_n PM_SKY130_FD_SC_LS__XNOR3_2%A_397_21#
x_PM_SKY130_FD_SC_LS__XNOR3_2%B N_B_M1018_g N_B_c_473_n N_B_c_474_n N_B_c_467_n
+ N_B_M1005_g N_B_c_477_n N_B_c_478_n N_B_c_468_n N_B_M1001_g N_B_c_480_n
+ N_B_c_481_n N_B_M1003_g N_B_c_483_n N_B_c_484_n N_B_M1014_g N_B_c_485_n
+ N_B_M1020_g N_B_c_486_n B N_B_c_471_n N_B_c_472_n
+ PM_SKY130_FD_SC_LS__XNOR3_2%B
x_PM_SKY130_FD_SC_LS__XNOR3_2%A_1027_48# N_A_1027_48#_M1010_s
+ N_A_1027_48#_M1017_s N_A_1027_48#_M1023_g N_A_1027_48#_c_604_n
+ N_A_1027_48#_M1021_g N_A_1027_48#_c_605_n N_A_1027_48#_c_606_n
+ N_A_1027_48#_c_611_n N_A_1027_48#_c_607_n N_A_1027_48#_c_608_n
+ N_A_1027_48#_c_613_n PM_SKY130_FD_SC_LS__XNOR3_2%A_1027_48#
x_PM_SKY130_FD_SC_LS__XNOR3_2%C N_C_c_679_n N_C_M1019_g N_C_c_680_n N_C_c_681_n
+ N_C_c_682_n N_C_c_683_n N_C_c_689_n N_C_M1016_g N_C_c_684_n N_C_c_685_n
+ N_C_M1010_g N_C_c_686_n N_C_M1017_g C N_C_c_687_n
+ PM_SKY130_FD_SC_LS__XNOR3_2%C
x_PM_SKY130_FD_SC_LS__XNOR3_2%A_1057_74# N_A_1057_74#_M1023_d
+ N_A_1057_74#_M1021_d N_A_1057_74#_c_772_n N_A_1057_74#_M1013_g
+ N_A_1057_74#_c_762_n N_A_1057_74#_M1006_g N_A_1057_74#_c_773_n
+ N_A_1057_74#_M1022_g N_A_1057_74#_c_763_n N_A_1057_74#_M1015_g
+ N_A_1057_74#_c_791_n N_A_1057_74#_c_764_n N_A_1057_74#_c_765_n
+ N_A_1057_74#_c_774_n N_A_1057_74#_c_766_n N_A_1057_74#_c_767_n
+ N_A_1057_74#_c_768_n N_A_1057_74#_c_862_p N_A_1057_74#_c_775_n
+ N_A_1057_74#_c_802_n N_A_1057_74#_c_804_n N_A_1057_74#_c_816_p
+ N_A_1057_74#_c_788_n N_A_1057_74#_c_776_n N_A_1057_74#_c_777_n
+ N_A_1057_74#_c_769_n N_A_1057_74#_c_770_n N_A_1057_74#_c_771_n
+ PM_SKY130_FD_SC_LS__XNOR3_2%A_1057_74#
x_PM_SKY130_FD_SC_LS__XNOR3_2%A_27_373# N_A_27_373#_M1009_s N_A_27_373#_M1002_d
+ N_A_27_373#_M1008_s N_A_27_373#_M1004_d N_A_27_373#_c_884_n
+ N_A_27_373#_c_885_n N_A_27_373#_c_886_n N_A_27_373#_c_887_n
+ N_A_27_373#_c_895_n N_A_27_373#_c_896_n N_A_27_373#_c_897_n
+ N_A_27_373#_c_888_n N_A_27_373#_c_898_n N_A_27_373#_c_889_n
+ N_A_27_373#_c_890_n N_A_27_373#_c_891_n N_A_27_373#_c_892_n
+ N_A_27_373#_c_893_n PM_SKY130_FD_SC_LS__XNOR3_2%A_27_373#
x_PM_SKY130_FD_SC_LS__XNOR3_2%VPWR N_VPWR_M1008_d N_VPWR_M1020_d N_VPWR_M1017_d
+ N_VPWR_M1022_s N_VPWR_c_990_n N_VPWR_c_991_n N_VPWR_c_992_n N_VPWR_c_993_n
+ N_VPWR_c_994_n VPWR N_VPWR_c_995_n N_VPWR_c_996_n N_VPWR_c_997_n
+ N_VPWR_c_998_n N_VPWR_c_999_n N_VPWR_c_1000_n N_VPWR_c_989_n
+ PM_SKY130_FD_SC_LS__XNOR3_2%VPWR
x_PM_SKY130_FD_SC_LS__XNOR3_2%A_332_373# N_A_332_373#_M1001_d
+ N_A_332_373#_M1019_d N_A_332_373#_M1005_d N_A_332_373#_M1021_s
+ N_A_332_373#_c_1083_n N_A_332_373#_c_1072_n N_A_332_373#_c_1073_n
+ N_A_332_373#_c_1074_n N_A_332_373#_c_1075_n N_A_332_373#_c_1076_n
+ N_A_332_373#_c_1077_n N_A_332_373#_c_1078_n N_A_332_373#_c_1087_n
+ N_A_332_373#_c_1079_n N_A_332_373#_c_1080_n N_A_332_373#_c_1081_n
+ N_A_332_373#_c_1082_n PM_SKY130_FD_SC_LS__XNOR3_2%A_332_373#
x_PM_SKY130_FD_SC_LS__XNOR3_2%A_329_81# N_A_329_81#_M1018_d N_A_329_81#_M1023_s
+ N_A_329_81#_M1003_d N_A_329_81#_M1016_d N_A_329_81#_c_1183_n
+ N_A_329_81#_c_1211_n N_A_329_81#_c_1189_n N_A_329_81#_c_1190_n
+ N_A_329_81#_c_1184_n N_A_329_81#_c_1185_n N_A_329_81#_c_1192_n
+ N_A_329_81#_c_1193_n N_A_329_81#_c_1186_n N_A_329_81#_c_1187_n
+ N_A_329_81#_c_1188_n N_A_329_81#_c_1246_n
+ PM_SKY130_FD_SC_LS__XNOR3_2%A_329_81#
x_PM_SKY130_FD_SC_LS__XNOR3_2%X N_X_M1006_d N_X_M1013_d N_X_c_1312_n
+ N_X_c_1313_n N_X_c_1310_n X X X PM_SKY130_FD_SC_LS__XNOR3_2%X
x_PM_SKY130_FD_SC_LS__XNOR3_2%VGND N_VGND_M1009_d N_VGND_M1014_d N_VGND_M1010_d
+ N_VGND_M1015_s N_VGND_c_1343_n N_VGND_c_1344_n N_VGND_c_1345_n N_VGND_c_1346_n
+ N_VGND_c_1347_n VGND N_VGND_c_1348_n N_VGND_c_1349_n N_VGND_c_1350_n
+ N_VGND_c_1351_n N_VGND_c_1352_n N_VGND_c_1353_n N_VGND_c_1354_n
+ PM_SKY130_FD_SC_LS__XNOR3_2%VGND
cc_1 VNB N_A_83_247#_c_175_n 0.0404635f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.79
cc_2 VNB N_A_83_247#_M1009_g 0.0240792f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=0.725
cc_3 VNB N_A_83_247#_c_177_n 0.00193372f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.36
cc_4 VNB N_A_83_247#_c_178_n 6.25663e-19 $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.4
cc_5 VNB N_A_83_247#_c_179_n 0.00535503f $X=-0.19 $Y=-0.245 $X2=1.095 $Y2=1.12
cc_6 VNB N_A_83_247#_c_180_n 0.00209465f $X=-0.19 $Y=-0.245 $X2=1.345 $Y2=0.34
cc_7 VNB N_A_83_247#_c_181_n 0.00538013f $X=-0.19 $Y=-0.245 $X2=3.365 $Y2=0.36
cc_8 VNB N_A_83_247#_c_182_n 0.0208851f $X=-0.19 $Y=-0.245 $X2=3.2 $Y2=0.35
cc_9 VNB N_A_M1007_g 0.0268525f $X=-0.19 $Y=-0.245 $X2=1.12 $Y2=1.865
cc_10 VNB N_A_c_304_n 0.0232609f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_c_305_n 0.00334759f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_397_21#_M1002_g 0.0385893f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_397_21#_c_346_n 0.0171761f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_397_21#_c_347_n 0.00877638f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_397_21#_c_348_n 0.0693021f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.235
cc_16 VNB N_A_397_21#_c_349_n 0.012806f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=0.725
cc_17 VNB N_A_397_21#_M1000_g 0.0373065f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.95
cc_18 VNB N_A_397_21#_c_351_n 0.033559f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.4
cc_19 VNB N_A_397_21#_c_352_n 8.62302e-19 $X=-0.19 $Y=-0.245 $X2=1.235 $Y2=2.12
cc_20 VNB N_A_397_21#_c_353_n 0.00521129f $X=-0.19 $Y=-0.245 $X2=3.2 $Y2=0.34
cc_21 VNB N_A_397_21#_c_354_n 0.00440373f $X=-0.19 $Y=-0.245 $X2=3.365 $Y2=0.35
cc_22 VNB N_A_397_21#_c_355_n 0.00404841f $X=-0.19 $Y=-0.245 $X2=3.2 $Y2=0.35
cc_23 VNB N_B_M1018_g 0.0344444f $X=-0.19 $Y=-0.245 $X2=1.12 $Y2=1.865
cc_24 VNB N_B_c_467_n 0.00920414f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_B_c_468_n 0.0135715f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.79
cc_26 VNB N_B_M1001_g 0.0212321f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.365
cc_27 VNB N_B_M1014_g 0.025787f $X=-0.19 $Y=-0.245 $X2=1.22 $Y2=0.425
cc_28 VNB N_B_c_471_n 0.0515765f $X=-0.19 $Y=-0.245 $X2=1.28 $Y2=2.115
cc_29 VNB N_B_c_472_n 0.0030506f $X=-0.19 $Y=-0.245 $X2=3.365 $Y2=0.35
cc_30 VNB N_A_1027_48#_M1023_g 0.0450805f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_1027_48#_c_604_n 0.0269945f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_1027_48#_c_605_n 0.00182968f $X=-0.19 $Y=-0.245 $X2=0.505
+ $Y2=2.365
cc_33 VNB N_A_1027_48#_c_606_n 0.00260252f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.36
cc_34 VNB N_A_1027_48#_c_607_n 0.00161761f $X=-0.19 $Y=-0.245 $X2=1.095
+ $Y2=2.035
cc_35 VNB N_A_1027_48#_c_608_n 9.42831e-19 $X=-0.19 $Y=-0.245 $X2=1.22 $Y2=1.035
cc_36 VNB N_C_c_679_n 0.0175588f $X=-0.19 $Y=-0.245 $X2=1.12 $Y2=0.405
cc_37 VNB N_C_c_680_n 0.0115589f $X=-0.19 $Y=-0.245 $X2=3.28 $Y2=1.865
cc_38 VNB N_C_c_681_n 0.00905308f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_C_c_682_n 0.0295931f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_C_c_683_n 0.00372515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_C_c_684_n 0.0409078f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_C_c_685_n 0.0222798f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.79
cc_43 VNB N_C_c_686_n 0.0351571f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.235
cc_44 VNB N_C_c_687_n 0.00330598f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=1.12
cc_45 VNB N_A_1057_74#_c_762_n 0.0170165f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_1057_74#_c_763_n 0.0188693f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.235
cc_47 VNB N_A_1057_74#_c_764_n 0.0163721f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.4
cc_48 VNB N_A_1057_74#_c_765_n 0.00383604f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.4
cc_49 VNB N_A_1057_74#_c_766_n 0.0104484f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=2.035
cc_50 VNB N_A_1057_74#_c_767_n 0.00552332f $X=-0.19 $Y=-0.245 $X2=1.22 $Y2=0.425
cc_51 VNB N_A_1057_74#_c_768_n 0.00315591f $X=-0.19 $Y=-0.245 $X2=1.22 $Y2=1.035
cc_52 VNB N_A_1057_74#_c_769_n 0.00443367f $X=-0.19 $Y=-0.245 $X2=3.51 $Y2=2.99
cc_53 VNB N_A_1057_74#_c_770_n 0.00228435f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.4
cc_54 VNB N_A_1057_74#_c_771_n 0.0649881f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_27_373#_c_884_n 0.0241546f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.365
cc_56 VNB N_A_27_373#_c_885_n 6.56034e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_27_373#_c_886_n 0.00263335f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.36
cc_58 VNB N_A_27_373#_c_887_n 0.00475524f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.95
cc_59 VNB N_A_27_373#_c_888_n 0.00770296f $X=-0.19 $Y=-0.245 $X2=1.22 $Y2=1.035
cc_60 VNB N_A_27_373#_c_889_n 0.00157907f $X=-0.19 $Y=-0.245 $X2=1.345 $Y2=0.34
cc_61 VNB N_A_27_373#_c_890_n 0.0203735f $X=-0.19 $Y=-0.245 $X2=1.235 $Y2=2.035
cc_62 VNB N_A_27_373#_c_891_n 0.0033312f $X=-0.19 $Y=-0.245 $X2=1.28 $Y2=2.115
cc_63 VNB N_A_27_373#_c_892_n 0.029419f $X=-0.19 $Y=-0.245 $X2=3.2 $Y2=0.35
cc_64 VNB N_A_27_373#_c_893_n 0.00459486f $X=-0.19 $Y=-0.245 $X2=3.51 $Y2=2.795
cc_65 VNB N_VPWR_c_989_n 0.362705f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_332_373#_c_1072_n 0.00567041f $X=-0.19 $Y=-0.245 $X2=0.535
+ $Y2=0.725
cc_67 VNB N_A_332_373#_c_1073_n 0.00249128f $X=-0.19 $Y=-0.245 $X2=0.535
+ $Y2=0.725
cc_68 VNB N_A_332_373#_c_1074_n 0.00300639f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_332_373#_c_1075_n 0.00255368f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.36
cc_70 VNB N_A_332_373#_c_1076_n 0.0112843f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.95
cc_71 VNB N_A_332_373#_c_1077_n 0.00652094f $X=-0.19 $Y=-0.245 $X2=1.095
+ $Y2=1.12
cc_72 VNB N_A_332_373#_c_1078_n 0.00257282f $X=-0.19 $Y=-0.245 $X2=1.22 $Y2=0.55
cc_73 VNB N_A_332_373#_c_1079_n 0.0262647f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.12
cc_74 VNB N_A_332_373#_c_1080_n 0.00286242f $X=-0.19 $Y=-0.245 $X2=1.235
+ $Y2=2.035
cc_75 VNB N_A_332_373#_c_1081_n 0.00185916f $X=-0.19 $Y=-0.245 $X2=3.365
+ $Y2=0.36
cc_76 VNB N_A_332_373#_c_1082_n 0.00202343f $X=-0.19 $Y=-0.245 $X2=3.51
+ $Y2=2.795
cc_77 VNB N_A_329_81#_c_1183_n 0.009648f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.365
cc_78 VNB N_A_329_81#_c_1184_n 0.0164249f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.4
cc_79 VNB N_A_329_81#_c_1185_n 0.0153705f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.4
cc_80 VNB N_A_329_81#_c_1186_n 0.00141657f $X=-0.19 $Y=-0.245 $X2=1.22 $Y2=0.55
cc_81 VNB N_A_329_81#_c_1187_n 0.00408737f $X=-0.19 $Y=-0.245 $X2=1.345 $Y2=0.34
cc_82 VNB N_A_329_81#_c_1188_n 6.99046e-19 $X=-0.19 $Y=-0.245 $X2=3.345 $Y2=2.99
cc_83 VNB N_X_c_1310_n 0.00115496f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.365
cc_84 VNB X 0.00279061f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.235
cc_85 VNB N_VGND_c_1343_n 0.0080712f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.365
cc_86 VNB N_VGND_c_1344_n 0.0123225f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1345_n 0.0566416f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.95
cc_88 VNB N_VGND_c_1346_n 0.010678f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.4
cc_89 VNB N_VGND_c_1347_n 0.0540788f $X=-0.19 $Y=-0.245 $X2=1.095 $Y2=1.12
cc_90 VNB N_VGND_c_1348_n 0.0184398f $X=-0.19 $Y=-0.245 $X2=1.22 $Y2=0.425
cc_91 VNB N_VGND_c_1349_n 0.0801099f $X=-0.19 $Y=-0.245 $X2=1.235 $Y2=2.905
cc_92 VNB N_VGND_c_1350_n 0.0197463f $X=-0.19 $Y=-0.245 $X2=3.365 $Y2=0.35
cc_93 VNB N_VGND_c_1351_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_VGND_c_1352_n 0.00631318f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.4
cc_95 VNB N_VGND_c_1353_n 0.0297566f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_VGND_c_1354_n 0.466708f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VPB N_A_83_247#_c_175_n 0.0272324f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.79
cc_98 VPB N_A_83_247#_c_178_n 0.00168018f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=1.4
cc_99 VPB N_A_83_247#_c_185_n 4.07879e-19 $X=-0.19 $Y=1.66 $X2=1.235 $Y2=2.905
cc_100 VPB N_A_83_247#_c_186_n 0.0344487f $X=-0.19 $Y=1.66 $X2=3.345 $Y2=2.99
cc_101 VPB N_A_83_247#_c_187_n 0.00288386f $X=-0.19 $Y=1.66 $X2=1.375 $Y2=2.99
cc_102 VPB N_A_83_247#_c_188_n 0.0087718f $X=-0.19 $Y=1.66 $X2=3.51 $Y2=2.795
cc_103 VPB N_A_c_304_n 0.0288224f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB N_A_c_305_n 0.0024708f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_105 VPB N_A_397_21#_c_347_n 0.00200104f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_A_397_21#_c_357_n 0.0211628f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.79
cc_107 VPB N_A_397_21#_c_351_n 0.0341272f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=1.4
cc_108 VPB N_A_397_21#_c_359_n 0.00272795f $X=-0.19 $Y=1.66 $X2=1.26 $Y2=0.55
cc_109 VPB N_A_397_21#_c_360_n 0.00318289f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=1.12
cc_110 VPB N_A_397_21#_c_354_n 0.00197208f $X=-0.19 $Y=1.66 $X2=3.365 $Y2=0.35
cc_111 VPB N_B_c_473_n 0.00917565f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_B_c_474_n 0.0148771f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_B_c_467_n 0.00872715f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_B_M1005_g 0.0100136f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_B_c_477_n 0.0602821f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_B_c_478_n 0.0140969f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_B_c_468_n 0.00813311f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.79
cc_118 VPB N_B_c_480_n 0.00677815f $X=-0.19 $Y=1.66 $X2=0.535 $Y2=0.725
cc_119 VPB N_B_c_481_n 0.0332401f $X=-0.19 $Y=1.66 $X2=0.535 $Y2=0.725
cc_120 VPB N_B_M1003_g 0.00832021f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=1.4
cc_121 VPB N_B_c_483_n 0.0788088f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=1.4
cc_122 VPB N_B_c_484_n 0.0795247f $X=-0.19 $Y=1.66 $X2=0.745 $Y2=1.12
cc_123 VPB N_B_c_485_n 0.0170968f $X=-0.19 $Y=1.66 $X2=1.22 $Y2=0.55
cc_124 VPB N_B_c_486_n 0.00898834f $X=-0.19 $Y=1.66 $X2=3.2 $Y2=0.34
cc_125 VPB N_B_c_471_n 0.0180797f $X=-0.19 $Y=1.66 $X2=1.28 $Y2=2.115
cc_126 VPB N_B_c_472_n 0.00376962f $X=-0.19 $Y=1.66 $X2=3.365 $Y2=0.35
cc_127 VPB N_A_1027_48#_c_604_n 0.050405f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_A_1027_48#_c_605_n 0.0093761f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.365
cc_129 VPB N_A_1027_48#_c_611_n 0.0116878f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=1.4
cc_130 VPB N_A_1027_48#_c_608_n 0.00702052f $X=-0.19 $Y=1.66 $X2=1.22 $Y2=1.035
cc_131 VPB N_A_1027_48#_c_613_n 0.00279714f $X=-0.19 $Y=1.66 $X2=1.22 $Y2=0.55
cc_132 VPB N_C_c_683_n 0.0102901f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_C_c_689_n 0.026501f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_C_c_686_n 0.0347077f $X=-0.19 $Y=1.66 $X2=0.535 $Y2=1.235
cc_135 VPB N_C_c_687_n 0.00528748f $X=-0.19 $Y=1.66 $X2=0.745 $Y2=1.12
cc_136 VPB N_A_1057_74#_c_772_n 0.0166918f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_A_1057_74#_c_773_n 0.0174317f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.79
cc_138 VPB N_A_1057_74#_c_774_n 0.0346042f $X=-0.19 $Y=1.66 $X2=1.095 $Y2=1.12
cc_139 VPB N_A_1057_74#_c_775_n 0.0137001f $X=-0.19 $Y=1.66 $X2=1.235 $Y2=2.905
cc_140 VPB N_A_1057_74#_c_776_n 0.00275108f $X=-0.19 $Y=1.66 $X2=3.365 $Y2=0.35
cc_141 VPB N_A_1057_74#_c_777_n 0.00987431f $X=-0.19 $Y=1.66 $X2=3.2 $Y2=0.35
cc_142 VPB N_A_1057_74#_c_769_n 8.15627e-19 $X=-0.19 $Y=1.66 $X2=3.51 $Y2=2.99
cc_143 VPB N_A_1057_74#_c_771_n 0.022501f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_144 VPB N_A_27_373#_c_886_n 0.00137656f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=1.36
cc_145 VPB N_A_27_373#_c_895_n 0.00764312f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=1.4
cc_146 VPB N_A_27_373#_c_896_n 4.01397e-19 $X=-0.19 $Y=1.66 $X2=0.58 $Y2=1.4
cc_147 VPB N_A_27_373#_c_897_n 4.52711e-19 $X=-0.19 $Y=1.66 $X2=1.095 $Y2=2.035
cc_148 VPB N_A_27_373#_c_898_n 0.0269797f $X=-0.19 $Y=1.66 $X2=1.235 $Y2=2.12
cc_149 VPB N_A_27_373#_c_892_n 0.0262582f $X=-0.19 $Y=1.66 $X2=3.2 $Y2=0.35
cc_150 VPB N_VPWR_c_990_n 0.0138363f $X=-0.19 $Y=1.66 $X2=0.535 $Y2=0.725
cc_151 VPB N_VPWR_c_991_n 0.0160933f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=1.95
cc_152 VPB N_VPWR_c_992_n 0.00831246f $X=-0.19 $Y=1.66 $X2=1.095 $Y2=1.12
cc_153 VPB N_VPWR_c_993_n 0.0104926f $X=-0.19 $Y=1.66 $X2=1.095 $Y2=2.035
cc_154 VPB N_VPWR_c_994_n 0.0587528f $X=-0.19 $Y=1.66 $X2=1.22 $Y2=0.425
cc_155 VPB N_VPWR_c_995_n 0.0877154f $X=-0.19 $Y=1.66 $X2=3.2 $Y2=0.34
cc_156 VPB N_VPWR_c_996_n 0.0667808f $X=-0.19 $Y=1.66 $X2=3.365 $Y2=0.36
cc_157 VPB N_VPWR_c_997_n 0.0204869f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_158 VPB N_VPWR_c_998_n 0.0257077f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_159 VPB N_VPWR_c_999_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_160 VPB N_VPWR_c_1000_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_161 VPB N_VPWR_c_989_n 0.104008f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_162 VPB N_A_332_373#_c_1083_n 0.00243376f $X=-0.19 $Y=1.66 $X2=0.505
+ $Y2=2.365
cc_163 VPB N_A_332_373#_c_1072_n 0.00320013f $X=-0.19 $Y=1.66 $X2=0.535
+ $Y2=0.725
cc_164 VPB N_A_332_373#_c_1073_n 4.66474e-19 $X=-0.19 $Y=1.66 $X2=0.535
+ $Y2=0.725
cc_165 VPB N_A_332_373#_c_1075_n 0.00496772f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=1.36
cc_166 VPB N_A_332_373#_c_1087_n 0.00582446f $X=-0.19 $Y=1.66 $X2=3.345 $Y2=2.99
cc_167 VPB N_A_329_81#_c_1189_n 0.00355392f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=1.95
cc_168 VPB N_A_329_81#_c_1190_n 7.38419e-19 $X=-0.19 $Y=1.66 $X2=0.62 $Y2=1.4
cc_169 VPB N_A_329_81#_c_1185_n 0.00366751f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=1.4
cc_170 VPB N_A_329_81#_c_1192_n 0.0124642f $X=-0.19 $Y=1.66 $X2=1.095 $Y2=1.12
cc_171 VPB N_A_329_81#_c_1193_n 0.00186348f $X=-0.19 $Y=1.66 $X2=1.22 $Y2=0.425
cc_172 VPB N_X_c_1312_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_173 VPB N_X_c_1313_n 9.54502e-19 $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.365
cc_174 VPB N_X_c_1310_n 9.68834e-19 $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.365
cc_175 N_A_83_247#_c_175_n N_A_M1007_g 0.00862331f $X=0.505 $Y=1.79 $X2=0 $Y2=0
cc_176 N_A_83_247#_M1009_g N_A_M1007_g 0.0220707f $X=0.535 $Y=0.725 $X2=0 $Y2=0
cc_177 N_A_83_247#_c_177_n N_A_M1007_g 0.00186641f $X=0.62 $Y=1.36 $X2=0 $Y2=0
cc_178 N_A_83_247#_c_179_n N_A_M1007_g 0.0139401f $X=1.095 $Y=1.12 $X2=0 $Y2=0
cc_179 N_A_83_247#_c_193_p N_A_M1007_g 0.00778962f $X=1.26 $Y=0.55 $X2=0 $Y2=0
cc_180 N_A_83_247#_c_180_n N_A_M1007_g 0.00383348f $X=1.345 $Y=0.34 $X2=0 $Y2=0
cc_181 N_A_83_247#_c_175_n N_A_c_304_n 0.0431097f $X=0.505 $Y=1.79 $X2=0 $Y2=0
cc_182 N_A_83_247#_c_178_n N_A_c_304_n 0.00589127f $X=0.58 $Y=1.4 $X2=0 $Y2=0
cc_183 N_A_83_247#_c_179_n N_A_c_304_n 0.00140382f $X=1.095 $Y=1.12 $X2=0 $Y2=0
cc_184 N_A_83_247#_c_198_p N_A_c_304_n 0.0116599f $X=1.095 $Y=2.035 $X2=0 $Y2=0
cc_185 N_A_83_247#_c_199_p N_A_c_304_n 0.00159742f $X=1.235 $Y=2.12 $X2=0 $Y2=0
cc_186 N_A_83_247#_c_185_n N_A_c_304_n 0.0127913f $X=1.235 $Y=2.905 $X2=0 $Y2=0
cc_187 N_A_83_247#_c_187_n N_A_c_304_n 0.00264858f $X=1.375 $Y=2.99 $X2=0 $Y2=0
cc_188 N_A_83_247#_c_175_n N_A_c_305_n 8.83049e-19 $X=0.505 $Y=1.79 $X2=0 $Y2=0
cc_189 N_A_83_247#_c_178_n N_A_c_305_n 0.0260663f $X=0.58 $Y=1.4 $X2=0 $Y2=0
cc_190 N_A_83_247#_c_179_n N_A_c_305_n 0.0225458f $X=1.095 $Y=1.12 $X2=0 $Y2=0
cc_191 N_A_83_247#_c_198_p N_A_c_305_n 0.00941924f $X=1.095 $Y=2.035 $X2=0 $Y2=0
cc_192 N_A_83_247#_c_199_p N_A_c_305_n 0.0161536f $X=1.235 $Y=2.12 $X2=0 $Y2=0
cc_193 N_A_83_247#_c_182_n N_A_397_21#_M1002_g 0.012253f $X=3.2 $Y=0.35 $X2=0
+ $Y2=0
cc_194 N_A_83_247#_c_186_n N_A_397_21#_c_357_n 4.1597e-19 $X=3.345 $Y=2.99 $X2=0
+ $Y2=0
cc_195 N_A_83_247#_c_182_n N_A_397_21#_c_348_n 0.0135339f $X=3.2 $Y=0.35 $X2=0
+ $Y2=0
cc_196 N_A_83_247#_c_181_n N_A_397_21#_M1000_g 8.00488e-19 $X=3.365 $Y=0.36
+ $X2=0 $Y2=0
cc_197 N_A_83_247#_c_182_n N_A_397_21#_M1000_g 0.0134669f $X=3.2 $Y=0.35 $X2=0
+ $Y2=0
cc_198 N_A_83_247#_c_186_n N_A_397_21#_c_351_n 0.00155688f $X=3.345 $Y=2.99
+ $X2=0 $Y2=0
cc_199 N_A_83_247#_c_188_n N_A_397_21#_c_351_n 0.00359571f $X=3.51 $Y=2.795
+ $X2=0 $Y2=0
cc_200 N_A_83_247#_M1012_d N_A_397_21#_c_359_n 0.00231783f $X=3.28 $Y=1.865
+ $X2=0 $Y2=0
cc_201 N_A_83_247#_M1000_d N_A_397_21#_c_352_n 0.00454958f $X=3.145 $Y=0.625
+ $X2=0 $Y2=0
cc_202 N_A_83_247#_M1012_d N_A_397_21#_c_371_n 0.00640721f $X=3.28 $Y=1.865
+ $X2=0 $Y2=0
cc_203 N_A_83_247#_M1012_d N_A_397_21#_c_360_n 0.00266017f $X=3.28 $Y=1.865
+ $X2=0 $Y2=0
cc_204 N_A_83_247#_M1000_d N_A_397_21#_c_355_n 0.00205319f $X=3.145 $Y=0.625
+ $X2=0 $Y2=0
cc_205 N_A_83_247#_c_179_n N_B_M1018_g 0.00412463f $X=1.095 $Y=1.12 $X2=0 $Y2=0
cc_206 N_A_83_247#_c_193_p N_B_M1018_g 0.00833237f $X=1.26 $Y=0.55 $X2=0 $Y2=0
cc_207 N_A_83_247#_c_182_n N_B_M1018_g 0.0145029f $X=3.2 $Y=0.35 $X2=0 $Y2=0
cc_208 N_A_83_247#_c_185_n N_B_c_473_n 0.00316116f $X=1.235 $Y=2.905 $X2=0 $Y2=0
cc_209 N_A_83_247#_c_186_n N_B_c_474_n 0.0152848f $X=3.345 $Y=2.99 $X2=0 $Y2=0
cc_210 N_A_83_247#_c_199_p N_B_M1005_g 0.00136921f $X=1.235 $Y=2.12 $X2=0 $Y2=0
cc_211 N_A_83_247#_c_185_n N_B_M1005_g 0.0056749f $X=1.235 $Y=2.905 $X2=0 $Y2=0
cc_212 N_A_83_247#_c_186_n N_B_c_477_n 0.0148918f $X=3.345 $Y=2.99 $X2=0 $Y2=0
cc_213 N_A_83_247#_c_182_n N_B_M1001_g 0.00116683f $X=3.2 $Y=0.35 $X2=0 $Y2=0
cc_214 N_A_83_247#_c_186_n N_B_c_481_n 0.0193481f $X=3.345 $Y=2.99 $X2=0 $Y2=0
cc_215 N_A_83_247#_c_188_n N_B_c_481_n 0.0023392f $X=3.51 $Y=2.795 $X2=0 $Y2=0
cc_216 N_A_83_247#_c_186_n N_B_c_483_n 0.00930692f $X=3.345 $Y=2.99 $X2=0 $Y2=0
cc_217 N_A_83_247#_c_188_n N_B_c_483_n 0.00889438f $X=3.51 $Y=2.795 $X2=0 $Y2=0
cc_218 N_A_83_247#_c_188_n N_B_c_484_n 0.0137952f $X=3.51 $Y=2.795 $X2=0 $Y2=0
cc_219 N_A_83_247#_c_181_n N_B_M1014_g 0.00356999f $X=3.365 $Y=0.36 $X2=0 $Y2=0
cc_220 N_A_83_247#_M1009_g N_A_27_373#_c_884_n 8.91276e-19 $X=0.535 $Y=0.725
+ $X2=0 $Y2=0
cc_221 N_A_83_247#_c_179_n N_A_27_373#_c_885_n 0.00266509f $X=1.095 $Y=1.12
+ $X2=0 $Y2=0
cc_222 N_A_83_247#_c_199_p N_A_27_373#_c_886_n 0.0134182f $X=1.235 $Y=2.12 $X2=0
+ $Y2=0
cc_223 N_A_83_247#_c_185_n N_A_27_373#_c_886_n 0.0324215f $X=1.235 $Y=2.905
+ $X2=0 $Y2=0
cc_224 N_A_83_247#_c_186_n N_A_27_373#_c_895_n 0.065451f $X=3.345 $Y=2.99 $X2=0
+ $Y2=0
cc_225 N_A_83_247#_c_185_n N_A_27_373#_c_896_n 0.0138427f $X=1.235 $Y=2.905
+ $X2=0 $Y2=0
cc_226 N_A_83_247#_c_186_n N_A_27_373#_c_896_n 0.0124042f $X=3.345 $Y=2.99 $X2=0
+ $Y2=0
cc_227 N_A_83_247#_c_177_n N_A_27_373#_c_888_n 0.00205386f $X=0.62 $Y=1.36 $X2=0
+ $Y2=0
cc_228 N_A_83_247#_c_175_n N_A_27_373#_c_898_n 0.00748541f $X=0.505 $Y=1.79
+ $X2=0 $Y2=0
cc_229 N_A_83_247#_c_185_n N_A_27_373#_c_898_n 3.6586e-19 $X=1.235 $Y=2.905
+ $X2=0 $Y2=0
cc_230 N_A_83_247#_c_175_n N_A_27_373#_c_890_n 0.00595161f $X=0.505 $Y=1.79
+ $X2=0 $Y2=0
cc_231 N_A_83_247#_M1009_g N_A_27_373#_c_890_n 0.00484232f $X=0.535 $Y=0.725
+ $X2=0 $Y2=0
cc_232 N_A_83_247#_c_177_n N_A_27_373#_c_890_n 0.0125183f $X=0.62 $Y=1.36 $X2=0
+ $Y2=0
cc_233 N_A_83_247#_c_178_n N_A_27_373#_c_890_n 0.0133627f $X=0.58 $Y=1.4 $X2=0
+ $Y2=0
cc_234 N_A_83_247#_c_179_n N_A_27_373#_c_890_n 0.0234041f $X=1.095 $Y=1.12 $X2=0
+ $Y2=0
cc_235 N_A_83_247#_c_198_p N_A_27_373#_c_890_n 0.00662056f $X=1.095 $Y=2.035
+ $X2=0 $Y2=0
cc_236 N_A_83_247#_c_199_p N_A_27_373#_c_890_n 0.00256823f $X=1.235 $Y=2.12
+ $X2=0 $Y2=0
cc_237 N_A_83_247#_c_175_n N_A_27_373#_c_891_n 0.00130928f $X=0.505 $Y=1.79
+ $X2=0 $Y2=0
cc_238 N_A_83_247#_M1009_g N_A_27_373#_c_891_n 0.00113427f $X=0.535 $Y=0.725
+ $X2=0 $Y2=0
cc_239 N_A_83_247#_c_177_n N_A_27_373#_c_891_n 0.00131456f $X=0.62 $Y=1.36 $X2=0
+ $Y2=0
cc_240 N_A_83_247#_c_178_n N_A_27_373#_c_891_n 0.00136538f $X=0.58 $Y=1.4 $X2=0
+ $Y2=0
cc_241 N_A_83_247#_c_175_n N_A_27_373#_c_892_n 0.0237585f $X=0.505 $Y=1.79 $X2=0
+ $Y2=0
cc_242 N_A_83_247#_M1009_g N_A_27_373#_c_892_n 0.00350179f $X=0.535 $Y=0.725
+ $X2=0 $Y2=0
cc_243 N_A_83_247#_c_177_n N_A_27_373#_c_892_n 0.0180374f $X=0.62 $Y=1.36 $X2=0
+ $Y2=0
cc_244 N_A_83_247#_c_178_n N_A_27_373#_c_892_n 0.0438299f $X=0.58 $Y=1.4 $X2=0
+ $Y2=0
cc_245 N_A_83_247#_c_259_p N_A_27_373#_c_892_n 0.0136905f $X=0.745 $Y=2.035
+ $X2=0 $Y2=0
cc_246 N_A_83_247#_c_179_n N_A_27_373#_c_893_n 6.39812e-19 $X=1.095 $Y=1.12
+ $X2=0 $Y2=0
cc_247 N_A_83_247#_c_178_n N_VPWR_M1008_d 0.00106255f $X=0.58 $Y=1.4 $X2=-0.19
+ $Y2=-0.245
cc_248 N_A_83_247#_c_198_p N_VPWR_M1008_d 0.00542485f $X=1.095 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_249 N_A_83_247#_c_259_p N_VPWR_M1008_d 0.00153028f $X=0.745 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_250 N_A_83_247#_c_175_n N_VPWR_c_990_n 0.00609674f $X=0.505 $Y=1.79 $X2=0
+ $Y2=0
cc_251 N_A_83_247#_c_198_p N_VPWR_c_990_n 0.0127971f $X=1.095 $Y=2.035 $X2=0
+ $Y2=0
cc_252 N_A_83_247#_c_259_p N_VPWR_c_990_n 0.00833394f $X=0.745 $Y=2.035 $X2=0
+ $Y2=0
cc_253 N_A_83_247#_c_185_n N_VPWR_c_990_n 0.0235f $X=1.235 $Y=2.905 $X2=0 $Y2=0
cc_254 N_A_83_247#_c_187_n N_VPWR_c_990_n 0.0144537f $X=1.375 $Y=2.99 $X2=0
+ $Y2=0
cc_255 N_A_83_247#_c_186_n N_VPWR_c_995_n 0.1258f $X=3.345 $Y=2.99 $X2=0 $Y2=0
cc_256 N_A_83_247#_c_187_n N_VPWR_c_995_n 0.0200723f $X=1.375 $Y=2.99 $X2=0
+ $Y2=0
cc_257 N_A_83_247#_c_188_n N_VPWR_c_995_n 0.0213919f $X=3.51 $Y=2.795 $X2=0
+ $Y2=0
cc_258 N_A_83_247#_c_175_n N_VPWR_c_998_n 0.00497687f $X=0.505 $Y=1.79 $X2=0
+ $Y2=0
cc_259 N_A_83_247#_c_175_n N_VPWR_c_989_n 0.00515964f $X=0.505 $Y=1.79 $X2=0
+ $Y2=0
cc_260 N_A_83_247#_c_186_n N_VPWR_c_989_n 0.0663994f $X=3.345 $Y=2.99 $X2=0
+ $Y2=0
cc_261 N_A_83_247#_c_187_n N_VPWR_c_989_n 0.0108858f $X=1.375 $Y=2.99 $X2=0
+ $Y2=0
cc_262 N_A_83_247#_c_188_n N_VPWR_c_989_n 0.0110564f $X=3.51 $Y=2.795 $X2=0
+ $Y2=0
cc_263 N_A_83_247#_M1000_d N_A_332_373#_c_1079_n 0.00275472f $X=3.145 $Y=0.625
+ $X2=0 $Y2=0
cc_264 N_A_83_247#_c_182_n N_A_329_81#_M1018_d 0.00221108f $X=3.2 $Y=0.35
+ $X2=-0.19 $Y2=-0.245
cc_265 N_A_83_247#_M1000_d N_A_329_81#_c_1183_n 0.00880418f $X=3.145 $Y=0.625
+ $X2=0 $Y2=0
cc_266 N_A_83_247#_c_181_n N_A_329_81#_c_1183_n 0.022946f $X=3.365 $Y=0.36 $X2=0
+ $Y2=0
cc_267 N_A_83_247#_c_182_n N_A_329_81#_c_1183_n 0.0296435f $X=3.2 $Y=0.35 $X2=0
+ $Y2=0
cc_268 N_A_83_247#_M1012_d N_A_329_81#_c_1189_n 0.00744972f $X=3.28 $Y=1.865
+ $X2=0 $Y2=0
cc_269 N_A_83_247#_c_186_n N_A_329_81#_c_1189_n 0.0063494f $X=3.345 $Y=2.99
+ $X2=0 $Y2=0
cc_270 N_A_83_247#_c_188_n N_A_329_81#_c_1189_n 0.0247866f $X=3.51 $Y=2.795
+ $X2=0 $Y2=0
cc_271 N_A_83_247#_c_186_n N_A_329_81#_c_1190_n 0.0137218f $X=3.345 $Y=2.99
+ $X2=0 $Y2=0
cc_272 N_A_83_247#_c_193_p N_A_329_81#_c_1186_n 0.0207307f $X=1.26 $Y=0.55 $X2=0
+ $Y2=0
cc_273 N_A_83_247#_c_182_n N_A_329_81#_c_1186_n 0.0198438f $X=3.2 $Y=0.35 $X2=0
+ $Y2=0
cc_274 N_A_83_247#_c_182_n N_A_329_81#_c_1187_n 0.0530595f $X=3.2 $Y=0.35 $X2=0
+ $Y2=0
cc_275 N_A_83_247#_c_177_n N_VGND_M1009_d 8.63167e-19 $X=0.62 $Y=1.36 $X2=-0.19
+ $Y2=-0.245
cc_276 N_A_83_247#_c_179_n N_VGND_M1009_d 0.00177524f $X=1.095 $Y=1.12 $X2=-0.19
+ $Y2=-0.245
cc_277 N_A_83_247#_c_175_n N_VGND_c_1343_n 5.55578e-19 $X=0.505 $Y=1.79 $X2=0
+ $Y2=0
cc_278 N_A_83_247#_M1009_g N_VGND_c_1343_n 0.0146489f $X=0.535 $Y=0.725 $X2=0
+ $Y2=0
cc_279 N_A_83_247#_c_177_n N_VGND_c_1343_n 0.00852004f $X=0.62 $Y=1.36 $X2=0
+ $Y2=0
cc_280 N_A_83_247#_c_179_n N_VGND_c_1343_n 0.0127781f $X=1.095 $Y=1.12 $X2=0
+ $Y2=0
cc_281 N_A_83_247#_c_180_n N_VGND_c_1343_n 0.0129079f $X=1.345 $Y=0.34 $X2=0
+ $Y2=0
cc_282 N_A_83_247#_M1009_g N_VGND_c_1348_n 0.0045897f $X=0.535 $Y=0.725 $X2=0
+ $Y2=0
cc_283 N_A_83_247#_c_180_n N_VGND_c_1349_n 0.0179217f $X=1.345 $Y=0.34 $X2=0
+ $Y2=0
cc_284 N_A_83_247#_c_182_n N_VGND_c_1349_n 0.139665f $X=3.2 $Y=0.35 $X2=0 $Y2=0
cc_285 N_A_83_247#_M1000_d N_VGND_c_1354_n 0.00251887f $X=3.145 $Y=0.625 $X2=0
+ $Y2=0
cc_286 N_A_83_247#_M1009_g N_VGND_c_1354_n 0.0044912f $X=0.535 $Y=0.725 $X2=0
+ $Y2=0
cc_287 N_A_83_247#_c_180_n N_VGND_c_1354_n 0.00971942f $X=1.345 $Y=0.34 $X2=0
+ $Y2=0
cc_288 N_A_83_247#_c_182_n N_VGND_c_1354_n 0.0773214f $X=3.2 $Y=0.35 $X2=0 $Y2=0
cc_289 N_A_M1007_g N_B_M1018_g 0.0218506f $X=1.045 $Y=0.725 $X2=0 $Y2=0
cc_290 N_A_c_304_n N_B_M1018_g 0.0196651f $X=1.045 $Y=1.79 $X2=0 $Y2=0
cc_291 N_A_c_305_n N_B_M1018_g 0.00253548f $X=1.12 $Y=1.54 $X2=0 $Y2=0
cc_292 N_A_c_304_n N_B_c_473_n 0.00482393f $X=1.045 $Y=1.79 $X2=0 $Y2=0
cc_293 N_A_c_304_n N_B_c_467_n 0.00253898f $X=1.045 $Y=1.79 $X2=0 $Y2=0
cc_294 N_A_c_304_n N_B_M1005_g 0.0168148f $X=1.045 $Y=1.79 $X2=0 $Y2=0
cc_295 N_A_M1007_g N_A_27_373#_c_885_n 0.00146258f $X=1.045 $Y=0.725 $X2=0 $Y2=0
cc_296 N_A_c_305_n N_A_27_373#_c_885_n 2.43113e-19 $X=1.12 $Y=1.54 $X2=0 $Y2=0
cc_297 N_A_c_304_n N_A_27_373#_c_886_n 0.00158086f $X=1.045 $Y=1.79 $X2=0 $Y2=0
cc_298 N_A_c_305_n N_A_27_373#_c_886_n 0.0238695f $X=1.12 $Y=1.54 $X2=0 $Y2=0
cc_299 N_A_M1007_g N_A_27_373#_c_890_n 0.00523989f $X=1.045 $Y=0.725 $X2=0 $Y2=0
cc_300 N_A_c_305_n N_A_27_373#_c_890_n 0.0103716f $X=1.12 $Y=1.54 $X2=0 $Y2=0
cc_301 N_A_c_305_n N_A_27_373#_c_893_n 8.6259e-19 $X=1.12 $Y=1.54 $X2=0 $Y2=0
cc_302 N_A_c_304_n N_VPWR_c_990_n 0.00434996f $X=1.045 $Y=1.79 $X2=0 $Y2=0
cc_303 N_A_c_304_n N_VPWR_c_995_n 0.00438247f $X=1.045 $Y=1.79 $X2=0 $Y2=0
cc_304 N_A_c_304_n N_VPWR_c_989_n 0.0042997f $X=1.045 $Y=1.79 $X2=0 $Y2=0
cc_305 N_A_M1007_g N_VGND_c_1343_n 0.00352423f $X=1.045 $Y=0.725 $X2=0 $Y2=0
cc_306 N_A_M1007_g N_VGND_c_1349_n 0.0047553f $X=1.045 $Y=0.725 $X2=0 $Y2=0
cc_307 N_A_M1007_g N_VGND_c_1354_n 0.00445555f $X=1.045 $Y=0.725 $X2=0 $Y2=0
cc_308 N_A_397_21#_M1002_g N_B_M1018_g 0.0348758f $X=2.06 $Y=1.055 $X2=0 $Y2=0
cc_309 N_A_397_21#_c_347_n N_B_M1018_g 2.98053e-19 $X=2.195 $Y=1.7 $X2=0 $Y2=0
cc_310 N_A_397_21#_c_347_n N_B_c_467_n 0.00678918f $X=2.195 $Y=1.7 $X2=0 $Y2=0
cc_311 N_A_397_21#_c_357_n N_B_M1005_g 0.0135936f $X=2.195 $Y=1.79 $X2=0 $Y2=0
cc_312 N_A_397_21#_c_357_n N_B_c_477_n 0.00313361f $X=2.195 $Y=1.79 $X2=0 $Y2=0
cc_313 N_A_397_21#_c_347_n N_B_c_468_n 0.0161249f $X=2.195 $Y=1.7 $X2=0 $Y2=0
cc_314 N_A_397_21#_c_351_n N_B_c_468_n 0.0140229f $X=3.205 $Y=1.79 $X2=0 $Y2=0
cc_315 N_A_397_21#_c_354_n N_B_c_468_n 2.81659e-19 $X=3.32 $Y=1.54 $X2=0 $Y2=0
cc_316 N_A_397_21#_M1002_g N_B_M1001_g 0.022321f $X=2.06 $Y=1.055 $X2=0 $Y2=0
cc_317 N_A_397_21#_c_346_n N_B_M1001_g 0.0101362f $X=2.195 $Y=1.49 $X2=0 $Y2=0
cc_318 N_A_397_21#_c_348_n N_B_M1001_g 0.00737859f $X=2.995 $Y=0.18 $X2=0 $Y2=0
cc_319 N_A_397_21#_M1000_g N_B_M1001_g 0.0245034f $X=3.07 $Y=0.945 $X2=0 $Y2=0
cc_320 N_A_397_21#_c_357_n N_B_c_480_n 0.00222081f $X=2.195 $Y=1.79 $X2=0 $Y2=0
cc_321 N_A_397_21#_c_351_n N_B_c_480_n 0.00736303f $X=3.205 $Y=1.79 $X2=0 $Y2=0
cc_322 N_A_397_21#_c_357_n N_B_M1003_g 0.00551715f $X=2.195 $Y=1.79 $X2=0 $Y2=0
cc_323 N_A_397_21#_c_351_n N_B_M1003_g 0.0105677f $X=3.205 $Y=1.79 $X2=0 $Y2=0
cc_324 N_A_397_21#_c_351_n N_B_c_483_n 0.00737859f $X=3.205 $Y=1.79 $X2=0 $Y2=0
cc_325 N_A_397_21#_c_351_n N_B_c_484_n 0.0259158f $X=3.205 $Y=1.79 $X2=0 $Y2=0
cc_326 N_A_397_21#_c_360_n N_B_c_484_n 0.0149371f $X=4.09 $Y=2.115 $X2=0 $Y2=0
cc_327 N_A_397_21#_c_354_n N_B_c_484_n 0.00342023f $X=3.32 $Y=1.54 $X2=0 $Y2=0
cc_328 N_A_397_21#_c_353_n N_B_M1014_g 0.00383817f $X=3.925 $Y=1.04 $X2=0 $Y2=0
cc_329 N_A_397_21#_c_355_n N_B_M1014_g 0.00357912f $X=3.36 $Y=1.375 $X2=0 $Y2=0
cc_330 N_A_397_21#_c_360_n N_B_c_485_n 0.00388282f $X=4.09 $Y=2.115 $X2=0 $Y2=0
cc_331 N_A_397_21#_M1000_g N_B_c_471_n 4.40661e-19 $X=3.07 $Y=0.945 $X2=0 $Y2=0
cc_332 N_A_397_21#_c_351_n N_B_c_471_n 0.0181869f $X=3.205 $Y=1.79 $X2=0 $Y2=0
cc_333 N_A_397_21#_c_353_n N_B_c_471_n 0.00237277f $X=3.925 $Y=1.04 $X2=0 $Y2=0
cc_334 N_A_397_21#_c_360_n N_B_c_471_n 0.00187046f $X=4.09 $Y=2.115 $X2=0 $Y2=0
cc_335 N_A_397_21#_c_355_n N_B_c_471_n 0.00342023f $X=3.36 $Y=1.375 $X2=0 $Y2=0
cc_336 N_A_397_21#_c_351_n N_B_c_472_n 3.47661e-19 $X=3.205 $Y=1.79 $X2=0 $Y2=0
cc_337 N_A_397_21#_c_353_n N_B_c_472_n 0.0145936f $X=3.925 $Y=1.04 $X2=0 $Y2=0
cc_338 N_A_397_21#_c_360_n N_B_c_472_n 0.0385923f $X=4.09 $Y=2.115 $X2=0 $Y2=0
cc_339 N_A_397_21#_c_355_n N_B_c_472_n 0.0356463f $X=3.36 $Y=1.375 $X2=0 $Y2=0
cc_340 N_A_397_21#_c_346_n N_A_27_373#_c_886_n 0.00200088f $X=2.195 $Y=1.49
+ $X2=0 $Y2=0
cc_341 N_A_397_21#_c_347_n N_A_27_373#_c_886_n 0.00138386f $X=2.195 $Y=1.7 $X2=0
+ $Y2=0
cc_342 N_A_397_21#_c_357_n N_A_27_373#_c_886_n 6.75198e-19 $X=2.195 $Y=1.79
+ $X2=0 $Y2=0
cc_343 N_A_397_21#_M1002_g N_A_27_373#_c_887_n 0.00808752f $X=2.06 $Y=1.055
+ $X2=0 $Y2=0
cc_344 N_A_397_21#_c_346_n N_A_27_373#_c_887_n 0.00253261f $X=2.195 $Y=1.49
+ $X2=0 $Y2=0
cc_345 N_A_397_21#_c_357_n N_A_27_373#_c_895_n 0.0110237f $X=2.195 $Y=1.79 $X2=0
+ $Y2=0
cc_346 N_A_397_21#_c_351_n N_A_27_373#_c_895_n 4.54131e-19 $X=3.205 $Y=1.79
+ $X2=0 $Y2=0
cc_347 N_A_397_21#_c_357_n N_A_27_373#_c_897_n 8.89727e-19 $X=2.195 $Y=1.79
+ $X2=0 $Y2=0
cc_348 N_A_397_21#_M1002_g N_A_27_373#_c_889_n 0.00115834f $X=2.06 $Y=1.055
+ $X2=0 $Y2=0
cc_349 N_A_397_21#_c_346_n N_A_27_373#_c_889_n 0.00618395f $X=2.195 $Y=1.49
+ $X2=0 $Y2=0
cc_350 N_A_397_21#_c_346_n N_A_27_373#_c_893_n 5.07152e-19 $X=2.195 $Y=1.49
+ $X2=0 $Y2=0
cc_351 N_A_397_21#_c_357_n N_A_332_373#_c_1083_n 0.00512528f $X=2.195 $Y=1.79
+ $X2=0 $Y2=0
cc_352 N_A_397_21#_c_347_n N_A_332_373#_c_1072_n 0.00638935f $X=2.195 $Y=1.7
+ $X2=0 $Y2=0
cc_353 N_A_397_21#_c_357_n N_A_332_373#_c_1072_n 0.00799422f $X=2.195 $Y=1.79
+ $X2=0 $Y2=0
cc_354 N_A_397_21#_c_351_n N_A_332_373#_c_1072_n 7.31148e-19 $X=3.205 $Y=1.79
+ $X2=0 $Y2=0
cc_355 N_A_397_21#_c_359_n N_A_332_373#_c_1072_n 4.14392e-19 $X=3.48 $Y=1.95
+ $X2=0 $Y2=0
cc_356 N_A_397_21#_c_354_n N_A_332_373#_c_1072_n 0.00629057f $X=3.32 $Y=1.54
+ $X2=0 $Y2=0
cc_357 N_A_397_21#_c_346_n N_A_332_373#_c_1073_n 0.00373139f $X=2.195 $Y=1.49
+ $X2=0 $Y2=0
cc_358 N_A_397_21#_c_347_n N_A_332_373#_c_1073_n 0.00177444f $X=2.195 $Y=1.7
+ $X2=0 $Y2=0
cc_359 N_A_397_21#_c_357_n N_A_332_373#_c_1073_n 2.27799e-19 $X=2.195 $Y=1.79
+ $X2=0 $Y2=0
cc_360 N_A_397_21#_M1000_g N_A_332_373#_c_1078_n 3.44089e-19 $X=3.07 $Y=0.945
+ $X2=0 $Y2=0
cc_361 N_A_397_21#_c_355_n N_A_332_373#_c_1078_n 0.00301081f $X=3.36 $Y=1.375
+ $X2=0 $Y2=0
cc_362 N_A_397_21#_M1000_g N_A_332_373#_c_1079_n 0.00695074f $X=3.07 $Y=0.945
+ $X2=0 $Y2=0
cc_363 N_A_397_21#_c_351_n N_A_332_373#_c_1079_n 3.48429e-19 $X=3.205 $Y=1.79
+ $X2=0 $Y2=0
cc_364 N_A_397_21#_c_353_n N_A_332_373#_c_1079_n 0.018201f $X=3.925 $Y=1.04
+ $X2=0 $Y2=0
cc_365 N_A_397_21#_c_360_n N_A_332_373#_c_1079_n 0.00714987f $X=4.09 $Y=2.115
+ $X2=0 $Y2=0
cc_366 N_A_397_21#_c_354_n N_A_332_373#_c_1079_n 0.00904642f $X=3.32 $Y=1.54
+ $X2=0 $Y2=0
cc_367 N_A_397_21#_c_355_n N_A_332_373#_c_1079_n 0.0193866f $X=3.36 $Y=1.375
+ $X2=0 $Y2=0
cc_368 N_A_397_21#_M1000_g N_A_332_373#_c_1080_n 7.21505e-19 $X=3.07 $Y=0.945
+ $X2=0 $Y2=0
cc_369 N_A_397_21#_c_354_n N_A_332_373#_c_1080_n 8.91892e-19 $X=3.32 $Y=1.54
+ $X2=0 $Y2=0
cc_370 N_A_397_21#_c_355_n N_A_332_373#_c_1080_n 4.32441e-19 $X=3.36 $Y=1.375
+ $X2=0 $Y2=0
cc_371 N_A_397_21#_c_346_n N_A_332_373#_c_1081_n 0.00119995f $X=2.195 $Y=1.49
+ $X2=0 $Y2=0
cc_372 N_A_397_21#_M1000_g N_A_332_373#_c_1081_n 0.00178826f $X=3.07 $Y=0.945
+ $X2=0 $Y2=0
cc_373 N_A_397_21#_c_354_n N_A_332_373#_c_1081_n 0.00645185f $X=3.32 $Y=1.54
+ $X2=0 $Y2=0
cc_374 N_A_397_21#_c_355_n N_A_332_373#_c_1081_n 0.00139636f $X=3.36 $Y=1.375
+ $X2=0 $Y2=0
cc_375 N_A_397_21#_M1014_s N_A_329_81#_c_1183_n 0.00698754f $X=3.78 $Y=0.445
+ $X2=0 $Y2=0
cc_376 N_A_397_21#_M1000_g N_A_329_81#_c_1183_n 0.0140287f $X=3.07 $Y=0.945
+ $X2=0 $Y2=0
cc_377 N_A_397_21#_c_351_n N_A_329_81#_c_1183_n 0.00133872f $X=3.205 $Y=1.79
+ $X2=0 $Y2=0
cc_378 N_A_397_21#_c_352_n N_A_329_81#_c_1183_n 0.01346f $X=3.565 $Y=1.04 $X2=0
+ $Y2=0
cc_379 N_A_397_21#_c_353_n N_A_329_81#_c_1183_n 0.0328652f $X=3.925 $Y=1.04
+ $X2=0 $Y2=0
cc_380 N_A_397_21#_c_354_n N_A_329_81#_c_1183_n 0.00253746f $X=3.32 $Y=1.54
+ $X2=0 $Y2=0
cc_381 N_A_397_21#_c_351_n N_A_329_81#_c_1211_n 0.0125403f $X=3.205 $Y=1.79
+ $X2=0 $Y2=0
cc_382 N_A_397_21#_c_359_n N_A_329_81#_c_1211_n 0.0040702f $X=3.48 $Y=1.95 $X2=0
+ $Y2=0
cc_383 N_A_397_21#_c_371_n N_A_329_81#_c_1211_n 0.0152791f $X=3.565 $Y=2.075
+ $X2=0 $Y2=0
cc_384 N_A_397_21#_M1020_s N_A_329_81#_c_1189_n 0.00684634f $X=3.95 $Y=1.84
+ $X2=0 $Y2=0
cc_385 N_A_397_21#_c_351_n N_A_329_81#_c_1189_n 0.0115837f $X=3.205 $Y=1.79
+ $X2=0 $Y2=0
cc_386 N_A_397_21#_c_371_n N_A_329_81#_c_1189_n 0.0137412f $X=3.565 $Y=2.075
+ $X2=0 $Y2=0
cc_387 N_A_397_21#_c_360_n N_A_329_81#_c_1189_n 0.0468706f $X=4.09 $Y=2.115
+ $X2=0 $Y2=0
cc_388 N_A_397_21#_c_354_n N_A_329_81#_c_1189_n 0.0049788f $X=3.32 $Y=1.54 $X2=0
+ $Y2=0
cc_389 N_A_397_21#_c_351_n N_A_329_81#_c_1190_n 4.28378e-19 $X=3.205 $Y=1.79
+ $X2=0 $Y2=0
cc_390 N_A_397_21#_c_353_n N_A_329_81#_c_1184_n 3.53781e-19 $X=3.925 $Y=1.04
+ $X2=0 $Y2=0
cc_391 N_A_397_21#_c_353_n N_A_329_81#_c_1185_n 0.00564206f $X=3.925 $Y=1.04
+ $X2=0 $Y2=0
cc_392 N_A_397_21#_c_360_n N_A_329_81#_c_1185_n 0.0116682f $X=4.09 $Y=2.115
+ $X2=0 $Y2=0
cc_393 N_A_397_21#_M1002_g N_A_329_81#_c_1186_n 0.0033689f $X=2.06 $Y=1.055
+ $X2=0 $Y2=0
cc_394 N_A_397_21#_M1002_g N_A_329_81#_c_1187_n 0.0109418f $X=2.06 $Y=1.055
+ $X2=0 $Y2=0
cc_395 N_A_397_21#_c_346_n N_A_329_81#_c_1187_n 4.49394e-19 $X=2.195 $Y=1.49
+ $X2=0 $Y2=0
cc_396 N_A_397_21#_M1000_g N_A_329_81#_c_1188_n 4.77048e-19 $X=3.07 $Y=0.945
+ $X2=0 $Y2=0
cc_397 N_A_397_21#_c_349_n N_VGND_c_1349_n 0.0250991f $X=2.135 $Y=0.18 $X2=0
+ $Y2=0
cc_398 N_A_397_21#_c_348_n N_VGND_c_1354_n 0.0262914f $X=2.995 $Y=0.18 $X2=0
+ $Y2=0
cc_399 N_A_397_21#_c_349_n N_VGND_c_1354_n 0.00604517f $X=2.135 $Y=0.18 $X2=0
+ $Y2=0
cc_400 N_B_M1018_g N_A_27_373#_c_885_n 0.0126155f $X=1.57 $Y=0.725 $X2=0 $Y2=0
cc_401 N_B_M1018_g N_A_27_373#_c_886_n 0.00273704f $X=1.57 $Y=0.725 $X2=0 $Y2=0
cc_402 N_B_c_467_n N_A_27_373#_c_886_n 0.00863201f $X=1.585 $Y=1.79 $X2=0 $Y2=0
cc_403 N_B_M1005_g N_A_27_373#_c_886_n 0.0204145f $X=1.585 $Y=2.285 $X2=0 $Y2=0
cc_404 N_B_c_480_n N_A_27_373#_c_895_n 0.00353132f $X=2.665 $Y=2.67 $X2=0 $Y2=0
cc_405 N_B_c_481_n N_A_27_373#_c_895_n 0.00341288f $X=2.665 $Y=3.075 $X2=0 $Y2=0
cc_406 N_B_M1003_g N_A_27_373#_c_895_n 3.18186e-19 $X=2.665 $Y=2.185 $X2=0 $Y2=0
cc_407 N_B_c_473_n N_A_27_373#_c_896_n 4.31853e-19 $X=1.585 $Y=2.87 $X2=0 $Y2=0
cc_408 N_B_M1005_g N_A_27_373#_c_896_n 0.00798502f $X=1.585 $Y=2.285 $X2=0 $Y2=0
cc_409 N_B_c_468_n N_A_27_373#_c_897_n 4.34797e-19 $X=2.57 $Y=1.505 $X2=0 $Y2=0
cc_410 N_B_M1003_g N_A_27_373#_c_897_n 0.00828225f $X=2.665 $Y=2.185 $X2=0 $Y2=0
cc_411 N_B_M1001_g N_A_27_373#_c_889_n 0.00345094f $X=2.57 $Y=0.945 $X2=0 $Y2=0
cc_412 N_B_M1018_g N_A_27_373#_c_890_n 0.00425614f $X=1.57 $Y=0.725 $X2=0 $Y2=0
cc_413 N_B_M1018_g N_A_27_373#_c_893_n 0.00193489f $X=1.57 $Y=0.725 $X2=0 $Y2=0
cc_414 N_B_c_474_n N_VPWR_c_990_n 2.90675e-19 $X=1.585 $Y=3.075 $X2=0 $Y2=0
cc_415 N_B_c_478_n N_VPWR_c_990_n 0.00242213f $X=1.675 $Y=3.15 $X2=0 $Y2=0
cc_416 N_B_c_484_n N_VPWR_c_991_n 0.0027703f $X=3.8 $Y=3.075 $X2=0 $Y2=0
cc_417 N_B_c_485_n N_VPWR_c_991_n 0.0147276f $X=4.315 $Y=1.765 $X2=0 $Y2=0
cc_418 N_B_c_478_n N_VPWR_c_995_n 0.0540846f $X=1.675 $Y=3.15 $X2=0 $Y2=0
cc_419 N_B_c_485_n N_VPWR_c_995_n 0.00461464f $X=4.315 $Y=1.765 $X2=0 $Y2=0
cc_420 N_B_c_477_n N_VPWR_c_989_n 0.0211783f $X=2.575 $Y=3.15 $X2=0 $Y2=0
cc_421 N_B_c_478_n N_VPWR_c_989_n 0.00675277f $X=1.675 $Y=3.15 $X2=0 $Y2=0
cc_422 N_B_c_483_n N_VPWR_c_989_n 0.0301174f $X=3.725 $Y=3.15 $X2=0 $Y2=0
cc_423 N_B_c_485_n N_VPWR_c_989_n 0.00457124f $X=4.315 $Y=1.765 $X2=0 $Y2=0
cc_424 N_B_c_486_n N_VPWR_c_989_n 0.00442127f $X=2.665 $Y=3.15 $X2=0 $Y2=0
cc_425 N_B_c_467_n N_A_332_373#_c_1083_n 2.33109e-19 $X=1.585 $Y=1.79 $X2=0
+ $Y2=0
cc_426 N_B_M1005_g N_A_332_373#_c_1083_n 0.00199937f $X=1.585 $Y=2.285 $X2=0
+ $Y2=0
cc_427 N_B_c_468_n N_A_332_373#_c_1072_n 0.0158183f $X=2.57 $Y=1.505 $X2=0 $Y2=0
cc_428 N_B_c_467_n N_A_332_373#_c_1073_n 6.85032e-19 $X=1.585 $Y=1.79 $X2=0
+ $Y2=0
cc_429 N_B_c_468_n N_A_332_373#_c_1078_n 4.47675e-19 $X=2.57 $Y=1.505 $X2=0
+ $Y2=0
cc_430 N_B_M1001_g N_A_332_373#_c_1078_n 0.00588367f $X=2.57 $Y=0.945 $X2=0
+ $Y2=0
cc_431 N_B_M1014_g N_A_332_373#_c_1079_n 0.00592452f $X=4.14 $Y=0.815 $X2=0
+ $Y2=0
cc_432 N_B_c_471_n N_A_332_373#_c_1079_n 0.00595754f $X=4.24 $Y=1.515 $X2=0
+ $Y2=0
cc_433 N_B_c_472_n N_A_332_373#_c_1079_n 0.0255335f $X=4.24 $Y=1.515 $X2=0 $Y2=0
cc_434 N_B_M1001_g N_A_332_373#_c_1080_n 0.00173286f $X=2.57 $Y=0.945 $X2=0
+ $Y2=0
cc_435 N_B_c_468_n N_A_332_373#_c_1081_n 0.00384975f $X=2.57 $Y=1.505 $X2=0
+ $Y2=0
cc_436 N_B_M1001_g N_A_332_373#_c_1081_n 0.005578f $X=2.57 $Y=0.945 $X2=0 $Y2=0
cc_437 N_B_M1014_g N_A_329_81#_c_1183_n 0.0169621f $X=4.14 $Y=0.815 $X2=0 $Y2=0
cc_438 N_B_c_471_n N_A_329_81#_c_1183_n 7.96102e-19 $X=4.24 $Y=1.515 $X2=0 $Y2=0
cc_439 N_B_c_472_n N_A_329_81#_c_1183_n 0.00378334f $X=4.24 $Y=1.515 $X2=0 $Y2=0
cc_440 N_B_M1003_g N_A_329_81#_c_1211_n 0.00473045f $X=2.665 $Y=2.185 $X2=0
+ $Y2=0
cc_441 N_B_c_484_n N_A_329_81#_c_1211_n 9.53238e-19 $X=3.8 $Y=3.075 $X2=0 $Y2=0
cc_442 N_B_c_483_n N_A_329_81#_c_1189_n 9.96978e-19 $X=3.725 $Y=3.15 $X2=0 $Y2=0
cc_443 N_B_c_484_n N_A_329_81#_c_1189_n 0.013112f $X=3.8 $Y=3.075 $X2=0 $Y2=0
cc_444 N_B_c_485_n N_A_329_81#_c_1189_n 0.0159691f $X=4.315 $Y=1.765 $X2=0 $Y2=0
cc_445 N_B_c_472_n N_A_329_81#_c_1189_n 0.00378789f $X=4.24 $Y=1.515 $X2=0 $Y2=0
cc_446 N_B_c_480_n N_A_329_81#_c_1190_n 3.6329e-19 $X=2.665 $Y=2.67 $X2=0 $Y2=0
cc_447 N_B_M1003_g N_A_329_81#_c_1190_n 0.00202095f $X=2.665 $Y=2.185 $X2=0
+ $Y2=0
cc_448 N_B_M1014_g N_A_329_81#_c_1184_n 0.00981436f $X=4.14 $Y=0.815 $X2=0 $Y2=0
cc_449 N_B_M1014_g N_A_329_81#_c_1185_n 0.00795796f $X=4.14 $Y=0.815 $X2=0 $Y2=0
cc_450 N_B_c_485_n N_A_329_81#_c_1185_n 0.0164961f $X=4.315 $Y=1.765 $X2=0 $Y2=0
cc_451 N_B_c_471_n N_A_329_81#_c_1185_n 0.0100866f $X=4.24 $Y=1.515 $X2=0 $Y2=0
cc_452 N_B_c_472_n N_A_329_81#_c_1185_n 0.0324535f $X=4.24 $Y=1.515 $X2=0 $Y2=0
cc_453 N_B_M1018_g N_A_329_81#_c_1186_n 0.00561682f $X=1.57 $Y=0.725 $X2=0 $Y2=0
cc_454 N_B_M1001_g N_A_329_81#_c_1187_n 0.00493879f $X=2.57 $Y=0.945 $X2=0 $Y2=0
cc_455 N_B_M1001_g N_A_329_81#_c_1188_n 0.00621366f $X=2.57 $Y=0.945 $X2=0 $Y2=0
cc_456 N_B_c_485_n N_A_329_81#_c_1246_n 0.00100036f $X=4.315 $Y=1.765 $X2=0
+ $Y2=0
cc_457 N_B_M1014_g N_VGND_c_1344_n 0.00546687f $X=4.14 $Y=0.815 $X2=0 $Y2=0
cc_458 N_B_M1018_g N_VGND_c_1349_n 9.15902e-19 $X=1.57 $Y=0.725 $X2=0 $Y2=0
cc_459 N_B_M1014_g N_VGND_c_1349_n 0.00399972f $X=4.14 $Y=0.815 $X2=0 $Y2=0
cc_460 N_B_M1014_g N_VGND_c_1354_n 0.0052212f $X=4.14 $Y=0.815 $X2=0 $Y2=0
cc_461 N_A_1027_48#_M1023_g N_C_c_679_n 0.0203498f $X=5.21 $Y=0.69 $X2=-0.19
+ $Y2=-0.245
cc_462 N_A_1027_48#_c_604_n N_C_c_681_n 0.0010582f $X=5.395 $Y=1.92 $X2=0 $Y2=0
cc_463 N_A_1027_48#_c_605_n N_C_c_681_n 0.00175105f $X=6.39 $Y=1.64 $X2=0 $Y2=0
cc_464 N_A_1027_48#_M1023_g N_C_c_682_n 0.00501499f $X=5.21 $Y=0.69 $X2=0 $Y2=0
cc_465 N_A_1027_48#_c_604_n N_C_c_682_n 0.0158957f $X=5.395 $Y=1.92 $X2=0 $Y2=0
cc_466 N_A_1027_48#_c_605_n N_C_c_682_n 0.00706975f $X=6.39 $Y=1.64 $X2=0 $Y2=0
cc_467 N_A_1027_48#_c_606_n N_C_c_682_n 0.00100186f $X=6.532 $Y=1.475 $X2=0
+ $Y2=0
cc_468 N_A_1027_48#_c_607_n N_C_c_682_n 8.39659e-19 $X=6.555 $Y=1.085 $X2=0
+ $Y2=0
cc_469 N_A_1027_48#_c_604_n N_C_c_683_n 0.00400946f $X=5.395 $Y=1.92 $X2=0 $Y2=0
cc_470 N_A_1027_48#_c_605_n N_C_c_683_n 0.0148889f $X=6.39 $Y=1.64 $X2=0 $Y2=0
cc_471 N_A_1027_48#_c_613_n N_C_c_683_n 0.00310748f $X=6.687 $Y=1.95 $X2=0 $Y2=0
cc_472 N_A_1027_48#_c_604_n N_C_c_689_n 0.0241798f $X=5.395 $Y=1.92 $X2=0 $Y2=0
cc_473 N_A_1027_48#_c_611_n N_C_c_689_n 0.00108764f $X=6.687 $Y=2.132 $X2=0
+ $Y2=0
cc_474 N_A_1027_48#_c_613_n N_C_c_689_n 0.00148353f $X=6.687 $Y=1.95 $X2=0 $Y2=0
cc_475 N_A_1027_48#_c_605_n N_C_c_684_n 0.0156516f $X=6.39 $Y=1.64 $X2=0 $Y2=0
cc_476 N_A_1027_48#_c_606_n N_C_c_684_n 0.0149313f $X=6.532 $Y=1.475 $X2=0 $Y2=0
cc_477 N_A_1027_48#_c_611_n N_C_c_684_n 6.80956e-19 $X=6.687 $Y=2.132 $X2=0
+ $Y2=0
cc_478 N_A_1027_48#_c_608_n N_C_c_684_n 0.00752536f $X=6.532 $Y=1.64 $X2=0 $Y2=0
cc_479 N_A_1027_48#_c_606_n N_C_c_685_n 0.00373839f $X=6.532 $Y=1.475 $X2=0
+ $Y2=0
cc_480 N_A_1027_48#_c_607_n N_C_c_685_n 0.00308441f $X=6.555 $Y=1.085 $X2=0
+ $Y2=0
cc_481 N_A_1027_48#_c_611_n N_C_c_686_n 0.0113116f $X=6.687 $Y=2.132 $X2=0 $Y2=0
cc_482 N_A_1027_48#_c_608_n N_C_c_686_n 0.00431019f $X=6.532 $Y=1.64 $X2=0 $Y2=0
cc_483 N_A_1027_48#_c_613_n N_C_c_686_n 0.00447616f $X=6.687 $Y=1.95 $X2=0 $Y2=0
cc_484 N_A_1027_48#_c_606_n N_C_c_687_n 0.00923975f $X=6.532 $Y=1.475 $X2=0
+ $Y2=0
cc_485 N_A_1027_48#_c_611_n N_C_c_687_n 0.0020105f $X=6.687 $Y=2.132 $X2=0 $Y2=0
cc_486 N_A_1027_48#_c_608_n N_C_c_687_n 0.0260181f $X=6.532 $Y=1.64 $X2=0 $Y2=0
cc_487 N_A_1027_48#_M1023_g N_A_1057_74#_c_765_n 0.00359689f $X=5.21 $Y=0.69
+ $X2=0 $Y2=0
cc_488 N_A_1027_48#_c_611_n N_A_1057_74#_c_774_n 0.0140322f $X=6.687 $Y=2.132
+ $X2=0 $Y2=0
cc_489 N_A_1027_48#_M1010_s N_A_1057_74#_c_767_n 0.0013543f $X=6.41 $Y=0.81
+ $X2=0 $Y2=0
cc_490 N_A_1027_48#_c_607_n N_A_1057_74#_c_767_n 0.0127928f $X=6.555 $Y=1.085
+ $X2=0 $Y2=0
cc_491 N_A_1027_48#_M1010_s N_A_1057_74#_c_768_n 9.85725e-19 $X=6.41 $Y=0.81
+ $X2=0 $Y2=0
cc_492 N_A_1027_48#_c_605_n N_A_1057_74#_c_768_n 0.00180192f $X=6.39 $Y=1.64
+ $X2=0 $Y2=0
cc_493 N_A_1027_48#_c_607_n N_A_1057_74#_c_768_n 0.00977295f $X=6.555 $Y=1.085
+ $X2=0 $Y2=0
cc_494 N_A_1027_48#_c_611_n N_A_1057_74#_c_775_n 0.0283041f $X=6.687 $Y=2.132
+ $X2=0 $Y2=0
cc_495 N_A_1027_48#_c_611_n N_A_1057_74#_c_788_n 0.0138654f $X=6.687 $Y=2.132
+ $X2=0 $Y2=0
cc_496 N_A_1027_48#_c_604_n N_A_1057_74#_c_777_n 0.00666738f $X=5.395 $Y=1.92
+ $X2=0 $Y2=0
cc_497 N_A_1027_48#_c_604_n N_VPWR_c_991_n 0.0058266f $X=5.395 $Y=1.92 $X2=0
+ $Y2=0
cc_498 N_A_1027_48#_c_604_n N_VPWR_c_996_n 0.00490845f $X=5.395 $Y=1.92 $X2=0
+ $Y2=0
cc_499 N_A_1027_48#_c_604_n N_VPWR_c_989_n 0.00506877f $X=5.395 $Y=1.92 $X2=0
+ $Y2=0
cc_500 N_A_1027_48#_M1023_g N_A_332_373#_c_1074_n 0.00376703f $X=5.21 $Y=0.69
+ $X2=0 $Y2=0
cc_501 N_A_1027_48#_M1023_g N_A_332_373#_c_1075_n 0.00796217f $X=5.21 $Y=0.69
+ $X2=0 $Y2=0
cc_502 N_A_1027_48#_c_604_n N_A_332_373#_c_1075_n 0.0177876f $X=5.395 $Y=1.92
+ $X2=0 $Y2=0
cc_503 N_A_1027_48#_c_605_n N_A_332_373#_c_1075_n 0.0255168f $X=6.39 $Y=1.64
+ $X2=0 $Y2=0
cc_504 N_A_1027_48#_M1023_g N_A_332_373#_c_1076_n 0.0134853f $X=5.21 $Y=0.69
+ $X2=0 $Y2=0
cc_505 N_A_1027_48#_c_604_n N_A_332_373#_c_1076_n 0.00879145f $X=5.395 $Y=1.92
+ $X2=0 $Y2=0
cc_506 N_A_1027_48#_c_605_n N_A_332_373#_c_1076_n 0.0663436f $X=6.39 $Y=1.64
+ $X2=0 $Y2=0
cc_507 N_A_1027_48#_c_607_n N_A_332_373#_c_1076_n 0.0120264f $X=6.555 $Y=1.085
+ $X2=0 $Y2=0
cc_508 N_A_1027_48#_M1023_g N_A_332_373#_c_1077_n 2.07613e-19 $X=5.21 $Y=0.69
+ $X2=0 $Y2=0
cc_509 N_A_1027_48#_c_607_n N_A_332_373#_c_1077_n 0.00906723f $X=6.555 $Y=1.085
+ $X2=0 $Y2=0
cc_510 N_A_1027_48#_c_604_n N_A_332_373#_c_1087_n 0.0113899f $X=5.395 $Y=1.92
+ $X2=0 $Y2=0
cc_511 N_A_1027_48#_c_605_n N_A_332_373#_c_1087_n 7.34818e-19 $X=6.39 $Y=1.64
+ $X2=0 $Y2=0
cc_512 N_A_1027_48#_M1023_g N_A_332_373#_c_1082_n 0.00454209f $X=5.21 $Y=0.69
+ $X2=0 $Y2=0
cc_513 N_A_1027_48#_M1023_g N_A_329_81#_c_1184_n 0.00727684f $X=5.21 $Y=0.69
+ $X2=0 $Y2=0
cc_514 N_A_1027_48#_M1023_g N_A_329_81#_c_1185_n 0.00688376f $X=5.21 $Y=0.69
+ $X2=0 $Y2=0
cc_515 N_A_1027_48#_c_604_n N_A_329_81#_c_1185_n 0.0024425f $X=5.395 $Y=1.92
+ $X2=0 $Y2=0
cc_516 N_A_1027_48#_c_604_n N_A_329_81#_c_1192_n 0.0196114f $X=5.395 $Y=1.92
+ $X2=0 $Y2=0
cc_517 N_A_1027_48#_c_605_n N_A_329_81#_c_1192_n 0.0192543f $X=6.39 $Y=1.64
+ $X2=0 $Y2=0
cc_518 N_A_1027_48#_c_611_n N_A_329_81#_c_1192_n 0.00862204f $X=6.687 $Y=2.132
+ $X2=0 $Y2=0
cc_519 N_A_1027_48#_c_604_n N_A_329_81#_c_1193_n 0.00184464f $X=5.395 $Y=1.92
+ $X2=0 $Y2=0
cc_520 N_A_1027_48#_c_605_n N_A_329_81#_c_1193_n 0.0217552f $X=6.39 $Y=1.64
+ $X2=0 $Y2=0
cc_521 N_A_1027_48#_c_611_n N_A_329_81#_c_1193_n 0.0318581f $X=6.687 $Y=2.132
+ $X2=0 $Y2=0
cc_522 N_A_1027_48#_c_604_n N_A_329_81#_c_1246_n 6.80962e-19 $X=5.395 $Y=1.92
+ $X2=0 $Y2=0
cc_523 N_A_1027_48#_M1023_g N_VGND_c_1344_n 0.00294228f $X=5.21 $Y=0.69 $X2=0
+ $Y2=0
cc_524 N_A_1027_48#_M1023_g N_VGND_c_1345_n 0.00433139f $X=5.21 $Y=0.69 $X2=0
+ $Y2=0
cc_525 N_A_1027_48#_M1023_g N_VGND_c_1354_n 0.00823312f $X=5.21 $Y=0.69 $X2=0
+ $Y2=0
cc_526 N_C_c_686_n N_A_1057_74#_c_772_n 0.0105426f $X=7.01 $Y=1.765 $X2=0 $Y2=0
cc_527 N_C_c_679_n N_A_1057_74#_c_791_n 0.00798135f $X=5.71 $Y=1.085 $X2=0 $Y2=0
cc_528 N_C_c_679_n N_A_1057_74#_c_764_n 0.0120726f $X=5.71 $Y=1.085 $X2=0 $Y2=0
cc_529 N_C_c_680_n N_A_1057_74#_c_764_n 7.03833e-19 $X=5.95 $Y=1.16 $X2=0 $Y2=0
cc_530 N_C_c_679_n N_A_1057_74#_c_765_n 0.00188363f $X=5.71 $Y=1.085 $X2=0 $Y2=0
cc_531 N_C_c_689_n N_A_1057_74#_c_774_n 0.00814435f $X=6.01 $Y=1.92 $X2=0 $Y2=0
cc_532 N_C_c_686_n N_A_1057_74#_c_774_n 0.0037979f $X=7.01 $Y=1.765 $X2=0 $Y2=0
cc_533 N_C_c_679_n N_A_1057_74#_c_766_n 0.00264822f $X=5.71 $Y=1.085 $X2=0 $Y2=0
cc_534 N_C_c_684_n N_A_1057_74#_c_767_n 3.54962e-19 $X=6.695 $Y=1.425 $X2=0
+ $Y2=0
cc_535 N_C_c_685_n N_A_1057_74#_c_767_n 0.0160581f $X=6.77 $Y=1.35 $X2=0 $Y2=0
cc_536 N_C_c_684_n N_A_1057_74#_c_768_n 0.0014427f $X=6.695 $Y=1.425 $X2=0 $Y2=0
cc_537 N_C_c_686_n N_A_1057_74#_c_775_n 0.0157293f $X=7.01 $Y=1.765 $X2=0 $Y2=0
cc_538 N_C_c_686_n N_A_1057_74#_c_802_n 7.98687e-19 $X=7.01 $Y=1.765 $X2=0 $Y2=0
cc_539 N_C_c_687_n N_A_1057_74#_c_802_n 0.00860034f $X=7.01 $Y=1.515 $X2=0 $Y2=0
cc_540 N_C_c_686_n N_A_1057_74#_c_804_n 0.00126265f $X=7.01 $Y=1.765 $X2=0 $Y2=0
cc_541 N_C_c_687_n N_A_1057_74#_c_804_n 0.0135553f $X=7.01 $Y=1.515 $X2=0 $Y2=0
cc_542 N_C_c_686_n N_A_1057_74#_c_788_n 0.00601579f $X=7.01 $Y=1.765 $X2=0 $Y2=0
cc_543 N_C_c_687_n N_A_1057_74#_c_788_n 0.00901545f $X=7.01 $Y=1.515 $X2=0 $Y2=0
cc_544 N_C_c_686_n N_A_1057_74#_c_776_n 0.00354611f $X=7.01 $Y=1.765 $X2=0 $Y2=0
cc_545 N_C_c_689_n N_A_1057_74#_c_777_n 0.00508269f $X=6.01 $Y=1.92 $X2=0 $Y2=0
cc_546 N_C_c_686_n N_A_1057_74#_c_769_n 0.00221788f $X=7.01 $Y=1.765 $X2=0 $Y2=0
cc_547 N_C_c_687_n N_A_1057_74#_c_769_n 0.026846f $X=7.01 $Y=1.515 $X2=0 $Y2=0
cc_548 N_C_c_685_n N_A_1057_74#_c_770_n 0.00377046f $X=6.77 $Y=1.35 $X2=0 $Y2=0
cc_549 N_C_c_686_n N_A_1057_74#_c_771_n 0.018609f $X=7.01 $Y=1.765 $X2=0 $Y2=0
cc_550 N_C_c_687_n N_A_1057_74#_c_771_n 3.96458e-19 $X=7.01 $Y=1.515 $X2=0 $Y2=0
cc_551 N_C_c_686_n N_VPWR_c_992_n 8.98963e-19 $X=7.01 $Y=1.765 $X2=0 $Y2=0
cc_552 N_C_c_689_n N_VPWR_c_996_n 7.17276e-19 $X=6.01 $Y=1.92 $X2=0 $Y2=0
cc_553 N_C_c_680_n N_A_332_373#_c_1076_n 0.00532259f $X=5.95 $Y=1.16 $X2=0 $Y2=0
cc_554 N_C_c_681_n N_A_332_373#_c_1076_n 0.0108015f $X=5.785 $Y=1.16 $X2=0 $Y2=0
cc_555 N_C_c_682_n N_A_332_373#_c_1076_n 0.00787214f $X=6.01 $Y=1.59 $X2=0 $Y2=0
cc_556 N_C_c_679_n N_A_332_373#_c_1077_n 0.0111838f $X=5.71 $Y=1.085 $X2=0 $Y2=0
cc_557 N_C_c_680_n N_A_332_373#_c_1077_n 0.00410159f $X=5.95 $Y=1.16 $X2=0 $Y2=0
cc_558 N_C_c_682_n N_A_332_373#_c_1077_n 0.00456415f $X=6.01 $Y=1.59 $X2=0 $Y2=0
cc_559 N_C_c_685_n N_A_332_373#_c_1077_n 0.0035702f $X=6.77 $Y=1.35 $X2=0 $Y2=0
cc_560 N_C_c_689_n N_A_332_373#_c_1087_n 0.00108608f $X=6.01 $Y=1.92 $X2=0 $Y2=0
cc_561 N_C_c_689_n N_A_329_81#_c_1192_n 0.0150092f $X=6.01 $Y=1.92 $X2=0 $Y2=0
cc_562 N_C_c_686_n N_A_329_81#_c_1192_n 0.00285906f $X=7.01 $Y=1.765 $X2=0 $Y2=0
cc_563 N_C_c_689_n N_A_329_81#_c_1193_n 0.0100539f $X=6.01 $Y=1.92 $X2=0 $Y2=0
cc_564 N_C_c_684_n N_A_329_81#_c_1193_n 9.00942e-19 $X=6.695 $Y=1.425 $X2=0
+ $Y2=0
cc_565 N_C_c_686_n N_X_c_1313_n 3.05758e-19 $X=7.01 $Y=1.765 $X2=0 $Y2=0
cc_566 N_C_c_679_n N_VGND_c_1345_n 0.00278247f $X=5.71 $Y=1.085 $X2=0 $Y2=0
cc_567 N_C_c_685_n N_VGND_c_1345_n 5.51389e-19 $X=6.77 $Y=1.35 $X2=0 $Y2=0
cc_568 N_C_c_685_n N_VGND_c_1353_n 7.18285e-19 $X=6.77 $Y=1.35 $X2=0 $Y2=0
cc_569 N_C_c_679_n N_VGND_c_1354_n 0.00359137f $X=5.71 $Y=1.085 $X2=0 $Y2=0
cc_570 N_A_1057_74#_c_775_n N_VPWR_M1017_d 0.00429932f $X=7.125 $Y=2.905 $X2=0
+ $Y2=0
cc_571 N_A_1057_74#_c_816_p N_VPWR_M1017_d 0.0190037f $X=7.41 $Y=2.035 $X2=0
+ $Y2=0
cc_572 N_A_1057_74#_c_788_n N_VPWR_M1017_d 0.00191279f $X=7.21 $Y=2.035 $X2=0
+ $Y2=0
cc_573 N_A_1057_74#_c_776_n N_VPWR_M1017_d 0.00223887f $X=7.495 $Y=1.95 $X2=0
+ $Y2=0
cc_574 N_A_1057_74#_c_772_n N_VPWR_c_992_n 0.00674914f $X=7.69 $Y=1.765 $X2=0
+ $Y2=0
cc_575 N_A_1057_74#_c_774_n N_VPWR_c_992_n 0.0142847f $X=7.04 $Y=2.99 $X2=0
+ $Y2=0
cc_576 N_A_1057_74#_c_775_n N_VPWR_c_992_n 0.0451978f $X=7.125 $Y=2.905 $X2=0
+ $Y2=0
cc_577 N_A_1057_74#_c_816_p N_VPWR_c_992_n 0.0148103f $X=7.41 $Y=2.035 $X2=0
+ $Y2=0
cc_578 N_A_1057_74#_c_771_n N_VPWR_c_992_n 3.98939e-19 $X=8.14 $Y=1.552 $X2=0
+ $Y2=0
cc_579 N_A_1057_74#_c_773_n N_VPWR_c_994_n 0.00981831f $X=8.14 $Y=1.765 $X2=0
+ $Y2=0
cc_580 N_A_1057_74#_c_774_n N_VPWR_c_996_n 0.0878491f $X=7.04 $Y=2.99 $X2=0
+ $Y2=0
cc_581 N_A_1057_74#_c_777_n N_VPWR_c_996_n 0.0223379f $X=5.7 $Y=2.82 $X2=0 $Y2=0
cc_582 N_A_1057_74#_c_772_n N_VPWR_c_997_n 0.00445602f $X=7.69 $Y=1.765 $X2=0
+ $Y2=0
cc_583 N_A_1057_74#_c_773_n N_VPWR_c_997_n 0.00428607f $X=8.14 $Y=1.765 $X2=0
+ $Y2=0
cc_584 N_A_1057_74#_c_772_n N_VPWR_c_989_n 0.00862391f $X=7.69 $Y=1.765 $X2=0
+ $Y2=0
cc_585 N_A_1057_74#_c_773_n N_VPWR_c_989_n 0.00806037f $X=8.14 $Y=1.765 $X2=0
+ $Y2=0
cc_586 N_A_1057_74#_c_774_n N_VPWR_c_989_n 0.0507826f $X=7.04 $Y=2.99 $X2=0
+ $Y2=0
cc_587 N_A_1057_74#_c_777_n N_VPWR_c_989_n 0.0125334f $X=5.7 $Y=2.82 $X2=0 $Y2=0
cc_588 N_A_1057_74#_c_764_n N_A_332_373#_M1019_d 0.00349202f $X=6.33 $Y=0.34
+ $X2=0 $Y2=0
cc_589 N_A_1057_74#_c_791_n N_A_332_373#_c_1076_n 0.0239462f $X=5.495 $Y=0.495
+ $X2=0 $Y2=0
cc_590 N_A_1057_74#_c_764_n N_A_332_373#_c_1077_n 0.0242638f $X=6.33 $Y=0.34
+ $X2=0 $Y2=0
cc_591 N_A_1057_74#_c_766_n N_A_332_373#_c_1077_n 0.00511588f $X=6.415 $Y=0.66
+ $X2=0 $Y2=0
cc_592 N_A_1057_74#_c_768_n N_A_332_373#_c_1077_n 0.0150383f $X=6.5 $Y=0.745
+ $X2=0 $Y2=0
cc_593 N_A_1057_74#_c_765_n N_A_329_81#_c_1184_n 0.00373319f $X=5.66 $Y=0.34
+ $X2=0 $Y2=0
cc_594 N_A_1057_74#_M1021_d N_A_329_81#_c_1192_n 0.0113203f $X=5.47 $Y=1.995
+ $X2=0 $Y2=0
cc_595 N_A_1057_74#_c_774_n N_A_329_81#_c_1192_n 0.0233426f $X=7.04 $Y=2.99
+ $X2=0 $Y2=0
cc_596 N_A_1057_74#_c_777_n N_A_329_81#_c_1192_n 0.0244725f $X=5.7 $Y=2.82 $X2=0
+ $Y2=0
cc_597 N_A_1057_74#_c_772_n N_X_c_1312_n 0.012186f $X=7.69 $Y=1.765 $X2=0 $Y2=0
cc_598 N_A_1057_74#_c_773_n N_X_c_1312_n 0.0119183f $X=8.14 $Y=1.765 $X2=0 $Y2=0
cc_599 N_A_1057_74#_c_775_n N_X_c_1312_n 0.00508722f $X=7.125 $Y=2.905 $X2=0
+ $Y2=0
cc_600 N_A_1057_74#_c_772_n N_X_c_1313_n 0.00234892f $X=7.69 $Y=1.765 $X2=0
+ $Y2=0
cc_601 N_A_1057_74#_c_773_n N_X_c_1313_n 0.00195791f $X=8.14 $Y=1.765 $X2=0
+ $Y2=0
cc_602 N_A_1057_74#_c_771_n N_X_c_1313_n 0.00374722f $X=8.14 $Y=1.552 $X2=0
+ $Y2=0
cc_603 N_A_1057_74#_c_762_n N_X_c_1310_n 9.57805e-19 $X=7.715 $Y=1.34 $X2=0
+ $Y2=0
cc_604 N_A_1057_74#_c_773_n N_X_c_1310_n 0.00342409f $X=8.14 $Y=1.765 $X2=0
+ $Y2=0
cc_605 N_A_1057_74#_c_763_n N_X_c_1310_n 0.00556338f $X=8.145 $Y=1.34 $X2=0
+ $Y2=0
cc_606 N_A_1057_74#_c_776_n N_X_c_1310_n 0.005496f $X=7.495 $Y=1.95 $X2=0 $Y2=0
cc_607 N_A_1057_74#_c_769_n N_X_c_1310_n 0.0238938f $X=7.59 $Y=1.505 $X2=0 $Y2=0
cc_608 N_A_1057_74#_c_770_n N_X_c_1310_n 0.00546742f $X=7.582 $Y=1.34 $X2=0
+ $Y2=0
cc_609 N_A_1057_74#_c_771_n N_X_c_1310_n 0.0317044f $X=8.14 $Y=1.552 $X2=0 $Y2=0
cc_610 N_A_1057_74#_c_762_n X 0.0123221f $X=7.715 $Y=1.34 $X2=0 $Y2=0
cc_611 N_A_1057_74#_c_763_n X 0.00701411f $X=8.145 $Y=1.34 $X2=0 $Y2=0
cc_612 N_A_1057_74#_c_762_n X 0.00258445f $X=7.715 $Y=1.34 $X2=0 $Y2=0
cc_613 N_A_1057_74#_c_763_n X 0.00180034f $X=8.145 $Y=1.34 $X2=0 $Y2=0
cc_614 N_A_1057_74#_c_802_n X 0.0123899f $X=7.41 $Y=1.095 $X2=0 $Y2=0
cc_615 N_A_1057_74#_c_771_n X 0.00131295f $X=8.14 $Y=1.552 $X2=0 $Y2=0
cc_616 N_A_1057_74#_c_767_n N_VGND_M1010_d 0.00352419f $X=6.89 $Y=0.745 $X2=0
+ $Y2=0
cc_617 N_A_1057_74#_c_862_p N_VGND_M1010_d 0.00320933f $X=6.975 $Y=1.01 $X2=0
+ $Y2=0
cc_618 N_A_1057_74#_c_802_n N_VGND_M1010_d 0.0227231f $X=7.41 $Y=1.095 $X2=0
+ $Y2=0
cc_619 N_A_1057_74#_c_804_n N_VGND_M1010_d 0.00276146f $X=7.06 $Y=1.095 $X2=0
+ $Y2=0
cc_620 N_A_1057_74#_c_770_n N_VGND_M1010_d 0.00133582f $X=7.582 $Y=1.34 $X2=0
+ $Y2=0
cc_621 N_A_1057_74#_c_764_n N_VGND_c_1345_n 0.0547745f $X=6.33 $Y=0.34 $X2=0
+ $Y2=0
cc_622 N_A_1057_74#_c_765_n N_VGND_c_1345_n 0.0236456f $X=5.66 $Y=0.34 $X2=0
+ $Y2=0
cc_623 N_A_1057_74#_c_767_n N_VGND_c_1345_n 0.00691154f $X=6.89 $Y=0.745 $X2=0
+ $Y2=0
cc_624 N_A_1057_74#_c_763_n N_VGND_c_1347_n 0.00595876f $X=8.145 $Y=1.34 $X2=0
+ $Y2=0
cc_625 N_A_1057_74#_c_762_n N_VGND_c_1350_n 0.00472938f $X=7.715 $Y=1.34 $X2=0
+ $Y2=0
cc_626 N_A_1057_74#_c_763_n N_VGND_c_1350_n 0.00472938f $X=8.145 $Y=1.34 $X2=0
+ $Y2=0
cc_627 N_A_1057_74#_c_762_n N_VGND_c_1353_n 0.0115709f $X=7.715 $Y=1.34 $X2=0
+ $Y2=0
cc_628 N_A_1057_74#_c_764_n N_VGND_c_1353_n 0.0087818f $X=6.33 $Y=0.34 $X2=0
+ $Y2=0
cc_629 N_A_1057_74#_c_766_n N_VGND_c_1353_n 0.00301349f $X=6.415 $Y=0.66 $X2=0
+ $Y2=0
cc_630 N_A_1057_74#_c_767_n N_VGND_c_1353_n 0.0280097f $X=6.89 $Y=0.745 $X2=0
+ $Y2=0
cc_631 N_A_1057_74#_c_862_p N_VGND_c_1353_n 7.35861e-19 $X=6.975 $Y=1.01 $X2=0
+ $Y2=0
cc_632 N_A_1057_74#_c_802_n N_VGND_c_1353_n 0.0358553f $X=7.41 $Y=1.095 $X2=0
+ $Y2=0
cc_633 N_A_1057_74#_c_771_n N_VGND_c_1353_n 6.33745e-19 $X=8.14 $Y=1.552 $X2=0
+ $Y2=0
cc_634 N_A_1057_74#_c_762_n N_VGND_c_1354_n 0.00508379f $X=7.715 $Y=1.34 $X2=0
+ $Y2=0
cc_635 N_A_1057_74#_c_763_n N_VGND_c_1354_n 0.00508379f $X=8.145 $Y=1.34 $X2=0
+ $Y2=0
cc_636 N_A_1057_74#_c_764_n N_VGND_c_1354_n 0.0311946f $X=6.33 $Y=0.34 $X2=0
+ $Y2=0
cc_637 N_A_1057_74#_c_765_n N_VGND_c_1354_n 0.0127298f $X=5.66 $Y=0.34 $X2=0
+ $Y2=0
cc_638 N_A_1057_74#_c_767_n N_VGND_c_1354_n 0.0119702f $X=6.89 $Y=0.745 $X2=0
+ $Y2=0
cc_639 N_A_27_373#_c_898_n N_VPWR_c_990_n 0.0394805f $X=0.28 $Y=2.375 $X2=0
+ $Y2=0
cc_640 N_A_27_373#_c_898_n N_VPWR_c_998_n 0.0114601f $X=0.28 $Y=2.375 $X2=0
+ $Y2=0
cc_641 N_A_27_373#_c_898_n N_VPWR_c_989_n 0.0124049f $X=0.28 $Y=2.375 $X2=0
+ $Y2=0
cc_642 N_A_27_373#_c_895_n N_A_332_373#_M1005_d 0.00760845f $X=2.275 $Y=2.65
+ $X2=0 $Y2=0
cc_643 N_A_27_373#_c_886_n N_A_332_373#_c_1083_n 0.0310635f $X=1.63 $Y=2.565
+ $X2=0 $Y2=0
cc_644 N_A_27_373#_c_895_n N_A_332_373#_c_1083_n 0.0161276f $X=2.275 $Y=2.65
+ $X2=0 $Y2=0
cc_645 N_A_27_373#_c_887_n N_A_332_373#_c_1072_n 0.00203691f $X=2.135 $Y=1.272
+ $X2=0 $Y2=0
cc_646 N_A_27_373#_c_897_n N_A_332_373#_c_1072_n 0.0221295f $X=2.44 $Y=2.01
+ $X2=0 $Y2=0
cc_647 N_A_27_373#_c_889_n N_A_332_373#_c_1072_n 0.0190342f $X=2.275 $Y=1.11
+ $X2=0 $Y2=0
cc_648 N_A_27_373#_c_886_n N_A_332_373#_c_1073_n 0.0143553f $X=1.63 $Y=2.565
+ $X2=0 $Y2=0
cc_649 N_A_27_373#_c_887_n N_A_332_373#_c_1073_n 0.0184143f $X=2.135 $Y=1.272
+ $X2=0 $Y2=0
cc_650 N_A_27_373#_c_889_n N_A_332_373#_c_1078_n 0.0240865f $X=2.275 $Y=1.11
+ $X2=0 $Y2=0
cc_651 N_A_27_373#_M1002_d N_A_332_373#_c_1080_n 7.00965e-19 $X=2.135 $Y=0.845
+ $X2=0 $Y2=0
cc_652 N_A_27_373#_c_897_n N_A_332_373#_c_1080_n 3.54735e-19 $X=2.44 $Y=2.01
+ $X2=0 $Y2=0
cc_653 N_A_27_373#_c_889_n N_A_332_373#_c_1080_n 0.00607915f $X=2.275 $Y=1.11
+ $X2=0 $Y2=0
cc_654 N_A_27_373#_c_889_n N_A_332_373#_c_1081_n 0.00608382f $X=2.275 $Y=1.11
+ $X2=0 $Y2=0
cc_655 N_A_27_373#_c_887_n N_A_329_81#_M1018_d 0.00206654f $X=2.135 $Y=1.272
+ $X2=-0.19 $Y2=-0.245
cc_656 N_A_27_373#_c_897_n N_A_329_81#_c_1211_n 0.029367f $X=2.44 $Y=2.01 $X2=0
+ $Y2=0
cc_657 N_A_27_373#_c_895_n N_A_329_81#_c_1190_n 0.00347496f $X=2.275 $Y=2.65
+ $X2=0 $Y2=0
cc_658 N_A_27_373#_c_897_n N_A_329_81#_c_1190_n 0.0125953f $X=2.44 $Y=2.01 $X2=0
+ $Y2=0
cc_659 N_A_27_373#_c_885_n N_A_329_81#_c_1186_n 0.00510362f $X=1.63 $Y=1.38
+ $X2=0 $Y2=0
cc_660 N_A_27_373#_c_887_n N_A_329_81#_c_1186_n 0.0160417f $X=2.135 $Y=1.272
+ $X2=0 $Y2=0
cc_661 N_A_27_373#_c_893_n N_A_329_81#_c_1186_n 0.00154277f $X=1.68 $Y=1.295
+ $X2=0 $Y2=0
cc_662 N_A_27_373#_M1002_d N_A_329_81#_c_1187_n 0.00349911f $X=2.135 $Y=0.845
+ $X2=0 $Y2=0
cc_663 N_A_27_373#_c_887_n N_A_329_81#_c_1187_n 0.00580419f $X=2.135 $Y=1.272
+ $X2=0 $Y2=0
cc_664 N_A_27_373#_c_889_n N_A_329_81#_c_1187_n 0.0172834f $X=2.275 $Y=1.11
+ $X2=0 $Y2=0
cc_665 N_A_27_373#_c_884_n N_VGND_c_1343_n 0.0179595f $X=0.32 $Y=0.55 $X2=0
+ $Y2=0
cc_666 N_A_27_373#_c_890_n N_VGND_c_1343_n 8.78751e-19 $X=1.535 $Y=1.295 $X2=0
+ $Y2=0
cc_667 N_A_27_373#_c_884_n N_VGND_c_1348_n 0.0124374f $X=0.32 $Y=0.55 $X2=0
+ $Y2=0
cc_668 N_A_27_373#_c_884_n N_VGND_c_1354_n 0.0114937f $X=0.32 $Y=0.55 $X2=0
+ $Y2=0
cc_669 N_VPWR_M1020_d N_A_329_81#_c_1189_n 0.00694562f $X=4.39 $Y=1.84 $X2=0
+ $Y2=0
cc_670 N_VPWR_c_991_n N_A_329_81#_c_1189_n 0.00908439f $X=4.62 $Y=2.9 $X2=0
+ $Y2=0
cc_671 N_VPWR_c_989_n N_A_329_81#_c_1189_n 0.0273817f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_672 N_VPWR_M1020_d N_A_329_81#_c_1185_n 0.0170324f $X=4.39 $Y=1.84 $X2=0
+ $Y2=0
cc_673 N_VPWR_c_991_n N_A_329_81#_c_1192_n 0.00232914f $X=4.62 $Y=2.9 $X2=0
+ $Y2=0
cc_674 N_VPWR_c_989_n N_A_329_81#_c_1192_n 0.0284422f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_675 N_VPWR_M1020_d N_A_329_81#_c_1246_n 0.00448587f $X=4.39 $Y=1.84 $X2=0
+ $Y2=0
cc_676 N_VPWR_c_991_n N_A_329_81#_c_1246_n 0.0147528f $X=4.62 $Y=2.9 $X2=0 $Y2=0
cc_677 N_VPWR_c_989_n N_A_329_81#_c_1246_n 6.89689e-19 $X=8.4 $Y=3.33 $X2=0
+ $Y2=0
cc_678 N_VPWR_c_992_n N_X_c_1312_n 0.045127f $X=7.465 $Y=2.455 $X2=0 $Y2=0
cc_679 N_VPWR_c_997_n N_X_c_1312_n 0.0151764f $X=8.28 $Y=3.33 $X2=0 $Y2=0
cc_680 N_VPWR_c_989_n N_X_c_1312_n 0.0124607f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_681 N_VPWR_c_994_n N_X_c_1310_n 0.0829236f $X=8.365 $Y=1.985 $X2=0 $Y2=0
cc_682 N_VPWR_c_994_n N_VGND_c_1347_n 0.00977564f $X=8.365 $Y=1.985 $X2=0 $Y2=0
cc_683 N_A_332_373#_M1001_d N_A_329_81#_c_1183_n 0.00218533f $X=2.645 $Y=0.625
+ $X2=0 $Y2=0
cc_684 N_A_332_373#_c_1079_n N_A_329_81#_c_1183_n 0.0256726f $X=4.895 $Y=1.295
+ $X2=0 $Y2=0
cc_685 N_A_332_373#_c_1078_n N_A_329_81#_c_1211_n 0.00277093f $X=2.8 $Y=1.12
+ $X2=0 $Y2=0
cc_686 N_A_332_373#_c_1079_n N_A_329_81#_c_1211_n 0.0088124f $X=4.895 $Y=1.295
+ $X2=0 $Y2=0
cc_687 N_A_332_373#_c_1074_n N_A_329_81#_c_1184_n 0.0169928f $X=5.04 $Y=1.305
+ $X2=0 $Y2=0
cc_688 N_A_332_373#_c_1076_n N_A_329_81#_c_1184_n 3.08288e-19 $X=5.83 $Y=1.22
+ $X2=0 $Y2=0
cc_689 N_A_332_373#_c_1079_n N_A_329_81#_c_1184_n 0.00643723f $X=4.895 $Y=1.295
+ $X2=0 $Y2=0
cc_690 N_A_332_373#_c_1082_n N_A_329_81#_c_1184_n 0.0032994f $X=5.04 $Y=1.295
+ $X2=0 $Y2=0
cc_691 N_A_332_373#_c_1074_n N_A_329_81#_c_1185_n 0.0126364f $X=5.04 $Y=1.305
+ $X2=0 $Y2=0
cc_692 N_A_332_373#_c_1075_n N_A_329_81#_c_1185_n 0.0505384f $X=5.04 $Y=1.975
+ $X2=0 $Y2=0
cc_693 N_A_332_373#_c_1087_n N_A_329_81#_c_1185_n 0.0197685f $X=5.17 $Y=2.14
+ $X2=0 $Y2=0
cc_694 N_A_332_373#_c_1079_n N_A_329_81#_c_1185_n 0.0264059f $X=4.895 $Y=1.295
+ $X2=0 $Y2=0
cc_695 N_A_332_373#_c_1082_n N_A_329_81#_c_1185_n 0.0026622f $X=5.04 $Y=1.295
+ $X2=0 $Y2=0
cc_696 N_A_332_373#_M1021_s N_A_329_81#_c_1192_n 0.00776593f $X=5.03 $Y=1.995
+ $X2=0 $Y2=0
cc_697 N_A_332_373#_c_1087_n N_A_329_81#_c_1192_n 0.0265436f $X=5.17 $Y=2.14
+ $X2=0 $Y2=0
cc_698 N_A_332_373#_c_1080_n N_A_329_81#_c_1187_n 0.00180844f $X=2.785 $Y=1.295
+ $X2=0 $Y2=0
cc_699 N_A_332_373#_M1001_d N_A_329_81#_c_1188_n 2.36577e-19 $X=2.645 $Y=0.625
+ $X2=0 $Y2=0
cc_700 N_A_332_373#_c_1078_n N_A_329_81#_c_1188_n 0.0233474f $X=2.8 $Y=1.12
+ $X2=0 $Y2=0
cc_701 N_A_332_373#_c_1080_n N_A_329_81#_c_1188_n 0.00102588f $X=2.785 $Y=1.295
+ $X2=0 $Y2=0
cc_702 N_A_329_81#_c_1183_n N_VGND_M1014_d 0.00993346f $X=4.585 $Y=0.7 $X2=0
+ $Y2=0
cc_703 N_A_329_81#_c_1183_n N_VGND_c_1344_n 0.0237317f $X=4.585 $Y=0.7 $X2=0
+ $Y2=0
cc_704 N_A_329_81#_c_1184_n N_VGND_c_1344_n 0.00764375f $X=4.67 $Y=0.965 $X2=0
+ $Y2=0
cc_705 N_A_329_81#_c_1184_n N_VGND_c_1345_n 0.0193145f $X=4.67 $Y=0.965 $X2=0
+ $Y2=0
cc_706 N_A_329_81#_c_1183_n N_VGND_c_1349_n 0.0126356f $X=4.585 $Y=0.7 $X2=0
+ $Y2=0
cc_707 N_A_329_81#_c_1183_n N_VGND_c_1354_n 0.0244914f $X=4.585 $Y=0.7 $X2=0
+ $Y2=0
cc_708 N_A_329_81#_c_1184_n N_VGND_c_1354_n 0.0191643f $X=4.67 $Y=0.965 $X2=0
+ $Y2=0
cc_709 X N_VGND_c_1347_n 0.0316671f $X=7.835 $Y=0.47 $X2=0 $Y2=0
cc_710 X N_VGND_c_1350_n 0.0105983f $X=7.835 $Y=0.47 $X2=0 $Y2=0
cc_711 X N_VGND_c_1353_n 0.0165965f $X=7.835 $Y=0.47 $X2=0 $Y2=0
cc_712 X N_VGND_c_1354_n 0.0113894f $X=7.835 $Y=0.47 $X2=0 $Y2=0
