* File: sky130_fd_sc_ls__nand4b_1.spice
* Created: Wed Sep  2 11:13:07 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__nand4b_1.pex.spice"
.subckt sky130_fd_sc_ls__nand4b_1  VNB VPB A_N D C B VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B	B
* C	C
* D	D
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1007 N_VGND_M1007_d N_A_N_M1007_g N_A_27_112#_M1007_s VNB NSHORT L=0.15 W=0.55
+ AD=0.114946 AS=0.2695 PD=0.963566 PS=2.08 NRD=23.988 NRS=0 M=1 R=3.66667
+ SA=75000.4 SB=75002.4 A=0.0825 P=1.4 MULT=1
MM1008 A_263_74# N_D_M1008_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.74 AD=0.0888
+ AS=0.154654 PD=0.98 PS=1.29643 NRD=10.536 NRS=0.804 M=1 R=4.93333 SA=75000.8
+ SB=75001.8 A=0.111 P=1.78 MULT=1
MM1009 A_341_74# N_C_M1009_g A_263_74# VNB NSHORT L=0.15 W=0.74 AD=0.1332
+ AS=0.0888 PD=1.1 PS=0.98 NRD=20.268 NRS=10.536 M=1 R=4.93333 SA=75001.2
+ SB=75001.4 A=0.111 P=1.78 MULT=1
MM1001 A_443_74# N_B_M1001_g A_341_74# VNB NSHORT L=0.15 W=0.74 AD=0.1443
+ AS=0.1332 PD=1.13 PS=1.1 NRD=22.692 NRS=20.268 M=1 R=4.93333 SA=75001.7
+ SB=75000.9 A=0.111 P=1.78 MULT=1
MM1002 N_Y_M1002_d N_A_27_112#_M1002_g A_443_74# VNB NSHORT L=0.15 W=0.74
+ AD=0.3404 AS=0.1443 PD=2.4 PS=1.13 NRD=15.396 NRS=22.692 M=1 R=4.93333
+ SA=75002.2 SB=75000.4 A=0.111 P=1.78 MULT=1
MM1000 N_VPWR_M1000_d N_A_N_M1000_g N_A_27_112#_M1000_s VPB PHIGHVT L=0.15
+ W=0.84 AD=0.198 AS=0.2478 PD=1.33286 PS=2.27 NRD=22.261 NRS=2.3443 M=1 R=5.6
+ SA=75000.2 SB=75002.3 A=0.126 P=1.98 MULT=1
MM1003 N_Y_M1003_d N_D_M1003_g N_VPWR_M1000_d VPB PHIGHVT L=0.15 W=1.12 AD=0.168
+ AS=0.264 PD=1.42 PS=1.77714 NRD=1.7533 NRS=10.5395 M=1 R=7.46667 SA=75000.7
+ SB=75001.7 A=0.168 P=2.54 MULT=1
MM1005 N_VPWR_M1005_d N_C_M1005_g N_Y_M1003_d VPB PHIGHVT L=0.15 W=1.12
+ AD=0.2352 AS=0.168 PD=1.54 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75001.3 A=0.168 P=2.54 MULT=1
MM1004 N_Y_M1004_d N_B_M1004_g N_VPWR_M1005_d VPB PHIGHVT L=0.15 W=1.12 AD=0.168
+ AS=0.2352 PD=1.42 PS=1.54 NRD=1.7533 NRS=14.0658 M=1 R=7.46667 SA=75001.7
+ SB=75000.7 A=0.168 P=2.54 MULT=1
MM1006 N_VPWR_M1006_d N_A_27_112#_M1006_g N_Y_M1004_d VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3864 AS=0.168 PD=2.93 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75002.1 SB=75000.3 A=0.168 P=2.54 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9564 P=11.2
*
.include "sky130_fd_sc_ls__nand4b_1.pxi.spice"
*
.ends
*
*
