* File: sky130_fd_sc_ls__dlxbp_1.pxi.spice
* Created: Wed Sep  2 11:04:33 2020
* 
x_PM_SKY130_FD_SC_LS__DLXBP_1%D N_D_c_143_n N_D_M1003_g N_D_c_148_n N_D_M1017_g
+ D N_D_c_145_n N_D_c_146_n PM_SKY130_FD_SC_LS__DLXBP_1%D
x_PM_SKY130_FD_SC_LS__DLXBP_1%GATE N_GATE_M1001_g N_GATE_c_183_n N_GATE_c_188_n
+ N_GATE_M1021_g GATE N_GATE_c_185_n N_GATE_c_186_n
+ PM_SKY130_FD_SC_LS__DLXBP_1%GATE
x_PM_SKY130_FD_SC_LS__DLXBP_1%A_231_74# N_A_231_74#_M1001_d N_A_231_74#_M1021_d
+ N_A_231_74#_M1016_g N_A_231_74#_c_234_n N_A_231_74#_M1014_g
+ N_A_231_74#_c_235_n N_A_231_74#_M1000_g N_A_231_74#_c_236_n
+ N_A_231_74#_c_237_n N_A_231_74#_M1002_g N_A_231_74#_c_239_n
+ N_A_231_74#_c_225_n N_A_231_74#_c_226_n N_A_231_74#_c_227_n
+ N_A_231_74#_c_228_n N_A_231_74#_c_229_n N_A_231_74#_c_230_n
+ N_A_231_74#_c_231_n N_A_231_74#_c_232_n N_A_231_74#_c_233_n
+ PM_SKY130_FD_SC_LS__DLXBP_1%A_231_74#
x_PM_SKY130_FD_SC_LS__DLXBP_1%A_27_413# N_A_27_413#_M1003_s N_A_27_413#_M1017_s
+ N_A_27_413#_c_357_n N_A_27_413#_M1012_g N_A_27_413#_M1010_g
+ N_A_27_413#_c_363_n N_A_27_413#_c_364_n N_A_27_413#_c_365_n
+ N_A_27_413#_c_366_n N_A_27_413#_c_367_n N_A_27_413#_c_368_n
+ N_A_27_413#_c_359_n N_A_27_413#_c_360_n N_A_27_413#_c_370_n
+ N_A_27_413#_c_361_n PM_SKY130_FD_SC_LS__DLXBP_1%A_27_413#
x_PM_SKY130_FD_SC_LS__DLXBP_1%A_373_82# N_A_373_82#_M1016_s N_A_373_82#_M1014_s
+ N_A_373_82#_M1009_g N_A_373_82#_c_458_n N_A_373_82#_M1005_g
+ N_A_373_82#_c_452_n N_A_373_82#_c_471_n N_A_373_82#_c_453_n
+ N_A_373_82#_c_460_n N_A_373_82#_c_461_n N_A_373_82#_c_454_n
+ N_A_373_82#_c_462_n N_A_373_82#_c_455_n N_A_373_82#_c_456_n
+ N_A_373_82#_c_490_n N_A_373_82#_c_457_n PM_SKY130_FD_SC_LS__DLXBP_1%A_373_82#
x_PM_SKY130_FD_SC_LS__DLXBP_1%A_863_98# N_A_863_98#_M1006_d N_A_863_98#_M1011_d
+ N_A_863_98#_M1018_g N_A_863_98#_c_578_n N_A_863_98#_c_579_n
+ N_A_863_98#_c_580_n N_A_863_98#_M1007_g N_A_863_98#_c_581_n
+ N_A_863_98#_M1019_g N_A_863_98#_M1013_g N_A_863_98#_c_568_n
+ N_A_863_98#_c_569_n N_A_863_98#_c_584_n N_A_863_98#_M1020_g
+ N_A_863_98#_M1015_g N_A_863_98#_c_571_n N_A_863_98#_c_585_n
+ N_A_863_98#_c_572_n N_A_863_98#_c_573_n N_A_863_98#_c_574_n
+ N_A_863_98#_c_587_n N_A_863_98#_c_575_n N_A_863_98#_c_576_n
+ N_A_863_98#_c_588_n PM_SKY130_FD_SC_LS__DLXBP_1%A_863_98#
x_PM_SKY130_FD_SC_LS__DLXBP_1%A_664_392# N_A_664_392#_M1009_d
+ N_A_664_392#_M1000_d N_A_664_392#_M1006_g N_A_664_392#_c_685_n
+ N_A_664_392#_M1011_g N_A_664_392#_c_696_n N_A_664_392#_c_692_n
+ N_A_664_392#_c_686_n N_A_664_392#_c_687_n N_A_664_392#_c_688_n
+ N_A_664_392#_c_689_n N_A_664_392#_c_690_n N_A_664_392#_c_708_n
+ PM_SKY130_FD_SC_LS__DLXBP_1%A_664_392#
x_PM_SKY130_FD_SC_LS__DLXBP_1%A_1347_424# N_A_1347_424#_M1015_d
+ N_A_1347_424#_M1020_d N_A_1347_424#_c_775_n N_A_1347_424#_M1004_g
+ N_A_1347_424#_M1008_g N_A_1347_424#_c_770_n N_A_1347_424#_c_771_n
+ N_A_1347_424#_c_772_n N_A_1347_424#_c_773_n N_A_1347_424#_c_774_n
+ PM_SKY130_FD_SC_LS__DLXBP_1%A_1347_424#
x_PM_SKY130_FD_SC_LS__DLXBP_1%VPWR N_VPWR_M1017_d N_VPWR_M1014_d N_VPWR_M1007_d
+ N_VPWR_M1019_d N_VPWR_M1004_s N_VPWR_c_814_n N_VPWR_c_815_n N_VPWR_c_816_n
+ N_VPWR_c_817_n N_VPWR_c_818_n N_VPWR_c_819_n N_VPWR_c_820_n N_VPWR_c_821_n
+ N_VPWR_c_822_n N_VPWR_c_823_n VPWR N_VPWR_c_824_n N_VPWR_c_825_n
+ N_VPWR_c_813_n N_VPWR_c_827_n N_VPWR_c_828_n N_VPWR_c_829_n
+ PM_SKY130_FD_SC_LS__DLXBP_1%VPWR
x_PM_SKY130_FD_SC_LS__DLXBP_1%Q N_Q_M1013_s N_Q_M1019_s N_Q_c_912_n N_Q_c_913_n
+ N_Q_c_909_n Q Q Q PM_SKY130_FD_SC_LS__DLXBP_1%Q
x_PM_SKY130_FD_SC_LS__DLXBP_1%Q_N N_Q_N_M1008_d N_Q_N_M1004_d Q_N Q_N Q_N Q_N
+ Q_N Q_N Q_N PM_SKY130_FD_SC_LS__DLXBP_1%Q_N
x_PM_SKY130_FD_SC_LS__DLXBP_1%VGND N_VGND_M1003_d N_VGND_M1016_d N_VGND_M1018_d
+ N_VGND_M1013_d N_VGND_M1008_s N_VGND_c_962_n N_VGND_c_963_n N_VGND_c_964_n
+ N_VGND_c_965_n N_VGND_c_966_n N_VGND_c_967_n VGND N_VGND_c_968_n
+ N_VGND_c_969_n N_VGND_c_970_n N_VGND_c_971_n N_VGND_c_972_n N_VGND_c_973_n
+ N_VGND_c_974_n N_VGND_c_975_n N_VGND_c_976_n PM_SKY130_FD_SC_LS__DLXBP_1%VGND
cc_1 VNB N_D_c_143_n 0.0192767f $X=-0.19 $Y=-0.245 $X2=0.587 $Y2=1.713
cc_2 VNB D 0.0038285f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_3 VNB N_D_c_145_n 0.0199975f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.385
cc_4 VNB N_D_c_146_n 0.0220891f $X=-0.19 $Y=-0.245 $X2=0.587 $Y2=1.22
cc_5 VNB N_GATE_c_183_n 0.00677649f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.835
cc_6 VNB GATE 0.00380422f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_7 VNB N_GATE_c_185_n 0.034476f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.385
cc_8 VNB N_GATE_c_186_n 0.0229286f $X=-0.19 $Y=-0.245 $X2=0.587 $Y2=1.22
cc_9 VNB N_A_231_74#_M1016_g 0.0363558f $X=-0.19 $Y=-0.245 $X2=0.587 $Y2=1.385
cc_10 VNB N_A_231_74#_M1002_g 0.0409372f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_231_74#_c_225_n 0.0100597f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_231_74#_c_226_n 0.0098903f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_231_74#_c_227_n 0.0017069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_231_74#_c_228_n 0.00127767f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_231_74#_c_229_n 0.036619f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_231_74#_c_230_n 0.00163443f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_231_74#_c_231_n 0.0102682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_231_74#_c_232_n 0.0439804f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_231_74#_c_233_n 0.0197237f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_27_413#_c_357_n 0.0228467f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.485
cc_21 VNB N_A_27_413#_M1010_g 0.0345878f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.385
cc_22 VNB N_A_27_413#_c_359_n 0.00282947f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_27_413#_c_360_n 0.0239006f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_27_413#_c_361_n 0.0281735f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_373_82#_c_452_n 0.0136924f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.385
cc_26 VNB N_A_373_82#_c_453_n 0.0037425f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_373_82#_c_454_n 0.00494001f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_373_82#_c_455_n 0.00686485f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_373_82#_c_456_n 0.0317275f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_373_82#_c_457_n 0.0154994f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_863_98#_M1018_g 0.0457697f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_32 VNB N_A_863_98#_M1013_g 0.0266486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_863_98#_c_568_n 0.0453248f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_863_98#_c_569_n 6.02304e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_863_98#_M1015_g 0.0250484f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_863_98#_c_571_n 0.0726176f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_863_98#_c_572_n 0.0115916f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_863_98#_c_573_n 0.007198f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_863_98#_c_574_n 7.02248e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_863_98#_c_575_n 0.00268063f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_863_98#_c_576_n 0.00432868f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_664_392#_M1006_g 0.0237086f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_43 VNB N_A_664_392#_c_685_n 0.052845f $X=-0.19 $Y=-0.245 $X2=0.587 $Y2=1.385
cc_44 VNB N_A_664_392#_c_686_n 0.00766084f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_664_392#_c_687_n 0.00246517f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_664_392#_c_688_n 0.00590121f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_664_392#_c_689_n 0.0131066f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_664_392#_c_690_n 0.00452768f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_1347_424#_M1008_g 0.0308289f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.385
cc_50 VNB N_A_1347_424#_c_770_n 0.06715f $X=-0.19 $Y=-0.245 $X2=0.587 $Y2=1.22
cc_51 VNB N_A_1347_424#_c_771_n 0.0178423f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.555
cc_52 VNB N_A_1347_424#_c_772_n 0.0118603f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_1347_424#_c_773_n 8.08981e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_1347_424#_c_774_n 0.00137047f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VPWR_c_813_n 0.342803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_Q_c_909_n 0.0020064f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.555
cc_57 VNB Q 0.0116039f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB Q 0.0038237f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.555
cc_59 VNB Q_N 0.0547467f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.485
cc_60 VNB N_VGND_c_962_n 0.0168478f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_963_n 0.0130264f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_964_n 0.0228469f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_965_n 0.0248337f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_966_n 0.0406978f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_967_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_968_n 0.0202939f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_969_n 0.0537058f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_970_n 0.0446163f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_971_n 0.0217644f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_972_n 0.0194307f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_973_n 0.483602f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_974_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_975_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_976_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VPB N_D_c_143_n 0.0307775f $X=-0.19 $Y=1.66 $X2=0.587 $Y2=1.713
cc_76 VPB N_D_c_148_n 0.0208017f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=1.99
cc_77 VPB D 0.00311708f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_78 VPB N_GATE_c_183_n 0.0147712f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=0.835
cc_79 VPB N_GATE_c_188_n 0.0278544f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=1.99
cc_80 VPB N_A_231_74#_c_234_n 0.0215962f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.385
cc_81 VPB N_A_231_74#_c_235_n 0.0159597f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 VPB N_A_231_74#_c_236_n 0.0440897f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 VPB N_A_231_74#_c_237_n 0.0107407f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_84 VPB N_A_231_74#_M1002_g 0.00162933f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_A_231_74#_c_239_n 0.00638477f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_A_231_74#_c_227_n 0.0121105f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_A_231_74#_c_228_n 0.00629739f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_A_231_74#_c_229_n 0.0345267f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_A_27_413#_c_357_n 0.0387839f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=2.485
cc_90 VPB N_A_27_413#_c_363_n 0.0121024f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.555
cc_91 VPB N_A_27_413#_c_364_n 0.00829651f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_92 VPB N_A_27_413#_c_365_n 0.0185378f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_A_27_413#_c_366_n 0.0078818f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB N_A_27_413#_c_367_n 0.00510726f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_95 VPB N_A_27_413#_c_368_n 0.00355124f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB N_A_27_413#_c_359_n 0.00134076f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_A_27_413#_c_370_n 0.0127813f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_A_27_413#_c_361_n 0.0188032f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB N_A_373_82#_c_458_n 0.0628053f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 VPB N_A_373_82#_c_453_n 0.00203232f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB N_A_373_82#_c_460_n 0.00213586f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_102 VPB N_A_373_82#_c_461_n 0.00298682f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 VPB N_A_373_82#_c_462_n 0.00333779f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB N_A_863_98#_M1018_g 0.00740385f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_105 VPB N_A_863_98#_c_578_n 0.0223095f $X=-0.19 $Y=1.66 $X2=0.587 $Y2=1.385
cc_106 VPB N_A_863_98#_c_579_n 0.0130956f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.385
cc_107 VPB N_A_863_98#_c_580_n 0.0446367f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.385
cc_108 VPB N_A_863_98#_c_581_n 0.0199799f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_109 VPB N_A_863_98#_c_568_n 0.00828604f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_110 VPB N_A_863_98#_c_569_n 0.0197826f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_A_863_98#_c_584_n 0.0255838f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_A_863_98#_c_585_n 0.00710108f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_A_863_98#_c_574_n 0.00339006f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_A_863_98#_c_587_n 0.00863439f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_A_863_98#_c_588_n 0.00297449f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_A_664_392#_c_685_n 0.0302f $X=-0.19 $Y=1.66 $X2=0.587 $Y2=1.385
cc_117 VPB N_A_664_392#_c_692_n 0.00481761f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_A_664_392#_c_687_n 2.13046e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_A_664_392#_c_689_n 0.0126135f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_A_1347_424#_c_775_n 0.0209167f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=2.485
cc_121 VPB N_A_1347_424#_c_771_n 0.00929219f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.555
cc_122 VPB N_A_1347_424#_c_773_n 0.0161066f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_814_n 0.0114238f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_815_n 0.014534f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_816_n 0.0511904f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_817_n 0.00885874f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_818_n 0.00969119f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_819_n 0.0223007f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_820_n 0.0346731f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_821_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_VPWR_c_822_n 0.020445f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_VPWR_c_823_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_824_n 0.0389828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_VPWR_c_825_n 0.019908f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_VPWR_c_813_n 0.129232f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_VPWR_c_827_n 0.0254774f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_VPWR_c_828_n 0.00631927f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_829_n 0.0102767f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_Q_c_912_n 0.0114864f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_140 VPB N_Q_c_913_n 0.0033481f $X=-0.19 $Y=1.66 $X2=0.587 $Y2=1.22
cc_141 VPB N_Q_c_909_n 0.00146455f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.555
cc_142 VPB Q_N 0.0538644f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=2.485
cc_143 N_D_c_143_n N_GATE_c_183_n 0.0189015f $X=0.587 $Y=1.713 $X2=0 $Y2=0
cc_144 D N_GATE_c_183_n 0.00329252f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_145 N_D_c_148_n N_GATE_c_188_n 0.0246328f $X=0.5 $Y=1.99 $X2=0 $Y2=0
cc_146 D GATE 0.0265692f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_147 N_D_c_145_n GATE 3.62319e-19 $X=0.6 $Y=1.385 $X2=0 $Y2=0
cc_148 N_D_c_146_n GATE 2.19319e-19 $X=0.587 $Y=1.22 $X2=0 $Y2=0
cc_149 D N_GATE_c_185_n 0.00202361f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_150 N_D_c_145_n N_GATE_c_185_n 0.0173771f $X=0.6 $Y=1.385 $X2=0 $Y2=0
cc_151 N_D_c_146_n N_GATE_c_186_n 0.0173684f $X=0.587 $Y=1.22 $X2=0 $Y2=0
cc_152 N_D_c_143_n N_A_231_74#_c_239_n 4.43209e-19 $X=0.587 $Y=1.713 $X2=0 $Y2=0
cc_153 N_D_c_148_n N_A_231_74#_c_239_n 0.00169291f $X=0.5 $Y=1.99 $X2=0 $Y2=0
cc_154 D N_A_231_74#_c_227_n 0.014445f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_155 N_D_c_148_n N_A_27_413#_c_363_n 0.00888398f $X=0.5 $Y=1.99 $X2=0 $Y2=0
cc_156 N_D_c_143_n N_A_27_413#_c_364_n 0.00293531f $X=0.587 $Y=1.713 $X2=0 $Y2=0
cc_157 N_D_c_148_n N_A_27_413#_c_364_n 0.0114522f $X=0.5 $Y=1.99 $X2=0 $Y2=0
cc_158 D N_A_27_413#_c_364_n 0.00982509f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_159 N_D_c_148_n N_A_27_413#_c_365_n 0.00508662f $X=0.5 $Y=1.99 $X2=0 $Y2=0
cc_160 D N_A_27_413#_c_360_n 0.00115262f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_161 N_D_c_146_n N_A_27_413#_c_360_n 0.0093194f $X=0.587 $Y=1.22 $X2=0 $Y2=0
cc_162 N_D_c_143_n N_A_27_413#_c_370_n 8.09327e-19 $X=0.587 $Y=1.713 $X2=0 $Y2=0
cc_163 N_D_c_148_n N_A_27_413#_c_370_n 0.00422419f $X=0.5 $Y=1.99 $X2=0 $Y2=0
cc_164 N_D_c_148_n N_A_27_413#_c_361_n 6.75098e-19 $X=0.5 $Y=1.99 $X2=0 $Y2=0
cc_165 D N_A_27_413#_c_361_n 0.0511216f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_166 N_D_c_145_n N_A_27_413#_c_361_n 0.0192748f $X=0.6 $Y=1.385 $X2=0 $Y2=0
cc_167 N_D_c_146_n N_A_27_413#_c_361_n 0.00413599f $X=0.587 $Y=1.22 $X2=0 $Y2=0
cc_168 N_D_c_148_n N_VPWR_c_814_n 0.00358041f $X=0.5 $Y=1.99 $X2=0 $Y2=0
cc_169 N_D_c_148_n N_VPWR_c_813_n 0.00528353f $X=0.5 $Y=1.99 $X2=0 $Y2=0
cc_170 N_D_c_148_n N_VPWR_c_827_n 0.00408232f $X=0.5 $Y=1.99 $X2=0 $Y2=0
cc_171 D N_VGND_c_962_n 0.0153407f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_172 N_D_c_145_n N_VGND_c_962_n 0.00350987f $X=0.6 $Y=1.385 $X2=0 $Y2=0
cc_173 N_D_c_146_n N_VGND_c_962_n 0.00610345f $X=0.587 $Y=1.22 $X2=0 $Y2=0
cc_174 N_D_c_146_n N_VGND_c_968_n 0.0043356f $X=0.587 $Y=1.22 $X2=0 $Y2=0
cc_175 N_D_c_146_n N_VGND_c_973_n 0.00487769f $X=0.587 $Y=1.22 $X2=0 $Y2=0
cc_176 N_GATE_c_183_n N_A_231_74#_c_239_n 2.96086e-19 $X=1.11 $Y=1.9 $X2=0 $Y2=0
cc_177 N_GATE_c_188_n N_A_231_74#_c_239_n 0.0129401f $X=1.11 $Y=1.99 $X2=0 $Y2=0
cc_178 GATE N_A_231_74#_c_225_n 0.0219228f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_179 N_GATE_c_185_n N_A_231_74#_c_225_n 0.00560294f $X=1.17 $Y=1.385 $X2=0
+ $Y2=0
cc_180 N_GATE_c_186_n N_A_231_74#_c_225_n 0.00357954f $X=1.17 $Y=1.22 $X2=0
+ $Y2=0
cc_181 N_GATE_c_183_n N_A_231_74#_c_227_n 0.00850028f $X=1.11 $Y=1.9 $X2=0 $Y2=0
cc_182 GATE N_A_231_74#_c_227_n 0.0205767f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_183 N_GATE_c_185_n N_A_231_74#_c_227_n 0.00166135f $X=1.17 $Y=1.385 $X2=0
+ $Y2=0
cc_184 N_GATE_c_183_n N_A_231_74#_c_229_n 0.00532741f $X=1.11 $Y=1.9 $X2=0 $Y2=0
cc_185 N_GATE_c_185_n N_A_231_74#_c_229_n 0.00282164f $X=1.17 $Y=1.385 $X2=0
+ $Y2=0
cc_186 GATE N_A_231_74#_c_233_n 0.0150231f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_187 N_GATE_c_185_n N_A_231_74#_c_233_n 0.00110094f $X=1.17 $Y=1.385 $X2=0
+ $Y2=0
cc_188 N_GATE_c_186_n N_A_231_74#_c_233_n 0.0081842f $X=1.17 $Y=1.22 $X2=0 $Y2=0
cc_189 N_GATE_c_188_n N_A_27_413#_c_364_n 0.0182894f $X=1.11 $Y=1.99 $X2=0 $Y2=0
cc_190 N_GATE_c_188_n N_A_27_413#_c_365_n 7.56151e-19 $X=1.11 $Y=1.99 $X2=0
+ $Y2=0
cc_191 N_GATE_c_188_n N_A_27_413#_c_366_n 0.00412999f $X=1.11 $Y=1.99 $X2=0
+ $Y2=0
cc_192 N_GATE_c_188_n N_A_27_413#_c_368_n 3.46389e-19 $X=1.11 $Y=1.99 $X2=0
+ $Y2=0
cc_193 N_GATE_c_186_n N_A_27_413#_c_360_n 2.77589e-19 $X=1.17 $Y=1.22 $X2=0
+ $Y2=0
cc_194 N_GATE_c_188_n N_A_27_413#_c_370_n 0.00212662f $X=1.11 $Y=1.99 $X2=0
+ $Y2=0
cc_195 N_GATE_c_188_n N_VPWR_c_814_n 0.00433999f $X=1.11 $Y=1.99 $X2=0 $Y2=0
cc_196 N_GATE_c_188_n N_VPWR_c_824_n 0.0041044f $X=1.11 $Y=1.99 $X2=0 $Y2=0
cc_197 N_GATE_c_188_n N_VPWR_c_813_n 0.00528353f $X=1.11 $Y=1.99 $X2=0 $Y2=0
cc_198 N_GATE_c_186_n N_VGND_c_962_n 0.00984417f $X=1.17 $Y=1.22 $X2=0 $Y2=0
cc_199 N_GATE_c_186_n N_VGND_c_969_n 0.00434272f $X=1.17 $Y=1.22 $X2=0 $Y2=0
cc_200 N_GATE_c_186_n N_VGND_c_973_n 0.00830058f $X=1.17 $Y=1.22 $X2=0 $Y2=0
cc_201 N_A_231_74#_c_234_n N_A_27_413#_c_357_n 0.0244395f $X=2.24 $Y=1.885 $X2=0
+ $Y2=0
cc_202 N_A_231_74#_c_235_n N_A_27_413#_c_357_n 0.0633746f $X=3.245 $Y=1.885
+ $X2=0 $Y2=0
cc_203 N_A_231_74#_c_237_n N_A_27_413#_c_357_n 0.0119882f $X=3.335 $Y=1.765
+ $X2=0 $Y2=0
cc_204 N_A_231_74#_c_228_n N_A_27_413#_c_357_n 0.00127781f $X=2.165 $Y=1.635
+ $X2=0 $Y2=0
cc_205 N_A_231_74#_c_229_n N_A_27_413#_c_357_n 0.0226139f $X=2.165 $Y=1.635
+ $X2=0 $Y2=0
cc_206 N_A_231_74#_M1016_g N_A_27_413#_M1010_g 0.0290125f $X=2.225 $Y=0.78 $X2=0
+ $Y2=0
cc_207 N_A_231_74#_c_226_n N_A_27_413#_M1010_g 0.00947503f $X=2.91 $Y=0.665
+ $X2=0 $Y2=0
cc_208 N_A_231_74#_c_230_n N_A_27_413#_M1010_g 0.0102057f $X=3.08 $Y=0.382 $X2=0
+ $Y2=0
cc_209 N_A_231_74#_c_231_n N_A_27_413#_M1010_g 2.4614e-19 $X=3.91 $Y=0.345 $X2=0
+ $Y2=0
cc_210 N_A_231_74#_M1021_d N_A_27_413#_c_364_n 0.00824855f $X=1.185 $Y=2.065
+ $X2=0 $Y2=0
cc_211 N_A_231_74#_c_239_n N_A_27_413#_c_364_n 0.0153777f $X=1.335 $Y=2.21 $X2=0
+ $Y2=0
cc_212 N_A_231_74#_c_227_n N_A_27_413#_c_364_n 0.00518908f $X=1.675 $Y=1.68
+ $X2=0 $Y2=0
cc_213 N_A_231_74#_c_234_n N_A_27_413#_c_366_n 0.00476969f $X=2.24 $Y=1.885
+ $X2=0 $Y2=0
cc_214 N_A_231_74#_c_239_n N_A_27_413#_c_366_n 0.0110004f $X=1.335 $Y=2.21 $X2=0
+ $Y2=0
cc_215 N_A_231_74#_c_234_n N_A_27_413#_c_367_n 0.013393f $X=2.24 $Y=1.885 $X2=0
+ $Y2=0
cc_216 N_A_231_74#_c_228_n N_A_27_413#_c_367_n 0.0418056f $X=2.165 $Y=1.635
+ $X2=0 $Y2=0
cc_217 N_A_231_74#_c_229_n N_A_27_413#_c_367_n 0.00209357f $X=2.165 $Y=1.635
+ $X2=0 $Y2=0
cc_218 N_A_231_74#_c_239_n N_A_27_413#_c_368_n 0.0145075f $X=1.335 $Y=2.21 $X2=0
+ $Y2=0
cc_219 N_A_231_74#_c_227_n N_A_27_413#_c_368_n 0.00794178f $X=1.675 $Y=1.68
+ $X2=0 $Y2=0
cc_220 N_A_231_74#_c_228_n N_A_27_413#_c_368_n 0.00758469f $X=2.165 $Y=1.635
+ $X2=0 $Y2=0
cc_221 N_A_231_74#_c_229_n N_A_27_413#_c_368_n 6.3956e-19 $X=2.165 $Y=1.635
+ $X2=0 $Y2=0
cc_222 N_A_231_74#_c_234_n N_A_27_413#_c_359_n 0.00401056f $X=2.24 $Y=1.885
+ $X2=0 $Y2=0
cc_223 N_A_231_74#_c_228_n N_A_27_413#_c_359_n 0.0280182f $X=2.165 $Y=1.635
+ $X2=0 $Y2=0
cc_224 N_A_231_74#_c_229_n N_A_27_413#_c_359_n 7.60564e-19 $X=2.165 $Y=1.635
+ $X2=0 $Y2=0
cc_225 N_A_231_74#_c_226_n N_A_373_82#_M1016_s 0.00711247f $X=2.91 $Y=0.665
+ $X2=-0.19 $Y2=-0.245
cc_226 N_A_231_74#_c_235_n N_A_373_82#_c_458_n 0.0315019f $X=3.245 $Y=1.885
+ $X2=0 $Y2=0
cc_227 N_A_231_74#_c_236_n N_A_373_82#_c_458_n 0.0247276f $X=3.925 $Y=1.765
+ $X2=0 $Y2=0
cc_228 N_A_231_74#_M1016_g N_A_373_82#_c_452_n 0.00987474f $X=2.225 $Y=0.78
+ $X2=0 $Y2=0
cc_229 N_A_231_74#_c_226_n N_A_373_82#_c_452_n 0.0309272f $X=2.91 $Y=0.665 $X2=0
+ $Y2=0
cc_230 N_A_231_74#_c_228_n N_A_373_82#_c_452_n 0.00769137f $X=2.165 $Y=1.635
+ $X2=0 $Y2=0
cc_231 N_A_231_74#_c_229_n N_A_373_82#_c_452_n 6.90333e-19 $X=2.165 $Y=1.635
+ $X2=0 $Y2=0
cc_232 N_A_231_74#_c_230_n N_A_373_82#_c_452_n 0.0041614f $X=3.08 $Y=0.382 $X2=0
+ $Y2=0
cc_233 N_A_231_74#_c_234_n N_A_373_82#_c_471_n 0.0105718f $X=2.24 $Y=1.885 $X2=0
+ $Y2=0
cc_234 N_A_231_74#_c_235_n N_A_373_82#_c_453_n 0.0110894f $X=3.245 $Y=1.885
+ $X2=0 $Y2=0
cc_235 N_A_231_74#_c_237_n N_A_373_82#_c_453_n 0.00574342f $X=3.335 $Y=1.765
+ $X2=0 $Y2=0
cc_236 N_A_231_74#_c_235_n N_A_373_82#_c_460_n 0.0112302f $X=3.245 $Y=1.885
+ $X2=0 $Y2=0
cc_237 N_A_231_74#_c_236_n N_A_373_82#_c_460_n 0.00313621f $X=3.925 $Y=1.765
+ $X2=0 $Y2=0
cc_238 N_A_231_74#_c_235_n N_A_373_82#_c_461_n 5.46839e-19 $X=3.245 $Y=1.885
+ $X2=0 $Y2=0
cc_239 N_A_231_74#_c_236_n N_A_373_82#_c_461_n 0.00108254f $X=3.925 $Y=1.765
+ $X2=0 $Y2=0
cc_240 N_A_231_74#_M1016_g N_A_373_82#_c_454_n 0.00460645f $X=2.225 $Y=0.78
+ $X2=0 $Y2=0
cc_241 N_A_231_74#_c_226_n N_A_373_82#_c_454_n 0.0203885f $X=2.91 $Y=0.665 $X2=0
+ $Y2=0
cc_242 N_A_231_74#_c_228_n N_A_373_82#_c_454_n 0.0178644f $X=2.165 $Y=1.635
+ $X2=0 $Y2=0
cc_243 N_A_231_74#_c_229_n N_A_373_82#_c_454_n 0.00640006f $X=2.165 $Y=1.635
+ $X2=0 $Y2=0
cc_244 N_A_231_74#_c_233_n N_A_373_82#_c_454_n 0.0220228f $X=1.295 $Y=0.52 $X2=0
+ $Y2=0
cc_245 N_A_231_74#_c_234_n N_A_373_82#_c_462_n 0.00635803f $X=2.24 $Y=1.885
+ $X2=0 $Y2=0
cc_246 N_A_231_74#_c_237_n N_A_373_82#_c_455_n 0.00123761f $X=3.335 $Y=1.765
+ $X2=0 $Y2=0
cc_247 N_A_231_74#_M1002_g N_A_373_82#_c_455_n 8.02895e-19 $X=4 $Y=0.83 $X2=0
+ $Y2=0
cc_248 N_A_231_74#_c_230_n N_A_373_82#_c_455_n 0.00206098f $X=3.08 $Y=0.382
+ $X2=0 $Y2=0
cc_249 N_A_231_74#_c_231_n N_A_373_82#_c_455_n 0.00566193f $X=3.91 $Y=0.345
+ $X2=0 $Y2=0
cc_250 N_A_231_74#_c_237_n N_A_373_82#_c_456_n 0.0212694f $X=3.335 $Y=1.765
+ $X2=0 $Y2=0
cc_251 N_A_231_74#_M1002_g N_A_373_82#_c_456_n 0.00843671f $X=4 $Y=0.83 $X2=0
+ $Y2=0
cc_252 N_A_231_74#_c_235_n N_A_373_82#_c_490_n 0.00351296f $X=3.245 $Y=1.885
+ $X2=0 $Y2=0
cc_253 N_A_231_74#_M1002_g N_A_373_82#_c_457_n 0.0109435f $X=4 $Y=0.83 $X2=0
+ $Y2=0
cc_254 N_A_231_74#_c_230_n N_A_373_82#_c_457_n 0.00451102f $X=3.08 $Y=0.382
+ $X2=0 $Y2=0
cc_255 N_A_231_74#_c_231_n N_A_373_82#_c_457_n 0.0139998f $X=3.91 $Y=0.345 $X2=0
+ $Y2=0
cc_256 N_A_231_74#_c_232_n N_A_373_82#_c_457_n 0.00643136f $X=3.91 $Y=0.345
+ $X2=0 $Y2=0
cc_257 N_A_231_74#_c_232_n N_A_863_98#_M1018_g 0.0350251f $X=3.91 $Y=0.345 $X2=0
+ $Y2=0
cc_258 N_A_231_74#_M1002_g N_A_863_98#_c_578_n 0.0350251f $X=4 $Y=0.83 $X2=0
+ $Y2=0
cc_259 N_A_231_74#_c_231_n N_A_664_392#_M1009_d 0.00228312f $X=3.91 $Y=0.345
+ $X2=-0.19 $Y2=-0.245
cc_260 N_A_231_74#_M1002_g N_A_664_392#_c_696_n 0.00664769f $X=4 $Y=0.83 $X2=0
+ $Y2=0
cc_261 N_A_231_74#_c_230_n N_A_664_392#_c_696_n 0.00426955f $X=3.08 $Y=0.382
+ $X2=0 $Y2=0
cc_262 N_A_231_74#_c_231_n N_A_664_392#_c_696_n 0.0403154f $X=3.91 $Y=0.345
+ $X2=0 $Y2=0
cc_263 N_A_231_74#_c_232_n N_A_664_392#_c_696_n 0.00398671f $X=3.91 $Y=0.345
+ $X2=0 $Y2=0
cc_264 N_A_231_74#_c_235_n N_A_664_392#_c_692_n 0.00244936f $X=3.245 $Y=1.885
+ $X2=0 $Y2=0
cc_265 N_A_231_74#_c_236_n N_A_664_392#_c_692_n 0.00501013f $X=3.925 $Y=1.765
+ $X2=0 $Y2=0
cc_266 N_A_231_74#_c_237_n N_A_664_392#_c_692_n 0.00102991f $X=3.335 $Y=1.765
+ $X2=0 $Y2=0
cc_267 N_A_231_74#_c_236_n N_A_664_392#_c_686_n 0.0092899f $X=3.925 $Y=1.765
+ $X2=0 $Y2=0
cc_268 N_A_231_74#_c_236_n N_A_664_392#_c_687_n 0.004769f $X=3.925 $Y=1.765
+ $X2=0 $Y2=0
cc_269 N_A_231_74#_M1002_g N_A_664_392#_c_688_n 0.0235251f $X=4 $Y=0.83 $X2=0
+ $Y2=0
cc_270 N_A_231_74#_c_236_n N_A_664_392#_c_689_n 0.00361813f $X=3.925 $Y=1.765
+ $X2=0 $Y2=0
cc_271 N_A_231_74#_M1002_g N_A_664_392#_c_689_n 0.00631498f $X=4 $Y=0.83 $X2=0
+ $Y2=0
cc_272 N_A_231_74#_c_236_n N_A_664_392#_c_708_n 0.00657304f $X=3.925 $Y=1.765
+ $X2=0 $Y2=0
cc_273 N_A_231_74#_M1002_g N_A_664_392#_c_708_n 9.83002e-19 $X=4 $Y=0.83 $X2=0
+ $Y2=0
cc_274 N_A_231_74#_c_234_n N_VPWR_c_815_n 0.00358937f $X=2.24 $Y=1.885 $X2=0
+ $Y2=0
cc_275 N_A_231_74#_c_235_n N_VPWR_c_816_n 0.00335042f $X=3.245 $Y=1.885 $X2=0
+ $Y2=0
cc_276 N_A_231_74#_c_234_n N_VPWR_c_824_n 0.00366035f $X=2.24 $Y=1.885 $X2=0
+ $Y2=0
cc_277 N_A_231_74#_c_234_n N_VPWR_c_813_n 0.0049649f $X=2.24 $Y=1.885 $X2=0
+ $Y2=0
cc_278 N_A_231_74#_c_235_n N_VPWR_c_813_n 0.00435185f $X=3.245 $Y=1.885 $X2=0
+ $Y2=0
cc_279 N_A_231_74#_c_226_n N_VGND_M1016_d 0.0101073f $X=2.91 $Y=0.665 $X2=0
+ $Y2=0
cc_280 N_A_231_74#_c_233_n N_VGND_c_962_n 0.0275297f $X=1.295 $Y=0.52 $X2=0
+ $Y2=0
cc_281 N_A_231_74#_c_231_n N_VGND_c_963_n 0.0102942f $X=3.91 $Y=0.345 $X2=0
+ $Y2=0
cc_282 N_A_231_74#_c_232_n N_VGND_c_963_n 0.00296924f $X=3.91 $Y=0.345 $X2=0
+ $Y2=0
cc_283 N_A_231_74#_M1016_g N_VGND_c_969_n 0.00811784f $X=2.225 $Y=0.78 $X2=0
+ $Y2=0
cc_284 N_A_231_74#_c_226_n N_VGND_c_969_n 0.041047f $X=2.91 $Y=0.665 $X2=0 $Y2=0
cc_285 N_A_231_74#_c_230_n N_VGND_c_969_n 0.0114424f $X=3.08 $Y=0.382 $X2=0
+ $Y2=0
cc_286 N_A_231_74#_c_233_n N_VGND_c_969_n 0.0241214f $X=1.295 $Y=0.52 $X2=0
+ $Y2=0
cc_287 N_A_231_74#_c_226_n N_VGND_c_970_n 0.00276577f $X=2.91 $Y=0.665 $X2=0
+ $Y2=0
cc_288 N_A_231_74#_c_230_n N_VGND_c_970_n 0.0117598f $X=3.08 $Y=0.382 $X2=0
+ $Y2=0
cc_289 N_A_231_74#_c_231_n N_VGND_c_970_n 0.0649228f $X=3.91 $Y=0.345 $X2=0
+ $Y2=0
cc_290 N_A_231_74#_c_232_n N_VGND_c_970_n 0.00653686f $X=3.91 $Y=0.345 $X2=0
+ $Y2=0
cc_291 N_A_231_74#_M1016_g N_VGND_c_973_n 0.00533081f $X=2.225 $Y=0.78 $X2=0
+ $Y2=0
cc_292 N_A_231_74#_c_226_n N_VGND_c_973_n 0.0270618f $X=2.91 $Y=0.665 $X2=0
+ $Y2=0
cc_293 N_A_231_74#_c_230_n N_VGND_c_973_n 0.00647831f $X=3.08 $Y=0.382 $X2=0
+ $Y2=0
cc_294 N_A_231_74#_c_231_n N_VGND_c_973_n 0.0362374f $X=3.91 $Y=0.345 $X2=0
+ $Y2=0
cc_295 N_A_231_74#_c_232_n N_VGND_c_973_n 0.0102677f $X=3.91 $Y=0.345 $X2=0
+ $Y2=0
cc_296 N_A_231_74#_c_233_n N_VGND_c_973_n 0.019925f $X=1.295 $Y=0.52 $X2=0 $Y2=0
cc_297 N_A_231_74#_c_230_n A_589_80# 0.00384904f $X=3.08 $Y=0.382 $X2=-0.19
+ $Y2=-0.245
cc_298 N_A_231_74#_c_231_n A_589_80# 0.0011484f $X=3.91 $Y=0.345 $X2=-0.19
+ $Y2=-0.245
cc_299 N_A_27_413#_c_367_n N_A_373_82#_M1014_s 0.00733516f $X=2.545 $Y=2.145
+ $X2=0 $Y2=0
cc_300 N_A_27_413#_c_357_n N_A_373_82#_c_452_n 0.00157896f $X=2.855 $Y=1.885
+ $X2=0 $Y2=0
cc_301 N_A_27_413#_M1010_g N_A_373_82#_c_452_n 0.0133358f $X=2.87 $Y=0.72 $X2=0
+ $Y2=0
cc_302 N_A_27_413#_c_359_n N_A_373_82#_c_452_n 0.0176986f $X=2.71 $Y=1.635 $X2=0
+ $Y2=0
cc_303 N_A_27_413#_c_357_n N_A_373_82#_c_471_n 0.0150034f $X=2.855 $Y=1.885
+ $X2=0 $Y2=0
cc_304 N_A_27_413#_c_367_n N_A_373_82#_c_471_n 0.0368491f $X=2.545 $Y=2.145
+ $X2=0 $Y2=0
cc_305 N_A_27_413#_c_357_n N_A_373_82#_c_453_n 0.0135537f $X=2.855 $Y=1.885
+ $X2=0 $Y2=0
cc_306 N_A_27_413#_c_367_n N_A_373_82#_c_453_n 0.0133618f $X=2.545 $Y=2.145
+ $X2=0 $Y2=0
cc_307 N_A_27_413#_M1010_g N_A_373_82#_c_454_n 5.18311e-19 $X=2.87 $Y=0.72 $X2=0
+ $Y2=0
cc_308 N_A_27_413#_c_357_n N_A_373_82#_c_462_n 0.00101548f $X=2.855 $Y=1.885
+ $X2=0 $Y2=0
cc_309 N_A_27_413#_c_364_n N_A_373_82#_c_462_n 0.0145003f $X=1.59 $Y=2.63 $X2=0
+ $Y2=0
cc_310 N_A_27_413#_c_366_n N_A_373_82#_c_462_n 0.0110004f $X=1.675 $Y=2.545
+ $X2=0 $Y2=0
cc_311 N_A_27_413#_c_367_n N_A_373_82#_c_462_n 0.0148773f $X=2.545 $Y=2.145
+ $X2=0 $Y2=0
cc_312 N_A_27_413#_M1010_g N_A_373_82#_c_455_n 0.00727424f $X=2.87 $Y=0.72 $X2=0
+ $Y2=0
cc_313 N_A_27_413#_c_359_n N_A_373_82#_c_455_n 0.0441572f $X=2.71 $Y=1.635 $X2=0
+ $Y2=0
cc_314 N_A_27_413#_c_357_n N_A_373_82#_c_456_n 0.0318813f $X=2.855 $Y=1.885
+ $X2=0 $Y2=0
cc_315 N_A_27_413#_M1010_g N_A_373_82#_c_457_n 0.0318813f $X=2.87 $Y=0.72 $X2=0
+ $Y2=0
cc_316 N_A_27_413#_M1010_g N_A_664_392#_c_696_n 5.45644e-19 $X=2.87 $Y=0.72
+ $X2=0 $Y2=0
cc_317 N_A_27_413#_c_364_n N_VPWR_M1017_d 0.0138739f $X=1.59 $Y=2.63 $X2=-0.19
+ $Y2=-0.245
cc_318 N_A_27_413#_c_367_n N_VPWR_M1014_d 0.0116894f $X=2.545 $Y=2.145 $X2=0
+ $Y2=0
cc_319 N_A_27_413#_c_359_n N_VPWR_M1014_d 0.00147061f $X=2.71 $Y=1.635 $X2=0
+ $Y2=0
cc_320 N_A_27_413#_c_364_n N_VPWR_c_814_n 0.024844f $X=1.59 $Y=2.63 $X2=0 $Y2=0
cc_321 N_A_27_413#_c_365_n N_VPWR_c_814_n 0.00279174f $X=0.44 $Y=2.63 $X2=0
+ $Y2=0
cc_322 N_A_27_413#_c_357_n N_VPWR_c_815_n 0.0109005f $X=2.855 $Y=1.885 $X2=0
+ $Y2=0
cc_323 N_A_27_413#_c_357_n N_VPWR_c_816_n 0.00335072f $X=2.855 $Y=1.885 $X2=0
+ $Y2=0
cc_324 N_A_27_413#_c_364_n N_VPWR_c_824_n 0.0138915f $X=1.59 $Y=2.63 $X2=0 $Y2=0
cc_325 N_A_27_413#_c_357_n N_VPWR_c_813_n 0.00438657f $X=2.855 $Y=1.885 $X2=0
+ $Y2=0
cc_326 N_A_27_413#_c_364_n N_VPWR_c_813_n 0.0303192f $X=1.59 $Y=2.63 $X2=0 $Y2=0
cc_327 N_A_27_413#_c_365_n N_VPWR_c_813_n 0.01229f $X=0.44 $Y=2.63 $X2=0 $Y2=0
cc_328 N_A_27_413#_c_364_n N_VPWR_c_827_n 0.00302772f $X=1.59 $Y=2.63 $X2=0
+ $Y2=0
cc_329 N_A_27_413#_c_365_n N_VPWR_c_827_n 0.0125402f $X=0.44 $Y=2.63 $X2=0 $Y2=0
cc_330 N_A_27_413#_c_360_n N_VGND_c_962_n 0.017794f $X=0.285 $Y=0.795 $X2=0
+ $Y2=0
cc_331 N_A_27_413#_c_360_n N_VGND_c_968_n 0.00868052f $X=0.285 $Y=0.795 $X2=0
+ $Y2=0
cc_332 N_A_27_413#_M1010_g N_VGND_c_969_n 0.00150827f $X=2.87 $Y=0.72 $X2=0
+ $Y2=0
cc_333 N_A_27_413#_M1010_g N_VGND_c_970_n 0.00347067f $X=2.87 $Y=0.72 $X2=0
+ $Y2=0
cc_334 N_A_27_413#_M1010_g N_VGND_c_973_n 0.00414706f $X=2.87 $Y=0.72 $X2=0
+ $Y2=0
cc_335 N_A_27_413#_c_360_n N_VGND_c_973_n 0.0113795f $X=0.285 $Y=0.795 $X2=0
+ $Y2=0
cc_336 N_A_373_82#_c_458_n N_A_863_98#_c_579_n 0.0167612f $X=3.775 $Y=2.465
+ $X2=0 $Y2=0
cc_337 N_A_373_82#_c_461_n N_A_863_98#_c_579_n 3.40059e-19 $X=3.935 $Y=2.215
+ $X2=0 $Y2=0
cc_338 N_A_373_82#_c_458_n N_A_863_98#_c_580_n 0.0195728f $X=3.775 $Y=2.465
+ $X2=0 $Y2=0
cc_339 N_A_373_82#_c_460_n N_A_863_98#_c_580_n 0.00348668f $X=3.77 $Y=2.525
+ $X2=0 $Y2=0
cc_340 N_A_373_82#_c_461_n N_A_863_98#_c_580_n 0.00178992f $X=3.935 $Y=2.215
+ $X2=0 $Y2=0
cc_341 N_A_373_82#_c_458_n N_A_863_98#_c_585_n 9.85724e-19 $X=3.775 $Y=2.465
+ $X2=0 $Y2=0
cc_342 N_A_373_82#_c_461_n N_A_863_98#_c_585_n 0.0177431f $X=3.935 $Y=2.215
+ $X2=0 $Y2=0
cc_343 N_A_373_82#_c_455_n N_A_664_392#_M1009_d 0.00156514f $X=3.28 $Y=1.105
+ $X2=-0.19 $Y2=-0.245
cc_344 N_A_373_82#_c_460_n N_A_664_392#_M1000_d 0.00786329f $X=3.77 $Y=2.525
+ $X2=0 $Y2=0
cc_345 N_A_373_82#_c_455_n N_A_664_392#_c_696_n 0.0114609f $X=3.28 $Y=1.105
+ $X2=0 $Y2=0
cc_346 N_A_373_82#_c_456_n N_A_664_392#_c_696_n 8.1443e-19 $X=3.35 $Y=1.315
+ $X2=0 $Y2=0
cc_347 N_A_373_82#_c_457_n N_A_664_392#_c_696_n 0.00657958f $X=3.35 $Y=1.15
+ $X2=0 $Y2=0
cc_348 N_A_373_82#_c_458_n N_A_664_392#_c_692_n 0.00191279f $X=3.775 $Y=2.465
+ $X2=0 $Y2=0
cc_349 N_A_373_82#_c_453_n N_A_664_392#_c_692_n 0.0316328f $X=3.13 $Y=2.44 $X2=0
+ $Y2=0
cc_350 N_A_373_82#_c_460_n N_A_664_392#_c_692_n 0.0135656f $X=3.77 $Y=2.525
+ $X2=0 $Y2=0
cc_351 N_A_373_82#_c_461_n N_A_664_392#_c_692_n 0.0135564f $X=3.935 $Y=2.215
+ $X2=0 $Y2=0
cc_352 N_A_373_82#_c_458_n N_A_664_392#_c_686_n 4.19696e-19 $X=3.775 $Y=2.465
+ $X2=0 $Y2=0
cc_353 N_A_373_82#_c_460_n N_A_664_392#_c_686_n 0.00535267f $X=3.77 $Y=2.525
+ $X2=0 $Y2=0
cc_354 N_A_373_82#_c_461_n N_A_664_392#_c_686_n 5.02386e-19 $X=3.935 $Y=2.215
+ $X2=0 $Y2=0
cc_355 N_A_373_82#_c_453_n N_A_664_392#_c_687_n 0.0132811f $X=3.13 $Y=2.44 $X2=0
+ $Y2=0
cc_356 N_A_373_82#_c_455_n N_A_664_392#_c_687_n 0.011103f $X=3.28 $Y=1.105 $X2=0
+ $Y2=0
cc_357 N_A_373_82#_c_456_n N_A_664_392#_c_687_n 4.7393e-19 $X=3.35 $Y=1.315
+ $X2=0 $Y2=0
cc_358 N_A_373_82#_c_453_n N_A_664_392#_c_688_n 0.00553075f $X=3.13 $Y=2.44
+ $X2=0 $Y2=0
cc_359 N_A_373_82#_c_455_n N_A_664_392#_c_688_n 0.0260074f $X=3.28 $Y=1.105
+ $X2=0 $Y2=0
cc_360 N_A_373_82#_c_456_n N_A_664_392#_c_688_n 0.0024439f $X=3.35 $Y=1.315
+ $X2=0 $Y2=0
cc_361 N_A_373_82#_c_457_n N_A_664_392#_c_688_n 0.00321011f $X=3.35 $Y=1.15
+ $X2=0 $Y2=0
cc_362 N_A_373_82#_c_458_n N_A_664_392#_c_689_n 3.12388e-19 $X=3.775 $Y=2.465
+ $X2=0 $Y2=0
cc_363 N_A_373_82#_c_461_n N_A_664_392#_c_689_n 0.00882513f $X=3.935 $Y=2.215
+ $X2=0 $Y2=0
cc_364 N_A_373_82#_c_458_n N_A_664_392#_c_708_n 2.0477e-19 $X=3.775 $Y=2.465
+ $X2=0 $Y2=0
cc_365 N_A_373_82#_c_461_n N_A_664_392#_c_708_n 0.0110761f $X=3.935 $Y=2.215
+ $X2=0 $Y2=0
cc_366 N_A_373_82#_c_471_n N_VPWR_M1014_d 0.00868895f $X=3.045 $Y=2.525 $X2=0
+ $Y2=0
cc_367 N_A_373_82#_c_471_n N_VPWR_c_815_n 0.0256243f $X=3.045 $Y=2.525 $X2=0
+ $Y2=0
cc_368 N_A_373_82#_c_462_n N_VPWR_c_815_n 0.0027161f $X=2.055 $Y=2.525 $X2=0
+ $Y2=0
cc_369 N_A_373_82#_c_458_n N_VPWR_c_816_n 0.00335018f $X=3.775 $Y=2.465 $X2=0
+ $Y2=0
cc_370 N_A_373_82#_c_471_n N_VPWR_c_816_n 0.00394293f $X=3.045 $Y=2.525 $X2=0
+ $Y2=0
cc_371 N_A_373_82#_c_460_n N_VPWR_c_816_n 0.01183f $X=3.77 $Y=2.525 $X2=0 $Y2=0
cc_372 N_A_373_82#_c_490_n N_VPWR_c_816_n 0.0022032f $X=3.13 $Y=2.525 $X2=0
+ $Y2=0
cc_373 N_A_373_82#_c_458_n N_VPWR_c_817_n 0.00210477f $X=3.775 $Y=2.465 $X2=0
+ $Y2=0
cc_374 N_A_373_82#_c_460_n N_VPWR_c_817_n 0.00293123f $X=3.77 $Y=2.525 $X2=0
+ $Y2=0
cc_375 N_A_373_82#_c_471_n N_VPWR_c_824_n 0.00237993f $X=3.045 $Y=2.525 $X2=0
+ $Y2=0
cc_376 N_A_373_82#_c_462_n N_VPWR_c_824_n 0.0064234f $X=2.055 $Y=2.525 $X2=0
+ $Y2=0
cc_377 N_A_373_82#_c_458_n N_VPWR_c_813_n 0.00437239f $X=3.775 $Y=2.465 $X2=0
+ $Y2=0
cc_378 N_A_373_82#_c_471_n N_VPWR_c_813_n 0.0147491f $X=3.045 $Y=2.525 $X2=0
+ $Y2=0
cc_379 N_A_373_82#_c_460_n N_VPWR_c_813_n 0.0228673f $X=3.77 $Y=2.525 $X2=0
+ $Y2=0
cc_380 N_A_373_82#_c_462_n N_VPWR_c_813_n 0.00806222f $X=2.055 $Y=2.525 $X2=0
+ $Y2=0
cc_381 N_A_373_82#_c_490_n N_VPWR_c_813_n 0.00459893f $X=3.13 $Y=2.525 $X2=0
+ $Y2=0
cc_382 N_A_373_82#_c_471_n A_586_392# 0.0032623f $X=3.045 $Y=2.525 $X2=-0.19
+ $Y2=-0.245
cc_383 N_A_373_82#_c_453_n A_586_392# 0.0045678f $X=3.13 $Y=2.44 $X2=-0.19
+ $Y2=-0.245
cc_384 N_A_373_82#_c_490_n A_586_392# 0.00134166f $X=3.13 $Y=2.525 $X2=-0.19
+ $Y2=-0.245
cc_385 N_A_373_82#_c_460_n A_770_508# 0.00487517f $X=3.77 $Y=2.525 $X2=-0.19
+ $Y2=-0.245
cc_386 N_A_373_82#_c_452_n N_VGND_M1016_d 0.00557246f $X=3.045 $Y=1.105 $X2=0
+ $Y2=0
cc_387 N_A_373_82#_c_457_n N_VGND_c_970_n 9.29978e-19 $X=3.35 $Y=1.15 $X2=0
+ $Y2=0
cc_388 N_A_373_82#_c_452_n A_589_80# 6.09291e-19 $X=3.045 $Y=1.105 $X2=-0.19
+ $Y2=-0.245
cc_389 N_A_373_82#_c_455_n A_589_80# 0.00141443f $X=3.28 $Y=1.105 $X2=-0.19
+ $Y2=-0.245
cc_390 N_A_863_98#_M1018_g N_A_664_392#_M1006_g 0.0165523f $X=4.39 $Y=0.83 $X2=0
+ $Y2=0
cc_391 N_A_863_98#_c_572_n N_A_664_392#_M1006_g 0.00627138f $X=5.185 $Y=0.515
+ $X2=0 $Y2=0
cc_392 N_A_863_98#_c_573_n N_A_664_392#_M1006_g 0.00716244f $X=5.29 $Y=1.32
+ $X2=0 $Y2=0
cc_393 N_A_863_98#_c_575_n N_A_664_392#_M1006_g 0.00261068f $X=5.197 $Y=1.07
+ $X2=0 $Y2=0
cc_394 N_A_863_98#_M1018_g N_A_664_392#_c_685_n 0.0217295f $X=4.39 $Y=0.83 $X2=0
+ $Y2=0
cc_395 N_A_863_98#_c_578_n N_A_664_392#_c_685_n 0.0139039f $X=4.48 $Y=1.975
+ $X2=0 $Y2=0
cc_396 N_A_863_98#_c_580_n N_A_664_392#_c_685_n 0.0128465f $X=4.43 $Y=2.465
+ $X2=0 $Y2=0
cc_397 N_A_863_98#_c_571_n N_A_664_392#_c_685_n 0.0176287f $X=6.065 $Y=1.485
+ $X2=0 $Y2=0
cc_398 N_A_863_98#_c_585_n N_A_664_392#_c_685_n 0.0232029f $X=5.205 $Y=2.155
+ $X2=0 $Y2=0
cc_399 N_A_863_98#_c_574_n N_A_664_392#_c_685_n 0.00947816f $X=5.37 $Y=1.985
+ $X2=0 $Y2=0
cc_400 N_A_863_98#_c_587_n N_A_664_392#_c_685_n 0.0118819f $X=5.37 $Y=2.815
+ $X2=0 $Y2=0
cc_401 N_A_863_98#_c_575_n N_A_664_392#_c_685_n 0.0051475f $X=5.197 $Y=1.07
+ $X2=0 $Y2=0
cc_402 N_A_863_98#_c_576_n N_A_664_392#_c_685_n 0.00700952f $X=5.61 $Y=1.485
+ $X2=0 $Y2=0
cc_403 N_A_863_98#_c_588_n N_A_664_392#_c_685_n 9.46256e-19 $X=5.37 $Y=2.155
+ $X2=0 $Y2=0
cc_404 N_A_863_98#_M1018_g N_A_664_392#_c_696_n 4.97999e-19 $X=4.39 $Y=0.83
+ $X2=0 $Y2=0
cc_405 N_A_863_98#_M1018_g N_A_664_392#_c_688_n 0.00357066f $X=4.39 $Y=0.83
+ $X2=0 $Y2=0
cc_406 N_A_863_98#_M1018_g N_A_664_392#_c_689_n 0.0134413f $X=4.39 $Y=0.83 $X2=0
+ $Y2=0
cc_407 N_A_863_98#_c_578_n N_A_664_392#_c_689_n 0.00818075f $X=4.48 $Y=1.975
+ $X2=0 $Y2=0
cc_408 N_A_863_98#_c_585_n N_A_664_392#_c_689_n 0.0558787f $X=5.205 $Y=2.155
+ $X2=0 $Y2=0
cc_409 N_A_863_98#_c_574_n N_A_664_392#_c_689_n 0.0142966f $X=5.37 $Y=1.985
+ $X2=0 $Y2=0
cc_410 N_A_863_98#_M1018_g N_A_664_392#_c_690_n 0.00406012f $X=4.39 $Y=0.83
+ $X2=0 $Y2=0
cc_411 N_A_863_98#_c_573_n N_A_664_392#_c_690_n 0.00601245f $X=5.29 $Y=1.32
+ $X2=0 $Y2=0
cc_412 N_A_863_98#_c_575_n N_A_664_392#_c_690_n 0.00109211f $X=5.197 $Y=1.07
+ $X2=0 $Y2=0
cc_413 N_A_863_98#_c_576_n N_A_664_392#_c_690_n 0.0265744f $X=5.61 $Y=1.485
+ $X2=0 $Y2=0
cc_414 N_A_863_98#_c_568_n N_A_1347_424#_c_770_n 0.0183347f $X=6.66 $Y=1.65
+ $X2=0 $Y2=0
cc_415 N_A_863_98#_M1013_g N_A_1347_424#_c_772_n 6.67726e-19 $X=6.175 $Y=0.76
+ $X2=0 $Y2=0
cc_416 N_A_863_98#_M1015_g N_A_1347_424#_c_772_n 0.017438f $X=6.675 $Y=0.855
+ $X2=0 $Y2=0
cc_417 N_A_863_98#_c_581_n N_A_1347_424#_c_773_n 0.00111647f $X=6.155 $Y=1.765
+ $X2=0 $Y2=0
cc_418 N_A_863_98#_c_568_n N_A_1347_424#_c_773_n 4.36622e-19 $X=6.66 $Y=1.65
+ $X2=0 $Y2=0
cc_419 N_A_863_98#_c_569_n N_A_1347_424#_c_773_n 0.0121493f $X=6.66 $Y=1.955
+ $X2=0 $Y2=0
cc_420 N_A_863_98#_c_584_n N_A_1347_424#_c_773_n 0.0187565f $X=6.66 $Y=2.045
+ $X2=0 $Y2=0
cc_421 N_A_863_98#_c_568_n N_A_1347_424#_c_774_n 0.013973f $X=6.66 $Y=1.65 $X2=0
+ $Y2=0
cc_422 N_A_863_98#_c_585_n N_VPWR_M1007_d 0.0056852f $X=5.205 $Y=2.155 $X2=0
+ $Y2=0
cc_423 N_A_863_98#_c_580_n N_VPWR_c_816_n 0.00413917f $X=4.43 $Y=2.465 $X2=0
+ $Y2=0
cc_424 N_A_863_98#_c_580_n N_VPWR_c_817_n 0.0249383f $X=4.43 $Y=2.465 $X2=0
+ $Y2=0
cc_425 N_A_863_98#_c_585_n N_VPWR_c_817_n 0.0338401f $X=5.205 $Y=2.155 $X2=0
+ $Y2=0
cc_426 N_A_863_98#_c_587_n N_VPWR_c_817_n 0.017175f $X=5.37 $Y=2.815 $X2=0 $Y2=0
cc_427 N_A_863_98#_c_581_n N_VPWR_c_818_n 0.00639895f $X=6.155 $Y=1.765 $X2=0
+ $Y2=0
cc_428 N_A_863_98#_c_568_n N_VPWR_c_818_n 0.00843419f $X=6.66 $Y=1.65 $X2=0
+ $Y2=0
cc_429 N_A_863_98#_c_584_n N_VPWR_c_818_n 0.00777948f $X=6.66 $Y=2.045 $X2=0
+ $Y2=0
cc_430 N_A_863_98#_c_569_n N_VPWR_c_819_n 8.61266e-19 $X=6.66 $Y=1.955 $X2=0
+ $Y2=0
cc_431 N_A_863_98#_c_584_n N_VPWR_c_819_n 0.00466055f $X=6.66 $Y=2.045 $X2=0
+ $Y2=0
cc_432 N_A_863_98#_c_581_n N_VPWR_c_820_n 0.00411612f $X=6.155 $Y=1.765 $X2=0
+ $Y2=0
cc_433 N_A_863_98#_c_587_n N_VPWR_c_820_n 0.0145938f $X=5.37 $Y=2.815 $X2=0
+ $Y2=0
cc_434 N_A_863_98#_c_584_n N_VPWR_c_822_n 0.00445602f $X=6.66 $Y=2.045 $X2=0
+ $Y2=0
cc_435 N_A_863_98#_c_580_n N_VPWR_c_813_n 0.0085718f $X=4.43 $Y=2.465 $X2=0
+ $Y2=0
cc_436 N_A_863_98#_c_581_n N_VPWR_c_813_n 0.00752835f $X=6.155 $Y=1.765 $X2=0
+ $Y2=0
cc_437 N_A_863_98#_c_584_n N_VPWR_c_813_n 0.00862336f $X=6.66 $Y=2.045 $X2=0
+ $Y2=0
cc_438 N_A_863_98#_c_587_n N_VPWR_c_813_n 0.0120466f $X=5.37 $Y=2.815 $X2=0
+ $Y2=0
cc_439 N_A_863_98#_c_581_n N_Q_c_912_n 0.0140359f $X=6.155 $Y=1.765 $X2=0 $Y2=0
cc_440 N_A_863_98#_c_584_n N_Q_c_912_n 3.87665e-19 $X=6.66 $Y=2.045 $X2=0 $Y2=0
cc_441 N_A_863_98#_c_587_n N_Q_c_912_n 0.0447573f $X=5.37 $Y=2.815 $X2=0 $Y2=0
cc_442 N_A_863_98#_c_581_n N_Q_c_913_n 0.00401482f $X=6.155 $Y=1.765 $X2=0 $Y2=0
cc_443 N_A_863_98#_c_584_n N_Q_c_913_n 6.39334e-19 $X=6.66 $Y=2.045 $X2=0 $Y2=0
cc_444 N_A_863_98#_c_571_n N_Q_c_913_n 0.00593917f $X=6.065 $Y=1.485 $X2=0 $Y2=0
cc_445 N_A_863_98#_c_574_n N_Q_c_913_n 0.0115034f $X=5.37 $Y=1.985 $X2=0 $Y2=0
cc_446 N_A_863_98#_c_576_n N_Q_c_913_n 7.59e-19 $X=5.61 $Y=1.485 $X2=0 $Y2=0
cc_447 N_A_863_98#_c_588_n N_Q_c_913_n 0.0237215f $X=5.37 $Y=2.155 $X2=0 $Y2=0
cc_448 N_A_863_98#_c_581_n N_Q_c_909_n 0.00218881f $X=6.155 $Y=1.765 $X2=0 $Y2=0
cc_449 N_A_863_98#_M1013_g N_Q_c_909_n 0.00641464f $X=6.175 $Y=0.76 $X2=0 $Y2=0
cc_450 N_A_863_98#_c_568_n N_Q_c_909_n 0.0164053f $X=6.66 $Y=1.65 $X2=0 $Y2=0
cc_451 N_A_863_98#_c_569_n N_Q_c_909_n 6.39334e-19 $X=6.66 $Y=1.955 $X2=0 $Y2=0
cc_452 N_A_863_98#_c_571_n N_Q_c_909_n 0.0132825f $X=6.065 $Y=1.485 $X2=0 $Y2=0
cc_453 N_A_863_98#_c_573_n N_Q_c_909_n 0.00385371f $X=5.29 $Y=1.32 $X2=0 $Y2=0
cc_454 N_A_863_98#_c_574_n N_Q_c_909_n 0.00509287f $X=5.37 $Y=1.985 $X2=0 $Y2=0
cc_455 N_A_863_98#_c_576_n N_Q_c_909_n 0.02351f $X=5.61 $Y=1.485 $X2=0 $Y2=0
cc_456 N_A_863_98#_M1013_g Q 0.00815919f $X=6.175 $Y=0.76 $X2=0 $Y2=0
cc_457 N_A_863_98#_M1015_g Q 6.83062e-19 $X=6.675 $Y=0.855 $X2=0 $Y2=0
cc_458 N_A_863_98#_c_572_n Q 0.0173558f $X=5.185 $Y=0.515 $X2=0 $Y2=0
cc_459 N_A_863_98#_M1013_g Q 0.00207147f $X=6.175 $Y=0.76 $X2=0 $Y2=0
cc_460 N_A_863_98#_c_571_n Q 0.00479624f $X=6.065 $Y=1.485 $X2=0 $Y2=0
cc_461 N_A_863_98#_c_575_n Q 0.0173558f $X=5.197 $Y=1.07 $X2=0 $Y2=0
cc_462 N_A_863_98#_M1018_g N_VGND_c_963_n 0.00629296f $X=4.39 $Y=0.83 $X2=0
+ $Y2=0
cc_463 N_A_863_98#_c_572_n N_VGND_c_963_n 0.0276929f $X=5.185 $Y=0.515 $X2=0
+ $Y2=0
cc_464 N_A_863_98#_M1013_g N_VGND_c_964_n 0.00780298f $X=6.175 $Y=0.76 $X2=0
+ $Y2=0
cc_465 N_A_863_98#_c_568_n N_VGND_c_964_n 0.00755502f $X=6.66 $Y=1.65 $X2=0
+ $Y2=0
cc_466 N_A_863_98#_M1015_g N_VGND_c_964_n 0.00406495f $X=6.675 $Y=0.855 $X2=0
+ $Y2=0
cc_467 N_A_863_98#_M1015_g N_VGND_c_965_n 0.00401509f $X=6.675 $Y=0.855 $X2=0
+ $Y2=0
cc_468 N_A_863_98#_M1013_g N_VGND_c_966_n 0.00537471f $X=6.175 $Y=0.76 $X2=0
+ $Y2=0
cc_469 N_A_863_98#_c_572_n N_VGND_c_966_n 0.0157133f $X=5.185 $Y=0.515 $X2=0
+ $Y2=0
cc_470 N_A_863_98#_M1018_g N_VGND_c_970_n 0.00417968f $X=4.39 $Y=0.83 $X2=0
+ $Y2=0
cc_471 N_A_863_98#_M1015_g N_VGND_c_971_n 0.0041935f $X=6.675 $Y=0.855 $X2=0
+ $Y2=0
cc_472 N_A_863_98#_M1018_g N_VGND_c_973_n 0.00470816f $X=4.39 $Y=0.83 $X2=0
+ $Y2=0
cc_473 N_A_863_98#_M1013_g N_VGND_c_973_n 0.00539454f $X=6.175 $Y=0.76 $X2=0
+ $Y2=0
cc_474 N_A_863_98#_M1015_g N_VGND_c_973_n 0.00482046f $X=6.675 $Y=0.855 $X2=0
+ $Y2=0
cc_475 N_A_863_98#_c_572_n N_VGND_c_973_n 0.012935f $X=5.185 $Y=0.515 $X2=0
+ $Y2=0
cc_476 N_A_664_392#_c_685_n N_VPWR_c_817_n 0.00720002f $X=5.145 $Y=1.765 $X2=0
+ $Y2=0
cc_477 N_A_664_392#_c_685_n N_VPWR_c_820_n 0.00445602f $X=5.145 $Y=1.765 $X2=0
+ $Y2=0
cc_478 N_A_664_392#_c_685_n N_VPWR_c_813_n 0.00863697f $X=5.145 $Y=1.765 $X2=0
+ $Y2=0
cc_479 N_A_664_392#_c_685_n N_Q_c_913_n 0.00220962f $X=5.145 $Y=1.765 $X2=0
+ $Y2=0
cc_480 N_A_664_392#_M1006_g N_VGND_c_963_n 0.0109443f $X=4.97 $Y=0.74 $X2=0
+ $Y2=0
cc_481 N_A_664_392#_c_685_n N_VGND_c_963_n 0.00108892f $X=5.145 $Y=1.765 $X2=0
+ $Y2=0
cc_482 N_A_664_392#_c_688_n N_VGND_c_963_n 0.00295015f $X=3.865 $Y=1.65 $X2=0
+ $Y2=0
cc_483 N_A_664_392#_c_689_n N_VGND_c_963_n 0.0061936f $X=4.705 $Y=1.735 $X2=0
+ $Y2=0
cc_484 N_A_664_392#_c_690_n N_VGND_c_963_n 0.0113399f $X=4.87 $Y=1.405 $X2=0
+ $Y2=0
cc_485 N_A_664_392#_M1006_g N_VGND_c_966_n 0.00434272f $X=4.97 $Y=0.74 $X2=0
+ $Y2=0
cc_486 N_A_664_392#_M1006_g N_VGND_c_973_n 0.00830058f $X=4.97 $Y=0.74 $X2=0
+ $Y2=0
cc_487 N_A_1347_424#_c_773_n N_VPWR_c_818_n 0.0337457f $X=6.885 $Y=2.265 $X2=0
+ $Y2=0
cc_488 N_A_1347_424#_c_775_n N_VPWR_c_819_n 0.0100009f $X=7.66 $Y=1.765 $X2=0
+ $Y2=0
cc_489 N_A_1347_424#_c_770_n N_VPWR_c_819_n 0.0099853f $X=7.57 $Y=1.485 $X2=0
+ $Y2=0
cc_490 N_A_1347_424#_c_773_n N_VPWR_c_819_n 0.07899f $X=6.885 $Y=2.265 $X2=0
+ $Y2=0
cc_491 N_A_1347_424#_c_774_n N_VPWR_c_819_n 0.00413233f $X=7.155 $Y=1.485 $X2=0
+ $Y2=0
cc_492 N_A_1347_424#_c_773_n N_VPWR_c_822_n 0.0145938f $X=6.885 $Y=2.265 $X2=0
+ $Y2=0
cc_493 N_A_1347_424#_c_775_n N_VPWR_c_825_n 0.00439937f $X=7.66 $Y=1.765 $X2=0
+ $Y2=0
cc_494 N_A_1347_424#_c_775_n N_VPWR_c_813_n 0.00847525f $X=7.66 $Y=1.765 $X2=0
+ $Y2=0
cc_495 N_A_1347_424#_c_773_n N_VPWR_c_813_n 0.0120466f $X=6.885 $Y=2.265 $X2=0
+ $Y2=0
cc_496 N_A_1347_424#_c_772_n N_Q_c_909_n 0.00441678f $X=6.89 $Y=0.855 $X2=0
+ $Y2=0
cc_497 N_A_1347_424#_c_773_n N_Q_c_909_n 0.0118796f $X=6.885 $Y=2.265 $X2=0
+ $Y2=0
cc_498 N_A_1347_424#_c_774_n N_Q_c_909_n 0.00875204f $X=7.155 $Y=1.485 $X2=0
+ $Y2=0
cc_499 N_A_1347_424#_c_775_n Q_N 0.016982f $X=7.66 $Y=1.765 $X2=0 $Y2=0
cc_500 N_A_1347_424#_M1008_g Q_N 0.0187771f $X=7.665 $Y=0.74 $X2=0 $Y2=0
cc_501 N_A_1347_424#_c_771_n Q_N 0.0206976f $X=7.66 $Y=1.542 $X2=0 $Y2=0
cc_502 N_A_1347_424#_c_772_n Q_N 0.00536073f $X=6.89 $Y=0.855 $X2=0 $Y2=0
cc_503 N_A_1347_424#_c_773_n Q_N 0.00475831f $X=6.885 $Y=2.265 $X2=0 $Y2=0
cc_504 N_A_1347_424#_c_774_n Q_N 0.0131263f $X=7.155 $Y=1.485 $X2=0 $Y2=0
cc_505 N_A_1347_424#_c_772_n N_VGND_c_964_n 0.0231643f $X=6.89 $Y=0.855 $X2=0
+ $Y2=0
cc_506 N_A_1347_424#_M1008_g N_VGND_c_965_n 0.00647412f $X=7.665 $Y=0.74 $X2=0
+ $Y2=0
cc_507 N_A_1347_424#_c_770_n N_VGND_c_965_n 0.0100916f $X=7.57 $Y=1.485 $X2=0
+ $Y2=0
cc_508 N_A_1347_424#_c_772_n N_VGND_c_965_n 0.0376813f $X=6.89 $Y=0.855 $X2=0
+ $Y2=0
cc_509 N_A_1347_424#_c_774_n N_VGND_c_965_n 0.00263736f $X=7.155 $Y=1.485 $X2=0
+ $Y2=0
cc_510 N_A_1347_424#_c_772_n N_VGND_c_971_n 0.00787778f $X=6.89 $Y=0.855 $X2=0
+ $Y2=0
cc_511 N_A_1347_424#_M1008_g N_VGND_c_972_n 0.00434272f $X=7.665 $Y=0.74 $X2=0
+ $Y2=0
cc_512 N_A_1347_424#_M1008_g N_VGND_c_973_n 0.00828941f $X=7.665 $Y=0.74 $X2=0
+ $Y2=0
cc_513 N_A_1347_424#_c_772_n N_VGND_c_973_n 0.0106412f $X=6.89 $Y=0.855 $X2=0
+ $Y2=0
cc_514 N_VPWR_c_818_n N_Q_c_912_n 0.0673472f $X=6.38 $Y=2.265 $X2=0 $Y2=0
cc_515 N_VPWR_c_820_n N_Q_c_912_n 0.0158428f $X=6.295 $Y=3.33 $X2=0 $Y2=0
cc_516 N_VPWR_c_813_n N_Q_c_912_n 0.0130099f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_517 N_VPWR_c_819_n Q_N 0.0794554f $X=7.435 $Y=1.985 $X2=0 $Y2=0
cc_518 N_VPWR_c_825_n Q_N 0.014802f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_519 N_VPWR_c_813_n Q_N 0.0122072f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_520 Q N_VGND_c_964_n 0.0307458f $X=5.915 $Y=0.47 $X2=0 $Y2=0
cc_521 Q N_VGND_c_966_n 0.0134772f $X=5.915 $Y=0.47 $X2=0 $Y2=0
cc_522 Q N_VGND_c_973_n 0.0119466f $X=5.915 $Y=0.47 $X2=0 $Y2=0
cc_523 Q_N N_VGND_c_965_n 0.0294766f $X=7.835 $Y=0.47 $X2=0 $Y2=0
cc_524 Q_N N_VGND_c_972_n 0.014787f $X=7.835 $Y=0.47 $X2=0 $Y2=0
cc_525 Q_N N_VGND_c_973_n 0.012183f $X=7.835 $Y=0.47 $X2=0 $Y2=0
