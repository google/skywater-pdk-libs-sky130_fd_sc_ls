* File: sky130_fd_sc_ls__or4_1.pex.spice
* Created: Fri Aug 28 13:59:33 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__OR4_1%D 3 5 7 8 12
r26 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.485
+ $Y=1.585 $X2=0.485 $Y2=1.585
r27 8 12 7.84301 $w=3.58e-07 $l=2.45e-07 $layer=LI1_cond $X=0.24 $Y=1.6
+ $X2=0.485 $Y2=1.6
r28 5 11 61.7771 $w=2.82e-07 $l=3.45543e-07 $layer=POLY_cond $X=0.59 $Y=1.885
+ $X2=0.492 $Y2=1.585
r29 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.59 $Y=1.885
+ $X2=0.59 $Y2=2.46
r30 1 11 38.7026 $w=2.82e-07 $l=1.98167e-07 $layer=POLY_cond $X=0.565 $Y=1.42
+ $X2=0.492 $Y2=1.585
r31 1 3 299.968 $w=1.5e-07 $l=5.85e-07 $layer=POLY_cond $X=0.565 $Y=1.42
+ $X2=0.565 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_LS__OR4_1%C 3 5 7 8
r29 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.085
+ $Y=1.585 $X2=1.085 $Y2=1.585
r30 8 12 3.68142 $w=3.58e-07 $l=1.15e-07 $layer=LI1_cond $X=1.2 $Y=1.6 $X2=1.085
+ $Y2=1.6
r31 5 11 61.4066 $w=2.86e-07 $l=3.3541e-07 $layer=POLY_cond $X=1.01 $Y=1.885
+ $X2=1.085 $Y2=1.585
r32 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.01 $Y=1.885
+ $X2=1.01 $Y2=2.46
r33 1 11 38.6549 $w=2.86e-07 $l=2.05122e-07 $layer=POLY_cond $X=0.995 $Y=1.42
+ $X2=1.085 $Y2=1.585
r34 1 3 299.968 $w=1.5e-07 $l=5.85e-07 $layer=POLY_cond $X=0.995 $Y=1.42
+ $X2=0.995 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_LS__OR4_1%B 1 3 6 8
r29 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.655
+ $Y=1.585 $X2=1.655 $Y2=1.585
r30 4 11 38.6549 $w=2.86e-07 $l=1.98997e-07 $layer=POLY_cond $X=1.73 $Y=1.42
+ $X2=1.655 $Y2=1.585
r31 4 6 299.968 $w=1.5e-07 $l=5.85e-07 $layer=POLY_cond $X=1.73 $Y=1.42 $X2=1.73
+ $Y2=0.835
r32 1 11 61.4066 $w=2.86e-07 $l=3.3541e-07 $layer=POLY_cond $X=1.58 $Y=1.885
+ $X2=1.655 $Y2=1.585
r33 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.58 $Y=1.885
+ $X2=1.58 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_LS__OR4_1%A 1 3 6 8 12
c35 1 0 1.09557e-19 $X=2.15 $Y=1.885
r36 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.225
+ $Y=1.515 $X2=2.225 $Y2=1.515
r37 8 12 5.01062 $w=3.43e-07 $l=1.5e-07 $layer=LI1_cond $X=2.217 $Y=1.665
+ $X2=2.217 $Y2=1.515
r38 4 11 38.8084 $w=2.75e-07 $l=2.06325e-07 $layer=POLY_cond $X=2.32 $Y=1.35
+ $X2=2.227 $Y2=1.515
r39 4 6 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=2.32 $Y=1.35 $X2=2.32
+ $Y2=0.835
r40 1 11 74.7393 $w=2.75e-07 $l=4.06682e-07 $layer=POLY_cond $X=2.15 $Y=1.885
+ $X2=2.227 $Y2=1.515
r41 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.15 $Y=1.885
+ $X2=2.15 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_LS__OR4_1%A_44_392# 1 2 3 12 14 16 17 19 21 25 27 28 31
+ 33 35 36 39
r95 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.77
+ $Y=1.465 $X2=2.77 $Y2=1.465
r96 35 42 9.06394 $w=2.79e-07 $l=2.09893e-07 $layer=LI1_cond $X=2.645 $Y=1.63
+ $X2=2.747 $Y2=1.465
r97 35 36 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2.645 $Y=1.63
+ $X2=2.645 $Y2=1.95
r98 34 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.19 $Y=1.095
+ $X2=2.025 $Y2=1.095
r99 33 42 16.1792 $w=2.79e-07 $l=4.53971e-07 $layer=LI1_cond $X=2.56 $Y=1.095
+ $X2=2.747 $Y2=1.465
r100 33 34 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.56 $Y=1.095
+ $X2=2.19 $Y2=1.095
r101 29 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.025 $Y=1.01
+ $X2=2.025 $Y2=1.095
r102 29 31 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=2.025 $Y=1.01
+ $X2=2.025 $Y2=0.835
r103 27 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.86 $Y=1.095
+ $X2=2.025 $Y2=1.095
r104 27 28 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=1.86 $Y=1.095
+ $X2=0.945 $Y2=1.095
r105 23 28 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.78 $Y=1.01
+ $X2=0.945 $Y2=1.095
r106 23 25 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=0.78 $Y=1.01
+ $X2=0.78 $Y2=0.835
r107 22 38 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.53 $Y=2.035
+ $X2=0.365 $Y2=2.035
r108 21 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.56 $Y=2.035
+ $X2=2.645 $Y2=1.95
r109 21 22 132.439 $w=1.68e-07 $l=2.03e-06 $layer=LI1_cond $X=2.56 $Y=2.035
+ $X2=0.53 $Y2=2.035
r110 17 38 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.365 $Y=2.12
+ $X2=0.365 $Y2=2.035
r111 17 19 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=0.365 $Y=2.12
+ $X2=0.365 $Y2=2.815
r112 14 43 61.4066 $w=2.86e-07 $l=3.33167e-07 $layer=POLY_cond $X=2.84 $Y=1.765
+ $X2=2.77 $Y2=1.465
r113 14 16 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.84 $Y=1.765
+ $X2=2.84 $Y2=2.4
r114 10 43 38.6549 $w=2.86e-07 $l=1.92678e-07 $layer=POLY_cond $X=2.83 $Y=1.3
+ $X2=2.77 $Y2=1.465
r115 10 12 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.83 $Y=1.3
+ $X2=2.83 $Y2=0.74
r116 3 38 400 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=1 $X=0.22
+ $Y=1.96 $X2=0.365 $Y2=2.115
r117 3 19 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.22
+ $Y=1.96 $X2=0.365 $Y2=2.815
r118 2 31 182 $w=1.7e-07 $l=3.68951e-07 $layer=licon1_NDIFF $count=1 $X=1.805
+ $Y=0.56 $X2=2.025 $Y2=0.835
r119 1 25 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=0.64
+ $Y=0.56 $X2=0.78 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_LS__OR4_1%VPWR 1 6 8 10 17 18 21
r27 21 22 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r28 18 22 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.16 $Y2=3.33
r29 17 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r30 15 21 10.0494 $w=1.7e-07 $l=2.08e-07 $layer=LI1_cond $X=2.565 $Y=3.33
+ $X2=2.357 $Y2=3.33
r31 15 17 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=2.565 $Y=3.33
+ $X2=3.12 $Y2=3.33
r32 12 13 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r33 10 21 10.0494 $w=1.7e-07 $l=2.07e-07 $layer=LI1_cond $X=2.15 $Y=3.33
+ $X2=2.357 $Y2=3.33
r34 10 12 124.61 $w=1.68e-07 $l=1.91e-06 $layer=LI1_cond $X=2.15 $Y=3.33
+ $X2=0.24 $Y2=3.33
r35 8 22 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r36 8 13 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.24 $Y2=3.33
r37 4 21 1.57254 $w=4.15e-07 $l=8.5e-08 $layer=LI1_cond $X=2.357 $Y=3.245
+ $X2=2.357 $Y2=3.33
r38 4 6 21.9381 $w=4.13e-07 $l=7.9e-07 $layer=LI1_cond $X=2.357 $Y=3.245
+ $X2=2.357 $Y2=2.455
r39 1 6 300 $w=1.7e-07 $l=5.65044e-07 $layer=licon1_PDIFF $count=2 $X=2.225
+ $Y=1.96 $X2=2.375 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_LS__OR4_1%X 1 2 9 13 14 15 16 23 32
c23 14 0 1.09557e-19 $X=3.035 $Y=1.95
r24 21 23 0.860491 $w=3.73e-07 $l=2.8e-08 $layer=LI1_cond $X=3.087 $Y=2.007
+ $X2=3.087 $Y2=2.035
r25 15 16 11.3708 $w=3.73e-07 $l=3.7e-07 $layer=LI1_cond $X=3.087 $Y=2.405
+ $X2=3.087 $Y2=2.775
r26 14 21 0.891223 $w=3.73e-07 $l=2.9e-08 $layer=LI1_cond $X=3.087 $Y=1.978
+ $X2=3.087 $Y2=2.007
r27 14 32 8.33934 $w=3.73e-07 $l=1.58e-07 $layer=LI1_cond $X=3.087 $Y=1.978
+ $X2=3.087 $Y2=1.82
r28 14 15 10.5103 $w=3.73e-07 $l=3.42e-07 $layer=LI1_cond $X=3.087 $Y=2.063
+ $X2=3.087 $Y2=2.405
r29 14 23 0.860491 $w=3.73e-07 $l=2.8e-08 $layer=LI1_cond $X=3.087 $Y=2.063
+ $X2=3.087 $Y2=2.035
r30 13 32 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.19 $Y=1.13 $X2=3.19
+ $Y2=1.82
r31 7 13 8.16989 $w=3.13e-07 $l=1.57e-07 $layer=LI1_cond $X=3.117 $Y=0.973
+ $X2=3.117 $Y2=1.13
r32 7 9 16.7562 $w=3.13e-07 $l=4.58e-07 $layer=LI1_cond $X=3.117 $Y=0.973
+ $X2=3.117 $Y2=0.515
r33 2 14 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.915
+ $Y=1.84 $X2=3.065 $Y2=1.985
r34 2 16 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.915
+ $Y=1.84 $X2=3.065 $Y2=2.815
r35 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.905
+ $Y=0.37 $X2=3.045 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__OR4_1%VGND 1 2 3 10 12 14 18 22 24 26 33 34 40 43
r46 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r47 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r48 38 41 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r49 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r50 34 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r51 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r52 31 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.78 $Y=0 $X2=2.615
+ $Y2=0
r53 31 33 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.78 $Y=0 $X2=3.12
+ $Y2=0
r54 30 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r55 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r56 27 40 10.9443 $w=1.7e-07 $l=2.38e-07 $layer=LI1_cond $X=1.6 $Y=0 $X2=1.362
+ $Y2=0
r57 27 29 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.6 $Y=0 $X2=2.16
+ $Y2=0
r58 26 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.45 $Y=0 $X2=2.615
+ $Y2=0
r59 26 29 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=2.45 $Y=0 $X2=2.16
+ $Y2=0
r60 24 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r61 24 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r62 20 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.615 $Y=0.085
+ $X2=2.615 $Y2=0
r63 20 22 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=2.615 $Y=0.085
+ $X2=2.615 $Y2=0.675
r64 16 40 1.94084 $w=4.75e-07 $l=8.5e-08 $layer=LI1_cond $X=1.362 $Y=0.085
+ $X2=1.362 $Y2=0
r65 16 18 14.8566 $w=4.73e-07 $l=5.9e-07 $layer=LI1_cond $X=1.362 $Y=0.085
+ $X2=1.362 $Y2=0.675
r66 15 37 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.222
+ $Y2=0
r67 14 40 10.9443 $w=1.7e-07 $l=2.37e-07 $layer=LI1_cond $X=1.125 $Y=0 $X2=1.362
+ $Y2=0
r68 14 15 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.125 $Y=0 $X2=0.445
+ $Y2=0
r69 10 37 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.222 $Y2=0
r70 10 12 26.1919 $w=3.28e-07 $l=7.5e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.28 $Y2=0.835
r71 3 22 182 $w=1.7e-07 $l=2.71477e-07 $layer=licon1_NDIFF $count=1 $X=2.395
+ $Y=0.56 $X2=2.615 $Y2=0.675
r72 2 18 182 $w=1.7e-07 $l=3.4271e-07 $layer=licon1_NDIFF $count=1 $X=1.07
+ $Y=0.56 $X2=1.36 $Y2=0.675
r73 1 12 182 $w=1.7e-07 $l=3.67083e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.56 $X2=0.35 $Y2=0.835
.ends

