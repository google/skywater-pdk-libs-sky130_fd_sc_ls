* File: sky130_fd_sc_ls__a2111oi_1.pex.spice
* Created: Fri Aug 28 12:48:11 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__A2111OI_1%D1 1 3 6 8 12
r24 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.63
+ $Y=1.515 $X2=0.63 $Y2=1.515
r25 8 12 4.67207 $w=3.68e-07 $l=1.5e-07 $layer=LI1_cond $X=0.65 $Y=1.665
+ $X2=0.65 $Y2=1.515
r26 4 11 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=0.72 $Y=1.35
+ $X2=0.63 $Y2=1.515
r27 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.72 $Y=1.35 $X2=0.72
+ $Y2=0.74
r28 1 11 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=0.705 $Y=1.765
+ $X2=0.63 $Y2=1.515
r29 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.705 $Y=1.765
+ $X2=0.705 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__A2111OI_1%C1 1 3 6 8 12
c32 1 0 1.48944e-19 $X=1.095 $Y=1.765
r33 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.17
+ $Y=1.515 $X2=1.17 $Y2=1.515
r34 8 12 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.17 $Y=1.665
+ $X2=1.17 $Y2=1.515
r35 4 11 38.5562 $w=2.99e-07 $l=1.74714e-07 $layer=POLY_cond $X=1.15 $Y=1.35
+ $X2=1.17 $Y2=1.515
r36 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.15 $Y=1.35 $X2=1.15
+ $Y2=0.74
r37 1 11 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=1.095 $Y=1.765
+ $X2=1.17 $Y2=1.515
r38 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.095 $Y=1.765
+ $X2=1.095 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__A2111OI_1%B1 1 3 6 8 12
r30 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.71
+ $Y=1.515 $X2=1.71 $Y2=1.515
r31 8 12 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.71 $Y=1.665
+ $X2=1.71 $Y2=1.515
r32 4 11 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=1.8 $Y=1.35
+ $X2=1.71 $Y2=1.515
r33 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.8 $Y=1.35 $X2=1.8
+ $Y2=0.74
r34 1 11 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=1.635 $Y=1.765
+ $X2=1.71 $Y2=1.515
r35 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.635 $Y=1.765
+ $X2=1.635 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__A2111OI_1%A1 1 3 6 8 12
r31 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.25
+ $Y=1.515 $X2=2.25 $Y2=1.515
r32 8 12 4.67207 $w=3.68e-07 $l=1.5e-07 $layer=LI1_cond $X=2.23 $Y=1.665
+ $X2=2.23 $Y2=1.515
r33 4 11 38.5562 $w=2.99e-07 $l=1.74714e-07 $layer=POLY_cond $X=2.23 $Y=1.35
+ $X2=2.25 $Y2=1.515
r34 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.23 $Y=1.35 $X2=2.23
+ $Y2=0.74
r35 1 11 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=2.175 $Y=1.765
+ $X2=2.25 $Y2=1.515
r36 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.175 $Y=1.765
+ $X2=2.175 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__A2111OI_1%A2 1 3 4 6 7
r25 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.79
+ $Y=1.385 $X2=2.79 $Y2=1.385
r26 7 11 10.2785 $w=3.68e-07 $l=3.3e-07 $layer=LI1_cond $X=3.12 $Y=1.365
+ $X2=2.79 $Y2=1.365
r27 4 10 77.2841 $w=2.7e-07 $l=4.15812e-07 $layer=POLY_cond $X=2.715 $Y=1.765
+ $X2=2.79 $Y2=1.385
r28 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.715 $Y=1.765
+ $X2=2.715 $Y2=2.4
r29 1 10 38.9026 $w=2.7e-07 $l=2.05122e-07 $layer=POLY_cond $X=2.7 $Y=1.22
+ $X2=2.79 $Y2=1.385
r30 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.7 $Y=1.22 $X2=2.7
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__A2111OI_1%Y 1 2 3 11 12 13 16 18 22 24 25 27 29
r58 27 29 5.68544 $w=1.028e-06 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=2.465
+ $X2=1.2 $Y2=2.465
r59 27 43 2.84272 $w=1.028e-06 $l=2.4e-07 $layer=LI1_cond $X=0.72 $Y=2.465
+ $X2=0.48 $Y2=2.465
r60 25 43 2.84272 $w=1.028e-06 $l=2.4e-07 $layer=LI1_cond $X=0.24 $Y=2.465
+ $X2=0.48 $Y2=2.465
r61 25 37 0.35534 $w=1.028e-06 $l=3e-08 $layer=LI1_cond $X=0.24 $Y=2.465
+ $X2=0.21 $Y2=2.465
r62 20 22 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=2.015 $Y=1.01
+ $X2=2.015 $Y2=0.515
r63 19 24 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.1 $Y=1.095
+ $X2=0.975 $Y2=1.095
r64 18 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.85 $Y=1.095
+ $X2=2.015 $Y2=1.01
r65 18 19 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=1.85 $Y=1.095
+ $X2=1.1 $Y2=1.095
r66 14 24 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.975 $Y=1.01
+ $X2=0.975 $Y2=1.095
r67 14 16 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=0.975 $Y=1.01
+ $X2=0.975 $Y2=0.515
r68 12 24 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.85 $Y=1.095
+ $X2=0.975 $Y2=1.095
r69 12 13 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=0.85 $Y=1.095
+ $X2=0.295 $Y2=1.095
r70 11 37 11.9281 $w=1.7e-07 $l=5.15e-07 $layer=LI1_cond $X=0.21 $Y=1.95
+ $X2=0.21 $Y2=2.465
r71 10 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.21 $Y=1.18
+ $X2=0.295 $Y2=1.095
r72 10 11 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=0.21 $Y=1.18
+ $X2=0.21 $Y2=1.95
r73 3 43 400 $w=1.7e-07 $l=1.03562e-06 $layer=licon1_PDIFF $count=1 $X=0.355
+ $Y=1.84 $X2=0.48 $Y2=2.815
r74 3 43 400 $w=1.7e-07 $l=2.498e-07 $layer=licon1_PDIFF $count=1 $X=0.355
+ $Y=1.84 $X2=0.48 $Y2=2.035
r75 2 22 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.875
+ $Y=0.37 $X2=2.015 $Y2=0.515
r76 1 16 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.795
+ $Y=0.37 $X2=0.935 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__A2111OI_1%A_342_368# 1 2 7 9 11 13 15
c27 7 0 1.48944e-19 $X=1.88 $Y=2.12
r28 13 20 3.0656 $w=3.3e-07 $l=1.5e-07 $layer=LI1_cond $X=2.94 $Y=2.12 $X2=2.94
+ $Y2=1.97
r29 13 15 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=2.94 $Y=2.12
+ $X2=2.94 $Y2=2.815
r30 12 18 5.55669 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=2.065 $Y=2.035
+ $X2=1.88 $Y2=2.035
r31 11 20 4.70058 $w=1.7e-07 $l=1.94808e-07 $layer=LI1_cond $X=2.775 $Y=2.035
+ $X2=2.94 $Y2=1.97
r32 11 12 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=2.775 $Y=2.035
+ $X2=2.065 $Y2=2.035
r33 7 18 2.55307 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.88 $Y=2.12 $X2=1.88
+ $Y2=2.035
r34 7 9 9.81134 $w=3.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.88 $Y=2.12 $X2=1.88
+ $Y2=2.435
r35 2 20 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.79
+ $Y=1.84 $X2=2.94 $Y2=1.985
r36 2 15 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.79
+ $Y=1.84 $X2=2.94 $Y2=2.815
r37 1 18 600 $w=1.7e-07 $l=2.66786e-07 $layer=licon1_PDIFF $count=1 $X=1.71
+ $Y=1.84 $X2=1.88 $Y2=2.035
r38 1 9 300 $w=1.7e-07 $l=6.74667e-07 $layer=licon1_PDIFF $count=2 $X=1.71
+ $Y=1.84 $X2=1.88 $Y2=2.435
.ends

.subckt PM_SKY130_FD_SC_LS__A2111OI_1%VPWR 1 6 9 10 11 21 22
r29 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r30 19 22 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r31 18 19 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r32 14 18 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=2.16 $Y2=3.33
r33 14 15 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r34 11 19 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r35 11 15 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.24 $Y2=3.33
r36 9 18 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=2.235 $Y=3.33
+ $X2=2.16 $Y2=3.33
r37 9 10 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=2.235 $Y=3.33
+ $X2=2.42 $Y2=3.33
r38 8 21 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=2.605 $Y=3.33
+ $X2=3.12 $Y2=3.33
r39 8 10 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=2.605 $Y=3.33
+ $X2=2.42 $Y2=3.33
r40 4 10 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.42 $Y=3.245 $X2=2.42
+ $Y2=3.33
r41 4 6 26.0078 $w=3.68e-07 $l=8.35e-07 $layer=LI1_cond $X=2.42 $Y=3.245
+ $X2=2.42 $Y2=2.41
r42 1 6 300 $w=1.7e-07 $l=6.49461e-07 $layer=licon1_PDIFF $count=2 $X=2.25
+ $Y=1.84 $X2=2.42 $Y2=2.41
.ends

.subckt PM_SKY130_FD_SC_LS__A2111OI_1%VGND 1 2 3 12 16 20 23 24 26 27 28 29 30
+ 31 48
r41 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r42 45 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r43 44 45 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r44 41 44 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r45 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r46 35 39 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r47 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r48 31 45 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r49 31 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r50 31 41 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r51 29 44 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=2.75 $Y=0 $X2=2.64
+ $Y2=0
r52 29 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.75 $Y=0 $X2=2.915
+ $Y2=0
r53 28 47 2.87059 $w=1.7e-07 $l=4e-08 $layer=LI1_cond $X=3.08 $Y=0 $X2=3.12
+ $Y2=0
r54 28 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.08 $Y=0 $X2=2.915
+ $Y2=0
r55 27 41 9.97069 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=1.475 $Y=0 $X2=1.68
+ $Y2=0
r56 26 38 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=1.27 $Y=0 $X2=1.2
+ $Y2=0
r57 26 27 9.97069 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=1.27 $Y=0 $X2=1.475
+ $Y2=0
r58 23 34 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=0.34 $Y=0 $X2=0.24
+ $Y2=0
r59 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.34 $Y=0 $X2=0.505
+ $Y2=0
r60 22 38 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=0.67 $Y=0 $X2=1.2
+ $Y2=0
r61 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.67 $Y=0 $X2=0.505
+ $Y2=0
r62 18 30 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.915 $Y=0.085
+ $X2=2.915 $Y2=0
r63 18 20 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.915 $Y=0.085
+ $X2=2.915 $Y2=0.515
r64 14 27 1.53834 $w=4.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.475 $Y=0.085
+ $X2=1.475 $Y2=0
r65 14 16 16.5839 $w=4.08e-07 $l=5.9e-07 $layer=LI1_cond $X=1.475 $Y=0.085
+ $X2=1.475 $Y2=0.675
r66 10 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.505 $Y=0.085
+ $X2=0.505 $Y2=0
r67 10 12 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=0.505 $Y=0.085
+ $X2=0.505 $Y2=0.675
r68 3 20 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.775
+ $Y=0.37 $X2=2.915 $Y2=0.515
r69 2 16 182 $w=1.7e-07 $l=4.1143e-07 $layer=licon1_NDIFF $count=1 $X=1.225
+ $Y=0.37 $X2=1.475 $Y2=0.675
r70 1 12 182 $w=1.7e-07 $l=3.62146e-07 $layer=licon1_NDIFF $count=1 $X=0.38
+ $Y=0.37 $X2=0.505 $Y2=0.675
.ends

