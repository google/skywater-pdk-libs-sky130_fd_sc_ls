* File: sky130_fd_sc_ls__clkbuf_4.pex.spice
* Created: Wed Sep  2 10:57:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__CLKBUF_4%A_83_270# 1 2 7 9 12 16 18 20 23 25 27 30
+ 32 34 35 40 44 49 53 54 58 68
c113 53 0 5.35093e-20 $X=1.885 $Y=1.55
r114 68 69 1.95405 $w=3.7e-07 $l=1.5e-08 $layer=POLY_cond $X=1.84 $Y=1.557
+ $X2=1.855 $Y2=1.557
r115 65 66 4.55946 $w=3.7e-07 $l=3.5e-08 $layer=POLY_cond $X=1.37 $Y=1.557
+ $X2=1.405 $Y2=1.557
r116 62 63 1.95405 $w=3.7e-07 $l=1.5e-08 $layer=POLY_cond $X=0.94 $Y=1.557
+ $X2=0.955 $Y2=1.557
r117 61 62 56.0162 $w=3.7e-07 $l=4.3e-07 $layer=POLY_cond $X=0.51 $Y=1.557
+ $X2=0.94 $Y2=1.557
r118 60 61 0.651351 $w=3.7e-07 $l=5e-09 $layer=POLY_cond $X=0.505 $Y=1.557
+ $X2=0.51 $Y2=1.557
r119 56 58 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=2.59 $Y=0.645
+ $X2=2.71 $Y2=0.645
r120 52 68 15.6324 $w=3.7e-07 $l=1.2e-07 $layer=POLY_cond $X=1.72 $Y=1.557
+ $X2=1.84 $Y2=1.557
r121 52 66 41.0351 $w=3.7e-07 $l=3.15e-07 $layer=POLY_cond $X=1.72 $Y=1.557
+ $X2=1.405 $Y2=1.557
r122 51 53 8.64761 $w=3.98e-07 $l=1.65e-07 $layer=LI1_cond $X=1.72 $Y=1.55
+ $X2=1.885 $Y2=1.55
r123 51 52 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.72
+ $Y=1.515 $X2=1.72 $Y2=1.515
r124 49 54 3.40559 $w=2.75e-07 $l=1.41244e-07 $layer=LI1_cond $X=2.71 $Y=1.58
+ $X2=2.605 $Y2=1.665
r125 48 58 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.71 $Y=0.81
+ $X2=2.71 $Y2=0.645
r126 48 49 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=2.71 $Y=0.81
+ $X2=2.71 $Y2=1.58
r127 44 46 25.1718 $w=3.78e-07 $l=8.3e-07 $layer=LI1_cond $X=2.605 $Y=1.985
+ $X2=2.605 $Y2=2.815
r128 42 54 3.40559 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=2.605 $Y=1.75
+ $X2=2.605 $Y2=1.665
r129 42 44 7.12695 $w=3.78e-07 $l=2.35e-07 $layer=LI1_cond $X=2.605 $Y=1.75
+ $X2=2.605 $Y2=1.985
r130 40 54 3.11956 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.415 $Y=1.665
+ $X2=2.605 $Y2=1.665
r131 40 53 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=2.415 $Y=1.665
+ $X2=1.885 $Y2=1.665
r132 38 65 42.9892 $w=3.7e-07 $l=3.3e-07 $layer=POLY_cond $X=1.04 $Y=1.557
+ $X2=1.37 $Y2=1.557
r133 38 63 11.073 $w=3.7e-07 $l=8.5e-08 $layer=POLY_cond $X=1.04 $Y=1.557
+ $X2=0.955 $Y2=1.557
r134 37 38 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.04
+ $Y=1.515 $X2=1.04 $Y2=1.515
r135 35 51 1.00839 $w=3.98e-07 $l=3.5e-08 $layer=LI1_cond $X=1.685 $Y=1.55
+ $X2=1.72 $Y2=1.55
r136 35 37 18.5831 $w=3.98e-07 $l=6.45e-07 $layer=LI1_cond $X=1.685 $Y=1.55
+ $X2=1.04 $Y2=1.55
r137 32 69 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.855 $Y=1.765
+ $X2=1.855 $Y2=1.557
r138 32 34 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.855 $Y=1.765
+ $X2=1.855 $Y2=2.4
r139 28 68 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.84 $Y=1.35
+ $X2=1.84 $Y2=1.557
r140 28 30 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=1.84 $Y=1.35
+ $X2=1.84 $Y2=0.58
r141 25 66 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.405 $Y=1.765
+ $X2=1.405 $Y2=1.557
r142 25 27 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.405 $Y=1.765
+ $X2=1.405 $Y2=2.4
r143 21 65 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.37 $Y=1.35
+ $X2=1.37 $Y2=1.557
r144 21 23 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=1.37 $Y=1.35
+ $X2=1.37 $Y2=0.58
r145 18 63 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.955 $Y=1.765
+ $X2=0.955 $Y2=1.557
r146 18 20 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.955 $Y=1.765
+ $X2=0.955 $Y2=2.4
r147 14 62 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.94 $Y=1.35
+ $X2=0.94 $Y2=1.557
r148 14 16 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=0.94 $Y=1.35
+ $X2=0.94 $Y2=0.58
r149 10 61 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.51 $Y=1.35
+ $X2=0.51 $Y2=1.557
r150 10 12 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=0.51 $Y=1.35
+ $X2=0.51 $Y2=0.58
r151 7 60 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=1.557
r152 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.4
r153 2 46 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.43
+ $Y=1.84 $X2=2.58 $Y2=2.815
r154 2 44 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.43
+ $Y=1.84 $X2=2.58 $Y2=1.985
r155 1 56 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=2.445
+ $Y=0.37 $X2=2.59 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_LS__CLKBUF_4%A 2 3 5 8 10 13 14
c40 13 0 5.35093e-20 $X=2.32 $Y=1.245
r41 13 16 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.32 $Y=1.245
+ $X2=2.32 $Y2=1.41
r42 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.32 $Y=1.245
+ $X2=2.32 $Y2=1.08
r43 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.32
+ $Y=1.245 $X2=2.32 $Y2=1.245
r44 10 14 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=2.16 $Y=1.245
+ $X2=2.32 $Y2=1.245
r45 8 15 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=2.37 $Y=0.58 $X2=2.37
+ $Y2=1.08
r46 3 5 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.355 $Y=1.765
+ $X2=2.355 $Y2=2.4
r47 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.355 $Y=1.675 $X2=2.355
+ $Y2=1.765
r48 2 16 103.008 $w=1.8e-07 $l=2.65e-07 $layer=POLY_cond $X=2.355 $Y=1.675
+ $X2=2.355 $Y2=1.41
.ends

.subckt PM_SKY130_FD_SC_LS__CLKBUF_4%VPWR 1 2 3 10 12 18 22 27 28 29 35 41 42 48
r44 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r45 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r46 42 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r47 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r48 39 48 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.245 $Y=3.33
+ $X2=2.12 $Y2=3.33
r49 39 41 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=2.245 $Y=3.33
+ $X2=2.64 $Y2=3.33
r50 38 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r51 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r52 35 48 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.995 $Y=3.33
+ $X2=2.12 $Y2=3.33
r53 35 37 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.995 $Y=3.33
+ $X2=1.68 $Y2=3.33
r54 34 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r55 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r56 31 45 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.182 $Y2=3.33
r57 31 33 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.72 $Y2=3.33
r58 29 38 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.68 $Y2=3.33
r59 29 34 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=0.72 $Y2=3.33
r60 27 33 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.015 $Y=3.33
+ $X2=0.72 $Y2=3.33
r61 27 28 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.015 $Y=3.33
+ $X2=1.14 $Y2=3.33
r62 26 37 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=1.265 $Y=3.33
+ $X2=1.68 $Y2=3.33
r63 26 28 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.265 $Y=3.33
+ $X2=1.14 $Y2=3.33
r64 22 25 33.6513 $w=2.48e-07 $l=7.3e-07 $layer=LI1_cond $X=2.12 $Y=2.085
+ $X2=2.12 $Y2=2.815
r65 20 48 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.12 $Y=3.245
+ $X2=2.12 $Y2=3.33
r66 20 25 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=2.12 $Y=3.245
+ $X2=2.12 $Y2=2.815
r67 16 28 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=3.245
+ $X2=1.14 $Y2=3.33
r68 16 18 37.8001 $w=2.48e-07 $l=8.2e-07 $layer=LI1_cond $X=1.14 $Y=3.245
+ $X2=1.14 $Y2=2.425
r69 12 15 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=0.24 $Y=1.985
+ $X2=0.24 $Y2=2.815
r70 10 45 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.182 $Y2=3.33
r71 10 15 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.24 $Y2=2.815
r72 3 25 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.93
+ $Y=1.84 $X2=2.08 $Y2=2.815
r73 3 22 400 $w=1.7e-07 $l=3.11087e-07 $layer=licon1_PDIFF $count=1 $X=1.93
+ $Y=1.84 $X2=2.08 $Y2=2.085
r74 2 18 300 $w=1.7e-07 $l=6.55725e-07 $layer=licon1_PDIFF $count=2 $X=1.03
+ $Y=1.84 $X2=1.18 $Y2=2.425
r75 1 15 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r76 1 12 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_LS__CLKBUF_4%X 1 2 3 4 14 17 19 21 25 27 29 32 35 36 47
r67 40 47 1.92074 $w=3.28e-07 $l=5.5e-08 $layer=LI1_cond $X=0.725 $Y=0.98
+ $X2=0.725 $Y2=0.925
r68 36 40 3.70735 $w=2.5e-07 $l=9.12688e-08 $layer=LI1_cond $X=0.712 $Y=1.065
+ $X2=0.725 $Y2=0.98
r69 36 47 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=0.725 $Y=0.91
+ $X2=0.725 $Y2=0.925
r70 35 36 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=0.725 $Y=0.555
+ $X2=0.725 $Y2=0.91
r71 27 34 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.63 $Y=2.09 $X2=1.63
+ $Y2=2.005
r72 27 29 25.3188 $w=3.28e-07 $l=7.25e-07 $layer=LI1_cond $X=1.63 $Y=2.09
+ $X2=1.63 $Y2=2.815
r73 23 25 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=1.585 $Y=0.98 $X2=1.585
+ $Y2=0.58
r74 22 36 2.76166 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=0.89 $Y=1.065
+ $X2=0.712 $Y2=1.065
r75 21 23 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.42 $Y=1.065
+ $X2=1.585 $Y2=0.98
r76 21 22 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.42 $Y=1.065
+ $X2=0.89 $Y2=1.065
r77 20 32 2.36881 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=0.815 $Y=2.005
+ $X2=0.675 $Y2=2.005
r78 19 34 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.465 $Y=2.005
+ $X2=1.63 $Y2=2.005
r79 19 20 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.465 $Y=2.005
+ $X2=0.815 $Y2=2.005
r80 15 32 4.06715 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=0.675 $Y=2.09
+ $X2=0.675 $Y2=2.005
r81 15 17 29.84 $w=2.78e-07 $l=7.25e-07 $layer=LI1_cond $X=0.675 $Y=2.09
+ $X2=0.675 $Y2=2.815
r82 14 32 4.06715 $w=2.25e-07 $l=1.09087e-07 $layer=LI1_cond $X=0.62 $Y=1.92
+ $X2=0.675 $Y2=2.005
r83 13 36 3.70735 $w=2.5e-07 $l=1.27609e-07 $layer=LI1_cond $X=0.62 $Y=1.15
+ $X2=0.712 $Y2=1.065
r84 13 14 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=0.62 $Y=1.15
+ $X2=0.62 $Y2=1.92
r85 4 34 400 $w=1.7e-07 $l=3.11087e-07 $layer=licon1_PDIFF $count=1 $X=1.48
+ $Y=1.84 $X2=1.63 $Y2=2.085
r86 4 29 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.48
+ $Y=1.84 $X2=1.63 $Y2=2.815
r87 3 32 400 $w=1.7e-07 $l=3.11087e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.84 $X2=0.73 $Y2=2.085
r88 3 17 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.84 $X2=0.73 $Y2=2.815
r89 2 25 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.445
+ $Y=0.37 $X2=1.585 $Y2=0.58
r90 1 35 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.585
+ $Y=0.37 $X2=0.725 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_LS__CLKBUF_4%VGND 1 2 3 10 12 16 20 23 24 25 31 37 38 44
r40 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r41 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r42 38 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r43 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r44 35 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.25 $Y=0 $X2=2.085
+ $Y2=0
r45 35 37 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=2.25 $Y=0 $X2=2.64
+ $Y2=0
r46 34 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r47 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r48 31 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.92 $Y=0 $X2=2.085
+ $Y2=0
r49 31 33 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r50 30 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r51 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r52 27 41 3.99177 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.38 $Y=0 $X2=0.19
+ $Y2=0
r53 27 29 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.38 $Y=0 $X2=0.72
+ $Y2=0
r54 25 34 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.68
+ $Y2=0
r55 25 30 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=0.72
+ $Y2=0
r56 23 29 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.07 $Y=0 $X2=0.72
+ $Y2=0
r57 23 24 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.07 $Y=0 $X2=1.155
+ $Y2=0
r58 22 33 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=1.24 $Y=0 $X2=1.68
+ $Y2=0
r59 22 24 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.24 $Y=0 $X2=1.155
+ $Y2=0
r60 18 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.085 $Y=0.085
+ $X2=2.085 $Y2=0
r61 18 20 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=2.085 $Y=0.085
+ $X2=2.085 $Y2=0.58
r62 14 24 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.155 $Y=0.085
+ $X2=1.155 $Y2=0
r63 14 16 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=1.155 $Y=0.085
+ $X2=1.155 $Y2=0.58
r64 10 41 3.1514 $w=2.5e-07 $l=1.12916e-07 $layer=LI1_cond $X=0.255 $Y=0.085
+ $X2=0.19 $Y2=0
r65 10 12 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=0.255 $Y=0.085
+ $X2=0.255 $Y2=0.58
r66 3 20 182 $w=1.7e-07 $l=2.82489e-07 $layer=licon1_NDIFF $count=1 $X=1.915
+ $Y=0.37 $X2=2.085 $Y2=0.58
r67 2 16 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.015
+ $Y=0.37 $X2=1.155 $Y2=0.58
r68 1 12 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.15
+ $Y=0.37 $X2=0.295 $Y2=0.58
.ends

