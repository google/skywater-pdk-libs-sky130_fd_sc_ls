* File: sky130_fd_sc_ls__a21oi_4.pxi.spice
* Created: Fri Aug 28 12:52:22 2020
* 
x_PM_SKY130_FD_SC_LS__A21OI_4%A2 N_A2_c_100_n N_A2_M1002_g N_A2_M1001_g
+ N_A2_c_101_n N_A2_M1003_g N_A2_M1013_g N_A2_c_102_n N_A2_M1005_g N_A2_M1014_g
+ N_A2_c_103_n N_A2_M1018_g N_A2_M1015_g A2 A2 A2 N_A2_c_99_n
+ PM_SKY130_FD_SC_LS__A21OI_4%A2
x_PM_SKY130_FD_SC_LS__A21OI_4%A1 N_A1_M1009_g N_A1_c_186_n N_A1_M1000_g
+ N_A1_M1012_g N_A1_c_187_n N_A1_M1006_g N_A1_M1020_g N_A1_c_188_n N_A1_M1010_g
+ N_A1_M1021_g N_A1_c_189_n N_A1_M1016_g A1 A1 N_A1_c_184_n N_A1_c_185_n
+ PM_SKY130_FD_SC_LS__A21OI_4%A1
x_PM_SKY130_FD_SC_LS__A21OI_4%B1 N_B1_c_273_n N_B1_M1004_g N_B1_c_274_n
+ N_B1_M1007_g N_B1_M1008_g N_B1_c_275_n N_B1_M1011_g N_B1_M1019_g N_B1_c_269_n
+ N_B1_c_270_n N_B1_c_278_n N_B1_M1017_g N_B1_c_271_n B1 B1 N_B1_c_272_n
+ PM_SKY130_FD_SC_LS__A21OI_4%B1
x_PM_SKY130_FD_SC_LS__A21OI_4%A_69_368# N_A_69_368#_M1002_d N_A_69_368#_M1003_d
+ N_A_69_368#_M1018_d N_A_69_368#_M1006_d N_A_69_368#_M1016_d
+ N_A_69_368#_M1007_s N_A_69_368#_M1017_s N_A_69_368#_c_332_n
+ N_A_69_368#_c_333_n N_A_69_368#_c_344_n N_A_69_368#_c_334_n
+ N_A_69_368#_c_352_n N_A_69_368#_c_356_n N_A_69_368#_c_358_n
+ N_A_69_368#_c_335_n N_A_69_368#_c_367_n N_A_69_368#_c_370_n
+ N_A_69_368#_c_372_n N_A_69_368#_c_373_n N_A_69_368#_c_336_n
+ N_A_69_368#_c_337_n N_A_69_368#_c_430_p N_A_69_368#_c_338_n
+ N_A_69_368#_c_339_n N_A_69_368#_c_361_n N_A_69_368#_c_365_n
+ N_A_69_368#_c_340_n N_A_69_368#_c_341_n PM_SKY130_FD_SC_LS__A21OI_4%A_69_368#
x_PM_SKY130_FD_SC_LS__A21OI_4%VPWR N_VPWR_M1002_s N_VPWR_M1005_s N_VPWR_M1000_s
+ N_VPWR_M1010_s N_VPWR_c_440_n N_VPWR_c_441_n N_VPWR_c_442_n N_VPWR_c_443_n
+ N_VPWR_c_444_n N_VPWR_c_445_n N_VPWR_c_446_n N_VPWR_c_447_n N_VPWR_c_448_n
+ VPWR N_VPWR_c_449_n N_VPWR_c_450_n N_VPWR_c_439_n N_VPWR_c_452_n
+ N_VPWR_c_453_n PM_SKY130_FD_SC_LS__A21OI_4%VPWR
x_PM_SKY130_FD_SC_LS__A21OI_4%Y N_Y_M1009_s N_Y_M1020_s N_Y_M1008_s N_Y_M1019_s
+ N_Y_M1004_d N_Y_M1011_d N_Y_c_537_n N_Y_c_542_n N_Y_c_525_n N_Y_c_526_n
+ N_Y_c_527_n N_Y_c_568_n N_Y_c_528_n N_Y_c_549_n N_Y_c_529_n N_Y_c_580_n Y Y Y
+ N_Y_c_557_n PM_SKY130_FD_SC_LS__A21OI_4%Y
x_PM_SKY130_FD_SC_LS__A21OI_4%A_84_74# N_A_84_74#_M1001_d N_A_84_74#_M1013_d
+ N_A_84_74#_M1015_d N_A_84_74#_M1012_d N_A_84_74#_M1021_d N_A_84_74#_c_626_n
+ N_A_84_74#_c_627_n N_A_84_74#_c_628_n N_A_84_74#_c_629_n N_A_84_74#_c_630_n
+ N_A_84_74#_c_631_n N_A_84_74#_c_632_n N_A_84_74#_c_633_n N_A_84_74#_c_634_n
+ N_A_84_74#_c_635_n N_A_84_74#_c_636_n PM_SKY130_FD_SC_LS__A21OI_4%A_84_74#
x_PM_SKY130_FD_SC_LS__A21OI_4%VGND N_VGND_M1001_s N_VGND_M1014_s N_VGND_M1008_d
+ N_VGND_c_698_n N_VGND_c_699_n N_VGND_c_700_n N_VGND_c_701_n N_VGND_c_702_n
+ N_VGND_c_703_n VGND N_VGND_c_704_n N_VGND_c_705_n N_VGND_c_706_n
+ N_VGND_c_707_n N_VGND_c_708_n PM_SKY130_FD_SC_LS__A21OI_4%VGND
cc_1 VNB N_A2_M1001_g 0.0318708f $X=-0.19 $Y=-0.245 $X2=0.76 $Y2=0.74
cc_2 VNB N_A2_M1013_g 0.0224899f $X=-0.19 $Y=-0.245 $X2=1.19 $Y2=0.74
cc_3 VNB N_A2_M1014_g 0.0224899f $X=-0.19 $Y=-0.245 $X2=1.62 $Y2=0.74
cc_4 VNB N_A2_M1015_g 0.0229394f $X=-0.19 $Y=-0.245 $X2=2.05 $Y2=0.74
cc_5 VNB A2 0.00342206f $X=-0.19 $Y=-0.245 $X2=2.075 $Y2=1.58
cc_6 VNB N_A2_c_99_n 0.081021f $X=-0.19 $Y=-0.245 $X2=2.045 $Y2=1.557
cc_7 VNB N_A1_M1009_g 0.0222136f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=2.4
cc_8 VNB N_A1_M1012_g 0.0221267f $X=-0.19 $Y=-0.245 $X2=1.145 $Y2=2.4
cc_9 VNB N_A1_M1020_g 0.022172f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=2.4
cc_10 VNB N_A1_M1021_g 0.030436f $X=-0.19 $Y=-0.245 $X2=2.045 $Y2=2.4
cc_11 VNB N_A1_c_184_n 0.0707007f $X=-0.19 $Y=-0.245 $X2=1.62 $Y2=1.557
cc_12 VNB N_A1_c_185_n 0.0024641f $X=-0.19 $Y=-0.245 $X2=1.97 $Y2=1.557
cc_13 VNB N_B1_M1008_g 0.0301827f $X=-0.19 $Y=-0.245 $X2=1.145 $Y2=2.4
cc_14 VNB N_B1_M1019_g 0.0318708f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=2.4
cc_15 VNB N_B1_c_269_n 0.0104672f $X=-0.19 $Y=-0.245 $X2=1.62 $Y2=1.35
cc_16 VNB N_B1_c_270_n 0.0629807f $X=-0.19 $Y=-0.245 $X2=1.62 $Y2=0.74
cc_17 VNB N_B1_c_271_n 0.0185831f $X=-0.19 $Y=-0.245 $X2=2.045 $Y2=2.4
cc_18 VNB N_B1_c_272_n 0.0024641f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=1.557
cc_19 VNB N_VPWR_c_439_n 0.263193f $X=-0.19 $Y=-0.245 $X2=2.16 $Y2=1.565
cc_20 VNB N_Y_c_525_n 0.0312951f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_Y_c_526_n 0.00857879f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_22 VNB N_Y_c_527_n 0.0138829f $X=-0.19 $Y=-0.245 $X2=2.075 $Y2=1.58
cc_23 VNB N_Y_c_528_n 0.0270834f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=1.515
cc_24 VNB N_Y_c_529_n 0.00215725f $X=-0.19 $Y=-0.245 $X2=1.97 $Y2=1.557
cc_25 VNB Y 9.59717e-19 $X=-0.19 $Y=-0.245 $X2=2.045 $Y2=1.557
cc_26 VNB Y 0.00160528f $X=-0.19 $Y=-0.245 $X2=2.05 $Y2=1.557
cc_27 VNB N_A_84_74#_c_626_n 0.0270834f $X=-0.19 $Y=-0.245 $X2=1.62 $Y2=1.35
cc_28 VNB N_A_84_74#_c_627_n 0.00326872f $X=-0.19 $Y=-0.245 $X2=1.62 $Y2=0.74
cc_29 VNB N_A_84_74#_c_628_n 0.0126777f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_84_74#_c_629_n 0.00178908f $X=-0.19 $Y=-0.245 $X2=2.045 $Y2=2.4
cc_31 VNB N_A_84_74#_c_630_n 0.00766679f $X=-0.19 $Y=-0.245 $X2=2.05 $Y2=0.74
cc_32 VNB N_A_84_74#_c_631_n 0.00237811f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_84_74#_c_632_n 0.00211517f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_84_74#_c_633_n 0.00199363f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_84_74#_c_634_n 0.00127131f $X=-0.19 $Y=-0.245 $X2=0.76 $Y2=1.557
cc_36 VNB N_A_84_74#_c_635_n 0.00202435f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=1.557
cc_37 VNB N_A_84_74#_c_636_n 0.00757932f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.557
cc_38 VNB N_VGND_c_698_n 0.00323505f $X=-0.19 $Y=-0.245 $X2=1.19 $Y2=0.74
cc_39 VNB N_VGND_c_699_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_700_n 0.00323505f $X=-0.19 $Y=-0.245 $X2=1.62 $Y2=1.35
cc_41 VNB N_VGND_c_701_n 0.00396467f $X=-0.19 $Y=-0.245 $X2=2.045 $Y2=1.765
cc_42 VNB N_VGND_c_702_n 0.0258237f $X=-0.19 $Y=-0.245 $X2=2.045 $Y2=2.4
cc_43 VNB N_VGND_c_703_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=2.05 $Y2=1.35
cc_44 VNB N_VGND_c_704_n 0.068654f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_705_n 0.0344157f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.557
cc_46 VNB N_VGND_c_706_n 0.383272f $X=-0.19 $Y=-0.245 $X2=1.62 $Y2=1.557
cc_47 VNB N_VGND_c_707_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=1.97 $Y2=1.515
cc_48 VNB N_VGND_c_708_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=1.565
cc_49 VPB N_A2_c_100_n 0.0199141f $X=-0.19 $Y=1.66 $X2=0.695 $Y2=1.765
cc_50 VPB N_A2_c_101_n 0.0155119f $X=-0.19 $Y=1.66 $X2=1.145 $Y2=1.765
cc_51 VPB N_A2_c_102_n 0.0155127f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.765
cc_52 VPB N_A2_c_103_n 0.0157789f $X=-0.19 $Y=1.66 $X2=2.045 $Y2=1.765
cc_53 VPB A2 0.0106654f $X=-0.19 $Y=1.66 $X2=2.075 $Y2=1.58
cc_54 VPB N_A2_c_99_n 0.0493136f $X=-0.19 $Y=1.66 $X2=2.045 $Y2=1.557
cc_55 VPB N_A1_c_186_n 0.015103f $X=-0.19 $Y=1.66 $X2=0.76 $Y2=0.74
cc_56 VPB N_A1_c_187_n 0.0155429f $X=-0.19 $Y=1.66 $X2=1.19 $Y2=0.74
cc_57 VPB N_A1_c_188_n 0.0155109f $X=-0.19 $Y=1.66 $X2=1.62 $Y2=0.74
cc_58 VPB N_A1_c_189_n 0.0152455f $X=-0.19 $Y=1.66 $X2=2.05 $Y2=0.74
cc_59 VPB N_A1_c_184_n 0.0465532f $X=-0.19 $Y=1.66 $X2=1.62 $Y2=1.557
cc_60 VPB N_A1_c_185_n 0.006683f $X=-0.19 $Y=1.66 $X2=1.97 $Y2=1.557
cc_61 VPB N_B1_c_273_n 0.0148631f $X=-0.19 $Y=1.66 $X2=0.695 $Y2=1.765
cc_62 VPB N_B1_c_274_n 0.014664f $X=-0.19 $Y=1.66 $X2=0.76 $Y2=1.35
cc_63 VPB N_B1_c_275_n 0.0147175f $X=-0.19 $Y=1.66 $X2=1.19 $Y2=1.35
cc_64 VPB N_B1_c_269_n 0.00694608f $X=-0.19 $Y=1.66 $X2=1.62 $Y2=1.35
cc_65 VPB N_B1_c_270_n 0.0327409f $X=-0.19 $Y=1.66 $X2=1.62 $Y2=0.74
cc_66 VPB N_B1_c_278_n 0.018444f $X=-0.19 $Y=1.66 $X2=1.62 $Y2=0.74
cc_67 VPB N_B1_c_271_n 0.00972066f $X=-0.19 $Y=1.66 $X2=2.045 $Y2=2.4
cc_68 VPB N_B1_c_272_n 0.00575485f $X=-0.19 $Y=1.66 $X2=0.95 $Y2=1.557
cc_69 VPB N_A_69_368#_c_332_n 0.0183334f $X=-0.19 $Y=1.66 $X2=2.045 $Y2=1.765
cc_70 VPB N_A_69_368#_c_333_n 0.0345863f $X=-0.19 $Y=1.66 $X2=2.045 $Y2=2.4
cc_71 VPB N_A_69_368#_c_334_n 0.00257348f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.58
cc_72 VPB N_A_69_368#_c_335_n 0.00216998f $X=-0.19 $Y=1.66 $X2=0.95 $Y2=1.515
cc_73 VPB N_A_69_368#_c_336_n 0.0030474f $X=-0.19 $Y=1.66 $X2=2.05 $Y2=1.557
cc_74 VPB N_A_69_368#_c_337_n 0.00171072f $X=-0.19 $Y=1.66 $X2=0.95 $Y2=1.565
cc_75 VPB N_A_69_368#_c_338_n 0.0124466f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_A_69_368#_c_339_n 0.051057f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_A_69_368#_c_340_n 0.00257417f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_A_69_368#_c_341_n 0.00123754f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_440_n 0.00571271f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.765
cc_80 VPB N_VPWR_c_441_n 0.00734662f $X=-0.19 $Y=1.66 $X2=1.62 $Y2=0.74
cc_81 VPB N_VPWR_c_442_n 0.00514362f $X=-0.19 $Y=1.66 $X2=2.045 $Y2=2.4
cc_82 VPB N_VPWR_c_443_n 0.0206041f $X=-0.19 $Y=1.66 $X2=2.05 $Y2=1.35
cc_83 VPB N_VPWR_c_444_n 0.00769929f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_84 VPB N_VPWR_c_445_n 0.0240735f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_446_n 0.00460249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_447_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0.695 $Y2=1.557
cc_87 VPB N_VPWR_c_448_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0.76 $Y2=1.557
cc_88 VPB N_VPWR_c_449_n 0.0185253f $X=-0.19 $Y=1.66 $X2=1.97 $Y2=1.515
cc_89 VPB N_VPWR_c_450_n 0.0621431f $X=-0.19 $Y=1.66 $X2=1.97 $Y2=1.565
cc_90 VPB N_VPWR_c_439_n 0.0975399f $X=-0.19 $Y=1.66 $X2=2.16 $Y2=1.565
cc_91 VPB N_VPWR_c_452_n 0.00460249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_453_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB Y 0.00116984f $X=-0.19 $Y=1.66 $X2=2.05 $Y2=1.557
cc_94 N_A2_M1015_g N_A1_M1009_g 0.0179032f $X=2.05 $Y=0.74 $X2=0 $Y2=0
cc_95 N_A2_c_103_n N_A1_c_186_n 0.0114143f $X=2.045 $Y=1.765 $X2=0 $Y2=0
cc_96 A2 N_A1_c_184_n 0.00390446f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_97 N_A2_c_99_n N_A1_c_184_n 0.0194052f $X=2.045 $Y=1.557 $X2=0 $Y2=0
cc_98 N_A2_c_100_n N_A_69_368#_c_332_n 0.00314968f $X=0.695 $Y=1.765 $X2=0 $Y2=0
cc_99 N_A2_c_100_n N_A_69_368#_c_333_n 0.00526798f $X=0.695 $Y=1.765 $X2=0 $Y2=0
cc_100 N_A2_c_100_n N_A_69_368#_c_344_n 0.017123f $X=0.695 $Y=1.765 $X2=0 $Y2=0
cc_101 N_A2_c_101_n N_A_69_368#_c_344_n 0.0120074f $X=1.145 $Y=1.765 $X2=0 $Y2=0
cc_102 A2 N_A_69_368#_c_344_n 0.0289213f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_103 N_A2_c_99_n N_A_69_368#_c_344_n 0.00130859f $X=2.045 $Y=1.557 $X2=0 $Y2=0
cc_104 N_A2_c_100_n N_A_69_368#_c_334_n 6.69308e-19 $X=0.695 $Y=1.765 $X2=0
+ $Y2=0
cc_105 N_A2_c_101_n N_A_69_368#_c_334_n 0.0105452f $X=1.145 $Y=1.765 $X2=0 $Y2=0
cc_106 N_A2_c_102_n N_A_69_368#_c_334_n 0.0103431f $X=1.595 $Y=1.765 $X2=0 $Y2=0
cc_107 N_A2_c_103_n N_A_69_368#_c_334_n 6.45594e-19 $X=2.045 $Y=1.765 $X2=0
+ $Y2=0
cc_108 N_A2_c_102_n N_A_69_368#_c_352_n 0.0119563f $X=1.595 $Y=1.765 $X2=0 $Y2=0
cc_109 N_A2_c_103_n N_A_69_368#_c_352_n 0.0120074f $X=2.045 $Y=1.765 $X2=0 $Y2=0
cc_110 A2 N_A_69_368#_c_352_n 0.0393875f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_111 N_A2_c_99_n N_A_69_368#_c_352_n 0.00130859f $X=2.045 $Y=1.557 $X2=0 $Y2=0
cc_112 N_A2_c_103_n N_A_69_368#_c_356_n 4.27055e-19 $X=2.045 $Y=1.765 $X2=0
+ $Y2=0
cc_113 A2 N_A_69_368#_c_356_n 0.012322f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_114 N_A2_c_102_n N_A_69_368#_c_358_n 4.35991e-19 $X=1.595 $Y=1.765 $X2=0
+ $Y2=0
cc_115 N_A2_c_103_n N_A_69_368#_c_358_n 0.00294319f $X=2.045 $Y=1.765 $X2=0
+ $Y2=0
cc_116 N_A2_c_103_n N_A_69_368#_c_335_n 0.00559111f $X=2.045 $Y=1.765 $X2=0
+ $Y2=0
cc_117 N_A2_c_101_n N_A_69_368#_c_361_n 4.27055e-19 $X=1.145 $Y=1.765 $X2=0
+ $Y2=0
cc_118 N_A2_c_102_n N_A_69_368#_c_361_n 4.27055e-19 $X=1.595 $Y=1.765 $X2=0
+ $Y2=0
cc_119 A2 N_A_69_368#_c_361_n 0.0237598f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_120 N_A2_c_99_n N_A_69_368#_c_361_n 0.00144162f $X=2.045 $Y=1.557 $X2=0 $Y2=0
cc_121 N_A2_c_103_n N_A_69_368#_c_365_n 0.0017329f $X=2.045 $Y=1.765 $X2=0 $Y2=0
cc_122 N_A2_c_100_n N_VPWR_c_440_n 0.0135832f $X=0.695 $Y=1.765 $X2=0 $Y2=0
cc_123 N_A2_c_101_n N_VPWR_c_440_n 0.00526215f $X=1.145 $Y=1.765 $X2=0 $Y2=0
cc_124 N_A2_c_102_n N_VPWR_c_441_n 0.00486623f $X=1.595 $Y=1.765 $X2=0 $Y2=0
cc_125 N_A2_c_103_n N_VPWR_c_441_n 0.00366463f $X=2.045 $Y=1.765 $X2=0 $Y2=0
cc_126 N_A2_c_103_n N_VPWR_c_442_n 4.52895e-19 $X=2.045 $Y=1.765 $X2=0 $Y2=0
cc_127 N_A2_c_100_n N_VPWR_c_445_n 0.00413917f $X=0.695 $Y=1.765 $X2=0 $Y2=0
cc_128 N_A2_c_101_n N_VPWR_c_447_n 0.00445602f $X=1.145 $Y=1.765 $X2=0 $Y2=0
cc_129 N_A2_c_102_n N_VPWR_c_447_n 0.00445602f $X=1.595 $Y=1.765 $X2=0 $Y2=0
cc_130 N_A2_c_103_n N_VPWR_c_449_n 0.00445602f $X=2.045 $Y=1.765 $X2=0 $Y2=0
cc_131 N_A2_c_100_n N_VPWR_c_439_n 0.00821701f $X=0.695 $Y=1.765 $X2=0 $Y2=0
cc_132 N_A2_c_101_n N_VPWR_c_439_n 0.00857589f $X=1.145 $Y=1.765 $X2=0 $Y2=0
cc_133 N_A2_c_102_n N_VPWR_c_439_n 0.00857589f $X=1.595 $Y=1.765 $X2=0 $Y2=0
cc_134 N_A2_c_103_n N_VPWR_c_439_n 0.00857673f $X=2.045 $Y=1.765 $X2=0 $Y2=0
cc_135 N_A2_c_103_n Y 8.01844e-19 $X=2.045 $Y=1.765 $X2=0 $Y2=0
cc_136 N_A2_M1015_g Y 8.33311e-19 $X=2.05 $Y=0.74 $X2=0 $Y2=0
cc_137 A2 Y 0.0263961f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_138 N_A2_c_99_n Y 3.58658e-19 $X=2.045 $Y=1.557 $X2=0 $Y2=0
cc_139 N_A2_M1001_g N_A_84_74#_c_626_n 0.00159319f $X=0.76 $Y=0.74 $X2=0 $Y2=0
cc_140 N_A2_M1001_g N_A_84_74#_c_627_n 0.0166797f $X=0.76 $Y=0.74 $X2=0 $Y2=0
cc_141 N_A2_M1013_g N_A_84_74#_c_627_n 0.0130918f $X=1.19 $Y=0.74 $X2=0 $Y2=0
cc_142 A2 N_A_84_74#_c_627_n 0.0402557f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_143 N_A2_c_99_n N_A_84_74#_c_627_n 0.00450756f $X=2.045 $Y=1.557 $X2=0 $Y2=0
cc_144 N_A2_c_99_n N_A_84_74#_c_628_n 0.00116678f $X=2.045 $Y=1.557 $X2=0 $Y2=0
cc_145 N_A2_M1013_g N_A_84_74#_c_629_n 3.92313e-19 $X=1.19 $Y=0.74 $X2=0 $Y2=0
cc_146 N_A2_M1014_g N_A_84_74#_c_629_n 3.92313e-19 $X=1.62 $Y=0.74 $X2=0 $Y2=0
cc_147 N_A2_M1014_g N_A_84_74#_c_630_n 0.0130453f $X=1.62 $Y=0.74 $X2=0 $Y2=0
cc_148 N_A2_M1015_g N_A_84_74#_c_630_n 0.0128967f $X=2.05 $Y=0.74 $X2=0 $Y2=0
cc_149 A2 N_A_84_74#_c_630_n 0.0604918f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_150 N_A2_c_99_n N_A_84_74#_c_630_n 0.00247712f $X=2.045 $Y=1.557 $X2=0 $Y2=0
cc_151 N_A2_M1015_g N_A_84_74#_c_632_n 9.48753e-19 $X=2.05 $Y=0.74 $X2=0 $Y2=0
cc_152 A2 N_A_84_74#_c_634_n 0.0146029f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_153 N_A2_c_99_n N_A_84_74#_c_634_n 0.00232957f $X=2.045 $Y=1.557 $X2=0 $Y2=0
cc_154 N_A2_M1001_g N_VGND_c_698_n 0.0133724f $X=0.76 $Y=0.74 $X2=0 $Y2=0
cc_155 N_A2_M1013_g N_VGND_c_698_n 0.0103289f $X=1.19 $Y=0.74 $X2=0 $Y2=0
cc_156 N_A2_M1014_g N_VGND_c_698_n 4.71636e-19 $X=1.62 $Y=0.74 $X2=0 $Y2=0
cc_157 N_A2_M1013_g N_VGND_c_699_n 0.00383152f $X=1.19 $Y=0.74 $X2=0 $Y2=0
cc_158 N_A2_M1014_g N_VGND_c_699_n 0.00383152f $X=1.62 $Y=0.74 $X2=0 $Y2=0
cc_159 N_A2_M1013_g N_VGND_c_700_n 4.71636e-19 $X=1.19 $Y=0.74 $X2=0 $Y2=0
cc_160 N_A2_M1014_g N_VGND_c_700_n 0.0103289f $X=1.62 $Y=0.74 $X2=0 $Y2=0
cc_161 N_A2_M1015_g N_VGND_c_700_n 0.00968343f $X=2.05 $Y=0.74 $X2=0 $Y2=0
cc_162 N_A2_M1001_g N_VGND_c_702_n 0.00383152f $X=0.76 $Y=0.74 $X2=0 $Y2=0
cc_163 N_A2_M1015_g N_VGND_c_704_n 0.00383152f $X=2.05 $Y=0.74 $X2=0 $Y2=0
cc_164 N_A2_M1001_g N_VGND_c_706_n 0.00761822f $X=0.76 $Y=0.74 $X2=0 $Y2=0
cc_165 N_A2_M1013_g N_VGND_c_706_n 0.0075754f $X=1.19 $Y=0.74 $X2=0 $Y2=0
cc_166 N_A2_M1014_g N_VGND_c_706_n 0.0075754f $X=1.62 $Y=0.74 $X2=0 $Y2=0
cc_167 N_A2_M1015_g N_VGND_c_706_n 0.00757637f $X=2.05 $Y=0.74 $X2=0 $Y2=0
cc_168 N_A1_c_189_n N_B1_c_273_n 0.0270425f $X=3.845 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_169 N_A1_c_184_n N_B1_c_270_n 0.0173183f $X=3.77 $Y=1.515 $X2=0 $Y2=0
cc_170 N_A1_c_185_n N_B1_c_270_n 7.08318e-19 $X=3.77 $Y=1.515 $X2=0 $Y2=0
cc_171 N_A1_c_184_n N_B1_c_272_n 5.21393e-19 $X=3.77 $Y=1.515 $X2=0 $Y2=0
cc_172 N_A1_c_185_n N_B1_c_272_n 0.0229482f $X=3.77 $Y=1.515 $X2=0 $Y2=0
cc_173 N_A1_c_186_n N_A_69_368#_c_335_n 0.00285725f $X=2.495 $Y=1.765 $X2=0
+ $Y2=0
cc_174 N_A1_c_186_n N_A_69_368#_c_367_n 0.0156331f $X=2.495 $Y=1.765 $X2=0 $Y2=0
cc_175 N_A1_c_187_n N_A_69_368#_c_367_n 0.011796f $X=2.945 $Y=1.765 $X2=0 $Y2=0
cc_176 N_A1_c_184_n N_A_69_368#_c_367_n 5.17185e-19 $X=3.77 $Y=1.515 $X2=0 $Y2=0
cc_177 N_A1_c_188_n N_A_69_368#_c_370_n 0.0117449f $X=3.395 $Y=1.765 $X2=0 $Y2=0
cc_178 N_A1_c_189_n N_A_69_368#_c_370_n 0.011796f $X=3.845 $Y=1.765 $X2=0 $Y2=0
cc_179 N_A1_c_189_n N_A_69_368#_c_372_n 4.27055e-19 $X=3.845 $Y=1.765 $X2=0
+ $Y2=0
cc_180 N_A1_c_188_n N_A_69_368#_c_373_n 5.42473e-19 $X=3.395 $Y=1.765 $X2=0
+ $Y2=0
cc_181 N_A1_c_189_n N_A_69_368#_c_373_n 0.00574124f $X=3.845 $Y=1.765 $X2=0
+ $Y2=0
cc_182 N_A1_c_189_n N_A_69_368#_c_337_n 0.0032261f $X=3.845 $Y=1.765 $X2=0 $Y2=0
cc_183 N_A1_c_186_n N_A_69_368#_c_340_n 5.8779e-19 $X=2.495 $Y=1.765 $X2=0 $Y2=0
cc_184 N_A1_c_187_n N_A_69_368#_c_340_n 0.00750758f $X=2.945 $Y=1.765 $X2=0
+ $Y2=0
cc_185 N_A1_c_188_n N_A_69_368#_c_340_n 0.00730551f $X=3.395 $Y=1.765 $X2=0
+ $Y2=0
cc_186 N_A1_c_189_n N_A_69_368#_c_340_n 5.64076e-19 $X=3.845 $Y=1.765 $X2=0
+ $Y2=0
cc_187 N_A1_c_186_n N_VPWR_c_442_n 0.00732722f $X=2.495 $Y=1.765 $X2=0 $Y2=0
cc_188 N_A1_c_187_n N_VPWR_c_442_n 0.00409001f $X=2.945 $Y=1.765 $X2=0 $Y2=0
cc_189 N_A1_c_187_n N_VPWR_c_443_n 0.00445602f $X=2.945 $Y=1.765 $X2=0 $Y2=0
cc_190 N_A1_c_188_n N_VPWR_c_443_n 0.00445602f $X=3.395 $Y=1.765 $X2=0 $Y2=0
cc_191 N_A1_c_188_n N_VPWR_c_444_n 0.00379374f $X=3.395 $Y=1.765 $X2=0 $Y2=0
cc_192 N_A1_c_189_n N_VPWR_c_444_n 0.00224402f $X=3.845 $Y=1.765 $X2=0 $Y2=0
cc_193 N_A1_c_186_n N_VPWR_c_449_n 0.00413917f $X=2.495 $Y=1.765 $X2=0 $Y2=0
cc_194 N_A1_c_189_n N_VPWR_c_450_n 0.0044313f $X=3.845 $Y=1.765 $X2=0 $Y2=0
cc_195 N_A1_c_186_n N_VPWR_c_439_n 0.0081781f $X=2.495 $Y=1.765 $X2=0 $Y2=0
cc_196 N_A1_c_187_n N_VPWR_c_439_n 0.00857589f $X=2.945 $Y=1.765 $X2=0 $Y2=0
cc_197 N_A1_c_188_n N_VPWR_c_439_n 0.00857589f $X=3.395 $Y=1.765 $X2=0 $Y2=0
cc_198 N_A1_c_189_n N_VPWR_c_439_n 0.00853445f $X=3.845 $Y=1.765 $X2=0 $Y2=0
cc_199 N_A1_c_187_n N_Y_c_537_n 0.0124117f $X=2.945 $Y=1.765 $X2=0 $Y2=0
cc_200 N_A1_c_188_n N_Y_c_537_n 0.0107319f $X=3.395 $Y=1.765 $X2=0 $Y2=0
cc_201 N_A1_c_189_n N_Y_c_537_n 0.0106809f $X=3.845 $Y=1.765 $X2=0 $Y2=0
cc_202 N_A1_c_184_n N_Y_c_537_n 0.0056763f $X=3.77 $Y=1.515 $X2=0 $Y2=0
cc_203 N_A1_c_185_n N_Y_c_537_n 0.0689808f $X=3.77 $Y=1.515 $X2=0 $Y2=0
cc_204 N_A1_c_186_n N_Y_c_542_n 0.00476412f $X=2.495 $Y=1.765 $X2=0 $Y2=0
cc_205 N_A1_M1012_g N_Y_c_525_n 0.0175675f $X=2.91 $Y=0.74 $X2=0 $Y2=0
cc_206 N_A1_M1020_g N_Y_c_525_n 0.0139916f $X=3.34 $Y=0.74 $X2=0 $Y2=0
cc_207 N_A1_M1021_g N_Y_c_525_n 0.0176112f $X=3.77 $Y=0.74 $X2=0 $Y2=0
cc_208 N_A1_c_184_n N_Y_c_525_n 0.0069026f $X=3.77 $Y=1.515 $X2=0 $Y2=0
cc_209 N_A1_c_185_n N_Y_c_525_n 0.0794462f $X=3.77 $Y=1.515 $X2=0 $Y2=0
cc_210 N_A1_M1021_g N_Y_c_526_n 0.00455139f $X=3.77 $Y=0.74 $X2=0 $Y2=0
cc_211 N_A1_c_189_n N_Y_c_549_n 7.3898e-19 $X=3.845 $Y=1.765 $X2=0 $Y2=0
cc_212 N_A1_M1009_g Y 0.00466718f $X=2.48 $Y=0.74 $X2=0 $Y2=0
cc_213 N_A1_M1009_g Y 0.00447162f $X=2.48 $Y=0.74 $X2=0 $Y2=0
cc_214 N_A1_c_186_n Y 0.0050736f $X=2.495 $Y=1.765 $X2=0 $Y2=0
cc_215 N_A1_M1012_g Y 0.00414079f $X=2.91 $Y=0.74 $X2=0 $Y2=0
cc_216 N_A1_c_187_n Y 0.00411977f $X=2.945 $Y=1.765 $X2=0 $Y2=0
cc_217 N_A1_c_184_n Y 0.0237693f $X=3.77 $Y=1.515 $X2=0 $Y2=0
cc_218 N_A1_c_185_n Y 0.0336392f $X=3.77 $Y=1.515 $X2=0 $Y2=0
cc_219 N_A1_M1009_g N_Y_c_557_n 0.0040538f $X=2.48 $Y=0.74 $X2=0 $Y2=0
cc_220 N_A1_M1009_g N_A_84_74#_c_630_n 5.67309e-19 $X=2.48 $Y=0.74 $X2=0 $Y2=0
cc_221 N_A1_M1009_g N_A_84_74#_c_631_n 0.0118512f $X=2.48 $Y=0.74 $X2=0 $Y2=0
cc_222 N_A1_M1012_g N_A_84_74#_c_631_n 0.00799819f $X=2.91 $Y=0.74 $X2=0 $Y2=0
cc_223 N_A1_M1020_g N_A_84_74#_c_633_n 0.00804476f $X=3.34 $Y=0.74 $X2=0 $Y2=0
cc_224 N_A1_M1021_g N_A_84_74#_c_633_n 0.00807644f $X=3.77 $Y=0.74 $X2=0 $Y2=0
cc_225 N_A1_M1009_g N_A_84_74#_c_635_n 6.64397e-19 $X=2.48 $Y=0.74 $X2=0 $Y2=0
cc_226 N_A1_M1012_g N_A_84_74#_c_635_n 0.00704884f $X=2.91 $Y=0.74 $X2=0 $Y2=0
cc_227 N_A1_M1020_g N_A_84_74#_c_635_n 0.00766985f $X=3.34 $Y=0.74 $X2=0 $Y2=0
cc_228 N_A1_M1021_g N_A_84_74#_c_635_n 9.18514e-19 $X=3.77 $Y=0.74 $X2=0 $Y2=0
cc_229 N_A1_M1020_g N_A_84_74#_c_636_n 9.18514e-19 $X=3.34 $Y=0.74 $X2=0 $Y2=0
cc_230 N_A1_M1021_g N_A_84_74#_c_636_n 0.00862162f $X=3.77 $Y=0.74 $X2=0 $Y2=0
cc_231 N_A1_M1009_g N_VGND_c_704_n 0.00278271f $X=2.48 $Y=0.74 $X2=0 $Y2=0
cc_232 N_A1_M1012_g N_VGND_c_704_n 0.00279469f $X=2.91 $Y=0.74 $X2=0 $Y2=0
cc_233 N_A1_M1020_g N_VGND_c_704_n 0.00279469f $X=3.34 $Y=0.74 $X2=0 $Y2=0
cc_234 N_A1_M1021_g N_VGND_c_704_n 0.00279469f $X=3.77 $Y=0.74 $X2=0 $Y2=0
cc_235 N_A1_M1009_g N_VGND_c_706_n 0.00353526f $X=2.48 $Y=0.74 $X2=0 $Y2=0
cc_236 N_A1_M1012_g N_VGND_c_706_n 0.00352518f $X=2.91 $Y=0.74 $X2=0 $Y2=0
cc_237 N_A1_M1020_g N_VGND_c_706_n 0.00352518f $X=3.34 $Y=0.74 $X2=0 $Y2=0
cc_238 N_A1_M1021_g N_VGND_c_706_n 0.00357517f $X=3.77 $Y=0.74 $X2=0 $Y2=0
cc_239 N_B1_c_273_n N_A_69_368#_c_336_n 0.0128006f $X=4.295 $Y=1.765 $X2=0 $Y2=0
cc_240 N_B1_c_274_n N_A_69_368#_c_336_n 0.0128349f $X=4.745 $Y=1.765 $X2=0 $Y2=0
cc_241 N_B1_c_275_n N_A_69_368#_c_338_n 0.0128349f $X=5.195 $Y=1.765 $X2=0 $Y2=0
cc_242 N_B1_c_278_n N_A_69_368#_c_338_n 0.0137046f $X=5.645 $Y=1.765 $X2=0 $Y2=0
cc_243 N_B1_c_278_n N_A_69_368#_c_339_n 0.010383f $X=5.645 $Y=1.765 $X2=0 $Y2=0
cc_244 N_B1_c_273_n N_VPWR_c_450_n 0.00278271f $X=4.295 $Y=1.765 $X2=0 $Y2=0
cc_245 N_B1_c_274_n N_VPWR_c_450_n 0.00278271f $X=4.745 $Y=1.765 $X2=0 $Y2=0
cc_246 N_B1_c_275_n N_VPWR_c_450_n 0.00278271f $X=5.195 $Y=1.765 $X2=0 $Y2=0
cc_247 N_B1_c_278_n N_VPWR_c_450_n 0.00278271f $X=5.645 $Y=1.765 $X2=0 $Y2=0
cc_248 N_B1_c_273_n N_VPWR_c_439_n 0.00353907f $X=4.295 $Y=1.765 $X2=0 $Y2=0
cc_249 N_B1_c_274_n N_VPWR_c_439_n 0.00353823f $X=4.745 $Y=1.765 $X2=0 $Y2=0
cc_250 N_B1_c_275_n N_VPWR_c_439_n 0.00353823f $X=5.195 $Y=1.765 $X2=0 $Y2=0
cc_251 N_B1_c_278_n N_VPWR_c_439_n 0.00357579f $X=5.645 $Y=1.765 $X2=0 $Y2=0
cc_252 N_B1_c_273_n N_Y_c_537_n 0.0123471f $X=4.295 $Y=1.765 $X2=0 $Y2=0
cc_253 N_B1_c_272_n N_Y_c_537_n 0.00872169f $X=5.08 $Y=1.515 $X2=0 $Y2=0
cc_254 N_B1_c_270_n N_Y_c_525_n 0.00476181f $X=5.285 $Y=1.605 $X2=0 $Y2=0
cc_255 N_B1_c_272_n N_Y_c_525_n 0.0131745f $X=5.08 $Y=1.515 $X2=0 $Y2=0
cc_256 N_B1_M1008_g N_Y_c_526_n 0.00159319f $X=4.78 $Y=0.74 $X2=0 $Y2=0
cc_257 N_B1_M1008_g N_Y_c_527_n 0.0139178f $X=4.78 $Y=0.74 $X2=0 $Y2=0
cc_258 N_B1_M1019_g N_Y_c_527_n 0.0148472f $X=5.21 $Y=0.74 $X2=0 $Y2=0
cc_259 N_B1_c_269_n N_Y_c_527_n 0.0101416f $X=5.555 $Y=1.605 $X2=0 $Y2=0
cc_260 N_B1_c_270_n N_Y_c_527_n 0.00362717f $X=5.285 $Y=1.605 $X2=0 $Y2=0
cc_261 N_B1_c_272_n N_Y_c_527_n 0.0446327f $X=5.08 $Y=1.515 $X2=0 $Y2=0
cc_262 N_B1_c_274_n N_Y_c_568_n 0.0120074f $X=4.745 $Y=1.765 $X2=0 $Y2=0
cc_263 N_B1_c_275_n N_Y_c_568_n 0.0122823f $X=5.195 $Y=1.765 $X2=0 $Y2=0
cc_264 N_B1_c_270_n N_Y_c_568_n 0.00130859f $X=5.285 $Y=1.605 $X2=0 $Y2=0
cc_265 N_B1_c_272_n N_Y_c_568_n 0.0386917f $X=5.08 $Y=1.515 $X2=0 $Y2=0
cc_266 N_B1_M1019_g N_Y_c_528_n 0.00159319f $X=5.21 $Y=0.74 $X2=0 $Y2=0
cc_267 N_B1_c_273_n N_Y_c_549_n 0.0089645f $X=4.295 $Y=1.765 $X2=0 $Y2=0
cc_268 N_B1_c_274_n N_Y_c_549_n 0.00891808f $X=4.745 $Y=1.765 $X2=0 $Y2=0
cc_269 N_B1_c_275_n N_Y_c_549_n 5.7112e-19 $X=5.195 $Y=1.765 $X2=0 $Y2=0
cc_270 N_B1_c_270_n N_Y_c_549_n 0.00145364f $X=5.285 $Y=1.605 $X2=0 $Y2=0
cc_271 N_B1_c_272_n N_Y_c_549_n 0.0237598f $X=5.08 $Y=1.515 $X2=0 $Y2=0
cc_272 N_B1_c_270_n N_Y_c_529_n 0.00582391f $X=5.285 $Y=1.605 $X2=0 $Y2=0
cc_273 N_B1_c_272_n N_Y_c_529_n 0.0214728f $X=5.08 $Y=1.515 $X2=0 $Y2=0
cc_274 N_B1_c_274_n N_Y_c_580_n 5.7112e-19 $X=4.745 $Y=1.765 $X2=0 $Y2=0
cc_275 N_B1_c_275_n N_Y_c_580_n 0.00944195f $X=5.195 $Y=1.765 $X2=0 $Y2=0
cc_276 N_B1_c_269_n N_Y_c_580_n 0.00811534f $X=5.555 $Y=1.605 $X2=0 $Y2=0
cc_277 N_B1_c_278_n N_Y_c_580_n 0.0101179f $X=5.645 $Y=1.765 $X2=0 $Y2=0
cc_278 N_B1_M1008_g N_A_84_74#_c_636_n 0.00301154f $X=4.78 $Y=0.74 $X2=0 $Y2=0
cc_279 N_B1_M1008_g N_VGND_c_701_n 0.0133724f $X=4.78 $Y=0.74 $X2=0 $Y2=0
cc_280 N_B1_M1019_g N_VGND_c_701_n 0.0133724f $X=5.21 $Y=0.74 $X2=0 $Y2=0
cc_281 N_B1_M1008_g N_VGND_c_704_n 0.00383152f $X=4.78 $Y=0.74 $X2=0 $Y2=0
cc_282 N_B1_M1019_g N_VGND_c_705_n 0.00383152f $X=5.21 $Y=0.74 $X2=0 $Y2=0
cc_283 N_B1_M1008_g N_VGND_c_706_n 0.00762539f $X=4.78 $Y=0.74 $X2=0 $Y2=0
cc_284 N_B1_M1019_g N_VGND_c_706_n 0.00762539f $X=5.21 $Y=0.74 $X2=0 $Y2=0
cc_285 N_A_69_368#_c_344_n N_VPWR_M1002_s 0.00384138f $X=1.205 $Y=2.035
+ $X2=-0.19 $Y2=1.66
cc_286 N_A_69_368#_c_352_n N_VPWR_M1005_s 0.00408911f $X=2.105 $Y=2.035 $X2=0
+ $Y2=0
cc_287 N_A_69_368#_c_367_n N_VPWR_M1000_s 0.00402919f $X=3.005 $Y=2.375 $X2=0
+ $Y2=0
cc_288 N_A_69_368#_c_370_n N_VPWR_M1010_s 0.00428955f $X=3.905 $Y=2.375 $X2=0
+ $Y2=0
cc_289 N_A_69_368#_c_333_n N_VPWR_c_440_n 0.0453479f $X=0.47 $Y=2.4 $X2=0 $Y2=0
cc_290 N_A_69_368#_c_344_n N_VPWR_c_440_n 0.0154248f $X=1.205 $Y=2.035 $X2=0
+ $Y2=0
cc_291 N_A_69_368#_c_334_n N_VPWR_c_440_n 0.0462948f $X=1.37 $Y=2.815 $X2=0
+ $Y2=0
cc_292 N_A_69_368#_c_334_n N_VPWR_c_441_n 0.0449718f $X=1.37 $Y=2.815 $X2=0
+ $Y2=0
cc_293 N_A_69_368#_c_352_n N_VPWR_c_441_n 0.0136682f $X=2.105 $Y=2.035 $X2=0
+ $Y2=0
cc_294 N_A_69_368#_c_335_n N_VPWR_c_441_n 0.0331533f $X=2.27 $Y=2.465 $X2=0
+ $Y2=0
cc_295 N_A_69_368#_c_365_n N_VPWR_c_441_n 0.0117758f $X=2.23 $Y=2.375 $X2=0
+ $Y2=0
cc_296 N_A_69_368#_c_335_n N_VPWR_c_442_n 0.0230171f $X=2.27 $Y=2.465 $X2=0
+ $Y2=0
cc_297 N_A_69_368#_c_367_n N_VPWR_c_442_n 0.0154248f $X=3.005 $Y=2.375 $X2=0
+ $Y2=0
cc_298 N_A_69_368#_c_340_n N_VPWR_c_442_n 0.0234974f $X=3.17 $Y=2.455 $X2=0
+ $Y2=0
cc_299 N_A_69_368#_c_340_n N_VPWR_c_443_n 0.0145674f $X=3.17 $Y=2.455 $X2=0
+ $Y2=0
cc_300 N_A_69_368#_c_370_n N_VPWR_c_444_n 0.0136682f $X=3.905 $Y=2.375 $X2=0
+ $Y2=0
cc_301 N_A_69_368#_c_373_n N_VPWR_c_444_n 0.0175037f $X=4.03 $Y=2.905 $X2=0
+ $Y2=0
cc_302 N_A_69_368#_c_337_n N_VPWR_c_444_n 0.0119328f $X=4.155 $Y=2.99 $X2=0
+ $Y2=0
cc_303 N_A_69_368#_c_340_n N_VPWR_c_444_n 0.0228252f $X=3.17 $Y=2.455 $X2=0
+ $Y2=0
cc_304 N_A_69_368#_c_333_n N_VPWR_c_445_n 0.011066f $X=0.47 $Y=2.4 $X2=0 $Y2=0
cc_305 N_A_69_368#_c_334_n N_VPWR_c_447_n 0.014552f $X=1.37 $Y=2.815 $X2=0 $Y2=0
cc_306 N_A_69_368#_c_335_n N_VPWR_c_449_n 0.0110241f $X=2.27 $Y=2.465 $X2=0
+ $Y2=0
cc_307 N_A_69_368#_c_336_n N_VPWR_c_450_n 0.0460938f $X=4.885 $Y=2.99 $X2=0
+ $Y2=0
cc_308 N_A_69_368#_c_337_n N_VPWR_c_450_n 0.017869f $X=4.155 $Y=2.99 $X2=0 $Y2=0
cc_309 N_A_69_368#_c_338_n N_VPWR_c_450_n 0.0640155f $X=5.785 $Y=2.99 $X2=0
+ $Y2=0
cc_310 N_A_69_368#_c_341_n N_VPWR_c_450_n 0.0121867f $X=4.97 $Y=2.99 $X2=0 $Y2=0
cc_311 N_A_69_368#_c_333_n N_VPWR_c_439_n 0.00915947f $X=0.47 $Y=2.4 $X2=0 $Y2=0
cc_312 N_A_69_368#_c_334_n N_VPWR_c_439_n 0.0119791f $X=1.37 $Y=2.815 $X2=0
+ $Y2=0
cc_313 N_A_69_368#_c_335_n N_VPWR_c_439_n 0.00909194f $X=2.27 $Y=2.465 $X2=0
+ $Y2=0
cc_314 N_A_69_368#_c_336_n N_VPWR_c_439_n 0.0260732f $X=4.885 $Y=2.99 $X2=0
+ $Y2=0
cc_315 N_A_69_368#_c_337_n N_VPWR_c_439_n 0.00965079f $X=4.155 $Y=2.99 $X2=0
+ $Y2=0
cc_316 N_A_69_368#_c_338_n N_VPWR_c_439_n 0.0357926f $X=5.785 $Y=2.99 $X2=0
+ $Y2=0
cc_317 N_A_69_368#_c_340_n N_VPWR_c_439_n 0.0119851f $X=3.17 $Y=2.455 $X2=0
+ $Y2=0
cc_318 N_A_69_368#_c_341_n N_VPWR_c_439_n 0.00660921f $X=4.97 $Y=2.99 $X2=0
+ $Y2=0
cc_319 N_A_69_368#_c_336_n N_Y_M1004_d 0.00197722f $X=4.885 $Y=2.99 $X2=0 $Y2=0
cc_320 N_A_69_368#_c_338_n N_Y_M1011_d 0.00197722f $X=5.785 $Y=2.99 $X2=0 $Y2=0
cc_321 N_A_69_368#_M1006_d N_Y_c_537_n 0.00359365f $X=3.02 $Y=1.84 $X2=0 $Y2=0
cc_322 N_A_69_368#_M1016_d N_Y_c_537_n 0.00929435f $X=3.92 $Y=1.84 $X2=0 $Y2=0
cc_323 N_A_69_368#_c_367_n N_Y_c_537_n 0.0132929f $X=3.005 $Y=2.375 $X2=0 $Y2=0
cc_324 N_A_69_368#_c_370_n N_Y_c_537_n 0.0317427f $X=3.905 $Y=2.375 $X2=0 $Y2=0
cc_325 N_A_69_368#_c_372_n N_Y_c_537_n 0.0155823f $X=4.03 $Y=2.46 $X2=0 $Y2=0
cc_326 N_A_69_368#_c_340_n N_Y_c_537_n 0.0173542f $X=3.17 $Y=2.455 $X2=0 $Y2=0
cc_327 N_A_69_368#_c_356_n N_Y_c_542_n 0.0148585f $X=2.23 $Y=2.12 $X2=0 $Y2=0
cc_328 N_A_69_368#_c_367_n N_Y_c_542_n 0.0137548f $X=3.005 $Y=2.375 $X2=0 $Y2=0
cc_329 N_A_69_368#_M1007_s N_Y_c_568_n 0.00408911f $X=4.82 $Y=1.84 $X2=0 $Y2=0
cc_330 N_A_69_368#_c_430_p N_Y_c_568_n 0.0136682f $X=4.97 $Y=2.455 $X2=0 $Y2=0
cc_331 N_A_69_368#_c_372_n N_Y_c_549_n 0.0123817f $X=4.03 $Y=2.46 $X2=0 $Y2=0
cc_332 N_A_69_368#_c_373_n N_Y_c_549_n 0.0184049f $X=4.03 $Y=2.905 $X2=0 $Y2=0
cc_333 N_A_69_368#_c_336_n N_Y_c_549_n 0.0160777f $X=4.885 $Y=2.99 $X2=0 $Y2=0
cc_334 N_A_69_368#_c_430_p N_Y_c_549_n 0.0289859f $X=4.97 $Y=2.455 $X2=0 $Y2=0
cc_335 N_A_69_368#_c_430_p N_Y_c_580_n 0.0289859f $X=4.97 $Y=2.455 $X2=0 $Y2=0
cc_336 N_A_69_368#_c_338_n N_Y_c_580_n 0.0160777f $X=5.785 $Y=2.99 $X2=0 $Y2=0
cc_337 N_A_69_368#_c_339_n N_Y_c_580_n 0.0533059f $X=5.87 $Y=1.985 $X2=0 $Y2=0
cc_338 N_A_69_368#_c_332_n N_A_84_74#_c_628_n 0.00646892f $X=0.43 $Y=2.12 $X2=0
+ $Y2=0
cc_339 N_VPWR_M1000_s N_Y_c_537_n 0.00132153f $X=2.57 $Y=1.84 $X2=0 $Y2=0
cc_340 N_VPWR_M1010_s N_Y_c_537_n 0.00359847f $X=3.47 $Y=1.84 $X2=0 $Y2=0
cc_341 N_VPWR_M1000_s N_Y_c_542_n 0.00140887f $X=2.57 $Y=1.84 $X2=0 $Y2=0
cc_342 N_VPWR_M1000_s Y 0.00127015f $X=2.57 $Y=1.84 $X2=0 $Y2=0
cc_343 N_Y_c_525_n N_A_84_74#_M1012_d 0.00179574f $X=4.4 $Y=1.03 $X2=0 $Y2=0
cc_344 N_Y_c_525_n N_A_84_74#_M1021_d 0.00379734f $X=4.4 $Y=1.03 $X2=0 $Y2=0
cc_345 Y N_A_84_74#_c_630_n 0.0101919f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_346 N_Y_M1009_s N_A_84_74#_c_631_n 0.00176461f $X=2.555 $Y=0.37 $X2=0 $Y2=0
cc_347 N_Y_c_525_n N_A_84_74#_c_631_n 0.00397126f $X=4.4 $Y=1.03 $X2=0 $Y2=0
cc_348 N_Y_c_557_n N_A_84_74#_c_631_n 0.0146809f $X=2.652 $Y=0.88 $X2=0 $Y2=0
cc_349 N_Y_M1020_s N_A_84_74#_c_633_n 0.00285125f $X=3.415 $Y=0.37 $X2=0 $Y2=0
cc_350 N_Y_c_525_n N_A_84_74#_c_633_n 0.0140305f $X=4.4 $Y=1.03 $X2=0 $Y2=0
cc_351 N_Y_c_525_n N_A_84_74#_c_635_n 0.0172179f $X=4.4 $Y=1.03 $X2=0 $Y2=0
cc_352 N_Y_c_525_n N_A_84_74#_c_636_n 0.0221161f $X=4.4 $Y=1.03 $X2=0 $Y2=0
cc_353 N_Y_c_526_n N_A_84_74#_c_636_n 0.0224421f $X=4.565 $Y=0.515 $X2=0 $Y2=0
cc_354 N_Y_c_527_n N_VGND_M1008_d 0.00176461f $X=5.34 $Y=1.095 $X2=0 $Y2=0
cc_355 N_Y_c_526_n N_VGND_c_701_n 0.0182902f $X=4.565 $Y=0.515 $X2=0 $Y2=0
cc_356 N_Y_c_527_n N_VGND_c_701_n 0.0171619f $X=5.34 $Y=1.095 $X2=0 $Y2=0
cc_357 N_Y_c_528_n N_VGND_c_701_n 0.0182902f $X=5.425 $Y=0.515 $X2=0 $Y2=0
cc_358 N_Y_c_526_n N_VGND_c_704_n 0.011066f $X=4.565 $Y=0.515 $X2=0 $Y2=0
cc_359 N_Y_c_528_n N_VGND_c_705_n 0.011066f $X=5.425 $Y=0.515 $X2=0 $Y2=0
cc_360 N_Y_c_526_n N_VGND_c_706_n 0.00915947f $X=4.565 $Y=0.515 $X2=0 $Y2=0
cc_361 N_Y_c_528_n N_VGND_c_706_n 0.00915947f $X=5.425 $Y=0.515 $X2=0 $Y2=0
cc_362 N_A_84_74#_c_627_n N_VGND_M1001_s 0.00176461f $X=1.32 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_363 N_A_84_74#_c_630_n N_VGND_M1014_s 0.00176461f $X=2.18 $Y=1.095 $X2=0
+ $Y2=0
cc_364 N_A_84_74#_c_626_n N_VGND_c_698_n 0.0182902f $X=0.545 $Y=0.515 $X2=0
+ $Y2=0
cc_365 N_A_84_74#_c_627_n N_VGND_c_698_n 0.0171619f $X=1.32 $Y=1.095 $X2=0 $Y2=0
cc_366 N_A_84_74#_c_629_n N_VGND_c_698_n 0.0182488f $X=1.405 $Y=0.515 $X2=0
+ $Y2=0
cc_367 N_A_84_74#_c_629_n N_VGND_c_699_n 0.00749631f $X=1.405 $Y=0.515 $X2=0
+ $Y2=0
cc_368 N_A_84_74#_c_629_n N_VGND_c_700_n 0.0182488f $X=1.405 $Y=0.515 $X2=0
+ $Y2=0
cc_369 N_A_84_74#_c_630_n N_VGND_c_700_n 0.0171619f $X=2.18 $Y=1.095 $X2=0 $Y2=0
cc_370 N_A_84_74#_c_632_n N_VGND_c_700_n 0.0112234f $X=2.35 $Y=0.34 $X2=0 $Y2=0
cc_371 N_A_84_74#_c_626_n N_VGND_c_702_n 0.011066f $X=0.545 $Y=0.515 $X2=0 $Y2=0
cc_372 N_A_84_74#_c_631_n N_VGND_c_704_n 0.0384655f $X=2.96 $Y=0.34 $X2=0 $Y2=0
cc_373 N_A_84_74#_c_632_n N_VGND_c_704_n 0.0121867f $X=2.35 $Y=0.34 $X2=0 $Y2=0
cc_374 N_A_84_74#_c_633_n N_VGND_c_704_n 0.033414f $X=3.82 $Y=0.34 $X2=0 $Y2=0
cc_375 N_A_84_74#_c_635_n N_VGND_c_704_n 0.0226572f $X=3.125 $Y=0.34 $X2=0 $Y2=0
cc_376 N_A_84_74#_c_636_n N_VGND_c_704_n 0.0227371f $X=3.985 $Y=0.34 $X2=0 $Y2=0
cc_377 N_A_84_74#_c_626_n N_VGND_c_706_n 0.00915947f $X=0.545 $Y=0.515 $X2=0
+ $Y2=0
cc_378 N_A_84_74#_c_629_n N_VGND_c_706_n 0.0062048f $X=1.405 $Y=0.515 $X2=0
+ $Y2=0
cc_379 N_A_84_74#_c_631_n N_VGND_c_706_n 0.0216792f $X=2.96 $Y=0.34 $X2=0 $Y2=0
cc_380 N_A_84_74#_c_632_n N_VGND_c_706_n 0.00660921f $X=2.35 $Y=0.34 $X2=0 $Y2=0
cc_381 N_A_84_74#_c_633_n N_VGND_c_706_n 0.0187892f $X=3.82 $Y=0.34 $X2=0 $Y2=0
cc_382 N_A_84_74#_c_635_n N_VGND_c_706_n 0.0124022f $X=3.125 $Y=0.34 $X2=0 $Y2=0
cc_383 N_A_84_74#_c_636_n N_VGND_c_706_n 0.0125119f $X=3.985 $Y=0.34 $X2=0 $Y2=0
