# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ls__sdfbbp_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ls__sdfbbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  15.84000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.455000 1.525000 1.765000 1.855000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.530100 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 15.395000 0.350000 15.735000 2.980000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.518900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.770000 0.350000 14.275000 1.050000 ;
        RECT 13.870000 1.720000 14.275000 2.890000 ;
        RECT 14.105000 1.050000 14.275000 1.720000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.065000 1.180000 13.360000 1.550000 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.125000 0.550000 2.135000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.805000 1.550000 1.285000 2.095000 ;
    END
  END SCE
  PIN SET_B
    ANTENNAGATEAREA  0.469500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  7.045000 1.410000  7.375000 1.655000 ;
        RECT  7.095000 1.655000  7.265000 2.905000 ;
        RECT  7.095000 2.905000  8.105000 3.075000 ;
        RECT  7.935000 2.165000  9.025000 2.335000 ;
        RECT  7.935000 2.335000  8.105000 2.905000 ;
        RECT  8.855000 2.335000  9.025000 2.905000 ;
        RECT  8.855000 2.905000 10.265000 3.075000 ;
        RECT 10.095000 2.015000 10.295000 2.185000 ;
        RECT 10.095000 2.185000 10.265000 2.905000 ;
        RECT 10.125000 1.690000 11.385000 1.800000 ;
        RECT 10.125000 1.800000 11.365000 1.860000 ;
        RECT 10.125000 1.860000 10.295000 2.015000 ;
        RECT 11.055000 1.520000 11.385000 1.690000 ;
        RECT 11.055000 1.860000 11.365000 2.150000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.430000 1.180000 3.760000 1.670000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 15.840000 0.085000 ;
        RECT  0.140000  0.085000  0.470000 0.955000 ;
        RECT  1.830000  0.085000  2.080000 1.015000 ;
        RECT  3.850000  0.085000  4.180000 0.490000 ;
        RECT  6.490000  0.085000  6.885000 0.560000 ;
        RECT  9.025000  0.085000  9.275000 1.050000 ;
        RECT 10.900000  0.085000 11.150000 1.010000 ;
        RECT 13.295000  0.085000 13.590000 1.000000 ;
        RECT 14.895000  0.085000 15.225000 0.940000 ;
      LAYER mcon ;
        RECT  0.155000 -0.085000  0.325000 0.085000 ;
        RECT  0.635000 -0.085000  0.805000 0.085000 ;
        RECT  1.115000 -0.085000  1.285000 0.085000 ;
        RECT  1.595000 -0.085000  1.765000 0.085000 ;
        RECT  2.075000 -0.085000  2.245000 0.085000 ;
        RECT  2.555000 -0.085000  2.725000 0.085000 ;
        RECT  3.035000 -0.085000  3.205000 0.085000 ;
        RECT  3.515000 -0.085000  3.685000 0.085000 ;
        RECT  3.995000 -0.085000  4.165000 0.085000 ;
        RECT  4.475000 -0.085000  4.645000 0.085000 ;
        RECT  4.955000 -0.085000  5.125000 0.085000 ;
        RECT  5.435000 -0.085000  5.605000 0.085000 ;
        RECT  5.915000 -0.085000  6.085000 0.085000 ;
        RECT  6.395000 -0.085000  6.565000 0.085000 ;
        RECT  6.875000 -0.085000  7.045000 0.085000 ;
        RECT  7.355000 -0.085000  7.525000 0.085000 ;
        RECT  7.835000 -0.085000  8.005000 0.085000 ;
        RECT  8.315000 -0.085000  8.485000 0.085000 ;
        RECT  8.795000 -0.085000  8.965000 0.085000 ;
        RECT  9.275000 -0.085000  9.445000 0.085000 ;
        RECT  9.755000 -0.085000  9.925000 0.085000 ;
        RECT 10.235000 -0.085000 10.405000 0.085000 ;
        RECT 10.715000 -0.085000 10.885000 0.085000 ;
        RECT 11.195000 -0.085000 11.365000 0.085000 ;
        RECT 11.675000 -0.085000 11.845000 0.085000 ;
        RECT 12.155000 -0.085000 12.325000 0.085000 ;
        RECT 12.635000 -0.085000 12.805000 0.085000 ;
        RECT 13.115000 -0.085000 13.285000 0.085000 ;
        RECT 13.595000 -0.085000 13.765000 0.085000 ;
        RECT 14.075000 -0.085000 14.245000 0.085000 ;
        RECT 14.555000 -0.085000 14.725000 0.085000 ;
        RECT 15.035000 -0.085000 15.205000 0.085000 ;
        RECT 15.515000 -0.085000 15.685000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 15.840000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 3.245000 15.840000 3.415000 ;
        RECT  0.615000 2.645000  0.945000 3.245000 ;
        RECT  2.505000 2.520000  2.755000 3.245000 ;
        RECT  4.045000 2.180000  4.215000 3.245000 ;
        RECT  6.595000 2.075000  6.925000 3.245000 ;
        RECT  8.315000 2.505000  8.685000 3.245000 ;
        RECT 10.435000 2.660000 11.150000 3.245000 ;
        RECT 12.295000 2.480000 12.625000 3.245000 ;
        RECT 13.340000 2.480000 13.670000 3.245000 ;
        RECT 14.945000 2.115000 15.205000 3.245000 ;
      LAYER mcon ;
        RECT  0.155000 3.245000  0.325000 3.415000 ;
        RECT  0.635000 3.245000  0.805000 3.415000 ;
        RECT  1.115000 3.245000  1.285000 3.415000 ;
        RECT  1.595000 3.245000  1.765000 3.415000 ;
        RECT  2.075000 3.245000  2.245000 3.415000 ;
        RECT  2.555000 3.245000  2.725000 3.415000 ;
        RECT  3.035000 3.245000  3.205000 3.415000 ;
        RECT  3.515000 3.245000  3.685000 3.415000 ;
        RECT  3.995000 3.245000  4.165000 3.415000 ;
        RECT  4.475000 3.245000  4.645000 3.415000 ;
        RECT  4.955000 3.245000  5.125000 3.415000 ;
        RECT  5.435000 3.245000  5.605000 3.415000 ;
        RECT  5.915000 3.245000  6.085000 3.415000 ;
        RECT  6.395000 3.245000  6.565000 3.415000 ;
        RECT  6.875000 3.245000  7.045000 3.415000 ;
        RECT  7.355000 3.245000  7.525000 3.415000 ;
        RECT  7.835000 3.245000  8.005000 3.415000 ;
        RECT  8.315000 3.245000  8.485000 3.415000 ;
        RECT  8.795000 3.245000  8.965000 3.415000 ;
        RECT  9.275000 3.245000  9.445000 3.415000 ;
        RECT  9.755000 3.245000  9.925000 3.415000 ;
        RECT 10.235000 3.245000 10.405000 3.415000 ;
        RECT 10.715000 3.245000 10.885000 3.415000 ;
        RECT 11.195000 3.245000 11.365000 3.415000 ;
        RECT 11.675000 3.245000 11.845000 3.415000 ;
        RECT 12.155000 3.245000 12.325000 3.415000 ;
        RECT 12.635000 3.245000 12.805000 3.415000 ;
        RECT 13.115000 3.245000 13.285000 3.415000 ;
        RECT 13.595000 3.245000 13.765000 3.415000 ;
        RECT 14.075000 3.245000 14.245000 3.415000 ;
        RECT 14.555000 3.245000 14.725000 3.415000 ;
        RECT 15.035000 3.245000 15.205000 3.415000 ;
        RECT 15.515000 3.245000 15.685000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 15.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.115000 2.305000  1.285000 2.475000 ;
      RECT  0.115000 2.475000  0.445000 2.980000 ;
      RECT  1.040000 0.575000  1.370000 1.185000 ;
      RECT  1.040000 1.185000  2.420000 1.355000 ;
      RECT  1.115000 2.475000  1.285000 2.905000 ;
      RECT  1.115000 2.905000  2.275000 3.075000 ;
      RECT  1.495000 2.025000  2.105000 2.195000 ;
      RECT  1.495000 2.195000  1.745000 2.735000 ;
      RECT  1.935000 1.355000  2.105000 2.025000 ;
      RECT  1.945000 2.520000  2.275000 2.905000 ;
      RECT  2.250000 0.255000  3.680000 0.425000 ;
      RECT  2.250000 0.425000  2.420000 1.185000 ;
      RECT  2.275000 1.830000  2.780000 2.180000 ;
      RECT  2.275000 2.180000  3.285000 2.350000 ;
      RECT  2.610000 0.595000  2.860000 1.035000 ;
      RECT  2.610000 1.035000  2.780000 1.830000 ;
      RECT  2.955000 2.350000  3.285000 2.980000 ;
      RECT  3.090000 0.595000  3.340000 1.010000 ;
      RECT  3.090000 1.010000  3.260000 1.840000 ;
      RECT  3.090000 1.840000  4.245000 2.010000 ;
      RECT  3.510000 0.425000  3.680000 0.660000 ;
      RECT  3.510000 0.660000  5.335000 0.830000 ;
      RECT  3.515000 2.010000  3.845000 2.980000 ;
      RECT  4.075000 1.340000  4.565000 1.670000 ;
      RECT  4.075000 1.670000  4.245000 1.840000 ;
      RECT  4.360000 1.000000  4.905000 1.170000 ;
      RECT  4.415000 1.840000  4.905000 2.980000 ;
      RECT  4.735000 1.170000  4.905000 1.365000 ;
      RECT  4.735000 1.365000  5.445000 1.695000 ;
      RECT  4.735000 1.695000  4.905000 1.840000 ;
      RECT  5.005000 0.460000  5.335000 0.660000 ;
      RECT  5.075000 1.865000  5.785000 2.035000 ;
      RECT  5.075000 2.035000  5.405000 2.755000 ;
      RECT  5.165000 0.830000  5.335000 1.025000 ;
      RECT  5.165000 1.025000  5.785000 1.195000 ;
      RECT  5.505000 0.460000  5.835000 0.685000 ;
      RECT  5.505000 0.685000  6.125000 0.855000 ;
      RECT  5.575000 2.205000  6.125000 2.535000 ;
      RECT  5.615000 1.195000  5.785000 1.865000 ;
      RECT  5.955000 0.855000  6.125000 1.655000 ;
      RECT  5.955000 1.655000  6.875000 1.825000 ;
      RECT  5.955000 1.825000  6.125000 2.205000 ;
      RECT  6.295000 0.730000  8.855000 0.900000 ;
      RECT  6.295000 0.900000  6.535000 1.485000 ;
      RECT  6.705000 1.070000  7.915000 1.240000 ;
      RECT  6.705000 1.240000  6.875000 1.655000 ;
      RECT  7.145000 0.310000  8.715000 0.480000 ;
      RECT  7.145000 0.480000  7.640000 0.560000 ;
      RECT  7.435000 1.825000  9.015000 1.995000 ;
      RECT  7.435000 1.995000  7.765000 2.735000 ;
      RECT  7.585000 1.240000  7.915000 1.585000 ;
      RECT  7.820000 0.655000  8.150000 0.730000 ;
      RECT  8.125000 1.180000  8.515000 1.585000 ;
      RECT  8.330000 0.480000  8.715000 0.560000 ;
      RECT  8.685000 0.900000  8.855000 1.335000 ;
      RECT  8.685000 1.335000  9.015000 1.825000 ;
      RECT  9.255000 1.335000  9.615000 1.505000 ;
      RECT  9.255000 1.505000  9.585000 1.940000 ;
      RECT  9.375000 2.110000  9.925000 2.735000 ;
      RECT  9.445000 0.255000 10.485000 0.425000 ;
      RECT  9.445000 0.425000  9.615000 1.335000 ;
      RECT  9.755000 1.675000  9.955000 1.845000 ;
      RECT  9.755000 1.845000  9.925000 2.110000 ;
      RECT  9.785000 0.595000  9.985000 1.350000 ;
      RECT  9.785000 1.350000 10.885000 1.520000 ;
      RECT  9.785000 1.520000  9.955000 1.675000 ;
      RECT 10.155000 0.425000 10.485000 1.180000 ;
      RECT 10.465000 2.030000 10.795000 2.320000 ;
      RECT 10.465000 2.320000 11.785000 2.490000 ;
      RECT 10.715000 1.180000 11.875000 1.350000 ;
      RECT 11.330000 0.255000 12.555000 0.425000 ;
      RECT 11.330000 0.425000 11.660000 1.010000 ;
      RECT 11.535000 1.970000 12.215000 2.140000 ;
      RECT 11.535000 2.140000 13.700000 2.310000 ;
      RECT 11.535000 2.310000 11.785000 2.320000 ;
      RECT 11.535000 2.490000 11.785000 2.980000 ;
      RECT 11.595000 1.350000 11.875000 1.550000 ;
      RECT 11.870000 0.595000 12.215000 1.010000 ;
      RECT 12.045000 1.010000 12.215000 1.970000 ;
      RECT 12.385000 0.425000 12.555000 1.010000 ;
      RECT 12.445000 1.180000 12.895000 1.720000 ;
      RECT 12.725000 0.670000 13.115000 1.010000 ;
      RECT 12.725000 1.010000 12.895000 1.180000 ;
      RECT 12.725000 1.720000 13.155000 1.970000 ;
      RECT 13.530000 1.220000 13.915000 1.550000 ;
      RECT 13.530000 1.550000 13.700000 2.140000 ;
      RECT 14.445000 0.350000 14.715000 1.355000 ;
      RECT 14.445000 1.355000 14.845000 1.685000 ;
      RECT 14.445000 1.685000 14.775000 2.980000 ;
    LAYER mcon ;
      RECT  8.315000 1.210000  8.485000 1.380000 ;
      RECT 12.635000 1.210000 12.805000 1.380000 ;
    LAYER met1 ;
      RECT  8.255000 1.180000  8.545000 1.225000 ;
      RECT  8.255000 1.225000 12.865000 1.365000 ;
      RECT  8.255000 1.365000  8.545000 1.410000 ;
      RECT 12.575000 1.180000 12.865000 1.225000 ;
      RECT 12.575000 1.365000 12.865000 1.410000 ;
  END
END sky130_fd_sc_ls__sdfbbp_1
