* File: sky130_fd_sc_ls__and2b_4.pxi.spice
* Created: Fri Aug 28 13:03:40 2020
* 
x_PM_SKY130_FD_SC_LS__AND2B_4%A_N N_A_N_c_109_n N_A_N_M1017_g N_A_N_M1009_g A_N
+ PM_SKY130_FD_SC_LS__AND2B_4%A_N
x_PM_SKY130_FD_SC_LS__AND2B_4%B N_B_M1007_g N_B_c_149_n N_B_M1002_g N_B_c_150_n
+ N_B_c_151_n N_B_c_143_n N_B_c_153_n N_B_M1008_g N_B_M1015_g N_B_c_154_n
+ N_B_c_145_n N_B_c_156_n N_B_c_146_n B B N_B_c_148_n
+ PM_SKY130_FD_SC_LS__AND2B_4%B
x_PM_SKY130_FD_SC_LS__AND2B_4%A_27_392# N_A_27_392#_M1009_s N_A_27_392#_M1017_s
+ N_A_27_392#_c_256_n N_A_27_392#_M1003_g N_A_27_392#_c_257_n
+ N_A_27_392#_c_258_n N_A_27_392#_c_259_n N_A_27_392#_M1010_g
+ N_A_27_392#_c_247_n N_A_27_392#_M1005_g N_A_27_392#_c_248_n
+ N_A_27_392#_c_249_n N_A_27_392#_M1014_g N_A_27_392#_c_261_n
+ N_A_27_392#_c_250_n N_A_27_392#_c_262_n N_A_27_392#_c_263_n
+ N_A_27_392#_c_251_n N_A_27_392#_c_252_n N_A_27_392#_c_253_n
+ N_A_27_392#_c_254_n N_A_27_392#_c_255_n PM_SKY130_FD_SC_LS__AND2B_4%A_27_392#
x_PM_SKY130_FD_SC_LS__AND2B_4%A_218_424# N_A_218_424#_M1005_d
+ N_A_218_424#_M1003_d N_A_218_424#_M1002_d N_A_218_424#_M1000_g
+ N_A_218_424#_c_353_n N_A_218_424#_M1001_g N_A_218_424#_M1006_g
+ N_A_218_424#_c_354_n N_A_218_424#_M1004_g N_A_218_424#_c_355_n
+ N_A_218_424#_M1011_g N_A_218_424#_c_345_n N_A_218_424#_M1012_g
+ N_A_218_424#_c_346_n N_A_218_424#_c_347_n N_A_218_424#_c_348_n
+ N_A_218_424#_M1013_g N_A_218_424#_c_349_n N_A_218_424#_c_358_n
+ N_A_218_424#_M1016_g N_A_218_424#_c_350_n N_A_218_424#_c_359_n
+ N_A_218_424#_c_360_n N_A_218_424#_c_365_n N_A_218_424#_c_382_n
+ N_A_218_424#_c_361_n N_A_218_424#_c_362_n N_A_218_424#_c_351_n
+ N_A_218_424#_c_363_n N_A_218_424#_c_458_p N_A_218_424#_c_397_n
+ N_A_218_424#_c_352_n PM_SKY130_FD_SC_LS__AND2B_4%A_218_424#
x_PM_SKY130_FD_SC_LS__AND2B_4%VPWR N_VPWR_M1017_d N_VPWR_M1010_s N_VPWR_M1008_s
+ N_VPWR_M1004_d N_VPWR_M1016_d N_VPWR_c_520_n N_VPWR_c_521_n N_VPWR_c_522_n
+ N_VPWR_c_523_n N_VPWR_c_524_n N_VPWR_c_525_n N_VPWR_c_526_n N_VPWR_c_527_n
+ VPWR N_VPWR_c_528_n N_VPWR_c_529_n N_VPWR_c_530_n N_VPWR_c_531_n
+ N_VPWR_c_532_n N_VPWR_c_533_n N_VPWR_c_534_n N_VPWR_c_519_n
+ PM_SKY130_FD_SC_LS__AND2B_4%VPWR
x_PM_SKY130_FD_SC_LS__AND2B_4%X N_X_M1000_s N_X_M1012_s N_X_M1001_s N_X_M1011_s
+ N_X_c_598_n N_X_c_607_n N_X_c_608_n N_X_c_599_n N_X_c_600_n N_X_c_609_n
+ N_X_c_601_n N_X_c_610_n N_X_c_611_n N_X_c_602_n N_X_c_603_n N_X_c_604_n
+ N_X_c_605_n N_X_c_653_n X PM_SKY130_FD_SC_LS__AND2B_4%X
x_PM_SKY130_FD_SC_LS__AND2B_4%VGND N_VGND_M1009_d N_VGND_M1015_s N_VGND_M1006_d
+ N_VGND_M1013_d N_VGND_c_681_n N_VGND_c_682_n N_VGND_c_683_n N_VGND_c_684_n
+ N_VGND_c_685_n VGND N_VGND_c_686_n N_VGND_c_687_n N_VGND_c_688_n
+ N_VGND_c_689_n N_VGND_c_690_n N_VGND_c_691_n N_VGND_c_692_n
+ PM_SKY130_FD_SC_LS__AND2B_4%VGND
x_PM_SKY130_FD_SC_LS__AND2B_4%A_233_74# N_A_233_74#_M1007_d N_A_233_74#_M1014_s
+ N_A_233_74#_c_754_n N_A_233_74#_c_750_n N_A_233_74#_c_751_n
+ PM_SKY130_FD_SC_LS__AND2B_4%A_233_74#
cc_1 VNB N_A_N_c_109_n 0.0197733f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.885
cc_2 VNB N_A_N_M1009_g 0.0425761f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=0.69
cc_3 VNB A_N 0.00184438f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_4 VNB N_B_M1007_g 0.030296f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.46
cc_5 VNB N_B_c_143_n 0.00618265f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.615
cc_6 VNB N_B_M1015_g 0.0236056f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_B_c_145_n 0.00619883f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_B_c_146_n 0.0253169f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB B 0.00880776f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_B_c_148_n 0.0329693f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_27_392#_c_247_n 0.0176057f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.615
cc_12 VNB N_A_27_392#_c_248_n 0.0123802f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_392#_c_249_n 0.0173846f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_392#_c_250_n 0.0368859f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_392#_c_251_n 0.0179929f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_27_392#_c_252_n 0.0154055f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_27_392#_c_253_n 0.0189908f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_27_392#_c_254_n 0.00357485f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_27_392#_c_255_n 0.0432998f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_218_424#_M1000_g 0.0212213f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.615
cc_21 VNB N_A_218_424#_M1006_g 0.0218136f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_218_424#_c_345_n 0.0151946f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_218_424#_c_346_n 0.0084015f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_218_424#_c_347_n 0.0751846f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_218_424#_c_348_n 0.0170341f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_218_424#_c_349_n 0.0141907f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_218_424#_c_350_n 0.0120521f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_218_424#_c_351_n 0.00151958f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_218_424#_c_352_n 0.00204131f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VPWR_c_519_n 0.203486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_X_c_598_n 0.00179817f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.615
cc_32 VNB N_X_c_599_n 0.00296071f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_X_c_600_n 0.00151717f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_X_c_601_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_X_c_602_n 0.00879366f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_X_c_603_n 0.0127874f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_X_c_604_n 0.00248839f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_X_c_605_n 0.00212146f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB X 0.0161443f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_681_n 0.00641543f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_682_n 0.00568769f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_683_n 0.00420532f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_684_n 0.0125057f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_685_n 0.0262963f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_686_n 0.0383162f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_687_n 0.0155668f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_688_n 0.0183662f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_689_n 0.027356f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_690_n 0.00613614f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_691_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_692_n 0.275826f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_233_74#_c_750_n 0.00250269f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=1.615
cc_53 VNB N_A_233_74#_c_751_n 0.00513172f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.615
cc_54 VPB N_A_N_c_109_n 0.0444206f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.885
cc_55 VPB A_N 0.0017388f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_56 VPB N_B_c_149_n 0.0156453f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=0.69
cc_57 VPB N_B_c_150_n 0.013158f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_58 VPB N_B_c_151_n 0.0100007f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_B_c_143_n 0.0146326f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=1.615
cc_60 VPB N_B_c_153_n 0.0156453f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=1.615
cc_61 VPB N_B_c_154_n 0.00811706f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_B_c_145_n 0.00562027f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_B_c_156_n 0.00327454f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_B_c_146_n 0.00489863f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB B 0.00399067f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_A_27_392#_c_256_n 0.0160881f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_A_27_392#_c_257_n 0.0137572f $X=-0.19 $Y=1.66 $X2=0.575 $Y2=1.615
cc_68 VPB N_A_27_392#_c_258_n 0.0104187f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=1.615
cc_69 VPB N_A_27_392#_c_259_n 0.0156461f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=1.615
cc_70 VPB N_A_27_392#_c_248_n 0.0180254f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_A_27_392#_c_261_n 0.0132346f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_A_27_392#_c_262_n 0.00932683f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_A_27_392#_c_263_n 0.0367128f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_A_27_392#_c_253_n 0.0139518f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_A_218_424#_c_353_n 0.0154065f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_A_218_424#_c_354_n 0.0148772f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_A_218_424#_c_355_n 0.0148649f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_A_218_424#_c_347_n 0.019561f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 VPB N_A_218_424#_c_349_n 0.00117364f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 VPB N_A_218_424#_c_358_n 0.0274153f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_A_218_424#_c_359_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 VPB N_A_218_424#_c_360_n 0.00167726f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 VPB N_A_218_424#_c_361_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_84 VPB N_A_218_424#_c_362_n 7.68838e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_A_218_424#_c_363_n 0.00136909f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_520_n 0.00811085f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_521_n 0.0202859f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_522_n 0.0089291f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_523_n 0.0199421f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_524_n 0.00591275f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_525_n 0.00261791f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_526_n 0.0116916f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_527_n 0.0566911f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_528_n 0.0175529f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_529_n 0.0164465f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_530_n 0.0164465f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_531_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_532_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_533_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_534_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_519_n 0.0754071f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_102 VPB N_X_c_607_n 0.00118063f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 VPB N_X_c_608_n 0.00180921f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB N_X_c_609_n 0.00305019f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_105 VPB N_X_c_610_n 0.00288841f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_X_c_611_n 0.00180921f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 N_A_N_M1009_g N_B_M1007_g 0.0251047f $X=0.59 $Y=0.69 $X2=0 $Y2=0
cc_108 N_A_N_c_109_n N_B_c_156_n 0.00115407f $X=0.495 $Y=1.885 $X2=0 $Y2=0
cc_109 A_N N_B_c_156_n 0.0267667f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_110 N_A_N_c_109_n N_B_c_146_n 0.0130918f $X=0.495 $Y=1.885 $X2=0 $Y2=0
cc_111 N_A_N_M1009_g N_B_c_146_n 0.00456823f $X=0.59 $Y=0.69 $X2=0 $Y2=0
cc_112 A_N N_B_c_146_n 0.00140103f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_113 N_A_N_c_109_n N_A_27_392#_c_256_n 0.017168f $X=0.495 $Y=1.885 $X2=0 $Y2=0
cc_114 N_A_N_c_109_n N_A_27_392#_c_258_n 0.00573773f $X=0.495 $Y=1.885 $X2=0
+ $Y2=0
cc_115 N_A_N_M1009_g N_A_27_392#_c_250_n 0.0117205f $X=0.59 $Y=0.69 $X2=0 $Y2=0
cc_116 N_A_N_c_109_n N_A_27_392#_c_262_n 0.00687876f $X=0.495 $Y=1.885 $X2=0
+ $Y2=0
cc_117 N_A_N_c_109_n N_A_27_392#_c_251_n 0.00177632f $X=0.495 $Y=1.885 $X2=0
+ $Y2=0
cc_118 N_A_N_M1009_g N_A_27_392#_c_251_n 0.0115584f $X=0.59 $Y=0.69 $X2=0 $Y2=0
cc_119 A_N N_A_27_392#_c_251_n 0.0184339f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_120 N_A_N_c_109_n N_A_27_392#_c_252_n 0.00334367f $X=0.495 $Y=1.885 $X2=0
+ $Y2=0
cc_121 N_A_N_M1009_g N_A_27_392#_c_252_n 0.00449058f $X=0.59 $Y=0.69 $X2=0 $Y2=0
cc_122 A_N N_A_27_392#_c_252_n 0.00898631f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_123 N_A_N_c_109_n N_A_27_392#_c_253_n 0.0136014f $X=0.495 $Y=1.885 $X2=0
+ $Y2=0
cc_124 N_A_N_M1009_g N_A_27_392#_c_253_n 0.00572006f $X=0.59 $Y=0.69 $X2=0 $Y2=0
cc_125 A_N N_A_27_392#_c_253_n 0.0250408f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_126 N_A_N_c_109_n N_A_218_424#_c_359_n 2.87917e-19 $X=0.495 $Y=1.885 $X2=0
+ $Y2=0
cc_127 N_A_N_c_109_n N_A_218_424#_c_365_n 5.59215e-19 $X=0.495 $Y=1.885 $X2=0
+ $Y2=0
cc_128 N_A_N_c_109_n N_VPWR_c_520_n 0.0217429f $X=0.495 $Y=1.885 $X2=0 $Y2=0
cc_129 A_N N_VPWR_c_520_n 0.0112377f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_130 N_A_N_c_109_n N_VPWR_c_528_n 0.00413917f $X=0.495 $Y=1.885 $X2=0 $Y2=0
cc_131 N_A_N_c_109_n N_VPWR_c_519_n 0.00821187f $X=0.495 $Y=1.885 $X2=0 $Y2=0
cc_132 N_A_N_M1009_g N_VGND_c_681_n 0.00615346f $X=0.59 $Y=0.69 $X2=0 $Y2=0
cc_133 N_A_N_M1009_g N_VGND_c_689_n 0.00434272f $X=0.59 $Y=0.69 $X2=0 $Y2=0
cc_134 N_A_N_M1009_g N_VGND_c_692_n 0.00824713f $X=0.59 $Y=0.69 $X2=0 $Y2=0
cc_135 N_B_c_145_n N_A_27_392#_c_257_n 0.00594459f $X=2.045 $Y=1.705 $X2=0 $Y2=0
cc_136 N_B_c_156_n N_A_27_392#_c_258_n 0.00408361f $X=1.14 $Y=1.52 $X2=0 $Y2=0
cc_137 N_B_c_146_n N_A_27_392#_c_258_n 0.0208602f $X=1.14 $Y=1.52 $X2=0 $Y2=0
cc_138 N_B_c_149_n N_A_27_392#_c_259_n 0.0178573f $X=1.985 $Y=2.045 $X2=0 $Y2=0
cc_139 N_B_M1007_g N_A_27_392#_c_247_n 0.0251644f $X=1.09 $Y=0.69 $X2=0 $Y2=0
cc_140 N_B_c_145_n N_A_27_392#_c_248_n 0.0118894f $X=2.045 $Y=1.705 $X2=0 $Y2=0
cc_141 N_B_c_156_n N_A_27_392#_c_248_n 4.97671e-19 $X=1.14 $Y=1.52 $X2=0 $Y2=0
cc_142 B N_A_27_392#_c_248_n 0.0040484f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_143 N_B_c_148_n N_A_27_392#_c_248_n 0.00646392f $X=2.47 $Y=1.385 $X2=0 $Y2=0
cc_144 N_B_M1015_g N_A_27_392#_c_249_n 0.0283032f $X=2.47 $Y=0.69 $X2=0 $Y2=0
cc_145 N_B_c_151_n N_A_27_392#_c_261_n 0.00993433f $X=2.06 $Y=1.97 $X2=0 $Y2=0
cc_146 N_B_M1007_g N_A_27_392#_c_250_n 7.4234e-19 $X=1.09 $Y=0.69 $X2=0 $Y2=0
cc_147 N_B_M1007_g N_A_27_392#_c_251_n 0.0149394f $X=1.09 $Y=0.69 $X2=0 $Y2=0
cc_148 N_B_c_145_n N_A_27_392#_c_251_n 0.00950432f $X=2.045 $Y=1.705 $X2=0 $Y2=0
cc_149 N_B_c_156_n N_A_27_392#_c_251_n 0.0243488f $X=1.14 $Y=1.52 $X2=0 $Y2=0
cc_150 N_B_c_146_n N_A_27_392#_c_251_n 0.00446668f $X=1.14 $Y=1.52 $X2=0 $Y2=0
cc_151 N_B_M1007_g N_A_27_392#_c_254_n 6.47392e-19 $X=1.09 $Y=0.69 $X2=0 $Y2=0
cc_152 N_B_M1015_g N_A_27_392#_c_254_n 2.55667e-19 $X=2.47 $Y=0.69 $X2=0 $Y2=0
cc_153 N_B_c_145_n N_A_27_392#_c_254_n 0.0243539f $X=2.045 $Y=1.705 $X2=0 $Y2=0
cc_154 N_B_c_156_n N_A_27_392#_c_254_n 9.50602e-19 $X=1.14 $Y=1.52 $X2=0 $Y2=0
cc_155 N_B_c_146_n N_A_27_392#_c_254_n 6.23084e-19 $X=1.14 $Y=1.52 $X2=0 $Y2=0
cc_156 B N_A_27_392#_c_254_n 0.0192912f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_157 N_B_c_151_n N_A_27_392#_c_255_n 0.0026999f $X=2.06 $Y=1.97 $X2=0 $Y2=0
cc_158 N_B_c_145_n N_A_27_392#_c_255_n 0.00607751f $X=2.045 $Y=1.705 $X2=0 $Y2=0
cc_159 N_B_c_156_n N_A_27_392#_c_255_n 0.00118989f $X=1.14 $Y=1.52 $X2=0 $Y2=0
cc_160 N_B_c_146_n N_A_27_392#_c_255_n 0.0214109f $X=1.14 $Y=1.52 $X2=0 $Y2=0
cc_161 B N_A_27_392#_c_255_n 0.00619253f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_162 N_B_c_148_n N_A_27_392#_c_255_n 0.00703692f $X=2.47 $Y=1.385 $X2=0 $Y2=0
cc_163 N_B_M1015_g N_A_218_424#_M1000_g 0.0220476f $X=2.47 $Y=0.69 $X2=0 $Y2=0
cc_164 B N_A_218_424#_M1000_g 3.49507e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_165 N_B_c_148_n N_A_218_424#_M1000_g 0.0127101f $X=2.47 $Y=1.385 $X2=0 $Y2=0
cc_166 N_B_c_143_n N_A_218_424#_c_353_n 0.00303511f $X=2.38 $Y=1.895 $X2=0 $Y2=0
cc_167 N_B_c_153_n N_A_218_424#_c_353_n 0.0184437f $X=2.435 $Y=2.045 $X2=0 $Y2=0
cc_168 N_B_c_154_n N_A_218_424#_c_353_n 0.00495829f $X=2.415 $Y=1.97 $X2=0 $Y2=0
cc_169 N_B_c_143_n N_A_218_424#_c_347_n 0.00573697f $X=2.38 $Y=1.895 $X2=0 $Y2=0
cc_170 B N_A_218_424#_c_347_n 7.65992e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_171 N_B_c_148_n N_A_218_424#_c_347_n 0.00443805f $X=2.47 $Y=1.385 $X2=0 $Y2=0
cc_172 N_B_c_149_n N_A_218_424#_c_359_n 6.92185e-19 $X=1.985 $Y=2.045 $X2=0
+ $Y2=0
cc_173 N_B_c_149_n N_A_218_424#_c_360_n 0.00817723f $X=1.985 $Y=2.045 $X2=0
+ $Y2=0
cc_174 N_B_c_151_n N_A_218_424#_c_360_n 0.00325231f $X=2.06 $Y=1.97 $X2=0 $Y2=0
cc_175 N_B_c_145_n N_A_218_424#_c_360_n 0.0460131f $X=2.045 $Y=1.705 $X2=0 $Y2=0
cc_176 N_B_c_145_n N_A_218_424#_c_365_n 0.00794883f $X=2.045 $Y=1.705 $X2=0
+ $Y2=0
cc_177 N_B_c_156_n N_A_218_424#_c_365_n 0.019374f $X=1.14 $Y=1.52 $X2=0 $Y2=0
cc_178 N_B_c_146_n N_A_218_424#_c_365_n 2.06523e-19 $X=1.14 $Y=1.52 $X2=0 $Y2=0
cc_179 N_B_M1015_g N_A_218_424#_c_382_n 0.0129721f $X=2.47 $Y=0.69 $X2=0 $Y2=0
cc_180 B N_A_218_424#_c_382_n 0.0275877f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_181 N_B_c_148_n N_A_218_424#_c_382_n 0.00178839f $X=2.47 $Y=1.385 $X2=0 $Y2=0
cc_182 N_B_c_149_n N_A_218_424#_c_361_n 0.0124504f $X=1.985 $Y=2.045 $X2=0 $Y2=0
cc_183 N_B_c_153_n N_A_218_424#_c_361_n 0.0124325f $X=2.435 $Y=2.045 $X2=0 $Y2=0
cc_184 N_B_c_153_n N_A_218_424#_c_362_n 0.00817723f $X=2.435 $Y=2.045 $X2=0
+ $Y2=0
cc_185 N_B_c_154_n N_A_218_424#_c_362_n 0.0041504f $X=2.415 $Y=1.97 $X2=0 $Y2=0
cc_186 B N_A_218_424#_c_362_n 0.0165376f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_187 N_B_c_148_n N_A_218_424#_c_362_n 0.00178207f $X=2.47 $Y=1.385 $X2=0 $Y2=0
cc_188 N_B_M1015_g N_A_218_424#_c_351_n 0.0052622f $X=2.47 $Y=0.69 $X2=0 $Y2=0
cc_189 B N_A_218_424#_c_351_n 0.0110703f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_190 N_B_c_148_n N_A_218_424#_c_351_n 6.31866e-19 $X=2.47 $Y=1.385 $X2=0 $Y2=0
cc_191 N_B_c_143_n N_A_218_424#_c_363_n 0.00233554f $X=2.38 $Y=1.895 $X2=0 $Y2=0
cc_192 N_B_c_154_n N_A_218_424#_c_363_n 0.00137158f $X=2.415 $Y=1.97 $X2=0 $Y2=0
cc_193 B N_A_218_424#_c_363_n 0.0115106f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_194 N_B_c_149_n N_A_218_424#_c_397_n 0.00104176f $X=1.985 $Y=2.045 $X2=0
+ $Y2=0
cc_195 N_B_c_150_n N_A_218_424#_c_397_n 0.00647252f $X=2.305 $Y=1.97 $X2=0 $Y2=0
cc_196 N_B_c_151_n N_A_218_424#_c_397_n 2.12488e-19 $X=2.06 $Y=1.97 $X2=0 $Y2=0
cc_197 N_B_c_153_n N_A_218_424#_c_397_n 0.00104176f $X=2.435 $Y=2.045 $X2=0
+ $Y2=0
cc_198 N_B_c_154_n N_A_218_424#_c_397_n 0.00157192f $X=2.415 $Y=1.97 $X2=0 $Y2=0
cc_199 B N_A_218_424#_c_397_n 0.0286849f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_200 N_B_c_143_n N_A_218_424#_c_352_n 3.22534e-19 $X=2.38 $Y=1.895 $X2=0 $Y2=0
cc_201 B N_A_218_424#_c_352_n 0.029241f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_202 N_B_c_148_n N_A_218_424#_c_352_n 0.00166039f $X=2.47 $Y=1.385 $X2=0 $Y2=0
cc_203 N_B_c_149_n N_VPWR_c_522_n 0.00663333f $X=1.985 $Y=2.045 $X2=0 $Y2=0
cc_204 N_B_c_149_n N_VPWR_c_523_n 0.00445602f $X=1.985 $Y=2.045 $X2=0 $Y2=0
cc_205 N_B_c_153_n N_VPWR_c_523_n 0.00445602f $X=2.435 $Y=2.045 $X2=0 $Y2=0
cc_206 N_B_c_153_n N_VPWR_c_524_n 0.00678915f $X=2.435 $Y=2.045 $X2=0 $Y2=0
cc_207 N_B_c_149_n N_VPWR_c_519_n 0.00858041f $X=1.985 $Y=2.045 $X2=0 $Y2=0
cc_208 N_B_c_153_n N_VPWR_c_519_n 0.00858041f $X=2.435 $Y=2.045 $X2=0 $Y2=0
cc_209 N_B_M1007_g N_VGND_c_681_n 0.0102293f $X=1.09 $Y=0.69 $X2=0 $Y2=0
cc_210 N_B_M1015_g N_VGND_c_682_n 0.00303986f $X=2.47 $Y=0.69 $X2=0 $Y2=0
cc_211 N_B_M1007_g N_VGND_c_686_n 0.00383152f $X=1.09 $Y=0.69 $X2=0 $Y2=0
cc_212 N_B_M1015_g N_VGND_c_686_n 0.00336923f $X=2.47 $Y=0.69 $X2=0 $Y2=0
cc_213 N_B_M1007_g N_VGND_c_692_n 0.00758251f $X=1.09 $Y=0.69 $X2=0 $Y2=0
cc_214 N_B_M1015_g N_VGND_c_692_n 0.00439691f $X=2.47 $Y=0.69 $X2=0 $Y2=0
cc_215 N_B_M1007_g N_A_233_74#_c_750_n 7.34787e-19 $X=1.09 $Y=0.69 $X2=0 $Y2=0
cc_216 N_B_M1015_g N_A_233_74#_c_751_n 0.0026545f $X=2.47 $Y=0.69 $X2=0 $Y2=0
cc_217 N_A_27_392#_c_256_n N_A_218_424#_c_359_n 0.0109401f $X=1.015 $Y=2.045
+ $X2=0 $Y2=0
cc_218 N_A_27_392#_c_259_n N_A_218_424#_c_359_n 0.0126119f $X=1.465 $Y=2.045
+ $X2=0 $Y2=0
cc_219 N_A_27_392#_c_259_n N_A_218_424#_c_360_n 0.00817723f $X=1.465 $Y=2.045
+ $X2=0 $Y2=0
cc_220 N_A_27_392#_c_261_n N_A_218_424#_c_360_n 0.00765867f $X=1.59 $Y=1.97
+ $X2=0 $Y2=0
cc_221 N_A_27_392#_c_256_n N_A_218_424#_c_365_n 0.00234049f $X=1.015 $Y=2.045
+ $X2=0 $Y2=0
cc_222 N_A_27_392#_c_257_n N_A_218_424#_c_365_n 0.00715034f $X=1.39 $Y=1.97
+ $X2=0 $Y2=0
cc_223 N_A_27_392#_c_258_n N_A_218_424#_c_365_n 0.00184982f $X=1.09 $Y=1.97
+ $X2=0 $Y2=0
cc_224 N_A_27_392#_c_259_n N_A_218_424#_c_365_n 0.00104176f $X=1.465 $Y=2.045
+ $X2=0 $Y2=0
cc_225 N_A_27_392#_c_261_n N_A_218_424#_c_365_n 2.21804e-19 $X=1.59 $Y=1.97
+ $X2=0 $Y2=0
cc_226 N_A_27_392#_c_247_n N_A_218_424#_c_382_n 0.00237855f $X=1.59 $Y=1.12
+ $X2=0 $Y2=0
cc_227 N_A_27_392#_c_249_n N_A_218_424#_c_382_n 0.0113406f $X=2.02 $Y=1.12 $X2=0
+ $Y2=0
cc_228 N_A_27_392#_c_254_n N_A_218_424#_c_382_n 0.0137945f $X=1.68 $Y=1.18 $X2=0
+ $Y2=0
cc_229 N_A_27_392#_c_255_n N_A_218_424#_c_382_n 9.53947e-19 $X=1.68 $Y=1.285
+ $X2=0 $Y2=0
cc_230 N_A_27_392#_c_259_n N_A_218_424#_c_361_n 6.13839e-19 $X=1.465 $Y=2.045
+ $X2=0 $Y2=0
cc_231 N_A_27_392#_c_256_n N_VPWR_c_520_n 0.00792774f $X=1.015 $Y=2.045 $X2=0
+ $Y2=0
cc_232 N_A_27_392#_c_263_n N_VPWR_c_520_n 0.0593822f $X=0.27 $Y=2.115 $X2=0
+ $Y2=0
cc_233 N_A_27_392#_c_256_n N_VPWR_c_521_n 0.00445602f $X=1.015 $Y=2.045 $X2=0
+ $Y2=0
cc_234 N_A_27_392#_c_259_n N_VPWR_c_521_n 0.00445602f $X=1.465 $Y=2.045 $X2=0
+ $Y2=0
cc_235 N_A_27_392#_c_259_n N_VPWR_c_522_n 0.00533971f $X=1.465 $Y=2.045 $X2=0
+ $Y2=0
cc_236 N_A_27_392#_c_261_n N_VPWR_c_522_n 3.72025e-19 $X=1.59 $Y=1.97 $X2=0
+ $Y2=0
cc_237 N_A_27_392#_c_263_n N_VPWR_c_528_n 0.0119584f $X=0.27 $Y=2.115 $X2=0
+ $Y2=0
cc_238 N_A_27_392#_c_256_n N_VPWR_c_519_n 0.00858041f $X=1.015 $Y=2.045 $X2=0
+ $Y2=0
cc_239 N_A_27_392#_c_259_n N_VPWR_c_519_n 0.00858265f $X=1.465 $Y=2.045 $X2=0
+ $Y2=0
cc_240 N_A_27_392#_c_263_n N_VPWR_c_519_n 0.00989813f $X=0.27 $Y=2.115 $X2=0
+ $Y2=0
cc_241 N_A_27_392#_c_247_n N_VGND_c_681_n 5.74073e-19 $X=1.59 $Y=1.12 $X2=0
+ $Y2=0
cc_242 N_A_27_392#_c_250_n N_VGND_c_681_n 0.0234524f $X=0.375 $Y=0.515 $X2=0
+ $Y2=0
cc_243 N_A_27_392#_c_251_n N_VGND_c_681_n 0.0238718f $X=1.515 $Y=1.18 $X2=0
+ $Y2=0
cc_244 N_A_27_392#_c_247_n N_VGND_c_686_n 0.00289603f $X=1.59 $Y=1.12 $X2=0
+ $Y2=0
cc_245 N_A_27_392#_c_249_n N_VGND_c_686_n 0.00289603f $X=2.02 $Y=1.12 $X2=0
+ $Y2=0
cc_246 N_A_27_392#_c_250_n N_VGND_c_689_n 0.0201415f $X=0.375 $Y=0.515 $X2=0
+ $Y2=0
cc_247 N_A_27_392#_c_247_n N_VGND_c_692_n 0.0035835f $X=1.59 $Y=1.12 $X2=0 $Y2=0
cc_248 N_A_27_392#_c_249_n N_VGND_c_692_n 0.00357919f $X=2.02 $Y=1.12 $X2=0
+ $Y2=0
cc_249 N_A_27_392#_c_250_n N_VGND_c_692_n 0.016615f $X=0.375 $Y=0.515 $X2=0
+ $Y2=0
cc_250 N_A_27_392#_c_251_n N_A_233_74#_c_754_n 0.0201258f $X=1.515 $Y=1.18 $X2=0
+ $Y2=0
cc_251 N_A_27_392#_c_247_n N_A_233_74#_c_751_n 0.0127013f $X=1.59 $Y=1.12 $X2=0
+ $Y2=0
cc_252 N_A_27_392#_c_249_n N_A_233_74#_c_751_n 0.0103014f $X=2.02 $Y=1.12 $X2=0
+ $Y2=0
cc_253 N_A_27_392#_c_254_n N_A_233_74#_c_751_n 0.00374521f $X=1.68 $Y=1.18 $X2=0
+ $Y2=0
cc_254 N_A_218_424#_c_360_n N_VPWR_M1010_s 0.00296906f $X=2.045 $Y=2.045 $X2=0
+ $Y2=0
cc_255 N_A_218_424#_c_362_n N_VPWR_M1008_s 0.00755397f $X=2.755 $Y=2.045 $X2=0
+ $Y2=0
cc_256 N_A_218_424#_c_363_n N_VPWR_M1008_s 0.00148303f $X=2.84 $Y=1.96 $X2=0
+ $Y2=0
cc_257 N_A_218_424#_c_359_n N_VPWR_c_520_n 0.0298716f $X=1.24 $Y=2.265 $X2=0
+ $Y2=0
cc_258 N_A_218_424#_c_365_n N_VPWR_c_520_n 0.00188899f $X=1.405 $Y=2.045 $X2=0
+ $Y2=0
cc_259 N_A_218_424#_c_359_n N_VPWR_c_521_n 0.014552f $X=1.24 $Y=2.265 $X2=0
+ $Y2=0
cc_260 N_A_218_424#_c_359_n N_VPWR_c_522_n 0.0456243f $X=1.24 $Y=2.265 $X2=0
+ $Y2=0
cc_261 N_A_218_424#_c_360_n N_VPWR_c_522_n 0.0200955f $X=2.045 $Y=2.045 $X2=0
+ $Y2=0
cc_262 N_A_218_424#_c_361_n N_VPWR_c_522_n 0.0240409f $X=2.21 $Y=2.265 $X2=0
+ $Y2=0
cc_263 N_A_218_424#_c_361_n N_VPWR_c_523_n 0.014552f $X=2.21 $Y=2.265 $X2=0
+ $Y2=0
cc_264 N_A_218_424#_c_353_n N_VPWR_c_524_n 0.0109116f $X=2.955 $Y=1.765 $X2=0
+ $Y2=0
cc_265 N_A_218_424#_c_354_n N_VPWR_c_524_n 5.32946e-19 $X=3.405 $Y=1.765 $X2=0
+ $Y2=0
cc_266 N_A_218_424#_c_361_n N_VPWR_c_524_n 0.0240709f $X=2.21 $Y=2.265 $X2=0
+ $Y2=0
cc_267 N_A_218_424#_c_362_n N_VPWR_c_524_n 0.0224876f $X=2.755 $Y=2.045 $X2=0
+ $Y2=0
cc_268 N_A_218_424#_c_353_n N_VPWR_c_525_n 5.75502e-19 $X=2.955 $Y=1.765 $X2=0
+ $Y2=0
cc_269 N_A_218_424#_c_354_n N_VPWR_c_525_n 0.0136211f $X=3.405 $Y=1.765 $X2=0
+ $Y2=0
cc_270 N_A_218_424#_c_355_n N_VPWR_c_525_n 0.0136211f $X=3.855 $Y=1.765 $X2=0
+ $Y2=0
cc_271 N_A_218_424#_c_358_n N_VPWR_c_525_n 5.75502e-19 $X=4.305 $Y=1.765 $X2=0
+ $Y2=0
cc_272 N_A_218_424#_c_355_n N_VPWR_c_527_n 6.868e-19 $X=3.855 $Y=1.765 $X2=0
+ $Y2=0
cc_273 N_A_218_424#_c_358_n N_VPWR_c_527_n 0.0186135f $X=4.305 $Y=1.765 $X2=0
+ $Y2=0
cc_274 N_A_218_424#_c_353_n N_VPWR_c_529_n 0.00413917f $X=2.955 $Y=1.765 $X2=0
+ $Y2=0
cc_275 N_A_218_424#_c_354_n N_VPWR_c_529_n 0.00413917f $X=3.405 $Y=1.765 $X2=0
+ $Y2=0
cc_276 N_A_218_424#_c_355_n N_VPWR_c_530_n 0.00413917f $X=3.855 $Y=1.765 $X2=0
+ $Y2=0
cc_277 N_A_218_424#_c_358_n N_VPWR_c_530_n 0.00413917f $X=4.305 $Y=1.765 $X2=0
+ $Y2=0
cc_278 N_A_218_424#_c_353_n N_VPWR_c_519_n 0.00817726f $X=2.955 $Y=1.765 $X2=0
+ $Y2=0
cc_279 N_A_218_424#_c_354_n N_VPWR_c_519_n 0.00817726f $X=3.405 $Y=1.765 $X2=0
+ $Y2=0
cc_280 N_A_218_424#_c_355_n N_VPWR_c_519_n 0.00817726f $X=3.855 $Y=1.765 $X2=0
+ $Y2=0
cc_281 N_A_218_424#_c_358_n N_VPWR_c_519_n 0.00817726f $X=4.305 $Y=1.765 $X2=0
+ $Y2=0
cc_282 N_A_218_424#_c_359_n N_VPWR_c_519_n 0.0119791f $X=1.24 $Y=2.265 $X2=0
+ $Y2=0
cc_283 N_A_218_424#_c_361_n N_VPWR_c_519_n 0.0119791f $X=2.21 $Y=2.265 $X2=0
+ $Y2=0
cc_284 N_A_218_424#_M1000_g N_X_c_598_n 0.00497662f $X=2.955 $Y=0.74 $X2=0 $Y2=0
cc_285 N_A_218_424#_M1006_g N_X_c_598_n 4.02861e-19 $X=3.395 $Y=0.74 $X2=0 $Y2=0
cc_286 N_A_218_424#_c_382_n N_X_c_598_n 0.0133617f $X=2.755 $Y=0.84 $X2=0 $Y2=0
cc_287 N_A_218_424#_c_351_n N_X_c_598_n 0.00379102f $X=2.84 $Y=1.32 $X2=0 $Y2=0
cc_288 N_A_218_424#_c_353_n N_X_c_607_n 7.2962e-19 $X=2.955 $Y=1.765 $X2=0 $Y2=0
cc_289 N_A_218_424#_c_347_n N_X_c_607_n 0.00419691f $X=3.945 $Y=1.26 $X2=0 $Y2=0
cc_290 N_A_218_424#_c_362_n N_X_c_607_n 0.00262209f $X=2.755 $Y=2.045 $X2=0
+ $Y2=0
cc_291 N_A_218_424#_c_363_n N_X_c_607_n 0.0110509f $X=2.84 $Y=1.96 $X2=0 $Y2=0
cc_292 N_A_218_424#_c_458_p N_X_c_607_n 0.0143367f $X=3.725 $Y=1.485 $X2=0 $Y2=0
cc_293 N_A_218_424#_c_353_n N_X_c_608_n 0.0061328f $X=2.955 $Y=1.765 $X2=0 $Y2=0
cc_294 N_A_218_424#_c_354_n N_X_c_608_n 0.00617886f $X=3.405 $Y=1.765 $X2=0
+ $Y2=0
cc_295 N_A_218_424#_c_362_n N_X_c_608_n 0.0109673f $X=2.755 $Y=2.045 $X2=0 $Y2=0
cc_296 N_A_218_424#_M1006_g N_X_c_599_n 0.0128363f $X=3.395 $Y=0.74 $X2=0 $Y2=0
cc_297 N_A_218_424#_c_345_n N_X_c_599_n 0.01254f $X=3.86 $Y=1.185 $X2=0 $Y2=0
cc_298 N_A_218_424#_c_347_n N_X_c_599_n 0.00302677f $X=3.945 $Y=1.26 $X2=0 $Y2=0
cc_299 N_A_218_424#_c_458_p N_X_c_599_n 0.0413425f $X=3.725 $Y=1.485 $X2=0 $Y2=0
cc_300 N_A_218_424#_M1000_g N_X_c_600_n 8.1288e-19 $X=2.955 $Y=0.74 $X2=0 $Y2=0
cc_301 N_A_218_424#_c_347_n N_X_c_600_n 0.00256252f $X=3.945 $Y=1.26 $X2=0 $Y2=0
cc_302 N_A_218_424#_c_351_n N_X_c_600_n 0.0134877f $X=2.84 $Y=1.32 $X2=0 $Y2=0
cc_303 N_A_218_424#_c_458_p N_X_c_600_n 0.0143379f $X=3.725 $Y=1.485 $X2=0 $Y2=0
cc_304 N_A_218_424#_c_354_n N_X_c_609_n 0.0128248f $X=3.405 $Y=1.765 $X2=0 $Y2=0
cc_305 N_A_218_424#_c_355_n N_X_c_609_n 0.0143722f $X=3.855 $Y=1.765 $X2=0 $Y2=0
cc_306 N_A_218_424#_c_347_n N_X_c_609_n 0.00980221f $X=3.945 $Y=1.26 $X2=0 $Y2=0
cc_307 N_A_218_424#_c_458_p N_X_c_609_n 0.0413195f $X=3.725 $Y=1.485 $X2=0 $Y2=0
cc_308 N_A_218_424#_M1006_g N_X_c_601_n 6.54757e-19 $X=3.395 $Y=0.74 $X2=0 $Y2=0
cc_309 N_A_218_424#_c_345_n N_X_c_601_n 0.00939704f $X=3.86 $Y=1.185 $X2=0 $Y2=0
cc_310 N_A_218_424#_c_348_n N_X_c_601_n 3.97481e-19 $X=4.29 $Y=1.185 $X2=0 $Y2=0
cc_311 N_A_218_424#_c_355_n N_X_c_610_n 0.00128638f $X=3.855 $Y=1.765 $X2=0
+ $Y2=0
cc_312 N_A_218_424#_c_347_n N_X_c_610_n 0.00274694f $X=3.945 $Y=1.26 $X2=0 $Y2=0
cc_313 N_A_218_424#_c_349_n N_X_c_610_n 0.00274264f $X=4.305 $Y=1.675 $X2=0
+ $Y2=0
cc_314 N_A_218_424#_c_358_n N_X_c_610_n 0.00128638f $X=4.305 $Y=1.765 $X2=0
+ $Y2=0
cc_315 N_A_218_424#_c_355_n N_X_c_611_n 0.00617886f $X=3.855 $Y=1.765 $X2=0
+ $Y2=0
cc_316 N_A_218_424#_c_358_n N_X_c_611_n 0.0034263f $X=4.305 $Y=1.765 $X2=0 $Y2=0
cc_317 N_A_218_424#_c_348_n N_X_c_602_n 0.0148509f $X=4.29 $Y=1.185 $X2=0 $Y2=0
cc_318 N_A_218_424#_c_350_n N_X_c_602_n 7.8992e-19 $X=4.215 $Y=1.185 $X2=0 $Y2=0
cc_319 N_A_218_424#_c_349_n N_X_c_603_n 0.0176895f $X=4.305 $Y=1.675 $X2=0 $Y2=0
cc_320 N_A_218_424#_c_346_n N_X_c_604_n 0.00208718f $X=4.215 $Y=1.26 $X2=0 $Y2=0
cc_321 N_A_218_424#_c_347_n N_X_c_604_n 0.00167782f $X=3.945 $Y=1.26 $X2=0 $Y2=0
cc_322 N_A_218_424#_c_458_p N_X_c_604_n 0.015065f $X=3.725 $Y=1.485 $X2=0 $Y2=0
cc_323 N_A_218_424#_c_345_n N_X_c_605_n 0.0015557f $X=3.86 $Y=1.185 $X2=0 $Y2=0
cc_324 N_A_218_424#_c_346_n N_X_c_605_n 0.00276997f $X=4.215 $Y=1.26 $X2=0 $Y2=0
cc_325 N_A_218_424#_c_358_n N_X_c_653_n 8.33339e-19 $X=4.305 $Y=1.765 $X2=0
+ $Y2=0
cc_326 N_A_218_424#_c_348_n X 0.00806324f $X=4.29 $Y=1.185 $X2=0 $Y2=0
cc_327 N_A_218_424#_c_350_n X 0.00418807f $X=4.215 $Y=1.185 $X2=0 $Y2=0
cc_328 N_A_218_424#_c_458_p X 0.00476845f $X=3.725 $Y=1.485 $X2=0 $Y2=0
cc_329 N_A_218_424#_c_382_n N_VGND_M1015_s 0.00728075f $X=2.755 $Y=0.84 $X2=0
+ $Y2=0
cc_330 N_A_218_424#_c_351_n N_VGND_M1015_s 0.00219581f $X=2.84 $Y=1.32 $X2=0
+ $Y2=0
cc_331 N_A_218_424#_M1000_g N_VGND_c_682_n 0.00650608f $X=2.955 $Y=0.74 $X2=0
+ $Y2=0
cc_332 N_A_218_424#_M1006_g N_VGND_c_682_n 3.97853e-19 $X=3.395 $Y=0.74 $X2=0
+ $Y2=0
cc_333 N_A_218_424#_c_382_n N_VGND_c_682_n 0.0194555f $X=2.755 $Y=0.84 $X2=0
+ $Y2=0
cc_334 N_A_218_424#_M1000_g N_VGND_c_683_n 4.63452e-19 $X=2.955 $Y=0.74 $X2=0
+ $Y2=0
cc_335 N_A_218_424#_M1006_g N_VGND_c_683_n 0.00960479f $X=3.395 $Y=0.74 $X2=0
+ $Y2=0
cc_336 N_A_218_424#_c_345_n N_VGND_c_683_n 0.00347183f $X=3.86 $Y=1.185 $X2=0
+ $Y2=0
cc_337 N_A_218_424#_c_345_n N_VGND_c_685_n 5.14978e-19 $X=3.86 $Y=1.185 $X2=0
+ $Y2=0
cc_338 N_A_218_424#_c_348_n N_VGND_c_685_n 0.011928f $X=4.29 $Y=1.185 $X2=0
+ $Y2=0
cc_339 N_A_218_424#_c_382_n N_VGND_c_686_n 0.00199065f $X=2.755 $Y=0.84 $X2=0
+ $Y2=0
cc_340 N_A_218_424#_M1000_g N_VGND_c_687_n 0.00378853f $X=2.955 $Y=0.74 $X2=0
+ $Y2=0
cc_341 N_A_218_424#_M1006_g N_VGND_c_687_n 0.00383152f $X=3.395 $Y=0.74 $X2=0
+ $Y2=0
cc_342 N_A_218_424#_c_382_n N_VGND_c_687_n 3.38697e-19 $X=2.755 $Y=0.84 $X2=0
+ $Y2=0
cc_343 N_A_218_424#_c_345_n N_VGND_c_688_n 0.00434272f $X=3.86 $Y=1.185 $X2=0
+ $Y2=0
cc_344 N_A_218_424#_c_348_n N_VGND_c_688_n 0.00383152f $X=4.29 $Y=1.185 $X2=0
+ $Y2=0
cc_345 N_A_218_424#_M1000_g N_VGND_c_692_n 0.00706821f $X=2.955 $Y=0.74 $X2=0
+ $Y2=0
cc_346 N_A_218_424#_M1006_g N_VGND_c_692_n 0.0075764f $X=3.395 $Y=0.74 $X2=0
+ $Y2=0
cc_347 N_A_218_424#_c_345_n N_VGND_c_692_n 0.00821408f $X=3.86 $Y=1.185 $X2=0
+ $Y2=0
cc_348 N_A_218_424#_c_348_n N_VGND_c_692_n 0.0075754f $X=4.29 $Y=1.185 $X2=0
+ $Y2=0
cc_349 N_A_218_424#_c_382_n N_VGND_c_692_n 0.00675954f $X=2.755 $Y=0.84 $X2=0
+ $Y2=0
cc_350 N_A_218_424#_c_382_n N_A_233_74#_M1014_s 0.00423148f $X=2.755 $Y=0.84
+ $X2=0 $Y2=0
cc_351 N_A_218_424#_M1005_d N_A_233_74#_c_751_n 0.00168037f $X=1.665 $Y=0.37
+ $X2=0 $Y2=0
cc_352 N_A_218_424#_c_382_n N_A_233_74#_c_751_n 0.037476f $X=2.755 $Y=0.84 $X2=0
+ $Y2=0
cc_353 N_VPWR_c_524_n N_X_c_608_n 0.0443204f $X=2.73 $Y=2.465 $X2=0 $Y2=0
cc_354 N_VPWR_c_525_n N_X_c_608_n 0.0534396f $X=3.63 $Y=2.325 $X2=0 $Y2=0
cc_355 N_VPWR_c_529_n N_X_c_608_n 0.00749631f $X=3.465 $Y=3.33 $X2=0 $Y2=0
cc_356 N_VPWR_c_519_n N_X_c_608_n 0.0062048f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_357 N_VPWR_M1004_d N_X_c_609_n 0.00197722f $X=3.48 $Y=1.84 $X2=0 $Y2=0
cc_358 N_VPWR_c_525_n N_X_c_609_n 0.0171813f $X=3.63 $Y=2.325 $X2=0 $Y2=0
cc_359 N_VPWR_c_525_n N_X_c_611_n 0.0534396f $X=3.63 $Y=2.325 $X2=0 $Y2=0
cc_360 N_VPWR_c_527_n N_X_c_611_n 0.0644806f $X=4.53 $Y=1.985 $X2=0 $Y2=0
cc_361 N_VPWR_c_530_n N_X_c_611_n 0.00749631f $X=4.365 $Y=3.33 $X2=0 $Y2=0
cc_362 N_VPWR_c_519_n N_X_c_611_n 0.0062048f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_363 N_VPWR_c_527_n N_X_c_603_n 0.0279882f $X=4.53 $Y=1.985 $X2=0 $Y2=0
cc_364 N_VPWR_c_527_n N_X_c_653_n 0.0124177f $X=4.53 $Y=1.985 $X2=0 $Y2=0
cc_365 N_X_c_599_n N_VGND_M1006_d 0.00307253f $X=3.91 $Y=1.065 $X2=0 $Y2=0
cc_366 N_X_c_602_n N_VGND_M1013_d 0.00325695f $X=4.445 $Y=1.065 $X2=0 $Y2=0
cc_367 N_X_c_598_n N_VGND_c_682_n 0.0156353f $X=3.18 $Y=0.515 $X2=0 $Y2=0
cc_368 N_X_c_598_n N_VGND_c_683_n 0.0164868f $X=3.18 $Y=0.515 $X2=0 $Y2=0
cc_369 N_X_c_599_n N_VGND_c_683_n 0.015373f $X=3.91 $Y=1.065 $X2=0 $Y2=0
cc_370 N_X_c_601_n N_VGND_c_683_n 0.0286138f $X=4.075 $Y=0.515 $X2=0 $Y2=0
cc_371 N_X_c_601_n N_VGND_c_685_n 0.017215f $X=4.075 $Y=0.515 $X2=0 $Y2=0
cc_372 N_X_c_602_n N_VGND_c_685_n 0.023862f $X=4.445 $Y=1.065 $X2=0 $Y2=0
cc_373 N_X_c_598_n N_VGND_c_687_n 0.00749631f $X=3.18 $Y=0.515 $X2=0 $Y2=0
cc_374 N_X_c_601_n N_VGND_c_688_n 0.0109942f $X=4.075 $Y=0.515 $X2=0 $Y2=0
cc_375 N_X_c_598_n N_VGND_c_692_n 0.0062048f $X=3.18 $Y=0.515 $X2=0 $Y2=0
cc_376 N_X_c_601_n N_VGND_c_692_n 0.00904371f $X=4.075 $Y=0.515 $X2=0 $Y2=0
cc_377 N_VGND_c_681_n N_A_233_74#_c_750_n 0.0110102f $X=0.875 $Y=0.495 $X2=0
+ $Y2=0
cc_378 N_VGND_c_686_n N_A_233_74#_c_750_n 0.0122168f $X=2.57 $Y=0 $X2=0 $Y2=0
cc_379 N_VGND_c_692_n N_A_233_74#_c_750_n 0.00964373f $X=4.56 $Y=0 $X2=0 $Y2=0
cc_380 N_VGND_c_682_n N_A_233_74#_c_751_n 0.0118255f $X=2.735 $Y=0.5 $X2=0 $Y2=0
cc_381 N_VGND_c_686_n N_A_233_74#_c_751_n 0.0401098f $X=2.57 $Y=0 $X2=0 $Y2=0
cc_382 N_VGND_c_692_n N_A_233_74#_c_751_n 0.0321234f $X=4.56 $Y=0 $X2=0 $Y2=0
