* File: sky130_fd_sc_ls__a21oi_1.pex.spice
* Created: Wed Sep  2 10:48:48 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__A21OI_1%A2 1 3 4 6 7
c22 7 0 1.40395e-19 $X=0.24 $Y=1.295
r23 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.385 $X2=0.27 $Y2=1.385
r24 7 11 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.27 $Y=1.295 $X2=0.27
+ $Y2=1.385
r25 4 10 38.924 $w=3.61e-07 $l=2.33345e-07 $layer=POLY_cond $X=0.51 $Y=1.22
+ $X2=0.345 $Y2=1.385
r26 4 6 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.51 $Y=1.22 $X2=0.51
+ $Y2=0.74
r27 1 10 67.6304 $w=3.61e-07 $l=4.48776e-07 $layer=POLY_cond $X=0.495 $Y=1.765
+ $X2=0.345 $Y2=1.385
r28 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.495 $Y=1.765
+ $X2=0.495 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__A21OI_1%A1 3 5 7 8 12
c33 5 0 1.40395e-19 $X=0.975 $Y=1.765
r34 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.96
+ $Y=1.515 $X2=0.96 $Y2=1.515
r35 8 12 6.43224 $w=4.28e-07 $l=2.4e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=0.96 $Y2=1.565
r36 5 11 52.2586 $w=2.99e-07 $l=2.57391e-07 $layer=POLY_cond $X=0.975 $Y=1.765
+ $X2=0.96 $Y2=1.515
r37 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.975 $Y=1.765
+ $X2=0.975 $Y2=2.4
r38 1 11 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=0.87 $Y=1.35
+ $X2=0.96 $Y2=1.515
r39 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.87 $Y=1.35 $X2=0.87
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__A21OI_1%B1 1 3 4 6 7
r24 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.65
+ $Y=1.385 $X2=1.65 $Y2=1.385
r25 7 11 4.06745 $w=2.53e-07 $l=9e-08 $layer=LI1_cond $X=1.687 $Y=1.295
+ $X2=1.687 $Y2=1.385
r26 4 10 67.6304 $w=3.61e-07 $l=4.48776e-07 $layer=POLY_cond $X=1.425 $Y=1.765
+ $X2=1.575 $Y2=1.385
r27 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.425 $Y=1.765
+ $X2=1.425 $Y2=2.4
r28 1 10 38.924 $w=3.61e-07 $l=2.33345e-07 $layer=POLY_cond $X=1.41 $Y=1.22
+ $X2=1.575 $Y2=1.385
r29 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.41 $Y=1.22 $X2=1.41
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__A21OI_1%A_29_368# 1 2 7 9 11 18
r25 12 16 3.62238 $w=2.45e-07 $l=2.01879e-07 $layer=LI1_cond $X=0.435 $Y=2.107
+ $X2=0.27 $Y2=2.025
r26 11 18 18.9889 $w=2.45e-07 $l=3.67e-07 $layer=LI1_cond $X=0.833 $Y=2.107
+ $X2=1.2 $Y2=2.107
r27 11 12 18.7213 $w=2.43e-07 $l=3.98e-07 $layer=LI1_cond $X=0.833 $Y=2.107
+ $X2=0.435 $Y2=2.107
r28 7 16 3.2704 $w=2.95e-07 $l=2.13811e-07 $layer=LI1_cond $X=0.252 $Y=2.23
+ $X2=0.27 $Y2=2.025
r29 7 9 6.6412 $w=2.93e-07 $l=1.7e-07 $layer=LI1_cond $X=0.252 $Y=2.23 $X2=0.252
+ $Y2=2.4
r30 2 18 300 $w=1.7e-07 $l=4.53845e-07 $layer=licon1_PDIFF $count=2 $X=1.05
+ $Y=1.84 $X2=1.2 $Y2=2.225
r31 1 16 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.84 $X2=0.27 $Y2=1.985
r32 1 9 300 $w=1.7e-07 $l=6.19354e-07 $layer=licon1_PDIFF $count=2 $X=0.145
+ $Y=1.84 $X2=0.27 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__A21OI_1%VPWR 1 6 8 10 17 18 21
r25 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r26 17 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r27 15 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.9 $Y=3.33
+ $X2=0.735 $Y2=3.33
r28 15 17 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=0.9 $Y=3.33 $X2=1.68
+ $Y2=3.33
r29 13 22 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r30 12 13 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r31 10 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.57 $Y=3.33
+ $X2=0.735 $Y2=3.33
r32 10 12 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.57 $Y=3.33
+ $X2=0.24 $Y2=3.33
r33 8 18 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=1.68 $Y2=3.33
r34 8 22 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=0.72 $Y2=3.33
r35 4 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.735 $Y=3.245
+ $X2=0.735 $Y2=3.33
r36 4 6 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=0.735 $Y=3.245
+ $X2=0.735 $Y2=2.485
r37 1 6 300 $w=1.7e-07 $l=7.22807e-07 $layer=licon1_PDIFF $count=2 $X=0.57
+ $Y=1.84 $X2=0.735 $Y2=2.485
.ends

.subckt PM_SKY130_FD_SC_LS__A21OI_1%Y 1 2 9 12 13 14 16 18 19 20
r36 19 20 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=1.69 $Y=2.405
+ $X2=1.69 $Y2=2.775
r37 18 19 19.361 $w=2.48e-07 $l=4.2e-07 $layer=LI1_cond $X=1.69 $Y=1.985
+ $X2=1.69 $Y2=2.405
r38 17 18 4.37928 $w=2.48e-07 $l=9.5e-08 $layer=LI1_cond $X=1.69 $Y=1.89
+ $X2=1.69 $Y2=1.985
r39 15 16 8.69455 $w=3.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.155 $Y=1.01
+ $X2=1.155 $Y2=1.18
r40 13 17 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.565 $Y=1.805
+ $X2=1.69 $Y2=1.89
r41 13 14 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.565 $Y=1.805
+ $X2=1.39 $Y2=1.805
r42 12 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.305 $Y=1.72
+ $X2=1.39 $Y2=1.805
r43 12 16 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=1.305 $Y=1.72
+ $X2=1.305 $Y2=1.18
r44 9 15 15.4178 $w=3.68e-07 $l=4.95e-07 $layer=LI1_cond $X=1.105 $Y=0.515
+ $X2=1.105 $Y2=1.01
r45 2 20 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.5
+ $Y=1.84 $X2=1.65 $Y2=2.815
r46 2 18 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.5
+ $Y=1.84 $X2=1.65 $Y2=1.985
r47 1 9 91 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=2 $X=0.945
+ $Y=0.37 $X2=1.105 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__A21OI_1%VGND 1 2 7 9 11 13 15 17 27
r24 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r25 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r26 21 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r27 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r28 18 23 4.70058 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=0.46 $Y=0 $X2=0.23
+ $Y2=0
r29 18 20 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=0.46 $Y=0 $X2=1.2
+ $Y2=0
r30 17 26 3.82794 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=1.56 $Y=0 $X2=1.74
+ $Y2=0
r31 17 20 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=1.56 $Y=0 $X2=1.2
+ $Y2=0
r32 15 21 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=1.2
+ $Y2=0
r33 15 24 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=0.24
+ $Y2=0
r34 11 26 3.18995 $w=2.3e-07 $l=1.12916e-07 $layer=LI1_cond $X=1.675 $Y=0.085
+ $X2=1.74 $Y2=0
r35 11 13 21.5457 $w=2.28e-07 $l=4.3e-07 $layer=LI1_cond $X=1.675 $Y=0.085
+ $X2=1.675 $Y2=0.515
r36 7 23 3.0656 $w=3.3e-07 $l=1.12916e-07 $layer=LI1_cond $X=0.295 $Y=0.085
+ $X2=0.23 $Y2=0
r37 7 9 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.295 $Y=0.085
+ $X2=0.295 $Y2=0.515
r38 2 13 91 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=2 $X=1.485
+ $Y=0.37 $X2=1.645 $Y2=0.515
r39 1 9 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.17
+ $Y=0.37 $X2=0.295 $Y2=0.515
.ends

