* File: sky130_fd_sc_ls__nand4_2.pxi.spice
* Created: Wed Sep  2 11:12:54 2020
* 
x_PM_SKY130_FD_SC_LS__NAND4_2%D N_D_M1001_g N_D_c_84_n N_D_M1006_g N_D_c_85_n
+ N_D_M1009_g N_D_M1011_g D D N_D_c_82_n N_D_c_83_n
+ PM_SKY130_FD_SC_LS__NAND4_2%D
x_PM_SKY130_FD_SC_LS__NAND4_2%C N_C_M1007_g N_C_c_127_n N_C_M1000_g N_C_M1013_g
+ N_C_c_128_n N_C_M1014_g C C N_C_c_124_n N_C_c_125_n N_C_c_126_n
+ PM_SKY130_FD_SC_LS__NAND4_2%C
x_PM_SKY130_FD_SC_LS__NAND4_2%B N_B_c_180_n N_B_M1002_g N_B_M1004_g N_B_c_181_n
+ N_B_M1005_g N_B_M1012_g B B N_B_c_179_n PM_SKY130_FD_SC_LS__NAND4_2%B
x_PM_SKY130_FD_SC_LS__NAND4_2%A N_A_c_234_n N_A_M1003_g N_A_M1010_g N_A_c_235_n
+ N_A_M1008_g N_A_M1015_g A N_A_c_232_n N_A_c_233_n
+ PM_SKY130_FD_SC_LS__NAND4_2%A
x_PM_SKY130_FD_SC_LS__NAND4_2%VPWR N_VPWR_M1006_s N_VPWR_M1009_s N_VPWR_M1014_s
+ N_VPWR_M1005_s N_VPWR_M1008_s N_VPWR_c_279_n N_VPWR_c_280_n N_VPWR_c_281_n
+ N_VPWR_c_282_n N_VPWR_c_283_n N_VPWR_c_284_n N_VPWR_c_285_n N_VPWR_c_286_n
+ N_VPWR_c_287_n N_VPWR_c_288_n VPWR N_VPWR_c_289_n N_VPWR_c_290_n
+ N_VPWR_c_291_n N_VPWR_c_292_n N_VPWR_c_278_n PM_SKY130_FD_SC_LS__NAND4_2%VPWR
x_PM_SKY130_FD_SC_LS__NAND4_2%Y N_Y_M1010_d N_Y_M1006_d N_Y_M1000_d N_Y_M1002_d
+ N_Y_M1003_d N_Y_c_358_n N_Y_c_352_n N_Y_c_360_n N_Y_c_353_n N_Y_c_365_n
+ N_Y_c_354_n N_Y_c_375_n N_Y_c_355_n N_Y_c_386_n N_Y_c_388_n N_Y_c_349_n
+ N_Y_c_350_n N_Y_c_368_n N_Y_c_379_n N_Y_c_396_n Y Y Y
+ PM_SKY130_FD_SC_LS__NAND4_2%Y
x_PM_SKY130_FD_SC_LS__NAND4_2%A_27_74# N_A_27_74#_M1001_d N_A_27_74#_M1011_d
+ N_A_27_74#_M1013_s N_A_27_74#_c_436_n N_A_27_74#_c_437_n N_A_27_74#_c_438_n
+ N_A_27_74#_c_439_n N_A_27_74#_c_440_n N_A_27_74#_c_441_n
+ PM_SKY130_FD_SC_LS__NAND4_2%A_27_74#
x_PM_SKY130_FD_SC_LS__NAND4_2%VGND N_VGND_M1001_s N_VGND_c_473_n VGND
+ N_VGND_c_474_n N_VGND_c_475_n N_VGND_c_476_n N_VGND_c_477_n
+ PM_SKY130_FD_SC_LS__NAND4_2%VGND
x_PM_SKY130_FD_SC_LS__NAND4_2%A_304_74# N_A_304_74#_M1007_d N_A_304_74#_M1004_s
+ N_A_304_74#_c_516_n N_A_304_74#_c_514_n N_A_304_74#_c_515_n
+ N_A_304_74#_c_529_n PM_SKY130_FD_SC_LS__NAND4_2%A_304_74#
x_PM_SKY130_FD_SC_LS__NAND4_2%A_515_74# N_A_515_74#_M1004_d N_A_515_74#_M1012_d
+ N_A_515_74#_M1015_s N_A_515_74#_c_544_n N_A_515_74#_c_545_n
+ N_A_515_74#_c_546_n N_A_515_74#_c_547_n N_A_515_74#_c_548_n
+ N_A_515_74#_c_549_n N_A_515_74#_c_550_n PM_SKY130_FD_SC_LS__NAND4_2%A_515_74#
cc_1 VNB N_D_M1001_g 0.0338822f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_D_M1011_g 0.0242263f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=0.74
cc_3 VNB N_D_c_82_n 0.0192271f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.515
cc_4 VNB N_D_c_83_n 0.039755f $X=-0.19 $Y=-0.245 $X2=1 $Y2=1.557
cc_5 VNB N_C_M1007_g 0.0229341f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_6 VNB N_C_M1013_g 0.0304502f $X=-0.19 $Y=-0.245 $X2=1 $Y2=2.4
cc_7 VNB N_C_c_124_n 0.0341628f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.557
cc_8 VNB N_C_c_125_n 0.0257749f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.557
cc_9 VNB N_C_c_126_n 0.00219487f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.515
cc_10 VNB N_B_M1004_g 0.0304502f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.4
cc_11 VNB N_B_M1012_g 0.0229481f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=0.74
cc_12 VNB B 0.00974538f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_13 VNB N_B_c_179_n 0.0398922f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.515
cc_14 VNB N_A_M1010_g 0.0232431f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.4
cc_15 VNB N_A_M1015_g 0.0264271f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=0.74
cc_16 VNB N_A_c_232_n 0.00111586f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.557
cc_17 VNB N_A_c_233_n 0.0370006f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.515
cc_18 VNB N_VPWR_c_278_n 0.203486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_Y_c_349_n 0.0129996f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_Y_c_350_n 0.00289607f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB Y 0.0244237f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_27_74#_c_436_n 0.0277086f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=0.74
cc_23 VNB N_A_27_74#_c_437_n 0.0121125f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_27_74#_c_438_n 0.0104987f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_25 VNB N_A_27_74#_c_439_n 0.0073244f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.557
cc_26 VNB N_A_27_74#_c_440_n 0.00213827f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.557
cc_27 VNB N_A_27_74#_c_441_n 0.00465049f $X=-0.19 $Y=-0.245 $X2=1 $Y2=1.557
cc_28 VNB N_VGND_c_473_n 0.00662552f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.4
cc_29 VNB N_VGND_c_474_n 0.0191515f $X=-0.19 $Y=-0.245 $X2=1 $Y2=2.4
cc_30 VNB N_VGND_c_475_n 0.0928206f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.557
cc_31 VNB N_VGND_c_476_n 0.28314f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.557
cc_32 VNB N_VGND_c_477_n 0.00617641f $X=-0.19 $Y=-0.245 $X2=1 $Y2=1.557
cc_33 VNB N_A_304_74#_c_514_n 0.0269092f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=1.35
cc_34 VNB N_A_304_74#_c_515_n 0.00229834f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=0.74
cc_35 VNB N_A_515_74#_c_544_n 0.00437839f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=0.74
cc_36 VNB N_A_515_74#_c_545_n 0.0026202f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_515_74#_c_546_n 0.0038714f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_38 VNB N_A_515_74#_c_547_n 0.00228245f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_515_74#_c_548_n 0.0127105f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.557
cc_40 VNB N_A_515_74#_c_549_n 0.0167552f $X=-0.19 $Y=-0.245 $X2=1 $Y2=1.557
cc_41 VNB N_A_515_74#_c_550_n 0.00138314f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.565
cc_42 VPB N_D_c_84_n 0.0191345f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.765
cc_43 VPB N_D_c_85_n 0.0156616f $X=-0.19 $Y=1.66 $X2=1 $Y2=1.765
cc_44 VPB N_D_c_82_n 0.0140108f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.515
cc_45 VPB N_D_c_83_n 0.0222326f $X=-0.19 $Y=1.66 $X2=1 $Y2=1.557
cc_46 VPB N_C_c_127_n 0.0164204f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.765
cc_47 VPB N_C_c_128_n 0.0179368f $X=-0.19 $Y=1.66 $X2=1.015 $Y2=0.74
cc_48 VPB N_C_c_124_n 0.020992f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.557
cc_49 VPB N_C_c_125_n 0.0121782f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.557
cc_50 VPB N_C_c_126_n 0.00760803f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.515
cc_51 VPB N_B_c_180_n 0.0177772f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.35
cc_52 VPB N_B_c_181_n 0.0165483f $X=-0.19 $Y=1.66 $X2=1 $Y2=1.765
cc_53 VPB B 0.00788501f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_54 VPB N_B_c_179_n 0.024091f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.515
cc_55 VPB N_A_c_234_n 0.0165945f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.35
cc_56 VPB N_A_c_235_n 0.0172088f $X=-0.19 $Y=1.66 $X2=1 $Y2=1.765
cc_57 VPB N_A_c_232_n 0.00307804f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.557
cc_58 VPB N_A_c_233_n 0.0206484f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.515
cc_59 VPB N_VPWR_c_279_n 0.0121068f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_60 VPB N_VPWR_c_280_n 0.0484283f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_281_n 0.00606947f $X=-0.19 $Y=1.66 $X2=1 $Y2=1.557
cc_62 VPB N_VPWR_c_282_n 0.019013f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.565
cc_63 VPB N_VPWR_c_283_n 0.0125119f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_284_n 0.00900023f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_285_n 0.0139291f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_286_n 0.0335032f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_287_n 0.019013f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_288_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_289_n 0.0172955f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_290_n 0.0177745f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_291_n 0.00615051f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_292_n 0.0109379f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_278_n 0.0683221f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_Y_c_352_n 0.00266762f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_Y_c_353_n 0.00290151f $X=-0.19 $Y=1.66 $X2=1 $Y2=1.557
cc_76 VPB N_Y_c_354_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_Y_c_355_n 0.00247739f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB Y 0.0133105f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 VPB Y 0.0105887f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 N_D_M1011_g N_C_M1007_g 0.0129244f $X=1.015 $Y=0.74 $X2=0 $Y2=0
cc_81 N_D_c_85_n N_C_c_127_n 0.0212394f $X=1 $Y=1.765 $X2=0 $Y2=0
cc_82 N_D_c_82_n N_C_c_124_n 0.00184507f $X=0.925 $Y=1.515 $X2=0 $Y2=0
cc_83 N_D_c_83_n N_C_c_124_n 0.0235065f $X=1 $Y=1.557 $X2=0 $Y2=0
cc_84 N_D_c_82_n N_C_c_126_n 0.02073f $X=0.925 $Y=1.515 $X2=0 $Y2=0
cc_85 N_D_c_83_n N_C_c_126_n 4.9167e-19 $X=1 $Y=1.557 $X2=0 $Y2=0
cc_86 N_D_c_84_n N_VPWR_c_280_n 0.0153782f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_87 N_D_c_85_n N_VPWR_c_280_n 5.53867e-19 $X=1 $Y=1.765 $X2=0 $Y2=0
cc_88 N_D_c_82_n N_VPWR_c_280_n 0.0259599f $X=0.925 $Y=1.515 $X2=0 $Y2=0
cc_89 N_D_c_84_n N_VPWR_c_281_n 4.86642e-19 $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_90 N_D_c_85_n N_VPWR_c_281_n 0.00978105f $X=1 $Y=1.765 $X2=0 $Y2=0
cc_91 N_D_c_84_n N_VPWR_c_289_n 0.00413917f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_92 N_D_c_85_n N_VPWR_c_289_n 0.00444681f $X=1 $Y=1.765 $X2=0 $Y2=0
cc_93 N_D_c_84_n N_VPWR_c_278_n 0.00818099f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_94 N_D_c_85_n N_VPWR_c_278_n 0.00878088f $X=1 $Y=1.765 $X2=0 $Y2=0
cc_95 N_D_c_82_n N_Y_c_358_n 0.0216748f $X=0.925 $Y=1.515 $X2=0 $Y2=0
cc_96 N_D_c_83_n N_Y_c_358_n 0.00153038f $X=1 $Y=1.557 $X2=0 $Y2=0
cc_97 N_D_c_85_n N_Y_c_360_n 0.0130991f $X=1 $Y=1.765 $X2=0 $Y2=0
cc_98 N_D_c_82_n N_Y_c_360_n 0.012644f $X=0.925 $Y=1.515 $X2=0 $Y2=0
cc_99 N_D_M1001_g N_A_27_74#_c_436_n 0.0101727f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_100 N_D_M1011_g N_A_27_74#_c_436_n 9.49764e-19 $X=1.015 $Y=0.74 $X2=0 $Y2=0
cc_101 N_D_M1001_g N_A_27_74#_c_437_n 0.0116427f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_102 N_D_M1011_g N_A_27_74#_c_437_n 0.0138917f $X=1.015 $Y=0.74 $X2=0 $Y2=0
cc_103 N_D_c_82_n N_A_27_74#_c_437_n 0.0484156f $X=0.925 $Y=1.515 $X2=0 $Y2=0
cc_104 N_D_c_83_n N_A_27_74#_c_437_n 0.0042599f $X=1 $Y=1.557 $X2=0 $Y2=0
cc_105 N_D_M1001_g N_A_27_74#_c_438_n 0.00214722f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_106 N_D_c_82_n N_A_27_74#_c_438_n 0.0286342f $X=0.925 $Y=1.515 $X2=0 $Y2=0
cc_107 N_D_M1011_g N_A_27_74#_c_440_n 9.95577e-19 $X=1.015 $Y=0.74 $X2=0 $Y2=0
cc_108 N_D_M1001_g N_VGND_c_473_n 0.005861f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_109 N_D_M1011_g N_VGND_c_473_n 0.00844304f $X=1.015 $Y=0.74 $X2=0 $Y2=0
cc_110 N_D_M1001_g N_VGND_c_474_n 0.00434272f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_111 N_D_M1011_g N_VGND_c_475_n 0.00444681f $X=1.015 $Y=0.74 $X2=0 $Y2=0
cc_112 N_D_M1001_g N_VGND_c_476_n 0.00824548f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_113 N_D_M1011_g N_VGND_c_476_n 0.00877616f $X=1.015 $Y=0.74 $X2=0 $Y2=0
cc_114 N_C_c_128_n N_B_c_180_n 0.0103933f $X=1.96 $Y=1.765 $X2=-0.19 $Y2=-0.245
cc_115 N_C_c_125_n B 4.13265e-19 $X=2.275 $Y=1.515 $X2=0 $Y2=0
cc_116 N_C_c_126_n B 0.0279555f $X=2.275 $Y=1.515 $X2=0 $Y2=0
cc_117 N_C_c_124_n N_B_c_179_n 0.00104119f $X=2.05 $Y=1.515 $X2=0 $Y2=0
cc_118 N_C_c_125_n N_B_c_179_n 0.0183161f $X=2.275 $Y=1.515 $X2=0 $Y2=0
cc_119 N_C_c_126_n N_B_c_179_n 8.49051e-19 $X=2.275 $Y=1.515 $X2=0 $Y2=0
cc_120 N_C_c_127_n N_VPWR_c_281_n 0.00345866f $X=1.49 $Y=1.765 $X2=0 $Y2=0
cc_121 N_C_c_127_n N_VPWR_c_282_n 0.00461464f $X=1.49 $Y=1.765 $X2=0 $Y2=0
cc_122 N_C_c_128_n N_VPWR_c_282_n 0.00445602f $X=1.96 $Y=1.765 $X2=0 $Y2=0
cc_123 N_C_c_128_n N_VPWR_c_283_n 0.00404718f $X=1.96 $Y=1.765 $X2=0 $Y2=0
cc_124 N_C_c_127_n N_VPWR_c_278_n 0.00908452f $X=1.49 $Y=1.765 $X2=0 $Y2=0
cc_125 N_C_c_128_n N_VPWR_c_278_n 0.00859794f $X=1.96 $Y=1.765 $X2=0 $Y2=0
cc_126 N_C_c_127_n N_Y_c_360_n 0.0137341f $X=1.49 $Y=1.765 $X2=0 $Y2=0
cc_127 N_C_c_126_n N_Y_c_360_n 0.0100328f $X=2.275 $Y=1.515 $X2=0 $Y2=0
cc_128 N_C_c_128_n N_Y_c_353_n 0.0146573f $X=1.96 $Y=1.765 $X2=0 $Y2=0
cc_129 N_C_c_128_n N_Y_c_365_n 0.0132683f $X=1.96 $Y=1.765 $X2=0 $Y2=0
cc_130 N_C_c_125_n N_Y_c_365_n 0.00204715f $X=2.275 $Y=1.515 $X2=0 $Y2=0
cc_131 N_C_c_126_n N_Y_c_365_n 0.0400047f $X=2.275 $Y=1.515 $X2=0 $Y2=0
cc_132 N_C_c_128_n N_Y_c_368_n 4.27055e-19 $X=1.96 $Y=1.765 $X2=0 $Y2=0
cc_133 N_C_c_124_n N_Y_c_368_n 0.00156348f $X=2.05 $Y=1.515 $X2=0 $Y2=0
cc_134 N_C_c_126_n N_Y_c_368_n 0.0241316f $X=2.275 $Y=1.515 $X2=0 $Y2=0
cc_135 N_C_M1007_g N_A_27_74#_c_437_n 5.7448e-19 $X=1.445 $Y=0.74 $X2=0 $Y2=0
cc_136 N_C_M1007_g N_A_27_74#_c_439_n 0.0120041f $X=1.445 $Y=0.74 $X2=0 $Y2=0
cc_137 N_C_M1013_g N_A_27_74#_c_439_n 0.0123342f $X=1.875 $Y=0.74 $X2=0 $Y2=0
cc_138 N_C_M1007_g N_VGND_c_475_n 0.00278271f $X=1.445 $Y=0.74 $X2=0 $Y2=0
cc_139 N_C_M1013_g N_VGND_c_475_n 0.00278271f $X=1.875 $Y=0.74 $X2=0 $Y2=0
cc_140 N_C_M1007_g N_VGND_c_476_n 0.00353526f $X=1.445 $Y=0.74 $X2=0 $Y2=0
cc_141 N_C_M1013_g N_VGND_c_476_n 0.00358427f $X=1.875 $Y=0.74 $X2=0 $Y2=0
cc_142 N_C_M1007_g N_A_304_74#_c_516_n 0.00546155f $X=1.445 $Y=0.74 $X2=0 $Y2=0
cc_143 N_C_M1013_g N_A_304_74#_c_516_n 0.0111175f $X=1.875 $Y=0.74 $X2=0 $Y2=0
cc_144 N_C_M1013_g N_A_304_74#_c_514_n 0.0110459f $X=1.875 $Y=0.74 $X2=0 $Y2=0
cc_145 N_C_c_124_n N_A_304_74#_c_514_n 0.011317f $X=2.05 $Y=1.515 $X2=0 $Y2=0
cc_146 N_C_c_126_n N_A_304_74#_c_514_n 0.046634f $X=2.275 $Y=1.515 $X2=0 $Y2=0
cc_147 N_C_M1007_g N_A_304_74#_c_515_n 0.00359492f $X=1.445 $Y=0.74 $X2=0 $Y2=0
cc_148 N_C_M1013_g N_A_304_74#_c_515_n 0.00223461f $X=1.875 $Y=0.74 $X2=0 $Y2=0
cc_149 N_C_c_124_n N_A_304_74#_c_515_n 0.00231547f $X=2.05 $Y=1.515 $X2=0 $Y2=0
cc_150 N_C_c_126_n N_A_304_74#_c_515_n 0.0277843f $X=2.275 $Y=1.515 $X2=0 $Y2=0
cc_151 N_C_M1013_g N_A_515_74#_c_546_n 6.36929e-19 $X=1.875 $Y=0.74 $X2=0 $Y2=0
cc_152 N_B_c_181_n N_A_c_234_n 0.0312563f $X=3.22 $Y=1.765 $X2=-0.19 $Y2=-0.245
cc_153 B N_A_c_234_n 4.52698e-19 $X=3.515 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_154 N_B_M1012_g N_A_M1010_g 0.0169947f $X=3.365 $Y=0.74 $X2=0 $Y2=0
cc_155 B N_A_c_232_n 0.0360052f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_156 N_B_c_179_n N_A_c_232_n 2.12629e-19 $X=3.275 $Y=1.515 $X2=0 $Y2=0
cc_157 B N_A_c_233_n 0.00589605f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_158 N_B_c_179_n N_A_c_233_n 0.0193938f $X=3.275 $Y=1.515 $X2=0 $Y2=0
cc_159 N_B_c_180_n N_VPWR_c_283_n 0.00404718f $X=2.77 $Y=1.765 $X2=0 $Y2=0
cc_160 N_B_c_181_n N_VPWR_c_284_n 0.00747273f $X=3.22 $Y=1.765 $X2=0 $Y2=0
cc_161 N_B_c_180_n N_VPWR_c_287_n 0.00445602f $X=2.77 $Y=1.765 $X2=0 $Y2=0
cc_162 N_B_c_181_n N_VPWR_c_287_n 0.00445602f $X=3.22 $Y=1.765 $X2=0 $Y2=0
cc_163 N_B_c_180_n N_VPWR_c_278_n 0.00859604f $X=2.77 $Y=1.765 $X2=0 $Y2=0
cc_164 N_B_c_181_n N_VPWR_c_278_n 0.00857899f $X=3.22 $Y=1.765 $X2=0 $Y2=0
cc_165 N_B_c_180_n N_Y_c_365_n 0.0132683f $X=2.77 $Y=1.765 $X2=0 $Y2=0
cc_166 B N_Y_c_365_n 0.0104662f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_167 N_B_c_180_n N_Y_c_354_n 0.0146845f $X=2.77 $Y=1.765 $X2=0 $Y2=0
cc_168 N_B_c_181_n N_Y_c_354_n 0.0103688f $X=3.22 $Y=1.765 $X2=0 $Y2=0
cc_169 N_B_c_181_n N_Y_c_375_n 0.0124941f $X=3.22 $Y=1.765 $X2=0 $Y2=0
cc_170 B N_Y_c_375_n 0.0390626f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_171 N_B_c_179_n N_Y_c_375_n 6.23858e-19 $X=3.275 $Y=1.515 $X2=0 $Y2=0
cc_172 N_B_c_181_n N_Y_c_355_n 7.75925e-19 $X=3.22 $Y=1.765 $X2=0 $Y2=0
cc_173 N_B_c_180_n N_Y_c_379_n 4.27055e-19 $X=2.77 $Y=1.765 $X2=0 $Y2=0
cc_174 N_B_c_181_n N_Y_c_379_n 4.27055e-19 $X=3.22 $Y=1.765 $X2=0 $Y2=0
cc_175 B N_Y_c_379_n 0.0237598f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_176 N_B_c_179_n N_Y_c_379_n 0.00143667f $X=3.275 $Y=1.515 $X2=0 $Y2=0
cc_177 N_B_M1004_g N_A_27_74#_c_439_n 7.14966e-19 $X=2.935 $Y=0.74 $X2=0 $Y2=0
cc_178 N_B_M1004_g N_VGND_c_475_n 0.00278271f $X=2.935 $Y=0.74 $X2=0 $Y2=0
cc_179 N_B_M1012_g N_VGND_c_475_n 0.00278271f $X=3.365 $Y=0.74 $X2=0 $Y2=0
cc_180 N_B_M1004_g N_VGND_c_476_n 0.00358427f $X=2.935 $Y=0.74 $X2=0 $Y2=0
cc_181 N_B_M1012_g N_VGND_c_476_n 0.00353526f $X=3.365 $Y=0.74 $X2=0 $Y2=0
cc_182 N_B_M1004_g N_A_304_74#_c_514_n 0.0138209f $X=2.935 $Y=0.74 $X2=0 $Y2=0
cc_183 N_B_M1012_g N_A_304_74#_c_514_n 0.00448299f $X=3.365 $Y=0.74 $X2=0 $Y2=0
cc_184 B N_A_304_74#_c_514_n 0.0504811f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_185 N_B_c_179_n N_A_304_74#_c_514_n 0.00720209f $X=3.275 $Y=1.515 $X2=0 $Y2=0
cc_186 N_B_M1004_g N_A_304_74#_c_529_n 0.0097752f $X=2.935 $Y=0.74 $X2=0 $Y2=0
cc_187 N_B_M1012_g N_A_304_74#_c_529_n 0.00405156f $X=3.365 $Y=0.74 $X2=0 $Y2=0
cc_188 N_B_M1004_g N_A_515_74#_c_545_n 0.0122639f $X=2.935 $Y=0.74 $X2=0 $Y2=0
cc_189 N_B_M1012_g N_A_515_74#_c_545_n 0.012345f $X=3.365 $Y=0.74 $X2=0 $Y2=0
cc_190 N_B_M1012_g N_A_515_74#_c_547_n 3.98786e-19 $X=3.365 $Y=0.74 $X2=0 $Y2=0
cc_191 B N_A_515_74#_c_547_n 0.0141398f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_192 N_A_c_234_n N_VPWR_c_284_n 0.00592249f $X=3.78 $Y=1.765 $X2=0 $Y2=0
cc_193 N_A_c_234_n N_VPWR_c_286_n 5.10274e-19 $X=3.78 $Y=1.765 $X2=0 $Y2=0
cc_194 N_A_c_235_n N_VPWR_c_286_n 0.0112376f $X=4.23 $Y=1.765 $X2=0 $Y2=0
cc_195 N_A_c_234_n N_VPWR_c_290_n 0.00445602f $X=3.78 $Y=1.765 $X2=0 $Y2=0
cc_196 N_A_c_235_n N_VPWR_c_290_n 0.00429299f $X=4.23 $Y=1.765 $X2=0 $Y2=0
cc_197 N_A_c_234_n N_VPWR_c_278_n 0.00858123f $X=3.78 $Y=1.765 $X2=0 $Y2=0
cc_198 N_A_c_235_n N_VPWR_c_278_n 0.00847721f $X=4.23 $Y=1.765 $X2=0 $Y2=0
cc_199 N_A_c_234_n N_Y_c_354_n 9.0208e-19 $X=3.78 $Y=1.765 $X2=0 $Y2=0
cc_200 N_A_c_234_n N_Y_c_375_n 0.0162588f $X=3.78 $Y=1.765 $X2=0 $Y2=0
cc_201 N_A_c_234_n N_Y_c_355_n 0.00985127f $X=3.78 $Y=1.765 $X2=0 $Y2=0
cc_202 N_A_M1010_g N_Y_c_386_n 0.00405156f $X=3.795 $Y=0.74 $X2=0 $Y2=0
cc_203 N_A_M1015_g N_Y_c_386_n 0.00885725f $X=4.245 $Y=0.74 $X2=0 $Y2=0
cc_204 N_A_c_235_n N_Y_c_388_n 0.0182918f $X=4.23 $Y=1.765 $X2=0 $Y2=0
cc_205 N_A_c_232_n N_Y_c_388_n 0.00564925f $X=4.05 $Y=1.515 $X2=0 $Y2=0
cc_206 N_A_M1015_g N_Y_c_349_n 0.0148503f $X=4.245 $Y=0.74 $X2=0 $Y2=0
cc_207 N_A_c_232_n N_Y_c_349_n 0.00282611f $X=4.05 $Y=1.515 $X2=0 $Y2=0
cc_208 N_A_M1010_g N_Y_c_350_n 0.00543662f $X=3.795 $Y=0.74 $X2=0 $Y2=0
cc_209 N_A_M1015_g N_Y_c_350_n 0.00223195f $X=4.245 $Y=0.74 $X2=0 $Y2=0
cc_210 N_A_c_232_n N_Y_c_350_n 0.0244451f $X=4.05 $Y=1.515 $X2=0 $Y2=0
cc_211 N_A_c_233_n N_Y_c_350_n 9.25948e-19 $X=4.23 $Y=1.557 $X2=0 $Y2=0
cc_212 N_A_c_234_n N_Y_c_396_n 0.00158578f $X=3.78 $Y=1.765 $X2=0 $Y2=0
cc_213 N_A_c_232_n N_Y_c_396_n 0.0188362f $X=4.05 $Y=1.515 $X2=0 $Y2=0
cc_214 N_A_c_233_n N_Y_c_396_n 0.00132932f $X=4.23 $Y=1.557 $X2=0 $Y2=0
cc_215 N_A_c_235_n Y 0.0065067f $X=4.23 $Y=1.765 $X2=0 $Y2=0
cc_216 N_A_M1015_g Y 0.0173098f $X=4.245 $Y=0.74 $X2=0 $Y2=0
cc_217 N_A_c_232_n Y 0.0263509f $X=4.05 $Y=1.515 $X2=0 $Y2=0
cc_218 N_A_M1010_g N_VGND_c_475_n 0.00278271f $X=3.795 $Y=0.74 $X2=0 $Y2=0
cc_219 N_A_M1015_g N_VGND_c_475_n 0.00278271f $X=4.245 $Y=0.74 $X2=0 $Y2=0
cc_220 N_A_M1010_g N_VGND_c_476_n 0.00353723f $X=3.795 $Y=0.74 $X2=0 $Y2=0
cc_221 N_A_M1015_g N_VGND_c_476_n 0.00353836f $X=4.245 $Y=0.74 $X2=0 $Y2=0
cc_222 N_A_M1010_g N_A_515_74#_c_547_n 3.98786e-19 $X=3.795 $Y=0.74 $X2=0 $Y2=0
cc_223 N_A_M1010_g N_A_515_74#_c_548_n 0.012465f $X=3.795 $Y=0.74 $X2=0 $Y2=0
cc_224 N_A_M1015_g N_A_515_74#_c_548_n 0.0121365f $X=4.245 $Y=0.74 $X2=0 $Y2=0
cc_225 N_VPWR_c_280_n N_Y_c_352_n 0.0309446f $X=0.28 $Y=2.035 $X2=0 $Y2=0
cc_226 N_VPWR_c_281_n N_Y_c_352_n 0.0266551f $X=1.235 $Y=2.41 $X2=0 $Y2=0
cc_227 N_VPWR_c_289_n N_Y_c_352_n 0.0117353f $X=1.07 $Y=3.33 $X2=0 $Y2=0
cc_228 N_VPWR_c_278_n N_Y_c_352_n 0.00971347f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_229 N_VPWR_M1009_s N_Y_c_360_n 0.0110256f $X=1.075 $Y=1.84 $X2=0 $Y2=0
cc_230 N_VPWR_c_281_n N_Y_c_360_n 0.0186496f $X=1.235 $Y=2.41 $X2=0 $Y2=0
cc_231 N_VPWR_c_281_n N_Y_c_353_n 0.00158095f $X=1.235 $Y=2.41 $X2=0 $Y2=0
cc_232 N_VPWR_c_282_n N_Y_c_353_n 0.0145938f $X=2.08 $Y=3.33 $X2=0 $Y2=0
cc_233 N_VPWR_c_283_n N_Y_c_353_n 0.0255551f $X=2.545 $Y=2.455 $X2=0 $Y2=0
cc_234 N_VPWR_c_278_n N_Y_c_353_n 0.0120466f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_235 N_VPWR_M1014_s N_Y_c_365_n 0.0191728f $X=2.035 $Y=1.84 $X2=0 $Y2=0
cc_236 N_VPWR_c_283_n N_Y_c_365_n 0.0444218f $X=2.545 $Y=2.455 $X2=0 $Y2=0
cc_237 N_VPWR_c_283_n N_Y_c_354_n 0.0255551f $X=2.545 $Y=2.455 $X2=0 $Y2=0
cc_238 N_VPWR_c_284_n N_Y_c_354_n 0.0266809f $X=3.495 $Y=2.41 $X2=0 $Y2=0
cc_239 N_VPWR_c_287_n N_Y_c_354_n 0.014552f $X=3.33 $Y=3.33 $X2=0 $Y2=0
cc_240 N_VPWR_c_278_n N_Y_c_354_n 0.0119791f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_241 N_VPWR_M1005_s N_Y_c_375_n 0.00659271f $X=3.295 $Y=1.84 $X2=0 $Y2=0
cc_242 N_VPWR_c_284_n N_Y_c_375_n 0.0240821f $X=3.495 $Y=2.41 $X2=0 $Y2=0
cc_243 N_VPWR_c_284_n N_Y_c_355_n 0.0249406f $X=3.495 $Y=2.41 $X2=0 $Y2=0
cc_244 N_VPWR_c_286_n N_Y_c_355_n 0.0255379f $X=4.46 $Y=2.41 $X2=0 $Y2=0
cc_245 N_VPWR_c_290_n N_Y_c_355_n 0.0125859f $X=4.295 $Y=3.33 $X2=0 $Y2=0
cc_246 N_VPWR_c_278_n N_Y_c_355_n 0.0103846f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_247 N_VPWR_M1008_s N_Y_c_388_n 0.00406699f $X=4.305 $Y=1.84 $X2=0 $Y2=0
cc_248 N_VPWR_c_286_n N_Y_c_388_n 0.00744128f $X=4.46 $Y=2.41 $X2=0 $Y2=0
cc_249 N_VPWR_M1008_s Y 0.00210164f $X=4.305 $Y=1.84 $X2=0 $Y2=0
cc_250 N_VPWR_M1008_s Y 0.00341998f $X=4.305 $Y=1.84 $X2=0 $Y2=0
cc_251 N_VPWR_c_286_n Y 0.016108f $X=4.46 $Y=2.41 $X2=0 $Y2=0
cc_252 N_Y_c_350_n N_A_304_74#_c_514_n 0.00165751f $X=4.175 $Y=1.095 $X2=0 $Y2=0
cc_253 N_Y_c_349_n N_A_515_74#_M1015_s 0.00248296f $X=4.445 $Y=1.095 $X2=0 $Y2=0
cc_254 N_Y_c_350_n N_A_515_74#_c_547_n 0.00578498f $X=4.175 $Y=1.095 $X2=0 $Y2=0
cc_255 N_Y_M1010_d N_A_515_74#_c_548_n 0.00221305f $X=3.87 $Y=0.37 $X2=0 $Y2=0
cc_256 N_Y_c_386_n N_A_515_74#_c_548_n 0.0126288f $X=4.01 $Y=0.81 $X2=0 $Y2=0
cc_257 N_Y_c_349_n N_A_515_74#_c_548_n 0.00352022f $X=4.445 $Y=1.095 $X2=0 $Y2=0
cc_258 N_Y_c_349_n N_A_515_74#_c_549_n 0.0262099f $X=4.445 $Y=1.095 $X2=0 $Y2=0
cc_259 N_A_27_74#_c_437_n N_VGND_M1001_s 0.00277613f $X=1.145 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_260 N_A_27_74#_c_436_n N_VGND_c_473_n 0.0191765f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_261 N_A_27_74#_c_437_n N_VGND_c_473_n 0.0211325f $X=1.145 $Y=1.095 $X2=0
+ $Y2=0
cc_262 N_A_27_74#_c_440_n N_VGND_c_473_n 0.0103602f $X=1.315 $Y=0.34 $X2=0 $Y2=0
cc_263 N_A_27_74#_c_436_n N_VGND_c_474_n 0.0145639f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_264 N_A_27_74#_c_439_n N_VGND_c_475_n 0.0662638f $X=1.995 $Y=0.34 $X2=0 $Y2=0
cc_265 N_A_27_74#_c_440_n N_VGND_c_475_n 0.0121867f $X=1.315 $Y=0.34 $X2=0 $Y2=0
cc_266 N_A_27_74#_c_436_n N_VGND_c_476_n 0.0119984f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_267 N_A_27_74#_c_439_n N_VGND_c_476_n 0.0369729f $X=1.995 $Y=0.34 $X2=0 $Y2=0
cc_268 N_A_27_74#_c_440_n N_VGND_c_476_n 0.00660921f $X=1.315 $Y=0.34 $X2=0
+ $Y2=0
cc_269 N_A_27_74#_c_439_n N_A_304_74#_M1007_d 0.00176461f $X=1.995 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_270 N_A_27_74#_c_439_n N_A_304_74#_c_516_n 0.0158692f $X=1.995 $Y=0.34 $X2=0
+ $Y2=0
cc_271 N_A_27_74#_M1013_s N_A_304_74#_c_514_n 0.0024352f $X=1.95 $Y=0.37 $X2=0
+ $Y2=0
cc_272 N_A_27_74#_c_439_n N_A_304_74#_c_514_n 0.00304353f $X=1.995 $Y=0.34 $X2=0
+ $Y2=0
cc_273 N_A_27_74#_c_441_n N_A_304_74#_c_514_n 0.0258546f $X=2.16 $Y=0.595 $X2=0
+ $Y2=0
cc_274 N_A_27_74#_c_437_n N_A_304_74#_c_515_n 0.00997012f $X=1.145 $Y=1.095
+ $X2=0 $Y2=0
cc_275 N_A_27_74#_c_441_n N_A_515_74#_c_544_n 0.0274168f $X=2.16 $Y=0.595 $X2=0
+ $Y2=0
cc_276 N_A_27_74#_c_439_n N_A_515_74#_c_546_n 0.0128666f $X=1.995 $Y=0.34 $X2=0
+ $Y2=0
cc_277 N_VGND_c_475_n N_A_515_74#_c_545_n 0.0422287f $X=4.56 $Y=0 $X2=0 $Y2=0
cc_278 N_VGND_c_476_n N_A_515_74#_c_545_n 0.0238173f $X=4.56 $Y=0 $X2=0 $Y2=0
cc_279 N_VGND_c_475_n N_A_515_74#_c_546_n 0.0184296f $X=4.56 $Y=0 $X2=0 $Y2=0
cc_280 N_VGND_c_476_n N_A_515_74#_c_546_n 0.0100689f $X=4.56 $Y=0 $X2=0 $Y2=0
cc_281 N_VGND_c_475_n N_A_515_74#_c_548_n 0.0656196f $X=4.56 $Y=0 $X2=0 $Y2=0
cc_282 N_VGND_c_476_n N_A_515_74#_c_548_n 0.036597f $X=4.56 $Y=0 $X2=0 $Y2=0
cc_283 N_VGND_c_475_n N_A_515_74#_c_550_n 0.0136205f $X=4.56 $Y=0 $X2=0 $Y2=0
cc_284 N_VGND_c_476_n N_A_515_74#_c_550_n 0.00738676f $X=4.56 $Y=0 $X2=0 $Y2=0
cc_285 N_A_304_74#_c_514_n N_A_515_74#_M1004_d 0.0024352f $X=2.985 $Y=1.095
+ $X2=-0.19 $Y2=-0.245
cc_286 N_A_304_74#_c_514_n N_A_515_74#_c_544_n 0.0200155f $X=2.985 $Y=1.095
+ $X2=0 $Y2=0
cc_287 N_A_304_74#_M1004_s N_A_515_74#_c_545_n 0.00197509f $X=3.01 $Y=0.37 $X2=0
+ $Y2=0
cc_288 N_A_304_74#_c_514_n N_A_515_74#_c_545_n 0.00304353f $X=2.985 $Y=1.095
+ $X2=0 $Y2=0
cc_289 N_A_304_74#_c_529_n N_A_515_74#_c_545_n 0.0125343f $X=3.15 $Y=0.81 $X2=0
+ $Y2=0
cc_290 N_A_304_74#_c_514_n N_A_515_74#_c_547_n 0.00578498f $X=2.985 $Y=1.095
+ $X2=0 $Y2=0
