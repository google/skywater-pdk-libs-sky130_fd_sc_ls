* File: sky130_fd_sc_ls__einvp_8.pex.spice
* Created: Fri Aug 28 13:24:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__EINVP_8%A 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22 24
+ 25 27 28 30 31 33 34 36 37 39 40 42 43 45 46 48 49 50 51 52 53 89 91
c157 91 0 5.65346e-20 $X=3.65 $Y=1.492
c158 46 0 1.9142e-19 $X=3.925 $Y=1.22
c159 43 0 1.88567e-19 $X=3.65 $Y=1.765
c160 40 0 8.60601e-20 $X=3.425 $Y=1.22
c161 28 0 8.60601e-20 $X=2.425 $Y=1.22
c162 16 0 8.60869e-20 $X=1.425 $Y=1.22
r163 90 91 26.9107 $w=4.03e-07 $l=2.25e-07 $layer=POLY_cond $X=3.425 $Y=1.492
+ $X2=3.65 $Y2=1.492
r164 88 90 15.5484 $w=4.03e-07 $l=1.3e-07 $layer=POLY_cond $X=3.295 $Y=1.492
+ $X2=3.425 $Y2=1.492
r165 88 89 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.295
+ $Y=1.385 $X2=3.295 $Y2=1.385
r166 86 88 11.3623 $w=4.03e-07 $l=9.5e-08 $layer=POLY_cond $X=3.2 $Y=1.492
+ $X2=3.295 $Y2=1.492
r167 85 86 32.8908 $w=4.03e-07 $l=2.75e-07 $layer=POLY_cond $X=2.925 $Y=1.492
+ $X2=3.2 $Y2=1.492
r168 84 85 20.9305 $w=4.03e-07 $l=1.75e-07 $layer=POLY_cond $X=2.75 $Y=1.492
+ $X2=2.925 $Y2=1.492
r169 82 84 16.1464 $w=4.03e-07 $l=1.35e-07 $layer=POLY_cond $X=2.615 $Y=1.492
+ $X2=2.75 $Y2=1.492
r170 82 83 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.615
+ $Y=1.385 $X2=2.615 $Y2=1.385
r171 80 82 22.7246 $w=4.03e-07 $l=1.9e-07 $layer=POLY_cond $X=2.425 $Y=1.492
+ $X2=2.615 $Y2=1.492
r172 79 80 14.9504 $w=4.03e-07 $l=1.25e-07 $layer=POLY_cond $X=2.3 $Y=1.492
+ $X2=2.425 $Y2=1.492
r173 78 83 10.59 $w=3.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.275 $Y=1.365
+ $X2=2.615 $Y2=1.365
r174 77 79 2.99007 $w=4.03e-07 $l=2.5e-08 $layer=POLY_cond $X=2.275 $Y=1.492
+ $X2=2.3 $Y2=1.492
r175 77 78 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.275
+ $Y=1.385 $X2=2.275 $Y2=1.385
r176 75 77 41.861 $w=4.03e-07 $l=3.5e-07 $layer=POLY_cond $X=1.925 $Y=1.492
+ $X2=2.275 $Y2=1.492
r177 74 75 8.97022 $w=4.03e-07 $l=7.5e-08 $layer=POLY_cond $X=1.85 $Y=1.492
+ $X2=1.925 $Y2=1.492
r178 72 74 30.4988 $w=4.03e-07 $l=2.55e-07 $layer=POLY_cond $X=1.595 $Y=1.492
+ $X2=1.85 $Y2=1.492
r179 72 73 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.595
+ $Y=1.385 $X2=1.595 $Y2=1.385
r180 70 72 20.3325 $w=4.03e-07 $l=1.7e-07 $layer=POLY_cond $X=1.425 $Y=1.492
+ $X2=1.595 $Y2=1.492
r181 69 70 2.99007 $w=4.03e-07 $l=2.5e-08 $layer=POLY_cond $X=1.4 $Y=1.492
+ $X2=1.425 $Y2=1.492
r182 68 73 10.59 $w=3.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.255 $Y=1.365
+ $X2=1.595 $Y2=1.365
r183 67 69 17.3424 $w=4.03e-07 $l=1.45e-07 $layer=POLY_cond $X=1.255 $Y=1.492
+ $X2=1.4 $Y2=1.492
r184 67 68 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.255
+ $Y=1.385 $X2=1.255 $Y2=1.385
r185 65 67 36.4789 $w=4.03e-07 $l=3.05e-07 $layer=POLY_cond $X=0.95 $Y=1.492
+ $X2=1.255 $Y2=1.492
r186 64 65 2.99007 $w=4.03e-07 $l=2.5e-08 $layer=POLY_cond $X=0.925 $Y=1.492
+ $X2=0.95 $Y2=1.492
r187 62 64 1.19603 $w=4.03e-07 $l=1e-08 $layer=POLY_cond $X=0.915 $Y=1.492
+ $X2=0.925 $Y2=1.492
r188 62 63 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.915
+ $Y=1.385 $X2=0.915 $Y2=1.385
r189 60 62 49.6352 $w=4.03e-07 $l=4.15e-07 $layer=POLY_cond $X=0.5 $Y=1.492
+ $X2=0.915 $Y2=1.492
r190 59 60 0.598015 $w=4.03e-07 $l=5e-09 $layer=POLY_cond $X=0.495 $Y=1.492
+ $X2=0.5 $Y2=1.492
r191 53 89 5.45074 $w=3.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.12 $Y=1.365
+ $X2=3.295 $Y2=1.365
r192 52 53 14.9506 $w=3.68e-07 $l=4.8e-07 $layer=LI1_cond $X=2.64 $Y=1.365
+ $X2=3.12 $Y2=1.365
r193 52 83 0.778678 $w=3.68e-07 $l=2.5e-08 $layer=LI1_cond $X=2.64 $Y=1.365
+ $X2=2.615 $Y2=1.365
r194 51 78 3.58192 $w=3.68e-07 $l=1.15e-07 $layer=LI1_cond $X=2.16 $Y=1.365
+ $X2=2.275 $Y2=1.365
r195 50 51 14.9506 $w=3.68e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=1.365
+ $X2=2.16 $Y2=1.365
r196 50 73 2.6475 $w=3.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.68 $Y=1.365
+ $X2=1.595 $Y2=1.365
r197 49 68 1.71309 $w=3.68e-07 $l=5.5e-08 $layer=LI1_cond $X=1.2 $Y=1.365
+ $X2=1.255 $Y2=1.365
r198 49 63 8.87693 $w=3.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.2 $Y=1.365
+ $X2=0.915 $Y2=1.365
r199 46 91 32.8908 $w=4.03e-07 $l=3.87847e-07 $layer=POLY_cond $X=3.925 $Y=1.22
+ $X2=3.65 $Y2=1.492
r200 46 48 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.925 $Y=1.22
+ $X2=3.925 $Y2=0.74
r201 43 91 26.0447 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=3.65 $Y=1.765
+ $X2=3.65 $Y2=1.492
r202 43 45 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.65 $Y=1.765
+ $X2=3.65 $Y2=2.4
r203 40 90 26.0447 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=3.425 $Y=1.22
+ $X2=3.425 $Y2=1.492
r204 40 42 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.425 $Y=1.22
+ $X2=3.425 $Y2=0.74
r205 37 86 26.0447 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=3.2 $Y=1.765
+ $X2=3.2 $Y2=1.492
r206 37 39 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.2 $Y=1.765
+ $X2=3.2 $Y2=2.4
r207 34 85 26.0447 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=2.925 $Y=1.22
+ $X2=2.925 $Y2=1.492
r208 34 36 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.925 $Y=1.22
+ $X2=2.925 $Y2=0.74
r209 31 84 26.0447 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=2.75 $Y=1.765
+ $X2=2.75 $Y2=1.492
r210 31 33 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.75 $Y=1.765
+ $X2=2.75 $Y2=2.4
r211 28 80 26.0447 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=2.425 $Y=1.22
+ $X2=2.425 $Y2=1.492
r212 28 30 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.425 $Y=1.22
+ $X2=2.425 $Y2=0.74
r213 25 79 26.0447 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=2.3 $Y=1.765
+ $X2=2.3 $Y2=1.492
r214 25 27 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.3 $Y=1.765
+ $X2=2.3 $Y2=2.4
r215 22 75 26.0447 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=1.925 $Y=1.22
+ $X2=1.925 $Y2=1.492
r216 22 24 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.925 $Y=1.22
+ $X2=1.925 $Y2=0.74
r217 19 74 26.0447 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=1.85 $Y=1.765
+ $X2=1.85 $Y2=1.492
r218 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.85 $Y=1.765
+ $X2=1.85 $Y2=2.4
r219 16 70 26.0447 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=1.425 $Y=1.22
+ $X2=1.425 $Y2=1.492
r220 16 18 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.425 $Y=1.22
+ $X2=1.425 $Y2=0.74
r221 13 69 26.0447 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=1.4 $Y=1.765
+ $X2=1.4 $Y2=1.492
r222 13 15 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.4 $Y=1.765
+ $X2=1.4 $Y2=2.4
r223 10 65 26.0447 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=0.95 $Y=1.765
+ $X2=0.95 $Y2=1.492
r224 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.95 $Y=1.765
+ $X2=0.95 $Y2=2.4
r225 7 64 26.0447 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=0.925 $Y=1.22
+ $X2=0.925 $Y2=1.492
r226 7 9 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.925 $Y=1.22
+ $X2=0.925 $Y2=0.74
r227 4 60 26.0447 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=0.5 $Y=1.765
+ $X2=0.5 $Y2=1.492
r228 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.5 $Y=1.765 $X2=0.5
+ $Y2=2.4
r229 1 59 26.0447 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=0.495 $Y=1.22
+ $X2=0.495 $Y2=1.492
r230 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.495 $Y=1.22
+ $X2=0.495 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__EINVP_8%A_802_323# 1 2 7 9 10 11 12 14 15 17 19 20
+ 22 24 25 27 29 30 32 34 35 37 39 40 42 44 45 47 48 49 50 51 52 53 56 59 63 68
c180 56 0 3.05834e-20 $X=8.14 $Y=1.615
r181 68 70 17.9954 $w=4.48e-07 $l=4.95e-07 $layer=LI1_cond $X=8.28 $Y=0.515
+ $X2=8.28 $Y2=1.01
r182 63 66 0.249659 $w=7.33e-07 $l=1.5e-08 $layer=LI1_cond $X=8.17 $Y=2.8
+ $X2=8.17 $Y2=2.815
r183 63 64 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.94
+ $Y=2.8 $X2=7.94 $Y2=2.8
r184 61 63 13.5648 $w=7.33e-07 $l=8.15e-07 $layer=LI1_cond $X=8.17 $Y=1.985
+ $X2=8.17 $Y2=2.8
r185 59 64 178.359 $w=3.3e-07 $l=1.02e-06 $layer=POLY_cond $X=7.94 $Y=1.78
+ $X2=7.94 $Y2=2.8
r186 58 61 3.41201 $w=7.33e-07 $l=2.05e-07 $layer=LI1_cond $X=8.17 $Y=1.78
+ $X2=8.17 $Y2=1.985
r187 58 59 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.94
+ $Y=1.78 $X2=7.94 $Y2=1.78
r188 56 58 11.2359 $w=7.33e-07 $l=1.79374e-07 $layer=LI1_cond $X=8.14 $Y=1.615
+ $X2=8.17 $Y2=1.78
r189 56 70 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=8.14 $Y=1.615
+ $X2=8.14 $Y2=1.01
r190 54 59 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=7.94 $Y=1.765
+ $X2=7.94 $Y2=1.78
r191 46 53 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.325 $Y=1.69
+ $X2=7.25 $Y2=1.69
r192 45 54 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=7.775 $Y=1.69
+ $X2=7.94 $Y2=1.765
r193 45 46 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=7.775 $Y=1.69
+ $X2=7.325 $Y2=1.69
r194 42 53 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.25 $Y=1.765
+ $X2=7.25 $Y2=1.69
r195 42 44 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.25 $Y=1.765
+ $X2=7.25 $Y2=2.4
r196 41 52 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.875 $Y=1.69
+ $X2=6.8 $Y2=1.69
r197 40 53 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.175 $Y=1.69
+ $X2=7.25 $Y2=1.69
r198 40 41 153.83 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=7.175 $Y=1.69
+ $X2=6.875 $Y2=1.69
r199 37 52 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.8 $Y=1.765
+ $X2=6.8 $Y2=1.69
r200 37 39 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.8 $Y=1.765
+ $X2=6.8 $Y2=2.4
r201 36 51 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.425 $Y=1.69
+ $X2=6.35 $Y2=1.69
r202 35 52 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.725 $Y=1.69
+ $X2=6.8 $Y2=1.69
r203 35 36 153.83 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=6.725 $Y=1.69
+ $X2=6.425 $Y2=1.69
r204 32 51 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.35 $Y=1.765
+ $X2=6.35 $Y2=1.69
r205 32 34 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.35 $Y=1.765
+ $X2=6.35 $Y2=2.4
r206 31 50 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.975 $Y=1.69
+ $X2=5.9 $Y2=1.69
r207 30 51 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.275 $Y=1.69
+ $X2=6.35 $Y2=1.69
r208 30 31 153.83 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=6.275 $Y=1.69
+ $X2=5.975 $Y2=1.69
r209 27 50 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.9 $Y=1.765
+ $X2=5.9 $Y2=1.69
r210 27 29 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.9 $Y=1.765
+ $X2=5.9 $Y2=2.4
r211 26 49 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.525 $Y=1.69
+ $X2=5.45 $Y2=1.69
r212 25 50 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.825 $Y=1.69
+ $X2=5.9 $Y2=1.69
r213 25 26 153.83 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=5.825 $Y=1.69
+ $X2=5.525 $Y2=1.69
r214 22 49 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.45 $Y=1.765
+ $X2=5.45 $Y2=1.69
r215 22 24 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.45 $Y=1.765
+ $X2=5.45 $Y2=2.4
r216 21 48 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.075 $Y=1.69 $X2=5
+ $Y2=1.69
r217 20 49 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.375 $Y=1.69
+ $X2=5.45 $Y2=1.69
r218 20 21 153.83 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=5.375 $Y=1.69
+ $X2=5.075 $Y2=1.69
r219 17 48 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5 $Y=1.765 $X2=5
+ $Y2=1.69
r220 17 19 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5 $Y=1.765 $X2=5
+ $Y2=2.4
r221 16 47 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.625 $Y=1.69
+ $X2=4.55 $Y2=1.69
r222 15 48 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.925 $Y=1.69 $X2=5
+ $Y2=1.69
r223 15 16 153.83 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=4.925 $Y=1.69
+ $X2=4.625 $Y2=1.69
r224 12 47 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.55 $Y=1.765
+ $X2=4.55 $Y2=1.69
r225 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.55 $Y=1.765
+ $X2=4.55 $Y2=2.4
r226 10 47 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.475 $Y=1.69
+ $X2=4.55 $Y2=1.69
r227 10 11 153.83 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=4.475 $Y=1.69
+ $X2=4.175 $Y2=1.69
r228 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.1 $Y=1.765
+ $X2=4.175 $Y2=1.69
r229 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.1 $Y=1.765 $X2=4.1
+ $Y2=2.4
r230 2 66 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=8.265
+ $Y=1.84 $X2=8.4 $Y2=2.815
r231 2 61 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=8.265
+ $Y=1.84 $X2=8.4 $Y2=1.985
r232 1 68 91 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_NDIFF $count=2 $X=8.19
+ $Y=0.37 $X2=8.34 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__EINVP_8%TE 1 3 4 5 6 8 9 11 13 14 16 18 19 21 23 24
+ 26 28 29 31 33 34 36 38 39 41 43 44 46 47 48 49 50 51 52 53 54
c150 36 0 3.05834e-20 $X=7.505 $Y=1.22
c151 31 0 1.07496e-19 $X=7.005 $Y=1.22
c152 6 0 1.07496e-19 $X=4.855 $Y=1.22
c153 1 0 3.03515e-19 $X=4.355 $Y=1.22
r154 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.6
+ $Y=1.385 $X2=8.6 $Y2=1.385
r155 56 58 16.0667 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=8.6 $Y=1.295 $X2=8.6
+ $Y2=1.385
r156 54 59 10.9487 $w=3.12e-07 $l=2.8e-07 $layer=LI1_cond $X=8.88 $Y=1.365
+ $X2=8.6 $Y2=1.365
r157 44 58 77.2841 $w=2.7e-07 $l=3.92301e-07 $layer=POLY_cond $X=8.625 $Y=1.765
+ $X2=8.6 $Y2=1.385
r158 44 46 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.625 $Y=1.765
+ $X2=8.625 $Y2=2.4
r159 41 56 22.8359 $w=2.7e-07 $l=9.48683e-08 $layer=POLY_cond $X=8.555 $Y=1.22
+ $X2=8.6 $Y2=1.295
r160 41 43 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=8.555 $Y=1.22
+ $X2=8.555 $Y2=0.74
r161 40 53 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.58 $Y=1.295
+ $X2=7.505 $Y2=1.295
r162 39 56 16.5046 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.435 $Y=1.295
+ $X2=8.6 $Y2=1.295
r163 39 40 438.415 $w=1.5e-07 $l=8.55e-07 $layer=POLY_cond $X=8.435 $Y=1.295
+ $X2=7.58 $Y2=1.295
r164 36 53 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.505 $Y=1.22
+ $X2=7.505 $Y2=1.295
r165 36 38 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=7.505 $Y=1.22
+ $X2=7.505 $Y2=0.74
r166 35 52 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.08 $Y=1.295
+ $X2=7.005 $Y2=1.295
r167 34 53 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.43 $Y=1.295
+ $X2=7.505 $Y2=1.295
r168 34 35 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=7.43 $Y=1.295
+ $X2=7.08 $Y2=1.295
r169 31 52 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.005 $Y=1.22
+ $X2=7.005 $Y2=1.295
r170 31 33 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=7.005 $Y=1.22
+ $X2=7.005 $Y2=0.74
r171 30 51 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.65 $Y=1.295
+ $X2=6.575 $Y2=1.295
r172 29 52 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.93 $Y=1.295
+ $X2=7.005 $Y2=1.295
r173 29 30 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=6.93 $Y=1.295
+ $X2=6.65 $Y2=1.295
r174 26 51 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.575 $Y=1.22
+ $X2=6.575 $Y2=1.295
r175 26 28 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=6.575 $Y=1.22
+ $X2=6.575 $Y2=0.74
r176 25 50 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.22 $Y=1.295
+ $X2=6.145 $Y2=1.295
r177 24 51 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.5 $Y=1.295
+ $X2=6.575 $Y2=1.295
r178 24 25 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=6.5 $Y=1.295
+ $X2=6.22 $Y2=1.295
r179 21 50 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.145 $Y=1.22
+ $X2=6.145 $Y2=1.295
r180 21 23 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=6.145 $Y=1.22
+ $X2=6.145 $Y2=0.74
r181 20 49 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.79 $Y=1.295
+ $X2=5.715 $Y2=1.295
r182 19 50 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.07 $Y=1.295
+ $X2=6.145 $Y2=1.295
r183 19 20 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=6.07 $Y=1.295
+ $X2=5.79 $Y2=1.295
r184 16 49 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.715 $Y=1.22
+ $X2=5.715 $Y2=1.295
r185 16 18 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.715 $Y=1.22
+ $X2=5.715 $Y2=0.74
r186 15 48 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.36 $Y=1.295
+ $X2=5.285 $Y2=1.295
r187 14 49 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.64 $Y=1.295
+ $X2=5.715 $Y2=1.295
r188 14 15 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=5.64 $Y=1.295
+ $X2=5.36 $Y2=1.295
r189 11 48 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.285 $Y=1.22
+ $X2=5.285 $Y2=1.295
r190 11 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.285 $Y=1.22
+ $X2=5.285 $Y2=0.74
r191 10 47 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.93 $Y=1.295
+ $X2=4.855 $Y2=1.295
r192 9 48 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.21 $Y=1.295
+ $X2=5.285 $Y2=1.295
r193 9 10 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=5.21 $Y=1.295
+ $X2=4.93 $Y2=1.295
r194 6 47 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.855 $Y=1.22
+ $X2=4.855 $Y2=1.295
r195 6 8 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.855 $Y=1.22
+ $X2=4.855 $Y2=0.74
r196 4 47 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.78 $Y=1.295
+ $X2=4.855 $Y2=1.295
r197 4 5 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=4.78 $Y=1.295
+ $X2=4.43 $Y2=1.295
r198 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.355 $Y=1.22
+ $X2=4.43 $Y2=1.295
r199 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.355 $Y=1.22
+ $X2=4.355 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__EINVP_8%A_27_368# 1 2 3 4 5 6 7 8 9 30 34 35 38 40
+ 44 46 50 52 54 55 56 61 64 66 67 70 74 78 82 86 90 91 92 95 96 97
r163 86 88 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=7.435 $Y=1.985
+ $X2=7.435 $Y2=2.815
r164 84 86 12.2159 $w=2.48e-07 $l=2.65e-07 $layer=LI1_cond $X=7.435 $Y=1.72
+ $X2=7.435 $Y2=1.985
r165 83 97 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.66 $Y=1.635
+ $X2=6.535 $Y2=1.635
r166 82 84 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=7.31 $Y=1.635
+ $X2=7.435 $Y2=1.72
r167 82 83 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=7.31 $Y=1.635
+ $X2=6.66 $Y2=1.635
r168 78 80 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=6.535 $Y=1.985
+ $X2=6.535 $Y2=2.815
r169 76 97 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.535 $Y=1.72
+ $X2=6.535 $Y2=1.635
r170 76 78 12.2159 $w=2.48e-07 $l=2.65e-07 $layer=LI1_cond $X=6.535 $Y=1.72
+ $X2=6.535 $Y2=1.985
r171 75 96 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.76 $Y=1.635
+ $X2=5.635 $Y2=1.635
r172 74 97 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.41 $Y=1.635
+ $X2=6.535 $Y2=1.635
r173 74 75 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=6.41 $Y=1.635
+ $X2=5.76 $Y2=1.635
r174 70 72 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=5.635 $Y=1.985
+ $X2=5.635 $Y2=2.815
r175 68 96 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.635 $Y=1.72
+ $X2=5.635 $Y2=1.635
r176 68 70 12.2159 $w=2.48e-07 $l=2.65e-07 $layer=LI1_cond $X=5.635 $Y=1.72
+ $X2=5.635 $Y2=1.985
r177 66 96 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.51 $Y=1.635
+ $X2=5.635 $Y2=1.635
r178 66 67 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=5.51 $Y=1.635
+ $X2=4.94 $Y2=1.635
r179 62 95 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.815 $Y=2.23
+ $X2=4.815 $Y2=2.145
r180 62 64 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=4.815 $Y=2.23
+ $X2=4.815 $Y2=2.4
r181 59 95 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.815 $Y=2.06
+ $X2=4.815 $Y2=2.145
r182 59 61 3.45733 $w=2.48e-07 $l=7.5e-08 $layer=LI1_cond $X=4.815 $Y=2.06
+ $X2=4.815 $Y2=1.985
r183 58 67 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.815 $Y=1.72
+ $X2=4.94 $Y2=1.635
r184 58 61 12.2159 $w=2.48e-07 $l=2.65e-07 $layer=LI1_cond $X=4.815 $Y=1.72
+ $X2=4.815 $Y2=1.985
r185 57 94 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.96 $Y=2.145
+ $X2=3.875 $Y2=2.145
r186 56 95 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.69 $Y=2.145
+ $X2=4.815 $Y2=2.145
r187 56 57 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=4.69 $Y=2.145
+ $X2=3.96 $Y2=2.145
r188 54 94 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.875 $Y=2.23
+ $X2=3.875 $Y2=2.145
r189 54 55 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=3.875 $Y=2.23
+ $X2=3.875 $Y2=2.905
r190 53 92 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=3.075 $Y=2.99
+ $X2=2.975 $Y2=2.99
r191 52 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.79 $Y=2.99
+ $X2=3.875 $Y2=2.905
r192 52 53 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=3.79 $Y=2.99
+ $X2=3.075 $Y2=2.99
r193 48 92 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=2.975 $Y=2.905
+ $X2=2.975 $Y2=2.99
r194 48 50 37.7091 $w=1.98e-07 $l=6.8e-07 $layer=LI1_cond $X=2.975 $Y=2.905
+ $X2=2.975 $Y2=2.225
r195 47 91 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=2.19 $Y=2.99
+ $X2=2.08 $Y2=2.99
r196 46 92 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=2.875 $Y=2.99
+ $X2=2.975 $Y2=2.99
r197 46 47 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=2.875 $Y=2.99
+ $X2=2.19 $Y2=2.99
r198 42 91 0.432806 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=2.08 $Y=2.905
+ $X2=2.08 $Y2=2.99
r199 42 44 35.621 $w=2.18e-07 $l=6.8e-07 $layer=LI1_cond $X=2.08 $Y=2.905
+ $X2=2.08 $Y2=2.225
r200 41 90 6.01921 $w=1.7e-07 $l=1.03e-07 $layer=LI1_cond $X=1.275 $Y=2.99
+ $X2=1.172 $Y2=2.99
r201 40 91 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=1.97 $Y=2.99
+ $X2=2.08 $Y2=2.99
r202 40 41 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=1.97 $Y=2.99
+ $X2=1.275 $Y2=2.99
r203 36 90 0.677923 $w=2.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.172 $Y=2.905
+ $X2=1.172 $Y2=2.99
r204 36 38 36.7894 $w=2.03e-07 $l=6.8e-07 $layer=LI1_cond $X=1.172 $Y=2.905
+ $X2=1.172 $Y2=2.225
r205 34 90 6.01921 $w=1.7e-07 $l=1.02e-07 $layer=LI1_cond $X=1.07 $Y=2.99
+ $X2=1.172 $Y2=2.99
r206 34 35 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=1.07 $Y=2.99
+ $X2=0.375 $Y2=2.99
r207 30 33 36.0954 $w=2.63e-07 $l=8.3e-07 $layer=LI1_cond $X=0.242 $Y=1.985
+ $X2=0.242 $Y2=2.815
r208 28 35 7.24806 $w=1.7e-07 $l=1.70276e-07 $layer=LI1_cond $X=0.242 $Y=2.905
+ $X2=0.375 $Y2=2.99
r209 28 33 3.91396 $w=2.63e-07 $l=9e-08 $layer=LI1_cond $X=0.242 $Y=2.905
+ $X2=0.242 $Y2=2.815
r210 9 88 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=7.325
+ $Y=1.84 $X2=7.475 $Y2=2.815
r211 9 86 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=7.325
+ $Y=1.84 $X2=7.475 $Y2=1.985
r212 8 80 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=6.425
+ $Y=1.84 $X2=6.575 $Y2=2.815
r213 8 78 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=6.425
+ $Y=1.84 $X2=6.575 $Y2=1.985
r214 7 72 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=5.525
+ $Y=1.84 $X2=5.675 $Y2=2.815
r215 7 70 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=5.525
+ $Y=1.84 $X2=5.675 $Y2=1.985
r216 6 64 300 $w=1.7e-07 $l=6.30555e-07 $layer=licon1_PDIFF $count=2 $X=4.625
+ $Y=1.84 $X2=4.775 $Y2=2.4
r217 6 61 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=4.625
+ $Y=1.84 $X2=4.775 $Y2=1.985
r218 5 94 300 $w=1.7e-07 $l=4.53845e-07 $layer=licon1_PDIFF $count=2 $X=3.725
+ $Y=1.84 $X2=3.875 $Y2=2.225
r219 4 50 300 $w=1.7e-07 $l=4.53845e-07 $layer=licon1_PDIFF $count=2 $X=2.825
+ $Y=1.84 $X2=2.975 $Y2=2.225
r220 3 44 300 $w=1.7e-07 $l=4.53845e-07 $layer=licon1_PDIFF $count=2 $X=1.925
+ $Y=1.84 $X2=2.075 $Y2=2.225
r221 2 38 300 $w=1.7e-07 $l=4.53845e-07 $layer=licon1_PDIFF $count=2 $X=1.025
+ $Y=1.84 $X2=1.175 $Y2=2.225
r222 1 33 400 $w=1.7e-07 $l=1.04265e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.275 $Y2=2.815
r223 1 30 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.275 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_LS__EINVP_8%Z 1 2 3 4 5 6 7 8 27 33 34 37 41 47 51 53 57
+ 62 64 68 71 72 73 76 77 79 83
c130 79 0 1.86694e-19 $X=3.71 $Y=0.76
c131 62 0 1.16821e-19 $X=3.79 $Y=1.55
r132 83 86 13.6602 $w=2.59e-07 $l=2.9e-07 $layer=LI1_cond $X=4.08 $Y=1.72
+ $X2=3.79 $Y2=1.72
r133 81 82 5.66838 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=3.71 $Y=0.925
+ $X2=3.71 $Y2=1.01
r134 79 81 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.71 $Y=0.76
+ $X2=3.71 $Y2=0.925
r135 75 77 8.6272 $w=3.93e-07 $l=1.65e-07 $layer=LI1_cond $X=2.71 $Y=0.812
+ $X2=2.875 $Y2=0.812
r136 75 76 8.6272 $w=3.93e-07 $l=1.65e-07 $layer=LI1_cond $X=2.71 $Y=0.812
+ $X2=2.545 $Y2=0.812
r137 72 76 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.875 $Y=0.925
+ $X2=2.545 $Y2=0.925
r138 70 72 8.6272 $w=3.93e-07 $l=1.65e-07 $layer=LI1_cond $X=1.71 $Y=0.812
+ $X2=1.875 $Y2=0.812
r139 70 71 8.6272 $w=3.93e-07 $l=1.65e-07 $layer=LI1_cond $X=1.71 $Y=0.812
+ $X2=1.545 $Y2=0.812
r140 64 66 6.68417 $w=2.48e-07 $l=1.45e-07 $layer=LI1_cond $X=0.75 $Y=0.78
+ $X2=0.75 $Y2=0.925
r141 62 86 3.20129 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=3.79 $Y=1.55
+ $X2=3.79 $Y2=1.72
r142 62 82 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=3.79 $Y=1.55
+ $X2=3.79 $Y2=1.01
r143 57 59 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=3.425 $Y=1.97
+ $X2=3.425 $Y2=2.65
r144 55 86 17.1931 $w=2.59e-07 $l=3.65e-07 $layer=LI1_cond $X=3.425 $Y=1.72
+ $X2=3.79 $Y2=1.72
r145 55 57 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=3.425 $Y=1.89
+ $X2=3.425 $Y2=1.97
r146 53 81 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.545 $Y=0.925
+ $X2=3.71 $Y2=0.925
r147 53 77 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.545 $Y=0.925
+ $X2=2.875 $Y2=0.925
r148 52 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.69 $Y=1.805
+ $X2=2.525 $Y2=1.805
r149 51 55 9.21269 $w=2.59e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.26 $Y=1.805
+ $X2=3.425 $Y2=1.72
r150 51 52 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=3.26 $Y=1.805
+ $X2=2.69 $Y2=1.805
r151 47 49 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=2.525 $Y=1.97
+ $X2=2.525 $Y2=2.65
r152 45 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.525 $Y=1.89
+ $X2=2.525 $Y2=1.805
r153 45 47 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=2.525 $Y=1.89
+ $X2=2.525 $Y2=1.97
r154 42 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.79 $Y=1.805
+ $X2=1.625 $Y2=1.805
r155 41 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.36 $Y=1.805
+ $X2=2.525 $Y2=1.805
r156 41 42 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=2.36 $Y=1.805
+ $X2=1.79 $Y2=1.805
r157 37 39 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.625 $Y=1.97
+ $X2=1.625 $Y2=2.65
r158 35 68 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.625 $Y=1.89
+ $X2=1.625 $Y2=1.805
r159 35 37 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=1.625 $Y=1.89
+ $X2=1.625 $Y2=1.97
r160 33 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.46 $Y=1.805
+ $X2=1.625 $Y2=1.805
r161 33 34 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.46 $Y=1.805
+ $X2=0.89 $Y2=1.805
r162 32 66 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.875 $Y=0.925
+ $X2=0.75 $Y2=0.925
r163 32 71 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.875 $Y=0.925
+ $X2=1.545 $Y2=0.925
r164 27 29 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.725 $Y=1.97
+ $X2=0.725 $Y2=2.65
r165 25 34 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.725 $Y=1.89
+ $X2=0.89 $Y2=1.805
r166 25 27 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=0.725 $Y=1.89
+ $X2=0.725 $Y2=1.97
r167 8 59 400 $w=1.7e-07 $l=8.81816e-07 $layer=licon1_PDIFF $count=1 $X=3.275
+ $Y=1.84 $X2=3.425 $Y2=2.65
r168 8 57 400 $w=1.7e-07 $l=2.04939e-07 $layer=licon1_PDIFF $count=1 $X=3.275
+ $Y=1.84 $X2=3.425 $Y2=1.97
r169 7 49 400 $w=1.7e-07 $l=8.81816e-07 $layer=licon1_PDIFF $count=1 $X=2.375
+ $Y=1.84 $X2=2.525 $Y2=2.65
r170 7 47 400 $w=1.7e-07 $l=2.04939e-07 $layer=licon1_PDIFF $count=1 $X=2.375
+ $Y=1.84 $X2=2.525 $Y2=1.97
r171 6 39 400 $w=1.7e-07 $l=8.81816e-07 $layer=licon1_PDIFF $count=1 $X=1.475
+ $Y=1.84 $X2=1.625 $Y2=2.65
r172 6 37 400 $w=1.7e-07 $l=2.04939e-07 $layer=licon1_PDIFF $count=1 $X=1.475
+ $Y=1.84 $X2=1.625 $Y2=1.97
r173 5 29 400 $w=1.7e-07 $l=8.81816e-07 $layer=licon1_PDIFF $count=1 $X=0.575
+ $Y=1.84 $X2=0.725 $Y2=2.65
r174 5 27 400 $w=1.7e-07 $l=2.04939e-07 $layer=licon1_PDIFF $count=1 $X=0.575
+ $Y=1.84 $X2=0.725 $Y2=1.97
r175 4 79 182 $w=1.7e-07 $l=4.83735e-07 $layer=licon1_NDIFF $count=1 $X=3.5
+ $Y=0.37 $X2=3.71 $Y2=0.76
r176 3 75 182 $w=1.7e-07 $l=5.04182e-07 $layer=licon1_NDIFF $count=1 $X=2.5
+ $Y=0.37 $X2=2.71 $Y2=0.78
r177 2 70 182 $w=1.7e-07 $l=5.04182e-07 $layer=licon1_NDIFF $count=1 $X=1.5
+ $Y=0.37 $X2=1.71 $Y2=0.78
r178 1 64 182 $w=1.7e-07 $l=4.74868e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.78
.ends

.subckt PM_SKY130_FD_SC_LS__EINVP_8%VPWR 1 2 3 4 5 18 22 26 30 36 40 42 47 48 49
+ 50 51 63 68 77 80 84
c111 18 0 1.88567e-19 $X=4.325 $Y=2.485
r112 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r113 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r114 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r115 75 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=8.88 $Y2=3.33
r116 74 75 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r117 72 75 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=8.4 $Y2=3.33
r118 72 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6.96 $Y2=3.33
r119 71 74 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=7.44 $Y=3.33 $X2=8.4
+ $Y2=3.33
r120 71 72 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r121 69 80 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.11 $Y=3.33
+ $X2=6.985 $Y2=3.33
r122 69 71 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=7.11 $Y=3.33
+ $X2=7.44 $Y2=3.33
r123 68 83 4.02656 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=8.765 $Y=3.33
+ $X2=8.942 $Y2=3.33
r124 68 74 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=8.765 $Y=3.33
+ $X2=8.4 $Y2=3.33
r125 67 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6.96 $Y2=3.33
r126 67 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33 $X2=6
+ $Y2=3.33
r127 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r128 64 77 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.21 $Y=3.33
+ $X2=6.085 $Y2=3.33
r129 64 66 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=6.21 $Y=3.33
+ $X2=6.48 $Y2=3.33
r130 63 80 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.86 $Y=3.33
+ $X2=6.985 $Y2=3.33
r131 63 66 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=6.86 $Y=3.33
+ $X2=6.48 $Y2=3.33
r132 62 78 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33 $X2=6
+ $Y2=3.33
r133 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r134 58 59 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r135 55 59 1.07034 $w=4.9e-07 $l=3.84e-06 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=4.08 $Y2=3.33
r136 54 58 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=4.08 $Y2=3.33
r137 54 55 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r138 51 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r139 51 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r140 49 61 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=5.14 $Y=3.33 $X2=5.04
+ $Y2=3.33
r141 49 50 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.14 $Y=3.33
+ $X2=5.225 $Y2=3.33
r142 47 58 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=4.16 $Y=3.33 $X2=4.08
+ $Y2=3.33
r143 47 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.16 $Y=3.33
+ $X2=4.325 $Y2=3.33
r144 46 61 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=4.49 $Y=3.33
+ $X2=5.04 $Y2=3.33
r145 46 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.49 $Y=3.33
+ $X2=4.325 $Y2=3.33
r146 42 45 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=8.89 $Y=1.985
+ $X2=8.89 $Y2=2.815
r147 40 83 3.1166 $w=2.5e-07 $l=1.07912e-07 $layer=LI1_cond $X=8.89 $Y=3.245
+ $X2=8.942 $Y2=3.33
r148 40 45 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=8.89 $Y=3.245
+ $X2=8.89 $Y2=2.815
r149 36 39 35.0343 $w=2.48e-07 $l=7.6e-07 $layer=LI1_cond $X=6.985 $Y=2.055
+ $X2=6.985 $Y2=2.815
r150 34 80 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.985 $Y=3.245
+ $X2=6.985 $Y2=3.33
r151 34 39 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=6.985 $Y=3.245
+ $X2=6.985 $Y2=2.815
r152 30 33 35.0343 $w=2.48e-07 $l=7.6e-07 $layer=LI1_cond $X=6.085 $Y=2.055
+ $X2=6.085 $Y2=2.815
r153 28 77 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.085 $Y=3.245
+ $X2=6.085 $Y2=3.33
r154 28 33 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=6.085 $Y=3.245
+ $X2=6.085 $Y2=2.815
r155 27 50 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.31 $Y=3.33
+ $X2=5.225 $Y2=3.33
r156 26 77 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.96 $Y=3.33
+ $X2=6.085 $Y2=3.33
r157 26 27 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=5.96 $Y=3.33
+ $X2=5.31 $Y2=3.33
r158 22 25 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=5.225 $Y=2.055
+ $X2=5.225 $Y2=2.815
r159 20 50 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.225 $Y=3.245
+ $X2=5.225 $Y2=3.33
r160 20 25 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=5.225 $Y=3.245
+ $X2=5.225 $Y2=2.815
r161 16 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.325 $Y=3.245
+ $X2=4.325 $Y2=3.33
r162 16 18 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=4.325 $Y=3.245
+ $X2=4.325 $Y2=2.485
r163 5 45 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=8.7
+ $Y=1.84 $X2=8.85 $Y2=2.815
r164 5 42 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=8.7
+ $Y=1.84 $X2=8.85 $Y2=1.985
r165 4 39 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=6.875
+ $Y=1.84 $X2=7.025 $Y2=2.815
r166 4 36 400 $w=1.7e-07 $l=2.80134e-07 $layer=licon1_PDIFF $count=1 $X=6.875
+ $Y=1.84 $X2=7.025 $Y2=2.055
r167 3 33 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=5.975
+ $Y=1.84 $X2=6.125 $Y2=2.815
r168 3 30 400 $w=1.7e-07 $l=2.80134e-07 $layer=licon1_PDIFF $count=1 $X=5.975
+ $Y=1.84 $X2=6.125 $Y2=2.055
r169 2 25 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=5.075
+ $Y=1.84 $X2=5.225 $Y2=2.815
r170 2 22 400 $w=1.7e-07 $l=2.80134e-07 $layer=licon1_PDIFF $count=1 $X=5.075
+ $Y=1.84 $X2=5.225 $Y2=2.055
r171 1 18 300 $w=1.7e-07 $l=7.16083e-07 $layer=licon1_PDIFF $count=2 $X=4.175
+ $Y=1.84 $X2=4.325 $Y2=2.485
.ends

.subckt PM_SKY130_FD_SC_LS__EINVP_8%A_27_74# 1 2 3 4 5 6 7 8 9 30 32 33 34 36 38
+ 43 44 45 48 50 54 56 60 62 66 68 73 78 83 84 85
c172 85 0 1.07496e-19 $X=6.83 $Y=1.295
c173 83 0 1.07496e-19 $X=5.03 $Y=1.295
c174 45 0 5.65346e-20 $X=4.225 $Y=1.295
c175 36 0 8.60601e-20 $X=3.045 $Y=0.34
c176 34 0 8.60601e-20 $X=2.045 $Y=0.34
c177 32 0 8.60869e-20 $X=1.045 $Y=0.34
r178 78 81 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=3.21 $Y=0.34
+ $X2=3.21 $Y2=0.55
r179 73 76 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=2.21 $Y=0.34
+ $X2=2.21 $Y2=0.55
r180 68 71 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=1.21 $Y=0.34
+ $X2=1.21 $Y2=0.55
r181 64 66 32.0379 $w=2.48e-07 $l=6.95e-07 $layer=LI1_cond $X=7.76 $Y=1.21
+ $X2=7.76 $Y2=0.515
r182 63 85 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.955 $Y=1.295
+ $X2=6.83 $Y2=1.295
r183 62 64 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=7.635 $Y=1.295
+ $X2=7.76 $Y2=1.21
r184 62 63 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=7.635 $Y=1.295
+ $X2=6.955 $Y2=1.295
r185 58 85 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.83 $Y=1.21
+ $X2=6.83 $Y2=1.295
r186 58 60 32.0379 $w=2.48e-07 $l=6.95e-07 $layer=LI1_cond $X=6.83 $Y=1.21
+ $X2=6.83 $Y2=0.515
r187 57 84 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.015 $Y=1.295
+ $X2=5.93 $Y2=1.295
r188 56 85 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.705 $Y=1.295
+ $X2=6.83 $Y2=1.295
r189 56 57 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=6.705 $Y=1.295
+ $X2=6.015 $Y2=1.295
r190 52 84 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.93 $Y=1.21
+ $X2=5.93 $Y2=1.295
r191 52 54 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=5.93 $Y=1.21
+ $X2=5.93 $Y2=0.515
r192 51 83 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.155 $Y=1.295
+ $X2=5.03 $Y2=1.295
r193 50 84 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.845 $Y=1.295
+ $X2=5.93 $Y2=1.295
r194 50 51 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.845 $Y=1.295
+ $X2=5.155 $Y2=1.295
r195 46 83 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.03 $Y=1.21
+ $X2=5.03 $Y2=1.295
r196 46 48 32.0379 $w=2.48e-07 $l=6.95e-07 $layer=LI1_cond $X=5.03 $Y=1.21
+ $X2=5.03 $Y2=0.515
r197 44 83 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.905 $Y=1.295
+ $X2=5.03 $Y2=1.295
r198 44 45 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.905 $Y=1.295
+ $X2=4.225 $Y2=1.295
r199 41 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.14 $Y=1.21
+ $X2=4.225 $Y2=1.295
r200 41 43 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=4.14 $Y=1.21
+ $X2=4.14 $Y2=0.515
r201 40 43 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=4.14 $Y=0.425
+ $X2=4.14 $Y2=0.515
r202 39 78 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.375 $Y=0.34
+ $X2=3.21 $Y2=0.34
r203 38 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.055 $Y=0.34
+ $X2=4.14 $Y2=0.425
r204 38 39 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.055 $Y=0.34
+ $X2=3.375 $Y2=0.34
r205 37 73 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.375 $Y=0.34
+ $X2=2.21 $Y2=0.34
r206 36 78 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.045 $Y=0.34
+ $X2=3.21 $Y2=0.34
r207 36 37 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.045 $Y=0.34
+ $X2=2.375 $Y2=0.34
r208 35 68 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.375 $Y=0.34
+ $X2=1.21 $Y2=0.34
r209 34 73 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.045 $Y=0.34
+ $X2=2.21 $Y2=0.34
r210 34 35 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.045 $Y=0.34
+ $X2=1.375 $Y2=0.34
r211 32 68 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.045 $Y=0.34
+ $X2=1.21 $Y2=0.34
r212 32 33 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=1.045 $Y=0.34
+ $X2=0.445 $Y2=0.34
r213 28 33 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=0.425
+ $X2=0.445 $Y2=0.34
r214 28 30 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=0.28 $Y=0.425
+ $X2=0.28 $Y2=0.55
r215 9 66 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.58
+ $Y=0.37 $X2=7.72 $Y2=0.515
r216 8 60 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.65
+ $Y=0.37 $X2=6.79 $Y2=0.515
r217 7 54 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.79
+ $Y=0.37 $X2=5.93 $Y2=0.515
r218 6 48 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.93
+ $Y=0.37 $X2=5.07 $Y2=0.515
r219 5 43 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4 $Y=0.37
+ $X2=4.14 $Y2=0.515
r220 4 81 182 $w=1.7e-07 $l=2.86182e-07 $layer=licon1_NDIFF $count=1 $X=3
+ $Y=0.37 $X2=3.21 $Y2=0.55
r221 3 76 182 $w=1.7e-07 $l=2.86182e-07 $layer=licon1_NDIFF $count=1 $X=2
+ $Y=0.37 $X2=2.21 $Y2=0.55
r222 2 71 182 $w=1.7e-07 $l=2.86182e-07 $layer=licon1_NDIFF $count=1 $X=1
+ $Y=0.37 $X2=1.21 $Y2=0.55
r223 1 30 91 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_LS__EINVP_8%VGND 1 2 3 4 5 18 22 26 30 32 34 37 38 39 41
+ 49 58 62 68 71 74 78
c111 18 0 1.9142e-19 $X=4.57 $Y=0.515
r112 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r113 74 75 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r114 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r115 66 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=8.88
+ $Y2=0
r116 66 75 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=7.44
+ $Y2=0
r117 65 66 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r118 63 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.455 $Y=0 $X2=7.29
+ $Y2=0
r119 63 65 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=7.455 $Y=0 $X2=8.4
+ $Y2=0
r120 62 77 4.01281 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=8.675 $Y=0
+ $X2=8.897 $Y2=0
r121 62 65 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=8.675 $Y=0 $X2=8.4
+ $Y2=0
r122 61 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r123 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r124 58 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.125 $Y=0 $X2=7.29
+ $Y2=0
r125 58 60 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=7.125 $Y=0
+ $X2=6.96 $Y2=0
r126 57 61 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.96
+ $Y2=0
r127 57 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.52
+ $Y2=0
r128 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r129 54 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.665 $Y=0 $X2=5.5
+ $Y2=0
r130 54 56 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=5.665 $Y=0 $X2=6
+ $Y2=0
r131 53 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r132 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r133 50 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.735 $Y=0 $X2=4.57
+ $Y2=0
r134 50 52 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.735 $Y=0
+ $X2=5.04 $Y2=0
r135 49 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.335 $Y=0 $X2=5.5
+ $Y2=0
r136 49 52 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.335 $Y=0 $X2=5.04
+ $Y2=0
r137 47 48 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r138 44 48 1.07034 $w=4.9e-07 $l=3.84e-06 $layer=MET1_cond $X=0.24 $Y=0 $X2=4.08
+ $Y2=0
r139 43 47 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=4.08
+ $Y2=0
r140 43 44 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r141 41 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.405 $Y=0 $X2=4.57
+ $Y2=0
r142 41 47 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=4.405 $Y=0
+ $X2=4.08 $Y2=0
r143 39 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r144 39 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r145 39 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r146 37 56 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=6.195 $Y=0 $X2=6
+ $Y2=0
r147 37 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.195 $Y=0 $X2=6.36
+ $Y2=0
r148 36 60 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=6.525 $Y=0
+ $X2=6.96 $Y2=0
r149 36 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.525 $Y=0 $X2=6.36
+ $Y2=0
r150 32 77 3.19941 $w=2.6e-07 $l=1.27609e-07 $layer=LI1_cond $X=8.805 $Y=0.085
+ $X2=8.897 $Y2=0
r151 32 34 18.6164 $w=2.58e-07 $l=4.2e-07 $layer=LI1_cond $X=8.805 $Y=0.085
+ $X2=8.805 $Y2=0.505
r152 28 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.29 $Y=0.085
+ $X2=7.29 $Y2=0
r153 28 30 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=7.29 $Y=0.085
+ $X2=7.29 $Y2=0.515
r154 24 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.36 $Y=0.085
+ $X2=6.36 $Y2=0
r155 24 26 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=6.36 $Y=0.085
+ $X2=6.36 $Y2=0.515
r156 20 71 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.5 $Y=0.085 $X2=5.5
+ $Y2=0
r157 20 22 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=5.5 $Y=0.085
+ $X2=5.5 $Y2=0.515
r158 16 68 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.57 $Y=0.085
+ $X2=4.57 $Y2=0
r159 16 18 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=4.57 $Y=0.085
+ $X2=4.57 $Y2=0.515
r160 5 34 91 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=2 $X=8.63
+ $Y=0.37 $X2=8.77 $Y2=0.505
r161 4 30 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=7.08
+ $Y=0.37 $X2=7.29 $Y2=0.515
r162 3 26 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.22
+ $Y=0.37 $X2=6.36 $Y2=0.515
r163 2 22 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.36
+ $Y=0.37 $X2=5.5 $Y2=0.515
r164 1 18 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.43
+ $Y=0.37 $X2=4.57 $Y2=0.515
.ends

