* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
M1000 VPWR a_27_368# X VPB phighvt w=1.12e+06u l=150000u
+  ad=1.5282e+12p pd=9.39e+06u as=3.36e+11p ps=2.84e+06u
M1001 X a_27_368# VGND VNB nshort w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=7.498e+11p ps=6.7e+06u
M1002 a_195_74# B1 a_117_74# VNB nshort w=740000u l=150000u
+  ad=4.662e+11p pd=4.22e+06u as=1.776e+11p ps=1.96e+06u
M1003 VGND a_27_368# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR C1 a_27_368# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=5.95e+11p ps=5.19e+06u
M1005 VPWR A1 a_314_368# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=3.2e+11p ps=2.64e+06u
M1006 X a_27_368# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND A2 a_195_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_27_368# B1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_117_74# C1 a_27_368# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1010 a_195_74# A1 VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_314_368# A2 a_27_368# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
