* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__clkinv_16 A VGND VNB VPB VPWR Y
M1000 VPWR A Y VPB phighvt w=1.12e+06u l=150000u
+  ad=4.4688e+12p pd=3.71e+07u as=4.0992e+12p ps=3.42e+07u
M1001 Y A VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 VGND A Y VNB nshort w=420000u l=150000u
+  ad=1.83765e+12p pd=1.762e+07u as=9.408e+11p ps=1.12e+07u
M1003 Y A VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND A Y VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y A VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y A VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y A VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y A VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y A VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR A Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND A Y VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Y A VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR A Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR A Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y A VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Y A VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND A Y VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 Y A VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR A Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 Y A VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 Y A VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND A Y VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 Y A VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 Y A VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPWR A Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 Y A VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 Y A VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VPWR A Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VGND A Y VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VGND A Y VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 Y A VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 VPWR A Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VPWR A Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 VGND A Y VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 VPWR A Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 Y A VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 VPWR A Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 VPWR A Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 Y A VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
