* File: sky130_fd_sc_ls__a2111o_2.spice
* Created: Fri Aug 28 12:47:31 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__a2111o_2.pex.spice"
.subckt sky130_fd_sc_ls__a2111o_2  VNB VPB D1 C1 B1 A2 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A2	A2
* B1	B1
* C1	C1
* D1	D1
* VPB	VPB
* VNB	VNB
MM1005 N_VGND_M1005_d N_A_91_244#_M1005_g N_X_M1005_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1961 AS=0.1036 PD=2.01 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1006 N_VGND_M1006_d N_A_91_244#_M1006_g N_X_M1005_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1961 AS=0.1036 PD=2.01 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1013 N_VGND_M1013_d N_D1_M1013_g N_A_91_244#_M1013_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1184 AS=0.1961 PD=1.06 PS=2.01 NRD=3.24 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75002.2 A=0.111 P=1.78 MULT=1
MM1004 N_A_91_244#_M1004_d N_C1_M1004_g N_VGND_M1013_d VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1184 PD=1.02 PS=1.06 NRD=0 NRS=3.24 M=1 R=4.93333 SA=75000.7
+ SB=75001.7 A=0.111 P=1.78 MULT=1
MM1012 N_VGND_M1012_d N_B1_M1012_g N_A_91_244#_M1004_d VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=1.31 PS=1.02 NRD=27.564 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75001.3 A=0.111 P=1.78 MULT=1
MM1007 A_771_74# N_A2_M1007_g N_VGND_M1012_d VNB NSHORT L=0.15 W=0.74 AD=0.0777
+ AS=0.2109 PD=0.95 PS=1.31 NRD=8.1 NRS=19.452 M=1 R=4.93333 SA=75001.8
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1008 N_A_91_244#_M1008_d N_A1_M1008_g A_771_74# VNB NSHORT L=0.15 W=0.74
+ AD=0.1961 AS=0.0777 PD=2.01 PS=0.95 NRD=0 NRS=8.1 M=1 R=4.93333 SA=75002.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1009 N_X_M1009_d N_A_91_244#_M1009_g N_VPWR_M1009_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.308 PD=1.42 PS=2.79 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.6 A=0.168 P=2.54 MULT=1
MM1010 N_X_M1009_d N_A_91_244#_M1010_g N_VPWR_M1010_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.308 PD=1.42 PS=2.79 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.6 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1002 A_444_368# N_D1_M1002_g N_A_91_244#_M1002_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.1344 AS=0.308 PD=1.36 PS=2.79 NRD=11.426 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75002.2 A=0.168 P=2.54 MULT=1
MM1003 A_522_368# N_C1_M1003_g A_444_368# VPB PHIGHVT L=0.15 W=1.12 AD=0.2184
+ AS=0.1344 PD=1.51 PS=1.36 NRD=24.6053 NRS=11.426 M=1 R=7.46667 SA=75000.6
+ SB=75001.8 A=0.168 P=2.54 MULT=1
MM1001 N_A_630_368#_M1001_d N_B1_M1001_g A_522_368# VPB PHIGHVT L=0.15 W=1.12
+ AD=0.2184 AS=0.2184 PD=1.51 PS=1.51 NRD=5.2599 NRS=24.6053 M=1 R=7.46667
+ SA=75001.1 SB=75001.3 A=0.168 P=2.54 MULT=1
MM1011 N_VPWR_M1011_d N_A2_M1011_g N_A_630_368#_M1001_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.2184 AS=0.2184 PD=1.51 PS=1.51 NRD=5.2599 NRS=14.0658 M=1
+ R=7.46667 SA=75001.7 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1000 N_A_630_368#_M1000_d N_A1_M1000_g N_VPWR_M1011_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.308 AS=0.2184 PD=2.79 PS=1.51 NRD=1.7533 NRS=14.0658 M=1 R=7.46667
+ SA=75002.2 SB=75000.2 A=0.168 P=2.54 MULT=1
DX14_noxref VNB VPB NWDIODE A=9.6348 P=14.08
c_80 VPB 0 1.2388e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_ls__a2111o_2.pxi.spice"
*
.ends
*
*
