* NGSPICE file created from sky130_fd_sc_ls__sedfxtp_4.ext - technology: sky130A

.subckt sky130_fd_sc_ls__sedfxtp_4 CLK D DE SCD SCE VGND VNB VPB VPWR Q
M1000 a_135_74# D a_37_464# VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=2.373e+11p ps=2.81e+06u
M1001 a_661_113# SCE a_1044_125# VNB nshort w=420000u l=150000u
+  ad=5.502e+11p pd=5.14e+06u as=8.82e+10p ps=1.26e+06u
M1002 a_1943_53# a_1756_97# VPWR VPB phighvt w=840000u l=150000u
+  ad=2.31e+11p pd=2.23e+06u as=3.30785e+12p ps=2.82e+07u
M1003 VPWR a_2403_74# Q VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=6.72e+11p ps=5.68e+06u
M1004 VGND DE a_177_290# VNB nshort w=420000u l=150000u
+  ad=2.3264e+12p pd=2.159e+07u as=1.197e+11p ps=1.41e+06u
M1005 VPWR a_177_290# a_126_464# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1006 a_37_464# a_545_87# a_572_463# VPB phighvt w=640000u l=150000u
+  ad=3.808e+11p pd=3.75e+06u as=1.536e+11p ps=1.76e+06u
M1007 a_1044_125# SCD VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_2403_74# a_1313_74# a_2292_392# VPB phighvt w=1e+06u l=150000u
+  ad=3.049e+11p pd=2.72e+06u as=8.1e+11p ps=3.62e+06u
M1009 VPWR a_1943_53# a_1899_508# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.386e+11p ps=1.5e+06u
M1010 VPWR DE a_177_290# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.888e+11p ps=1.87e+06u
M1011 a_1510_74# a_1313_74# VGND VNB nshort w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1012 a_1071_455# SCD VPWR VPB phighvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1013 a_2498_74# a_1313_74# a_2403_74# VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=1.915e+11p ps=1.93e+06u
M1014 VGND a_545_87# a_2498_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_661_113# SCE a_37_464# VPB phighvt w=640000u l=150000u
+  ad=4.707e+11p pd=5.06e+06u as=0p ps=0u
M1016 a_545_87# a_2403_74# VGND VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1017 a_1510_74# a_1313_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.08e+11p pd=2.79e+06u as=0p ps=0u
M1018 a_1756_97# a_1510_74# a_661_113# VPB phighvt w=420000u l=150000u
+  ad=1.26e+11p pd=1.44e+06u as=0p ps=0u
M1019 Q a_2403_74# VGND VNB nshort w=740000u l=150000u
+  ad=4.255e+11p pd=4.11e+06u as=0p ps=0u
M1020 a_37_464# a_545_87# a_497_113# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1021 a_661_113# a_631_87# a_37_464# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_1313_74# CLK VGND VNB nshort w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1023 a_126_464# D a_37_464# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VPWR a_2403_74# Q VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_1899_508# a_1313_74# a_1756_97# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_2403_74# a_1510_74# a_2331_74# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=1.344e+11p ps=1.7e+06u
M1027 VGND a_1943_53# a_1858_79# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.785e+11p ps=1.69e+06u
M1028 a_572_463# DE VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VGND DE a_135_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VPWR a_545_87# a_2586_508# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1031 a_545_87# a_2403_74# VPWR VPB phighvt w=640000u l=150000u
+  ad=1.76e+11p pd=1.83e+06u as=0p ps=0u
M1032 a_1858_79# a_1510_74# a_1756_97# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.6695e+11p ps=1.74e+06u
M1033 Q a_2403_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_661_113# a_631_87# a_1071_455# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_497_113# a_177_290# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 VGND a_2403_74# Q VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_1756_97# a_1313_74# a_661_113# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 Q a_2403_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 Q a_2403_74# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1040 VGND a_2403_74# Q VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1041 a_1313_74# CLK VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.08e+11p pd=2.79e+06u as=0p ps=0u
M1042 VGND SCE a_631_87# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1043 a_2292_392# a_1943_53# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1044 VPWR SCE a_631_87# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1045 a_2586_508# a_1510_74# a_2403_74# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1046 a_1943_53# a_1756_97# VGND VNB nshort w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=0p ps=0u
M1047 a_2331_74# a_1943_53# VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

