* File: sky130_fd_sc_ls__o22ai_1.pxi.spice
* Created: Fri Aug 28 13:49:15 2020
* 
x_PM_SKY130_FD_SC_LS__O22AI_1%B1 N_B1_c_44_n N_B1_M1007_g N_B1_c_45_n
+ N_B1_M1000_g B1 PM_SKY130_FD_SC_LS__O22AI_1%B1
x_PM_SKY130_FD_SC_LS__O22AI_1%B2 N_B2_c_68_n N_B2_M1005_g N_B2_M1002_g B2
+ N_B2_c_70_n PM_SKY130_FD_SC_LS__O22AI_1%B2
x_PM_SKY130_FD_SC_LS__O22AI_1%A2 N_A2_c_95_n N_A2_M1006_g N_A2_M1001_g A2
+ N_A2_c_97_n PM_SKY130_FD_SC_LS__O22AI_1%A2
x_PM_SKY130_FD_SC_LS__O22AI_1%A1 N_A1_c_128_n N_A1_M1004_g N_A1_M1003_g A1 A1
+ N_A1_c_131_n PM_SKY130_FD_SC_LS__O22AI_1%A1
x_PM_SKY130_FD_SC_LS__O22AI_1%VPWR N_VPWR_M1000_s N_VPWR_M1004_d N_VPWR_c_155_n
+ N_VPWR_c_156_n N_VPWR_c_157_n N_VPWR_c_158_n N_VPWR_c_159_n N_VPWR_c_160_n
+ VPWR N_VPWR_c_154_n PM_SKY130_FD_SC_LS__O22AI_1%VPWR
x_PM_SKY130_FD_SC_LS__O22AI_1%Y N_Y_M1007_d N_Y_M1005_d N_Y_c_180_n Y Y
+ N_Y_c_182_n N_Y_c_181_n PM_SKY130_FD_SC_LS__O22AI_1%Y
x_PM_SKY130_FD_SC_LS__O22AI_1%A_27_74# N_A_27_74#_M1007_s N_A_27_74#_M1002_d
+ N_A_27_74#_M1003_d N_A_27_74#_c_207_n N_A_27_74#_c_208_n N_A_27_74#_c_209_n
+ N_A_27_74#_c_221_n N_A_27_74#_c_210_n N_A_27_74#_c_211_n N_A_27_74#_c_212_n
+ PM_SKY130_FD_SC_LS__O22AI_1%A_27_74#
x_PM_SKY130_FD_SC_LS__O22AI_1%VGND N_VGND_M1001_d N_VGND_c_248_n N_VGND_c_249_n
+ N_VGND_c_250_n VGND N_VGND_c_251_n N_VGND_c_252_n
+ PM_SKY130_FD_SC_LS__O22AI_1%VGND
cc_1 VNB N_B1_c_44_n 0.0245603f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.22
cc_2 VNB N_B1_c_45_n 0.0802438f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.765
cc_3 VNB B1 0.00820169f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_B2_c_68_n 0.0253517f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.22
cc_5 VNB N_B2_M1002_g 0.0285891f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=2.4
cc_6 VNB N_B2_c_70_n 0.00694829f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.295
cc_7 VNB N_A2_c_95_n 0.026988f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.22
cc_8 VNB N_A2_M1001_g 0.0268957f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=2.4
cc_9 VNB N_A2_c_97_n 0.00181735f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.295
cc_10 VNB N_A1_c_128_n 0.0199821f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.22
cc_11 VNB N_A1_M1003_g 0.0317431f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=2.4
cc_12 VNB A1 0.0177202f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.385
cc_13 VNB N_A1_c_131_n 0.0481093f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.385
cc_14 VNB N_VPWR_c_154_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_Y_c_180_n 0.00809472f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.385
cc_16 VNB N_Y_c_181_n 0.00612152f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_27_74#_c_207_n 0.0200157f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.295
cc_18 VNB N_A_27_74#_c_208_n 0.00778015f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_27_74#_c_209_n 0.00972033f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.385
cc_20 VNB N_A_27_74#_c_210_n 0.0168726f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_27_74#_c_211_n 0.00894964f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_27_74#_c_212_n 0.02581f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_248_n 0.0095417f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=2.4
cc_24 VNB N_VGND_c_249_n 0.0477009f $X=-0.19 $Y=-0.245 $X2=0.42 $Y2=1.385
cc_25 VNB N_VGND_c_250_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.385
cc_26 VNB N_VGND_c_251_n 0.0221746f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_252_n 0.188569f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VPB N_B1_c_45_n 0.0269271f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.765
cc_29 VPB N_B2_c_68_n 0.0275518f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.22
cc_30 VPB N_B2_c_70_n 0.00274883f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=1.295
cc_31 VPB N_A2_c_95_n 0.0293774f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.22
cc_32 VPB N_A2_c_97_n 0.00718364f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=1.295
cc_33 VPB N_A1_c_128_n 0.0275505f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.22
cc_34 VPB A1 0.0189556f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=1.385
cc_35 VPB N_VPWR_c_155_n 0.0125099f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_36 VPB N_VPWR_c_156_n 0.0594576f $X=-0.19 $Y=1.66 $X2=0.42 $Y2=1.385
cc_37 VPB N_VPWR_c_157_n 0.0485725f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=1.385
cc_38 VPB N_VPWR_c_158_n 0.0115308f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_39 VPB N_VPWR_c_159_n 0.0498348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_40 VPB N_VPWR_c_160_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_41 VPB N_VPWR_c_154_n 0.0792335f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_42 VPB N_Y_c_182_n 0.00628825f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_43 VPB N_Y_c_181_n 0.00130347f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_44 N_B1_c_45_n N_B2_c_68_n 0.0822463f $X=0.635 $Y=1.765 $X2=-0.19 $Y2=-0.245
cc_45 N_B1_c_44_n N_B2_M1002_g 0.0175332f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_46 N_B1_c_45_n N_B2_c_70_n 4.4696e-19 $X=0.635 $Y=1.765 $X2=0 $Y2=0
cc_47 N_B1_c_45_n N_VPWR_c_156_n 0.0315674f $X=0.635 $Y=1.765 $X2=0 $Y2=0
cc_48 B1 N_VPWR_c_156_n 0.0192059f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_49 N_B1_c_45_n N_VPWR_c_159_n 0.00366292f $X=0.635 $Y=1.765 $X2=0 $Y2=0
cc_50 N_B1_c_45_n N_VPWR_c_154_n 0.00605201f $X=0.635 $Y=1.765 $X2=0 $Y2=0
cc_51 N_B1_c_44_n N_Y_c_180_n 0.0041759f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_52 N_B1_c_45_n N_Y_c_180_n 3.73516e-19 $X=0.635 $Y=1.765 $X2=0 $Y2=0
cc_53 N_B1_c_45_n N_Y_c_182_n 0.0276669f $X=0.635 $Y=1.765 $X2=0 $Y2=0
cc_54 N_B1_c_44_n N_Y_c_181_n 0.00431169f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_55 N_B1_c_45_n N_Y_c_181_n 0.0235978f $X=0.635 $Y=1.765 $X2=0 $Y2=0
cc_56 B1 N_Y_c_181_n 0.0260309f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_57 N_B1_c_44_n N_A_27_74#_c_207_n 0.0118446f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_58 N_B1_c_45_n N_A_27_74#_c_207_n 0.00199342f $X=0.635 $Y=1.765 $X2=0 $Y2=0
cc_59 B1 N_A_27_74#_c_207_n 0.0261036f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_60 N_B1_c_44_n N_A_27_74#_c_208_n 0.0116366f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_61 N_B1_c_44_n N_A_27_74#_c_209_n 0.00167496f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_62 N_B1_c_44_n N_VGND_c_249_n 0.00286814f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_63 N_B1_c_44_n N_VGND_c_252_n 0.00361864f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_64 N_B2_c_68_n N_A2_c_95_n 0.0529063f $X=1.055 $Y=1.765 $X2=-0.19 $Y2=-0.245
cc_65 N_B2_c_70_n N_A2_c_95_n 0.00269474f $X=1.13 $Y=1.515 $X2=-0.19 $Y2=-0.245
cc_66 N_B2_M1002_g N_A2_M1001_g 0.0250863f $X=1.22 $Y=0.74 $X2=0 $Y2=0
cc_67 N_B2_c_68_n N_A2_c_97_n 5.32787e-19 $X=1.055 $Y=1.765 $X2=0 $Y2=0
cc_68 N_B2_c_70_n N_A2_c_97_n 0.0282656f $X=1.13 $Y=1.515 $X2=0 $Y2=0
cc_69 N_B2_c_68_n N_VPWR_c_159_n 0.00291513f $X=1.055 $Y=1.765 $X2=0 $Y2=0
cc_70 N_B2_c_68_n N_VPWR_c_154_n 0.00360271f $X=1.055 $Y=1.765 $X2=0 $Y2=0
cc_71 N_B2_c_68_n N_Y_c_180_n 7.13242e-19 $X=1.055 $Y=1.765 $X2=0 $Y2=0
cc_72 N_B2_M1002_g N_Y_c_180_n 0.00587202f $X=1.22 $Y=0.74 $X2=0 $Y2=0
cc_73 N_B2_c_70_n N_Y_c_180_n 0.00676358f $X=1.13 $Y=1.515 $X2=0 $Y2=0
cc_74 N_B2_c_68_n N_Y_c_182_n 0.0459731f $X=1.055 $Y=1.765 $X2=0 $Y2=0
cc_75 N_B2_c_70_n N_Y_c_182_n 0.0266535f $X=1.13 $Y=1.515 $X2=0 $Y2=0
cc_76 N_B2_c_68_n N_Y_c_181_n 0.00488074f $X=1.055 $Y=1.765 $X2=0 $Y2=0
cc_77 N_B2_M1002_g N_Y_c_181_n 0.00318696f $X=1.22 $Y=0.74 $X2=0 $Y2=0
cc_78 N_B2_c_70_n N_Y_c_181_n 0.0325254f $X=1.13 $Y=1.515 $X2=0 $Y2=0
cc_79 N_B2_M1002_g N_A_27_74#_c_208_n 0.0157492f $X=1.22 $Y=0.74 $X2=0 $Y2=0
cc_80 N_B2_M1002_g N_A_27_74#_c_211_n 0.00100357f $X=1.22 $Y=0.74 $X2=0 $Y2=0
cc_81 N_B2_M1002_g N_VGND_c_249_n 0.00286838f $X=1.22 $Y=0.74 $X2=0 $Y2=0
cc_82 N_B2_M1002_g N_VGND_c_252_n 0.0035893f $X=1.22 $Y=0.74 $X2=0 $Y2=0
cc_83 N_A2_c_95_n N_A1_c_128_n 0.0556315f $X=1.625 $Y=1.765 $X2=-0.19 $Y2=-0.245
cc_84 N_A2_M1001_g N_A1_c_128_n 0.00181425f $X=1.72 $Y=0.74 $X2=-0.19 $Y2=-0.245
cc_85 N_A2_c_97_n N_A1_c_128_n 6.98729e-19 $X=1.7 $Y=1.515 $X2=-0.19 $Y2=-0.245
cc_86 N_A2_M1001_g N_A1_M1003_g 0.0250949f $X=1.72 $Y=0.74 $X2=0 $Y2=0
cc_87 N_A2_c_95_n A1 0.00247461f $X=1.625 $Y=1.765 $X2=0 $Y2=0
cc_88 N_A2_M1001_g A1 0.00123883f $X=1.72 $Y=0.74 $X2=0 $Y2=0
cc_89 N_A2_c_97_n A1 0.0350656f $X=1.7 $Y=1.515 $X2=0 $Y2=0
cc_90 N_A2_c_95_n N_VPWR_c_157_n 0.00512579f $X=1.625 $Y=1.765 $X2=0 $Y2=0
cc_91 N_A2_c_95_n N_VPWR_c_159_n 0.00461464f $X=1.625 $Y=1.765 $X2=0 $Y2=0
cc_92 N_A2_c_95_n N_VPWR_c_154_n 0.00911823f $X=1.625 $Y=1.765 $X2=0 $Y2=0
cc_93 N_A2_c_95_n N_Y_c_182_n 0.00741073f $X=1.625 $Y=1.765 $X2=0 $Y2=0
cc_94 N_A2_M1001_g N_A_27_74#_c_208_n 0.00272067f $X=1.72 $Y=0.74 $X2=0 $Y2=0
cc_95 N_A2_M1001_g N_A_27_74#_c_221_n 0.00730256f $X=1.72 $Y=0.74 $X2=0 $Y2=0
cc_96 N_A2_c_95_n N_A_27_74#_c_210_n 4.60538e-19 $X=1.625 $Y=1.765 $X2=0 $Y2=0
cc_97 N_A2_M1001_g N_A_27_74#_c_210_n 0.0120407f $X=1.72 $Y=0.74 $X2=0 $Y2=0
cc_98 N_A2_c_97_n N_A_27_74#_c_210_n 0.0118018f $X=1.7 $Y=1.515 $X2=0 $Y2=0
cc_99 N_A2_c_95_n N_A_27_74#_c_211_n 8.2764e-19 $X=1.625 $Y=1.765 $X2=0 $Y2=0
cc_100 N_A2_M1001_g N_A_27_74#_c_211_n 0.00102901f $X=1.72 $Y=0.74 $X2=0 $Y2=0
cc_101 N_A2_c_97_n N_A_27_74#_c_211_n 0.00940645f $X=1.7 $Y=1.515 $X2=0 $Y2=0
cc_102 N_A2_M1001_g N_A_27_74#_c_212_n 6.18925e-19 $X=1.72 $Y=0.74 $X2=0 $Y2=0
cc_103 N_A2_M1001_g N_VGND_c_248_n 0.00522681f $X=1.72 $Y=0.74 $X2=0 $Y2=0
cc_104 N_A2_M1001_g N_VGND_c_249_n 0.00432337f $X=1.72 $Y=0.74 $X2=0 $Y2=0
cc_105 N_A2_M1001_g N_VGND_c_252_n 0.00817838f $X=1.72 $Y=0.74 $X2=0 $Y2=0
cc_106 N_A1_c_128_n N_VPWR_c_157_n 0.0270384f $X=2.195 $Y=1.765 $X2=0 $Y2=0
cc_107 A1 N_VPWR_c_157_n 0.0265674f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_108 N_A1_c_128_n N_VPWR_c_159_n 0.00413917f $X=2.195 $Y=1.765 $X2=0 $Y2=0
cc_109 N_A1_c_128_n N_VPWR_c_154_n 0.00818781f $X=2.195 $Y=1.765 $X2=0 $Y2=0
cc_110 N_A1_M1003_g N_A_27_74#_c_221_n 5.91875e-19 $X=2.29 $Y=0.74 $X2=0 $Y2=0
cc_111 N_A1_c_128_n N_A_27_74#_c_210_n 0.00286524f $X=2.195 $Y=1.765 $X2=0 $Y2=0
cc_112 N_A1_M1003_g N_A_27_74#_c_210_n 0.0129307f $X=2.29 $Y=0.74 $X2=0 $Y2=0
cc_113 A1 N_A_27_74#_c_210_n 0.0509938f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_114 N_A1_c_131_n N_A_27_74#_c_210_n 0.00708493f $X=2.61 $Y=1.465 $X2=0 $Y2=0
cc_115 N_A1_M1003_g N_A_27_74#_c_212_n 0.00981823f $X=2.29 $Y=0.74 $X2=0 $Y2=0
cc_116 N_A1_M1003_g N_VGND_c_248_n 0.00592235f $X=2.29 $Y=0.74 $X2=0 $Y2=0
cc_117 N_A1_M1003_g N_VGND_c_251_n 0.00434272f $X=2.29 $Y=0.74 $X2=0 $Y2=0
cc_118 N_A1_M1003_g N_VGND_c_252_n 0.00825253f $X=2.29 $Y=0.74 $X2=0 $Y2=0
cc_119 N_VPWR_c_159_n N_Y_c_182_n 0.0404856f $X=2.255 $Y=3.33 $X2=0 $Y2=0
cc_120 N_VPWR_c_154_n N_Y_c_182_n 0.0329608f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_121 N_VPWR_c_156_n N_Y_c_181_n 0.0945277f $X=0.29 $Y=1.985 $X2=0 $Y2=0
cc_122 A_142_368# N_Y_c_182_n 0.00577415f $X=0.71 $Y=1.84 $X2=1.335 $Y2=2.115
cc_123 A_142_368# N_Y_c_181_n 7.03062e-19 $X=0.71 $Y=1.84 $X2=1.087 $Y2=1.95
cc_124 N_Y_M1007_d N_A_27_74#_c_208_n 0.00691776f $X=0.57 $Y=0.37 $X2=0 $Y2=0
cc_125 N_Y_c_180_n N_A_27_74#_c_208_n 0.0331049f $X=0.855 $Y=0.84 $X2=0 $Y2=0
cc_126 N_Y_c_180_n N_A_27_74#_c_211_n 0.00568934f $X=0.855 $Y=0.84 $X2=0 $Y2=0
cc_127 N_A_27_74#_c_210_n N_VGND_M1001_d 0.00374767f $X=2.34 $Y=1.045 $X2=-0.19
+ $Y2=-0.245
cc_128 N_A_27_74#_c_208_n N_VGND_c_248_n 0.0094172f $X=1.34 $Y=0.4 $X2=0 $Y2=0
cc_129 N_A_27_74#_c_210_n N_VGND_c_248_n 0.0248957f $X=2.34 $Y=1.045 $X2=0 $Y2=0
cc_130 N_A_27_74#_c_212_n N_VGND_c_248_n 0.0173003f $X=2.505 $Y=0.515 $X2=0
+ $Y2=0
cc_131 N_A_27_74#_c_208_n N_VGND_c_249_n 0.0581922f $X=1.34 $Y=0.4 $X2=0 $Y2=0
cc_132 N_A_27_74#_c_209_n N_VGND_c_249_n 0.0170692f $X=0.445 $Y=0.4 $X2=0 $Y2=0
cc_133 N_A_27_74#_c_212_n N_VGND_c_251_n 0.0145639f $X=2.505 $Y=0.515 $X2=0
+ $Y2=0
cc_134 N_A_27_74#_c_208_n N_VGND_c_252_n 0.0434237f $X=1.34 $Y=0.4 $X2=0 $Y2=0
cc_135 N_A_27_74#_c_209_n N_VGND_c_252_n 0.0123284f $X=0.445 $Y=0.4 $X2=0 $Y2=0
cc_136 N_A_27_74#_c_212_n N_VGND_c_252_n 0.0119984f $X=2.505 $Y=0.515 $X2=0
+ $Y2=0
