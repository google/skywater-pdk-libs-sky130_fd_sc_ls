* File: sky130_fd_sc_ls__ebufn_2.pex.spice
* Created: Wed Sep  2 11:05:59 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__EBUFN_2%A_84_48# 1 2 9 11 13 16 18 20 21 27 28 29 32
+ 36 40 42 43 48
c112 36 0 1.50682e-19 $X=4.04 $Y=2.715
r113 47 48 13.7358 $w=3.86e-07 $l=1.1e-07 $layer=POLY_cond $X=0.925 $Y=1.532
+ $X2=1.035 $Y2=1.532
r114 46 47 48.6995 $w=3.86e-07 $l=3.9e-07 $layer=POLY_cond $X=0.535 $Y=1.532
+ $X2=0.925 $Y2=1.532
r115 45 46 4.99482 $w=3.86e-07 $l=4e-08 $layer=POLY_cond $X=0.495 $Y=1.532
+ $X2=0.535 $Y2=1.532
r116 42 44 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=4.04 $Y=2.035
+ $X2=4.04 $Y2=2.325
r117 42 43 5.66838 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=4.04 $Y=2.035
+ $X2=4.04 $Y2=1.95
r118 40 43 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=4.12 $Y=1.03
+ $X2=4.12 $Y2=1.95
r119 34 44 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=4.04 $Y=2.41
+ $X2=4.04 $Y2=2.325
r120 34 36 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=4.04 $Y=2.41
+ $X2=4.04 $Y2=2.715
r121 30 40 9.06106 $w=3.63e-07 $l=1.82e-07 $layer=LI1_cond $X=4.022 $Y=0.848
+ $X2=4.022 $Y2=1.03
r122 30 32 10.5141 $w=3.63e-07 $l=3.33e-07 $layer=LI1_cond $X=4.022 $Y=0.848
+ $X2=4.022 $Y2=0.515
r123 28 44 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.875 $Y=2.325
+ $X2=4.04 $Y2=2.325
r124 28 29 113.519 $w=1.68e-07 $l=1.74e-06 $layer=LI1_cond $X=3.875 $Y=2.325
+ $X2=2.135 $Y2=2.325
r125 27 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.05 $Y=2.24
+ $X2=2.135 $Y2=2.325
r126 26 27 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=2.05 $Y=1.63
+ $X2=2.05 $Y2=2.24
r127 24 48 0.624352 $w=3.86e-07 $l=5e-09 $layer=POLY_cond $X=1.04 $Y=1.532
+ $X2=1.035 $Y2=1.532
r128 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.04
+ $Y=1.465 $X2=1.04 $Y2=1.465
r129 21 26 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.965 $Y=1.465
+ $X2=2.05 $Y2=1.63
r130 21 23 32.3033 $w=3.28e-07 $l=9.25e-07 $layer=LI1_cond $X=1.965 $Y=1.465
+ $X2=1.04 $Y2=1.465
r131 18 48 24.9932 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=1.035 $Y=1.765
+ $X2=1.035 $Y2=1.532
r132 18 20 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.035 $Y=1.765
+ $X2=1.035 $Y2=2.4
r133 14 47 24.9932 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=0.925 $Y=1.3
+ $X2=0.925 $Y2=1.532
r134 14 16 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.925 $Y=1.3
+ $X2=0.925 $Y2=0.74
r135 11 46 24.9932 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=0.535 $Y=1.765
+ $X2=0.535 $Y2=1.532
r136 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.535 $Y=1.765
+ $X2=0.535 $Y2=2.4
r137 7 45 24.9932 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=0.495 $Y=1.3
+ $X2=0.495 $Y2=1.532
r138 7 9 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.495 $Y=1.3
+ $X2=0.495 $Y2=0.74
r139 2 42 400 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=3.89
+ $Y=1.84 $X2=4.04 $Y2=2.035
r140 2 36 400 $w=1.7e-07 $l=9.47035e-07 $layer=licon1_PDIFF $count=1 $X=3.89
+ $Y=1.84 $X2=4.04 $Y2=2.715
r141 1 32 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.865
+ $Y=0.37 $X2=4.005 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__EBUFN_2%A_283_48# 1 2 7 9 10 11 12 14 15 17 22 24 26
+ 30 33
c72 15 0 6.40996e-20 $X=2.395 $Y=1.26
c73 7 0 1.83135e-19 $X=1.49 $Y=1.185
r74 29 33 7.77014 $w=6.83e-07 $l=4.45e-07 $layer=LI1_cond $X=2.56 $Y=0.667
+ $X2=3.005 $Y2=0.667
r75 29 30 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.56
+ $Y=0.49 $X2=2.56 $Y2=0.49
r76 24 26 9.91101 $w=2.48e-07 $l=2.15e-07 $layer=LI1_cond $X=2.725 $Y=1.945
+ $X2=2.94 $Y2=1.945
r77 23 30 118.906 $w=3.3e-07 $l=6.8e-07 $layer=POLY_cond $X=2.56 $Y=1.17
+ $X2=2.56 $Y2=0.49
r78 22 23 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.56
+ $Y=1.17 $X2=2.56 $Y2=1.17
r79 20 24 6.98653 $w=2.5e-07 $l=2.18746e-07 $layer=LI1_cond $X=2.56 $Y=1.82
+ $X2=2.725 $Y2=1.945
r80 20 22 22.6996 $w=3.28e-07 $l=6.5e-07 $layer=LI1_cond $X=2.56 $Y=1.82
+ $X2=2.56 $Y2=1.17
r81 19 29 5.02295 $w=3.3e-07 $l=3.43e-07 $layer=LI1_cond $X=2.56 $Y=1.01
+ $X2=2.56 $Y2=0.667
r82 19 22 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=2.56 $Y=1.01 $X2=2.56
+ $Y2=1.17
r83 18 23 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=2.56 $Y=1.185
+ $X2=2.56 $Y2=1.17
r84 16 17 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2 $Y=1.26 $X2=1.925
+ $Y2=1.26
r85 15 18 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=2.395 $Y=1.26
+ $X2=2.56 $Y2=1.185
r86 15 16 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.395 $Y=1.26 $X2=2
+ $Y2=1.26
r87 12 17 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.925 $Y=1.185
+ $X2=1.925 $Y2=1.26
r88 12 14 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.925 $Y=1.185
+ $X2=1.925 $Y2=0.74
r89 10 17 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.85 $Y=1.26
+ $X2=1.925 $Y2=1.26
r90 10 11 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.85 $Y=1.26
+ $X2=1.565 $Y2=1.26
r91 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.49 $Y=1.185
+ $X2=1.565 $Y2=1.26
r92 7 9 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.49 $Y=1.185
+ $X2=1.49 $Y2=0.74
r93 2 26 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=2.795
+ $Y=1.84 $X2=2.94 $Y2=1.985
r94 1 33 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=2.86
+ $Y=0.37 $X2=3.005 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__EBUFN_2%TE_B 1 3 4 5 6 8 9 11 13 16 18 19
c85 19 0 6.40996e-20 $X=3.12 $Y=1.295
c86 11 0 1.50682e-19 $X=3.165 $Y=1.765
c87 1 0 8.35221e-20 $X=1.535 $Y=1.765
r88 22 24 25.1677 $w=3.16e-07 $l=1.65e-07 $layer=POLY_cond $X=3.13 $Y=1.485
+ $X2=3.13 $Y2=1.65
r89 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.13
+ $Y=1.485 $X2=3.13 $Y2=1.485
r90 19 23 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=3.13 $Y=1.295
+ $X2=3.13 $Y2=1.485
r91 14 22 38.5382 $w=3.16e-07 $l=2.05122e-07 $layer=POLY_cond $X=3.22 $Y=1.32
+ $X2=3.13 $Y2=1.485
r92 14 16 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=3.22 $Y=1.32
+ $X2=3.22 $Y2=0.69
r93 11 24 30.9117 $w=3.16e-07 $l=1.31339e-07 $layer=POLY_cond $X=3.165 $Y=1.765
+ $X2=3.13 $Y2=1.65
r94 11 13 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.165 $Y=1.765
+ $X2=3.165 $Y2=2.34
r95 10 18 20.4101 $w=1.5e-07 $l=9.94987e-08 $layer=POLY_cond $X=2.245 $Y=1.65
+ $X2=2.155 $Y2=1.67
r96 9 24 20.1942 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.965 $Y=1.65
+ $X2=3.13 $Y2=1.65
r97 9 10 369.191 $w=1.5e-07 $l=7.2e-07 $layer=POLY_cond $X=2.965 $Y=1.65
+ $X2=2.245 $Y2=1.65
r98 6 18 5.30422 $w=1.5e-07 $l=9.5e-08 $layer=POLY_cond $X=2.155 $Y=1.765
+ $X2=2.155 $Y2=1.67
r99 6 8 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.155 $Y=1.765
+ $X2=2.155 $Y2=2.4
r100 4 18 20.4101 $w=1.5e-07 $l=9.94987e-08 $layer=POLY_cond $X=2.065 $Y=1.65
+ $X2=2.155 $Y2=1.67
r101 4 5 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=2.065 $Y=1.65
+ $X2=1.625 $Y2=1.65
r102 1 5 26.9307 $w=1.5e-07 $l=1.53542e-07 $layer=POLY_cond $X=1.535 $Y=1.765
+ $X2=1.625 $Y2=1.65
r103 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.535 $Y=1.765
+ $X2=1.535 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__EBUFN_2%A 3 5 7 8 12
r31 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.7
+ $Y=1.515 $X2=3.7 $Y2=1.515
r32 8 12 4.54912 $w=3.78e-07 $l=1.5e-07 $layer=LI1_cond $X=3.675 $Y=1.665
+ $X2=3.675 $Y2=1.515
r33 5 11 50.9845 $w=3.31e-07 $l=2.93684e-07 $layer=POLY_cond $X=3.815 $Y=1.765
+ $X2=3.72 $Y2=1.515
r34 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.815 $Y=1.765
+ $X2=3.815 $Y2=2.34
r35 1 11 38.6069 $w=3.31e-07 $l=1.96914e-07 $layer=POLY_cond $X=3.79 $Y=1.35
+ $X2=3.72 $Y2=1.515
r36 1 3 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.79 $Y=1.35 $X2=3.79
+ $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_LS__EBUFN_2%A_33_368# 1 2 3 12 14 15 16 19 24
c44 14 0 8.35221e-20 $X=1.145 $Y=2.99
r45 24 27 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=2.38 $Y=2.665
+ $X2=2.38 $Y2=2.78
r46 21 22 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=1.31 $Y=2.665
+ $X2=1.31 $Y2=2.99
r47 19 21 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=1.31 $Y=2.44
+ $X2=1.31 $Y2=2.665
r48 17 21 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.475 $Y=2.665
+ $X2=1.31 $Y2=2.665
r49 16 24 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.215 $Y=2.665
+ $X2=2.38 $Y2=2.665
r50 16 17 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=2.215 $Y=2.665
+ $X2=1.475 $Y2=2.665
r51 14 22 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.145 $Y=2.99
+ $X2=1.31 $Y2=2.99
r52 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.145 $Y=2.99
+ $X2=0.475 $Y2=2.99
r53 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.31 $Y=2.905
+ $X2=0.475 $Y2=2.99
r54 10 12 22.6996 $w=3.28e-07 $l=6.5e-07 $layer=LI1_cond $X=0.31 $Y=2.905
+ $X2=0.31 $Y2=2.255
r55 3 27 600 $w=1.7e-07 $l=1.01223e-06 $layer=licon1_PDIFF $count=1 $X=2.23
+ $Y=1.84 $X2=2.38 $Y2=2.78
r56 2 19 300 $w=1.7e-07 $l=6.9282e-07 $layer=licon1_PDIFF $count=2 $X=1.11
+ $Y=1.84 $X2=1.31 $Y2=2.44
r57 1 12 300 $w=1.7e-07 $l=4.82079e-07 $layer=licon1_PDIFF $count=2 $X=0.165
+ $Y=1.84 $X2=0.31 $Y2=2.255
.ends

.subckt PM_SKY130_FD_SC_LS__EBUFN_2%Z 1 2 9 12 15 17 20 21 22
c40 17 0 1.11307e-19 $X=0.705 $Y=1.13
c41 9 0 7.18276e-20 $X=0.71 $Y=0.78
r42 21 22 15.8049 $w=3.48e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.975
+ $X2=1.68 $Y2=1.975
r43 18 21 7.40856 $w=3.48e-07 $l=2.25e-07 $layer=LI1_cond $X=0.975 $Y=1.975
+ $X2=1.2 $Y2=1.975
r44 18 20 0.164012 $w=3.5e-07 $l=5.20192e-07 $layer=LI1_cond $X=0.975 $Y=1.975
+ $X2=0.535 $Y2=1.8
r45 13 20 6.76825 $w=2.5e-07 $l=4.67707e-07 $layer=LI1_cond $X=0.81 $Y=2.15
+ $X2=0.535 $Y2=1.8
r46 13 15 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=0.81 $Y=2.15 $X2=0.81
+ $Y2=2.65
r47 12 20 6.76825 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.62 $Y=1.8 $X2=0.535
+ $Y2=1.8
r48 12 17 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.62 $Y=1.8 $X2=0.62
+ $Y2=1.13
r49 7 17 8.64139 $w=3.38e-07 $l=1.7e-07 $layer=LI1_cond $X=0.705 $Y=0.96
+ $X2=0.705 $Y2=1.13
r50 7 9 6.10117 $w=3.38e-07 $l=1.8e-07 $layer=LI1_cond $X=0.705 $Y=0.96
+ $X2=0.705 $Y2=0.78
r51 2 20 400 $w=1.7e-07 $l=2.56905e-07 $layer=licon1_PDIFF $count=1 $X=0.61
+ $Y=1.84 $X2=0.81 $Y2=1.97
r52 2 15 400 $w=1.7e-07 $l=9.04489e-07 $layer=licon1_PDIFF $count=1 $X=0.61
+ $Y=1.84 $X2=0.81 $Y2=2.65
r53 1 9 182 $w=1.7e-07 $l=4.74868e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.78
.ends

.subckt PM_SKY130_FD_SC_LS__EBUFN_2%VPWR 1 2 9 11 13 18 28 29 32 39
r47 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r48 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r49 32 35 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=1.845 $Y=3.005
+ $X2=1.845 $Y2=3.33
r50 29 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r51 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r52 26 39 11.015 $w=1.7e-07 $l=2.4e-07 $layer=LI1_cond $X=3.705 $Y=3.33
+ $X2=3.465 $Y2=3.33
r53 26 28 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=3.705 $Y=3.33
+ $X2=4.08 $Y2=3.33
r54 25 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r55 24 25 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r56 21 24 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=3.33 $X2=3.12
+ $Y2=3.33
r57 19 35 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.01 $Y=3.33
+ $X2=1.845 $Y2=3.33
r58 19 21 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=2.01 $Y=3.33 $X2=2.16
+ $Y2=3.33
r59 18 39 11.015 $w=1.7e-07 $l=2.4e-07 $layer=LI1_cond $X=3.225 $Y=3.33
+ $X2=3.465 $Y2=3.33
r60 18 24 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=3.225 $Y=3.33
+ $X2=3.12 $Y2=3.33
r61 16 36 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.68 $Y2=3.33
r62 15 16 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r63 13 35 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.68 $Y=3.33
+ $X2=1.845 $Y2=3.33
r64 13 15 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.68 $Y=3.33
+ $X2=0.24 $Y2=3.33
r65 11 25 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r66 11 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r67 11 21 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r68 7 39 1.96841 $w=4.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.465 $Y=3.245
+ $X2=3.465 $Y2=3.33
r69 7 9 13.7051 $w=4.78e-07 $l=5.5e-07 $layer=LI1_cond $X=3.465 $Y=3.245
+ $X2=3.465 $Y2=2.695
r70 2 9 600 $w=1.7e-07 $l=9.60937e-07 $layer=licon1_PDIFF $count=1 $X=3.24
+ $Y=1.84 $X2=3.465 $Y2=2.695
r71 1 32 600 $w=1.7e-07 $l=1.27711e-06 $layer=licon1_PDIFF $count=1 $X=1.61
+ $Y=1.84 $X2=1.845 $Y2=3.005
.ends

.subckt PM_SKY130_FD_SC_LS__EBUFN_2%A_27_74# 1 2 3 12 14 15 20 21 24
r41 22 24 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=2.1 $Y=0.96 $X2=2.1
+ $Y2=0.515
r42 20 22 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.975 $Y=1.045
+ $X2=2.1 $Y2=0.96
r43 20 21 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=1.975 $Y=1.045
+ $X2=1.375 $Y2=1.045
r44 17 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.21 $Y=0.96
+ $X2=1.375 $Y2=1.045
r45 17 19 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=1.21 $Y=0.96
+ $X2=1.21 $Y2=0.515
r46 16 19 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=1.21 $Y=0.425 $X2=1.21
+ $Y2=0.515
r47 14 16 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.045 $Y=0.34
+ $X2=1.21 $Y2=0.425
r48 14 15 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.045 $Y=0.34
+ $X2=0.365 $Y2=0.34
r49 10 15 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.24 $Y=0.425
+ $X2=0.365 $Y2=0.34
r50 10 12 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=0.24 $Y=0.425 $X2=0.24
+ $Y2=0.515
r51 3 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2 $Y=0.37
+ $X2=2.14 $Y2=0.515
r52 2 19 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=1 $Y=0.37
+ $X2=1.21 $Y2=0.515
r53 1 12 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__EBUFN_2%VGND 1 2 9 13 16 17 18 20 36 37 40
r46 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r47 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r48 34 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r49 33 34 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r50 30 33 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r51 28 40 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.795 $Y=0 $X2=1.67
+ $Y2=0
r52 28 30 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.795 $Y=0 $X2=2.16
+ $Y2=0
r53 27 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r54 26 27 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r55 23 27 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r56 22 26 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r57 22 23 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r58 20 40 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.545 $Y=0 $X2=1.67
+ $Y2=0
r59 20 26 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.545 $Y=0 $X2=1.2
+ $Y2=0
r60 18 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r61 18 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r62 18 30 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r63 16 33 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=3.34 $Y=0 $X2=3.12
+ $Y2=0
r64 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.34 $Y=0 $X2=3.505
+ $Y2=0
r65 15 36 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=3.67 $Y=0 $X2=4.08
+ $Y2=0
r66 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.67 $Y=0 $X2=3.505
+ $Y2=0
r67 11 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.505 $Y=0.085
+ $X2=3.505 $Y2=0
r68 11 13 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.505 $Y=0.085
+ $X2=3.505 $Y2=0.515
r69 7 40 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.67 $Y=0.085
+ $X2=1.67 $Y2=0
r70 7 9 24.8928 $w=2.48e-07 $l=5.4e-07 $layer=LI1_cond $X=1.67 $Y=0.085 $X2=1.67
+ $Y2=0.625
r71 2 13 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=3.295
+ $Y=0.37 $X2=3.505 $Y2=0.515
r72 1 9 182 $w=1.7e-07 $l=3.19374e-07 $layer=licon1_NDIFF $count=1 $X=1.565
+ $Y=0.37 $X2=1.71 $Y2=0.625
.ends

