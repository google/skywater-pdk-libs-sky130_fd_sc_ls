* File: sky130_fd_sc_ls__nand4_1.pex.spice
* Created: Fri Aug 28 13:34:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__NAND4_1%D 1 3 4 6 7
r26 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.74
+ $Y=1.385 $X2=0.74 $Y2=1.385
r27 7 11 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.74 $Y=1.295 $X2=0.74
+ $Y2=1.385
r28 4 10 38.9026 $w=2.7e-07 $l=2.05122e-07 $layer=POLY_cond $X=0.83 $Y=1.22
+ $X2=0.74 $Y2=1.385
r29 4 6 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.83 $Y=1.22 $X2=0.83
+ $Y2=0.74
r30 1 10 77.2841 $w=2.7e-07 $l=4.15812e-07 $layer=POLY_cond $X=0.815 $Y=1.765
+ $X2=0.74 $Y2=1.385
r31 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.815 $Y=1.765
+ $X2=0.815 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__NAND4_1%C 1 3 4 6 7 11
c29 11 0 1.64093e-19 $X=1.31 $Y=1.385
c30 1 0 3.78555e-20 $X=1.22 $Y=1.22
r31 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.31
+ $Y=1.385 $X2=1.31 $Y2=1.385
r32 7 11 3.42618 $w=3.68e-07 $l=1.1e-07 $layer=LI1_cond $X=1.2 $Y=1.365 $X2=1.31
+ $Y2=1.365
r33 4 10 77.2841 $w=2.7e-07 $l=4.01871e-07 $layer=POLY_cond $X=1.265 $Y=1.765
+ $X2=1.31 $Y2=1.385
r34 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.265 $Y=1.765
+ $X2=1.265 $Y2=2.4
r35 1 10 38.9026 $w=2.7e-07 $l=2.05122e-07 $layer=POLY_cond $X=1.22 $Y=1.22
+ $X2=1.31 $Y2=1.385
r36 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.22 $Y=1.22 $X2=1.22
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__NAND4_1%B 1 3 4 6 7
c31 7 0 3.78555e-20 $X=2.16 $Y=1.295
c32 1 0 1.64093e-19 $X=1.79 $Y=1.22
r33 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.88
+ $Y=1.385 $X2=1.88 $Y2=1.385
r34 7 11 8.72119 $w=3.68e-07 $l=2.8e-07 $layer=LI1_cond $X=2.16 $Y=1.365
+ $X2=1.88 $Y2=1.365
r35 4 10 77.2841 $w=2.7e-07 $l=3.82492e-07 $layer=POLY_cond $X=1.875 $Y=1.765
+ $X2=1.88 $Y2=1.385
r36 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.875 $Y=1.765
+ $X2=1.875 $Y2=2.4
r37 1 10 38.9026 $w=2.7e-07 $l=2.05122e-07 $layer=POLY_cond $X=1.79 $Y=1.22
+ $X2=1.88 $Y2=1.385
r38 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.79 $Y=1.22 $X2=1.79
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__NAND4_1%A 1 3 4 6 7
r21 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.61
+ $Y=1.385 $X2=2.61 $Y2=1.385
r22 7 11 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=2.61 $Y=1.295 $X2=2.61
+ $Y2=1.385
r23 4 10 67.2473 $w=3.67e-07 $l=4.50888e-07 $layer=POLY_cond $X=2.375 $Y=1.765
+ $X2=2.53 $Y2=1.385
r24 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.375 $Y=1.765
+ $X2=2.375 $Y2=2.4
r25 1 10 39.0103 $w=3.67e-07 $l=2.38642e-07 $layer=POLY_cond $X=2.36 $Y=1.22
+ $X2=2.53 $Y2=1.385
r26 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.36 $Y=1.22 $X2=2.36
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__NAND4_1%VPWR 1 2 3 12 18 20 22 27 28 30 31 32 41 47
c39 1 0 1.38338e-19 $X=0.395 $Y=1.84
r40 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r41 44 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r42 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r43 41 46 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=2.435 $Y=3.33
+ $X2=2.657 $Y2=3.33
r44 41 43 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.435 $Y=3.33
+ $X2=2.16 $Y2=3.33
r45 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r46 36 40 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r47 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r48 32 44 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=2.16 $Y2=3.33
r49 32 40 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.2 $Y2=3.33
r50 30 39 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=1.4 $Y=3.33 $X2=1.2
+ $Y2=3.33
r51 30 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.4 $Y=3.33
+ $X2=1.565 $Y2=3.33
r52 29 43 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=1.73 $Y=3.33
+ $X2=2.16 $Y2=3.33
r53 29 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.73 $Y=3.33
+ $X2=1.565 $Y2=3.33
r54 27 35 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=0.375 $Y=3.33
+ $X2=0.24 $Y2=3.33
r55 27 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.375 $Y=3.33
+ $X2=0.54 $Y2=3.33
r56 26 39 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=0.705 $Y=3.33
+ $X2=1.2 $Y2=3.33
r57 26 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.705 $Y=3.33
+ $X2=0.54 $Y2=3.33
r58 22 25 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=2.6 $Y=1.985 $X2=2.6
+ $Y2=2.815
r59 20 46 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=2.6 $Y=3.245
+ $X2=2.657 $Y2=3.33
r60 20 25 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.6 $Y=3.245 $X2=2.6
+ $Y2=2.815
r61 16 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.565 $Y=3.245
+ $X2=1.565 $Y2=3.33
r62 16 18 29.3349 $w=3.28e-07 $l=8.4e-07 $layer=LI1_cond $X=1.565 $Y=3.245
+ $X2=1.565 $Y2=2.405
r63 12 15 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.54 $Y=2.145
+ $X2=0.54 $Y2=2.825
r64 10 28 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.54 $Y=3.245
+ $X2=0.54 $Y2=3.33
r65 10 15 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=0.54 $Y=3.245
+ $X2=0.54 $Y2=2.825
r66 3 25 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.45
+ $Y=1.84 $X2=2.6 $Y2=2.815
r67 3 22 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.45
+ $Y=1.84 $X2=2.6 $Y2=1.985
r68 2 18 300 $w=1.7e-07 $l=6.68094e-07 $layer=licon1_PDIFF $count=2 $X=1.34
+ $Y=1.84 $X2=1.565 $Y2=2.405
r69 1 15 400 $w=1.7e-07 $l=1.05501e-06 $layer=licon1_PDIFF $count=1 $X=0.395
+ $Y=1.84 $X2=0.54 $Y2=2.825
r70 1 12 400 $w=1.7e-07 $l=3.70473e-07 $layer=licon1_PDIFF $count=1 $X=0.395
+ $Y=1.84 $X2=0.54 $Y2=2.145
.ends

.subckt PM_SKY130_FD_SC_LS__NAND4_1%Y 1 2 3 11 12 13 14 15 18 20 22 26 30 31 34
c73 15 0 1.38338e-19 $X=0.405 $Y=1.805
r74 31 34 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=1.935 $Y=1.985
+ $X2=1.68 $Y2=1.985
r75 31 33 3.40825 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=1.935 $Y=1.985
+ $X2=2.1 $Y2=1.985
r76 28 34 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=1.205 $Y=1.985
+ $X2=1.68 $Y2=1.985
r77 28 30 6.46576 $w=2.5e-07 $l=1.88348e-07 $layer=LI1_cond $X=1.205 $Y=1.985
+ $X2=1.04 $Y2=1.935
r78 24 26 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=2.575 $Y=0.84
+ $X2=2.575 $Y2=0.515
r79 20 33 3.40825 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=2.1 $Y=2.15 $X2=2.1
+ $Y2=1.985
r80 20 22 23.2235 $w=3.28e-07 $l=6.65e-07 $layer=LI1_cond $X=2.1 $Y=2.15 $X2=2.1
+ $Y2=2.815
r81 16 30 0.364692 $w=3.3e-07 $l=2.15e-07 $layer=LI1_cond $X=1.04 $Y=2.15
+ $X2=1.04 $Y2=1.935
r82 16 18 23.2235 $w=3.28e-07 $l=6.65e-07 $layer=LI1_cond $X=1.04 $Y=2.15
+ $X2=1.04 $Y2=2.815
r83 14 30 6.46576 $w=2.5e-07 $l=2.20624e-07 $layer=LI1_cond $X=0.875 $Y=1.805
+ $X2=1.04 $Y2=1.935
r84 14 15 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=0.875 $Y=1.805
+ $X2=0.405 $Y2=1.805
r85 12 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.41 $Y=0.925
+ $X2=2.575 $Y2=0.84
r86 12 13 130.807 $w=1.68e-07 $l=2.005e-06 $layer=LI1_cond $X=2.41 $Y=0.925
+ $X2=0.405 $Y2=0.925
r87 11 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.32 $Y=1.72
+ $X2=0.405 $Y2=1.805
r88 10 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.32 $Y=1.01
+ $X2=0.405 $Y2=0.925
r89 10 11 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=0.32 $Y=1.01
+ $X2=0.32 $Y2=1.72
r90 3 33 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.95
+ $Y=1.84 $X2=2.1 $Y2=1.985
r91 3 22 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.95
+ $Y=1.84 $X2=2.1 $Y2=2.815
r92 2 30 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=0.89
+ $Y=1.84 $X2=1.04 $Y2=1.985
r93 2 18 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=0.89
+ $Y=1.84 $X2=1.04 $Y2=2.815
r94 1 26 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.435
+ $Y=0.37 $X2=2.575 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__NAND4_1%VGND 1 4 8 9 12
r20 13 15 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r21 12 17 8.95014 $w=7.02e-07 $l=5.15e-07 $layer=LI1_cond $X=0.392 $Y=0
+ $X2=0.392 $Y2=0.515
r22 12 15 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r23 12 13 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r24 8 9 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r25 6 12 9.34032 $w=1.7e-07 $l=3.93e-07 $layer=LI1_cond $X=0.785 $Y=0 $X2=0.392
+ $Y2=0
r26 6 8 121.021 $w=1.68e-07 $l=1.855e-06 $layer=LI1_cond $X=0.785 $Y=0 $X2=2.64
+ $Y2=0
r27 4 9 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.44 $Y=0 $X2=2.64
+ $Y2=0
r28 4 15 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=0.72
+ $Y2=0
r29 1 17 91 $w=1.7e-07 $l=5.47723e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.615 $Y2=0.515
.ends

