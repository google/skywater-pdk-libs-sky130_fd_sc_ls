# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ls__dfsbp_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ls__dfsbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  12.00000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.475000 1.010000 0.805000 2.020000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.555000 0.350000 11.885000 1.050000 ;
        RECT 11.555000 1.820000 11.885000 2.980000 ;
        RECT 11.715000 1.050000 11.885000 1.820000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  9.985000 0.350000 10.315000 1.130000 ;
        RECT 10.120000 1.130000 10.315000 1.180000 ;
        RECT 10.120000 1.180000 10.435000 2.980000 ;
    END
  END Q_N
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.405000 1.550000 5.695000 1.955000 ;
        RECT 8.285000 1.180000 8.670000 1.780000 ;
      LAYER mcon ;
        RECT 5.435000 1.580000 5.605000 1.750000 ;
        RECT 8.315000 1.580000 8.485000 1.750000 ;
      LAYER met1 ;
        RECT 5.375000 1.550000 5.665000 1.595000 ;
        RECT 5.375000 1.595000 8.545000 1.735000 ;
        RECT 5.375000 1.735000 5.665000 1.780000 ;
        RECT 8.255000 1.550000 8.545000 1.595000 ;
        RECT 8.255000 1.735000 8.545000 1.780000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.315000 1.180000 1.795000 1.550000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 12.000000 0.085000 ;
        RECT  0.545000  0.085000  0.795000 0.840000 ;
        RECT  1.605000  0.085000  1.865000 1.010000 ;
        RECT  4.105000  0.085000  4.435000 0.715000 ;
        RECT  5.855000  0.085000  6.185000 0.950000 ;
        RECT  8.065000  0.085000  8.755000 0.670000 ;
        RECT  9.485000  0.085000  9.815000 0.670000 ;
        RECT 11.055000  0.085000 11.385000 0.940000 ;
      LAYER mcon ;
        RECT  0.155000 -0.085000  0.325000 0.085000 ;
        RECT  0.635000 -0.085000  0.805000 0.085000 ;
        RECT  1.115000 -0.085000  1.285000 0.085000 ;
        RECT  1.595000 -0.085000  1.765000 0.085000 ;
        RECT  2.075000 -0.085000  2.245000 0.085000 ;
        RECT  2.555000 -0.085000  2.725000 0.085000 ;
        RECT  3.035000 -0.085000  3.205000 0.085000 ;
        RECT  3.515000 -0.085000  3.685000 0.085000 ;
        RECT  3.995000 -0.085000  4.165000 0.085000 ;
        RECT  4.475000 -0.085000  4.645000 0.085000 ;
        RECT  4.955000 -0.085000  5.125000 0.085000 ;
        RECT  5.435000 -0.085000  5.605000 0.085000 ;
        RECT  5.915000 -0.085000  6.085000 0.085000 ;
        RECT  6.395000 -0.085000  6.565000 0.085000 ;
        RECT  6.875000 -0.085000  7.045000 0.085000 ;
        RECT  7.355000 -0.085000  7.525000 0.085000 ;
        RECT  7.835000 -0.085000  8.005000 0.085000 ;
        RECT  8.315000 -0.085000  8.485000 0.085000 ;
        RECT  8.795000 -0.085000  8.965000 0.085000 ;
        RECT  9.275000 -0.085000  9.445000 0.085000 ;
        RECT  9.755000 -0.085000  9.925000 0.085000 ;
        RECT 10.235000 -0.085000 10.405000 0.085000 ;
        RECT 10.715000 -0.085000 10.885000 0.085000 ;
        RECT 11.195000 -0.085000 11.365000 0.085000 ;
        RECT 11.675000 -0.085000 11.845000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 12.000000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 3.245000 12.000000 3.415000 ;
        RECT  0.565000 2.590000  0.895000 3.245000 ;
        RECT  1.575000 2.530000  1.905000 3.245000 ;
        RECT  4.045000 2.505000  4.440000 3.245000 ;
        RECT  5.710000 2.465000  6.050000 3.245000 ;
        RECT  8.070000 2.650000  8.240000 3.245000 ;
        RECT  9.560000 2.730000  9.910000 3.245000 ;
        RECT 11.050000 1.995000 11.380000 3.245000 ;
      LAYER mcon ;
        RECT  0.155000 3.245000  0.325000 3.415000 ;
        RECT  0.635000 3.245000  0.805000 3.415000 ;
        RECT  1.115000 3.245000  1.285000 3.415000 ;
        RECT  1.595000 3.245000  1.765000 3.415000 ;
        RECT  2.075000 3.245000  2.245000 3.415000 ;
        RECT  2.555000 3.245000  2.725000 3.415000 ;
        RECT  3.035000 3.245000  3.205000 3.415000 ;
        RECT  3.515000 3.245000  3.685000 3.415000 ;
        RECT  3.995000 3.245000  4.165000 3.415000 ;
        RECT  4.475000 3.245000  4.645000 3.415000 ;
        RECT  4.955000 3.245000  5.125000 3.415000 ;
        RECT  5.435000 3.245000  5.605000 3.415000 ;
        RECT  5.915000 3.245000  6.085000 3.415000 ;
        RECT  6.395000 3.245000  6.565000 3.415000 ;
        RECT  6.875000 3.245000  7.045000 3.415000 ;
        RECT  7.355000 3.245000  7.525000 3.415000 ;
        RECT  7.835000 3.245000  8.005000 3.415000 ;
        RECT  8.315000 3.245000  8.485000 3.415000 ;
        RECT  8.795000 3.245000  8.965000 3.415000 ;
        RECT  9.275000 3.245000  9.445000 3.415000 ;
        RECT  9.755000 3.245000  9.925000 3.415000 ;
        RECT 10.235000 3.245000 10.405000 3.415000 ;
        RECT 10.715000 3.245000 10.885000 3.415000 ;
        RECT 11.195000 3.245000 11.365000 3.415000 ;
        RECT 11.675000 3.245000 11.845000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 12.000000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.115000 0.380000  0.365000 0.840000 ;
      RECT  0.115000 0.840000  0.285000 2.190000 ;
      RECT  0.115000 2.190000  2.695000 2.230000 ;
      RECT  0.115000 2.230000  1.795000 2.360000 ;
      RECT  0.115000 2.360000  0.365000 2.980000 ;
      RECT  0.975000 0.350000  1.435000 1.010000 ;
      RECT  0.975000 1.010000  1.145000 1.720000 ;
      RECT  0.975000 1.720000  2.355000 1.890000 ;
      RECT  0.975000 1.890000  1.455000 2.020000 ;
      RECT  1.625000 2.060000  2.695000 2.190000 ;
      RECT  2.025000 1.300000  2.355000 1.720000 ;
      RECT  2.045000 0.255000  3.195000 0.425000 ;
      RECT  2.045000 0.425000  2.295000 1.130000 ;
      RECT  2.105000 2.400000  2.355000 2.905000 ;
      RECT  2.105000 2.905000  3.875000 3.075000 ;
      RECT  2.525000 0.595000  2.855000 0.845000 ;
      RECT  2.525000 0.845000  2.695000 2.060000 ;
      RECT  2.525000 2.230000  2.695000 2.295000 ;
      RECT  2.525000 2.295000  3.005000 2.735000 ;
      RECT  2.865000 1.435000  3.195000 2.105000 ;
      RECT  3.025000 0.425000  3.195000 1.435000 ;
      RECT  3.175000 2.295000  3.535000 2.735000 ;
      RECT  3.365000 0.385000  3.615000 0.885000 ;
      RECT  3.365000 0.885000  4.285000 1.055000 ;
      RECT  3.365000 1.055000  3.535000 2.295000 ;
      RECT  3.705000 1.360000  3.945000 2.165000 ;
      RECT  3.705000 2.165000  4.780000 2.335000 ;
      RECT  3.705000 2.335000  3.875000 2.905000 ;
      RECT  4.115000 1.055000  4.285000 1.435000 ;
      RECT  4.115000 1.435000  5.235000 1.605000 ;
      RECT  4.230000 1.775000  5.200000 1.995000 ;
      RECT  4.455000 0.885000  4.775000 1.265000 ;
      RECT  4.605000 0.435000  5.180000 0.885000 ;
      RECT  4.610000 2.335000  4.780000 2.905000 ;
      RECT  4.610000 2.905000  5.540000 3.075000 ;
      RECT  4.950000 1.055000  5.235000 1.120000 ;
      RECT  4.950000 1.120000  6.265000 1.290000 ;
      RECT  4.950000 1.290000  5.235000 1.435000 ;
      RECT  4.950000 1.995000  5.200000 2.735000 ;
      RECT  5.370000 2.125000  6.035000 2.295000 ;
      RECT  5.370000 2.295000  5.540000 2.905000 ;
      RECT  5.865000 1.620000  6.605000 1.790000 ;
      RECT  5.865000 1.790000  6.035000 2.125000 ;
      RECT  5.935000 1.290000  6.265000 1.450000 ;
      RECT  6.435000 0.255000  7.560000 0.425000 ;
      RECT  6.435000 0.425000  6.605000 1.120000 ;
      RECT  6.435000 1.120000  6.880000 1.450000 ;
      RECT  6.435000 1.450000  6.605000 1.620000 ;
      RECT  6.760000 1.960000  7.010000 2.480000 ;
      RECT  6.760000 2.480000  7.900000 2.650000 ;
      RECT  6.760000 2.650000  7.450000 2.905000 ;
      RECT  6.775000 0.595000  7.220000 0.925000 ;
      RECT  6.840000 1.680000  7.220000 1.850000 ;
      RECT  6.840000 1.850000  7.010000 1.960000 ;
      RECT  7.050000 0.925000  7.220000 1.680000 ;
      RECT  7.230000 2.020000  7.560000 2.310000 ;
      RECT  7.390000 0.425000  7.560000 2.020000 ;
      RECT  7.730000 2.050000  9.395000 2.220000 ;
      RECT  7.730000 2.220000  8.770000 2.480000 ;
      RECT  7.770000 0.840000  9.735000 1.010000 ;
      RECT  7.770000 1.010000  8.100000 1.880000 ;
      RECT  8.440000 2.480000  8.770000 2.980000 ;
      RECT  8.925000 0.415000  9.255000 0.840000 ;
      RECT  9.000000 2.390000  9.735000 2.560000 ;
      RECT  9.000000 2.560000  9.330000 2.980000 ;
      RECT  9.065000 1.210000  9.395000 2.050000 ;
      RECT  9.565000 1.010000  9.735000 2.390000 ;
      RECT 10.545000 0.350000 10.875000 0.940000 ;
      RECT 10.680000 0.940000 10.875000 1.220000 ;
      RECT 10.680000 1.220000 11.540000 1.550000 ;
      RECT 10.680000 1.550000 10.850000 2.875000 ;
  END
END sky130_fd_sc_ls__dfsbp_1
