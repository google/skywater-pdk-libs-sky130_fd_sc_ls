* File: sky130_fd_sc_ls__a31o_1.pex.spice
* Created: Fri Aug 28 12:58:36 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__A31O_1%A_81_270# 1 2 7 9 10 12 13 17 19 23 27 31
r73 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.59
+ $Y=1.515 $X2=0.59 $Y2=1.515
r74 27 29 10.4785 $w=3.26e-07 $l=2.8e-07 $layer=LI1_cond $X=0.625 $Y=1.235
+ $X2=0.625 $Y2=1.515
r75 23 25 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=2.97 $Y=2.105
+ $X2=2.97 $Y2=2.815
r76 21 23 36.1867 $w=2.48e-07 $l=7.85e-07 $layer=LI1_cond $X=2.97 $Y=1.32
+ $X2=2.97 $Y2=2.105
r77 20 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.61 $Y=1.235
+ $X2=2.445 $Y2=1.235
r78 19 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.845 $Y=1.235
+ $X2=2.97 $Y2=1.32
r79 19 20 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=2.845 $Y=1.235
+ $X2=2.61 $Y2=1.235
r80 15 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.445 $Y=1.15
+ $X2=2.445 $Y2=1.235
r81 15 17 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=2.445 $Y=1.15
+ $X2=2.445 $Y2=0.955
r82 14 27 4.55145 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=0.825 $Y=1.235
+ $X2=0.625 $Y2=1.235
r83 13 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.28 $Y=1.235
+ $X2=2.445 $Y2=1.235
r84 13 14 94.9251 $w=1.68e-07 $l=1.455e-06 $layer=LI1_cond $X=2.28 $Y=1.235
+ $X2=0.825 $Y2=1.235
r85 10 30 38.5363 $w=3.15e-07 $l=1.96914e-07 $layer=POLY_cond $X=0.51 $Y=1.35
+ $X2=0.58 $Y2=1.515
r86 10 12 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.51 $Y=1.35 $X2=0.51
+ $Y2=0.87
r87 7 30 51.5426 $w=3.15e-07 $l=2.89396e-07 $layer=POLY_cond $X=0.495 $Y=1.765
+ $X2=0.58 $Y2=1.515
r88 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.495 $Y=1.765
+ $X2=0.495 $Y2=2.4
r89 2 25 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=2.78
+ $Y=1.96 $X2=2.93 $Y2=2.815
r90 2 23 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.78
+ $Y=1.96 $X2=2.93 $Y2=2.105
r91 1 17 182 $w=1.7e-07 $l=4.36348e-07 $layer=licon1_NDIFF $count=1 $X=2.225
+ $Y=0.615 $X2=2.445 $Y2=0.955
.ends

.subckt PM_SKY130_FD_SC_LS__A31O_1%A3 1 3 6 8
r32 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.16
+ $Y=1.635 $X2=1.16 $Y2=1.635
r33 4 11 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=1.25 $Y=1.47
+ $X2=1.16 $Y2=1.635
r34 4 6 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.25 $Y=1.47 $X2=1.25
+ $Y2=0.92
r35 1 11 52.2586 $w=2.99e-07 $l=2.57391e-07 $layer=POLY_cond $X=1.175 $Y=1.885
+ $X2=1.16 $Y2=1.635
r36 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.175 $Y=1.885
+ $X2=1.175 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_LS__A31O_1%A2 3 5 7 8
r30 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.7
+ $Y=1.635 $X2=1.7 $Y2=1.635
r31 5 11 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=1.625 $Y=1.885
+ $X2=1.7 $Y2=1.635
r32 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.625 $Y=1.885
+ $X2=1.625 $Y2=2.46
r33 1 11 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=1.61 $Y=1.47
+ $X2=1.7 $Y2=1.635
r34 1 3 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.61 $Y=1.47 $X2=1.61
+ $Y2=0.92
.ends

.subckt PM_SKY130_FD_SC_LS__A31O_1%A1 3 5 7 8
r33 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.24
+ $Y=1.635 $X2=2.24 $Y2=1.635
r34 5 11 52.2586 $w=2.99e-07 $l=2.57391e-07 $layer=POLY_cond $X=2.255 $Y=1.885
+ $X2=2.24 $Y2=1.635
r35 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.255 $Y=1.885
+ $X2=2.255 $Y2=2.46
r36 1 11 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=2.15 $Y=1.47
+ $X2=2.24 $Y2=1.635
r37 1 3 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=2.15 $Y=1.47 $X2=2.15
+ $Y2=0.935
.ends

.subckt PM_SKY130_FD_SC_LS__A31O_1%B1 2 3 5 9 11 12 13 14 19 20
r41 19 22 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.65 $Y=0.34
+ $X2=2.65 $Y2=0.505
r42 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.65
+ $Y=0.34 $X2=2.65 $Y2=0.34
r43 14 20 0.299336 $w=3.83e-07 $l=1e-08 $layer=LI1_cond $X=2.64 $Y=0.447
+ $X2=2.65 $Y2=0.447
r44 13 14 14.3681 $w=3.83e-07 $l=4.8e-07 $layer=LI1_cond $X=2.16 $Y=0.447
+ $X2=2.64 $Y2=0.447
r45 12 13 14.3681 $w=3.83e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=0.447
+ $X2=2.16 $Y2=0.447
r46 10 11 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=2.715 $Y=1.435
+ $X2=2.715 $Y2=1.585
r47 9 10 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=2.74 $Y=0.935 $X2=2.74
+ $Y2=1.435
r48 9 22 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.74 $Y=0.935
+ $X2=2.74 $Y2=0.505
r49 3 5 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.705 $Y=1.885
+ $X2=2.705 $Y2=2.46
r50 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.705 $Y=1.795 $X2=2.705
+ $Y2=1.885
r51 2 11 81.629 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=2.705 $Y=1.795
+ $X2=2.705 $Y2=1.585
.ends

.subckt PM_SKY130_FD_SC_LS__A31O_1%X 1 2 9 13 14 15 16 23 32
r22 21 23 0.329269 $w=3.48e-07 $l=1e-08 $layer=LI1_cond $X=0.26 $Y=2.025
+ $X2=0.26 $Y2=2.035
r23 15 16 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.26 $Y=2.405
+ $X2=0.26 $Y2=2.775
r24 14 21 1.25122 $w=3.48e-07 $l=3.8e-08 $layer=LI1_cond $X=0.26 $Y=1.987
+ $X2=0.26 $Y2=2.025
r25 14 32 7.56653 $w=3.48e-07 $l=1.37e-07 $layer=LI1_cond $X=0.26 $Y=1.987
+ $X2=0.26 $Y2=1.85
r26 14 15 10.9647 $w=3.48e-07 $l=3.33e-07 $layer=LI1_cond $X=0.26 $Y=2.072
+ $X2=0.26 $Y2=2.405
r27 14 23 1.2183 $w=3.48e-07 $l=3.7e-08 $layer=LI1_cond $X=0.26 $Y=2.072
+ $X2=0.26 $Y2=2.035
r28 13 32 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.17 $Y=1.18
+ $X2=0.17 $Y2=1.85
r29 7 13 9.06106 $w=3.63e-07 $l=1.82e-07 $layer=LI1_cond $X=0.267 $Y=0.998
+ $X2=0.267 $Y2=1.18
r30 7 9 11.1455 $w=3.63e-07 $l=3.53e-07 $layer=LI1_cond $X=0.267 $Y=0.998
+ $X2=0.267 $Y2=0.645
r31 2 14 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.84 $X2=0.27 $Y2=2.015
r32 2 16 400 $w=1.7e-07 $l=1.03562e-06 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.84 $X2=0.27 $Y2=2.815
r33 1 9 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.17 $Y=0.5
+ $X2=0.295 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_LS__A31O_1%VPWR 1 2 9 15 18 19 20 22 35 36 39
r40 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r41 35 36 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r42 33 36 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r43 32 35 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=3.33 $X2=3.12
+ $Y2=3.33
r44 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r45 27 39 10.7288 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=1.065 $Y=3.33
+ $X2=0.835 $Y2=3.33
r46 27 29 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=1.065 $Y=3.33
+ $X2=1.68 $Y2=3.33
r47 25 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r48 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r49 22 39 10.7288 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=0.605 $Y=3.33
+ $X2=0.835 $Y2=3.33
r50 22 24 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.605 $Y=3.33
+ $X2=0.24 $Y2=3.33
r51 20 33 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r52 20 40 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r53 20 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r54 18 29 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=1.735 $Y=3.33
+ $X2=1.68 $Y2=3.33
r55 18 19 9.97069 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=1.735 $Y=3.33
+ $X2=1.94 $Y2=3.33
r56 17 32 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=2.145 $Y=3.33
+ $X2=2.16 $Y2=3.33
r57 17 19 9.97069 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=2.145 $Y=3.33
+ $X2=1.94 $Y2=3.33
r58 13 19 1.53834 $w=4.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.94 $Y=3.245
+ $X2=1.94 $Y2=3.33
r59 13 15 23.1894 $w=4.08e-07 $l=8.25e-07 $layer=LI1_cond $X=1.94 $Y=3.245
+ $X2=1.94 $Y2=2.42
r60 9 12 17.6812 $w=4.58e-07 $l=6.8e-07 $layer=LI1_cond $X=0.835 $Y=2.135
+ $X2=0.835 $Y2=2.815
r61 7 39 1.85547 $w=4.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.835 $Y=3.245
+ $X2=0.835 $Y2=3.33
r62 7 12 11.1807 $w=4.58e-07 $l=4.3e-07 $layer=LI1_cond $X=0.835 $Y=3.245
+ $X2=0.835 $Y2=2.815
r63 2 15 300 $w=1.7e-07 $l=5.6745e-07 $layer=licon1_PDIFF $count=2 $X=1.7
+ $Y=1.96 $X2=1.94 $Y2=2.42
r64 1 12 400 $w=1.7e-07 $l=1.09955e-06 $layer=licon1_PDIFF $count=1 $X=0.57
+ $Y=1.84 $X2=0.835 $Y2=2.815
r65 1 9 400 $w=1.7e-07 $l=4.06448e-07 $layer=licon1_PDIFF $count=1 $X=0.57
+ $Y=1.84 $X2=0.835 $Y2=2.135
.ends

.subckt PM_SKY130_FD_SC_LS__A31O_1%A_250_392# 1 2 7 9 11 13 15
r34 13 20 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.48 $Y=2.14 $X2=2.48
+ $Y2=2.055
r35 13 15 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.48 $Y=2.14
+ $X2=2.48 $Y2=2.815
r36 12 18 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.565 $Y=2.055
+ $X2=1.4 $Y2=2.055
r37 11 20 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.315 $Y=2.055
+ $X2=2.48 $Y2=2.055
r38 11 12 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=2.315 $Y=2.055
+ $X2=1.565 $Y2=2.055
r39 7 18 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.4 $Y=2.14 $X2=1.4
+ $Y2=2.055
r40 7 9 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=1.4 $Y=2.14 $X2=1.4
+ $Y2=2.815
r41 2 20 400 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=1 $X=2.33
+ $Y=1.96 $X2=2.48 $Y2=2.135
r42 2 15 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=2.33
+ $Y=1.96 $X2=2.48 $Y2=2.815
r43 1 18 400 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=1 $X=1.25
+ $Y=1.96 $X2=1.4 $Y2=2.135
r44 1 9 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=1.25
+ $Y=1.96 $X2=1.4 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_LS__A31O_1%VGND 1 2 9 11 12 16 18 20 25 34 38
r38 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r39 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r40 32 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r41 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r42 29 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r43 28 34 12.3201 $w=1.7e-07 $l=2.9e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=0.91
+ $Y2=0
r44 28 31 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r45 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r46 25 37 3.40825 $w=1.7e-07 $l=1.87e-07 $layer=LI1_cond $X=2.985 $Y=0 $X2=3.172
+ $Y2=0
r47 25 31 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.985 $Y=0 $X2=2.64
+ $Y2=0
r48 23 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r49 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r50 20 34 12.3201 $w=1.7e-07 $l=2.9e-07 $layer=LI1_cond $X=0.62 $Y=0 $X2=0.91
+ $Y2=0
r51 20 22 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=0.62 $Y=0 $X2=0.24
+ $Y2=0
r52 18 32 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r53 18 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r54 14 16 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=2.955 $Y=0.895
+ $X2=3.07 $Y2=0.895
r55 12 16 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.07 $Y=0.81
+ $X2=3.07 $Y2=0.895
r56 11 37 3.40825 $w=1.7e-07 $l=1.38109e-07 $layer=LI1_cond $X=3.07 $Y=0.085
+ $X2=3.172 $Y2=0
r57 11 12 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=3.07 $Y=0.085
+ $X2=3.07 $Y2=0.81
r58 7 34 2.44113 $w=5.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.91 $Y=0.085 $X2=0.91
+ $Y2=0
r59 7 9 11.1359 $w=5.78e-07 $l=5.4e-07 $layer=LI1_cond $X=0.91 $Y=0.085 $X2=0.91
+ $Y2=0.625
r60 2 14 182 $w=1.7e-07 $l=3.42929e-07 $layer=licon1_NDIFF $count=1 $X=2.815
+ $Y=0.615 $X2=2.955 $Y2=0.895
r61 1 9 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=0.585
+ $Y=0.5 $X2=0.725 $Y2=0.625
.ends

