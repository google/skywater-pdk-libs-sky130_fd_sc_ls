* File: sky130_fd_sc_ls__dfrbp_1.pex.spice
* Created: Fri Aug 28 13:13:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__DFRBP_1%D 1 3 6 8 9 10 11 17 20 21
r34 20 22 45.79 $w=4.05e-07 $l=1.65e-07 $layer=POLY_cond $X=0.422 $Y=1.165
+ $X2=0.422 $Y2=1
r35 20 21 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.165 $X2=0.385 $Y2=1.165
r36 17 18 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.845 $X2=0.385 $Y2=1.845
r37 15 20 5.08091 $w=4.05e-07 $l=3.7e-08 $layer=POLY_cond $X=0.422 $Y=1.202
+ $X2=0.422 $Y2=1.165
r38 15 17 88.298 $w=4.05e-07 $l=6.43e-07 $layer=POLY_cond $X=0.422 $Y=1.202
+ $X2=0.422 $Y2=1.845
r39 11 18 5.5434 $w=3.93e-07 $l=1.9e-07 $layer=LI1_cond $X=0.322 $Y=2.035
+ $X2=0.322 $Y2=1.845
r40 10 18 5.25164 $w=3.93e-07 $l=1.8e-07 $layer=LI1_cond $X=0.322 $Y=1.665
+ $X2=0.322 $Y2=1.845
r41 9 10 10.795 $w=3.93e-07 $l=3.7e-07 $layer=LI1_cond $X=0.322 $Y=1.295
+ $X2=0.322 $Y2=1.665
r42 9 21 3.79285 $w=3.93e-07 $l=1.3e-07 $layer=LI1_cond $X=0.322 $Y=1.295
+ $X2=0.322 $Y2=1.165
r43 8 17 41.6085 $w=4.05e-07 $l=3.03e-07 $layer=POLY_cond $X=0.422 $Y=2.148
+ $X2=0.422 $Y2=1.845
r44 6 22 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=0.55 $Y=0.6 $X2=0.55
+ $Y2=1
r45 1 8 47.3046 $w=3.23e-07 $l=3.5609e-07 $layer=POLY_cond $X=0.505 $Y=2.465
+ $X2=0.422 $Y2=2.148
r46 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.505 $Y=2.465
+ $X2=0.505 $Y2=2.75
.ends

.subckt PM_SKY130_FD_SC_LS__DFRBP_1%CLK 3 7 8 11 13
c48 13 0 3.22254e-19 $X=1.962 $Y=1.41
r49 11 14 46.504 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=1.962 $Y=1.61
+ $X2=1.962 $Y2=1.775
r50 11 13 52.1932 $w=3.55e-07 $l=2e-07 $layer=POLY_cond $X=1.962 $Y=1.61
+ $X2=1.962 $Y2=1.41
r51 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.975
+ $Y=1.61 $X2=1.975 $Y2=1.61
r52 8 12 5.28571 $w=4.27e-07 $l=1.85e-07 $layer=LI1_cond $X=2.16 $Y=1.545
+ $X2=1.975 $Y2=1.545
r53 7 13 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.97 $Y=0.965
+ $X2=1.97 $Y2=1.41
r54 3 14 351.245 $w=1.5e-07 $l=6.85e-07 $layer=POLY_cond $X=1.965 $Y=2.46
+ $X2=1.965 $Y2=1.775
.ends

.subckt PM_SKY130_FD_SC_LS__DFRBP_1%A_500_392# 1 2 7 8 11 12 15 18 19 21 22 23
+ 24 26 27 28 29 30 37 38 41 42 43 45 46 47 50 52 53 55 58 64 67 68
c205 68 0 1.81428e-19 $X=3.052 $Y=1.39
c206 58 0 9.20497e-20 $X=2.862 $Y=0.34
c207 52 0 1.08581e-19 $X=6.735 $Y=1.865
c208 47 0 1.02732e-19 $X=6.255 $Y=1.065
c209 43 0 1.61434e-19 $X=4.52 $Y=0.665
c210 37 0 1.94586e-20 $X=3.067 $Y=1.575
c211 28 0 3.00656e-19 $X=4.05 $Y=1.09
c212 7 0 2.61274e-19 $X=3.462 $Y=1.985
r213 67 68 11.1834 $w=1.83e-07 $l=1.85e-07 $layer=LI1_cond $X=3.052 $Y=1.205
+ $X2=3.052 $Y2=1.39
r214 65 69 29.2361 $w=3.05e-07 $l=1.85e-07 $layer=POLY_cond $X=3.385 $Y=1.82
+ $X2=3.385 $Y2=1.635
r215 64 65 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.385
+ $Y=1.82 $X2=3.385 $Y2=1.82
r216 62 67 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=3.03 $Y=0.805
+ $X2=3.03 $Y2=1.205
r217 61 62 7.65311 $w=5.03e-07 $l=8.5e-08 $layer=LI1_cond $X=2.862 $Y=0.72
+ $X2=2.862 $Y2=0.805
r218 58 61 9.00019 $w=5.03e-07 $l=3.8e-07 $layer=LI1_cond $X=2.862 $Y=0.34
+ $X2=2.862 $Y2=0.72
r219 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.205
+ $Y=2.03 $X2=7.205 $Y2=2.03
r220 53 55 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=6.82 $Y=2.03
+ $X2=7.205 $Y2=2.03
r221 52 53 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.735 $Y=1.865
+ $X2=6.82 $Y2=2.03
r222 51 52 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=6.735 $Y=1.23
+ $X2=6.735 $Y2=1.865
r223 50 73 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=6.645 $Y=1.065
+ $X2=6.645 $Y2=1.16
r224 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.645
+ $Y=1.065 $X2=6.645 $Y2=1.065
r225 47 49 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=6.255 $Y=1.065
+ $X2=6.645 $Y2=1.065
r226 46 51 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.65 $Y=1.065
+ $X2=6.735 $Y2=1.23
r227 46 49 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=6.65 $Y=1.065
+ $X2=6.645 $Y2=1.065
r228 45 47 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.17 $Y=0.9
+ $X2=6.255 $Y2=1.065
r229 44 45 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=6.17 $Y=0.75
+ $X2=6.17 $Y2=0.9
r230 42 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.085 $Y=0.665
+ $X2=6.17 $Y2=0.75
r231 42 43 102.102 $w=1.68e-07 $l=1.565e-06 $layer=LI1_cond $X=6.085 $Y=0.665
+ $X2=4.52 $Y2=0.665
r232 41 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.435 $Y=0.58
+ $X2=4.52 $Y2=0.665
r233 40 41 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=4.435 $Y=0.425
+ $X2=4.435 $Y2=0.58
r234 39 58 7.21919 $w=1.7e-07 $l=2.53e-07 $layer=LI1_cond $X=3.115 $Y=0.34
+ $X2=2.862 $Y2=0.34
r235 38 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.35 $Y=0.34
+ $X2=4.435 $Y2=0.425
r236 38 39 80.5722 $w=1.68e-07 $l=1.235e-06 $layer=LI1_cond $X=4.35 $Y=0.34
+ $X2=3.115 $Y2=0.34
r237 37 64 11.05 $w=3.91e-07 $l=3.07124e-07 $layer=LI1_cond $X=3.067 $Y=1.575
+ $X2=3.207 $Y2=1.82
r238 37 68 11.0909 $w=1.83e-07 $l=1.85e-07 $layer=LI1_cond $X=3.067 $Y=1.575
+ $X2=3.067 $Y2=1.39
r239 30 64 7.23887 $w=3.91e-07 $l=3.91162e-07 $layer=LI1_cond $X=2.915 $Y=2.052
+ $X2=3.207 $Y2=1.82
r240 30 32 8.45125 $w=3.73e-07 $l=2.75e-07 $layer=LI1_cond $X=2.915 $Y=2.052
+ $X2=2.64 $Y2=2.052
r241 28 29 43.7534 $w=2.2e-07 $l=1.5e-07 $layer=POLY_cond $X=4.05 $Y=1.09
+ $X2=4.05 $Y2=1.24
r242 24 56 52.2586 $w=2.99e-07 $l=2.7157e-07 $layer=POLY_cond $X=7.25 $Y=2.28
+ $X2=7.205 $Y2=2.03
r243 24 26 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.25 $Y=2.28
+ $X2=7.25 $Y2=2.565
r244 22 73 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.48 $Y=1.16
+ $X2=6.645 $Y2=1.16
r245 22 23 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=6.48 $Y=1.16
+ $X2=6.12 $Y2=1.16
r246 19 23 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.045 $Y=1.085
+ $X2=6.12 $Y2=1.16
r247 19 21 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=6.045 $Y=1.085
+ $X2=6.045 $Y2=0.69
r248 18 28 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.085 $Y=0.805
+ $X2=4.085 $Y2=1.09
r249 15 29 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.015 $Y=1.56
+ $X2=4.015 $Y2=1.24
r250 13 69 19.3576 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.55 $Y=1.635
+ $X2=3.385 $Y2=1.635
r251 12 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.94 $Y=1.635
+ $X2=4.015 $Y2=1.56
r252 12 13 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=3.94 $Y=1.635
+ $X2=3.55 $Y2=1.635
r253 11 27 101.22 $w=1.5e-07 $l=3.15e-07 $layer=POLY_cond $X=3.45 $Y=2.525
+ $X2=3.45 $Y2=2.21
r254 8 27 36.4084 $w=1.75e-07 $l=8.7e-08 $layer=POLY_cond $X=3.462 $Y=2.123
+ $X2=3.462 $Y2=2.21
r255 7 65 34.7586 $w=3.05e-07 $l=1.99825e-07 $layer=POLY_cond $X=3.462 $Y=1.985
+ $X2=3.385 $Y2=1.82
r256 7 8 55.1746 $w=1.75e-07 $l=1.38e-07 $layer=POLY_cond $X=3.462 $Y=1.985
+ $X2=3.462 $Y2=2.123
r257 2 32 600 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_PDIFF $count=1 $X=2.5
+ $Y=1.96 $X2=2.64 $Y2=2.155
r258 1 61 182 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_NDIFF $count=1 $X=2.625
+ $Y=0.595 $X2=2.775 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_LS__DFRBP_1%A_841_401# 1 2 7 9 12 14 19 20 22 23 24 25
+ 26 27 30
c111 23 0 5.58686e-20 $X=4.63 $Y=1.005
c112 12 0 3.41044e-19 $X=4.475 $Y=0.805
c113 7 0 2.19701e-19 $X=4.295 $Y=2.24
r114 30 32 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=6.355 $Y=1.88
+ $X2=6.355 $Y2=2.59
r115 28 30 14.2903 $w=2.48e-07 $l=3.1e-07 $layer=LI1_cond $X=6.355 $Y=1.57
+ $X2=6.355 $Y2=1.88
r116 26 28 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.23 $Y=1.485
+ $X2=6.355 $Y2=1.57
r117 26 27 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=6.23 $Y=1.485
+ $X2=5.915 $Y2=1.485
r118 25 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.83 $Y=1.4
+ $X2=5.915 $Y2=1.485
r119 24 35 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.83 $Y=1.09
+ $X2=5.83 $Y2=1.005
r120 24 25 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=5.83 $Y=1.09
+ $X2=5.83 $Y2=1.4
r121 22 35 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.745 $Y=1.005
+ $X2=5.83 $Y2=1.005
r122 22 23 72.7433 $w=1.68e-07 $l=1.115e-06 $layer=LI1_cond $X=5.745 $Y=1.005
+ $X2=4.63 $Y2=1.005
r123 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.465
+ $Y=1.65 $X2=4.465 $Y2=1.65
r124 17 23 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=4.49 $Y=1.09
+ $X2=4.63 $Y2=1.005
r125 17 19 23.0489 $w=2.78e-07 $l=5.6e-07 $layer=LI1_cond $X=4.49 $Y=1.09
+ $X2=4.49 $Y2=1.65
r126 16 20 38.0424 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.465 $Y=1.485
+ $X2=4.465 $Y2=1.65
r127 14 20 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=4.465 $Y=2.005
+ $X2=4.465 $Y2=1.65
r128 12 16 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=4.475 $Y=0.805
+ $X2=4.475 $Y2=1.485
r129 7 14 33.7113 $w=3.36e-07 $l=3.08504e-07 $layer=POLY_cond $X=4.295 $Y=2.24
+ $X2=4.465 $Y2=2.005
r130 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.295 $Y=2.24
+ $X2=4.295 $Y2=2.525
r131 2 32 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=6.165
+ $Y=1.735 $X2=6.315 $Y2=2.59
r132 2 30 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=6.165
+ $Y=1.735 $X2=6.315 $Y2=1.88
r133 1 35 182 $w=1.7e-07 $l=7.36834e-07 $layer=licon1_NDIFF $count=1 $X=5.53
+ $Y=0.37 $X2=5.75 $Y2=1.005
.ends

.subckt PM_SKY130_FD_SC_LS__DFRBP_1%RESET_B 4 6 8 9 11 12 13 17 19 20 22 25 27
+ 29 31 33 34 35 36 37 42 45 48 49 52 53 56 61
c212 53 0 4.15557e-20 $X=1.165 $Y=1.295
c213 52 0 1.03964e-19 $X=1.165 $Y=1.295
c214 42 0 6.85463e-20 $X=7.92 $Y=2.035
c215 34 0 1.81428e-19 $X=5.375 $Y=2.035
c216 12 0 4.00428e-20 $X=4.79 $Y=0.18
r217 60 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.135
+ $Y=2 $X2=8.135 $Y2=2
r218 56 58 41.4566 $w=4.65e-07 $l=1.65e-07 $layer=POLY_cond $X=1.097 $Y=1.975
+ $X2=1.097 $Y2=2.14
r219 56 57 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.165
+ $Y=1.975 $X2=1.165 $Y2=1.975
r220 53 57 29.0245 $w=2.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.165 $Y=1.295
+ $X2=1.165 $Y2=1.975
r221 52 54 47.3569 $w=4.65e-07 $l=1.65e-07 $layer=POLY_cond $X=1.097 $Y=1.295
+ $X2=1.097 $Y2=1.13
r222 52 53 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.165
+ $Y=1.295 $X2=1.165 $Y2=1.295
r223 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.395
+ $Y=1.99 $X2=5.395 $Y2=1.99
r224 45 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=2.035
+ $X2=1.2 $Y2=2.035
r225 43 61 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=7.92 $Y=2
+ $X2=8.135 $Y2=2
r226 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=2.035
+ $X2=7.92 $Y2=2.035
r227 39 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=2.035
+ $X2=5.52 $Y2=2.035
r228 37 39 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.665 $Y=2.035
+ $X2=5.52 $Y2=2.035
r229 36 42 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.775 $Y=2.035
+ $X2=7.92 $Y2=2.035
r230 36 37 2.61138 $w=1.4e-07 $l=2.11e-06 $layer=MET1_cond $X=7.775 $Y=2.035
+ $X2=5.665 $Y2=2.035
r231 35 45 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.345 $Y=2.035
+ $X2=1.2 $Y2=2.035
r232 34 39 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.375 $Y=2.035
+ $X2=5.52 $Y2=2.035
r233 34 35 4.98761 $w=1.4e-07 $l=4.03e-06 $layer=MET1_cond $X=5.375 $Y=2.035
+ $X2=1.345 $Y2=2.035
r234 32 48 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=5.02 $Y=1.99
+ $X2=5.395 $Y2=1.99
r235 32 33 5.03009 $w=3.3e-07 $l=1.08995e-07 $layer=POLY_cond $X=5.02 $Y=1.99
+ $X2=4.93 $Y2=2.032
r236 30 31 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=4.89 $Y=1.09 $X2=4.89
+ $Y2=1.24
r237 27 60 57.6553 $w=2.91e-07 $l=3.01662e-07 $layer=POLY_cond $X=8.18 $Y=2.28
+ $X2=8.135 $Y2=2
r238 27 29 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=8.18 $Y=2.28
+ $X2=8.18 $Y2=2.565
r239 23 60 38.6072 $w=2.91e-07 $l=2.05122e-07 $layer=POLY_cond $X=8.045 $Y=1.835
+ $X2=8.135 $Y2=2
r240 23 25 643.521 $w=1.5e-07 $l=1.255e-06 $layer=POLY_cond $X=8.045 $Y=1.835
+ $X2=8.045 $Y2=0.58
r241 20 33 37.0704 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=4.93 $Y=2.24
+ $X2=4.93 $Y2=2.032
r242 20 22 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.93 $Y=2.24
+ $X2=4.93 $Y2=2.525
r243 19 33 37.0704 $w=1.5e-07 $l=2.14369e-07 $layer=POLY_cond $X=4.915 $Y=1.825
+ $X2=4.93 $Y2=2.032
r244 19 31 299.968 $w=1.5e-07 $l=5.85e-07 $layer=POLY_cond $X=4.915 $Y=1.825
+ $X2=4.915 $Y2=1.24
r245 17 30 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.865 $Y=0.805
+ $X2=4.865 $Y2=1.09
r246 14 17 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=4.865 $Y=0.255
+ $X2=4.865 $Y2=0.805
r247 12 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.79 $Y=0.18
+ $X2=4.865 $Y2=0.255
r248 12 13 1935.69 $w=1.5e-07 $l=3.775e-06 $layer=POLY_cond $X=4.79 $Y=0.18
+ $X2=1.015 $Y2=0.18
r249 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.955 $Y=2.465
+ $X2=0.955 $Y2=2.75
r250 8 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.955 $Y=2.375
+ $X2=0.955 $Y2=2.465
r251 8 58 91.3468 $w=1.8e-07 $l=2.35e-07 $layer=POLY_cond $X=0.955 $Y=2.375
+ $X2=0.955 $Y2=2.14
r252 6 56 8.0134 $w=4.65e-07 $l=6.7e-08 $layer=POLY_cond $X=1.097 $Y=1.908
+ $X2=1.097 $Y2=1.975
r253 5 52 8.0134 $w=4.65e-07 $l=6.7e-08 $layer=POLY_cond $X=1.097 $Y=1.362
+ $X2=1.097 $Y2=1.295
r254 5 6 65.3032 $w=4.65e-07 $l=5.46e-07 $layer=POLY_cond $X=1.097 $Y=1.362
+ $X2=1.097 $Y2=1.908
r255 4 54 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.94 $Y=0.6 $X2=0.94
+ $Y2=1.13
r256 1 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.94 $Y=0.255
+ $X2=1.015 $Y2=0.18
r257 1 4 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=0.94 $Y=0.255
+ $X2=0.94 $Y2=0.6
.ends

.subckt PM_SKY130_FD_SC_LS__DFRBP_1%A_705_463# 1 2 3 12 14 16 18 19 25 28 32 34
+ 35 38 41 42
c128 38 0 1.55214e-19 $X=4.975 $Y=1.45
c129 35 0 1.25323e-19 $X=4.14 $Y=2.325
c130 32 0 1.09016e-19 $X=4.095 $Y=0.812
c131 28 0 1.98111e-19 $X=4.975 $Y=2.28
c132 19 0 7.95804e-20 $X=4.01 $Y=2.61
c133 14 0 2.11313e-19 $X=6 $Y=1.54
r134 42 44 6.65782 $w=3.39e-07 $l=1.85e-07 $layer=LI1_cond $X=4.975 $Y=2.48
+ $X2=5.16 $Y2=2.48
r135 41 47 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.395 $Y=1.45
+ $X2=5.395 $Y2=1.54
r136 41 46 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.395 $Y=1.45
+ $X2=5.395 $Y2=1.285
r137 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.395
+ $Y=1.45 $X2=5.395 $Y2=1.45
r138 38 40 20.6613 $w=2.48e-07 $l=4.2e-07 $layer=LI1_cond $X=4.975 $Y=1.45
+ $X2=5.395 $Y2=1.45
r139 34 36 8.86495 $w=2.58e-07 $l=2e-07 $layer=LI1_cond $X=4.14 $Y=2.41 $X2=4.14
+ $Y2=2.61
r140 34 35 5.14764 $w=2.58e-07 $l=8.5e-08 $layer=LI1_cond $X=4.14 $Y=2.41
+ $X2=4.14 $Y2=2.325
r141 30 32 5.96091 $w=4.33e-07 $l=2.25e-07 $layer=LI1_cond $X=3.87 $Y=0.812
+ $X2=4.095 $Y2=0.812
r142 28 42 4.78362 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=4.975 $Y=2.28
+ $X2=4.975 $Y2=2.48
r143 27 38 2.94836 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.975 $Y=1.615
+ $X2=4.975 $Y2=1.45
r144 27 28 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=4.975 $Y=1.615
+ $X2=4.975 $Y2=2.28
r145 26 34 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.27 $Y=2.41
+ $X2=4.14 $Y2=2.41
r146 25 42 6.08812 $w=3.39e-07 $l=1.14782e-07 $layer=LI1_cond $X=4.89 $Y=2.41
+ $X2=4.975 $Y2=2.48
r147 25 26 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=4.89 $Y=2.41
+ $X2=4.27 $Y2=2.41
r148 23 32 6.29128 $w=1.7e-07 $l=2.18e-07 $layer=LI1_cond $X=4.095 $Y=1.03
+ $X2=4.095 $Y2=0.812
r149 23 35 84.4866 $w=1.68e-07 $l=1.295e-06 $layer=LI1_cond $X=4.095 $Y=1.03
+ $X2=4.095 $Y2=2.325
r150 19 36 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.01 $Y=2.61
+ $X2=4.14 $Y2=2.61
r151 19 21 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=4.01 $Y=2.61
+ $X2=3.68 $Y2=2.61
r152 16 18 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.09 $Y=1.66
+ $X2=6.09 $Y2=2.235
r153 15 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.56 $Y=1.54
+ $X2=5.395 $Y2=1.54
r154 14 16 26.9307 $w=1.5e-07 $l=1.58745e-07 $layer=POLY_cond $X=6 $Y=1.54
+ $X2=6.09 $Y2=1.66
r155 14 15 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=6 $Y=1.54 $X2=5.56
+ $Y2=1.54
r156 12 46 305.096 $w=1.5e-07 $l=5.95e-07 $layer=POLY_cond $X=5.455 $Y=0.69
+ $X2=5.455 $Y2=1.285
r157 3 44 600 $w=1.7e-07 $l=2.66458e-07 $layer=licon1_PDIFF $count=1 $X=5.005
+ $Y=2.315 $X2=5.16 $Y2=2.515
r158 2 21 600 $w=1.7e-07 $l=3.64349e-07 $layer=licon1_PDIFF $count=1 $X=3.525
+ $Y=2.315 $X2=3.68 $Y2=2.61
r159 1 30 182 $w=1.7e-07 $l=3.02283e-07 $layer=licon1_NDIFF $count=1 $X=3.66
+ $Y=0.595 $X2=3.87 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_LS__DFRBP_1%A_319_392# 1 2 9 11 13 15 16 17 18 19 22 24
+ 25 26 28 29 31 32 36 37 38 41 43 45 46 49 54 55
c192 54 0 1.03964e-19 $X=1.92 $Y=0.867
c193 49 0 2.58586e-19 $X=2.61 $Y=1.49
c194 22 0 1.58258e-20 $X=3.585 $Y=0.805
c195 19 0 1.41973e-19 $X=3.145 $Y=1.275
c196 18 0 1.25323e-19 $X=3.51 $Y=1.275
c197 15 0 7.95804e-20 $X=2.935 $Y=3.075
c198 11 0 1.94586e-20 $X=2.55 $Y=1.41
c199 9 0 4.7274e-20 $X=2.425 $Y=2.46
r200 60 64 39.3878 $w=3.61e-07 $l=2.95e-07 $layer=POLY_cond $X=2.64 $Y=1.487
+ $X2=2.935 $Y2=1.487
r201 59 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.64
+ $Y=1.61 $X2=2.64 $Y2=1.61
r202 55 57 6.52312 $w=3.46e-07 $l=1.85e-07 $layer=LI1_cond $X=1.555 $Y=2.057
+ $X2=1.74 $Y2=2.057
r203 53 54 9.79992 $w=5.43e-07 $l=1.65e-07 $layer=LI1_cond $X=1.755 $Y=0.867
+ $X2=1.92 $Y2=0.867
r204 50 53 4.38928 $w=5.43e-07 $l=2e-07 $layer=LI1_cond $X=1.555 $Y=0.867
+ $X2=1.755 $Y2=0.867
r205 49 59 4.33136 $w=3.38e-07 $l=1.27279e-07 $layer=LI1_cond $X=2.61 $Y=1.49
+ $X2=2.625 $Y2=1.61
r206 48 49 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=2.61 $Y=1.14
+ $X2=2.61 $Y2=1.49
r207 46 48 15.37 $w=1.26e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.445 $Y=1.055
+ $X2=2.61 $Y2=1.14
r208 46 54 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=2.445 $Y=1.055
+ $X2=1.92 $Y2=1.055
r209 45 55 4.90539 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=1.555 $Y=1.865
+ $X2=1.555 $Y2=2.057
r210 44 50 7.70116 $w=1.7e-07 $l=2.73e-07 $layer=LI1_cond $X=1.555 $Y=1.14
+ $X2=1.555 $Y2=0.867
r211 44 45 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=1.555 $Y=1.14
+ $X2=1.555 $Y2=1.865
r212 39 41 458.926 $w=1.5e-07 $l=8.95e-07 $layer=POLY_cond $X=7.095 $Y=1.475
+ $X2=7.095 $Y2=0.58
r213 37 39 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.02 $Y=1.55
+ $X2=7.095 $Y2=1.475
r214 37 38 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=7.02 $Y=1.55
+ $X2=6.63 $Y2=1.55
r215 34 36 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.54 $Y=2.81
+ $X2=6.54 $Y2=2.235
r216 33 38 26.9307 $w=1.5e-07 $l=1.48324e-07 $layer=POLY_cond $X=6.54 $Y=1.66
+ $X2=6.63 $Y2=1.55
r217 33 36 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.54 $Y=1.66
+ $X2=6.54 $Y2=2.235
r218 31 34 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.54 $Y=2.9 $X2=6.54
+ $Y2=2.81
r219 31 32 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=6.54 $Y=2.9
+ $X2=6.54 $Y2=3.075
r220 30 43 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.995 $Y=3.15
+ $X2=3.905 $Y2=3.15
r221 29 32 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=6.45 $Y=3.15
+ $X2=6.54 $Y2=3.075
r222 29 30 1258.84 $w=1.5e-07 $l=2.455e-06 $layer=POLY_cond $X=6.45 $Y=3.15
+ $X2=3.995 $Y2=3.15
r223 26 28 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.905 $Y=2.81
+ $X2=3.905 $Y2=2.525
r224 25 43 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=3.905 $Y=3.075
+ $X2=3.905 $Y2=3.15
r225 24 26 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.905 $Y=2.9
+ $X2=3.905 $Y2=2.81
r226 24 25 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=3.905 $Y=2.9
+ $X2=3.905 $Y2=3.075
r227 20 22 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.585 $Y=1.2
+ $X2=3.585 $Y2=0.805
r228 19 64 44.9323 $w=3.61e-07 $l=2.99105e-07 $layer=POLY_cond $X=3.145 $Y=1.275
+ $X2=2.935 $Y2=1.487
r229 18 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.51 $Y=1.275
+ $X2=3.585 $Y2=1.2
r230 18 19 187.16 $w=1.5e-07 $l=3.65e-07 $layer=POLY_cond $X=3.51 $Y=1.275
+ $X2=3.145 $Y2=1.275
r231 16 43 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.815 $Y=3.15
+ $X2=3.905 $Y2=3.15
r232 16 17 412.777 $w=1.5e-07 $l=8.05e-07 $layer=POLY_cond $X=3.815 $Y=3.15
+ $X2=3.01 $Y2=3.15
r233 15 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.935 $Y=3.075
+ $X2=3.01 $Y2=3.15
r234 14 64 23.3725 $w=1.5e-07 $l=2.88e-07 $layer=POLY_cond $X=2.935 $Y=1.775
+ $X2=2.935 $Y2=1.487
r235 14 15 666.596 $w=1.5e-07 $l=1.3e-06 $layer=POLY_cond $X=2.935 $Y=1.775
+ $X2=2.935 $Y2=3.075
r236 11 60 12.0166 $w=3.61e-07 $l=9e-08 $layer=POLY_cond $X=2.55 $Y=1.487
+ $X2=2.64 $Y2=1.487
r237 11 61 16.6898 $w=3.61e-07 $l=1.25e-07 $layer=POLY_cond $X=2.55 $Y=1.487
+ $X2=2.425 $Y2=1.487
r238 11 13 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.55 $Y=1.41
+ $X2=2.55 $Y2=0.965
r239 7 61 23.3725 $w=1.5e-07 $l=2.88e-07 $layer=POLY_cond $X=2.425 $Y=1.775
+ $X2=2.425 $Y2=1.487
r240 7 9 351.245 $w=1.5e-07 $l=6.85e-07 $layer=POLY_cond $X=2.425 $Y=1.775
+ $X2=2.425 $Y2=2.46
r241 2 57 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.595
+ $Y=1.96 $X2=1.74 $Y2=2.085
r242 1 53 182 $w=1.7e-07 $l=3.85746e-07 $layer=licon1_NDIFF $count=1 $X=1.61
+ $Y=0.595 $X2=1.755 $Y2=0.915
.ends

.subckt PM_SKY130_FD_SC_LS__DFRBP_1%A_1482_48# 1 2 7 9 11 12 14 15 18 21 24 25
+ 38 40 44
c95 38 0 6.85463e-20 $X=8.885 $Y=1.85
c96 15 0 1.98491e-19 $X=8.485 $Y=0.985
r97 36 38 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=8.555 $Y=1.85
+ $X2=8.885 $Y2=1.85
r98 29 44 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=7.595 $Y=1.065
+ $X2=7.67 $Y2=1.065
r99 29 41 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=7.595 $Y=1.065
+ $X2=7.485 $Y2=1.065
r100 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.595
+ $Y=1.065 $X2=7.595 $Y2=1.065
r101 25 28 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=7.595 $Y=0.985
+ $X2=7.595 $Y2=1.065
r102 24 38 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.885 $Y=1.765
+ $X2=8.885 $Y2=1.85
r103 23 40 2.90768 $w=3.27e-07 $l=1.95944e-07 $layer=LI1_cond $X=8.885 $Y=1.07
+ $X2=8.727 $Y2=0.985
r104 23 24 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=8.885 $Y=1.07
+ $X2=8.885 $Y2=1.765
r105 19 40 2.90768 $w=3.27e-07 $l=8.5e-08 $layer=LI1_cond $X=8.727 $Y=0.9
+ $X2=8.727 $Y2=0.985
r106 19 21 7.89165 $w=4.83e-07 $l=3.2e-07 $layer=LI1_cond $X=8.727 $Y=0.9
+ $X2=8.727 $Y2=0.58
r107 18 32 4.37637 $w=3.93e-07 $l=1.5e-07 $layer=LI1_cond $X=8.555 $Y=2.532
+ $X2=8.405 $Y2=2.532
r108 17 36 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.555 $Y=1.935
+ $X2=8.555 $Y2=1.85
r109 17 18 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=8.555 $Y=1.935
+ $X2=8.555 $Y2=2.335
r110 16 25 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.76 $Y=0.985
+ $X2=7.595 $Y2=0.985
r111 15 40 3.78066 $w=1.7e-07 $l=2.42e-07 $layer=LI1_cond $X=8.485 $Y=0.985
+ $X2=8.727 $Y2=0.985
r112 15 16 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=8.485 $Y=0.985
+ $X2=7.76 $Y2=0.985
r113 12 14 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.67 $Y=2.28
+ $X2=7.67 $Y2=2.565
r114 11 12 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=7.67 $Y=2.19 $X2=7.67
+ $Y2=2.28
r115 10 44 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.67 $Y=1.23
+ $X2=7.67 $Y2=1.065
r116 10 11 373.161 $w=1.8e-07 $l=9.6e-07 $layer=POLY_cond $X=7.67 $Y=1.23
+ $X2=7.67 $Y2=2.19
r117 7 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.485 $Y=0.9
+ $X2=7.485 $Y2=1.065
r118 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=7.485 $Y=0.9
+ $X2=7.485 $Y2=0.58
r119 2 32 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=8.255
+ $Y=2.355 $X2=8.405 $Y2=2.565
r120 1 21 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=8.51
+ $Y=0.37 $X2=8.65 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_LS__DFRBP_1%A_1224_74# 1 2 9 12 13 15 16 17 18 20 23 25
+ 28 29 31 34 37 38 42 47 48 49 51 52 54 56
c164 51 0 1.04385e-19 $X=7.58 $Y=2.365
c165 29 0 1.79977e-19 $X=10.5 $Y=2.045
c166 17 0 1.98491e-19 $X=8.72 $Y=1.43
r167 57 64 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=8.495 $Y=1.43
+ $X2=8.63 $Y2=1.43
r168 57 61 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=8.495 $Y=1.43
+ $X2=8.435 $Y2=1.43
r169 56 59 3.07318 $w=2.98e-07 $l=8e-08 $layer=LI1_cond $X=8.48 $Y=1.43 $X2=8.48
+ $Y2=1.51
r170 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.495
+ $Y=1.43 $X2=8.495 $Y2=1.43
r171 53 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.665 $Y=1.51
+ $X2=7.58 $Y2=1.51
r172 52 59 4.061 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=8.33 $Y=1.51 $X2=8.48
+ $Y2=1.51
r173 52 53 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=8.33 $Y=1.51
+ $X2=7.665 $Y2=1.51
r174 50 54 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.58 $Y=1.595
+ $X2=7.58 $Y2=1.51
r175 50 51 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=7.58 $Y=1.595
+ $X2=7.58 $Y2=2.365
r176 48 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.495 $Y=1.51
+ $X2=7.58 $Y2=1.51
r177 48 49 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=7.495 $Y=1.51
+ $X2=7.16 $Y2=1.51
r178 47 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.075 $Y=1.425
+ $X2=7.16 $Y2=1.51
r179 46 47 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=7.075 $Y=0.73
+ $X2=7.075 $Y2=1.425
r180 42 51 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.495 $Y=2.53
+ $X2=7.58 $Y2=2.365
r181 42 44 21.1281 $w=3.28e-07 $l=6.05e-07 $layer=LI1_cond $X=7.495 $Y=2.53
+ $X2=6.89 $Y2=2.53
r182 38 46 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.99 $Y=0.565
+ $X2=7.075 $Y2=0.73
r183 38 40 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=6.99 $Y=0.565
+ $X2=6.695 $Y2=0.565
r184 32 37 34.7346 $w=1.65e-07 $l=1.72337e-07 $layer=POLY_cond $X=10.515
+ $Y=1.265 $X2=10.5 $Y2=1.43
r185 32 34 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=10.515 $Y=1.265
+ $X2=10.515 $Y2=0.645
r186 29 31 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=10.5 $Y=2.045
+ $X2=10.5 $Y2=2.54
r187 28 29 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=10.5 $Y=1.955
+ $X2=10.5 $Y2=2.045
r188 27 37 34.7346 $w=1.65e-07 $l=1.65e-07 $layer=POLY_cond $X=10.5 $Y=1.595
+ $X2=10.5 $Y2=1.43
r189 27 28 139.935 $w=1.8e-07 $l=3.6e-07 $layer=POLY_cond $X=10.5 $Y=1.595
+ $X2=10.5 $Y2=1.955
r190 26 36 5.16599 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=9.515 $Y=1.43
+ $X2=9.285 $Y2=1.43
r191 25 37 3.90195 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=10.41 $Y=1.43
+ $X2=10.5 $Y2=1.43
r192 25 26 156.501 $w=3.3e-07 $l=8.95e-07 $layer=POLY_cond $X=10.41 $Y=1.43
+ $X2=9.515 $Y2=1.43
r193 21 36 38.9663 $w=3.64e-07 $l=2.29783e-07 $layer=POLY_cond $X=9.44 $Y=1.265
+ $X2=9.285 $Y2=1.43
r194 21 23 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=9.44 $Y=1.265
+ $X2=9.44 $Y2=0.74
r195 18 36 61.4773 $w=3.64e-07 $l=3.98905e-07 $layer=POLY_cond $X=9.145 $Y=1.765
+ $X2=9.285 $Y2=1.43
r196 18 20 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=9.145 $Y=1.765
+ $X2=9.145 $Y2=2.4
r197 17 64 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=8.72 $Y=1.43 $X2=8.63
+ $Y2=1.43
r198 16 36 5.16599 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=9.055 $Y=1.43
+ $X2=9.285 $Y2=1.43
r199 16 17 58.5785 $w=3.3e-07 $l=3.35e-07 $layer=POLY_cond $X=9.055 $Y=1.43
+ $X2=8.72 $Y2=1.43
r200 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=8.63 $Y=2.28
+ $X2=8.63 $Y2=2.565
r201 12 13 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=8.63 $Y=2.19 $X2=8.63
+ $Y2=2.28
r202 11 64 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=8.63 $Y=1.595
+ $X2=8.63 $Y2=1.43
r203 11 12 231.282 $w=1.8e-07 $l=5.95e-07 $layer=POLY_cond $X=8.63 $Y=1.595
+ $X2=8.63 $Y2=2.19
r204 7 61 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.435 $Y=1.265
+ $X2=8.435 $Y2=1.43
r205 7 9 351.245 $w=1.5e-07 $l=6.85e-07 $layer=POLY_cond $X=8.435 $Y=1.265
+ $X2=8.435 $Y2=0.58
r206 2 44 600 $w=1.7e-07 $l=9.22307e-07 $layer=licon1_PDIFF $count=1 $X=6.615
+ $Y=1.735 $X2=6.89 $Y2=2.53
r207 1 40 182 $w=1.7e-07 $l=6.65395e-07 $layer=licon1_NDIFF $count=1 $X=6.12
+ $Y=0.37 $X2=6.695 $Y2=0.565
.ends

.subckt PM_SKY130_FD_SC_LS__DFRBP_1%A_2026_424# 1 2 9 11 13 16 20 24 27
r50 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.965
+ $Y=1.465 $X2=10.965 $Y2=1.465
r51 22 27 0.364692 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=10.44 $Y=1.465
+ $X2=10.315 $Y2=1.465
r52 22 24 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=10.44 $Y=1.465
+ $X2=10.965 $Y2=1.465
r53 18 27 6.46576 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=10.315 $Y=1.63
+ $X2=10.315 $Y2=1.465
r54 18 20 29.5025 $w=2.48e-07 $l=6.4e-07 $layer=LI1_cond $X=10.315 $Y=1.63
+ $X2=10.315 $Y2=2.27
r55 14 27 6.46576 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=10.315 $Y=1.3
+ $X2=10.315 $Y2=1.465
r56 14 16 30.4245 $w=2.48e-07 $l=6.6e-07 $layer=LI1_cond $X=10.315 $Y=1.3
+ $X2=10.315 $Y2=0.64
r57 11 25 61.4066 $w=2.86e-07 $l=3.24037e-07 $layer=POLY_cond $X=11.015 $Y=1.765
+ $X2=10.965 $Y2=1.465
r58 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=11.015 $Y=1.765
+ $X2=11.015 $Y2=2.4
r59 7 25 38.6549 $w=2.86e-07 $l=1.88348e-07 $layer=POLY_cond $X=11.015 $Y=1.3
+ $X2=10.965 $Y2=1.465
r60 7 9 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=11.015 $Y=1.3
+ $X2=11.015 $Y2=0.74
r61 2 20 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=10.13
+ $Y=2.12 $X2=10.275 $Y2=2.27
r62 1 16 182 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_NDIFF $count=1 $X=10.155
+ $Y=0.37 $X2=10.3 $Y2=0.64
.ends

.subckt PM_SKY130_FD_SC_LS__DFRBP_1%VPWR 1 2 3 4 5 6 7 8 25 27 31 35 39 43 49 51
+ 55 59 63 65 70 75 83 88 93 103 104 110 113 116 119 122 125 128
r155 128 129 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r156 125 126 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r157 123 126 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.88 $Y2=3.33
r158 122 123 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r159 119 120 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r160 116 117 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r161 113 114 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r162 110 111 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r163 107 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r164 104 129 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=10.8 $Y2=3.33
r165 103 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r166 101 128 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=10.905 $Y=3.33
+ $X2=10.757 $Y2=3.33
r167 101 103 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=10.905 $Y=3.33
+ $X2=11.28 $Y2=3.33
r168 100 129 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=10.8 $Y2=3.33
r169 99 100 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r170 97 100 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=10.32 $Y2=3.33
r171 97 126 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=8.88 $Y2=3.33
r172 96 99 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=9.36 $Y=3.33
+ $X2=10.32 $Y2=3.33
r173 96 97 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r174 94 125 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=9.025 $Y=3.33
+ $X2=8.917 $Y2=3.33
r175 94 96 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=9.025 $Y=3.33
+ $X2=9.36 $Y2=3.33
r176 93 128 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=10.61 $Y=3.33
+ $X2=10.757 $Y2=3.33
r177 93 99 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=10.61 $Y=3.33
+ $X2=10.32 $Y2=3.33
r178 92 123 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r179 92 120 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6 $Y2=3.33
r180 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r181 89 119 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.03 $Y=3.33
+ $X2=5.905 $Y2=3.33
r182 89 91 91.9893 $w=1.68e-07 $l=1.41e-06 $layer=LI1_cond $X=6.03 $Y=3.33
+ $X2=7.44 $Y2=3.33
r183 88 122 6.47928 $w=1.7e-07 $l=1.12e-07 $layer=LI1_cond $X=7.835 $Y=3.33
+ $X2=7.947 $Y2=3.33
r184 88 91 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=7.835 $Y=3.33
+ $X2=7.44 $Y2=3.33
r185 87 117 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=4.56 $Y2=3.33
r186 86 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r187 84 116 8.88104 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=4.785 $Y=3.33
+ $X2=4.612 $Y2=3.33
r188 84 86 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=4.785 $Y=3.33
+ $X2=5.52 $Y2=3.33
r189 83 119 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.78 $Y=3.33
+ $X2=5.905 $Y2=3.33
r190 83 86 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=5.78 $Y=3.33
+ $X2=5.52 $Y2=3.33
r191 82 117 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r192 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r193 79 82 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=4.08 $Y2=3.33
r194 79 114 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r195 78 81 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.64 $Y=3.33
+ $X2=4.08 $Y2=3.33
r196 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r197 76 113 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.355 $Y=3.33
+ $X2=2.19 $Y2=3.33
r198 76 78 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.355 $Y=3.33
+ $X2=2.64 $Y2=3.33
r199 75 116 8.88104 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=4.44 $Y=3.33
+ $X2=4.612 $Y2=3.33
r200 75 81 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=4.44 $Y=3.33
+ $X2=4.08 $Y2=3.33
r201 74 114 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r202 74 111 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r203 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r204 71 110 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.345 $Y=3.33
+ $X2=1.18 $Y2=3.33
r205 71 73 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.345 $Y=3.33
+ $X2=1.68 $Y2=3.33
r206 70 113 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.025 $Y=3.33
+ $X2=2.19 $Y2=3.33
r207 70 73 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.025 $Y=3.33
+ $X2=1.68 $Y2=3.33
r208 69 111 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r209 69 108 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r210 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r211 66 107 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.182 $Y2=3.33
r212 66 68 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.72 $Y2=3.33
r213 65 110 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.015 $Y=3.33
+ $X2=1.18 $Y2=3.33
r214 65 68 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.015 $Y=3.33
+ $X2=0.72 $Y2=3.33
r215 63 120 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=5.76 $Y=3.33
+ $X2=6 $Y2=3.33
r216 63 87 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=5.76 $Y=3.33
+ $X2=5.52 $Y2=3.33
r217 59 62 16.2123 $w=2.93e-07 $l=4.15e-07 $layer=LI1_cond $X=10.757 $Y=1.985
+ $X2=10.757 $Y2=2.4
r218 57 128 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=10.757 $Y=3.245
+ $X2=10.757 $Y2=3.33
r219 57 62 33.0107 $w=2.93e-07 $l=8.45e-07 $layer=LI1_cond $X=10.757 $Y=3.245
+ $X2=10.757 $Y2=2.4
r220 53 125 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=8.917 $Y=3.245
+ $X2=8.917 $Y2=3.33
r221 53 55 52.262 $w=2.13e-07 $l=9.75e-07 $layer=LI1_cond $X=8.917 $Y=3.245
+ $X2=8.917 $Y2=2.27
r222 52 122 6.47928 $w=1.7e-07 $l=1.13e-07 $layer=LI1_cond $X=8.06 $Y=3.33
+ $X2=7.947 $Y2=3.33
r223 51 125 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=8.81 $Y=3.33
+ $X2=8.917 $Y2=3.33
r224 51 52 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=8.81 $Y=3.33
+ $X2=8.06 $Y2=3.33
r225 47 122 0.355529 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=7.947 $Y=3.245
+ $X2=7.947 $Y2=3.33
r226 47 49 34.8294 $w=2.23e-07 $l=6.8e-07 $layer=LI1_cond $X=7.947 $Y=3.245
+ $X2=7.947 $Y2=2.565
r227 43 46 31.5769 $w=2.48e-07 $l=6.85e-07 $layer=LI1_cond $X=5.905 $Y=1.905
+ $X2=5.905 $Y2=2.59
r228 41 119 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.905 $Y=3.245
+ $X2=5.905 $Y2=3.33
r229 41 46 30.194 $w=2.48e-07 $l=6.55e-07 $layer=LI1_cond $X=5.905 $Y=3.245
+ $X2=5.905 $Y2=2.59
r230 37 116 1.03204 $w=3.45e-07 $l=8.5e-08 $layer=LI1_cond $X=4.612 $Y=3.245
+ $X2=4.612 $Y2=3.33
r231 37 39 16.5351 $w=3.43e-07 $l=4.95e-07 $layer=LI1_cond $X=4.612 $Y=3.245
+ $X2=4.612 $Y2=2.75
r232 33 113 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.19 $Y=3.245
+ $X2=2.19 $Y2=3.33
r233 33 35 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=2.19 $Y=3.245
+ $X2=2.19 $Y2=2.835
r234 29 110 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.18 $Y=3.245
+ $X2=1.18 $Y2=3.33
r235 29 31 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=1.18 $Y=3.245
+ $X2=1.18 $Y2=2.835
r236 25 107 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.182 $Y2=3.33
r237 25 27 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.24 $Y2=2.75
r238 8 62 300 $w=1.7e-07 $l=3.60832e-07 $layer=licon1_PDIFF $count=2 $X=10.575
+ $Y=2.12 $X2=10.76 $Y2=2.4
r239 8 59 600 $w=1.7e-07 $l=2.74317e-07 $layer=licon1_PDIFF $count=1 $X=10.575
+ $Y=2.12 $X2=10.79 $Y2=1.985
r240 7 55 300 $w=1.7e-07 $l=2.53969e-07 $layer=licon1_PDIFF $count=2 $X=8.705
+ $Y=2.355 $X2=8.92 $Y2=2.27
r241 6 49 600 $w=1.7e-07 $l=2.84341e-07 $layer=licon1_PDIFF $count=1 $X=7.745
+ $Y=2.355 $X2=7.92 $Y2=2.565
r242 5 46 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=5.72
+ $Y=1.735 $X2=5.865 $Y2=2.59
r243 5 43 400 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_PDIFF $count=1 $X=5.72
+ $Y=1.735 $X2=5.865 $Y2=1.905
r244 4 39 600 $w=1.7e-07 $l=5.41872e-07 $layer=licon1_PDIFF $count=1 $X=4.37
+ $Y=2.315 $X2=4.61 $Y2=2.75
r245 3 35 600 $w=1.7e-07 $l=9.47035e-07 $layer=licon1_PDIFF $count=1 $X=2.04
+ $Y=1.96 $X2=2.19 $Y2=2.835
r246 2 31 600 $w=1.7e-07 $l=3.62319e-07 $layer=licon1_PDIFF $count=1 $X=1.03
+ $Y=2.54 $X2=1.18 $Y2=2.835
r247 1 27 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.54 $X2=0.28 $Y2=2.75
.ends

.subckt PM_SKY130_FD_SC_LS__DFRBP_1%A_38_78# 1 2 3 4 13 17 20 21 25 29 32 33 36
+ 38 42 43 44 46 49 52
c130 52 0 1.41973e-19 $X=3.755 $Y=1.285
c131 49 0 1.78683e-19 $X=3.41 $Y=1.035
c132 44 0 4.7274e-20 $X=1.965 $Y=2.5
c133 33 0 2.12927e-19 $X=3.67 $Y=2.27
c134 29 0 1.21972e-19 $X=3.37 $Y=0.81
r135 46 48 1.5 $w=2.44e-07 $l=3e-08 $layer=LI1_cond $X=3.205 $Y=2.495 $X2=3.205
+ $Y2=2.525
r136 45 46 11.25 $w=2.44e-07 $l=2.25e-07 $layer=LI1_cond $X=3.205 $Y=2.27
+ $X2=3.205 $Y2=2.495
r137 43 44 4.62121 $w=1.78e-07 $l=7.5e-08 $layer=LI1_cond $X=1.89 $Y=2.5
+ $X2=1.965 $Y2=2.5
r138 38 40 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=0.335 $Y=0.6
+ $X2=0.335 $Y2=0.745
r139 35 52 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.755 $Y=1.37
+ $X2=3.755 $Y2=1.285
r140 35 36 53.1711 $w=1.68e-07 $l=8.15e-07 $layer=LI1_cond $X=3.755 $Y=1.37
+ $X2=3.755 $Y2=2.185
r141 34 45 2.85362 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=3.345 $Y=2.27
+ $X2=3.205 $Y2=2.27
r142 33 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.67 $Y=2.27
+ $X2=3.755 $Y2=2.185
r143 33 34 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=3.67 $Y=2.27
+ $X2=3.345 $Y2=2.27
r144 32 52 21.0727 $w=1.68e-07 $l=3.23e-07 $layer=LI1_cond $X=3.432 $Y=1.285
+ $X2=3.755 $Y2=1.285
r145 32 49 8.92683 $w=2.03e-07 $l=1.65e-07 $layer=LI1_cond $X=3.432 $Y=1.2
+ $X2=3.432 $Y2=1.035
r146 27 49 6.16968 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=3.41 $Y=0.91
+ $X2=3.41 $Y2=1.035
r147 27 29 4.60977 $w=2.48e-07 $l=1e-07 $layer=LI1_cond $X=3.41 $Y=0.91 $X2=3.41
+ $Y2=0.81
r148 25 46 2.85362 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=3.065 $Y=2.495
+ $X2=3.205 $Y2=2.495
r149 25 44 71.7647 $w=1.68e-07 $l=1.1e-06 $layer=LI1_cond $X=3.065 $Y=2.495
+ $X2=1.965 $Y2=2.495
r150 24 43 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=1.53 $Y=2.505
+ $X2=1.89 $Y2=2.505
r151 22 42 0.695019 $w=2.7e-07 $l=3.60555e-07 $layer=LI1_cond $X=0.89 $Y=2.445
+ $X2=0.565 $Y2=2.52
r152 21 24 7.78061 $w=1.96e-07 $l=1.52069e-07 $layer=LI1_cond $X=1.405 $Y=2.445
+ $X2=1.53 $Y2=2.505
r153 21 22 21.9818 $w=2.68e-07 $l=5.15e-07 $layer=LI1_cond $X=1.405 $Y=2.445
+ $X2=0.89 $Y2=2.445
r154 20 42 5.99569 $w=2.25e-07 $l=2.96985e-07 $layer=LI1_cond $X=0.775 $Y=2.31
+ $X2=0.565 $Y2=2.52
r155 19 20 96.5562 $w=1.68e-07 $l=1.48e-06 $layer=LI1_cond $X=0.775 $Y=0.83
+ $X2=0.775 $Y2=2.31
r156 15 42 5.99569 $w=2.25e-07 $l=1.87083e-07 $layer=LI1_cond $X=0.705 $Y=2.63
+ $X2=0.565 $Y2=2.52
r157 15 17 4.93904 $w=2.78e-07 $l=1.2e-07 $layer=LI1_cond $X=0.705 $Y=2.63
+ $X2=0.705 $Y2=2.75
r158 14 40 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.5 $Y=0.745
+ $X2=0.335 $Y2=0.745
r159 13 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.69 $Y=0.745
+ $X2=0.775 $Y2=0.83
r160 13 14 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=0.69 $Y=0.745
+ $X2=0.5 $Y2=0.745
r161 4 48 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=3.085
+ $Y=2.315 $X2=3.23 $Y2=2.525
r162 3 17 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=2.54 $X2=0.73 $Y2=2.75
r163 2 29 182 $w=1.7e-07 $l=2.82046e-07 $layer=licon1_NDIFF $count=1 $X=3.215
+ $Y=0.595 $X2=3.37 $Y2=0.81
r164 1 38 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.19
+ $Y=0.39 $X2=0.335 $Y2=0.6
.ends

.subckt PM_SKY130_FD_SC_LS__DFRBP_1%Q_N 1 2 9 11 12 13 26
c24 12 0 1.79977e-19 $X=9.84 $Y=2.405
r25 26 27 5.27602 $w=6.88e-07 $l=1.75e-07 $layer=LI1_cond $X=9.605 $Y=1.985
+ $X2=9.605 $Y2=1.81
r26 13 23 0.693379 $w=6.88e-07 $l=4e-08 $layer=LI1_cond $X=9.605 $Y=2.775
+ $X2=9.605 $Y2=2.815
r27 12 13 6.41375 $w=6.88e-07 $l=3.7e-07 $layer=LI1_cond $X=9.605 $Y=2.405
+ $X2=9.605 $Y2=2.775
r28 12 17 4.33362 $w=6.88e-07 $l=2.5e-07 $layer=LI1_cond $X=9.605 $Y=2.405
+ $X2=9.605 $Y2=2.155
r29 11 17 2.08014 $w=6.88e-07 $l=1.2e-07 $layer=LI1_cond $X=9.605 $Y=2.035
+ $X2=9.605 $Y2=2.155
r30 11 26 0.866723 $w=6.88e-07 $l=5e-08 $layer=LI1_cond $X=9.605 $Y=2.035
+ $X2=9.605 $Y2=1.985
r31 9 27 38.267 $w=3.88e-07 $l=1.295e-06 $layer=LI1_cond $X=9.755 $Y=0.515
+ $X2=9.755 $Y2=1.81
r32 2 26 200 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=3 $X=9.22
+ $Y=1.84 $X2=9.37 $Y2=1.985
r33 2 23 200 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=3 $X=9.22
+ $Y=1.84 $X2=9.37 $Y2=2.815
r34 1 9 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=9.515
+ $Y=0.37 $X2=9.725 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__DFRBP_1%Q 1 2 9 10 11 24 27 35
r22 33 35 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=11.35 $Y=1.13
+ $X2=11.35 $Y2=1.82
r23 25 27 1.12043 $w=3.58e-07 $l=3.5e-08 $layer=LI1_cond $X=11.255 $Y=2
+ $X2=11.255 $Y2=2.035
r24 17 24 0.622942 $w=3.68e-07 $l=2e-08 $layer=LI1_cond $X=11.25 $Y=0.945
+ $X2=11.25 $Y2=0.925
r25 11 25 0.800308 $w=3.58e-07 $l=2.5e-08 $layer=LI1_cond $X=11.255 $Y=1.975
+ $X2=11.255 $Y2=2
r26 11 35 8.1909 $w=3.58e-07 $l=1.55e-07 $layer=LI1_cond $X=11.255 $Y=1.975
+ $X2=11.255 $Y2=1.82
r27 11 30 24.1693 $w=3.58e-07 $l=7.55e-07 $layer=LI1_cond $X=11.255 $Y=2.06
+ $X2=11.255 $Y2=2.815
r28 11 27 0.800308 $w=3.58e-07 $l=2.5e-08 $layer=LI1_cond $X=11.255 $Y=2.06
+ $X2=11.255 $Y2=2.035
r29 10 33 8.16504 $w=3.68e-07 $l=1.53e-07 $layer=LI1_cond $X=11.25 $Y=0.977
+ $X2=11.25 $Y2=1.13
r30 10 17 0.996707 $w=3.68e-07 $l=3.2e-08 $layer=LI1_cond $X=11.25 $Y=0.977
+ $X2=11.25 $Y2=0.945
r31 10 24 1.02785 $w=3.68e-07 $l=3.3e-08 $layer=LI1_cond $X=11.25 $Y=0.892
+ $X2=11.25 $Y2=0.925
r32 9 10 11.7425 $w=3.68e-07 $l=3.77e-07 $layer=LI1_cond $X=11.25 $Y=0.515
+ $X2=11.25 $Y2=0.892
r33 2 11 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=11.09
+ $Y=1.84 $X2=11.24 $Y2=1.985
r34 2 30 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=11.09
+ $Y=1.84 $X2=11.24 $Y2=2.815
r35 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=11.09
+ $Y=0.37 $X2=11.23 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__DFRBP_1%VGND 1 2 3 4 5 6 21 23 27 31 35 39 43 45 50
+ 55 63 68 75 76 79 82 86 92 95 98
c114 76 0 1.90308e-19 $X=11.28 $Y=0
r115 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=0 $X2=10.8
+ $Y2=0
r116 95 96 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r117 92 93 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r118 86 89 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=5.16 $Y=0 $X2=5.16
+ $Y2=0.325
r119 86 87 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r120 82 83 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r121 80 83 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r122 79 80 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r123 76 99 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=10.8 $Y2=0
r124 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r125 73 98 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.895 $Y=0
+ $X2=10.77 $Y2=0
r126 73 75 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=10.895 $Y=0
+ $X2=11.28 $Y2=0
r127 72 99 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=10.8 $Y2=0
r128 72 96 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=9.36 $Y2=0
r129 71 72 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r130 69 95 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.39 $Y=0 $X2=9.265
+ $Y2=0
r131 69 71 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=9.39 $Y=0 $X2=10.32
+ $Y2=0
r132 68 98 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.645 $Y=0
+ $X2=10.77 $Y2=0
r133 68 71 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=10.645 $Y=0
+ $X2=10.32 $Y2=0
r134 67 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=9.36
+ $Y2=0
r135 67 93 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=7.92
+ $Y2=0
r136 66 67 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r137 64 92 10.7288 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=7.995 $Y=0 $X2=7.765
+ $Y2=0
r138 64 66 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=7.995 $Y=0 $X2=8.88
+ $Y2=0
r139 63 95 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.14 $Y=0 $X2=9.265
+ $Y2=0
r140 63 66 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=9.14 $Y=0 $X2=8.88
+ $Y2=0
r141 62 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=7.92
+ $Y2=0
r142 61 62 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r143 59 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r144 58 61 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=5.52 $Y=0 $X2=7.44
+ $Y2=0
r145 58 59 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r146 56 86 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.325 $Y=0 $X2=5.16
+ $Y2=0
r147 56 58 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=5.325 $Y=0
+ $X2=5.52 $Y2=0
r148 55 92 10.7288 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=7.535 $Y=0 $X2=7.765
+ $Y2=0
r149 55 61 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=7.535 $Y=0 $X2=7.44
+ $Y2=0
r150 54 87 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=2.64 $Y=0 $X2=5.04
+ $Y2=0
r151 54 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r152 53 54 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r153 51 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.42 $Y=0 $X2=2.255
+ $Y2=0
r154 51 53 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=2.42 $Y=0 $X2=2.64
+ $Y2=0
r155 50 86 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.995 $Y=0 $X2=5.16
+ $Y2=0
r156 50 53 153.642 $w=1.68e-07 $l=2.355e-06 $layer=LI1_cond $X=4.995 $Y=0
+ $X2=2.64 $Y2=0
r157 48 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r158 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r159 45 79 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.03 $Y=0 $X2=1.155
+ $Y2=0
r160 45 47 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1.03 $Y=0 $X2=0.72
+ $Y2=0
r161 43 62 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=5.76 $Y=0
+ $X2=7.44 $Y2=0
r162 43 59 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=5.76 $Y=0
+ $X2=5.52 $Y2=0
r163 39 41 20.744 $w=2.48e-07 $l=4.5e-07 $layer=LI1_cond $X=10.77 $Y=0.515
+ $X2=10.77 $Y2=0.965
r164 37 98 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=10.77 $Y=0.085
+ $X2=10.77 $Y2=0
r165 37 39 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=10.77 $Y=0.085
+ $X2=10.77 $Y2=0.515
r166 33 95 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.265 $Y=0.085
+ $X2=9.265 $Y2=0
r167 33 35 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=9.265 $Y=0.085
+ $X2=9.265 $Y2=0.515
r168 29 92 1.85547 $w=4.6e-07 $l=8.5e-08 $layer=LI1_cond $X=7.765 $Y=0.085
+ $X2=7.765 $Y2=0
r169 29 31 12.2208 $w=4.58e-07 $l=4.7e-07 $layer=LI1_cond $X=7.765 $Y=0.085
+ $X2=7.765 $Y2=0.555
r170 25 82 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.255 $Y=0.085
+ $X2=2.255 $Y2=0
r171 25 27 22.0012 $w=3.28e-07 $l=6.3e-07 $layer=LI1_cond $X=2.255 $Y=0.085
+ $X2=2.255 $Y2=0.715
r172 24 79 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.28 $Y=0 $X2=1.155
+ $Y2=0
r173 23 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.09 $Y=0 $X2=2.255
+ $Y2=0
r174 23 24 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=2.09 $Y=0 $X2=1.28
+ $Y2=0
r175 19 79 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.155 $Y=0.085
+ $X2=1.155 $Y2=0
r176 19 21 23.7403 $w=2.48e-07 $l=5.15e-07 $layer=LI1_cond $X=1.155 $Y=0.085
+ $X2=1.155 $Y2=0.6
r177 6 41 182 $w=1.7e-07 $l=6.87768e-07 $layer=licon1_NDIFF $count=1 $X=10.59
+ $Y=0.37 $X2=10.79 $Y2=0.965
r178 6 39 182 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_NDIFF $count=1 $X=10.59
+ $Y=0.37 $X2=10.79 $Y2=0.515
r179 5 35 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=9.08
+ $Y=0.37 $X2=9.225 $Y2=0.515
r180 4 31 182 $w=1.7e-07 $l=2.82754e-07 $layer=licon1_NDIFF $count=1 $X=7.56
+ $Y=0.37 $X2=7.765 $Y2=0.555
r181 3 89 182 $w=1.7e-07 $l=3.63731e-07 $layer=licon1_NDIFF $count=1 $X=4.94
+ $Y=0.595 $X2=5.16 $Y2=0.325
r182 2 27 182 $w=1.7e-07 $l=2.63249e-07 $layer=licon1_NDIFF $count=1 $X=2.045
+ $Y=0.595 $X2=2.255 $Y2=0.715
r183 1 21 182 $w=1.7e-07 $l=2.86182e-07 $layer=licon1_NDIFF $count=1 $X=1.015
+ $Y=0.39 $X2=1.195 $Y2=0.6
.ends

