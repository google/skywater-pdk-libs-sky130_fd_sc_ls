# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ls__buf_8
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ls__buf_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.760000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.837000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.350000 1.430000 1.780000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  2.249300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.960000 0.350000 2.130000 0.960000 ;
        RECT 1.960000 0.960000 5.145000 1.130000 ;
        RECT 1.970000 1.800000 5.155000 1.970000 ;
        RECT 1.970000 1.970000 2.300000 2.980000 ;
        RECT 2.810000 0.350000 3.140000 0.960000 ;
        RECT 2.920000 1.970000 3.250000 2.980000 ;
        RECT 3.810000 0.350000 4.140000 0.960000 ;
        RECT 3.870000 1.970000 4.200000 2.980000 ;
        RECT 4.810000 0.350000 5.145000 0.960000 ;
        RECT 4.820000 1.970000 5.155000 2.980000 ;
        RECT 4.975000 1.130000 5.145000 1.800000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 5.760000 0.085000 ;
        RECT 0.545000  0.085000 0.875000 0.840000 ;
        RECT 1.450000  0.085000 1.780000 0.840000 ;
        RECT 2.310000  0.085000 2.640000 0.790000 ;
        RECT 3.310000  0.085000 3.640000 0.790000 ;
        RECT 4.310000  0.085000 4.640000 0.790000 ;
        RECT 5.315000  0.085000 5.645000 1.130000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.760000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 5.760000 3.415000 ;
        RECT 0.650000 2.290000 0.820000 3.245000 ;
        RECT 1.550000 2.290000 1.800000 3.245000 ;
        RECT 2.500000 2.140000 2.750000 3.245000 ;
        RECT 3.450000 2.140000 3.700000 3.245000 ;
        RECT 4.400000 2.140000 4.650000 3.245000 ;
        RECT 5.350000 1.820000 5.600000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 5.760000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.115000 0.350000 0.365000 1.010000 ;
      RECT 0.115000 1.010000 1.770000 1.180000 ;
      RECT 0.120000 1.950000 1.770000 2.120000 ;
      RECT 0.120000 2.120000 0.450000 2.980000 ;
      RECT 1.020000 2.120000 1.350000 2.980000 ;
      RECT 1.100000 0.350000 1.270000 1.010000 ;
      RECT 1.600000 1.180000 1.770000 1.300000 ;
      RECT 1.600000 1.300000 4.805000 1.630000 ;
      RECT 1.600000 1.630000 1.770000 1.950000 ;
  END
END sky130_fd_sc_ls__buf_8
