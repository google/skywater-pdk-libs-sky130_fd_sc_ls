* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__bufbuf_16 A VGND VNB VPB VPWR X
M1000 a_588_74# a_203_74# VGND VNB nshort w=740000u l=150000u
+  ad=6.216e+11p pd=6.12e+06u as=3.3855e+12p ps=2.987e+07u
M1001 a_203_74# a_27_368# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=6.664e+11p pd=5.67e+06u as=4.7712e+12p ps=3.988e+07u
M1002 VGND a_588_74# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=1.6576e+12p ps=1.632e+07u
M1003 X a_588_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=2.744e+12p pd=2.282e+07u as=0p ps=0u
M1004 X a_588_74# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR a_203_74# a_588_74# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=1.008e+12p ps=8.52e+06u
M1006 VGND a_203_74# a_588_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_588_74# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_588_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 X a_588_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 X a_588_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 X a_588_74# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND a_588_74# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 X a_588_74# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND a_588_74# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR a_588_74# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_588_74# a_203_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR a_588_74# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 X a_588_74# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR a_588_74# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR a_588_74# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 X a_588_74# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND a_588_74# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VGND a_203_74# a_588_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND a_588_74# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VGND a_27_368# a_203_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=4.181e+11p ps=4.09e+06u
M1026 VPWR a_588_74# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_588_74# a_203_74# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VPWR a_203_74# a_588_74# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_203_74# a_27_368# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VPWR A a_27_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.304e+11p ps=2.83e+06u
M1031 a_203_74# a_27_368# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_588_74# a_203_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 X a_588_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 X a_588_74# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 X a_588_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 VPWR a_203_74# a_588_74# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 VGND a_588_74# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 X a_588_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 X a_588_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1040 VGND a_588_74# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1041 a_588_74# a_203_74# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1042 VGND a_588_74# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1043 VPWR a_27_368# a_203_74# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1044 VPWR a_588_74# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1045 X a_588_74# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1046 a_588_74# a_203_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1047 VPWR a_588_74# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1048 VGND a_203_74# a_588_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1049 VGND A a_27_368# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1050 a_203_74# a_27_368# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1051 VPWR a_588_74# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
