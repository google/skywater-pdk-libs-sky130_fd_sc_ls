* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__o41a_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
M1000 X a_110_48# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=6.72e+11p pd=5.68e+06u as=1.6953e+12p ps=1.387e+07u
M1001 a_523_124# A4 VGND VNB nshort w=640000u l=150000u
+  ad=1.1456e+12p pd=1.126e+07u as=1.69995e+12p ps=1.463e+07u
M1002 a_523_124# A3 VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_523_124# B1 a_110_48# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1004 VPWR a_110_48# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_523_124# A2 VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 X a_110_48# VGND VNB nshort w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=0p ps=0u
M1007 a_523_124# A1 VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_1213_368# A1 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=7.28e+11p pd=5.78e+06u as=0p ps=0u
M1009 VGND A1 a_523_124# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_110_48# B1 VPWR VPB phighvt w=840000u l=150000u
+  ad=5.992e+11p pd=5.14e+06u as=0p ps=0u
M1011 a_110_48# B1 a_523_124# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 X a_110_48# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND A3 a_523_124# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 X a_110_48# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_762_368# A3 a_851_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=1.0528e+12p pd=8.6e+06u as=6.72e+11p ps=5.68e+06u
M1016 VGND a_110_48# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_762_368# A2 a_1213_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR B1 a_110_48# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_851_368# A3 a_762_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND A2 a_523_124# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPWR a_110_48# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_851_368# A4 a_110_48# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_1213_368# A2 a_762_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND a_110_48# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_110_48# A4 a_851_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VGND A4 a_523_124# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VPWR A1 a_1213_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
