* File: sky130_fd_sc_ls__nor4_2.spice
* Created: Wed Sep  2 11:15:29 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__nor4_2.pex.spice"
.subckt sky130_fd_sc_ls__nor4_2  VNB VPB C D B A Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A	A
* B	B
* D	D
* C	C
* VPB	VPB
* VNB	VNB
MM1007 N_Y_M1007_d N_D_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.74 AD=0.1184
+ AS=0.3329 PD=1.06 PS=3 NRD=6.48 NRS=4.86 M=1 R=4.93333 SA=75000.4 SB=75001.8
+ A=0.111 P=1.78 MULT=1
MM1004 N_VGND_M1004_d N_C_M1004_g N_Y_M1007_d VNB NSHORT L=0.15 W=0.74 AD=0.1554
+ AS=0.1184 PD=1.16 PS=1.06 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.8 SB=75001.3
+ A=0.111 P=1.78 MULT=1
MM1010 N_Y_M1010_d N_B_M1010_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.74 AD=0.1036
+ AS=0.1554 PD=1.02 PS=1.16 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.4 SB=75000.7
+ A=0.111 P=1.78 MULT=1
MM1000 N_VGND_M1000_d N_A_M1000_g N_Y_M1010_d VNB NSHORT L=0.15 W=0.74 AD=0.2627
+ AS=0.1036 PD=2.19 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.8 SB=75000.3
+ A=0.111 P=1.78 MULT=1
MM1001 N_A_27_368#_M1001_d N_C_M1001_g N_A_116_368#_M1001_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.3304 AS=0.1764 PD=2.83 PS=1.435 NRD=1.7533 NRS=2.6201 M=1
+ R=7.46667 SA=75000.2 SB=75003.5 A=0.168 P=2.54 MULT=1
MM1003 N_Y_M1003_d N_D_M1003_g N_A_116_368#_M1001_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.182 AS=0.1764 PD=1.445 PS=1.435 NRD=3.5066 NRS=3.5066 M=1 R=7.46667
+ SA=75000.7 SB=75003.1 A=0.168 P=2.54 MULT=1
MM1011 N_Y_M1003_d N_D_M1011_g N_A_116_368#_M1011_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.182 AS=0.168 PD=1.445 PS=1.42 NRD=4.3931 NRS=1.7533 M=1 R=7.46667
+ SA=75001.2 SB=75002.6 A=0.168 P=2.54 MULT=1
MM1006 N_A_27_368#_M1006_d N_C_M1006_g N_A_116_368#_M1011_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.1848 AS=0.168 PD=1.45 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.6 SB=75002.1 A=0.168 P=2.54 MULT=1
MM1008 N_A_27_368#_M1006_d N_B_M1008_g N_A_490_368#_M1008_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.1848 AS=0.2184 PD=1.45 PS=1.51 NRD=7.0329 NRS=8.7862 M=1 R=7.46667
+ SA=75002.1 SB=75001.7 A=0.168 P=2.54 MULT=1
MM1002 N_VPWR_M1002_d N_A_M1002_g N_A_490_368#_M1008_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.2184 PD=1.42 PS=1.51 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75002.6 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1005 N_VPWR_M1002_d N_A_M1005_g N_A_490_368#_M1005_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75003.1 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1009 N_A_27_368#_M1009_d N_B_M1009_g N_A_490_368#_M1005_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75003.5 SB=75000.2 A=0.168 P=2.54 MULT=1
DX12_noxref VNB VPB NWDIODE A=8.742 P=13.12
*
.include "sky130_fd_sc_ls__nor4_2.pxi.spice"
*
.ends
*
*
