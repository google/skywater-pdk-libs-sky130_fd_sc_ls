* File: sky130_fd_sc_ls__o311ai_1.pex.spice
* Created: Fri Aug 28 13:51:51 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__O311AI_1%A1 3 5 7 8 12
r23 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.54
+ $Y=1.515 $X2=0.54 $Y2=1.515
r24 8 12 8.0403 $w=4.28e-07 $l=3e-07 $layer=LI1_cond $X=0.24 $Y=1.565 $X2=0.54
+ $Y2=1.565
r25 5 11 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=0.615 $Y=1.765
+ $X2=0.54 $Y2=1.515
r26 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.615 $Y=1.765
+ $X2=0.615 $Y2=2.4
r27 1 11 38.5562 $w=2.99e-07 $l=1.77059e-07 $layer=POLY_cond $X=0.565 $Y=1.35
+ $X2=0.54 $Y2=1.515
r28 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.565 $Y=1.35
+ $X2=0.565 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__O311AI_1%A2 3 5 7 8 9 10 11 18
r33 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.11
+ $Y=1.515 $X2=1.11 $Y2=1.515
r34 10 11 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.13 $Y=2.405
+ $X2=1.13 $Y2=2.775
r35 9 10 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.13 $Y=2.035
+ $X2=1.13 $Y2=2.405
r36 8 9 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.13 $Y=1.665 $X2=1.13
+ $Y2=2.035
r37 8 18 4.67207 $w=3.68e-07 $l=1.5e-07 $layer=LI1_cond $X=1.13 $Y=1.665
+ $X2=1.13 $Y2=1.515
r38 5 17 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=1.035 $Y=1.765
+ $X2=1.11 $Y2=1.515
r39 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.035 $Y=1.765
+ $X2=1.035 $Y2=2.4
r40 1 17 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=1.02 $Y=1.35
+ $X2=1.11 $Y2=1.515
r41 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.02 $Y=1.35 $X2=1.02
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__O311AI_1%A3 1 3 4 6 7
c28 7 0 4.01776e-20 $X=1.68 $Y=1.295
r29 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.68
+ $Y=1.385 $X2=1.68 $Y2=1.385
r30 7 11 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=1.68 $Y=1.295 $X2=1.68
+ $Y2=1.385
r31 4 10 38.9026 $w=2.7e-07 $l=2.05122e-07 $layer=POLY_cond $X=1.77 $Y=1.22
+ $X2=1.68 $Y2=1.385
r32 4 6 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.77 $Y=1.22 $X2=1.77
+ $Y2=0.74
r33 1 10 77.2841 $w=2.7e-07 $l=4.15812e-07 $layer=POLY_cond $X=1.605 $Y=1.765
+ $X2=1.68 $Y2=1.385
r34 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.605 $Y=1.765
+ $X2=1.605 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__O311AI_1%B1 1 3 4 6 7
c30 7 0 1.2348e-19 $X=2.16 $Y=1.295
c31 4 0 1.48672e-19 $X=2.27 $Y=1.22
r32 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.25
+ $Y=1.385 $X2=2.25 $Y2=1.385
r33 7 11 2.80324 $w=3.68e-07 $l=9e-08 $layer=LI1_cond $X=2.23 $Y=1.295 $X2=2.23
+ $Y2=1.385
r34 4 10 38.9026 $w=2.7e-07 $l=1.74714e-07 $layer=POLY_cond $X=2.27 $Y=1.22
+ $X2=2.25 $Y2=1.385
r35 4 6 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.27 $Y=1.22 $X2=2.27
+ $Y2=0.74
r36 1 10 77.2841 $w=2.7e-07 $l=4.15812e-07 $layer=POLY_cond $X=2.175 $Y=1.765
+ $X2=2.25 $Y2=1.385
r37 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.175 $Y=1.765
+ $X2=2.175 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__O311AI_1%C1 1 3 4 6 7
c23 1 0 2.8952e-19 $X=2.73 $Y=1.22
r24 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.09
+ $Y=1.385 $X2=3.09 $Y2=1.385
r25 7 11 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=3.09 $Y=1.295 $X2=3.09
+ $Y2=1.385
r26 4 10 64.1863 $w=4.34e-07 $l=4.73498e-07 $layer=POLY_cond $X=2.745 $Y=1.765
+ $X2=2.955 $Y2=1.385
r27 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.745 $Y=1.765
+ $X2=2.745 $Y2=2.4
r28 1 10 40.3085 $w=4.34e-07 $l=2.96226e-07 $layer=POLY_cond $X=2.73 $Y=1.22
+ $X2=2.955 $Y2=1.385
r29 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.73 $Y=1.22 $X2=2.73
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__O311AI_1%VPWR 1 2 7 9 15 20 21 22 32 33
r35 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r36 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r37 30 33 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r38 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r39 27 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r40 26 29 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.72 $Y=3.33
+ $X2=2.16 $Y2=3.33
r41 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r42 24 36 4.53571 $w=1.7e-07 $l=2.78e-07 $layer=LI1_cond $X=0.555 $Y=3.33
+ $X2=0.277 $Y2=3.33
r43 24 26 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=0.555 $Y=3.33
+ $X2=0.72 $Y2=3.33
r44 22 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r45 22 27 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r46 20 29 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.285 $Y=3.33
+ $X2=2.16 $Y2=3.33
r47 20 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.285 $Y=3.33
+ $X2=2.45 $Y2=3.33
r48 19 32 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=2.615 $Y=3.33
+ $X2=3.12 $Y2=3.33
r49 19 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.615 $Y=3.33
+ $X2=2.45 $Y2=3.33
r50 15 18 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=2.45 $Y=2.145
+ $X2=2.45 $Y2=2.825
r51 13 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.45 $Y=3.245
+ $X2=2.45 $Y2=3.33
r52 13 18 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=2.45 $Y=3.245
+ $X2=2.45 $Y2=2.825
r53 9 12 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=0.39 $Y=2.115 $X2=0.39
+ $Y2=2.815
r54 7 36 3.23047 $w=3.3e-07 $l=1.49579e-07 $layer=LI1_cond $X=0.39 $Y=3.245
+ $X2=0.277 $Y2=3.33
r55 7 12 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.39 $Y=3.245
+ $X2=0.39 $Y2=2.815
r56 2 18 400 $w=1.7e-07 $l=1.08038e-06 $layer=licon1_PDIFF $count=1 $X=2.25
+ $Y=1.84 $X2=2.45 $Y2=2.825
r57 2 15 400 $w=1.7e-07 $l=3.9246e-07 $layer=licon1_PDIFF $count=1 $X=2.25
+ $Y=1.84 $X2=2.45 $Y2=2.145
r58 1 12 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.245
+ $Y=1.84 $X2=0.39 $Y2=2.815
r59 1 9 400 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.245
+ $Y=1.84 $X2=0.39 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_LS__O311AI_1%Y 1 2 3 12 16 17 19 21 25 26 27 28 33
c48 19 0 1.08494e-19 $X=2.67 $Y=1.72
r49 28 41 1.07204 $w=4.28e-07 $l=4e-08 $layer=LI1_cond $X=3.02 $Y=2.775 $X2=3.02
+ $Y2=2.815
r50 27 28 9.91637 $w=4.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.02 $Y=2.405
+ $X2=3.02 $Y2=2.775
r51 26 27 9.91637 $w=4.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.02 $Y=2.035
+ $X2=3.02 $Y2=2.405
r52 26 33 1.34005 $w=4.28e-07 $l=5e-08 $layer=LI1_cond $X=3.02 $Y=2.035 $X2=3.02
+ $Y2=1.985
r53 24 33 2.54609 $w=4.28e-07 $l=9.5e-08 $layer=LI1_cond $X=3.02 $Y=1.89
+ $X2=3.02 $Y2=1.985
r54 24 25 3.14896 $w=3e-07 $l=1.46458e-07 $layer=LI1_cond $X=3.02 $Y=1.89
+ $X2=2.91 $Y2=1.805
r55 21 23 17.191 $w=5.23e-07 $l=4.95e-07 $layer=LI1_cond $X=2.847 $Y=0.515
+ $X2=2.847 $Y2=1.01
r56 19 25 3.14896 $w=3e-07 $l=2.79285e-07 $layer=LI1_cond $X=2.67 $Y=1.72
+ $X2=2.91 $Y2=1.805
r57 19 23 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=2.67 $Y=1.72
+ $X2=2.67 $Y2=1.01
r58 16 25 3.44808 $w=1.7e-07 $l=3.25e-07 $layer=LI1_cond $X=2.585 $Y=1.805
+ $X2=2.91 $Y2=1.805
r59 16 17 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=2.585 $Y=1.805
+ $X2=2.115 $Y2=1.805
r60 12 14 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=1.95 $Y=1.985
+ $X2=1.95 $Y2=2.815
r61 10 17 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.95 $Y=1.89
+ $X2=2.115 $Y2=1.805
r62 10 12 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=1.95 $Y=1.89
+ $X2=1.95 $Y2=1.985
r63 3 41 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.82
+ $Y=1.84 $X2=2.97 $Y2=2.815
r64 3 33 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.82
+ $Y=1.84 $X2=2.97 $Y2=1.985
r65 2 14 400 $w=1.7e-07 $l=1.10176e-06 $layer=licon1_PDIFF $count=1 $X=1.68
+ $Y=1.84 $X2=1.95 $Y2=2.815
r66 2 12 400 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_PDIFF $count=1 $X=1.68
+ $Y=1.84 $X2=1.95 $Y2=1.985
r67 1 21 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.805
+ $Y=0.37 $X2=2.945 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__O311AI_1%VGND 1 2 7 9 13 15 17 27 28 34
r35 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r36 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r37 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r38 24 27 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.68 $Y=0 $X2=3.12
+ $Y2=0
r39 22 34 12.0744 $w=1.7e-07 $l=2.8e-07 $layer=LI1_cond $X=1.675 $Y=0 $X2=1.395
+ $Y2=0
r40 22 24 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=1.675 $Y=0 $X2=1.68
+ $Y2=0
r41 21 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r42 21 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r43 20 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r44 18 31 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.222
+ $Y2=0
r45 18 20 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.72
+ $Y2=0
r46 17 34 12.0744 $w=1.7e-07 $l=2.8e-07 $layer=LI1_cond $X=1.115 $Y=0 $X2=1.395
+ $Y2=0
r47 17 20 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.115 $Y=0 $X2=0.72
+ $Y2=0
r48 15 28 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=0 $X2=3.12
+ $Y2=0
r49 15 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r50 15 24 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r51 11 34 2.35715 $w=5.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.395 $Y=0.085
+ $X2=1.395 $Y2=0
r52 11 13 9.18417 $w=5.58e-07 $l=4.3e-07 $layer=LI1_cond $X=1.395 $Y=0.085
+ $X2=1.395 $Y2=0.515
r53 7 31 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.222 $Y2=0
r54 7 9 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.28 $Y=0.085 $X2=0.28
+ $Y2=0.515
r55 2 13 182 $w=1.7e-07 $l=3.75566e-07 $layer=licon1_NDIFF $count=1 $X=1.095
+ $Y=0.37 $X2=1.405 $Y2=0.515
r56 1 9 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__O311AI_1%A_128_74# 1 2 9 11 12 13 15
c34 13 0 1.6604e-19 $X=2.055 $Y=0.84
r35 13 18 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.055 $Y=0.84
+ $X2=2.055 $Y2=0.925
r36 13 15 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=2.055 $Y=0.84
+ $X2=2.055 $Y2=0.495
r37 11 18 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.89 $Y=0.925
+ $X2=2.055 $Y2=0.925
r38 11 12 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=1.89 $Y=0.925
+ $X2=0.945 $Y2=0.925
r39 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.78 $Y=0.84
+ $X2=0.945 $Y2=0.925
r40 7 9 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=0.78 $Y=0.84 $X2=0.78
+ $Y2=0.515
r41 2 18 182 $w=1.7e-07 $l=6.51594e-07 $layer=licon1_NDIFF $count=1 $X=1.845
+ $Y=0.37 $X2=2.055 $Y2=0.925
r42 2 15 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=1.845
+ $Y=0.37 $X2=2.055 $Y2=0.495
r43 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.64
+ $Y=0.37 $X2=0.78 $Y2=0.515
.ends

