* File: sky130_fd_sc_ls__ebufn_4.spice
* Created: Fri Aug 28 13:22:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__ebufn_4.pex.spice"
.subckt sky130_fd_sc_ls__ebufn_4  VNB VPB A TE_B VPWR Z VGND
* 
* VGND	VGND
* Z	Z
* VPWR	VPWR
* TE_B	TE_B
* A	A
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_A_M1003_g N_A_27_368#_M1003_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1011 N_A_208_74#_M1011_d N_TE_B_M1011_g N_VGND_M1003_d VNB NSHORT L=0.15
+ W=0.74 AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1005 N_VGND_M1005_d N_A_208_74#_M1005_g N_A_378_74#_M1005_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.2072 PD=1.02 PS=2.04 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75003.2 A=0.111 P=1.78 MULT=1
MM1006 N_VGND_M1005_d N_A_208_74#_M1006_g N_A_378_74#_M1006_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75002.8 A=0.111 P=1.78 MULT=1
MM1010 N_VGND_M1010_d N_A_208_74#_M1010_g N_A_378_74#_M1006_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.1 SB=75002.4 A=0.111 P=1.78 MULT=1
MM1016 N_VGND_M1010_d N_A_208_74#_M1016_g N_A_378_74#_M1016_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.5 SB=75001.9 A=0.111 P=1.78 MULT=1
MM1004 N_A_378_74#_M1016_s N_A_27_368#_M1004_g N_Z_M1004_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.9 SB=75001.5 A=0.111 P=1.78 MULT=1
MM1013 N_A_378_74#_M1013_d N_A_27_368#_M1013_g N_Z_M1004_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75002.4 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1014 N_A_378_74#_M1013_d N_A_27_368#_M1014_g N_Z_M1014_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.111 PD=1.02 PS=1.04 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.8
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1018 N_A_378_74#_M1018_d N_A_27_368#_M1018_g N_Z_M1014_s VNB NSHORT L=0.15
+ W=0.74 AD=0.2035 AS=0.111 PD=2.03 PS=1.04 NRD=0 NRS=3.24 M=1 R=4.93333
+ SA=75003.2 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1015 N_VPWR_M1015_d N_A_M1015_g N_A_27_368#_M1015_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.182 AS=0.3304 PD=1.445 PS=2.83 NRD=3.5066 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1000 N_A_208_74#_M1000_d N_TE_B_M1000_g N_VPWR_M1015_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.3304 AS=0.182 PD=2.83 PS=1.445 NRD=1.7533 NRS=4.3931 M=1 R=7.46667
+ SA=75000.7 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1001 N_A_348_368#_M1001_d N_TE_B_M1001_g N_VPWR_M1001_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75003.4 A=0.168 P=2.54 MULT=1
MM1007 N_A_348_368#_M1007_d N_TE_B_M1007_g N_VPWR_M1001_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75002.9 A=0.168 P=2.54 MULT=1
MM1009 N_A_348_368#_M1007_d N_TE_B_M1009_g N_VPWR_M1009_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75002.5 A=0.168 P=2.54 MULT=1
MM1012 N_A_348_368#_M1012_d N_TE_B_M1012_g N_VPWR_M1009_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.6 SB=75002 A=0.168 P=2.54 MULT=1
MM1002 N_Z_M1002_d N_A_27_368#_M1002_g N_A_348_368#_M1012_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1008 N_Z_M1002_d N_A_27_368#_M1008_g N_A_348_368#_M1008_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.5 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1017 N_Z_M1017_d N_A_27_368#_M1017_g N_A_348_368#_M1008_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.9 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1019 N_Z_M1017_d N_A_27_368#_M1019_g N_A_348_368#_M1019_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.3248 PD=1.42 PS=2.82 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75003.4 SB=75000.2 A=0.168 P=2.54 MULT=1
DX20_noxref VNB VPB NWDIODE A=11.4204 P=16
*
.include "sky130_fd_sc_ls__ebufn_4.pxi.spice"
*
.ends
*
*
