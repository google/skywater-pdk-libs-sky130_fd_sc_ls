* NGSPICE file created from sky130_fd_sc_ls__nor3b_2.ext - technology: sky130A

.subckt sky130_fd_sc_ls__nor3b_2 A B C_N VGND VNB VPB VPWR Y
M1000 VGND a_27_392# Y VNB nshort w=740000u l=150000u
+  ad=1.6739e+12p pd=1.049e+07u as=6.697e+11p ps=6.25e+06u
M1001 a_227_368# a_27_392# Y VPB phighvt w=1.12e+06u l=150000u
+  ad=9.856e+11p pd=8.48e+06u as=3.36e+11p ps=2.84e+06u
M1002 Y B VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPWR A a_495_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=9.396e+11p pd=8.22e+06u as=6.72e+11p ps=5.68e+06u
M1004 Y A VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND A Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_495_368# B a_227_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND C_N a_27_392# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1008 a_227_368# B a_495_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y a_27_392# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND B Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR C_N a_27_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1012 Y a_27_392# a_227_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_495_368# A VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

