* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__or4_4 A B C D VGND VNB VPB VPWR X
M1000 VGND a_83_264# X VNB nshort w=740000u l=150000u
+  ad=2.2402e+12p pd=1.413e+07u as=6.549e+11p ps=4.73e+06u
M1001 VPWR a_83_264# X VPB phighvt w=1.12e+06u l=150000u
+  ad=1.2968e+12p pd=1.11e+07u as=6.72e+11p ps=5.68e+06u
M1002 a_962_392# D a_83_264# VPB phighvt w=1e+06u l=150000u
+  ad=6.5e+11p pd=5.3e+06u as=3e+11p ps=2.6e+06u
M1003 a_83_264# B VGND VNB nshort w=740000u l=150000u
+  ad=4.662e+11p pd=4.22e+06u as=0p ps=0u
M1004 X a_83_264# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND D a_83_264# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_499_392# C a_962_392# VPB phighvt w=1e+06u l=150000u
+  ad=9.9e+11p pd=7.98e+06u as=0p ps=0u
M1007 X a_83_264# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND a_83_264# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_588_392# B a_499_392# VPB phighvt w=1e+06u l=150000u
+  ad=6.2e+11p pd=5.24e+06u as=0p ps=0u
M1010 VGND A a_83_264# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 X a_83_264# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR a_83_264# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_83_264# C VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_499_392# B a_588_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR A a_588_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 X a_83_264# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_962_392# C a_499_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_588_392# A VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_83_264# D a_962_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
