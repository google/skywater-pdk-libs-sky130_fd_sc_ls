* File: sky130_fd_sc_ls__a31oi_4.pex.spice
* Created: Fri Aug 28 12:59:40 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__A31OI_4%A3 1 3 6 10 12 14 17 19 21 22 24 27 29 30 31
+ 46 47
c80 27 0 1.69199e-19 $X=1.87 $Y=0.74
r81 47 48 1.95405 $w=3.7e-07 $l=1.5e-08 $layer=POLY_cond $X=1.855 $Y=1.557
+ $X2=1.87 $Y2=1.557
r82 45 47 30.6135 $w=3.7e-07 $l=2.35e-07 $layer=POLY_cond $X=1.62 $Y=1.557
+ $X2=1.855 $Y2=1.557
r83 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.62
+ $Y=1.515 $X2=1.62 $Y2=1.515
r84 43 45 28.0081 $w=3.7e-07 $l=2.15e-07 $layer=POLY_cond $X=1.405 $Y=1.557
+ $X2=1.62 $Y2=1.557
r85 42 43 4.55946 $w=3.7e-07 $l=3.5e-08 $layer=POLY_cond $X=1.37 $Y=1.557
+ $X2=1.405 $Y2=1.557
r86 41 42 54.0622 $w=3.7e-07 $l=4.15e-07 $layer=POLY_cond $X=0.955 $Y=1.557
+ $X2=1.37 $Y2=1.557
r87 40 41 1.95405 $w=3.7e-07 $l=1.5e-08 $layer=POLY_cond $X=0.94 $Y=1.557
+ $X2=0.955 $Y2=1.557
r88 38 40 44.2919 $w=3.7e-07 $l=3.4e-07 $layer=POLY_cond $X=0.6 $Y=1.557
+ $X2=0.94 $Y2=1.557
r89 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.6
+ $Y=1.515 $X2=0.6 $Y2=1.515
r90 36 38 11.7243 $w=3.7e-07 $l=9e-08 $layer=POLY_cond $X=0.51 $Y=1.557 $X2=0.6
+ $Y2=1.557
r91 35 36 0.651351 $w=3.7e-07 $l=5e-09 $layer=POLY_cond $X=0.505 $Y=1.557
+ $X2=0.51 $Y2=1.557
r92 31 46 11.2564 $w=4.28e-07 $l=4.2e-07 $layer=LI1_cond $X=1.2 $Y=1.565
+ $X2=1.62 $Y2=1.565
r93 30 31 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=1.2 $Y2=1.565
r94 30 39 3.21612 $w=4.28e-07 $l=1.2e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=0.6 $Y2=1.565
r95 29 39 9.64836 $w=4.28e-07 $l=3.6e-07 $layer=LI1_cond $X=0.24 $Y=1.565
+ $X2=0.6 $Y2=1.565
r96 25 48 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.87 $Y=1.35
+ $X2=1.87 $Y2=1.557
r97 25 27 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.87 $Y=1.35
+ $X2=1.87 $Y2=0.74
r98 22 47 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.855 $Y=1.765
+ $X2=1.855 $Y2=1.557
r99 22 24 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.855 $Y=1.765
+ $X2=1.855 $Y2=2.4
r100 19 43 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.405 $Y=1.765
+ $X2=1.405 $Y2=1.557
r101 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.405 $Y=1.765
+ $X2=1.405 $Y2=2.4
r102 15 42 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.37 $Y=1.35
+ $X2=1.37 $Y2=1.557
r103 15 17 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.37 $Y=1.35
+ $X2=1.37 $Y2=0.74
r104 12 41 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.955 $Y=1.765
+ $X2=0.955 $Y2=1.557
r105 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.955 $Y=1.765
+ $X2=0.955 $Y2=2.4
r106 8 40 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.94 $Y=1.35
+ $X2=0.94 $Y2=1.557
r107 8 10 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.94 $Y=1.35
+ $X2=0.94 $Y2=0.74
r108 4 36 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.51 $Y=1.35
+ $X2=0.51 $Y2=1.557
r109 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.51 $Y=1.35 $X2=0.51
+ $Y2=0.74
r110 1 35 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=1.557
r111 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__A31OI_4%A2 3 5 7 10 12 14 17 19 21 24 26 28 29 30 31
+ 32 49
c90 32 0 1.0093e-20 $X=4.08 $Y=1.665
c91 26 0 9.21447e-20 $X=3.755 $Y=1.765
r92 49 50 1.98626 $w=3.64e-07 $l=1.5e-08 $layer=POLY_cond $X=3.74 $Y=1.557
+ $X2=3.755 $Y2=1.557
r93 47 49 23.8352 $w=3.64e-07 $l=1.8e-07 $layer=POLY_cond $X=3.56 $Y=1.557
+ $X2=3.74 $Y2=1.557
r94 47 48 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.56
+ $Y=1.515 $X2=3.56 $Y2=1.515
r95 45 47 40.3874 $w=3.64e-07 $l=3.05e-07 $layer=POLY_cond $X=3.255 $Y=1.557
+ $X2=3.56 $Y2=1.557
r96 44 45 11.2555 $w=3.64e-07 $l=8.5e-08 $layer=POLY_cond $X=3.17 $Y=1.557
+ $X2=3.255 $Y2=1.557
r97 43 44 48.3324 $w=3.64e-07 $l=3.65e-07 $layer=POLY_cond $X=2.805 $Y=1.557
+ $X2=3.17 $Y2=1.557
r98 42 43 8.60714 $w=3.64e-07 $l=6.5e-08 $layer=POLY_cond $X=2.74 $Y=1.557
+ $X2=2.805 $Y2=1.557
r99 40 42 26.4835 $w=3.64e-07 $l=2e-07 $layer=POLY_cond $X=2.54 $Y=1.557
+ $X2=2.74 $Y2=1.557
r100 40 41 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.54
+ $Y=1.515 $X2=2.54 $Y2=1.515
r101 38 40 31.1181 $w=3.64e-07 $l=2.35e-07 $layer=POLY_cond $X=2.305 $Y=1.557
+ $X2=2.54 $Y2=1.557
r102 37 38 0.662088 $w=3.64e-07 $l=5e-09 $layer=POLY_cond $X=2.3 $Y=1.557
+ $X2=2.305 $Y2=1.557
r103 31 32 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=3.6 $Y=1.565
+ $X2=4.08 $Y2=1.565
r104 31 48 1.07204 $w=4.28e-07 $l=4e-08 $layer=LI1_cond $X=3.6 $Y=1.565 $X2=3.56
+ $Y2=1.565
r105 30 48 11.7924 $w=4.28e-07 $l=4.4e-07 $layer=LI1_cond $X=3.12 $Y=1.565
+ $X2=3.56 $Y2=1.565
r106 29 30 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=2.64 $Y=1.565
+ $X2=3.12 $Y2=1.565
r107 29 41 2.6801 $w=4.28e-07 $l=1e-07 $layer=LI1_cond $X=2.64 $Y=1.565 $X2=2.54
+ $Y2=1.565
r108 26 50 23.572 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.755 $Y=1.765
+ $X2=3.755 $Y2=1.557
r109 26 28 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.755 $Y=1.765
+ $X2=3.755 $Y2=2.4
r110 22 49 23.572 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.74 $Y=1.35
+ $X2=3.74 $Y2=1.557
r111 22 24 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.74 $Y=1.35
+ $X2=3.74 $Y2=0.74
r112 19 45 23.572 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.255 $Y=1.765
+ $X2=3.255 $Y2=1.557
r113 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.255 $Y=1.765
+ $X2=3.255 $Y2=2.4
r114 15 44 23.572 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.17 $Y=1.35
+ $X2=3.17 $Y2=1.557
r115 15 17 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.17 $Y=1.35
+ $X2=3.17 $Y2=0.74
r116 12 43 23.572 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.805 $Y=1.765
+ $X2=2.805 $Y2=1.557
r117 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.805 $Y=1.765
+ $X2=2.805 $Y2=2.4
r118 8 42 23.572 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.74 $Y=1.35
+ $X2=2.74 $Y2=1.557
r119 8 10 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.74 $Y=1.35
+ $X2=2.74 $Y2=0.74
r120 5 38 23.572 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.305 $Y=1.765
+ $X2=2.305 $Y2=1.557
r121 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.305 $Y=1.765
+ $X2=2.305 $Y2=2.4
r122 1 37 23.572 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.3 $Y=1.35 $X2=2.3
+ $Y2=1.557
r123 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.3 $Y=1.35 $X2=2.3
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__A31OI_4%A1 1 3 4 5 8 10 12 13 17 19 21 24 26 28 31
+ 33 34 35 36 49
c109 36 0 1.82133e-19 $X=6 $Y=1.665
c110 26 0 1.55065e-19 $X=6.285 $Y=1.765
c111 10 0 1.41876e-19 $X=4.755 $Y=1.765
r112 48 49 42.3378 $w=3.7e-07 $l=3.25e-07 $layer=POLY_cond $X=5.96 $Y=1.542
+ $X2=6.285 $Y2=1.542
r113 46 48 11.7243 $w=3.7e-07 $l=9e-08 $layer=POLY_cond $X=5.87 $Y=1.542
+ $X2=5.96 $Y2=1.542
r114 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.87
+ $Y=1.515 $X2=5.87 $Y2=1.515
r115 44 46 17.5865 $w=3.7e-07 $l=1.35e-07 $layer=POLY_cond $X=5.735 $Y=1.542
+ $X2=5.87 $Y2=1.542
r116 43 47 9.11234 $w=4.28e-07 $l=3.4e-07 $layer=LI1_cond $X=5.53 $Y=1.565
+ $X2=5.87 $Y2=1.565
r117 42 44 26.7054 $w=3.7e-07 $l=2.05e-07 $layer=POLY_cond $X=5.53 $Y=1.542
+ $X2=5.735 $Y2=1.542
r118 42 43 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.53
+ $Y=1.515 $X2=5.53 $Y2=1.515
r119 40 42 9.11892 $w=3.7e-07 $l=7e-08 $layer=POLY_cond $X=5.46 $Y=1.542
+ $X2=5.53 $Y2=1.542
r120 36 47 3.48413 $w=4.28e-07 $l=1.3e-07 $layer=LI1_cond $X=6 $Y=1.565 $X2=5.87
+ $Y2=1.565
r121 35 43 0.26801 $w=4.28e-07 $l=1e-08 $layer=LI1_cond $X=5.52 $Y=1.565
+ $X2=5.53 $Y2=1.565
r122 34 35 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=5.04 $Y=1.565
+ $X2=5.52 $Y2=1.565
r123 29 49 13.6784 $w=3.7e-07 $l=2.69433e-07 $layer=POLY_cond $X=6.39 $Y=1.32
+ $X2=6.285 $Y2=1.542
r124 29 31 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.39 $Y=1.32
+ $X2=6.39 $Y2=0.74
r125 26 49 23.9667 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=6.285 $Y=1.765
+ $X2=6.285 $Y2=1.542
r126 26 28 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.285 $Y=1.765
+ $X2=6.285 $Y2=2.4
r127 22 48 23.9667 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=5.96 $Y=1.32
+ $X2=5.96 $Y2=1.542
r128 22 24 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=5.96 $Y=1.32
+ $X2=5.96 $Y2=0.74
r129 19 44 23.9667 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=5.735 $Y=1.765
+ $X2=5.735 $Y2=1.542
r130 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.735 $Y=1.765
+ $X2=5.735 $Y2=2.4
r131 15 40 23.9667 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=5.46 $Y=1.32
+ $X2=5.46 $Y2=1.542
r132 15 17 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=5.46 $Y=1.32
+ $X2=5.46 $Y2=0.74
r133 14 33 6.33988 $w=3.6e-07 $l=1.08995e-07 $layer=POLY_cond $X=4.845 $Y=1.5
+ $X2=4.755 $Y2=1.542
r134 13 40 9.77027 $w=3.7e-07 $l=9.3675e-08 $layer=POLY_cond $X=5.385 $Y=1.5
+ $X2=5.46 $Y2=1.542
r135 13 14 86.5563 $w=3.6e-07 $l=5.4e-07 $layer=POLY_cond $X=5.385 $Y=1.5
+ $X2=4.845 $Y2=1.5
r136 10 33 18.972 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=4.755 $Y=1.765
+ $X2=4.755 $Y2=1.542
r137 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.755 $Y=1.765
+ $X2=4.755 $Y2=2.4
r138 6 33 18.972 $w=1.5e-07 $l=2.29377e-07 $layer=POLY_cond $X=4.74 $Y=1.32
+ $X2=4.755 $Y2=1.542
r139 6 8 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=4.74 $Y=1.32 $X2=4.74
+ $Y2=0.74
r140 4 33 6.33988 $w=1.5e-07 $l=1.87681e-07 $layer=POLY_cond $X=4.665 $Y=1.69
+ $X2=4.755 $Y2=1.542
r141 4 5 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=4.665 $Y=1.69
+ $X2=4.33 $Y2=1.69
r142 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.255 $Y=1.765
+ $X2=4.33 $Y2=1.69
r143 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.255 $Y=1.765
+ $X2=4.255 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__A31OI_4%B1 1 3 6 8 10 11 13 14 16 19 21 22 23 24 25
+ 41
c60 41 0 1.82133e-19 $X=8.135 $Y=1.557
c61 25 0 1.55065e-19 $X=8.4 $Y=1.665
c62 6 0 1.25471e-19 $X=6.89 $Y=0.74
r63 41 42 1.30978 $w=3.68e-07 $l=1e-08 $layer=POLY_cond $X=8.135 $Y=1.557
+ $X2=8.145 $Y2=1.557
r64 40 41 58.9402 $w=3.68e-07 $l=4.5e-07 $layer=POLY_cond $X=7.685 $Y=1.557
+ $X2=8.135 $Y2=1.557
r65 38 40 21.6114 $w=3.68e-07 $l=1.65e-07 $layer=POLY_cond $X=7.52 $Y=1.557
+ $X2=7.685 $Y2=1.557
r66 38 39 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=7.52
+ $Y=1.515 $X2=7.52 $Y2=1.515
r67 36 38 37.3288 $w=3.68e-07 $l=2.85e-07 $layer=POLY_cond $X=7.235 $Y=1.557
+ $X2=7.52 $Y2=1.557
r68 35 36 45.1875 $w=3.68e-07 $l=3.45e-07 $layer=POLY_cond $X=6.89 $Y=1.557
+ $X2=7.235 $Y2=1.557
r69 33 35 6.54891 $w=3.68e-07 $l=5e-08 $layer=POLY_cond $X=6.84 $Y=1.557
+ $X2=6.89 $Y2=1.557
r70 33 34 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=6.84
+ $Y=1.515 $X2=6.84 $Y2=1.515
r71 31 33 9.82337 $w=3.68e-07 $l=7.5e-08 $layer=POLY_cond $X=6.765 $Y=1.557
+ $X2=6.84 $Y2=1.557
r72 24 25 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=7.92 $Y=1.565
+ $X2=8.4 $Y2=1.565
r73 24 39 10.7204 $w=4.28e-07 $l=4e-07 $layer=LI1_cond $X=7.92 $Y=1.565 $X2=7.52
+ $Y2=1.565
r74 23 39 2.14408 $w=4.28e-07 $l=8e-08 $layer=LI1_cond $X=7.44 $Y=1.565 $X2=7.52
+ $Y2=1.565
r75 22 23 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=6.96 $Y=1.565
+ $X2=7.44 $Y2=1.565
r76 22 34 3.21612 $w=4.28e-07 $l=1.2e-07 $layer=LI1_cond $X=6.96 $Y=1.565
+ $X2=6.84 $Y2=1.565
r77 21 34 9.64836 $w=4.28e-07 $l=3.6e-07 $layer=LI1_cond $X=6.48 $Y=1.565
+ $X2=6.84 $Y2=1.565
r78 17 42 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=8.145 $Y=1.35
+ $X2=8.145 $Y2=1.557
r79 17 19 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=8.145 $Y=1.35
+ $X2=8.145 $Y2=0.74
r80 14 41 23.8357 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=8.135 $Y=1.765
+ $X2=8.135 $Y2=1.557
r81 14 16 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.135 $Y=1.765
+ $X2=8.135 $Y2=2.4
r82 11 40 23.8357 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=7.685 $Y=1.765
+ $X2=7.685 $Y2=1.557
r83 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.685 $Y=1.765
+ $X2=7.685 $Y2=2.4
r84 8 36 23.8357 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=7.235 $Y=1.765
+ $X2=7.235 $Y2=1.557
r85 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.235 $Y=1.765
+ $X2=7.235 $Y2=2.4
r86 4 35 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.89 $Y=1.35
+ $X2=6.89 $Y2=1.557
r87 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.89 $Y=1.35 $X2=6.89
+ $Y2=0.74
r88 1 31 23.8357 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=6.765 $Y=1.765
+ $X2=6.765 $Y2=1.557
r89 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.765 $Y=1.765
+ $X2=6.765 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__A31OI_4%A_27_368# 1 2 3 4 5 6 7 8 9 28 30 32 36 38
+ 40 42 44 48 50 52 53 58 60 61 62 63 66 68 72 79 85 89 92 93 96
c120 85 0 9.21447e-20 $X=3.03 $Y=2.035
c121 52 0 1.31783e-19 $X=4.03 $Y=2.12
c122 40 0 1.06564e-19 $X=2.08 $Y=2.15
r123 91 93 10.4169 $w=6.38e-07 $l=1.65e-07 $layer=LI1_cond $X=5.51 $Y=2.61
+ $X2=5.675 $Y2=2.61
r124 91 92 19.3874 $w=6.38e-07 $l=6.45e-07 $layer=LI1_cond $X=5.51 $Y=2.61
+ $X2=4.865 $Y2=2.61
r125 82 83 0.563077 $w=3.25e-07 $l=1.5e-08 $layer=LI1_cond $X=2.08 $Y=2.035
+ $X2=2.08 $Y2=2.05
r126 81 82 2.62769 $w=3.25e-07 $l=7e-08 $layer=LI1_cond $X=2.08 $Y=1.965
+ $X2=2.08 $Y2=2.035
r127 72 75 29.8782 $w=2.68e-07 $l=7e-07 $layer=LI1_cond $X=8.39 $Y=2.115
+ $X2=8.39 $Y2=2.815
r128 70 75 3.84148 $w=2.68e-07 $l=9e-08 $layer=LI1_cond $X=8.39 $Y=2.905
+ $X2=8.39 $Y2=2.815
r129 69 96 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=7.575 $Y=2.99
+ $X2=7.475 $Y2=2.99
r130 68 70 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=8.255 $Y=2.99
+ $X2=8.39 $Y2=2.905
r131 68 69 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=8.255 $Y=2.99
+ $X2=7.575 $Y2=2.99
r132 64 96 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=7.475 $Y=2.905
+ $X2=7.475 $Y2=2.99
r133 64 66 24.9545 $w=1.98e-07 $l=4.5e-07 $layer=LI1_cond $X=7.475 $Y=2.905
+ $X2=7.475 $Y2=2.455
r134 62 96 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=7.375 $Y=2.99
+ $X2=7.475 $Y2=2.99
r135 62 63 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=7.375 $Y=2.99
+ $X2=6.675 $Y2=2.99
r136 61 63 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.51 $Y=2.905
+ $X2=6.675 $Y2=2.99
r137 60 95 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.51 $Y=2.46 $X2=6.51
+ $Y2=2.375
r138 60 61 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=6.51 $Y=2.46
+ $X2=6.51 $Y2=2.905
r139 58 95 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.345 $Y=2.375
+ $X2=6.51 $Y2=2.375
r140 58 93 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.345 $Y=2.375
+ $X2=5.675 $Y2=2.375
r141 57 89 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.195 $Y=2.375
+ $X2=4.03 $Y2=2.375
r142 57 92 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.195 $Y=2.375
+ $X2=4.865 $Y2=2.375
r143 53 89 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.03 $Y=2.29
+ $X2=4.03 $Y2=2.375
r144 52 87 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.03 $Y=2.12 $X2=4.03
+ $Y2=2.035
r145 52 53 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=4.03 $Y=2.12
+ $X2=4.03 $Y2=2.29
r146 51 85 8.10876 $w=1.85e-07 $l=1.72337e-07 $layer=LI1_cond $X=3.195 $Y=2.035
+ $X2=3.03 $Y2=2.05
r147 50 87 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.865 $Y=2.035
+ $X2=4.03 $Y2=2.035
r148 50 51 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.865 $Y=2.035
+ $X2=3.195 $Y2=2.035
r149 46 85 0.63164 $w=3.3e-07 $l=1e-07 $layer=LI1_cond $X=3.03 $Y=2.15 $X2=3.03
+ $Y2=2.05
r150 46 48 23.2235 $w=3.28e-07 $l=6.65e-07 $layer=LI1_cond $X=3.03 $Y=2.15
+ $X2=3.03 $Y2=2.815
r151 45 83 3.57764 $w=2e-07 $l=1.65e-07 $layer=LI1_cond $X=2.245 $Y=2.05
+ $X2=2.08 $Y2=2.05
r152 44 85 8.10876 $w=1.85e-07 $l=1.65e-07 $layer=LI1_cond $X=2.865 $Y=2.05
+ $X2=3.03 $Y2=2.05
r153 44 45 34.3818 $w=1.98e-07 $l=6.2e-07 $layer=LI1_cond $X=2.865 $Y=2.05
+ $X2=2.245 $Y2=2.05
r154 40 83 4.8124 $w=3.25e-07 $l=1e-07 $layer=LI1_cond $X=2.08 $Y=2.15 $X2=2.08
+ $Y2=2.05
r155 40 42 10.7728 $w=2.28e-07 $l=2.15e-07 $layer=LI1_cond $X=2.08 $Y=2.15
+ $X2=2.08 $Y2=2.365
r156 39 79 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=1.295 $Y=2.035
+ $X2=1.18 $Y2=2.035
r157 38 82 4.53325 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.915 $Y=2.035
+ $X2=2.08 $Y2=2.035
r158 38 39 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=1.915 $Y=2.035
+ $X2=1.295 $Y2=2.035
r159 34 79 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.18 $Y=2.12
+ $X2=1.18 $Y2=2.035
r160 34 36 14.0297 $w=2.28e-07 $l=2.8e-07 $layer=LI1_cond $X=1.18 $Y=2.12
+ $X2=1.18 $Y2=2.4
r161 33 77 4.57959 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=0.395 $Y=2.035
+ $X2=0.255 $Y2=2.035
r162 32 79 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=1.065 $Y=2.035
+ $X2=1.18 $Y2=2.035
r163 32 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.065 $Y=2.035
+ $X2=0.395 $Y2=2.035
r164 28 77 2.78046 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.255 $Y=2.12
+ $X2=0.255 $Y2=2.035
r165 28 30 12.965 $w=2.78e-07 $l=3.15e-07 $layer=LI1_cond $X=0.255 $Y=2.12
+ $X2=0.255 $Y2=2.435
r166 9 75 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=8.21
+ $Y=1.84 $X2=8.36 $Y2=2.815
r167 9 72 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=8.21
+ $Y=1.84 $X2=8.36 $Y2=2.115
r168 8 66 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=7.31
+ $Y=1.84 $X2=7.46 $Y2=2.455
r169 7 95 300 $w=1.7e-07 $l=6.05372e-07 $layer=licon1_PDIFF $count=2 $X=6.36
+ $Y=1.84 $X2=6.51 $Y2=2.375
r170 6 91 150 $w=1.7e-07 $l=9.08955e-07 $layer=licon1_PDIFF $count=4 $X=4.83
+ $Y=1.84 $X2=5.51 $Y2=2.375
r171 5 89 300 $w=1.7e-07 $l=6.9282e-07 $layer=licon1_PDIFF $count=2 $X=3.83
+ $Y=1.84 $X2=4.03 $Y2=2.44
r172 5 87 600 $w=1.7e-07 $l=2.81069e-07 $layer=licon1_PDIFF $count=1 $X=3.83
+ $Y=1.84 $X2=4.03 $Y2=2.035
r173 4 85 400 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=2.88
+ $Y=1.84 $X2=3.03 $Y2=2.035
r174 4 48 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.88
+ $Y=1.84 $X2=3.03 $Y2=2.815
r175 3 81 600 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_PDIFF $count=1 $X=1.93
+ $Y=1.84 $X2=2.08 $Y2=1.965
r176 3 42 300 $w=1.7e-07 $l=5.95294e-07 $layer=licon1_PDIFF $count=2 $X=1.93
+ $Y=1.84 $X2=2.08 $Y2=2.365
r177 2 79 600 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=1.03
+ $Y=1.84 $X2=1.18 $Y2=2.035
r178 2 36 300 $w=1.7e-07 $l=6.30555e-07 $layer=licon1_PDIFF $count=2 $X=1.03
+ $Y=1.84 $X2=1.18 $Y2=2.4
r179 1 77 600 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.035
r180 1 30 300 $w=1.7e-07 $l=6.63551e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.435
.ends

.subckt PM_SKY130_FD_SC_LS__A31OI_4%VPWR 1 2 3 4 5 6 21 25 29 33 37 41 44 45 46
+ 48 53 62 66 71 81 82 85 88 91 94 97
r111 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r112 94 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r113 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r114 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r115 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r116 81 82 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r117 79 82 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=8.4 $Y2=3.33
r118 79 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33 $X2=6
+ $Y2=3.33
r119 78 81 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=6.48 $Y=3.33
+ $X2=8.4 $Y2=3.33
r120 78 79 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r121 76 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.175 $Y=3.33
+ $X2=6.01 $Y2=3.33
r122 76 78 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=6.175 $Y=3.33
+ $X2=6.48 $Y2=3.33
r123 75 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33 $X2=6
+ $Y2=3.33
r124 75 95 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=4.56 $Y2=3.33
r125 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r126 72 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.695 $Y=3.33
+ $X2=4.53 $Y2=3.33
r127 72 74 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=4.695 $Y=3.33
+ $X2=5.52 $Y2=3.33
r128 71 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.845 $Y=3.33
+ $X2=6.01 $Y2=3.33
r129 71 74 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=5.845 $Y=3.33
+ $X2=5.52 $Y2=3.33
r130 70 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r131 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r132 67 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.695 $Y=3.33
+ $X2=3.53 $Y2=3.33
r133 67 69 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=3.695 $Y=3.33
+ $X2=4.08 $Y2=3.33
r134 66 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.365 $Y=3.33
+ $X2=4.53 $Y2=3.33
r135 66 69 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=4.365 $Y=3.33
+ $X2=4.08 $Y2=3.33
r136 65 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r137 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r138 62 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.365 $Y=3.33
+ $X2=3.53 $Y2=3.33
r139 62 64 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=3.365 $Y=3.33
+ $X2=3.12 $Y2=3.33
r140 61 65 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r141 61 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r142 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r143 58 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.795 $Y=3.33
+ $X2=1.63 $Y2=3.33
r144 58 60 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.795 $Y=3.33
+ $X2=2.16 $Y2=3.33
r145 57 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r146 57 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r147 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r148 54 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=0.73 $Y2=3.33
r149 54 56 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=1.2 $Y2=3.33
r150 53 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.465 $Y=3.33
+ $X2=1.63 $Y2=3.33
r151 53 56 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.465 $Y=3.33
+ $X2=1.2 $Y2=3.33
r152 51 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r153 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r154 48 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.73 $Y2=3.33
r155 48 50 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.24 $Y2=3.33
r156 46 95 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=3.33
+ $X2=4.56 $Y2=3.33
r157 46 70 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=3.33
+ $X2=4.08 $Y2=3.33
r158 44 60 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=2.365 $Y=3.33
+ $X2=2.16 $Y2=3.33
r159 44 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.365 $Y=3.33
+ $X2=2.53 $Y2=3.33
r160 43 64 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=2.695 $Y=3.33
+ $X2=3.12 $Y2=3.33
r161 43 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.695 $Y=3.33
+ $X2=2.53 $Y2=3.33
r162 39 97 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.01 $Y=3.245
+ $X2=6.01 $Y2=3.33
r163 39 41 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=6.01 $Y=3.245
+ $X2=6.01 $Y2=2.765
r164 35 94 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.53 $Y=3.245
+ $X2=4.53 $Y2=3.33
r165 35 37 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=4.53 $Y=3.245
+ $X2=4.53 $Y2=2.765
r166 31 91 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.53 $Y=3.245
+ $X2=3.53 $Y2=3.33
r167 31 33 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=3.53 $Y=3.245
+ $X2=3.53 $Y2=2.375
r168 27 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.53 $Y=3.245
+ $X2=2.53 $Y2=3.33
r169 27 29 29.3349 $w=3.28e-07 $l=8.4e-07 $layer=LI1_cond $X=2.53 $Y=3.245
+ $X2=2.53 $Y2=2.405
r170 23 88 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.63 $Y=3.245
+ $X2=1.63 $Y2=3.33
r171 23 25 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=1.63 $Y=3.245
+ $X2=1.63 $Y2=2.375
r172 19 85 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=3.33
r173 19 21 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=2.375
r174 6 41 600 $w=1.7e-07 $l=1.02011e-06 $layer=licon1_PDIFF $count=1 $X=5.81
+ $Y=1.84 $X2=6.01 $Y2=2.765
r175 5 37 600 $w=1.7e-07 $l=1.02011e-06 $layer=licon1_PDIFF $count=1 $X=4.33
+ $Y=1.84 $X2=4.53 $Y2=2.765
r176 4 33 300 $w=1.7e-07 $l=6.27077e-07 $layer=licon1_PDIFF $count=2 $X=3.33
+ $Y=1.84 $X2=3.53 $Y2=2.375
r177 3 29 300 $w=1.7e-07 $l=6.3559e-07 $layer=licon1_PDIFF $count=2 $X=2.38
+ $Y=1.84 $X2=2.53 $Y2=2.405
r178 2 25 300 $w=1.7e-07 $l=6.05372e-07 $layer=licon1_PDIFF $count=2 $X=1.48
+ $Y=1.84 $X2=1.63 $Y2=2.375
r179 1 21 300 $w=1.7e-07 $l=6.05372e-07 $layer=licon1_PDIFF $count=2 $X=0.58
+ $Y=1.84 $X2=0.73 $Y2=2.375
.ends

.subckt PM_SKY130_FD_SC_LS__A31OI_4%Y 1 2 3 4 5 6 19 21 22 25 27 31 33 37 43 45
+ 49 50 52 54 55 56
r111 55 56 17.4042 $w=2.43e-07 $l=3.7e-07 $layer=LI1_cond $X=4.567 $Y=1.295
+ $X2=4.567 $Y2=1.665
r112 48 56 13.406 $w=2.43e-07 $l=2.85e-07 $layer=LI1_cond $X=4.567 $Y=1.95
+ $X2=4.567 $Y2=1.665
r113 45 55 5.40943 $w=2.43e-07 $l=1.15e-07 $layer=LI1_cond $X=4.567 $Y=1.18
+ $X2=4.567 $Y2=1.295
r114 45 47 3.32808 $w=2.45e-07 $l=2.27288e-07 $layer=LI1_cond $X=4.567 $Y=1.18
+ $X2=4.52 $Y2=0.975
r115 41 43 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=8.36 $Y=1.01
+ $X2=8.36 $Y2=0.515
r116 38 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.175 $Y=2.035
+ $X2=7.01 $Y2=2.035
r117 37 54 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.745 $Y=2.035
+ $X2=7.91 $Y2=2.035
r118 37 38 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=7.745 $Y=2.035
+ $X2=7.175 $Y2=2.035
r119 34 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.84 $Y=1.095
+ $X2=6.675 $Y2=1.095
r120 33 41 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.195 $Y=1.095
+ $X2=8.36 $Y2=1.01
r121 33 34 88.4011 $w=1.68e-07 $l=1.355e-06 $layer=LI1_cond $X=8.195 $Y=1.095
+ $X2=6.84 $Y2=1.095
r122 29 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.675 $Y=1.01
+ $X2=6.675 $Y2=1.095
r123 29 31 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=6.675 $Y=1.01
+ $X2=6.675 $Y2=0.515
r124 28 49 7.87875 $w=1.92e-07 $l=1.76125e-07 $layer=LI1_cond $X=5.84 $Y=1.095
+ $X2=5.675 $Y2=1.072
r125 27 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.51 $Y=1.095
+ $X2=6.675 $Y2=1.095
r126 27 28 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.51 $Y=1.095
+ $X2=5.84 $Y2=1.095
r127 23 49 0.50483 $w=3.3e-07 $l=1.07e-07 $layer=LI1_cond $X=5.675 $Y=0.965
+ $X2=5.675 $Y2=1.072
r128 23 25 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=5.675 $Y=0.965
+ $X2=5.675 $Y2=0.76
r129 22 48 7.11011 $w=1.7e-07 $l=1.5995e-07 $layer=LI1_cond $X=4.69 $Y=2.035
+ $X2=4.567 $Y2=1.95
r130 21 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.845 $Y=2.035
+ $X2=7.01 $Y2=2.035
r131 21 22 140.594 $w=1.68e-07 $l=2.155e-06 $layer=LI1_cond $X=6.845 $Y=2.035
+ $X2=4.69 $Y2=2.035
r132 20 47 3.52619 $w=2.15e-07 $l=2.13049e-07 $layer=LI1_cond $X=4.69 $Y=1.072
+ $X2=4.52 $Y2=0.975
r133 19 49 7.87875 $w=1.92e-07 $l=1.65e-07 $layer=LI1_cond $X=5.51 $Y=1.072
+ $X2=5.675 $Y2=1.072
r134 19 20 43.9536 $w=2.13e-07 $l=8.2e-07 $layer=LI1_cond $X=5.51 $Y=1.072
+ $X2=4.69 $Y2=1.072
r135 6 54 300 $w=1.7e-07 $l=2.90474e-07 $layer=licon1_PDIFF $count=2 $X=7.76
+ $Y=1.84 $X2=7.91 $Y2=2.065
r136 5 52 300 $w=1.7e-07 $l=2.98119e-07 $layer=licon1_PDIFF $count=2 $X=6.84
+ $Y=1.84 $X2=7.01 $Y2=2.065
r137 4 43 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.22
+ $Y=0.37 $X2=8.36 $Y2=0.515
r138 3 31 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=6.465
+ $Y=0.37 $X2=6.675 $Y2=0.515
r139 2 25 182 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_NDIFF $count=1 $X=5.535
+ $Y=0.37 $X2=5.675 $Y2=0.76
r140 1 47 182 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_NDIFF $count=1 $X=4.37
+ $Y=0.82 $X2=4.52 $Y2=0.965
.ends

.subckt PM_SKY130_FD_SC_LS__A31OI_4%A_30_74# 1 2 3 4 5 18 20 21 24 26 30 32 36
+ 38 42 44 45 46
c77 26 0 1.06564e-19 $X=1.92 $Y=1.095
r78 40 42 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=3.955 $Y=1.01
+ $X2=3.955 $Y2=0.76
r79 39 46 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=3.12 $Y=1.095
+ $X2=2.972 $Y2=1.095
r80 38 40 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.79 $Y=1.095
+ $X2=3.955 $Y2=1.01
r81 38 39 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.79 $Y=1.095
+ $X2=3.12 $Y2=1.095
r82 34 46 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=2.972 $Y=1.01
+ $X2=2.972 $Y2=1.095
r83 34 36 9.76647 $w=2.93e-07 $l=2.5e-07 $layer=LI1_cond $X=2.972 $Y=1.01
+ $X2=2.972 $Y2=0.76
r84 33 45 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.17 $Y=1.095
+ $X2=2.045 $Y2=1.095
r85 32 46 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=2.825 $Y=1.095
+ $X2=2.972 $Y2=1.095
r86 32 33 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=2.825 $Y=1.095
+ $X2=2.17 $Y2=1.095
r87 28 45 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.045 $Y=1.01
+ $X2=2.045 $Y2=1.095
r88 28 30 23.7403 $w=2.48e-07 $l=5.15e-07 $layer=LI1_cond $X=2.045 $Y=1.01
+ $X2=2.045 $Y2=0.495
r89 27 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.24 $Y=1.095
+ $X2=1.155 $Y2=1.095
r90 26 45 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.92 $Y=1.095
+ $X2=2.045 $Y2=1.095
r91 26 27 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.92 $Y=1.095
+ $X2=1.24 $Y2=1.095
r92 22 44 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.155 $Y=1.01
+ $X2=1.155 $Y2=1.095
r93 22 24 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=1.155 $Y=1.01
+ $X2=1.155 $Y2=0.515
r94 20 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.07 $Y=1.095
+ $X2=1.155 $Y2=1.095
r95 20 21 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.07 $Y=1.095
+ $X2=0.38 $Y2=1.095
r96 16 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.255 $Y=1.01
+ $X2=0.38 $Y2=1.095
r97 16 18 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=0.255 $Y=1.01
+ $X2=0.255 $Y2=0.515
r98 5 42 182 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_NDIFF $count=1 $X=3.815
+ $Y=0.37 $X2=3.955 $Y2=0.76
r99 4 36 182 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_NDIFF $count=1 $X=2.815
+ $Y=0.37 $X2=2.955 $Y2=0.76
r100 3 30 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.945
+ $Y=0.37 $X2=2.085 $Y2=0.495
r101 2 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.015
+ $Y=0.37 $X2=1.155 $Y2=0.515
r102 1 18 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.15
+ $Y=0.37 $X2=0.295 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__A31OI_4%VGND 1 2 3 12 16 18 20 25 37 38 41 44 48 54
r82 53 54 11.4973 $w=9.23e-07 $l=9.5e-08 $layer=LI1_cond $X=7.93 $Y=0.377
+ $X2=8.025 $Y2=0.377
r83 50 53 0.131892 $w=9.23e-07 $l=1e-08 $layer=LI1_cond $X=7.92 $Y=0.377
+ $X2=7.93 $Y2=0.377
r84 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r85 47 50 10.7492 $w=9.23e-07 $l=8.15e-07 $layer=LI1_cond $X=7.105 $Y=0.377
+ $X2=7.92 $Y2=0.377
r86 47 48 11.4973 $w=9.23e-07 $l=9.5e-08 $layer=LI1_cond $X=7.105 $Y=0.377
+ $X2=7.01 $Y2=0.377
r87 44 45 1.55 $w=1.7e-07 $l=1.02e-06 $layer=mcon $count=6 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r88 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r89 38 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=7.92
+ $Y2=0
r90 37 54 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=8.4 $Y=0 $X2=8.025
+ $Y2=0
r91 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r92 34 51 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.92
+ $Y2=0
r93 33 48 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=6.96 $Y=0 $X2=7.01
+ $Y2=0
r94 33 34 1.55 $w=1.7e-07 $l=1.02e-06 $layer=mcon $count=6 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r95 31 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.75 $Y=0 $X2=1.585
+ $Y2=0
r96 31 33 339.904 $w=1.68e-07 $l=5.21e-06 $layer=LI1_cond $X=1.75 $Y=0 $X2=6.96
+ $Y2=0
r97 29 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r98 29 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r99 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r100 26 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.89 $Y=0 $X2=0.725
+ $Y2=0
r101 26 28 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.89 $Y=0 $X2=1.2
+ $Y2=0
r102 25 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.42 $Y=0 $X2=1.585
+ $Y2=0
r103 25 28 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=1.42 $Y=0 $X2=1.2
+ $Y2=0
r104 23 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r105 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r106 20 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.56 $Y=0 $X2=0.725
+ $Y2=0
r107 20 22 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.56 $Y=0 $X2=0.24
+ $Y2=0
r108 18 34 0.73586 $w=4.9e-07 $l=2.64e-06 $layer=MET1_cond $X=4.32 $Y=0 $X2=6.96
+ $Y2=0
r109 18 45 0.73586 $w=4.9e-07 $l=2.64e-06 $layer=MET1_cond $X=4.32 $Y=0 $X2=1.68
+ $Y2=0
r110 14 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.585 $Y=0.085
+ $X2=1.585 $Y2=0
r111 14 16 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=1.585 $Y=0.085
+ $X2=1.585 $Y2=0.675
r112 10 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.725 $Y=0.085
+ $X2=0.725 $Y2=0
r113 10 12 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=0.725 $Y=0.085
+ $X2=0.725 $Y2=0.675
r114 3 53 121.333 $w=1.7e-07 $l=1.10705e-06 $layer=licon1_NDIFF $count=1
+ $X=6.965 $Y=0.37 $X2=7.93 $Y2=0.675
r115 3 47 121.333 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1
+ $X=6.965 $Y=0.37 $X2=7.105 $Y2=0.675
r116 2 16 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=1.445
+ $Y=0.37 $X2=1.585 $Y2=0.675
r117 1 12 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=0.585
+ $Y=0.37 $X2=0.725 $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_LS__A31OI_4%A_475_74# 1 2 3 4 15 17 18 21 23 27 29 33 35
+ 36
c62 33 0 1.25471e-19 $X=6.175 $Y=0.675
c63 15 0 1.69199e-19 $X=2.52 $Y=0.675
r64 31 33 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=6.175 $Y=0.425
+ $X2=6.175 $Y2=0.675
r65 30 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.265 $Y=0.34
+ $X2=5.1 $Y2=0.34
r66 29 31 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.01 $Y=0.34
+ $X2=6.175 $Y2=0.425
r67 29 30 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=6.01 $Y=0.34
+ $X2=5.265 $Y2=0.34
r68 25 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.1 $Y=0.425 $X2=5.1
+ $Y2=0.34
r69 25 27 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=5.1 $Y=0.425
+ $X2=5.1 $Y2=0.63
r70 24 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.62 $Y=0.34
+ $X2=3.455 $Y2=0.34
r71 23 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.935 $Y=0.34
+ $X2=5.1 $Y2=0.34
r72 23 24 85.7914 $w=1.68e-07 $l=1.315e-06 $layer=LI1_cond $X=4.935 $Y=0.34
+ $X2=3.62 $Y2=0.34
r73 19 35 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.455 $Y=0.425
+ $X2=3.455 $Y2=0.34
r74 19 21 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=3.455 $Y=0.425
+ $X2=3.455 $Y2=0.675
r75 17 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.29 $Y=0.34
+ $X2=3.455 $Y2=0.34
r76 17 18 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=3.29 $Y=0.34
+ $X2=2.655 $Y2=0.34
r77 13 18 7.55824 $w=1.7e-07 $l=1.90825e-07 $layer=LI1_cond $X=2.502 $Y=0.425
+ $X2=2.655 $Y2=0.34
r78 13 15 9.44625 $w=3.03e-07 $l=2.5e-07 $layer=LI1_cond $X=2.502 $Y=0.425
+ $X2=2.502 $Y2=0.675
r79 4 33 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=6.035
+ $Y=0.37 $X2=6.175 $Y2=0.675
r80 3 27 182 $w=1.7e-07 $l=3.94113e-07 $layer=licon1_NDIFF $count=1 $X=4.815
+ $Y=0.37 $X2=5.1 $Y2=0.63
r81 2 21 182 $w=1.7e-07 $l=3.96327e-07 $layer=licon1_NDIFF $count=1 $X=3.245
+ $Y=0.37 $X2=3.455 $Y2=0.675
r82 1 15 182 $w=1.7e-07 $l=3.70473e-07 $layer=licon1_NDIFF $count=1 $X=2.375
+ $Y=0.37 $X2=2.52 $Y2=0.675
.ends

