* NGSPICE file created from sky130_fd_sc_ls__dlrtn_4.ext - technology: sky130A

.subckt sky130_fd_sc_ls__dlrtn_4 D GATE_N RESET_B VGND VNB VPB VPWR Q
M1000 a_1035_74# RESET_B VGND VNB nshort w=640000u l=150000u
+  ad=5.44e+11p pd=5.54e+06u as=2.1144e+12p ps=1.632e+07u
M1001 a_888_406# a_639_392# VPWR VPB phighvt w=840000u l=150000u
+  ad=5.628e+11p pd=4.7e+06u as=2.7364e+12p ps=2.028e+07u
M1002 a_232_98# GATE_N VGND VNB nshort w=740000u l=150000u
+  ad=2.886e+11p pd=2.26e+06u as=0p ps=0u
M1003 VGND a_888_406# Q VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=4.144e+11p ps=4.08e+06u
M1004 VPWR a_888_406# Q VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=7.84e+11p ps=5.88e+06u
M1005 a_747_504# a_232_98# a_639_392# VPB phighvt w=420000u l=150000u
+  ad=3.024e+11p pd=2.28e+06u as=3.371e+11p ps=2.78e+06u
M1006 a_561_392# a_27_136# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.4e+11p pd=2.48e+06u as=0p ps=0u
M1007 a_839_74# a_348_392# a_639_392# VNB nshort w=420000u l=150000u
+  ad=1.155e+11p pd=1.39e+06u as=1.915e+11p ps=1.93e+06u
M1008 VPWR a_639_392# a_888_406# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR RESET_B a_888_406# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_1035_74# a_639_392# a_888_406# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1011 Q a_888_406# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR a_232_98# a_348_392# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=2.478e+11p ps=2.27e+06u
M1013 Q a_888_406# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR D a_27_136# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=2.478e+11p ps=2.27e+06u
M1015 a_888_406# RESET_B VPWR VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND a_888_406# a_839_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_639_392# a_232_98# a_666_74# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=1.536e+11p ps=1.76e+06u
M1018 a_666_74# a_27_136# VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_639_392# a_348_392# a_561_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR a_888_406# a_747_504# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND a_232_98# a_348_392# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1022 VPWR a_888_406# Q VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VGND RESET_B a_1035_74# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 Q a_888_406# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VGND D a_27_136# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1026 a_888_406# a_639_392# a_1035_74# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_232_98# GATE_N VPWR VPB phighvt w=840000u l=150000u
+  ad=2.478e+11p pd=2.27e+06u as=0p ps=0u
M1028 Q a_888_406# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VGND a_888_406# Q VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

