# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ls__or2b_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ls__or2b_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.760000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525000 1.450000 3.235000 1.780000 ;
    END
  END A
  PIN B_N
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.905000 1.120000 5.235000 1.790000 ;
    END
  END B_N
  PIN X
    ANTENNADIFFAREA  1.104900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.180000 0.775000 1.410000 ;
        RECT 0.545000 0.350000 0.795000 0.960000 ;
        RECT 0.545000 0.960000 1.805000 1.130000 ;
        RECT 0.545000 1.130000 0.775000 1.180000 ;
        RECT 0.605000 1.410000 0.775000 1.800000 ;
        RECT 0.605000 1.800000 1.785000 1.970000 ;
        RECT 0.605000 1.970000 0.805000 2.980000 ;
        RECT 1.455000 1.970000 1.785000 2.980000 ;
        RECT 1.475000 0.350000 1.805000 0.960000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 5.760000 0.085000 ;
        RECT 0.115000  0.085000 0.365000 1.010000 ;
        RECT 0.975000  0.085000 1.305000 0.765000 ;
        RECT 1.975000  0.085000 2.305000 0.940000 ;
        RECT 3.005000  0.085000 3.335000 0.940000 ;
        RECT 3.935000  0.085000 4.265000 1.030000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.760000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 5.760000 3.415000 ;
        RECT 0.105000 1.820000 0.435000 3.245000 ;
        RECT 1.005000 2.140000 1.255000 3.245000 ;
        RECT 1.985000 1.940000 2.235000 3.245000 ;
        RECT 2.960000 2.290000 3.210000 3.245000 ;
        RECT 4.875000 1.960000 5.205000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 5.760000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.945000 1.300000 2.145000 1.630000 ;
      RECT 1.975000 1.110000 3.755000 1.280000 ;
      RECT 1.975000 1.280000 2.145000 1.300000 ;
      RECT 2.430000 1.950000 3.675000 2.120000 ;
      RECT 2.430000 2.120000 2.760000 2.980000 ;
      RECT 2.475000 0.350000 2.805000 1.110000 ;
      RECT 3.425000 1.915000 3.675000 1.950000 ;
      RECT 3.425000 2.120000 3.675000 2.905000 ;
      RECT 3.425000 2.905000 4.655000 3.075000 ;
      RECT 3.505000 0.350000 3.755000 1.110000 ;
      RECT 3.505000 1.280000 4.125000 1.450000 ;
      RECT 3.875000 1.450000 4.125000 2.735000 ;
      RECT 4.295000 1.445000 4.625000 1.775000 ;
      RECT 4.325000 1.945000 4.655000 2.905000 ;
      RECT 4.435000 0.350000 5.655000 0.950000 ;
      RECT 4.435000 0.950000 4.625000 1.445000 ;
      RECT 5.405000 0.950000 5.655000 2.980000 ;
  END
END sky130_fd_sc_ls__or2b_4
