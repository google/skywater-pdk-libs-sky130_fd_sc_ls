* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__sedfxtp_2 CLK D DE SCD SCE VGND VNB VPB VPWR Q
M1000 a_1736_97# a_1538_74# a_693_113# VPB phighvt w=420000u l=150000u
+  ad=1.26e+11p pd=1.44e+06u as=4.983e+11p ps=5.16e+06u
M1001 VPWR a_1979_71# a_1936_508# VPB phighvt w=420000u l=150000u
+  ad=3.08865e+12p pd=2.56e+07u as=1.68e+11p ps=1.64e+06u
M1002 a_693_113# SCE a_40_464# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=3.808e+11p ps=3.75e+06u
M1003 VPWR SCE a_663_87# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.856e+11p ps=1.86e+06u
M1004 a_693_113# SCE a_1068_125# VNB nshort w=420000u l=150000u
+  ad=3.885e+11p pd=4.37e+06u as=8.82e+10p ps=1.26e+06u
M1005 a_138_74# D a_40_464# VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=2.982e+11p ps=3.1e+06u
M1006 a_2657_508# a_1538_74# a_2474_74# VPB phighvt w=420000u l=150000u
+  ad=1.134e+11p pd=1.38e+06u as=3.175e+11p ps=2.78e+06u
M1007 a_1936_508# a_1340_74# a_1736_97# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Q a_2474_74# VGND VNB nshort w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=2.2744e+12p ps=1.998e+07u
M1009 a_129_464# D a_40_464# VPB phighvt w=640000u l=150000u
+  ad=1.728e+11p pd=1.82e+06u as=0p ps=0u
M1010 a_693_113# a_663_87# a_1079_455# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1011 a_1340_74# CLK VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=0p ps=0u
M1012 a_1736_97# a_1340_74# a_693_113# VNB nshort w=420000u l=150000u
+  ad=2.226e+11p pd=1.9e+06u as=0p ps=0u
M1013 VGND DE a_180_290# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1014 a_575_463# DE VPWR VPB phighvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1015 a_500_113# a_180_290# VGND VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1016 a_1872_97# a_1538_74# a_1736_97# VNB nshort w=420000u l=150000u
+  ad=2.247e+11p pd=1.91e+06u as=0p ps=0u
M1017 a_1979_71# a_1736_97# VGND VNB nshort w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=0p ps=0u
M1018 a_1079_455# SCD VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND a_1979_71# a_1872_97# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_2569_74# a_1340_74# a_2474_74# VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=1.915e+11p ps=1.93e+06u
M1021 VGND a_548_87# a_2569_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPWR a_2474_74# Q VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.528e+11p ps=2.87e+06u
M1023 a_548_87# a_2474_74# VGND VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1024 a_1538_74# a_1340_74# VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1025 a_40_464# a_548_87# a_500_113# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_693_113# a_663_87# a_40_464# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 Q a_2474_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_2357_392# a_1979_71# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=8.1e+11p pd=3.62e+06u as=0p ps=0u
M1029 VGND DE a_138_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_1979_71# a_1736_97# VPWR VPB phighvt w=840000u l=150000u
+  ad=2.478e+11p pd=2.27e+06u as=0p ps=0u
M1031 VGND SCE a_663_87# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1032 a_40_464# a_548_87# a_575_463# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_1538_74# a_1340_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=0p ps=0u
M1034 VPWR a_180_290# a_129_464# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_548_87# a_2474_74# VPWR VPB phighvt w=640000u l=150000u
+  ad=1.888e+11p pd=1.87e+06u as=0p ps=0u
M1036 VGND a_2474_74# Q VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 VPWR a_548_87# a_2657_508# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 VPWR DE a_180_290# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.888e+11p ps=1.87e+06u
M1039 a_2402_74# a_1979_71# VGND VNB nshort w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1040 a_2474_74# a_1538_74# a_2402_74# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1041 a_1068_125# SCD VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1042 a_1340_74# CLK VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1043 a_2474_74# a_1340_74# a_2357_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
