* NGSPICE file created from sky130_fd_sc_ls__dlrtp_4.ext - technology: sky130A

.subckt sky130_fd_sc_ls__dlrtp_4 D GATE RESET_B VGND VNB VPB VPWR Q
M1000 a_240_394# GATE VPWR VPB phighvt w=840000u l=150000u
+  ad=2.94e+11p pd=2.38e+06u as=2.7109e+12p ps=2.052e+07u
M1001 a_562_392# a_27_126# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.4e+11p pd=2.48e+06u as=0p ps=0u
M1002 a_240_394# GATE VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=1.6158e+12p ps=1.463e+07u
M1003 a_797_48# a_640_74# a_938_74# VNB nshort w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=5.44e+11p ps=5.54e+06u
M1004 VPWR D a_27_126# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=2.478e+11p ps=2.27e+06u
M1005 Q a_797_48# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=7.504e+11p pd=5.82e+06u as=0p ps=0u
M1006 Q a_797_48# VGND VNB nshort w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=0p ps=0u
M1007 a_797_48# a_640_74# VPWR VPB phighvt w=840000u l=150000u
+  ad=5.46e+11p pd=4.66e+06u as=0p ps=0u
M1008 Q a_797_48# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR a_640_74# a_797_48# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR a_797_48# a_747_508# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.995e+11p ps=1.79e+06u
M1011 VPWR a_797_48# Q VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_640_74# a_240_394# a_562_392# VPB phighvt w=1e+06u l=150000u
+  ad=3.328e+11p pd=2.77e+06u as=0p ps=0u
M1013 VPWR a_797_48# Q VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND D a_27_126# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1015 a_797_48# RESET_B VPWR VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND RESET_B a_938_74# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND a_797_48# Q VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND a_240_394# a_364_120# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.294e+11p ps=2.1e+06u
M1019 Q a_797_48# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND a_797_48# a_755_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1021 VPWR a_240_394# a_364_120# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=2.478e+11p ps=2.27e+06u
M1022 VPWR RESET_B a_797_48# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_747_508# a_364_120# a_640_74# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_640_74# a_364_120# a_559_74# VNB nshort w=640000u l=150000u
+  ad=2.555e+11p pd=2.13e+06u as=1.632e+11p ps=1.79e+06u
M1025 a_938_74# RESET_B VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VGND a_797_48# Q VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_938_74# a_640_74# a_797_48# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_559_74# a_27_126# VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_755_74# a_240_394# a_640_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

