* NGSPICE file created from sky130_fd_sc_ls__dlrtn_1.ext - technology: sky130A

.subckt sky130_fd_sc_ls__dlrtn_1 D GATE_N RESET_B VGND VNB VPB VPWR Q
M1000 VPWR D a_27_136# VPB phighvt w=840000u l=150000u
+  ad=1.81275e+12p pd=1.271e+07u as=2.478e+11p ps=2.27e+06u
M1001 a_232_98# GATE_N VGND VNB nshort w=740000u l=150000u
+  ad=1.961e+11p pd=2.01e+06u as=1.64835e+12p ps=1.063e+07u
M1002 a_654_392# a_357_392# a_570_392# VPB phighvt w=1e+06u l=150000u
+  ad=4.029e+11p pd=3.09e+06u as=2.7e+11p ps=2.54e+06u
M1003 a_793_508# a_232_98# a_654_392# VPB phighvt w=420000u l=150000u
+  ad=2.247e+11p pd=1.91e+06u as=0p ps=0u
M1004 VGND a_897_406# a_854_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.155e+11p ps=1.39e+06u
M1005 a_570_392# a_27_136# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Q a_897_406# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=0p ps=0u
M1007 a_854_74# a_357_392# a_654_392# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.915e+11p ps=1.93e+06u
M1008 VGND RESET_B a_1139_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=1.776e+11p ps=1.96e+06u
M1009 VPWR a_232_98# a_357_392# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=2.478e+11p ps=2.27e+06u
M1010 a_897_406# a_654_392# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=4.7e+11p pd=2.94e+06u as=0p ps=0u
M1011 a_681_74# a_27_136# VGND VNB nshort w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1012 VGND D a_27_136# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1013 a_1139_74# a_654_392# a_897_406# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1014 Q a_897_406# VGND VNB nshort w=740000u l=150000u
+  ad=2.701e+11p pd=2.21e+06u as=0p ps=0u
M1015 VGND a_232_98# a_357_392# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1016 VPWR RESET_B a_897_406# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_654_392# a_232_98# a_681_74# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR a_897_406# a_793_508# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_232_98# GATE_N VPWR VPB phighvt w=840000u l=150000u
+  ad=2.478e+11p pd=2.27e+06u as=0p ps=0u
.ends

