* File: sky130_fd_sc_ls__o21ba_2.spice
* Created: Wed Sep  2 11:18:39 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__o21ba_2.pex.spice"
.subckt sky130_fd_sc_ls__o21ba_2  VNB VPB B1_N A2 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A2	A2
* B1_N	B1_N
* VPB	VPB
* VNB	VNB
MM1002 N_VGND_M1002_d N_B1_N_M1002_g N_A_27_74#_M1002_s VNB NSHORT L=0.15 W=0.55
+ AD=0.0964632 AS=0.15125 PD=0.90814 PS=1.65 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75001.1 A=0.0825 P=1.4 MULT=1
MM1000 N_VGND_M1002_d N_A_177_48#_M1000_g N_X_M1000_s VNB NSHORT L=0.15 W=0.74
+ AD=0.129787 AS=0.1036 PD=1.22186 PS=1.02 NRD=7.296 NRS=0 M=1 R=4.93333
+ SA=75000.5 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1006 N_VGND_M1006_d N_A_177_48#_M1006_g N_X_M1000_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2035 AS=0.1036 PD=2.03 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1011 N_A_487_74#_M1011_d N_A_27_74#_M1011_g N_A_177_48#_M1011_s VNB NSHORT
+ L=0.15 W=0.74 AD=0.1036 AS=0.2035 PD=1.02 PS=2.03 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001.2 A=0.111 P=1.78 MULT=1
MM1001 N_VGND_M1001_d N_A2_M1001_g N_A_487_74#_M1011_d VNB NSHORT L=0.15 W=0.74
+ AD=0.1797 AS=0.1036 PD=1.34 PS=1.02 NRD=30.456 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75000.8 A=0.111 P=1.78 MULT=1
MM1007 N_A_487_74#_M1007_d N_A1_M1007_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.74
+ AD=0.1998 AS=0.1797 PD=2.02 PS=1.34 NRD=0 NRS=30.456 M=1 R=4.93333 SA=75001.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1003 N_VPWR_M1003_d N_B1_N_M1003_g N_A_27_74#_M1003_s VPB PHIGHVT L=0.15
+ W=0.84 AD=0.1788 AS=0.2478 PD=1.29857 PS=2.27 NRD=37.0163 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75003.1 A=0.126 P=1.98 MULT=1
MM1005 N_X_M1005_d N_A_177_48#_M1005_g N_VPWR_M1003_d VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.2384 PD=1.42 PS=1.73143 NRD=1.7533 NRS=3.5066 M=1 R=7.46667
+ SA=75000.6 SB=75002.3 A=0.168 P=2.54 MULT=1
MM1010 N_X_M1005_d N_A_177_48#_M1010_g N_VPWR_M1010_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.427291 PD=1.42 PS=1.96 NRD=1.7533 NRS=2.6201 M=1 R=7.46667
+ SA=75001.1 SB=75001.9 A=0.168 P=2.54 MULT=1
MM1004 N_A_177_48#_M1004_d N_A_27_74#_M1004_g N_VPWR_M1010_s VPB PHIGHVT L=0.15
+ W=1 AD=0.15 AS=0.381509 PD=1.3 PS=1.75 NRD=1.9503 NRS=19.7 M=1 R=6.66667
+ SA=75002 SB=75001.2 A=0.15 P=2.3 MULT=1
MM1008 A_582_368# N_A2_M1008_g N_A_177_48#_M1004_d VPB PHIGHVT L=0.15 W=1
+ AD=0.18 AS=0.15 PD=1.36 PS=1.3 NRD=24.6053 NRS=1.9503 M=1 R=6.66667 SA=75002.5
+ SB=75000.7 A=0.15 P=2.3 MULT=1
MM1009 N_VPWR_M1009_d N_A1_M1009_g A_582_368# VPB PHIGHVT L=0.15 W=1 AD=0.285
+ AS=0.18 PD=2.57 PS=1.36 NRD=1.9503 NRS=24.6053 M=1 R=6.66667 SA=75003
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8492 P=12.16
*
.include "sky130_fd_sc_ls__o21ba_2.pxi.spice"
*
.ends
*
*
