* File: sky130_fd_sc_ls__inv_16.pex.spice
* Created: Fri Aug 28 13:27:55 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__INV_16%A 1 3 6 8 10 13 15 17 20 22 24 27 29 31 34 38
+ 40 42 45 47 49 52 54 56 59 61 63 66 68 70 73 75 77 80 82 84 87 89 91 94 96 98
+ 101 103 105 108 110 112 113 116 118 120 123 130 137 143 149 156 163 201 209
c332 120 0 1.29621e-19 $X=6.745 $Y=1.515
c333 116 0 1.2274e-19 $X=7.595 $Y=1.557
c334 113 0 1.20571e-19 $X=7.09 $Y=1.515
c335 80 0 1.79483e-19 $X=5.575 $Y=0.74
c336 66 0 1.75317e-19 $X=4.645 $Y=0.74
r337 196 201 0.638396 $w=2.3e-07 $l=9.95e-07 $layer=MET1_cond $X=5.93 $Y=1.665
+ $X2=6.925 $Y2=1.665
r338 191 196 0.638396 $w=2.3e-07 $l=9.95e-07 $layer=MET1_cond $X=4.935 $Y=1.665
+ $X2=5.93 $Y2=1.665
r339 191 209 0.548572 $w=2.3e-07 $l=8.55e-07 $layer=MET1_cond $X=4.935 $Y=1.665
+ $X2=4.08 $Y2=1.665
r340 176 181 0.603108 $w=2.3e-07 $l=9.4e-07 $layer=MET1_cond $X=2.17 $Y=1.665
+ $X2=3.11 $Y2=1.665
r341 171 176 0.603108 $w=2.3e-07 $l=9.4e-07 $layer=MET1_cond $X=1.23 $Y=1.665
+ $X2=2.17 $Y2=1.665
r342 166 167 10.6226 $w=3.63e-07 $l=8e-08 $layer=POLY_cond $X=6.575 $Y=1.557
+ $X2=6.655 $Y2=1.557
r343 165 166 49.1295 $w=3.63e-07 $l=3.7e-07 $layer=POLY_cond $X=6.205 $Y=1.557
+ $X2=6.575 $Y2=1.557
r344 164 165 7.96694 $w=3.63e-07 $l=6e-08 $layer=POLY_cond $X=6.145 $Y=1.557
+ $X2=6.205 $Y2=1.557
r345 163 196 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.93 $Y=1.665
+ $X2=5.93 $Y2=1.665
r346 162 164 28.5482 $w=3.63e-07 $l=2.15e-07 $layer=POLY_cond $X=5.93 $Y=1.557
+ $X2=6.145 $Y2=1.557
r347 162 163 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.93
+ $Y=1.515 $X2=5.93 $Y2=1.515
r348 160 162 36.5152 $w=3.63e-07 $l=2.75e-07 $layer=POLY_cond $X=5.655 $Y=1.557
+ $X2=5.93 $Y2=1.557
r349 159 160 10.6226 $w=3.63e-07 $l=8e-08 $layer=POLY_cond $X=5.575 $Y=1.557
+ $X2=5.655 $Y2=1.557
r350 158 159 53.1129 $w=3.63e-07 $l=4e-07 $layer=POLY_cond $X=5.175 $Y=1.557
+ $X2=5.575 $Y2=1.557
r351 157 158 3.98347 $w=3.63e-07 $l=3e-08 $layer=POLY_cond $X=5.145 $Y=1.557
+ $X2=5.175 $Y2=1.557
r352 156 191 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.935 $Y=1.665
+ $X2=4.935 $Y2=1.665
r353 155 157 27.8843 $w=3.63e-07 $l=2.1e-07 $layer=POLY_cond $X=4.935 $Y=1.557
+ $X2=5.145 $Y2=1.557
r354 155 156 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.935
+ $Y=1.515 $X2=4.935 $Y2=1.515
r355 153 155 30.5399 $w=3.63e-07 $l=2.3e-07 $layer=POLY_cond $X=4.705 $Y=1.557
+ $X2=4.935 $Y2=1.557
r356 152 153 7.96694 $w=3.63e-07 $l=6e-08 $layer=POLY_cond $X=4.645 $Y=1.557
+ $X2=4.705 $Y2=1.557
r357 151 152 51.7851 $w=3.63e-07 $l=3.9e-07 $layer=POLY_cond $X=4.255 $Y=1.557
+ $X2=4.645 $Y2=1.557
r358 150 151 5.31129 $w=3.63e-07 $l=4e-08 $layer=POLY_cond $X=4.215 $Y=1.557
+ $X2=4.255 $Y2=1.557
r359 148 150 25.2287 $w=3.63e-07 $l=1.9e-07 $layer=POLY_cond $X=4.025 $Y=1.557
+ $X2=4.215 $Y2=1.557
r360 148 149 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.025
+ $Y=1.515 $X2=4.025 $Y2=1.515
r361 146 148 29.2121 $w=3.63e-07 $l=2.2e-07 $layer=POLY_cond $X=3.805 $Y=1.557
+ $X2=4.025 $Y2=1.557
r362 145 146 2.65565 $w=3.63e-07 $l=2e-08 $layer=POLY_cond $X=3.785 $Y=1.557
+ $X2=3.805 $Y2=1.557
r363 144 145 57.0964 $w=3.63e-07 $l=4.3e-07 $layer=POLY_cond $X=3.355 $Y=1.557
+ $X2=3.785 $Y2=1.557
r364 143 181 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.11 $Y=1.665
+ $X2=3.11 $Y2=1.665
r365 142 144 32.5317 $w=3.63e-07 $l=2.45e-07 $layer=POLY_cond $X=3.11 $Y=1.557
+ $X2=3.355 $Y2=1.557
r366 142 143 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.11
+ $Y=1.515 $X2=3.11 $Y2=1.515
r367 140 142 33.8595 $w=3.63e-07 $l=2.55e-07 $layer=POLY_cond $X=2.855 $Y=1.557
+ $X2=3.11 $Y2=1.557
r368 139 140 57.0964 $w=3.63e-07 $l=4.3e-07 $layer=POLY_cond $X=2.425 $Y=1.557
+ $X2=2.855 $Y2=1.557
r369 138 139 2.65565 $w=3.63e-07 $l=2e-08 $layer=POLY_cond $X=2.405 $Y=1.557
+ $X2=2.425 $Y2=1.557
r370 137 176 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.17 $Y=1.665
+ $X2=2.17 $Y2=1.665
r371 136 138 31.2039 $w=3.63e-07 $l=2.35e-07 $layer=POLY_cond $X=2.17 $Y=1.557
+ $X2=2.405 $Y2=1.557
r372 136 137 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.17
+ $Y=1.515 $X2=2.17 $Y2=1.515
r373 134 136 32.5317 $w=3.63e-07 $l=2.45e-07 $layer=POLY_cond $X=1.925 $Y=1.557
+ $X2=2.17 $Y2=1.557
r374 133 134 2.65565 $w=3.63e-07 $l=2e-08 $layer=POLY_cond $X=1.905 $Y=1.557
+ $X2=1.925 $Y2=1.557
r375 132 133 54.4408 $w=3.63e-07 $l=4.1e-07 $layer=POLY_cond $X=1.495 $Y=1.557
+ $X2=1.905 $Y2=1.557
r376 131 132 5.31129 $w=3.63e-07 $l=4e-08 $layer=POLY_cond $X=1.455 $Y=1.557
+ $X2=1.495 $Y2=1.557
r377 130 171 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.23 $Y=1.665
+ $X2=1.23 $Y2=1.665
r378 129 131 29.876 $w=3.63e-07 $l=2.25e-07 $layer=POLY_cond $X=1.23 $Y=1.557
+ $X2=1.455 $Y2=1.557
r379 129 130 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.23
+ $Y=1.515 $X2=1.23 $Y2=1.515
r380 127 129 31.2039 $w=3.63e-07 $l=2.35e-07 $layer=POLY_cond $X=0.995 $Y=1.557
+ $X2=1.23 $Y2=1.557
r381 126 127 5.31129 $w=3.63e-07 $l=4e-08 $layer=POLY_cond $X=0.955 $Y=1.557
+ $X2=0.995 $Y2=1.557
r382 125 126 51.7851 $w=3.63e-07 $l=3.9e-07 $layer=POLY_cond $X=0.565 $Y=1.557
+ $X2=0.955 $Y2=1.557
r383 124 125 7.96694 $w=3.63e-07 $l=6e-08 $layer=POLY_cond $X=0.505 $Y=1.557
+ $X2=0.565 $Y2=1.557
r384 123 201 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.925 $Y=1.665
+ $X2=6.925 $Y2=1.665
r385 122 123 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.925
+ $Y=1.515 $X2=6.925 $Y2=1.515
r386 120 167 12.4447 $w=3.63e-07 $l=1.08995e-07 $layer=POLY_cond $X=6.745
+ $Y=1.515 $X2=6.655 $Y2=1.557
r387 120 122 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=6.745 $Y=1.515
+ $X2=6.925 $Y2=1.515
r388 118 209 0.0352882 $w=2.3e-07 $l=5.5e-08 $layer=MET1_cond $X=4.025 $Y=1.665
+ $X2=4.08 $Y2=1.665
r389 118 181 0.587068 $w=2.3e-07 $l=9.15e-07 $layer=MET1_cond $X=4.025 $Y=1.665
+ $X2=3.11 $Y2=1.665
r390 118 149 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.025 $Y=1.665
+ $X2=4.025 $Y2=1.665
r391 116 117 7.69149 $w=3.76e-07 $l=6e-08 $layer=POLY_cond $X=7.595 $Y=1.557
+ $X2=7.655 $Y2=1.557
r392 115 116 49.9947 $w=3.76e-07 $l=3.9e-07 $layer=POLY_cond $X=7.205 $Y=1.557
+ $X2=7.595 $Y2=1.557
r393 114 115 5.12766 $w=3.76e-07 $l=4e-08 $layer=POLY_cond $X=7.165 $Y=1.557
+ $X2=7.205 $Y2=1.557
r394 113 122 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.09 $Y=1.515
+ $X2=6.925 $Y2=1.515
r395 113 114 10.4594 $w=3.76e-07 $l=9.3675e-08 $layer=POLY_cond $X=7.09 $Y=1.515
+ $X2=7.165 $Y2=1.557
r396 110 117 24.356 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=7.655 $Y=1.765
+ $X2=7.655 $Y2=1.557
r397 110 112 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.655 $Y=1.765
+ $X2=7.655 $Y2=2.4
r398 106 116 24.356 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.595 $Y=1.35
+ $X2=7.595 $Y2=1.557
r399 106 108 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.595 $Y=1.35
+ $X2=7.595 $Y2=0.74
r400 103 115 24.356 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=7.205 $Y=1.765
+ $X2=7.205 $Y2=1.557
r401 103 105 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.205 $Y=1.765
+ $X2=7.205 $Y2=2.4
r402 99 114 24.356 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.165 $Y=1.35
+ $X2=7.165 $Y2=1.557
r403 99 101 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.165 $Y=1.35
+ $X2=7.165 $Y2=0.74
r404 96 167 23.5056 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=6.655 $Y=1.765
+ $X2=6.655 $Y2=1.557
r405 96 98 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.655 $Y=1.765
+ $X2=6.655 $Y2=2.4
r406 92 166 23.5056 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.575 $Y=1.35
+ $X2=6.575 $Y2=1.557
r407 92 94 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.575 $Y=1.35
+ $X2=6.575 $Y2=0.74
r408 89 165 23.5056 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=6.205 $Y=1.765
+ $X2=6.205 $Y2=1.557
r409 89 91 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.205 $Y=1.765
+ $X2=6.205 $Y2=2.4
r410 85 164 23.5056 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.145 $Y=1.35
+ $X2=6.145 $Y2=1.557
r411 85 87 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.145 $Y=1.35
+ $X2=6.145 $Y2=0.74
r412 82 160 23.5056 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=5.655 $Y=1.765
+ $X2=5.655 $Y2=1.557
r413 82 84 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.655 $Y=1.765
+ $X2=5.655 $Y2=2.4
r414 78 159 23.5056 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.575 $Y=1.35
+ $X2=5.575 $Y2=1.557
r415 78 80 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.575 $Y=1.35
+ $X2=5.575 $Y2=0.74
r416 75 158 23.5056 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=5.175 $Y=1.765
+ $X2=5.175 $Y2=1.557
r417 75 77 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.175 $Y=1.765
+ $X2=5.175 $Y2=2.4
r418 71 157 23.5056 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.145 $Y=1.35
+ $X2=5.145 $Y2=1.557
r419 71 73 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.145 $Y=1.35
+ $X2=5.145 $Y2=0.74
r420 68 153 23.5056 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=4.705 $Y=1.765
+ $X2=4.705 $Y2=1.557
r421 68 70 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.705 $Y=1.765
+ $X2=4.705 $Y2=2.4
r422 64 152 23.5056 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.645 $Y=1.35
+ $X2=4.645 $Y2=1.557
r423 64 66 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.645 $Y=1.35
+ $X2=4.645 $Y2=0.74
r424 61 151 23.5056 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=4.255 $Y=1.765
+ $X2=4.255 $Y2=1.557
r425 61 63 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.255 $Y=1.765
+ $X2=4.255 $Y2=2.4
r426 57 150 23.5056 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.215 $Y=1.35
+ $X2=4.215 $Y2=1.557
r427 57 59 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.215 $Y=1.35
+ $X2=4.215 $Y2=0.74
r428 54 146 23.5056 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.805 $Y=1.765
+ $X2=3.805 $Y2=1.557
r429 54 56 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.805 $Y=1.765
+ $X2=3.805 $Y2=2.4
r430 50 145 23.5056 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.785 $Y=1.35
+ $X2=3.785 $Y2=1.557
r431 50 52 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.785 $Y=1.35
+ $X2=3.785 $Y2=0.74
r432 47 144 23.5056 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.355 $Y=1.765
+ $X2=3.355 $Y2=1.557
r433 47 49 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.355 $Y=1.765
+ $X2=3.355 $Y2=2.4
r434 43 144 23.5056 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.355 $Y=1.35
+ $X2=3.355 $Y2=1.557
r435 43 45 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.355 $Y=1.35
+ $X2=3.355 $Y2=0.74
r436 40 140 23.5056 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.855 $Y=1.765
+ $X2=2.855 $Y2=1.557
r437 40 42 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.855 $Y=1.765
+ $X2=2.855 $Y2=2.4
r438 36 140 23.5056 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.855 $Y=1.35
+ $X2=2.855 $Y2=1.557
r439 36 38 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.855 $Y=1.35
+ $X2=2.855 $Y2=0.74
r440 32 139 23.5056 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.425 $Y=1.35
+ $X2=2.425 $Y2=1.557
r441 32 34 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.425 $Y=1.35
+ $X2=2.425 $Y2=0.74
r442 29 138 23.5056 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.405 $Y=1.765
+ $X2=2.405 $Y2=1.557
r443 29 31 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.405 $Y=1.765
+ $X2=2.405 $Y2=2.4
r444 25 134 23.5056 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.925 $Y=1.35
+ $X2=1.925 $Y2=1.557
r445 25 27 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.925 $Y=1.35
+ $X2=1.925 $Y2=0.74
r446 22 133 23.5056 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.905 $Y=1.765
+ $X2=1.905 $Y2=1.557
r447 22 24 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.905 $Y=1.765
+ $X2=1.905 $Y2=2.4
r448 18 132 23.5056 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.495 $Y=1.35
+ $X2=1.495 $Y2=1.557
r449 18 20 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.495 $Y=1.35
+ $X2=1.495 $Y2=0.74
r450 15 131 23.5056 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.455 $Y=1.765
+ $X2=1.455 $Y2=1.557
r451 15 17 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.455 $Y=1.765
+ $X2=1.455 $Y2=2.4
r452 11 127 23.5056 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.995 $Y=1.35
+ $X2=0.995 $Y2=1.557
r453 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.995 $Y=1.35
+ $X2=0.995 $Y2=0.74
r454 8 126 23.5056 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.955 $Y=1.765
+ $X2=0.955 $Y2=1.557
r455 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.955 $Y=1.765
+ $X2=0.955 $Y2=2.4
r456 4 125 23.5056 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.565 $Y=1.35
+ $X2=0.565 $Y2=1.557
r457 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.565 $Y=1.35
+ $X2=0.565 $Y2=0.74
r458 1 124 23.5056 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=1.557
r459 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__INV_16%VPWR 1 2 3 4 5 6 7 8 9 28 30 36 42 48 54 60
+ 66 72 76 78 83 84 86 87 88 90 95 100 112 116 121 130 133 136 139 142 146
c146 72 0 1.2274e-19 $X=6.93 $Y=2.105
r147 145 146 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r148 142 143 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r149 139 140 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r150 136 137 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r151 133 134 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r152 130 131 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r153 127 128 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r154 125 146 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r155 125 143 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6.96 $Y2=3.33
r156 124 125 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r157 122 142 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.095 $Y=3.33
+ $X2=6.93 $Y2=3.33
r158 122 124 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=7.095 $Y=3.33
+ $X2=7.44 $Y2=3.33
r159 121 145 4.55093 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=7.735 $Y=3.33
+ $X2=7.947 $Y2=3.33
r160 121 124 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=7.735 $Y=3.33
+ $X2=7.44 $Y2=3.33
r161 120 143 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6.96 $Y2=3.33
r162 120 140 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6 $Y2=3.33
r163 119 120 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r164 117 139 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.095 $Y=3.33
+ $X2=5.93 $Y2=3.33
r165 117 119 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=6.095 $Y=3.33
+ $X2=6.48 $Y2=3.33
r166 116 142 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.765 $Y=3.33
+ $X2=6.93 $Y2=3.33
r167 116 119 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=6.765 $Y=3.33
+ $X2=6.48 $Y2=3.33
r168 115 140 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6 $Y2=3.33
r169 114 115 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r170 112 139 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.765 $Y=3.33
+ $X2=5.93 $Y2=3.33
r171 112 114 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=5.765 $Y=3.33
+ $X2=5.52 $Y2=3.33
r172 111 115 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r173 110 111 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r174 108 137 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r175 107 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r176 105 136 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.245 $Y=3.33
+ $X2=3.12 $Y2=3.33
r177 105 107 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=3.245 $Y=3.33
+ $X2=3.6 $Y2=3.33
r178 104 137 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r179 104 134 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r180 103 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r181 101 133 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.295 $Y=3.33
+ $X2=2.17 $Y2=3.33
r182 101 103 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.295 $Y=3.33
+ $X2=2.64 $Y2=3.33
r183 100 136 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.995 $Y=3.33
+ $X2=3.12 $Y2=3.33
r184 100 103 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=2.995 $Y=3.33
+ $X2=2.64 $Y2=3.33
r185 99 134 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r186 99 131 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r187 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r188 96 130 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=1.345 $Y=3.33
+ $X2=1.2 $Y2=3.33
r189 96 98 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.345 $Y=3.33
+ $X2=1.68 $Y2=3.33
r190 95 133 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.045 $Y=3.33
+ $X2=2.17 $Y2=3.33
r191 95 98 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.045 $Y=3.33
+ $X2=1.68 $Y2=3.33
r192 94 131 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r193 94 128 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r194 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r195 91 127 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.182 $Y2=3.33
r196 91 93 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.72 $Y2=3.33
r197 90 130 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=1.055 $Y=3.33
+ $X2=1.2 $Y2=3.33
r198 90 93 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.055 $Y=3.33
+ $X2=0.72 $Y2=3.33
r199 88 111 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r200 88 108 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r201 86 110 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=4.81 $Y=3.33
+ $X2=4.56 $Y2=3.33
r202 86 87 7.75133 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=4.81 $Y=3.33
+ $X2=4.952 $Y2=3.33
r203 85 114 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=5.095 $Y=3.33
+ $X2=5.52 $Y2=3.33
r204 85 87 7.75133 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=5.095 $Y=3.33
+ $X2=4.952 $Y2=3.33
r205 83 107 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=3.915 $Y=3.33
+ $X2=3.6 $Y2=3.33
r206 83 84 6.70225 $w=1.7e-07 $l=1.17e-07 $layer=LI1_cond $X=3.915 $Y=3.33
+ $X2=4.032 $Y2=3.33
r207 82 110 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=4.15 $Y=3.33
+ $X2=4.56 $Y2=3.33
r208 82 84 6.70225 $w=1.7e-07 $l=1.18e-07 $layer=LI1_cond $X=4.15 $Y=3.33
+ $X2=4.032 $Y2=3.33
r209 78 81 30.8557 $w=3.08e-07 $l=8.3e-07 $layer=LI1_cond $X=7.89 $Y=1.985
+ $X2=7.89 $Y2=2.815
r210 76 145 3.04826 $w=3.1e-07 $l=1.09864e-07 $layer=LI1_cond $X=7.89 $Y=3.245
+ $X2=7.947 $Y2=3.33
r211 76 81 15.9855 $w=3.08e-07 $l=4.3e-07 $layer=LI1_cond $X=7.89 $Y=3.245
+ $X2=7.89 $Y2=2.815
r212 72 75 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=6.93 $Y=2.105
+ $X2=6.93 $Y2=2.815
r213 70 142 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.93 $Y=3.245
+ $X2=6.93 $Y2=3.33
r214 70 75 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=6.93 $Y=3.245
+ $X2=6.93 $Y2=2.815
r215 66 69 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=5.93 $Y=2.105
+ $X2=5.93 $Y2=2.815
r216 64 139 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.93 $Y=3.245
+ $X2=5.93 $Y2=3.33
r217 64 69 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=5.93 $Y=3.245
+ $X2=5.93 $Y2=2.815
r218 60 63 28.71 $w=2.83e-07 $l=7.1e-07 $layer=LI1_cond $X=4.952 $Y=2.105
+ $X2=4.952 $Y2=2.815
r219 58 87 0.432977 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=4.952 $Y=3.245
+ $X2=4.952 $Y2=3.33
r220 58 63 17.3877 $w=2.83e-07 $l=4.3e-07 $layer=LI1_cond $X=4.952 $Y=3.245
+ $X2=4.952 $Y2=2.815
r221 54 57 34.8185 $w=2.33e-07 $l=7.1e-07 $layer=LI1_cond $X=4.032 $Y=2.105
+ $X2=4.032 $Y2=2.815
r222 52 84 0.207053 $w=2.35e-07 $l=8.5e-08 $layer=LI1_cond $X=4.032 $Y=3.245
+ $X2=4.032 $Y2=3.33
r223 52 57 21.0873 $w=2.33e-07 $l=4.3e-07 $layer=LI1_cond $X=4.032 $Y=3.245
+ $X2=4.032 $Y2=2.815
r224 48 51 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=3.12 $Y=2.105
+ $X2=3.12 $Y2=2.815
r225 46 136 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.12 $Y=3.245
+ $X2=3.12 $Y2=3.33
r226 46 51 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=3.12 $Y=3.245
+ $X2=3.12 $Y2=2.815
r227 42 45 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=2.17 $Y=2.105
+ $X2=2.17 $Y2=2.815
r228 40 133 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.17 $Y=3.245
+ $X2=2.17 $Y2=3.33
r229 40 45 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=2.17 $Y=3.245
+ $X2=2.17 $Y2=2.815
r230 36 39 28.215 $w=2.88e-07 $l=7.1e-07 $layer=LI1_cond $X=1.2 $Y=2.105 $X2=1.2
+ $Y2=2.815
r231 34 130 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=3.245
+ $X2=1.2 $Y2=3.33
r232 34 39 17.0879 $w=2.88e-07 $l=4.3e-07 $layer=LI1_cond $X=1.2 $Y=3.245
+ $X2=1.2 $Y2=2.815
r233 30 33 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=0.24 $Y=1.985
+ $X2=0.24 $Y2=2.815
r234 28 127 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.182 $Y2=3.33
r235 28 33 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.24 $Y2=2.815
r236 9 81 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=7.73
+ $Y=1.84 $X2=7.88 $Y2=2.815
r237 9 78 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=7.73
+ $Y=1.84 $X2=7.88 $Y2=1.985
r238 8 75 400 $w=1.7e-07 $l=1.07034e-06 $layer=licon1_PDIFF $count=1 $X=6.73
+ $Y=1.84 $X2=6.93 $Y2=2.815
r239 8 72 400 $w=1.7e-07 $l=3.51034e-07 $layer=licon1_PDIFF $count=1 $X=6.73
+ $Y=1.84 $X2=6.93 $Y2=2.105
r240 7 69 400 $w=1.7e-07 $l=1.07034e-06 $layer=licon1_PDIFF $count=1 $X=5.73
+ $Y=1.84 $X2=5.93 $Y2=2.815
r241 7 66 400 $w=1.7e-07 $l=3.51034e-07 $layer=licon1_PDIFF $count=1 $X=5.73
+ $Y=1.84 $X2=5.93 $Y2=2.105
r242 6 63 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=4.78
+ $Y=1.84 $X2=4.93 $Y2=2.815
r243 6 60 400 $w=1.7e-07 $l=3.31625e-07 $layer=licon1_PDIFF $count=1 $X=4.78
+ $Y=1.84 $X2=4.93 $Y2=2.105
r244 5 57 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=3.88
+ $Y=1.84 $X2=4.03 $Y2=2.815
r245 5 54 400 $w=1.7e-07 $l=3.31625e-07 $layer=licon1_PDIFF $count=1 $X=3.88
+ $Y=1.84 $X2=4.03 $Y2=2.105
r246 4 51 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.93
+ $Y=1.84 $X2=3.08 $Y2=2.815
r247 4 48 400 $w=1.7e-07 $l=3.31625e-07 $layer=licon1_PDIFF $count=1 $X=2.93
+ $Y=1.84 $X2=3.08 $Y2=2.105
r248 3 45 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.98
+ $Y=1.84 $X2=2.13 $Y2=2.815
r249 3 42 400 $w=1.7e-07 $l=3.31625e-07 $layer=licon1_PDIFF $count=1 $X=1.98
+ $Y=1.84 $X2=2.13 $Y2=2.105
r250 2 39 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.03
+ $Y=1.84 $X2=1.18 $Y2=2.815
r251 2 36 400 $w=1.7e-07 $l=3.31625e-07 $layer=licon1_PDIFF $count=1 $X=1.03
+ $Y=1.84 $X2=1.18 $Y2=2.105
r252 1 33 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r253 1 30 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_LS__INV_16%Y 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 51
+ 57 61 65 69 73 77 79 81 83 85 89 91 92 93 97 98 101 108 118 125 132 134 139
+ 144 149
c245 144 0 1.29621e-19 $X=2.63 $Y=1.985
c246 134 0 1.20571e-19 $X=7.43 $Y=2.035
c247 91 0 1.71499e-19 $X=0.725 $Y=1.49
c248 83 0 1.79483e-19 $X=6.36 $Y=1.015
c249 79 0 1.75317e-19 $X=5.37 $Y=1.025
r250 149 152 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.48 $Y=2.035
+ $X2=4.48 $Y2=2.035
r251 149 150 1.98543 $w=2.88e-07 $l=4.5e-08 $layer=LI1_cond $X=4.485 $Y=1.985
+ $X2=4.485 $Y2=1.94
r252 144 147 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.63 $Y=2.035
+ $X2=2.63 $Y2=2.035
r253 144 145 1.62839 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=2.63 $Y=1.985
+ $X2=2.63 $Y2=1.94
r254 142 147 0.609524 $w=2.3e-07 $l=9.5e-07 $layer=MET1_cond $X=1.68 $Y=2.035
+ $X2=2.63 $Y2=2.035
r255 139 142 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=2.035
+ $X2=1.68 $Y2=2.035
r256 139 140 3.16711 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=1.68 $Y=2.025
+ $X2=1.68 $Y2=1.94
r257 132 136 34.1617 $w=2.78e-07 $l=8.3e-07 $layer=LI1_cond $X=7.405 $Y=1.985
+ $X2=7.405 $Y2=2.815
r258 132 134 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.43 $Y=2.035
+ $X2=7.43 $Y2=2.035
r259 127 134 0.641604 $w=2.3e-07 $l=1e-06 $layer=MET1_cond $X=6.43 $Y=2.035
+ $X2=7.43 $Y2=2.035
r260 125 129 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=6.43 $Y=1.985
+ $X2=6.43 $Y2=2.815
r261 125 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.43 $Y=2.035
+ $X2=6.43 $Y2=2.035
r262 120 127 0.641604 $w=2.3e-07 $l=1e-06 $layer=MET1_cond $X=5.43 $Y=2.035
+ $X2=6.43 $Y2=2.035
r263 120 152 0.609524 $w=2.3e-07 $l=9.5e-07 $layer=MET1_cond $X=5.43 $Y=2.035
+ $X2=4.48 $Y2=2.035
r264 118 122 30.366 $w=3.13e-07 $l=8.3e-07 $layer=LI1_cond $X=5.422 $Y=1.985
+ $X2=5.422 $Y2=2.815
r265 118 120 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.43 $Y=2.035
+ $X2=5.43 $Y2=2.035
r266 113 147 0.609524 $w=2.3e-07 $l=9.5e-07 $layer=MET1_cond $X=3.58 $Y=2.035
+ $X2=2.63 $Y2=2.035
r267 111 115 32.4247 $w=2.93e-07 $l=8.3e-07 $layer=LI1_cond $X=3.562 $Y=1.985
+ $X2=3.562 $Y2=2.815
r268 111 113 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.58 $Y=2.035
+ $X2=3.58 $Y2=2.035
r269 108 111 57.4268 $w=2.93e-07 $l=1.47e-06 $layer=LI1_cond $X=3.562 $Y=0.515
+ $X2=3.562 $Y2=1.985
r270 103 142 0.609524 $w=2.3e-07 $l=9.5e-07 $layer=MET1_cond $X=0.73 $Y=2.035
+ $X2=1.68 $Y2=2.035
r271 101 105 29.8915 $w=3.18e-07 $l=8.3e-07 $layer=LI1_cond $X=0.725 $Y=1.985
+ $X2=0.725 $Y2=2.815
r272 101 103 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.73 $Y=2.035
+ $X2=0.73 $Y2=2.035
r273 98 152 0.256642 $w=2.3e-07 $l=4e-07 $layer=MET1_cond $X=4.08 $Y=2.035
+ $X2=4.48 $Y2=2.035
r274 98 113 0.320802 $w=2.3e-07 $l=5e-07 $layer=MET1_cond $X=4.08 $Y=2.035
+ $X2=3.58 $Y2=2.035
r275 97 132 35.1907 $w=2.78e-07 $l=8.55e-07 $layer=LI1_cond $X=7.405 $Y=1.13
+ $X2=7.405 $Y2=1.985
r276 95 125 18.6835 $w=3.28e-07 $l=5.35e-07 $layer=LI1_cond $X=6.43 $Y=1.45
+ $X2=6.43 $Y2=1.985
r277 94 118 19.8659 $w=3.13e-07 $l=5.43e-07 $layer=LI1_cond $X=5.422 $Y=1.442
+ $X2=5.422 $Y2=1.985
r278 92 93 8.53661 $w=2.68e-07 $l=2e-07 $layer=LI1_cond $X=0.75 $Y=1.33 $X2=0.75
+ $Y2=1.13
r279 91 101 17.8269 $w=3.18e-07 $l=4.95e-07 $layer=LI1_cond $X=0.725 $Y=1.49
+ $X2=0.725 $Y2=1.985
r280 91 92 6.07707 $w=3.18e-07 $l=1.6e-07 $layer=LI1_cond $X=0.725 $Y=1.49
+ $X2=0.725 $Y2=1.33
r281 87 97 6.05995 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.38 $Y=0.965
+ $X2=7.38 $Y2=1.13
r282 87 89 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=7.38 $Y=0.965
+ $X2=7.38 $Y2=0.515
r283 83 95 16.9553 $w=3.13e-07 $l=4.68695e-07 $layer=LI1_cond $X=6.36 $Y=1.015
+ $X2=6.43 $Y2=1.45
r284 83 85 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=6.36 $Y=1.015
+ $X2=6.36 $Y2=0.515
r285 79 94 17.0147 $w=2.99e-07 $l=4.42236e-07 $layer=LI1_cond $X=5.37 $Y=1.025
+ $X2=5.422 $Y2=1.442
r286 79 81 18.9595 $w=3.08e-07 $l=5.1e-07 $layer=LI1_cond $X=5.37 $Y=1.025
+ $X2=5.37 $Y2=0.515
r287 75 149 3.97394 $w=2.88e-07 $l=1e-07 $layer=LI1_cond $X=4.485 $Y=2.085
+ $X2=4.485 $Y2=1.985
r288 75 77 12.5179 $w=2.88e-07 $l=3.15e-07 $layer=LI1_cond $X=4.485 $Y=2.085
+ $X2=4.485 $Y2=2.4
r289 73 150 64.4012 $w=2.53e-07 $l=1.425e-06 $layer=LI1_cond $X=4.467 $Y=0.515
+ $X2=4.467 $Y2=1.94
r290 69 145 52.9752 $w=3.08e-07 $l=1.425e-06 $layer=LI1_cond $X=2.64 $Y=0.515
+ $X2=2.64 $Y2=1.94
r291 63 144 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=2.63 $Y=2.105
+ $X2=2.63 $Y2=1.985
r292 63 65 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.63 $Y=2.105
+ $X2=2.63 $Y2=2.4
r293 61 140 56.6287 $w=2.88e-07 $l=1.425e-06 $layer=LI1_cond $X=1.7 $Y=0.515
+ $X2=1.7 $Y2=1.94
r294 55 139 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=1.68 $Y=2.105
+ $X2=1.68 $Y2=2.025
r295 55 57 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=1.68 $Y=2.105
+ $X2=1.68 $Y2=2.815
r296 49 93 6.17723 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.78 $Y=0.965
+ $X2=0.78 $Y2=1.13
r297 49 51 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=0.78 $Y=0.965
+ $X2=0.78 $Y2=0.515
r298 16 136 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=7.28
+ $Y=1.84 $X2=7.43 $Y2=2.815
r299 16 132 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=7.28
+ $Y=1.84 $X2=7.43 $Y2=1.985
r300 15 129 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=6.28
+ $Y=1.84 $X2=6.43 $Y2=2.815
r301 15 125 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=6.28
+ $Y=1.84 $X2=6.43 $Y2=1.985
r302 14 122 400 $w=1.7e-07 $l=1.06119e-06 $layer=licon1_PDIFF $count=1 $X=5.25
+ $Y=1.84 $X2=5.43 $Y2=2.815
r303 14 118 400 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_PDIFF $count=1 $X=5.25
+ $Y=1.84 $X2=5.43 $Y2=1.985
r304 13 149 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=4.33
+ $Y=1.84 $X2=4.48 $Y2=1.985
r305 13 77 300 $w=1.7e-07 $l=6.30555e-07 $layer=licon1_PDIFF $count=2 $X=4.33
+ $Y=1.84 $X2=4.48 $Y2=2.4
r306 12 115 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=3.43
+ $Y=1.84 $X2=3.58 $Y2=2.815
r307 12 111 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=3.43
+ $Y=1.84 $X2=3.58 $Y2=1.985
r308 11 144 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.48
+ $Y=1.84 $X2=2.63 $Y2=1.985
r309 11 65 300 $w=1.7e-07 $l=6.30555e-07 $layer=licon1_PDIFF $count=2 $X=2.48
+ $Y=1.84 $X2=2.63 $Y2=2.4
r310 10 139 400 $w=1.7e-07 $l=2.48948e-07 $layer=licon1_PDIFF $count=1 $X=1.53
+ $Y=1.84 $X2=1.68 $Y2=2.025
r311 10 57 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.53
+ $Y=1.84 $X2=1.68 $Y2=2.815
r312 9 105 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.84 $X2=0.73 $Y2=2.815
r313 9 101 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.84 $X2=0.73 $Y2=1.985
r314 8 89 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.24
+ $Y=0.37 $X2=7.38 $Y2=0.515
r315 7 85 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.22
+ $Y=0.37 $X2=6.36 $Y2=0.515
r316 6 81 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.22
+ $Y=0.37 $X2=5.36 $Y2=0.515
r317 5 73 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.29
+ $Y=0.37 $X2=4.43 $Y2=0.515
r318 4 108 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.43
+ $Y=0.37 $X2=3.57 $Y2=0.515
r319 3 69 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.5
+ $Y=0.37 $X2=2.64 $Y2=0.515
r320 2 61 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.57
+ $Y=0.37 $X2=1.71 $Y2=0.515
r321 1 51 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.64
+ $Y=0.37 $X2=0.78 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__INV_16%VGND 1 2 3 4 5 6 7 8 9 28 30 34 38 42 46 50
+ 54 58 60 62 65 66 68 69 71 72 73 75 80 85 100 104 113 116 119 122 126
r136 125 126 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r137 122 123 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r138 119 120 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r139 116 117 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r140 113 114 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r141 110 111 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r142 108 126 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=7.92 $Y2=0
r143 108 123 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=6.96 $Y2=0
r144 107 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r145 105 122 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=7.045 $Y=0
+ $X2=6.875 $Y2=0
r146 105 107 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=7.045 $Y=0
+ $X2=7.44 $Y2=0
r147 104 125 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=7.715 $Y=0
+ $X2=7.937 $Y2=0
r148 104 107 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=7.715 $Y=0
+ $X2=7.44 $Y2=0
r149 103 123 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0
+ $X2=6.96 $Y2=0
r150 102 103 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r151 100 122 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=6.705 $Y=0
+ $X2=6.875 $Y2=0
r152 100 102 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=6.705 $Y=0
+ $X2=6.48 $Y2=0
r153 99 103 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0
+ $X2=6.48 $Y2=0
r154 98 99 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r155 96 99 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.52
+ $Y2=0
r156 95 96 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r157 93 120 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r158 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r159 90 119 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.245 $Y=0
+ $X2=3.11 $Y2=0
r160 90 92 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=3.245 $Y=0 $X2=3.6
+ $Y2=0
r161 89 120 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=3.12 $Y2=0
r162 89 117 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=2.16 $Y2=0
r163 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r164 86 116 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.305 $Y=0 $X2=2.165
+ $Y2=0
r165 86 88 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.305 $Y=0
+ $X2=2.64 $Y2=0
r166 85 119 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.975 $Y=0
+ $X2=3.11 $Y2=0
r167 85 88 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.975 $Y=0
+ $X2=2.64 $Y2=0
r168 84 117 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0
+ $X2=2.16 $Y2=0
r169 84 114 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r170 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r171 81 113 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.375 $Y=0
+ $X2=1.245 $Y2=0
r172 81 83 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.375 $Y=0
+ $X2=1.68 $Y2=0
r173 80 116 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.025 $Y=0 $X2=2.165
+ $Y2=0
r174 80 83 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.025 $Y=0 $X2=1.68
+ $Y2=0
r175 79 114 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r176 79 111 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0
+ $X2=0.24 $Y2=0
r177 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r178 76 110 4.01078 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=0
+ $X2=0.222 $Y2=0
r179 76 78 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=0
+ $X2=0.72 $Y2=0
r180 75 113 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.115 $Y=0
+ $X2=1.245 $Y2=0
r181 75 78 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.115 $Y=0
+ $X2=0.72 $Y2=0
r182 73 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r183 73 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r184 71 98 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=5.705 $Y=0
+ $X2=5.52 $Y2=0
r185 71 72 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=5.705 $Y=0 $X2=5.865
+ $Y2=0
r186 70 102 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=6.025 $Y=0
+ $X2=6.48 $Y2=0
r187 70 72 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=6.025 $Y=0 $X2=5.865
+ $Y2=0
r188 68 95 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=4.765 $Y=0
+ $X2=4.56 $Y2=0
r189 68 69 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.765 $Y=0 $X2=4.895
+ $Y2=0
r190 67 98 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=5.025 $Y=0
+ $X2=5.52 $Y2=0
r191 67 69 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.025 $Y=0 $X2=4.895
+ $Y2=0
r192 65 92 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=3.89 $Y=0 $X2=3.6
+ $Y2=0
r193 65 66 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.89 $Y=0 $X2=4.02
+ $Y2=0
r194 64 95 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=4.15 $Y=0 $X2=4.56
+ $Y2=0
r195 64 66 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.15 $Y=0 $X2=4.02
+ $Y2=0
r196 60 125 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=7.88 $Y=0.085
+ $X2=7.937 $Y2=0
r197 60 62 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=7.88 $Y=0.085
+ $X2=7.88 $Y2=0.515
r198 56 122 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=6.875 $Y=0.085
+ $X2=6.875 $Y2=0
r199 56 58 15.0834 $w=3.38e-07 $l=4.45e-07 $layer=LI1_cond $X=6.875 $Y=0.085
+ $X2=6.875 $Y2=0.53
r200 52 72 0.800721 $w=3.2e-07 $l=8.5e-08 $layer=LI1_cond $X=5.865 $Y=0.085
+ $X2=5.865 $Y2=0
r201 52 54 16.0262 $w=3.18e-07 $l=4.45e-07 $layer=LI1_cond $X=5.865 $Y=0.085
+ $X2=5.865 $Y2=0.53
r202 48 69 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=4.895 $Y=0.085
+ $X2=4.895 $Y2=0
r203 48 50 19.7245 $w=2.58e-07 $l=4.45e-07 $layer=LI1_cond $X=4.895 $Y=0.085
+ $X2=4.895 $Y2=0.53
r204 44 66 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=4.02 $Y=0.085
+ $X2=4.02 $Y2=0
r205 44 46 19.0596 $w=2.58e-07 $l=4.3e-07 $layer=LI1_cond $X=4.02 $Y=0.085
+ $X2=4.02 $Y2=0.515
r206 40 119 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.11 $Y=0.085
+ $X2=3.11 $Y2=0
r207 40 42 18.3537 $w=2.68e-07 $l=4.3e-07 $layer=LI1_cond $X=3.11 $Y=0.085
+ $X2=3.11 $Y2=0.515
r208 36 116 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.165 $Y=0.085
+ $X2=2.165 $Y2=0
r209 36 38 17.6982 $w=2.78e-07 $l=4.3e-07 $layer=LI1_cond $X=2.165 $Y=0.085
+ $X2=2.165 $Y2=0.515
r210 32 113 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.245 $Y=0.085
+ $X2=1.245 $Y2=0
r211 32 34 19.0596 $w=2.58e-07 $l=4.3e-07 $layer=LI1_cond $X=1.245 $Y=0.085
+ $X2=1.245 $Y2=0.515
r212 28 110 3.20143 $w=2.6e-07 $l=1.28662e-07 $layer=LI1_cond $X=0.315 $Y=0.085
+ $X2=0.222 $Y2=0
r213 28 30 19.0596 $w=2.58e-07 $l=4.3e-07 $layer=LI1_cond $X=0.315 $Y=0.085
+ $X2=0.315 $Y2=0.515
r214 9 62 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.67
+ $Y=0.37 $X2=7.81 $Y2=0.515
r215 8 58 91 $w=1.7e-07 $l=2.89137e-07 $layer=licon1_NDIFF $count=2 $X=6.65
+ $Y=0.37 $X2=6.87 $Y2=0.53
r216 7 54 91 $w=1.7e-07 $l=2.78747e-07 $layer=licon1_NDIFF $count=2 $X=5.65
+ $Y=0.37 $X2=5.86 $Y2=0.53
r217 6 50 91 $w=1.7e-07 $l=2.42126e-07 $layer=licon1_NDIFF $count=2 $X=4.72
+ $Y=0.37 $X2=4.895 $Y2=0.53
r218 5 46 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.86
+ $Y=0.37 $X2=4 $Y2=0.515
r219 4 42 91 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_NDIFF $count=2 $X=2.93
+ $Y=0.37 $X2=3.12 $Y2=0.515
r220 3 38 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2 $Y=0.37
+ $X2=2.14 $Y2=0.515
r221 2 34 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=1.07
+ $Y=0.37 $X2=1.28 $Y2=0.515
r222 1 30 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.225
+ $Y=0.37 $X2=0.35 $Y2=0.515
.ends

