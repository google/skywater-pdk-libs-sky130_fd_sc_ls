* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__bufbuf_16 A VGND VNB VPB VPWR X
X0 VGND a_588_74# X VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X1 X a_588_74# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X2 X a_588_74# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X3 a_588_74# a_203_74# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X4 a_588_74# a_203_74# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X5 a_588_74# a_203_74# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X6 VGND a_588_74# X VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X7 VPWR a_588_74# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X8 VGND a_588_74# X VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X9 a_203_74# a_27_368# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X10 X a_588_74# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X11 VPWR a_588_74# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X12 VGND a_27_368# a_203_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X13 VGND a_588_74# X VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X14 X a_588_74# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X15 VPWR a_588_74# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X16 VGND a_27_368# a_203_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X17 VGND a_203_74# a_588_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X18 VGND a_588_74# X VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X19 VPWR a_588_74# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X20 X a_588_74# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X21 VPWR a_588_74# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X22 VPWR a_588_74# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X23 X a_588_74# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X24 a_27_368# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X25 VPWR a_588_74# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X26 X a_588_74# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X27 a_203_74# a_27_368# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X28 VPWR a_203_74# a_588_74# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X29 VGND a_203_74# a_588_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X30 X a_588_74# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X31 VPWR a_203_74# a_588_74# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X32 a_588_74# a_203_74# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X33 X a_588_74# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X34 VPWR a_203_74# a_588_74# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X35 X a_588_74# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X36 VGND a_588_74# X VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X37 VPWR a_27_368# a_203_74# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X38 X a_588_74# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X39 a_588_74# a_203_74# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X40 X a_588_74# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X41 VPWR a_27_368# a_203_74# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X42 X a_588_74# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X43 X a_588_74# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X44 VGND a_203_74# a_588_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X45 a_27_368# A VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X46 a_588_74# a_203_74# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X47 X a_588_74# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X48 X a_588_74# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X49 VPWR a_588_74# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X50 VGND a_588_74# X VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X51 VGND a_588_74# X VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
.ends
