# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ls__mux4_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ls__mux4_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.56000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A0
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.315000 1.450000 3.685000 1.780000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.975000 1.450000 1.315000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.915000 1.180000 6.345000 1.780000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.855000 1.450000 4.195000 1.780000 ;
    END
  END A3
  PIN S0
    ANTENNAGATEAREA  0.768000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.435000 1.180000 1.655000 1.260000 ;
        RECT 0.435000 1.260000 1.845000 1.280000 ;
        RECT 0.435000 1.280000 0.805000 1.550000 ;
        RECT 0.635000 1.110000 1.655000 1.180000 ;
        RECT 1.485000 0.420000 3.105000 0.590000 ;
        RECT 1.485000 0.590000 1.655000 1.110000 ;
        RECT 1.485000 1.280000 1.845000 1.590000 ;
        RECT 2.835000 0.590000 3.105000 1.110000 ;
        RECT 2.835000 1.110000 5.745000 1.280000 ;
        RECT 2.835000 1.280000 3.105000 1.780000 ;
        RECT 4.395000 1.280000 4.725000 1.550000 ;
        RECT 5.475000 1.280000 5.745000 1.750000 ;
    END
  END S0
  PIN S1
    ANTENNAGATEAREA  0.507000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.900000 1.450000 7.555000 1.780000 ;
    END
  END S1
  PIN X
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.650000 0.440000  9.980000 1.820000 ;
        RECT 9.650000 1.820000 10.000000 2.980000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.560000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 10.560000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 10.560000 0.085000 ;
      RECT  0.000000  3.245000 10.560000 3.415000 ;
      RECT  0.095000  0.500000  0.465000 1.010000 ;
      RECT  0.095000  1.010000  0.265000 1.920000 ;
      RECT  0.095000  1.920000  0.585000 2.150000 ;
      RECT  0.255000  2.150000  0.585000 2.980000 ;
      RECT  0.755000  1.950000  1.085000 3.245000 ;
      RECT  0.820000  0.085000  1.150000 0.940000 ;
      RECT  1.850000  0.760000  2.665000 1.090000 ;
      RECT  2.045000  1.450000  2.325000 2.150000 ;
      RECT  2.495000  1.090000  2.665000 1.950000 ;
      RECT  2.495000  1.950000  4.285000 2.120000 ;
      RECT  2.495000  2.120000  3.445000 2.980000 ;
      RECT  3.445000  0.085000  3.925000 0.940000 ;
      RECT  3.615000  2.290000  3.945000 3.245000 ;
      RECT  4.115000  2.120000  4.285000 2.320000 ;
      RECT  4.115000  2.320000  5.605000 2.490000 ;
      RECT  4.530000  0.350000  5.105000 0.770000 ;
      RECT  4.530000  0.770000  8.015000 0.940000 ;
      RECT  4.925000  1.460000  5.265000 2.150000 ;
      RECT  5.055000  2.660000  5.945000 2.910000 ;
      RECT  5.435000  1.960000  7.080000 2.200000 ;
      RECT  5.435000  2.200000  5.605000 2.320000 ;
      RECT  5.775000  2.370000  7.980000 2.540000 ;
      RECT  5.775000  2.540000  5.945000 2.660000 ;
      RECT  6.140000  0.085000  6.470000 0.600000 ;
      RECT  6.165000  2.710000  6.495000 3.245000 ;
      RECT  6.560000  1.110000  7.955000 1.280000 ;
      RECT  6.560000  1.280000  6.730000 1.950000 ;
      RECT  6.560000  1.950000  7.080000 1.960000 ;
      RECT  6.690000  0.350000  6.940000 0.770000 ;
      RECT  7.120000  0.255000  9.130000 0.425000 ;
      RECT  7.120000  0.425000  7.450000 0.600000 ;
      RECT  7.200000  2.710000  7.530000 2.905000 ;
      RECT  7.200000  2.905000  9.130000 3.075000 ;
      RECT  7.650000  1.950000  7.980000 2.370000 ;
      RECT  7.725000  1.450000  8.450000 1.780000 ;
      RECT  7.810000  2.540000  7.980000 2.565000 ;
      RECT  7.810000  2.565000  8.790000 2.735000 ;
      RECT  7.845000  0.595000  8.790000 0.765000 ;
      RECT  7.845000  0.765000  8.015000 0.770000 ;
      RECT  8.185000  0.935000  8.450000 1.450000 ;
      RECT  8.200000  1.780000  8.450000 2.395000 ;
      RECT  8.620000  0.765000  8.790000 2.565000 ;
      RECT  8.960000  0.425000  9.130000 1.350000 ;
      RECT  8.960000  1.350000  9.385000 1.680000 ;
      RECT  8.960000  1.680000  9.130000 2.905000 ;
      RECT  9.300000  0.085000  9.470000 1.180000 ;
      RECT  9.300000  1.850000  9.470000 3.245000 ;
      RECT 10.160000  0.085000 10.410000 1.260000 ;
      RECT 10.200000  1.820000 10.450000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  1.950000  0.325000 2.120000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  1.950000  2.245000 2.120000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  1.950000  5.125000 2.120000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
    LAYER met1 ;
      RECT 0.095000 1.920000 0.385000 1.965000 ;
      RECT 0.095000 1.965000 5.185000 2.105000 ;
      RECT 0.095000 2.105000 0.385000 2.150000 ;
      RECT 2.015000 1.920000 2.305000 1.965000 ;
      RECT 2.015000 2.105000 2.305000 2.150000 ;
      RECT 4.895000 1.920000 5.185000 1.965000 ;
      RECT 4.895000 2.105000 5.185000 2.150000 ;
  END
END sky130_fd_sc_ls__mux4_2
END LIBRARY
