* File: sky130_fd_sc_ls__sdfxtp_2.pxi.spice
* Created: Fri Aug 28 14:05:42 2020
* 
x_PM_SKY130_FD_SC_LS__SDFXTP_2%A_27_74# N_A_27_74#_M1030_s N_A_27_74#_M1024_s
+ N_A_27_74#_M1014_g N_A_27_74#_c_234_n N_A_27_74#_M1006_g N_A_27_74#_c_230_n
+ N_A_27_74#_c_231_n N_A_27_74#_c_236_n N_A_27_74#_c_237_n N_A_27_74#_c_232_n
+ N_A_27_74#_c_233_n N_A_27_74#_c_239_n PM_SKY130_FD_SC_LS__SDFXTP_2%A_27_74#
x_PM_SKY130_FD_SC_LS__SDFXTP_2%SCE N_SCE_c_311_n N_SCE_c_320_n N_SCE_M1024_g
+ N_SCE_c_312_n N_SCE_M1030_g N_SCE_c_321_n N_SCE_c_322_n N_SCE_c_323_n
+ N_SCE_M1022_g N_SCE_c_313_n N_SCE_M1012_g N_SCE_c_314_n N_SCE_c_315_n SCE
+ N_SCE_c_316_n N_SCE_c_317_n N_SCE_c_318_n PM_SKY130_FD_SC_LS__SDFXTP_2%SCE
x_PM_SKY130_FD_SC_LS__SDFXTP_2%D N_D_c_398_n N_D_c_399_n N_D_M1013_g N_D_M1015_g
+ N_D_c_395_n N_D_c_401_n D N_D_c_396_n N_D_c_397_n
+ PM_SKY130_FD_SC_LS__SDFXTP_2%D
x_PM_SKY130_FD_SC_LS__SDFXTP_2%SCD N_SCD_M1000_g N_SCD_c_444_n N_SCD_M1017_g
+ N_SCD_c_441_n SCD SCD N_SCD_c_443_n PM_SKY130_FD_SC_LS__SDFXTP_2%SCD
x_PM_SKY130_FD_SC_LS__SDFXTP_2%CLK N_CLK_M1029_g N_CLK_c_486_n N_CLK_M1004_g CLK
+ N_CLK_c_484_n N_CLK_c_485_n PM_SKY130_FD_SC_LS__SDFXTP_2%CLK
x_PM_SKY130_FD_SC_LS__SDFXTP_2%A_846_74# N_A_846_74#_M1028_d N_A_846_74#_M1027_d
+ N_A_846_74#_c_548_n N_A_846_74#_M1026_g N_A_846_74#_M1002_g
+ N_A_846_74#_M1010_g N_A_846_74#_c_549_n N_A_846_74#_M1011_g
+ N_A_846_74#_c_550_n N_A_846_74#_c_529_n N_A_846_74#_c_530_n
+ N_A_846_74#_c_531_n N_A_846_74#_c_532_n N_A_846_74#_c_533_n
+ N_A_846_74#_c_534_n N_A_846_74#_c_535_n N_A_846_74#_c_536_n
+ N_A_846_74#_c_606_p N_A_846_74#_c_607_p N_A_846_74#_c_537_n
+ N_A_846_74#_c_538_n N_A_846_74#_c_539_n N_A_846_74#_c_540_n
+ N_A_846_74#_c_541_n N_A_846_74#_c_542_n N_A_846_74#_c_543_n
+ N_A_846_74#_c_639_p N_A_846_74#_c_544_n N_A_846_74#_c_545_n
+ N_A_846_74#_c_554_n N_A_846_74#_c_546_n N_A_846_74#_c_547_n
+ PM_SKY130_FD_SC_LS__SDFXTP_2%A_846_74#
x_PM_SKY130_FD_SC_LS__SDFXTP_2%A_634_74# N_A_634_74#_M1029_d N_A_634_74#_M1004_d
+ N_A_634_74#_c_720_n N_A_634_74#_M1028_g N_A_634_74#_c_736_n
+ N_A_634_74#_M1027_g N_A_634_74#_c_721_n N_A_634_74#_c_722_n
+ N_A_634_74#_M1033_g N_A_634_74#_c_724_n N_A_634_74#_c_725_n
+ N_A_634_74#_c_739_n N_A_634_74#_c_740_n N_A_634_74#_c_741_n
+ N_A_634_74#_M1031_g N_A_634_74#_c_726_n N_A_634_74#_M1025_g
+ N_A_634_74#_c_727_n N_A_634_74#_M1020_g N_A_634_74#_c_729_n
+ N_A_634_74#_c_730_n N_A_634_74#_c_731_n N_A_634_74#_c_744_n
+ N_A_634_74#_c_732_n N_A_634_74#_c_733_n N_A_634_74#_c_734_n
+ N_A_634_74#_c_746_n N_A_634_74#_c_820_p N_A_634_74#_c_747_n
+ N_A_634_74#_c_748_n N_A_634_74#_c_749_n N_A_634_74#_c_750_n
+ N_A_634_74#_c_735_n PM_SKY130_FD_SC_LS__SDFXTP_2%A_634_74#
x_PM_SKY130_FD_SC_LS__SDFXTP_2%A_1287_320# N_A_1287_320#_M1003_d
+ N_A_1287_320#_M1007_d N_A_1287_320#_c_943_n N_A_1287_320#_c_944_n
+ N_A_1287_320#_M1005_g N_A_1287_320#_M1008_g N_A_1287_320#_c_935_n
+ N_A_1287_320#_c_936_n N_A_1287_320#_c_937_n N_A_1287_320#_c_938_n
+ N_A_1287_320#_c_939_n N_A_1287_320#_c_940_n N_A_1287_320#_c_941_n
+ N_A_1287_320#_c_942_n PM_SKY130_FD_SC_LS__SDFXTP_2%A_1287_320#
x_PM_SKY130_FD_SC_LS__SDFXTP_2%A_1044_100# N_A_1044_100#_M1033_d
+ N_A_1044_100#_M1026_d N_A_1044_100#_c_1027_n N_A_1044_100#_M1007_g
+ N_A_1044_100#_c_1019_n N_A_1044_100#_M1003_g N_A_1044_100#_c_1020_n
+ N_A_1044_100#_c_1021_n N_A_1044_100#_c_1022_n N_A_1044_100#_c_1023_n
+ N_A_1044_100#_c_1024_n N_A_1044_100#_c_1029_n N_A_1044_100#_c_1030_n
+ N_A_1044_100#_c_1031_n N_A_1044_100#_c_1025_n N_A_1044_100#_c_1026_n
+ PM_SKY130_FD_SC_LS__SDFXTP_2%A_1044_100#
x_PM_SKY130_FD_SC_LS__SDFXTP_2%A_1829_398# N_A_1829_398#_M1016_d
+ N_A_1829_398#_M1018_d N_A_1829_398#_c_1124_n N_A_1829_398#_c_1137_n
+ N_A_1829_398#_c_1138_n N_A_1829_398#_M1032_g N_A_1829_398#_M1021_g
+ N_A_1829_398#_c_1126_n N_A_1829_398#_M1001_g N_A_1829_398#_c_1139_n
+ N_A_1829_398#_M1009_g N_A_1829_398#_c_1127_n N_A_1829_398#_M1023_g
+ N_A_1829_398#_c_1140_n N_A_1829_398#_M1019_g N_A_1829_398#_c_1128_n
+ N_A_1829_398#_c_1129_n N_A_1829_398#_c_1130_n N_A_1829_398#_c_1131_n
+ N_A_1829_398#_c_1132_n N_A_1829_398#_c_1133_n N_A_1829_398#_c_1134_n
+ N_A_1829_398#_c_1185_p N_A_1829_398#_c_1143_n N_A_1829_398#_c_1135_n
+ PM_SKY130_FD_SC_LS__SDFXTP_2%A_1829_398#
x_PM_SKY130_FD_SC_LS__SDFXTP_2%A_1592_424# N_A_1592_424#_M1010_d
+ N_A_1592_424#_M1025_d N_A_1592_424#_c_1227_n N_A_1592_424#_M1016_g
+ N_A_1592_424#_c_1228_n N_A_1592_424#_M1018_g N_A_1592_424#_c_1239_n
+ N_A_1592_424#_c_1229_n N_A_1592_424#_c_1234_n N_A_1592_424#_c_1235_n
+ N_A_1592_424#_c_1230_n N_A_1592_424#_c_1237_n N_A_1592_424#_c_1231_n
+ N_A_1592_424#_c_1238_n PM_SKY130_FD_SC_LS__SDFXTP_2%A_1592_424#
x_PM_SKY130_FD_SC_LS__SDFXTP_2%VPWR N_VPWR_M1024_d N_VPWR_M1017_d N_VPWR_M1027_s
+ N_VPWR_M1005_d N_VPWR_M1032_d N_VPWR_M1009_s N_VPWR_M1019_s N_VPWR_c_1316_n
+ N_VPWR_c_1317_n N_VPWR_c_1318_n N_VPWR_c_1319_n N_VPWR_c_1320_n
+ N_VPWR_c_1321_n N_VPWR_c_1322_n N_VPWR_c_1323_n N_VPWR_c_1324_n
+ N_VPWR_c_1325_n N_VPWR_c_1326_n VPWR N_VPWR_c_1327_n N_VPWR_c_1328_n
+ N_VPWR_c_1329_n N_VPWR_c_1330_n N_VPWR_c_1331_n N_VPWR_c_1332_n
+ N_VPWR_c_1333_n N_VPWR_c_1334_n N_VPWR_c_1335_n N_VPWR_c_1315_n
+ PM_SKY130_FD_SC_LS__SDFXTP_2%VPWR
x_PM_SKY130_FD_SC_LS__SDFXTP_2%A_300_453# N_A_300_453#_M1015_d
+ N_A_300_453#_M1033_s N_A_300_453#_M1013_d N_A_300_453#_M1026_s
+ N_A_300_453#_c_1452_n N_A_300_453#_c_1468_n N_A_300_453#_c_1453_n
+ N_A_300_453#_c_1454_n N_A_300_453#_c_1455_n N_A_300_453#_c_1456_n
+ N_A_300_453#_c_1462_n N_A_300_453#_c_1457_n N_A_300_453#_c_1458_n
+ N_A_300_453#_c_1514_n N_A_300_453#_c_1464_n N_A_300_453#_c_1459_n
+ N_A_300_453#_c_1465_n N_A_300_453#_c_1466_n N_A_300_453#_c_1508_n
+ N_A_300_453#_c_1544_n N_A_300_453#_c_1460_n
+ PM_SKY130_FD_SC_LS__SDFXTP_2%A_300_453#
x_PM_SKY130_FD_SC_LS__SDFXTP_2%Q N_Q_M1001_s N_Q_M1009_d N_Q_c_1590_n
+ N_Q_c_1596_n Q Q Q Q N_Q_c_1591_n PM_SKY130_FD_SC_LS__SDFXTP_2%Q
x_PM_SKY130_FD_SC_LS__SDFXTP_2%VGND N_VGND_M1030_d N_VGND_M1000_d N_VGND_M1028_s
+ N_VGND_M1008_d N_VGND_M1021_d N_VGND_M1001_d N_VGND_M1023_d N_VGND_c_1613_n
+ N_VGND_c_1614_n N_VGND_c_1615_n N_VGND_c_1616_n N_VGND_c_1617_n
+ N_VGND_c_1618_n N_VGND_c_1619_n N_VGND_c_1620_n N_VGND_c_1621_n
+ N_VGND_c_1622_n N_VGND_c_1623_n N_VGND_c_1624_n VGND N_VGND_c_1625_n
+ N_VGND_c_1626_n N_VGND_c_1627_n N_VGND_c_1628_n N_VGND_c_1629_n
+ N_VGND_c_1630_n N_VGND_c_1631_n N_VGND_c_1632_n N_VGND_c_1633_n
+ PM_SKY130_FD_SC_LS__SDFXTP_2%VGND
cc_1 VNB N_A_27_74#_M1014_g 0.0464673f $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=0.58
cc_2 VNB N_A_27_74#_c_230_n 0.0237434f $X=-0.19 $Y=-0.245 $X2=0.965 $Y2=1.635
cc_3 VNB N_A_27_74#_c_231_n 0.0317033f $X=-0.19 $Y=-0.245 $X2=0.17 $Y2=1.47
cc_4 VNB N_A_27_74#_c_232_n 0.0105324f $X=-0.19 $Y=-0.245 $X2=0.3 $Y2=0.555
cc_5 VNB N_A_27_74#_c_233_n 0.0101156f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=1.827
cc_6 VNB N_SCE_c_311_n 0.0257263f $X=-0.19 $Y=-0.245 $X2=0.135 $Y2=2.265
cc_7 VNB N_SCE_c_312_n 0.0225561f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_SCE_c_313_n 0.0190943f $X=-0.19 $Y=-0.245 $X2=0.965 $Y2=1.635
cc_9 VNB N_SCE_c_314_n 0.0204981f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_SCE_c_315_n 0.00565687f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=2.1
cc_11 VNB N_SCE_c_316_n 0.0490702f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.827
cc_12 VNB N_SCE_c_317_n 0.0363935f $X=-0.19 $Y=-0.245 $X2=2.045 $Y2=1.94
cc_13 VNB N_SCE_c_318_n 0.00826743f $X=-0.19 $Y=-0.245 $X2=2.045 $Y2=1.94
cc_14 VNB N_D_M1015_g 0.0337335f $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=0.58
cc_15 VNB N_D_c_395_n 0.0225791f $X=-0.19 $Y=-0.245 $X2=2.12 $Y2=2.585
cc_16 VNB N_D_c_396_n 0.0161693f $X=-0.19 $Y=-0.245 $X2=0.265 $Y2=2.185
cc_17 VNB N_D_c_397_n 0.0194658f $X=-0.19 $Y=-0.245 $X2=0.265 $Y2=2.41
cc_18 VNB N_SCD_M1000_g 0.0509958f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_SCD_c_441_n 0.00612749f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB SCD 0.00168234f $X=-0.19 $Y=-0.245 $X2=2.12 $Y2=2.19
cc_21 VNB N_SCD_c_443_n 0.0222454f $X=-0.19 $Y=-0.245 $X2=0.17 $Y2=1.47
cc_22 VNB N_CLK_M1029_g 0.0287628f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_CLK_c_484_n 0.0407916f $X=-0.19 $Y=-0.245 $X2=2.12 $Y2=2.19
cc_24 VNB N_CLK_c_485_n 0.00569067f $X=-0.19 $Y=-0.245 $X2=0.965 $Y2=1.635
cc_25 VNB N_A_846_74#_c_529_n 0.0110753f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_846_74#_c_530_n 0.0173473f $X=-0.19 $Y=-0.245 $X2=0.3 $Y2=0.555
cc_27 VNB N_A_846_74#_c_531_n 0.00279267f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_846_74#_c_532_n 0.00751998f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_846_74#_c_533_n 0.0241576f $X=-0.19 $Y=-0.245 $X2=0.265 $Y2=1.827
cc_30 VNB N_A_846_74#_c_534_n 7.97527e-19 $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.635
cc_31 VNB N_A_846_74#_c_535_n 0.00398981f $X=-0.19 $Y=-0.245 $X2=2.045 $Y2=1.94
cc_32 VNB N_A_846_74#_c_536_n 0.0351961f $X=-0.19 $Y=-0.245 $X2=2.045 $Y2=1.94
cc_33 VNB N_A_846_74#_c_537_n 0.00797819f $X=-0.19 $Y=-0.245 $X2=2.045 $Y2=1.94
cc_34 VNB N_A_846_74#_c_538_n 0.00246487f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_846_74#_c_539_n 0.00188696f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_846_74#_c_540_n 0.0105271f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_846_74#_c_541_n 0.00277883f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_846_74#_c_542_n 0.00701425f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_846_74#_c_543_n 0.00123754f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_846_74#_c_544_n 0.035006f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_846_74#_c_545_n 0.0066653f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_846_74#_c_546_n 0.0185456f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_846_74#_c_547_n 0.0209836f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_634_74#_c_720_n 0.0209609f $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=1.47
cc_45 VNB N_A_634_74#_c_721_n 0.0306611f $X=-0.19 $Y=-0.245 $X2=2.12 $Y2=2.585
cc_46 VNB N_A_634_74#_c_722_n 0.0913541f $X=-0.19 $Y=-0.245 $X2=0.965 $Y2=1.635
cc_47 VNB N_A_634_74#_M1033_g 0.0337086f $X=-0.19 $Y=-0.245 $X2=0.265 $Y2=2.185
cc_48 VNB N_A_634_74#_c_724_n 0.0354769f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.41
cc_49 VNB N_A_634_74#_c_725_n 0.0199077f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=2.1
cc_50 VNB N_A_634_74#_c_726_n 0.0161123f $X=-0.19 $Y=-0.245 $X2=0.17 $Y2=1.827
cc_51 VNB N_A_634_74#_c_727_n 0.026855f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.827
cc_52 VNB N_A_634_74#_M1020_g 0.0526436f $X=-0.19 $Y=-0.245 $X2=2.045 $Y2=1.94
cc_53 VNB N_A_634_74#_c_729_n 0.00487969f $X=-0.19 $Y=-0.245 $X2=2.045 $Y2=1.94
cc_54 VNB N_A_634_74#_c_730_n 0.00531483f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_634_74#_c_731_n 0.00653492f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_634_74#_c_732_n 0.0161092f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_634_74#_c_733_n 0.00162017f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_634_74#_c_734_n 3.8036e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_634_74#_c_735_n 0.00162437f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_1287_320#_M1008_g 0.0240304f $X=-0.19 $Y=-0.245 $X2=0.17 $Y2=1.47
cc_61 VNB N_A_1287_320#_c_935_n 0.0228992f $X=-0.19 $Y=-0.245 $X2=0.265 $Y2=2.41
cc_62 VNB N_A_1287_320#_c_936_n 0.00742455f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.41
cc_63 VNB N_A_1287_320#_c_937_n 0.0117738f $X=-0.19 $Y=-0.245 $X2=1.88 $Y2=2.1
cc_64 VNB N_A_1287_320#_c_938_n 0.00693555f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=2.1
cc_65 VNB N_A_1287_320#_c_939_n 0.0427778f $X=-0.19 $Y=-0.245 $X2=0.3 $Y2=0.515
cc_66 VNB N_A_1287_320#_c_940_n 0.0082105f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_1287_320#_c_941_n 0.00156076f $X=-0.19 $Y=-0.245 $X2=0.75
+ $Y2=1.635
cc_68 VNB N_A_1287_320#_c_942_n 0.0101f $X=-0.19 $Y=-0.245 $X2=2.045 $Y2=1.94
cc_69 VNB N_A_1044_100#_c_1019_n 0.0344813f $X=-0.19 $Y=-0.245 $X2=2.12 $Y2=2.19
cc_70 VNB N_A_1044_100#_c_1020_n 0.0203774f $X=-0.19 $Y=-0.245 $X2=0.17 $Y2=0.64
cc_71 VNB N_A_1044_100#_c_1021_n 0.0128169f $X=-0.19 $Y=-0.245 $X2=0.17 $Y2=1.47
cc_72 VNB N_A_1044_100#_c_1022_n 0.0166384f $X=-0.19 $Y=-0.245 $X2=0.265
+ $Y2=2.41
cc_73 VNB N_A_1044_100#_c_1023_n 0.0152439f $X=-0.19 $Y=-0.245 $X2=1.88 $Y2=2.1
cc_74 VNB N_A_1044_100#_c_1024_n 7.52377e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_1044_100#_c_1025_n 0.00236957f $X=-0.19 $Y=-0.245 $X2=0.75
+ $Y2=1.635
cc_76 VNB N_A_1044_100#_c_1026_n 0.0131463f $X=-0.19 $Y=-0.245 $X2=2.045 $Y2=2.1
cc_77 VNB N_A_1829_398#_c_1124_n 0.0122567f $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=1.47
cc_78 VNB N_A_1829_398#_M1021_g 0.0521092f $X=-0.19 $Y=-0.245 $X2=0.965
+ $Y2=1.635
cc_79 VNB N_A_1829_398#_c_1126_n 0.0192106f $X=-0.19 $Y=-0.245 $X2=0.17 $Y2=1.47
cc_80 VNB N_A_1829_398#_c_1127_n 0.0208149f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=2.1
cc_81 VNB N_A_1829_398#_c_1128_n 0.0646217f $X=-0.19 $Y=-0.245 $X2=0.17
+ $Y2=1.827
cc_82 VNB N_A_1829_398#_c_1129_n 0.0662148f $X=-0.19 $Y=-0.245 $X2=0.75
+ $Y2=1.827
cc_83 VNB N_A_1829_398#_c_1130_n 0.00292583f $X=-0.19 $Y=-0.245 $X2=2.045
+ $Y2=1.94
cc_84 VNB N_A_1829_398#_c_1131_n 0.00477515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_1829_398#_c_1132_n 0.00109972f $X=-0.19 $Y=-0.245 $X2=2.045
+ $Y2=2.1
cc_86 VNB N_A_1829_398#_c_1133_n 0.0140362f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_1829_398#_c_1134_n 0.0243141f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_1829_398#_c_1135_n 0.00206023f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_1592_424#_c_1227_n 0.0199771f $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=1.47
cc_90 VNB N_A_1592_424#_c_1228_n 0.0496836f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_1592_424#_c_1229_n 0.00586125f $X=-0.19 $Y=-0.245 $X2=0.17
+ $Y2=1.47
cc_92 VNB N_A_1592_424#_c_1230_n 0.00167757f $X=-0.19 $Y=-0.245 $X2=0.17
+ $Y2=0.515
cc_93 VNB N_A_1592_424#_c_1231_n 0.006113f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.635
cc_94 VNB N_VPWR_c_1315_n 0.502022f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_300_453#_c_1452_n 0.00687649f $X=-0.19 $Y=-0.245 $X2=2.12
+ $Y2=2.585
cc_96 VNB N_A_300_453#_c_1453_n 0.00203061f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_300_453#_c_1454_n 0.0114324f $X=-0.19 $Y=-0.245 $X2=1.88 $Y2=2.1
cc_98 VNB N_A_300_453#_c_1455_n 0.00530706f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=2.1
cc_99 VNB N_A_300_453#_c_1456_n 0.0032386f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_A_300_453#_c_1457_n 2.33396e-19 $X=-0.19 $Y=-0.245 $X2=0.17
+ $Y2=1.827
cc_101 VNB N_A_300_453#_c_1458_n 0.00559479f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_A_300_453#_c_1459_n 0.0056581f $X=-0.19 $Y=-0.245 $X2=0.915
+ $Y2=1.827
cc_103 VNB N_A_300_453#_c_1460_n 0.00724572f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_Q_c_1590_n 0.00280957f $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=0.58
cc_105 VNB N_Q_c_1591_n 0.0039544f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.635
cc_106 VNB N_VGND_c_1613_n 0.00649742f $X=-0.19 $Y=-0.245 $X2=0.3 $Y2=0.555
cc_107 VNB N_VGND_c_1614_n 0.00913749f $X=-0.19 $Y=-0.245 $X2=0.265 $Y2=1.827
cc_108 VNB N_VGND_c_1615_n 0.0140895f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=1.827
cc_109 VNB N_VGND_c_1616_n 0.0105681f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_1617_n 0.00751516f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_1618_n 0.011396f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_1619_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_1620_n 0.0543186f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_1621_n 0.0463653f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_VGND_c_1622_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_VGND_c_1623_n 0.0205017f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_VGND_c_1624_n 0.00634377f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_VGND_c_1625_n 0.0650416f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_VGND_c_1626_n 0.0568499f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_VGND_c_1627_n 0.0287187f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_VGND_c_1628_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_VGND_c_1629_n 0.0263788f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB N_VGND_c_1630_n 0.00631927f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_VGND_c_1631_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_1632_n 0.00519339f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_1633_n 0.652156f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VPB N_A_27_74#_c_234_n 0.0571826f $X=-0.19 $Y=1.66 $X2=2.12 $Y2=2.19
cc_128 VPB N_A_27_74#_c_230_n 0.0185473f $X=-0.19 $Y=1.66 $X2=0.965 $Y2=1.635
cc_129 VPB N_A_27_74#_c_236_n 0.0325133f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.41
cc_130 VPB N_A_27_74#_c_237_n 0.0239416f $X=-0.19 $Y=1.66 $X2=1.88 $Y2=2.1
cc_131 VPB N_A_27_74#_c_233_n 0.0243751f $X=-0.19 $Y=1.66 $X2=0.915 $Y2=1.827
cc_132 VPB N_A_27_74#_c_239_n 0.00536678f $X=-0.19 $Y=1.66 $X2=2.045 $Y2=1.94
cc_133 VPB N_SCE_c_311_n 0.0228022f $X=-0.19 $Y=1.66 $X2=0.135 $Y2=2.265
cc_134 VPB N_SCE_c_320_n 0.0191429f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_SCE_c_321_n 0.0203159f $X=-0.19 $Y=1.66 $X2=1.04 $Y2=0.58
cc_136 VPB N_SCE_c_322_n 0.0238116f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_SCE_c_323_n 0.0146453f $X=-0.19 $Y=1.66 $X2=2.12 $Y2=2.19
cc_138 VPB N_D_c_398_n 0.014901f $X=-0.19 $Y=1.66 $X2=0.135 $Y2=2.265
cc_139 VPB N_D_c_399_n 0.0223577f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_140 VPB N_D_c_395_n 0.00252529f $X=-0.19 $Y=1.66 $X2=2.12 $Y2=2.585
cc_141 VPB N_D_c_401_n 0.0157578f $X=-0.19 $Y=1.66 $X2=2.12 $Y2=2.585
cc_142 VPB N_D_c_397_n 0.0077491f $X=-0.19 $Y=1.66 $X2=0.265 $Y2=2.41
cc_143 VPB N_SCD_c_444_n 0.0167465f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_144 VPB N_SCD_c_441_n 0.048083f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_145 VPB SCD 0.00181008f $X=-0.19 $Y=1.66 $X2=2.12 $Y2=2.19
cc_146 VPB N_CLK_c_486_n 0.0192814f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_147 VPB N_CLK_c_484_n 0.0228698f $X=-0.19 $Y=1.66 $X2=2.12 $Y2=2.19
cc_148 VPB N_CLK_c_485_n 0.00418389f $X=-0.19 $Y=1.66 $X2=0.965 $Y2=1.635
cc_149 VPB N_A_846_74#_c_548_n 0.0189115f $X=-0.19 $Y=1.66 $X2=1.04 $Y2=1.47
cc_150 VPB N_A_846_74#_c_549_n 0.0635321f $X=-0.19 $Y=1.66 $X2=0.17 $Y2=1.47
cc_151 VPB N_A_846_74#_c_550_n 0.0518931f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_152 VPB N_A_846_74#_c_540_n 0.00506093f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_153 VPB N_A_846_74#_c_541_n 0.0143637f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_154 VPB N_A_846_74#_c_542_n 0.0325565f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_155 VPB N_A_846_74#_c_554_n 0.00382134f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_156 VPB N_A_634_74#_c_736_n 0.0208016f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_157 VPB N_A_634_74#_c_722_n 0.00856871f $X=-0.19 $Y=1.66 $X2=0.965 $Y2=1.635
cc_158 VPB N_A_634_74#_c_725_n 0.00394332f $X=-0.19 $Y=1.66 $X2=0.915 $Y2=2.1
cc_159 VPB N_A_634_74#_c_739_n 0.0329764f $X=-0.19 $Y=1.66 $X2=0.17 $Y2=0.515
cc_160 VPB N_A_634_74#_c_740_n 0.0188717f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_161 VPB N_A_634_74#_c_741_n 0.0434151f $X=-0.19 $Y=1.66 $X2=0.3 $Y2=0.515
cc_162 VPB N_A_634_74#_c_726_n 0.0503784f $X=-0.19 $Y=1.66 $X2=0.17 $Y2=1.827
cc_163 VPB N_A_634_74#_c_727_n 0.0340196f $X=-0.19 $Y=1.66 $X2=0.75 $Y2=1.827
cc_164 VPB N_A_634_74#_c_744_n 0.0119316f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_165 VPB N_A_634_74#_c_734_n 0.00489579f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_166 VPB N_A_634_74#_c_746_n 0.0161768f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_167 VPB N_A_634_74#_c_747_n 0.00450328f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_168 VPB N_A_634_74#_c_748_n 0.00171139f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_169 VPB N_A_634_74#_c_749_n 0.0015471f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_170 VPB N_A_634_74#_c_750_n 0.00593009f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_171 VPB N_A_634_74#_c_735_n 0.00356866f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_172 VPB N_A_1287_320#_c_943_n 0.0345231f $X=-0.19 $Y=1.66 $X2=1.04 $Y2=0.58
cc_173 VPB N_A_1287_320#_c_944_n 0.0246903f $X=-0.19 $Y=1.66 $X2=1.04 $Y2=0.58
cc_174 VPB N_A_1287_320#_c_936_n 0.00540297f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.41
cc_175 VPB N_A_1287_320#_c_940_n 0.00247539f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_176 VPB N_A_1044_100#_c_1027_n 0.0177828f $X=-0.19 $Y=1.66 $X2=1.04 $Y2=1.47
cc_177 VPB N_A_1044_100#_c_1023_n 0.00523956f $X=-0.19 $Y=1.66 $X2=1.88 $Y2=2.1
cc_178 VPB N_A_1044_100#_c_1029_n 8.77116e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_179 VPB N_A_1044_100#_c_1030_n 0.00526875f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_180 VPB N_A_1044_100#_c_1031_n 0.00684046f $X=-0.19 $Y=1.66 $X2=0.265
+ $Y2=1.827
cc_181 VPB N_A_1044_100#_c_1025_n 0.00249299f $X=-0.19 $Y=1.66 $X2=0.75
+ $Y2=1.635
cc_182 VPB N_A_1044_100#_c_1026_n 0.0560786f $X=-0.19 $Y=1.66 $X2=2.045 $Y2=2.1
cc_183 VPB N_A_1829_398#_c_1124_n 0.0395067f $X=-0.19 $Y=1.66 $X2=1.04 $Y2=1.47
cc_184 VPB N_A_1829_398#_c_1137_n 0.0147306f $X=-0.19 $Y=1.66 $X2=1.04 $Y2=0.58
cc_185 VPB N_A_1829_398#_c_1138_n 0.0265227f $X=-0.19 $Y=1.66 $X2=1.04 $Y2=0.58
cc_186 VPB N_A_1829_398#_c_1139_n 0.0165962f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.41
cc_187 VPB N_A_1829_398#_c_1140_n 0.0176406f $X=-0.19 $Y=1.66 $X2=0.3 $Y2=0.515
cc_188 VPB N_A_1829_398#_c_1129_n 0.0179937f $X=-0.19 $Y=1.66 $X2=0.75 $Y2=1.827
cc_189 VPB N_A_1829_398#_c_1130_n 0.00196261f $X=-0.19 $Y=1.66 $X2=2.045
+ $Y2=1.94
cc_190 VPB N_A_1829_398#_c_1143_n 0.00793483f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_191 VPB N_A_1829_398#_c_1135_n 0.0098712f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_192 VPB N_A_1592_424#_c_1228_n 0.0348307f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_193 VPB N_A_1592_424#_c_1229_n 0.00708854f $X=-0.19 $Y=1.66 $X2=0.17 $Y2=1.47
cc_194 VPB N_A_1592_424#_c_1234_n 0.00514681f $X=-0.19 $Y=1.66 $X2=0.265
+ $Y2=2.41
cc_195 VPB N_A_1592_424#_c_1235_n 0.0181622f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.41
cc_196 VPB N_A_1592_424#_c_1230_n 0.00112555f $X=-0.19 $Y=1.66 $X2=0.17
+ $Y2=0.515
cc_197 VPB N_A_1592_424#_c_1237_n 6.9017e-19 $X=-0.19 $Y=1.66 $X2=0.3 $Y2=0.555
cc_198 VPB N_A_1592_424#_c_1238_n 0.00143964f $X=-0.19 $Y=1.66 $X2=0.915
+ $Y2=1.827
cc_199 VPB N_VPWR_c_1316_n 0.010839f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_200 VPB N_VPWR_c_1317_n 0.0112503f $X=-0.19 $Y=1.66 $X2=0.17 $Y2=1.827
cc_201 VPB N_VPWR_c_1318_n 0.00796163f $X=-0.19 $Y=1.66 $X2=0.75 $Y2=1.635
cc_202 VPB N_VPWR_c_1319_n 0.0155378f $X=-0.19 $Y=1.66 $X2=2.045 $Y2=1.94
cc_203 VPB N_VPWR_c_1320_n 0.0229793f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_204 VPB N_VPWR_c_1321_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_205 VPB N_VPWR_c_1322_n 0.0645756f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_206 VPB N_VPWR_c_1323_n 0.0487271f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_207 VPB N_VPWR_c_1324_n 0.00862587f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_208 VPB N_VPWR_c_1325_n 0.0626084f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_209 VPB N_VPWR_c_1326_n 0.00460249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_210 VPB N_VPWR_c_1327_n 0.0191905f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_211 VPB N_VPWR_c_1328_n 0.0213889f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_212 VPB N_VPWR_c_1329_n 0.0649326f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_213 VPB N_VPWR_c_1330_n 0.0207499f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_214 VPB N_VPWR_c_1331_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_215 VPB N_VPWR_c_1332_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_216 VPB N_VPWR_c_1333_n 0.0219125f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_217 VPB N_VPWR_c_1334_n 0.012092f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_218 VPB N_VPWR_c_1335_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_219 VPB N_VPWR_c_1315_n 0.173093f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_220 VPB N_A_300_453#_c_1456_n 0.00221239f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_221 VPB N_A_300_453#_c_1462_n 0.00781763f $X=-0.19 $Y=1.66 $X2=0.3 $Y2=0.515
cc_222 VPB N_A_300_453#_c_1457_n 0.00162545f $X=-0.19 $Y=1.66 $X2=0.17 $Y2=1.827
cc_223 VPB N_A_300_453#_c_1464_n 0.00982402f $X=-0.19 $Y=1.66 $X2=0.75 $Y2=1.827
cc_224 VPB N_A_300_453#_c_1465_n 0.00767653f $X=-0.19 $Y=1.66 $X2=2.045 $Y2=1.94
cc_225 VPB N_A_300_453#_c_1466_n 0.00522047f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_226 VPB Q 0.00696915f $X=-0.19 $Y=1.66 $X2=0.965 $Y2=1.635
cc_227 VPB N_Q_c_1591_n 0.0025253f $X=-0.19 $Y=1.66 $X2=0.75 $Y2=1.635
cc_228 N_A_27_74#_M1014_g N_SCE_c_311_n 0.00365204f $X=1.04 $Y=0.58 $X2=0 $Y2=0
cc_229 N_A_27_74#_c_230_n N_SCE_c_311_n 0.0181319f $X=0.965 $Y=1.635 $X2=0 $Y2=0
cc_230 N_A_27_74#_c_231_n N_SCE_c_311_n 0.0150312f $X=0.17 $Y=1.47 $X2=0 $Y2=0
cc_231 N_A_27_74#_c_233_n N_SCE_c_311_n 0.0287559f $X=0.915 $Y=1.827 $X2=0 $Y2=0
cc_232 N_A_27_74#_c_236_n N_SCE_c_320_n 0.0105826f $X=0.28 $Y=2.41 $X2=0 $Y2=0
cc_233 N_A_27_74#_M1014_g N_SCE_c_312_n 0.015292f $X=1.04 $Y=0.58 $X2=0 $Y2=0
cc_234 N_A_27_74#_c_231_n N_SCE_c_312_n 0.00439162f $X=0.17 $Y=1.47 $X2=0 $Y2=0
cc_235 N_A_27_74#_c_232_n N_SCE_c_312_n 0.00316265f $X=0.3 $Y=0.555 $X2=0 $Y2=0
cc_236 N_A_27_74#_c_230_n N_SCE_c_321_n 0.0281061f $X=0.965 $Y=1.635 $X2=0 $Y2=0
cc_237 N_A_27_74#_c_237_n N_SCE_c_321_n 0.0113305f $X=1.88 $Y=2.1 $X2=0 $Y2=0
cc_238 N_A_27_74#_c_233_n N_SCE_c_321_n 0.0124644f $X=0.915 $Y=1.827 $X2=0 $Y2=0
cc_239 N_A_27_74#_c_236_n N_SCE_c_322_n 0.00703504f $X=0.28 $Y=2.41 $X2=0 $Y2=0
cc_240 N_A_27_74#_c_233_n N_SCE_c_322_n 0.0208969f $X=0.915 $Y=1.827 $X2=0 $Y2=0
cc_241 N_A_27_74#_c_236_n N_SCE_c_323_n 6.93314e-19 $X=0.28 $Y=2.41 $X2=0 $Y2=0
cc_242 N_A_27_74#_M1014_g N_SCE_c_314_n 0.0148534f $X=1.04 $Y=0.58 $X2=0 $Y2=0
cc_243 N_A_27_74#_c_230_n N_SCE_c_314_n 0.00283648f $X=0.965 $Y=1.635 $X2=0
+ $Y2=0
cc_244 N_A_27_74#_c_233_n N_SCE_c_314_n 0.00305183f $X=0.915 $Y=1.827 $X2=0
+ $Y2=0
cc_245 N_A_27_74#_c_234_n N_SCE_c_315_n 3.65439e-19 $X=2.12 $Y=2.19 $X2=0 $Y2=0
cc_246 N_A_27_74#_c_239_n N_SCE_c_315_n 0.00961704f $X=2.045 $Y=1.94 $X2=0 $Y2=0
cc_247 N_A_27_74#_M1014_g N_SCE_c_316_n 0.020149f $X=1.04 $Y=0.58 $X2=0 $Y2=0
cc_248 N_A_27_74#_c_230_n N_SCE_c_316_n 0.00889754f $X=0.965 $Y=1.635 $X2=0
+ $Y2=0
cc_249 N_A_27_74#_c_231_n N_SCE_c_316_n 0.00789794f $X=0.17 $Y=1.47 $X2=0 $Y2=0
cc_250 N_A_27_74#_c_232_n N_SCE_c_316_n 0.00501366f $X=0.3 $Y=0.555 $X2=0 $Y2=0
cc_251 N_A_27_74#_c_233_n N_SCE_c_316_n 0.00770903f $X=0.915 $Y=1.827 $X2=0
+ $Y2=0
cc_252 N_A_27_74#_c_234_n N_SCE_c_317_n 0.00551385f $X=2.12 $Y=2.19 $X2=0 $Y2=0
cc_253 N_A_27_74#_c_239_n N_SCE_c_317_n 3.97776e-19 $X=2.045 $Y=1.94 $X2=0 $Y2=0
cc_254 N_A_27_74#_M1014_g N_SCE_c_318_n 0.00557782f $X=1.04 $Y=0.58 $X2=0 $Y2=0
cc_255 N_A_27_74#_c_230_n N_SCE_c_318_n 0.00238461f $X=0.965 $Y=1.635 $X2=0
+ $Y2=0
cc_256 N_A_27_74#_c_231_n N_SCE_c_318_n 0.0324652f $X=0.17 $Y=1.47 $X2=0 $Y2=0
cc_257 N_A_27_74#_c_232_n N_SCE_c_318_n 0.00341317f $X=0.3 $Y=0.555 $X2=0 $Y2=0
cc_258 N_A_27_74#_c_233_n N_SCE_c_318_n 0.0263644f $X=0.915 $Y=1.827 $X2=0 $Y2=0
cc_259 N_A_27_74#_c_234_n N_D_c_398_n 0.00851487f $X=2.12 $Y=2.19 $X2=0 $Y2=0
cc_260 N_A_27_74#_c_237_n N_D_c_398_n 0.00624901f $X=1.88 $Y=2.1 $X2=0 $Y2=0
cc_261 N_A_27_74#_c_239_n N_D_c_398_n 9.91144e-19 $X=2.045 $Y=1.94 $X2=0 $Y2=0
cc_262 N_A_27_74#_c_234_n N_D_c_399_n 0.0183105f $X=2.12 $Y=2.19 $X2=0 $Y2=0
cc_263 N_A_27_74#_c_237_n N_D_c_399_n 0.0104204f $X=1.88 $Y=2.1 $X2=0 $Y2=0
cc_264 N_A_27_74#_M1014_g N_D_M1015_g 0.050486f $X=1.04 $Y=0.58 $X2=0 $Y2=0
cc_265 N_A_27_74#_c_230_n N_D_c_395_n 0.0186275f $X=0.965 $Y=1.635 $X2=0 $Y2=0
cc_266 N_A_27_74#_c_234_n N_D_c_401_n 0.00527201f $X=2.12 $Y=2.19 $X2=0 $Y2=0
cc_267 N_A_27_74#_c_237_n N_D_c_401_n 0.00396341f $X=1.88 $Y=2.1 $X2=0 $Y2=0
cc_268 N_A_27_74#_c_233_n N_D_c_401_n 0.00570978f $X=0.915 $Y=1.827 $X2=0 $Y2=0
cc_269 N_A_27_74#_c_239_n N_D_c_401_n 2.01112e-19 $X=2.045 $Y=1.94 $X2=0 $Y2=0
cc_270 N_A_27_74#_M1014_g N_D_c_396_n 0.0186275f $X=1.04 $Y=0.58 $X2=0 $Y2=0
cc_271 N_A_27_74#_M1014_g N_D_c_397_n 0.0147252f $X=1.04 $Y=0.58 $X2=0 $Y2=0
cc_272 N_A_27_74#_c_234_n N_D_c_397_n 2.42546e-19 $X=2.12 $Y=2.19 $X2=0 $Y2=0
cc_273 N_A_27_74#_c_230_n N_D_c_397_n 0.00914129f $X=0.965 $Y=1.635 $X2=0 $Y2=0
cc_274 N_A_27_74#_c_237_n N_D_c_397_n 0.0464516f $X=1.88 $Y=2.1 $X2=0 $Y2=0
cc_275 N_A_27_74#_c_233_n N_D_c_397_n 0.031591f $X=0.915 $Y=1.827 $X2=0 $Y2=0
cc_276 N_A_27_74#_c_239_n N_D_c_397_n 0.0045026f $X=2.045 $Y=1.94 $X2=0 $Y2=0
cc_277 N_A_27_74#_c_234_n N_SCD_c_444_n 0.0402063f $X=2.12 $Y=2.19 $X2=0 $Y2=0
cc_278 N_A_27_74#_c_234_n N_SCD_c_441_n 0.0213601f $X=2.12 $Y=2.19 $X2=0 $Y2=0
cc_279 N_A_27_74#_c_239_n N_SCD_c_441_n 0.00159042f $X=2.045 $Y=1.94 $X2=0 $Y2=0
cc_280 N_A_27_74#_c_234_n SCD 0.00136225f $X=2.12 $Y=2.19 $X2=0 $Y2=0
cc_281 N_A_27_74#_c_239_n SCD 0.0213355f $X=2.045 $Y=1.94 $X2=0 $Y2=0
cc_282 N_A_27_74#_c_236_n N_VPWR_c_1316_n 0.022465f $X=0.28 $Y=2.41 $X2=0 $Y2=0
cc_283 N_A_27_74#_c_233_n N_VPWR_c_1316_n 0.0247451f $X=0.915 $Y=1.827 $X2=0
+ $Y2=0
cc_284 N_A_27_74#_c_234_n N_VPWR_c_1323_n 0.00416979f $X=2.12 $Y=2.19 $X2=0
+ $Y2=0
cc_285 N_A_27_74#_c_236_n N_VPWR_c_1327_n 0.0130353f $X=0.28 $Y=2.41 $X2=0 $Y2=0
cc_286 N_A_27_74#_c_234_n N_VPWR_c_1315_n 0.00528353f $X=2.12 $Y=2.19 $X2=0
+ $Y2=0
cc_287 N_A_27_74#_c_236_n N_VPWR_c_1315_n 0.0127617f $X=0.28 $Y=2.41 $X2=0 $Y2=0
cc_288 N_A_27_74#_M1014_g N_A_300_453#_c_1452_n 0.00100617f $X=1.04 $Y=0.58
+ $X2=0 $Y2=0
cc_289 N_A_27_74#_c_234_n N_A_300_453#_c_1468_n 0.0121528f $X=2.12 $Y=2.19 $X2=0
+ $Y2=0
cc_290 N_A_27_74#_c_239_n N_A_300_453#_c_1468_n 0.0107328f $X=2.045 $Y=1.94
+ $X2=0 $Y2=0
cc_291 N_A_27_74#_c_234_n N_A_300_453#_c_1466_n 0.0191923f $X=2.12 $Y=2.19 $X2=0
+ $Y2=0
cc_292 N_A_27_74#_c_237_n N_A_300_453#_c_1466_n 0.0295592f $X=1.88 $Y=2.1 $X2=0
+ $Y2=0
cc_293 N_A_27_74#_c_239_n N_A_300_453#_c_1466_n 0.0129086f $X=2.045 $Y=1.94
+ $X2=0 $Y2=0
cc_294 N_A_27_74#_M1014_g N_VGND_c_1613_n 0.0091955f $X=1.04 $Y=0.58 $X2=0 $Y2=0
cc_295 N_A_27_74#_M1014_g N_VGND_c_1621_n 0.00383152f $X=1.04 $Y=0.58 $X2=0
+ $Y2=0
cc_296 N_A_27_74#_c_232_n N_VGND_c_1629_n 0.0132203f $X=0.3 $Y=0.555 $X2=0 $Y2=0
cc_297 N_A_27_74#_M1014_g N_VGND_c_1633_n 0.00385768f $X=1.04 $Y=0.58 $X2=0
+ $Y2=0
cc_298 N_A_27_74#_c_232_n N_VGND_c_1633_n 0.0139586f $X=0.3 $Y=0.555 $X2=0 $Y2=0
cc_299 N_SCE_c_321_n N_D_c_398_n 0.00830278f $X=0.93 $Y=2.115 $X2=0 $Y2=0
cc_300 N_SCE_c_323_n N_D_c_399_n 0.037892f $X=1.005 $Y=2.19 $X2=0 $Y2=0
cc_301 N_SCE_c_313_n N_D_M1015_g 0.0136155f $X=2.135 $Y=0.9 $X2=0 $Y2=0
cc_302 N_SCE_c_314_n N_D_M1015_g 0.0119168f $X=1.875 $Y=0.935 $X2=0 $Y2=0
cc_303 N_SCE_c_315_n N_D_M1015_g 0.00112165f $X=2.04 $Y=0.935 $X2=0 $Y2=0
cc_304 N_SCE_c_317_n N_D_M1015_g 0.00981569f $X=2.135 $Y=1.065 $X2=0 $Y2=0
cc_305 N_SCE_c_314_n N_D_c_396_n 0.00468585f $X=1.875 $Y=0.935 $X2=0 $Y2=0
cc_306 N_SCE_c_317_n N_D_c_396_n 0.00253031f $X=2.135 $Y=1.065 $X2=0 $Y2=0
cc_307 N_SCE_c_314_n N_D_c_397_n 0.0463166f $X=1.875 $Y=0.935 $X2=0 $Y2=0
cc_308 N_SCE_c_315_n N_D_c_397_n 0.0025934f $X=2.04 $Y=0.935 $X2=0 $Y2=0
cc_309 N_SCE_c_318_n N_D_c_397_n 0.00240592f $X=0.835 $Y=1.02 $X2=0 $Y2=0
cc_310 N_SCE_c_313_n N_SCD_M1000_g 0.0522534f $X=2.135 $Y=0.9 $X2=0 $Y2=0
cc_311 N_SCE_c_315_n N_SCD_M1000_g 4.19134e-19 $X=2.04 $Y=0.935 $X2=0 $Y2=0
cc_312 N_SCE_c_320_n N_VPWR_c_1316_n 0.00625754f $X=0.505 $Y=2.19 $X2=0 $Y2=0
cc_313 N_SCE_c_321_n N_VPWR_c_1316_n 0.0034144f $X=0.93 $Y=2.115 $X2=0 $Y2=0
cc_314 N_SCE_c_323_n N_VPWR_c_1316_n 0.0135831f $X=1.005 $Y=2.19 $X2=0 $Y2=0
cc_315 N_SCE_c_323_n N_VPWR_c_1323_n 0.0048289f $X=1.005 $Y=2.19 $X2=0 $Y2=0
cc_316 N_SCE_c_320_n N_VPWR_c_1327_n 0.00523995f $X=0.505 $Y=2.19 $X2=0 $Y2=0
cc_317 N_SCE_c_320_n N_VPWR_c_1315_n 0.00528353f $X=0.505 $Y=2.19 $X2=0 $Y2=0
cc_318 N_SCE_c_323_n N_VPWR_c_1315_n 0.0047904f $X=1.005 $Y=2.19 $X2=0 $Y2=0
cc_319 N_SCE_c_313_n N_A_300_453#_c_1452_n 0.0178483f $X=2.135 $Y=0.9 $X2=0
+ $Y2=0
cc_320 N_SCE_c_314_n N_A_300_453#_c_1452_n 0.0275614f $X=1.875 $Y=0.935 $X2=0
+ $Y2=0
cc_321 N_SCE_c_315_n N_A_300_453#_c_1452_n 0.0233279f $X=2.04 $Y=0.935 $X2=0
+ $Y2=0
cc_322 N_SCE_c_317_n N_A_300_453#_c_1452_n 0.00105893f $X=2.135 $Y=1.065 $X2=0
+ $Y2=0
cc_323 N_SCE_c_313_n N_A_300_453#_c_1453_n 0.00481728f $X=2.135 $Y=0.9 $X2=0
+ $Y2=0
cc_324 N_SCE_c_315_n N_A_300_453#_c_1453_n 0.0183381f $X=2.04 $Y=0.935 $X2=0
+ $Y2=0
cc_325 N_SCE_c_315_n N_A_300_453#_c_1455_n 0.0113849f $X=2.04 $Y=0.935 $X2=0
+ $Y2=0
cc_326 N_SCE_c_317_n N_A_300_453#_c_1455_n 8.92401e-19 $X=2.135 $Y=1.065 $X2=0
+ $Y2=0
cc_327 N_SCE_c_323_n N_A_300_453#_c_1466_n 0.00169591f $X=1.005 $Y=2.19 $X2=0
+ $Y2=0
cc_328 N_SCE_c_312_n N_VGND_c_1613_n 0.00504481f $X=0.54 $Y=0.9 $X2=0 $Y2=0
cc_329 N_SCE_c_314_n N_VGND_c_1613_n 0.00809823f $X=1.875 $Y=0.935 $X2=0 $Y2=0
cc_330 N_SCE_c_316_n N_VGND_c_1613_n 5.64633e-19 $X=0.54 $Y=1.065 $X2=0 $Y2=0
cc_331 N_SCE_c_318_n N_VGND_c_1613_n 0.0144474f $X=0.835 $Y=1.02 $X2=0 $Y2=0
cc_332 N_SCE_c_313_n N_VGND_c_1621_n 0.00291649f $X=2.135 $Y=0.9 $X2=0 $Y2=0
cc_333 N_SCE_c_312_n N_VGND_c_1629_n 0.00434051f $X=0.54 $Y=0.9 $X2=0 $Y2=0
cc_334 N_SCE_c_312_n N_VGND_c_1633_n 0.00444892f $X=0.54 $Y=0.9 $X2=0 $Y2=0
cc_335 N_SCE_c_313_n N_VGND_c_1633_n 0.0036095f $X=2.135 $Y=0.9 $X2=0 $Y2=0
cc_336 N_SCE_c_314_n N_VGND_c_1633_n 0.01609f $X=1.875 $Y=0.935 $X2=0 $Y2=0
cc_337 N_SCE_c_318_n N_VGND_c_1633_n 0.00638792f $X=0.835 $Y=1.02 $X2=0 $Y2=0
cc_338 N_D_c_399_n N_VPWR_c_1316_n 0.00213493f $X=1.425 $Y=2.19 $X2=0 $Y2=0
cc_339 N_D_c_399_n N_VPWR_c_1323_n 0.00523782f $X=1.425 $Y=2.19 $X2=0 $Y2=0
cc_340 N_D_c_399_n N_VPWR_c_1315_n 0.00528353f $X=1.425 $Y=2.19 $X2=0 $Y2=0
cc_341 N_D_M1015_g N_A_300_453#_c_1452_n 0.0122799f $X=1.43 $Y=0.58 $X2=0 $Y2=0
cc_342 N_D_c_399_n N_A_300_453#_c_1466_n 0.0212042f $X=1.425 $Y=2.19 $X2=0 $Y2=0
cc_343 N_D_M1015_g N_VGND_c_1613_n 0.00138367f $X=1.43 $Y=0.58 $X2=0 $Y2=0
cc_344 N_D_M1015_g N_VGND_c_1621_n 0.00433162f $X=1.43 $Y=0.58 $X2=0 $Y2=0
cc_345 N_D_M1015_g N_VGND_c_1633_n 0.00450914f $X=1.43 $Y=0.58 $X2=0 $Y2=0
cc_346 N_SCD_M1000_g N_CLK_M1029_g 0.023592f $X=2.525 $Y=0.58 $X2=0 $Y2=0
cc_347 N_SCD_c_444_n N_CLK_c_486_n 0.0125849f $X=2.54 $Y=2.19 $X2=0 $Y2=0
cc_348 N_SCD_c_441_n N_CLK_c_486_n 0.00799165f $X=2.615 $Y=1.94 $X2=0 $Y2=0
cc_349 N_SCD_c_441_n N_CLK_c_484_n 0.00184988f $X=2.615 $Y=1.94 $X2=0 $Y2=0
cc_350 SCD N_CLK_c_484_n 2.68407e-19 $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_351 N_SCD_c_443_n N_CLK_c_484_n 0.0129251f $X=2.615 $Y=1.6 $X2=0 $Y2=0
cc_352 N_SCD_M1000_g N_A_634_74#_c_730_n 3.49205e-19 $X=2.525 $Y=0.58 $X2=0
+ $Y2=0
cc_353 N_SCD_c_444_n N_VPWR_c_1317_n 0.00561084f $X=2.54 $Y=2.19 $X2=0 $Y2=0
cc_354 N_SCD_c_444_n N_VPWR_c_1323_n 0.00419287f $X=2.54 $Y=2.19 $X2=0 $Y2=0
cc_355 N_SCD_c_444_n N_VPWR_c_1315_n 0.00528353f $X=2.54 $Y=2.19 $X2=0 $Y2=0
cc_356 N_SCD_M1000_g N_A_300_453#_c_1452_n 0.00927742f $X=2.525 $Y=0.58 $X2=0
+ $Y2=0
cc_357 N_SCD_c_444_n N_A_300_453#_c_1468_n 0.0174367f $X=2.54 $Y=2.19 $X2=0
+ $Y2=0
cc_358 N_SCD_c_441_n N_A_300_453#_c_1468_n 8.24906e-19 $X=2.615 $Y=1.94 $X2=0
+ $Y2=0
cc_359 SCD N_A_300_453#_c_1468_n 0.0210048f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_360 N_SCD_M1000_g N_A_300_453#_c_1453_n 0.010612f $X=2.525 $Y=0.58 $X2=0
+ $Y2=0
cc_361 N_SCD_M1000_g N_A_300_453#_c_1454_n 0.00663453f $X=2.525 $Y=0.58 $X2=0
+ $Y2=0
cc_362 SCD N_A_300_453#_c_1454_n 0.0185361f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_363 N_SCD_c_443_n N_A_300_453#_c_1454_n 0.00124629f $X=2.615 $Y=1.6 $X2=0
+ $Y2=0
cc_364 N_SCD_M1000_g N_A_300_453#_c_1455_n 0.00402007f $X=2.525 $Y=0.58 $X2=0
+ $Y2=0
cc_365 SCD N_A_300_453#_c_1455_n 0.00798768f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_366 N_SCD_M1000_g N_A_300_453#_c_1456_n 0.0029973f $X=2.525 $Y=0.58 $X2=0
+ $Y2=0
cc_367 N_SCD_c_444_n N_A_300_453#_c_1456_n 0.00315112f $X=2.54 $Y=2.19 $X2=0
+ $Y2=0
cc_368 N_SCD_c_441_n N_A_300_453#_c_1456_n 9.09006e-19 $X=2.615 $Y=1.94 $X2=0
+ $Y2=0
cc_369 SCD N_A_300_453#_c_1456_n 0.0534381f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_370 N_SCD_c_443_n N_A_300_453#_c_1456_n 0.00474092f $X=2.615 $Y=1.6 $X2=0
+ $Y2=0
cc_371 N_SCD_c_444_n N_A_300_453#_c_1466_n 0.00139235f $X=2.54 $Y=2.19 $X2=0
+ $Y2=0
cc_372 N_SCD_M1000_g N_VGND_c_1614_n 0.00645761f $X=2.525 $Y=0.58 $X2=0 $Y2=0
cc_373 N_SCD_M1000_g N_VGND_c_1621_n 0.00353828f $X=2.525 $Y=0.58 $X2=0 $Y2=0
cc_374 N_SCD_M1000_g N_VGND_c_1633_n 0.00561756f $X=2.525 $Y=0.58 $X2=0 $Y2=0
cc_375 N_CLK_M1029_g N_A_634_74#_c_722_n 0.00276249f $X=3.095 $Y=0.74 $X2=0
+ $Y2=0
cc_376 N_CLK_c_484_n N_A_634_74#_c_722_n 0.0180073f $X=3.28 $Y=1.557 $X2=0 $Y2=0
cc_377 N_CLK_c_485_n N_A_634_74#_c_722_n 0.00187012f $X=3.455 $Y=1.515 $X2=0
+ $Y2=0
cc_378 N_CLK_M1029_g N_A_634_74#_c_730_n 0.0105679f $X=3.095 $Y=0.74 $X2=0 $Y2=0
cc_379 N_CLK_c_484_n N_A_634_74#_c_730_n 0.00469055f $X=3.28 $Y=1.557 $X2=0
+ $Y2=0
cc_380 N_CLK_c_485_n N_A_634_74#_c_730_n 0.0152412f $X=3.455 $Y=1.515 $X2=0
+ $Y2=0
cc_381 N_CLK_M1029_g N_A_634_74#_c_731_n 0.0053769f $X=3.095 $Y=0.74 $X2=0 $Y2=0
cc_382 N_CLK_c_486_n N_A_634_74#_c_744_n 0.00403724f $X=3.28 $Y=1.765 $X2=0
+ $Y2=0
cc_383 N_CLK_c_484_n N_A_634_74#_c_744_n 0.00134694f $X=3.28 $Y=1.557 $X2=0
+ $Y2=0
cc_384 N_CLK_c_485_n N_A_634_74#_c_744_n 0.0264522f $X=3.455 $Y=1.515 $X2=0
+ $Y2=0
cc_385 N_CLK_c_484_n N_A_634_74#_c_732_n 0.00101999f $X=3.28 $Y=1.557 $X2=0
+ $Y2=0
cc_386 N_CLK_c_485_n N_A_634_74#_c_732_n 0.0163452f $X=3.455 $Y=1.515 $X2=0
+ $Y2=0
cc_387 N_CLK_M1029_g N_A_634_74#_c_733_n 0.00140815f $X=3.095 $Y=0.74 $X2=0
+ $Y2=0
cc_388 N_CLK_c_485_n N_A_634_74#_c_733_n 0.00759441f $X=3.455 $Y=1.515 $X2=0
+ $Y2=0
cc_389 N_CLK_c_486_n N_A_634_74#_c_734_n 0.00407092f $X=3.28 $Y=1.765 $X2=0
+ $Y2=0
cc_390 N_CLK_c_484_n N_A_634_74#_c_734_n 8.20654e-19 $X=3.28 $Y=1.557 $X2=0
+ $Y2=0
cc_391 N_CLK_c_485_n N_A_634_74#_c_734_n 0.0272207f $X=3.455 $Y=1.515 $X2=0
+ $Y2=0
cc_392 N_CLK_c_486_n N_VPWR_c_1317_n 0.0101043f $X=3.28 $Y=1.765 $X2=0 $Y2=0
cc_393 N_CLK_c_486_n N_VPWR_c_1328_n 0.00334059f $X=3.28 $Y=1.765 $X2=0 $Y2=0
cc_394 N_CLK_c_486_n N_VPWR_c_1333_n 0.00781345f $X=3.28 $Y=1.765 $X2=0 $Y2=0
cc_395 N_CLK_c_486_n N_VPWR_c_1315_n 0.00441457f $X=3.28 $Y=1.765 $X2=0 $Y2=0
cc_396 N_CLK_M1029_g N_A_300_453#_c_1453_n 0.00131902f $X=3.095 $Y=0.74 $X2=0
+ $Y2=0
cc_397 N_CLK_M1029_g N_A_300_453#_c_1454_n 0.0137646f $X=3.095 $Y=0.74 $X2=0
+ $Y2=0
cc_398 N_CLK_M1029_g N_A_300_453#_c_1456_n 0.00452193f $X=3.095 $Y=0.74 $X2=0
+ $Y2=0
cc_399 N_CLK_c_486_n N_A_300_453#_c_1456_n 0.00954243f $X=3.28 $Y=1.765 $X2=0
+ $Y2=0
cc_400 N_CLK_c_484_n N_A_300_453#_c_1456_n 0.0125263f $X=3.28 $Y=1.557 $X2=0
+ $Y2=0
cc_401 N_CLK_c_485_n N_A_300_453#_c_1456_n 0.0314924f $X=3.455 $Y=1.515 $X2=0
+ $Y2=0
cc_402 N_CLK_c_486_n N_A_300_453#_c_1462_n 0.0186435f $X=3.28 $Y=1.765 $X2=0
+ $Y2=0
cc_403 N_CLK_c_485_n N_A_300_453#_c_1462_n 0.00113812f $X=3.455 $Y=1.515 $X2=0
+ $Y2=0
cc_404 N_CLK_c_486_n N_A_300_453#_c_1508_n 0.00322164f $X=3.28 $Y=1.765 $X2=0
+ $Y2=0
cc_405 N_CLK_M1029_g N_VGND_c_1614_n 0.00316386f $X=3.095 $Y=0.74 $X2=0 $Y2=0
cc_406 N_CLK_M1029_g N_VGND_c_1615_n 0.00319982f $X=3.095 $Y=0.74 $X2=0 $Y2=0
cc_407 N_CLK_M1029_g N_VGND_c_1623_n 0.00433834f $X=3.095 $Y=0.74 $X2=0 $Y2=0
cc_408 N_CLK_M1029_g N_VGND_c_1633_n 0.00826005f $X=3.095 $Y=0.74 $X2=0 $Y2=0
cc_409 N_A_846_74#_c_529_n N_A_634_74#_c_720_n 0.0158581f $X=4.37 $Y=0.515 $X2=0
+ $Y2=0
cc_410 N_A_846_74#_c_531_n N_A_634_74#_c_720_n 0.00469864f $X=4.535 $Y=0.34
+ $X2=0 $Y2=0
cc_411 N_A_846_74#_c_541_n N_A_634_74#_c_736_n 0.00238041f $X=5.21 $Y=1.775
+ $X2=0 $Y2=0
cc_412 N_A_846_74#_c_542_n N_A_634_74#_c_736_n 0.0070157f $X=5.21 $Y=1.775 $X2=0
+ $Y2=0
cc_413 N_A_846_74#_c_541_n N_A_634_74#_c_721_n 0.00734434f $X=5.21 $Y=1.775
+ $X2=0 $Y2=0
cc_414 N_A_846_74#_c_542_n N_A_634_74#_c_721_n 0.0182849f $X=5.21 $Y=1.775 $X2=0
+ $Y2=0
cc_415 N_A_846_74#_c_529_n N_A_634_74#_c_722_n 0.00605381f $X=4.37 $Y=0.515
+ $X2=0 $Y2=0
cc_416 N_A_846_74#_c_532_n N_A_634_74#_c_722_n 0.00417255f $X=5.27 $Y=1.61 $X2=0
+ $Y2=0
cc_417 N_A_846_74#_c_541_n N_A_634_74#_c_722_n 6.32683e-19 $X=5.21 $Y=1.775
+ $X2=0 $Y2=0
cc_418 N_A_846_74#_c_542_n N_A_634_74#_c_722_n 0.00366322f $X=5.21 $Y=1.775
+ $X2=0 $Y2=0
cc_419 N_A_846_74#_c_529_n N_A_634_74#_M1033_g 0.00312236f $X=4.37 $Y=0.515
+ $X2=0 $Y2=0
cc_420 N_A_846_74#_c_530_n N_A_634_74#_M1033_g 0.00881128f $X=5.185 $Y=0.34
+ $X2=0 $Y2=0
cc_421 N_A_846_74#_c_532_n N_A_634_74#_M1033_g 0.0254789f $X=5.27 $Y=1.61 $X2=0
+ $Y2=0
cc_422 N_A_846_74#_c_543_n N_A_634_74#_M1033_g 0.00208685f $X=5.27 $Y=0.34 $X2=0
+ $Y2=0
cc_423 N_A_846_74#_c_532_n N_A_634_74#_c_724_n 0.00859513f $X=5.27 $Y=1.61 $X2=0
+ $Y2=0
cc_424 N_A_846_74#_c_536_n N_A_634_74#_c_724_n 0.00878848f $X=6.11 $Y=1.195
+ $X2=0 $Y2=0
cc_425 N_A_846_74#_c_532_n N_A_634_74#_c_725_n 0.00152862f $X=5.27 $Y=1.61 $X2=0
+ $Y2=0
cc_426 N_A_846_74#_c_541_n N_A_634_74#_c_725_n 3.34039e-19 $X=5.21 $Y=1.775
+ $X2=0 $Y2=0
cc_427 N_A_846_74#_c_542_n N_A_634_74#_c_725_n 0.0181311f $X=5.21 $Y=1.775 $X2=0
+ $Y2=0
cc_428 N_A_846_74#_c_550_n N_A_634_74#_c_739_n 0.00165953f $X=5.21 $Y=2.13 $X2=0
+ $Y2=0
cc_429 N_A_846_74#_c_535_n N_A_634_74#_c_739_n 2.99613e-19 $X=6.11 $Y=1.195
+ $X2=0 $Y2=0
cc_430 N_A_846_74#_c_536_n N_A_634_74#_c_739_n 0.00847815f $X=6.11 $Y=1.195
+ $X2=0 $Y2=0
cc_431 N_A_846_74#_c_542_n N_A_634_74#_c_740_n 0.00418254f $X=5.21 $Y=1.775
+ $X2=0 $Y2=0
cc_432 N_A_846_74#_c_548_n N_A_634_74#_c_741_n 0.0101329f $X=5.525 $Y=2.465
+ $X2=0 $Y2=0
cc_433 N_A_846_74#_c_550_n N_A_634_74#_c_741_n 0.0148092f $X=5.21 $Y=2.13 $X2=0
+ $Y2=0
cc_434 N_A_846_74#_c_549_n N_A_634_74#_c_726_n 0.0227111f $X=8.445 $Y=2.405
+ $X2=0 $Y2=0
cc_435 N_A_846_74#_c_540_n N_A_634_74#_c_726_n 0.00240349f $X=8.37 $Y=1.99 $X2=0
+ $Y2=0
cc_436 N_A_846_74#_c_544_n N_A_634_74#_c_726_n 0.0182582f $X=8.26 $Y=1.195 $X2=0
+ $Y2=0
cc_437 N_A_846_74#_c_545_n N_A_634_74#_c_726_n 0.00194029f $X=8.37 $Y=1.195
+ $X2=0 $Y2=0
cc_438 N_A_846_74#_c_554_n N_A_634_74#_c_726_n 0.00265301f $X=8.58 $Y=2.155
+ $X2=0 $Y2=0
cc_439 N_A_846_74#_c_549_n N_A_634_74#_c_727_n 0.0221484f $X=8.445 $Y=2.405
+ $X2=0 $Y2=0
cc_440 N_A_846_74#_c_540_n N_A_634_74#_c_727_n 0.012144f $X=8.37 $Y=1.99 $X2=0
+ $Y2=0
cc_441 N_A_846_74#_c_545_n N_A_634_74#_c_727_n 2.07844e-19 $X=8.37 $Y=1.195
+ $X2=0 $Y2=0
cc_442 N_A_846_74#_c_554_n N_A_634_74#_c_727_n 0.00206412f $X=8.58 $Y=2.155
+ $X2=0 $Y2=0
cc_443 N_A_846_74#_c_540_n N_A_634_74#_M1020_g 0.00430768f $X=8.37 $Y=1.99 $X2=0
+ $Y2=0
cc_444 N_A_846_74#_c_545_n N_A_634_74#_M1020_g 0.00251517f $X=8.37 $Y=1.195
+ $X2=0 $Y2=0
cc_445 N_A_846_74#_c_547_n N_A_634_74#_M1020_g 0.0291315f $X=8.26 $Y=1.03 $X2=0
+ $Y2=0
cc_446 N_A_846_74#_c_532_n N_A_634_74#_c_729_n 0.00367699f $X=5.27 $Y=1.61 $X2=0
+ $Y2=0
cc_447 N_A_846_74#_c_529_n N_A_634_74#_c_733_n 0.00517805f $X=4.37 $Y=0.515
+ $X2=0 $Y2=0
cc_448 N_A_846_74#_c_549_n N_A_634_74#_c_747_n 5.21046e-19 $X=8.445 $Y=2.405
+ $X2=0 $Y2=0
cc_449 N_A_846_74#_c_549_n N_A_634_74#_c_749_n 0.00115715f $X=8.445 $Y=2.405
+ $X2=0 $Y2=0
cc_450 N_A_846_74#_c_540_n N_A_634_74#_c_749_n 0.0021476f $X=8.37 $Y=1.99 $X2=0
+ $Y2=0
cc_451 N_A_846_74#_c_554_n N_A_634_74#_c_749_n 0.0127458f $X=8.58 $Y=2.155 $X2=0
+ $Y2=0
cc_452 N_A_846_74#_c_540_n N_A_634_74#_c_735_n 0.0247243f $X=8.37 $Y=1.99 $X2=0
+ $Y2=0
cc_453 N_A_846_74#_c_545_n N_A_634_74#_c_735_n 0.00328136f $X=8.37 $Y=1.195
+ $X2=0 $Y2=0
cc_454 N_A_846_74#_c_537_n N_A_1287_320#_M1003_d 0.0104718f $X=8.06 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_455 N_A_846_74#_c_539_n N_A_1287_320#_M1003_d 0.00949439f $X=8.145 $Y=1.03
+ $X2=-0.19 $Y2=-0.245
cc_456 N_A_846_74#_c_533_n N_A_1287_320#_M1008_g 5.08947e-19 $X=5.945 $Y=0.34
+ $X2=0 $Y2=0
cc_457 N_A_846_74#_c_534_n N_A_1287_320#_M1008_g 0.00124396f $X=6.03 $Y=0.72
+ $X2=0 $Y2=0
cc_458 N_A_846_74#_c_535_n N_A_1287_320#_M1008_g 0.00337966f $X=6.11 $Y=1.195
+ $X2=0 $Y2=0
cc_459 N_A_846_74#_c_536_n N_A_1287_320#_M1008_g 0.00165335f $X=6.11 $Y=1.195
+ $X2=0 $Y2=0
cc_460 N_A_846_74#_c_606_p N_A_1287_320#_M1008_g 0.0145368f $X=7.22 $Y=0.805
+ $X2=0 $Y2=0
cc_461 N_A_846_74#_c_607_p N_A_1287_320#_M1008_g 0.00401876f $X=7.305 $Y=0.72
+ $X2=0 $Y2=0
cc_462 N_A_846_74#_c_546_n N_A_1287_320#_M1008_g 0.0161107f $X=6.11 $Y=1.03
+ $X2=0 $Y2=0
cc_463 N_A_846_74#_c_535_n N_A_1287_320#_c_937_n 3.74353e-19 $X=6.11 $Y=1.195
+ $X2=0 $Y2=0
cc_464 N_A_846_74#_c_536_n N_A_1287_320#_c_937_n 0.0189574f $X=6.11 $Y=1.195
+ $X2=0 $Y2=0
cc_465 N_A_846_74#_c_535_n N_A_1287_320#_c_938_n 0.0201369f $X=6.11 $Y=1.195
+ $X2=0 $Y2=0
cc_466 N_A_846_74#_c_536_n N_A_1287_320#_c_938_n 0.00103924f $X=6.11 $Y=1.195
+ $X2=0 $Y2=0
cc_467 N_A_846_74#_c_606_p N_A_1287_320#_c_938_n 0.0616788f $X=7.22 $Y=0.805
+ $X2=0 $Y2=0
cc_468 N_A_846_74#_c_606_p N_A_1287_320#_c_939_n 0.0108408f $X=7.22 $Y=0.805
+ $X2=0 $Y2=0
cc_469 N_A_846_74#_c_537_n N_A_1287_320#_c_941_n 0.020365f $X=8.06 $Y=0.34 $X2=0
+ $Y2=0
cc_470 N_A_846_74#_c_539_n N_A_1287_320#_c_941_n 0.0335581f $X=8.145 $Y=1.03
+ $X2=0 $Y2=0
cc_471 N_A_846_74#_c_545_n N_A_1287_320#_c_941_n 0.00241705f $X=8.37 $Y=1.195
+ $X2=0 $Y2=0
cc_472 N_A_846_74#_c_606_p N_A_1287_320#_c_942_n 0.00358083f $X=7.22 $Y=0.805
+ $X2=0 $Y2=0
cc_473 N_A_846_74#_c_537_n N_A_1287_320#_c_942_n 0.00370708f $X=8.06 $Y=0.34
+ $X2=0 $Y2=0
cc_474 N_A_846_74#_c_544_n N_A_1287_320#_c_942_n 8.61966e-19 $X=8.26 $Y=1.195
+ $X2=0 $Y2=0
cc_475 N_A_846_74#_c_545_n N_A_1287_320#_c_942_n 0.0198541f $X=8.37 $Y=1.195
+ $X2=0 $Y2=0
cc_476 N_A_846_74#_c_532_n N_A_1044_100#_M1033_d 0.00467191f $X=5.27 $Y=1.61
+ $X2=-0.19 $Y2=-0.245
cc_477 N_A_846_74#_c_544_n N_A_1044_100#_c_1019_n 0.00350562f $X=8.26 $Y=1.195
+ $X2=0 $Y2=0
cc_478 N_A_846_74#_c_545_n N_A_1044_100#_c_1019_n 0.00111253f $X=8.37 $Y=1.195
+ $X2=0 $Y2=0
cc_479 N_A_846_74#_c_537_n N_A_1044_100#_c_1020_n 0.0134983f $X=8.06 $Y=0.34
+ $X2=0 $Y2=0
cc_480 N_A_846_74#_c_539_n N_A_1044_100#_c_1020_n 0.00195086f $X=8.145 $Y=1.03
+ $X2=0 $Y2=0
cc_481 N_A_846_74#_c_547_n N_A_1044_100#_c_1020_n 0.00570247f $X=8.26 $Y=1.03
+ $X2=0 $Y2=0
cc_482 N_A_846_74#_c_544_n N_A_1044_100#_c_1021_n 0.00215159f $X=8.26 $Y=1.195
+ $X2=0 $Y2=0
cc_483 N_A_846_74#_c_545_n N_A_1044_100#_c_1021_n 2.47351e-19 $X=8.37 $Y=1.195
+ $X2=0 $Y2=0
cc_484 N_A_846_74#_c_532_n N_A_1044_100#_c_1022_n 0.0446664f $X=5.27 $Y=1.61
+ $X2=0 $Y2=0
cc_485 N_A_846_74#_c_536_n N_A_1044_100#_c_1022_n 0.00385914f $X=6.11 $Y=1.195
+ $X2=0 $Y2=0
cc_486 N_A_846_74#_c_541_n N_A_1044_100#_c_1022_n 0.00143774f $X=5.21 $Y=1.775
+ $X2=0 $Y2=0
cc_487 N_A_846_74#_c_535_n N_A_1044_100#_c_1023_n 0.0184576f $X=6.11 $Y=1.195
+ $X2=0 $Y2=0
cc_488 N_A_846_74#_c_536_n N_A_1044_100#_c_1023_n 0.00132041f $X=6.11 $Y=1.195
+ $X2=0 $Y2=0
cc_489 N_A_846_74#_c_532_n N_A_1044_100#_c_1024_n 0.0258589f $X=5.27 $Y=1.61
+ $X2=0 $Y2=0
cc_490 N_A_846_74#_c_533_n N_A_1044_100#_c_1024_n 0.0190961f $X=5.945 $Y=0.34
+ $X2=0 $Y2=0
cc_491 N_A_846_74#_c_534_n N_A_1044_100#_c_1024_n 0.0090117f $X=6.03 $Y=0.72
+ $X2=0 $Y2=0
cc_492 N_A_846_74#_c_535_n N_A_1044_100#_c_1024_n 0.0359115f $X=6.11 $Y=1.195
+ $X2=0 $Y2=0
cc_493 N_A_846_74#_c_639_p N_A_1044_100#_c_1024_n 0.0137306f $X=6.11 $Y=0.805
+ $X2=0 $Y2=0
cc_494 N_A_846_74#_c_546_n N_A_1044_100#_c_1024_n 0.00752036f $X=6.11 $Y=1.03
+ $X2=0 $Y2=0
cc_495 N_A_846_74#_c_541_n N_A_1044_100#_c_1029_n 0.013796f $X=5.21 $Y=1.775
+ $X2=0 $Y2=0
cc_496 N_A_846_74#_c_542_n N_A_1044_100#_c_1029_n 6.5394e-19 $X=5.21 $Y=1.775
+ $X2=0 $Y2=0
cc_497 N_A_846_74#_c_548_n N_A_1044_100#_c_1030_n 0.00682813f $X=5.525 $Y=2.465
+ $X2=0 $Y2=0
cc_498 N_A_846_74#_c_548_n N_A_1044_100#_c_1031_n 0.00102276f $X=5.525 $Y=2.465
+ $X2=0 $Y2=0
cc_499 N_A_846_74#_c_550_n N_A_1044_100#_c_1031_n 0.0139785f $X=5.21 $Y=2.13
+ $X2=0 $Y2=0
cc_500 N_A_846_74#_c_541_n N_A_1044_100#_c_1031_n 0.0361623f $X=5.21 $Y=1.775
+ $X2=0 $Y2=0
cc_501 N_A_846_74#_c_542_n N_A_1044_100#_c_1031_n 0.00117474f $X=5.21 $Y=1.775
+ $X2=0 $Y2=0
cc_502 N_A_846_74#_c_549_n N_A_1829_398#_c_1124_n 0.00805304f $X=8.445 $Y=2.405
+ $X2=0 $Y2=0
cc_503 N_A_846_74#_c_549_n N_A_1829_398#_c_1138_n 0.0124754f $X=8.445 $Y=2.405
+ $X2=0 $Y2=0
cc_504 N_A_846_74#_c_549_n N_A_1592_424#_c_1239_n 0.0173623f $X=8.445 $Y=2.405
+ $X2=0 $Y2=0
cc_505 N_A_846_74#_c_554_n N_A_1592_424#_c_1239_n 0.0279036f $X=8.58 $Y=2.155
+ $X2=0 $Y2=0
cc_506 N_A_846_74#_c_549_n N_A_1592_424#_c_1229_n 7.14051e-19 $X=8.445 $Y=2.405
+ $X2=0 $Y2=0
cc_507 N_A_846_74#_c_539_n N_A_1592_424#_c_1229_n 0.00394924f $X=8.145 $Y=1.03
+ $X2=0 $Y2=0
cc_508 N_A_846_74#_c_540_n N_A_1592_424#_c_1229_n 0.022699f $X=8.37 $Y=1.99
+ $X2=0 $Y2=0
cc_509 N_A_846_74#_c_544_n N_A_1592_424#_c_1229_n 3.46053e-19 $X=8.26 $Y=1.195
+ $X2=0 $Y2=0
cc_510 N_A_846_74#_c_545_n N_A_1592_424#_c_1229_n 0.0125435f $X=8.37 $Y=1.195
+ $X2=0 $Y2=0
cc_511 N_A_846_74#_c_554_n N_A_1592_424#_c_1229_n 0.00644238f $X=8.58 $Y=2.155
+ $X2=0 $Y2=0
cc_512 N_A_846_74#_c_547_n N_A_1592_424#_c_1229_n 7.20283e-19 $X=8.26 $Y=1.03
+ $X2=0 $Y2=0
cc_513 N_A_846_74#_c_549_n N_A_1592_424#_c_1234_n 0.00382531f $X=8.445 $Y=2.405
+ $X2=0 $Y2=0
cc_514 N_A_846_74#_c_554_n N_A_1592_424#_c_1234_n 0.00567093f $X=8.58 $Y=2.155
+ $X2=0 $Y2=0
cc_515 N_A_846_74#_c_549_n N_A_1592_424#_c_1237_n 0.00711213f $X=8.445 $Y=2.405
+ $X2=0 $Y2=0
cc_516 N_A_846_74#_c_537_n N_A_1592_424#_c_1231_n 0.00381206f $X=8.06 $Y=0.34
+ $X2=0 $Y2=0
cc_517 N_A_846_74#_c_545_n N_A_1592_424#_c_1231_n 0.00261887f $X=8.37 $Y=1.195
+ $X2=0 $Y2=0
cc_518 N_A_846_74#_c_547_n N_A_1592_424#_c_1231_n 0.00657447f $X=8.26 $Y=1.03
+ $X2=0 $Y2=0
cc_519 N_A_846_74#_c_549_n N_A_1592_424#_c_1238_n 0.00155529f $X=8.445 $Y=2.405
+ $X2=0 $Y2=0
cc_520 N_A_846_74#_c_554_n N_A_1592_424#_c_1238_n 0.0146828f $X=8.58 $Y=2.155
+ $X2=0 $Y2=0
cc_521 N_A_846_74#_c_548_n N_VPWR_c_1325_n 0.00411612f $X=5.525 $Y=2.465 $X2=0
+ $Y2=0
cc_522 N_A_846_74#_c_549_n N_VPWR_c_1329_n 0.0041293f $X=8.445 $Y=2.405 $X2=0
+ $Y2=0
cc_523 N_A_846_74#_c_548_n N_VPWR_c_1315_n 0.00753176f $X=5.525 $Y=2.465 $X2=0
+ $Y2=0
cc_524 N_A_846_74#_c_549_n N_VPWR_c_1315_n 0.00526787f $X=8.445 $Y=2.405 $X2=0
+ $Y2=0
cc_525 N_A_846_74#_c_550_n N_VPWR_c_1315_n 3.36114e-19 $X=5.21 $Y=2.13 $X2=0
+ $Y2=0
cc_526 N_A_846_74#_c_541_n N_A_300_453#_c_1457_n 0.0421436f $X=5.21 $Y=1.775
+ $X2=0 $Y2=0
cc_527 N_A_846_74#_c_542_n N_A_300_453#_c_1457_n 5.20094e-19 $X=5.21 $Y=1.775
+ $X2=0 $Y2=0
cc_528 N_A_846_74#_c_529_n N_A_300_453#_c_1458_n 0.003919f $X=4.37 $Y=0.515
+ $X2=0 $Y2=0
cc_529 N_A_846_74#_c_532_n N_A_300_453#_c_1458_n 0.00870834f $X=5.27 $Y=1.61
+ $X2=0 $Y2=0
cc_530 N_A_846_74#_c_541_n N_A_300_453#_c_1458_n 0.0116273f $X=5.21 $Y=1.775
+ $X2=0 $Y2=0
cc_531 N_A_846_74#_c_529_n N_A_300_453#_c_1514_n 0.0151548f $X=4.37 $Y=0.515
+ $X2=0 $Y2=0
cc_532 N_A_846_74#_M1027_d N_A_300_453#_c_1464_n 0.00830482f $X=4.59 $Y=1.84
+ $X2=0 $Y2=0
cc_533 N_A_846_74#_c_548_n N_A_300_453#_c_1464_n 0.00227377f $X=5.525 $Y=2.465
+ $X2=0 $Y2=0
cc_534 N_A_846_74#_c_550_n N_A_300_453#_c_1464_n 0.00321103f $X=5.21 $Y=2.13
+ $X2=0 $Y2=0
cc_535 N_A_846_74#_c_541_n N_A_300_453#_c_1464_n 0.0593436f $X=5.21 $Y=1.775
+ $X2=0 $Y2=0
cc_536 N_A_846_74#_c_529_n N_A_300_453#_c_1459_n 0.015064f $X=4.37 $Y=0.515
+ $X2=0 $Y2=0
cc_537 N_A_846_74#_c_532_n N_A_300_453#_c_1459_n 0.0161196f $X=5.27 $Y=1.61
+ $X2=0 $Y2=0
cc_538 N_A_846_74#_c_548_n N_A_300_453#_c_1465_n 0.00173049f $X=5.525 $Y=2.465
+ $X2=0 $Y2=0
cc_539 N_A_846_74#_c_529_n N_A_300_453#_c_1460_n 0.0285593f $X=4.37 $Y=0.515
+ $X2=0 $Y2=0
cc_540 N_A_846_74#_c_530_n N_A_300_453#_c_1460_n 0.0227483f $X=5.185 $Y=0.34
+ $X2=0 $Y2=0
cc_541 N_A_846_74#_c_532_n N_A_300_453#_c_1460_n 0.0124252f $X=5.27 $Y=1.61
+ $X2=0 $Y2=0
cc_542 N_A_846_74#_c_606_p N_VGND_M1008_d 0.0173766f $X=7.22 $Y=0.805 $X2=0
+ $Y2=0
cc_543 N_A_846_74#_c_607_p N_VGND_M1008_d 0.0052578f $X=7.305 $Y=0.72 $X2=0
+ $Y2=0
cc_544 N_A_846_74#_c_538_n N_VGND_M1008_d 6.57704e-19 $X=7.39 $Y=0.34 $X2=0
+ $Y2=0
cc_545 N_A_846_74#_c_531_n N_VGND_c_1615_n 0.011924f $X=4.535 $Y=0.34 $X2=0
+ $Y2=0
cc_546 N_A_846_74#_c_533_n N_VGND_c_1616_n 0.00618185f $X=5.945 $Y=0.34 $X2=0
+ $Y2=0
cc_547 N_A_846_74#_c_534_n N_VGND_c_1616_n 0.00238541f $X=6.03 $Y=0.72 $X2=0
+ $Y2=0
cc_548 N_A_846_74#_c_606_p N_VGND_c_1616_n 0.0255462f $X=7.22 $Y=0.805 $X2=0
+ $Y2=0
cc_549 N_A_846_74#_c_607_p N_VGND_c_1616_n 0.0095164f $X=7.305 $Y=0.72 $X2=0
+ $Y2=0
cc_550 N_A_846_74#_c_538_n N_VGND_c_1616_n 0.0148568f $X=7.39 $Y=0.34 $X2=0
+ $Y2=0
cc_551 N_A_846_74#_c_530_n N_VGND_c_1625_n 0.0418136f $X=5.185 $Y=0.34 $X2=0
+ $Y2=0
cc_552 N_A_846_74#_c_531_n N_VGND_c_1625_n 0.0235688f $X=4.535 $Y=0.34 $X2=0
+ $Y2=0
cc_553 N_A_846_74#_c_533_n N_VGND_c_1625_n 0.0501353f $X=5.945 $Y=0.34 $X2=0
+ $Y2=0
cc_554 N_A_846_74#_c_606_p N_VGND_c_1625_n 0.00556178f $X=7.22 $Y=0.805 $X2=0
+ $Y2=0
cc_555 N_A_846_74#_c_543_n N_VGND_c_1625_n 0.0121867f $X=5.27 $Y=0.34 $X2=0
+ $Y2=0
cc_556 N_A_846_74#_c_639_p N_VGND_c_1625_n 0.00227233f $X=6.11 $Y=0.805 $X2=0
+ $Y2=0
cc_557 N_A_846_74#_c_546_n N_VGND_c_1625_n 7.07447e-19 $X=6.11 $Y=1.03 $X2=0
+ $Y2=0
cc_558 N_A_846_74#_c_606_p N_VGND_c_1626_n 0.00246644f $X=7.22 $Y=0.805 $X2=0
+ $Y2=0
cc_559 N_A_846_74#_c_537_n N_VGND_c_1626_n 0.0548521f $X=8.06 $Y=0.34 $X2=0
+ $Y2=0
cc_560 N_A_846_74#_c_538_n N_VGND_c_1626_n 0.0121237f $X=7.39 $Y=0.34 $X2=0
+ $Y2=0
cc_561 N_A_846_74#_c_547_n N_VGND_c_1626_n 0.00433139f $X=8.26 $Y=1.03 $X2=0
+ $Y2=0
cc_562 N_A_846_74#_c_530_n N_VGND_c_1633_n 0.0244305f $X=5.185 $Y=0.34 $X2=0
+ $Y2=0
cc_563 N_A_846_74#_c_531_n N_VGND_c_1633_n 0.0127152f $X=4.535 $Y=0.34 $X2=0
+ $Y2=0
cc_564 N_A_846_74#_c_533_n N_VGND_c_1633_n 0.0287839f $X=5.945 $Y=0.34 $X2=0
+ $Y2=0
cc_565 N_A_846_74#_c_606_p N_VGND_c_1633_n 0.0176164f $X=7.22 $Y=0.805 $X2=0
+ $Y2=0
cc_566 N_A_846_74#_c_537_n N_VGND_c_1633_n 0.0311091f $X=8.06 $Y=0.34 $X2=0
+ $Y2=0
cc_567 N_A_846_74#_c_538_n N_VGND_c_1633_n 0.00659733f $X=7.39 $Y=0.34 $X2=0
+ $Y2=0
cc_568 N_A_846_74#_c_543_n N_VGND_c_1633_n 0.00660921f $X=5.27 $Y=0.34 $X2=0
+ $Y2=0
cc_569 N_A_846_74#_c_639_p N_VGND_c_1633_n 0.00453863f $X=6.11 $Y=0.805 $X2=0
+ $Y2=0
cc_570 N_A_846_74#_c_547_n N_VGND_c_1633_n 0.00821191f $X=8.26 $Y=1.03 $X2=0
+ $Y2=0
cc_571 N_A_846_74#_c_535_n A_1219_100# 3.83906e-19 $X=6.11 $Y=1.195 $X2=-0.19
+ $Y2=-0.245
cc_572 N_A_846_74#_c_606_p A_1219_100# 0.0108377f $X=7.22 $Y=0.805 $X2=-0.19
+ $Y2=-0.245
cc_573 N_A_846_74#_c_639_p A_1219_100# 0.0024378f $X=6.11 $Y=0.805 $X2=-0.19
+ $Y2=-0.245
cc_574 N_A_634_74#_c_747_n N_A_1287_320#_M1007_d 0.00963911f $X=7.685 $Y=2.99
+ $X2=0 $Y2=0
cc_575 N_A_634_74#_c_749_n N_A_1287_320#_M1007_d 0.00850114f $X=7.77 $Y=2.905
+ $X2=0 $Y2=0
cc_576 N_A_634_74#_c_740_n N_A_1287_320#_c_943_n 0.0186227f $X=6.055 $Y=2.13
+ $X2=0 $Y2=0
cc_577 N_A_634_74#_c_741_n N_A_1287_320#_c_943_n 0.00667645f $X=5.975 $Y=2.465
+ $X2=0 $Y2=0
cc_578 N_A_634_74#_c_746_n N_A_1287_320#_c_943_n 0.017876f $X=7.005 $Y=2.215
+ $X2=0 $Y2=0
cc_579 N_A_634_74#_c_820_p N_A_1287_320#_c_943_n 0.00290101f $X=7.09 $Y=2.905
+ $X2=0 $Y2=0
cc_580 N_A_634_74#_c_750_n N_A_1287_320#_c_943_n 0.00119336f $X=6.06 $Y=2.135
+ $X2=0 $Y2=0
cc_581 N_A_634_74#_c_741_n N_A_1287_320#_c_944_n 0.0177572f $X=5.975 $Y=2.465
+ $X2=0 $Y2=0
cc_582 N_A_634_74#_c_820_p N_A_1287_320#_c_944_n 0.00151708f $X=7.09 $Y=2.905
+ $X2=0 $Y2=0
cc_583 N_A_634_74#_c_748_n N_A_1287_320#_c_944_n 4.36296e-19 $X=7.175 $Y=2.99
+ $X2=0 $Y2=0
cc_584 N_A_634_74#_c_725_n N_A_1287_320#_c_936_n 0.00140785f $X=5.66 $Y=1.74
+ $X2=0 $Y2=0
cc_585 N_A_634_74#_c_739_n N_A_1287_320#_c_936_n 0.0186227f $X=6.055 $Y=1.89
+ $X2=0 $Y2=0
cc_586 N_A_634_74#_c_726_n N_A_1287_320#_c_940_n 0.00218584f $X=7.885 $Y=2.045
+ $X2=0 $Y2=0
cc_587 N_A_634_74#_c_746_n N_A_1287_320#_c_940_n 0.0133617f $X=7.005 $Y=2.215
+ $X2=0 $Y2=0
cc_588 N_A_634_74#_c_820_p N_A_1287_320#_c_940_n 0.0217294f $X=7.09 $Y=2.905
+ $X2=0 $Y2=0
cc_589 N_A_634_74#_c_747_n N_A_1287_320#_c_940_n 0.00795931f $X=7.685 $Y=2.99
+ $X2=0 $Y2=0
cc_590 N_A_634_74#_c_749_n N_A_1287_320#_c_940_n 0.0497825f $X=7.77 $Y=2.905
+ $X2=0 $Y2=0
cc_591 N_A_634_74#_c_735_n N_A_1287_320#_c_940_n 0.0254106f $X=7.95 $Y=1.765
+ $X2=0 $Y2=0
cc_592 N_A_634_74#_c_726_n N_A_1287_320#_c_942_n 0.00242456f $X=7.885 $Y=2.045
+ $X2=0 $Y2=0
cc_593 N_A_634_74#_c_735_n N_A_1287_320#_c_942_n 0.0100661f $X=7.95 $Y=1.765
+ $X2=0 $Y2=0
cc_594 N_A_634_74#_c_726_n N_A_1044_100#_c_1027_n 0.0142873f $X=7.885 $Y=2.045
+ $X2=0 $Y2=0
cc_595 N_A_634_74#_c_746_n N_A_1044_100#_c_1027_n 0.00569916f $X=7.005 $Y=2.215
+ $X2=0 $Y2=0
cc_596 N_A_634_74#_c_820_p N_A_1044_100#_c_1027_n 0.0162181f $X=7.09 $Y=2.905
+ $X2=0 $Y2=0
cc_597 N_A_634_74#_c_747_n N_A_1044_100#_c_1027_n 0.00981164f $X=7.685 $Y=2.99
+ $X2=0 $Y2=0
cc_598 N_A_634_74#_c_748_n N_A_1044_100#_c_1027_n 0.00287436f $X=7.175 $Y=2.99
+ $X2=0 $Y2=0
cc_599 N_A_634_74#_c_749_n N_A_1044_100#_c_1027_n 0.00302367f $X=7.77 $Y=2.905
+ $X2=0 $Y2=0
cc_600 N_A_634_74#_c_726_n N_A_1044_100#_c_1019_n 0.0181601f $X=7.885 $Y=2.045
+ $X2=0 $Y2=0
cc_601 N_A_634_74#_c_735_n N_A_1044_100#_c_1019_n 0.00234362f $X=7.95 $Y=1.765
+ $X2=0 $Y2=0
cc_602 N_A_634_74#_M1033_g N_A_1044_100#_c_1022_n 0.00144305f $X=5.145 $Y=0.71
+ $X2=0 $Y2=0
cc_603 N_A_634_74#_c_724_n N_A_1044_100#_c_1022_n 0.00943459f $X=5.585 $Y=1.295
+ $X2=0 $Y2=0
cc_604 N_A_634_74#_c_725_n N_A_1044_100#_c_1022_n 0.0108414f $X=5.66 $Y=1.74
+ $X2=0 $Y2=0
cc_605 N_A_634_74#_c_739_n N_A_1044_100#_c_1023_n 0.0171749f $X=6.055 $Y=1.89
+ $X2=0 $Y2=0
cc_606 N_A_634_74#_c_746_n N_A_1044_100#_c_1023_n 0.0281079f $X=7.005 $Y=2.215
+ $X2=0 $Y2=0
cc_607 N_A_634_74#_c_750_n N_A_1044_100#_c_1023_n 0.023546f $X=6.06 $Y=2.135
+ $X2=0 $Y2=0
cc_608 N_A_634_74#_M1033_g N_A_1044_100#_c_1024_n 0.00181773f $X=5.145 $Y=0.71
+ $X2=0 $Y2=0
cc_609 N_A_634_74#_c_724_n N_A_1044_100#_c_1024_n 0.00115095f $X=5.585 $Y=1.295
+ $X2=0 $Y2=0
cc_610 N_A_634_74#_c_725_n N_A_1044_100#_c_1029_n 0.00402552f $X=5.66 $Y=1.74
+ $X2=0 $Y2=0
cc_611 N_A_634_74#_c_739_n N_A_1044_100#_c_1029_n 0.004382f $X=6.055 $Y=1.89
+ $X2=0 $Y2=0
cc_612 N_A_634_74#_c_739_n N_A_1044_100#_c_1030_n 0.00389495f $X=6.055 $Y=1.89
+ $X2=0 $Y2=0
cc_613 N_A_634_74#_c_741_n N_A_1044_100#_c_1030_n 0.0109441f $X=5.975 $Y=2.465
+ $X2=0 $Y2=0
cc_614 N_A_634_74#_c_750_n N_A_1044_100#_c_1030_n 0.0011545f $X=6.06 $Y=2.135
+ $X2=0 $Y2=0
cc_615 N_A_634_74#_c_739_n N_A_1044_100#_c_1031_n 0.00811793f $X=6.055 $Y=1.89
+ $X2=0 $Y2=0
cc_616 N_A_634_74#_c_740_n N_A_1044_100#_c_1031_n 0.00790739f $X=6.055 $Y=2.13
+ $X2=0 $Y2=0
cc_617 N_A_634_74#_c_741_n N_A_1044_100#_c_1031_n 0.00112121f $X=5.975 $Y=2.465
+ $X2=0 $Y2=0
cc_618 N_A_634_74#_c_750_n N_A_1044_100#_c_1031_n 0.0247638f $X=6.06 $Y=2.135
+ $X2=0 $Y2=0
cc_619 N_A_634_74#_c_746_n N_A_1044_100#_c_1025_n 0.0231235f $X=7.005 $Y=2.215
+ $X2=0 $Y2=0
cc_620 N_A_634_74#_c_726_n N_A_1044_100#_c_1026_n 0.00301676f $X=7.885 $Y=2.045
+ $X2=0 $Y2=0
cc_621 N_A_634_74#_c_746_n N_A_1044_100#_c_1026_n 0.00186203f $X=7.005 $Y=2.215
+ $X2=0 $Y2=0
cc_622 N_A_634_74#_c_749_n N_A_1044_100#_c_1026_n 2.06351e-19 $X=7.77 $Y=2.905
+ $X2=0 $Y2=0
cc_623 N_A_634_74#_c_727_n N_A_1829_398#_c_1124_n 0.0376175f $X=8.785 $Y=1.675
+ $X2=0 $Y2=0
cc_624 N_A_634_74#_M1020_g N_A_1829_398#_M1021_g 0.0376175f $X=8.86 $Y=0.58
+ $X2=0 $Y2=0
cc_625 N_A_634_74#_M1020_g N_A_1829_398#_c_1130_n 4.71258e-19 $X=8.86 $Y=0.58
+ $X2=0 $Y2=0
cc_626 N_A_634_74#_c_727_n N_A_1592_424#_c_1229_n 0.00603578f $X=8.785 $Y=1.675
+ $X2=0 $Y2=0
cc_627 N_A_634_74#_M1020_g N_A_1592_424#_c_1229_n 0.0194763f $X=8.86 $Y=0.58
+ $X2=0 $Y2=0
cc_628 N_A_634_74#_c_726_n N_A_1592_424#_c_1237_n 0.0030559f $X=7.885 $Y=2.045
+ $X2=0 $Y2=0
cc_629 N_A_634_74#_c_747_n N_A_1592_424#_c_1237_n 0.0012115f $X=7.685 $Y=2.99
+ $X2=0 $Y2=0
cc_630 N_A_634_74#_c_749_n N_A_1592_424#_c_1237_n 0.0299969f $X=7.77 $Y=2.905
+ $X2=0 $Y2=0
cc_631 N_A_634_74#_c_735_n N_A_1592_424#_c_1237_n 0.00278637f $X=7.95 $Y=1.765
+ $X2=0 $Y2=0
cc_632 N_A_634_74#_M1020_g N_A_1592_424#_c_1231_n 0.0223895f $X=8.86 $Y=0.58
+ $X2=0 $Y2=0
cc_633 N_A_634_74#_c_744_n N_VPWR_M1027_s 0.00960989f $X=3.855 $Y=2.115 $X2=0
+ $Y2=0
cc_634 N_A_634_74#_c_734_n N_VPWR_M1027_s 0.00232415f $X=4 $Y=1.465 $X2=0 $Y2=0
cc_635 N_A_634_74#_c_746_n N_VPWR_M1005_d 0.00780352f $X=7.005 $Y=2.215 $X2=0
+ $Y2=0
cc_636 N_A_634_74#_c_820_p N_VPWR_M1005_d 0.00658543f $X=7.09 $Y=2.905 $X2=0
+ $Y2=0
cc_637 N_A_634_74#_c_748_n N_VPWR_M1005_d 5.2468e-19 $X=7.175 $Y=2.99 $X2=0
+ $Y2=0
cc_638 N_A_634_74#_c_741_n N_VPWR_c_1318_n 0.0019285f $X=5.975 $Y=2.465 $X2=0
+ $Y2=0
cc_639 N_A_634_74#_c_746_n N_VPWR_c_1318_n 0.0172937f $X=7.005 $Y=2.215 $X2=0
+ $Y2=0
cc_640 N_A_634_74#_c_820_p N_VPWR_c_1318_n 0.0287875f $X=7.09 $Y=2.905 $X2=0
+ $Y2=0
cc_641 N_A_634_74#_c_748_n N_VPWR_c_1318_n 0.0145682f $X=7.175 $Y=2.99 $X2=0
+ $Y2=0
cc_642 N_A_634_74#_c_736_n N_VPWR_c_1325_n 0.00334029f $X=4.515 $Y=1.765 $X2=0
+ $Y2=0
cc_643 N_A_634_74#_c_741_n N_VPWR_c_1325_n 0.00445602f $X=5.975 $Y=2.465 $X2=0
+ $Y2=0
cc_644 N_A_634_74#_c_726_n N_VPWR_c_1329_n 0.00406462f $X=7.885 $Y=2.045 $X2=0
+ $Y2=0
cc_645 N_A_634_74#_c_747_n N_VPWR_c_1329_n 0.0444882f $X=7.685 $Y=2.99 $X2=0
+ $Y2=0
cc_646 N_A_634_74#_c_748_n N_VPWR_c_1329_n 0.0120286f $X=7.175 $Y=2.99 $X2=0
+ $Y2=0
cc_647 N_A_634_74#_c_736_n N_VPWR_c_1333_n 0.0129364f $X=4.515 $Y=1.765 $X2=0
+ $Y2=0
cc_648 N_A_634_74#_c_736_n N_VPWR_c_1315_n 0.00441383f $X=4.515 $Y=1.765 $X2=0
+ $Y2=0
cc_649 N_A_634_74#_c_741_n N_VPWR_c_1315_n 0.0089717f $X=5.975 $Y=2.465 $X2=0
+ $Y2=0
cc_650 N_A_634_74#_c_726_n N_VPWR_c_1315_n 0.00749521f $X=7.885 $Y=2.045 $X2=0
+ $Y2=0
cc_651 N_A_634_74#_c_747_n N_VPWR_c_1315_n 0.0250882f $X=7.685 $Y=2.99 $X2=0
+ $Y2=0
cc_652 N_A_634_74#_c_748_n N_VPWR_c_1315_n 0.0064033f $X=7.175 $Y=2.99 $X2=0
+ $Y2=0
cc_653 N_A_634_74#_c_730_n N_A_300_453#_c_1453_n 0.00277283f $X=3.31 $Y=0.755
+ $X2=0 $Y2=0
cc_654 N_A_634_74#_c_730_n N_A_300_453#_c_1454_n 0.00711146f $X=3.31 $Y=0.755
+ $X2=0 $Y2=0
cc_655 N_A_634_74#_c_744_n N_A_300_453#_c_1456_n 0.0211068f $X=3.855 $Y=2.115
+ $X2=0 $Y2=0
cc_656 N_A_634_74#_M1004_d N_A_300_453#_c_1462_n 0.00810075f $X=3.355 $Y=1.84
+ $X2=0 $Y2=0
cc_657 N_A_634_74#_c_744_n N_A_300_453#_c_1462_n 0.059138f $X=3.855 $Y=2.115
+ $X2=0 $Y2=0
cc_658 N_A_634_74#_c_736_n N_A_300_453#_c_1457_n 0.0250759f $X=4.515 $Y=1.765
+ $X2=0 $Y2=0
cc_659 N_A_634_74#_c_722_n N_A_300_453#_c_1457_n 0.0184134f $X=4.605 $Y=1.295
+ $X2=0 $Y2=0
cc_660 N_A_634_74#_c_744_n N_A_300_453#_c_1457_n 0.0268482f $X=3.855 $Y=2.115
+ $X2=0 $Y2=0
cc_661 N_A_634_74#_c_734_n N_A_300_453#_c_1457_n 0.0360363f $X=4 $Y=1.465 $X2=0
+ $Y2=0
cc_662 N_A_634_74#_c_721_n N_A_300_453#_c_1458_n 0.00973978f $X=5.07 $Y=1.295
+ $X2=0 $Y2=0
cc_663 N_A_634_74#_c_722_n N_A_300_453#_c_1458_n 0.0120397f $X=4.605 $Y=1.295
+ $X2=0 $Y2=0
cc_664 N_A_634_74#_c_722_n N_A_300_453#_c_1514_n 0.00637908f $X=4.605 $Y=1.295
+ $X2=0 $Y2=0
cc_665 N_A_634_74#_c_733_n N_A_300_453#_c_1514_n 0.0113493f $X=4 $Y=1.445 $X2=0
+ $Y2=0
cc_666 N_A_634_74#_c_734_n N_A_300_453#_c_1514_n 0.00190953f $X=4 $Y=1.465 $X2=0
+ $Y2=0
cc_667 N_A_634_74#_c_736_n N_A_300_453#_c_1464_n 0.0127753f $X=4.515 $Y=1.765
+ $X2=0 $Y2=0
cc_668 N_A_634_74#_c_720_n N_A_300_453#_c_1459_n 0.00250911f $X=4.155 $Y=1.22
+ $X2=0 $Y2=0
cc_669 N_A_634_74#_c_721_n N_A_300_453#_c_1459_n 0.0095699f $X=5.07 $Y=1.295
+ $X2=0 $Y2=0
cc_670 N_A_634_74#_M1033_g N_A_300_453#_c_1459_n 0.00559554f $X=5.145 $Y=0.71
+ $X2=0 $Y2=0
cc_671 N_A_634_74#_c_736_n N_A_300_453#_c_1465_n 0.00871208f $X=4.515 $Y=1.765
+ $X2=0 $Y2=0
cc_672 N_A_634_74#_c_736_n N_A_300_453#_c_1544_n 0.0058649f $X=4.515 $Y=1.765
+ $X2=0 $Y2=0
cc_673 N_A_634_74#_c_720_n N_A_300_453#_c_1460_n 6.35404e-19 $X=4.155 $Y=1.22
+ $X2=0 $Y2=0
cc_674 N_A_634_74#_c_721_n N_A_300_453#_c_1460_n 0.00412678f $X=5.07 $Y=1.295
+ $X2=0 $Y2=0
cc_675 N_A_634_74#_M1033_g N_A_300_453#_c_1460_n 4.21674e-19 $X=5.145 $Y=0.71
+ $X2=0 $Y2=0
cc_676 N_A_634_74#_c_732_n N_VGND_M1028_s 0.00157836f $X=3.855 $Y=1.095 $X2=0
+ $Y2=0
cc_677 N_A_634_74#_c_733_n N_VGND_M1028_s 0.00213809f $X=4 $Y=1.445 $X2=0 $Y2=0
cc_678 N_A_634_74#_c_731_n N_VGND_c_1614_n 0.0174746f $X=3.31 $Y=0.495 $X2=0
+ $Y2=0
cc_679 N_A_634_74#_c_720_n N_VGND_c_1615_n 0.0123061f $X=4.155 $Y=1.22 $X2=0
+ $Y2=0
cc_680 N_A_634_74#_c_722_n N_VGND_c_1615_n 8.25268e-19 $X=4.605 $Y=1.295 $X2=0
+ $Y2=0
cc_681 N_A_634_74#_c_730_n N_VGND_c_1615_n 0.00575054f $X=3.31 $Y=0.755 $X2=0
+ $Y2=0
cc_682 N_A_634_74#_c_731_n N_VGND_c_1615_n 0.0286194f $X=3.31 $Y=0.495 $X2=0
+ $Y2=0
cc_683 N_A_634_74#_c_732_n N_VGND_c_1615_n 0.0121449f $X=3.855 $Y=1.095 $X2=0
+ $Y2=0
cc_684 N_A_634_74#_c_733_n N_VGND_c_1615_n 0.0151471f $X=4 $Y=1.445 $X2=0 $Y2=0
cc_685 N_A_634_74#_M1020_g N_VGND_c_1617_n 0.00153607f $X=8.86 $Y=0.58 $X2=0
+ $Y2=0
cc_686 N_A_634_74#_c_731_n N_VGND_c_1623_n 0.0157574f $X=3.31 $Y=0.495 $X2=0
+ $Y2=0
cc_687 N_A_634_74#_c_720_n N_VGND_c_1625_n 0.00430908f $X=4.155 $Y=1.22 $X2=0
+ $Y2=0
cc_688 N_A_634_74#_M1033_g N_VGND_c_1625_n 7.26171e-19 $X=5.145 $Y=0.71 $X2=0
+ $Y2=0
cc_689 N_A_634_74#_M1020_g N_VGND_c_1626_n 0.0032429f $X=8.86 $Y=0.58 $X2=0
+ $Y2=0
cc_690 N_A_634_74#_c_720_n N_VGND_c_1633_n 0.00825456f $X=4.155 $Y=1.22 $X2=0
+ $Y2=0
cc_691 N_A_634_74#_M1020_g N_VGND_c_1633_n 0.00411459f $X=8.86 $Y=0.58 $X2=0
+ $Y2=0
cc_692 N_A_634_74#_c_731_n N_VGND_c_1633_n 0.012116f $X=3.31 $Y=0.495 $X2=0
+ $Y2=0
cc_693 N_A_1287_320#_c_943_n N_A_1044_100#_c_1027_n 0.00852317f $X=6.525
+ $Y=2.375 $X2=0 $Y2=0
cc_694 N_A_1287_320#_c_944_n N_A_1044_100#_c_1027_n 0.00739406f $X=6.525
+ $Y=2.465 $X2=0 $Y2=0
cc_695 N_A_1287_320#_c_940_n N_A_1044_100#_c_1027_n 0.0041807f $X=7.43 $Y=2.41
+ $X2=0 $Y2=0
cc_696 N_A_1287_320#_c_940_n N_A_1044_100#_c_1019_n 0.0141225f $X=7.43 $Y=2.41
+ $X2=0 $Y2=0
cc_697 N_A_1287_320#_c_942_n N_A_1044_100#_c_1019_n 0.0112775f $X=7.345 $Y=1.06
+ $X2=0 $Y2=0
cc_698 N_A_1287_320#_c_941_n N_A_1044_100#_c_1020_n 0.00921118f $X=7.725
+ $Y=0.765 $X2=0 $Y2=0
cc_699 N_A_1287_320#_c_939_n N_A_1044_100#_c_1021_n 0.0181405f $X=6.99 $Y=1.225
+ $X2=0 $Y2=0
cc_700 N_A_1287_320#_c_941_n N_A_1044_100#_c_1021_n 0.0038152f $X=7.725 $Y=0.765
+ $X2=0 $Y2=0
cc_701 N_A_1287_320#_c_942_n N_A_1044_100#_c_1021_n 0.0086565f $X=7.345 $Y=1.06
+ $X2=0 $Y2=0
cc_702 N_A_1287_320#_c_936_n N_A_1044_100#_c_1022_n 4.23402e-19 $X=6.535 $Y=1.75
+ $X2=0 $Y2=0
cc_703 N_A_1287_320#_c_943_n N_A_1044_100#_c_1023_n 0.0052513f $X=6.525 $Y=2.375
+ $X2=0 $Y2=0
cc_704 N_A_1287_320#_c_936_n N_A_1044_100#_c_1023_n 0.0102739f $X=6.535 $Y=1.75
+ $X2=0 $Y2=0
cc_705 N_A_1287_320#_c_937_n N_A_1044_100#_c_1023_n 0.00458197f $X=6.575
+ $Y=1.225 $X2=0 $Y2=0
cc_706 N_A_1287_320#_c_938_n N_A_1044_100#_c_1023_n 0.0202979f $X=7.345 $Y=1.225
+ $X2=0 $Y2=0
cc_707 N_A_1287_320#_c_944_n N_A_1044_100#_c_1030_n 0.00141636f $X=6.525
+ $Y=2.465 $X2=0 $Y2=0
cc_708 N_A_1287_320#_c_943_n N_A_1044_100#_c_1025_n 0.00110089f $X=6.525
+ $Y=2.375 $X2=0 $Y2=0
cc_709 N_A_1287_320#_c_938_n N_A_1044_100#_c_1025_n 0.0188377f $X=7.345 $Y=1.225
+ $X2=0 $Y2=0
cc_710 N_A_1287_320#_c_939_n N_A_1044_100#_c_1025_n 0.00113929f $X=6.99 $Y=1.225
+ $X2=0 $Y2=0
cc_711 N_A_1287_320#_c_940_n N_A_1044_100#_c_1025_n 0.0235661f $X=7.43 $Y=2.41
+ $X2=0 $Y2=0
cc_712 N_A_1287_320#_c_943_n N_A_1044_100#_c_1026_n 0.015606f $X=6.525 $Y=2.375
+ $X2=0 $Y2=0
cc_713 N_A_1287_320#_c_936_n N_A_1044_100#_c_1026_n 0.00780769f $X=6.535 $Y=1.75
+ $X2=0 $Y2=0
cc_714 N_A_1287_320#_c_938_n N_A_1044_100#_c_1026_n 0.00732192f $X=7.345
+ $Y=1.225 $X2=0 $Y2=0
cc_715 N_A_1287_320#_c_939_n N_A_1044_100#_c_1026_n 0.016565f $X=6.99 $Y=1.225
+ $X2=0 $Y2=0
cc_716 N_A_1287_320#_c_940_n N_A_1044_100#_c_1026_n 0.0188151f $X=7.43 $Y=2.41
+ $X2=0 $Y2=0
cc_717 N_A_1287_320#_c_944_n N_VPWR_c_1318_n 0.0145822f $X=6.525 $Y=2.465 $X2=0
+ $Y2=0
cc_718 N_A_1287_320#_c_944_n N_VPWR_c_1325_n 0.00413917f $X=6.525 $Y=2.465 $X2=0
+ $Y2=0
cc_719 N_A_1287_320#_c_944_n N_VPWR_c_1315_n 0.00856462f $X=6.525 $Y=2.465 $X2=0
+ $Y2=0
cc_720 N_A_1287_320#_M1008_g N_VGND_c_1616_n 0.00467601f $X=6.59 $Y=0.71 $X2=0
+ $Y2=0
cc_721 N_A_1287_320#_M1008_g N_VGND_c_1625_n 0.00381137f $X=6.59 $Y=0.71 $X2=0
+ $Y2=0
cc_722 N_A_1287_320#_M1008_g N_VGND_c_1633_n 0.00505379f $X=6.59 $Y=0.71 $X2=0
+ $Y2=0
cc_723 N_A_1044_100#_c_1027_n N_VPWR_c_1318_n 0.00193557f $X=7.205 $Y=2.045
+ $X2=0 $Y2=0
cc_724 N_A_1044_100#_c_1030_n N_VPWR_c_1318_n 0.010809f $X=5.75 $Y=2.75 $X2=0
+ $Y2=0
cc_725 N_A_1044_100#_c_1030_n N_VPWR_c_1325_n 0.015569f $X=5.75 $Y=2.75 $X2=0
+ $Y2=0
cc_726 N_A_1044_100#_c_1027_n N_VPWR_c_1329_n 0.00278227f $X=7.205 $Y=2.045
+ $X2=0 $Y2=0
cc_727 N_A_1044_100#_c_1027_n N_VPWR_c_1315_n 0.00357373f $X=7.205 $Y=2.045
+ $X2=0 $Y2=0
cc_728 N_A_1044_100#_c_1030_n N_VPWR_c_1315_n 0.0128526f $X=5.75 $Y=2.75 $X2=0
+ $Y2=0
cc_729 N_A_1044_100#_c_1031_n N_A_300_453#_c_1464_n 0.0139222f $X=5.735 $Y=2.52
+ $X2=0 $Y2=0
cc_730 N_A_1044_100#_c_1030_n N_A_300_453#_c_1465_n 0.0275295f $X=5.75 $Y=2.75
+ $X2=0 $Y2=0
cc_731 N_A_1044_100#_c_1020_n N_VGND_c_1616_n 0.00140326f $X=7.49 $Y=0.995 $X2=0
+ $Y2=0
cc_732 N_A_1044_100#_c_1020_n N_VGND_c_1626_n 0.00278271f $X=7.49 $Y=0.995 $X2=0
+ $Y2=0
cc_733 N_A_1044_100#_c_1020_n N_VGND_c_1633_n 0.00361224f $X=7.49 $Y=0.995 $X2=0
+ $Y2=0
cc_734 N_A_1829_398#_M1021_g N_A_1592_424#_c_1227_n 0.0271894f $X=9.25 $Y=0.58
+ $X2=0 $Y2=0
cc_735 N_A_1829_398#_c_1131_n N_A_1592_424#_c_1227_n 0.00837726f $X=9.8 $Y=1.155
+ $X2=0 $Y2=0
cc_736 N_A_1829_398#_c_1133_n N_A_1592_424#_c_1227_n 0.0115382f $X=9.965
+ $Y=0.515 $X2=0 $Y2=0
cc_737 N_A_1829_398#_c_1134_n N_A_1592_424#_c_1227_n 0.00197213f $X=10.445
+ $Y=1.385 $X2=0 $Y2=0
cc_738 N_A_1829_398#_c_1124_n N_A_1592_424#_c_1228_n 0.0207424f $X=9.235 $Y=2.08
+ $X2=0 $Y2=0
cc_739 N_A_1829_398#_c_1138_n N_A_1592_424#_c_1228_n 0.00494332f $X=9.235
+ $Y=2.405 $X2=0 $Y2=0
cc_740 N_A_1829_398#_M1021_g N_A_1592_424#_c_1228_n 0.00518086f $X=9.25 $Y=0.58
+ $X2=0 $Y2=0
cc_741 N_A_1829_398#_c_1128_n N_A_1592_424#_c_1228_n 0.0112539f $X=10.93
+ $Y=1.385 $X2=0 $Y2=0
cc_742 N_A_1829_398#_c_1130_n N_A_1592_424#_c_1228_n 0.00625737f $X=9.37 $Y=1.74
+ $X2=0 $Y2=0
cc_743 N_A_1829_398#_c_1131_n N_A_1592_424#_c_1228_n 0.00547485f $X=9.8 $Y=1.155
+ $X2=0 $Y2=0
cc_744 N_A_1829_398#_c_1134_n N_A_1592_424#_c_1228_n 0.0134873f $X=10.445
+ $Y=1.385 $X2=0 $Y2=0
cc_745 N_A_1829_398#_c_1143_n N_A_1592_424#_c_1228_n 0.0136868f $X=10.26
+ $Y=2.665 $X2=0 $Y2=0
cc_746 N_A_1829_398#_c_1135_n N_A_1592_424#_c_1228_n 0.0200171f $X=10.27
+ $Y=2.415 $X2=0 $Y2=0
cc_747 N_A_1829_398#_c_1138_n N_A_1592_424#_c_1239_n 0.00423723f $X=9.235
+ $Y=2.405 $X2=0 $Y2=0
cc_748 N_A_1829_398#_c_1124_n N_A_1592_424#_c_1229_n 0.00207463f $X=9.235
+ $Y=2.08 $X2=0 $Y2=0
cc_749 N_A_1829_398#_M1021_g N_A_1592_424#_c_1229_n 0.0164674f $X=9.25 $Y=0.58
+ $X2=0 $Y2=0
cc_750 N_A_1829_398#_c_1130_n N_A_1592_424#_c_1229_n 0.0496022f $X=9.37 $Y=1.74
+ $X2=0 $Y2=0
cc_751 N_A_1829_398#_c_1132_n N_A_1592_424#_c_1229_n 0.0135848f $X=9.535
+ $Y=1.155 $X2=0 $Y2=0
cc_752 N_A_1829_398#_c_1137_n N_A_1592_424#_c_1234_n 0.00410845f $X=9.235
+ $Y=2.315 $X2=0 $Y2=0
cc_753 N_A_1829_398#_c_1138_n N_A_1592_424#_c_1234_n 0.00221096f $X=9.235
+ $Y=2.405 $X2=0 $Y2=0
cc_754 N_A_1829_398#_c_1124_n N_A_1592_424#_c_1235_n 0.00642866f $X=9.235
+ $Y=2.08 $X2=0 $Y2=0
cc_755 N_A_1829_398#_c_1137_n N_A_1592_424#_c_1235_n 0.0150636f $X=9.235
+ $Y=2.315 $X2=0 $Y2=0
cc_756 N_A_1829_398#_c_1130_n N_A_1592_424#_c_1235_n 0.0238629f $X=9.37 $Y=1.74
+ $X2=0 $Y2=0
cc_757 N_A_1829_398#_c_1143_n N_A_1592_424#_c_1235_n 7.0267e-19 $X=10.26
+ $Y=2.665 $X2=0 $Y2=0
cc_758 N_A_1829_398#_c_1135_n N_A_1592_424#_c_1235_n 0.0133619f $X=10.27
+ $Y=2.415 $X2=0 $Y2=0
cc_759 N_A_1829_398#_c_1124_n N_A_1592_424#_c_1230_n 0.00520692f $X=9.235
+ $Y=2.08 $X2=0 $Y2=0
cc_760 N_A_1829_398#_c_1130_n N_A_1592_424#_c_1230_n 0.0294108f $X=9.37 $Y=1.74
+ $X2=0 $Y2=0
cc_761 N_A_1829_398#_c_1131_n N_A_1592_424#_c_1230_n 0.00179416f $X=9.8 $Y=1.155
+ $X2=0 $Y2=0
cc_762 N_A_1829_398#_c_1134_n N_A_1592_424#_c_1230_n 0.0383463f $X=10.445
+ $Y=1.385 $X2=0 $Y2=0
cc_763 N_A_1829_398#_c_1135_n N_A_1592_424#_c_1230_n 0.0391131f $X=10.27
+ $Y=2.415 $X2=0 $Y2=0
cc_764 N_A_1829_398#_M1021_g N_A_1592_424#_c_1231_n 0.00213201f $X=9.25 $Y=0.58
+ $X2=0 $Y2=0
cc_765 N_A_1829_398#_c_1138_n N_VPWR_c_1319_n 0.0208784f $X=9.235 $Y=2.405 $X2=0
+ $Y2=0
cc_766 N_A_1829_398#_c_1143_n N_VPWR_c_1319_n 0.013366f $X=10.26 $Y=2.665 $X2=0
+ $Y2=0
cc_767 N_A_1829_398#_c_1139_n N_VPWR_c_1320_n 0.0100916f $X=11.045 $Y=1.765
+ $X2=0 $Y2=0
cc_768 N_A_1829_398#_c_1128_n N_VPWR_c_1320_n 0.00546342f $X=10.93 $Y=1.385
+ $X2=0 $Y2=0
cc_769 N_A_1829_398#_c_1185_p N_VPWR_c_1320_n 0.0148177f $X=10.88 $Y=1.385 $X2=0
+ $Y2=0
cc_770 N_A_1829_398#_c_1135_n N_VPWR_c_1320_n 0.0754487f $X=10.27 $Y=2.415 $X2=0
+ $Y2=0
cc_771 N_A_1829_398#_c_1140_n N_VPWR_c_1322_n 0.0100916f $X=11.495 $Y=1.765
+ $X2=0 $Y2=0
cc_772 N_A_1829_398#_c_1138_n N_VPWR_c_1329_n 0.00479724f $X=9.235 $Y=2.405
+ $X2=0 $Y2=0
cc_773 N_A_1829_398#_c_1143_n N_VPWR_c_1330_n 0.0123287f $X=10.26 $Y=2.665 $X2=0
+ $Y2=0
cc_774 N_A_1829_398#_c_1139_n N_VPWR_c_1331_n 0.00445602f $X=11.045 $Y=1.765
+ $X2=0 $Y2=0
cc_775 N_A_1829_398#_c_1140_n N_VPWR_c_1331_n 0.00445602f $X=11.495 $Y=1.765
+ $X2=0 $Y2=0
cc_776 N_A_1829_398#_c_1138_n N_VPWR_c_1315_n 0.00477621f $X=9.235 $Y=2.405
+ $X2=0 $Y2=0
cc_777 N_A_1829_398#_c_1139_n N_VPWR_c_1315_n 0.00862391f $X=11.045 $Y=1.765
+ $X2=0 $Y2=0
cc_778 N_A_1829_398#_c_1140_n N_VPWR_c_1315_n 0.00861084f $X=11.495 $Y=1.765
+ $X2=0 $Y2=0
cc_779 N_A_1829_398#_c_1143_n N_VPWR_c_1315_n 0.0122947f $X=10.26 $Y=2.665 $X2=0
+ $Y2=0
cc_780 N_A_1829_398#_c_1126_n N_Q_c_1590_n 0.00683953f $X=11.005 $Y=1.22 $X2=0
+ $Y2=0
cc_781 N_A_1829_398#_c_1127_n N_Q_c_1590_n 0.00293584f $X=11.48 $Y=1.22 $X2=0
+ $Y2=0
cc_782 N_A_1829_398#_c_1126_n N_Q_c_1596_n 0.00295571f $X=11.005 $Y=1.22 $X2=0
+ $Y2=0
cc_783 N_A_1829_398#_c_1129_n N_Q_c_1596_n 0.00217037f $X=11.48 $Y=1.492 $X2=0
+ $Y2=0
cc_784 N_A_1829_398#_c_1139_n Q 0.0144379f $X=11.045 $Y=1.765 $X2=0 $Y2=0
cc_785 N_A_1829_398#_c_1140_n Q 0.0144379f $X=11.495 $Y=1.765 $X2=0 $Y2=0
cc_786 N_A_1829_398#_c_1129_n Q 0.00164557f $X=11.48 $Y=1.492 $X2=0 $Y2=0
cc_787 N_A_1829_398#_c_1126_n N_Q_c_1591_n 0.00260601f $X=11.005 $Y=1.22 $X2=0
+ $Y2=0
cc_788 N_A_1829_398#_c_1140_n N_Q_c_1591_n 0.00172446f $X=11.495 $Y=1.765 $X2=0
+ $Y2=0
cc_789 N_A_1829_398#_c_1129_n N_Q_c_1591_n 0.0375743f $X=11.48 $Y=1.492 $X2=0
+ $Y2=0
cc_790 N_A_1829_398#_c_1185_p N_Q_c_1591_n 0.0249855f $X=10.88 $Y=1.385 $X2=0
+ $Y2=0
cc_791 N_A_1829_398#_c_1131_n N_VGND_M1021_d 0.00105556f $X=9.8 $Y=1.155 $X2=0
+ $Y2=0
cc_792 N_A_1829_398#_c_1132_n N_VGND_M1021_d 0.00147687f $X=9.535 $Y=1.155 $X2=0
+ $Y2=0
cc_793 N_A_1829_398#_M1021_g N_VGND_c_1617_n 0.0119193f $X=9.25 $Y=0.58 $X2=0
+ $Y2=0
cc_794 N_A_1829_398#_c_1131_n N_VGND_c_1617_n 0.00490389f $X=9.8 $Y=1.155 $X2=0
+ $Y2=0
cc_795 N_A_1829_398#_c_1132_n N_VGND_c_1617_n 0.0156223f $X=9.535 $Y=1.155 $X2=0
+ $Y2=0
cc_796 N_A_1829_398#_c_1133_n N_VGND_c_1617_n 0.0180508f $X=9.965 $Y=0.515 $X2=0
+ $Y2=0
cc_797 N_A_1829_398#_c_1126_n N_VGND_c_1618_n 0.00365549f $X=11.005 $Y=1.22
+ $X2=0 $Y2=0
cc_798 N_A_1829_398#_c_1128_n N_VGND_c_1618_n 0.00620972f $X=10.93 $Y=1.385
+ $X2=0 $Y2=0
cc_799 N_A_1829_398#_c_1133_n N_VGND_c_1618_n 0.0266944f $X=9.965 $Y=0.515 $X2=0
+ $Y2=0
cc_800 N_A_1829_398#_c_1185_p N_VGND_c_1618_n 0.0216379f $X=10.88 $Y=1.385 $X2=0
+ $Y2=0
cc_801 N_A_1829_398#_c_1127_n N_VGND_c_1620_n 0.00560767f $X=11.48 $Y=1.22 $X2=0
+ $Y2=0
cc_802 N_A_1829_398#_c_1129_n N_VGND_c_1620_n 0.00150639f $X=11.48 $Y=1.492
+ $X2=0 $Y2=0
cc_803 N_A_1829_398#_M1021_g N_VGND_c_1626_n 0.00383152f $X=9.25 $Y=0.58 $X2=0
+ $Y2=0
cc_804 N_A_1829_398#_c_1133_n N_VGND_c_1627_n 0.0145639f $X=9.965 $Y=0.515 $X2=0
+ $Y2=0
cc_805 N_A_1829_398#_c_1126_n N_VGND_c_1628_n 0.00434272f $X=11.005 $Y=1.22
+ $X2=0 $Y2=0
cc_806 N_A_1829_398#_c_1127_n N_VGND_c_1628_n 0.00460063f $X=11.48 $Y=1.22 $X2=0
+ $Y2=0
cc_807 N_A_1829_398#_M1021_g N_VGND_c_1633_n 0.0075725f $X=9.25 $Y=0.58 $X2=0
+ $Y2=0
cc_808 N_A_1829_398#_c_1126_n N_VGND_c_1633_n 0.00825492f $X=11.005 $Y=1.22
+ $X2=0 $Y2=0
cc_809 N_A_1829_398#_c_1127_n N_VGND_c_1633_n 0.00911274f $X=11.48 $Y=1.22 $X2=0
+ $Y2=0
cc_810 N_A_1829_398#_c_1133_n N_VGND_c_1633_n 0.0119984f $X=9.965 $Y=0.515 $X2=0
+ $Y2=0
cc_811 N_A_1592_424#_c_1235_n N_VPWR_M1032_d 0.00692596f $X=9.775 $Y=2.16 $X2=0
+ $Y2=0
cc_812 N_A_1592_424#_c_1230_n N_VPWR_M1032_d 0.00276332f $X=9.94 $Y=1.575 $X2=0
+ $Y2=0
cc_813 N_A_1592_424#_c_1228_n N_VPWR_c_1319_n 0.00419354f $X=10.035 $Y=1.825
+ $X2=0 $Y2=0
cc_814 N_A_1592_424#_c_1239_n N_VPWR_c_1319_n 0.00471635f $X=8.89 $Y=2.575 $X2=0
+ $Y2=0
cc_815 N_A_1592_424#_c_1235_n N_VPWR_c_1319_n 0.0287956f $X=9.775 $Y=2.16 $X2=0
+ $Y2=0
cc_816 N_A_1592_424#_c_1228_n N_VPWR_c_1320_n 0.00365662f $X=10.035 $Y=1.825
+ $X2=0 $Y2=0
cc_817 N_A_1592_424#_c_1239_n N_VPWR_c_1329_n 0.0119795f $X=8.89 $Y=2.575 $X2=0
+ $Y2=0
cc_818 N_A_1592_424#_c_1237_n N_VPWR_c_1329_n 0.00841934f $X=8.15 $Y=2.575 $X2=0
+ $Y2=0
cc_819 N_A_1592_424#_c_1228_n N_VPWR_c_1330_n 0.00520623f $X=10.035 $Y=1.825
+ $X2=0 $Y2=0
cc_820 N_A_1592_424#_c_1228_n N_VPWR_c_1315_n 0.00526787f $X=10.035 $Y=1.825
+ $X2=0 $Y2=0
cc_821 N_A_1592_424#_c_1239_n N_VPWR_c_1315_n 0.0219446f $X=8.89 $Y=2.575 $X2=0
+ $Y2=0
cc_822 N_A_1592_424#_c_1237_n N_VPWR_c_1315_n 0.00867391f $X=8.15 $Y=2.575 $X2=0
+ $Y2=0
cc_823 N_A_1592_424#_c_1239_n A_1704_496# 0.0210894f $X=8.89 $Y=2.575 $X2=-0.19
+ $Y2=-0.245
cc_824 N_A_1592_424#_c_1234_n A_1704_496# 3.02905e-19 $X=8.975 $Y=2.49 $X2=-0.19
+ $Y2=-0.245
cc_825 N_A_1592_424#_c_1227_n N_VGND_c_1617_n 0.00555396f $X=9.75 $Y=1.185 $X2=0
+ $Y2=0
cc_826 N_A_1592_424#_c_1231_n N_VGND_c_1617_n 0.0198687f $X=8.565 $Y=0.58 $X2=0
+ $Y2=0
cc_827 N_A_1592_424#_c_1231_n N_VGND_c_1626_n 0.0212211f $X=8.565 $Y=0.58 $X2=0
+ $Y2=0
cc_828 N_A_1592_424#_c_1227_n N_VGND_c_1627_n 0.00434272f $X=9.75 $Y=1.185 $X2=0
+ $Y2=0
cc_829 N_A_1592_424#_c_1227_n N_VGND_c_1633_n 0.00825771f $X=9.75 $Y=1.185 $X2=0
+ $Y2=0
cc_830 N_A_1592_424#_c_1231_n N_VGND_c_1633_n 0.0213723f $X=8.565 $Y=0.58 $X2=0
+ $Y2=0
cc_831 N_A_1592_424#_c_1231_n A_1787_74# 0.00272169f $X=8.565 $Y=0.58 $X2=-0.19
+ $Y2=-0.245
cc_832 N_VPWR_M1017_d N_A_300_453#_c_1468_n 0.0130974f $X=2.615 $Y=2.265 $X2=0
+ $Y2=0
cc_833 N_VPWR_c_1317_n N_A_300_453#_c_1468_n 0.0211438f $X=2.91 $Y=2.955 $X2=0
+ $Y2=0
cc_834 N_VPWR_c_1323_n N_A_300_453#_c_1468_n 0.0080152f $X=2.685 $Y=3.33 $X2=0
+ $Y2=0
cc_835 N_VPWR_c_1315_n N_A_300_453#_c_1468_n 0.0179485f $X=11.76 $Y=3.33 $X2=0
+ $Y2=0
cc_836 N_VPWR_M1017_d N_A_300_453#_c_1456_n 0.0142674f $X=2.615 $Y=2.265 $X2=0
+ $Y2=0
cc_837 N_VPWR_M1017_d N_A_300_453#_c_1462_n 0.00141021f $X=2.615 $Y=2.265 $X2=0
+ $Y2=0
cc_838 N_VPWR_M1027_s N_A_300_453#_c_1462_n 0.0160667f $X=3.92 $Y=1.84 $X2=0
+ $Y2=0
cc_839 N_VPWR_c_1317_n N_A_300_453#_c_1462_n 0.00105725f $X=2.91 $Y=2.955 $X2=0
+ $Y2=0
cc_840 N_VPWR_c_1328_n N_A_300_453#_c_1462_n 0.0106324f $X=3.9 $Y=3.33 $X2=0
+ $Y2=0
cc_841 N_VPWR_c_1333_n N_A_300_453#_c_1462_n 0.0322805f $X=4.135 $Y=2.955 $X2=0
+ $Y2=0
cc_842 N_VPWR_c_1315_n N_A_300_453#_c_1462_n 0.0216282f $X=11.76 $Y=3.33 $X2=0
+ $Y2=0
cc_843 N_VPWR_M1027_s N_A_300_453#_c_1457_n 0.0111284f $X=3.92 $Y=1.84 $X2=0
+ $Y2=0
cc_844 N_VPWR_c_1325_n N_A_300_453#_c_1464_n 0.00935318f $X=6.585 $Y=3.33 $X2=0
+ $Y2=0
cc_845 N_VPWR_c_1315_n N_A_300_453#_c_1464_n 0.0169876f $X=11.76 $Y=3.33 $X2=0
+ $Y2=0
cc_846 N_VPWR_c_1325_n N_A_300_453#_c_1465_n 0.010868f $X=6.585 $Y=3.33 $X2=0
+ $Y2=0
cc_847 N_VPWR_c_1315_n N_A_300_453#_c_1465_n 0.0090832f $X=11.76 $Y=3.33 $X2=0
+ $Y2=0
cc_848 N_VPWR_c_1316_n N_A_300_453#_c_1466_n 0.0179176f $X=0.78 $Y=2.44 $X2=0
+ $Y2=0
cc_849 N_VPWR_c_1317_n N_A_300_453#_c_1466_n 0.00464102f $X=2.91 $Y=2.955 $X2=0
+ $Y2=0
cc_850 N_VPWR_c_1323_n N_A_300_453#_c_1466_n 0.0221045f $X=2.685 $Y=3.33 $X2=0
+ $Y2=0
cc_851 N_VPWR_c_1315_n N_A_300_453#_c_1466_n 0.02058f $X=11.76 $Y=3.33 $X2=0
+ $Y2=0
cc_852 N_VPWR_M1017_d N_A_300_453#_c_1508_n 0.00415415f $X=2.615 $Y=2.265 $X2=0
+ $Y2=0
cc_853 N_VPWR_c_1317_n N_A_300_453#_c_1508_n 0.0145502f $X=2.91 $Y=2.955 $X2=0
+ $Y2=0
cc_854 N_VPWR_c_1315_n N_A_300_453#_c_1508_n 7.5402e-19 $X=11.76 $Y=3.33 $X2=0
+ $Y2=0
cc_855 N_VPWR_M1027_s N_A_300_453#_c_1544_n 8.28388e-19 $X=3.92 $Y=1.84 $X2=0
+ $Y2=0
cc_856 N_VPWR_c_1325_n N_A_300_453#_c_1544_n 0.00135165f $X=6.585 $Y=3.33 $X2=0
+ $Y2=0
cc_857 N_VPWR_c_1333_n N_A_300_453#_c_1544_n 0.00460666f $X=4.135 $Y=2.955 $X2=0
+ $Y2=0
cc_858 N_VPWR_c_1315_n N_A_300_453#_c_1544_n 0.00334631f $X=11.76 $Y=3.33 $X2=0
+ $Y2=0
cc_859 N_VPWR_c_1320_n Q 0.0778054f $X=10.82 $Y=1.985 $X2=0 $Y2=0
cc_860 N_VPWR_c_1322_n Q 0.0778054f $X=11.72 $Y=1.985 $X2=0 $Y2=0
cc_861 N_VPWR_c_1331_n Q 0.014552f $X=11.635 $Y=3.33 $X2=0 $Y2=0
cc_862 N_VPWR_c_1315_n Q 0.0119791f $X=11.76 $Y=3.33 $X2=0 $Y2=0
cc_863 N_A_300_453#_c_1468_n A_439_453# 0.00927389f $X=2.95 $Y=2.487 $X2=-0.19
+ $Y2=-0.245
cc_864 N_A_300_453#_c_1454_n N_VGND_M1000_d 0.00311051f $X=2.95 $Y=1.18 $X2=0
+ $Y2=0
cc_865 N_A_300_453#_c_1452_n N_VGND_c_1613_n 0.00971011f $X=2.375 $Y=0.515 $X2=0
+ $Y2=0
cc_866 N_A_300_453#_c_1452_n N_VGND_c_1614_n 0.0267569f $X=2.375 $Y=0.515 $X2=0
+ $Y2=0
cc_867 N_A_300_453#_c_1453_n N_VGND_c_1614_n 0.00943156f $X=2.46 $Y=1.095 $X2=0
+ $Y2=0
cc_868 N_A_300_453#_c_1454_n N_VGND_c_1614_n 0.0138324f $X=2.95 $Y=1.18 $X2=0
+ $Y2=0
cc_869 N_A_300_453#_c_1452_n N_VGND_c_1621_n 0.0445784f $X=2.375 $Y=0.515 $X2=0
+ $Y2=0
cc_870 N_A_300_453#_c_1452_n N_VGND_c_1633_n 0.0372402f $X=2.375 $Y=0.515 $X2=0
+ $Y2=0
cc_871 N_A_300_453#_c_1452_n A_442_74# 0.00442324f $X=2.375 $Y=0.515 $X2=-0.19
+ $Y2=-0.245
cc_872 N_A_300_453#_c_1453_n A_442_74# 0.00126008f $X=2.46 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_873 N_Q_c_1590_n N_VGND_c_1618_n 0.026995f $X=11.22 $Y=0.515 $X2=0 $Y2=0
cc_874 N_Q_c_1590_n N_VGND_c_1620_n 0.031377f $X=11.22 $Y=0.515 $X2=0 $Y2=0
cc_875 N_Q_c_1590_n N_VGND_c_1628_n 0.0145787f $X=11.22 $Y=0.515 $X2=0 $Y2=0
cc_876 N_Q_c_1590_n N_VGND_c_1633_n 0.0120042f $X=11.22 $Y=0.515 $X2=0 $Y2=0
