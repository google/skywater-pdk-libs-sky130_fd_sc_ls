* File: sky130_fd_sc_ls__dfrtp_1.spice
* Created: Wed Sep  2 11:01:06 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__dfrtp_1.pex.spice"
.subckt sky130_fd_sc_ls__dfrtp_1  VNB VPB D CLK RESET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* RESET_B	RESET_B
* CLK	CLK
* D	D
* VPB	VPB
* VNB	VNB
MM1020 A_117_78# N_D_M1020_g N_A_30_78#_M1020_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1008 N_VGND_M1008_d N_RESET_B_M1008_g A_117_78# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1030 N_VGND_M1030_d N_CLK_M1030_g N_A_306_96#_M1030_s VNB NSHORT L=0.15 W=0.74
+ AD=0.162375 AS=0.2646 PD=1.255 PS=2.4 NRD=9.72 NRS=5.268 M=1 R=4.93333
+ SA=75000.2 SB=75000.8 A=0.111 P=1.78 MULT=1
MM1025 N_A_490_390#_M1025_d N_A_306_96#_M1025_g N_VGND_M1030_d VNB NSHORT L=0.15
+ W=0.74 AD=0.2183 AS=0.162375 PD=2.07 PS=1.255 NRD=1.62 NRS=9.72 M=1 R=4.93333
+ SA=75000.8 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1031 N_A_695_457#_M1031_d N_A_306_96#_M1031_g N_A_30_78#_M1031_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0735 AS=0.1197 PD=0.77 PS=1.41 NRD=19.992 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75003.7 A=0.063 P=1.14 MULT=1
MM1027 A_816_138# N_A_490_390#_M1027_g N_A_695_457#_M1031_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.0735 PD=0.66 PS=0.77 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75000.7 SB=75003.2 A=0.063 P=1.14 MULT=1
MM1012 A_894_138# N_A_830_359#_M1012_g A_816_138# VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0504 PD=0.66 PS=0.66 NRD=18.564 NRS=18.564 M=1 R=2.8 SA=75001.1
+ SB=75002.8 A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_RESET_B_M1004_g A_894_138# VNB NSHORT L=0.15 W=0.42
+ AD=0.152965 AS=0.0504 PD=1.05 PS=0.66 NRD=88.332 NRS=18.564 M=1 R=2.8
+ SA=75001.5 SB=75002.4 A=0.063 P=1.14 MULT=1
MM1026 N_A_830_359#_M1026_d N_A_695_457#_M1026_g N_VGND_M1004_d VNB NSHORT
+ L=0.15 W=0.74 AD=0.24605 AS=0.26951 PD=1.405 PS=1.85 NRD=22.296 NRS=50.136 M=1
+ R=4.93333 SA=75001.4 SB=75002.3 A=0.111 P=1.78 MULT=1
MM1022 N_A_1266_74#_M1022_d N_A_490_390#_M1022_g N_A_830_359#_M1026_d VNB NSHORT
+ L=0.15 W=0.74 AD=0.292172 AS=0.24605 PD=2.09241 PS=1.405 NRD=2.424 NRS=8.916
+ M=1 R=4.93333 SA=75002.2 SB=75001.5 A=0.111 P=1.78 MULT=1
MM1016 A_1476_81# N_A_306_96#_M1016_g N_A_1266_74#_M1022_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.165828 PD=0.66 PS=1.18759 NRD=18.564 NRS=49.992 M=1
+ R=2.8 SA=75002.8 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1014 N_VGND_M1014_d N_A_1518_203#_M1014_g A_1476_81# VNB NSHORT L=0.15 W=0.42
+ AD=0.0756 AS=0.0504 PD=0.78 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75003.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1028 A_1656_81# N_RESET_B_M1028_g N_VGND_M1014_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0756 PD=0.63 PS=0.78 NRD=14.28 NRS=22.848 M=1 R=2.8 SA=75003.7
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1017 N_A_1518_203#_M1017_d N_A_1266_74#_M1017_g A_1656_81# VNB NSHORT L=0.15
+ W=0.42 AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8
+ SA=75004.1 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1023 N_A_1864_409#_M1023_d N_A_1266_74#_M1023_g N_VGND_M1023_s VNB NSHORT
+ L=0.15 W=0.55 AD=0.15675 AS=0.15675 PD=1.67 PS=1.67 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1002 N_VGND_M1002_d N_A_1864_409#_M1002_g N_Q_M1002_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.2109 PD=2.05 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1018 N_A_30_78#_M1018_d N_D_M1018_g N_VPWR_M1018_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.05985 AS=0.1197 PD=0.705 PS=1.41 NRD=2.3443 NRS=4.6886 M=1 R=2.8
+ SA=75000.2 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1000 N_VPWR_M1000_d N_RESET_B_M1000_g N_A_30_78#_M1018_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.05985 PD=1.37 PS=0.705 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1006 N_VPWR_M1006_d N_CLK_M1006_g N_A_306_96#_M1006_s VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.31 PD=1.3 PS=2.62 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75000.2
+ SB=75000.7 A=0.15 P=2.3 MULT=1
MM1011 N_A_490_390#_M1011_d N_A_306_96#_M1011_g N_VPWR_M1006_d VPB PHIGHVT
+ L=0.15 W=1 AD=0.285 AS=0.15 PD=2.57 PS=1.3 NRD=3.9203 NRS=1.9503 M=1 R=6.66667
+ SA=75000.7 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1009 N_A_695_457#_M1009_d N_A_490_390#_M1009_g N_A_30_78#_M1009_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.063 AS=0.1218 PD=0.72 PS=1.42 NRD=4.6886 NRS=4.6886 M=1
+ R=2.8 SA=75000.2 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1019 A_785_457# N_A_306_96#_M1019_g N_A_695_457#_M1009_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0504 AS=0.063 PD=0.66 PS=0.72 NRD=30.4759 NRS=4.6886 M=1 R=2.8
+ SA=75000.7 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1003 N_VPWR_M1003_d N_A_830_359#_M1003_g A_785_457# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.137125 AS=0.0504 PD=1.155 PS=0.66 NRD=127.341 NRS=30.4759 M=1 R=2.8
+ SA=75001.1 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1029 N_A_695_457#_M1029_d N_RESET_B_M1029_g N_VPWR_M1003_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1239 AS=0.137125 PD=1.43 PS=1.155 NRD=4.6886 NRS=127.341 M=1 R=2.8
+ SA=75001.7 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1005 N_A_830_359#_M1005_d N_A_695_457#_M1005_g N_VPWR_M1005_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.190625 AS=0.305 PD=1.505 PS=2.61 NRD=9.8303 NRS=3.9203 M=1
+ R=6.66667 SA=75000.2 SB=75001.4 A=0.15 P=2.3 MULT=1
MM1015 N_A_1266_74#_M1015_d N_A_306_96#_M1015_g N_A_830_359#_M1005_d VPB PHIGHVT
+ L=0.15 W=1 AD=0.324155 AS=0.190625 PD=2.43662 PS=1.505 NRD=8.8453 NRS=4.9053
+ M=1 R=6.66667 SA=75000.7 SB=75001.4 A=0.15 P=2.3 MULT=1
MM1001 A_1468_493# N_A_490_390#_M1001_g N_A_1266_74#_M1015_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0567 AS=0.136145 PD=0.69 PS=1.02338 NRD=37.5088 NRS=4.6886 M=1
+ R=2.8 SA=75001.4 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1024 N_VPWR_M1024_d N_A_1518_203#_M1024_g A_1468_493# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.08925 AS=0.0567 PD=0.845 PS=0.69 NRD=32.8202 NRS=37.5088 M=1 R=2.8
+ SA=75001.8 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1010 N_A_1518_203#_M1010_d N_RESET_B_M1010_g N_VPWR_M1024_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.063 AS=0.08925 PD=0.72 PS=0.845 NRD=4.6886 NRS=35.1645 M=1 R=2.8
+ SA=75002.4 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1021 N_VPWR_M1021_d N_A_1266_74#_M1021_g N_A_1518_203#_M1010_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0952 AS=0.063 PD=0.816667 PS=0.72 NRD=44.5417 NRS=4.6886
+ M=1 R=2.8 SA=75002.9 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1013 N_A_1864_409#_M1013_d N_A_1266_74#_M1013_g N_VPWR_M1021_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.2478 AS=0.1904 PD=2.27 PS=1.63333 NRD=2.3443 NRS=2.3443 M=1
+ R=5.6 SA=75001.8 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1007 N_VPWR_M1007_d N_A_1864_409#_M1007_g N_Q_M1007_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.336 AS=0.3808 PD=2.84 PS=2.92 NRD=2.6201 NRS=9.6727 M=1 R=7.46667
+ SA=75000.3 SB=75000.2 A=0.168 P=2.54 MULT=1
DX32_noxref VNB VPB NWDIODE A=21.2956 P=26.8
c_237 VPB 0 1.4888e-19 $X=0 $Y=3.085
c_1760 A_1468_493# 0 1.01622e-19 $X=7.34 $Y=2.465
*
.include "sky130_fd_sc_ls__dfrtp_1.pxi.spice"
*
.ends
*
*
