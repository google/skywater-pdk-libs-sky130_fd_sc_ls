* NGSPICE file created from sky130_fd_sc_ls__a32oi_2.ext - technology: sky130A

.subckt sky130_fd_sc_ls__a32oi_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
M1000 a_27_368# A2 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=2.3184e+12p pd=1.758e+07u as=1.6296e+12p ps=9.63e+06u
M1001 VPWR A2 a_27_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_771_74# A3 VGND VNB nshort w=740000u l=150000u
+  ad=4.995e+11p pd=4.31e+06u as=6.66e+11p ps=6.24e+06u
M1003 Y B1 a_27_74# VNB nshort w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=6.808e+11p ps=6.28e+06u
M1004 VPWR A1 a_27_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y A1 a_507_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=6.475e+11p ps=6.19e+06u
M1006 VGND A3 a_771_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y B2 a_27_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=7.784e+11p pd=5.87e+06u as=0p ps=0u
M1008 a_27_74# B1 Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_27_368# B2 Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_27_74# B2 VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR A3 a_27_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_27_368# A3 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_507_74# A2 a_771_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_771_74# A2 a_507_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y B1 a_27_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND B2 a_27_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_27_368# A1 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_507_74# A1 Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_27_368# B1 Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

