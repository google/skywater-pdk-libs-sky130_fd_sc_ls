* File: sky130_fd_sc_ls__dfsbp_1.spice
* Created: Fri Aug 28 13:14:58 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__dfsbp_1.pex.spice"
.subckt sky130_fd_sc_ls__dfsbp_1  VNB VPB D CLK SET_B VPWR Q_N Q VGND
* 
* VGND	VGND
* Q	Q
* Q_N	Q_N
* VPWR	VPWR
* SET_B	SET_B
* CLK	CLK
* D	D
* VPB	VPB
* VNB	VNB
MM1002 N_VGND_M1002_d N_D_M1002_g N_A_27_80#_M1002_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.1197 PD=1.41 PS=1.41 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1029 N_VGND_M1029_d N_CLK_M1029_g N_A_225_74#_M1029_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1012 N_A_398_74#_M1012_d N_A_225_74#_M1012_g N_VGND_M1029_d VNB NSHORT L=0.15
+ W=0.74 AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1003 N_A_596_81#_M1003_d N_A_225_74#_M1003_g N_A_27_80#_M1003_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.1281 AS=0.1197 PD=1.03 PS=1.41 NRD=94.284 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1019 A_748_81# N_A_398_74#_M1019_g N_A_596_81#_M1003_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.1281 PD=0.66 PS=1.03 NRD=18.564 NRS=0 M=1 R=2.8 SA=75001
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1007 N_VGND_M1007_d N_A_779_380#_M1007_g A_748_81# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1013 A_1061_74# N_A_596_81#_M1013_g N_A_779_380#_M1013_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.1113 PD=0.66 PS=1.37 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75003.9 A=0.063 P=1.14 MULT=1
MM1024 N_VGND_M1024_d N_SET_B_M1024_g A_1061_74# VNB NSHORT L=0.15 W=0.42
+ AD=0.102226 AS=0.0504 PD=0.87566 PS=0.66 NRD=53.568 NRS=18.564 M=1 R=2.8
+ SA=75000.6 SB=75003.5 A=0.063 P=1.14 MULT=1
MM1033 A_1262_74# N_A_596_81#_M1033_g N_VGND_M1024_d VNB NSHORT L=0.15 W=0.64
+ AD=0.1088 AS=0.155774 PD=0.98 PS=1.33434 NRD=21.552 NRS=0 M=1 R=4.26667
+ SA=75000.9 SB=75002.1 A=0.096 P=1.58 MULT=1
MM1014 N_A_1355_377#_M1014_d N_A_398_74#_M1014_g A_1262_74# VNB NSHORT L=0.15
+ W=0.64 AD=0.129147 AS=0.1088 PD=1.20755 PS=0.98 NRD=0 NRS=21.552 M=1 R=4.26667
+ SA=75001.3 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1027 A_1462_74# N_A_225_74#_M1027_g N_A_1355_377#_M1014_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.0847528 PD=0.66 PS=0.792453 NRD=18.564 NRS=24.276 M=1
+ R=2.8 SA=75002.2 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1026 A_1540_74# N_A_1510_48#_M1026_g A_1462_74# VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0504 PD=0.66 PS=0.66 NRD=18.564 NRS=18.564 M=1 R=2.8 SA=75002.6
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1022 N_VGND_M1022_d N_SET_B_M1022_g A_1540_74# VNB NSHORT L=0.15 W=0.42
+ AD=0.1491 AS=0.0504 PD=1.13 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75003
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1011 N_A_1510_48#_M1011_d N_A_1355_377#_M1011_g N_VGND_M1022_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.1197 AS=0.1491 PD=1.41 PS=1.13 NRD=0 NRS=19.992 M=1 R=2.8
+ SA=75003.8 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1010 N_Q_N_M1010_d N_A_1355_377#_M1010_g N_VGND_M1010_s VNB NSHORT L=0.15
+ W=0.74 AD=0.2109 AS=0.2627 PD=2.05 PS=2.19 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75000.3 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1023 N_VGND_M1023_d N_A_1355_377#_M1023_g N_A_2113_74#_M1023_s VNB NSHORT
+ L=0.15 W=0.55 AD=0.129591 AS=0.15675 PD=0.997674 PS=1.67 NRD=17.988 NRS=0 M=1
+ R=3.66667 SA=75000.2 SB=75000.8 A=0.0825 P=1.4 MULT=1
MM1018 N_Q_M1018_d N_A_2113_74#_M1018_g N_VGND_M1023_d VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.174359 PD=2.05 PS=1.34233 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75000.7 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1016 N_VPWR_M1016_d N_D_M1016_g N_A_27_80#_M1016_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1239 AS=0.1239 PD=1.43 PS=1.43 NRD=4.6886 NRS=4.6886 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1028 N_VPWR_M1028_d N_CLK_M1028_g N_A_225_74#_M1028_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1001 N_A_398_74#_M1001_d N_A_225_74#_M1001_g N_VPWR_M1028_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1000 N_A_596_81#_M1000_d N_A_398_74#_M1000_g N_A_27_80#_M1000_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0735 AS=0.1239 PD=0.77 PS=1.43 NRD=28.1316 NRS=4.6886 M=1
+ R=2.8 SA=75000.2 SB=75004.4 A=0.063 P=1.14 MULT=1
MM1004 A_728_463# N_A_225_74#_M1004_g N_A_596_81#_M1000_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0567 AS=0.0735 PD=0.69 PS=0.77 NRD=37.5088 NRS=4.6886 M=1 R=2.8
+ SA=75000.7 SB=75003.9 A=0.063 P=1.14 MULT=1
MM1032 N_VPWR_M1032_d N_A_779_380#_M1032_g A_728_463# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.15855 AS=0.0567 PD=1.175 PS=0.69 NRD=18.7544 NRS=37.5088 M=1 R=2.8
+ SA=75001.1 SB=75003.5 A=0.063 P=1.14 MULT=1
MM1008 N_A_779_380#_M1008_d N_A_596_81#_M1008_g N_VPWR_M1032_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0756 AS=0.15855 PD=0.78 PS=1.175 NRD=4.6886 NRS=204.033 M=1
+ R=2.8 SA=75002 SB=75002.6 A=0.063 P=1.14 MULT=1
MM1005 N_VPWR_M1005_d N_SET_B_M1005_g N_A_779_380#_M1008_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.131635 AS=0.0756 PD=1.01451 PS=0.78 NRD=105.533 NRS=32.8202 M=1
+ R=2.8 SA=75002.6 SB=75002.1 A=0.063 P=1.14 MULT=1
MM1006 A_1254_341# N_A_596_81#_M1006_g N_VPWR_M1005_d VPB PHIGHVT L=0.15 W=1
+ AD=0.19325 AS=0.313415 PD=1.535 PS=2.41549 NRD=27.2254 NRS=28.5453 M=1
+ R=6.66667 SA=75001.4 SB=75000.9 A=0.15 P=2.3 MULT=1
MM1020 N_A_1355_377#_M1020_d N_A_225_74#_M1020_g A_1254_341# VPB PHIGHVT L=0.15
+ W=1 AD=0.310423 AS=0.19325 PD=2.44366 PS=1.535 NRD=1.9503 NRS=27.2254 M=1
+ R=6.66667 SA=75001.8 SB=75000.8 A=0.15 P=2.3 MULT=1
MM1030 A_1517_508# N_A_398_74#_M1030_g N_A_1355_377#_M1020_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0567 AS=0.130377 PD=0.69 PS=1.02634 NRD=37.5088 NRS=4.6886 M=1
+ R=2.8 SA=75002.3 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1021 N_VPWR_M1021_d N_A_1510_48#_M1021_g A_1517_508# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.063 AS=0.0567 PD=0.72 PS=0.69 NRD=4.6886 NRS=37.5088 M=1 R=2.8 SA=75002.7
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1031 N_A_1355_377#_M1031_d N_SET_B_M1031_g N_VPWR_M1021_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1239 AS=0.063 PD=1.43 PS=0.72 NRD=4.6886 NRS=4.6886 M=1 R=2.8
+ SA=75003.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1009 N_VPWR_M1009_d N_A_1355_377#_M1009_g N_A_1510_48#_M1009_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0912545 AS=0.1596 PD=0.804545 PS=1.6 NRD=21.0987
+ NRS=44.5417 M=1 R=2.8 SA=75000.3 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1017 N_Q_N_M1017_d N_A_1355_377#_M1017_g N_VPWR_M1009_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.3304 AS=0.243345 PD=2.83 PS=2.14545 NRD=1.7533 NRS=5.2599 M=1
+ R=7.46667 SA=75000.4 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1025 N_VPWR_M1025_d N_A_1355_377#_M1025_g N_A_2113_74#_M1025_s VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.1596 AS=0.2478 PD=1.26429 PS=2.27 NRD=2.3443 NRS=2.3443 M=1
+ R=5.6 SA=75000.2 SB=75000.7 A=0.126 P=1.98 MULT=1
MM1015 N_Q_M1015_d N_A_2113_74#_M1015_g N_VPWR_M1025_d VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.2128 PD=2.83 PS=1.68571 NRD=1.7533 NRS=11.426 M=1 R=7.46667
+ SA=75000.6 SB=75000.2 A=0.168 P=2.54 MULT=1
DX34_noxref VNB VPB NWDIODE A=23.4027 P=28.75
c_1799 A_728_463# 0 1.69669e-19 $X=3.64 $Y=2.315
*
.include "sky130_fd_sc_ls__dfsbp_1.pxi.spice"
*
.ends
*
*
