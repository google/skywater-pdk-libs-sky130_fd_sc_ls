* File: sky130_fd_sc_ls__dfstp_1.spice
* Created: Fri Aug 28 13:15:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__dfstp_1.pex.spice"
.subckt sky130_fd_sc_ls__dfstp_1  VNB VPB D CLK SET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* SET_B	SET_B
* CLK	CLK
* D	D
* VPB	VPB
* VNB	VNB
MM1024 N_VGND_M1024_d N_D_M1024_g N_A_27_74#_M1024_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.1197 PD=1.41 PS=1.41 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1026 N_VGND_M1026_d N_CLK_M1026_g N_A_224_350#_M1026_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1015 N_A_398_74#_M1015_d N_A_224_350#_M1015_g N_VGND_M1026_d VNB NSHORT L=0.15
+ W=0.74 AD=0.1961 AS=0.1036 PD=2.01 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1010 N_A_604_74#_M1010_d N_A_224_350#_M1010_g N_A_27_74#_M1010_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.1113 AS=0.17595 PD=0.95 PS=1.76 NRD=71.424 NRS=24.276 M=1
+ R=2.8 SA=75000.3 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1022 A_740_74# N_A_398_74#_M1022_g N_A_604_74#_M1010_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.1113 PD=0.66 PS=0.95 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75000.9 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1017 N_VGND_M1017_d N_A_760_395#_M1017_g A_740_74# VNB NSHORT L=0.15 W=0.42
+ AD=0.1449 AS=0.0504 PD=1.53 PS=0.66 NRD=8.568 NRS=18.564 M=1 R=2.8 SA=75001.3
+ SB=75000.3 A=0.063 P=1.14 MULT=1
MM1009 A_1027_118# N_A_604_74#_M1009_g N_A_760_395#_M1009_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.1176 PD=0.63 PS=1.4 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.8 A=0.063 P=1.14 MULT=1
MM1008 N_VGND_M1008_d N_SET_B_M1008_g A_1027_118# VNB NSHORT L=0.15 W=0.42
+ AD=0.0964019 AS=0.0441 PD=0.847925 PS=0.63 NRD=43.56 NRS=14.28 M=1 R=2.8
+ SA=75000.6 SB=75002.4 A=0.063 P=1.14 MULT=1
MM1030 A_1215_74# N_A_604_74#_M1030_g N_VGND_M1008_d VNB NSHORT L=0.15 W=0.64
+ AD=0.12 AS=0.146898 PD=1.015 PS=1.29208 NRD=24.84 NRS=0 M=1 R=4.26667
+ SA=75000.8 SB=75002.3 A=0.096 P=1.58 MULT=1
MM1006 N_A_1298_392#_M1006_d N_A_398_74#_M1006_g A_1215_74# VNB NSHORT L=0.15
+ W=0.64 AD=0.129147 AS=0.12 PD=1.20755 PS=1.015 NRD=0 NRS=24.84 M=1 R=4.26667
+ SA=75001.3 SB=75001.8 A=0.096 P=1.58 MULT=1
MM1013 A_1422_74# N_A_224_350#_M1013_g N_A_1298_392#_M1006_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.0847528 PD=0.66 PS=0.792453 NRD=18.564 NRS=24.276 M=1
+ R=2.8 SA=75001.7 SB=75002.1 A=0.063 P=1.14 MULT=1
MM1014 A_1500_74# N_A_1470_48#_M1014_g A_1422_74# VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0504 PD=0.66 PS=0.66 NRD=18.564 NRS=18.564 M=1 R=2.8 SA=75002.1
+ SB=75001.7 A=0.063 P=1.14 MULT=1
MM1020 N_VGND_M1020_d N_SET_B_M1020_g A_1500_74# VNB NSHORT L=0.15 W=0.42
+ AD=0.19215 AS=0.0504 PD=1.335 PS=0.66 NRD=1.428 NRS=18.564 M=1 R=2.8
+ SA=75002.5 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1005 N_A_1470_48#_M1005_d N_A_1298_392#_M1005_g N_VGND_M1020_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.1197 AS=0.19215 PD=1.41 PS=1.335 NRD=0 NRS=19.992 M=1 R=2.8
+ SA=75003.5 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1023 N_VGND_M1023_d N_A_1298_392#_M1023_g N_A_1902_74#_M1023_s VNB NSHORT
+ L=0.15 W=0.55 AD=0.129591 AS=0.15675 PD=0.997674 PS=1.67 NRD=17.988 NRS=0 M=1
+ R=3.66667 SA=75000.2 SB=75000.8 A=0.0825 P=1.4 MULT=1
MM1012 N_Q_M1012_d N_A_1902_74#_M1012_g N_VGND_M1023_d VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.174359 PD=2.05 PS=1.34233 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75000.7 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1021 N_VPWR_M1021_d N_D_M1021_g N_A_27_74#_M1021_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1176 AS=0.1197 PD=1.4 PS=1.41 NRD=4.6886 NRS=4.6886 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1000 N_VPWR_M1000_d N_CLK_M1000_g N_A_224_350#_M1000_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.3192 PD=1.42 PS=2.81 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1011 N_A_398_74#_M1011_d N_A_224_350#_M1011_g N_VPWR_M1000_d VPB PHIGHVT
+ L=0.15 W=1.12 AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1
+ R=7.46667 SA=75000.7 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1027 N_A_604_74#_M1027_d N_A_398_74#_M1027_g N_A_27_74#_M1027_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0735 AS=0.1239 PD=0.77 PS=1.43 NRD=28.1316 NRS=4.6886 M=1
+ R=2.8 SA=75000.2 SB=75004.2 A=0.063 P=1.14 MULT=1
MM1007 A_709_463# N_A_224_350#_M1007_g N_A_604_74#_M1027_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0567 AS=0.0735 PD=0.69 PS=0.77 NRD=37.5088 NRS=4.6886 M=1 R=2.8
+ SA=75000.7 SB=75003.7 A=0.063 P=1.14 MULT=1
MM1028 N_VPWR_M1028_d N_A_760_395#_M1028_g A_709_463# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.14175 AS=0.0567 PD=1.095 PS=0.69 NRD=11.7215 NRS=37.5088 M=1 R=2.8
+ SA=75001.1 SB=75003.3 A=0.063 P=1.14 MULT=1
MM1029 N_A_760_395#_M1029_d N_A_604_74#_M1029_g N_VPWR_M1028_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.063 AS=0.14175 PD=0.72 PS=1.095 NRD=4.6886 NRS=173.537 M=1
+ R=2.8 SA=75002 SB=75002.5 A=0.063 P=1.14 MULT=1
MM1001 N_VPWR_M1001_d N_SET_B_M1001_g N_A_760_395#_M1029_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.139694 AS=0.063 PD=1.10028 PS=0.72 NRD=130.197 NRS=4.6886 M=1
+ R=2.8 SA=75002.4 SB=75002 A=0.063 P=1.14 MULT=1
MM1018 A_1197_341# N_A_604_74#_M1018_g N_VPWR_M1001_d VPB PHIGHVT L=0.15 W=1
+ AD=0.199812 AS=0.332606 PD=1.61 PS=2.61972 NRD=28.5256 NRS=54.6872 M=1
+ R=6.66667 SA=75001.3 SB=75000.9 A=0.15 P=2.3 MULT=1
MM1019 N_A_1298_392#_M1019_d N_A_224_350#_M1019_g A_1197_341# VPB PHIGHVT L=0.15
+ W=1 AD=0.305141 AS=0.199812 PD=2.3169 PS=1.61 NRD=2.2852 NRS=28.5256 M=1
+ R=6.66667 SA=75001.7 SB=75000.9 A=0.15 P=2.3 MULT=1
MM1002 A_1457_508# N_A_398_74#_M1002_g N_A_1298_392#_M1019_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0567 AS=0.128159 PD=0.69 PS=0.973099 NRD=37.5088 NRS=86.7588 M=1
+ R=2.8 SA=75002.4 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1025 N_VPWR_M1025_d N_A_1470_48#_M1025_g A_1457_508# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.063 AS=0.0567 PD=0.72 PS=0.69 NRD=4.6886 NRS=37.5088 M=1 R=2.8 SA=75002.8
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1003 N_A_1298_392#_M1003_d N_SET_B_M1003_g N_VPWR_M1025_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1155 AS=0.063 PD=1.39 PS=0.72 NRD=4.6886 NRS=4.6886 M=1 R=2.8
+ SA=75003.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1016 N_A_1470_48#_M1016_d N_A_1298_392#_M1016_g N_VPWR_M1016_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.1155 AS=0.1176 PD=1.39 PS=1.4 NRD=4.6886 NRS=4.6886 M=1
+ R=2.8 SA=75000.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1031 N_VPWR_M1031_d N_A_1298_392#_M1031_g N_A_1902_74#_M1031_s VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.1668 AS=0.231 PD=1.27714 PS=2.23 NRD=35.7555 NRS=0 M=1
+ R=5.6 SA=75000.2 SB=75000.7 A=0.126 P=1.98 MULT=1
MM1004 N_Q_M1004_d N_A_1902_74#_M1004_g N_VPWR_M1031_d VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3192 AS=0.2224 PD=2.81 PS=1.70286 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.6 SB=75000.2 A=0.168 P=2.54 MULT=1
DX32_noxref VNB VPB NWDIODE A=21.7821 P=26.83
c_1667 A_1197_341# 0 1.10875e-19 $X=5.985 $Y=1.705
*
.include "sky130_fd_sc_ls__dfstp_1.pxi.spice"
*
.ends
*
*
