* File: sky130_fd_sc_ls__a211oi_2.spice
* Created: Wed Sep  2 10:47:39 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__a211oi_2.pex.spice"
.subckt sky130_fd_sc_ls__a211oi_2  VNB VPB A1 A2 B1 C1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* C1	C1
* B1	B1
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1008 N_Y_M1008_d N_A1_M1008_g N_A_38_74#_M1008_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1961 PD=1.02 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1010 N_Y_M1008_d N_A1_M1010_g N_A_38_74#_M1010_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1001 N_A_38_74#_M1010_s N_A2_M1001_g N_VGND_M1001_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1184 PD=1.02 PS=1.06 NRD=0 NRS=3.24 M=1 R=4.93333 SA=75001.1
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1003 N_A_38_74#_M1003_d N_A2_M1003_g N_VGND_M1001_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2183 AS=0.1184 PD=2.07 PS=1.06 NRD=0 NRS=3.24 M=1 R=4.93333 SA=75001.5
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1002 N_Y_M1002_d N_B1_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2664 AS=0.1961 PD=1.46 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1006 N_VGND_M1006_d N_C1_M1006_g N_Y_M1002_d VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.2664 PD=2.05 PS=1.46 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.1
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1011 N_A_114_368#_M1011_d N_A1_M1011_g N_VPWR_M1011_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.308 PD=1.42 PS=2.79 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1012 N_A_114_368#_M1011_d N_A1_M1012_g N_VPWR_M1012_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.6 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1000 N_A_114_368#_M1000_d N_A2_M1000_g N_VPWR_M1012_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1005 N_A_114_368#_M1000_d N_A2_M1005_g N_VPWR_M1005_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.5 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1007 N_A_114_368#_M1007_d N_B1_M1007_g N_A_497_368#_M1007_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75001.5 A=0.168 P=2.54 MULT=1
MM1009 N_A_114_368#_M1007_d N_B1_M1009_g N_A_497_368#_M1009_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1004 N_A_497_368#_M1009_s N_C1_M1004_g N_Y_M1004_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75000.6 A=0.168 P=2.54 MULT=1
MM1013 N_A_497_368#_M1013_d N_C1_M1013_g N_Y_M1004_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.308 AS=0.168 PD=2.79 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.6 SB=75000.2 A=0.168 P=2.54 MULT=1
DX14_noxref VNB VPB NWDIODE A=9.6348 P=14.08
*
.include "sky130_fd_sc_ls__a211oi_2.pxi.spice"
*
.ends
*
*
