* File: sky130_fd_sc_ls__o31ai_2.spice
* Created: Fri Aug 28 13:53:37 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__o31ai_2.pex.spice"
.subckt sky130_fd_sc_ls__o31ai_2  VNB VPB A1 A2 A3 B1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1	B1
* A3	A3
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1012 N_VGND_M1012_d N_A1_M1012_g N_A_27_74#_M1012_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1554 AS=0.2109 PD=1.16 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75004 A=0.111 P=1.78 MULT=1
MM1014 N_VGND_M1012_d N_A1_M1014_g N_A_27_74#_M1014_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1554 AS=0.1036 PD=1.16 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.8
+ SB=75003.4 A=0.111 P=1.78 MULT=1
MM1004 N_VGND_M1004_d N_A2_M1004_g N_A_27_74#_M1014_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1554 AS=0.1036 PD=1.16 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75001.2
+ SB=75003 A=0.111 P=1.78 MULT=1
MM1011 N_VGND_M1004_d N_A2_M1011_g N_A_27_74#_M1011_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1554 AS=0.1036 PD=1.16 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75001.8
+ SB=75002.4 A=0.111 P=1.78 MULT=1
MM1001 N_VGND_M1001_d N_A3_M1001_g N_A_27_74#_M1011_s VNB NSHORT L=0.15 W=0.74
+ AD=0.32 AS=0.1036 PD=1.645 PS=1.02 NRD=61.2 NRS=0 M=1 R=4.93333 SA=75002.2
+ SB=75002 A=0.111 P=1.78 MULT=1
MM1002 N_VGND_M1001_d N_A3_M1002_g N_A_27_74#_M1002_s VNB NSHORT L=0.15 W=0.74
+ AD=0.32 AS=0.1036 PD=1.645 PS=1.02 NRD=61.2 NRS=0 M=1 R=4.93333 SA=75003.1
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1007 N_Y_M1007_d N_B1_M1007_g N_A_27_74#_M1002_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1221 AS=0.1036 PD=1.07 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75003.5
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1008 N_Y_M1007_d N_B1_M1008_g N_A_27_74#_M1008_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1221 AS=0.2257 PD=1.07 PS=2.09 NRD=8.1 NRS=3.24 M=1 R=4.93333 SA=75004
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1005 N_VPWR_M1005_d N_A1_M1005_g N_A_28_368#_M1005_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1006 N_VPWR_M1005_d N_A1_M1006_g N_A_28_368#_M1006_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1010 N_A_297_368#_M1010_d N_A2_M1010_g N_A_28_368#_M1006_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1015 N_A_297_368#_M1010_d N_A2_M1015_g N_A_28_368#_M1015_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.6 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1009 N_A_297_368#_M1009_d N_A3_M1009_g N_Y_M1009_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1013 N_A_297_368#_M1009_d N_A3_M1013_g N_Y_M1013_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75000.7 SB=75001.2 A=0.168 P=2.54 MULT=1
MM1000 N_VPWR_M1000_d N_B1_M1000_g N_Y_M1013_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.2 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1003 N_VPWR_M1000_d N_B1_M1003_g N_Y_M1003_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.6 SB=75000.2 A=0.168 P=2.54 MULT=1
DX16_noxref VNB VPB NWDIODE A=9.6348 P=14.08
c_80 VPB 0 1.34959e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_ls__o31ai_2.pxi.spice"
*
.ends
*
*
