* File: sky130_fd_sc_ls__xnor3_2.pex.spice
* Created: Fri Aug 28 14:09:40 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__XNOR3_2%A_83_247# 1 2 3 4 13 15 18 20 23 25 27 28 32
+ 33 34 36 37 38 43 44 47
c128 23 0 1.07216e-19 $X=0.58 $Y=1.4
r129 47 49 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=3.51 $Y=2.795
+ $X2=3.51 $Y2=2.99
r130 43 44 9.77977 $w=1.88e-07 $l=1.65e-07 $layer=LI1_cond $X=3.365 $Y=0.35
+ $X2=3.2 $Y2=0.35
r131 37 49 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.345 $Y=2.99
+ $X2=3.51 $Y2=2.99
r132 37 38 128.524 $w=1.68e-07 $l=1.97e-06 $layer=LI1_cond $X=3.345 $Y=2.99
+ $X2=1.375 $Y2=2.99
r133 36 44 121.021 $w=1.68e-07 $l=1.855e-06 $layer=LI1_cond $X=1.345 $Y=0.34
+ $X2=3.2 $Y2=0.34
r134 34 38 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=1.235 $Y=2.905
+ $X2=1.375 $Y2=2.99
r135 33 41 2.78046 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.235 $Y=2.12
+ $X2=1.235 $Y2=2.035
r136 33 34 32.3096 $w=2.78e-07 $l=7.85e-07 $layer=LI1_cond $X=1.235 $Y=2.12
+ $X2=1.235 $Y2=2.905
r137 30 32 22.3574 $w=2.48e-07 $l=4.85e-07 $layer=LI1_cond $X=1.22 $Y=1.035
+ $X2=1.22 $Y2=0.55
r138 29 36 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.22 $Y=0.425
+ $X2=1.345 $Y2=0.34
r139 29 32 5.76222 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=1.22 $Y=0.425
+ $X2=1.22 $Y2=0.55
r140 27 41 4.57959 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=1.095 $Y=2.035
+ $X2=1.235 $Y2=2.035
r141 27 28 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.095 $Y=2.035
+ $X2=0.745 $Y2=2.035
r142 26 39 1.68994 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.745 $Y=1.12
+ $X2=0.62 $Y2=1.12
r143 25 30 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.095 $Y=1.12
+ $X2=1.22 $Y2=1.035
r144 25 26 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.095 $Y=1.12
+ $X2=0.745 $Y2=1.12
r145 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.58
+ $Y=1.4 $X2=0.58 $Y2=1.4
r146 21 28 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.62 $Y=1.95
+ $X2=0.745 $Y2=2.035
r147 21 23 25.3537 $w=2.48e-07 $l=5.5e-07 $layer=LI1_cond $X=0.62 $Y=1.95
+ $X2=0.62 $Y2=1.4
r148 20 39 12.2351 $w=2.5e-07 $l=2.4e-07 $layer=LI1_cond $X=0.62 $Y=1.36
+ $X2=0.62 $Y2=1.12
r149 20 23 1.84391 $w=2.48e-07 $l=4e-08 $layer=LI1_cond $X=0.62 $Y=1.36 $X2=0.62
+ $Y2=1.4
r150 16 24 38.9235 $w=2.69e-07 $l=1.86145e-07 $layer=POLY_cond $X=0.535 $Y=1.235
+ $X2=0.58 $Y2=1.4
r151 16 18 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=0.535 $Y=1.235
+ $X2=0.535 $Y2=0.725
r152 13 24 79.2394 $w=2.69e-07 $l=4.25852e-07 $layer=POLY_cond $X=0.505 $Y=1.79
+ $X2=0.58 $Y2=1.4
r153 13 15 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.505 $Y=1.79
+ $X2=0.505 $Y2=2.365
r154 4 47 600 $w=1.7e-07 $l=1.03865e-06 $layer=licon1_PDIFF $count=1 $X=3.28
+ $Y=1.865 $X2=3.51 $Y2=2.795
r155 3 41 300 $w=1.7e-07 $l=3.20156e-07 $layer=licon1_PDIFF $count=2 $X=1.12
+ $Y=1.865 $X2=1.28 $Y2=2.115
r156 2 43 182 $w=1.7e-07 $l=3.58504e-07 $layer=licon1_NDIFF $count=1 $X=3.145
+ $Y=0.625 $X2=3.365 $Y2=0.36
r157 1 32 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.12
+ $Y=0.405 $X2=1.26 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_LS__XNOR3_2%A 3 5 7 8 12
c42 5 0 2.23227e-19 $X=1.045 $Y=1.79
c43 3 0 2.53685e-19 $X=1.045 $Y=0.725
r44 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.12
+ $Y=1.54 $X2=1.12 $Y2=1.54
r45 8 12 4.00154 $w=3.58e-07 $l=1.25e-07 $layer=LI1_cond $X=1.135 $Y=1.665
+ $X2=1.135 $Y2=1.54
r46 5 11 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=1.045 $Y=1.79
+ $X2=1.12 $Y2=1.54
r47 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.045 $Y=1.79
+ $X2=1.045 $Y2=2.365
r48 1 11 38.5562 $w=2.99e-07 $l=1.98997e-07 $layer=POLY_cond $X=1.045 $Y=1.375
+ $X2=1.12 $Y2=1.54
r49 1 3 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=1.045 $Y=1.375
+ $X2=1.045 $Y2=0.725
.ends

.subckt PM_SKY130_FD_SC_LS__XNOR3_2%A_397_21# 1 2 10 11 12 13 15 16 17 21 22 24
+ 32 33 35 37 39 42 44
c121 42 0 1.16185e-19 $X=3.32 $Y=1.54
c122 22 0 3.85518e-19 $X=3.205 $Y=1.79
c123 11 0 1.69141e-19 $X=2.195 $Y=1.49
c124 10 0 6.5827e-20 $X=2.06 $Y=1.055
r125 42 45 8.69073 $w=4.08e-07 $l=1.65e-07 $layer=LI1_cond $X=3.36 $Y=1.54
+ $X2=3.36 $Y2=1.705
r126 42 44 8.69073 $w=4.08e-07 $l=1.65e-07 $layer=LI1_cond $X=3.36 $Y=1.54
+ $X2=3.36 $Y2=1.375
r127 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.32
+ $Y=1.54 $X2=3.32 $Y2=1.54
r128 37 39 24.2013 $w=2.48e-07 $l=5.25e-07 $layer=LI1_cond $X=3.565 $Y=2.075
+ $X2=4.09 $Y2=2.075
r129 33 35 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=3.565 $Y=1.04
+ $X2=3.925 $Y2=1.04
r130 32 37 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.48 $Y=1.95
+ $X2=3.565 $Y2=2.075
r131 32 45 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=3.48 $Y=1.95
+ $X2=3.48 $Y2=1.705
r132 29 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.48 $Y=1.125
+ $X2=3.565 $Y2=1.04
r133 29 44 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.48 $Y=1.125
+ $X2=3.48 $Y2=1.375
r134 22 43 49.7466 $w=4.26e-07 $l=2.66927e-07 $layer=POLY_cond $X=3.205 $Y=1.79
+ $X2=3.24 $Y2=1.54
r135 22 24 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=3.205 $Y=1.79
+ $X2=3.205 $Y2=2.285
r136 19 43 40.1292 $w=4.26e-07 $l=2.38642e-07 $layer=POLY_cond $X=3.07 $Y=1.375
+ $X2=3.24 $Y2=1.54
r137 19 21 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.07 $Y=1.375
+ $X2=3.07 $Y2=0.945
r138 18 21 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.07 $Y=0.255
+ $X2=3.07 $Y2=0.945
r139 16 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.995 $Y=0.18
+ $X2=3.07 $Y2=0.255
r140 16 17 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=2.995 $Y=0.18
+ $X2=2.135 $Y2=0.18
r141 13 15 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.195 $Y=1.79
+ $X2=2.195 $Y2=2.185
r142 12 13 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.195 $Y=1.7
+ $X2=2.195 $Y2=1.79
r143 11 25 69.2234 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.195 $Y=1.415
+ $X2=2.06 $Y2=1.415
r144 11 12 81.629 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=2.195 $Y=1.49
+ $X2=2.195 $Y2=1.7
r145 8 25 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.06 $Y=1.34
+ $X2=2.06 $Y2=1.415
r146 8 10 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.06 $Y=1.34
+ $X2=2.06 $Y2=1.055
r147 7 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.06 $Y=0.255
+ $X2=2.135 $Y2=0.18
r148 7 10 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=2.06 $Y=0.255 $X2=2.06
+ $Y2=1.055
r149 2 39 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=3.95
+ $Y=1.84 $X2=4.09 $Y2=2.115
r150 1 35 182 $w=1.7e-07 $l=6.63551e-07 $layer=licon1_NDIFF $count=1 $X=3.78
+ $Y=0.445 $X2=3.925 $Y2=1.04
.ends

.subckt PM_SKY130_FD_SC_LS__XNOR3_2%B 3 5 6 7 10 11 12 13 15 17 18 22 23 26 29
+ 31 33 35 36 41 42
c137 15 0 1.16185e-19 $X=2.57 $Y=0.945
c138 13 0 2.64147e-20 $X=2.57 $Y=1.505
c139 3 0 2.86506e-20 $X=1.57 $Y=0.725
r140 41 43 10.2699 $w=3.52e-07 $l=7.5e-08 $layer=POLY_cond $X=4.24 $Y=1.557
+ $X2=4.315 $Y2=1.557
r141 41 42 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.24
+ $Y=1.515 $X2=4.24 $Y2=1.515
r142 39 41 13.6932 $w=3.52e-07 $l=1e-07 $layer=POLY_cond $X=4.14 $Y=1.557
+ $X2=4.24 $Y2=1.557
r143 36 42 2.67779 $w=6.68e-07 $l=1.5e-07 $layer=LI1_cond $X=4.07 $Y=1.665
+ $X2=4.07 $Y2=1.515
r144 31 43 22.7654 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=4.315 $Y=1.765
+ $X2=4.315 $Y2=1.557
r145 31 33 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.315 $Y=1.765
+ $X2=4.315 $Y2=2.4
r146 27 39 22.7654 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.14 $Y=1.35
+ $X2=4.14 $Y2=1.557
r147 27 29 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=4.14 $Y=1.35
+ $X2=4.14 $Y2=0.815
r148 25 39 46.5568 $w=3.52e-07 $l=3.4e-07 $layer=POLY_cond $X=3.8 $Y=1.557
+ $X2=4.14 $Y2=1.557
r149 25 26 715.309 $w=1.5e-07 $l=1.395e-06 $layer=POLY_cond $X=3.8 $Y=1.68
+ $X2=3.8 $Y2=3.075
r150 24 35 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.755 $Y=3.15
+ $X2=2.665 $Y2=3.15
r151 23 26 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.725 $Y=3.15
+ $X2=3.8 $Y2=3.075
r152 23 24 497.383 $w=1.5e-07 $l=9.7e-07 $layer=POLY_cond $X=3.725 $Y=3.15
+ $X2=2.755 $Y2=3.15
r153 20 22 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.665 $Y=2.58
+ $X2=2.665 $Y2=2.185
r154 19 22 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.665 $Y=1.79
+ $X2=2.665 $Y2=2.185
r155 18 35 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=2.665 $Y=3.075
+ $X2=2.665 $Y2=3.15
r156 17 20 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.665 $Y=2.67
+ $X2=2.665 $Y2=2.58
r157 17 18 157.427 $w=1.8e-07 $l=4.05e-07 $layer=POLY_cond $X=2.665 $Y=2.67
+ $X2=2.665 $Y2=3.075
r158 13 19 61.8784 $w=2.22e-07 $l=3.2909e-07 $layer=POLY_cond $X=2.57 $Y=1.505
+ $X2=2.665 $Y2=1.79
r159 13 15 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.57 $Y=1.505
+ $X2=2.57 $Y2=0.945
r160 11 35 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.575 $Y=3.15
+ $X2=2.665 $Y2=3.15
r161 11 12 461.489 $w=1.5e-07 $l=9e-07 $layer=POLY_cond $X=2.575 $Y=3.15
+ $X2=1.675 $Y2=3.15
r162 8 10 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.585 $Y=2.78
+ $X2=1.585 $Y2=2.285
r163 7 34 110.782 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=1.585 $Y=1.79
+ $X2=1.585 $Y2=1.505
r164 7 10 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.585 $Y=1.79
+ $X2=1.585 $Y2=2.285
r165 6 12 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=1.585 $Y=3.075
+ $X2=1.675 $Y2=3.15
r166 5 8 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.585 $Y=2.87 $X2=1.585
+ $Y2=2.78
r167 5 6 79.6855 $w=1.8e-07 $l=2.05e-07 $layer=POLY_cond $X=1.585 $Y=2.87
+ $X2=1.585 $Y2=3.075
r168 3 34 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=1.57 $Y=0.725
+ $X2=1.57 $Y2=1.505
.ends

.subckt PM_SKY130_FD_SC_LS__XNOR3_2%A_1027_48# 1 2 9 11 13 14 20 23 27 30 31
r76 27 29 3.21434 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=6.555 $Y=1.085
+ $X2=6.555 $Y2=1.17
r77 23 31 9.06106 $w=3.63e-07 $l=1.82e-07 $layer=LI1_cond $X=6.687 $Y=2.132
+ $X2=6.687 $Y2=1.95
r78 23 25 3.10849 $w=3.65e-07 $l=9.3e-08 $layer=LI1_cond $X=6.687 $Y=2.132
+ $X2=6.687 $Y2=2.225
r79 21 30 6.95506 $w=2.27e-07 $l=1.9182e-07 $layer=LI1_cond $X=6.59 $Y=1.805
+ $X2=6.532 $Y2=1.64
r80 21 31 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=6.59 $Y=1.805
+ $X2=6.59 $Y2=1.95
r81 20 30 6.95506 $w=2.27e-07 $l=1.65e-07 $layer=LI1_cond $X=6.532 $Y=1.475
+ $X2=6.532 $Y2=1.64
r82 20 29 12.3332 $w=2.83e-07 $l=3.05e-07 $layer=LI1_cond $X=6.532 $Y=1.475
+ $X2=6.532 $Y2=1.17
r83 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.49
+ $Y=1.64 $X2=5.49 $Y2=1.64
r84 14 30 0.0443336 $w=3.3e-07 $l=1.42e-07 $layer=LI1_cond $X=6.39 $Y=1.64
+ $X2=6.532 $Y2=1.64
r85 14 16 31.4303 $w=3.28e-07 $l=9e-07 $layer=LI1_cond $X=6.39 $Y=1.64 $X2=5.49
+ $Y2=1.64
r86 11 17 53.0942 $w=4.32e-07 $l=2.8e-07 $layer=POLY_cond $X=5.395 $Y=1.92
+ $X2=5.395 $Y2=1.64
r87 11 13 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=5.395 $Y=1.92
+ $X2=5.395 $Y2=2.415
r88 7 17 40.2632 $w=4.32e-07 $l=2.5446e-07 $layer=POLY_cond $X=5.21 $Y=1.475
+ $X2=5.395 $Y2=1.64
r89 7 9 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=5.21 $Y=1.475
+ $X2=5.21 $Y2=0.69
r90 2 25 600 $w=1.7e-07 $l=4.49583e-07 $layer=licon1_PDIFF $count=1 $X=6.645
+ $Y=1.84 $X2=6.785 $Y2=2.225
r91 1 27 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=6.41
+ $Y=0.81 $X2=6.555 $Y2=1.085
.ends

.subckt PM_SKY130_FD_SC_LS__XNOR3_2%C 1 3 4 5 6 7 8 10 11 13 15 16 18 21 26
c83 16 0 1.73622e-19 $X=7.01 $Y=1.765
c84 13 0 1.44369e-19 $X=6.77 $Y=1.35
c85 1 0 1.52403e-19 $X=5.71 $Y=1.085
r86 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.01
+ $Y=1.515 $X2=7.01 $Y2=1.515
r87 23 25 10.378 $w=4.18e-07 $l=9e-08 $layer=POLY_cond $X=6.935 $Y=1.425
+ $X2=6.935 $Y2=1.515
r88 21 26 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=7.01 $Y=1.665
+ $X2=7.01 $Y2=1.515
r89 16 25 49.7565 $w=4.18e-07 $l=2.85044e-07 $layer=POLY_cond $X=7.01 $Y=1.765
+ $X2=6.935 $Y2=1.515
r90 16 18 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=7.01 $Y=1.765
+ $X2=7.01 $Y2=2.16
r91 13 23 29.5771 $w=4.18e-07 $l=1.98997e-07 $layer=POLY_cond $X=6.77 $Y=1.35
+ $X2=6.935 $Y2=1.425
r92 13 15 106.04 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=6.77 $Y=1.35 $X2=6.77
+ $Y2=1.02
r93 12 20 3.61756 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=6.1 $Y=1.425 $X2=6.01
+ $Y2=1.425
r94 11 23 26.9416 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=6.695 $Y=1.425
+ $X2=6.935 $Y2=1.425
r95 11 12 305.096 $w=1.5e-07 $l=5.95e-07 $layer=POLY_cond $X=6.695 $Y=1.425
+ $X2=6.1 $Y2=1.425
r96 8 10 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=6.01 $Y=1.92 $X2=6.01
+ $Y2=2.415
r97 7 8 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.01 $Y=1.83 $X2=6.01
+ $Y2=1.92
r98 6 20 45.2467 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.01 $Y=1.59
+ $X2=6.01 $Y2=1.425
r99 6 7 93.2903 $w=1.8e-07 $l=2.4e-07 $layer=POLY_cond $X=6.01 $Y=1.59 $X2=6.01
+ $Y2=1.83
r100 4 20 82.4064 $w=1.55e-07 $l=2.65e-07 $layer=POLY_cond $X=6.01 $Y=1.16
+ $X2=6.01 $Y2=1.425
r101 4 5 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.95 $Y=1.16
+ $X2=5.785 $Y2=1.16
r102 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.71 $Y=1.085
+ $X2=5.785 $Y2=1.16
r103 1 3 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=5.71 $Y=1.085
+ $X2=5.71 $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_LS__XNOR3_2%A_1057_74# 1 2 7 9 10 12 13 15 16 18 21 23
+ 24 25 28 29 30 32 34 35 36 37 38 42 44 49 51 56
c122 56 0 1.44369e-19 $X=8.14 $Y=1.552
c123 49 0 1.38659e-19 $X=7.59 $Y=1.505
c124 7 0 1.92468e-19 $X=7.69 $Y=1.765
r125 56 57 0.68661 $w=3.51e-07 $l=5e-09 $layer=POLY_cond $X=8.14 $Y=1.552
+ $X2=8.145 $Y2=1.552
r126 55 56 58.3618 $w=3.51e-07 $l=4.25e-07 $layer=POLY_cond $X=7.715 $Y=1.552
+ $X2=8.14 $Y2=1.552
r127 54 55 3.43305 $w=3.51e-07 $l=2.5e-08 $layer=POLY_cond $X=7.69 $Y=1.552
+ $X2=7.715 $Y2=1.552
r128 50 54 13.7322 $w=3.51e-07 $l=1e-07 $layer=POLY_cond $X=7.59 $Y=1.552
+ $X2=7.69 $Y2=1.552
r129 49 52 8.4794 $w=3.43e-07 $l=1.65e-07 $layer=LI1_cond $X=7.582 $Y=1.505
+ $X2=7.582 $Y2=1.67
r130 49 51 8.4794 $w=3.43e-07 $l=1.65e-07 $layer=LI1_cond $X=7.582 $Y=1.505
+ $X2=7.582 $Y2=1.34
r131 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.59
+ $Y=1.505 $X2=7.59 $Y2=1.505
r132 44 46 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=5.7 $Y=2.82 $X2=5.7
+ $Y2=2.99
r133 42 52 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=7.495 $Y=1.95
+ $X2=7.495 $Y2=1.67
r134 39 51 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=7.495 $Y=1.18
+ $X2=7.495 $Y2=1.34
r135 37 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.41 $Y=2.035
+ $X2=7.495 $Y2=1.95
r136 37 38 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=7.41 $Y=2.035
+ $X2=7.21 $Y2=2.035
r137 35 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.41 $Y=1.095
+ $X2=7.495 $Y2=1.18
r138 35 36 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=7.41 $Y=1.095
+ $X2=7.06 $Y2=1.095
r139 33 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.125 $Y=2.12
+ $X2=7.21 $Y2=2.035
r140 33 34 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=7.125 $Y=2.12
+ $X2=7.125 $Y2=2.905
r141 32 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.975 $Y=1.01
+ $X2=7.06 $Y2=1.095
r142 31 32 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=6.975 $Y=0.83
+ $X2=6.975 $Y2=1.01
r143 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.89 $Y=0.745
+ $X2=6.975 $Y2=0.83
r144 29 30 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=6.89 $Y=0.745
+ $X2=6.5 $Y2=0.745
r145 28 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.415 $Y=0.66
+ $X2=6.5 $Y2=0.745
r146 27 28 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=6.415 $Y=0.425
+ $X2=6.415 $Y2=0.66
r147 26 46 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.865 $Y=2.99
+ $X2=5.7 $Y2=2.99
r148 25 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.04 $Y=2.99
+ $X2=7.125 $Y2=2.905
r149 25 26 76.6578 $w=1.68e-07 $l=1.175e-06 $layer=LI1_cond $X=7.04 $Y=2.99
+ $X2=5.865 $Y2=2.99
r150 23 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.33 $Y=0.34
+ $X2=6.415 $Y2=0.425
r151 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.33 $Y=0.34
+ $X2=5.66 $Y2=0.34
r152 19 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.495 $Y=0.425
+ $X2=5.66 $Y2=0.34
r153 19 21 2.44458 $w=3.28e-07 $l=7e-08 $layer=LI1_cond $X=5.495 $Y=0.425
+ $X2=5.495 $Y2=0.495
r154 16 57 22.6971 $w=1.5e-07 $l=2.12e-07 $layer=POLY_cond $X=8.145 $Y=1.34
+ $X2=8.145 $Y2=1.552
r155 16 18 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=8.145 $Y=1.34
+ $X2=8.145 $Y2=0.86
r156 13 56 22.6971 $w=1.5e-07 $l=2.13e-07 $layer=POLY_cond $X=8.14 $Y=1.765
+ $X2=8.14 $Y2=1.552
r157 13 15 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.14 $Y=1.765
+ $X2=8.14 $Y2=2.4
r158 10 55 22.6971 $w=1.5e-07 $l=2.12e-07 $layer=POLY_cond $X=7.715 $Y=1.34
+ $X2=7.715 $Y2=1.552
r159 10 12 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=7.715 $Y=1.34
+ $X2=7.715 $Y2=0.86
r160 7 54 22.6971 $w=1.5e-07 $l=2.13e-07 $layer=POLY_cond $X=7.69 $Y=1.765
+ $X2=7.69 $Y2=1.552
r161 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.69 $Y=1.765
+ $X2=7.69 $Y2=2.4
r162 2 44 600 $w=1.7e-07 $l=9.32939e-07 $layer=licon1_PDIFF $count=1 $X=5.47
+ $Y=1.995 $X2=5.7 $Y2=2.82
r163 1 21 91 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=2 $X=5.285
+ $Y=0.37 $X2=5.495 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LS__XNOR3_2%A_27_373# 1 2 3 4 15 19 20 21 23 24 27 30 33
+ 36 40 41 44 47
c105 47 0 1.46469e-19 $X=1.68 $Y=1.295
c106 40 0 2.76385e-20 $X=1.535 $Y=1.295
c107 36 0 1.9829e-20 $X=2.275 $Y=1.11
c108 33 0 1.86262e-19 $X=0.28 $Y=2.375
c109 27 0 1.90902e-19 $X=2.44 $Y=2.01
c110 19 0 9.32687e-21 $X=1.63 $Y=1.38
r111 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=1.295
+ $X2=1.68 $Y2=1.295
r112 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=1.295
+ $X2=0.24 $Y2=1.295
r113 41 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.385 $Y=1.295
+ $X2=0.24 $Y2=1.295
r114 40 47 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.535 $Y=1.295
+ $X2=1.68 $Y2=1.295
r115 40 41 1.42326 $w=1.4e-07 $l=1.15e-06 $layer=MET1_cond $X=1.535 $Y=1.295
+ $X2=0.385 $Y2=1.295
r116 36 38 7.46783 $w=2.48e-07 $l=1.62e-07 $layer=LI1_cond $X=2.26 $Y=1.11
+ $X2=2.26 $Y2=1.272
r117 34 44 47.7784 $w=2.38e-07 $l=9.95e-07 $layer=LI1_cond $X=0.205 $Y=2.29
+ $X2=0.205 $Y2=1.295
r118 33 34 4.00454 $w=3.58e-07 $l=8.5e-08 $layer=LI1_cond $X=0.265 $Y=2.375
+ $X2=0.265 $Y2=2.29
r119 30 44 11.0442 $w=2.38e-07 $l=2.3e-07 $layer=LI1_cond $X=0.205 $Y=1.065
+ $X2=0.205 $Y2=1.295
r120 25 27 19.382 $w=3.28e-07 $l=5.55e-07 $layer=LI1_cond $X=2.44 $Y=2.565
+ $X2=2.44 $Y2=2.01
r121 23 25 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.275 $Y=2.65
+ $X2=2.44 $Y2=2.565
r122 23 24 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=2.275 $Y=2.65
+ $X2=1.715 $Y2=2.65
r123 22 48 3.05574 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=1.715 $Y=1.272
+ $X2=1.63 $Y2=1.272
r124 21 38 1.64524 $w=2.15e-07 $l=1.25e-07 $layer=LI1_cond $X=2.135 $Y=1.272
+ $X2=2.26 $Y2=1.272
r125 21 22 22.5128 $w=2.13e-07 $l=4.2e-07 $layer=LI1_cond $X=2.135 $Y=1.272
+ $X2=1.715 $Y2=1.272
r126 20 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.63 $Y=2.565
+ $X2=1.715 $Y2=2.65
r127 19 48 3.88258 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=1.63 $Y=1.38
+ $X2=1.63 $Y2=1.272
r128 19 20 77.3102 $w=1.68e-07 $l=1.185e-06 $layer=LI1_cond $X=1.63 $Y=1.38
+ $X2=1.63 $Y2=2.565
r129 13 30 6.50835 $w=3.18e-07 $l=1.6e-07 $layer=LI1_cond $X=0.245 $Y=0.905
+ $X2=0.245 $Y2=1.065
r130 13 15 12.7849 $w=3.18e-07 $l=3.55e-07 $layer=LI1_cond $X=0.245 $Y=0.905
+ $X2=0.245 $Y2=0.55
r131 4 27 300 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_PDIFF $count=2 $X=2.27
+ $Y=1.865 $X2=2.44 $Y2=2.01
r132 3 33 300 $w=1.7e-07 $l=5.77971e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.865 $X2=0.28 $Y2=2.375
r133 2 36 182 $w=1.7e-07 $l=3.27605e-07 $layer=licon1_NDIFF $count=1 $X=2.135
+ $Y=0.845 $X2=2.275 $Y2=1.11
r134 1 15 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.175
+ $Y=0.405 $X2=0.32 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_LS__XNOR3_2%VPWR 1 2 3 4 17 21 25 27 29 33 35 43 48 54
+ 57 60 64
c83 43 0 1.73622e-19 $X=7.38 $Y=3.33
c84 2 0 3.71954e-20 $X=4.39 $Y=1.84
r85 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33 $X2=8.4
+ $Y2=3.33
r86 60 61 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r87 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r88 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r89 52 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r90 52 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=7.44 $Y2=3.33
r91 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r92 49 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.55 $Y=3.33
+ $X2=7.465 $Y2=3.33
r93 49 51 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=7.55 $Y=3.33 $X2=7.92
+ $Y2=3.33
r94 48 63 4.01803 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=8.28 $Y=3.33 $X2=8.46
+ $Y2=3.33
r95 48 51 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=8.28 $Y=3.33
+ $X2=7.92 $Y2=3.33
r96 47 61 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=7.44 $Y2=3.33
r97 47 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r98 46 47 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r99 44 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.785 $Y=3.33
+ $X2=4.62 $Y2=3.33
r100 44 46 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=4.785 $Y=3.33
+ $X2=5.04 $Y2=3.33
r101 43 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.38 $Y=3.33
+ $X2=7.465 $Y2=3.33
r102 43 46 152.663 $w=1.68e-07 $l=2.34e-06 $layer=LI1_cond $X=7.38 $Y=3.33
+ $X2=5.04 $Y2=3.33
r103 41 42 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r104 39 42 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=4.08 $Y2=3.33
r105 39 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r106 38 41 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=4.08 $Y2=3.33
r107 38 39 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r108 36 54 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=0.925 $Y=3.33
+ $X2=0.785 $Y2=3.33
r109 36 38 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.925 $Y=3.33
+ $X2=1.2 $Y2=3.33
r110 35 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.455 $Y=3.33
+ $X2=4.62 $Y2=3.33
r111 35 41 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=4.455 $Y=3.33
+ $X2=4.08 $Y2=3.33
r112 33 58 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=3.33
+ $X2=4.56 $Y2=3.33
r113 33 42 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=3.33
+ $X2=4.08 $Y2=3.33
r114 29 32 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=8.405 $Y=1.985
+ $X2=8.405 $Y2=2.815
r115 27 63 3.12513 $w=2.5e-07 $l=1.09087e-07 $layer=LI1_cond $X=8.405 $Y=3.245
+ $X2=8.46 $Y2=3.33
r116 27 32 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=8.405 $Y=3.245
+ $X2=8.405 $Y2=2.815
r117 23 60 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.465 $Y=3.245
+ $X2=7.465 $Y2=3.33
r118 23 25 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=7.465 $Y=3.245
+ $X2=7.465 $Y2=2.455
r119 19 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.62 $Y=3.245
+ $X2=4.62 $Y2=3.33
r120 19 21 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=4.62 $Y=3.245
+ $X2=4.62 $Y2=2.9
r121 15 54 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.785 $Y=3.245
+ $X2=0.785 $Y2=3.33
r122 15 17 29.84 $w=2.78e-07 $l=7.25e-07 $layer=LI1_cond $X=0.785 $Y=3.245
+ $X2=0.785 $Y2=2.52
r123 4 32 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=8.215
+ $Y=1.84 $X2=8.365 $Y2=2.815
r124 4 29 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=8.215
+ $Y=1.84 $X2=8.365 $Y2=1.985
r125 3 25 300 $w=1.7e-07 $l=7.82256e-07 $layer=licon1_PDIFF $count=2 $X=7.085
+ $Y=1.84 $X2=7.465 $Y2=2.455
r126 2 21 600 $w=1.7e-07 $l=1.16936e-06 $layer=licon1_PDIFF $count=1 $X=4.39
+ $Y=1.84 $X2=4.62 $Y2=2.9
r127 1 17 600 $w=1.7e-07 $l=7.32871e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.865 $X2=0.745 $Y2=2.52
.ends

.subckt PM_SKY130_FD_SC_LS__XNOR3_2%A_332_373# 1 2 3 4 15 17 18 19 20 21 25 31
+ 37 39 40 43 46
c111 43 0 1.94615e-19 $X=2.64 $Y=1.295
c112 40 0 1.95555e-19 $X=2.785 $Y=1.295
r113 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=1.295
+ $X2=5.04 $Y2=1.295
r114 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=1.295
+ $X2=2.64 $Y2=1.295
r115 40 42 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.785 $Y=1.295
+ $X2=2.64 $Y2=1.295
r116 39 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.895 $Y=1.295
+ $X2=5.04 $Y2=1.295
r117 39 40 2.61138 $w=1.4e-07 $l=2.11e-06 $layer=MET1_cond $X=4.895 $Y=1.295
+ $X2=2.785 $Y2=1.295
r118 34 37 5.9927 $w=2.48e-07 $l=1.3e-07 $layer=LI1_cond $X=5.04 $Y=2.1 $X2=5.17
+ $Y2=2.1
r119 33 43 14.1409 $w=1.98e-07 $l=2.55e-07 $layer=LI1_cond $X=2.655 $Y=1.55
+ $X2=2.655 $Y2=1.295
r120 28 43 0.554545 $w=1.98e-07 $l=1e-08 $layer=LI1_cond $X=2.655 $Y=1.285
+ $X2=2.655 $Y2=1.295
r121 27 31 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=2.655 $Y=1.12
+ $X2=2.8 $Y2=1.12
r122 27 28 3.66692 $w=2e-07 $l=1.65e-07 $layer=LI1_cond $X=2.655 $Y=1.12
+ $X2=2.655 $Y2=1.285
r123 23 25 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=5.995 $Y=1.135
+ $X2=5.995 $Y2=0.81
r124 22 47 4.03528 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=5.155 $Y=1.22
+ $X2=5.04 $Y2=1.22
r125 21 23 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.83 $Y=1.22
+ $X2=5.995 $Y2=1.135
r126 21 22 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=5.83 $Y=1.22
+ $X2=5.155 $Y2=1.22
r127 20 34 1.2199 $w=2.3e-07 $l=1.25e-07 $layer=LI1_cond $X=5.04 $Y=1.975
+ $X2=5.04 $Y2=2.1
r128 19 47 2.9826 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.04 $Y=1.305
+ $X2=5.04 $Y2=1.22
r129 19 20 33.5712 $w=2.28e-07 $l=6.7e-07 $layer=LI1_cond $X=5.04 $Y=1.305
+ $X2=5.04 $Y2=1.975
r130 17 33 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=2.555 $Y=1.635
+ $X2=2.655 $Y2=1.55
r131 17 18 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=2.555 $Y=1.635
+ $X2=2.105 $Y2=1.635
r132 13 18 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=1.995 $Y=1.72
+ $X2=2.105 $Y2=1.635
r133 13 15 20.9535 $w=2.18e-07 $l=4e-07 $layer=LI1_cond $X=1.995 $Y=1.72
+ $X2=1.995 $Y2=2.12
r134 4 37 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=5.03
+ $Y=1.995 $X2=5.17 $Y2=2.14
r135 3 15 600 $w=1.7e-07 $l=4.18509e-07 $layer=licon1_PDIFF $count=1 $X=1.66
+ $Y=1.865 $X2=1.97 $Y2=2.12
r136 2 25 182 $w=1.7e-07 $l=5.3479e-07 $layer=licon1_NDIFF $count=1 $X=5.785
+ $Y=0.37 $X2=5.995 $Y2=0.81
r137 1 31 182 $w=1.7e-07 $l=5.6723e-07 $layer=licon1_NDIFF $count=1 $X=2.645
+ $Y=0.625 $X2=2.8 $Y2=1.12
.ends

.subckt PM_SKY130_FD_SC_LS__XNOR3_2%A_329_81# 1 2 3 4 15 19 21 22 23 24 25 29 31
+ 36 37 41
c127 37 0 6.5827e-20 $X=2.725 $Y=0.69
c128 36 0 8.82162e-21 $X=2.555 $Y=0.69
c129 25 0 3.71954e-20 $X=6.07 $Y=2.48
c130 23 0 1.52403e-19 $X=4.67 $Y=0.965
r131 39 40 4.81237 $w=4.69e-07 $l=1.85e-07 $layer=LI1_cond $X=4.872 $Y=0.515
+ $X2=4.872 $Y2=0.7
r132 36 37 9.92344 $w=1.88e-07 $l=1.7e-07 $layer=LI1_cond $X=2.555 $Y=0.69
+ $X2=2.725 $Y2=0.69
r133 31 34 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=1.79 $Y=0.68
+ $X2=1.79 $Y2=0.8
r134 27 29 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=6.195 $Y=2.395
+ $X2=6.195 $Y2=2.14
r135 26 41 5.16603 $w=1.7e-07 $l=9.12688e-08 $layer=LI1_cond $X=4.755 $Y=2.48
+ $X2=4.67 $Y2=2.467
r136 25 27 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.07 $Y=2.48
+ $X2=6.195 $Y2=2.395
r137 25 26 85.7914 $w=1.68e-07 $l=1.315e-06 $layer=LI1_cond $X=6.07 $Y=2.48
+ $X2=4.755 $Y2=2.48
r138 24 41 1.34256 $w=1.7e-07 $l=9.7e-08 $layer=LI1_cond $X=4.67 $Y=2.37
+ $X2=4.67 $Y2=2.467
r139 23 40 12.1197 $w=4.69e-07 $l=3.51788e-07 $layer=LI1_cond $X=4.67 $Y=0.965
+ $X2=4.872 $Y2=0.7
r140 23 24 91.6631 $w=1.68e-07 $l=1.405e-06 $layer=LI1_cond $X=4.67 $Y=0.965
+ $X2=4.67 $Y2=2.37
r141 21 41 5.16603 $w=1.7e-07 $l=9.0802e-08 $layer=LI1_cond $X=4.585 $Y=2.455
+ $X2=4.67 $Y2=2.467
r142 21 22 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=4.585 $Y=2.455
+ $X2=3.145 $Y2=2.455
r143 17 22 10.2712 $w=1.77e-07 $l=1.92873e-07 $layer=LI1_cond $X=2.99 $Y=2.37
+ $X2=3.145 $Y2=2.455
r144 17 19 12.2679 $w=3.08e-07 $l=3.3e-07 $layer=LI1_cond $X=2.99 $Y=2.37
+ $X2=2.99 $Y2=2.04
r145 15 40 6.75673 $w=1.7e-07 $l=2.87e-07 $layer=LI1_cond $X=4.585 $Y=0.7
+ $X2=4.872 $Y2=0.7
r146 15 37 121.348 $w=1.68e-07 $l=1.86e-06 $layer=LI1_cond $X=4.585 $Y=0.7
+ $X2=2.725 $Y2=0.7
r147 14 31 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.955 $Y=0.68
+ $X2=1.79 $Y2=0.68
r148 14 36 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=1.955 $Y=0.68
+ $X2=2.555 $Y2=0.68
r149 4 29 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=6.085
+ $Y=1.995 $X2=6.235 $Y2=2.14
r150 3 19 300 $w=1.7e-07 $l=3.15595e-07 $layer=licon1_PDIFF $count=2 $X=2.74
+ $Y=1.865 $X2=2.98 $Y2=2.04
r151 2 39 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=4.85
+ $Y=0.37 $X2=4.995 $Y2=0.515
r152 1 34 182 $w=1.7e-07 $l=4.59701e-07 $layer=licon1_NDIFF $count=1 $X=1.645
+ $Y=0.405 $X2=1.785 $Y2=0.8
.ends

.subckt PM_SKY130_FD_SC_LS__XNOR3_2%X 1 2 9 14 15 16 17 28
c33 15 0 1.92468e-19 $X=7.922 $Y=1.84
r34 21 28 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=7.93 $Y=1.005 $X2=7.93
+ $Y2=0.925
r35 17 30 8.39233 $w=3.28e-07 $l=1.63e-07 $layer=LI1_cond $X=7.93 $Y=1.007
+ $X2=7.93 $Y2=1.17
r36 17 21 0.069845 $w=3.28e-07 $l=2e-09 $layer=LI1_cond $X=7.93 $Y=1.007
+ $X2=7.93 $Y2=1.005
r37 17 28 0.104768 $w=3.28e-07 $l=3e-09 $layer=LI1_cond $X=7.93 $Y=0.922
+ $X2=7.93 $Y2=0.925
r38 16 17 12.8166 $w=3.28e-07 $l=3.67e-07 $layer=LI1_cond $X=7.93 $Y=0.555
+ $X2=7.93 $Y2=0.922
r39 15 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.01 $Y=1.84
+ $X2=8.01 $Y2=1.17
r40 14 15 8.4794 $w=3.43e-07 $l=1.65e-07 $layer=LI1_cond $X=7.922 $Y=2.005
+ $X2=7.922 $Y2=1.84
r41 7 14 0.233829 $w=3.43e-07 $l=7e-09 $layer=LI1_cond $X=7.922 $Y=2.012
+ $X2=7.922 $Y2=2.005
r42 7 9 26.8235 $w=3.43e-07 $l=8.03e-07 $layer=LI1_cond $X=7.922 $Y=2.012
+ $X2=7.922 $Y2=2.815
r43 2 14 400 $w=1.7e-07 $l=2.2798e-07 $layer=licon1_PDIFF $count=1 $X=7.765
+ $Y=1.84 $X2=7.915 $Y2=2.005
r44 2 9 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=7.765
+ $Y=1.84 $X2=7.915 $Y2=2.815
r45 1 16 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.79
+ $Y=0.49 $X2=7.93 $Y2=0.635
.ends

.subckt PM_SKY130_FD_SC_LS__XNOR3_2%VGND 1 2 3 4 15 19 21 23 25 27 29 34 42 48
+ 51 54 62
c82 54 0 1.38659e-19 $X=6.96 $Y=0
r83 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r84 55 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r85 54 59 7.08036 $w=5.6e-07 $l=3.25e-07 $layer=LI1_cond $X=7.242 $Y=0 $X2=7.242
+ $Y2=0.325
r86 54 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r87 54 55 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r88 52 55 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=4.56 $Y=0 $X2=6.96
+ $Y2=0
r89 51 52 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r90 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r91 46 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.4
+ $Y2=0
r92 46 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=7.44
+ $Y2=0
r93 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r94 43 54 7.87414 $w=1.7e-07 $l=3.43e-07 $layer=LI1_cond $X=7.585 $Y=0 $X2=7.242
+ $Y2=0
r95 43 45 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=7.585 $Y=0 $X2=7.92
+ $Y2=0
r96 42 61 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=8.275 $Y=0 $X2=8.457
+ $Y2=0
r97 42 45 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=8.275 $Y=0 $X2=7.92
+ $Y2=0
r98 40 41 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r99 38 41 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=4.08
+ $Y2=0
r100 38 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r101 37 40 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=4.08
+ $Y2=0
r102 37 38 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=1.2 $Y=0
+ $X2=1.2 $Y2=0
r103 35 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.915 $Y=0 $X2=0.75
+ $Y2=0
r104 35 37 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.915 $Y=0 $X2=1.2
+ $Y2=0
r105 34 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.27 $Y=0 $X2=4.435
+ $Y2=0
r106 34 40 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=4.27 $Y=0 $X2=4.08
+ $Y2=0
r107 32 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r108 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r109 29 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.585 $Y=0 $X2=0.75
+ $Y2=0
r110 29 31 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.585 $Y=0 $X2=0.24
+ $Y2=0
r111 27 52 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=0
+ $X2=4.56 $Y2=0
r112 27 41 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=0
+ $X2=4.08 $Y2=0
r113 23 61 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=8.4 $Y=0.085
+ $X2=8.457 $Y2=0
r114 23 25 25.3537 $w=2.48e-07 $l=5.5e-07 $layer=LI1_cond $X=8.4 $Y=0.085
+ $X2=8.4 $Y2=0.635
r115 22 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.6 $Y=0 $X2=4.435
+ $Y2=0
r116 21 54 7.87414 $w=1.7e-07 $l=3.42e-07 $layer=LI1_cond $X=6.9 $Y=0 $X2=7.242
+ $Y2=0
r117 21 22 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=6.9 $Y=0 $X2=4.6
+ $Y2=0
r118 17 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.435 $Y=0.085
+ $X2=4.435 $Y2=0
r119 17 19 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=4.435 $Y=0.085
+ $X2=4.435 $Y2=0.36
r120 13 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=0.085
+ $X2=0.75 $Y2=0
r121 13 15 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=0.75 $Y=0.085
+ $X2=0.75 $Y2=0.78
r122 4 25 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.22
+ $Y=0.49 $X2=8.36 $Y2=0.635
r123 3 59 60.6667 $w=1.7e-07 $l=7.80705e-07 $layer=licon1_NDIFF $count=3
+ $X=6.845 $Y=0.81 $X2=7.42 $Y2=0.325
r124 2 19 182 $w=1.7e-07 $l=2.59037e-07 $layer=licon1_NDIFF $count=1 $X=4.215
+ $Y=0.445 $X2=4.435 $Y2=0.36
r125 1 15 182 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_NDIFF $count=1 $X=0.61
+ $Y=0.405 $X2=0.75 $Y2=0.78
.ends

