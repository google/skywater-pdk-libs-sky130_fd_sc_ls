* File: sky130_fd_sc_ls__dfstp_2.pxi.spice
* Created: Fri Aug 28 13:15:46 2020
* 
x_PM_SKY130_FD_SC_LS__DFSTP_2%D N_D_c_245_n N_D_c_250_n N_D_M1026_g N_D_c_251_n
+ N_D_M1018_g D D N_D_c_247_n N_D_c_248_n N_D_c_253_n
+ PM_SKY130_FD_SC_LS__DFSTP_2%D
x_PM_SKY130_FD_SC_LS__DFSTP_2%CLK N_CLK_c_279_n N_CLK_M1029_g N_CLK_c_280_n
+ N_CLK_M1028_g CLK PM_SKY130_FD_SC_LS__DFSTP_2%CLK
x_PM_SKY130_FD_SC_LS__DFSTP_2%A_398_74# N_A_398_74#_M1016_d N_A_398_74#_M1007_d
+ N_A_398_74#_c_312_n N_A_398_74#_c_331_n N_A_398_74#_c_332_n
+ N_A_398_74#_M1000_g N_A_398_74#_c_313_n N_A_398_74#_c_314_n
+ N_A_398_74#_M1014_g N_A_398_74#_M1032_g N_A_398_74#_c_335_n
+ N_A_398_74#_M1013_g N_A_398_74#_c_316_n N_A_398_74#_c_428_p
+ N_A_398_74#_c_317_n N_A_398_74#_c_318_n N_A_398_74#_c_336_n
+ N_A_398_74#_c_337_n N_A_398_74#_c_319_n N_A_398_74#_c_320_n
+ N_A_398_74#_c_340_n N_A_398_74#_c_341_n N_A_398_74#_c_342_n
+ N_A_398_74#_c_343_n N_A_398_74#_c_344_n N_A_398_74#_c_345_n
+ N_A_398_74#_c_376_p N_A_398_74#_c_366_p N_A_398_74#_c_321_n
+ N_A_398_74#_c_322_n N_A_398_74#_c_323_n N_A_398_74#_c_324_n
+ N_A_398_74#_c_325_n N_A_398_74#_c_326_n N_A_398_74#_c_348_n
+ N_A_398_74#_c_327_n N_A_398_74#_c_328_n N_A_398_74#_c_329_n
+ PM_SKY130_FD_SC_LS__DFSTP_2%A_398_74#
x_PM_SKY130_FD_SC_LS__DFSTP_2%A_767_384# N_A_767_384#_M1001_s
+ N_A_767_384#_M1004_d N_A_767_384#_c_584_n N_A_767_384#_M1033_g
+ N_A_767_384#_c_585_n N_A_767_384#_c_580_n N_A_767_384#_M1022_g
+ N_A_767_384#_c_586_n N_A_767_384#_c_587_n N_A_767_384#_c_588_n
+ N_A_767_384#_c_581_n N_A_767_384#_c_589_n N_A_767_384#_c_590_n
+ N_A_767_384#_c_582_n N_A_767_384#_c_583_n
+ PM_SKY130_FD_SC_LS__DFSTP_2%A_767_384#
x_PM_SKY130_FD_SC_LS__DFSTP_2%A_612_74# N_A_612_74#_M1019_d N_A_612_74#_M1000_d
+ N_A_612_74#_c_664_n N_A_612_74#_c_679_n N_A_612_74#_M1004_g
+ N_A_612_74#_M1001_g N_A_612_74#_c_666_n N_A_612_74#_M1005_g
+ N_A_612_74#_M1031_g N_A_612_74#_c_668_n N_A_612_74#_c_669_n
+ N_A_612_74#_c_670_n N_A_612_74#_c_671_n N_A_612_74#_c_672_n
+ N_A_612_74#_c_681_n N_A_612_74#_c_673_n N_A_612_74#_c_674_n
+ N_A_612_74#_c_675_n N_A_612_74#_c_683_n N_A_612_74#_c_676_n
+ N_A_612_74#_c_677_n PM_SKY130_FD_SC_LS__DFSTP_2%A_612_74#
x_PM_SKY130_FD_SC_LS__DFSTP_2%SET_B N_SET_B_c_801_n N_SET_B_M1008_g
+ N_SET_B_M1020_g N_SET_B_M1002_g N_SET_B_c_803_n N_SET_B_c_804_n
+ N_SET_B_M1021_g N_SET_B_c_798_n N_SET_B_c_806_n N_SET_B_c_807_n
+ N_SET_B_c_808_n N_SET_B_c_809_n SET_B N_SET_B_c_799_n N_SET_B_c_800_n
+ PM_SKY130_FD_SC_LS__DFSTP_2%SET_B
x_PM_SKY130_FD_SC_LS__DFSTP_2%A_225_74# N_A_225_74#_M1029_s N_A_225_74#_M1028_s
+ N_A_225_74#_M1016_g N_A_225_74#_c_921_n N_A_225_74#_M1007_g
+ N_A_225_74#_c_922_n N_A_225_74#_c_935_n N_A_225_74#_c_923_n
+ N_A_225_74#_c_924_n N_A_225_74#_c_936_n N_A_225_74#_c_937_n
+ N_A_225_74#_M1019_g N_A_225_74#_c_938_n N_A_225_74#_c_939_n
+ N_A_225_74#_c_940_n N_A_225_74#_M1010_g N_A_225_74#_c_941_n
+ N_A_225_74#_M1006_g N_A_225_74#_c_926_n N_A_225_74#_c_927_n
+ N_A_225_74#_M1009_g N_A_225_74#_c_929_n N_A_225_74#_c_930_n
+ N_A_225_74#_c_947_n N_A_225_74#_c_931_n N_A_225_74#_c_949_n
+ N_A_225_74#_c_950_n N_A_225_74#_c_951_n N_A_225_74#_c_932_n
+ N_A_225_74#_c_933_n N_A_225_74#_c_953_n PM_SKY130_FD_SC_LS__DFSTP_2%A_225_74#
x_PM_SKY130_FD_SC_LS__DFSTP_2%A_1566_92# N_A_1566_92#_M1024_d
+ N_A_1566_92#_M1030_d N_A_1566_92#_M1025_g N_A_1566_92#_c_1122_n
+ N_A_1566_92#_c_1123_n N_A_1566_92#_M1012_g N_A_1566_92#_c_1114_n
+ N_A_1566_92#_c_1124_n N_A_1566_92#_c_1115_n N_A_1566_92#_c_1116_n
+ N_A_1566_92#_c_1117_n N_A_1566_92#_c_1118_n N_A_1566_92#_c_1119_n
+ N_A_1566_92#_c_1120_n N_A_1566_92#_c_1121_n N_A_1566_92#_c_1127_n
+ PM_SKY130_FD_SC_LS__DFSTP_2%A_1566_92#
x_PM_SKY130_FD_SC_LS__DFSTP_2%A_1356_74# N_A_1356_74#_M1032_d
+ N_A_1356_74#_M1006_d N_A_1356_74#_M1021_d N_A_1356_74#_M1024_g
+ N_A_1356_74#_c_1207_n N_A_1356_74#_M1030_g N_A_1356_74#_c_1200_n
+ N_A_1356_74#_M1015_g N_A_1356_74#_c_1209_n N_A_1356_74#_M1027_g
+ N_A_1356_74#_c_1202_n N_A_1356_74#_c_1211_n N_A_1356_74#_c_1203_n
+ N_A_1356_74#_c_1213_n N_A_1356_74#_c_1204_n N_A_1356_74#_c_1233_n
+ N_A_1356_74#_c_1214_n N_A_1356_74#_c_1215_n N_A_1356_74#_c_1216_n
+ N_A_1356_74#_c_1217_n N_A_1356_74#_c_1205_n N_A_1356_74#_c_1219_n
+ N_A_1356_74#_c_1206_n N_A_1356_74#_c_1220_n N_A_1356_74#_c_1243_n
+ N_A_1356_74#_c_1221_n PM_SKY130_FD_SC_LS__DFSTP_2%A_1356_74#
x_PM_SKY130_FD_SC_LS__DFSTP_2%A_2022_94# N_A_2022_94#_M1015_s
+ N_A_2022_94#_M1027_s N_A_2022_94#_c_1363_n N_A_2022_94#_M1011_g
+ N_A_2022_94#_M1003_g N_A_2022_94#_M1023_g N_A_2022_94#_c_1364_n
+ N_A_2022_94#_M1017_g N_A_2022_94#_c_1359_n N_A_2022_94#_c_1365_n
+ N_A_2022_94#_c_1360_n N_A_2022_94#_c_1361_n N_A_2022_94#_c_1362_n
+ PM_SKY130_FD_SC_LS__DFSTP_2%A_2022_94#
x_PM_SKY130_FD_SC_LS__DFSTP_2%A_27_74# N_A_27_74#_M1026_s N_A_27_74#_M1019_s
+ N_A_27_74#_M1018_s N_A_27_74#_M1000_s N_A_27_74#_c_1425_n N_A_27_74#_c_1430_n
+ N_A_27_74#_c_1431_n N_A_27_74#_c_1432_n N_A_27_74#_c_1426_n
+ N_A_27_74#_c_1427_n N_A_27_74#_c_1434_n N_A_27_74#_c_1480_n
+ N_A_27_74#_c_1428_n PM_SKY130_FD_SC_LS__DFSTP_2%A_27_74#
x_PM_SKY130_FD_SC_LS__DFSTP_2%VPWR N_VPWR_M1018_d N_VPWR_M1028_d N_VPWR_M1033_d
+ N_VPWR_M1008_d N_VPWR_M1012_d N_VPWR_M1030_s N_VPWR_M1027_d N_VPWR_M1017_s
+ N_VPWR_c_1497_n N_VPWR_c_1498_n N_VPWR_c_1499_n N_VPWR_c_1500_n
+ N_VPWR_c_1501_n N_VPWR_c_1502_n N_VPWR_c_1503_n N_VPWR_c_1504_n
+ N_VPWR_c_1505_n N_VPWR_c_1506_n N_VPWR_c_1507_n N_VPWR_c_1508_n VPWR
+ N_VPWR_c_1509_n N_VPWR_c_1510_n N_VPWR_c_1511_n N_VPWR_c_1512_n
+ N_VPWR_c_1513_n N_VPWR_c_1514_n N_VPWR_c_1515_n N_VPWR_c_1516_n
+ N_VPWR_c_1517_n N_VPWR_c_1518_n N_VPWR_c_1519_n N_VPWR_c_1520_n
+ N_VPWR_c_1521_n N_VPWR_c_1496_n PM_SKY130_FD_SC_LS__DFSTP_2%VPWR
x_PM_SKY130_FD_SC_LS__DFSTP_2%Q N_Q_M1003_s N_Q_M1011_d N_Q_c_1652_n
+ N_Q_c_1655_n N_Q_c_1653_n N_Q_c_1654_n Q Q N_Q_c_1658_n
+ PM_SKY130_FD_SC_LS__DFSTP_2%Q
x_PM_SKY130_FD_SC_LS__DFSTP_2%VGND N_VGND_M1026_d N_VGND_M1029_d N_VGND_M1022_d
+ N_VGND_M1020_d N_VGND_M1002_d N_VGND_M1015_d N_VGND_M1023_d N_VGND_c_1690_n
+ N_VGND_c_1691_n N_VGND_c_1692_n N_VGND_c_1693_n N_VGND_c_1694_n
+ N_VGND_c_1695_n N_VGND_c_1696_n N_VGND_c_1697_n VGND N_VGND_c_1698_n
+ N_VGND_c_1699_n N_VGND_c_1700_n N_VGND_c_1701_n N_VGND_c_1702_n
+ N_VGND_c_1703_n N_VGND_c_1704_n N_VGND_c_1705_n N_VGND_c_1706_n
+ N_VGND_c_1707_n N_VGND_c_1708_n N_VGND_c_1709_n
+ PM_SKY130_FD_SC_LS__DFSTP_2%VGND
cc_1 VNB N_D_c_245_n 0.0447809f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.795
cc_2 VNB N_D_M1026_g 0.0288784f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.58
cc_3 VNB N_D_c_247_n 0.025337f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.145
cc_4 VNB N_D_c_248_n 0.00269121f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.145
cc_5 VNB N_CLK_c_279_n 0.019964f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.175
cc_6 VNB N_CLK_c_280_n 0.036162f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.375
cc_7 VNB CLK 0.00873773f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.58
cc_8 VNB N_A_398_74#_c_312_n 0.0168103f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.58
cc_9 VNB N_A_398_74#_c_313_n 0.0368422f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_10 VNB N_A_398_74#_c_314_n 0.0112016f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_398_74#_M1014_g 0.0507397f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.145
cc_12 VNB N_A_398_74#_c_316_n 0.00150841f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.295
cc_13 VNB N_A_398_74#_c_317_n 0.0158463f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_398_74#_c_318_n 0.00264685f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_398_74#_c_319_n 0.00190286f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_398_74#_c_320_n 0.0012865f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_398_74#_c_321_n 0.00247322f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_398_74#_c_322_n 0.00213614f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_398_74#_c_323_n 0.0230647f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_398_74#_c_324_n 0.00190332f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_398_74#_c_325_n 0.0153419f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_398_74#_c_326_n 0.00680136f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_398_74#_c_327_n 0.00734472f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_398_74#_c_328_n 0.031744f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_398_74#_c_329_n 0.0197653f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_767_384#_c_580_n 0.0195194f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_27 VNB N_A_767_384#_c_581_n 0.0240574f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_767_384#_c_582_n 0.0224227f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_767_384#_c_583_n 0.0535767f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_612_74#_c_664_n 0.00366225f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_612_74#_M1001_g 0.0241071f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_612_74#_c_666_n 0.0331869f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.145
cc_33 VNB N_A_612_74#_M1031_g 0.0253106f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.825
cc_34 VNB N_A_612_74#_c_668_n 0.00685615f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_612_74#_c_669_n 0.0205132f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_612_74#_c_670_n 0.00415803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_612_74#_c_671_n 0.00363794f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_612_74#_c_672_n 0.00239084f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_612_74#_c_673_n 0.00313488f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_612_74#_c_674_n 0.00482349f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_612_74#_c_675_n 0.00993512f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_612_74#_c_676_n 0.0192723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_612_74#_c_677_n 0.0304134f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_SET_B_M1020_g 0.0410395f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.58
cc_45 VNB N_SET_B_M1002_g 0.04772f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.75
cc_46 VNB N_SET_B_c_798_n 9.90083e-19 $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.98
cc_47 VNB N_SET_B_c_799_n 0.0178127f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.825
cc_48 VNB N_SET_B_c_800_n 0.00389433f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_225_74#_M1016_g 0.0224523f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.465
cc_50 VNB N_A_225_74#_c_921_n 0.0123708f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.75
cc_51 VNB N_A_225_74#_c_922_n 0.00808021f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_225_74#_c_923_n 0.0340583f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.145
cc_53 VNB N_A_225_74#_c_924_n 0.010226f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.98
cc_54 VNB N_A_225_74#_M1019_g 0.0265626f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.145
cc_55 VNB N_A_225_74#_c_926_n 0.0106772f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_225_74#_c_927_n 0.00106868f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_225_74#_M1009_g 0.0502374f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_225_74#_c_929_n 0.0195076f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_225_74#_c_930_n 0.00971956f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_225_74#_c_931_n 0.0104758f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_225_74#_c_932_n 0.00365457f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_225_74#_c_933_n 0.0133435f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_1566_92#_c_1114_n 0.0188877f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.145
cc_64 VNB N_A_1566_92#_c_1115_n 0.0161793f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.825
cc_65 VNB N_A_1566_92#_c_1116_n 0.0283476f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.99
cc_66 VNB N_A_1566_92#_c_1117_n 0.0447681f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_1566_92#_c_1118_n 0.00788489f $X=-0.19 $Y=-0.245 $X2=0.64
+ $Y2=1.295
cc_68 VNB N_A_1566_92#_c_1119_n 0.00499052f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_1566_92#_c_1120_n 0.00759688f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_1566_92#_c_1121_n 0.00570228f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_1356_74#_M1024_g 0.0604445f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_72 VNB N_A_1356_74#_c_1200_n 0.0264413f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.145
cc_73 VNB N_A_1356_74#_M1015_g 0.0460006f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.825
cc_74 VNB N_A_1356_74#_c_1202_n 0.0107945f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_1356_74#_c_1203_n 0.00337962f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_1356_74#_c_1204_n 0.00606384f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_1356_74#_c_1205_n 0.00342147f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_1356_74#_c_1206_n 0.00447039f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_2022_94#_M1003_g 0.0229692f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_80 VNB N_A_2022_94#_M1023_g 0.0260335f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.145
cc_81 VNB N_A_2022_94#_c_1359_n 0.0125258f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.99
cc_82 VNB N_A_2022_94#_c_1360_n 0.0084f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_2022_94#_c_1361_n 0.00309584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_2022_94#_c_1362_n 0.0737363f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_27_74#_c_1425_n 0.0420755f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_27_74#_c_1426_n 0.00574528f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.145
cc_87 VNB N_A_27_74#_c_1427_n 0.0137638f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.295
cc_88 VNB N_A_27_74#_c_1428_n 0.00619147f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_VPWR_c_1496_n 0.502022f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_Q_c_1652_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.465
cc_91 VNB N_Q_c_1653_n 0.00143777f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.145
cc_92 VNB N_Q_c_1654_n 0.00457514f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.145
cc_93 VNB N_VGND_c_1690_n 0.00619735f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.145
cc_94 VNB N_VGND_c_1691_n 0.0224525f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.295
cc_95 VNB N_VGND_c_1692_n 0.00559476f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.825
cc_96 VNB N_VGND_c_1693_n 0.0163103f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_VGND_c_1694_n 0.0214836f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_VGND_c_1695_n 0.0164768f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_VGND_c_1696_n 0.010678f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_VGND_c_1697_n 0.0505491f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_VGND_c_1698_n 0.0175546f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_VGND_c_1699_n 0.0636081f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_VGND_c_1700_n 0.0313742f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_VGND_c_1701_n 0.113496f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_VGND_c_1702_n 0.0357284f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_VGND_c_1703_n 0.0195351f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_VGND_c_1704_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_VGND_c_1705_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_VGND_c_1706_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_1707_n 0.0112736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_1708_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_1709_n 0.696385f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VPB N_D_c_245_n 0.0126976f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.795
cc_114 VPB N_D_c_250_n 0.0313518f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.375
cc_115 VPB N_D_c_251_n 0.0313209f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.465
cc_116 VPB N_D_c_248_n 0.00207792f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.145
cc_117 VPB N_D_c_253_n 0.0244664f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.825
cc_118 VPB N_CLK_c_280_n 0.0230735f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.375
cc_119 VPB N_A_398_74#_c_312_n 0.00525997f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.58
cc_120 VPB N_A_398_74#_c_331_n 0.0416235f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_A_398_74#_c_332_n 0.014641f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.465
cc_122 VPB N_A_398_74#_c_313_n 0.0258782f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_123 VPB N_A_398_74#_c_314_n 0.00803075f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_A_398_74#_c_335_n 0.0582781f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.825
cc_125 VPB N_A_398_74#_c_336_n 0.021907f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 VPB N_A_398_74#_c_337_n 0.00295783f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_127 VPB N_A_398_74#_c_319_n 0.00207712f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_A_398_74#_c_320_n 0.00587373f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_129 VPB N_A_398_74#_c_340_n 0.00334946f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_A_398_74#_c_341_n 0.00858286f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_A_398_74#_c_342_n 0.00469938f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_A_398_74#_c_343_n 0.0159882f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_A_398_74#_c_344_n 0.00428736f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_A_398_74#_c_345_n 0.00229911f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_A_398_74#_c_322_n 0.00419714f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_A_398_74#_c_325_n 0.01332f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_A_398_74#_c_348_n 2.61361e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_A_767_384#_c_584_n 0.0148273f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.58
cc_139 VPB N_A_767_384#_c_585_n 0.0150258f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.75
cc_140 VPB N_A_767_384#_c_586_n 0.0248545f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.145
cc_141 VPB N_A_767_384#_c_587_n 0.0134053f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=0.98
cc_142 VPB N_A_767_384#_c_588_n 0.0357903f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.825
cc_143 VPB N_A_767_384#_c_589_n 0.00155413f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_144 VPB N_A_767_384#_c_590_n 0.00168453f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_145 VPB N_A_767_384#_c_582_n 0.00840486f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_146 VPB N_A_612_74#_c_664_n 0.0285239f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_147 VPB N_A_612_74#_c_679_n 0.0228766f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.465
cc_148 VPB N_A_612_74#_c_666_n 0.0333093f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.145
cc_149 VPB N_A_612_74#_c_681_n 0.00504088f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_150 VPB N_A_612_74#_c_673_n 0.00808624f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_151 VPB N_A_612_74#_c_683_n 0.00253708f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_152 VPB N_A_612_74#_c_676_n 0.00168218f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_153 VPB N_SET_B_c_801_n 0.0561862f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.175
cc_154 VPB N_SET_B_M1020_g 0.0117516f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.58
cc_155 VPB N_SET_B_c_803_n 0.0152279f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_156 VPB N_SET_B_c_804_n 0.0240784f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_157 VPB N_SET_B_c_798_n 0.0229134f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=0.98
cc_158 VPB N_SET_B_c_806_n 0.0160157f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.825
cc_159 VPB N_SET_B_c_807_n 0.0178302f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.825
cc_160 VPB N_SET_B_c_808_n 4.31814e-19 $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.825
cc_161 VPB N_SET_B_c_809_n 0.0043956f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_162 VPB SET_B 0.00404524f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_163 VPB N_SET_B_c_800_n 0.00416461f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_164 VPB N_A_225_74#_c_921_n 0.0210337f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.75
cc_165 VPB N_A_225_74#_c_935_n 0.0754345f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.145
cc_166 VPB N_A_225_74#_c_936_n 0.0561762f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.825
cc_167 VPB N_A_225_74#_c_937_n 0.0125859f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.825
cc_168 VPB N_A_225_74#_c_938_n 0.00746259f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.295
cc_169 VPB N_A_225_74#_c_939_n 0.0164245f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_170 VPB N_A_225_74#_c_940_n 0.0141807f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.665
cc_171 VPB N_A_225_74#_c_941_n 0.244573f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_172 VPB N_A_225_74#_M1006_g 0.0102628f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_173 VPB N_A_225_74#_c_926_n 0.0399382f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_174 VPB N_A_225_74#_c_927_n 0.0150893f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_175 VPB N_A_225_74#_c_929_n 0.011123f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_176 VPB N_A_225_74#_c_930_n 5.35904e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_177 VPB N_A_225_74#_c_947_n 0.00898675f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_178 VPB N_A_225_74#_c_931_n 0.00236347f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_179 VPB N_A_225_74#_c_949_n 0.00592994f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_180 VPB N_A_225_74#_c_950_n 0.00539283f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_181 VPB N_A_225_74#_c_951_n 0.00468204f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_182 VPB N_A_225_74#_c_932_n 5.33031e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_183 VPB N_A_225_74#_c_953_n 8.57544e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_184 VPB N_A_1566_92#_c_1122_n 0.0136639f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.75
cc_185 VPB N_A_1566_92#_c_1123_n 0.0209384f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_186 VPB N_A_1566_92#_c_1124_n 0.00129748f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=0.98
cc_187 VPB N_A_1566_92#_c_1116_n 0.0232163f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.99
cc_188 VPB N_A_1566_92#_c_1120_n 0.0230925f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_189 VPB N_A_1566_92#_c_1127_n 0.0160359f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_190 VPB N_A_1356_74#_c_1207_n 0.0211924f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_191 VPB N_A_1356_74#_c_1200_n 0.0317157f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.145
cc_192 VPB N_A_1356_74#_c_1209_n 0.0178722f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.99
cc_193 VPB N_A_1356_74#_c_1202_n 0.0076044f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_194 VPB N_A_1356_74#_c_1211_n 0.0434221f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.665
cc_195 VPB N_A_1356_74#_c_1203_n 0.00539632f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_196 VPB N_A_1356_74#_c_1213_n 0.00201305f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_197 VPB N_A_1356_74#_c_1214_n 0.00335263f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_198 VPB N_A_1356_74#_c_1215_n 0.00291932f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_199 VPB N_A_1356_74#_c_1216_n 0.00685144f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_200 VPB N_A_1356_74#_c_1217_n 0.0163396f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_201 VPB N_A_1356_74#_c_1205_n 4.98981e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_202 VPB N_A_1356_74#_c_1219_n 0.0280862f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_203 VPB N_A_1356_74#_c_1220_n 0.00541621f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_204 VPB N_A_1356_74#_c_1221_n 0.00857572f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_205 VPB N_A_2022_94#_c_1363_n 0.0169085f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.58
cc_206 VPB N_A_2022_94#_c_1364_n 0.0173548f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.145
cc_207 VPB N_A_2022_94#_c_1365_n 0.0137341f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_208 VPB N_A_2022_94#_c_1362_n 0.016423f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_209 VPB N_A_27_74#_c_1425_n 0.0250181f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_210 VPB N_A_27_74#_c_1430_n 0.0274899f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.145
cc_211 VPB N_A_27_74#_c_1431_n 0.0257471f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=0.98
cc_212 VPB N_A_27_74#_c_1432_n 0.0143569f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.825
cc_213 VPB N_A_27_74#_c_1426_n 0.00273955f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.145
cc_214 VPB N_A_27_74#_c_1434_n 0.0109364f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_215 VPB N_VPWR_c_1497_n 0.017335f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_216 VPB N_VPWR_c_1498_n 0.0065563f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_217 VPB N_VPWR_c_1499_n 0.00509177f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_218 VPB N_VPWR_c_1500_n 0.0066771f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_219 VPB N_VPWR_c_1501_n 0.00666708f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_220 VPB N_VPWR_c_1502_n 0.00996541f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_221 VPB N_VPWR_c_1503_n 0.0104462f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_222 VPB N_VPWR_c_1504_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_223 VPB N_VPWR_c_1505_n 0.063793f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_224 VPB N_VPWR_c_1506_n 0.00553856f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_225 VPB N_VPWR_c_1507_n 0.0549518f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_226 VPB N_VPWR_c_1508_n 0.006142f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_227 VPB N_VPWR_c_1509_n 0.0180274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_228 VPB N_VPWR_c_1510_n 0.0215753f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_229 VPB N_VPWR_c_1511_n 0.0523685f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_230 VPB N_VPWR_c_1512_n 0.0384523f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_231 VPB N_VPWR_c_1513_n 0.01948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_232 VPB N_VPWR_c_1514_n 0.0342956f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_233 VPB N_VPWR_c_1515_n 0.0180566f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_234 VPB N_VPWR_c_1516_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_235 VPB N_VPWR_c_1517_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_236 VPB N_VPWR_c_1518_n 0.00223285f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_237 VPB N_VPWR_c_1519_n 0.00330333f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_238 VPB N_VPWR_c_1520_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_239 VPB N_VPWR_c_1521_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_240 VPB N_VPWR_c_1496_n 0.12454f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_241 VPB N_Q_c_1655_n 0.0024312f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_242 VPB N_Q_c_1653_n 0.00104928f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.145
cc_243 VPB Q 0.00161434f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=0.98
cc_244 VPB N_Q_c_1658_n 0.00274714f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.825
cc_245 N_D_c_247_n N_CLK_c_279_n 0.00223659f $X=0.64 $Y=1.145 $X2=-0.19
+ $Y2=-0.245
cc_246 N_D_c_245_n N_CLK_c_280_n 0.00972409f $X=0.61 $Y=1.795 $X2=0 $Y2=0
cc_247 N_D_c_245_n N_A_225_74#_c_931_n 0.00357638f $X=0.61 $Y=1.795 $X2=0 $Y2=0
cc_248 N_D_c_245_n N_A_225_74#_c_950_n 0.00302188f $X=0.61 $Y=1.795 $X2=0 $Y2=0
cc_249 N_D_c_250_n N_A_225_74#_c_950_n 9.40485e-19 $X=0.505 $Y=2.375 $X2=0 $Y2=0
cc_250 N_D_c_248_n N_A_225_74#_c_950_n 0.0224944f $X=0.64 $Y=1.145 $X2=0 $Y2=0
cc_251 N_D_M1026_g N_A_225_74#_c_933_n 0.00721478f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_252 N_D_c_247_n N_A_225_74#_c_933_n 0.00357638f $X=0.64 $Y=1.145 $X2=0 $Y2=0
cc_253 N_D_c_248_n N_A_225_74#_c_933_n 0.0556869f $X=0.64 $Y=1.145 $X2=0 $Y2=0
cc_254 N_D_M1026_g N_A_27_74#_c_1425_n 0.00743437f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_255 N_D_c_247_n N_A_27_74#_c_1425_n 0.0320429f $X=0.64 $Y=1.145 $X2=0 $Y2=0
cc_256 N_D_c_248_n N_A_27_74#_c_1425_n 0.0697394f $X=0.64 $Y=1.145 $X2=0 $Y2=0
cc_257 N_D_c_250_n N_A_27_74#_c_1430_n 0.00433476f $X=0.505 $Y=2.375 $X2=0 $Y2=0
cc_258 N_D_c_251_n N_A_27_74#_c_1430_n 0.00528173f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_259 N_D_c_250_n N_A_27_74#_c_1431_n 0.0216554f $X=0.505 $Y=2.375 $X2=0 $Y2=0
cc_260 N_D_c_248_n N_A_27_74#_c_1431_n 0.0227191f $X=0.64 $Y=1.145 $X2=0 $Y2=0
cc_261 N_D_c_253_n N_A_27_74#_c_1431_n 0.00140505f $X=0.64 $Y=1.825 $X2=0 $Y2=0
cc_262 N_D_c_251_n N_VPWR_c_1497_n 0.0138303f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_263 N_D_c_251_n N_VPWR_c_1509_n 0.00413917f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_264 N_D_c_251_n N_VPWR_c_1496_n 0.00859049f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_265 N_D_M1026_g N_VGND_c_1690_n 0.0140619f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_266 N_D_c_247_n N_VGND_c_1690_n 0.00150697f $X=0.64 $Y=1.145 $X2=0 $Y2=0
cc_267 N_D_c_248_n N_VGND_c_1690_n 0.0158023f $X=0.64 $Y=1.145 $X2=0 $Y2=0
cc_268 N_D_M1026_g N_VGND_c_1698_n 0.00383152f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_269 N_D_M1026_g N_VGND_c_1709_n 0.00761198f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_270 N_CLK_c_279_n N_A_225_74#_M1016_g 0.0131399f $X=1.485 $Y=1.22 $X2=0 $Y2=0
cc_271 N_CLK_c_280_n N_A_225_74#_M1016_g 0.0210236f $X=1.515 $Y=1.715 $X2=0
+ $Y2=0
cc_272 CLK N_A_225_74#_M1016_g 0.00369616f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_273 N_CLK_c_280_n N_A_225_74#_c_921_n 0.0477833f $X=1.515 $Y=1.715 $X2=0
+ $Y2=0
cc_274 N_CLK_c_279_n N_A_225_74#_c_931_n 0.00321998f $X=1.485 $Y=1.22 $X2=0
+ $Y2=0
cc_275 N_CLK_c_280_n N_A_225_74#_c_931_n 0.0065169f $X=1.515 $Y=1.715 $X2=0
+ $Y2=0
cc_276 CLK N_A_225_74#_c_931_n 0.0286813f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_277 N_CLK_c_280_n N_A_225_74#_c_949_n 0.00313913f $X=1.515 $Y=1.715 $X2=0
+ $Y2=0
cc_278 N_CLK_c_280_n N_A_225_74#_c_951_n 0.00952984f $X=1.515 $Y=1.715 $X2=0
+ $Y2=0
cc_279 N_CLK_c_280_n N_A_225_74#_c_932_n 0.00111203f $X=1.515 $Y=1.715 $X2=0
+ $Y2=0
cc_280 CLK N_A_225_74#_c_932_n 0.0203335f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_281 N_CLK_c_279_n N_A_225_74#_c_933_n 0.00791767f $X=1.485 $Y=1.22 $X2=0
+ $Y2=0
cc_282 N_CLK_c_280_n N_A_225_74#_c_933_n 0.00114511f $X=1.515 $Y=1.715 $X2=0
+ $Y2=0
cc_283 CLK N_A_225_74#_c_933_n 0.00762435f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_284 N_CLK_c_280_n N_A_225_74#_c_953_n 0.00477306f $X=1.515 $Y=1.715 $X2=0
+ $Y2=0
cc_285 CLK N_A_225_74#_c_953_n 0.0353587f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_286 N_CLK_c_280_n N_A_27_74#_c_1431_n 0.0161052f $X=1.515 $Y=1.715 $X2=0
+ $Y2=0
cc_287 CLK N_A_27_74#_c_1426_n 0.00323107f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_288 N_CLK_c_280_n N_VPWR_c_1497_n 0.0127906f $X=1.515 $Y=1.715 $X2=0 $Y2=0
cc_289 N_CLK_c_280_n N_VPWR_c_1498_n 0.0238569f $X=1.515 $Y=1.715 $X2=0 $Y2=0
cc_290 N_CLK_c_280_n N_VPWR_c_1510_n 0.0048608f $X=1.515 $Y=1.715 $X2=0 $Y2=0
cc_291 N_CLK_c_280_n N_VPWR_c_1496_n 0.00480464f $X=1.515 $Y=1.715 $X2=0 $Y2=0
cc_292 N_CLK_c_279_n N_VGND_c_1690_n 0.00295547f $X=1.485 $Y=1.22 $X2=0 $Y2=0
cc_293 N_CLK_c_279_n N_VGND_c_1691_n 0.00434272f $X=1.485 $Y=1.22 $X2=0 $Y2=0
cc_294 N_CLK_c_279_n N_VGND_c_1692_n 0.00294833f $X=1.485 $Y=1.22 $X2=0 $Y2=0
cc_295 CLK N_VGND_c_1692_n 0.013855f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_296 N_CLK_c_279_n N_VGND_c_1709_n 0.00825381f $X=1.485 $Y=1.22 $X2=0 $Y2=0
cc_297 N_A_398_74#_c_320_n N_A_767_384#_c_584_n 0.00181075f $X=3.77 $Y=1.545
+ $X2=0 $Y2=0
cc_298 N_A_398_74#_c_340_n N_A_767_384#_c_584_n 0.00225077f $X=3.71 $Y=2.89
+ $X2=0 $Y2=0
cc_299 N_A_398_74#_c_341_n N_A_767_384#_c_584_n 0.0100039f $X=4.745 $Y=2.325
+ $X2=0 $Y2=0
cc_300 N_A_398_74#_c_348_n N_A_767_384#_c_584_n 0.00403791f $X=3.77 $Y=2.325
+ $X2=0 $Y2=0
cc_301 N_A_398_74#_c_341_n N_A_767_384#_c_585_n 0.0138336f $X=4.745 $Y=2.325
+ $X2=0 $Y2=0
cc_302 N_A_398_74#_M1014_g N_A_767_384#_c_580_n 0.043019f $X=3.83 $Y=0.58 $X2=0
+ $Y2=0
cc_303 N_A_398_74#_c_331_n N_A_767_384#_c_586_n 0.00118696f $X=2.95 $Y=1.885
+ $X2=0 $Y2=0
cc_304 N_A_398_74#_c_314_n N_A_767_384#_c_586_n 0.00675415f $X=3.83 $Y=1.38
+ $X2=0 $Y2=0
cc_305 N_A_398_74#_c_320_n N_A_767_384#_c_586_n 0.0157854f $X=3.77 $Y=1.545
+ $X2=0 $Y2=0
cc_306 N_A_398_74#_c_341_n N_A_767_384#_c_586_n 6.41468e-19 $X=4.745 $Y=2.325
+ $X2=0 $Y2=0
cc_307 N_A_398_74#_c_320_n N_A_767_384#_c_587_n 0.0165446f $X=3.77 $Y=1.545
+ $X2=0 $Y2=0
cc_308 N_A_398_74#_c_341_n N_A_767_384#_c_587_n 0.0544703f $X=4.745 $Y=2.325
+ $X2=0 $Y2=0
cc_309 N_A_398_74#_c_320_n N_A_767_384#_c_588_n 0.00117498f $X=3.77 $Y=1.545
+ $X2=0 $Y2=0
cc_310 N_A_398_74#_M1014_g N_A_767_384#_c_581_n 6.56857e-19 $X=3.83 $Y=0.58
+ $X2=0 $Y2=0
cc_311 N_A_398_74#_c_342_n N_A_767_384#_c_589_n 0.0119623f $X=4.83 $Y=2.89 $X2=0
+ $Y2=0
cc_312 N_A_398_74#_c_343_n N_A_767_384#_c_589_n 0.020429f $X=5.52 $Y=2.975 $X2=0
+ $Y2=0
cc_313 N_A_398_74#_c_345_n N_A_767_384#_c_589_n 0.0167159f $X=5.605 $Y=2.89
+ $X2=0 $Y2=0
cc_314 N_A_398_74#_c_366_p N_A_767_384#_c_589_n 0.0137878f $X=5.69 $Y=2.405
+ $X2=0 $Y2=0
cc_315 N_A_398_74#_c_341_n N_A_767_384#_c_590_n 0.00778912f $X=4.745 $Y=2.325
+ $X2=0 $Y2=0
cc_316 N_A_398_74#_c_314_n N_A_767_384#_c_582_n 0.00809956f $X=3.83 $Y=1.38
+ $X2=0 $Y2=0
cc_317 N_A_398_74#_c_320_n N_A_767_384#_c_582_n 0.00165073f $X=3.77 $Y=1.545
+ $X2=0 $Y2=0
cc_318 N_A_398_74#_M1014_g N_A_767_384#_c_583_n 0.00534415f $X=3.83 $Y=0.58
+ $X2=0 $Y2=0
cc_319 N_A_398_74#_c_341_n N_A_612_74#_c_679_n 0.00343009f $X=4.745 $Y=2.325
+ $X2=0 $Y2=0
cc_320 N_A_398_74#_c_342_n N_A_612_74#_c_679_n 0.00905109f $X=4.83 $Y=2.89 $X2=0
+ $Y2=0
cc_321 N_A_398_74#_c_343_n N_A_612_74#_c_679_n 0.00364277f $X=5.52 $Y=2.975
+ $X2=0 $Y2=0
cc_322 N_A_398_74#_c_345_n N_A_612_74#_c_679_n 4.26354e-19 $X=5.605 $Y=2.89
+ $X2=0 $Y2=0
cc_323 N_A_398_74#_c_345_n N_A_612_74#_c_666_n 0.00293952f $X=5.605 $Y=2.89
+ $X2=0 $Y2=0
cc_324 N_A_398_74#_c_376_p N_A_612_74#_c_666_n 0.0115077f $X=6.415 $Y=2.405
+ $X2=0 $Y2=0
cc_325 N_A_398_74#_c_322_n N_A_612_74#_c_666_n 0.0169858f $X=6.5 $Y=2.32 $X2=0
+ $Y2=0
cc_326 N_A_398_74#_c_328_n N_A_612_74#_c_666_n 0.0283335f $X=6.795 $Y=1.285
+ $X2=0 $Y2=0
cc_327 N_A_398_74#_c_321_n N_A_612_74#_M1031_g 0.00450375f $X=6.5 $Y=1.12 $X2=0
+ $Y2=0
cc_328 N_A_398_74#_c_324_n N_A_612_74#_M1031_g 0.0010322f $X=6.585 $Y=0.365
+ $X2=0 $Y2=0
cc_329 N_A_398_74#_c_327_n N_A_612_74#_M1031_g 0.00497904f $X=6.795 $Y=1.285
+ $X2=0 $Y2=0
cc_330 N_A_398_74#_c_329_n N_A_612_74#_M1031_g 0.0283335f $X=6.795 $Y=1.12 $X2=0
+ $Y2=0
cc_331 N_A_398_74#_M1014_g N_A_612_74#_c_668_n 0.0143447f $X=3.83 $Y=0.58 $X2=0
+ $Y2=0
cc_332 N_A_398_74#_c_326_n N_A_612_74#_c_668_n 0.0343771f $X=2.95 $Y=1.38 $X2=0
+ $Y2=0
cc_333 N_A_398_74#_c_313_n N_A_612_74#_c_669_n 0.0013004f $X=3.755 $Y=1.545
+ $X2=0 $Y2=0
cc_334 N_A_398_74#_c_314_n N_A_612_74#_c_669_n 8.52337e-19 $X=3.83 $Y=1.38 $X2=0
+ $Y2=0
cc_335 N_A_398_74#_M1014_g N_A_612_74#_c_669_n 0.0169962f $X=3.83 $Y=0.58 $X2=0
+ $Y2=0
cc_336 N_A_398_74#_c_320_n N_A_612_74#_c_669_n 0.0224126f $X=3.77 $Y=1.545 $X2=0
+ $Y2=0
cc_337 N_A_398_74#_M1014_g N_A_612_74#_c_670_n 0.0020456f $X=3.83 $Y=0.58 $X2=0
+ $Y2=0
cc_338 N_A_398_74#_c_320_n N_A_612_74#_c_670_n 0.00145075f $X=3.77 $Y=1.545
+ $X2=0 $Y2=0
cc_339 N_A_398_74#_c_314_n N_A_612_74#_c_671_n 0.00187189f $X=3.83 $Y=1.38 $X2=0
+ $Y2=0
cc_340 N_A_398_74#_c_320_n N_A_612_74#_c_671_n 0.0142106f $X=3.77 $Y=1.545 $X2=0
+ $Y2=0
cc_341 N_A_398_74#_c_341_n N_A_612_74#_c_671_n 0.00453594f $X=4.745 $Y=2.325
+ $X2=0 $Y2=0
cc_342 N_A_398_74#_c_332_n N_A_612_74#_c_681_n 0.00257632f $X=3.005 $Y=2.205
+ $X2=0 $Y2=0
cc_343 N_A_398_74#_c_313_n N_A_612_74#_c_681_n 0.00478473f $X=3.755 $Y=1.545
+ $X2=0 $Y2=0
cc_344 N_A_398_74#_c_336_n N_A_612_74#_c_681_n 0.0261466f $X=3.625 $Y=2.975
+ $X2=0 $Y2=0
cc_345 N_A_398_74#_c_340_n N_A_612_74#_c_681_n 0.0124001f $X=3.71 $Y=2.89 $X2=0
+ $Y2=0
cc_346 N_A_398_74#_c_331_n N_A_612_74#_c_673_n 0.00909258f $X=2.95 $Y=1.885
+ $X2=0 $Y2=0
cc_347 N_A_398_74#_c_332_n N_A_612_74#_c_673_n 5.65712e-19 $X=3.005 $Y=2.205
+ $X2=0 $Y2=0
cc_348 N_A_398_74#_c_313_n N_A_612_74#_c_673_n 0.022329f $X=3.755 $Y=1.545 $X2=0
+ $Y2=0
cc_349 N_A_398_74#_M1014_g N_A_612_74#_c_673_n 0.00339481f $X=3.83 $Y=0.58 $X2=0
+ $Y2=0
cc_350 N_A_398_74#_c_320_n N_A_612_74#_c_673_n 0.0645348f $X=3.77 $Y=1.545 $X2=0
+ $Y2=0
cc_351 N_A_398_74#_c_326_n N_A_612_74#_c_673_n 0.0617327f $X=2.95 $Y=1.38 $X2=0
+ $Y2=0
cc_352 N_A_398_74#_c_348_n N_A_612_74#_c_673_n 0.00814612f $X=3.77 $Y=2.325
+ $X2=0 $Y2=0
cc_353 N_A_398_74#_c_313_n N_A_612_74#_c_674_n 0.00711061f $X=3.755 $Y=1.545
+ $X2=0 $Y2=0
cc_354 N_A_398_74#_c_326_n N_A_612_74#_c_674_n 0.0143569f $X=2.95 $Y=1.38 $X2=0
+ $Y2=0
cc_355 N_A_398_74#_c_322_n N_A_612_74#_c_683_n 0.00950869f $X=6.5 $Y=2.32 $X2=0
+ $Y2=0
cc_356 N_A_398_74#_c_327_n N_A_612_74#_c_683_n 0.0204128f $X=6.795 $Y=1.285
+ $X2=0 $Y2=0
cc_357 N_A_398_74#_c_343_n N_SET_B_c_801_n 0.00292991f $X=5.52 $Y=2.975
+ $X2=-0.19 $Y2=-0.245
cc_358 N_A_398_74#_c_345_n N_SET_B_c_801_n 0.00942707f $X=5.605 $Y=2.89
+ $X2=-0.19 $Y2=-0.245
cc_359 N_A_398_74#_c_376_p N_SET_B_c_801_n 4.19495e-19 $X=6.415 $Y=2.405
+ $X2=-0.19 $Y2=-0.245
cc_360 N_A_398_74#_c_366_p N_SET_B_c_801_n 0.00662706f $X=5.69 $Y=2.405
+ $X2=-0.19 $Y2=-0.245
cc_361 N_A_398_74#_c_335_n N_SET_B_c_807_n 5.05992e-19 $X=7.53 $Y=2.465 $X2=0
+ $Y2=0
cc_362 N_A_398_74#_c_376_p N_SET_B_c_807_n 0.010574f $X=6.415 $Y=2.405 $X2=0
+ $Y2=0
cc_363 N_A_398_74#_c_322_n N_SET_B_c_807_n 0.0176826f $X=6.5 $Y=2.32 $X2=0 $Y2=0
cc_364 N_A_398_74#_c_325_n N_SET_B_c_807_n 0.026653f $X=7.575 $Y=1.98 $X2=0
+ $Y2=0
cc_365 N_A_398_74#_c_327_n N_SET_B_c_807_n 0.00748379f $X=6.795 $Y=1.285 $X2=0
+ $Y2=0
cc_366 N_A_398_74#_c_328_n N_SET_B_c_807_n 0.00149631f $X=6.795 $Y=1.285 $X2=0
+ $Y2=0
cc_367 N_A_398_74#_c_376_p N_SET_B_c_808_n 0.00857725f $X=6.415 $Y=2.405 $X2=0
+ $Y2=0
cc_368 N_A_398_74#_c_322_n N_SET_B_c_808_n 0.0024765f $X=6.5 $Y=2.32 $X2=0 $Y2=0
cc_369 N_A_398_74#_c_376_p N_SET_B_c_809_n 0.0297221f $X=6.415 $Y=2.405 $X2=0
+ $Y2=0
cc_370 N_A_398_74#_c_366_p N_SET_B_c_809_n 0.0118997f $X=5.69 $Y=2.405 $X2=0
+ $Y2=0
cc_371 N_A_398_74#_c_322_n N_SET_B_c_809_n 0.0154685f $X=6.5 $Y=2.32 $X2=0 $Y2=0
cc_372 N_A_398_74#_c_325_n SET_B 4.96175e-19 $X=7.575 $Y=1.98 $X2=0 $Y2=0
cc_373 N_A_398_74#_c_325_n N_SET_B_c_800_n 3.31672e-19 $X=7.575 $Y=1.98 $X2=0
+ $Y2=0
cc_374 N_A_398_74#_c_316_n N_A_225_74#_M1016_g 0.00164183f $X=2.13 $Y=0.515
+ $X2=0 $Y2=0
cc_375 N_A_398_74#_c_318_n N_A_225_74#_M1016_g 0.00266901f $X=2.215 $Y=0.34
+ $X2=0 $Y2=0
cc_376 N_A_398_74#_c_428_p N_A_225_74#_c_921_n 0.00418454f $X=2.19 $Y=2.665
+ $X2=0 $Y2=0
cc_377 N_A_398_74#_c_337_n N_A_225_74#_c_921_n 0.00144647f $X=2.275 $Y=2.975
+ $X2=0 $Y2=0
cc_378 N_A_398_74#_c_326_n N_A_225_74#_c_922_n 8.19668e-19 $X=2.95 $Y=1.38 $X2=0
+ $Y2=0
cc_379 N_A_398_74#_c_331_n N_A_225_74#_c_935_n 0.0244246f $X=2.95 $Y=1.885 $X2=0
+ $Y2=0
cc_380 N_A_398_74#_c_332_n N_A_225_74#_c_935_n 0.0136783f $X=3.005 $Y=2.205
+ $X2=0 $Y2=0
cc_381 N_A_398_74#_c_428_p N_A_225_74#_c_935_n 0.00602998f $X=2.19 $Y=2.665
+ $X2=0 $Y2=0
cc_382 N_A_398_74#_c_336_n N_A_225_74#_c_935_n 0.0108241f $X=3.625 $Y=2.975
+ $X2=0 $Y2=0
cc_383 N_A_398_74#_c_319_n N_A_225_74#_c_935_n 3.78496e-19 $X=2.95 $Y=1.545
+ $X2=0 $Y2=0
cc_384 N_A_398_74#_c_312_n N_A_225_74#_c_923_n 0.0147005f $X=2.95 $Y=1.71 $X2=0
+ $Y2=0
cc_385 N_A_398_74#_c_317_n N_A_225_74#_c_923_n 0.00256866f $X=2.945 $Y=0.34
+ $X2=0 $Y2=0
cc_386 N_A_398_74#_c_319_n N_A_225_74#_c_923_n 0.00105733f $X=2.95 $Y=1.545
+ $X2=0 $Y2=0
cc_387 N_A_398_74#_c_326_n N_A_225_74#_c_923_n 0.0074497f $X=2.95 $Y=1.38 $X2=0
+ $Y2=0
cc_388 N_A_398_74#_c_316_n N_A_225_74#_c_924_n 0.00127231f $X=2.13 $Y=0.515
+ $X2=0 $Y2=0
cc_389 N_A_398_74#_c_317_n N_A_225_74#_c_924_n 9.7974e-19 $X=2.945 $Y=0.34 $X2=0
+ $Y2=0
cc_390 N_A_398_74#_c_332_n N_A_225_74#_c_936_n 0.00716579f $X=3.005 $Y=2.205
+ $X2=0 $Y2=0
cc_391 N_A_398_74#_c_336_n N_A_225_74#_c_936_n 0.0133272f $X=3.625 $Y=2.975
+ $X2=0 $Y2=0
cc_392 N_A_398_74#_M1014_g N_A_225_74#_M1019_g 0.0087307f $X=3.83 $Y=0.58 $X2=0
+ $Y2=0
cc_393 N_A_398_74#_c_316_n N_A_225_74#_M1019_g 0.00387291f $X=2.13 $Y=0.515
+ $X2=0 $Y2=0
cc_394 N_A_398_74#_c_317_n N_A_225_74#_M1019_g 0.0106029f $X=2.945 $Y=0.34 $X2=0
+ $Y2=0
cc_395 N_A_398_74#_c_326_n N_A_225_74#_M1019_g 0.021296f $X=2.95 $Y=1.38 $X2=0
+ $Y2=0
cc_396 N_A_398_74#_c_332_n N_A_225_74#_c_938_n 0.00215978f $X=3.005 $Y=2.205
+ $X2=0 $Y2=0
cc_397 N_A_398_74#_c_340_n N_A_225_74#_c_938_n 0.00374862f $X=3.71 $Y=2.89 $X2=0
+ $Y2=0
cc_398 N_A_398_74#_c_336_n N_A_225_74#_c_939_n 0.0182504f $X=3.625 $Y=2.975
+ $X2=0 $Y2=0
cc_399 N_A_398_74#_c_331_n N_A_225_74#_c_940_n 0.00177603f $X=2.95 $Y=1.885
+ $X2=0 $Y2=0
cc_400 N_A_398_74#_c_332_n N_A_225_74#_c_940_n 0.0105971f $X=3.005 $Y=2.205
+ $X2=0 $Y2=0
cc_401 N_A_398_74#_c_313_n N_A_225_74#_c_940_n 0.0056641f $X=3.755 $Y=1.545
+ $X2=0 $Y2=0
cc_402 N_A_398_74#_c_320_n N_A_225_74#_c_940_n 6.4886e-19 $X=3.77 $Y=1.545 $X2=0
+ $Y2=0
cc_403 N_A_398_74#_c_340_n N_A_225_74#_c_940_n 0.00266173f $X=3.71 $Y=2.89 $X2=0
+ $Y2=0
cc_404 N_A_398_74#_c_348_n N_A_225_74#_c_940_n 8.62673e-19 $X=3.77 $Y=2.325
+ $X2=0 $Y2=0
cc_405 N_A_398_74#_c_335_n N_A_225_74#_c_941_n 0.0013954f $X=7.53 $Y=2.465 $X2=0
+ $Y2=0
cc_406 N_A_398_74#_c_336_n N_A_225_74#_c_941_n 0.00485499f $X=3.625 $Y=2.975
+ $X2=0 $Y2=0
cc_407 N_A_398_74#_c_341_n N_A_225_74#_c_941_n 0.0048983f $X=4.745 $Y=2.325
+ $X2=0 $Y2=0
cc_408 N_A_398_74#_c_343_n N_A_225_74#_c_941_n 0.0134765f $X=5.52 $Y=2.975 $X2=0
+ $Y2=0
cc_409 N_A_398_74#_c_344_n N_A_225_74#_c_941_n 0.00417961f $X=4.915 $Y=2.975
+ $X2=0 $Y2=0
cc_410 N_A_398_74#_c_376_p N_A_225_74#_c_941_n 0.0117359f $X=6.415 $Y=2.405
+ $X2=0 $Y2=0
cc_411 N_A_398_74#_c_335_n N_A_225_74#_M1006_g 0.00790409f $X=7.53 $Y=2.465
+ $X2=0 $Y2=0
cc_412 N_A_398_74#_c_376_p N_A_225_74#_M1006_g 0.0016067f $X=6.415 $Y=2.405
+ $X2=0 $Y2=0
cc_413 N_A_398_74#_c_322_n N_A_225_74#_M1006_g 0.00332936f $X=6.5 $Y=2.32 $X2=0
+ $Y2=0
cc_414 N_A_398_74#_c_325_n N_A_225_74#_M1006_g 4.58926e-19 $X=7.575 $Y=1.98
+ $X2=0 $Y2=0
cc_415 N_A_398_74#_c_335_n N_A_225_74#_c_926_n 0.00860205f $X=7.53 $Y=2.465
+ $X2=0 $Y2=0
cc_416 N_A_398_74#_c_325_n N_A_225_74#_c_926_n 0.00260094f $X=7.575 $Y=1.98
+ $X2=0 $Y2=0
cc_417 N_A_398_74#_c_322_n N_A_225_74#_c_927_n 0.00217336f $X=6.5 $Y=2.32 $X2=0
+ $Y2=0
cc_418 N_A_398_74#_c_325_n N_A_225_74#_c_927_n 3.00547e-19 $X=7.575 $Y=1.98
+ $X2=0 $Y2=0
cc_419 N_A_398_74#_c_327_n N_A_225_74#_c_927_n 0.00130377f $X=6.795 $Y=1.285
+ $X2=0 $Y2=0
cc_420 N_A_398_74#_c_328_n N_A_225_74#_c_927_n 0.0196747f $X=6.795 $Y=1.285
+ $X2=0 $Y2=0
cc_421 N_A_398_74#_c_323_n N_A_225_74#_M1009_g 0.00697755f $X=7.49 $Y=0.365
+ $X2=0 $Y2=0
cc_422 N_A_398_74#_c_325_n N_A_225_74#_M1009_g 0.0129179f $X=7.575 $Y=1.98 $X2=0
+ $Y2=0
cc_423 N_A_398_74#_c_327_n N_A_225_74#_M1009_g 3.37207e-19 $X=6.795 $Y=1.285
+ $X2=0 $Y2=0
cc_424 N_A_398_74#_c_328_n N_A_225_74#_M1009_g 0.0118136f $X=6.795 $Y=1.285
+ $X2=0 $Y2=0
cc_425 N_A_398_74#_c_329_n N_A_225_74#_M1009_g 0.0128826f $X=6.795 $Y=1.12 $X2=0
+ $Y2=0
cc_426 N_A_398_74#_c_316_n N_A_225_74#_c_929_n 0.00106057f $X=2.13 $Y=0.515
+ $X2=0 $Y2=0
cc_427 N_A_398_74#_c_312_n N_A_225_74#_c_930_n 0.0196818f $X=2.95 $Y=1.71 $X2=0
+ $Y2=0
cc_428 N_A_398_74#_c_319_n N_A_225_74#_c_930_n 3.78496e-19 $X=2.95 $Y=1.545
+ $X2=0 $Y2=0
cc_429 N_A_398_74#_M1007_d N_A_225_74#_c_951_n 0.00293855f $X=2.04 $Y=1.79 $X2=0
+ $Y2=0
cc_430 N_A_398_74#_c_316_n N_A_225_74#_c_932_n 0.0147852f $X=2.13 $Y=0.515 $X2=0
+ $Y2=0
cc_431 N_A_398_74#_c_335_n N_A_1566_92#_c_1122_n 0.0180148f $X=7.53 $Y=2.465
+ $X2=0 $Y2=0
cc_432 N_A_398_74#_c_325_n N_A_1566_92#_c_1122_n 0.00132197f $X=7.575 $Y=1.98
+ $X2=0 $Y2=0
cc_433 N_A_398_74#_c_335_n N_A_1566_92#_c_1123_n 0.0281869f $X=7.53 $Y=2.465
+ $X2=0 $Y2=0
cc_434 N_A_398_74#_c_325_n N_A_1566_92#_c_1114_n 0.013857f $X=7.575 $Y=1.98
+ $X2=0 $Y2=0
cc_435 N_A_398_74#_c_325_n N_A_1566_92#_c_1124_n 0.0656794f $X=7.575 $Y=1.98
+ $X2=0 $Y2=0
cc_436 N_A_398_74#_c_325_n N_A_1566_92#_c_1115_n 0.00795872f $X=7.575 $Y=1.98
+ $X2=0 $Y2=0
cc_437 N_A_398_74#_c_325_n N_A_1566_92#_c_1118_n 0.0135436f $X=7.575 $Y=1.98
+ $X2=0 $Y2=0
cc_438 N_A_398_74#_c_335_n N_A_1566_92#_c_1127_n 0.00529714f $X=7.53 $Y=2.465
+ $X2=0 $Y2=0
cc_439 N_A_398_74#_c_325_n N_A_1566_92#_c_1127_n 0.00154377f $X=7.575 $Y=1.98
+ $X2=0 $Y2=0
cc_440 N_A_398_74#_c_323_n N_A_1356_74#_M1032_d 0.00227017f $X=7.49 $Y=0.365
+ $X2=-0.19 $Y2=-0.245
cc_441 N_A_398_74#_c_335_n N_A_1356_74#_c_1213_n 0.00461908f $X=7.53 $Y=2.465
+ $X2=0 $Y2=0
cc_442 N_A_398_74#_c_376_p N_A_1356_74#_c_1213_n 0.0107348f $X=6.415 $Y=2.405
+ $X2=0 $Y2=0
cc_443 N_A_398_74#_c_322_n N_A_1356_74#_c_1213_n 0.0285495f $X=6.5 $Y=2.32 $X2=0
+ $Y2=0
cc_444 N_A_398_74#_c_325_n N_A_1356_74#_c_1213_n 0.0313601f $X=7.575 $Y=1.98
+ $X2=0 $Y2=0
cc_445 N_A_398_74#_c_321_n N_A_1356_74#_c_1204_n 0.00444057f $X=6.5 $Y=1.12
+ $X2=0 $Y2=0
cc_446 N_A_398_74#_c_322_n N_A_1356_74#_c_1204_n 0.00556347f $X=6.5 $Y=2.32
+ $X2=0 $Y2=0
cc_447 N_A_398_74#_c_325_n N_A_1356_74#_c_1204_n 0.0456192f $X=7.575 $Y=1.98
+ $X2=0 $Y2=0
cc_448 N_A_398_74#_c_327_n N_A_1356_74#_c_1204_n 0.0236708f $X=6.795 $Y=1.285
+ $X2=0 $Y2=0
cc_449 N_A_398_74#_c_328_n N_A_1356_74#_c_1204_n 0.00110295f $X=6.795 $Y=1.285
+ $X2=0 $Y2=0
cc_450 N_A_398_74#_c_329_n N_A_1356_74#_c_1204_n 0.00140588f $X=6.795 $Y=1.12
+ $X2=0 $Y2=0
cc_451 N_A_398_74#_c_335_n N_A_1356_74#_c_1233_n 0.00820781f $X=7.53 $Y=2.465
+ $X2=0 $Y2=0
cc_452 N_A_398_74#_c_325_n N_A_1356_74#_c_1233_n 0.00180543f $X=7.575 $Y=1.98
+ $X2=0 $Y2=0
cc_453 N_A_398_74#_c_335_n N_A_1356_74#_c_1215_n 0.00413826f $X=7.53 $Y=2.465
+ $X2=0 $Y2=0
cc_454 N_A_398_74#_c_325_n N_A_1356_74#_c_1215_n 0.00449885f $X=7.575 $Y=1.98
+ $X2=0 $Y2=0
cc_455 N_A_398_74#_c_322_n N_A_1356_74#_c_1206_n 0.0103198f $X=6.5 $Y=2.32 $X2=0
+ $Y2=0
cc_456 N_A_398_74#_c_325_n N_A_1356_74#_c_1206_n 0.014742f $X=7.575 $Y=1.98
+ $X2=0 $Y2=0
cc_457 N_A_398_74#_c_327_n N_A_1356_74#_c_1206_n 0.0101698f $X=6.795 $Y=1.285
+ $X2=0 $Y2=0
cc_458 N_A_398_74#_c_328_n N_A_1356_74#_c_1206_n 7.38251e-19 $X=6.795 $Y=1.285
+ $X2=0 $Y2=0
cc_459 N_A_398_74#_c_335_n N_A_1356_74#_c_1220_n 0.0078896f $X=7.53 $Y=2.465
+ $X2=0 $Y2=0
cc_460 N_A_398_74#_c_325_n N_A_1356_74#_c_1220_n 0.0204053f $X=7.575 $Y=1.98
+ $X2=0 $Y2=0
cc_461 N_A_398_74#_c_323_n N_A_1356_74#_c_1243_n 0.0330935f $X=7.49 $Y=0.365
+ $X2=0 $Y2=0
cc_462 N_A_398_74#_c_327_n N_A_1356_74#_c_1243_n 0.00999825f $X=6.795 $Y=1.285
+ $X2=0 $Y2=0
cc_463 N_A_398_74#_c_328_n N_A_1356_74#_c_1243_n 0.00304494f $X=6.795 $Y=1.285
+ $X2=0 $Y2=0
cc_464 N_A_398_74#_c_317_n N_A_27_74#_M1019_s 0.00404388f $X=2.945 $Y=0.34 $X2=0
+ $Y2=0
cc_465 N_A_398_74#_M1007_d N_A_27_74#_c_1432_n 0.00598015f $X=2.04 $Y=1.79 $X2=0
+ $Y2=0
cc_466 N_A_398_74#_c_331_n N_A_27_74#_c_1432_n 0.0030474f $X=2.95 $Y=1.885 $X2=0
+ $Y2=0
cc_467 N_A_398_74#_c_332_n N_A_27_74#_c_1432_n 0.00630881f $X=3.005 $Y=2.205
+ $X2=0 $Y2=0
cc_468 N_A_398_74#_c_428_p N_A_27_74#_c_1432_n 0.0381703f $X=2.19 $Y=2.665 $X2=0
+ $Y2=0
cc_469 N_A_398_74#_c_336_n N_A_27_74#_c_1432_n 0.042362f $X=3.625 $Y=2.975 $X2=0
+ $Y2=0
cc_470 N_A_398_74#_c_319_n N_A_27_74#_c_1432_n 0.0116371f $X=2.95 $Y=1.545 $X2=0
+ $Y2=0
cc_471 N_A_398_74#_c_312_n N_A_27_74#_c_1426_n 0.0038721f $X=2.95 $Y=1.71 $X2=0
+ $Y2=0
cc_472 N_A_398_74#_c_316_n N_A_27_74#_c_1426_n 0.0116911f $X=2.13 $Y=0.515 $X2=0
+ $Y2=0
cc_473 N_A_398_74#_c_319_n N_A_27_74#_c_1426_n 0.0502423f $X=2.95 $Y=1.545 $X2=0
+ $Y2=0
cc_474 N_A_398_74#_c_326_n N_A_27_74#_c_1426_n 0.0201904f $X=2.95 $Y=1.38 $X2=0
+ $Y2=0
cc_475 N_A_398_74#_c_316_n N_A_27_74#_c_1428_n 0.0206593f $X=2.13 $Y=0.515 $X2=0
+ $Y2=0
cc_476 N_A_398_74#_c_317_n N_A_27_74#_c_1428_n 0.0239262f $X=2.945 $Y=0.34 $X2=0
+ $Y2=0
cc_477 N_A_398_74#_c_326_n N_A_27_74#_c_1428_n 0.0244211f $X=2.95 $Y=1.38 $X2=0
+ $Y2=0
cc_478 N_A_398_74#_c_341_n N_VPWR_M1033_d 0.0133836f $X=4.745 $Y=2.325 $X2=0
+ $Y2=0
cc_479 N_A_398_74#_c_342_n N_VPWR_M1033_d 0.0103108f $X=4.83 $Y=2.89 $X2=0 $Y2=0
cc_480 N_A_398_74#_c_345_n N_VPWR_M1008_d 0.00295815f $X=5.605 $Y=2.89 $X2=0
+ $Y2=0
cc_481 N_A_398_74#_c_376_p N_VPWR_M1008_d 0.010565f $X=6.415 $Y=2.405 $X2=0
+ $Y2=0
cc_482 N_A_398_74#_c_366_p N_VPWR_M1008_d 5.98664e-19 $X=5.69 $Y=2.405 $X2=0
+ $Y2=0
cc_483 N_A_398_74#_c_428_p N_VPWR_c_1498_n 0.0234171f $X=2.19 $Y=2.665 $X2=0
+ $Y2=0
cc_484 N_A_398_74#_c_337_n N_VPWR_c_1498_n 0.0127362f $X=2.275 $Y=2.975 $X2=0
+ $Y2=0
cc_485 N_A_398_74#_c_336_n N_VPWR_c_1499_n 0.00905466f $X=3.625 $Y=2.975 $X2=0
+ $Y2=0
cc_486 N_A_398_74#_c_344_n N_VPWR_c_1499_n 0.0059477f $X=4.915 $Y=2.975 $X2=0
+ $Y2=0
cc_487 N_A_398_74#_c_343_n N_VPWR_c_1500_n 0.0146305f $X=5.52 $Y=2.975 $X2=0
+ $Y2=0
cc_488 N_A_398_74#_c_345_n N_VPWR_c_1500_n 0.017418f $X=5.605 $Y=2.89 $X2=0
+ $Y2=0
cc_489 N_A_398_74#_c_376_p N_VPWR_c_1500_n 0.0189842f $X=6.415 $Y=2.405 $X2=0
+ $Y2=0
cc_490 N_A_398_74#_c_336_n N_VPWR_c_1506_n 0.00124242f $X=3.625 $Y=2.975 $X2=0
+ $Y2=0
cc_491 N_A_398_74#_c_340_n N_VPWR_c_1506_n 0.0147011f $X=3.71 $Y=2.89 $X2=0
+ $Y2=0
cc_492 N_A_398_74#_c_341_n N_VPWR_c_1506_n 0.038593f $X=4.745 $Y=2.325 $X2=0
+ $Y2=0
cc_493 N_A_398_74#_c_342_n N_VPWR_c_1506_n 0.0250726f $X=4.83 $Y=2.89 $X2=0
+ $Y2=0
cc_494 N_A_398_74#_c_344_n N_VPWR_c_1506_n 0.00174131f $X=4.915 $Y=2.975 $X2=0
+ $Y2=0
cc_495 N_A_398_74#_c_335_n N_VPWR_c_1507_n 0.00319296f $X=7.53 $Y=2.465 $X2=0
+ $Y2=0
cc_496 N_A_398_74#_c_336_n N_VPWR_c_1511_n 0.0896378f $X=3.625 $Y=2.975 $X2=0
+ $Y2=0
cc_497 N_A_398_74#_c_337_n N_VPWR_c_1511_n 0.0111058f $X=2.275 $Y=2.975 $X2=0
+ $Y2=0
cc_498 N_A_398_74#_c_343_n N_VPWR_c_1512_n 0.0466947f $X=5.52 $Y=2.975 $X2=0
+ $Y2=0
cc_499 N_A_398_74#_c_344_n N_VPWR_c_1512_n 0.0111256f $X=4.915 $Y=2.975 $X2=0
+ $Y2=0
cc_500 N_A_398_74#_c_335_n N_VPWR_c_1496_n 0.0040313f $X=7.53 $Y=2.465 $X2=0
+ $Y2=0
cc_501 N_A_398_74#_c_336_n N_VPWR_c_1496_n 0.051041f $X=3.625 $Y=2.975 $X2=0
+ $Y2=0
cc_502 N_A_398_74#_c_337_n N_VPWR_c_1496_n 0.0065564f $X=2.275 $Y=2.975 $X2=0
+ $Y2=0
cc_503 N_A_398_74#_c_343_n N_VPWR_c_1496_n 0.0260024f $X=5.52 $Y=2.975 $X2=0
+ $Y2=0
cc_504 N_A_398_74#_c_344_n N_VPWR_c_1496_n 0.00588338f $X=4.915 $Y=2.975 $X2=0
+ $Y2=0
cc_505 N_A_398_74#_c_376_p N_VPWR_c_1496_n 0.0209521f $X=6.415 $Y=2.405 $X2=0
+ $Y2=0
cc_506 N_A_398_74#_c_340_n A_716_456# 0.00127677f $X=3.71 $Y=2.89 $X2=-0.19
+ $Y2=-0.245
cc_507 N_A_398_74#_c_376_p A_1266_341# 0.00464741f $X=6.415 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_508 N_A_398_74#_c_322_n A_1266_341# 0.0161564f $X=6.5 $Y=2.32 $X2=-0.19
+ $Y2=-0.245
cc_509 N_A_398_74#_c_318_n N_VGND_c_1692_n 0.0109685f $X=2.215 $Y=0.34 $X2=0
+ $Y2=0
cc_510 N_A_398_74#_M1014_g N_VGND_c_1693_n 0.00175448f $X=3.83 $Y=0.58 $X2=0
+ $Y2=0
cc_511 N_A_398_74#_c_321_n N_VGND_c_1694_n 0.02453f $X=6.5 $Y=1.12 $X2=0 $Y2=0
cc_512 N_A_398_74#_c_324_n N_VGND_c_1694_n 0.0111625f $X=6.585 $Y=0.365 $X2=0
+ $Y2=0
cc_513 N_A_398_74#_c_329_n N_VGND_c_1694_n 5.00668e-19 $X=6.795 $Y=1.12 $X2=0
+ $Y2=0
cc_514 N_A_398_74#_M1014_g N_VGND_c_1699_n 0.00461464f $X=3.83 $Y=0.58 $X2=0
+ $Y2=0
cc_515 N_A_398_74#_c_317_n N_VGND_c_1699_n 0.0586507f $X=2.945 $Y=0.34 $X2=0
+ $Y2=0
cc_516 N_A_398_74#_c_318_n N_VGND_c_1699_n 0.0121867f $X=2.215 $Y=0.34 $X2=0
+ $Y2=0
cc_517 N_A_398_74#_c_323_n N_VGND_c_1701_n 0.0604764f $X=7.49 $Y=0.365 $X2=0
+ $Y2=0
cc_518 N_A_398_74#_c_324_n N_VGND_c_1701_n 0.0105206f $X=6.585 $Y=0.365 $X2=0
+ $Y2=0
cc_519 N_A_398_74#_c_329_n N_VGND_c_1701_n 0.00281891f $X=6.795 $Y=1.12 $X2=0
+ $Y2=0
cc_520 N_A_398_74#_M1014_g N_VGND_c_1709_n 0.00911847f $X=3.83 $Y=0.58 $X2=0
+ $Y2=0
cc_521 N_A_398_74#_c_317_n N_VGND_c_1709_n 0.0333627f $X=2.945 $Y=0.34 $X2=0
+ $Y2=0
cc_522 N_A_398_74#_c_318_n N_VGND_c_1709_n 0.00660921f $X=2.215 $Y=0.34 $X2=0
+ $Y2=0
cc_523 N_A_398_74#_c_323_n N_VGND_c_1709_n 0.0393398f $X=7.49 $Y=0.365 $X2=0
+ $Y2=0
cc_524 N_A_398_74#_c_324_n N_VGND_c_1709_n 0.00652894f $X=6.585 $Y=0.365 $X2=0
+ $Y2=0
cc_525 N_A_398_74#_c_329_n N_VGND_c_1709_n 0.00358754f $X=6.795 $Y=1.12 $X2=0
+ $Y2=0
cc_526 N_A_398_74#_c_321_n A_1278_74# 0.00221695f $X=6.5 $Y=1.12 $X2=-0.19
+ $Y2=-0.245
cc_527 N_A_398_74#_c_325_n A_1489_118# 0.00846132f $X=7.575 $Y=1.98 $X2=-0.19
+ $Y2=-0.245
cc_528 N_A_767_384#_c_587_n N_A_612_74#_c_664_n 0.0216132f $X=5.085 $Y=1.905
+ $X2=0 $Y2=0
cc_529 N_A_767_384#_c_588_n N_A_612_74#_c_664_n 0.0127717f $X=4.395 $Y=1.905
+ $X2=0 $Y2=0
cc_530 N_A_767_384#_c_590_n N_A_612_74#_c_664_n 0.00210237f $X=5.217 $Y=2.32
+ $X2=0 $Y2=0
cc_531 N_A_767_384#_c_589_n N_A_612_74#_c_679_n 0.00484379f $X=5.265 $Y=2.52
+ $X2=0 $Y2=0
cc_532 N_A_767_384#_c_590_n N_A_612_74#_c_679_n 0.00785968f $X=5.217 $Y=2.32
+ $X2=0 $Y2=0
cc_533 N_A_767_384#_c_581_n N_A_612_74#_M1001_g 0.0137077f $X=4.575 $Y=1.065
+ $X2=0 $Y2=0
cc_534 N_A_767_384#_c_583_n N_A_612_74#_M1001_g 0.00740402f $X=4.485 $Y=1.065
+ $X2=0 $Y2=0
cc_535 N_A_767_384#_c_581_n N_A_612_74#_c_669_n 0.0144466f $X=4.575 $Y=1.065
+ $X2=0 $Y2=0
cc_536 N_A_767_384#_c_583_n N_A_612_74#_c_669_n 0.00990744f $X=4.485 $Y=1.065
+ $X2=0 $Y2=0
cc_537 N_A_767_384#_c_581_n N_A_612_74#_c_670_n 0.00147785f $X=4.575 $Y=1.065
+ $X2=0 $Y2=0
cc_538 N_A_767_384#_c_583_n N_A_612_74#_c_670_n 0.00411471f $X=4.485 $Y=1.065
+ $X2=0 $Y2=0
cc_539 N_A_767_384#_c_585_n N_A_612_74#_c_671_n 0.00298868f $X=4.23 $Y=1.995
+ $X2=0 $Y2=0
cc_540 N_A_767_384#_c_587_n N_A_612_74#_c_671_n 0.00206546f $X=5.085 $Y=1.905
+ $X2=0 $Y2=0
cc_541 N_A_767_384#_c_588_n N_A_612_74#_c_671_n 2.83197e-19 $X=4.395 $Y=1.905
+ $X2=0 $Y2=0
cc_542 N_A_767_384#_c_587_n N_A_612_74#_c_672_n 0.0146716f $X=5.085 $Y=1.905
+ $X2=0 $Y2=0
cc_543 N_A_767_384#_c_581_n N_A_612_74#_c_672_n 0.0178654f $X=4.575 $Y=1.065
+ $X2=0 $Y2=0
cc_544 N_A_767_384#_c_582_n N_A_612_74#_c_672_n 9.72701e-19 $X=4.395 $Y=1.74
+ $X2=0 $Y2=0
cc_545 N_A_767_384#_c_586_n N_A_612_74#_c_673_n 8.04382e-19 $X=3.925 $Y=1.995
+ $X2=0 $Y2=0
cc_546 N_A_767_384#_c_587_n N_A_612_74#_c_675_n 0.0633465f $X=5.085 $Y=1.905
+ $X2=0 $Y2=0
cc_547 N_A_767_384#_c_588_n N_A_612_74#_c_675_n 0.00165087f $X=4.395 $Y=1.905
+ $X2=0 $Y2=0
cc_548 N_A_767_384#_c_581_n N_A_612_74#_c_675_n 0.0347181f $X=4.575 $Y=1.065
+ $X2=0 $Y2=0
cc_549 N_A_767_384#_c_582_n N_A_612_74#_c_675_n 0.0118646f $X=4.395 $Y=1.74
+ $X2=0 $Y2=0
cc_550 N_A_767_384#_c_583_n N_A_612_74#_c_675_n 0.00436216f $X=4.485 $Y=1.065
+ $X2=0 $Y2=0
cc_551 N_A_767_384#_c_587_n N_A_612_74#_c_677_n 9.26944e-19 $X=5.085 $Y=1.905
+ $X2=0 $Y2=0
cc_552 N_A_767_384#_c_581_n N_A_612_74#_c_677_n 0.00500011f $X=4.575 $Y=1.065
+ $X2=0 $Y2=0
cc_553 N_A_767_384#_c_582_n N_A_612_74#_c_677_n 0.0127717f $X=4.395 $Y=1.74
+ $X2=0 $Y2=0
cc_554 N_A_767_384#_c_583_n N_A_612_74#_c_677_n 6.53703e-19 $X=4.485 $Y=1.065
+ $X2=0 $Y2=0
cc_555 N_A_767_384#_c_587_n N_SET_B_c_801_n 0.0020735f $X=5.085 $Y=1.905
+ $X2=-0.19 $Y2=-0.245
cc_556 N_A_767_384#_c_589_n N_SET_B_c_801_n 0.00131208f $X=5.265 $Y=2.52
+ $X2=-0.19 $Y2=-0.245
cc_557 N_A_767_384#_c_590_n N_SET_B_c_801_n 0.00409522f $X=5.217 $Y=2.32
+ $X2=-0.19 $Y2=-0.245
cc_558 N_A_767_384#_c_587_n N_SET_B_M1020_g 0.00127041f $X=5.085 $Y=1.905 $X2=0
+ $Y2=0
cc_559 N_A_767_384#_c_581_n N_SET_B_M1020_g 0.0013988f $X=4.575 $Y=1.065 $X2=0
+ $Y2=0
cc_560 N_A_767_384#_c_587_n N_SET_B_c_808_n 5.40656e-19 $X=5.085 $Y=1.905 $X2=0
+ $Y2=0
cc_561 N_A_767_384#_c_590_n N_SET_B_c_808_n 2.51551e-19 $X=5.217 $Y=2.32 $X2=0
+ $Y2=0
cc_562 N_A_767_384#_c_587_n N_SET_B_c_809_n 0.0245674f $X=5.085 $Y=1.905 $X2=0
+ $Y2=0
cc_563 N_A_767_384#_c_590_n N_SET_B_c_809_n 0.00614145f $X=5.217 $Y=2.32 $X2=0
+ $Y2=0
cc_564 N_A_767_384#_c_584_n N_A_225_74#_c_938_n 0.00222191f $X=3.925 $Y=2.205
+ $X2=0 $Y2=0
cc_565 N_A_767_384#_c_584_n N_A_225_74#_c_940_n 0.021981f $X=3.925 $Y=2.205
+ $X2=0 $Y2=0
cc_566 N_A_767_384#_c_586_n N_A_225_74#_c_940_n 0.00249025f $X=3.925 $Y=1.995
+ $X2=0 $Y2=0
cc_567 N_A_767_384#_c_584_n N_A_225_74#_c_941_n 0.00850438f $X=3.925 $Y=2.205
+ $X2=0 $Y2=0
cc_568 N_A_767_384#_c_584_n N_VPWR_c_1506_n 0.00602275f $X=3.925 $Y=2.205 $X2=0
+ $Y2=0
cc_569 N_A_767_384#_c_584_n N_VPWR_c_1496_n 9.51552e-19 $X=3.925 $Y=2.205 $X2=0
+ $Y2=0
cc_570 N_A_767_384#_c_580_n N_VGND_c_1693_n 0.0129647f $X=4.22 $Y=0.9 $X2=0
+ $Y2=0
cc_571 N_A_767_384#_c_581_n N_VGND_c_1693_n 0.0271148f $X=4.575 $Y=1.065 $X2=0
+ $Y2=0
cc_572 N_A_767_384#_c_583_n N_VGND_c_1693_n 0.00527761f $X=4.485 $Y=1.065 $X2=0
+ $Y2=0
cc_573 N_A_767_384#_c_581_n N_VGND_c_1694_n 0.015698f $X=4.575 $Y=1.065 $X2=0
+ $Y2=0
cc_574 N_A_767_384#_c_580_n N_VGND_c_1699_n 0.00383152f $X=4.22 $Y=0.9 $X2=0
+ $Y2=0
cc_575 N_A_767_384#_c_581_n N_VGND_c_1700_n 0.00880728f $X=4.575 $Y=1.065 $X2=0
+ $Y2=0
cc_576 N_A_767_384#_c_580_n N_VGND_c_1709_n 0.0075725f $X=4.22 $Y=0.9 $X2=0
+ $Y2=0
cc_577 N_A_767_384#_c_581_n N_VGND_c_1709_n 0.012195f $X=4.575 $Y=1.065 $X2=0
+ $Y2=0
cc_578 N_A_612_74#_c_664_n N_SET_B_c_801_n 0.0184979f $X=5.04 $Y=2.115 $X2=-0.19
+ $Y2=-0.245
cc_579 N_A_612_74#_c_679_n N_SET_B_c_801_n 0.00927723f $X=5.04 $Y=2.205
+ $X2=-0.19 $Y2=-0.245
cc_580 N_A_612_74#_c_666_n N_SET_B_c_801_n 0.0191623f $X=6.255 $Y=1.63 $X2=-0.19
+ $Y2=-0.245
cc_581 N_A_612_74#_c_676_n N_SET_B_c_801_n 0.00537596f $X=5.915 $Y=1.392
+ $X2=-0.19 $Y2=-0.245
cc_582 N_A_612_74#_c_664_n N_SET_B_M1020_g 0.00824355f $X=5.04 $Y=2.115 $X2=0
+ $Y2=0
cc_583 N_A_612_74#_M1001_g N_SET_B_M1020_g 0.0572199f $X=5.21 $Y=0.8 $X2=0 $Y2=0
cc_584 N_A_612_74#_c_666_n N_SET_B_M1020_g 0.025215f $X=6.255 $Y=1.63 $X2=0
+ $Y2=0
cc_585 N_A_612_74#_M1031_g N_SET_B_M1020_g 0.00913306f $X=6.315 $Y=0.69 $X2=0
+ $Y2=0
cc_586 N_A_612_74#_c_676_n N_SET_B_M1020_g 0.0211117f $X=5.915 $Y=1.392 $X2=0
+ $Y2=0
cc_587 N_A_612_74#_c_666_n N_SET_B_c_807_n 0.00991712f $X=6.255 $Y=1.63 $X2=0
+ $Y2=0
cc_588 N_A_612_74#_c_683_n N_SET_B_c_807_n 0.00338559f $X=6.08 $Y=1.38 $X2=0
+ $Y2=0
cc_589 N_A_612_74#_c_666_n N_SET_B_c_808_n 0.00164794f $X=6.255 $Y=1.63 $X2=0
+ $Y2=0
cc_590 N_A_612_74#_c_683_n N_SET_B_c_808_n 0.00128918f $X=6.08 $Y=1.38 $X2=0
+ $Y2=0
cc_591 N_A_612_74#_c_676_n N_SET_B_c_808_n 0.00154953f $X=5.915 $Y=1.392 $X2=0
+ $Y2=0
cc_592 N_A_612_74#_c_664_n N_SET_B_c_809_n 3.53369e-19 $X=5.04 $Y=2.115 $X2=0
+ $Y2=0
cc_593 N_A_612_74#_c_666_n N_SET_B_c_809_n 0.00524035f $X=6.255 $Y=1.63 $X2=0
+ $Y2=0
cc_594 N_A_612_74#_c_676_n N_SET_B_c_809_n 0.0443631f $X=5.915 $Y=1.392 $X2=0
+ $Y2=0
cc_595 N_A_612_74#_c_674_n N_A_225_74#_c_923_n 4.37445e-19 $X=3.45 $Y=1.125
+ $X2=0 $Y2=0
cc_596 N_A_612_74#_c_668_n N_A_225_74#_M1019_g 0.00255027f $X=3.45 $Y=0.585
+ $X2=0 $Y2=0
cc_597 N_A_612_74#_c_681_n N_A_225_74#_c_938_n 4.27465e-19 $X=3.28 $Y=2.49 $X2=0
+ $Y2=0
cc_598 N_A_612_74#_c_681_n N_A_225_74#_c_940_n 0.00583751f $X=3.28 $Y=2.49 $X2=0
+ $Y2=0
cc_599 N_A_612_74#_c_673_n N_A_225_74#_c_940_n 0.00245035f $X=3.285 $Y=2.26
+ $X2=0 $Y2=0
cc_600 N_A_612_74#_c_679_n N_A_225_74#_c_941_n 0.00716579f $X=5.04 $Y=2.205
+ $X2=0 $Y2=0
cc_601 N_A_612_74#_c_666_n N_A_225_74#_c_941_n 0.00862445f $X=6.255 $Y=1.63
+ $X2=0 $Y2=0
cc_602 N_A_612_74#_c_666_n N_A_225_74#_M1006_g 0.0292179f $X=6.255 $Y=1.63 $X2=0
+ $Y2=0
cc_603 N_A_612_74#_c_666_n N_A_225_74#_c_927_n 0.00651444f $X=6.255 $Y=1.63
+ $X2=0 $Y2=0
cc_604 N_A_612_74#_c_666_n N_A_1356_74#_c_1213_n 6.29517e-19 $X=6.255 $Y=1.63
+ $X2=0 $Y2=0
cc_605 N_A_612_74#_c_666_n N_A_1356_74#_c_1220_n 0.00130593f $X=6.255 $Y=1.63
+ $X2=0 $Y2=0
cc_606 N_A_612_74#_c_681_n N_A_27_74#_c_1432_n 0.0200861f $X=3.28 $Y=2.49 $X2=0
+ $Y2=0
cc_607 N_A_612_74#_c_673_n N_A_27_74#_c_1432_n 0.00626921f $X=3.285 $Y=2.26
+ $X2=0 $Y2=0
cc_608 N_A_612_74#_c_673_n N_A_27_74#_c_1426_n 2.70958e-19 $X=3.285 $Y=2.26
+ $X2=0 $Y2=0
cc_609 N_A_612_74#_c_666_n N_VPWR_c_1500_n 0.0051214f $X=6.255 $Y=1.63 $X2=0
+ $Y2=0
cc_610 N_A_612_74#_c_666_n N_VPWR_c_1496_n 9.49986e-19 $X=6.255 $Y=1.63 $X2=0
+ $Y2=0
cc_611 N_A_612_74#_M1001_g N_VGND_c_1693_n 0.00304548f $X=5.21 $Y=0.8 $X2=0
+ $Y2=0
cc_612 N_A_612_74#_c_668_n N_VGND_c_1693_n 0.00823525f $X=3.45 $Y=0.585 $X2=0
+ $Y2=0
cc_613 N_A_612_74#_M1001_g N_VGND_c_1694_n 0.00183638f $X=5.21 $Y=0.8 $X2=0
+ $Y2=0
cc_614 N_A_612_74#_c_666_n N_VGND_c_1694_n 0.00776361f $X=6.255 $Y=1.63 $X2=0
+ $Y2=0
cc_615 N_A_612_74#_M1031_g N_VGND_c_1694_n 0.0162104f $X=6.315 $Y=0.69 $X2=0
+ $Y2=0
cc_616 N_A_612_74#_c_683_n N_VGND_c_1694_n 0.0261475f $X=6.08 $Y=1.38 $X2=0
+ $Y2=0
cc_617 N_A_612_74#_c_676_n N_VGND_c_1694_n 0.021427f $X=5.915 $Y=1.392 $X2=0
+ $Y2=0
cc_618 N_A_612_74#_c_668_n N_VGND_c_1699_n 0.0118117f $X=3.45 $Y=0.585 $X2=0
+ $Y2=0
cc_619 N_A_612_74#_M1001_g N_VGND_c_1700_n 0.00416964f $X=5.21 $Y=0.8 $X2=0
+ $Y2=0
cc_620 N_A_612_74#_M1031_g N_VGND_c_1701_n 0.00444681f $X=6.315 $Y=0.69 $X2=0
+ $Y2=0
cc_621 N_A_612_74#_M1001_g N_VGND_c_1709_n 0.00479212f $X=5.21 $Y=0.8 $X2=0
+ $Y2=0
cc_622 N_A_612_74#_M1031_g N_VGND_c_1709_n 0.00877228f $X=6.315 $Y=0.69 $X2=0
+ $Y2=0
cc_623 N_A_612_74#_c_668_n N_VGND_c_1709_n 0.011742f $X=3.45 $Y=0.585 $X2=0
+ $Y2=0
cc_624 N_SET_B_c_801_n N_A_225_74#_c_941_n 0.00718133f $X=5.49 $Y=2.205 $X2=0
+ $Y2=0
cc_625 N_SET_B_c_807_n N_A_225_74#_M1006_g 0.00851485f $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_626 N_SET_B_c_807_n N_A_225_74#_c_926_n 0.00682877f $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_627 N_SET_B_c_807_n N_A_225_74#_c_927_n 3.57752e-19 $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_628 N_SET_B_c_806_n N_A_1566_92#_c_1122_n 0.00614889f $X=8.565 $Y=2.15 $X2=0
+ $Y2=0
cc_629 SET_B N_A_1566_92#_c_1122_n 3.05387e-19 $X=8.315 $Y=1.95 $X2=0 $Y2=0
cc_630 N_SET_B_c_803_n N_A_1566_92#_c_1123_n 0.00614889f $X=8.49 $Y=2.375 $X2=0
+ $Y2=0
cc_631 N_SET_B_c_804_n N_A_1566_92#_c_1123_n 0.0115888f $X=8.49 $Y=2.465 $X2=0
+ $Y2=0
cc_632 N_SET_B_M1002_g N_A_1566_92#_c_1114_n 0.0205048f $X=8.475 $Y=0.8 $X2=0
+ $Y2=0
cc_633 N_SET_B_M1002_g N_A_1566_92#_c_1124_n 0.00149238f $X=8.475 $Y=0.8 $X2=0
+ $Y2=0
cc_634 N_SET_B_c_807_n N_A_1566_92#_c_1124_n 0.027726f $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_635 SET_B N_A_1566_92#_c_1124_n 0.00213174f $X=8.315 $Y=1.95 $X2=0 $Y2=0
cc_636 N_SET_B_c_799_n N_A_1566_92#_c_1124_n 7.54692e-19 $X=8.565 $Y=1.645 $X2=0
+ $Y2=0
cc_637 N_SET_B_c_800_n N_A_1566_92#_c_1124_n 0.0495655f $X=8.565 $Y=1.645 $X2=0
+ $Y2=0
cc_638 N_SET_B_M1002_g N_A_1566_92#_c_1115_n 0.0182739f $X=8.475 $Y=0.8 $X2=0
+ $Y2=0
cc_639 SET_B N_A_1566_92#_c_1116_n 7.33174e-19 $X=8.315 $Y=1.95 $X2=0 $Y2=0
cc_640 N_SET_B_c_799_n N_A_1566_92#_c_1116_n 0.0182739f $X=8.565 $Y=1.645 $X2=0
+ $Y2=0
cc_641 N_SET_B_c_800_n N_A_1566_92#_c_1116_n 0.0038385f $X=8.565 $Y=1.645 $X2=0
+ $Y2=0
cc_642 N_SET_B_M1002_g N_A_1566_92#_c_1117_n 0.0165527f $X=8.475 $Y=0.8 $X2=0
+ $Y2=0
cc_643 N_SET_B_c_799_n N_A_1566_92#_c_1117_n 0.00116081f $X=8.565 $Y=1.645 $X2=0
+ $Y2=0
cc_644 N_SET_B_c_800_n N_A_1566_92#_c_1117_n 0.0252292f $X=8.565 $Y=1.645 $X2=0
+ $Y2=0
cc_645 N_SET_B_c_798_n N_A_1566_92#_c_1127_n 0.0182739f $X=8.565 $Y=1.985 $X2=0
+ $Y2=0
cc_646 N_SET_B_c_807_n N_A_1566_92#_c_1127_n 0.00323607f $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_647 SET_B N_A_1566_92#_c_1127_n 4.08782e-19 $X=8.315 $Y=1.95 $X2=0 $Y2=0
cc_648 N_SET_B_c_807_n N_A_1356_74#_M1006_d 0.00115767f $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_649 N_SET_B_c_799_n N_A_1356_74#_M1024_g 0.00259971f $X=8.565 $Y=1.645 $X2=0
+ $Y2=0
cc_650 N_SET_B_c_800_n N_A_1356_74#_M1024_g 6.32828e-19 $X=8.565 $Y=1.645 $X2=0
+ $Y2=0
cc_651 N_SET_B_c_799_n N_A_1356_74#_c_1202_n 0.00494777f $X=8.565 $Y=1.645 $X2=0
+ $Y2=0
cc_652 N_SET_B_c_800_n N_A_1356_74#_c_1202_n 0.0024583f $X=8.565 $Y=1.645 $X2=0
+ $Y2=0
cc_653 N_SET_B_c_803_n N_A_1356_74#_c_1211_n 0.00328286f $X=8.49 $Y=2.375 $X2=0
+ $Y2=0
cc_654 N_SET_B_c_806_n N_A_1356_74#_c_1211_n 0.00494777f $X=8.565 $Y=2.15 $X2=0
+ $Y2=0
cc_655 N_SET_B_c_807_n N_A_1356_74#_c_1213_n 0.0144054f $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_656 N_SET_B_c_807_n N_A_1356_74#_c_1233_n 0.00350245f $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_657 N_SET_B_c_803_n N_A_1356_74#_c_1214_n 0.00534918f $X=8.49 $Y=2.375 $X2=0
+ $Y2=0
cc_658 N_SET_B_c_804_n N_A_1356_74#_c_1214_n 0.0129101f $X=8.49 $Y=2.465 $X2=0
+ $Y2=0
cc_659 N_SET_B_c_806_n N_A_1356_74#_c_1214_n 3.53728e-19 $X=8.565 $Y=2.15 $X2=0
+ $Y2=0
cc_660 N_SET_B_c_807_n N_A_1356_74#_c_1214_n 0.00640638f $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_661 SET_B N_A_1356_74#_c_1214_n 0.00471918f $X=8.315 $Y=1.95 $X2=0 $Y2=0
cc_662 N_SET_B_c_800_n N_A_1356_74#_c_1214_n 0.0215664f $X=8.565 $Y=1.645 $X2=0
+ $Y2=0
cc_663 N_SET_B_c_804_n N_A_1356_74#_c_1215_n 6.15967e-19 $X=8.49 $Y=2.465 $X2=0
+ $Y2=0
cc_664 N_SET_B_c_807_n N_A_1356_74#_c_1215_n 0.00403539f $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_665 N_SET_B_c_804_n N_A_1356_74#_c_1216_n 0.00524508f $X=8.49 $Y=2.465 $X2=0
+ $Y2=0
cc_666 N_SET_B_c_803_n N_A_1356_74#_c_1205_n 0.00157501f $X=8.49 $Y=2.375 $X2=0
+ $Y2=0
cc_667 SET_B N_A_1356_74#_c_1205_n 0.00107107f $X=8.315 $Y=1.95 $X2=0 $Y2=0
cc_668 N_SET_B_c_799_n N_A_1356_74#_c_1205_n 0.00225352f $X=8.565 $Y=1.645 $X2=0
+ $Y2=0
cc_669 N_SET_B_c_800_n N_A_1356_74#_c_1205_n 0.018807f $X=8.565 $Y=1.645 $X2=0
+ $Y2=0
cc_670 N_SET_B_c_798_n N_A_1356_74#_c_1219_n 0.00494777f $X=8.565 $Y=1.985 $X2=0
+ $Y2=0
cc_671 N_SET_B_c_807_n N_A_1356_74#_c_1206_n 0.0111047f $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_672 N_SET_B_c_807_n N_A_1356_74#_c_1220_n 0.0108359f $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_673 N_SET_B_c_806_n N_A_1356_74#_c_1221_n 7.69224e-19 $X=8.565 $Y=2.15 $X2=0
+ $Y2=0
cc_674 N_SET_B_c_800_n N_A_1356_74#_c_1221_n 0.00879631f $X=8.565 $Y=1.645 $X2=0
+ $Y2=0
cc_675 N_SET_B_c_807_n N_VPWR_M1008_d 6.35591e-19 $X=8.255 $Y=2.035 $X2=0 $Y2=0
cc_676 N_SET_B_c_808_n N_VPWR_M1008_d 0.00306855f $X=6.145 $Y=2.035 $X2=0 $Y2=0
cc_677 N_SET_B_c_809_n N_VPWR_M1008_d 0.00961121f $X=6 $Y=2.035 $X2=0 $Y2=0
cc_678 N_SET_B_c_801_n N_VPWR_c_1500_n 5.2853e-19 $X=5.49 $Y=2.205 $X2=0 $Y2=0
cc_679 N_SET_B_c_804_n N_VPWR_c_1501_n 0.00951807f $X=8.49 $Y=2.465 $X2=0 $Y2=0
cc_680 N_SET_B_c_804_n N_VPWR_c_1502_n 0.00325258f $X=8.49 $Y=2.465 $X2=0 $Y2=0
cc_681 N_SET_B_c_804_n N_VPWR_c_1513_n 0.00413917f $X=8.49 $Y=2.465 $X2=0 $Y2=0
cc_682 N_SET_B_c_804_n N_VPWR_c_1496_n 0.00405713f $X=8.49 $Y=2.465 $X2=0 $Y2=0
cc_683 N_SET_B_c_807_n A_1266_341# 0.00775606f $X=8.255 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_684 N_SET_B_M1020_g N_VGND_c_1694_n 0.0149224f $X=5.6 $Y=0.8 $X2=0 $Y2=0
cc_685 N_SET_B_M1020_g N_VGND_c_1700_n 0.00360926f $X=5.6 $Y=0.8 $X2=0 $Y2=0
cc_686 N_SET_B_M1002_g N_VGND_c_1701_n 0.0172888f $X=8.475 $Y=0.8 $X2=0 $Y2=0
cc_687 N_SET_B_M1020_g N_VGND_c_1709_n 0.00402538f $X=5.6 $Y=0.8 $X2=0 $Y2=0
cc_688 N_SET_B_M1002_g N_VGND_c_1709_n 0.00402538f $X=8.475 $Y=0.8 $X2=0 $Y2=0
cc_689 N_A_225_74#_M1009_g N_A_1566_92#_c_1114_n 0.0158751f $X=7.37 $Y=0.8 $X2=0
+ $Y2=0
cc_690 N_A_225_74#_c_926_n N_A_1566_92#_c_1115_n 0.0158751f $X=7.295 $Y=1.735
+ $X2=0 $Y2=0
cc_691 N_A_225_74#_M1006_g N_A_1356_74#_c_1213_n 0.00895465f $X=6.76 $Y=2.46
+ $X2=0 $Y2=0
cc_692 N_A_225_74#_c_926_n N_A_1356_74#_c_1213_n 0.00672058f $X=7.295 $Y=1.735
+ $X2=0 $Y2=0
cc_693 N_A_225_74#_c_927_n N_A_1356_74#_c_1213_n 0.00307469f $X=6.85 $Y=1.735
+ $X2=0 $Y2=0
cc_694 N_A_225_74#_c_926_n N_A_1356_74#_c_1204_n 0.0015047f $X=7.295 $Y=1.735
+ $X2=0 $Y2=0
cc_695 N_A_225_74#_M1009_g N_A_1356_74#_c_1204_n 0.0149235f $X=7.37 $Y=0.8 $X2=0
+ $Y2=0
cc_696 N_A_225_74#_c_926_n N_A_1356_74#_c_1206_n 0.0155989f $X=7.295 $Y=1.735
+ $X2=0 $Y2=0
cc_697 N_A_225_74#_c_927_n N_A_1356_74#_c_1206_n 0.00183668f $X=6.85 $Y=1.735
+ $X2=0 $Y2=0
cc_698 N_A_225_74#_M1009_g N_A_1356_74#_c_1206_n 0.00131824f $X=7.37 $Y=0.8
+ $X2=0 $Y2=0
cc_699 N_A_225_74#_c_941_n N_A_1356_74#_c_1220_n 3.80133e-19 $X=6.67 $Y=3.15
+ $X2=0 $Y2=0
cc_700 N_A_225_74#_M1006_g N_A_1356_74#_c_1220_n 0.0172017f $X=6.76 $Y=2.46
+ $X2=0 $Y2=0
cc_701 N_A_225_74#_M1009_g N_A_1356_74#_c_1243_n 0.00926501f $X=7.37 $Y=0.8
+ $X2=0 $Y2=0
cc_702 N_A_225_74#_M1028_s N_A_27_74#_c_1431_n 0.0126187f $X=1.145 $Y=1.79 $X2=0
+ $Y2=0
cc_703 N_A_225_74#_c_949_n N_A_27_74#_c_1431_n 0.0190006f $X=1.305 $Y=1.87 $X2=0
+ $Y2=0
cc_704 N_A_225_74#_c_950_n N_A_27_74#_c_1431_n 0.0142272f $X=1.145 $Y=1.87 $X2=0
+ $Y2=0
cc_705 N_A_225_74#_c_951_n N_A_27_74#_c_1431_n 0.0057885f $X=1.945 $Y=1.805
+ $X2=0 $Y2=0
cc_706 N_A_225_74#_c_921_n N_A_27_74#_c_1432_n 0.014987f $X=1.965 $Y=1.715 $X2=0
+ $Y2=0
cc_707 N_A_225_74#_c_935_n N_A_27_74#_c_1432_n 0.0265478f $X=2.485 $Y=3.075
+ $X2=0 $Y2=0
cc_708 N_A_225_74#_c_929_n N_A_27_74#_c_1432_n 0.00492213f $X=2.41 $Y=1.465
+ $X2=0 $Y2=0
cc_709 N_A_225_74#_c_951_n N_A_27_74#_c_1432_n 0.0278803f $X=1.945 $Y=1.805
+ $X2=0 $Y2=0
cc_710 N_A_225_74#_M1016_g N_A_27_74#_c_1426_n 7.54241e-19 $X=1.915 $Y=0.74
+ $X2=0 $Y2=0
cc_711 N_A_225_74#_c_921_n N_A_27_74#_c_1426_n 0.00116731f $X=1.965 $Y=1.715
+ $X2=0 $Y2=0
cc_712 N_A_225_74#_c_922_n N_A_27_74#_c_1426_n 0.00518646f $X=2.485 $Y=1.3 $X2=0
+ $Y2=0
cc_713 N_A_225_74#_c_935_n N_A_27_74#_c_1426_n 0.00991345f $X=2.485 $Y=3.075
+ $X2=0 $Y2=0
cc_714 N_A_225_74#_c_923_n N_A_27_74#_c_1426_n 0.00578804f $X=2.91 $Y=1.065
+ $X2=0 $Y2=0
cc_715 N_A_225_74#_c_924_n N_A_27_74#_c_1426_n 0.00450019f $X=2.56 $Y=1.065
+ $X2=0 $Y2=0
cc_716 N_A_225_74#_M1019_g N_A_27_74#_c_1426_n 0.00115087f $X=2.985 $Y=0.58
+ $X2=0 $Y2=0
cc_717 N_A_225_74#_c_930_n N_A_27_74#_c_1426_n 0.0101071f $X=2.485 $Y=1.465
+ $X2=0 $Y2=0
cc_718 N_A_225_74#_c_951_n N_A_27_74#_c_1426_n 0.0135406f $X=1.945 $Y=1.805
+ $X2=0 $Y2=0
cc_719 N_A_225_74#_c_932_n N_A_27_74#_c_1426_n 0.0302859f $X=2.11 $Y=1.465 $X2=0
+ $Y2=0
cc_720 N_A_225_74#_c_921_n N_A_27_74#_c_1480_n 0.00185704f $X=1.965 $Y=1.715
+ $X2=0 $Y2=0
cc_721 N_A_225_74#_c_951_n N_A_27_74#_c_1480_n 0.0112057f $X=1.945 $Y=1.805
+ $X2=0 $Y2=0
cc_722 N_A_225_74#_c_923_n N_A_27_74#_c_1428_n 0.00669646f $X=2.91 $Y=1.065
+ $X2=0 $Y2=0
cc_723 N_A_225_74#_c_924_n N_A_27_74#_c_1428_n 0.00134438f $X=2.56 $Y=1.065
+ $X2=0 $Y2=0
cc_724 N_A_225_74#_M1019_g N_A_27_74#_c_1428_n 0.0066603f $X=2.985 $Y=0.58 $X2=0
+ $Y2=0
cc_725 N_A_225_74#_c_951_n N_VPWR_M1028_d 0.00196757f $X=1.945 $Y=1.805 $X2=0
+ $Y2=0
cc_726 N_A_225_74#_c_921_n N_VPWR_c_1498_n 0.00746756f $X=1.965 $Y=1.715 $X2=0
+ $Y2=0
cc_727 N_A_225_74#_c_935_n N_VPWR_c_1498_n 0.00346889f $X=2.485 $Y=3.075 $X2=0
+ $Y2=0
cc_728 N_A_225_74#_c_939_n N_VPWR_c_1499_n 0.00103154f $X=3.505 $Y=3.075 $X2=0
+ $Y2=0
cc_729 N_A_225_74#_c_941_n N_VPWR_c_1499_n 0.0160168f $X=6.67 $Y=3.15 $X2=0
+ $Y2=0
cc_730 N_A_225_74#_c_941_n N_VPWR_c_1500_n 0.0220021f $X=6.67 $Y=3.15 $X2=0
+ $Y2=0
cc_731 N_A_225_74#_M1006_g N_VPWR_c_1500_n 0.00504437f $X=6.76 $Y=2.46 $X2=0
+ $Y2=0
cc_732 N_A_225_74#_c_939_n N_VPWR_c_1506_n 2.53362e-19 $X=3.505 $Y=3.075 $X2=0
+ $Y2=0
cc_733 N_A_225_74#_c_941_n N_VPWR_c_1506_n 0.00817058f $X=6.67 $Y=3.15 $X2=0
+ $Y2=0
cc_734 N_A_225_74#_c_941_n N_VPWR_c_1507_n 0.0262434f $X=6.67 $Y=3.15 $X2=0
+ $Y2=0
cc_735 N_A_225_74#_c_921_n N_VPWR_c_1511_n 0.0048608f $X=1.965 $Y=1.715 $X2=0
+ $Y2=0
cc_736 N_A_225_74#_c_937_n N_VPWR_c_1511_n 0.0396626f $X=2.56 $Y=3.15 $X2=0
+ $Y2=0
cc_737 N_A_225_74#_c_941_n N_VPWR_c_1512_n 0.0386563f $X=6.67 $Y=3.15 $X2=0
+ $Y2=0
cc_738 N_A_225_74#_c_921_n N_VPWR_c_1496_n 0.00480464f $X=1.965 $Y=1.715 $X2=0
+ $Y2=0
cc_739 N_A_225_74#_c_936_n N_VPWR_c_1496_n 0.0201442f $X=3.415 $Y=3.15 $X2=0
+ $Y2=0
cc_740 N_A_225_74#_c_937_n N_VPWR_c_1496_n 0.00604809f $X=2.56 $Y=3.15 $X2=0
+ $Y2=0
cc_741 N_A_225_74#_c_941_n N_VPWR_c_1496_n 0.0906242f $X=6.67 $Y=3.15 $X2=0
+ $Y2=0
cc_742 N_A_225_74#_c_947_n N_VPWR_c_1496_n 0.00441963f $X=3.505 $Y=3.15 $X2=0
+ $Y2=0
cc_743 N_A_225_74#_c_933_n N_VGND_c_1690_n 0.0327823f $X=1.27 $Y=0.51 $X2=0
+ $Y2=0
cc_744 N_A_225_74#_c_933_n N_VGND_c_1691_n 0.0203368f $X=1.27 $Y=0.51 $X2=0
+ $Y2=0
cc_745 N_A_225_74#_M1016_g N_VGND_c_1692_n 0.0115598f $X=1.915 $Y=0.74 $X2=0
+ $Y2=0
cc_746 N_A_225_74#_c_933_n N_VGND_c_1692_n 0.0256161f $X=1.27 $Y=0.51 $X2=0
+ $Y2=0
cc_747 N_A_225_74#_M1016_g N_VGND_c_1699_n 0.00383152f $X=1.915 $Y=0.74 $X2=0
+ $Y2=0
cc_748 N_A_225_74#_M1019_g N_VGND_c_1699_n 0.00278159f $X=2.985 $Y=0.58 $X2=0
+ $Y2=0
cc_749 N_A_225_74#_M1016_g N_VGND_c_1709_n 0.00762539f $X=1.915 $Y=0.74 $X2=0
+ $Y2=0
cc_750 N_A_225_74#_M1019_g N_VGND_c_1709_n 0.00361237f $X=2.985 $Y=0.58 $X2=0
+ $Y2=0
cc_751 N_A_225_74#_c_933_n N_VGND_c_1709_n 0.0167889f $X=1.27 $Y=0.51 $X2=0
+ $Y2=0
cc_752 N_A_1566_92#_c_1117_n N_A_1356_74#_M1024_g 0.0152849f $X=9.53 $Y=1.155
+ $X2=0 $Y2=0
cc_753 N_A_1566_92#_c_1119_n N_A_1356_74#_M1024_g 0.0121665f $X=9.695 $Y=0.8
+ $X2=0 $Y2=0
cc_754 N_A_1566_92#_c_1120_n N_A_1356_74#_M1024_g 0.0147061f $X=9.725 $Y=2.75
+ $X2=0 $Y2=0
cc_755 N_A_1566_92#_c_1121_n N_A_1356_74#_M1024_g 0.00513932f $X=9.71 $Y=1.155
+ $X2=0 $Y2=0
cc_756 N_A_1566_92#_c_1120_n N_A_1356_74#_c_1207_n 0.00713854f $X=9.725 $Y=2.75
+ $X2=0 $Y2=0
cc_757 N_A_1566_92#_c_1120_n N_A_1356_74#_c_1200_n 0.0188128f $X=9.725 $Y=2.75
+ $X2=0 $Y2=0
cc_758 N_A_1566_92#_c_1120_n N_A_1356_74#_M1015_g 0.0014319f $X=9.725 $Y=2.75
+ $X2=0 $Y2=0
cc_759 N_A_1566_92#_c_1121_n N_A_1356_74#_M1015_g 6.25308e-19 $X=9.71 $Y=1.155
+ $X2=0 $Y2=0
cc_760 N_A_1566_92#_c_1120_n N_A_1356_74#_c_1209_n 0.00440805f $X=9.725 $Y=2.75
+ $X2=0 $Y2=0
cc_761 N_A_1566_92#_c_1117_n N_A_1356_74#_c_1202_n 0.00155183f $X=9.53 $Y=1.155
+ $X2=0 $Y2=0
cc_762 N_A_1566_92#_c_1123_n N_A_1356_74#_c_1233_n 2.25853e-19 $X=7.95 $Y=2.465
+ $X2=0 $Y2=0
cc_763 N_A_1566_92#_c_1122_n N_A_1356_74#_c_1214_n 0.00301856f $X=7.95 $Y=2.375
+ $X2=0 $Y2=0
cc_764 N_A_1566_92#_c_1123_n N_A_1356_74#_c_1214_n 0.00709151f $X=7.95 $Y=2.465
+ $X2=0 $Y2=0
cc_765 N_A_1566_92#_c_1124_n N_A_1356_74#_c_1214_n 0.0141202f $X=7.995 $Y=1.285
+ $X2=0 $Y2=0
cc_766 N_A_1566_92#_c_1127_n N_A_1356_74#_c_1214_n 0.00139354f $X=7.995 $Y=2.13
+ $X2=0 $Y2=0
cc_767 N_A_1566_92#_c_1122_n N_A_1356_74#_c_1215_n 0.0017867f $X=7.95 $Y=2.375
+ $X2=0 $Y2=0
cc_768 N_A_1566_92#_c_1123_n N_A_1356_74#_c_1215_n 0.00872981f $X=7.95 $Y=2.465
+ $X2=0 $Y2=0
cc_769 N_A_1566_92#_c_1124_n N_A_1356_74#_c_1215_n 0.00668502f $X=7.995 $Y=1.285
+ $X2=0 $Y2=0
cc_770 N_A_1566_92#_c_1127_n N_A_1356_74#_c_1215_n 2.12417e-19 $X=7.995 $Y=2.13
+ $X2=0 $Y2=0
cc_771 N_A_1566_92#_c_1120_n N_A_1356_74#_c_1217_n 0.0139292f $X=9.725 $Y=2.75
+ $X2=0 $Y2=0
cc_772 N_A_1566_92#_c_1117_n N_A_1356_74#_c_1205_n 0.0142071f $X=9.53 $Y=1.155
+ $X2=0 $Y2=0
cc_773 N_A_1566_92#_c_1120_n N_A_1356_74#_c_1205_n 0.0538751f $X=9.725 $Y=2.75
+ $X2=0 $Y2=0
cc_774 N_A_1566_92#_c_1120_n N_A_1356_74#_c_1219_n 0.0185789f $X=9.725 $Y=2.75
+ $X2=0 $Y2=0
cc_775 N_A_1566_92#_c_1123_n N_A_1356_74#_c_1220_n 7.42617e-19 $X=7.95 $Y=2.465
+ $X2=0 $Y2=0
cc_776 N_A_1566_92#_c_1119_n N_A_2022_94#_c_1359_n 0.0324928f $X=9.695 $Y=0.8
+ $X2=0 $Y2=0
cc_777 N_A_1566_92#_c_1120_n N_A_2022_94#_c_1359_n 0.00429293f $X=9.725 $Y=2.75
+ $X2=0 $Y2=0
cc_778 N_A_1566_92#_c_1121_n N_A_2022_94#_c_1359_n 0.0134078f $X=9.71 $Y=1.155
+ $X2=0 $Y2=0
cc_779 N_A_1566_92#_c_1120_n N_A_2022_94#_c_1365_n 0.088949f $X=9.725 $Y=2.75
+ $X2=0 $Y2=0
cc_780 N_A_1566_92#_c_1120_n N_A_2022_94#_c_1361_n 0.0253904f $X=9.725 $Y=2.75
+ $X2=0 $Y2=0
cc_781 N_A_1566_92#_c_1123_n N_VPWR_c_1501_n 0.00682814f $X=7.95 $Y=2.465 $X2=0
+ $Y2=0
cc_782 N_A_1566_92#_c_1120_n N_VPWR_c_1502_n 0.0214859f $X=9.725 $Y=2.75 $X2=0
+ $Y2=0
cc_783 N_A_1566_92#_c_1123_n N_VPWR_c_1507_n 0.00411349f $X=7.95 $Y=2.465 $X2=0
+ $Y2=0
cc_784 N_A_1566_92#_c_1120_n N_VPWR_c_1514_n 0.011066f $X=9.725 $Y=2.75 $X2=0
+ $Y2=0
cc_785 N_A_1566_92#_c_1123_n N_VPWR_c_1496_n 0.00432531f $X=7.95 $Y=2.465 $X2=0
+ $Y2=0
cc_786 N_A_1566_92#_c_1120_n N_VPWR_c_1496_n 0.00915947f $X=9.725 $Y=2.75 $X2=0
+ $Y2=0
cc_787 N_A_1566_92#_c_1114_n N_VGND_c_1701_n 0.00633226f $X=7.995 $Y=1.12 $X2=0
+ $Y2=0
cc_788 N_A_1566_92#_c_1117_n N_VGND_c_1701_n 0.0656301f $X=9.53 $Y=1.155 $X2=0
+ $Y2=0
cc_789 N_A_1566_92#_c_1119_n N_VGND_c_1702_n 0.00636076f $X=9.695 $Y=0.8 $X2=0
+ $Y2=0
cc_790 N_A_1566_92#_c_1114_n N_VGND_c_1709_n 0.00479212f $X=7.995 $Y=1.12 $X2=0
+ $Y2=0
cc_791 N_A_1566_92#_c_1119_n N_VGND_c_1709_n 0.010804f $X=9.695 $Y=0.8 $X2=0
+ $Y2=0
cc_792 N_A_1356_74#_c_1209_n N_A_2022_94#_c_1363_n 0.0210645f $X=10.51 $Y=1.765
+ $X2=0 $Y2=0
cc_793 N_A_1356_74#_M1015_g N_A_2022_94#_M1003_g 0.0194305f $X=10.47 $Y=0.79
+ $X2=0 $Y2=0
cc_794 N_A_1356_74#_M1024_g N_A_2022_94#_c_1359_n 0.00555362f $X=9.48 $Y=0.8
+ $X2=0 $Y2=0
cc_795 N_A_1356_74#_M1015_g N_A_2022_94#_c_1359_n 0.0151436f $X=10.47 $Y=0.79
+ $X2=0 $Y2=0
cc_796 N_A_1356_74#_c_1200_n N_A_2022_94#_c_1365_n 0.0120472f $X=10.395 $Y=1.69
+ $X2=0 $Y2=0
cc_797 N_A_1356_74#_c_1209_n N_A_2022_94#_c_1365_n 0.0157206f $X=10.51 $Y=1.765
+ $X2=0 $Y2=0
cc_798 N_A_1356_74#_c_1203_n N_A_2022_94#_c_1365_n 0.00308043f $X=10.497 $Y=1.69
+ $X2=0 $Y2=0
cc_799 N_A_1356_74#_M1015_g N_A_2022_94#_c_1360_n 0.0107422f $X=10.47 $Y=0.79
+ $X2=0 $Y2=0
cc_800 N_A_1356_74#_c_1203_n N_A_2022_94#_c_1360_n 0.0084622f $X=10.497 $Y=1.69
+ $X2=0 $Y2=0
cc_801 N_A_1356_74#_c_1200_n N_A_2022_94#_c_1361_n 0.00584559f $X=10.395 $Y=1.69
+ $X2=0 $Y2=0
cc_802 N_A_1356_74#_M1015_g N_A_2022_94#_c_1361_n 0.00952755f $X=10.47 $Y=0.79
+ $X2=0 $Y2=0
cc_803 N_A_1356_74#_M1015_g N_A_2022_94#_c_1362_n 0.0153086f $X=10.47 $Y=0.79
+ $X2=0 $Y2=0
cc_804 N_A_1356_74#_c_1203_n N_A_2022_94#_c_1362_n 0.00603519f $X=10.497 $Y=1.69
+ $X2=0 $Y2=0
cc_805 N_A_1356_74#_c_1214_n N_VPWR_M1012_d 0.00308164f $X=8.63 $Y=2.435 $X2=0
+ $Y2=0
cc_806 N_A_1356_74#_c_1214_n N_VPWR_c_1501_n 0.0212032f $X=8.63 $Y=2.435 $X2=0
+ $Y2=0
cc_807 N_A_1356_74#_c_1215_n N_VPWR_c_1501_n 7.39924e-19 $X=7.93 $Y=2.435 $X2=0
+ $Y2=0
cc_808 N_A_1356_74#_c_1216_n N_VPWR_c_1501_n 0.0174628f $X=8.715 $Y=2.75 $X2=0
+ $Y2=0
cc_809 N_A_1356_74#_c_1220_n N_VPWR_c_1501_n 0.00722955f $X=7.47 $Y=2.765 $X2=0
+ $Y2=0
cc_810 N_A_1356_74#_c_1207_n N_VPWR_c_1502_n 0.0111174f $X=9.5 $Y=2.465 $X2=0
+ $Y2=0
cc_811 N_A_1356_74#_c_1211_n N_VPWR_c_1502_n 0.0012294f $X=9.365 $Y=2.06 $X2=0
+ $Y2=0
cc_812 N_A_1356_74#_c_1216_n N_VPWR_c_1502_n 0.0211299f $X=8.715 $Y=2.75 $X2=0
+ $Y2=0
cc_813 N_A_1356_74#_c_1217_n N_VPWR_c_1502_n 0.0264432f $X=9.14 $Y=2.405 $X2=0
+ $Y2=0
cc_814 N_A_1356_74#_c_1209_n N_VPWR_c_1503_n 0.00797697f $X=10.51 $Y=1.765 $X2=0
+ $Y2=0
cc_815 N_A_1356_74#_c_1233_n N_VPWR_c_1507_n 0.00486764f $X=7.76 $Y=2.64 $X2=0
+ $Y2=0
cc_816 N_A_1356_74#_c_1215_n N_VPWR_c_1507_n 0.00277491f $X=7.93 $Y=2.435 $X2=0
+ $Y2=0
cc_817 N_A_1356_74#_c_1220_n N_VPWR_c_1507_n 0.0278413f $X=7.47 $Y=2.765 $X2=0
+ $Y2=0
cc_818 N_A_1356_74#_c_1216_n N_VPWR_c_1513_n 0.0110419f $X=8.715 $Y=2.75 $X2=0
+ $Y2=0
cc_819 N_A_1356_74#_c_1207_n N_VPWR_c_1514_n 0.00413917f $X=9.5 $Y=2.465 $X2=0
+ $Y2=0
cc_820 N_A_1356_74#_c_1209_n N_VPWR_c_1514_n 0.00481995f $X=10.51 $Y=1.765 $X2=0
+ $Y2=0
cc_821 N_A_1356_74#_c_1207_n N_VPWR_c_1496_n 0.00730566f $X=9.5 $Y=2.465 $X2=0
+ $Y2=0
cc_822 N_A_1356_74#_c_1209_n N_VPWR_c_1496_n 0.00508379f $X=10.51 $Y=1.765 $X2=0
+ $Y2=0
cc_823 N_A_1356_74#_c_1211_n N_VPWR_c_1496_n 3.7828e-19 $X=9.365 $Y=2.06 $X2=0
+ $Y2=0
cc_824 N_A_1356_74#_c_1233_n N_VPWR_c_1496_n 0.00785195f $X=7.76 $Y=2.64 $X2=0
+ $Y2=0
cc_825 N_A_1356_74#_c_1214_n N_VPWR_c_1496_n 0.0133813f $X=8.63 $Y=2.435 $X2=0
+ $Y2=0
cc_826 N_A_1356_74#_c_1215_n N_VPWR_c_1496_n 0.00484018f $X=7.93 $Y=2.435 $X2=0
+ $Y2=0
cc_827 N_A_1356_74#_c_1216_n N_VPWR_c_1496_n 0.00915013f $X=8.715 $Y=2.75 $X2=0
+ $Y2=0
cc_828 N_A_1356_74#_c_1217_n N_VPWR_c_1496_n 0.0101254f $X=9.14 $Y=2.405 $X2=0
+ $Y2=0
cc_829 N_A_1356_74#_c_1220_n N_VPWR_c_1496_n 0.0234183f $X=7.47 $Y=2.765 $X2=0
+ $Y2=0
cc_830 N_A_1356_74#_c_1233_n A_1521_508# 0.00378641f $X=7.76 $Y=2.64 $X2=-0.19
+ $Y2=-0.245
cc_831 N_A_1356_74#_c_1215_n A_1521_508# 0.00153468f $X=7.93 $Y=2.435 $X2=-0.19
+ $Y2=-0.245
cc_832 N_A_1356_74#_c_1209_n N_Q_c_1658_n 0.00321103f $X=10.51 $Y=1.765 $X2=0
+ $Y2=0
cc_833 N_A_1356_74#_M1015_g N_VGND_c_1695_n 0.00744268f $X=10.47 $Y=0.79 $X2=0
+ $Y2=0
cc_834 N_A_1356_74#_M1024_g N_VGND_c_1701_n 0.0120948f $X=9.48 $Y=0.8 $X2=0
+ $Y2=0
cc_835 N_A_1356_74#_M1024_g N_VGND_c_1702_n 0.00418347f $X=9.48 $Y=0.8 $X2=0
+ $Y2=0
cc_836 N_A_1356_74#_M1015_g N_VGND_c_1702_n 0.00485498f $X=10.47 $Y=0.79 $X2=0
+ $Y2=0
cc_837 N_A_1356_74#_M1024_g N_VGND_c_1709_n 0.00479212f $X=9.48 $Y=0.8 $X2=0
+ $Y2=0
cc_838 N_A_1356_74#_M1015_g N_VGND_c_1709_n 0.00514438f $X=10.47 $Y=0.79 $X2=0
+ $Y2=0
cc_839 N_A_2022_94#_c_1363_n N_VPWR_c_1503_n 0.0115759f $X=11.045 $Y=1.765 $X2=0
+ $Y2=0
cc_840 N_A_2022_94#_c_1364_n N_VPWR_c_1503_n 5.28947e-19 $X=11.495 $Y=1.765
+ $X2=0 $Y2=0
cc_841 N_A_2022_94#_c_1365_n N_VPWR_c_1503_n 0.0365588f $X=10.285 $Y=1.985 $X2=0
+ $Y2=0
cc_842 N_A_2022_94#_c_1364_n N_VPWR_c_1505_n 0.00822761f $X=11.495 $Y=1.765
+ $X2=0 $Y2=0
cc_843 N_A_2022_94#_c_1365_n N_VPWR_c_1514_n 0.0106977f $X=10.285 $Y=1.985 $X2=0
+ $Y2=0
cc_844 N_A_2022_94#_c_1363_n N_VPWR_c_1515_n 0.00413917f $X=11.045 $Y=1.765
+ $X2=0 $Y2=0
cc_845 N_A_2022_94#_c_1364_n N_VPWR_c_1515_n 0.00411612f $X=11.495 $Y=1.765
+ $X2=0 $Y2=0
cc_846 N_A_2022_94#_c_1363_n N_VPWR_c_1496_n 0.00817726f $X=11.045 $Y=1.765
+ $X2=0 $Y2=0
cc_847 N_A_2022_94#_c_1364_n N_VPWR_c_1496_n 0.00751023f $X=11.495 $Y=1.765
+ $X2=0 $Y2=0
cc_848 N_A_2022_94#_c_1365_n N_VPWR_c_1496_n 0.0122155f $X=10.285 $Y=1.985 $X2=0
+ $Y2=0
cc_849 N_A_2022_94#_M1003_g N_Q_c_1652_n 0.00735215f $X=11.05 $Y=0.74 $X2=0
+ $Y2=0
cc_850 N_A_2022_94#_M1023_g N_Q_c_1652_n 0.00930275f $X=11.48 $Y=0.74 $X2=0
+ $Y2=0
cc_851 N_A_2022_94#_c_1363_n N_Q_c_1655_n 3.89491e-19 $X=11.045 $Y=1.765 $X2=0
+ $Y2=0
cc_852 N_A_2022_94#_c_1364_n N_Q_c_1655_n 0.0111066f $X=11.495 $Y=1.765 $X2=0
+ $Y2=0
cc_853 N_A_2022_94#_M1003_g N_Q_c_1653_n 0.00247818f $X=11.05 $Y=0.74 $X2=0
+ $Y2=0
cc_854 N_A_2022_94#_M1023_g N_Q_c_1653_n 0.00892862f $X=11.48 $Y=0.74 $X2=0
+ $Y2=0
cc_855 N_A_2022_94#_c_1364_n N_Q_c_1653_n 0.0030228f $X=11.495 $Y=1.765 $X2=0
+ $Y2=0
cc_856 N_A_2022_94#_c_1360_n N_Q_c_1653_n 0.0249855f $X=10.975 $Y=1.465 $X2=0
+ $Y2=0
cc_857 N_A_2022_94#_c_1362_n N_Q_c_1653_n 0.0353622f $X=11.48 $Y=1.532 $X2=0
+ $Y2=0
cc_858 N_A_2022_94#_M1003_g N_Q_c_1654_n 0.00245603f $X=11.05 $Y=0.74 $X2=0
+ $Y2=0
cc_859 N_A_2022_94#_M1023_g N_Q_c_1654_n 0.00259764f $X=11.48 $Y=0.74 $X2=0
+ $Y2=0
cc_860 N_A_2022_94#_c_1360_n N_Q_c_1654_n 0.00191579f $X=10.975 $Y=1.465 $X2=0
+ $Y2=0
cc_861 N_A_2022_94#_c_1362_n N_Q_c_1654_n 0.0035553f $X=11.48 $Y=1.532 $X2=0
+ $Y2=0
cc_862 N_A_2022_94#_c_1364_n Q 0.00422024f $X=11.495 $Y=1.765 $X2=0 $Y2=0
cc_863 N_A_2022_94#_c_1362_n Q 0.00632057f $X=11.48 $Y=1.532 $X2=0 $Y2=0
cc_864 N_A_2022_94#_c_1363_n N_Q_c_1658_n 0.0177743f $X=11.045 $Y=1.765 $X2=0
+ $Y2=0
cc_865 N_A_2022_94#_c_1365_n N_Q_c_1658_n 0.0212716f $X=10.285 $Y=1.985 $X2=0
+ $Y2=0
cc_866 N_A_2022_94#_c_1360_n N_Q_c_1658_n 0.0319354f $X=10.975 $Y=1.465 $X2=0
+ $Y2=0
cc_867 N_A_2022_94#_c_1362_n N_Q_c_1658_n 0.00519695f $X=11.48 $Y=1.532 $X2=0
+ $Y2=0
cc_868 N_A_2022_94#_M1003_g N_VGND_c_1695_n 0.00946427f $X=11.05 $Y=0.74 $X2=0
+ $Y2=0
cc_869 N_A_2022_94#_c_1359_n N_VGND_c_1695_n 0.0258905f $X=10.255 $Y=0.615 $X2=0
+ $Y2=0
cc_870 N_A_2022_94#_c_1360_n N_VGND_c_1695_n 0.0285241f $X=10.975 $Y=1.465 $X2=0
+ $Y2=0
cc_871 N_A_2022_94#_c_1362_n N_VGND_c_1695_n 0.00277218f $X=11.48 $Y=1.532 $X2=0
+ $Y2=0
cc_872 N_A_2022_94#_M1023_g N_VGND_c_1697_n 0.00842499f $X=11.48 $Y=0.74 $X2=0
+ $Y2=0
cc_873 N_A_2022_94#_c_1359_n N_VGND_c_1702_n 0.0103491f $X=10.255 $Y=0.615 $X2=0
+ $Y2=0
cc_874 N_A_2022_94#_M1003_g N_VGND_c_1703_n 0.00434272f $X=11.05 $Y=0.74 $X2=0
+ $Y2=0
cc_875 N_A_2022_94#_M1023_g N_VGND_c_1703_n 0.00394617f $X=11.48 $Y=0.74 $X2=0
+ $Y2=0
cc_876 N_A_2022_94#_M1003_g N_VGND_c_1709_n 0.00825059f $X=11.05 $Y=0.74 $X2=0
+ $Y2=0
cc_877 N_A_2022_94#_M1023_g N_VGND_c_1709_n 0.00696181f $X=11.48 $Y=0.74 $X2=0
+ $Y2=0
cc_878 N_A_2022_94#_c_1359_n N_VGND_c_1709_n 0.0113354f $X=10.255 $Y=0.615 $X2=0
+ $Y2=0
cc_879 N_A_27_74#_c_1432_n N_VPWR_M1028_d 0.00134035f $X=2.445 $Y=2.145 $X2=0
+ $Y2=0
cc_880 N_A_27_74#_c_1480_n N_VPWR_M1028_d 0.00532631f $X=1.71 $Y=2.145 $X2=0
+ $Y2=0
cc_881 N_A_27_74#_c_1430_n N_VPWR_c_1497_n 0.0302173f $X=0.28 $Y=2.75 $X2=0
+ $Y2=0
cc_882 N_A_27_74#_c_1431_n N_VPWR_c_1497_n 0.0275301f $X=1.625 $Y=2.275 $X2=0
+ $Y2=0
cc_883 N_A_27_74#_c_1431_n N_VPWR_c_1498_n 0.00106645f $X=1.625 $Y=2.275 $X2=0
+ $Y2=0
cc_884 N_A_27_74#_c_1432_n N_VPWR_c_1498_n 0.00270804f $X=2.445 $Y=2.145 $X2=0
+ $Y2=0
cc_885 N_A_27_74#_c_1480_n N_VPWR_c_1498_n 0.0124964f $X=1.71 $Y=2.145 $X2=0
+ $Y2=0
cc_886 N_A_27_74#_c_1430_n N_VPWR_c_1509_n 0.011066f $X=0.28 $Y=2.75 $X2=0 $Y2=0
cc_887 N_A_27_74#_c_1430_n N_VPWR_c_1496_n 0.00915947f $X=0.28 $Y=2.75 $X2=0
+ $Y2=0
cc_888 N_A_27_74#_c_1427_n N_VGND_c_1698_n 0.00897649f $X=0.28 $Y=0.58 $X2=0
+ $Y2=0
cc_889 N_A_27_74#_c_1427_n N_VGND_c_1709_n 0.00884022f $X=0.28 $Y=0.58 $X2=0
+ $Y2=0
cc_890 N_VPWR_c_1503_n N_Q_c_1655_n 0.0255478f $X=10.82 $Y=2.405 $X2=0 $Y2=0
cc_891 N_VPWR_c_1505_n N_Q_c_1655_n 0.0627709f $X=11.72 $Y=1.985 $X2=0 $Y2=0
cc_892 N_VPWR_c_1515_n N_Q_c_1655_n 0.0136117f $X=11.635 $Y=3.33 $X2=0 $Y2=0
cc_893 N_VPWR_c_1496_n N_Q_c_1655_n 0.0111632f $X=11.76 $Y=3.33 $X2=0 $Y2=0
cc_894 N_VPWR_c_1505_n Q 0.0266814f $X=11.72 $Y=1.985 $X2=0 $Y2=0
cc_895 N_VPWR_M1027_d N_Q_c_1658_n 0.00726973f $X=10.585 $Y=1.84 $X2=0 $Y2=0
cc_896 N_VPWR_c_1503_n N_Q_c_1658_n 0.0204928f $X=10.82 $Y=2.405 $X2=0 $Y2=0
cc_897 N_Q_c_1652_n N_VGND_c_1695_n 0.0312654f $X=11.265 $Y=0.515 $X2=0 $Y2=0
cc_898 N_Q_c_1652_n N_VGND_c_1697_n 0.0597505f $X=11.265 $Y=0.515 $X2=0 $Y2=0
cc_899 N_Q_c_1652_n N_VGND_c_1703_n 0.0159493f $X=11.265 $Y=0.515 $X2=0 $Y2=0
cc_900 N_Q_c_1652_n N_VGND_c_1709_n 0.0130065f $X=11.265 $Y=0.515 $X2=0 $Y2=0
