* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
M1000 a_398_392# B1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.7e+11p pd=2.54e+06u as=1.5868e+12p ps=7.35e+06u
M1001 a_572_392# A2 a_83_260# VPB phighvt w=1e+06u l=150000u
+  ad=3.9e+11p pd=2.78e+06u as=3e+11p ps=2.6e+06u
M1002 a_299_139# A1 VGND VNB nshort w=640000u l=150000u
+  ad=5.3175e+11p pd=5.54e+06u as=5.00375e+11p ps=4.3e+06u
M1003 a_83_260# B1 a_299_139# VNB nshort w=640000u l=150000u
+  ad=2.048e+11p pd=1.92e+06u as=0p ps=0u
M1004 VPWR A1 a_572_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND A2 a_299_139# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR a_83_260# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.304e+11p ps=2.83e+06u
M1007 a_299_139# B2 a_83_260# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_83_260# B2 a_398_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND a_83_260# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
.ends
