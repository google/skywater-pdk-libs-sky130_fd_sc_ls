* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__einvp_4 A TE VGND VNB VPB VPWR Z
X0 a_27_74# A Z VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X1 VGND TE a_27_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X2 a_27_368# a_473_323# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X3 Z A a_27_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X4 a_27_74# TE VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X5 Z A a_27_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X6 a_473_323# TE VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X7 a_473_323# TE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X8 VGND TE a_27_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X9 a_27_368# a_473_323# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X10 a_27_368# A Z VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X11 Z A a_27_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X12 VPWR a_473_323# a_27_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X13 VPWR a_473_323# a_27_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X14 a_27_368# A Z VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X15 a_27_74# A Z VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X16 Z A a_27_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X17 a_27_74# TE VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
.ends
