* NGSPICE file created from sky130_fd_sc_ls__a31oi_1.ext - technology: sky130A

.subckt sky130_fd_sc_ls__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
M1000 Y A1 a_223_74# VNB nshort w=740000u l=150000u
+  ad=3.108e+11p pd=2.32e+06u as=3.108e+11p ps=2.32e+06u
M1001 a_136_368# A1 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=7.28e+11p pd=5.78e+06u as=9.8e+11p ps=6.23e+06u
M1002 a_223_74# A2 a_145_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=1.776e+11p ps=1.96e+06u
M1003 VGND B1 Y VNB nshort w=740000u l=150000u
+  ad=5.291e+11p pd=4.39e+06u as=0p ps=0u
M1004 Y B1 a_136_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=0p ps=0u
M1005 VPWR A2 a_136_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_136_368# A3 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_145_74# A3 VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

