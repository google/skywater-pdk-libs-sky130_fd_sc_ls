* File: sky130_fd_sc_ls__a31oi_2.spice
* Created: Fri Aug 28 12:59:31 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__a31oi_2.pex.spice"
.subckt sky130_fd_sc_ls__a31oi_2  VNB VPB A3 A2 B1 A1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A1	A1
* B1	B1
* A2	A2
* A3	A3
* VPB	VPB
* VNB	VNB
MM1008 N_VGND_M1008_d N_A3_M1008_g N_A_114_74#_M1008_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75003.5 A=0.111 P=1.78 MULT=1
MM1010 N_A_114_74#_M1008_s N_A2_M1010_g N_A_200_74#_M1010_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75000.6 SB=75003.1 A=0.111 P=1.78 MULT=1
MM1013 N_A_114_74#_M1013_d N_A2_M1013_g N_A_200_74#_M1010_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1295 AS=0.1295 PD=1.09 PS=1.09 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75001.1 SB=75002.6 A=0.111 P=1.78 MULT=1
MM1012 N_VGND_M1012_d N_A3_M1012_g N_A_114_74#_M1013_d VNB NSHORT L=0.15 W=0.74
+ AD=0.1554 AS=0.1295 PD=1.16 PS=1.09 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75001.6
+ SB=75002.1 A=0.111 P=1.78 MULT=1
MM1002 N_Y_M1002_d N_B1_M1002_g N_VGND_M1012_d VNB NSHORT L=0.15 W=0.74
+ AD=0.24605 AS=0.1554 PD=1.405 PS=1.16 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75002.2
+ SB=75001.5 A=0.111 P=1.78 MULT=1
MM1005 N_Y_M1002_d N_A1_M1005_g N_A_200_74#_M1005_s VNB NSHORT L=0.15 W=0.74
+ AD=0.24605 AS=0.10915 PD=1.405 PS=1.035 NRD=0 NRS=2.424 M=1 R=4.93333 SA=75003
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1014 N_Y_M1014_d N_A1_M1014_g N_A_200_74#_M1005_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2627 AS=0.10915 PD=2.19 PS=1.035 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75003.5
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1000 N_A_27_368#_M1000_d N_A3_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.1736 PD=2.83 PS=1.43 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75003.5 A=0.168 P=2.54 MULT=1
MM1004 N_A_27_368#_M1004_d N_A2_M1004_g N_VPWR_M1000_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.1904 AS=0.1736 PD=1.46 PS=1.43 NRD=8.7862 NRS=3.5066 M=1 R=7.46667
+ SA=75000.7 SB=75003.1 A=0.168 P=2.54 MULT=1
MM1011 N_A_27_368#_M1004_d N_A2_M1011_g N_VPWR_M1011_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.1904 AS=0.196 PD=1.46 PS=1.47 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.2 SB=75002.6 A=0.168 P=2.54 MULT=1
MM1007 N_A_27_368#_M1007_d N_A3_M1007_g N_VPWR_M1011_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.1736 AS=0.196 PD=1.43 PS=1.47 NRD=2.6201 NRS=10.5395 M=1 R=7.46667
+ SA=75001.7 SB=75002.1 A=0.168 P=2.54 MULT=1
MM1001 N_Y_M1001_d N_B1_M1001_g N_A_27_368#_M1007_d VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.1736 PD=1.42 PS=1.43 NRD=1.7533 NRS=2.6201 M=1 R=7.46667
+ SA=75002.1 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1003 N_Y_M1001_d N_B1_M1003_g N_A_27_368#_M1003_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75002.6 SB=75001.2 A=0.168 P=2.54 MULT=1
MM1006 N_VPWR_M1006_d N_A1_M1006_g N_A_27_368#_M1003_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75003.1 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1009 N_VPWR_M1006_d N_A1_M1009_g N_A_27_368#_M1009_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75003.5 SB=75000.2 A=0.168 P=2.54 MULT=1
DX15_noxref VNB VPB NWDIODE A=8.742 P=13.12
*
.include "sky130_fd_sc_ls__a31oi_2.pxi.spice"
*
.ends
*
*
