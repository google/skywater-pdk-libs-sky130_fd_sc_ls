* File: sky130_fd_sc_ls__clkdlyinv5sd2_1.pex.spice
* Created: Wed Sep  2 10:58:22 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__CLKDLYINV5SD2_1%A 3 6 7 9 10 11 15
r38 15 18 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.57 $Y=1.355
+ $X2=0.57 $Y2=1.52
r39 15 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.57 $Y=1.355
+ $X2=0.57 $Y2=1.19
r40 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.57
+ $Y=1.355 $X2=0.57 $Y2=1.355
r41 11 16 5.88547 $w=6.28e-07 $l=3.1e-07 $layer=LI1_cond $X=0.415 $Y=1.665
+ $X2=0.415 $Y2=1.355
r42 10 16 1.13912 $w=6.28e-07 $l=6e-08 $layer=LI1_cond $X=0.415 $Y=1.295
+ $X2=0.415 $Y2=1.355
r43 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.495 $Y=1.765
+ $X2=0.495 $Y2=2.4
r44 6 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.495 $Y=1.675 $X2=0.495
+ $Y2=1.765
r45 6 18 60.25 $w=1.8e-07 $l=1.55e-07 $layer=POLY_cond $X=0.495 $Y=1.675
+ $X2=0.495 $Y2=1.52
r46 3 17 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.48 $Y=0.58 $X2=0.48
+ $Y2=1.19
.ends

.subckt PM_SKY130_FD_SC_LS__CLKDLYINV5SD2_1%A_28_74# 1 2 9 13 17 19 21 23 25 26
+ 30 37
r62 36 37 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=1.32 $Y=1.295 $X2=1.35
+ $Y2=1.295
r63 31 36 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=1.14 $Y=1.295
+ $X2=1.32 $Y2=1.295
r64 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.14
+ $Y=1.295 $X2=1.14 $Y2=1.295
r65 28 30 25.668 $w=3.28e-07 $l=7.35e-07 $layer=LI1_cond $X=1.14 $Y=2.03
+ $X2=1.14 $Y2=1.295
r66 27 30 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.14 $Y=1.02
+ $X2=1.14 $Y2=1.295
r67 25 27 7.36389 $w=2e-07 $l=2.09105e-07 $layer=LI1_cond $X=0.975 $Y=0.92
+ $X2=1.14 $Y2=1.02
r68 25 26 31.3318 $w=1.98e-07 $l=5.65e-07 $layer=LI1_cond $X=0.975 $Y=0.92
+ $X2=0.41 $Y2=0.92
r69 24 33 4.75367 $w=1.75e-07 $l=1.53e-07 $layer=LI1_cond $X=0.4 $Y=2.117
+ $X2=0.247 $Y2=2.117
r70 23 28 7.68689 $w=1.75e-07 $l=2.03912e-07 $layer=LI1_cond $X=0.975 $Y=2.117
+ $X2=1.14 $Y2=2.03
r71 23 24 36.4416 $w=1.73e-07 $l=5.75e-07 $layer=LI1_cond $X=0.975 $Y=2.117
+ $X2=0.4 $Y2=2.117
r72 19 33 2.73414 $w=3.05e-07 $l=8.8e-08 $layer=LI1_cond $X=0.247 $Y=2.205
+ $X2=0.247 $Y2=2.117
r73 19 21 13.4137 $w=3.03e-07 $l=3.55e-07 $layer=LI1_cond $X=0.247 $Y=2.205
+ $X2=0.247 $Y2=2.56
r74 15 26 7.26812 $w=2e-07 $l=2.01901e-07 $layer=LI1_cond $X=0.252 $Y=0.82
+ $X2=0.41 $Y2=0.92
r75 15 17 8.78052 $w=3.13e-07 $l=2.4e-07 $layer=LI1_cond $X=0.252 $Y=0.82
+ $X2=0.252 $Y2=0.58
r76 11 37 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.35 $Y=1.13
+ $X2=1.35 $Y2=1.295
r77 11 13 213.79 $w=1.8e-07 $l=5.5e-07 $layer=POLY_cond $X=1.35 $Y=1.13 $X2=1.35
+ $Y2=0.58
r78 7 36 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.32 $Y=1.46
+ $X2=1.32 $Y2=1.295
r79 7 9 248.454 $w=2.5e-07 $l=1e-06 $layer=POLY_cond $X=1.32 $Y=1.46 $X2=1.32
+ $Y2=2.46
r80 2 33 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=0.14
+ $Y=1.84 $X2=0.265 $Y2=2.115
r81 2 21 600 $w=1.7e-07 $l=7.8e-07 $layer=licon1_PDIFF $count=1 $X=0.14 $Y=1.84
+ $X2=0.265 $Y2=2.56
r82 1 17 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.14
+ $Y=0.37 $X2=0.265 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_LS__CLKDLYINV5SD2_1%A_288_74# 1 2 9 13 17 22 25 29 32 36
r43 35 36 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=2.62 $Y=1.305
+ $X2=2.655 $Y2=1.305
r44 29 30 6.17723 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.58 $Y=2.815
+ $X2=1.58 $Y2=2.65
r45 26 35 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=2.425 $Y=1.305
+ $X2=2.62 $Y2=1.305
r46 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.425
+ $Y=1.305 $X2=2.425 $Y2=1.305
r47 23 32 0.466467 $w=3.3e-07 $l=1.35e-07 $layer=LI1_cond $X=1.745 $Y=1.305
+ $X2=1.61 $Y2=1.305
r48 23 25 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.745 $Y=1.305
+ $X2=2.425 $Y2=1.305
r49 22 30 23.2623 $w=2.68e-07 $l=5.45e-07 $layer=LI1_cond $X=1.61 $Y=2.105
+ $X2=1.61 $Y2=2.65
r50 19 32 6.31733 $w=2.57e-07 $l=1.65e-07 $layer=LI1_cond $X=1.61 $Y=1.47
+ $X2=1.61 $Y2=1.305
r51 19 22 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.61 $Y=1.47
+ $X2=1.61 $Y2=2.105
r52 15 32 6.31733 $w=2.57e-07 $l=1.71377e-07 $layer=LI1_cond $X=1.597 $Y=1.14
+ $X2=1.61 $Y2=1.305
r53 15 17 26.3416 $w=2.43e-07 $l=5.6e-07 $layer=LI1_cond $X=1.597 $Y=1.14
+ $X2=1.597 $Y2=0.58
r54 11 36 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.655 $Y=1.14
+ $X2=2.655 $Y2=1.305
r55 11 13 217.677 $w=1.8e-07 $l=5.6e-07 $layer=POLY_cond $X=2.655 $Y=1.14
+ $X2=2.655 $Y2=0.58
r56 7 35 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.62 $Y=1.47
+ $X2=2.62 $Y2=1.305
r57 7 9 245.969 $w=2.5e-07 $l=9.9e-07 $layer=POLY_cond $X=2.62 $Y=1.47 $X2=2.62
+ $Y2=2.46
r58 2 29 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.445
+ $Y=1.96 $X2=1.58 $Y2=2.815
r59 2 22 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=1.445
+ $Y=1.96 $X2=1.58 $Y2=2.105
r60 1 17 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.44
+ $Y=0.37 $X2=1.58 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_LS__CLKDLYINV5SD2_1%A_549_74# 1 2 9 13 17 21 27 30 32
c48 27 0 6.34885e-20 $X=3.84 $Y=1.305
r49 32 33 5.87805 $w=3.28e-07 $l=4e-08 $layer=POLY_cond $X=4.045 $Y=1.305
+ $X2=4.085 $Y2=1.305
r50 28 32 30.125 $w=3.28e-07 $l=2.05e-07 $layer=POLY_cond $X=3.84 $Y=1.305
+ $X2=4.045 $Y2=1.305
r51 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.84
+ $Y=1.305 $X2=3.84 $Y2=1.305
r52 25 30 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.97 $Y=1.305
+ $X2=2.885 $Y2=1.305
r53 25 27 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=2.97 $Y=1.305
+ $X2=3.84 $Y2=1.305
r54 21 23 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=2.885 $Y=2.105
+ $X2=2.885 $Y2=2.815
r55 19 30 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.885 $Y=1.39
+ $X2=2.885 $Y2=1.305
r56 19 21 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=2.885 $Y=1.39
+ $X2=2.885 $Y2=2.105
r57 15 30 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.885 $Y=1.22
+ $X2=2.885 $Y2=1.305
r58 15 17 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=2.885 $Y=1.22
+ $X2=2.885 $Y2=0.58
r59 11 33 16.7902 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.085 $Y=1.14
+ $X2=4.085 $Y2=1.305
r60 11 13 217.677 $w=1.8e-07 $l=5.6e-07 $layer=POLY_cond $X=4.085 $Y=1.14
+ $X2=4.085 $Y2=0.58
r61 7 32 9.20465 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.045 $Y=1.47
+ $X2=4.045 $Y2=1.305
r62 7 9 245.969 $w=2.5e-07 $l=9.9e-07 $layer=POLY_cond $X=4.045 $Y=1.47
+ $X2=4.045 $Y2=2.46
r63 2 23 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=2.745
+ $Y=1.96 $X2=2.885 $Y2=2.815
r64 2 21 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.745
+ $Y=1.96 $X2=2.885 $Y2=2.105
r65 1 17 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.745
+ $Y=0.37 $X2=2.885 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_LS__CLKDLYINV5SD2_1%A_682_74# 1 2 9 11 13 16 20 24 25 26
+ 27 31
c56 9 0 6.34885e-20 $X=4.71 $Y=0.58
r57 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.67
+ $Y=1.46 $X2=4.67 $Y2=1.46
r58 29 31 5.12197 $w=2.23e-07 $l=1e-07 $layer=LI1_cond $X=4.642 $Y=1.56
+ $X2=4.642 $Y2=1.46
r59 28 31 21.0001 $w=2.23e-07 $l=4.1e-07 $layer=LI1_cond $X=4.642 $Y=1.05
+ $X2=4.642 $Y2=1.46
r60 26 28 9.89123 $w=1.39e-07 $l=1.4854e-07 $layer=LI1_cond $X=4.53 $Y=0.965
+ $X2=4.642 $Y2=1.05
r61 26 27 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=4.53 $Y=0.965
+ $X2=3.7 $Y2=0.965
r62 24 29 6.9898 $w=1.7e-07 $l=1.4854e-07 $layer=LI1_cond $X=4.53 $Y=1.645
+ $X2=4.642 $Y2=1.56
r63 24 25 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=4.53 $Y=1.645
+ $X2=3.655 $Y2=1.645
r64 20 22 34.0931 $w=2.38e-07 $l=7.1e-07 $layer=LI1_cond $X=3.535 $Y=2.105
+ $X2=3.535 $Y2=2.815
r65 18 25 7.07814 $w=1.7e-07 $l=1.56844e-07 $layer=LI1_cond $X=3.535 $Y=1.73
+ $X2=3.655 $Y2=1.645
r66 18 20 18.0069 $w=2.38e-07 $l=3.75e-07 $layer=LI1_cond $X=3.535 $Y=1.73
+ $X2=3.535 $Y2=2.105
r67 14 27 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.535 $Y=0.88
+ $X2=3.7 $Y2=0.965
r68 14 16 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=3.535 $Y=0.88
+ $X2=3.535 $Y2=0.565
r69 11 32 62.3432 $w=2.85e-07 $l=3.29052e-07 $layer=POLY_cond $X=4.72 $Y=1.765
+ $X2=4.67 $Y2=1.46
r70 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.72 $Y=1.765
+ $X2=4.72 $Y2=2.4
r71 7 32 38.666 $w=2.85e-07 $l=1.83916e-07 $layer=POLY_cond $X=4.71 $Y=1.295
+ $X2=4.67 $Y2=1.46
r72 7 9 366.628 $w=1.5e-07 $l=7.15e-07 $layer=POLY_cond $X=4.71 $Y=1.295
+ $X2=4.71 $Y2=0.58
r73 2 22 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=3.41
+ $Y=1.96 $X2=3.535 $Y2=2.815
r74 2 20 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=3.41
+ $Y=1.96 $X2=3.535 $Y2=2.105
r75 1 16 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=3.41
+ $Y=0.37 $X2=3.535 $Y2=0.565
.ends

.subckt PM_SKY130_FD_SC_LS__CLKDLYINV5SD2_1%VPWR 1 2 3 12 16 22 26 28 33 38 48
+ 49 52 55 58 65
r50 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r51 56 65 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.92 $Y2=3.33
r52 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r53 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r54 49 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r55 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r56 46 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.66 $Y=3.33
+ $X2=4.495 $Y2=3.33
r57 46 48 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=4.66 $Y=3.33
+ $X2=5.04 $Y2=3.33
r58 45 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r59 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r60 41 44 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.64 $Y=3.33
+ $X2=4.08 $Y2=3.33
r61 39 55 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=2.265 $Y=3.33
+ $X2=2.09 $Y2=3.33
r62 39 41 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=2.265 $Y=3.33
+ $X2=2.64 $Y2=3.33
r63 38 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.33 $Y=3.33
+ $X2=4.495 $Y2=3.33
r64 38 44 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=4.33 $Y=3.33
+ $X2=4.08 $Y2=3.33
r65 37 65 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.92 $Y2=3.33
r66 37 53 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r67 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r68 34 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.905 $Y=3.33
+ $X2=0.74 $Y2=3.33
r69 34 36 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=0.905 $Y=3.33
+ $X2=1.68 $Y2=3.33
r70 33 55 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=1.915 $Y=3.33
+ $X2=2.09 $Y2=3.33
r71 33 36 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=1.915 $Y=3.33
+ $X2=1.68 $Y2=3.33
r72 31 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r73 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r74 28 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.575 $Y=3.33
+ $X2=0.74 $Y2=3.33
r75 28 30 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.575 $Y=3.33
+ $X2=0.24 $Y2=3.33
r76 26 45 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=4.08 $Y2=3.33
r77 26 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r78 26 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r79 22 25 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=4.495 $Y=1.985
+ $X2=4.495 $Y2=2.415
r80 20 58 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.495 $Y=3.245
+ $X2=4.495 $Y2=3.33
r81 20 25 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=4.495 $Y=3.245
+ $X2=4.495 $Y2=2.415
r82 16 19 23.3781 $w=3.48e-07 $l=7.1e-07 $layer=LI1_cond $X=2.09 $Y=2.105
+ $X2=2.09 $Y2=2.815
r83 14 55 1.07557 $w=3.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.09 $Y=3.245
+ $X2=2.09 $Y2=3.33
r84 14 19 14.1586 $w=3.48e-07 $l=4.3e-07 $layer=LI1_cond $X=2.09 $Y=3.245
+ $X2=2.09 $Y2=2.815
r85 10 52 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.74 $Y=3.245
+ $X2=0.74 $Y2=3.33
r86 10 12 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=0.74 $Y=3.245
+ $X2=0.74 $Y2=2.465
r87 3 25 300 $w=1.7e-07 $l=5.95735e-07 $layer=licon1_PDIFF $count=2 $X=4.17
+ $Y=1.96 $X2=4.495 $Y2=2.415
r88 3 22 600 $w=1.7e-07 $l=3.37268e-07 $layer=licon1_PDIFF $count=1 $X=4.17
+ $Y=1.96 $X2=4.495 $Y2=1.985
r89 2 19 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=1.975
+ $Y=1.96 $X2=2.1 $Y2=2.815
r90 2 16 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.975
+ $Y=1.96 $X2=2.1 $Y2=2.105
r91 1 12 300 $w=1.7e-07 $l=7.04894e-07 $layer=licon1_PDIFF $count=2 $X=0.57
+ $Y=1.84 $X2=0.74 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LS__CLKDLYINV5SD2_1%Y 1 2 7 8 9 10 11 12 13 47
r17 42 43 6.10729 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=5.01 $Y=0.59
+ $X2=5.01 $Y2=0.755
r18 30 47 1.44055 $w=3.58e-07 $l=4.5e-08 $layer=LI1_cond $X=5.01 $Y=2.08
+ $X2=5.01 $Y2=2.035
r19 13 45 10.2198 $w=2.63e-07 $l=2.35e-07 $layer=LI1_cond $X=5.057 $Y=1.665
+ $X2=5.057 $Y2=1.9
r20 11 12 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=5.01 $Y=2.405
+ $X2=5.01 $Y2=2.775
r21 10 47 0.640246 $w=3.58e-07 $l=2e-08 $layer=LI1_cond $X=5.01 $Y=2.015
+ $X2=5.01 $Y2=2.035
r22 10 45 4.50667 $w=3.58e-07 $l=1.15e-07 $layer=LI1_cond $X=5.01 $Y=2.015
+ $X2=5.01 $Y2=1.9
r23 10 11 9.76375 $w=3.58e-07 $l=3.05e-07 $layer=LI1_cond $X=5.01 $Y=2.1
+ $X2=5.01 $Y2=2.405
r24 10 30 0.640246 $w=3.58e-07 $l=2e-08 $layer=LI1_cond $X=5.01 $Y=2.1 $X2=5.01
+ $Y2=2.08
r25 9 13 16.0907 $w=2.63e-07 $l=3.7e-07 $layer=LI1_cond $X=5.057 $Y=1.295
+ $X2=5.057 $Y2=1.665
r26 8 9 16.0907 $w=2.63e-07 $l=3.7e-07 $layer=LI1_cond $X=5.057 $Y=0.925
+ $X2=5.057 $Y2=1.295
r27 8 43 7.39303 $w=2.63e-07 $l=1.7e-07 $layer=LI1_cond $X=5.057 $Y=0.925
+ $X2=5.057 $Y2=0.755
r28 7 42 1.12043 $w=3.58e-07 $l=3.5e-08 $layer=LI1_cond $X=5.01 $Y=0.555
+ $X2=5.01 $Y2=0.59
r29 2 47 400 $w=1.7e-07 $l=2.92404e-07 $layer=licon1_PDIFF $count=1 $X=4.795
+ $Y=1.84 $X2=4.95 $Y2=2.065
r30 2 12 400 $w=1.7e-07 $l=1.04463e-06 $layer=licon1_PDIFF $count=1 $X=4.795
+ $Y=1.84 $X2=4.95 $Y2=2.81
r31 1 42 182 $w=1.7e-07 $l=2.81425e-07 $layer=licon1_NDIFF $count=1 $X=4.785
+ $Y=0.37 $X2=4.925 $Y2=0.59
.ends

.subckt PM_SKY130_FD_SC_LS__CLKDLYINV5SD2_1%VGND 1 2 3 12 16 20 22 24 29 34 44
+ 45 48 51 54 61
r48 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r49 52 61 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.92
+ $Y2=0
r50 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r51 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r52 45 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.56
+ $Y2=0
r53 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r54 42 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.66 $Y=0 $X2=4.495
+ $Y2=0
r55 42 44 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=4.66 $Y=0 $X2=5.04
+ $Y2=0
r56 41 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r57 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r58 37 40 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.64 $Y=0 $X2=4.08
+ $Y2=0
r59 35 51 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=2.265 $Y=0 $X2=2.09
+ $Y2=0
r60 35 37 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=2.265 $Y=0 $X2=2.64
+ $Y2=0
r61 34 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.33 $Y=0 $X2=4.495
+ $Y2=0
r62 34 40 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=4.33 $Y=0 $X2=4.08
+ $Y2=0
r63 33 61 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.92
+ $Y2=0
r64 33 49 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r65 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r66 30 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.915 $Y=0 $X2=0.75
+ $Y2=0
r67 30 32 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=0.915 $Y=0 $X2=1.68
+ $Y2=0
r68 29 51 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=1.915 $Y=0 $X2=2.09
+ $Y2=0
r69 29 32 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=1.915 $Y=0 $X2=1.68
+ $Y2=0
r70 27 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r71 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r72 24 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.585 $Y=0 $X2=0.75
+ $Y2=0
r73 24 26 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.585 $Y=0 $X2=0.24
+ $Y2=0
r74 22 41 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.64 $Y=0 $X2=4.08
+ $Y2=0
r75 22 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r76 22 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r77 18 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.495 $Y=0.085
+ $X2=4.495 $Y2=0
r78 18 20 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=4.495 $Y=0.085
+ $X2=4.495 $Y2=0.585
r79 14 51 1.07557 $w=3.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.09 $Y=0.085
+ $X2=2.09 $Y2=0
r80 14 16 16.2988 $w=3.48e-07 $l=4.95e-07 $layer=LI1_cond $X=2.09 $Y=0.085
+ $X2=2.09 $Y2=0.58
r81 10 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=0.085
+ $X2=0.75 $Y2=0
r82 10 12 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.75 $Y=0.085
+ $X2=0.75 $Y2=0.565
r83 3 20 182 $w=1.7e-07 $l=4.13763e-07 $layer=licon1_NDIFF $count=1 $X=4.175
+ $Y=0.37 $X2=4.495 $Y2=0.585
r84 2 16 182 $w=1.7e-07 $l=2.67208e-07 $layer=licon1_NDIFF $count=1 $X=1.975
+ $Y=0.37 $X2=2.105 $Y2=0.58
r85 1 12 182 $w=1.7e-07 $l=2.75772e-07 $layer=licon1_NDIFF $count=1 $X=0.555
+ $Y=0.37 $X2=0.75 $Y2=0.565
.ends

