* File: sky130_fd_sc_ls__clkinv_1.spice
* Created: Fri Aug 28 13:10:37 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__clkinv_1.pex.spice"
.subckt sky130_fd_sc_ls__clkinv_1  VNB VPB A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1000 N_Y_M1000_d N_A_M1000_g N_VGND_M1000_s VNB NSHORT L=0.15 W=0.42
+ AD=0.22535 AS=0.1491 PD=2.17 PS=1.55 NRD=0 NRS=19.992 M=1 R=2.8 SA=75000.3
+ SB=75000.5 A=0.063 P=1.14 MULT=1
MM1001 N_Y_M1001_d N_A_M1001_g N_VPWR_M1001_s VPB PHIGHVT L=0.15 W=0.84 AD=0.126
+ AS=0.2394 PD=1.14 PS=2.25 NRD=2.3443 NRS=2.3443 M=1 R=5.6 SA=75000.2
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1002 N_Y_M1001_d N_A_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=0.15 W=0.84 AD=0.126
+ AS=0.2394 PD=1.14 PS=2.25 NRD=2.3443 NRS=2.3443 M=1 R=5.6 SA=75000.7
+ SB=75000.2 A=0.126 P=1.98 MULT=1
DX3_noxref VNB VPB NWDIODE A=3.3852 P=7.36
*
.include "sky130_fd_sc_ls__clkinv_1.pxi.spice"
*
.ends
*
*
