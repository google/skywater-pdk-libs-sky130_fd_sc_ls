* File: sky130_fd_sc_ls__buf_16.pex.spice
* Created: Wed Sep  2 10:56:24 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__BUF_16%A_83_260# 1 2 3 4 5 6 19 21 24 28 30 32 35 37
+ 39 42 44 46 49 51 53 56 58 60 63 65 67 70 72 74 77 79 81 84 86 88 91 93 95 98
+ 100 102 105 107 109 112 114 116 117 119 122 124 126 129 131 132 133 134 137
+ 141 143 145 149 153 155 157 159 161 165 170 171 173 174 200 201 209 216 223
+ 230 237 244 251 254
c457 254 0 2.68688e-20 $X=7.305 $Y=1.532
c458 200 0 8.59108e-19 $X=7.505 $Y=1.665
r459 254 255 9.38961 $w=3.85e-07 $l=7.5e-08 $layer=POLY_cond $X=7.305 $Y=1.532
+ $X2=7.38 $Y2=1.532
r460 253 254 44.4442 $w=3.85e-07 $l=3.55e-07 $layer=POLY_cond $X=6.95 $Y=1.532
+ $X2=7.305 $Y2=1.532
r461 252 253 11.8935 $w=3.85e-07 $l=9.5e-08 $layer=POLY_cond $X=6.855 $Y=1.532
+ $X2=6.95 $Y2=1.532
r462 250 252 23.787 $w=3.85e-07 $l=1.9e-07 $layer=POLY_cond $X=6.665 $Y=1.532
+ $X2=6.855 $Y2=1.532
r463 250 251 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.665
+ $Y=1.465 $X2=6.665 $Y2=1.465
r464 248 250 32.5506 $w=3.85e-07 $l=2.6e-07 $layer=POLY_cond $X=6.405 $Y=1.532
+ $X2=6.665 $Y2=1.532
r465 247 248 3.12987 $w=3.85e-07 $l=2.5e-08 $layer=POLY_cond $X=6.38 $Y=1.532
+ $X2=6.405 $Y2=1.532
r466 246 247 53.2078 $w=3.85e-07 $l=4.25e-07 $layer=POLY_cond $X=5.955 $Y=1.532
+ $X2=6.38 $Y2=1.532
r467 245 246 0.625974 $w=3.85e-07 $l=5e-09 $layer=POLY_cond $X=5.95 $Y=1.532
+ $X2=5.955 $Y2=1.532
r468 243 245 26.2909 $w=3.85e-07 $l=2.1e-07 $layer=POLY_cond $X=5.74 $Y=1.532
+ $X2=5.95 $Y2=1.532
r469 243 244 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.74
+ $Y=1.465 $X2=5.74 $Y2=1.465
r470 241 243 29.4208 $w=3.85e-07 $l=2.35e-07 $layer=POLY_cond $X=5.505 $Y=1.532
+ $X2=5.74 $Y2=1.532
r471 240 241 15.6494 $w=3.85e-07 $l=1.25e-07 $layer=POLY_cond $X=5.38 $Y=1.532
+ $X2=5.505 $Y2=1.532
r472 239 240 40.6883 $w=3.85e-07 $l=3.25e-07 $layer=POLY_cond $X=5.055 $Y=1.532
+ $X2=5.38 $Y2=1.532
r473 238 239 13.1455 $w=3.85e-07 $l=1.05e-07 $layer=POLY_cond $X=4.95 $Y=1.532
+ $X2=5.055 $Y2=1.532
r474 236 238 28.7948 $w=3.85e-07 $l=2.3e-07 $layer=POLY_cond $X=4.72 $Y=1.532
+ $X2=4.95 $Y2=1.532
r475 236 237 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.72
+ $Y=1.465 $X2=4.72 $Y2=1.465
r476 234 236 14.3974 $w=3.85e-07 $l=1.15e-07 $layer=POLY_cond $X=4.605 $Y=1.532
+ $X2=4.72 $Y2=1.532
r477 233 234 28.1688 $w=3.85e-07 $l=2.25e-07 $layer=POLY_cond $X=4.38 $Y=1.532
+ $X2=4.605 $Y2=1.532
r478 232 233 28.1688 $w=3.85e-07 $l=2.25e-07 $layer=POLY_cond $X=4.155 $Y=1.532
+ $X2=4.38 $Y2=1.532
r479 231 232 25.6649 $w=3.85e-07 $l=2.05e-07 $layer=POLY_cond $X=3.95 $Y=1.532
+ $X2=4.155 $Y2=1.532
r480 229 231 11.2675 $w=3.85e-07 $l=9e-08 $layer=POLY_cond $X=3.86 $Y=1.532
+ $X2=3.95 $Y2=1.532
r481 229 230 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.86
+ $Y=1.465 $X2=3.86 $Y2=1.465
r482 227 229 19.4052 $w=3.85e-07 $l=1.55e-07 $layer=POLY_cond $X=3.705 $Y=1.532
+ $X2=3.86 $Y2=1.532
r483 226 227 23.161 $w=3.85e-07 $l=1.85e-07 $layer=POLY_cond $X=3.52 $Y=1.532
+ $X2=3.705 $Y2=1.532
r484 225 226 33.1766 $w=3.85e-07 $l=2.65e-07 $layer=POLY_cond $X=3.255 $Y=1.532
+ $X2=3.52 $Y2=1.532
r485 224 225 20.6571 $w=3.85e-07 $l=1.65e-07 $layer=POLY_cond $X=3.09 $Y=1.532
+ $X2=3.255 $Y2=1.532
r486 222 224 11.8935 $w=3.85e-07 $l=9.5e-08 $layer=POLY_cond $X=2.995 $Y=1.532
+ $X2=3.09 $Y2=1.532
r487 222 223 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.995
+ $Y=1.465 $X2=2.995 $Y2=1.465
r488 220 222 23.787 $w=3.85e-07 $l=1.9e-07 $layer=POLY_cond $X=2.805 $Y=1.532
+ $X2=2.995 $Y2=1.532
r489 219 220 18.1532 $w=3.85e-07 $l=1.45e-07 $layer=POLY_cond $X=2.66 $Y=1.532
+ $X2=2.805 $Y2=1.532
r490 218 219 38.1844 $w=3.85e-07 $l=3.05e-07 $layer=POLY_cond $X=2.355 $Y=1.532
+ $X2=2.66 $Y2=1.532
r491 217 218 15.6494 $w=3.85e-07 $l=1.25e-07 $layer=POLY_cond $X=2.23 $Y=1.532
+ $X2=2.355 $Y2=1.532
r492 215 217 24.413 $w=3.85e-07 $l=1.95e-07 $layer=POLY_cond $X=2.035 $Y=1.532
+ $X2=2.23 $Y2=1.532
r493 215 216 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.035
+ $Y=1.465 $X2=2.035 $Y2=1.465
r494 213 215 22.5351 $w=3.85e-07 $l=1.8e-07 $layer=POLY_cond $X=1.855 $Y=1.532
+ $X2=2.035 $Y2=1.532
r495 212 213 6.88571 $w=3.85e-07 $l=5.5e-08 $layer=POLY_cond $X=1.8 $Y=1.532
+ $X2=1.855 $Y2=1.532
r496 211 212 49.4519 $w=3.85e-07 $l=3.95e-07 $layer=POLY_cond $X=1.405 $Y=1.532
+ $X2=1.8 $Y2=1.532
r497 210 211 4.38182 $w=3.85e-07 $l=3.5e-08 $layer=POLY_cond $X=1.37 $Y=1.532
+ $X2=1.405 $Y2=1.532
r498 208 210 27.5429 $w=3.85e-07 $l=2.2e-07 $layer=POLY_cond $X=1.15 $Y=1.532
+ $X2=1.37 $Y2=1.532
r499 208 209 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.15
+ $Y=1.465 $X2=1.15 $Y2=1.465
r500 206 208 24.413 $w=3.85e-07 $l=1.95e-07 $layer=POLY_cond $X=0.955 $Y=1.532
+ $X2=1.15 $Y2=1.532
r501 205 206 1.87792 $w=3.85e-07 $l=1.5e-08 $layer=POLY_cond $X=0.94 $Y=1.532
+ $X2=0.955 $Y2=1.532
r502 204 205 53.8338 $w=3.85e-07 $l=4.3e-07 $layer=POLY_cond $X=0.51 $Y=1.532
+ $X2=0.94 $Y2=1.532
r503 203 204 0.625974 $w=3.85e-07 $l=5e-09 $layer=POLY_cond $X=0.505 $Y=1.532
+ $X2=0.51 $Y2=1.532
r504 200 201 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.505 $Y=1.665
+ $X2=7.505 $Y2=1.665
r505 198 251 7.43512 $w=3.08e-07 $l=2e-07 $layer=LI1_cond $X=6.655 $Y=1.665
+ $X2=6.655 $Y2=1.465
r506 197 200 0.548572 $w=2.3e-07 $l=8.55e-07 $layer=MET1_cond $X=6.65 $Y=1.665
+ $X2=7.505 $Y2=1.665
r507 197 198 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.65 $Y=1.665
+ $X2=6.65 $Y2=1.665
r508 195 244 7.43512 $w=3.08e-07 $l=2e-07 $layer=LI1_cond $X=5.735 $Y=1.665
+ $X2=5.735 $Y2=1.465
r509 194 197 0.587068 $w=2.3e-07 $l=9.15e-07 $layer=MET1_cond $X=5.735 $Y=1.665
+ $X2=6.65 $Y2=1.665
r510 194 195 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.735 $Y=1.665
+ $X2=5.735 $Y2=1.665
r511 192 237 8.21549 $w=2.97e-07 $l=2e-07 $layer=LI1_cond $X=4.71 $Y=1.665
+ $X2=4.71 $Y2=1.465
r512 191 194 0.622356 $w=2.3e-07 $l=9.7e-07 $layer=MET1_cond $X=4.765 $Y=1.665
+ $X2=5.735 $Y2=1.665
r513 191 192 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.765 $Y=1.665
+ $X2=4.765 $Y2=1.665
r514 189 230 6.61247 $w=3.69e-07 $l=2e-07 $layer=LI1_cond $X=3.85 $Y=1.665
+ $X2=3.85 $Y2=1.465
r515 188 191 0.564612 $w=2.3e-07 $l=8.8e-07 $layer=MET1_cond $X=3.885 $Y=1.665
+ $X2=4.765 $Y2=1.665
r516 188 189 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.885 $Y=1.665
+ $X2=3.885 $Y2=1.665
r517 186 223 7.81317 $w=2.93e-07 $l=2e-07 $layer=LI1_cond $X=2.992 $Y=1.665
+ $X2=2.992 $Y2=1.465
r518 185 188 0.571028 $w=2.3e-07 $l=8.9e-07 $layer=MET1_cond $X=2.995 $Y=1.665
+ $X2=3.885 $Y2=1.665
r519 185 186 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.995 $Y=1.665
+ $X2=2.995 $Y2=1.665
r520 183 216 8.08732 $w=2.83e-07 $l=2e-07 $layer=LI1_cond $X=2.032 $Y=1.665
+ $X2=2.032 $Y2=1.465
r521 182 185 0.61594 $w=2.3e-07 $l=9.6e-07 $layer=MET1_cond $X=2.035 $Y=1.665
+ $X2=2.995 $Y2=1.665
r522 182 183 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.035 $Y=1.665
+ $X2=2.035 $Y2=1.665
r523 179 209 7.43512 $w=3.08e-07 $l=2e-07 $layer=LI1_cond $X=1.14 $Y=1.665
+ $X2=1.14 $Y2=1.465
r524 178 182 0.574236 $w=2.3e-07 $l=8.95e-07 $layer=MET1_cond $X=1.14 $Y=1.665
+ $X2=2.035 $Y2=1.665
r525 178 179 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.14 $Y=1.665
+ $X2=1.14 $Y2=1.665
r526 168 201 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=7.505 $Y=1.95
+ $X2=7.505 $Y2=1.665
r527 167 201 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=7.505 $Y=1.18
+ $X2=7.505 $Y2=1.665
r528 163 165 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=9.82 $Y=1.01
+ $X2=9.82 $Y2=0.515
r529 159 176 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.83 $Y=2.12
+ $X2=9.83 $Y2=2.035
r530 159 161 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=9.83 $Y=2.12
+ $X2=9.83 $Y2=2.815
r531 158 173 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.095 $Y=2.035
+ $X2=8.93 $Y2=2.035
r532 157 176 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.665 $Y=2.035
+ $X2=9.83 $Y2=2.035
r533 157 158 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=9.665 $Y=2.035
+ $X2=9.095 $Y2=2.035
r534 156 174 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.97 $Y=1.095
+ $X2=8.885 $Y2=1.095
r535 155 163 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=9.695 $Y=1.095
+ $X2=9.82 $Y2=1.01
r536 155 156 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=9.695 $Y=1.095
+ $X2=8.97 $Y2=1.095
r537 151 174 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.885 $Y=1.01
+ $X2=8.885 $Y2=1.095
r538 151 153 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=8.885 $Y=1.01
+ $X2=8.885 $Y2=0.515
r539 147 173 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.93 $Y=2.12
+ $X2=8.93 $Y2=2.035
r540 147 149 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=8.93 $Y=2.12
+ $X2=8.93 $Y2=2.815
r541 146 170 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.195 $Y=2.035
+ $X2=8.03 $Y2=2.035
r542 145 173 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.765 $Y=2.035
+ $X2=8.93 $Y2=2.035
r543 145 146 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=8.765 $Y=2.035
+ $X2=8.195 $Y2=2.035
r544 144 171 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.11 $Y=1.095
+ $X2=8.025 $Y2=1.095
r545 143 174 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.8 $Y=1.095
+ $X2=8.885 $Y2=1.095
r546 143 144 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=8.8 $Y=1.095
+ $X2=8.11 $Y2=1.095
r547 139 171 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.025 $Y=1.01
+ $X2=8.025 $Y2=1.095
r548 139 141 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=8.025 $Y=1.01
+ $X2=8.025 $Y2=0.515
r549 135 170 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.03 $Y=2.12
+ $X2=8.03 $Y2=2.035
r550 135 137 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=8.03 $Y=2.12
+ $X2=8.03 $Y2=2.815
r551 134 168 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.59 $Y=2.035
+ $X2=7.505 $Y2=1.95
r552 133 170 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.865 $Y=2.035
+ $X2=8.03 $Y2=2.035
r553 133 134 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=7.865 $Y=2.035
+ $X2=7.59 $Y2=2.035
r554 132 167 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.59 $Y=1.095
+ $X2=7.505 $Y2=1.18
r555 131 171 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.94 $Y=1.095
+ $X2=8.025 $Y2=1.095
r556 131 132 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=7.94 $Y=1.095
+ $X2=7.59 $Y2=1.095
r557 127 255 24.9301 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=7.38 $Y=1.3
+ $X2=7.38 $Y2=1.532
r558 127 129 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=7.38 $Y=1.3
+ $X2=7.38 $Y2=0.74
r559 124 254 24.9301 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=7.305 $Y=1.765
+ $X2=7.305 $Y2=1.532
r560 124 126 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.305 $Y=1.765
+ $X2=7.305 $Y2=2.4
r561 120 253 24.9301 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=6.95 $Y=1.3
+ $X2=6.95 $Y2=1.532
r562 120 122 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=6.95 $Y=1.3
+ $X2=6.95 $Y2=0.74
r563 117 252 24.9301 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=6.855 $Y=1.765
+ $X2=6.855 $Y2=1.532
r564 117 119 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.855 $Y=1.765
+ $X2=6.855 $Y2=2.4
r565 114 248 24.9301 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=6.405 $Y=1.765
+ $X2=6.405 $Y2=1.532
r566 114 116 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.405 $Y=1.765
+ $X2=6.405 $Y2=2.4
r567 110 247 24.9301 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=6.38 $Y=1.3
+ $X2=6.38 $Y2=1.532
r568 110 112 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=6.38 $Y=1.3
+ $X2=6.38 $Y2=0.74
r569 107 246 24.9301 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=5.955 $Y=1.765
+ $X2=5.955 $Y2=1.532
r570 107 109 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.955 $Y=1.765
+ $X2=5.955 $Y2=2.4
r571 103 245 24.9301 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=5.95 $Y=1.3
+ $X2=5.95 $Y2=1.532
r572 103 105 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=5.95 $Y=1.3
+ $X2=5.95 $Y2=0.74
r573 100 241 24.9301 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=5.505 $Y=1.765
+ $X2=5.505 $Y2=1.532
r574 100 102 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.505 $Y=1.765
+ $X2=5.505 $Y2=2.4
r575 96 240 24.9301 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=5.38 $Y=1.3
+ $X2=5.38 $Y2=1.532
r576 96 98 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=5.38 $Y=1.3
+ $X2=5.38 $Y2=0.74
r577 93 239 24.9301 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=5.055 $Y=1.765
+ $X2=5.055 $Y2=1.532
r578 93 95 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.055 $Y=1.765
+ $X2=5.055 $Y2=2.4
r579 89 238 24.9301 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=4.95 $Y=1.3
+ $X2=4.95 $Y2=1.532
r580 89 91 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.95 $Y=1.3
+ $X2=4.95 $Y2=0.74
r581 86 234 24.9301 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=4.605 $Y=1.765
+ $X2=4.605 $Y2=1.532
r582 86 88 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.605 $Y=1.765
+ $X2=4.605 $Y2=2.4
r583 82 233 24.9301 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=4.38 $Y=1.3
+ $X2=4.38 $Y2=1.532
r584 82 84 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.38 $Y=1.3
+ $X2=4.38 $Y2=0.74
r585 79 232 24.9301 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=4.155 $Y=1.765
+ $X2=4.155 $Y2=1.532
r586 79 81 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.155 $Y=1.765
+ $X2=4.155 $Y2=2.4
r587 75 231 24.9301 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=3.95 $Y=1.3
+ $X2=3.95 $Y2=1.532
r588 75 77 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.95 $Y=1.3
+ $X2=3.95 $Y2=0.74
r589 72 227 24.9301 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=3.705 $Y=1.765
+ $X2=3.705 $Y2=1.532
r590 72 74 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.705 $Y=1.765
+ $X2=3.705 $Y2=2.4
r591 68 226 24.9301 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=3.52 $Y=1.3
+ $X2=3.52 $Y2=1.532
r592 68 70 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.52 $Y=1.3
+ $X2=3.52 $Y2=0.74
r593 65 225 24.9301 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=3.255 $Y=1.765
+ $X2=3.255 $Y2=1.532
r594 65 67 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.255 $Y=1.765
+ $X2=3.255 $Y2=2.4
r595 61 224 24.9301 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=3.09 $Y=1.3
+ $X2=3.09 $Y2=1.532
r596 61 63 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.09 $Y=1.3
+ $X2=3.09 $Y2=0.74
r597 58 220 24.9301 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=2.805 $Y=1.765
+ $X2=2.805 $Y2=1.532
r598 58 60 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.805 $Y=1.765
+ $X2=2.805 $Y2=2.4
r599 54 219 24.9301 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=2.66 $Y=1.3
+ $X2=2.66 $Y2=1.532
r600 54 56 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.66 $Y=1.3
+ $X2=2.66 $Y2=0.74
r601 51 218 24.9301 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=2.355 $Y=1.765
+ $X2=2.355 $Y2=1.532
r602 51 53 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.355 $Y=1.765
+ $X2=2.355 $Y2=2.4
r603 47 217 24.9301 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=2.23 $Y=1.3
+ $X2=2.23 $Y2=1.532
r604 47 49 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.23 $Y=1.3
+ $X2=2.23 $Y2=0.74
r605 44 213 24.9301 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=1.855 $Y=1.765
+ $X2=1.855 $Y2=1.532
r606 44 46 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.855 $Y=1.765
+ $X2=1.855 $Y2=2.4
r607 40 212 24.9301 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=1.8 $Y=1.3
+ $X2=1.8 $Y2=1.532
r608 40 42 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.8 $Y=1.3 $X2=1.8
+ $Y2=0.74
r609 37 211 24.9301 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=1.405 $Y=1.765
+ $X2=1.405 $Y2=1.532
r610 37 39 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.405 $Y=1.765
+ $X2=1.405 $Y2=2.4
r611 33 210 24.9301 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=1.37 $Y=1.3
+ $X2=1.37 $Y2=1.532
r612 33 35 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.37 $Y=1.3
+ $X2=1.37 $Y2=0.74
r613 30 206 24.9301 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=0.955 $Y=1.765
+ $X2=0.955 $Y2=1.532
r614 30 32 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.955 $Y=1.765
+ $X2=0.955 $Y2=2.4
r615 26 205 24.9301 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=0.94 $Y=1.3
+ $X2=0.94 $Y2=1.532
r616 26 28 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.94 $Y=1.3
+ $X2=0.94 $Y2=0.74
r617 22 204 24.9301 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=0.51 $Y=1.3
+ $X2=0.51 $Y2=1.532
r618 22 24 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.51 $Y=1.3
+ $X2=0.51 $Y2=0.74
r619 19 203 24.9301 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=1.532
r620 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.4
r621 6 176 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=9.68
+ $Y=1.84 $X2=9.83 $Y2=2.115
r622 6 161 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=9.68
+ $Y=1.84 $X2=9.83 $Y2=2.815
r623 5 173 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=8.78
+ $Y=1.84 $X2=8.93 $Y2=2.115
r624 5 149 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=8.78
+ $Y=1.84 $X2=8.93 $Y2=2.815
r625 4 170 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=7.88
+ $Y=1.84 $X2=8.03 $Y2=2.115
r626 4 137 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=7.88
+ $Y=1.84 $X2=8.03 $Y2=2.815
r627 3 165 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.64
+ $Y=0.37 $X2=9.78 $Y2=0.515
r628 2 153 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.745
+ $Y=0.37 $X2=8.885 $Y2=0.515
r629 1 141 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.885
+ $Y=0.37 $X2=8.025 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__BUF_16%A 1 3 6 10 12 14 17 19 21 24 26 28 31 33 35
+ 36 38 41 43 44 45 46 47 69
c125 69 0 1.18608e-19 $X=10.055 $Y=1.557
c126 1 0 1.43649e-19 $X=7.805 $Y=1.765
r127 69 70 1.31335 $w=3.67e-07 $l=1e-08 $layer=POLY_cond $X=10.055 $Y=1.557
+ $X2=10.065 $Y2=1.557
r128 67 69 9.85014 $w=3.67e-07 $l=7.5e-08 $layer=POLY_cond $X=9.98 $Y=1.557
+ $X2=10.055 $Y2=1.557
r129 67 68 41.5086 $w=1.7e-07 $l=5.95e-07 $layer=licon1_POLY $count=3 $X=9.98
+ $Y=1.515 $X2=9.98 $Y2=1.515
r130 65 67 49.2507 $w=3.67e-07 $l=3.75e-07 $layer=POLY_cond $X=9.605 $Y=1.557
+ $X2=9.98 $Y2=1.557
r131 64 65 5.25341 $w=3.67e-07 $l=4e-08 $layer=POLY_cond $X=9.565 $Y=1.557
+ $X2=9.605 $Y2=1.557
r132 63 64 53.8474 $w=3.67e-07 $l=4.1e-07 $layer=POLY_cond $X=9.155 $Y=1.557
+ $X2=9.565 $Y2=1.557
r133 62 63 7.22343 $w=3.67e-07 $l=5.5e-08 $layer=POLY_cond $X=9.1 $Y=1.557
+ $X2=9.155 $Y2=1.557
r134 61 62 51.8774 $w=3.67e-07 $l=3.95e-07 $layer=POLY_cond $X=8.705 $Y=1.557
+ $X2=9.1 $Y2=1.557
r135 60 61 4.59673 $w=3.67e-07 $l=3.5e-08 $layer=POLY_cond $X=8.67 $Y=1.557
+ $X2=8.705 $Y2=1.557
r136 59 60 54.5041 $w=3.67e-07 $l=4.15e-07 $layer=POLY_cond $X=8.255 $Y=1.557
+ $X2=8.67 $Y2=1.557
r137 58 59 1.97003 $w=3.67e-07 $l=1.5e-08 $layer=POLY_cond $X=8.24 $Y=1.557
+ $X2=8.255 $Y2=1.557
r138 56 58 39.4005 $w=3.67e-07 $l=3e-07 $layer=POLY_cond $X=7.94 $Y=1.557
+ $X2=8.24 $Y2=1.557
r139 56 57 41.5086 $w=1.7e-07 $l=5.95e-07 $layer=licon1_POLY $count=3 $X=7.94
+ $Y=1.515 $X2=7.94 $Y2=1.515
r140 54 56 17.0736 $w=3.67e-07 $l=1.3e-07 $layer=POLY_cond $X=7.81 $Y=1.557
+ $X2=7.94 $Y2=1.557
r141 53 54 0.656676 $w=3.67e-07 $l=5e-09 $layer=POLY_cond $X=7.805 $Y=1.557
+ $X2=7.81 $Y2=1.557
r142 47 68 9.11234 $w=4.28e-07 $l=3.4e-07 $layer=LI1_cond $X=10.32 $Y=1.565
+ $X2=9.98 $Y2=1.565
r143 46 68 3.75214 $w=4.28e-07 $l=1.4e-07 $layer=LI1_cond $X=9.84 $Y=1.565
+ $X2=9.98 $Y2=1.565
r144 45 46 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=9.36 $Y=1.565
+ $X2=9.84 $Y2=1.565
r145 44 45 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=8.88 $Y=1.565
+ $X2=9.36 $Y2=1.565
r146 43 44 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=8.4 $Y=1.565
+ $X2=8.88 $Y2=1.565
r147 43 57 12.3285 $w=4.28e-07 $l=4.6e-07 $layer=LI1_cond $X=8.4 $Y=1.565
+ $X2=7.94 $Y2=1.565
r148 39 70 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=10.065 $Y=1.35
+ $X2=10.065 $Y2=1.557
r149 39 41 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=10.065 $Y=1.35
+ $X2=10.065 $Y2=0.74
r150 36 69 23.77 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=10.055 $Y=1.765
+ $X2=10.055 $Y2=1.557
r151 36 38 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=10.055 $Y=1.765
+ $X2=10.055 $Y2=2.4
r152 33 65 23.77 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=9.605 $Y=1.765
+ $X2=9.605 $Y2=1.557
r153 33 35 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=9.605 $Y=1.765
+ $X2=9.605 $Y2=2.4
r154 29 64 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=9.565 $Y=1.35
+ $X2=9.565 $Y2=1.557
r155 29 31 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=9.565 $Y=1.35
+ $X2=9.565 $Y2=0.74
r156 26 63 23.77 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=9.155 $Y=1.765
+ $X2=9.155 $Y2=1.557
r157 26 28 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=9.155 $Y=1.765
+ $X2=9.155 $Y2=2.4
r158 22 62 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=9.1 $Y=1.35 $X2=9.1
+ $Y2=1.557
r159 22 24 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=9.1 $Y=1.35 $X2=9.1
+ $Y2=0.74
r160 19 61 23.77 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=8.705 $Y=1.765
+ $X2=8.705 $Y2=1.557
r161 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.705 $Y=1.765
+ $X2=8.705 $Y2=2.4
r162 15 60 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=8.67 $Y=1.35
+ $X2=8.67 $Y2=1.557
r163 15 17 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=8.67 $Y=1.35
+ $X2=8.67 $Y2=0.74
r164 12 59 23.77 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=8.255 $Y=1.765
+ $X2=8.255 $Y2=1.557
r165 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.255 $Y=1.765
+ $X2=8.255 $Y2=2.4
r166 8 58 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=8.24 $Y=1.35 $X2=8.24
+ $Y2=1.557
r167 8 10 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=8.24 $Y=1.35
+ $X2=8.24 $Y2=0.74
r168 4 54 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.81 $Y=1.35 $X2=7.81
+ $Y2=1.557
r169 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.81 $Y=1.35 $X2=7.81
+ $Y2=0.74
r170 1 53 23.77 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=7.805 $Y=1.765
+ $X2=7.805 $Y2=1.557
r171 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.805 $Y=1.765
+ $X2=7.805 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__BUF_16%VPWR 1 2 3 4 5 6 7 8 9 10 11 12 37 39 45 51
+ 57 63 69 75 81 87 89 93 95 99 101 103 108 109 111 112 114 115 117 118 120 121
+ 123 124 126 127 128 129 130 157 166 169 173
c190 87 0 2.68688e-20 $X=7.53 $Y=2.455
c191 81 0 1.71822e-19 $X=6.63 $Y=2.13
c192 75 0 1.71822e-19 $X=5.73 $Y=2.13
c193 63 0 1.71822e-19 $X=3.93 $Y=2.13
c194 57 0 1.71822e-19 $X=3.03 $Y=2.13
c195 45 0 1.71822e-19 $X=1.18 $Y=2.13
r196 172 173 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r197 169 170 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r198 167 170 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=9.36 $Y2=3.33
r199 166 167 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r200 163 164 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r201 161 173 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=10.32 $Y2=3.33
r202 161 170 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=9.36 $Y2=3.33
r203 160 161 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r204 158 169 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.465 $Y=3.33
+ $X2=9.38 $Y2=3.33
r205 158 160 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=9.465 $Y=3.33
+ $X2=9.84 $Y2=3.33
r206 157 172 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=10.195 $Y=3.33
+ $X2=10.377 $Y2=3.33
r207 157 160 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=10.195 $Y=3.33
+ $X2=9.84 $Y2=3.33
r208 156 167 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=8.4 $Y2=3.33
r209 155 156 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r210 153 156 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=7.44 $Y2=3.33
r211 152 153 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r212 150 153 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6.48 $Y2=3.33
r213 149 150 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r214 146 147 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r215 144 147 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r216 143 144 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r217 141 144 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r218 140 141 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r219 138 141 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r220 137 138 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r221 135 138 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r222 135 164 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r223 134 135 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r224 132 163 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.182 $Y2=3.33
r225 132 134 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.72 $Y2=3.33
r226 130 150 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=5.28 $Y=3.33
+ $X2=5.52 $Y2=3.33
r227 130 147 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=5.28 $Y=3.33
+ $X2=4.56 $Y2=3.33
r228 128 155 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=7.445 $Y=3.33
+ $X2=7.44 $Y2=3.33
r229 128 129 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.445 $Y=3.33
+ $X2=7.57 $Y2=3.33
r230 126 152 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=6.545 $Y=3.33
+ $X2=6.48 $Y2=3.33
r231 126 127 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.545 $Y=3.33
+ $X2=6.63 $Y2=3.33
r232 125 155 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=6.715 $Y=3.33
+ $X2=7.44 $Y2=3.33
r233 125 127 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.715 $Y=3.33
+ $X2=6.63 $Y2=3.33
r234 123 149 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=5.645 $Y=3.33
+ $X2=5.52 $Y2=3.33
r235 123 124 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.645 $Y=3.33
+ $X2=5.73 $Y2=3.33
r236 122 152 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=5.815 $Y=3.33
+ $X2=6.48 $Y2=3.33
r237 122 124 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.815 $Y=3.33
+ $X2=5.73 $Y2=3.33
r238 120 146 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=4.745 $Y=3.33
+ $X2=4.56 $Y2=3.33
r239 120 121 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.745 $Y=3.33
+ $X2=4.83 $Y2=3.33
r240 119 149 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=4.915 $Y=3.33
+ $X2=5.52 $Y2=3.33
r241 119 121 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.915 $Y=3.33
+ $X2=4.83 $Y2=3.33
r242 117 143 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=3.845 $Y=3.33
+ $X2=3.6 $Y2=3.33
r243 117 118 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.845 $Y=3.33
+ $X2=3.93 $Y2=3.33
r244 116 146 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=4.015 $Y=3.33
+ $X2=4.56 $Y2=3.33
r245 116 118 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.015 $Y=3.33
+ $X2=3.93 $Y2=3.33
r246 114 140 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.945 $Y=3.33
+ $X2=2.64 $Y2=3.33
r247 114 115 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.945 $Y=3.33
+ $X2=3.03 $Y2=3.33
r248 113 143 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=3.115 $Y=3.33
+ $X2=3.6 $Y2=3.33
r249 113 115 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.115 $Y=3.33
+ $X2=3.03 $Y2=3.33
r250 111 137 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.965 $Y=3.33
+ $X2=1.68 $Y2=3.33
r251 111 112 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.965 $Y=3.33
+ $X2=2.09 $Y2=3.33
r252 110 140 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=2.215 $Y=3.33
+ $X2=2.64 $Y2=3.33
r253 110 112 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.215 $Y=3.33
+ $X2=2.09 $Y2=3.33
r254 108 134 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.095 $Y=3.33
+ $X2=0.72 $Y2=3.33
r255 108 109 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.095 $Y=3.33
+ $X2=1.18 $Y2=3.33
r256 107 137 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=1.265 $Y=3.33
+ $X2=1.68 $Y2=3.33
r257 107 109 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.265 $Y=3.33
+ $X2=1.18 $Y2=3.33
r258 103 106 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=10.32 $Y=2.115
+ $X2=10.32 $Y2=2.815
r259 101 172 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=10.32 $Y=3.245
+ $X2=10.377 $Y2=3.33
r260 101 106 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=10.32 $Y=3.245
+ $X2=10.32 $Y2=2.815
r261 97 169 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.38 $Y=3.245
+ $X2=9.38 $Y2=3.33
r262 97 99 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=9.38 $Y=3.245
+ $X2=9.38 $Y2=2.455
r263 96 166 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.565 $Y=3.33
+ $X2=8.48 $Y2=3.33
r264 95 169 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.295 $Y=3.33
+ $X2=9.38 $Y2=3.33
r265 95 96 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=9.295 $Y=3.33
+ $X2=8.565 $Y2=3.33
r266 91 166 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.48 $Y=3.245
+ $X2=8.48 $Y2=3.33
r267 91 93 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=8.48 $Y=3.245
+ $X2=8.48 $Y2=2.455
r268 90 129 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.695 $Y=3.33
+ $X2=7.57 $Y2=3.33
r269 89 166 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.395 $Y=3.33
+ $X2=8.48 $Y2=3.33
r270 89 90 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=8.395 $Y=3.33
+ $X2=7.695 $Y2=3.33
r271 85 129 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.57 $Y=3.245
+ $X2=7.57 $Y2=3.33
r272 85 87 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=7.57 $Y=3.245
+ $X2=7.57 $Y2=2.455
r273 81 84 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=6.63 $Y=2.13
+ $X2=6.63 $Y2=2.815
r274 79 127 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.63 $Y=3.245
+ $X2=6.63 $Y2=3.33
r275 79 84 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=6.63 $Y=3.245
+ $X2=6.63 $Y2=2.815
r276 75 78 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=5.73 $Y=2.13
+ $X2=5.73 $Y2=2.81
r277 73 124 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.73 $Y=3.245
+ $X2=5.73 $Y2=3.33
r278 73 78 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=5.73 $Y=3.245
+ $X2=5.73 $Y2=2.81
r279 69 72 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=4.83 $Y=2.13
+ $X2=4.83 $Y2=2.815
r280 67 121 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.83 $Y=3.245
+ $X2=4.83 $Y2=3.33
r281 67 72 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=4.83 $Y=3.245
+ $X2=4.83 $Y2=2.815
r282 63 66 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.93 $Y=2.13
+ $X2=3.93 $Y2=2.81
r283 61 118 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.93 $Y=3.245
+ $X2=3.93 $Y2=3.33
r284 61 66 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=3.93 $Y=3.245
+ $X2=3.93 $Y2=2.81
r285 57 60 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=3.03 $Y=2.13
+ $X2=3.03 $Y2=2.815
r286 55 115 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.03 $Y=3.245
+ $X2=3.03 $Y2=3.33
r287 55 60 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=3.03 $Y=3.245
+ $X2=3.03 $Y2=2.815
r288 51 54 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=2.09 $Y=2.13
+ $X2=2.09 $Y2=2.81
r289 49 112 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.09 $Y=3.245
+ $X2=2.09 $Y2=3.33
r290 49 54 20.0525 $w=2.48e-07 $l=4.35e-07 $layer=LI1_cond $X=2.09 $Y=3.245
+ $X2=2.09 $Y2=2.81
r291 45 48 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.18 $Y=2.13
+ $X2=1.18 $Y2=2.81
r292 43 109 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.18 $Y=3.245
+ $X2=1.18 $Y2=3.33
r293 43 48 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=1.18 $Y=3.245
+ $X2=1.18 $Y2=2.81
r294 39 42 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=0.24 $Y=1.985
+ $X2=0.24 $Y2=2.815
r295 37 163 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.182 $Y2=3.33
r296 37 42 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.24 $Y2=2.815
r297 12 106 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=10.13
+ $Y=1.84 $X2=10.28 $Y2=2.815
r298 12 103 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=10.13
+ $Y=1.84 $X2=10.28 $Y2=2.115
r299 11 99 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=9.23
+ $Y=1.84 $X2=9.38 $Y2=2.455
r300 10 93 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=8.33
+ $Y=1.84 $X2=8.48 $Y2=2.455
r301 9 87 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=7.38
+ $Y=1.84 $X2=7.53 $Y2=2.455
r302 8 84 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=6.48
+ $Y=1.84 $X2=6.63 $Y2=2.815
r303 8 81 400 $w=1.7e-07 $l=3.57211e-07 $layer=licon1_PDIFF $count=1 $X=6.48
+ $Y=1.84 $X2=6.63 $Y2=2.13
r304 7 78 400 $w=1.7e-07 $l=1.04231e-06 $layer=licon1_PDIFF $count=1 $X=5.58
+ $Y=1.84 $X2=5.73 $Y2=2.81
r305 7 75 400 $w=1.7e-07 $l=3.57211e-07 $layer=licon1_PDIFF $count=1 $X=5.58
+ $Y=1.84 $X2=5.73 $Y2=2.13
r306 6 72 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=4.68
+ $Y=1.84 $X2=4.83 $Y2=2.815
r307 6 69 400 $w=1.7e-07 $l=3.57211e-07 $layer=licon1_PDIFF $count=1 $X=4.68
+ $Y=1.84 $X2=4.83 $Y2=2.13
r308 5 66 400 $w=1.7e-07 $l=1.04231e-06 $layer=licon1_PDIFF $count=1 $X=3.78
+ $Y=1.84 $X2=3.93 $Y2=2.81
r309 5 63 400 $w=1.7e-07 $l=3.57211e-07 $layer=licon1_PDIFF $count=1 $X=3.78
+ $Y=1.84 $X2=3.93 $Y2=2.13
r310 4 60 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.88
+ $Y=1.84 $X2=3.03 $Y2=2.815
r311 4 57 400 $w=1.7e-07 $l=3.57211e-07 $layer=licon1_PDIFF $count=1 $X=2.88
+ $Y=1.84 $X2=3.03 $Y2=2.13
r312 3 54 400 $w=1.7e-07 $l=1.06532e-06 $layer=licon1_PDIFF $count=1 $X=1.93
+ $Y=1.84 $X2=2.13 $Y2=2.81
r313 3 51 400 $w=1.7e-07 $l=3.76962e-07 $layer=licon1_PDIFF $count=1 $X=1.93
+ $Y=1.84 $X2=2.13 $Y2=2.13
r314 2 48 400 $w=1.7e-07 $l=1.04231e-06 $layer=licon1_PDIFF $count=1 $X=1.03
+ $Y=1.84 $X2=1.18 $Y2=2.81
r315 2 45 400 $w=1.7e-07 $l=3.57211e-07 $layer=licon1_PDIFF $count=1 $X=1.03
+ $Y=1.84 $X2=1.18 $Y2=2.13
r316 1 42 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r317 1 39 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_LS__BUF_16%X 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 51
+ 55 61 67 71 75 77 79 83 84 85 86 87 90 92 94 97 107 117 124 131 138 145 147
+ 152 153
c259 147 0 1.43649e-19 $X=7.11 $Y=2.035
c260 145 0 1.0264e-19 $X=7.08 $Y=1.985
c261 131 0 1.02687e-19 $X=5.28 $Y=1.985
c262 117 0 1.02631e-19 $X=2.58 $Y=1.985
r263 152 155 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.385 $Y=2.035
+ $X2=4.385 $Y2=2.035
r264 152 153 5.66838 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=4.38 $Y=1.985
+ $X2=4.38 $Y2=1.9
r265 145 149 36.0954 $w=2.63e-07 $l=8.3e-07 $layer=LI1_cond $X=7.112 $Y=1.985
+ $X2=7.112 $Y2=2.815
r266 145 147 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.11 $Y=2.035
+ $X2=7.11 $Y2=2.035
r267 140 147 0.596692 $w=2.3e-07 $l=9.3e-07 $layer=MET1_cond $X=6.18 $Y=2.035
+ $X2=7.11 $Y2=2.035
r268 138 142 35.427 $w=2.68e-07 $l=8.3e-07 $layer=LI1_cond $X=6.195 $Y=1.985
+ $X2=6.195 $Y2=2.815
r269 138 140 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.18 $Y=2.035
+ $X2=6.18 $Y2=2.035
r270 133 140 0.577444 $w=2.3e-07 $l=9e-07 $layer=MET1_cond $X=5.28 $Y=2.035
+ $X2=6.18 $Y2=2.035
r271 133 155 0.574236 $w=2.3e-07 $l=8.95e-07 $layer=MET1_cond $X=5.28 $Y=2.035
+ $X2=4.385 $Y2=2.035
r272 131 135 32.4247 $w=2.93e-07 $l=8.3e-07 $layer=LI1_cond $X=5.262 $Y=1.985
+ $X2=5.262 $Y2=2.815
r273 131 133 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.28 $Y=2.035
+ $X2=5.28 $Y2=2.035
r274 124 128 37.5109 $w=2.53e-07 $l=8.3e-07 $layer=LI1_cond $X=3.437 $Y=1.985
+ $X2=3.437 $Y2=2.815
r275 124 126 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.445 $Y=2.035
+ $X2=3.445 $Y2=2.035
r276 119 126 0.571028 $w=2.3e-07 $l=8.9e-07 $layer=MET1_cond $X=2.555 $Y=2.035
+ $X2=3.445 $Y2=2.035
r277 117 121 36.7895 $w=2.58e-07 $l=8.3e-07 $layer=LI1_cond $X=2.545 $Y=1.985
+ $X2=2.545 $Y2=2.815
r278 117 119 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.555 $Y=2.035
+ $X2=2.555 $Y2=2.035
r279 112 119 0.612732 $w=2.3e-07 $l=9.55e-07 $layer=MET1_cond $X=1.6 $Y=2.035
+ $X2=2.555 $Y2=2.035
r280 110 114 37.5109 $w=2.53e-07 $l=8.3e-07 $layer=LI1_cond $X=1.592 $Y=1.985
+ $X2=1.592 $Y2=2.815
r281 110 112 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.6 $Y=2.035
+ $X2=1.6 $Y2=2.035
r282 107 110 66.435 $w=2.53e-07 $l=1.47e-06 $layer=LI1_cond $X=1.592 $Y=0.515
+ $X2=1.592 $Y2=1.985
r283 102 112 0.564612 $w=2.3e-07 $l=8.8e-07 $layer=MET1_cond $X=0.72 $Y=2.035
+ $X2=1.6 $Y2=2.035
r284 100 104 37.5109 $w=2.53e-07 $l=8.3e-07 $layer=LI1_cond $X=0.687 $Y=1.985
+ $X2=0.687 $Y2=2.815
r285 100 102 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=2.035
+ $X2=0.72 $Y2=2.035
r286 97 100 66.435 $w=2.53e-07 $l=1.47e-06 $layer=LI1_cond $X=0.687 $Y=0.515
+ $X2=0.687 $Y2=1.985
r287 94 155 0.301554 $w=2.3e-07 $l=4.7e-07 $layer=MET1_cond $X=3.915 $Y=2.035
+ $X2=4.385 $Y2=2.035
r288 94 126 0.301554 $w=2.3e-07 $l=4.7e-07 $layer=MET1_cond $X=3.915 $Y=2.035
+ $X2=3.445 $Y2=2.035
r289 93 145 26.2235 $w=2.63e-07 $l=6.03e-07 $layer=LI1_cond $X=7.112 $Y=1.382
+ $X2=7.112 $Y2=1.985
r290 92 138 36.494 $w=2.68e-07 $l=8.55e-07 $layer=LI1_cond $X=6.195 $Y=1.13
+ $X2=6.195 $Y2=1.985
r291 90 131 23.8302 $w=2.93e-07 $l=6.1e-07 $layer=LI1_cond $X=5.262 $Y=1.375
+ $X2=5.262 $Y2=1.985
r292 89 90 5.22441 $w=3.73e-07 $l=1.7e-07 $layer=LI1_cond $X=5.222 $Y=1.205
+ $X2=5.222 $Y2=1.375
r293 87 153 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=4.3 $Y=1.13
+ $X2=4.3 $Y2=1.9
r294 85 124 1.71737 $w=2.53e-07 $l=3.8e-08 $layer=LI1_cond $X=3.437 $Y=1.947
+ $X2=3.437 $Y2=1.985
r295 85 86 7.02311 $w=2.53e-07 $l=1.27e-07 $layer=LI1_cond $X=3.437 $Y=1.947
+ $X2=3.437 $Y2=1.82
r296 84 86 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.395 $Y=1.13
+ $X2=3.395 $Y2=1.82
r297 83 117 27.9246 $w=2.58e-07 $l=6.3e-07 $layer=LI1_cond $X=2.545 $Y=1.355
+ $X2=2.545 $Y2=1.985
r298 82 83 7.39303 $w=2.63e-07 $l=1.7e-07 $layer=LI1_cond $X=2.51 $Y=1.185
+ $X2=2.51 $Y2=1.355
r299 77 93 12.2 $w=2.57e-07 $l=2.6342e-07 $layer=LI1_cond $X=7.125 $Y=1.125
+ $X2=7.112 $Y2=1.382
r300 77 79 28.1196 $w=2.48e-07 $l=6.1e-07 $layer=LI1_cond $X=7.125 $Y=1.125
+ $X2=7.125 $Y2=0.515
r301 73 92 6.17723 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=6.165 $Y=0.965
+ $X2=6.165 $Y2=1.13
r302 73 75 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=6.165 $Y=0.965
+ $X2=6.165 $Y2=0.515
r303 71 89 26.9554 $w=2.93e-07 $l=6.9e-07 $layer=LI1_cond $X=5.182 $Y=0.515
+ $X2=5.182 $Y2=1.205
r304 65 152 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=4.38 $Y=2.065
+ $X2=4.38 $Y2=1.985
r305 65 67 26.1919 $w=3.28e-07 $l=7.5e-07 $layer=LI1_cond $X=4.38 $Y=2.065
+ $X2=4.38 $Y2=2.815
r306 59 87 9.39714 $w=3.83e-07 $l=1.92e-07 $layer=LI1_cond $X=4.192 $Y=0.938
+ $X2=4.192 $Y2=1.13
r307 59 61 12.6619 $w=3.83e-07 $l=4.23e-07 $layer=LI1_cond $X=4.192 $Y=0.938
+ $X2=4.192 $Y2=0.515
r308 53 84 7.14225 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=3.35 $Y=1 $X2=3.35
+ $Y2=1.13
r309 53 55 21.4975 $w=2.58e-07 $l=4.85e-07 $layer=LI1_cond $X=3.35 $Y=1 $X2=3.35
+ $Y2=0.515
r310 51 82 29.1372 $w=2.63e-07 $l=6.7e-07 $layer=LI1_cond $X=2.477 $Y=0.515
+ $X2=2.477 $Y2=1.185
r311 16 149 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=6.93
+ $Y=1.84 $X2=7.08 $Y2=2.815
r312 16 145 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=6.93
+ $Y=1.84 $X2=7.08 $Y2=1.985
r313 15 142 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=6.03
+ $Y=1.84 $X2=6.18 $Y2=2.815
r314 15 138 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=6.03
+ $Y=1.84 $X2=6.18 $Y2=1.985
r315 14 135 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=5.13
+ $Y=1.84 $X2=5.28 $Y2=2.815
r316 14 131 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=5.13
+ $Y=1.84 $X2=5.28 $Y2=1.985
r317 13 152 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=4.23
+ $Y=1.84 $X2=4.38 $Y2=1.985
r318 13 67 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=4.23
+ $Y=1.84 $X2=4.38 $Y2=2.815
r319 12 128 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=3.33
+ $Y=1.84 $X2=3.48 $Y2=2.815
r320 12 124 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=3.33
+ $Y=1.84 $X2=3.48 $Y2=1.985
r321 11 121 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.43
+ $Y=1.84 $X2=2.58 $Y2=2.815
r322 11 117 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.43
+ $Y=1.84 $X2=2.58 $Y2=1.985
r323 10 114 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.48
+ $Y=1.84 $X2=1.63 $Y2=2.815
r324 10 110 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.48
+ $Y=1.84 $X2=1.63 $Y2=1.985
r325 9 104 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.84 $X2=0.73 $Y2=2.815
r326 9 100 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.84 $X2=0.73 $Y2=1.985
r327 8 79 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.025
+ $Y=0.37 $X2=7.165 $Y2=0.515
r328 7 75 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.025
+ $Y=0.37 $X2=6.165 $Y2=0.515
r329 6 71 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.025
+ $Y=0.37 $X2=5.165 $Y2=0.515
r330 5 61 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.025
+ $Y=0.37 $X2=4.165 $Y2=0.515
r331 4 55 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.165
+ $Y=0.37 $X2=3.305 $Y2=0.515
r332 3 51 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.305
+ $Y=0.37 $X2=2.445 $Y2=0.515
r333 2 107 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.445
+ $Y=0.37 $X2=1.585 $Y2=0.515
r334 1 97 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.585
+ $Y=0.37 $X2=0.725 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__BUF_16%VGND 1 2 3 4 5 6 7 8 9 10 11 12 37 39 43 47
+ 51 55 57 61 63 67 71 73 77 81 85 87 89 92 93 95 96 97 98 99 100 101 103 122
+ 127 132 141 144 147 150 153 156 160
c185 89 0 1.18608e-19 $X=10.28 $Y=0.515
r186 159 160 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r187 156 157 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r188 153 154 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r189 150 151 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r190 147 148 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r191 144 145 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r192 141 142 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r193 138 139 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r194 136 160 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=10.32 $Y2=0
r195 136 157 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=9.36 $Y2=0
r196 135 136 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0
+ $X2=9.84 $Y2=0
r197 133 156 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.48 $Y=0
+ $X2=9.315 $Y2=0
r198 133 135 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=9.48 $Y=0
+ $X2=9.84 $Y2=0
r199 132 159 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=10.115 $Y=0
+ $X2=10.337 $Y2=0
r200 132 135 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=10.115 $Y=0
+ $X2=9.84 $Y2=0
r201 131 157 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0
+ $X2=9.36 $Y2=0
r202 131 154 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0
+ $X2=8.4 $Y2=0
r203 130 131 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r204 128 153 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.62 $Y=0
+ $X2=8.455 $Y2=0
r205 128 130 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=8.62 $Y=0
+ $X2=8.88 $Y2=0
r206 127 156 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.15 $Y=0
+ $X2=9.315 $Y2=0
r207 127 130 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=9.15 $Y=0 $X2=8.88
+ $Y2=0
r208 126 154 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0
+ $X2=8.4 $Y2=0
r209 126 151 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0
+ $X2=7.44 $Y2=0
r210 125 126 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r211 123 150 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.76 $Y=0
+ $X2=7.595 $Y2=0
r212 123 125 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=7.76 $Y=0
+ $X2=7.92 $Y2=0
r213 122 153 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.29 $Y=0
+ $X2=8.455 $Y2=0
r214 122 125 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=8.29 $Y=0 $X2=7.92
+ $Y2=0
r215 121 151 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=0
+ $X2=7.44 $Y2=0
r216 121 148 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=0
+ $X2=5.52 $Y2=0
r217 120 121 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r218 118 147 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.83 $Y=0
+ $X2=5.665 $Y2=0
r219 118 120 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=5.83 $Y=0
+ $X2=6.48 $Y2=0
r220 117 145 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0
+ $X2=4.56 $Y2=0
r221 116 117 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r222 114 117 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=3.6 $Y2=0
r223 113 114 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r224 111 114 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0
+ $X2=2.64 $Y2=0
r225 111 142 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0
+ $X2=1.2 $Y2=0
r226 110 111 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0
+ $X2=1.68 $Y2=0
r227 108 141 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=1.285 $Y=0
+ $X2=1.137 $Y2=0
r228 108 110 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.285 $Y=0
+ $X2=1.68 $Y2=0
r229 107 142 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0
+ $X2=1.2 $Y2=0
r230 107 139 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0
+ $X2=0.24 $Y2=0
r231 106 107 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0
+ $X2=0.72 $Y2=0
r232 104 138 3.99177 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.38 $Y=0 $X2=0.19
+ $Y2=0
r233 104 106 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.38 $Y=0
+ $X2=0.72 $Y2=0
r234 103 141 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=0.99 $Y=0
+ $X2=1.137 $Y2=0
r235 103 106 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.99 $Y=0 $X2=0.72
+ $Y2=0
r236 101 148 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=5.28 $Y=0
+ $X2=5.52 $Y2=0
r237 101 145 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=5.28 $Y=0
+ $X2=4.56 $Y2=0
r238 99 120 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=6.5 $Y=0 $X2=6.48
+ $Y2=0
r239 99 100 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.5 $Y=0 $X2=6.665
+ $Y2=0
r240 97 116 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=3.65 $Y=0 $X2=3.6
+ $Y2=0
r241 97 98 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.65 $Y=0 $X2=3.735
+ $Y2=0
r242 95 113 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=2.79 $Y=0 $X2=2.64
+ $Y2=0
r243 95 96 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.79 $Y=0 $X2=2.875
+ $Y2=0
r244 94 116 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=2.96 $Y=0 $X2=3.6
+ $Y2=0
r245 94 96 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.96 $Y=0 $X2=2.875
+ $Y2=0
r246 92 110 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.895 $Y=0
+ $X2=1.68 $Y2=0
r247 92 93 6.01921 $w=1.7e-07 $l=1.02e-07 $layer=LI1_cond $X=1.895 $Y=0
+ $X2=1.997 $Y2=0
r248 91 113 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=2.1 $Y=0 $X2=2.64
+ $Y2=0
r249 91 93 6.01921 $w=1.7e-07 $l=1.03e-07 $layer=LI1_cond $X=2.1 $Y=0 $X2=1.997
+ $Y2=0
r250 87 159 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=10.28 $Y=0.085
+ $X2=10.337 $Y2=0
r251 87 89 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=10.28 $Y=0.085
+ $X2=10.28 $Y2=0.515
r252 83 156 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.315 $Y=0.085
+ $X2=9.315 $Y2=0
r253 83 85 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=9.315 $Y=0.085
+ $X2=9.315 $Y2=0.675
r254 79 153 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.455 $Y=0.085
+ $X2=8.455 $Y2=0
r255 79 81 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=8.455 $Y=0.085
+ $X2=8.455 $Y2=0.675
r256 75 150 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.595 $Y=0.085
+ $X2=7.595 $Y2=0
r257 75 77 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=7.595 $Y=0.085
+ $X2=7.595 $Y2=0.675
r258 74 100 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.83 $Y=0
+ $X2=6.665 $Y2=0
r259 73 150 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.43 $Y=0
+ $X2=7.595 $Y2=0
r260 73 74 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=7.43 $Y=0 $X2=6.83
+ $Y2=0
r261 69 100 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.665 $Y=0.085
+ $X2=6.665 $Y2=0
r262 69 71 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=6.665 $Y=0.085
+ $X2=6.665 $Y2=0.495
r263 65 147 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.665 $Y=0.085
+ $X2=5.665 $Y2=0
r264 65 67 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=5.665 $Y=0.085
+ $X2=5.665 $Y2=0.495
r265 64 144 7.54988 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=4.83 $Y=0
+ $X2=4.692 $Y2=0
r266 63 147 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.5 $Y=0 $X2=5.665
+ $Y2=0
r267 63 64 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.5 $Y=0 $X2=4.83
+ $Y2=0
r268 59 144 0.316938 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=4.692 $Y=0.085
+ $X2=4.692 $Y2=0
r269 59 61 17.1819 $w=2.73e-07 $l=4.1e-07 $layer=LI1_cond $X=4.692 $Y=0.085
+ $X2=4.692 $Y2=0.495
r270 58 98 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.82 $Y=0 $X2=3.735
+ $Y2=0
r271 57 144 7.54988 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=4.555 $Y=0
+ $X2=4.692 $Y2=0
r272 57 58 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=4.555 $Y=0
+ $X2=3.82 $Y2=0
r273 53 98 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.735 $Y=0.085
+ $X2=3.735 $Y2=0
r274 53 55 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=3.735 $Y=0.085
+ $X2=3.735 $Y2=0.495
r275 49 96 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.875 $Y=0.085
+ $X2=2.875 $Y2=0
r276 49 51 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=2.875 $Y=0.085
+ $X2=2.875 $Y2=0.495
r277 45 93 0.677923 $w=2.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.997 $Y=0.085
+ $X2=1.997 $Y2=0
r278 45 47 22.1818 $w=2.03e-07 $l=4.1e-07 $layer=LI1_cond $X=1.997 $Y=0.085
+ $X2=1.997 $Y2=0.495
r279 41 141 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=1.137 $Y=0.085
+ $X2=1.137 $Y2=0
r280 41 43 16.017 $w=2.93e-07 $l=4.1e-07 $layer=LI1_cond $X=1.137 $Y=0.085
+ $X2=1.137 $Y2=0.495
r281 37 138 3.1514 $w=2.5e-07 $l=1.12916e-07 $layer=LI1_cond $X=0.255 $Y=0.085
+ $X2=0.19 $Y2=0
r282 37 39 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.255 $Y=0.085
+ $X2=0.255 $Y2=0.515
r283 12 89 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.14
+ $Y=0.37 $X2=10.28 $Y2=0.515
r284 11 85 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=9.175
+ $Y=0.37 $X2=9.315 $Y2=0.675
r285 10 81 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=8.315
+ $Y=0.37 $X2=8.455 $Y2=0.675
r286 9 77 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=7.455
+ $Y=0.37 $X2=7.595 $Y2=0.675
r287 8 71 91 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=2 $X=6.455
+ $Y=0.37 $X2=6.665 $Y2=0.495
r288 7 67 91 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=2 $X=5.455
+ $Y=0.37 $X2=5.665 $Y2=0.495
r289 6 61 91 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=2 $X=4.455
+ $Y=0.37 $X2=4.665 $Y2=0.495
r290 5 55 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=3.595
+ $Y=0.37 $X2=3.735 $Y2=0.495
r291 4 51 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=2.735
+ $Y=0.37 $X2=2.875 $Y2=0.495
r292 3 47 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.875
+ $Y=0.37 $X2=2.015 $Y2=0.495
r293 2 43 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.015
+ $Y=0.37 $X2=1.155 $Y2=0.495
r294 1 39 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.15
+ $Y=0.37 $X2=0.295 $Y2=0.515
.ends

