# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ls__sdfrtn_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ls__sdfrtn_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  13.92000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.780000 1.980000 2.120000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.546900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.475000 0.350000 13.805000 2.980000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.411000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  3.405000 1.355000  3.735000 2.025000 ;
        RECT  7.685000 1.470000  8.035000 1.800000 ;
        RECT 10.995000 1.210000 11.395000 1.540000 ;
        RECT 11.195000 1.540000 11.395000 1.780000 ;
      LAYER mcon ;
        RECT  3.515000 1.580000  3.685000 1.750000 ;
        RECT  7.835000 1.580000  8.005000 1.750000 ;
        RECT 11.195000 1.580000 11.365000 1.750000 ;
      LAYER met1 ;
        RECT  3.455000 1.550000  3.745000 1.595000 ;
        RECT  3.455000 1.595000 11.425000 1.735000 ;
        RECT  3.455000 1.735000  3.745000 1.780000 ;
        RECT  7.775000 1.550000  8.065000 1.595000 ;
        RECT  7.775000 1.735000  8.065000 1.780000 ;
        RECT 11.135000 1.550000 11.425000 1.595000 ;
        RECT 11.135000 1.735000 11.425000 1.780000 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.800000 1.525000 3.235000 2.150000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 1.410000 2.045000 1.580000 ;
        RECT 0.535000 1.580000 0.865000 2.080000 ;
        RECT 1.875000 0.955000 2.550000 1.410000 ;
    END
  END SCE
  PIN CLK_N
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 4.275000 1.210000 4.675000 1.550000 ;
    END
  END CLK_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 13.920000 0.085000 ;
        RECT  0.615000  0.085000  0.945000 0.880000 ;
        RECT  3.575000  0.085000  4.065000 0.360000 ;
        RECT  4.805000  0.085000  5.165000 0.360000 ;
        RECT  7.890000  0.085000  8.220000 0.620000 ;
        RECT 10.730000  0.085000 11.200000 0.680000 ;
        RECT 12.975000  0.085000 13.305000 1.130000 ;
      LAYER mcon ;
        RECT  0.155000 -0.085000  0.325000 0.085000 ;
        RECT  0.635000 -0.085000  0.805000 0.085000 ;
        RECT  1.115000 -0.085000  1.285000 0.085000 ;
        RECT  1.595000 -0.085000  1.765000 0.085000 ;
        RECT  2.075000 -0.085000  2.245000 0.085000 ;
        RECT  2.555000 -0.085000  2.725000 0.085000 ;
        RECT  3.035000 -0.085000  3.205000 0.085000 ;
        RECT  3.515000 -0.085000  3.685000 0.085000 ;
        RECT  3.995000 -0.085000  4.165000 0.085000 ;
        RECT  4.475000 -0.085000  4.645000 0.085000 ;
        RECT  4.955000 -0.085000  5.125000 0.085000 ;
        RECT  5.435000 -0.085000  5.605000 0.085000 ;
        RECT  5.915000 -0.085000  6.085000 0.085000 ;
        RECT  6.395000 -0.085000  6.565000 0.085000 ;
        RECT  6.875000 -0.085000  7.045000 0.085000 ;
        RECT  7.355000 -0.085000  7.525000 0.085000 ;
        RECT  7.835000 -0.085000  8.005000 0.085000 ;
        RECT  8.315000 -0.085000  8.485000 0.085000 ;
        RECT  8.795000 -0.085000  8.965000 0.085000 ;
        RECT  9.275000 -0.085000  9.445000 0.085000 ;
        RECT  9.755000 -0.085000  9.925000 0.085000 ;
        RECT 10.235000 -0.085000 10.405000 0.085000 ;
        RECT 10.715000 -0.085000 10.885000 0.085000 ;
        RECT 11.195000 -0.085000 11.365000 0.085000 ;
        RECT 11.675000 -0.085000 11.845000 0.085000 ;
        RECT 12.155000 -0.085000 12.325000 0.085000 ;
        RECT 12.635000 -0.085000 12.805000 0.085000 ;
        RECT 13.115000 -0.085000 13.285000 0.085000 ;
        RECT 13.595000 -0.085000 13.765000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 13.920000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 3.245000 13.920000 3.415000 ;
        RECT  0.565000 2.630000  0.895000 3.245000 ;
        RECT  2.815000 2.970000  3.145000 3.245000 ;
        RECT  4.780000 2.500000  5.110000 3.245000 ;
        RECT  7.225000 2.380000  7.395000 3.245000 ;
        RECT  8.295000 2.310000  8.625000 3.245000 ;
        RECT 10.605000 2.650000 11.210000 3.245000 ;
        RECT 11.880000 2.630000 12.210000 3.245000 ;
        RECT 12.975000 1.820000 13.305000 3.245000 ;
      LAYER mcon ;
        RECT  0.155000 3.245000  0.325000 3.415000 ;
        RECT  0.635000 3.245000  0.805000 3.415000 ;
        RECT  1.115000 3.245000  1.285000 3.415000 ;
        RECT  1.595000 3.245000  1.765000 3.415000 ;
        RECT  2.075000 3.245000  2.245000 3.415000 ;
        RECT  2.555000 3.245000  2.725000 3.415000 ;
        RECT  3.035000 3.245000  3.205000 3.415000 ;
        RECT  3.515000 3.245000  3.685000 3.415000 ;
        RECT  3.995000 3.245000  4.165000 3.415000 ;
        RECT  4.475000 3.245000  4.645000 3.415000 ;
        RECT  4.955000 3.245000  5.125000 3.415000 ;
        RECT  5.435000 3.245000  5.605000 3.415000 ;
        RECT  5.915000 3.245000  6.085000 3.415000 ;
        RECT  6.395000 3.245000  6.565000 3.415000 ;
        RECT  6.875000 3.245000  7.045000 3.415000 ;
        RECT  7.355000 3.245000  7.525000 3.415000 ;
        RECT  7.835000 3.245000  8.005000 3.415000 ;
        RECT  8.315000 3.245000  8.485000 3.415000 ;
        RECT  8.795000 3.245000  8.965000 3.415000 ;
        RECT  9.275000 3.245000  9.445000 3.415000 ;
        RECT  9.755000 3.245000  9.925000 3.415000 ;
        RECT 10.235000 3.245000 10.405000 3.415000 ;
        RECT 10.715000 3.245000 10.885000 3.415000 ;
        RECT 11.195000 3.245000 11.365000 3.415000 ;
        RECT 11.675000 3.245000 11.845000 3.415000 ;
        RECT 12.155000 3.245000 12.325000 3.415000 ;
        RECT 12.635000 3.245000 12.805000 3.415000 ;
        RECT 13.115000 3.245000 13.285000 3.415000 ;
        RECT 13.595000 3.245000 13.765000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 13.920000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.115000 0.420000  0.445000 1.050000 ;
      RECT  0.115000 1.050000  1.620000 1.240000 ;
      RECT  0.115000 1.240000  0.365000 2.290000 ;
      RECT  0.115000 2.290000  2.545000 2.460000 ;
      RECT  0.115000 2.460000  0.365000 2.980000 ;
      RECT  1.165000 0.255000  3.390000 0.425000 ;
      RECT  1.165000 0.425000  1.495000 0.765000 ;
      RECT  1.290000 0.935000  1.620000 1.050000 ;
      RECT  1.405000 2.630000  3.680000 2.800000 ;
      RECT  1.405000 2.800000  2.220000 2.960000 ;
      RECT  1.955000 0.595000  2.890000 0.765000 ;
      RECT  2.215000 1.580000  2.545000 2.290000 ;
      RECT  2.720000 0.765000  2.890000 1.015000 ;
      RECT  2.720000 1.015000  4.075000 1.185000 ;
      RECT  3.060000 0.425000  3.390000 0.845000 ;
      RECT  3.430000 2.195000  6.115000 2.330000 ;
      RECT  3.430000 2.330000  4.720000 2.340000 ;
      RECT  3.430000 2.340000  4.700000 2.350000 ;
      RECT  3.430000 2.350000  4.645000 2.395000 ;
      RECT  3.430000 2.395000  3.680000 2.630000 ;
      RECT  3.430000 2.800000  3.680000 2.980000 ;
      RECT  3.905000 0.530000  6.155000 0.700000 ;
      RECT  3.905000 0.700000  4.075000 1.015000 ;
      RECT  3.905000 1.185000  4.075000 2.170000 ;
      RECT  3.905000 2.170000  6.115000 2.195000 ;
      RECT  4.245000 0.870000  5.165000 1.040000 ;
      RECT  4.255000 1.820000  5.030000 1.990000 ;
      RECT  4.255000 1.990000  4.600000 2.000000 ;
      RECT  4.660000 2.160000  6.115000 2.170000 ;
      RECT  4.845000 1.040000  5.165000 1.235000 ;
      RECT  4.845000 1.235000  5.255000 1.605000 ;
      RECT  4.845000 1.605000  5.030000 1.820000 ;
      RECT  5.230000 1.775000  6.715000 1.990000 ;
      RECT  5.345000 0.870000  5.675000 1.085000 ;
      RECT  5.425000 1.085000  5.675000 1.265000 ;
      RECT  5.425000 1.265000  6.495000 1.465000 ;
      RECT  5.425000 1.465000  5.675000 1.735000 ;
      RECT  5.425000 1.735000  6.715000 1.775000 ;
      RECT  5.855000 2.330000  6.115000 2.735000 ;
      RECT  5.905000 0.700000  6.155000 1.095000 ;
      RECT  6.285000 2.235000  7.055000 2.445000 ;
      RECT  6.285000 2.445000  6.570000 2.735000 ;
      RECT  6.325000 0.255000  7.720000 0.545000 ;
      RECT  6.325000 0.545000  6.495000 1.265000 ;
      RECT  6.495000 1.990000  6.715000 2.065000 ;
      RECT  6.665000 0.725000  7.055000 1.095000 ;
      RECT  6.885000 1.095000  7.055000 2.040000 ;
      RECT  6.885000 2.040000  8.520000 2.140000 ;
      RECT  6.885000 2.140000  7.950000 2.210000 ;
      RECT  6.885000 2.210000  7.055000 2.235000 ;
      RECT  7.225000 1.130000  9.010000 1.300000 ;
      RECT  7.225000 1.300000  7.475000 1.870000 ;
      RECT  7.495000 0.545000  7.720000 0.790000 ;
      RECT  7.495000 0.790000  9.825000 0.960000 ;
      RECT  7.575000 2.210000  7.950000 2.735000 ;
      RECT  7.645000 1.970000  8.520000 2.040000 ;
      RECT  8.225000 1.470000  8.520000 1.970000 ;
      RECT  8.690000 1.300000  8.860000 1.970000 ;
      RECT  8.690000 1.970000  9.565000 2.140000 ;
      RECT  8.795000 2.140000  9.565000 2.980000 ;
      RECT  9.030000 1.470000 10.395000 1.540000 ;
      RECT  9.030000 1.540000  9.350000 1.800000 ;
      RECT  9.180000 1.370000 10.395000 1.470000 ;
      RECT  9.190000 0.290000 10.165000 0.620000 ;
      RECT  9.495000 0.960000  9.825000 1.200000 ;
      RECT  9.735000 1.710000 11.025000 1.880000 ;
      RECT  9.735000 1.880000 10.065000 2.980000 ;
      RECT  9.995000 0.620000 10.165000 0.870000 ;
      RECT  9.995000 0.870000 11.895000 1.040000 ;
      RECT 10.065000 1.225000 10.395000 1.370000 ;
      RECT 10.435000 2.050000 10.685000 2.290000 ;
      RECT 10.435000 2.290000 12.235000 2.460000 ;
      RECT 10.855000 1.880000 11.025000 1.950000 ;
      RECT 10.855000 1.950000 11.895000 2.120000 ;
      RECT 11.380000 2.460000 11.710000 2.980000 ;
      RECT 11.565000 1.040000 11.895000 1.950000 ;
      RECT 11.690000 0.450000 12.235000 0.700000 ;
      RECT 12.065000 0.700000 12.235000 2.290000 ;
      RECT 12.440000 0.350000 12.795000 1.355000 ;
      RECT 12.440000 1.355000 12.810000 1.685000 ;
      RECT 12.440000 1.685000 12.795000 2.980000 ;
  END
END sky130_fd_sc_ls__sdfrtn_1
