# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ls__dlrtp_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ls__dlrtp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.720000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.208500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.300000 0.375000 1.780000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.100000 0.350000 6.635000 0.840000 ;
        RECT 6.275000 1.820000 6.635000 2.980000 ;
        RECT 6.465000 0.840000 6.635000 1.820000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.435000 1.350000 5.765000 1.780000 ;
    END
  END RESET_B
  PIN GATE
    ANTENNAGATEAREA  0.237000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.930000 1.450000 1.285000 1.780000 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 6.720000 0.085000 ;
        RECT 0.885000  0.085000 1.055000 1.130000 ;
        RECT 2.295000  0.085000 2.680000 0.600000 ;
        RECT 4.210000  0.085000 4.540000 0.810000 ;
        RECT 5.590000  0.085000 5.920000 0.840000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
        RECT 6.395000 -0.085000 6.565000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.720000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 6.720000 3.415000 ;
        RECT 0.615000 2.730000 0.945000 3.245000 ;
        RECT 2.330000 2.730000 2.705000 3.245000 ;
        RECT 4.435000 2.650000 5.075000 3.245000 ;
        RECT 5.745000 1.950000 6.075000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
        RECT 6.395000 3.245000 6.565000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 6.720000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.115000 2.100000 0.715000 2.390000 ;
      RECT 0.115000 2.390000 2.695000 2.560000 ;
      RECT 0.115000 2.560000 0.445000 2.980000 ;
      RECT 0.220000 0.540000 0.715000 1.130000 ;
      RECT 0.545000 1.130000 0.715000 2.100000 ;
      RECT 1.150000 1.970000 1.625000 2.220000 ;
      RECT 1.235000 0.350000 1.625000 0.770000 ;
      RECT 1.235000 0.770000 3.020000 0.940000 ;
      RECT 1.235000 0.940000 1.625000 1.130000 ;
      RECT 1.455000 1.130000 1.625000 1.450000 ;
      RECT 1.455000 1.450000 1.830000 1.780000 ;
      RECT 1.455000 1.780000 1.625000 1.970000 ;
      RECT 1.795000 1.110000 3.325000 1.280000 ;
      RECT 1.795000 2.020000 2.170000 2.220000 ;
      RECT 2.000000 1.280000 2.170000 2.020000 ;
      RECT 2.525000 1.470000 2.855000 1.800000 ;
      RECT 2.525000 1.800000 2.695000 2.390000 ;
      RECT 2.850000 0.255000 4.005000 0.425000 ;
      RECT 2.850000 0.425000 3.020000 0.770000 ;
      RECT 2.905000 1.970000 3.195000 2.140000 ;
      RECT 2.905000 2.140000 3.075000 2.905000 ;
      RECT 2.905000 2.905000 4.045000 3.075000 ;
      RECT 3.025000 1.280000 3.325000 1.450000 ;
      RECT 3.025000 1.450000 3.195000 1.970000 ;
      RECT 3.190000 0.595000 3.665000 0.925000 ;
      RECT 3.245000 2.405000 3.535000 2.735000 ;
      RECT 3.365000 1.725000 4.925000 1.895000 ;
      RECT 3.365000 1.895000 3.535000 2.405000 ;
      RECT 3.495000 0.925000 3.665000 1.725000 ;
      RECT 3.715000 2.065000 4.045000 2.905000 ;
      RECT 3.835000 0.425000 4.005000 1.225000 ;
      RECT 3.835000 1.225000 4.095000 1.555000 ;
      RECT 4.305000 2.065000 5.575000 2.380000 ;
      RECT 4.665000 1.470000 4.925000 1.725000 ;
      RECT 4.770000 0.350000 5.100000 1.010000 ;
      RECT 4.770000 1.010000 6.295000 1.180000 ;
      RECT 5.095000 1.180000 5.265000 1.950000 ;
      RECT 5.095000 1.950000 5.575000 2.065000 ;
      RECT 5.245000 2.380000 5.575000 2.980000 ;
      RECT 5.975000 1.180000 6.295000 1.550000 ;
  END
END sky130_fd_sc_ls__dlrtp_1
