* File: sky130_fd_sc_ls__a221o_1.pxi.spice
* Created: Fri Aug 28 12:52:39 2020
* 
x_PM_SKY130_FD_SC_LS__A221O_1%A_148_260# N_A_148_260#_M1003_d
+ N_A_148_260#_M1001_d N_A_148_260#_M1009_d N_A_148_260#_c_69_n
+ N_A_148_260#_M1007_g N_A_148_260#_M1004_g N_A_148_260#_c_71_n
+ N_A_148_260#_c_72_n N_A_148_260#_c_73_n N_A_148_260#_c_74_n
+ N_A_148_260#_c_75_n N_A_148_260#_c_76_n N_A_148_260#_c_77_n
+ PM_SKY130_FD_SC_LS__A221O_1%A_148_260#
x_PM_SKY130_FD_SC_LS__A221O_1%A2 N_A2_c_151_n N_A2_M1008_g N_A2_c_152_n
+ N_A2_c_153_n N_A2_M1002_g A2 PM_SKY130_FD_SC_LS__A221O_1%A2
x_PM_SKY130_FD_SC_LS__A221O_1%A1 N_A1_c_193_n N_A1_M1010_g N_A1_M1003_g A1
+ N_A1_c_192_n PM_SKY130_FD_SC_LS__A221O_1%A1
x_PM_SKY130_FD_SC_LS__A221O_1%B1 N_B1_c_229_n N_B1_M1011_g N_B1_M1005_g B1
+ N_B1_c_231_n PM_SKY130_FD_SC_LS__A221O_1%B1
x_PM_SKY130_FD_SC_LS__A221O_1%B2 N_B2_M1006_g N_B2_c_263_n N_B2_M1000_g B2
+ PM_SKY130_FD_SC_LS__A221O_1%B2
x_PM_SKY130_FD_SC_LS__A221O_1%C1 N_C1_M1001_g N_C1_c_296_n N_C1_c_297_n
+ N_C1_c_301_n N_C1_M1009_g C1 N_C1_c_298_n N_C1_c_299_n
+ PM_SKY130_FD_SC_LS__A221O_1%C1
x_PM_SKY130_FD_SC_LS__A221O_1%X N_X_M1004_s N_X_M1007_s N_X_c_325_n X X X
+ N_X_c_327_n N_X_c_326_n PM_SKY130_FD_SC_LS__A221O_1%X
x_PM_SKY130_FD_SC_LS__A221O_1%VPWR N_VPWR_M1007_d N_VPWR_M1010_d N_VPWR_c_345_n
+ N_VPWR_c_346_n VPWR N_VPWR_c_347_n N_VPWR_c_348_n N_VPWR_c_349_n
+ N_VPWR_c_344_n N_VPWR_c_351_n N_VPWR_c_352_n PM_SKY130_FD_SC_LS__A221O_1%VPWR
x_PM_SKY130_FD_SC_LS__A221O_1%A_310_392# N_A_310_392#_M1008_d
+ N_A_310_392#_M1011_d N_A_310_392#_c_389_n N_A_310_392#_c_390_n
+ N_A_310_392#_c_391_n N_A_310_392#_c_392_n
+ PM_SKY130_FD_SC_LS__A221O_1%A_310_392#
x_PM_SKY130_FD_SC_LS__A221O_1%A_509_392# N_A_509_392#_M1011_s
+ N_A_509_392#_M1000_d N_A_509_392#_c_421_n N_A_509_392#_c_422_n
+ N_A_509_392#_c_423_n N_A_509_392#_c_424_n
+ PM_SKY130_FD_SC_LS__A221O_1%A_509_392#
x_PM_SKY130_FD_SC_LS__A221O_1%VGND N_VGND_M1004_d N_VGND_M1006_d N_VGND_c_445_n
+ VGND N_VGND_c_446_n N_VGND_c_447_n N_VGND_c_448_n N_VGND_c_449_n
+ N_VGND_c_450_n N_VGND_c_451_n PM_SKY130_FD_SC_LS__A221O_1%VGND
cc_1 VNB N_A_148_260#_c_69_n 0.0359115f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=1.765
cc_2 VNB N_A_148_260#_M1004_g 0.0272723f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_3 VNB N_A_148_260#_c_71_n 0.00606973f $X=-0.19 $Y=-0.245 $X2=2.42 $Y2=1.095
cc_4 VNB N_A_148_260#_c_72_n 0.0146376f $X=-0.19 $Y=-0.245 $X2=1.205 $Y2=1.095
cc_5 VNB N_A_148_260#_c_73_n 0.00351237f $X=-0.19 $Y=-0.245 $X2=2.64 $Y2=0.52
cc_6 VNB N_A_148_260#_c_74_n 0.0155437f $X=-0.19 $Y=-0.245 $X2=3.86 $Y2=1.2
cc_7 VNB N_A_148_260#_c_75_n 0.016015f $X=-0.19 $Y=-0.245 $X2=4.05 $Y2=2.105
cc_8 VNB N_A_148_260#_c_76_n 0.00697255f $X=-0.19 $Y=-0.245 $X2=2.42 $Y2=1.01
cc_9 VNB N_A_148_260#_c_77_n 0.018536f $X=-0.19 $Y=-0.245 $X2=4.025 $Y2=1.005
cc_10 VNB N_A2_c_151_n 0.0427115f $X=-0.19 $Y=-0.245 $X2=2.445 $Y2=0.395
cc_11 VNB N_A2_c_152_n 0.0278546f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A2_c_153_n 0.0158993f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB A2 0.00382554f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A1_M1003_g 0.0360321f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB A1 0.00325885f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A1_c_192_n 0.0280825f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=2.4
cc_17 VNB N_B1_c_229_n 0.0160825f $X=-0.19 $Y=-0.245 $X2=2.445 $Y2=0.395
cc_18 VNB N_B1_M1005_g 0.0314209f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_B1_c_231_n 0.00393964f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=2.4
cc_20 VNB N_B2_M1006_g 0.0312467f $X=-0.19 $Y=-0.245 $X2=3.9 $Y2=1.96
cc_21 VNB N_B2_c_263_n 0.0162046f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB B2 0.00431791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_C1_M1001_g 0.0117153f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_C1_c_296_n 0.00721292f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_C1_c_297_n 0.015492f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_C1_c_298_n 0.0650756f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_C1_c_299_n 0.00655821f $X=-0.19 $Y=-0.245 $X2=2.42 $Y2=1.095
cc_28 VNB N_X_c_325_n 0.0653482f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=2.4
cc_29 VNB N_X_c_326_n 0.0329591f $X=-0.19 $Y=-0.245 $X2=4.05 $Y2=2.815
cc_30 VNB N_VPWR_c_344_n 0.183584f $X=-0.19 $Y=-0.245 $X2=2.42 $Y2=1.01
cc_31 VNB N_VGND_c_445_n 0.00920632f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_446_n 0.0397973f $X=-0.19 $Y=-0.245 $X2=1.205 $Y2=1.095
cc_33 VNB N_VGND_c_447_n 0.0188832f $X=-0.19 $Y=-0.245 $X2=4.05 $Y2=2.815
cc_34 VNB N_VGND_c_448_n 0.269269f $X=-0.19 $Y=-0.245 $X2=4.05 $Y2=2.815
cc_35 VNB N_VGND_c_449_n 0.0294689f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.465
cc_36 VNB N_VGND_c_450_n 0.0280769f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_451_n 0.00711538f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VPB N_A_148_260#_c_69_n 0.0284372f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=1.765
cc_39 VPB N_A_148_260#_c_75_n 0.0547501f $X=-0.19 $Y=1.66 $X2=4.05 $Y2=2.105
cc_40 VPB N_A2_c_151_n 0.034894f $X=-0.19 $Y=1.66 $X2=2.445 $Y2=0.395
cc_41 VPB A2 0.00443709f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_42 VPB N_A1_c_193_n 0.0194376f $X=-0.19 $Y=1.66 $X2=2.445 $Y2=0.395
cc_43 VPB A1 0.00258775f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_44 VPB N_A1_c_192_n 0.0340961f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=2.4
cc_45 VPB N_B1_c_229_n 0.0383639f $X=-0.19 $Y=1.66 $X2=2.445 $Y2=0.395
cc_46 VPB N_B1_c_231_n 0.00281847f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=2.4
cc_47 VPB N_B2_c_263_n 0.0341959f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 VPB B2 0.00411652f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 VPB N_C1_c_297_n 0.00860859f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_C1_c_301_n 0.0276533f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_51 VPB N_X_c_327_n 0.0853596f $X=-0.19 $Y=1.66 $X2=4.05 $Y2=2.105
cc_52 VPB N_X_c_326_n 0.0102153f $X=-0.19 $Y=1.66 $X2=4.05 $Y2=2.815
cc_53 VPB N_VPWR_c_345_n 0.00873403f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_346_n 0.0119493f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=0.74
cc_55 VPB N_VPWR_c_347_n 0.0311089f $X=-0.19 $Y=1.66 $X2=2.64 $Y2=1.01
cc_56 VPB N_VPWR_c_348_n 0.018048f $X=-0.19 $Y=1.66 $X2=2.86 $Y2=1.2
cc_57 VPB N_VPWR_c_349_n 0.0520118f $X=-0.19 $Y=1.66 $X2=0.905 $Y2=1.465
cc_58 VPB N_VPWR_c_344_n 0.0803342f $X=-0.19 $Y=1.66 $X2=2.42 $Y2=1.01
cc_59 VPB N_VPWR_c_351_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_352_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0.905 $Y2=1.465
cc_61 VPB N_A_310_392#_c_389_n 0.00184202f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_A_310_392#_c_390_n 0.00216998f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_A_310_392#_c_391_n 0.0134249f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=2.4
cc_64 VPB N_A_310_392#_c_392_n 0.00417513f $X=-0.19 $Y=1.66 $X2=1.205 $Y2=1.095
cc_65 VPB N_A_509_392#_c_421_n 0.00568f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_A_509_392#_c_422_n 0.00580134f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=2.4
cc_67 VPB N_A_509_392#_c_423_n 0.00398658f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=2.4
cc_68 VPB N_A_509_392#_c_424_n 0.00185469f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=0.74
cc_69 N_A_148_260#_c_69_n N_A2_c_151_n 0.0268948f $X=0.96 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_70 N_A_148_260#_M1004_g N_A2_c_151_n 0.0250238f $X=0.995 $Y=0.74 $X2=-0.19
+ $Y2=-0.245
cc_71 N_A_148_260#_c_71_n N_A2_c_151_n 0.0128506f $X=2.42 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_72 N_A_148_260#_c_72_n N_A2_c_151_n 0.00598031f $X=1.205 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_73 N_A_148_260#_c_71_n N_A2_c_152_n 0.0141544f $X=2.42 $Y=1.095 $X2=0 $Y2=0
cc_74 N_A_148_260#_c_71_n N_A2_c_153_n 0.0103411f $X=2.42 $Y=1.095 $X2=0 $Y2=0
cc_75 N_A_148_260#_c_73_n N_A2_c_153_n 0.00210649f $X=2.64 $Y=0.52 $X2=0 $Y2=0
cc_76 N_A_148_260#_c_69_n A2 0.00260476f $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_77 N_A_148_260#_c_71_n A2 0.031704f $X=2.42 $Y=1.095 $X2=0 $Y2=0
cc_78 N_A_148_260#_c_72_n A2 0.0233111f $X=1.205 $Y=1.095 $X2=0 $Y2=0
cc_79 N_A_148_260#_c_71_n N_A1_M1003_g 0.0142322f $X=2.42 $Y=1.095 $X2=0 $Y2=0
cc_80 N_A_148_260#_c_73_n N_A1_M1003_g 0.0109036f $X=2.64 $Y=0.52 $X2=0 $Y2=0
cc_81 N_A_148_260#_c_76_n N_A1_M1003_g 0.00743095f $X=2.42 $Y=1.01 $X2=0 $Y2=0
cc_82 N_A_148_260#_c_71_n A1 0.0161399f $X=2.42 $Y=1.095 $X2=0 $Y2=0
cc_83 N_A_148_260#_c_71_n N_A1_c_192_n 0.00228749f $X=2.42 $Y=1.095 $X2=0 $Y2=0
cc_84 N_A_148_260#_c_76_n N_B1_c_229_n 0.00429782f $X=2.42 $Y=1.01 $X2=-0.19
+ $Y2=-0.245
cc_85 N_A_148_260#_c_73_n N_B1_M1005_g 0.0107522f $X=2.64 $Y=0.52 $X2=0 $Y2=0
cc_86 N_A_148_260#_c_74_n N_B1_M1005_g 0.0106483f $X=3.86 $Y=1.2 $X2=0 $Y2=0
cc_87 N_A_148_260#_c_76_n N_B1_M1005_g 0.00634212f $X=2.42 $Y=1.01 $X2=0 $Y2=0
cc_88 N_A_148_260#_c_74_n N_B1_c_231_n 0.00888173f $X=3.86 $Y=1.2 $X2=0 $Y2=0
cc_89 N_A_148_260#_c_76_n N_B1_c_231_n 0.0286449f $X=2.42 $Y=1.01 $X2=0 $Y2=0
cc_90 N_A_148_260#_c_73_n N_B2_M1006_g 0.00186941f $X=2.64 $Y=0.52 $X2=0 $Y2=0
cc_91 N_A_148_260#_c_74_n N_B2_M1006_g 0.0143581f $X=3.86 $Y=1.2 $X2=0 $Y2=0
cc_92 N_A_148_260#_c_75_n N_B2_M1006_g 5.28813e-19 $X=4.05 $Y=2.105 $X2=0 $Y2=0
cc_93 N_A_148_260#_c_76_n N_B2_M1006_g 5.21288e-19 $X=2.42 $Y=1.01 $X2=0 $Y2=0
cc_94 N_A_148_260#_c_77_n N_B2_M1006_g 6.52731e-19 $X=4.025 $Y=1.005 $X2=0 $Y2=0
cc_95 N_A_148_260#_c_74_n N_B2_c_263_n 0.00437633f $X=3.86 $Y=1.2 $X2=0 $Y2=0
cc_96 N_A_148_260#_c_75_n N_B2_c_263_n 0.00134953f $X=4.05 $Y=2.105 $X2=0 $Y2=0
cc_97 N_A_148_260#_c_74_n B2 0.0392571f $X=3.86 $Y=1.2 $X2=0 $Y2=0
cc_98 N_A_148_260#_c_75_n B2 0.0266398f $X=4.05 $Y=2.105 $X2=0 $Y2=0
cc_99 N_A_148_260#_c_74_n N_C1_M1001_g 0.0160646f $X=3.86 $Y=1.2 $X2=0 $Y2=0
cc_100 N_A_148_260#_c_75_n N_C1_M1001_g 0.00196628f $X=4.05 $Y=2.105 $X2=0 $Y2=0
cc_101 N_A_148_260#_c_77_n N_C1_M1001_g 0.00871597f $X=4.025 $Y=1.005 $X2=0
+ $Y2=0
cc_102 N_A_148_260#_c_75_n N_C1_c_296_n 0.00434931f $X=4.05 $Y=2.105 $X2=0 $Y2=0
cc_103 N_A_148_260#_c_75_n N_C1_c_297_n 0.0120954f $X=4.05 $Y=2.105 $X2=0 $Y2=0
cc_104 N_A_148_260#_c_75_n N_C1_c_301_n 0.0176364f $X=4.05 $Y=2.105 $X2=0 $Y2=0
cc_105 N_A_148_260#_c_77_n N_C1_c_298_n 0.00152775f $X=4.025 $Y=1.005 $X2=0
+ $Y2=0
cc_106 N_A_148_260#_M1001_d N_C1_c_299_n 0.00226737f $X=3.885 $Y=0.615 $X2=0
+ $Y2=0
cc_107 N_A_148_260#_c_77_n N_C1_c_299_n 0.0229409f $X=4.025 $Y=1.005 $X2=0 $Y2=0
cc_108 N_A_148_260#_c_69_n N_X_c_325_n 9.8857e-19 $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_109 N_A_148_260#_M1004_g N_X_c_325_n 0.00202121f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_110 N_A_148_260#_c_72_n N_X_c_325_n 0.0164255f $X=1.205 $Y=1.095 $X2=0 $Y2=0
cc_111 N_A_148_260#_c_69_n N_X_c_327_n 0.0171322f $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_112 N_A_148_260#_c_72_n N_X_c_327_n 0.0123231f $X=1.205 $Y=1.095 $X2=0 $Y2=0
cc_113 N_A_148_260#_c_69_n N_X_c_326_n 0.00815006f $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_114 N_A_148_260#_M1004_g N_X_c_326_n 0.00297287f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_115 N_A_148_260#_c_72_n N_X_c_326_n 0.0266447f $X=1.205 $Y=1.095 $X2=0 $Y2=0
cc_116 N_A_148_260#_c_69_n N_VPWR_c_345_n 0.00653855f $X=0.96 $Y=1.765 $X2=0
+ $Y2=0
cc_117 N_A_148_260#_c_72_n N_VPWR_c_345_n 0.00602121f $X=1.205 $Y=1.095 $X2=0
+ $Y2=0
cc_118 N_A_148_260#_c_69_n N_VPWR_c_347_n 0.00445602f $X=0.96 $Y=1.765 $X2=0
+ $Y2=0
cc_119 N_A_148_260#_c_75_n N_VPWR_c_349_n 0.0145938f $X=4.05 $Y=2.105 $X2=0
+ $Y2=0
cc_120 N_A_148_260#_c_69_n N_VPWR_c_344_n 0.00863027f $X=0.96 $Y=1.765 $X2=0
+ $Y2=0
cc_121 N_A_148_260#_c_75_n N_VPWR_c_344_n 0.0120466f $X=4.05 $Y=2.105 $X2=0
+ $Y2=0
cc_122 N_A_148_260#_c_74_n N_A_310_392#_c_392_n 0.00682195f $X=3.86 $Y=1.2 $X2=0
+ $Y2=0
cc_123 N_A_148_260#_c_75_n N_A_509_392#_c_422_n 0.00549849f $X=4.05 $Y=2.105
+ $X2=0 $Y2=0
cc_124 N_A_148_260#_c_75_n N_A_509_392#_c_424_n 0.0629452f $X=4.05 $Y=2.105
+ $X2=0 $Y2=0
cc_125 N_A_148_260#_c_71_n N_VGND_M1004_d 0.00740749f $X=2.42 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_126 N_A_148_260#_c_72_n N_VGND_M1004_d 8.62855e-19 $X=1.205 $Y=1.095
+ $X2=-0.19 $Y2=-0.245
cc_127 N_A_148_260#_c_74_n N_VGND_M1006_d 0.00228244f $X=3.86 $Y=1.2 $X2=0 $Y2=0
cc_128 N_A_148_260#_c_73_n N_VGND_c_445_n 0.0196681f $X=2.64 $Y=0.52 $X2=0 $Y2=0
cc_129 N_A_148_260#_c_74_n N_VGND_c_445_n 0.0265066f $X=3.86 $Y=1.2 $X2=0 $Y2=0
cc_130 N_A_148_260#_c_73_n N_VGND_c_446_n 0.0176208f $X=2.64 $Y=0.52 $X2=0 $Y2=0
cc_131 N_A_148_260#_M1004_g N_VGND_c_448_n 0.00757924f $X=0.995 $Y=0.74 $X2=0
+ $Y2=0
cc_132 N_A_148_260#_c_73_n N_VGND_c_448_n 0.0158894f $X=2.64 $Y=0.52 $X2=0 $Y2=0
cc_133 N_A_148_260#_c_77_n N_VGND_c_448_n 0.0015257f $X=4.025 $Y=1.005 $X2=0
+ $Y2=0
cc_134 N_A_148_260#_M1004_g N_VGND_c_449_n 0.00383152f $X=0.995 $Y=0.74 $X2=0
+ $Y2=0
cc_135 N_A_148_260#_M1004_g N_VGND_c_450_n 0.0170948f $X=0.995 $Y=0.74 $X2=0
+ $Y2=0
cc_136 N_A_148_260#_c_71_n N_VGND_c_450_n 0.0567101f $X=2.42 $Y=1.095 $X2=0
+ $Y2=0
cc_137 N_A_148_260#_c_72_n N_VGND_c_450_n 0.00900333f $X=1.205 $Y=1.095 $X2=0
+ $Y2=0
cc_138 N_A_148_260#_c_73_n N_VGND_c_450_n 0.0169741f $X=2.64 $Y=0.52 $X2=0 $Y2=0
cc_139 N_A_148_260#_c_71_n A_417_79# 0.00366293f $X=2.42 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_140 N_A2_c_151_n N_A1_c_193_n 0.00837512f $X=1.475 $Y=1.885 $X2=-0.19
+ $Y2=-0.245
cc_141 N_A2_c_151_n N_A1_M1003_g 0.00353069f $X=1.475 $Y=1.885 $X2=0 $Y2=0
cc_142 N_A2_c_153_n N_A1_M1003_g 0.0598892f $X=2.01 $Y=1.11 $X2=0 $Y2=0
cc_143 A2 N_A1_M1003_g 0.00226541f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_144 N_A2_c_151_n A1 3.32859e-19 $X=1.475 $Y=1.885 $X2=0 $Y2=0
cc_145 N_A2_c_152_n A1 5.06846e-19 $X=1.935 $Y=1.185 $X2=0 $Y2=0
cc_146 A2 A1 0.0250482f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_147 N_A2_c_151_n N_A1_c_192_n 0.0238621f $X=1.475 $Y=1.885 $X2=0 $Y2=0
cc_148 N_A2_c_152_n N_A1_c_192_n 0.0170914f $X=1.935 $Y=1.185 $X2=0 $Y2=0
cc_149 A2 N_A1_c_192_n 0.00263634f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_150 N_A2_c_151_n N_X_c_327_n 8.60374e-19 $X=1.475 $Y=1.885 $X2=0 $Y2=0
cc_151 N_A2_c_151_n N_VPWR_c_345_n 0.00941688f $X=1.475 $Y=1.885 $X2=0 $Y2=0
cc_152 N_A2_c_151_n N_VPWR_c_346_n 5.47162e-19 $X=1.475 $Y=1.885 $X2=0 $Y2=0
cc_153 N_A2_c_151_n N_VPWR_c_348_n 0.00445602f $X=1.475 $Y=1.885 $X2=0 $Y2=0
cc_154 N_A2_c_151_n N_VPWR_c_344_n 0.00857973f $X=1.475 $Y=1.885 $X2=0 $Y2=0
cc_155 N_A2_c_151_n N_A_310_392#_c_389_n 0.00302753f $X=1.475 $Y=1.885 $X2=0
+ $Y2=0
cc_156 A2 N_A_310_392#_c_389_n 0.0223454f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_157 N_A2_c_151_n N_A_310_392#_c_390_n 0.00863729f $X=1.475 $Y=1.885 $X2=0
+ $Y2=0
cc_158 A2 N_A_310_392#_c_391_n 6.34813e-19 $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_159 N_A2_c_153_n N_VGND_c_446_n 0.00446421f $X=2.01 $Y=1.11 $X2=0 $Y2=0
cc_160 N_A2_c_153_n N_VGND_c_448_n 0.00430282f $X=2.01 $Y=1.11 $X2=0 $Y2=0
cc_161 N_A2_c_151_n N_VGND_c_450_n 0.00269777f $X=1.475 $Y=1.885 $X2=0 $Y2=0
cc_162 N_A2_c_153_n N_VGND_c_450_n 0.0158598f $X=2.01 $Y=1.11 $X2=0 $Y2=0
cc_163 N_A1_M1003_g N_B1_c_229_n 0.0212847f $X=2.37 $Y=0.715 $X2=-0.19
+ $Y2=-0.245
cc_164 A1 N_B1_c_229_n 3.42046e-19 $X=2.075 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_165 N_A1_c_192_n N_B1_c_229_n 8.1341e-19 $X=2.13 $Y=1.635 $X2=-0.19
+ $Y2=-0.245
cc_166 N_A1_M1003_g N_B1_M1005_g 0.0176935f $X=2.37 $Y=0.715 $X2=0 $Y2=0
cc_167 N_A1_M1003_g N_B1_c_231_n 0.00303956f $X=2.37 $Y=0.715 $X2=0 $Y2=0
cc_168 A1 N_B1_c_231_n 0.0201161f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_169 N_A1_c_193_n N_VPWR_c_346_n 0.0119223f $X=1.925 $Y=1.885 $X2=0 $Y2=0
cc_170 N_A1_c_193_n N_VPWR_c_348_n 0.00413917f $X=1.925 $Y=1.885 $X2=0 $Y2=0
cc_171 N_A1_c_193_n N_VPWR_c_344_n 0.0081781f $X=1.925 $Y=1.885 $X2=0 $Y2=0
cc_172 N_A1_c_193_n N_A_310_392#_c_389_n 4.701e-19 $X=1.925 $Y=1.885 $X2=0 $Y2=0
cc_173 N_A1_c_193_n N_A_310_392#_c_390_n 0.00598833f $X=1.925 $Y=1.885 $X2=0
+ $Y2=0
cc_174 N_A1_c_193_n N_A_310_392#_c_391_n 0.0178341f $X=1.925 $Y=1.885 $X2=0
+ $Y2=0
cc_175 A1 N_A_310_392#_c_391_n 0.0222046f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_176 N_A1_c_192_n N_A_310_392#_c_391_n 0.00813866f $X=2.13 $Y=1.635 $X2=0
+ $Y2=0
cc_177 N_A1_c_193_n N_A_509_392#_c_423_n 5.75404e-19 $X=1.925 $Y=1.885 $X2=0
+ $Y2=0
cc_178 N_A1_M1003_g N_VGND_c_446_n 0.00534051f $X=2.37 $Y=0.715 $X2=0 $Y2=0
cc_179 N_A1_M1003_g N_VGND_c_448_n 0.00537853f $X=2.37 $Y=0.715 $X2=0 $Y2=0
cc_180 N_A1_M1003_g N_VGND_c_450_n 0.00181914f $X=2.37 $Y=0.715 $X2=0 $Y2=0
cc_181 N_B1_M1005_g N_B2_M1006_g 0.0463342f $X=2.91 $Y=0.715 $X2=0 $Y2=0
cc_182 N_B1_c_229_n N_B2_c_263_n 0.0714128f $X=2.895 $Y=1.885 $X2=0 $Y2=0
cc_183 N_B1_c_231_n N_B2_c_263_n 4.06919e-19 $X=2.82 $Y=1.615 $X2=0 $Y2=0
cc_184 N_B1_c_229_n B2 4.06298e-19 $X=2.895 $Y=1.885 $X2=0 $Y2=0
cc_185 N_B1_c_231_n B2 0.0219204f $X=2.82 $Y=1.615 $X2=0 $Y2=0
cc_186 N_B1_c_229_n N_VPWR_c_346_n 8.71134e-19 $X=2.895 $Y=1.885 $X2=0 $Y2=0
cc_187 N_B1_c_229_n N_VPWR_c_349_n 0.00278271f $X=2.895 $Y=1.885 $X2=0 $Y2=0
cc_188 N_B1_c_229_n N_VPWR_c_344_n 0.00358708f $X=2.895 $Y=1.885 $X2=0 $Y2=0
cc_189 N_B1_c_229_n N_A_310_392#_c_391_n 0.0172584f $X=2.895 $Y=1.885 $X2=0
+ $Y2=0
cc_190 N_B1_c_231_n N_A_310_392#_c_391_n 0.0274068f $X=2.82 $Y=1.615 $X2=0 $Y2=0
cc_191 N_B1_c_229_n N_A_310_392#_c_392_n 0.0149088f $X=2.895 $Y=1.885 $X2=0
+ $Y2=0
cc_192 N_B1_c_231_n N_A_310_392#_c_392_n 0.00245955f $X=2.82 $Y=1.615 $X2=0
+ $Y2=0
cc_193 N_B1_c_229_n N_A_509_392#_c_422_n 0.0136535f $X=2.895 $Y=1.885 $X2=0
+ $Y2=0
cc_194 N_B1_M1005_g N_VGND_c_445_n 0.00210079f $X=2.91 $Y=0.715 $X2=0 $Y2=0
cc_195 N_B1_M1005_g N_VGND_c_446_n 0.00534051f $X=2.91 $Y=0.715 $X2=0 $Y2=0
cc_196 N_B1_M1005_g N_VGND_c_448_n 0.00537853f $X=2.91 $Y=0.715 $X2=0 $Y2=0
cc_197 N_B2_c_263_n N_C1_c_297_n 0.0241402f $X=3.345 $Y=1.885 $X2=0 $Y2=0
cc_198 B2 N_C1_c_297_n 0.0024298f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_199 N_B2_c_263_n N_C1_c_301_n 0.0070726f $X=3.345 $Y=1.885 $X2=0 $Y2=0
cc_200 N_B2_M1006_g N_C1_c_298_n 0.0241579f $X=3.27 $Y=0.715 $X2=0 $Y2=0
cc_201 N_B2_c_263_n N_VPWR_c_349_n 0.00278271f $X=3.345 $Y=1.885 $X2=0 $Y2=0
cc_202 N_B2_c_263_n N_VPWR_c_344_n 0.00354253f $X=3.345 $Y=1.885 $X2=0 $Y2=0
cc_203 N_B2_c_263_n N_A_310_392#_c_392_n 0.0120529f $X=3.345 $Y=1.885 $X2=0
+ $Y2=0
cc_204 B2 N_A_310_392#_c_392_n 0.00751427f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_205 N_B2_c_263_n N_A_509_392#_c_422_n 0.0125894f $X=3.345 $Y=1.885 $X2=0
+ $Y2=0
cc_206 N_B2_c_263_n N_A_509_392#_c_424_n 0.0069352f $X=3.345 $Y=1.885 $X2=0
+ $Y2=0
cc_207 B2 N_A_509_392#_c_424_n 0.0173356f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_208 N_B2_M1006_g N_VGND_c_445_n 0.0135704f $X=3.27 $Y=0.715 $X2=0 $Y2=0
cc_209 N_B2_M1006_g N_VGND_c_446_n 0.00465077f $X=3.27 $Y=0.715 $X2=0 $Y2=0
cc_210 N_B2_M1006_g N_VGND_c_448_n 0.00451796f $X=3.27 $Y=0.715 $X2=0 $Y2=0
cc_211 N_C1_c_301_n N_VPWR_c_349_n 0.00445602f $X=3.825 $Y=1.885 $X2=0 $Y2=0
cc_212 N_C1_c_301_n N_VPWR_c_344_n 0.00862158f $X=3.825 $Y=1.885 $X2=0 $Y2=0
cc_213 N_C1_c_301_n N_A_509_392#_c_422_n 0.00345421f $X=3.825 $Y=1.885 $X2=0
+ $Y2=0
cc_214 N_C1_c_301_n N_A_509_392#_c_424_n 0.0031718f $X=3.825 $Y=1.885 $X2=0
+ $Y2=0
cc_215 N_C1_c_298_n N_VGND_c_445_n 0.0089245f $X=4.03 $Y=0.34 $X2=0 $Y2=0
cc_216 N_C1_c_299_n N_VGND_c_445_n 0.0300657f $X=4.03 $Y=0.34 $X2=0 $Y2=0
cc_217 N_C1_c_298_n N_VGND_c_447_n 0.0108828f $X=4.03 $Y=0.34 $X2=0 $Y2=0
cc_218 N_C1_c_299_n N_VGND_c_447_n 0.0215843f $X=4.03 $Y=0.34 $X2=0 $Y2=0
cc_219 N_C1_c_298_n N_VGND_c_448_n 0.0176737f $X=4.03 $Y=0.34 $X2=0 $Y2=0
cc_220 N_C1_c_299_n N_VGND_c_448_n 0.0110944f $X=4.03 $Y=0.34 $X2=0 $Y2=0
cc_221 N_X_c_327_n N_VPWR_c_345_n 0.0730738f $X=0.735 $Y=1.985 $X2=0 $Y2=0
cc_222 N_X_c_327_n N_VPWR_c_347_n 0.0344501f $X=0.735 $Y=1.985 $X2=0 $Y2=0
cc_223 N_X_c_327_n N_VPWR_c_344_n 0.0284819f $X=0.735 $Y=1.985 $X2=0 $Y2=0
cc_224 N_X_c_325_n N_VGND_c_448_n 0.0273142f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_225 N_X_c_325_n N_VGND_c_449_n 0.0328875f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_226 N_X_c_325_n N_VGND_c_450_n 0.0205275f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_227 N_VPWR_c_345_n N_A_310_392#_c_389_n 0.00770453f $X=1.185 $Y=2.115 $X2=0
+ $Y2=0
cc_228 N_VPWR_c_345_n N_A_310_392#_c_390_n 0.0289071f $X=1.185 $Y=2.115 $X2=0
+ $Y2=0
cc_229 N_VPWR_c_346_n N_A_310_392#_c_390_n 0.0449538f $X=2.15 $Y=2.475 $X2=0
+ $Y2=0
cc_230 N_VPWR_c_348_n N_A_310_392#_c_390_n 0.0110241f $X=1.985 $Y=3.33 $X2=0
+ $Y2=0
cc_231 N_VPWR_c_344_n N_A_310_392#_c_390_n 0.00909194f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_232 N_VPWR_M1010_d N_A_310_392#_c_391_n 0.00497391f $X=2 $Y=1.96 $X2=0 $Y2=0
cc_233 N_VPWR_c_346_n N_A_310_392#_c_391_n 0.0220544f $X=2.15 $Y=2.475 $X2=0
+ $Y2=0
cc_234 N_VPWR_c_346_n N_A_509_392#_c_421_n 0.0452163f $X=2.15 $Y=2.475 $X2=0
+ $Y2=0
cc_235 N_VPWR_c_349_n N_A_509_392#_c_422_n 0.0584986f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_236 N_VPWR_c_344_n N_A_509_392#_c_422_n 0.0327208f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_237 N_VPWR_c_346_n N_A_509_392#_c_423_n 0.0139f $X=2.15 $Y=2.475 $X2=0 $Y2=0
cc_238 N_VPWR_c_349_n N_A_509_392#_c_423_n 0.0200723f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_239 N_VPWR_c_344_n N_A_509_392#_c_423_n 0.0108858f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_240 N_A_310_392#_c_391_n N_A_509_392#_M1011_s 0.00537906f $X=2.955 $Y=2.055
+ $X2=-0.19 $Y2=1.66
cc_241 N_A_310_392#_c_391_n N_A_509_392#_c_421_n 0.0210301f $X=2.955 $Y=2.055
+ $X2=0 $Y2=0
cc_242 N_A_310_392#_M1011_d N_A_509_392#_c_422_n 0.00197722f $X=2.97 $Y=1.96
+ $X2=0 $Y2=0
cc_243 N_A_310_392#_c_392_n N_A_509_392#_c_422_n 0.0160777f $X=3.12 $Y=2.115
+ $X2=0 $Y2=0
cc_244 N_A_310_392#_c_392_n N_A_509_392#_c_424_n 0.0524457f $X=3.12 $Y=2.115
+ $X2=0 $Y2=0
