* File: sky130_fd_sc_ls__dlrtp_2.pex.spice
* Created: Fri Aug 28 13:19:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__DLRTP_2%D 1 3 6 8 12
c28 6 0 1.60049e-19 $X=0.52 $Y=0.835
r29 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.615 $X2=0.385 $Y2=1.615
r30 8 12 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=0.24 $Y=1.615
+ $X2=0.385 $Y2=1.615
r31 4 11 38.5818 $w=3.27e-07 $l=2.14173e-07 $layer=POLY_cond $X=0.52 $Y=1.45
+ $X2=0.407 $Y2=1.615
r32 4 6 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=0.52 $Y=1.45 $X2=0.52
+ $Y2=0.835
r33 1 11 54.0589 $w=3.27e-07 $l=3.15214e-07 $layer=POLY_cond $X=0.505 $Y=1.885
+ $X2=0.407 $Y2=1.615
r34 1 3 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.505 $Y=1.885
+ $X2=0.505 $Y2=2.38
.ends

.subckt PM_SKY130_FD_SC_LS__DLRTP_2%GATE 3 5 6 8 9 12 14
c43 9 0 2.85504e-19 $X=1.2 $Y=1.295
r44 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.155 $Y=1.385
+ $X2=1.155 $Y2=1.55
r45 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.155 $Y=1.385
+ $X2=1.155 $Y2=1.22
r46 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.155
+ $Y=1.385 $X2=1.155 $Y2=1.385
r47 9 13 3.98923 $w=2.58e-07 $l=9e-08 $layer=LI1_cond $X=1.155 $Y=1.295
+ $X2=1.155 $Y2=1.385
r48 6 8 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.125 $Y=1.885
+ $X2=1.125 $Y2=2.38
r49 5 6 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.125 $Y=1.795 $X2=1.125
+ $Y2=1.885
r50 5 15 95.2339 $w=1.8e-07 $l=2.45e-07 $layer=POLY_cond $X=1.125 $Y=1.795
+ $X2=1.125 $Y2=1.55
r51 3 14 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.1 $Y=0.74 $X2=1.1
+ $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_LS__DLRTP_2%A_235_74# 1 2 7 9 12 14 16 17 18 21 24 26 28
+ 29 32 33 34 38 45 50 54 55 56
c151 33 0 1.78997e-19 $X=3.92 $Y=0.34
c152 24 0 1.25456e-19 $X=2.045 $Y=1.585
c153 21 0 1.18818e-19 $X=3.845 $Y=0.615
c154 18 0 3.77203e-19 $X=3.26 $Y=1.735
c155 17 0 1.64562e-19 $X=3.76 $Y=1.735
c156 7 0 1.86781e-19 $X=2.135 $Y=1.885
r157 54 56 8.65224 $w=2.63e-07 $l=1.65e-07 $layer=LI1_cond $X=3.957 $Y=1.425
+ $X2=3.957 $Y2=1.26
r158 54 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.925
+ $Y=1.425 $X2=3.925 $Y2=1.425
r159 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.725
+ $Y=1.585 $X2=1.725 $Y2=1.585
r160 47 50 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=1.54 $Y=1.585
+ $X2=1.725 $Y2=1.585
r161 43 45 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=1.35 $Y=2.105
+ $X2=1.54 $Y2=2.105
r162 40 41 13.8993 $w=4.73e-07 $l=3.45e-07 $layer=LI1_cond $X=1.387 $Y=0.665
+ $X2=1.387 $Y2=1.01
r163 38 40 3.77709 $w=4.73e-07 $l=1.5e-07 $layer=LI1_cond $X=1.387 $Y=0.515
+ $X2=1.387 $Y2=0.665
r164 35 56 54.4759 $w=1.68e-07 $l=8.35e-07 $layer=LI1_cond $X=4.005 $Y=0.425
+ $X2=4.005 $Y2=1.26
r165 33 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.92 $Y=0.34
+ $X2=4.005 $Y2=0.425
r166 33 34 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=3.92 $Y=0.34
+ $X2=2.975 $Y2=0.34
r167 31 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.89 $Y=0.425
+ $X2=2.975 $Y2=0.34
r168 31 32 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=2.89 $Y=0.425
+ $X2=2.89 $Y2=0.58
r169 30 40 6.83586 $w=1.7e-07 $l=2.38e-07 $layer=LI1_cond $X=1.625 $Y=0.665
+ $X2=1.387 $Y2=0.665
r170 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.805 $Y=0.665
+ $X2=2.89 $Y2=0.58
r171 29 30 76.984 $w=1.68e-07 $l=1.18e-06 $layer=LI1_cond $X=2.805 $Y=0.665
+ $X2=1.625 $Y2=0.665
r172 28 45 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.54 $Y=1.94
+ $X2=1.54 $Y2=2.105
r173 27 47 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.54 $Y=1.75
+ $X2=1.54 $Y2=1.585
r174 27 28 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.54 $Y=1.75
+ $X2=1.54 $Y2=1.94
r175 26 47 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.54 $Y=1.42
+ $X2=1.54 $Y2=1.585
r176 26 41 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=1.54 $Y=1.42
+ $X2=1.54 $Y2=1.01
r177 24 51 55.9556 $w=3.3e-07 $l=3.2e-07 $layer=POLY_cond $X=2.045 $Y=1.585
+ $X2=1.725 $Y2=1.585
r178 19 55 39.2009 $w=2.58e-07 $l=2.0106e-07 $layer=POLY_cond $X=3.845 $Y=1.26
+ $X2=3.925 $Y2=1.425
r179 19 21 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=3.845 $Y=1.26
+ $X2=3.845 $Y2=0.615
r180 17 55 57.9147 $w=2.58e-07 $l=3.83732e-07 $layer=POLY_cond $X=3.76 $Y=1.735
+ $X2=3.925 $Y2=1.425
r181 17 18 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=3.76 $Y=1.735
+ $X2=3.26 $Y2=1.735
r182 14 18 26.9307 $w=1.5e-07 $l=1.89737e-07 $layer=POLY_cond $X=3.17 $Y=1.885
+ $X2=3.26 $Y2=1.735
r183 14 16 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.17 $Y=1.885
+ $X2=3.17 $Y2=2.46
r184 10 24 44.4105 $w=1.88e-07 $l=1.78452e-07 $layer=POLY_cond $X=2.175 $Y=1.42
+ $X2=2.147 $Y2=1.585
r185 10 12 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.175 $Y=1.42
+ $X2=2.175 $Y2=0.86
r186 7 24 79.0222 $w=1.88e-07 $l=3.05941e-07 $layer=POLY_cond $X=2.135 $Y=1.885
+ $X2=2.147 $Y2=1.585
r187 7 9 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.135 $Y=1.885
+ $X2=2.135 $Y2=2.38
r188 2 43 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.2
+ $Y=1.96 $X2=1.35 $Y2=2.105
r189 1 38 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.175
+ $Y=0.37 $X2=1.315 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__DLRTP_2%A_27_392# 1 2 7 9 12 16 18 19 21 22 25 27 30
c97 30 0 1.66318e-19 $X=2.675 $Y=1.605
c98 25 0 1.12738e-19 $X=2.595 $Y=2.44
r99 30 33 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.675 $Y=1.605
+ $X2=2.675 $Y2=1.77
r100 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.675
+ $Y=1.605 $X2=2.675 $Y2=1.605
r101 27 28 7.80343 $w=6.41e-07 $l=4.1e-07 $layer=LI1_cond $X=0.485 $Y=2.115
+ $X2=0.485 $Y2=2.525
r102 25 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.595 $Y=2.44
+ $X2=2.595 $Y2=1.77
r103 23 28 8.74498 $w=1.7e-07 $l=3.7e-07 $layer=LI1_cond $X=0.855 $Y=2.525
+ $X2=0.485 $Y2=2.525
r104 22 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.51 $Y=2.525
+ $X2=2.595 $Y2=2.44
r105 22 23 107.973 $w=1.68e-07 $l=1.655e-06 $layer=LI1_cond $X=2.51 $Y=2.525
+ $X2=0.855 $Y2=2.525
r106 21 27 10.6318 $w=6.41e-07 $l=3.5812e-07 $layer=LI1_cond $X=0.77 $Y=1.95
+ $X2=0.485 $Y2=2.115
r107 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.77 $Y=1.28
+ $X2=0.77 $Y2=1.95
r108 18 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.685 $Y=1.195
+ $X2=0.77 $Y2=1.28
r109 18 19 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=0.685 $Y=1.195
+ $X2=0.47 $Y2=1.195
r110 14 19 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.305 $Y=1.11
+ $X2=0.47 $Y2=1.195
r111 14 16 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=0.305 $Y=1.11
+ $X2=0.305 $Y2=0.835
r112 10 31 38.6072 $w=2.91e-07 $l=2.05122e-07 $layer=POLY_cond $X=2.765 $Y=1.44
+ $X2=2.675 $Y2=1.605
r113 10 12 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=2.765 $Y=1.44
+ $X2=2.765 $Y2=0.69
r114 7 31 57.6553 $w=2.91e-07 $l=3.15278e-07 $layer=POLY_cond $X=2.75 $Y=1.885
+ $X2=2.675 $Y2=1.605
r115 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.75 $Y=1.885
+ $X2=2.75 $Y2=2.46
r116 2 27 300 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.96 $X2=0.28 $Y2=2.115
r117 1 16 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=0.16
+ $Y=0.56 $X2=0.305 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_LS__DLRTP_2%A_347_98# 1 2 9 10 12 14 15 18 20 21 22 25
+ 32 36 40 46 49 51
c115 46 0 3.48291e-20 $X=3.215 $Y=1.285
c116 40 0 1.32977e-19 $X=3.135 $Y=2.025
c117 32 0 1.86781e-19 $X=2.23 $Y=1.085
c118 25 0 1.64562e-19 $X=3.895 $Y=2.215
r119 46 49 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.215 $Y=1.285
+ $X2=3.215 $Y2=1.12
r120 45 47 8.65224 $w=2.63e-07 $l=1.65e-07 $layer=LI1_cond $X=3.182 $Y=1.285
+ $X2=3.182 $Y2=1.45
r121 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.215
+ $Y=1.285 $X2=3.215 $Y2=1.285
r122 38 40 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=2.975 $Y=2.025
+ $X2=3.135 $Y2=2.025
r123 34 36 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=1.91 $Y=2.105
+ $X2=2.145 $Y2=2.105
r124 31 32 5.66838 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=2.145 $Y=1.085
+ $X2=2.23 $Y2=1.085
r125 29 31 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=1.88 $Y=1.085
+ $X2=2.145 $Y2=1.085
r126 26 51 25.1593 $w=3.64e-07 $l=1.9e-07 $layer=POLY_cond $X=3.895 $Y=2.257
+ $X2=3.705 $Y2=2.257
r127 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.895
+ $Y=2.215 $X2=3.895 $Y2=2.215
r128 23 25 24.0965 $w=3.28e-07 $l=6.9e-07 $layer=LI1_cond $X=3.895 $Y=2.905
+ $X2=3.895 $Y2=2.215
r129 21 23 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.73 $Y=2.99
+ $X2=3.895 $Y2=2.905
r130 21 22 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.73 $Y=2.99
+ $X2=3.06 $Y2=2.99
r131 20 40 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.135 $Y=1.94
+ $X2=3.135 $Y2=2.025
r132 20 47 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=3.135 $Y=1.94
+ $X2=3.135 $Y2=1.45
r133 18 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.975 $Y=2.905
+ $X2=3.06 $Y2=2.99
r134 17 38 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.975 $Y=2.11
+ $X2=2.975 $Y2=2.025
r135 17 18 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=2.975 $Y=2.11
+ $X2=2.975 $Y2=2.905
r136 15 45 5.21861 $w=2.63e-07 $l=1.2e-07 $layer=LI1_cond $X=3.182 $Y=1.165
+ $X2=3.182 $Y2=1.285
r137 15 32 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=3.05 $Y=1.165
+ $X2=2.23 $Y2=1.165
r138 14 36 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.145 $Y=1.94
+ $X2=2.145 $Y2=2.105
r139 13 31 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.145 $Y=1.25
+ $X2=2.145 $Y2=1.085
r140 13 14 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.145 $Y=1.25
+ $X2=2.145 $Y2=1.94
r141 10 51 23.572 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.705 $Y=2.465
+ $X2=3.705 $Y2=2.257
r142 10 12 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.705 $Y=2.465
+ $X2=3.705 $Y2=2.75
r143 9 49 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.155 $Y=0.69
+ $X2=3.155 $Y2=1.12
r144 2 34 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.765
+ $Y=1.96 $X2=1.91 $Y2=2.105
r145 1 29 182 $w=1.7e-07 $l=6.63551e-07 $layer=licon1_NDIFF $count=1 $X=1.735
+ $Y=0.49 $X2=1.88 $Y2=1.085
.ends

.subckt PM_SKY130_FD_SC_LS__DLRTP_2%A_832_55# 1 2 7 9 11 12 14 15 17 20 24 26 28
+ 31 33 40 46 48 50 52 55 56 57 70
c131 70 0 1.0789e-19 $X=6.645 $Y=1.532
c132 57 0 3.83707e-20 $X=5.34 $Y=1.72
c133 48 0 7.28255e-20 $X=6.05 $Y=1.805
c134 26 0 1.68639e-19 $X=6.66 $Y=1.765
r135 70 71 1.8491 $w=3.91e-07 $l=1.5e-08 $layer=POLY_cond $X=6.645 $Y=1.532
+ $X2=6.66 $Y2=1.532
r136 67 68 1.23274 $w=3.91e-07 $l=1e-08 $layer=POLY_cond $X=6.195 $Y=1.532
+ $X2=6.205 $Y2=1.532
r137 60 61 4.69791 $w=4.88e-07 $l=1.4e-07 $layer=LI1_cond $X=5.34 $Y=2.24
+ $X2=5.34 $Y2=2.38
r138 59 60 6.22449 $w=4.88e-07 $l=2.55e-07 $layer=LI1_cond $X=5.34 $Y=1.985
+ $X2=5.34 $Y2=2.24
r139 56 59 4.39376 $w=4.88e-07 $l=1.8e-07 $layer=LI1_cond $X=5.34 $Y=1.805
+ $X2=5.34 $Y2=1.985
r140 56 57 7.50345 $w=4.88e-07 $l=8.5e-08 $layer=LI1_cond $X=5.34 $Y=1.805
+ $X2=5.34 $Y2=1.72
r141 55 57 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=5.18 $Y=1.13
+ $X2=5.18 $Y2=1.72
r142 53 70 11.0946 $w=3.91e-07 $l=9e-08 $layer=POLY_cond $X=6.555 $Y=1.532
+ $X2=6.645 $Y2=1.532
r143 53 68 43.1458 $w=3.91e-07 $l=3.5e-07 $layer=POLY_cond $X=6.555 $Y=1.532
+ $X2=6.205 $Y2=1.532
r144 52 53 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.555
+ $Y=1.465 $X2=6.555 $Y2=1.465
r145 50 64 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=6.135 $Y=1.465
+ $X2=6.135 $Y2=1.805
r146 50 52 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=6.22 $Y=1.465
+ $X2=6.555 $Y2=1.465
r147 49 56 7.03003 $w=1.7e-07 $l=2.45e-07 $layer=LI1_cond $X=5.585 $Y=1.805
+ $X2=5.34 $Y2=1.805
r148 48 64 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.05 $Y=1.805
+ $X2=6.135 $Y2=1.805
r149 48 49 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=6.05 $Y=1.805
+ $X2=5.585 $Y2=1.805
r150 46 61 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=5.42 $Y=2.815
+ $X2=5.42 $Y2=2.38
r151 38 55 9.97136 $w=4.18e-07 $l=2.1e-07 $layer=LI1_cond $X=5.055 $Y=0.92
+ $X2=5.055 $Y2=1.13
r152 38 40 11.1128 $w=4.18e-07 $l=4.05e-07 $layer=LI1_cond $X=5.055 $Y=0.92
+ $X2=5.055 $Y2=0.515
r153 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.465
+ $Y=2.215 $X2=4.465 $Y2=2.215
r154 33 60 4.01183 $w=2.8e-07 $l=2.45e-07 $layer=LI1_cond $X=5.095 $Y=2.24
+ $X2=5.34 $Y2=2.24
r155 33 35 25.93 $w=2.78e-07 $l=6.3e-07 $layer=LI1_cond $X=5.095 $Y=2.24
+ $X2=4.465 $Y2=2.24
r156 29 31 71.7872 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=4.235 $Y=0.975
+ $X2=4.375 $Y2=0.975
r157 26 71 25.3065 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=6.66 $Y=1.765
+ $X2=6.66 $Y2=1.532
r158 26 28 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.66 $Y=1.765
+ $X2=6.66 $Y2=2.4
r159 22 70 25.3065 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=6.645 $Y=1.3
+ $X2=6.645 $Y2=1.532
r160 22 24 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=6.645 $Y=1.3
+ $X2=6.645 $Y2=0.74
r161 18 68 25.3065 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=6.205 $Y=1.3
+ $X2=6.205 $Y2=1.532
r162 18 20 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=6.205 $Y=1.3
+ $X2=6.205 $Y2=0.74
r163 15 67 25.3065 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=6.195 $Y=1.765
+ $X2=6.195 $Y2=1.532
r164 15 17 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.195 $Y=1.765
+ $X2=6.195 $Y2=2.4
r165 12 36 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=4.39 $Y=2.465
+ $X2=4.465 $Y2=2.215
r166 12 14 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.39 $Y=2.465
+ $X2=4.39 $Y2=2.75
r167 11 36 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=4.375 $Y=2.05
+ $X2=4.465 $Y2=2.215
r168 10 31 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.375 $Y=1.05
+ $X2=4.375 $Y2=0.975
r169 10 11 512.766 $w=1.5e-07 $l=1e-06 $layer=POLY_cond $X=4.375 $Y=1.05
+ $X2=4.375 $Y2=2.05
r170 7 29 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.235 $Y=0.9
+ $X2=4.235 $Y2=0.975
r171 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.235 $Y=0.9 $X2=4.235
+ $Y2=0.615
r172 2 59 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=5.27
+ $Y=1.84 $X2=5.42 $Y2=1.985
r173 2 46 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=5.27
+ $Y=1.84 $X2=5.42 $Y2=2.815
r174 1 40 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=4.865
+ $Y=0.37 $X2=5.01 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__DLRTP_2%A_646_74# 1 2 7 9 12 14 15 16 22 23 27 31 32
+ 34
c89 15 0 2.6214e-20 $X=5.105 $Y=1.35
c90 7 0 4.66116e-20 $X=5.195 $Y=1.765
r91 31 32 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.395 $Y=2.57
+ $X2=3.395 $Y2=2.405
r92 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.825
+ $Y=1.515 $X2=4.825 $Y2=1.515
r93 25 27 10.6547 $w=2.63e-07 $l=2.45e-07 $layer=LI1_cond $X=4.792 $Y=1.76
+ $X2=4.792 $Y2=1.515
r94 24 34 1.34256 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=3.655 $Y=1.845
+ $X2=3.522 $Y2=1.845
r95 23 25 7.24806 $w=1.7e-07 $l=1.69245e-07 $layer=LI1_cond $X=4.66 $Y=1.845
+ $X2=4.792 $Y2=1.76
r96 23 24 65.5668 $w=1.68e-07 $l=1.005e-06 $layer=LI1_cond $X=4.66 $Y=1.845
+ $X2=3.655 $Y2=1.845
r97 22 34 5.16603 $w=1.7e-07 $l=1.06325e-07 $layer=LI1_cond $X=3.57 $Y=1.76
+ $X2=3.522 $Y2=1.845
r98 21 22 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=3.57 $Y=0.845
+ $X2=3.57 $Y2=1.76
r99 19 34 5.16603 $w=1.7e-07 $l=1.05924e-07 $layer=LI1_cond $X=3.475 $Y=1.93
+ $X2=3.522 $Y2=1.845
r100 19 32 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=3.475 $Y=1.93
+ $X2=3.475 $Y2=2.405
r101 16 21 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.485 $Y=0.72
+ $X2=3.57 $Y2=0.845
r102 16 18 1.22 $w=2.5e-07 $l=2.5e-08 $layer=LI1_cond $X=3.485 $Y=0.72 $X2=3.46
+ $Y2=0.72
r103 14 28 48.9612 $w=3.3e-07 $l=2.8e-07 $layer=POLY_cond $X=5.105 $Y=1.515
+ $X2=4.825 $Y2=1.515
r104 14 15 5.03009 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.105 $Y=1.515
+ $X2=5.105 $Y2=1.35
r105 10 15 37.0704 $w=1.5e-07 $l=1.2e-07 $layer=POLY_cond $X=5.225 $Y=1.35
+ $X2=5.105 $Y2=1.35
r106 10 12 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.225 $Y=1.35
+ $X2=5.225 $Y2=0.74
r107 7 15 37.0704 $w=1.5e-07 $l=4.57794e-07 $layer=POLY_cond $X=5.195 $Y=1.765
+ $X2=5.105 $Y2=1.35
r108 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.195 $Y=1.765
+ $X2=5.195 $Y2=2.4
r109 2 31 600 $w=1.7e-07 $l=6.80882e-07 $layer=licon1_PDIFF $count=1 $X=3.245
+ $Y=1.96 $X2=3.395 $Y2=2.57
r110 1 18 182 $w=1.7e-07 $l=4.09145e-07 $layer=licon1_NDIFF $count=1 $X=3.23
+ $Y=0.37 $X2=3.46 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_LS__DLRTP_2%RESET_B 1 3 4 6 7 11
c35 1 0 3.83707e-20 $X=5.615 $Y=1.22
r36 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.675
+ $Y=1.385 $X2=5.675 $Y2=1.385
r37 7 11 4.8278 $w=3.68e-07 $l=1.55e-07 $layer=LI1_cond $X=5.52 $Y=1.365
+ $X2=5.675 $Y2=1.365
r38 4 10 77.2841 $w=2.7e-07 $l=3.94715e-07 $layer=POLY_cond $X=5.645 $Y=1.765
+ $X2=5.675 $Y2=1.385
r39 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.645 $Y=1.765
+ $X2=5.645 $Y2=2.4
r40 1 10 38.9026 $w=2.7e-07 $l=1.92678e-07 $layer=POLY_cond $X=5.615 $Y=1.22
+ $X2=5.675 $Y2=1.385
r41 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.615 $Y=1.22 $X2=5.615
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__DLRTP_2%VPWR 1 2 3 4 5 20 24 28 32 34 37 38 39 48 55
+ 60 66 69 76 80
c84 28 0 1.0789e-19 $X=5.92 $Y=2.145
r85 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r86 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r87 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r88 64 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6.96 $Y2=3.33
r89 64 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33 $X2=6
+ $Y2=3.33
r90 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r91 61 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.085 $Y=3.33
+ $X2=5.92 $Y2=3.33
r92 61 63 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=6.085 $Y=3.33
+ $X2=6.48 $Y2=3.33
r93 60 79 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=6.755 $Y=3.33
+ $X2=6.977 $Y2=3.33
r94 60 63 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.755 $Y=3.33
+ $X2=6.48 $Y2=3.33
r95 59 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33 $X2=6
+ $Y2=3.33
r96 59 73 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=4.56 $Y2=3.33
r97 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r98 56 58 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=5.085 $Y=3.33
+ $X2=5.52 $Y2=3.33
r99 55 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.755 $Y=3.33
+ $X2=5.92 $Y2=3.33
r100 55 58 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=5.755 $Y=3.33
+ $X2=5.52 $Y2=3.33
r101 54 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r102 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r103 50 53 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.64 $Y=3.33
+ $X2=4.08 $Y2=3.33
r104 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r105 48 56 8.68381 $w=1.7e-07 $l=3.18e-07 $layer=LI1_cond $X=4.767 $Y=3.33
+ $X2=5.085 $Y2=3.33
r106 48 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r107 48 69 9.70048 $w=6.33e-07 $l=5.15e-07 $layer=LI1_cond $X=4.767 $Y=3.33
+ $X2=4.767 $Y2=2.815
r108 48 53 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=4.45 $Y=3.33
+ $X2=4.08 $Y2=3.33
r109 47 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r110 46 47 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r111 44 47 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r112 44 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r113 43 46 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r114 43 44 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r115 41 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.98 $Y=3.33
+ $X2=0.815 $Y2=3.33
r116 41 43 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.98 $Y=3.33
+ $X2=1.2 $Y2=3.33
r117 39 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r118 39 51 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=2.64 $Y2=3.33
r119 37 46 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=2.28 $Y=3.33
+ $X2=2.16 $Y2=3.33
r120 37 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.28 $Y=3.33
+ $X2=2.445 $Y2=3.33
r121 36 50 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=2.61 $Y=3.33 $X2=2.64
+ $Y2=3.33
r122 36 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.61 $Y=3.33
+ $X2=2.445 $Y2=3.33
r123 32 79 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=6.92 $Y=3.245
+ $X2=6.977 $Y2=3.33
r124 32 34 32.8272 $w=3.28e-07 $l=9.4e-07 $layer=LI1_cond $X=6.92 $Y=3.245
+ $X2=6.92 $Y2=2.305
r125 28 31 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=5.92 $Y=2.145
+ $X2=5.92 $Y2=2.825
r126 26 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.92 $Y=3.245
+ $X2=5.92 $Y2=3.33
r127 26 31 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=5.92 $Y=3.245
+ $X2=5.92 $Y2=2.825
r128 22 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.445 $Y=3.245
+ $X2=2.445 $Y2=3.33
r129 22 24 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=2.445 $Y=3.245
+ $X2=2.445 $Y2=2.945
r130 18 66 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=3.245
+ $X2=0.815 $Y2=3.33
r131 18 20 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=0.815 $Y=3.245
+ $X2=0.815 $Y2=2.945
r132 5 34 300 $w=1.7e-07 $l=5.49773e-07 $layer=licon1_PDIFF $count=2 $X=6.735
+ $Y=1.84 $X2=6.92 $Y2=2.305
r133 4 31 400 $w=1.7e-07 $l=1.08038e-06 $layer=licon1_PDIFF $count=1 $X=5.72
+ $Y=1.84 $X2=5.92 $Y2=2.825
r134 4 28 400 $w=1.7e-07 $l=3.9246e-07 $layer=licon1_PDIFF $count=1 $X=5.72
+ $Y=1.84 $X2=5.92 $Y2=2.145
r135 3 69 600 $w=1.7e-07 $l=4.15331e-07 $layer=licon1_PDIFF $count=1 $X=4.465
+ $Y=2.54 $X2=4.765 $Y2=2.815
r136 2 24 600 $w=1.7e-07 $l=1.09622e-06 $layer=licon1_PDIFF $count=1 $X=2.21
+ $Y=1.96 $X2=2.445 $Y2=2.945
r137 1 20 600 $w=1.7e-07 $l=1.09622e-06 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.96 $X2=0.815 $Y2=2.945
.ends

.subckt PM_SKY130_FD_SC_LS__DLRTP_2%Q 1 2 9 11 13 15 16 17 24
c44 13 0 1.68639e-19 $X=6.42 $Y=2.825
r45 23 24 25.3036 $w=2.28e-07 $l=5.05e-07 $layer=LI1_cond $X=6.96 $Y=1.8
+ $X2=6.96 $Y2=1.295
r46 22 24 8.26753 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=6.96 $Y=1.13
+ $X2=6.96 $Y2=1.295
r47 19 21 13.6724 $w=2.32e-07 $l=2.6e-07 $layer=LI1_cond $X=6.42 $Y=1.885
+ $X2=6.42 $Y2=2.145
r48 18 19 2.55969 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.585 $Y=1.885
+ $X2=6.42 $Y2=1.885
r49 17 23 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=6.845 $Y=1.885
+ $X2=6.96 $Y2=1.8
r50 17 18 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=6.845 $Y=1.885
+ $X2=6.585 $Y2=1.885
r51 15 22 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=6.845 $Y=1.045
+ $X2=6.96 $Y2=1.13
r52 15 16 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=6.845 $Y=1.045
+ $X2=6.585 $Y2=1.045
r53 11 21 4.04823 $w=3.3e-07 $l=8e-08 $layer=LI1_cond $X=6.42 $Y=2.225 $X2=6.42
+ $Y2=2.145
r54 11 13 20.9535 $w=3.28e-07 $l=6e-07 $layer=LI1_cond $X=6.42 $Y=2.225 $X2=6.42
+ $Y2=2.825
r55 7 16 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.42 $Y=0.96
+ $X2=6.585 $Y2=1.045
r56 7 9 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=6.42 $Y=0.96 $X2=6.42
+ $Y2=0.515
r57 2 21 400 $w=1.7e-07 $l=3.72525e-07 $layer=licon1_PDIFF $count=1 $X=6.27
+ $Y=1.84 $X2=6.42 $Y2=2.145
r58 2 13 400 $w=1.7e-07 $l=1.05734e-06 $layer=licon1_PDIFF $count=1 $X=6.27
+ $Y=1.84 $X2=6.42 $Y2=2.825
r59 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.28
+ $Y=0.37 $X2=6.42 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__DLRTP_2%VGND 1 2 3 4 5 20 24 28 30 32 34 35 41 50 57
+ 62 68 71 74 78
c80 24 0 1.18818e-19 $X=4.45 $Y=0.615
r81 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r82 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r83 71 72 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r84 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r85 66 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6.96
+ $Y2=0
r86 66 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r87 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r88 63 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.085 $Y=0 $X2=5.92
+ $Y2=0
r89 63 65 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=6.085 $Y=0 $X2=6.48
+ $Y2=0
r90 62 77 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=6.755 $Y=0 $X2=6.977
+ $Y2=0
r91 62 65 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.755 $Y=0 $X2=6.48
+ $Y2=0
r92 61 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r93 61 72 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=4.56
+ $Y2=0
r94 60 61 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r95 58 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.615 $Y=0 $X2=4.45
+ $Y2=0
r96 58 60 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=4.615 $Y=0 $X2=5.52
+ $Y2=0
r97 57 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.755 $Y=0 $X2=5.92
+ $Y2=0
r98 57 60 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=5.755 $Y=0 $X2=5.52
+ $Y2=0
r99 56 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r100 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r101 52 55 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.64 $Y=0 $X2=4.08
+ $Y2=0
r102 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r103 50 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.285 $Y=0 $X2=4.45
+ $Y2=0
r104 50 55 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=4.285 $Y=0
+ $X2=4.08 $Y2=0
r105 49 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r106 48 49 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r107 46 49 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r108 46 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r109 45 48 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r110 45 46 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r111 43 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.98 $Y=0 $X2=0.815
+ $Y2=0
r112 43 45 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.98 $Y=0 $X2=1.2
+ $Y2=0
r113 41 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r114 41 53 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=2.64
+ $Y2=0
r115 37 52 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=2.635 $Y=0 $X2=2.64
+ $Y2=0
r116 35 48 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=2.305 $Y=0
+ $X2=2.16 $Y2=0
r117 34 39 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=2.47 $Y=0 $X2=2.47
+ $Y2=0.325
r118 34 37 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.47 $Y=0 $X2=2.635
+ $Y2=0
r119 34 35 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.47 $Y=0 $X2=2.305
+ $Y2=0
r120 30 77 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=6.92 $Y=0.085
+ $X2=6.977 $Y2=0
r121 30 32 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=6.92 $Y=0.085
+ $X2=6.92 $Y2=0.625
r122 26 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.92 $Y=0.085
+ $X2=5.92 $Y2=0
r123 26 28 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=5.92 $Y=0.085
+ $X2=5.92 $Y2=0.515
r124 22 71 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.45 $Y=0.085
+ $X2=4.45 $Y2=0
r125 22 24 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=4.45 $Y=0.085
+ $X2=4.45 $Y2=0.615
r126 18 68 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=0.085
+ $X2=0.815 $Y2=0
r127 18 20 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.815 $Y=0.085
+ $X2=0.815 $Y2=0.515
r128 5 32 182 $w=1.7e-07 $l=3.40624e-07 $layer=licon1_NDIFF $count=1 $X=6.72
+ $Y=0.37 $X2=6.92 $Y2=0.625
r129 4 28 91 $w=1.7e-07 $l=2.93684e-07 $layer=licon1_NDIFF $count=2 $X=5.69
+ $Y=0.37 $X2=5.92 $Y2=0.515
r130 3 24 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.31
+ $Y=0.405 $X2=4.45 $Y2=0.615
r131 2 39 182 $w=1.7e-07 $l=2.91033e-07 $layer=licon1_NDIFF $count=1 $X=2.25
+ $Y=0.49 $X2=2.47 $Y2=0.325
r132 1 20 91 $w=1.7e-07 $l=2.41454e-07 $layer=licon1_NDIFF $count=2 $X=0.595
+ $Y=0.56 $X2=0.815 $Y2=0.515
.ends

