* File: sky130_fd_sc_ls__and3b_1.pex.spice
* Created: Fri Aug 28 13:04:24 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__AND3B_1%A_N 3 9 12 13 14 15 16 17 21 22
r31 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.405
+ $Y=1.275 $X2=0.405 $Y2=1.275
r32 16 17 9.58211 $w=4.43e-07 $l=3.7e-07 $layer=LI1_cond $X=0.347 $Y=1.295
+ $X2=0.347 $Y2=1.665
r33 16 22 0.517952 $w=4.43e-07 $l=2e-08 $layer=LI1_cond $X=0.347 $Y=1.295
+ $X2=0.347 $Y2=1.275
r34 14 15 45.74 $w=1.65e-07 $l=1.05e-07 $layer=POLY_cond $X=0.502 $Y=1.94
+ $X2=0.502 $Y2=2.045
r35 13 14 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=0.495 $Y=1.78
+ $X2=0.495 $Y2=1.94
r36 12 21 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.405 $Y=1.615
+ $X2=0.405 $Y2=1.275
r37 12 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.405 $Y=1.615
+ $X2=0.405 $Y2=1.78
r38 11 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.405 $Y=1.11
+ $X2=0.405 $Y2=1.275
r39 9 15 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.51 $Y=2.54 $X2=0.51
+ $Y2=2.045
r40 3 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.495 $Y=0.645
+ $X2=0.495 $Y2=1.11
.ends

.subckt PM_SKY130_FD_SC_LS__AND3B_1%A_114_74# 1 2 9 12 13 15 16 18 19 22 26 28
+ 29 34 35 36
c68 34 0 7.864e-20 $X=0.975 $Y=1.195
r69 35 36 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=0.86 $Y=2.1 $X2=0.86
+ $Y2=1.7
r70 33 34 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.975
+ $Y=1.195 $X2=0.975 $Y2=1.195
r71 29 36 9.06106 $w=3.63e-07 $l=1.82e-07 $layer=LI1_cond $X=0.957 $Y=1.518
+ $X2=0.957 $Y2=1.7
r72 28 33 0.870046 $w=3.65e-07 $l=8.80909e-08 $layer=LI1_cond $X=0.957 $Y=1.212
+ $X2=0.877 $Y2=1.195
r73 28 29 9.66158 $w=3.63e-07 $l=3.06e-07 $layer=LI1_cond $X=0.957 $Y=1.212
+ $X2=0.957 $Y2=1.518
r74 26 35 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.78 $Y=2.265
+ $X2=0.78 $Y2=2.1
r75 20 33 15.5822 $w=3.3e-07 $l=4.65983e-07 $layer=LI1_cond $X=0.78 $Y=0.775
+ $X2=0.877 $Y2=1.195
r76 20 22 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=0.78 $Y=0.775
+ $X2=0.78 $Y2=0.645
r77 16 18 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.7 $Y=1.765 $X2=1.7
+ $Y2=2.26
r78 13 19 18.8402 $w=1.65e-07 $l=8e-08 $layer=POLY_cond $X=1.69 $Y=1.185
+ $X2=1.61 $Y2=1.185
r79 13 15 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.69 $Y=1.185
+ $X2=1.69 $Y2=0.79
r80 12 16 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.7 $Y=1.675 $X2=1.7
+ $Y2=1.765
r81 11 19 18.8402 $w=1.65e-07 $l=2.81425e-07 $layer=POLY_cond $X=1.7 $Y=1.425
+ $X2=1.61 $Y2=1.185
r82 11 12 97.1774 $w=1.8e-07 $l=2.5e-07 $layer=POLY_cond $X=1.7 $Y=1.425 $X2=1.7
+ $Y2=1.675
r83 10 34 19.7453 $w=1.5e-07 $l=2.00237e-07 $layer=POLY_cond $X=1.14 $Y=1.26
+ $X2=0.975 $Y2=1.182
r84 9 19 6.66866 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.61 $Y=1.26 $X2=1.61
+ $Y2=1.185
r85 9 10 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=1.61 $Y=1.26 $X2=1.14
+ $Y2=1.26
r86 2 26 300 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=2.12 $X2=0.78 $Y2=2.265
r87 1 22 182 $w=1.7e-07 $l=3.65205e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.78 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_LS__AND3B_1%B 3 5 7 8 12
r33 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.17
+ $Y=1.515 $X2=2.17 $Y2=1.515
r34 8 12 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=2.17 $Y=1.665
+ $X2=2.17 $Y2=1.515
r35 5 11 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=2.245 $Y=1.765
+ $X2=2.17 $Y2=1.515
r36 5 7 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.245 $Y=1.765
+ $X2=2.245 $Y2=2.26
r37 1 11 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=2.08 $Y=1.35
+ $X2=2.17 $Y2=1.515
r38 1 3 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.08 $Y=1.35 $X2=2.08
+ $Y2=0.79
.ends

.subckt PM_SKY130_FD_SC_LS__AND3B_1%C 3 5 7 8 12
c28 3 0 4.57304e-20 $X=2.62 $Y=0.79
r29 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.71
+ $Y=1.515 $X2=2.71 $Y2=1.515
r30 8 12 4.93904 $w=3.48e-07 $l=1.5e-07 $layer=LI1_cond $X=2.7 $Y=1.665 $X2=2.7
+ $Y2=1.515
r31 5 11 52.2586 $w=2.99e-07 $l=2.54951e-07 $layer=POLY_cond $X=2.7 $Y=1.765
+ $X2=2.71 $Y2=1.515
r32 5 7 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.7 $Y=1.765 $X2=2.7
+ $Y2=2.26
r33 1 11 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=2.62 $Y=1.35
+ $X2=2.71 $Y2=1.515
r34 1 3 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.62 $Y=1.35 $X2=2.62
+ $Y2=0.79
.ends

.subckt PM_SKY130_FD_SC_LS__AND3B_1%A_266_94# 1 2 3 10 12 15 19 22 25 27 31 33
+ 35
c86 19 0 7.864e-20 $X=1.475 $Y=0.615
c87 10 0 3.95737e-20 $X=3.285 $Y=1.765
r88 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.25
+ $Y=1.465 $X2=3.25 $Y2=1.465
r89 28 33 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.64 $Y=2.035
+ $X2=1.475 $Y2=2.035
r90 27 35 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.31 $Y=2.035
+ $X2=2.475 $Y2=2.035
r91 27 28 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.31 $Y=2.035
+ $X2=1.64 $Y2=2.035
r92 26 31 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.64 $Y=1.135
+ $X2=1.475 $Y2=1.135
r93 25 38 14.2261 $w=2.83e-07 $l=4.1225e-07 $layer=LI1_cond $X=3.045 $Y=1.135
+ $X2=3.23 $Y2=1.465
r94 25 26 91.6631 $w=1.68e-07 $l=1.405e-06 $layer=LI1_cond $X=3.045 $Y=1.135
+ $X2=1.64 $Y2=1.135
r95 22 33 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.475 $Y=1.95
+ $X2=1.475 $Y2=2.035
r96 21 31 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.475 $Y=1.22
+ $X2=1.475 $Y2=1.135
r97 21 22 25.4934 $w=3.28e-07 $l=7.3e-07 $layer=LI1_cond $X=1.475 $Y=1.22
+ $X2=1.475 $Y2=1.95
r98 17 31 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.475 $Y=1.05
+ $X2=1.475 $Y2=1.135
r99 17 19 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=1.475 $Y=1.05
+ $X2=1.475 $Y2=0.615
r100 13 39 38.6549 $w=2.86e-07 $l=2.03101e-07 $layer=POLY_cond $X=3.335 $Y=1.3
+ $X2=3.25 $Y2=1.465
r101 13 15 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.335 $Y=1.3
+ $X2=3.335 $Y2=0.74
r102 10 39 61.4066 $w=2.86e-07 $l=3.17017e-07 $layer=POLY_cond $X=3.285 $Y=1.765
+ $X2=3.25 $Y2=1.465
r103 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.285 $Y=1.765
+ $X2=3.285 $Y2=2.4
r104 3 35 300 $w=1.7e-07 $l=3.43875e-07 $layer=licon1_PDIFF $count=2 $X=2.32
+ $Y=1.84 $X2=2.475 $Y2=2.115
r105 2 33 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=1.33
+ $Y=1.84 $X2=1.475 $Y2=1.985
r106 1 19 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=1.33
+ $Y=0.47 $X2=1.475 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_LS__AND3B_1%VPWR 1 2 3 10 12 16 20 23 24 26 27 28 41 42
r45 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r46 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r47 39 42 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r48 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r49 35 36 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r50 33 36 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r51 33 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r52 32 35 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=3.33 $X2=1.68
+ $Y2=3.33
r53 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r54 30 45 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.222 $Y2=3.33
r55 30 32 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.72 $Y2=3.33
r56 28 39 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.64 $Y2=3.33
r57 28 36 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r58 26 38 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=2.845 $Y=3.33
+ $X2=2.64 $Y2=3.33
r59 26 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.845 $Y=3.33
+ $X2=3.01 $Y2=3.33
r60 25 41 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=3.175 $Y=3.33
+ $X2=3.6 $Y2=3.33
r61 25 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.175 $Y=3.33
+ $X2=3.01 $Y2=3.33
r62 23 35 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=1.81 $Y=3.33
+ $X2=1.68 $Y2=3.33
r63 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.81 $Y=3.33
+ $X2=1.975 $Y2=3.33
r64 22 38 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=2.14 $Y=3.33 $X2=2.64
+ $Y2=3.33
r65 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.14 $Y=3.33
+ $X2=1.975 $Y2=3.33
r66 18 27 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.01 $Y=3.245
+ $X2=3.01 $Y2=3.33
r67 18 20 39.4624 $w=3.28e-07 $l=1.13e-06 $layer=LI1_cond $X=3.01 $Y=3.245
+ $X2=3.01 $Y2=2.115
r68 14 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.975 $Y=3.245
+ $X2=1.975 $Y2=3.33
r69 14 16 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=1.975 $Y=3.245
+ $X2=1.975 $Y2=2.455
r70 10 45 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.222 $Y2=3.33
r71 10 12 34.2241 $w=3.28e-07 $l=9.8e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.28 $Y2=2.265
r72 3 20 300 $w=1.7e-07 $l=3.745e-07 $layer=licon1_PDIFF $count=2 $X=2.775
+ $Y=1.84 $X2=3.01 $Y2=2.115
r73 2 16 600 $w=1.7e-07 $l=7.07972e-07 $layer=licon1_PDIFF $count=1 $X=1.775
+ $Y=1.84 $X2=1.975 $Y2=2.455
r74 1 12 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.12 $X2=0.28 $Y2=2.265
.ends

.subckt PM_SKY130_FD_SC_LS__AND3B_1%X 1 2 9 13 14 15 16 23 33 34
c23 13 0 8.53041e-20 $X=3.57 $Y=1.13
r24 33 34 8.69073 $w=4.08e-07 $l=1.65e-07 $layer=LI1_cond $X=3.55 $Y=1.985
+ $X2=3.55 $Y2=1.82
r25 21 23 0.281084 $w=4.08e-07 $l=1e-08 $layer=LI1_cond $X=3.55 $Y=2.025
+ $X2=3.55 $Y2=2.035
r26 16 30 1.12433 $w=4.08e-07 $l=4e-08 $layer=LI1_cond $X=3.55 $Y=2.775 $X2=3.55
+ $Y2=2.815
r27 15 16 10.4001 $w=4.08e-07 $l=3.7e-07 $layer=LI1_cond $X=3.55 $Y=2.405
+ $X2=3.55 $Y2=2.775
r28 14 21 1.06812 $w=4.08e-07 $l=3.8e-08 $layer=LI1_cond $X=3.55 $Y=1.987
+ $X2=3.55 $Y2=2.025
r29 14 33 0.0562167 $w=4.08e-07 $l=2e-09 $layer=LI1_cond $X=3.55 $Y=1.987
+ $X2=3.55 $Y2=1.985
r30 14 15 9.36009 $w=4.08e-07 $l=3.33e-07 $layer=LI1_cond $X=3.55 $Y=2.072
+ $X2=3.55 $Y2=2.405
r31 14 23 1.04001 $w=4.08e-07 $l=3.7e-08 $layer=LI1_cond $X=3.55 $Y=2.072
+ $X2=3.55 $Y2=2.035
r32 13 34 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.67 $Y=1.13 $X2=3.67
+ $Y2=1.82
r33 7 13 9.16175 $w=3.68e-07 $l=1.85e-07 $layer=LI1_cond $X=3.57 $Y=0.945
+ $X2=3.57 $Y2=1.13
r34 7 9 13.3933 $w=3.68e-07 $l=4.3e-07 $layer=LI1_cond $X=3.57 $Y=0.945 $X2=3.57
+ $Y2=0.515
r35 2 33 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=3.36
+ $Y=1.84 $X2=3.51 $Y2=1.985
r36 2 30 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=3.36
+ $Y=1.84 $X2=3.51 $Y2=2.815
r37 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.41
+ $Y=0.37 $X2=3.55 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__AND3B_1%VGND 1 2 7 9 13 15 17 24 25 31
r35 32 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r36 31 34 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r37 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r38 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r39 25 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r40 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r41 22 31 12.4404 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=3.215 $Y=0 $X2=2.92
+ $Y2=0
r42 22 24 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=3.215 $Y=0 $X2=3.6
+ $Y2=0
r43 21 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r44 20 21 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r45 18 28 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.222
+ $Y2=0
r46 18 20 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.72
+ $Y2=0
r47 17 31 12.4404 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=2.625 $Y=0 $X2=2.92
+ $Y2=0
r48 17 20 124.283 $w=1.68e-07 $l=1.905e-06 $layer=LI1_cond $X=2.625 $Y=0
+ $X2=0.72 $Y2=0
r49 15 34 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.64
+ $Y2=0
r50 15 21 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.92 $Y=0 $X2=0.72
+ $Y2=0
r51 11 31 2.48142 $w=5.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.92 $Y=0.085
+ $X2=2.92 $Y2=0
r52 11 13 8.31173 $w=5.88e-07 $l=4.1e-07 $layer=LI1_cond $X=2.92 $Y=0.085
+ $X2=2.92 $Y2=0.495
r53 7 28 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.222 $Y2=0
r54 7 9 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=0.28 $Y=0.085 $X2=0.28
+ $Y2=0.645
r55 2 13 91 $w=1.7e-07 $l=4.37321e-07 $layer=licon1_NDIFF $count=2 $X=2.695
+ $Y=0.47 $X2=3.12 $Y2=0.495
r56 1 9 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.645
.ends

