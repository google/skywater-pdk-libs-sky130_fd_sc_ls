* File: sky130_fd_sc_ls__or4_2.pxi.spice
* Created: Fri Aug 28 13:59:44 2020
* 
x_PM_SKY130_FD_SC_LS__OR4_2%D N_D_M1004_g N_D_c_67_n N_D_M1000_g D
+ PM_SKY130_FD_SC_LS__OR4_2%D
x_PM_SKY130_FD_SC_LS__OR4_2%C N_C_M1007_g N_C_c_98_n N_C_c_102_n N_C_M1011_g C C
+ C C N_C_c_99_n N_C_c_100_n PM_SKY130_FD_SC_LS__OR4_2%C
x_PM_SKY130_FD_SC_LS__OR4_2%B N_B_c_142_n N_B_M1009_g N_B_M1001_g B B B B
+ N_B_c_144_n PM_SKY130_FD_SC_LS__OR4_2%B
x_PM_SKY130_FD_SC_LS__OR4_2%A N_A_c_178_n N_A_M1003_g N_A_M1006_g A N_A_c_180_n
+ PM_SKY130_FD_SC_LS__OR4_2%A
x_PM_SKY130_FD_SC_LS__OR4_2%A_85_392# N_A_85_392#_M1004_d N_A_85_392#_M1001_d
+ N_A_85_392#_M1000_s N_A_85_392#_c_220_n N_A_85_392#_M1005_g
+ N_A_85_392#_M1002_g N_A_85_392#_c_221_n N_A_85_392#_M1010_g
+ N_A_85_392#_M1008_g N_A_85_392#_c_213_n N_A_85_392#_c_229_n
+ N_A_85_392#_c_214_n N_A_85_392#_c_223_n N_A_85_392#_c_215_n
+ N_A_85_392#_c_241_n N_A_85_392#_c_216_n N_A_85_392#_c_217_n
+ N_A_85_392#_c_224_n N_A_85_392#_c_236_n N_A_85_392#_c_218_n
+ N_A_85_392#_c_219_n PM_SKY130_FD_SC_LS__OR4_2%A_85_392#
x_PM_SKY130_FD_SC_LS__OR4_2%VPWR N_VPWR_M1003_d N_VPWR_M1010_s N_VPWR_c_325_n
+ N_VPWR_c_326_n N_VPWR_c_327_n N_VPWR_c_328_n N_VPWR_c_329_n VPWR
+ N_VPWR_c_330_n N_VPWR_c_324_n PM_SKY130_FD_SC_LS__OR4_2%VPWR
x_PM_SKY130_FD_SC_LS__OR4_2%X N_X_M1002_d N_X_M1005_d N_X_c_366_n N_X_c_362_n
+ N_X_c_367_n N_X_c_368_n N_X_c_363_n N_X_c_364_n X X
+ PM_SKY130_FD_SC_LS__OR4_2%X
x_PM_SKY130_FD_SC_LS__OR4_2%VGND N_VGND_M1004_s N_VGND_M1007_d N_VGND_M1006_d
+ N_VGND_M1008_s N_VGND_c_403_n N_VGND_c_404_n N_VGND_c_405_n N_VGND_c_406_n
+ N_VGND_c_407_n N_VGND_c_408_n N_VGND_c_409_n VGND N_VGND_c_410_n
+ N_VGND_c_411_n N_VGND_c_412_n N_VGND_c_413_n N_VGND_c_414_n
+ PM_SKY130_FD_SC_LS__OR4_2%VGND
cc_1 VNB N_D_M1004_g 0.0374614f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=0.69
cc_2 VNB N_D_c_67_n 0.021515f $X=-0.19 $Y=-0.245 $X2=0.795 $Y2=1.885
cc_3 VNB D 0.00789517f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_4 VNB N_C_M1007_g 0.0228946f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=0.69
cc_5 VNB N_C_c_98_n 0.00776858f $X=-0.19 $Y=-0.245 $X2=0.795 $Y2=2.46
cc_6 VNB N_C_c_99_n 0.0352858f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_C_c_100_n 0.00391066f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_B_c_142_n 0.0274531f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.44
cc_9 VNB N_B_M1001_g 0.0326694f $X=-0.19 $Y=-0.245 $X2=0.795 $Y2=2.46
cc_10 VNB N_B_c_144_n 0.00238742f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_c_178_n 0.0252743f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.44
cc_12 VNB N_A_M1006_g 0.0315486f $X=-0.19 $Y=-0.245 $X2=0.795 $Y2=2.46
cc_13 VNB N_A_c_180_n 0.00428428f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.605
cc_14 VNB N_A_85_392#_M1002_g 0.0237774f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_85_392#_M1008_g 0.0232511f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_85_392#_c_213_n 0.0315891f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_85_392#_c_214_n 0.00803133f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_85_392#_c_215_n 0.00239958f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_85_392#_c_216_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_85_392#_c_217_n 0.0209257f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_85_392#_c_218_n 0.00754266f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_85_392#_c_219_n 0.0551076f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VPWR_c_324_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_X_c_362_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_X_c_363_n 0.00895476f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_X_c_364_n 0.00250148f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB X 0.0271747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_403_n 0.013467f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.295
cc_29 VNB N_VGND_c_404_n 0.0250687f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_405_n 0.0193312f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_406_n 0.0111136f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_407_n 0.0100164f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_408_n 0.0120272f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_409_n 0.0251975f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_410_n 0.019013f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_411_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_412_n 0.00923268f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_413_n 0.00836712f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_414_n 0.221765f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VPB N_D_c_67_n 0.0520901f $X=-0.19 $Y=1.66 $X2=0.795 $Y2=1.885
cc_41 VPB D 4.86891e-19 $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_42 VPB N_C_c_98_n 0.00605085f $X=-0.19 $Y=1.66 $X2=0.795 $Y2=2.46
cc_43 VPB N_C_c_102_n 0.0197198f $X=-0.19 $Y=1.66 $X2=0.795 $Y2=2.46
cc_44 VPB N_C_c_100_n 0.00453059f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_45 VPB N_B_c_142_n 0.0344136f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.44
cc_46 VPB N_B_c_144_n 0.00311922f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB N_A_c_178_n 0.0377374f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.44
cc_48 VPB N_A_c_180_n 0.0079905f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.605
cc_49 VPB N_A_85_392#_c_220_n 0.0166035f $X=-0.19 $Y=1.66 $X2=0.655 $Y2=1.605
cc_50 VPB N_A_85_392#_c_221_n 0.016419f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_51 VPB N_A_85_392#_c_213_n 0.0142037f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_A_85_392#_c_223_n 0.0358679f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_A_85_392#_c_224_n 0.0280007f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_A_85_392#_c_219_n 0.0141822f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_325_n 0.00936647f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_326_n 0.0133073f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.295
cc_57 VPB N_VPWR_c_327_n 0.0438947f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_328_n 0.0703865f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_329_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_330_n 0.0186948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_324_n 0.0968228f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_X_c_366_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_X_c_367_n 0.0105469f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_X_c_368_n 0.00220939f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB X 0.00739632f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 N_D_M1004_g N_C_M1007_g 0.0252464f $X=0.64 $Y=0.69 $X2=0 $Y2=0
cc_67 N_D_c_67_n N_C_c_98_n 0.0154464f $X=0.795 $Y=1.885 $X2=0 $Y2=0
cc_68 D N_C_c_98_n 7.37299e-19 $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_69 N_D_c_67_n N_C_c_102_n 0.0525551f $X=0.795 $Y=1.885 $X2=0 $Y2=0
cc_70 N_D_c_67_n N_C_c_99_n 0.0028993f $X=0.795 $Y=1.885 $X2=0 $Y2=0
cc_71 D N_C_c_99_n 0.00212694f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_72 N_D_M1004_g N_C_c_100_n 3.59156e-19 $X=0.64 $Y=0.69 $X2=0 $Y2=0
cc_73 N_D_c_67_n N_C_c_100_n 0.0125974f $X=0.795 $Y=1.885 $X2=0 $Y2=0
cc_74 D N_C_c_100_n 0.0484939f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_75 N_D_M1004_g N_A_85_392#_c_213_n 0.00675107f $X=0.64 $Y=0.69 $X2=0 $Y2=0
cc_76 N_D_c_67_n N_A_85_392#_c_213_n 0.0133259f $X=0.795 $Y=1.885 $X2=0 $Y2=0
cc_77 D N_A_85_392#_c_213_n 0.0461938f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_78 N_D_M1004_g N_A_85_392#_c_229_n 0.0103047f $X=0.64 $Y=0.69 $X2=0 $Y2=0
cc_79 N_D_c_67_n N_A_85_392#_c_229_n 4.63018e-19 $X=0.795 $Y=1.885 $X2=0 $Y2=0
cc_80 D N_A_85_392#_c_229_n 0.0175441f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_81 N_D_c_67_n N_A_85_392#_c_223_n 0.0112378f $X=0.795 $Y=1.885 $X2=0 $Y2=0
cc_82 N_D_M1004_g N_A_85_392#_c_215_n 0.0111125f $X=0.64 $Y=0.69 $X2=0 $Y2=0
cc_83 N_D_c_67_n N_A_85_392#_c_224_n 0.0111403f $X=0.795 $Y=1.885 $X2=0 $Y2=0
cc_84 D N_A_85_392#_c_224_n 0.0243567f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_85 N_D_M1004_g N_A_85_392#_c_236_n 7.30818e-19 $X=0.64 $Y=0.69 $X2=0 $Y2=0
cc_86 D N_A_85_392#_c_236_n 0.00964857f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_87 N_D_c_67_n N_VPWR_c_328_n 0.00445602f $X=0.795 $Y=1.885 $X2=0 $Y2=0
cc_88 N_D_c_67_n N_VPWR_c_324_n 0.00862959f $X=0.795 $Y=1.885 $X2=0 $Y2=0
cc_89 N_D_M1004_g N_VGND_c_404_n 0.0106017f $X=0.64 $Y=0.69 $X2=0 $Y2=0
cc_90 N_D_M1004_g N_VGND_c_405_n 0.00434272f $X=0.64 $Y=0.69 $X2=0 $Y2=0
cc_91 N_D_M1004_g N_VGND_c_414_n 0.00446102f $X=0.64 $Y=0.69 $X2=0 $Y2=0
cc_92 N_C_c_98_n N_B_c_142_n 0.0201388f $X=1.215 $Y=1.795 $X2=-0.19 $Y2=-0.245
cc_93 N_C_c_102_n N_B_c_142_n 0.0578169f $X=1.215 $Y=1.885 $X2=-0.19 $Y2=-0.245
cc_94 N_C_c_99_n N_B_c_142_n 0.00887637f $X=1.17 $Y=1.33 $X2=-0.19 $Y2=-0.245
cc_95 N_C_c_100_n N_B_c_142_n 0.0037741f $X=1.17 $Y=1.33 $X2=-0.19 $Y2=-0.245
cc_96 N_C_M1007_g N_B_M1001_g 0.015666f $X=1.07 $Y=0.69 $X2=0 $Y2=0
cc_97 N_C_c_99_n N_B_M1001_g 0.00602707f $X=1.17 $Y=1.33 $X2=0 $Y2=0
cc_98 N_C_c_100_n N_B_M1001_g 0.00103009f $X=1.17 $Y=1.33 $X2=0 $Y2=0
cc_99 N_C_c_98_n N_B_c_144_n 4.73511e-19 $X=1.215 $Y=1.795 $X2=0 $Y2=0
cc_100 N_C_c_102_n N_B_c_144_n 8.85319e-19 $X=1.215 $Y=1.885 $X2=0 $Y2=0
cc_101 N_C_c_99_n N_B_c_144_n 5.07843e-19 $X=1.17 $Y=1.33 $X2=0 $Y2=0
cc_102 N_C_c_100_n N_B_c_144_n 0.0408537f $X=1.17 $Y=1.33 $X2=0 $Y2=0
cc_103 N_C_c_102_n N_A_85_392#_c_223_n 0.00111334f $X=1.215 $Y=1.885 $X2=0 $Y2=0
cc_104 N_C_c_100_n N_A_85_392#_c_223_n 0.0424697f $X=1.17 $Y=1.33 $X2=0 $Y2=0
cc_105 N_C_M1007_g N_A_85_392#_c_215_n 0.0111125f $X=1.07 $Y=0.69 $X2=0 $Y2=0
cc_106 N_C_M1007_g N_A_85_392#_c_241_n 0.00969478f $X=1.07 $Y=0.69 $X2=0 $Y2=0
cc_107 N_C_c_99_n N_A_85_392#_c_241_n 0.00119292f $X=1.17 $Y=1.33 $X2=0 $Y2=0
cc_108 N_C_c_100_n N_A_85_392#_c_241_n 0.022264f $X=1.17 $Y=1.33 $X2=0 $Y2=0
cc_109 N_C_c_100_n N_A_85_392#_c_224_n 0.0096832f $X=1.17 $Y=1.33 $X2=0 $Y2=0
cc_110 N_C_M1007_g N_A_85_392#_c_236_n 0.00105683f $X=1.07 $Y=0.69 $X2=0 $Y2=0
cc_111 N_C_c_100_n N_A_85_392#_c_236_n 0.00118071f $X=1.17 $Y=1.33 $X2=0 $Y2=0
cc_112 N_C_c_100_n N_A_85_392#_c_218_n 4.4735e-19 $X=1.17 $Y=1.33 $X2=0 $Y2=0
cc_113 N_C_c_100_n A_174_392# 0.0105191f $X=1.17 $Y=1.33 $X2=-0.19 $Y2=-0.245
cc_114 N_C_c_102_n N_VPWR_c_328_n 0.00303293f $X=1.215 $Y=1.885 $X2=0 $Y2=0
cc_115 N_C_c_100_n N_VPWR_c_328_n 0.00865352f $X=1.17 $Y=1.33 $X2=0 $Y2=0
cc_116 N_C_c_102_n N_VPWR_c_324_n 0.00371687f $X=1.215 $Y=1.885 $X2=0 $Y2=0
cc_117 N_C_c_100_n N_VPWR_c_324_n 0.0106888f $X=1.17 $Y=1.33 $X2=0 $Y2=0
cc_118 N_C_M1007_g N_VGND_c_405_n 0.00434272f $X=1.07 $Y=0.69 $X2=0 $Y2=0
cc_119 N_C_M1007_g N_VGND_c_406_n 0.00601649f $X=1.07 $Y=0.69 $X2=0 $Y2=0
cc_120 N_C_M1007_g N_VGND_c_414_n 0.00444353f $X=1.07 $Y=0.69 $X2=0 $Y2=0
cc_121 N_B_c_142_n N_A_c_178_n 0.0514021f $X=1.635 $Y=1.885 $X2=-0.19 $Y2=-0.245
cc_122 N_B_c_144_n N_A_c_178_n 0.0133798f $X=1.71 $Y=1.515 $X2=-0.19 $Y2=-0.245
cc_123 N_B_M1001_g N_A_M1006_g 0.0217822f $X=1.81 $Y=0.69 $X2=0 $Y2=0
cc_124 N_B_c_142_n N_A_c_180_n 0.00236361f $X=1.635 $Y=1.885 $X2=0 $Y2=0
cc_125 N_B_c_144_n N_A_c_180_n 0.0350381f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_126 N_B_c_142_n N_A_85_392#_c_241_n 9.55021e-19 $X=1.635 $Y=1.885 $X2=0 $Y2=0
cc_127 N_B_M1001_g N_A_85_392#_c_241_n 0.0110935f $X=1.81 $Y=0.69 $X2=0 $Y2=0
cc_128 N_B_c_144_n N_A_85_392#_c_241_n 0.0124554f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_129 N_B_M1001_g N_A_85_392#_c_216_n 0.0111125f $X=1.81 $Y=0.69 $X2=0 $Y2=0
cc_130 N_B_M1001_g N_A_85_392#_c_218_n 0.0112764f $X=1.81 $Y=0.69 $X2=0 $Y2=0
cc_131 N_B_c_144_n N_A_85_392#_c_218_n 0.00110046f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_132 N_B_c_144_n A_342_392# 0.0143476f $X=1.71 $Y=1.515 $X2=-0.19 $Y2=-0.245
cc_133 N_B_c_144_n N_VPWR_c_325_n 0.0346485f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_134 N_B_c_142_n N_VPWR_c_328_n 0.00303293f $X=1.635 $Y=1.885 $X2=0 $Y2=0
cc_135 N_B_c_144_n N_VPWR_c_328_n 0.00909385f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_136 N_B_c_142_n N_VPWR_c_324_n 0.00373008f $X=1.635 $Y=1.885 $X2=0 $Y2=0
cc_137 N_B_c_144_n N_VPWR_c_324_n 0.0106888f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_138 N_B_M1001_g N_VGND_c_406_n 0.00601649f $X=1.81 $Y=0.69 $X2=0 $Y2=0
cc_139 N_B_M1001_g N_VGND_c_410_n 0.00434272f $X=1.81 $Y=0.69 $X2=0 $Y2=0
cc_140 N_B_M1001_g N_VGND_c_414_n 0.00444353f $X=1.81 $Y=0.69 $X2=0 $Y2=0
cc_141 N_A_c_178_n N_A_85_392#_c_220_n 0.0260756f $X=2.215 $Y=1.885 $X2=0 $Y2=0
cc_142 N_A_c_180_n N_A_85_392#_c_220_n 3.41323e-19 $X=2.29 $Y=1.515 $X2=0 $Y2=0
cc_143 N_A_M1006_g N_A_85_392#_M1002_g 0.015669f $X=2.24 $Y=0.69 $X2=0 $Y2=0
cc_144 N_A_M1006_g N_A_85_392#_c_216_n 0.00540115f $X=2.24 $Y=0.69 $X2=0 $Y2=0
cc_145 N_A_c_178_n N_A_85_392#_c_217_n 0.00276349f $X=2.215 $Y=1.885 $X2=0 $Y2=0
cc_146 N_A_M1006_g N_A_85_392#_c_217_n 0.0160107f $X=2.24 $Y=0.69 $X2=0 $Y2=0
cc_147 N_A_c_180_n N_A_85_392#_c_217_n 0.0429165f $X=2.29 $Y=1.515 $X2=0 $Y2=0
cc_148 N_A_c_178_n N_A_85_392#_c_218_n 3.13347e-19 $X=2.215 $Y=1.885 $X2=0 $Y2=0
cc_149 N_A_M1006_g N_A_85_392#_c_218_n 0.0073033f $X=2.24 $Y=0.69 $X2=0 $Y2=0
cc_150 N_A_c_180_n N_A_85_392#_c_218_n 0.012571f $X=2.29 $Y=1.515 $X2=0 $Y2=0
cc_151 N_A_c_178_n N_A_85_392#_c_219_n 0.0184557f $X=2.215 $Y=1.885 $X2=0 $Y2=0
cc_152 N_A_M1006_g N_A_85_392#_c_219_n 0.00129529f $X=2.24 $Y=0.69 $X2=0 $Y2=0
cc_153 N_A_c_180_n N_A_85_392#_c_219_n 0.00261926f $X=2.29 $Y=1.515 $X2=0 $Y2=0
cc_154 N_A_c_178_n N_VPWR_c_325_n 0.0191498f $X=2.215 $Y=1.885 $X2=0 $Y2=0
cc_155 N_A_c_180_n N_VPWR_c_325_n 0.00829271f $X=2.29 $Y=1.515 $X2=0 $Y2=0
cc_156 N_A_c_178_n N_VPWR_c_328_n 0.00461464f $X=2.215 $Y=1.885 $X2=0 $Y2=0
cc_157 N_A_c_178_n N_VPWR_c_324_n 0.00911352f $X=2.215 $Y=1.885 $X2=0 $Y2=0
cc_158 N_A_M1006_g N_X_c_362_n 6.55935e-19 $X=2.24 $Y=0.69 $X2=0 $Y2=0
cc_159 N_A_c_178_n N_X_c_368_n 6.76073e-19 $X=2.215 $Y=1.885 $X2=0 $Y2=0
cc_160 N_A_M1006_g N_X_c_364_n 2.87707e-19 $X=2.24 $Y=0.69 $X2=0 $Y2=0
cc_161 N_A_M1006_g N_VGND_c_407_n 0.00699865f $X=2.24 $Y=0.69 $X2=0 $Y2=0
cc_162 N_A_M1006_g N_VGND_c_410_n 0.00434272f $X=2.24 $Y=0.69 $X2=0 $Y2=0
cc_163 N_A_M1006_g N_VGND_c_414_n 0.00822102f $X=2.24 $Y=0.69 $X2=0 $Y2=0
cc_164 N_A_85_392#_c_220_n N_VPWR_c_325_n 0.00849498f $X=2.8 $Y=1.765 $X2=0
+ $Y2=0
cc_165 N_A_85_392#_c_217_n N_VPWR_c_325_n 0.00311314f $X=2.625 $Y=1.095 $X2=0
+ $Y2=0
cc_166 N_A_85_392#_c_221_n N_VPWR_c_327_n 0.0198182f $X=3.25 $Y=1.765 $X2=0
+ $Y2=0
cc_167 N_A_85_392#_c_223_n N_VPWR_c_328_n 0.0145938f $X=0.57 $Y=2.815 $X2=0
+ $Y2=0
cc_168 N_A_85_392#_c_220_n N_VPWR_c_330_n 0.00445602f $X=2.8 $Y=1.765 $X2=0
+ $Y2=0
cc_169 N_A_85_392#_c_221_n N_VPWR_c_330_n 0.00445602f $X=3.25 $Y=1.765 $X2=0
+ $Y2=0
cc_170 N_A_85_392#_c_220_n N_VPWR_c_324_n 0.0085808f $X=2.8 $Y=1.765 $X2=0 $Y2=0
cc_171 N_A_85_392#_c_221_n N_VPWR_c_324_n 0.00860661f $X=3.25 $Y=1.765 $X2=0
+ $Y2=0
cc_172 N_A_85_392#_c_223_n N_VPWR_c_324_n 0.0120466f $X=0.57 $Y=2.815 $X2=0
+ $Y2=0
cc_173 N_A_85_392#_c_220_n N_X_c_366_n 0.0107497f $X=2.8 $Y=1.765 $X2=0 $Y2=0
cc_174 N_A_85_392#_c_221_n N_X_c_366_n 0.0165744f $X=3.25 $Y=1.765 $X2=0 $Y2=0
cc_175 N_A_85_392#_M1002_g N_X_c_362_n 0.00876649f $X=2.915 $Y=0.74 $X2=0 $Y2=0
cc_176 N_A_85_392#_M1008_g N_X_c_362_n 3.97481e-19 $X=3.345 $Y=0.74 $X2=0 $Y2=0
cc_177 N_A_85_392#_c_221_n N_X_c_367_n 0.0154459f $X=3.25 $Y=1.765 $X2=0 $Y2=0
cc_178 N_A_85_392#_c_219_n N_X_c_367_n 0.00256871f $X=3.25 $Y=1.532 $X2=0 $Y2=0
cc_179 N_A_85_392#_c_220_n N_X_c_368_n 0.00412323f $X=2.8 $Y=1.765 $X2=0 $Y2=0
cc_180 N_A_85_392#_c_221_n N_X_c_368_n 0.0011347f $X=3.25 $Y=1.765 $X2=0 $Y2=0
cc_181 N_A_85_392#_c_217_n N_X_c_368_n 0.0151863f $X=2.625 $Y=1.095 $X2=0 $Y2=0
cc_182 N_A_85_392#_c_219_n N_X_c_368_n 0.00600344f $X=3.25 $Y=1.532 $X2=0 $Y2=0
cc_183 N_A_85_392#_M1008_g N_X_c_363_n 0.0156857f $X=3.345 $Y=0.74 $X2=0 $Y2=0
cc_184 N_A_85_392#_M1002_g N_X_c_364_n 0.00302365f $X=2.915 $Y=0.74 $X2=0 $Y2=0
cc_185 N_A_85_392#_c_217_n N_X_c_364_n 0.0121973f $X=2.625 $Y=1.095 $X2=0 $Y2=0
cc_186 N_A_85_392#_c_219_n N_X_c_364_n 0.00306094f $X=3.25 $Y=1.532 $X2=0 $Y2=0
cc_187 N_A_85_392#_c_221_n X 0.0012197f $X=3.25 $Y=1.765 $X2=0 $Y2=0
cc_188 N_A_85_392#_M1008_g X 0.0117876f $X=3.345 $Y=0.74 $X2=0 $Y2=0
cc_189 N_A_85_392#_c_217_n X 0.0125557f $X=2.625 $Y=1.095 $X2=0 $Y2=0
cc_190 N_A_85_392#_c_219_n X 0.0103954f $X=3.25 $Y=1.532 $X2=0 $Y2=0
cc_191 N_A_85_392#_c_213_n N_VGND_M1004_s 2.73857e-19 $X=0.17 $Y=1.94 $X2=-0.19
+ $Y2=-0.245
cc_192 N_A_85_392#_c_229_n N_VGND_M1004_s 0.0111118f $X=0.69 $Y=0.91 $X2=-0.19
+ $Y2=-0.245
cc_193 N_A_85_392#_c_214_n N_VGND_M1004_s 0.00243753f $X=0.255 $Y=0.91 $X2=-0.19
+ $Y2=-0.245
cc_194 N_A_85_392#_c_241_n N_VGND_M1007_d 0.0178395f $X=1.86 $Y=0.91 $X2=0 $Y2=0
cc_195 N_A_85_392#_c_217_n N_VGND_M1006_d 0.0032429f $X=2.625 $Y=1.095 $X2=0
+ $Y2=0
cc_196 N_A_85_392#_c_229_n N_VGND_c_404_n 0.0200716f $X=0.69 $Y=0.91 $X2=0 $Y2=0
cc_197 N_A_85_392#_c_214_n N_VGND_c_404_n 0.0122781f $X=0.255 $Y=0.91 $X2=0
+ $Y2=0
cc_198 N_A_85_392#_c_215_n N_VGND_c_404_n 0.0117117f $X=0.855 $Y=0.515 $X2=0
+ $Y2=0
cc_199 N_A_85_392#_c_215_n N_VGND_c_405_n 0.0144369f $X=0.855 $Y=0.515 $X2=0
+ $Y2=0
cc_200 N_A_85_392#_c_215_n N_VGND_c_406_n 0.0117351f $X=0.855 $Y=0.515 $X2=0
+ $Y2=0
cc_201 N_A_85_392#_c_241_n N_VGND_c_406_n 0.0378283f $X=1.86 $Y=0.91 $X2=0 $Y2=0
cc_202 N_A_85_392#_c_216_n N_VGND_c_406_n 0.0117351f $X=2.025 $Y=0.515 $X2=0
+ $Y2=0
cc_203 N_A_85_392#_M1002_g N_VGND_c_407_n 0.0054327f $X=2.915 $Y=0.74 $X2=0
+ $Y2=0
cc_204 N_A_85_392#_c_216_n N_VGND_c_407_n 0.0186098f $X=2.025 $Y=0.515 $X2=0
+ $Y2=0
cc_205 N_A_85_392#_c_217_n N_VGND_c_407_n 0.0332559f $X=2.625 $Y=1.095 $X2=0
+ $Y2=0
cc_206 N_A_85_392#_c_219_n N_VGND_c_407_n 3.32959e-19 $X=3.25 $Y=1.532 $X2=0
+ $Y2=0
cc_207 N_A_85_392#_M1002_g N_VGND_c_409_n 4.98425e-19 $X=2.915 $Y=0.74 $X2=0
+ $Y2=0
cc_208 N_A_85_392#_M1008_g N_VGND_c_409_n 0.0107998f $X=3.345 $Y=0.74 $X2=0
+ $Y2=0
cc_209 N_A_85_392#_c_216_n N_VGND_c_410_n 0.0144922f $X=2.025 $Y=0.515 $X2=0
+ $Y2=0
cc_210 N_A_85_392#_M1002_g N_VGND_c_411_n 0.00434272f $X=2.915 $Y=0.74 $X2=0
+ $Y2=0
cc_211 N_A_85_392#_M1008_g N_VGND_c_411_n 0.00383152f $X=3.345 $Y=0.74 $X2=0
+ $Y2=0
cc_212 N_A_85_392#_M1002_g N_VGND_c_414_n 0.00822005f $X=2.915 $Y=0.74 $X2=0
+ $Y2=0
cc_213 N_A_85_392#_M1008_g N_VGND_c_414_n 0.0075754f $X=3.345 $Y=0.74 $X2=0
+ $Y2=0
cc_214 N_A_85_392#_c_229_n N_VGND_c_414_n 0.00625727f $X=0.69 $Y=0.91 $X2=0
+ $Y2=0
cc_215 N_A_85_392#_c_214_n N_VGND_c_414_n 0.00175584f $X=0.255 $Y=0.91 $X2=0
+ $Y2=0
cc_216 N_A_85_392#_c_215_n N_VGND_c_414_n 0.0118609f $X=0.855 $Y=0.515 $X2=0
+ $Y2=0
cc_217 N_A_85_392#_c_241_n N_VGND_c_414_n 0.0124314f $X=1.86 $Y=0.91 $X2=0 $Y2=0
cc_218 N_A_85_392#_c_216_n N_VGND_c_414_n 0.0118826f $X=2.025 $Y=0.515 $X2=0
+ $Y2=0
cc_219 N_VPWR_c_325_n N_X_c_366_n 0.0386506f $X=2.525 $Y=2.115 $X2=0 $Y2=0
cc_220 N_VPWR_c_327_n N_X_c_366_n 0.0323093f $X=3.525 $Y=2.225 $X2=0 $Y2=0
cc_221 N_VPWR_c_330_n N_X_c_366_n 0.014552f $X=3.36 $Y=3.33 $X2=0 $Y2=0
cc_222 N_VPWR_c_324_n N_X_c_366_n 0.0119791f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_223 N_VPWR_M1010_s N_X_c_367_n 0.0043188f $X=3.325 $Y=1.84 $X2=0 $Y2=0
cc_224 N_VPWR_c_327_n N_X_c_367_n 0.0268036f $X=3.525 $Y=2.225 $X2=0 $Y2=0
cc_225 N_X_c_363_n N_VGND_M1008_s 0.00347278f $X=3.485 $Y=1.045 $X2=0 $Y2=0
cc_226 N_X_c_362_n N_VGND_c_407_n 0.0179049f $X=3.13 $Y=0.515 $X2=0 $Y2=0
cc_227 N_X_c_362_n N_VGND_c_409_n 0.0159605f $X=3.13 $Y=0.515 $X2=0 $Y2=0
cc_228 N_X_c_363_n N_VGND_c_409_n 0.0217412f $X=3.485 $Y=1.045 $X2=0 $Y2=0
cc_229 N_X_c_362_n N_VGND_c_411_n 0.0109942f $X=3.13 $Y=0.515 $X2=0 $Y2=0
cc_230 N_X_c_362_n N_VGND_c_414_n 0.00904371f $X=3.13 $Y=0.515 $X2=0 $Y2=0
