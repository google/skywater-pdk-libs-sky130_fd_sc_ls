* File: sky130_fd_sc_ls__or4_1.pxi.spice
* Created: Fri Aug 28 13:59:33 2020
* 
x_PM_SKY130_FD_SC_LS__OR4_1%D N_D_M1002_g N_D_c_59_n N_D_M1000_g D N_D_c_60_n
+ PM_SKY130_FD_SC_LS__OR4_1%D
x_PM_SKY130_FD_SC_LS__OR4_1%C N_C_M1001_g N_C_c_85_n N_C_M1007_g C
+ PM_SKY130_FD_SC_LS__OR4_1%C
x_PM_SKY130_FD_SC_LS__OR4_1%B N_B_c_113_n N_B_M1009_g N_B_M1004_g B
+ PM_SKY130_FD_SC_LS__OR4_1%B
x_PM_SKY130_FD_SC_LS__OR4_1%A N_A_c_142_n N_A_M1005_g N_A_M1003_g A N_A_c_144_n
+ PM_SKY130_FD_SC_LS__OR4_1%A
x_PM_SKY130_FD_SC_LS__OR4_1%A_44_392# N_A_44_392#_M1002_d N_A_44_392#_M1004_d
+ N_A_44_392#_M1000_s N_A_44_392#_M1006_g N_A_44_392#_c_178_n
+ N_A_44_392#_M1008_g N_A_44_392#_c_188_n N_A_44_392#_c_189_n
+ N_A_44_392#_c_190_n N_A_44_392#_c_179_n N_A_44_392#_c_180_n
+ N_A_44_392#_c_181_n N_A_44_392#_c_182_n N_A_44_392#_c_183_n
+ N_A_44_392#_c_184_n N_A_44_392#_c_185_n N_A_44_392#_c_186_n
+ PM_SKY130_FD_SC_LS__OR4_1%A_44_392#
x_PM_SKY130_FD_SC_LS__OR4_1%VPWR N_VPWR_M1005_d N_VPWR_c_276_n VPWR
+ N_VPWR_c_277_n N_VPWR_c_278_n N_VPWR_c_275_n N_VPWR_c_280_n
+ PM_SKY130_FD_SC_LS__OR4_1%VPWR
x_PM_SKY130_FD_SC_LS__OR4_1%X N_X_M1006_d N_X_M1008_d N_X_c_302_n N_X_c_303_n X
+ X X X N_X_c_304_n PM_SKY130_FD_SC_LS__OR4_1%X
x_PM_SKY130_FD_SC_LS__OR4_1%VGND N_VGND_M1002_s N_VGND_M1001_d N_VGND_M1003_d
+ N_VGND_c_325_n N_VGND_c_326_n N_VGND_c_327_n N_VGND_c_328_n N_VGND_c_329_n
+ VGND N_VGND_c_330_n N_VGND_c_331_n N_VGND_c_332_n N_VGND_c_333_n
+ N_VGND_c_334_n PM_SKY130_FD_SC_LS__OR4_1%VGND
cc_1 VNB N_D_M1002_g 0.0360698f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.835
cc_2 VNB N_D_c_59_n 0.0241911f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.885
cc_3 VNB N_D_c_60_n 0.0135797f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.585
cc_4 VNB N_C_M1001_g 0.0312133f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.835
cc_5 VNB N_C_c_85_n 0.0188573f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.885
cc_6 VNB C 0.00378948f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_7 VNB N_B_c_113_n 0.0220247f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.42
cc_8 VNB N_B_M1004_g 0.0332829f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=2.46
cc_9 VNB B 0.00187616f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_10 VNB N_A_c_142_n 0.0252463f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.42
cc_11 VNB N_A_M1003_g 0.0262449f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=2.46
cc_12 VNB N_A_c_144_n 0.00426371f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.585
cc_13 VNB N_A_44_392#_M1006_g 0.0287893f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.585
cc_14 VNB N_A_44_392#_c_178_n 0.0356542f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_44_392#_c_179_n 0.00325236f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_44_392#_c_180_n 0.0116367f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_44_392#_c_181_n 0.0106209f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_44_392#_c_182_n 0.00430793f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_44_392#_c_183_n 0.00595784f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_44_392#_c_184_n 0.0103286f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_44_392#_c_185_n 3.93303e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_44_392#_c_186_n 0.00857761f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VPWR_c_275_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_X_c_302_n 0.0279492f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_X_c_303_n 0.012405f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.6
cc_26 VNB N_X_c_304_n 0.0247746f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_325_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0.492 $Y2=1.585
cc_28 VNB N_VGND_c_326_n 0.0551753f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.585
cc_29 VNB N_VGND_c_327_n 0.0198125f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_328_n 0.0288416f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_329_n 0.0135712f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_330_n 0.0252222f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_331_n 0.0179969f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_332_n 0.222079f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_333_n 0.00913651f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_334_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VPB N_D_c_59_n 0.0446231f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.885
cc_38 VPB N_D_c_60_n 0.0110488f $X=-0.19 $Y=1.66 $X2=0.485 $Y2=1.585
cc_39 VPB N_C_c_85_n 0.0351009f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.885
cc_40 VPB C 0.00346319f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_41 VPB N_B_c_113_n 0.0379428f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=1.42
cc_42 VPB B 0.00159046f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_43 VPB N_A_c_142_n 0.0363925f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=1.42
cc_44 VPB N_A_c_144_n 0.00303074f $X=-0.19 $Y=1.66 $X2=0.485 $Y2=1.585
cc_45 VPB N_A_44_392#_c_178_n 0.0304508f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_A_44_392#_c_188_n 0.00942361f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB N_A_44_392#_c_189_n 0.035396f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 VPB N_A_44_392#_c_190_n 0.0307924f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 VPB N_A_44_392#_c_185_n 0.0029843f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_276_n 0.00701163f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=2.46
cc_51 VPB N_VPWR_c_277_n 0.0678403f $X=-0.19 $Y=1.66 $X2=0.492 $Y2=1.585
cc_52 VPB N_VPWR_c_278_n 0.0245279f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_275_n 0.106073f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_280_n 0.0076819f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB X 0.0146542f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB X 0.042262f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_X_c_304_n 0.00758423f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 N_D_M1002_g N_C_M1001_g 0.027997f $X=0.565 $Y=0.835 $X2=0 $Y2=0
cc_59 N_D_c_59_n N_C_c_85_n 0.0809994f $X=0.59 $Y=1.885 $X2=0 $Y2=0
cc_60 N_D_c_60_n N_C_c_85_n 4.57439e-19 $X=0.485 $Y=1.585 $X2=0 $Y2=0
cc_61 N_D_c_59_n C 5.19757e-19 $X=0.59 $Y=1.885 $X2=0 $Y2=0
cc_62 N_D_c_60_n C 0.0195595f $X=0.485 $Y=1.585 $X2=0 $Y2=0
cc_63 N_D_c_59_n N_A_44_392#_c_188_n 0.00240296f $X=0.59 $Y=1.885 $X2=0 $Y2=0
cc_64 N_D_c_60_n N_A_44_392#_c_188_n 0.029179f $X=0.485 $Y=1.585 $X2=0 $Y2=0
cc_65 N_D_c_59_n N_A_44_392#_c_189_n 0.0154541f $X=0.59 $Y=1.885 $X2=0 $Y2=0
cc_66 N_D_c_59_n N_A_44_392#_c_190_n 0.0121603f $X=0.59 $Y=1.885 $X2=0 $Y2=0
cc_67 N_D_c_60_n N_A_44_392#_c_190_n 0.00859598f $X=0.485 $Y=1.585 $X2=0 $Y2=0
cc_68 N_D_M1002_g N_A_44_392#_c_179_n 0.0065178f $X=0.565 $Y=0.835 $X2=0 $Y2=0
cc_69 N_D_M1002_g N_A_44_392#_c_181_n 0.00581878f $X=0.565 $Y=0.835 $X2=0 $Y2=0
cc_70 N_D_c_59_n N_A_44_392#_c_181_n 7.3211e-19 $X=0.59 $Y=1.885 $X2=0 $Y2=0
cc_71 N_D_c_60_n N_A_44_392#_c_181_n 0.00216782f $X=0.485 $Y=1.585 $X2=0 $Y2=0
cc_72 N_D_c_59_n N_VPWR_c_277_n 0.00445602f $X=0.59 $Y=1.885 $X2=0 $Y2=0
cc_73 N_D_c_59_n N_VPWR_c_275_n 0.00861901f $X=0.59 $Y=1.885 $X2=0 $Y2=0
cc_74 N_D_M1002_g N_VGND_c_326_n 0.00867578f $X=0.565 $Y=0.835 $X2=0 $Y2=0
cc_75 N_D_c_59_n N_VGND_c_326_n 0.0026975f $X=0.59 $Y=1.885 $X2=0 $Y2=0
cc_76 N_D_c_60_n N_VGND_c_326_n 0.0190298f $X=0.485 $Y=1.585 $X2=0 $Y2=0
cc_77 N_D_M1002_g N_VGND_c_327_n 0.0043356f $X=0.565 $Y=0.835 $X2=0 $Y2=0
cc_78 N_D_M1002_g N_VGND_c_332_n 0.00487769f $X=0.565 $Y=0.835 $X2=0 $Y2=0
cc_79 N_C_c_85_n N_B_c_113_n 0.0630662f $X=1.01 $Y=1.885 $X2=-0.19 $Y2=-0.245
cc_80 C N_B_c_113_n 0.00223685f $X=1.115 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_81 N_C_M1001_g N_B_M1004_g 0.0175401f $X=0.995 $Y=0.835 $X2=0 $Y2=0
cc_82 N_C_c_85_n B 4.12227e-19 $X=1.01 $Y=1.885 $X2=0 $Y2=0
cc_83 C B 0.0259384f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_84 N_C_c_85_n N_A_44_392#_c_189_n 0.00413008f $X=1.01 $Y=1.885 $X2=0 $Y2=0
cc_85 N_C_c_85_n N_A_44_392#_c_190_n 0.0174443f $X=1.01 $Y=1.885 $X2=0 $Y2=0
cc_86 C N_A_44_392#_c_190_n 0.0286231f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_87 N_C_M1001_g N_A_44_392#_c_179_n 0.0121196f $X=0.995 $Y=0.835 $X2=0 $Y2=0
cc_88 N_C_M1001_g N_A_44_392#_c_180_n 0.0124559f $X=0.995 $Y=0.835 $X2=0 $Y2=0
cc_89 N_C_c_85_n N_A_44_392#_c_180_n 0.00392723f $X=1.01 $Y=1.885 $X2=0 $Y2=0
cc_90 C N_A_44_392#_c_180_n 0.0201443f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_91 N_C_M1001_g N_A_44_392#_c_181_n 0.00256575f $X=0.995 $Y=0.835 $X2=0 $Y2=0
cc_92 C N_A_44_392#_c_181_n 0.00151542f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_93 N_C_c_85_n N_VPWR_c_277_n 0.00461464f $X=1.01 $Y=1.885 $X2=0 $Y2=0
cc_94 N_C_c_85_n N_VPWR_c_275_n 0.00910574f $X=1.01 $Y=1.885 $X2=0 $Y2=0
cc_95 N_C_M1001_g N_VGND_c_327_n 0.0043356f $X=0.995 $Y=0.835 $X2=0 $Y2=0
cc_96 N_C_M1001_g N_VGND_c_328_n 0.00598528f $X=0.995 $Y=0.835 $X2=0 $Y2=0
cc_97 N_C_M1001_g N_VGND_c_332_n 0.00487769f $X=0.995 $Y=0.835 $X2=0 $Y2=0
cc_98 N_B_c_113_n N_A_c_142_n 0.0589024f $X=1.58 $Y=1.885 $X2=-0.19 $Y2=-0.245
cc_99 N_B_M1004_g N_A_c_142_n 0.00324793f $X=1.73 $Y=0.835 $X2=-0.19 $Y2=-0.245
cc_100 B N_A_c_142_n 5.27828e-19 $X=1.595 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_101 N_B_M1004_g N_A_M1003_g 0.0208052f $X=1.73 $Y=0.835 $X2=0 $Y2=0
cc_102 N_B_c_113_n N_A_c_144_n 0.00210886f $X=1.58 $Y=1.885 $X2=0 $Y2=0
cc_103 N_B_M1004_g N_A_c_144_n 0.00151003f $X=1.73 $Y=0.835 $X2=0 $Y2=0
cc_104 B N_A_c_144_n 0.0233207f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_105 N_B_c_113_n N_A_44_392#_c_190_n 0.0181897f $X=1.58 $Y=1.885 $X2=0 $Y2=0
cc_106 B N_A_44_392#_c_190_n 0.0249968f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_107 N_B_c_113_n N_A_44_392#_c_180_n 0.00115496f $X=1.58 $Y=1.885 $X2=0 $Y2=0
cc_108 N_B_M1004_g N_A_44_392#_c_180_n 0.0171248f $X=1.73 $Y=0.835 $X2=0 $Y2=0
cc_109 B N_A_44_392#_c_180_n 0.0186612f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_110 N_B_M1004_g N_A_44_392#_c_182_n 0.00299671f $X=1.73 $Y=0.835 $X2=0 $Y2=0
cc_111 N_B_c_113_n N_VPWR_c_276_n 0.00397122f $X=1.58 $Y=1.885 $X2=0 $Y2=0
cc_112 N_B_c_113_n N_VPWR_c_277_n 0.00461464f $X=1.58 $Y=1.885 $X2=0 $Y2=0
cc_113 N_B_c_113_n N_VPWR_c_275_n 0.00911823f $X=1.58 $Y=1.885 $X2=0 $Y2=0
cc_114 N_B_M1004_g N_VGND_c_328_n 0.00601282f $X=1.73 $Y=0.835 $X2=0 $Y2=0
cc_115 N_B_M1004_g N_VGND_c_330_n 0.00451272f $X=1.73 $Y=0.835 $X2=0 $Y2=0
cc_116 N_B_M1004_g N_VGND_c_332_n 0.00487769f $X=1.73 $Y=0.835 $X2=0 $Y2=0
cc_117 N_A_M1003_g N_A_44_392#_M1006_g 0.0183187f $X=2.32 $Y=0.835 $X2=0 $Y2=0
cc_118 N_A_c_142_n N_A_44_392#_c_178_n 0.0180457f $X=2.15 $Y=1.885 $X2=0 $Y2=0
cc_119 N_A_M1003_g N_A_44_392#_c_178_n 0.0204349f $X=2.32 $Y=0.835 $X2=0 $Y2=0
cc_120 N_A_c_144_n N_A_44_392#_c_178_n 3.1599e-19 $X=2.225 $Y=1.515 $X2=0 $Y2=0
cc_121 N_A_c_142_n N_A_44_392#_c_190_n 0.0162645f $X=2.15 $Y=1.885 $X2=0 $Y2=0
cc_122 N_A_c_144_n N_A_44_392#_c_190_n 0.0265723f $X=2.225 $Y=1.515 $X2=0 $Y2=0
cc_123 N_A_M1003_g N_A_44_392#_c_182_n 0.00299671f $X=2.32 $Y=0.835 $X2=0 $Y2=0
cc_124 N_A_c_142_n N_A_44_392#_c_183_n 3.81366e-19 $X=2.15 $Y=1.885 $X2=0 $Y2=0
cc_125 N_A_M1003_g N_A_44_392#_c_183_n 0.0158031f $X=2.32 $Y=0.835 $X2=0 $Y2=0
cc_126 N_A_c_144_n N_A_44_392#_c_183_n 0.0147621f $X=2.225 $Y=1.515 $X2=0 $Y2=0
cc_127 N_A_M1003_g N_A_44_392#_c_184_n 0.00539948f $X=2.32 $Y=0.835 $X2=0 $Y2=0
cc_128 N_A_c_144_n N_A_44_392#_c_184_n 0.0225675f $X=2.225 $Y=1.515 $X2=0 $Y2=0
cc_129 N_A_c_142_n N_A_44_392#_c_185_n 0.00385701f $X=2.15 $Y=1.885 $X2=0 $Y2=0
cc_130 N_A_c_144_n N_A_44_392#_c_185_n 0.0116888f $X=2.225 $Y=1.515 $X2=0 $Y2=0
cc_131 N_A_c_142_n N_A_44_392#_c_186_n 0.00100681f $X=2.15 $Y=1.885 $X2=0 $Y2=0
cc_132 N_A_c_144_n N_A_44_392#_c_186_n 0.0124267f $X=2.225 $Y=1.515 $X2=0 $Y2=0
cc_133 N_A_c_142_n N_VPWR_c_276_n 0.024208f $X=2.15 $Y=1.885 $X2=0 $Y2=0
cc_134 N_A_c_142_n N_VPWR_c_277_n 0.00229331f $X=2.15 $Y=1.885 $X2=0 $Y2=0
cc_135 N_A_c_142_n N_VPWR_c_275_n 0.00458846f $X=2.15 $Y=1.885 $X2=0 $Y2=0
cc_136 N_A_c_142_n X 8.41746e-19 $X=2.15 $Y=1.885 $X2=0 $Y2=0
cc_137 N_A_M1003_g N_VGND_c_329_n 0.00475377f $X=2.32 $Y=0.835 $X2=0 $Y2=0
cc_138 N_A_M1003_g N_VGND_c_330_n 0.00451272f $X=2.32 $Y=0.835 $X2=0 $Y2=0
cc_139 N_A_M1003_g N_VGND_c_332_n 0.00487769f $X=2.32 $Y=0.835 $X2=0 $Y2=0
cc_140 N_A_44_392#_c_190_n A_133_392# 0.00595227f $X=2.56 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_141 N_A_44_392#_c_190_n A_217_392# 0.0122036f $X=2.56 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_142 N_A_44_392#_c_190_n A_331_392# 0.0122036f $X=2.56 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_143 N_A_44_392#_c_190_n N_VPWR_M1005_d 0.0146043f $X=2.56 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_144 N_A_44_392#_c_185_n N_VPWR_M1005_d 0.00231635f $X=2.645 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_145 N_A_44_392#_c_178_n N_VPWR_c_276_n 0.00988355f $X=2.84 $Y=1.765 $X2=0
+ $Y2=0
cc_146 N_A_44_392#_c_190_n N_VPWR_c_276_n 0.028176f $X=2.56 $Y=2.035 $X2=0 $Y2=0
cc_147 N_A_44_392#_c_189_n N_VPWR_c_277_n 0.0145938f $X=0.365 $Y=2.815 $X2=0
+ $Y2=0
cc_148 N_A_44_392#_c_178_n N_VPWR_c_278_n 0.00445602f $X=2.84 $Y=1.765 $X2=0
+ $Y2=0
cc_149 N_A_44_392#_c_178_n N_VPWR_c_275_n 0.0086373f $X=2.84 $Y=1.765 $X2=0
+ $Y2=0
cc_150 N_A_44_392#_c_189_n N_VPWR_c_275_n 0.0120466f $X=0.365 $Y=2.815 $X2=0
+ $Y2=0
cc_151 N_A_44_392#_M1006_g N_X_c_302_n 0.00205928f $X=2.83 $Y=0.74 $X2=0 $Y2=0
cc_152 N_A_44_392#_c_184_n N_X_c_303_n 0.00135284f $X=2.645 $Y=1.63 $X2=0 $Y2=0
cc_153 N_A_44_392#_c_178_n X 0.00290257f $X=2.84 $Y=1.765 $X2=0 $Y2=0
cc_154 N_A_44_392#_c_184_n X 0.00258446f $X=2.645 $Y=1.63 $X2=0 $Y2=0
cc_155 N_A_44_392#_c_185_n X 0.00568912f $X=2.645 $Y=1.95 $X2=0 $Y2=0
cc_156 N_A_44_392#_c_178_n X 0.0158482f $X=2.84 $Y=1.765 $X2=0 $Y2=0
cc_157 N_A_44_392#_M1006_g N_X_c_304_n 0.00244983f $X=2.83 $Y=0.74 $X2=0 $Y2=0
cc_158 N_A_44_392#_c_178_n N_X_c_304_n 0.00537395f $X=2.84 $Y=1.765 $X2=0 $Y2=0
cc_159 N_A_44_392#_c_184_n N_X_c_304_n 0.0303927f $X=2.645 $Y=1.63 $X2=0 $Y2=0
cc_160 N_A_44_392#_c_185_n N_X_c_304_n 0.00605514f $X=2.645 $Y=1.95 $X2=0 $Y2=0
cc_161 N_A_44_392#_c_180_n N_VGND_M1001_d 0.00623975f $X=1.86 $Y=1.095 $X2=0
+ $Y2=0
cc_162 N_A_44_392#_c_183_n N_VGND_M1003_d 0.00113743f $X=2.56 $Y=1.095 $X2=0
+ $Y2=0
cc_163 N_A_44_392#_c_184_n N_VGND_M1003_d 0.00214042f $X=2.645 $Y=1.63 $X2=0
+ $Y2=0
cc_164 N_A_44_392#_c_179_n N_VGND_c_326_n 0.0183885f $X=0.78 $Y=0.835 $X2=0
+ $Y2=0
cc_165 N_A_44_392#_c_181_n N_VGND_c_326_n 0.00584871f $X=0.945 $Y=1.095 $X2=0
+ $Y2=0
cc_166 N_A_44_392#_c_179_n N_VGND_c_327_n 0.00805448f $X=0.78 $Y=0.835 $X2=0
+ $Y2=0
cc_167 N_A_44_392#_c_179_n N_VGND_c_328_n 0.0115546f $X=0.78 $Y=0.835 $X2=0
+ $Y2=0
cc_168 N_A_44_392#_c_180_n N_VGND_c_328_n 0.0383199f $X=1.86 $Y=1.095 $X2=0
+ $Y2=0
cc_169 N_A_44_392#_c_182_n N_VGND_c_328_n 0.00120817f $X=2.025 $Y=0.835 $X2=0
+ $Y2=0
cc_170 N_A_44_392#_M1006_g N_VGND_c_329_n 0.0155432f $X=2.83 $Y=0.74 $X2=0 $Y2=0
cc_171 N_A_44_392#_c_178_n N_VGND_c_329_n 4.70665e-19 $X=2.84 $Y=1.765 $X2=0
+ $Y2=0
cc_172 N_A_44_392#_c_182_n N_VGND_c_329_n 0.00117493f $X=2.025 $Y=0.835 $X2=0
+ $Y2=0
cc_173 N_A_44_392#_c_183_n N_VGND_c_329_n 0.00875025f $X=2.56 $Y=1.095 $X2=0
+ $Y2=0
cc_174 N_A_44_392#_c_184_n N_VGND_c_329_n 0.0136978f $X=2.645 $Y=1.63 $X2=0
+ $Y2=0
cc_175 N_A_44_392#_c_182_n N_VGND_c_330_n 0.00817062f $X=2.025 $Y=0.835 $X2=0
+ $Y2=0
cc_176 N_A_44_392#_M1006_g N_VGND_c_331_n 0.00383152f $X=2.83 $Y=0.74 $X2=0
+ $Y2=0
cc_177 N_A_44_392#_M1006_g N_VGND_c_332_n 0.00761312f $X=2.83 $Y=0.74 $X2=0
+ $Y2=0
cc_178 N_A_44_392#_c_179_n N_VGND_c_332_n 0.0105848f $X=0.78 $Y=0.835 $X2=0
+ $Y2=0
cc_179 N_A_44_392#_c_182_n N_VGND_c_332_n 0.010638f $X=2.025 $Y=0.835 $X2=0
+ $Y2=0
cc_180 N_VPWR_c_276_n X 0.0327496f $X=2.375 $Y=2.455 $X2=0 $Y2=0
cc_181 N_VPWR_c_278_n X 0.0166018f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_182 N_VPWR_c_275_n X 0.0137086f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_183 N_X_c_302_n N_VGND_c_329_n 0.0183161f $X=3.045 $Y=0.515 $X2=0 $Y2=0
cc_184 N_X_c_302_n N_VGND_c_331_n 0.0139663f $X=3.045 $Y=0.515 $X2=0 $Y2=0
cc_185 N_X_c_302_n N_VGND_c_332_n 0.0115601f $X=3.045 $Y=0.515 $X2=0 $Y2=0
