* File: sky130_fd_sc_ls__sdfrtp_4.spice
* Created: Fri Aug 28 14:03:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__sdfrtp_4.pex.spice"
.subckt sky130_fd_sc_ls__sdfrtp_4  VNB VPB SCE D SCD CLK RESET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* RESET_B	RESET_B
* CLK	CLK
* SCD	SCD
* D	D
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1036 N_VGND_M1036_d N_SCE_M1036_g N_A_27_74#_M1036_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.1197 PD=1.41 PS=1.41 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1005 noxref_25 N_A_27_74#_M1005_g N_noxref_24_M1005_s VNB NSHORT L=0.15 W=0.42
+ AD=0.07665 AS=0.1197 PD=0.785 PS=1.41 NRD=36.42 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.3 A=0.063 P=1.14 MULT=1
MM1006 N_A_415_81#_M1006_d N_D_M1006_g noxref_25 VNB NSHORT L=0.15 W=0.42
+ AD=0.13335 AS=0.07665 PD=1.055 PS=0.785 NRD=81.42 NRS=36.42 M=1 R=2.8
+ SA=75000.7 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1037 noxref_26 N_SCE_M1037_g N_A_415_81#_M1006_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.13335 PD=0.63 PS=1.055 NRD=14.28 NRS=19.992 M=1 R=2.8
+ SA=75001.5 SB=75001 A=0.063 P=1.14 MULT=1
MM1040 N_noxref_24_M1040_d N_SCD_M1040_g noxref_26 VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.9
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1012 N_VGND_M1012_d N_RESET_B_M1012_g N_noxref_24_M1040_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75002.3
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1010 N_VGND_M1010_d N_CLK_M1010_g N_A_837_98#_M1010_s VNB NSHORT L=0.15 W=0.74
+ AD=0.161125 AS=0.242325 PD=1.245 PS=2.38 NRD=10.536 NRS=10.536 M=1 R=4.93333
+ SA=75000.2 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1013 N_A_1034_392#_M1013_d N_A_837_98#_M1013_g N_VGND_M1010_d VNB NSHORT
+ L=0.15 W=0.74 AD=0.1961 AS=0.161125 PD=2.01 PS=1.245 NRD=0 NRS=10.536 M=1
+ R=4.93333 SA=75000.8 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1032 N_A_1236_138#_M1032_d N_A_837_98#_M1032_g N_A_415_81#_M1032_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75003.2 A=0.063 P=1.14 MULT=1
MM1041 A_1322_138# N_A_1034_392#_M1041_g N_A_1236_138#_M1032_d VNB NSHORT L=0.15
+ W=0.42 AD=0.04725 AS=0.0588 PD=0.645 PS=0.7 NRD=16.428 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75002.8 A=0.063 P=1.14 MULT=1
MM1044 A_1397_138# N_A_1367_112#_M1044_g A_1322_138# VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.04725 PD=0.66 PS=0.645 NRD=18.564 NRS=16.428 M=1 R=2.8 SA=75001
+ SB=75002.4 A=0.063 P=1.14 MULT=1
MM1024 N_VGND_M1024_d N_RESET_B_M1024_g A_1397_138# VNB NSHORT L=0.15 W=0.42
+ AD=0.20551 AS=0.0504 PD=1.19845 PS=0.66 NRD=124.08 NRS=18.564 M=1 R=2.8
+ SA=75001.4 SB=75002 A=0.063 P=1.14 MULT=1
MM1019 N_A_1367_112#_M1019_d N_A_1236_138#_M1019_g N_VGND_M1024_d VNB NSHORT
+ L=0.15 W=0.74 AD=0.124942 AS=0.36209 PD=1.14217 PS=2.11155 NRD=0 NRS=70.428
+ M=1 R=4.93333 SA=75001.5 SB=75002 A=0.111 P=1.78 MULT=1
MM1003 N_A_1745_74#_M1003_d N_A_1034_392#_M1003_g N_A_1367_112#_M1019_d VNB
+ NSHORT L=0.15 W=0.64 AD=0.261434 AS=0.108058 PD=1.85962 PS=0.987826
+ NRD=101.244 NRS=0 M=1 R=4.26667 SA=75001.9 SB=75001.8 A=0.096 P=1.58 MULT=1
MM1027 A_1955_74# N_A_837_98#_M1027_g N_A_1745_74#_M1003_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.171566 PD=0.66 PS=1.22038 NRD=18.564 NRS=22.848 M=1
+ R=2.8 SA=75002.5 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1021 N_VGND_M1021_d N_A_2003_48#_M1021_g A_1955_74# VNB NSHORT L=0.15 W=0.42
+ AD=0.0819 AS=0.0504 PD=0.81 PS=0.66 NRD=15.708 NRS=18.564 M=1 R=2.8 SA=75002.9
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1038 A_2141_74# N_RESET_B_M1038_g N_VGND_M1021_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0819 PD=0.63 PS=0.81 NRD=14.28 NRS=15.708 M=1 R=2.8 SA=75003.4
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1020 N_A_2003_48#_M1020_d N_A_1745_74#_M1020_g A_2141_74# VNB NSHORT L=0.15
+ W=0.42 AD=0.1512 AS=0.0441 PD=1.56 PS=0.63 NRD=9.996 NRS=14.28 M=1 R=2.8
+ SA=75003.8 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1011 N_VGND_M1011_d N_A_1745_74#_M1011_g N_A_2339_74#_M1011_s VNB NSHORT
+ L=0.15 W=0.74 AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75002.5 A=0.111 P=1.78 MULT=1
MM1007 N_VGND_M1011_d N_A_2339_74#_M1007_g N_Q_M1007_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75002.1 A=0.111 P=1.78 MULT=1
MM1016 N_VGND_M1016_d N_A_2339_74#_M1016_g N_Q_M1007_s VNB NSHORT L=0.15 W=0.74
+ AD=0.3293 AS=0.1036 PD=1.63 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75001.7 A=0.111 P=1.78 MULT=1
MM1022 N_VGND_M1016_d N_A_2339_74#_M1022_g N_Q_M1022_s VNB NSHORT L=0.15 W=0.74
+ AD=0.3293 AS=0.1036 PD=1.63 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.1
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1028 N_VGND_M1028_d N_A_2339_74#_M1028_g N_Q_M1022_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.5
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1023 N_VPWR_M1023_d N_SCE_M1023_g N_A_27_74#_M1023_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.3104 AS=0.1888 PD=1.61 PS=1.87 NRD=18.4589 NRS=3.0732 M=1 R=4.26667
+ SA=75000.2 SB=75003.3 A=0.096 P=1.58 MULT=1
MM1026 A_340_464# N_SCE_M1026_g N_VPWR_M1023_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0864 AS=0.3104 PD=0.91 PS=1.61 NRD=24.625 NRS=3.0732 M=1 R=4.26667
+ SA=75001.3 SB=75002.2 A=0.096 P=1.58 MULT=1
MM1002 N_A_415_81#_M1002_d N_D_M1002_g A_340_464# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.096 AS=0.0864 PD=0.94 PS=0.91 NRD=3.0732 NRS=24.625 M=1 R=4.26667
+ SA=75001.8 SB=75001.8 A=0.096 P=1.58 MULT=1
MM1014 A_514_464# N_A_27_74#_M1014_g N_A_415_81#_M1002_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1248 AS=0.096 PD=1.03 PS=0.94 NRD=43.0839 NRS=3.0732 M=1 R=4.26667
+ SA=75002.2 SB=75001.3 A=0.096 P=1.58 MULT=1
MM1029 N_VPWR_M1029_d N_SCD_M1029_g A_514_464# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1344 AS=0.1248 PD=1.06 PS=1.03 NRD=3.0732 NRS=43.0839 M=1 R=4.26667
+ SA=75002.8 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1045 N_A_415_81#_M1045_d N_RESET_B_M1045_g N_VPWR_M1029_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1888 AS=0.1344 PD=1.87 PS=1.06 NRD=3.0732 NRS=40.0107 M=1
+ R=4.26667 SA=75003.3 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1030 N_VPWR_M1030_d N_CLK_M1030_g N_A_837_98#_M1030_s VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.295 PD=1.3 PS=2.59 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75000.2
+ SB=75000.7 A=0.15 P=2.3 MULT=1
MM1034 N_A_1034_392#_M1034_d N_A_837_98#_M1034_g N_VPWR_M1030_d VPB PHIGHVT
+ L=0.15 W=1 AD=0.295 AS=0.15 PD=2.59 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75000.7 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1000 N_A_1236_138#_M1000_d N_A_1034_392#_M1000_g N_A_415_81#_M1000_s VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.0735 AS=0.1239 PD=0.77 PS=1.43 NRD=28.1316
+ NRS=4.6886 M=1 R=2.8 SA=75000.2 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1008 A_1342_463# N_A_837_98#_M1008_g N_A_1236_138#_M1000_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0504 AS=0.0735 PD=0.66 PS=0.77 NRD=30.4759 NRS=4.6886 M=1 R=2.8
+ SA=75000.7 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1009 N_VPWR_M1009_d N_A_1367_112#_M1009_g A_1342_463# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.139325 AS=0.0504 PD=1.145 PS=0.66 NRD=129.784 NRS=30.4759 M=1
+ R=2.8 SA=75001.1 SB=75000.9 A=0.063 P=1.14 MULT=1
MM1001 N_A_1236_138#_M1001_d N_RESET_B_M1001_g N_VPWR_M1009_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1239 AS=0.139325 PD=1.43 PS=1.145 NRD=4.6886 NRS=129.784 M=1 R=2.8
+ SA=75001.7 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1031 N_A_1367_112#_M1031_d N_A_1236_138#_M1031_g N_VPWR_M1031_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.15 AS=0.295 PD=1.3 PS=2.59 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75001.5 A=0.15 P=2.3 MULT=1
MM1042 N_A_1745_74#_M1042_d N_A_837_98#_M1042_g N_A_1367_112#_M1031_d VPB
+ PHIGHVT L=0.15 W=1 AD=0.301602 AS=0.15 PD=2.51408 PS=1.3 NRD=36.445 NRS=1.9503
+ M=1 R=6.66667 SA=75000.7 SB=75001.1 A=0.15 P=2.3 MULT=1
MM1018 A_1982_508# N_A_1034_392#_M1018_g N_A_1745_74#_M1042_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0567 AS=0.126673 PD=0.69 PS=1.05592 NRD=37.5088 NRS=46.886 M=1
+ R=2.8 SA=75000.9 SB=75002.8 A=0.063 P=1.14 MULT=1
MM1043 N_VPWR_M1043_d N_A_2003_48#_M1043_g A_1982_508# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.11235 AS=0.0567 PD=0.955 PS=0.69 NRD=75.0373 NRS=37.5088 M=1 R=2.8
+ SA=75001.3 SB=75002.4 A=0.063 P=1.14 MULT=1
MM1015 N_A_2003_48#_M1015_d N_RESET_B_M1015_g N_VPWR_M1043_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.08085 AS=0.11235 PD=0.805 PS=0.955 NRD=4.6886 NRS=44.5417 M=1
+ R=2.8 SA=75002 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1035 N_VPWR_M1035_d N_A_1745_74#_M1035_g N_A_2003_48#_M1015_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.1197 AS=0.08085 PD=1.02333 PS=0.805 NRD=60.9715 NRS=44.5417
+ M=1 R=2.8 SA=75002.5 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1033 N_A_2339_74#_M1033_d N_A_1745_74#_M1033_g N_VPWR_M1035_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.126 AS=0.2394 PD=1.14 PS=2.04667 NRD=2.3443 NRS=2.3443 M=1
+ R=5.6 SA=75000.8 SB=75002.6 A=0.126 P=1.98 MULT=1
MM1046 N_A_2339_74#_M1033_d N_A_1745_74#_M1046_g N_VPWR_M1046_s VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.126 AS=0.174 PD=1.14 PS=1.29 NRD=2.3443 NRS=22.261 M=1
+ R=5.6 SA=75001.2 SB=75002.1 A=0.126 P=1.98 MULT=1
MM1004 N_VPWR_M1046_s N_A_2339_74#_M1004_g N_Q_M1004_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.232 AS=0.168 PD=1.72 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.4 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1017 N_VPWR_M1017_d N_A_2339_74#_M1017_g N_Q_M1004_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.8 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1025 N_VPWR_M1017_d N_A_2339_74#_M1025_g N_Q_M1025_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.3 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1039 N_VPWR_M1039_d N_A_2339_74#_M1039_g N_Q_M1025_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.7 SB=75000.2 A=0.168 P=2.54 MULT=1
DX47_noxref VNB VPB NWDIODE A=28.3212 P=34.69
c_156 VNB 0 1.59743e-19 $X=0 $Y=0
c_2243 A_1342_463# 0 9.53373e-20 $X=6.71 $Y=2.315
c_2491 A_1397_138# 0 1.57165e-19 $X=6.985 $Y=0.69
*
.include "sky130_fd_sc_ls__sdfrtp_4.pxi.spice"
*
.ends
*
*
