* File: sky130_fd_sc_ls__nor3_2.pxi.spice
* Created: Fri Aug 28 13:38:28 2020
* 
x_PM_SKY130_FD_SC_LS__NOR3_2%C N_C_c_57_n N_C_M1006_g N_C_c_60_n N_C_M1003_g
+ N_C_c_61_n N_C_M1004_g C N_C_c_59_n PM_SKY130_FD_SC_LS__NOR3_2%C
x_PM_SKY130_FD_SC_LS__NOR3_2%B N_B_c_97_n N_B_M1002_g N_B_c_98_n N_B_M1008_g
+ N_B_c_99_n N_B_M1005_g N_B_c_100_n N_B_c_101_n B PM_SKY130_FD_SC_LS__NOR3_2%B
x_PM_SKY130_FD_SC_LS__NOR3_2%A N_A_c_160_n N_A_c_171_n N_A_M1000_g N_A_c_161_n
+ N_A_M1007_g N_A_c_162_n N_A_c_163_n N_A_c_173_n N_A_M1001_g N_A_c_164_n
+ N_A_c_165_n N_A_c_166_n N_A_c_167_n A N_A_c_169_n PM_SKY130_FD_SC_LS__NOR3_2%A
x_PM_SKY130_FD_SC_LS__NOR3_2%A_27_368# N_A_27_368#_M1003_d N_A_27_368#_M1004_d
+ N_A_27_368#_M1005_d N_A_27_368#_c_222_n N_A_27_368#_c_223_n
+ N_A_27_368#_c_224_n N_A_27_368#_c_233_n N_A_27_368#_c_225_n
+ N_A_27_368#_c_226_n N_A_27_368#_c_227_n PM_SKY130_FD_SC_LS__NOR3_2%A_27_368#
x_PM_SKY130_FD_SC_LS__NOR3_2%Y N_Y_M1006_s N_Y_M1008_d N_Y_M1003_s N_Y_c_274_n
+ N_Y_c_281_n N_Y_c_284_n N_Y_c_270_n Y Y Y Y N_Y_c_276_n Y
+ PM_SKY130_FD_SC_LS__NOR3_2%Y
x_PM_SKY130_FD_SC_LS__NOR3_2%A_306_368# N_A_306_368#_M1002_s
+ N_A_306_368#_M1001_d N_A_306_368#_c_317_n N_A_306_368#_c_315_n
+ N_A_306_368#_c_322_n N_A_306_368#_c_319_n N_A_306_368#_c_316_n
+ PM_SKY130_FD_SC_LS__NOR3_2%A_306_368#
x_PM_SKY130_FD_SC_LS__NOR3_2%VPWR N_VPWR_M1000_s N_VPWR_c_343_n VPWR
+ N_VPWR_c_344_n N_VPWR_c_345_n N_VPWR_c_342_n N_VPWR_c_347_n
+ PM_SKY130_FD_SC_LS__NOR3_2%VPWR
x_PM_SKY130_FD_SC_LS__NOR3_2%VGND N_VGND_M1006_d N_VGND_M1007_d N_VGND_c_378_n
+ N_VGND_c_379_n VGND N_VGND_c_380_n N_VGND_c_381_n N_VGND_c_382_n
+ N_VGND_c_383_n N_VGND_c_384_n PM_SKY130_FD_SC_LS__NOR3_2%VGND
cc_1 VNB N_C_c_57_n 0.0238316f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.22
cc_2 VNB C 0.0064001f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_3 VNB N_C_c_59_n 0.061852f $X=-0.19 $Y=-0.245 $X2=0.81 $Y2=1.385
cc_4 VNB N_B_c_97_n 0.0371541f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.22
cc_5 VNB N_B_c_98_n 0.0218521f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_6 VNB N_B_c_99_n 0.063754f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.765
cc_7 VNB N_B_c_100_n 0.0196703f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_8 VNB N_B_c_101_n 0.00315176f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_9 VNB B 0.00742405f $X=-0.19 $Y=-0.245 $X2=0.79 $Y2=1.295
cc_10 VNB N_A_c_160_n 0.0159305f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_11 VNB N_A_c_161_n 0.0171724f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_12 VNB N_A_c_162_n 0.00880223f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.4
cc_13 VNB N_A_c_163_n 0.0176973f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.22
cc_14 VNB N_A_c_164_n 0.0171751f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.492
cc_15 VNB N_A_c_165_n 0.009551f $X=-0.19 $Y=-0.245 $X2=0.79 $Y2=1.295
cc_16 VNB N_A_c_166_n 0.0169193f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_c_167_n 0.029959f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB A 0.0323167f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_c_169_n 0.0558262f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_Y_c_270_n 0.00280505f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB Y 0.0212531f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB Y 0.00704942f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB Y 0.033575f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VPWR_c_342_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0.79 $Y2=1.385
cc_25 VNB N_VGND_c_378_n 0.0185359f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.765
cc_26 VNB N_VGND_c_379_n 0.0188688f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_380_n 0.0252139f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_381_n 0.206462f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_382_n 0.0191515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_383_n 0.0280581f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_384_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VPB N_C_c_60_n 0.0175858f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_33 VPB N_C_c_61_n 0.0149425f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.765
cc_34 VPB N_C_c_59_n 0.0235519f $X=-0.19 $Y=1.66 $X2=0.81 $Y2=1.385
cc_35 VPB N_B_c_97_n 0.0219408f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.22
cc_36 VPB N_B_c_99_n 0.0328261f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.765
cc_37 VPB N_A_c_160_n 7.98165e-19 $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_38 VPB N_A_c_171_n 0.0211753f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_39 VPB N_A_c_163_n 7.82107e-19 $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.22
cc_40 VPB N_A_c_173_n 0.0202511f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_41 VPB N_A_27_368#_c_222_n 0.0322259f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.22
cc_42 VPB N_A_27_368#_c_223_n 0.00552368f $X=-0.19 $Y=1.66 $X2=0.81 $Y2=1.385
cc_43 VPB N_A_27_368#_c_224_n 0.00982439f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.492
cc_44 VPB N_A_27_368#_c_225_n 0.0151346f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_45 VPB N_A_27_368#_c_226_n 0.00752119f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_A_27_368#_c_227_n 0.0432125f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB N_Y_c_274_n 0.00202686f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_48 VPB Y 0.00293411f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 VPB N_Y_c_276_n 0.00767133f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_A_306_368#_c_315_n 0.00296428f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.4
cc_51 VPB N_A_306_368#_c_316_n 0.00247909f $X=-0.19 $Y=1.66 $X2=0.81 $Y2=1.385
cc_52 VPB N_VPWR_c_343_n 0.00653303f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_53 VPB N_VPWR_c_344_n 0.0520079f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_54 VPB N_VPWR_c_345_n 0.0298982f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_342_n 0.0647115f $X=-0.19 $Y=1.66 $X2=0.79 $Y2=1.385
cc_56 VPB N_VPWR_c_347_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 N_C_c_61_n N_B_c_97_n 0.00918779f $X=1.005 $Y=1.765 $X2=-0.19 $Y2=-0.245
cc_58 C N_B_c_97_n 9.60045e-19 $X=0.635 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_59 N_C_c_59_n N_B_c_97_n 0.0339258f $X=0.81 $Y=1.385 $X2=-0.19 $Y2=-0.245
cc_60 C N_B_c_98_n 0.00107469f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_61 C N_B_c_101_n 0.0146852f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_62 N_C_c_59_n N_B_c_101_n 0.00140882f $X=0.81 $Y=1.385 $X2=0 $Y2=0
cc_63 N_C_c_60_n N_A_27_368#_c_222_n 0.00975493f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_64 N_C_c_61_n N_A_27_368#_c_222_n 5.33746e-19 $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_65 N_C_c_60_n N_A_27_368#_c_223_n 0.0111147f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_66 N_C_c_61_n N_A_27_368#_c_223_n 0.012733f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_67 N_C_c_60_n N_A_27_368#_c_224_n 0.00262934f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_68 N_C_c_61_n N_A_27_368#_c_233_n 0.00616696f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_69 N_C_c_61_n N_A_27_368#_c_226_n 8.70506e-19 $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_70 N_C_c_59_n N_A_27_368#_c_226_n 4.57296e-19 $X=0.81 $Y=1.385 $X2=0 $Y2=0
cc_71 N_C_c_60_n N_Y_c_274_n 0.0122042f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_72 N_C_c_61_n N_Y_c_274_n 0.00230202f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_73 C N_Y_c_274_n 0.0274789f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_74 N_C_c_59_n N_Y_c_274_n 0.0207066f $X=0.81 $Y=1.385 $X2=0 $Y2=0
cc_75 N_C_c_57_n N_Y_c_281_n 0.0112f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_76 C N_Y_c_281_n 0.028324f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_77 N_C_c_59_n N_Y_c_281_n 0.0075351f $X=0.81 $Y=1.385 $X2=0 $Y2=0
cc_78 N_C_c_61_n N_Y_c_284_n 0.00875043f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_79 N_C_c_57_n Y 0.0124397f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_80 N_C_c_57_n Y 8.87593e-19 $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_81 N_C_c_57_n Y 0.01042f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_82 C Y 0.0225409f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_83 N_C_c_59_n Y 0.0056331f $X=0.81 $Y=1.385 $X2=0 $Y2=0
cc_84 N_C_c_60_n N_VPWR_c_344_n 0.00278257f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_85 N_C_c_61_n N_VPWR_c_344_n 0.00278271f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_86 N_C_c_60_n N_VPWR_c_342_n 0.00357777f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_87 N_C_c_61_n N_VPWR_c_342_n 0.00354368f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_88 N_C_c_57_n N_VGND_c_381_n 0.00453471f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_89 N_C_c_57_n N_VGND_c_382_n 0.00434272f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_90 N_C_c_57_n N_VGND_c_383_n 0.0110054f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_91 N_B_c_97_n N_A_c_160_n 0.0101827f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_92 N_B_c_100_n N_A_c_160_n 0.0129333f $X=2.925 $Y=1.465 $X2=0 $Y2=0
cc_93 N_B_c_97_n N_A_c_171_n 0.0113418f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_94 N_B_c_98_n N_A_c_161_n 0.0179489f $X=1.53 $Y=1.22 $X2=0 $Y2=0
cc_95 N_B_c_100_n N_A_c_162_n 0.00380862f $X=2.925 $Y=1.465 $X2=0 $Y2=0
cc_96 N_B_c_99_n N_A_c_163_n 0.0167686f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_97 N_B_c_100_n N_A_c_163_n 0.0129019f $X=2.925 $Y=1.465 $X2=0 $Y2=0
cc_98 B N_A_c_163_n 3.6606e-19 $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_99 N_B_c_99_n N_A_c_173_n 0.0130706f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_100 B N_A_c_164_n 0.00159669f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_101 N_B_c_97_n N_A_c_165_n 0.0221136f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_102 N_B_c_98_n N_A_c_165_n 0.00228878f $X=1.53 $Y=1.22 $X2=0 $Y2=0
cc_103 N_B_c_101_n N_A_c_165_n 0.0011932f $X=1.47 $Y=1.385 $X2=0 $Y2=0
cc_104 N_B_c_99_n N_A_c_166_n 0.00713314f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_105 N_B_c_100_n N_A_c_166_n 0.00855379f $X=2.925 $Y=1.465 $X2=0 $Y2=0
cc_106 B N_A_c_166_n 8.70735e-19 $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_107 N_B_c_99_n N_A_c_167_n 0.00549703f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_108 N_B_c_100_n N_A_c_167_n 0.00317985f $X=2.925 $Y=1.465 $X2=0 $Y2=0
cc_109 B N_A_c_167_n 3.63484e-19 $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_110 N_B_c_99_n A 0.0018366f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_111 N_B_c_100_n A 0.0114949f $X=2.925 $Y=1.465 $X2=0 $Y2=0
cc_112 B A 0.0242925f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_113 N_B_c_97_n N_A_27_368#_c_223_n 0.00318326f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_114 N_B_c_97_n N_A_27_368#_c_233_n 0.00616454f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_115 N_B_c_97_n N_A_27_368#_c_225_n 0.0158205f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_116 N_B_c_99_n N_A_27_368#_c_225_n 0.0214915f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_117 N_B_c_100_n N_A_27_368#_c_225_n 0.093824f $X=2.925 $Y=1.465 $X2=0 $Y2=0
cc_118 N_B_c_101_n N_A_27_368#_c_225_n 0.0233821f $X=1.47 $Y=1.385 $X2=0 $Y2=0
cc_119 B N_A_27_368#_c_225_n 0.0262111f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_120 N_B_c_101_n N_A_27_368#_c_226_n 7.62703e-19 $X=1.47 $Y=1.385 $X2=0 $Y2=0
cc_121 N_B_c_99_n N_A_27_368#_c_227_n 0.00143254f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_122 N_B_c_97_n N_Y_c_281_n 8.5738e-19 $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_123 N_B_c_98_n N_Y_c_281_n 0.0142961f $X=1.53 $Y=1.22 $X2=0 $Y2=0
cc_124 N_B_c_100_n N_Y_c_281_n 0.0144587f $X=2.925 $Y=1.465 $X2=0 $Y2=0
cc_125 N_B_c_101_n N_Y_c_281_n 0.0176193f $X=1.47 $Y=1.385 $X2=0 $Y2=0
cc_126 N_B_c_98_n N_Y_c_270_n 0.00261686f $X=1.53 $Y=1.22 $X2=0 $Y2=0
cc_127 N_B_c_97_n N_A_306_368#_c_317_n 0.00193585f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_128 N_B_c_97_n N_A_306_368#_c_315_n 0.00816586f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_129 N_B_c_99_n N_A_306_368#_c_319_n 0.0019041f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_130 N_B_c_99_n N_A_306_368#_c_316_n 0.00831152f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_131 N_B_c_99_n N_VPWR_c_343_n 6.55355e-19 $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_132 N_B_c_97_n N_VPWR_c_344_n 0.00445475f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_133 N_B_c_99_n N_VPWR_c_345_n 0.00445475f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_134 N_B_c_97_n N_VPWR_c_342_n 0.00858688f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_135 N_B_c_99_n N_VPWR_c_342_n 0.00861836f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_136 N_B_c_98_n N_VGND_c_378_n 0.00383152f $X=1.53 $Y=1.22 $X2=0 $Y2=0
cc_137 N_B_c_100_n N_VGND_c_379_n 0.0204916f $X=2.925 $Y=1.465 $X2=0 $Y2=0
cc_138 N_B_c_98_n N_VGND_c_381_n 0.00383029f $X=1.53 $Y=1.22 $X2=0 $Y2=0
cc_139 N_B_c_98_n N_VGND_c_383_n 0.00924883f $X=1.53 $Y=1.22 $X2=0 $Y2=0
cc_140 N_A_c_171_n N_A_27_368#_c_225_n 0.0118692f $X=1.935 $Y=1.765 $X2=0 $Y2=0
cc_141 N_A_c_173_n N_A_27_368#_c_225_n 0.0117043f $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_142 N_A_c_161_n N_Y_c_281_n 0.00265815f $X=2.03 $Y=1.185 $X2=0 $Y2=0
cc_143 N_A_c_165_n N_Y_c_281_n 0.00305887f $X=1.975 $Y=1.26 $X2=0 $Y2=0
cc_144 N_A_c_161_n N_Y_c_270_n 0.0055158f $X=2.03 $Y=1.185 $X2=0 $Y2=0
cc_145 N_A_c_171_n N_A_306_368#_c_315_n 2.60538e-19 $X=1.935 $Y=1.765 $X2=0
+ $Y2=0
cc_146 N_A_c_171_n N_A_306_368#_c_322_n 0.0132272f $X=1.935 $Y=1.765 $X2=0 $Y2=0
cc_147 N_A_c_173_n N_A_306_368#_c_322_n 0.012799f $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_148 N_A_c_173_n N_A_306_368#_c_316_n 2.3414e-19 $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_149 N_A_c_171_n N_VPWR_c_343_n 0.00318166f $X=1.935 $Y=1.765 $X2=0 $Y2=0
cc_150 N_A_c_173_n N_VPWR_c_343_n 0.00934717f $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_151 N_A_c_171_n N_VPWR_c_344_n 0.00461464f $X=1.935 $Y=1.765 $X2=0 $Y2=0
cc_152 N_A_c_173_n N_VPWR_c_345_n 0.00413917f $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_153 N_A_c_171_n N_VPWR_c_342_n 0.00908143f $X=1.935 $Y=1.765 $X2=0 $Y2=0
cc_154 N_A_c_173_n N_VPWR_c_342_n 0.0081781f $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_155 N_A_c_161_n N_VGND_c_378_n 0.00434272f $X=2.03 $Y=1.185 $X2=0 $Y2=0
cc_156 N_A_c_161_n N_VGND_c_379_n 0.0080629f $X=2.03 $Y=1.185 $X2=0 $Y2=0
cc_157 N_A_c_162_n N_VGND_c_379_n 0.00793039f $X=2.315 $Y=1.26 $X2=0 $Y2=0
cc_158 A N_VGND_c_379_n 0.0553698f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_159 N_A_c_169_n N_VGND_c_379_n 0.0117383f $X=2.815 $Y=0.475 $X2=0 $Y2=0
cc_160 A N_VGND_c_380_n 0.0298314f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_161 N_A_c_169_n N_VGND_c_380_n 0.0120882f $X=2.815 $Y=0.475 $X2=0 $Y2=0
cc_162 N_A_c_161_n N_VGND_c_381_n 0.00825771f $X=2.03 $Y=1.185 $X2=0 $Y2=0
cc_163 A N_VGND_c_381_n 0.0218461f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_164 N_A_c_169_n N_VGND_c_381_n 0.0154157f $X=2.815 $Y=0.475 $X2=0 $Y2=0
cc_165 N_A_c_161_n N_VGND_c_383_n 4.24281e-19 $X=2.03 $Y=1.185 $X2=0 $Y2=0
cc_166 N_A_27_368#_c_223_n N_Y_M1003_s 0.00250873f $X=1.145 $Y=2.99 $X2=0 $Y2=0
cc_167 N_A_27_368#_c_222_n N_Y_c_274_n 0.00245231f $X=0.28 $Y=2.145 $X2=0 $Y2=0
cc_168 N_A_27_368#_c_226_n N_Y_c_274_n 0.0132705f $X=1.315 $Y=1.805 $X2=0 $Y2=0
cc_169 N_A_27_368#_c_223_n N_Y_c_284_n 0.018923f $X=1.145 $Y=2.99 $X2=0 $Y2=0
cc_170 N_A_27_368#_c_233_n N_Y_c_284_n 0.0549755f $X=1.23 $Y=1.985 $X2=0 $Y2=0
cc_171 N_A_27_368#_M1003_d N_Y_c_276_n 0.00271132f $X=0.135 $Y=1.84 $X2=0 $Y2=0
cc_172 N_A_27_368#_c_222_n N_Y_c_276_n 0.0216158f $X=0.28 $Y=2.145 $X2=0 $Y2=0
cc_173 N_A_27_368#_c_225_n N_A_306_368#_M1002_s 0.00229612f $X=2.965 $Y=1.805
+ $X2=-0.19 $Y2=1.66
cc_174 N_A_27_368#_c_225_n N_A_306_368#_M1001_d 0.00197722f $X=2.965 $Y=1.805
+ $X2=0 $Y2=0
cc_175 N_A_27_368#_c_233_n N_A_306_368#_c_317_n 0.0117758f $X=1.23 $Y=1.985
+ $X2=0 $Y2=0
cc_176 N_A_27_368#_c_225_n N_A_306_368#_c_317_n 0.018674f $X=2.965 $Y=1.805
+ $X2=0 $Y2=0
cc_177 N_A_27_368#_c_223_n N_A_306_368#_c_315_n 0.0062448f $X=1.145 $Y=2.99
+ $X2=0 $Y2=0
cc_178 N_A_27_368#_c_233_n N_A_306_368#_c_315_n 0.0439022f $X=1.23 $Y=1.985
+ $X2=0 $Y2=0
cc_179 N_A_27_368#_c_225_n N_A_306_368#_c_322_n 0.0352288f $X=2.965 $Y=1.805
+ $X2=0 $Y2=0
cc_180 N_A_27_368#_c_225_n N_A_306_368#_c_319_n 0.0162332f $X=2.965 $Y=1.805
+ $X2=0 $Y2=0
cc_181 N_A_27_368#_c_227_n N_A_306_368#_c_316_n 0.0281768f $X=3.08 $Y=1.985
+ $X2=0 $Y2=0
cc_182 N_A_27_368#_c_225_n N_VPWR_M1000_s 0.00219516f $X=2.965 $Y=1.805
+ $X2=-0.19 $Y2=1.66
cc_183 N_A_27_368#_c_223_n N_VPWR_c_344_n 0.0563945f $X=1.145 $Y=2.99 $X2=0
+ $Y2=0
cc_184 N_A_27_368#_c_224_n N_VPWR_c_344_n 0.0235677f $X=0.445 $Y=2.99 $X2=0
+ $Y2=0
cc_185 N_A_27_368#_c_227_n N_VPWR_c_345_n 0.0124046f $X=3.08 $Y=1.985 $X2=0
+ $Y2=0
cc_186 N_A_27_368#_c_223_n N_VPWR_c_342_n 0.0316233f $X=1.145 $Y=2.99 $X2=0
+ $Y2=0
cc_187 N_A_27_368#_c_224_n N_VPWR_c_342_n 0.0127557f $X=0.445 $Y=2.99 $X2=0
+ $Y2=0
cc_188 N_A_27_368#_c_227_n N_VPWR_c_342_n 0.0102675f $X=3.08 $Y=1.985 $X2=0
+ $Y2=0
cc_189 N_Y_c_281_n N_VGND_M1006_d 0.0266486f $X=1.65 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_190 N_Y_c_270_n N_VGND_c_378_n 0.0145947f $X=1.815 $Y=0.515 $X2=0 $Y2=0
cc_191 N_Y_c_270_n N_VGND_c_379_n 0.0191389f $X=1.815 $Y=0.515 $X2=0 $Y2=0
cc_192 N_Y_c_281_n N_VGND_c_381_n 0.0128359f $X=1.65 $Y=0.925 $X2=0 $Y2=0
cc_193 N_Y_c_270_n N_VGND_c_381_n 0.0120104f $X=1.815 $Y=0.515 $X2=0 $Y2=0
cc_194 Y N_VGND_c_381_n 0.011995f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_195 Y N_VGND_c_382_n 0.0145556f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_196 N_Y_c_281_n N_VGND_c_383_n 0.0573941f $X=1.65 $Y=0.925 $X2=0 $Y2=0
cc_197 N_Y_c_270_n N_VGND_c_383_n 0.0133889f $X=1.815 $Y=0.515 $X2=0 $Y2=0
cc_198 Y N_VGND_c_383_n 0.0121582f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_199 N_A_306_368#_c_322_n N_VPWR_M1000_s 0.00438498f $X=2.515 $Y=2.145
+ $X2=-0.19 $Y2=1.66
cc_200 N_A_306_368#_c_315_n N_VPWR_c_343_n 0.00241304f $X=1.68 $Y=2.485 $X2=0
+ $Y2=0
cc_201 N_A_306_368#_c_322_n N_VPWR_c_343_n 0.0177842f $X=2.515 $Y=2.145 $X2=0
+ $Y2=0
cc_202 N_A_306_368#_c_316_n N_VPWR_c_343_n 0.0233151f $X=2.63 $Y=2.485 $X2=0
+ $Y2=0
cc_203 N_A_306_368#_c_315_n N_VPWR_c_344_n 0.0152042f $X=1.68 $Y=2.485 $X2=0
+ $Y2=0
cc_204 N_A_306_368#_c_316_n N_VPWR_c_345_n 0.01288f $X=2.63 $Y=2.485 $X2=0 $Y2=0
cc_205 N_A_306_368#_c_315_n N_VPWR_c_342_n 0.0121192f $X=1.68 $Y=2.485 $X2=0
+ $Y2=0
cc_206 N_A_306_368#_c_316_n N_VPWR_c_342_n 0.0102615f $X=2.63 $Y=2.485 $X2=0
+ $Y2=0
