* File: sky130_fd_sc_ls__clkbuf_16.pxi.spice
* Created: Fri Aug 28 13:08:23 2020
* 
x_PM_SKY130_FD_SC_LS__CLKBUF_16%A N_A_M1022_g N_A_c_202_n N_A_M1020_g
+ N_A_M1029_g N_A_c_203_n N_A_M1021_g N_A_M1030_g N_A_c_204_n N_A_M1025_g
+ N_A_M1036_g N_A_c_205_n N_A_M1038_g A A A A N_A_c_201_n
+ PM_SKY130_FD_SC_LS__CLKBUF_16%A
x_PM_SKY130_FD_SC_LS__CLKBUF_16%A_114_74# N_A_114_74#_M1022_s
+ N_A_114_74#_M1030_s N_A_114_74#_M1020_d N_A_114_74#_M1025_d
+ N_A_114_74#_M1003_g N_A_114_74#_c_285_n N_A_114_74#_c_334_n
+ N_A_114_74#_M1000_g N_A_114_74#_M1005_g N_A_114_74#_c_287_n
+ N_A_114_74#_c_336_n N_A_114_74#_M1001_g N_A_114_74#_M1008_g
+ N_A_114_74#_c_289_n N_A_114_74#_c_338_n N_A_114_74#_M1002_g
+ N_A_114_74#_M1010_g N_A_114_74#_c_291_n N_A_114_74#_c_340_n
+ N_A_114_74#_M1004_g N_A_114_74#_M1012_g N_A_114_74#_c_293_n
+ N_A_114_74#_c_342_n N_A_114_74#_M1006_g N_A_114_74#_M1013_g
+ N_A_114_74#_c_295_n N_A_114_74#_c_344_n N_A_114_74#_M1007_g
+ N_A_114_74#_M1014_g N_A_114_74#_c_297_n N_A_114_74#_c_346_n
+ N_A_114_74#_M1009_g N_A_114_74#_M1015_g N_A_114_74#_c_299_n
+ N_A_114_74#_c_348_n N_A_114_74#_M1011_g N_A_114_74#_M1018_g
+ N_A_114_74#_c_301_n N_A_114_74#_c_350_n N_A_114_74#_M1016_g
+ N_A_114_74#_M1019_g N_A_114_74#_c_303_n N_A_114_74#_c_352_n
+ N_A_114_74#_M1017_g N_A_114_74#_c_304_n N_A_114_74#_M1027_g
+ N_A_114_74#_c_354_n N_A_114_74#_M1023_g N_A_114_74#_M1028_g
+ N_A_114_74#_c_307_n N_A_114_74#_c_356_n N_A_114_74#_M1024_g
+ N_A_114_74#_c_308_n N_A_114_74#_c_358_n N_A_114_74#_M1026_g
+ N_A_114_74#_M1031_g N_A_114_74#_c_310_n N_A_114_74#_c_360_n
+ N_A_114_74#_M1033_g N_A_114_74#_M1032_g N_A_114_74#_c_312_n
+ N_A_114_74#_c_362_n N_A_114_74#_M1034_g N_A_114_74#_M1037_g
+ N_A_114_74#_c_314_n N_A_114_74#_c_364_n N_A_114_74#_M1035_g
+ N_A_114_74#_M1039_g N_A_114_74#_c_316_n N_A_114_74#_c_372_n
+ N_A_114_74#_c_365_n N_A_114_74#_c_317_n N_A_114_74#_c_318_n
+ N_A_114_74#_c_386_n N_A_114_74#_c_319_n N_A_114_74#_c_366_n
+ N_A_114_74#_c_320_n N_A_114_74#_c_321_n N_A_114_74#_c_322_n
+ N_A_114_74#_c_323_n N_A_114_74#_c_408_n N_A_114_74#_c_324_n
+ N_A_114_74#_c_325_n N_A_114_74#_c_326_n N_A_114_74#_c_327_n
+ N_A_114_74#_c_328_n N_A_114_74#_c_329_n N_A_114_74#_c_330_n
+ N_A_114_74#_c_331_n N_A_114_74#_c_332_n
+ PM_SKY130_FD_SC_LS__CLKBUF_16%A_114_74#
x_PM_SKY130_FD_SC_LS__CLKBUF_16%VPWR N_VPWR_M1020_s N_VPWR_M1021_s
+ N_VPWR_M1038_s N_VPWR_M1001_s N_VPWR_M1004_s N_VPWR_M1007_s N_VPWR_M1011_s
+ N_VPWR_M1017_s N_VPWR_M1024_s N_VPWR_M1033_s N_VPWR_M1035_s N_VPWR_c_755_n
+ N_VPWR_c_756_n N_VPWR_c_757_n N_VPWR_c_758_n N_VPWR_c_759_n N_VPWR_c_760_n
+ N_VPWR_c_761_n N_VPWR_c_762_n N_VPWR_c_763_n N_VPWR_c_764_n N_VPWR_c_765_n
+ N_VPWR_c_766_n N_VPWR_c_767_n N_VPWR_c_768_n N_VPWR_c_769_n N_VPWR_c_770_n
+ N_VPWR_c_771_n N_VPWR_c_772_n N_VPWR_c_773_n N_VPWR_c_774_n N_VPWR_c_775_n
+ N_VPWR_c_776_n N_VPWR_c_777_n N_VPWR_c_778_n VPWR N_VPWR_c_779_n
+ N_VPWR_c_780_n N_VPWR_c_781_n N_VPWR_c_782_n N_VPWR_c_783_n N_VPWR_c_784_n
+ N_VPWR_c_785_n N_VPWR_c_786_n N_VPWR_c_754_n
+ PM_SKY130_FD_SC_LS__CLKBUF_16%VPWR
x_PM_SKY130_FD_SC_LS__CLKBUF_16%X N_X_M1003_d N_X_M1008_d N_X_M1012_d
+ N_X_M1014_d N_X_M1018_d N_X_M1027_d N_X_M1031_d N_X_M1037_d N_X_M1000_d
+ N_X_M1002_d N_X_M1006_d N_X_M1009_d N_X_M1016_d N_X_M1023_d N_X_M1026_d
+ N_X_M1034_d N_X_c_946_n N_X_c_956_n N_X_c_947_n N_X_c_948_n N_X_c_949_n
+ N_X_c_950_n N_X_c_951_n N_X_c_962_n N_X_c_952_n N_X_c_964_n N_X_c_953_n
+ N_X_c_954_n N_X_c_966_n N_X_c_967_n N_X_c_968_n N_X_c_969_n N_X_c_970_n X
+ N_X_c_971_n N_X_c_972_n N_X_c_973_n N_X_c_974_n N_X_c_975_n N_X_c_976_n
+ N_X_c_977_n N_X_c_1105_n N_X_c_1132_n PM_SKY130_FD_SC_LS__CLKBUF_16%X
x_PM_SKY130_FD_SC_LS__CLKBUF_16%VGND N_VGND_M1022_d N_VGND_M1029_d
+ N_VGND_M1036_d N_VGND_M1005_s N_VGND_M1010_s N_VGND_M1013_s N_VGND_M1015_s
+ N_VGND_M1019_s N_VGND_M1028_s N_VGND_M1032_s N_VGND_M1039_s N_VGND_c_1212_n
+ N_VGND_c_1213_n N_VGND_c_1214_n N_VGND_c_1215_n N_VGND_c_1216_n
+ N_VGND_c_1217_n N_VGND_c_1218_n N_VGND_c_1219_n N_VGND_c_1220_n
+ N_VGND_c_1221_n N_VGND_c_1222_n N_VGND_c_1223_n N_VGND_c_1224_n
+ N_VGND_c_1225_n N_VGND_c_1226_n N_VGND_c_1227_n N_VGND_c_1228_n
+ N_VGND_c_1229_n N_VGND_c_1230_n N_VGND_c_1231_n N_VGND_c_1232_n
+ N_VGND_c_1233_n VGND N_VGND_c_1234_n N_VGND_c_1235_n N_VGND_c_1236_n
+ N_VGND_c_1237_n N_VGND_c_1238_n N_VGND_c_1239_n N_VGND_c_1240_n
+ N_VGND_c_1241_n N_VGND_c_1242_n N_VGND_c_1243_n N_VGND_c_1244_n
+ PM_SKY130_FD_SC_LS__CLKBUF_16%VGND
cc_1 VNB N_A_M1022_g 0.0550782f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.58
cc_2 VNB N_A_M1029_g 0.0383342f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.58
cc_3 VNB N_A_M1030_g 0.0382364f $X=-0.19 $Y=-0.245 $X2=1.375 $Y2=0.58
cc_4 VNB N_A_M1036_g 0.0401024f $X=-0.19 $Y=-0.245 $X2=1.805 $Y2=0.58
cc_5 VNB A 0.0197254f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_6 VNB N_A_c_201_n 0.074705f $X=-0.19 $Y=-0.245 $X2=1.805 $Y2=1.557
cc_7 VNB N_A_114_74#_M1003_g 0.0338011f $X=-0.19 $Y=-0.245 $X2=1.375 $Y2=1.35
cc_8 VNB N_A_114_74#_c_285_n 0.00707624f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_114_74#_M1005_g 0.0316604f $X=-0.19 $Y=-0.245 $X2=1.805 $Y2=0.58
cc_10 VNB N_A_114_74#_c_287_n 0.00734506f $X=-0.19 $Y=-0.245 $X2=1.86 $Y2=2.4
cc_11 VNB N_A_114_74#_M1008_g 0.03169f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_114_74#_c_289_n 0.00680742f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_114_74#_M1010_g 0.0316814f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.557
cc_14 VNB N_A_114_74#_c_291_n 0.00734745f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=1.557
cc_15 VNB N_A_114_74#_M1012_g 0.0316038f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.565
cc_16 VNB N_A_114_74#_c_293_n 0.00680951f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.565
cc_17 VNB N_A_114_74#_M1013_g 0.0324981f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=1.565
cc_18 VNB N_A_114_74#_c_295_n 0.00734966f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_114_74#_M1014_g 0.0315189f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_114_74#_c_297_n 0.00681093f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_114_74#_M1015_g 0.0324679f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_114_74#_c_299_n 0.00734891f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_114_74#_M1018_g 0.0315167f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_114_74#_c_301_n 0.00681063f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_114_74#_M1019_g 0.0324679f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_114_74#_c_303_n 0.00734826f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_114_74#_c_304_n 0.00680992f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_114_74#_M1027_g 0.0315167f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_114_74#_M1028_g 0.0324679f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_114_74#_c_307_n 0.00734788f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_114_74#_c_308_n 0.00680906f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_114_74#_M1031_g 0.0315167f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_114_74#_c_310_n 0.00746164f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_114_74#_M1032_g 0.0324679f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_114_74#_c_312_n 0.00692273f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_114_74#_M1037_g 0.0315167f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_114_74#_c_314_n 0.0116517f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_114_74#_M1039_g 0.0449212f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_114_74#_c_316_n 0.00360655f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_114_74#_c_317_n 0.00956284f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_114_74#_c_318_n 0.00189788f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_114_74#_c_319_n 0.00380649f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_114_74#_c_320_n 0.00390804f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_114_74#_c_321_n 0.0101323f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_114_74#_c_322_n 0.00455461f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_114_74#_c_323_n 0.00189788f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_114_74#_c_324_n 0.00194085f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_114_74#_c_325_n 0.00189558f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_114_74#_c_326_n 0.00238431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_114_74#_c_327_n 0.00250109f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_114_74#_c_328_n 0.00250109f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_114_74#_c_329_n 0.00250109f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_114_74#_c_330_n 0.0568387f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_114_74#_c_331_n 0.00275453f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_114_74#_c_332_n 0.358908f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VPWR_c_754_n 0.40251f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_X_c_946_n 0.0124197f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.565
cc_58 VNB N_X_c_947_n 0.0120395f $X=-0.19 $Y=-0.245 $X2=1.605 $Y2=1.565
cc_59 VNB N_X_c_948_n 0.00757647f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_X_c_949_n 0.00760885f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_X_c_950_n 0.00759431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_X_c_951_n 0.00758503f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_X_c_952_n 0.00754993f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_X_c_953_n 0.00219225f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_X_c_954_n 0.00921522f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_1212_n 0.010678f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_1213_n 0.0320442f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_1214_n 0.00626911f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.515
cc_69 VNB N_VGND_c_1215_n 0.00869356f $X=-0.19 $Y=-0.245 $X2=1.375 $Y2=1.557
cc_70 VNB N_VGND_c_1216_n 0.00730898f $X=-0.19 $Y=-0.245 $X2=1.605 $Y2=1.515
cc_71 VNB N_VGND_c_1217_n 0.00715012f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1218_n 0.0172943f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.565
cc_73 VNB N_VGND_c_1219_n 0.0050287f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1220_n 0.00494723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1221_n 0.00494723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1222_n 0.00494723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1223_n 0.00494723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1224_n 0.0120272f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1225_n 0.0243692f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1226_n 0.0172524f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1227_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1228_n 0.0178889f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1229_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1230_n 0.0194689f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1231_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1232_n 0.0184013f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1233_n 0.00432782f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1234_n 0.0170705f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1235_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1236_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_VGND_c_1237_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_VGND_c_1238_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_VGND_c_1239_n 0.00606636f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_VGND_c_1240_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_VGND_c_1241_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_VGND_c_1242_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_VGND_c_1243_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_VGND_c_1244_n 0.508369f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VPB N_A_c_202_n 0.0179811f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.765
cc_100 VPB N_A_c_203_n 0.0155127f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=1.765
cc_101 VPB N_A_c_204_n 0.0155094f $X=-0.19 $Y=1.66 $X2=1.41 $Y2=1.765
cc_102 VPB N_A_c_205_n 0.0159315f $X=-0.19 $Y=1.66 $X2=1.86 $Y2=1.765
cc_103 VPB A 0.0185625f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.58
cc_104 VPB N_A_c_201_n 0.0478109f $X=-0.19 $Y=1.66 $X2=1.805 $Y2=1.557
cc_105 VPB N_A_114_74#_c_285_n 7.12715e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_A_114_74#_c_334_n 0.0204155f $X=-0.19 $Y=1.66 $X2=1.41 $Y2=1.765
cc_107 VPB N_A_114_74#_c_287_n 7.3979e-19 $X=-0.19 $Y=1.66 $X2=1.86 $Y2=2.4
cc_108 VPB N_A_114_74#_c_336_n 0.0208317f $X=-0.19 $Y=1.66 $X2=1.86 $Y2=2.4
cc_109 VPB N_A_114_74#_c_289_n 6.85639e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_110 VPB N_A_114_74#_c_338_n 0.0200162f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.557
cc_111 VPB N_A_114_74#_c_291_n 7.40031e-19 $X=-0.19 $Y=1.66 $X2=1.41 $Y2=1.557
cc_112 VPB N_A_114_74#_c_340_n 0.0208318f $X=-0.19 $Y=1.66 $X2=1.605 $Y2=1.557
cc_113 VPB N_A_114_74#_c_293_n 6.8585e-19 $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.565
cc_114 VPB N_A_114_74#_c_342_n 0.0200167f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.565
cc_115 VPB N_A_114_74#_c_295_n 7.40253e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_A_114_74#_c_344_n 0.0208201f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_A_114_74#_c_297_n 6.85993e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_A_114_74#_c_346_n 0.0200126f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_A_114_74#_c_299_n 7.40178e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_A_114_74#_c_348_n 0.0208228f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_A_114_74#_c_301_n 6.85962e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_A_114_74#_c_350_n 0.0200127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_A_114_74#_c_303_n 7.40112e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_A_114_74#_c_352_n 0.0208316f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_A_114_74#_c_304_n 6.85891e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 VPB N_A_114_74#_c_354_n 0.0200161f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_127 VPB N_A_114_74#_c_307_n 7.40074e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_A_114_74#_c_356_n 0.0208332f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_129 VPB N_A_114_74#_c_308_n 6.85805e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_A_114_74#_c_358_n 0.0202682f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_A_114_74#_c_310_n 7.51532e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_A_114_74#_c_360_n 0.0210662f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_A_114_74#_c_312_n 6.97253e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_A_114_74#_c_362_n 0.0213194f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_A_114_74#_c_314_n 0.00117356f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_A_114_74#_c_364_n 0.0276327f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_A_114_74#_c_365_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_A_114_74#_c_366_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_A_114_74#_c_322_n 0.00312895f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_140 VPB N_VPWR_c_755_n 0.0107598f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_756_n 0.0495498f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_142 VPB N_VPWR_c_757_n 0.00799266f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.557
cc_143 VPB N_VPWR_c_758_n 0.00516214f $X=-0.19 $Y=1.66 $X2=1.605 $Y2=1.557
cc_144 VPB N_VPWR_c_759_n 0.00263129f $X=-0.19 $Y=1.66 $X2=1.86 $Y2=1.557
cc_145 VPB N_VPWR_c_760_n 0.00261791f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_146 VPB N_VPWR_c_761_n 0.00261791f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_147 VPB N_VPWR_c_762_n 0.00261791f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_148 VPB N_VPWR_c_763_n 0.0161731f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_149 VPB N_VPWR_c_764_n 0.00261791f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_150 VPB N_VPWR_c_765_n 0.00261791f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_151 VPB N_VPWR_c_766_n 0.00505013f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_152 VPB N_VPWR_c_767_n 0.0121701f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_153 VPB N_VPWR_c_768_n 0.0455354f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_154 VPB N_VPWR_c_769_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_155 VPB N_VPWR_c_770_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_156 VPB N_VPWR_c_771_n 0.016296f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_157 VPB N_VPWR_c_772_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_158 VPB N_VPWR_c_773_n 0.0161731f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_159 VPB N_VPWR_c_774_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_160 VPB N_VPWR_c_775_n 0.0162121f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_161 VPB N_VPWR_c_776_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_162 VPB N_VPWR_c_777_n 0.016134f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_163 VPB N_VPWR_c_778_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_164 VPB N_VPWR_c_779_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_165 VPB N_VPWR_c_780_n 0.0161731f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_166 VPB N_VPWR_c_781_n 0.016134f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_167 VPB N_VPWR_c_782_n 0.0167991f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_168 VPB N_VPWR_c_783_n 0.00461173f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_169 VPB N_VPWR_c_784_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_170 VPB N_VPWR_c_785_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_171 VPB N_VPWR_c_786_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_172 VPB N_VPWR_c_754_n 0.103017f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_173 VPB N_X_c_946_n 0.0018252f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.565
cc_174 VPB N_X_c_956_n 0.00233969f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.565
cc_175 VPB N_X_c_947_n 2.50902e-19 $X=-0.19 $Y=1.66 $X2=1.605 $Y2=1.565
cc_176 VPB N_X_c_948_n 2.81093e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_177 VPB N_X_c_949_n 2.79936e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_178 VPB N_X_c_950_n 2.76924e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_179 VPB N_X_c_951_n 2.75001e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_180 VPB N_X_c_962_n 0.00222879f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_181 VPB N_X_c_952_n 4.26117e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_182 VPB N_X_c_964_n 0.00216056f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_183 VPB N_X_c_954_n 2.73116e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_184 VPB N_X_c_966_n 0.00219508f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_185 VPB N_X_c_967_n 0.00250782f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_186 VPB N_X_c_968_n 0.00232284f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_187 VPB N_X_c_969_n 0.00205843f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_188 VPB N_X_c_970_n 0.00220836f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_189 VPB N_X_c_971_n 0.00211605f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_190 VPB N_X_c_972_n 0.00207077f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_191 VPB N_X_c_973_n 0.00216153f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_192 VPB N_X_c_974_n 0.00211605f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_193 VPB N_X_c_975_n 0.00211605f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_194 VPB N_X_c_976_n 0.00216153f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_195 VPB N_X_c_977_n 0.00225625f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_196 N_A_M1036_g N_A_114_74#_M1003_g 0.0270312f $X=1.805 $Y=0.58 $X2=0 $Y2=0
cc_197 N_A_c_205_n N_A_114_74#_c_334_n 0.0212204f $X=1.86 $Y=1.765 $X2=0 $Y2=0
cc_198 N_A_M1022_g N_A_114_74#_c_316_n 0.0145444f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_199 N_A_M1029_g N_A_114_74#_c_316_n 0.00268841f $X=0.925 $Y=0.58 $X2=0 $Y2=0
cc_200 N_A_c_202_n N_A_114_74#_c_372_n 0.00203651f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_201 N_A_c_203_n N_A_114_74#_c_372_n 4.27055e-19 $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_202 A N_A_114_74#_c_372_n 0.0237598f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_203 N_A_c_201_n N_A_114_74#_c_372_n 0.00144162f $X=1.805 $Y=1.557 $X2=0 $Y2=0
cc_204 N_A_c_202_n N_A_114_74#_c_365_n 0.00960826f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_205 N_A_c_203_n N_A_114_74#_c_365_n 0.0103431f $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_206 N_A_c_204_n N_A_114_74#_c_365_n 6.45594e-19 $X=1.41 $Y=1.765 $X2=0 $Y2=0
cc_207 N_A_M1029_g N_A_114_74#_c_317_n 0.0146415f $X=0.925 $Y=0.58 $X2=0 $Y2=0
cc_208 N_A_M1030_g N_A_114_74#_c_317_n 0.0114202f $X=1.375 $Y=0.58 $X2=0 $Y2=0
cc_209 A N_A_114_74#_c_317_n 0.0416557f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_210 N_A_c_201_n N_A_114_74#_c_317_n 0.0026381f $X=1.805 $Y=1.557 $X2=0 $Y2=0
cc_211 N_A_M1022_g N_A_114_74#_c_318_n 0.010444f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_212 A N_A_114_74#_c_318_n 0.0188918f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_213 N_A_c_201_n N_A_114_74#_c_318_n 0.00229418f $X=1.805 $Y=1.557 $X2=0 $Y2=0
cc_214 N_A_c_203_n N_A_114_74#_c_386_n 0.0120074f $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_215 N_A_c_204_n N_A_114_74#_c_386_n 0.0120074f $X=1.41 $Y=1.765 $X2=0 $Y2=0
cc_216 A N_A_114_74#_c_386_n 0.0608989f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_217 N_A_c_201_n N_A_114_74#_c_386_n 0.00131001f $X=1.805 $Y=1.557 $X2=0 $Y2=0
cc_218 N_A_M1029_g N_A_114_74#_c_319_n 7.00296e-19 $X=0.925 $Y=0.58 $X2=0 $Y2=0
cc_219 N_A_M1030_g N_A_114_74#_c_319_n 0.0106356f $X=1.375 $Y=0.58 $X2=0 $Y2=0
cc_220 N_A_M1036_g N_A_114_74#_c_319_n 0.00476228f $X=1.805 $Y=0.58 $X2=0 $Y2=0
cc_221 N_A_c_203_n N_A_114_74#_c_366_n 6.46364e-19 $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_222 N_A_c_204_n N_A_114_74#_c_366_n 0.0104016f $X=1.41 $Y=1.765 $X2=0 $Y2=0
cc_223 N_A_c_205_n N_A_114_74#_c_366_n 0.0105164f $X=1.86 $Y=1.765 $X2=0 $Y2=0
cc_224 N_A_M1036_g N_A_114_74#_c_320_n 0.016885f $X=1.805 $Y=0.58 $X2=0 $Y2=0
cc_225 A N_A_114_74#_c_320_n 0.0078649f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_226 N_A_c_201_n N_A_114_74#_c_320_n 0.00270984f $X=1.805 $Y=1.557 $X2=0 $Y2=0
cc_227 N_A_M1036_g N_A_114_74#_c_321_n 0.00435841f $X=1.805 $Y=0.58 $X2=0 $Y2=0
cc_228 A N_A_114_74#_c_321_n 0.00414156f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_229 N_A_c_201_n N_A_114_74#_c_321_n 4.75687e-19 $X=1.805 $Y=1.557 $X2=0 $Y2=0
cc_230 N_A_c_205_n N_A_114_74#_c_322_n 0.00214468f $X=1.86 $Y=1.765 $X2=0 $Y2=0
cc_231 A N_A_114_74#_c_322_n 0.0294048f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_232 N_A_c_201_n N_A_114_74#_c_322_n 0.00323859f $X=1.805 $Y=1.557 $X2=0 $Y2=0
cc_233 N_A_M1030_g N_A_114_74#_c_323_n 0.00277828f $X=1.375 $Y=0.58 $X2=0 $Y2=0
cc_234 A N_A_114_74#_c_323_n 0.0188918f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_235 N_A_c_201_n N_A_114_74#_c_323_n 0.00229418f $X=1.805 $Y=1.557 $X2=0 $Y2=0
cc_236 N_A_c_204_n N_A_114_74#_c_408_n 4.54092e-19 $X=1.41 $Y=1.765 $X2=0 $Y2=0
cc_237 N_A_c_205_n N_A_114_74#_c_408_n 0.0161722f $X=1.86 $Y=1.765 $X2=0 $Y2=0
cc_238 N_A_c_201_n N_A_114_74#_c_408_n 0.00130859f $X=1.805 $Y=1.557 $X2=0 $Y2=0
cc_239 N_A_M1036_g N_A_114_74#_c_330_n 0.00366588f $X=1.805 $Y=0.58 $X2=0 $Y2=0
cc_240 A N_A_114_74#_c_330_n 0.00180161f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_241 N_A_c_201_n N_A_114_74#_c_330_n 0.00120791f $X=1.805 $Y=1.557 $X2=0 $Y2=0
cc_242 N_A_c_201_n N_A_114_74#_c_332_n 0.0175059f $X=1.805 $Y=1.557 $X2=0 $Y2=0
cc_243 N_A_c_202_n N_VPWR_c_756_n 0.00831454f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_244 A N_VPWR_c_756_n 0.0215956f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_245 N_A_c_203_n N_VPWR_c_757_n 0.00486623f $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_246 N_A_c_204_n N_VPWR_c_757_n 0.00486623f $X=1.41 $Y=1.765 $X2=0 $Y2=0
cc_247 N_A_c_205_n N_VPWR_c_758_n 0.00527858f $X=1.86 $Y=1.765 $X2=0 $Y2=0
cc_248 N_A_c_202_n N_VPWR_c_769_n 0.00445602f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_249 N_A_c_203_n N_VPWR_c_769_n 0.00445602f $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_250 N_A_c_204_n N_VPWR_c_779_n 0.00445602f $X=1.41 $Y=1.765 $X2=0 $Y2=0
cc_251 N_A_c_205_n N_VPWR_c_779_n 0.00445602f $X=1.86 $Y=1.765 $X2=0 $Y2=0
cc_252 N_A_c_202_n N_VPWR_c_754_n 0.008611f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_253 N_A_c_203_n N_VPWR_c_754_n 0.00857589f $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_254 N_A_c_204_n N_VPWR_c_754_n 0.00857589f $X=1.41 $Y=1.765 $X2=0 $Y2=0
cc_255 N_A_c_205_n N_VPWR_c_754_n 0.00857762f $X=1.86 $Y=1.765 $X2=0 $Y2=0
cc_256 N_A_c_205_n N_X_c_946_n 2.98438e-19 $X=1.86 $Y=1.765 $X2=0 $Y2=0
cc_257 N_A_M1022_g N_VGND_c_1213_n 0.00453696f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_258 A N_VGND_c_1213_n 0.00964677f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_259 N_A_M1022_g N_VGND_c_1214_n 5.07062e-19 $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_260 N_A_M1029_g N_VGND_c_1214_n 0.00935764f $X=0.925 $Y=0.58 $X2=0 $Y2=0
cc_261 N_A_M1030_g N_VGND_c_1214_n 0.00328886f $X=1.375 $Y=0.58 $X2=0 $Y2=0
cc_262 N_A_M1030_g N_VGND_c_1215_n 5.0842e-19 $X=1.375 $Y=0.58 $X2=0 $Y2=0
cc_263 N_A_M1036_g N_VGND_c_1215_n 0.00983752f $X=1.805 $Y=0.58 $X2=0 $Y2=0
cc_264 N_A_M1022_g N_VGND_c_1226_n 0.00434272f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_265 N_A_M1029_g N_VGND_c_1226_n 0.00383152f $X=0.925 $Y=0.58 $X2=0 $Y2=0
cc_266 N_A_M1030_g N_VGND_c_1228_n 0.00434272f $X=1.375 $Y=0.58 $X2=0 $Y2=0
cc_267 N_A_M1036_g N_VGND_c_1228_n 0.00383152f $X=1.805 $Y=0.58 $X2=0 $Y2=0
cc_268 N_A_M1022_g N_VGND_c_1244_n 0.00823942f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_269 N_A_M1029_g N_VGND_c_1244_n 0.0075754f $X=0.925 $Y=0.58 $X2=0 $Y2=0
cc_270 N_A_M1030_g N_VGND_c_1244_n 0.00820929f $X=1.375 $Y=0.58 $X2=0 $Y2=0
cc_271 N_A_M1036_g N_VGND_c_1244_n 0.0075754f $X=1.805 $Y=0.58 $X2=0 $Y2=0
cc_272 N_A_114_74#_c_386_n N_VPWR_M1021_s 0.00408911f $X=1.47 $Y=2.035 $X2=0
+ $Y2=0
cc_273 N_A_114_74#_c_322_n N_VPWR_M1038_s 0.00157395f $X=2.05 $Y=1.95 $X2=0
+ $Y2=0
cc_274 N_A_114_74#_c_408_n N_VPWR_M1038_s 0.00390109f $X=2.05 $Y=2.035 $X2=0
+ $Y2=0
cc_275 N_A_114_74#_c_372_n N_VPWR_c_756_n 0.0121024f $X=0.735 $Y=2.12 $X2=0
+ $Y2=0
cc_276 N_A_114_74#_c_365_n N_VPWR_c_756_n 0.0576605f $X=0.735 $Y=2.815 $X2=0
+ $Y2=0
cc_277 N_A_114_74#_c_365_n N_VPWR_c_757_n 0.0449718f $X=0.735 $Y=2.815 $X2=0
+ $Y2=0
cc_278 N_A_114_74#_c_386_n N_VPWR_c_757_n 0.0136682f $X=1.47 $Y=2.035 $X2=0
+ $Y2=0
cc_279 N_A_114_74#_c_366_n N_VPWR_c_757_n 0.0449718f $X=1.635 $Y=2.815 $X2=0
+ $Y2=0
cc_280 N_A_114_74#_c_334_n N_VPWR_c_758_n 0.00936797f $X=2.32 $Y=1.765 $X2=0
+ $Y2=0
cc_281 N_A_114_74#_c_336_n N_VPWR_c_758_n 5.08089e-19 $X=2.77 $Y=1.765 $X2=0
+ $Y2=0
cc_282 N_A_114_74#_c_366_n N_VPWR_c_758_n 0.0462948f $X=1.635 $Y=2.815 $X2=0
+ $Y2=0
cc_283 N_A_114_74#_c_408_n N_VPWR_c_758_n 0.0108656f $X=2.05 $Y=2.035 $X2=0
+ $Y2=0
cc_284 N_A_114_74#_c_334_n N_VPWR_c_759_n 5.62467e-19 $X=2.32 $Y=1.765 $X2=0
+ $Y2=0
cc_285 N_A_114_74#_c_336_n N_VPWR_c_759_n 0.0130723f $X=2.77 $Y=1.765 $X2=0
+ $Y2=0
cc_286 N_A_114_74#_c_338_n N_VPWR_c_759_n 0.0133915f $X=3.22 $Y=1.765 $X2=0
+ $Y2=0
cc_287 N_A_114_74#_c_340_n N_VPWR_c_759_n 6.31378e-19 $X=3.67 $Y=1.765 $X2=0
+ $Y2=0
cc_288 N_A_114_74#_c_324_n N_VPWR_c_759_n 0.00454065f $X=2.975 $Y=1.295 $X2=0
+ $Y2=0
cc_289 N_A_114_74#_c_330_n N_VPWR_c_759_n 6.60284e-19 $X=8.39 $Y=1.295 $X2=0
+ $Y2=0
cc_290 N_A_114_74#_c_332_n N_VPWR_c_759_n 4.10401e-19 $X=9.105 $Y=1.355 $X2=0
+ $Y2=0
cc_291 N_A_114_74#_c_338_n N_VPWR_c_760_n 6.39281e-19 $X=3.22 $Y=1.765 $X2=0
+ $Y2=0
cc_292 N_A_114_74#_c_340_n N_VPWR_c_760_n 0.0133415f $X=3.67 $Y=1.765 $X2=0
+ $Y2=0
cc_293 N_A_114_74#_c_342_n N_VPWR_c_760_n 0.0131805f $X=4.12 $Y=1.765 $X2=0
+ $Y2=0
cc_294 N_A_114_74#_c_344_n N_VPWR_c_760_n 6.15498e-19 $X=4.57 $Y=1.765 $X2=0
+ $Y2=0
cc_295 N_A_114_74#_c_325_n N_VPWR_c_760_n 0.00455004f $X=3.835 $Y=1.295 $X2=0
+ $Y2=0
cc_296 N_A_114_74#_c_330_n N_VPWR_c_760_n 6.3322e-19 $X=8.39 $Y=1.295 $X2=0
+ $Y2=0
cc_297 N_A_114_74#_c_332_n N_VPWR_c_760_n 4.08665e-19 $X=9.105 $Y=1.355 $X2=0
+ $Y2=0
cc_298 N_A_114_74#_c_342_n N_VPWR_c_761_n 6.62843e-19 $X=4.12 $Y=1.765 $X2=0
+ $Y2=0
cc_299 N_A_114_74#_c_344_n N_VPWR_c_761_n 0.0136433f $X=4.57 $Y=1.765 $X2=0
+ $Y2=0
cc_300 N_A_114_74#_c_346_n N_VPWR_c_761_n 0.0133915f $X=5.02 $Y=1.765 $X2=0
+ $Y2=0
cc_301 N_A_114_74#_c_348_n N_VPWR_c_761_n 6.31378e-19 $X=5.47 $Y=1.765 $X2=0
+ $Y2=0
cc_302 N_A_114_74#_c_326_n N_VPWR_c_761_n 0.0035092f $X=4.675 $Y=1.295 $X2=0
+ $Y2=0
cc_303 N_A_114_74#_c_330_n N_VPWR_c_761_n 8.68299e-19 $X=8.39 $Y=1.295 $X2=0
+ $Y2=0
cc_304 N_A_114_74#_c_332_n N_VPWR_c_761_n 4.05431e-19 $X=9.105 $Y=1.355 $X2=0
+ $Y2=0
cc_305 N_A_114_74#_c_346_n N_VPWR_c_762_n 6.31378e-19 $X=5.02 $Y=1.765 $X2=0
+ $Y2=0
cc_306 N_A_114_74#_c_348_n N_VPWR_c_762_n 0.0132247f $X=5.47 $Y=1.765 $X2=0
+ $Y2=0
cc_307 N_A_114_74#_c_350_n N_VPWR_c_762_n 0.0133915f $X=5.92 $Y=1.765 $X2=0
+ $Y2=0
cc_308 N_A_114_74#_c_352_n N_VPWR_c_762_n 6.31378e-19 $X=6.37 $Y=1.765 $X2=0
+ $Y2=0
cc_309 N_A_114_74#_c_327_n N_VPWR_c_762_n 0.00378069f $X=5.59 $Y=1.295 $X2=0
+ $Y2=0
cc_310 N_A_114_74#_c_330_n N_VPWR_c_762_n 8.0953e-19 $X=8.39 $Y=1.295 $X2=0
+ $Y2=0
cc_311 N_A_114_74#_c_332_n N_VPWR_c_762_n 4.11269e-19 $X=9.105 $Y=1.355 $X2=0
+ $Y2=0
cc_312 N_A_114_74#_c_350_n N_VPWR_c_763_n 0.00413917f $X=5.92 $Y=1.765 $X2=0
+ $Y2=0
cc_313 N_A_114_74#_c_352_n N_VPWR_c_763_n 0.00413917f $X=6.37 $Y=1.765 $X2=0
+ $Y2=0
cc_314 N_A_114_74#_c_350_n N_VPWR_c_764_n 6.39281e-19 $X=5.92 $Y=1.765 $X2=0
+ $Y2=0
cc_315 N_A_114_74#_c_352_n N_VPWR_c_764_n 0.0133415f $X=6.37 $Y=1.765 $X2=0
+ $Y2=0
cc_316 N_A_114_74#_c_354_n N_VPWR_c_764_n 0.0134974f $X=6.82 $Y=1.765 $X2=0
+ $Y2=0
cc_317 N_A_114_74#_c_356_n N_VPWR_c_764_n 6.39281e-19 $X=7.27 $Y=1.765 $X2=0
+ $Y2=0
cc_318 N_A_114_74#_c_328_n N_VPWR_c_764_n 0.00448005f $X=6.53 $Y=1.295 $X2=0
+ $Y2=0
cc_319 N_A_114_74#_c_330_n N_VPWR_c_764_n 6.5281e-19 $X=8.39 $Y=1.295 $X2=0
+ $Y2=0
cc_320 N_A_114_74#_c_332_n N_VPWR_c_764_n 4.12137e-19 $X=9.105 $Y=1.355 $X2=0
+ $Y2=0
cc_321 N_A_114_74#_c_354_n N_VPWR_c_765_n 6.31378e-19 $X=6.82 $Y=1.765 $X2=0
+ $Y2=0
cc_322 N_A_114_74#_c_356_n N_VPWR_c_765_n 0.0132356f $X=7.27 $Y=1.765 $X2=0
+ $Y2=0
cc_323 N_A_114_74#_c_358_n N_VPWR_c_765_n 0.0133915f $X=7.72 $Y=1.765 $X2=0
+ $Y2=0
cc_324 N_A_114_74#_c_360_n N_VPWR_c_765_n 6.31378e-19 $X=8.17 $Y=1.765 $X2=0
+ $Y2=0
cc_325 N_A_114_74#_c_329_n N_VPWR_c_765_n 0.00489996f $X=7.46 $Y=1.295 $X2=0
+ $Y2=0
cc_326 N_A_114_74#_c_330_n N_VPWR_c_765_n 5.35271e-19 $X=8.39 $Y=1.295 $X2=0
+ $Y2=0
cc_327 N_A_114_74#_c_332_n N_VPWR_c_765_n 4.12137e-19 $X=9.105 $Y=1.355 $X2=0
+ $Y2=0
cc_328 N_A_114_74#_c_358_n N_VPWR_c_766_n 6.31378e-19 $X=7.72 $Y=1.765 $X2=0
+ $Y2=0
cc_329 N_A_114_74#_c_360_n N_VPWR_c_766_n 0.0130897f $X=8.17 $Y=1.765 $X2=0
+ $Y2=0
cc_330 N_A_114_74#_c_362_n N_VPWR_c_766_n 0.00231512f $X=8.64 $Y=1.765 $X2=0
+ $Y2=0
cc_331 N_A_114_74#_c_330_n N_VPWR_c_766_n 3.24741e-19 $X=8.39 $Y=1.295 $X2=0
+ $Y2=0
cc_332 N_A_114_74#_c_331_n N_VPWR_c_766_n 0.00540191f $X=8.39 $Y=1.295 $X2=0
+ $Y2=0
cc_333 N_A_114_74#_c_332_n N_VPWR_c_766_n 5.03723e-19 $X=9.105 $Y=1.355 $X2=0
+ $Y2=0
cc_334 N_A_114_74#_c_362_n N_VPWR_c_768_n 5.9062e-19 $X=8.64 $Y=1.765 $X2=0
+ $Y2=0
cc_335 N_A_114_74#_c_364_n N_VPWR_c_768_n 0.0146808f $X=9.09 $Y=1.765 $X2=0
+ $Y2=0
cc_336 N_A_114_74#_c_365_n N_VPWR_c_769_n 0.014552f $X=0.735 $Y=2.815 $X2=0
+ $Y2=0
cc_337 N_A_114_74#_c_334_n N_VPWR_c_771_n 0.00444681f $X=2.32 $Y=1.765 $X2=0
+ $Y2=0
cc_338 N_A_114_74#_c_336_n N_VPWR_c_771_n 0.00413917f $X=2.77 $Y=1.765 $X2=0
+ $Y2=0
cc_339 N_A_114_74#_c_338_n N_VPWR_c_773_n 0.00413917f $X=3.22 $Y=1.765 $X2=0
+ $Y2=0
cc_340 N_A_114_74#_c_340_n N_VPWR_c_773_n 0.00413917f $X=3.67 $Y=1.765 $X2=0
+ $Y2=0
cc_341 N_A_114_74#_c_342_n N_VPWR_c_775_n 0.00413917f $X=4.12 $Y=1.765 $X2=0
+ $Y2=0
cc_342 N_A_114_74#_c_344_n N_VPWR_c_775_n 0.00413917f $X=4.57 $Y=1.765 $X2=0
+ $Y2=0
cc_343 N_A_114_74#_c_346_n N_VPWR_c_777_n 0.00413917f $X=5.02 $Y=1.765 $X2=0
+ $Y2=0
cc_344 N_A_114_74#_c_348_n N_VPWR_c_777_n 0.00413917f $X=5.47 $Y=1.765 $X2=0
+ $Y2=0
cc_345 N_A_114_74#_c_366_n N_VPWR_c_779_n 0.014552f $X=1.635 $Y=2.815 $X2=0
+ $Y2=0
cc_346 N_A_114_74#_c_354_n N_VPWR_c_780_n 0.00413917f $X=6.82 $Y=1.765 $X2=0
+ $Y2=0
cc_347 N_A_114_74#_c_356_n N_VPWR_c_780_n 0.00413917f $X=7.27 $Y=1.765 $X2=0
+ $Y2=0
cc_348 N_A_114_74#_c_358_n N_VPWR_c_781_n 0.00413917f $X=7.72 $Y=1.765 $X2=0
+ $Y2=0
cc_349 N_A_114_74#_c_360_n N_VPWR_c_781_n 0.00413917f $X=8.17 $Y=1.765 $X2=0
+ $Y2=0
cc_350 N_A_114_74#_c_362_n N_VPWR_c_782_n 0.00461464f $X=8.64 $Y=1.765 $X2=0
+ $Y2=0
cc_351 N_A_114_74#_c_364_n N_VPWR_c_782_n 0.00413917f $X=9.09 $Y=1.765 $X2=0
+ $Y2=0
cc_352 N_A_114_74#_c_334_n N_VPWR_c_754_n 0.00877716f $X=2.32 $Y=1.765 $X2=0
+ $Y2=0
cc_353 N_A_114_74#_c_336_n N_VPWR_c_754_n 0.00817726f $X=2.77 $Y=1.765 $X2=0
+ $Y2=0
cc_354 N_A_114_74#_c_338_n N_VPWR_c_754_n 0.00817726f $X=3.22 $Y=1.765 $X2=0
+ $Y2=0
cc_355 N_A_114_74#_c_340_n N_VPWR_c_754_n 0.00817726f $X=3.67 $Y=1.765 $X2=0
+ $Y2=0
cc_356 N_A_114_74#_c_342_n N_VPWR_c_754_n 0.00817726f $X=4.12 $Y=1.765 $X2=0
+ $Y2=0
cc_357 N_A_114_74#_c_344_n N_VPWR_c_754_n 0.00817726f $X=4.57 $Y=1.765 $X2=0
+ $Y2=0
cc_358 N_A_114_74#_c_346_n N_VPWR_c_754_n 0.00817726f $X=5.02 $Y=1.765 $X2=0
+ $Y2=0
cc_359 N_A_114_74#_c_348_n N_VPWR_c_754_n 0.00817726f $X=5.47 $Y=1.765 $X2=0
+ $Y2=0
cc_360 N_A_114_74#_c_350_n N_VPWR_c_754_n 0.00817726f $X=5.92 $Y=1.765 $X2=0
+ $Y2=0
cc_361 N_A_114_74#_c_352_n N_VPWR_c_754_n 0.00817726f $X=6.37 $Y=1.765 $X2=0
+ $Y2=0
cc_362 N_A_114_74#_c_354_n N_VPWR_c_754_n 0.00817726f $X=6.82 $Y=1.765 $X2=0
+ $Y2=0
cc_363 N_A_114_74#_c_356_n N_VPWR_c_754_n 0.00817726f $X=7.27 $Y=1.765 $X2=0
+ $Y2=0
cc_364 N_A_114_74#_c_358_n N_VPWR_c_754_n 0.00817726f $X=7.72 $Y=1.765 $X2=0
+ $Y2=0
cc_365 N_A_114_74#_c_360_n N_VPWR_c_754_n 0.00817726f $X=8.17 $Y=1.765 $X2=0
+ $Y2=0
cc_366 N_A_114_74#_c_362_n N_VPWR_c_754_n 0.00907797f $X=8.64 $Y=1.765 $X2=0
+ $Y2=0
cc_367 N_A_114_74#_c_364_n N_VPWR_c_754_n 0.00817726f $X=9.09 $Y=1.765 $X2=0
+ $Y2=0
cc_368 N_A_114_74#_c_365_n N_VPWR_c_754_n 0.0119791f $X=0.735 $Y=2.815 $X2=0
+ $Y2=0
cc_369 N_A_114_74#_c_366_n N_VPWR_c_754_n 0.0119791f $X=1.635 $Y=2.815 $X2=0
+ $Y2=0
cc_370 N_A_114_74#_M1003_g N_X_c_946_n 0.00713733f $X=2.305 $Y=0.58 $X2=0 $Y2=0
cc_371 N_A_114_74#_c_285_n N_X_c_946_n 0.00334203f $X=2.32 $Y=1.675 $X2=0 $Y2=0
cc_372 N_A_114_74#_c_334_n N_X_c_946_n 0.00513385f $X=2.32 $Y=1.765 $X2=0 $Y2=0
cc_373 N_A_114_74#_M1005_g N_X_c_946_n 0.00626885f $X=2.735 $Y=0.58 $X2=0 $Y2=0
cc_374 N_A_114_74#_c_287_n N_X_c_946_n 0.00352584f $X=2.77 $Y=1.675 $X2=0 $Y2=0
cc_375 N_A_114_74#_c_336_n N_X_c_946_n 0.00259422f $X=2.77 $Y=1.765 $X2=0 $Y2=0
cc_376 N_A_114_74#_c_321_n N_X_c_946_n 0.0278146f $X=2.05 $Y=1.41 $X2=0 $Y2=0
cc_377 N_A_114_74#_c_322_n N_X_c_946_n 0.0288522f $X=2.05 $Y=1.95 $X2=0 $Y2=0
cc_378 N_A_114_74#_c_408_n N_X_c_946_n 0.00744542f $X=2.05 $Y=2.035 $X2=0 $Y2=0
cc_379 N_A_114_74#_c_324_n N_X_c_946_n 0.0216971f $X=2.975 $Y=1.295 $X2=0 $Y2=0
cc_380 N_A_114_74#_c_330_n N_X_c_946_n 0.0338855f $X=8.39 $Y=1.295 $X2=0 $Y2=0
cc_381 N_A_114_74#_c_332_n N_X_c_946_n 0.0187914f $X=9.105 $Y=1.355 $X2=0 $Y2=0
cc_382 N_A_114_74#_c_334_n N_X_c_956_n 5.0205e-19 $X=2.32 $Y=1.765 $X2=0 $Y2=0
cc_383 N_A_114_74#_c_366_n N_X_c_956_n 0.0020949f $X=1.635 $Y=2.815 $X2=0 $Y2=0
cc_384 N_A_114_74#_c_287_n N_X_c_947_n 3.65363e-19 $X=2.77 $Y=1.675 $X2=0 $Y2=0
cc_385 N_A_114_74#_M1008_g N_X_c_947_n 0.00569263f $X=3.165 $Y=0.58 $X2=0 $Y2=0
cc_386 N_A_114_74#_c_289_n N_X_c_947_n 0.00433879f $X=3.22 $Y=1.675 $X2=0 $Y2=0
cc_387 N_A_114_74#_c_338_n N_X_c_947_n 3.97013e-19 $X=3.22 $Y=1.765 $X2=0 $Y2=0
cc_388 N_A_114_74#_M1010_g N_X_c_947_n 0.00608793f $X=3.595 $Y=0.58 $X2=0 $Y2=0
cc_389 N_A_114_74#_c_291_n N_X_c_947_n 0.00219426f $X=3.67 $Y=1.675 $X2=0 $Y2=0
cc_390 N_A_114_74#_c_324_n N_X_c_947_n 0.0222153f $X=2.975 $Y=1.295 $X2=0 $Y2=0
cc_391 N_A_114_74#_c_325_n N_X_c_947_n 0.0223522f $X=3.835 $Y=1.295 $X2=0 $Y2=0
cc_392 N_A_114_74#_c_330_n N_X_c_947_n 0.0288519f $X=8.39 $Y=1.295 $X2=0 $Y2=0
cc_393 N_A_114_74#_c_332_n N_X_c_947_n 0.0180435f $X=9.105 $Y=1.355 $X2=0 $Y2=0
cc_394 N_A_114_74#_M1013_g N_X_c_948_n 0.00212827f $X=4.455 $Y=0.58 $X2=0 $Y2=0
cc_395 N_A_114_74#_c_295_n N_X_c_948_n 5.68186e-19 $X=4.57 $Y=1.675 $X2=0 $Y2=0
cc_396 N_A_114_74#_M1014_g N_X_c_948_n 0.0154435f $X=4.955 $Y=0.58 $X2=0 $Y2=0
cc_397 N_A_114_74#_c_297_n N_X_c_948_n 0.00454319f $X=5.02 $Y=1.675 $X2=0 $Y2=0
cc_398 N_A_114_74#_c_346_n N_X_c_948_n 4.15716e-19 $X=5.02 $Y=1.765 $X2=0 $Y2=0
cc_399 N_A_114_74#_M1015_g N_X_c_948_n 0.0103156f $X=5.385 $Y=0.58 $X2=0 $Y2=0
cc_400 N_A_114_74#_c_299_n N_X_c_948_n 0.00391785f $X=5.47 $Y=1.675 $X2=0 $Y2=0
cc_401 N_A_114_74#_c_326_n N_X_c_948_n 0.020555f $X=4.675 $Y=1.295 $X2=0 $Y2=0
cc_402 N_A_114_74#_c_327_n N_X_c_948_n 0.0223666f $X=5.59 $Y=1.295 $X2=0 $Y2=0
cc_403 N_A_114_74#_c_330_n N_X_c_948_n 0.0295687f $X=8.39 $Y=1.295 $X2=0 $Y2=0
cc_404 N_A_114_74#_c_332_n N_X_c_948_n 0.0175276f $X=9.105 $Y=1.355 $X2=0 $Y2=0
cc_405 N_A_114_74#_M1015_g N_X_c_949_n 0.00245886f $X=5.385 $Y=0.58 $X2=0 $Y2=0
cc_406 N_A_114_74#_c_299_n N_X_c_949_n 5.56186e-19 $X=5.47 $Y=1.675 $X2=0 $Y2=0
cc_407 N_A_114_74#_M1018_g N_X_c_949_n 0.017286f $X=5.885 $Y=0.58 $X2=0 $Y2=0
cc_408 N_A_114_74#_c_301_n N_X_c_949_n 0.00455914f $X=5.92 $Y=1.675 $X2=0 $Y2=0
cc_409 N_A_114_74#_c_350_n N_X_c_949_n 4.17176e-19 $X=5.92 $Y=1.765 $X2=0 $Y2=0
cc_410 N_A_114_74#_M1019_g N_X_c_949_n 0.0104774f $X=6.315 $Y=0.58 $X2=0 $Y2=0
cc_411 N_A_114_74#_c_303_n N_X_c_949_n 0.00413224f $X=6.37 $Y=1.675 $X2=0 $Y2=0
cc_412 N_A_114_74#_c_327_n N_X_c_949_n 0.0211765f $X=5.59 $Y=1.295 $X2=0 $Y2=0
cc_413 N_A_114_74#_c_328_n N_X_c_949_n 0.0211765f $X=6.53 $Y=1.295 $X2=0 $Y2=0
cc_414 N_A_114_74#_c_330_n N_X_c_949_n 0.0318386f $X=8.39 $Y=1.295 $X2=0 $Y2=0
cc_415 N_A_114_74#_c_332_n N_X_c_949_n 0.018957f $X=9.105 $Y=1.355 $X2=0 $Y2=0
cc_416 N_A_114_74#_M1019_g N_X_c_950_n 0.00245886f $X=6.315 $Y=0.58 $X2=0 $Y2=0
cc_417 N_A_114_74#_c_303_n N_X_c_950_n 5.26607e-19 $X=6.37 $Y=1.675 $X2=0 $Y2=0
cc_418 N_A_114_74#_c_304_n N_X_c_950_n 0.00431332f $X=6.82 $Y=1.675 $X2=0 $Y2=0
cc_419 N_A_114_74#_M1027_g N_X_c_950_n 0.017286f $X=6.815 $Y=0.58 $X2=0 $Y2=0
cc_420 N_A_114_74#_c_354_n N_X_c_950_n 3.94683e-19 $X=6.82 $Y=1.765 $X2=0 $Y2=0
cc_421 N_A_114_74#_M1028_g N_X_c_950_n 0.0104774f $X=7.245 $Y=0.58 $X2=0 $Y2=0
cc_422 N_A_114_74#_c_307_n N_X_c_950_n 0.00429008f $X=7.27 $Y=1.675 $X2=0 $Y2=0
cc_423 N_A_114_74#_c_328_n N_X_c_950_n 0.0224219f $X=6.53 $Y=1.295 $X2=0 $Y2=0
cc_424 N_A_114_74#_c_329_n N_X_c_950_n 0.0211765f $X=7.46 $Y=1.295 $X2=0 $Y2=0
cc_425 N_A_114_74#_c_330_n N_X_c_950_n 0.0317626f $X=8.39 $Y=1.295 $X2=0 $Y2=0
cc_426 N_A_114_74#_c_332_n N_X_c_950_n 0.0189283f $X=9.105 $Y=1.355 $X2=0 $Y2=0
cc_427 N_A_114_74#_M1028_g N_X_c_951_n 0.00245886f $X=7.245 $Y=0.58 $X2=0 $Y2=0
cc_428 N_A_114_74#_c_307_n N_X_c_951_n 4.9893e-19 $X=7.27 $Y=1.675 $X2=0 $Y2=0
cc_429 N_A_114_74#_c_308_n N_X_c_951_n 0.00406073f $X=7.72 $Y=1.675 $X2=0 $Y2=0
cc_430 N_A_114_74#_c_358_n N_X_c_951_n 3.53114e-19 $X=7.72 $Y=1.765 $X2=0 $Y2=0
cc_431 N_A_114_74#_M1031_g N_X_c_951_n 0.017286f $X=7.745 $Y=0.58 $X2=0 $Y2=0
cc_432 N_A_114_74#_c_310_n N_X_c_951_n 0.00445575f $X=8.17 $Y=1.675 $X2=0 $Y2=0
cc_433 N_A_114_74#_M1032_g N_X_c_951_n 0.0104774f $X=8.175 $Y=0.58 $X2=0 $Y2=0
cc_434 N_A_114_74#_c_329_n N_X_c_951_n 0.0224219f $X=7.46 $Y=1.295 $X2=0 $Y2=0
cc_435 N_A_114_74#_c_330_n N_X_c_951_n 0.0318049f $X=8.39 $Y=1.295 $X2=0 $Y2=0
cc_436 N_A_114_74#_c_331_n N_X_c_951_n 0.0211765f $X=8.39 $Y=1.295 $X2=0 $Y2=0
cc_437 N_A_114_74#_c_332_n N_X_c_951_n 0.0189283f $X=9.105 $Y=1.355 $X2=0 $Y2=0
cc_438 N_A_114_74#_c_362_n N_X_c_962_n 0.0029347f $X=8.64 $Y=1.765 $X2=0 $Y2=0
cc_439 N_A_114_74#_c_364_n N_X_c_962_n 0.00356881f $X=9.09 $Y=1.765 $X2=0 $Y2=0
cc_440 N_A_114_74#_c_310_n N_X_c_952_n 8.05453e-19 $X=8.17 $Y=1.675 $X2=0 $Y2=0
cc_441 N_A_114_74#_M1032_g N_X_c_952_n 0.00242366f $X=8.175 $Y=0.58 $X2=0 $Y2=0
cc_442 N_A_114_74#_c_312_n N_X_c_952_n 0.00401977f $X=8.64 $Y=1.675 $X2=0 $Y2=0
cc_443 N_A_114_74#_c_362_n N_X_c_952_n 7.80255e-19 $X=8.64 $Y=1.765 $X2=0 $Y2=0
cc_444 N_A_114_74#_M1037_g N_X_c_952_n 0.0171618f $X=8.675 $Y=0.58 $X2=0 $Y2=0
cc_445 N_A_114_74#_c_314_n N_X_c_952_n 0.00491374f $X=9.09 $Y=1.675 $X2=0 $Y2=0
cc_446 N_A_114_74#_M1039_g N_X_c_952_n 0.0105222f $X=9.105 $Y=0.58 $X2=0 $Y2=0
cc_447 N_A_114_74#_c_330_n N_X_c_952_n 0.00755956f $X=8.39 $Y=1.295 $X2=0 $Y2=0
cc_448 N_A_114_74#_c_331_n N_X_c_952_n 0.0214654f $X=8.39 $Y=1.295 $X2=0 $Y2=0
cc_449 N_A_114_74#_c_332_n N_X_c_952_n 0.0303236f $X=9.105 $Y=1.355 $X2=0 $Y2=0
cc_450 N_A_114_74#_c_336_n N_X_c_964_n 6.50844e-19 $X=2.77 $Y=1.765 $X2=0 $Y2=0
cc_451 N_A_114_74#_c_338_n N_X_c_964_n 0.0052228f $X=3.22 $Y=1.765 $X2=0 $Y2=0
cc_452 N_A_114_74#_c_340_n N_X_c_964_n 0.00357375f $X=3.67 $Y=1.765 $X2=0 $Y2=0
cc_453 N_A_114_74#_c_330_n N_X_c_964_n 0.00144258f $X=8.39 $Y=1.295 $X2=0 $Y2=0
cc_454 N_A_114_74#_M1012_g N_X_c_953_n 0.00533114f $X=4.025 $Y=0.58 $X2=0 $Y2=0
cc_455 N_A_114_74#_M1013_g N_X_c_953_n 0.00995023f $X=4.455 $Y=0.58 $X2=0 $Y2=0
cc_456 N_A_114_74#_c_330_n N_X_c_953_n 0.00355816f $X=8.39 $Y=1.295 $X2=0 $Y2=0
cc_457 N_A_114_74#_c_291_n N_X_c_954_n 3.75323e-19 $X=3.67 $Y=1.675 $X2=0 $Y2=0
cc_458 N_A_114_74#_M1012_g N_X_c_954_n 0.00547607f $X=4.025 $Y=0.58 $X2=0 $Y2=0
cc_459 N_A_114_74#_c_293_n N_X_c_954_n 0.00428916f $X=4.12 $Y=1.675 $X2=0 $Y2=0
cc_460 N_A_114_74#_c_342_n N_X_c_954_n 3.92472e-19 $X=4.12 $Y=1.765 $X2=0 $Y2=0
cc_461 N_A_114_74#_c_295_n N_X_c_954_n 0.00362785f $X=4.57 $Y=1.675 $X2=0 $Y2=0
cc_462 N_A_114_74#_c_325_n N_X_c_954_n 0.0221713f $X=3.835 $Y=1.295 $X2=0 $Y2=0
cc_463 N_A_114_74#_c_326_n N_X_c_954_n 0.0221713f $X=4.675 $Y=1.295 $X2=0 $Y2=0
cc_464 N_A_114_74#_c_330_n N_X_c_954_n 0.0229117f $X=8.39 $Y=1.295 $X2=0 $Y2=0
cc_465 N_A_114_74#_c_332_n N_X_c_954_n 0.0150486f $X=9.105 $Y=1.355 $X2=0 $Y2=0
cc_466 N_A_114_74#_c_340_n N_X_c_966_n 6.6474e-19 $X=3.67 $Y=1.765 $X2=0 $Y2=0
cc_467 N_A_114_74#_c_342_n N_X_c_966_n 0.00534703f $X=4.12 $Y=1.765 $X2=0 $Y2=0
cc_468 N_A_114_74#_c_344_n N_X_c_966_n 0.00853484f $X=4.57 $Y=1.765 $X2=0 $Y2=0
cc_469 N_A_114_74#_c_330_n N_X_c_966_n 0.00291795f $X=8.39 $Y=1.295 $X2=0 $Y2=0
cc_470 N_A_114_74#_c_332_n N_X_c_966_n 0.00241927f $X=9.105 $Y=1.355 $X2=0 $Y2=0
cc_471 N_A_114_74#_c_344_n N_X_c_967_n 8.80793e-19 $X=4.57 $Y=1.765 $X2=0 $Y2=0
cc_472 N_A_114_74#_c_346_n N_X_c_967_n 0.00660033f $X=5.02 $Y=1.765 $X2=0 $Y2=0
cc_473 N_A_114_74#_c_348_n N_X_c_967_n 0.00359744f $X=5.47 $Y=1.765 $X2=0 $Y2=0
cc_474 N_A_114_74#_c_330_n N_X_c_967_n 0.00308188f $X=8.39 $Y=1.295 $X2=0 $Y2=0
cc_475 N_A_114_74#_c_332_n N_X_c_967_n 0.00169349f $X=9.105 $Y=1.355 $X2=0 $Y2=0
cc_476 N_A_114_74#_c_348_n N_X_c_968_n 8.61484e-19 $X=5.47 $Y=1.765 $X2=0 $Y2=0
cc_477 N_A_114_74#_c_350_n N_X_c_968_n 0.00627939f $X=5.92 $Y=1.765 $X2=0 $Y2=0
cc_478 N_A_114_74#_c_352_n N_X_c_968_n 0.00361089f $X=6.37 $Y=1.765 $X2=0 $Y2=0
cc_479 N_A_114_74#_c_330_n N_X_c_968_n 0.00193437f $X=8.39 $Y=1.295 $X2=0 $Y2=0
cc_480 N_A_114_74#_c_332_n N_X_c_968_n 2.41927e-19 $X=9.105 $Y=1.355 $X2=0 $Y2=0
cc_481 N_A_114_74#_c_352_n N_X_c_969_n 8.18167e-19 $X=6.37 $Y=1.765 $X2=0 $Y2=0
cc_482 N_A_114_74#_c_354_n N_X_c_969_n 0.00553316f $X=6.82 $Y=1.765 $X2=0 $Y2=0
cc_483 N_A_114_74#_c_356_n N_X_c_969_n 0.00365581f $X=7.27 $Y=1.765 $X2=0 $Y2=0
cc_484 N_A_114_74#_c_330_n N_X_c_969_n 0.00111472f $X=8.39 $Y=1.295 $X2=0 $Y2=0
cc_485 N_A_114_74#_c_356_n N_X_c_970_n 4.9893e-19 $X=7.27 $Y=1.765 $X2=0 $Y2=0
cc_486 N_A_114_74#_c_358_n N_X_c_970_n 0.00349903f $X=7.72 $Y=1.765 $X2=0 $Y2=0
cc_487 N_A_114_74#_c_360_n N_X_c_970_n 0.00366932f $X=8.17 $Y=1.765 $X2=0 $Y2=0
cc_488 N_A_114_74#_c_338_n N_X_c_971_n 0.00149334f $X=3.22 $Y=1.765 $X2=0 $Y2=0
cc_489 N_A_114_74#_c_342_n N_X_c_972_n 0.00150774f $X=4.12 $Y=1.765 $X2=0 $Y2=0
cc_490 N_A_114_74#_c_346_n N_X_c_973_n 0.00149701f $X=5.02 $Y=1.765 $X2=0 $Y2=0
cc_491 N_A_114_74#_c_350_n N_X_c_974_n 0.00149334f $X=5.92 $Y=1.765 $X2=0 $Y2=0
cc_492 N_A_114_74#_c_354_n N_X_c_975_n 0.00148425f $X=6.82 $Y=1.765 $X2=0 $Y2=0
cc_493 N_A_114_74#_c_358_n N_X_c_976_n 0.00149701f $X=7.72 $Y=1.765 $X2=0 $Y2=0
cc_494 N_A_114_74#_c_362_n N_X_c_977_n 0.00154509f $X=8.64 $Y=1.765 $X2=0 $Y2=0
cc_495 N_A_114_74#_c_364_n N_X_c_977_n 0.00150412f $X=9.09 $Y=1.765 $X2=0 $Y2=0
cc_496 N_A_114_74#_c_334_n N_X_c_1105_n 0.00232795f $X=2.32 $Y=1.765 $X2=0 $Y2=0
cc_497 N_A_114_74#_c_336_n N_X_c_1105_n 0.00883571f $X=2.77 $Y=1.765 $X2=0 $Y2=0
cc_498 N_A_114_74#_c_338_n N_X_c_1105_n 0.00842306f $X=3.22 $Y=1.765 $X2=0 $Y2=0
cc_499 N_A_114_74#_c_340_n N_X_c_1105_n 0.00850408f $X=3.67 $Y=1.765 $X2=0 $Y2=0
cc_500 N_A_114_74#_c_342_n N_X_c_1105_n 0.00838023f $X=4.12 $Y=1.765 $X2=0 $Y2=0
cc_501 N_A_114_74#_c_344_n N_X_c_1105_n 0.00820054f $X=4.57 $Y=1.765 $X2=0 $Y2=0
cc_502 N_A_114_74#_c_346_n N_X_c_1105_n 0.00803959f $X=5.02 $Y=1.765 $X2=0 $Y2=0
cc_503 N_A_114_74#_c_348_n N_X_c_1105_n 0.00825583f $X=5.47 $Y=1.765 $X2=0 $Y2=0
cc_504 N_A_114_74#_c_350_n N_X_c_1105_n 0.00811628f $X=5.92 $Y=1.765 $X2=0 $Y2=0
cc_505 N_A_114_74#_c_352_n N_X_c_1105_n 0.00847805f $X=6.37 $Y=1.765 $X2=0 $Y2=0
cc_506 N_A_114_74#_c_354_n N_X_c_1105_n 0.00834861f $X=6.82 $Y=1.765 $X2=0 $Y2=0
cc_507 N_A_114_74#_c_356_n N_X_c_1105_n 0.00863197f $X=7.27 $Y=1.765 $X2=0 $Y2=0
cc_508 N_A_114_74#_c_358_n N_X_c_1105_n 0.00856111f $X=7.72 $Y=1.765 $X2=0 $Y2=0
cc_509 N_A_114_74#_c_360_n N_X_c_1105_n 0.00878814f $X=8.17 $Y=1.765 $X2=0 $Y2=0
cc_510 N_A_114_74#_c_362_n N_X_c_1105_n 0.0113911f $X=8.64 $Y=1.765 $X2=0 $Y2=0
cc_511 N_A_114_74#_c_364_n N_X_c_1105_n 0.0123353f $X=9.09 $Y=1.765 $X2=0 $Y2=0
cc_512 N_A_114_74#_c_366_n N_X_c_1105_n 6.20324e-19 $X=1.635 $Y=2.815 $X2=0
+ $Y2=0
cc_513 N_A_114_74#_c_322_n N_X_c_1105_n 8.22299e-19 $X=2.05 $Y=1.95 $X2=0 $Y2=0
cc_514 N_A_114_74#_c_408_n N_X_c_1105_n 0.00479786f $X=2.05 $Y=2.035 $X2=0 $Y2=0
cc_515 N_A_114_74#_c_324_n N_X_c_1105_n 0.00274866f $X=2.975 $Y=1.295 $X2=0
+ $Y2=0
cc_516 N_A_114_74#_c_325_n N_X_c_1105_n 0.0040494f $X=3.835 $Y=1.295 $X2=0 $Y2=0
cc_517 N_A_114_74#_c_326_n N_X_c_1105_n 0.0047356f $X=4.675 $Y=1.295 $X2=0 $Y2=0
cc_518 N_A_114_74#_c_327_n N_X_c_1105_n 0.00456405f $X=5.59 $Y=1.295 $X2=0 $Y2=0
cc_519 N_A_114_74#_c_328_n N_X_c_1105_n 0.00410658f $X=6.53 $Y=1.295 $X2=0 $Y2=0
cc_520 N_A_114_74#_c_329_n N_X_c_1105_n 0.00376348f $X=7.46 $Y=1.295 $X2=0 $Y2=0
cc_521 N_A_114_74#_c_330_n N_X_c_1105_n 0.294859f $X=8.39 $Y=1.295 $X2=0 $Y2=0
cc_522 N_A_114_74#_c_331_n N_X_c_1105_n 0.00342038f $X=8.39 $Y=1.295 $X2=0 $Y2=0
cc_523 N_A_114_74#_c_334_n N_X_c_1132_n 9.40403e-19 $X=2.32 $Y=1.765 $X2=0 $Y2=0
cc_524 N_A_114_74#_c_316_n N_VGND_c_1213_n 0.0172562f $X=0.71 $Y=0.58 $X2=0
+ $Y2=0
cc_525 N_A_114_74#_c_316_n N_VGND_c_1214_n 0.0172562f $X=0.71 $Y=0.58 $X2=0
+ $Y2=0
cc_526 N_A_114_74#_c_317_n N_VGND_c_1214_n 0.0207473f $X=1.425 $Y=1.065 $X2=0
+ $Y2=0
cc_527 N_A_114_74#_c_319_n N_VGND_c_1214_n 0.0302714f $X=1.59 $Y=0.58 $X2=0
+ $Y2=0
cc_528 N_A_114_74#_M1003_g N_VGND_c_1215_n 0.00564006f $X=2.305 $Y=0.58 $X2=0
+ $Y2=0
cc_529 N_A_114_74#_c_319_n N_VGND_c_1215_n 0.0179429f $X=1.59 $Y=0.58 $X2=0
+ $Y2=0
cc_530 N_A_114_74#_c_320_n N_VGND_c_1215_n 0.00884164f $X=1.965 $Y=1.065 $X2=0
+ $Y2=0
cc_531 N_A_114_74#_c_321_n N_VGND_c_1215_n 0.0167244f $X=2.05 $Y=1.41 $X2=0
+ $Y2=0
cc_532 N_A_114_74#_c_330_n N_VGND_c_1215_n 0.00132171f $X=8.39 $Y=1.295 $X2=0
+ $Y2=0
cc_533 N_A_114_74#_M1005_g N_VGND_c_1216_n 0.00275427f $X=2.735 $Y=0.58 $X2=0
+ $Y2=0
cc_534 N_A_114_74#_M1008_g N_VGND_c_1216_n 0.0015425f $X=3.165 $Y=0.58 $X2=0
+ $Y2=0
cc_535 N_A_114_74#_c_324_n N_VGND_c_1216_n 0.00321205f $X=2.975 $Y=1.295 $X2=0
+ $Y2=0
cc_536 N_A_114_74#_c_330_n N_VGND_c_1216_n 0.00397428f $X=8.39 $Y=1.295 $X2=0
+ $Y2=0
cc_537 N_A_114_74#_c_332_n N_VGND_c_1216_n 6.62917e-19 $X=9.105 $Y=1.355 $X2=0
+ $Y2=0
cc_538 N_A_114_74#_M1010_g N_VGND_c_1217_n 0.00176998f $X=3.595 $Y=0.58 $X2=0
+ $Y2=0
cc_539 N_A_114_74#_M1012_g N_VGND_c_1217_n 0.00156717f $X=4.025 $Y=0.58 $X2=0
+ $Y2=0
cc_540 N_A_114_74#_c_325_n N_VGND_c_1217_n 0.00411715f $X=3.835 $Y=1.295 $X2=0
+ $Y2=0
cc_541 N_A_114_74#_c_330_n N_VGND_c_1217_n 0.00544071f $X=8.39 $Y=1.295 $X2=0
+ $Y2=0
cc_542 N_A_114_74#_c_332_n N_VGND_c_1217_n 6.77384e-19 $X=9.105 $Y=1.355 $X2=0
+ $Y2=0
cc_543 N_A_114_74#_M1012_g N_VGND_c_1218_n 0.00434272f $X=4.025 $Y=0.58 $X2=0
+ $Y2=0
cc_544 N_A_114_74#_M1013_g N_VGND_c_1218_n 0.00398535f $X=4.455 $Y=0.58 $X2=0
+ $Y2=0
cc_545 N_A_114_74#_M1012_g N_VGND_c_1219_n 4.58529e-19 $X=4.025 $Y=0.58 $X2=0
+ $Y2=0
cc_546 N_A_114_74#_M1013_g N_VGND_c_1219_n 0.0083302f $X=4.455 $Y=0.58 $X2=0
+ $Y2=0
cc_547 N_A_114_74#_M1014_g N_VGND_c_1219_n 0.00372052f $X=4.955 $Y=0.58 $X2=0
+ $Y2=0
cc_548 N_A_114_74#_c_326_n N_VGND_c_1219_n 0.00638102f $X=4.675 $Y=1.295 $X2=0
+ $Y2=0
cc_549 N_A_114_74#_c_330_n N_VGND_c_1219_n 0.00786623f $X=8.39 $Y=1.295 $X2=0
+ $Y2=0
cc_550 N_A_114_74#_c_332_n N_VGND_c_1219_n 0.00116186f $X=9.105 $Y=1.355 $X2=0
+ $Y2=0
cc_551 N_A_114_74#_M1014_g N_VGND_c_1220_n 4.49641e-19 $X=4.955 $Y=0.58 $X2=0
+ $Y2=0
cc_552 N_A_114_74#_M1015_g N_VGND_c_1220_n 0.00807893f $X=5.385 $Y=0.58 $X2=0
+ $Y2=0
cc_553 N_A_114_74#_M1018_g N_VGND_c_1220_n 0.0034049f $X=5.885 $Y=0.58 $X2=0
+ $Y2=0
cc_554 N_A_114_74#_c_327_n N_VGND_c_1220_n 0.00539651f $X=5.59 $Y=1.295 $X2=0
+ $Y2=0
cc_555 N_A_114_74#_c_330_n N_VGND_c_1220_n 0.00782376f $X=8.39 $Y=1.295 $X2=0
+ $Y2=0
cc_556 N_A_114_74#_c_332_n N_VGND_c_1220_n 0.00112643f $X=9.105 $Y=1.355 $X2=0
+ $Y2=0
cc_557 N_A_114_74#_M1018_g N_VGND_c_1221_n 4.49641e-19 $X=5.885 $Y=0.58 $X2=0
+ $Y2=0
cc_558 N_A_114_74#_M1019_g N_VGND_c_1221_n 0.00807893f $X=6.315 $Y=0.58 $X2=0
+ $Y2=0
cc_559 N_A_114_74#_M1027_g N_VGND_c_1221_n 0.0034049f $X=6.815 $Y=0.58 $X2=0
+ $Y2=0
cc_560 N_A_114_74#_c_328_n N_VGND_c_1221_n 0.00547196f $X=6.53 $Y=1.295 $X2=0
+ $Y2=0
cc_561 N_A_114_74#_c_330_n N_VGND_c_1221_n 0.00766033f $X=8.39 $Y=1.295 $X2=0
+ $Y2=0
cc_562 N_A_114_74#_c_332_n N_VGND_c_1221_n 0.00112718f $X=9.105 $Y=1.355 $X2=0
+ $Y2=0
cc_563 N_A_114_74#_M1027_g N_VGND_c_1222_n 4.49641e-19 $X=6.815 $Y=0.58 $X2=0
+ $Y2=0
cc_564 N_A_114_74#_M1028_g N_VGND_c_1222_n 0.00807893f $X=7.245 $Y=0.58 $X2=0
+ $Y2=0
cc_565 N_A_114_74#_M1031_g N_VGND_c_1222_n 0.0034049f $X=7.745 $Y=0.58 $X2=0
+ $Y2=0
cc_566 N_A_114_74#_c_329_n N_VGND_c_1222_n 0.00547196f $X=7.46 $Y=1.295 $X2=0
+ $Y2=0
cc_567 N_A_114_74#_c_330_n N_VGND_c_1222_n 0.00766033f $X=8.39 $Y=1.295 $X2=0
+ $Y2=0
cc_568 N_A_114_74#_c_332_n N_VGND_c_1222_n 0.00112718f $X=9.105 $Y=1.355 $X2=0
+ $Y2=0
cc_569 N_A_114_74#_M1031_g N_VGND_c_1223_n 4.49641e-19 $X=7.745 $Y=0.58 $X2=0
+ $Y2=0
cc_570 N_A_114_74#_M1032_g N_VGND_c_1223_n 0.00807893f $X=8.175 $Y=0.58 $X2=0
+ $Y2=0
cc_571 N_A_114_74#_M1037_g N_VGND_c_1223_n 0.0034049f $X=8.675 $Y=0.58 $X2=0
+ $Y2=0
cc_572 N_A_114_74#_c_330_n N_VGND_c_1223_n 0.00766033f $X=8.39 $Y=1.295 $X2=0
+ $Y2=0
cc_573 N_A_114_74#_c_331_n N_VGND_c_1223_n 0.00547196f $X=8.39 $Y=1.295 $X2=0
+ $Y2=0
cc_574 N_A_114_74#_c_332_n N_VGND_c_1223_n 0.00112804f $X=9.105 $Y=1.355 $X2=0
+ $Y2=0
cc_575 N_A_114_74#_M1037_g N_VGND_c_1225_n 4.69038e-19 $X=8.675 $Y=0.58 $X2=0
+ $Y2=0
cc_576 N_A_114_74#_M1039_g N_VGND_c_1225_n 0.010727f $X=9.105 $Y=0.58 $X2=0
+ $Y2=0
cc_577 N_A_114_74#_c_316_n N_VGND_c_1226_n 0.0109942f $X=0.71 $Y=0.58 $X2=0
+ $Y2=0
cc_578 N_A_114_74#_c_319_n N_VGND_c_1228_n 0.0109942f $X=1.59 $Y=0.58 $X2=0
+ $Y2=0
cc_579 N_A_114_74#_M1003_g N_VGND_c_1230_n 0.00461464f $X=2.305 $Y=0.58 $X2=0
+ $Y2=0
cc_580 N_A_114_74#_M1005_g N_VGND_c_1230_n 0.00461464f $X=2.735 $Y=0.58 $X2=0
+ $Y2=0
cc_581 N_A_114_74#_M1008_g N_VGND_c_1232_n 0.00461464f $X=3.165 $Y=0.58 $X2=0
+ $Y2=0
cc_582 N_A_114_74#_M1010_g N_VGND_c_1232_n 0.00460063f $X=3.595 $Y=0.58 $X2=0
+ $Y2=0
cc_583 N_A_114_74#_M1014_g N_VGND_c_1234_n 0.00456932f $X=4.955 $Y=0.58 $X2=0
+ $Y2=0
cc_584 N_A_114_74#_M1015_g N_VGND_c_1234_n 0.00383152f $X=5.385 $Y=0.58 $X2=0
+ $Y2=0
cc_585 N_A_114_74#_M1018_g N_VGND_c_1235_n 0.00434272f $X=5.885 $Y=0.58 $X2=0
+ $Y2=0
cc_586 N_A_114_74#_M1019_g N_VGND_c_1235_n 0.00383152f $X=6.315 $Y=0.58 $X2=0
+ $Y2=0
cc_587 N_A_114_74#_M1027_g N_VGND_c_1236_n 0.00434272f $X=6.815 $Y=0.58 $X2=0
+ $Y2=0
cc_588 N_A_114_74#_M1028_g N_VGND_c_1236_n 0.00383152f $X=7.245 $Y=0.58 $X2=0
+ $Y2=0
cc_589 N_A_114_74#_M1031_g N_VGND_c_1237_n 0.00434272f $X=7.745 $Y=0.58 $X2=0
+ $Y2=0
cc_590 N_A_114_74#_M1032_g N_VGND_c_1237_n 0.00383152f $X=8.175 $Y=0.58 $X2=0
+ $Y2=0
cc_591 N_A_114_74#_M1037_g N_VGND_c_1238_n 0.00434272f $X=8.675 $Y=0.58 $X2=0
+ $Y2=0
cc_592 N_A_114_74#_M1039_g N_VGND_c_1238_n 0.00383152f $X=9.105 $Y=0.58 $X2=0
+ $Y2=0
cc_593 N_A_114_74#_M1003_g N_VGND_c_1244_n 0.0090882f $X=2.305 $Y=0.58 $X2=0
+ $Y2=0
cc_594 N_A_114_74#_M1005_g N_VGND_c_1244_n 0.00908333f $X=2.735 $Y=0.58 $X2=0
+ $Y2=0
cc_595 N_A_114_74#_M1008_g N_VGND_c_1244_n 0.00908333f $X=3.165 $Y=0.58 $X2=0
+ $Y2=0
cc_596 N_A_114_74#_M1010_g N_VGND_c_1244_n 0.009071f $X=3.595 $Y=0.58 $X2=0
+ $Y2=0
cc_597 N_A_114_74#_M1012_g N_VGND_c_1244_n 0.00820284f $X=4.025 $Y=0.58 $X2=0
+ $Y2=0
cc_598 N_A_114_74#_M1013_g N_VGND_c_1244_n 0.00787535f $X=4.455 $Y=0.58 $X2=0
+ $Y2=0
cc_599 N_A_114_74#_M1014_g N_VGND_c_1244_n 0.00890307f $X=4.955 $Y=0.58 $X2=0
+ $Y2=0
cc_600 N_A_114_74#_M1015_g N_VGND_c_1244_n 0.0075754f $X=5.385 $Y=0.58 $X2=0
+ $Y2=0
cc_601 N_A_114_74#_M1018_g N_VGND_c_1244_n 0.00820718f $X=5.885 $Y=0.58 $X2=0
+ $Y2=0
cc_602 N_A_114_74#_M1019_g N_VGND_c_1244_n 0.0075754f $X=6.315 $Y=0.58 $X2=0
+ $Y2=0
cc_603 N_A_114_74#_M1027_g N_VGND_c_1244_n 0.00820718f $X=6.815 $Y=0.58 $X2=0
+ $Y2=0
cc_604 N_A_114_74#_M1028_g N_VGND_c_1244_n 0.0075754f $X=7.245 $Y=0.58 $X2=0
+ $Y2=0
cc_605 N_A_114_74#_M1031_g N_VGND_c_1244_n 0.00820718f $X=7.745 $Y=0.58 $X2=0
+ $Y2=0
cc_606 N_A_114_74#_M1032_g N_VGND_c_1244_n 0.0075754f $X=8.175 $Y=0.58 $X2=0
+ $Y2=0
cc_607 N_A_114_74#_M1037_g N_VGND_c_1244_n 0.00820718f $X=8.675 $Y=0.58 $X2=0
+ $Y2=0
cc_608 N_A_114_74#_M1039_g N_VGND_c_1244_n 0.0075754f $X=9.105 $Y=0.58 $X2=0
+ $Y2=0
cc_609 N_A_114_74#_c_316_n N_VGND_c_1244_n 0.00904371f $X=0.71 $Y=0.58 $X2=0
+ $Y2=0
cc_610 N_A_114_74#_c_319_n N_VGND_c_1244_n 0.00904371f $X=1.59 $Y=0.58 $X2=0
+ $Y2=0
cc_611 N_VPWR_c_758_n N_X_c_956_n 0.0244192f $X=2.085 $Y=2.455 $X2=0 $Y2=0
cc_612 N_VPWR_c_771_n N_X_c_956_n 0.0101736f $X=2.83 $Y=3.33 $X2=0 $Y2=0
cc_613 N_VPWR_c_754_n N_X_c_956_n 0.0084208f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_614 N_VPWR_c_759_n N_X_c_971_n 0.0361395f $X=2.995 $Y=2.115 $X2=0 $Y2=0
cc_615 N_VPWR_c_760_n N_X_c_971_n 0.0353169f $X=3.895 $Y=2.115 $X2=0 $Y2=0
cc_616 N_VPWR_c_773_n N_X_c_971_n 0.00905805f $X=3.73 $Y=3.33 $X2=0 $Y2=0
cc_617 N_VPWR_c_754_n N_X_c_971_n 0.00749747f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_618 N_VPWR_c_760_n N_X_c_972_n 0.0379186f $X=3.895 $Y=2.115 $X2=0 $Y2=0
cc_619 N_VPWR_c_761_n N_X_c_972_n 0.0615238f $X=4.795 $Y=2.115 $X2=0 $Y2=0
cc_620 N_VPWR_c_775_n N_X_c_972_n 0.00883494f $X=4.63 $Y=3.33 $X2=0 $Y2=0
cc_621 N_VPWR_c_754_n N_X_c_972_n 0.0073128f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_622 N_VPWR_c_761_n N_X_c_973_n 0.0361436f $X=4.795 $Y=2.115 $X2=0 $Y2=0
cc_623 N_VPWR_c_762_n N_X_c_973_n 0.0361436f $X=5.695 $Y=2.115 $X2=0 $Y2=0
cc_624 N_VPWR_c_777_n N_X_c_973_n 0.00928115f $X=5.53 $Y=3.33 $X2=0 $Y2=0
cc_625 N_VPWR_c_754_n N_X_c_973_n 0.00768213f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_626 N_VPWR_c_762_n N_X_c_974_n 0.0361395f $X=5.695 $Y=2.115 $X2=0 $Y2=0
cc_627 N_VPWR_c_763_n N_X_c_974_n 0.00905805f $X=6.43 $Y=3.33 $X2=0 $Y2=0
cc_628 N_VPWR_c_764_n N_X_c_974_n 0.0353169f $X=6.595 $Y=2.115 $X2=0 $Y2=0
cc_629 N_VPWR_c_754_n N_X_c_974_n 0.00749747f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_630 N_VPWR_c_764_n N_X_c_975_n 0.0353169f $X=6.595 $Y=2.115 $X2=0 $Y2=0
cc_631 N_VPWR_c_765_n N_X_c_975_n 0.0361395f $X=7.495 $Y=2.115 $X2=0 $Y2=0
cc_632 N_VPWR_c_780_n N_X_c_975_n 0.00905805f $X=7.33 $Y=3.33 $X2=0 $Y2=0
cc_633 N_VPWR_c_754_n N_X_c_975_n 0.00749747f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_634 N_VPWR_c_765_n N_X_c_976_n 0.0361436f $X=7.495 $Y=2.115 $X2=0 $Y2=0
cc_635 N_VPWR_c_766_n N_X_c_976_n 0.0361436f $X=8.395 $Y=2.115 $X2=0 $Y2=0
cc_636 N_VPWR_c_781_n N_X_c_976_n 0.00928115f $X=8.23 $Y=3.33 $X2=0 $Y2=0
cc_637 N_VPWR_c_754_n N_X_c_976_n 0.00768213f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_638 N_VPWR_c_766_n N_X_c_977_n 0.00526404f $X=8.395 $Y=2.115 $X2=0 $Y2=0
cc_639 N_VPWR_c_768_n N_X_c_977_n 0.0357471f $X=9.315 $Y=2.115 $X2=0 $Y2=0
cc_640 N_VPWR_c_782_n N_X_c_977_n 0.00972736f $X=9.15 $Y=3.33 $X2=0 $Y2=0
cc_641 N_VPWR_c_754_n N_X_c_977_n 0.00805147f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_642 N_VPWR_M1001_s N_X_c_1105_n 0.00271617f $X=2.845 $Y=1.84 $X2=0 $Y2=0
cc_643 N_VPWR_M1004_s N_X_c_1105_n 0.00274277f $X=3.745 $Y=1.84 $X2=0 $Y2=0
cc_644 N_VPWR_M1007_s N_X_c_1105_n 0.0030481f $X=4.645 $Y=1.84 $X2=0 $Y2=0
cc_645 N_VPWR_M1011_s N_X_c_1105_n 0.00298216f $X=5.545 $Y=1.84 $X2=0 $Y2=0
cc_646 N_VPWR_M1017_s N_X_c_1105_n 0.00276937f $X=6.445 $Y=1.84 $X2=0 $Y2=0
cc_647 N_VPWR_M1024_s N_X_c_1105_n 0.00260978f $X=7.345 $Y=1.84 $X2=0 $Y2=0
cc_648 N_VPWR_M1033_s N_X_c_1105_n 0.00270414f $X=8.245 $Y=1.84 $X2=0 $Y2=0
cc_649 N_VPWR_c_759_n N_X_c_1105_n 0.029332f $X=2.995 $Y=2.115 $X2=0 $Y2=0
cc_650 N_VPWR_c_760_n N_X_c_1105_n 0.0294061f $X=3.895 $Y=2.115 $X2=0 $Y2=0
cc_651 N_VPWR_c_761_n N_X_c_1105_n 0.0302679f $X=4.795 $Y=2.115 $X2=0 $Y2=0
cc_652 N_VPWR_c_762_n N_X_c_1105_n 0.0299699f $X=5.695 $Y=2.115 $X2=0 $Y2=0
cc_653 N_VPWR_c_764_n N_X_c_1105_n 0.0295568f $X=6.595 $Y=2.115 $X2=0 $Y2=0
cc_654 N_VPWR_c_765_n N_X_c_1105_n 0.0291491f $X=7.495 $Y=2.115 $X2=0 $Y2=0
cc_655 N_VPWR_c_766_n N_X_c_1105_n 0.0290535f $X=8.395 $Y=2.115 $X2=0 $Y2=0
cc_656 N_VPWR_c_768_n N_X_c_1105_n 0.00404225f $X=9.315 $Y=2.115 $X2=0 $Y2=0
cc_657 N_VPWR_c_759_n N_X_c_1132_n 0.037934f $X=2.995 $Y=2.115 $X2=0 $Y2=0
cc_658 N_X_c_946_n N_VGND_c_1215_n 0.00273037f $X=2.52 $Y=0.58 $X2=0 $Y2=0
cc_659 N_X_c_946_n N_VGND_c_1216_n 0.0117358f $X=2.52 $Y=0.58 $X2=0 $Y2=0
cc_660 N_X_c_947_n N_VGND_c_1216_n 0.00114748f $X=3.38 $Y=0.58 $X2=0 $Y2=0
cc_661 N_X_c_947_n N_VGND_c_1217_n 0.0154288f $X=3.38 $Y=0.58 $X2=0 $Y2=0
cc_662 N_X_c_953_n N_VGND_c_1217_n 0.0137127f $X=4.24 $Y=0.58 $X2=0 $Y2=0
cc_663 N_X_c_953_n N_VGND_c_1218_n 0.0115088f $X=4.24 $Y=0.58 $X2=0 $Y2=0
cc_664 N_X_c_948_n N_VGND_c_1219_n 0.0133947f $X=5.17 $Y=0.58 $X2=0 $Y2=0
cc_665 N_X_c_953_n N_VGND_c_1219_n 0.0153642f $X=4.24 $Y=0.58 $X2=0 $Y2=0
cc_666 N_X_c_948_n N_VGND_c_1220_n 0.0125465f $X=5.17 $Y=0.58 $X2=0 $Y2=0
cc_667 N_X_c_949_n N_VGND_c_1220_n 0.0126571f $X=6.1 $Y=0.58 $X2=0 $Y2=0
cc_668 N_X_c_949_n N_VGND_c_1221_n 0.0125556f $X=6.1 $Y=0.58 $X2=0 $Y2=0
cc_669 N_X_c_950_n N_VGND_c_1221_n 0.0126571f $X=7.03 $Y=0.58 $X2=0 $Y2=0
cc_670 N_X_c_950_n N_VGND_c_1222_n 0.0125556f $X=7.03 $Y=0.58 $X2=0 $Y2=0
cc_671 N_X_c_951_n N_VGND_c_1222_n 0.0126571f $X=7.96 $Y=0.58 $X2=0 $Y2=0
cc_672 N_X_c_951_n N_VGND_c_1223_n 0.0125556f $X=7.96 $Y=0.58 $X2=0 $Y2=0
cc_673 N_X_c_952_n N_VGND_c_1223_n 0.0126571f $X=8.89 $Y=0.58 $X2=0 $Y2=0
cc_674 N_X_c_952_n N_VGND_c_1225_n 0.0148853f $X=8.89 $Y=0.58 $X2=0 $Y2=0
cc_675 N_X_c_946_n N_VGND_c_1230_n 0.0119584f $X=2.52 $Y=0.58 $X2=0 $Y2=0
cc_676 N_X_c_947_n N_VGND_c_1232_n 0.00995046f $X=3.38 $Y=0.58 $X2=0 $Y2=0
cc_677 N_X_c_948_n N_VGND_c_1234_n 0.0101616f $X=5.17 $Y=0.58 $X2=0 $Y2=0
cc_678 N_X_c_949_n N_VGND_c_1235_n 0.0109942f $X=6.1 $Y=0.58 $X2=0 $Y2=0
cc_679 N_X_c_950_n N_VGND_c_1236_n 0.0109942f $X=7.03 $Y=0.58 $X2=0 $Y2=0
cc_680 N_X_c_951_n N_VGND_c_1237_n 0.0109942f $X=7.96 $Y=0.58 $X2=0 $Y2=0
cc_681 N_X_c_952_n N_VGND_c_1238_n 0.0109942f $X=8.89 $Y=0.58 $X2=0 $Y2=0
cc_682 N_X_c_946_n N_VGND_c_1244_n 0.00989813f $X=2.52 $Y=0.58 $X2=0 $Y2=0
cc_683 N_X_c_947_n N_VGND_c_1244_n 0.00823613f $X=3.38 $Y=0.58 $X2=0 $Y2=0
cc_684 N_X_c_948_n N_VGND_c_1244_n 0.00840151f $X=5.17 $Y=0.58 $X2=0 $Y2=0
cc_685 N_X_c_949_n N_VGND_c_1244_n 0.00904371f $X=6.1 $Y=0.58 $X2=0 $Y2=0
cc_686 N_X_c_950_n N_VGND_c_1244_n 0.00904371f $X=7.03 $Y=0.58 $X2=0 $Y2=0
cc_687 N_X_c_951_n N_VGND_c_1244_n 0.00904371f $X=7.96 $Y=0.58 $X2=0 $Y2=0
cc_688 N_X_c_952_n N_VGND_c_1244_n 0.00904371f $X=8.89 $Y=0.58 $X2=0 $Y2=0
cc_689 N_X_c_953_n N_VGND_c_1244_n 0.00953689f $X=4.24 $Y=0.58 $X2=0 $Y2=0
