* NGSPICE file created from sky130_fd_sc_ls__o21ba_2.ext - technology: sky130A

.subckt sky130_fd_sc_ls__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
M1000 VGND a_177_48# X VNB nshort w=740000u l=150000u
+  ad=7.8915e+11p pd=6.84e+06u as=2.072e+11p ps=2.04e+06u
M1001 VGND A2 a_487_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=4.07e+11p ps=4.06e+06u
M1002 VGND B1_N a_27_74# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=1.5125e+11p ps=1.65e+06u
M1003 VPWR B1_N a_27_74# VPB phighvt w=840000u l=150000u
+  ad=1.511e+12p pd=9.31e+06u as=2.478e+11p ps=2.27e+06u
M1004 a_177_48# a_27_74# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=3e+11p pd=2.6e+06u as=0p ps=0u
M1005 X a_177_48# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=0p ps=0u
M1006 X a_177_48# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_487_74# A1 VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_582_368# A2 a_177_48# VPB phighvt w=1e+06u l=150000u
+  ad=3.6e+11p pd=2.72e+06u as=0p ps=0u
M1009 VPWR A1 a_582_368# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR a_177_48# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_487_74# a_27_74# a_177_48# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.035e+11p ps=2.03e+06u
.ends

