* File: sky130_fd_sc_ls__a2bb2o_1.spice
* Created: Fri Aug 28 12:56:10 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__a2bb2o_1.pex.spice"
.subckt sky130_fd_sc_ls__a2bb2o_1  VNB VPB A1_N A2_N B2 B1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* B1	B1
* B2	B2
* A2_N	A2_N
* A1_N	A1_N
* VPB	VPB
* VNB	VNB
MM1007 N_VGND_M1007_d N_A_93_264#_M1007_g N_X_M1007_s VNB NSHORT L=0.15 W=0.74
+ AD=0.136154 AS=0.1961 PD=1.23907 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75002.2 A=0.111 P=1.78 MULT=1
MM1003 N_A_257_126#_M1003_d N_A1_N_M1003_g N_VGND_M1007_d VNB NSHORT L=0.15
+ W=0.55 AD=0.077 AS=0.101196 PD=0.83 PS=0.92093 NRD=0 NRS=13.632 M=1 R=3.66667
+ SA=75000.7 SB=75002.5 A=0.0825 P=1.4 MULT=1
MM1005 N_VGND_M1005_d N_A2_N_M1005_g N_A_257_126#_M1003_d VNB NSHORT L=0.15
+ W=0.55 AD=0.195966 AS=0.077 PD=1.26639 PS=0.83 NRD=15.264 NRS=0 M=1 R=3.66667
+ SA=75001.1 SB=75002 A=0.0825 P=1.4 MULT=1
MM1001 N_A_93_264#_M1001_d N_A_257_126#_M1001_g N_VGND_M1005_d VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.228034 PD=0.92 PS=1.47361 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.7 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1002 A_605_126# N_B2_M1002_g N_A_93_264#_M1001_d VNB NSHORT L=0.15 W=0.64
+ AD=0.1248 AS=0.0896 PD=1.03 PS=0.92 NRD=26.244 NRS=0 M=1 R=4.26667 SA=75002.2
+ SB=75000.7 A=0.096 P=1.58 MULT=1
MM1008 N_VGND_M1008_d N_B1_M1008_g A_605_126# VNB NSHORT L=0.15 W=0.64 AD=0.1696
+ AS=0.1248 PD=1.81 PS=1.03 NRD=0 NRS=26.244 M=1 R=4.26667 SA=75002.7 SB=75000.2
+ A=0.096 P=1.58 MULT=1
MM1010 N_VPWR_M1010_d N_A_93_264#_M1010_g N_X_M1010_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.210264 AS=0.308 PD=1.56906 PS=2.79 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75001 A=0.168 P=2.54 MULT=1
MM1011 A_258_392# N_A1_N_M1011_g N_VPWR_M1010_d VPB PHIGHVT L=0.15 W=1 AD=0.12
+ AS=0.187736 PD=1.24 PS=1.40094 NRD=12.7853 NRS=14.7553 M=1 R=6.66667
+ SA=75000.7 SB=75000.6 A=0.15 P=2.3 MULT=1
MM1006 N_A_257_126#_M1006_d N_A2_N_M1006_g A_258_392# VPB PHIGHVT L=0.15 W=1
+ AD=0.275 AS=0.12 PD=2.55 PS=1.24 NRD=1.9503 NRS=12.7853 M=1 R=6.66667
+ SA=75001.1 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1004 N_A_530_392#_M1004_d N_A_257_126#_M1004_g N_A_93_264#_M1004_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.15 AS=0.275 PD=1.3 PS=2.55 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75001.1 A=0.15 P=2.3 MULT=1
MM1000 N_VPWR_M1000_d N_B2_M1000_g N_A_530_392#_M1004_d VPB PHIGHVT L=0.15 W=1
+ AD=0.165 AS=0.15 PD=1.33 PS=1.3 NRD=4.9053 NRS=1.9503 M=1 R=6.66667 SA=75000.6
+ SB=75000.7 A=0.15 P=2.3 MULT=1
MM1009 N_A_530_392#_M1009_d N_B1_M1009_g N_VPWR_M1000_d VPB PHIGHVT L=0.15 W=1
+ AD=0.275 AS=0.165 PD=2.55 PS=1.33 NRD=1.9503 NRS=4.9053 M=1 R=6.66667
+ SA=75001.1 SB=75000.2 A=0.15 P=2.3 MULT=1
DX12_noxref VNB VPB NWDIODE A=8.742 P=13.12
*
.include "sky130_fd_sc_ls__a2bb2o_1.pxi.spice"
*
.ends
*
*
