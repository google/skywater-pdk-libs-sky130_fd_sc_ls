* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
M1000 VPWR B1 a_820_392# VPB phighvt w=1e+06u l=150000u
+  ad=1.6808e+12p pd=1.385e+07u as=1.15e+12p ps=1.03e+07u
M1001 VGND a_162_48# X VNB nshort w=740000u l=150000u
+  ad=1.6403e+12p pd=1.199e+07u as=4.144e+11p ps=4.08e+06u
M1002 a_1009_74# B2 a_162_48# VNB nshort w=640000u l=150000u
+  ad=5.184e+11p pd=5.46e+06u as=3.753e+11p ps=3.85e+06u
M1003 X a_162_48# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=6.72e+11p pd=5.68e+06u as=0p ps=0u
M1004 a_586_94# A2_N a_583_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=3.08e+11p pd=2.79e+06u as=2.688e+11p ps=2.72e+06u
M1005 a_820_392# B1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_162_48# a_586_94# a_820_392# VPB phighvt w=1e+06u l=150000u
+  ad=3e+11p pd=2.6e+06u as=0p ps=0u
M1007 a_1009_74# B1 VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR a_162_48# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND B1 a_1009_74# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 X a_162_48# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 X a_162_48# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_162_48# B2 a_1009_74# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_586_94# A1_N VGND VNB nshort w=640000u l=150000u
+  ad=1.792e+11p pd=1.84e+06u as=0p ps=0u
M1014 a_820_392# a_586_94# a_162_48# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_162_48# a_586_94# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR B2 a_820_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 X a_162_48# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_583_368# A1_N VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND a_162_48# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_820_392# B2 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND A2_N a_586_94# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPWR a_162_48# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
