* File: sky130_fd_sc_ls__sdfsbp_2.pxi.spice
* Created: Wed Sep  2 11:27:45 2020
* 
x_PM_SKY130_FD_SC_LS__SDFSBP_2%A_27_74# N_A_27_74#_M1044_s N_A_27_74#_M1008_s
+ N_A_27_74#_M1035_g N_A_27_74#_c_379_n N_A_27_74#_M1042_g N_A_27_74#_c_373_n
+ N_A_27_74#_c_374_n N_A_27_74#_c_381_n N_A_27_74#_c_375_n N_A_27_74#_c_376_n
+ N_A_27_74#_c_382_n N_A_27_74#_c_377_n N_A_27_74#_c_383_n N_A_27_74#_c_384_n
+ N_A_27_74#_c_378_n PM_SKY130_FD_SC_LS__SDFSBP_2%A_27_74#
x_PM_SKY130_FD_SC_LS__SDFSBP_2%SCE N_SCE_M1044_g N_SCE_c_458_n N_SCE_c_459_n
+ N_SCE_M1008_g N_SCE_c_460_n N_SCE_c_461_n N_SCE_M1006_g N_SCE_M1017_g
+ N_SCE_c_451_n N_SCE_c_452_n N_SCE_c_453_n N_SCE_c_454_n SCE N_SCE_c_455_n
+ N_SCE_c_456_n N_SCE_c_457_n PM_SKY130_FD_SC_LS__SDFSBP_2%SCE
x_PM_SKY130_FD_SC_LS__SDFSBP_2%D N_D_c_534_n N_D_c_535_n N_D_c_541_n N_D_M1048_g
+ N_D_M1036_g N_D_c_536_n D D N_D_c_538_n N_D_c_539_n
+ PM_SKY130_FD_SC_LS__SDFSBP_2%D
x_PM_SKY130_FD_SC_LS__SDFSBP_2%SCD N_SCD_c_589_n N_SCD_c_590_n N_SCD_M1030_g
+ N_SCD_c_591_n N_SCD_c_592_n N_SCD_M1018_g N_SCD_c_584_n N_SCD_c_585_n
+ N_SCD_c_586_n SCD N_SCD_c_588_n PM_SKY130_FD_SC_LS__SDFSBP_2%SCD
x_PM_SKY130_FD_SC_LS__SDFSBP_2%CLK N_CLK_c_635_n N_CLK_M1026_g N_CLK_c_636_n
+ N_CLK_M1039_g CLK PM_SKY130_FD_SC_LS__SDFSBP_2%CLK
x_PM_SKY130_FD_SC_LS__SDFSBP_2%A_871_74# N_A_871_74#_M1033_d N_A_871_74#_M1015_d
+ N_A_871_74#_c_692_n N_A_871_74#_c_693_n N_A_871_74#_M1031_g
+ N_A_871_74#_c_669_n N_A_871_74#_c_670_n N_A_871_74#_M1027_g
+ N_A_871_74#_M1032_g N_A_871_74#_M1037_g N_A_871_74#_c_674_n
+ N_A_871_74#_c_675_n N_A_871_74#_c_676_n N_A_871_74#_c_677_n
+ N_A_871_74#_c_695_n N_A_871_74#_M1047_g N_A_871_74#_c_696_n
+ N_A_871_74#_c_678_n N_A_871_74#_c_697_n N_A_871_74#_c_679_n
+ N_A_871_74#_c_680_n N_A_871_74#_c_698_n N_A_871_74#_c_699_n
+ N_A_871_74#_c_681_n N_A_871_74#_c_682_n N_A_871_74#_c_683_n
+ N_A_871_74#_c_684_n N_A_871_74#_c_703_n N_A_871_74#_c_704_n
+ N_A_871_74#_c_705_n N_A_871_74#_c_706_n N_A_871_74#_c_707_n
+ N_A_871_74#_c_708_n N_A_871_74#_c_709_n N_A_871_74#_c_710_n
+ N_A_871_74#_c_685_n N_A_871_74#_c_686_n N_A_871_74#_c_687_n
+ N_A_871_74#_c_688_n N_A_871_74#_c_689_n N_A_871_74#_c_712_n
+ N_A_871_74#_c_690_n N_A_871_74#_c_691_n PM_SKY130_FD_SC_LS__SDFSBP_2%A_871_74#
x_PM_SKY130_FD_SC_LS__SDFSBP_2%A_1252_376# N_A_1252_376#_M1012_s
+ N_A_1252_376#_M1016_d N_A_1252_376#_c_947_n N_A_1252_376#_M1034_g
+ N_A_1252_376#_c_948_n N_A_1252_376#_c_941_n N_A_1252_376#_M1024_g
+ N_A_1252_376#_c_949_n N_A_1252_376#_c_950_n N_A_1252_376#_c_951_n
+ N_A_1252_376#_c_942_n N_A_1252_376#_c_943_n N_A_1252_376#_c_944_n
+ N_A_1252_376#_c_952_n N_A_1252_376#_c_953_n N_A_1252_376#_c_945_n
+ N_A_1252_376#_c_946_n PM_SKY130_FD_SC_LS__SDFSBP_2%A_1252_376#
x_PM_SKY130_FD_SC_LS__SDFSBP_2%A_1069_81# N_A_1069_81#_M1019_d
+ N_A_1069_81#_M1031_d N_A_1069_81#_c_1032_n N_A_1069_81#_c_1053_n
+ N_A_1069_81#_M1016_g N_A_1069_81#_M1012_g N_A_1069_81#_c_1034_n
+ N_A_1069_81#_c_1035_n N_A_1069_81#_c_1055_n N_A_1069_81#_M1002_g
+ N_A_1069_81#_M1001_g N_A_1069_81#_c_1036_n N_A_1069_81#_c_1037_n
+ N_A_1069_81#_c_1057_n N_A_1069_81#_M1043_g N_A_1069_81#_M1009_g
+ N_A_1069_81#_c_1039_n N_A_1069_81#_c_1040_n N_A_1069_81#_c_1041_n
+ N_A_1069_81#_c_1074_n N_A_1069_81#_c_1078_n N_A_1069_81#_c_1042_n
+ N_A_1069_81#_c_1043_n N_A_1069_81#_c_1044_n N_A_1069_81#_c_1045_n
+ N_A_1069_81#_c_1046_n N_A_1069_81#_c_1047_n N_A_1069_81#_c_1048_n
+ N_A_1069_81#_c_1058_n N_A_1069_81#_c_1049_n N_A_1069_81#_c_1050_n
+ N_A_1069_81#_c_1051_n PM_SKY130_FD_SC_LS__SDFSBP_2%A_1069_81#
x_PM_SKY130_FD_SC_LS__SDFSBP_2%SET_B N_SET_B_c_1229_n N_SET_B_c_1230_n
+ N_SET_B_M1029_g N_SET_B_M1013_g N_SET_B_M1021_g N_SET_B_c_1231_n
+ N_SET_B_c_1232_n N_SET_B_M1014_g N_SET_B_c_1221_n N_SET_B_c_1234_n
+ N_SET_B_c_1222_n N_SET_B_c_1223_n N_SET_B_c_1224_n SET_B N_SET_B_c_1226_n
+ N_SET_B_c_1227_n N_SET_B_c_1228_n PM_SKY130_FD_SC_LS__SDFSBP_2%SET_B
x_PM_SKY130_FD_SC_LS__SDFSBP_2%A_619_368# N_A_619_368#_M1039_s
+ N_A_619_368#_M1026_s N_A_619_368#_M1033_g N_A_619_368#_c_1387_n
+ N_A_619_368#_M1015_g N_A_619_368#_c_1370_n N_A_619_368#_c_1388_n
+ N_A_619_368#_c_1371_n N_A_619_368#_c_1372_n N_A_619_368#_c_1389_n
+ N_A_619_368#_c_1390_n N_A_619_368#_c_1373_n N_A_619_368#_M1019_g
+ N_A_619_368#_c_1391_n N_A_619_368#_c_1392_n N_A_619_368#_c_1393_n
+ N_A_619_368#_M1040_g N_A_619_368#_c_1394_n N_A_619_368#_c_1395_n
+ N_A_619_368#_c_1396_n N_A_619_368#_M1005_g N_A_619_368#_c_1397_n
+ N_A_619_368#_c_1398_n N_A_619_368#_c_1399_n N_A_619_368#_M1046_g
+ N_A_619_368#_c_1400_n N_A_619_368#_c_1401_n N_A_619_368#_c_1402_n
+ N_A_619_368#_c_1403_n N_A_619_368#_c_1374_n N_A_619_368#_c_1375_n
+ N_A_619_368#_c_1376_n N_A_619_368#_M1007_g N_A_619_368#_c_1377_n
+ N_A_619_368#_c_1378_n N_A_619_368#_c_1379_n N_A_619_368#_c_1408_n
+ N_A_619_368#_c_1409_n N_A_619_368#_c_1380_n N_A_619_368#_c_1381_n
+ N_A_619_368#_c_1382_n N_A_619_368#_c_1411_n N_A_619_368#_c_1383_n
+ N_A_619_368#_c_1413_n N_A_619_368#_c_1384_n N_A_619_368#_c_1414_n
+ N_A_619_368#_c_1385_n N_A_619_368#_c_1386_n N_A_619_368#_c_1416_n
+ PM_SKY130_FD_SC_LS__SDFSBP_2%A_619_368#
x_PM_SKY130_FD_SC_LS__SDFSBP_2%A_2513_258# N_A_2513_258#_M1038_d
+ N_A_2513_258#_M1041_s N_A_2513_258#_c_1654_n N_A_2513_258#_c_1655_n
+ N_A_2513_258#_M1003_g N_A_2513_258#_M1020_g N_A_2513_258#_c_1646_n
+ N_A_2513_258#_c_1657_n N_A_2513_258#_c_1647_n N_A_2513_258#_c_1648_n
+ N_A_2513_258#_c_1649_n N_A_2513_258#_c_1650_n N_A_2513_258#_c_1651_n
+ N_A_2513_258#_c_1652_n N_A_2513_258#_c_1653_n N_A_2513_258#_c_1660_n
+ PM_SKY130_FD_SC_LS__SDFSBP_2%A_2513_258#
x_PM_SKY130_FD_SC_LS__SDFSBP_2%A_2067_74# N_A_2067_74#_M1032_s
+ N_A_2067_74#_M1007_s N_A_2067_74#_M1005_s N_A_2067_74#_M1047_d
+ N_A_2067_74#_M1014_d N_A_2067_74#_M1038_g N_A_2067_74#_c_1749_n
+ N_A_2067_74#_c_1768_n N_A_2067_74#_c_1769_n N_A_2067_74#_c_1770_n
+ N_A_2067_74#_M1041_g N_A_2067_74#_M1022_g N_A_2067_74#_c_1751_n
+ N_A_2067_74#_c_1772_n N_A_2067_74#_M1000_g N_A_2067_74#_c_1752_n
+ N_A_2067_74#_M1025_g N_A_2067_74#_c_1754_n N_A_2067_74#_c_1774_n
+ N_A_2067_74#_M1045_g N_A_2067_74#_c_1755_n N_A_2067_74#_c_1756_n
+ N_A_2067_74#_c_1776_n N_A_2067_74#_M1004_g N_A_2067_74#_M1010_g
+ N_A_2067_74#_c_1758_n N_A_2067_74#_c_1777_n N_A_2067_74#_c_1759_n
+ N_A_2067_74#_c_1760_n N_A_2067_74#_c_1761_n N_A_2067_74#_c_1804_n
+ N_A_2067_74#_c_1778_n N_A_2067_74#_c_1805_n N_A_2067_74#_c_1762_n
+ N_A_2067_74#_c_1841_n N_A_2067_74#_c_1763_n N_A_2067_74#_c_1779_n
+ N_A_2067_74#_c_1780_n N_A_2067_74#_c_1781_n N_A_2067_74#_c_1782_n
+ N_A_2067_74#_c_1764_n N_A_2067_74#_c_1765_n N_A_2067_74#_c_1766_n
+ N_A_2067_74#_c_1784_n N_A_2067_74#_c_1767_n
+ PM_SKY130_FD_SC_LS__SDFSBP_2%A_2067_74#
x_PM_SKY130_FD_SC_LS__SDFSBP_2%A_3177_368# N_A_3177_368#_M1010_s
+ N_A_3177_368#_M1004_s N_A_3177_368#_c_1995_n N_A_3177_368#_M1011_g
+ N_A_3177_368#_M1023_g N_A_3177_368#_c_1996_n N_A_3177_368#_M1028_g
+ N_A_3177_368#_M1049_g N_A_3177_368#_c_1990_n N_A_3177_368#_c_1991_n
+ N_A_3177_368#_c_1992_n N_A_3177_368#_c_1993_n N_A_3177_368#_c_1994_n
+ PM_SKY130_FD_SC_LS__SDFSBP_2%A_3177_368#
x_PM_SKY130_FD_SC_LS__SDFSBP_2%VPWR N_VPWR_M1008_d N_VPWR_M1030_d N_VPWR_M1026_d
+ N_VPWR_M1034_d N_VPWR_M1029_d N_VPWR_M1002_s N_VPWR_M1003_d N_VPWR_M1041_d
+ N_VPWR_M1045_s N_VPWR_M1004_d N_VPWR_M1028_s N_VPWR_c_2058_n N_VPWR_c_2059_n
+ N_VPWR_c_2060_n N_VPWR_c_2061_n N_VPWR_c_2062_n N_VPWR_c_2063_n
+ N_VPWR_c_2064_n N_VPWR_c_2065_n N_VPWR_c_2066_n N_VPWR_c_2067_n
+ N_VPWR_c_2068_n N_VPWR_c_2069_n N_VPWR_c_2070_n N_VPWR_c_2071_n
+ N_VPWR_c_2072_n N_VPWR_c_2073_n N_VPWR_c_2074_n N_VPWR_c_2075_n
+ N_VPWR_c_2076_n N_VPWR_c_2077_n VPWR N_VPWR_c_2078_n N_VPWR_c_2079_n
+ N_VPWR_c_2080_n N_VPWR_c_2081_n N_VPWR_c_2082_n N_VPWR_c_2083_n
+ N_VPWR_c_2084_n N_VPWR_c_2085_n N_VPWR_c_2086_n N_VPWR_c_2087_n
+ N_VPWR_c_2088_n N_VPWR_c_2089_n N_VPWR_c_2057_n
+ PM_SKY130_FD_SC_LS__SDFSBP_2%VPWR
x_PM_SKY130_FD_SC_LS__SDFSBP_2%A_304_464# N_A_304_464#_M1036_d
+ N_A_304_464#_M1019_s N_A_304_464#_M1048_d N_A_304_464#_M1031_s
+ N_A_304_464#_c_2260_n N_A_304_464#_c_2257_n N_A_304_464#_c_2262_n
+ N_A_304_464#_c_2263_n N_A_304_464#_c_2264_n N_A_304_464#_c_2279_n
+ N_A_304_464#_c_2298_n N_A_304_464#_c_2300_n N_A_304_464#_c_2258_n
+ N_A_304_464#_c_2265_n N_A_304_464#_c_2259_n
+ PM_SKY130_FD_SC_LS__SDFSBP_2%A_304_464#
x_PM_SKY130_FD_SC_LS__SDFSBP_2%A_1789_424# N_A_1789_424#_M1002_d
+ N_A_1789_424#_M1043_d N_A_1789_424#_M1046_d N_A_1789_424#_c_2379_n
+ N_A_1789_424#_c_2373_n N_A_1789_424#_c_2382_n N_A_1789_424#_c_2374_n
+ N_A_1789_424#_c_2375_n N_A_1789_424#_c_2376_n N_A_1789_424#_c_2377_n
+ PM_SKY130_FD_SC_LS__SDFSBP_2%A_1789_424#
x_PM_SKY130_FD_SC_LS__SDFSBP_2%A_2277_455# N_A_2277_455#_M1047_s
+ N_A_2277_455#_M1003_s N_A_2277_455#_c_2427_n N_A_2277_455#_c_2428_n
+ N_A_2277_455#_c_2429_n N_A_2277_455#_c_2430_n
+ PM_SKY130_FD_SC_LS__SDFSBP_2%A_2277_455#
x_PM_SKY130_FD_SC_LS__SDFSBP_2%Q_N N_Q_N_M1022_d N_Q_N_M1000_d N_Q_N_c_2459_n
+ Q_N Q_N Q_N N_Q_N_c_2460_n Q_N PM_SKY130_FD_SC_LS__SDFSBP_2%Q_N
x_PM_SKY130_FD_SC_LS__SDFSBP_2%Q N_Q_M1023_d N_Q_M1011_d N_Q_c_2490_n
+ N_Q_c_2491_n N_Q_c_2487_n Q Q Q PM_SKY130_FD_SC_LS__SDFSBP_2%Q
x_PM_SKY130_FD_SC_LS__SDFSBP_2%VGND N_VGND_M1044_d N_VGND_M1018_d N_VGND_M1039_d
+ N_VGND_M1024_d N_VGND_M1013_d N_VGND_M1001_d N_VGND_M1021_d N_VGND_M1022_s
+ N_VGND_M1025_s N_VGND_M1010_d N_VGND_M1049_s N_VGND_c_2517_n N_VGND_c_2518_n
+ N_VGND_c_2519_n N_VGND_c_2520_n N_VGND_c_2521_n N_VGND_c_2522_n
+ N_VGND_c_2523_n N_VGND_c_2524_n N_VGND_c_2525_n N_VGND_c_2526_n
+ N_VGND_c_2527_n N_VGND_c_2528_n N_VGND_c_2529_n N_VGND_c_2530_n
+ N_VGND_c_2531_n N_VGND_c_2532_n N_VGND_c_2533_n N_VGND_c_2534_n
+ N_VGND_c_2535_n N_VGND_c_2536_n N_VGND_c_2537_n N_VGND_c_2538_n VGND
+ N_VGND_c_2539_n N_VGND_c_2540_n N_VGND_c_2541_n N_VGND_c_2542_n
+ N_VGND_c_2543_n N_VGND_c_2544_n N_VGND_c_2545_n N_VGND_c_2546_n
+ N_VGND_c_2547_n N_VGND_c_2548_n N_VGND_c_2549_n N_VGND_c_2550_n
+ PM_SKY130_FD_SC_LS__SDFSBP_2%VGND
x_PM_SKY130_FD_SC_LS__SDFSBP_2%A_1794_74# N_A_1794_74#_M1001_s
+ N_A_1794_74#_M1009_s N_A_1794_74#_M1037_d N_A_1794_74#_c_2704_n
+ N_A_1794_74#_c_2705_n N_A_1794_74#_c_2706_n N_A_1794_74#_c_2714_n
+ N_A_1794_74#_c_2707_n N_A_1794_74#_c_2708_n N_A_1794_74#_c_2709_n
+ PM_SKY130_FD_SC_LS__SDFSBP_2%A_1794_74#
cc_1 VNB N_A_27_74#_c_373_n 0.0250407f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=0.58
cc_2 VNB N_A_27_74#_c_374_n 0.0202447f $X=-0.19 $Y=-0.245 $X2=0.17 $Y2=1.97
cc_3 VNB N_A_27_74#_c_375_n 0.00761332f $X=-0.19 $Y=-0.245 $X2=0.98 $Y2=1.065
cc_4 VNB N_A_27_74#_c_376_n 0.0300878f $X=-0.19 $Y=-0.245 $X2=0.98 $Y2=1.065
cc_5 VNB N_A_27_74#_c_377_n 0.0219083f $X=-0.19 $Y=-0.245 $X2=0.265 $Y2=1.065
cc_6 VNB N_A_27_74#_c_378_n 0.0178945f $X=-0.19 $Y=-0.245 $X2=0.98 $Y2=0.9
cc_7 VNB N_SCE_M1044_g 0.0623069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_SCE_c_451_n 0.0331355f $X=-0.19 $Y=-0.245 $X2=0.275 $Y2=2.465
cc_9 VNB N_SCE_c_452_n 0.00270489f $X=-0.19 $Y=-0.245 $X2=0.445 $Y2=1.065
cc_10 VNB N_SCE_c_453_n 0.0319242f $X=-0.19 $Y=-0.245 $X2=0.98 $Y2=1.065
cc_11 VNB N_SCE_c_454_n 0.00219979f $X=-0.19 $Y=-0.245 $X2=0.98 $Y2=1.065
cc_12 VNB N_SCE_c_455_n 0.0798121f $X=-0.19 $Y=-0.245 $X2=1.94 $Y2=1.975
cc_13 VNB N_SCE_c_456_n 0.00307321f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_SCE_c_457_n 0.0216104f $X=-0.19 $Y=-0.245 $X2=1.94 $Y2=2.055
cc_15 VNB N_D_c_534_n 0.00539996f $X=-0.19 $Y=-0.245 $X2=0.135 $Y2=0.37
cc_16 VNB N_D_c_535_n 0.00813295f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=2.32
cc_17 VNB N_D_c_536_n 0.0190815f $X=-0.19 $Y=-0.245 $X2=2.015 $Y2=2.64
cc_18 VNB D 0.00579289f $X=-0.19 $Y=-0.245 $X2=2.015 $Y2=2.64
cc_19 VNB N_D_c_538_n 0.0316793f $X=-0.19 $Y=-0.245 $X2=0.17 $Y2=1.23
cc_20 VNB N_D_c_539_n 0.0221915f $X=-0.19 $Y=-0.245 $X2=0.275 $Y2=2.14
cc_21 VNB N_SCD_M1018_g 0.0227695f $X=-0.19 $Y=-0.245 $X2=2.015 $Y2=2.245
cc_22 VNB N_SCD_c_584_n 0.0189523f $X=-0.19 $Y=-0.245 $X2=0.265 $Y2=0.9
cc_23 VNB N_SCD_c_585_n 0.00249185f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=0.58
cc_24 VNB N_SCD_c_586_n 0.0251837f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB SCD 0.00682024f $X=-0.19 $Y=-0.245 $X2=0.17 $Y2=1.23
cc_26 VNB N_SCD_c_588_n 0.0246471f $X=-0.19 $Y=-0.245 $X2=0.275 $Y2=2.465
cc_27 VNB N_CLK_c_635_n 0.0643171f $X=-0.19 $Y=-0.245 $X2=0.135 $Y2=0.37
cc_28 VNB N_CLK_c_636_n 0.0194708f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB CLK 0.00951065f $X=-0.19 $Y=-0.245 $X2=1.07 $Y2=0.9
cc_30 VNB N_A_871_74#_c_669_n 0.0346908f $X=-0.19 $Y=-0.245 $X2=2.015 $Y2=2.64
cc_31 VNB N_A_871_74#_c_670_n 0.0157874f $X=-0.19 $Y=-0.245 $X2=0.265 $Y2=0.9
cc_32 VNB N_A_871_74#_M1027_g 0.0207425f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_871_74#_M1032_g 0.0204977f $X=-0.19 $Y=-0.245 $X2=0.275 $Y2=2.465
cc_34 VNB N_A_871_74#_M1037_g 0.0284098f $X=-0.19 $Y=-0.245 $X2=0.98 $Y2=1.065
cc_35 VNB N_A_871_74#_c_674_n 0.028453f $X=-0.19 $Y=-0.245 $X2=0.98 $Y2=1.065
cc_36 VNB N_A_871_74#_c_675_n 0.0466008f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_871_74#_c_676_n 0.0332744f $X=-0.19 $Y=-0.245 $X2=1.775 $Y2=2.055
cc_38 VNB N_A_871_74#_c_677_n 0.00269371f $X=-0.19 $Y=-0.245 $X2=0.275 $Y2=2.055
cc_39 VNB N_A_871_74#_c_678_n 0.00620399f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_871_74#_c_679_n 0.0173245f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_871_74#_c_680_n 0.00279267f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_871_74#_c_681_n 0.00319375f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_871_74#_c_682_n 0.0172406f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_871_74#_c_683_n 0.00181342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_871_74#_c_684_n 0.0689707f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_871_74#_c_685_n 0.00513279f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_871_74#_c_686_n 0.00422606f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_871_74#_c_687_n 2.07961e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_871_74#_c_688_n 0.00317624f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_871_74#_c_689_n 0.00914437f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_871_74#_c_690_n 0.0200525f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_871_74#_c_691_n 0.0263125f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_1252_376#_c_941_n 0.0167981f $X=-0.19 $Y=-0.245 $X2=2.015 $Y2=2.64
cc_54 VNB N_A_1252_376#_c_942_n 0.0137517f $X=-0.19 $Y=-0.245 $X2=0.98 $Y2=1.065
cc_55 VNB N_A_1252_376#_c_943_n 0.00892759f $X=-0.19 $Y=-0.245 $X2=1.775
+ $Y2=2.055
cc_56 VNB N_A_1252_376#_c_944_n 0.00356983f $X=-0.19 $Y=-0.245 $X2=1.94
+ $Y2=1.975
cc_57 VNB N_A_1252_376#_c_945_n 0.0230627f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_1252_376#_c_946_n 0.0502327f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_1069_81#_c_1032_n 0.00122075f $X=-0.19 $Y=-0.245 $X2=1.07 $Y2=0.58
cc_60 VNB N_A_1069_81#_M1012_g 0.034972f $X=-0.19 $Y=-0.245 $X2=0.265 $Y2=0.58
cc_61 VNB N_A_1069_81#_c_1034_n 0.0250974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_1069_81#_c_1035_n 0.0181656f $X=-0.19 $Y=-0.245 $X2=0.275 $Y2=2.14
cc_63 VNB N_A_1069_81#_c_1036_n 0.00951082f $X=-0.19 $Y=-0.245 $X2=0.98
+ $Y2=1.065
cc_64 VNB N_A_1069_81#_c_1037_n 0.0155475f $X=-0.19 $Y=-0.245 $X2=0.465
+ $Y2=2.055
cc_65 VNB N_A_1069_81#_M1009_g 0.0215209f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_1069_81#_c_1039_n 0.015267f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_1069_81#_c_1040_n 0.0179261f $X=-0.19 $Y=-0.245 $X2=0.98 $Y2=1.065
cc_68 VNB N_A_1069_81#_c_1041_n 0.00574168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_1069_81#_c_1042_n 0.00683698f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_1069_81#_c_1043_n 0.0100682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_1069_81#_c_1044_n 0.00368108f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_1069_81#_c_1045_n 0.00596292f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_1069_81#_c_1046_n 0.0124499f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_1069_81#_c_1047_n 0.00977247f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_1069_81#_c_1048_n 0.0449671f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_1069_81#_c_1049_n 0.0115114f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_1069_81#_c_1050_n 0.00148462f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_1069_81#_c_1051_n 0.0540624f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_SET_B_M1013_g 0.0580087f $X=-0.19 $Y=-0.245 $X2=1.07 $Y2=0.58
cc_80 VNB N_SET_B_M1021_g 0.0375934f $X=-0.19 $Y=-0.245 $X2=2.015 $Y2=2.64
cc_81 VNB N_SET_B_c_1221_n 0.0107422f $X=-0.19 $Y=-0.245 $X2=0.3 $Y2=2.465
cc_82 VNB N_SET_B_c_1222_n 0.0186488f $X=-0.19 $Y=-0.245 $X2=0.445 $Y2=1.065
cc_83 VNB N_SET_B_c_1223_n 0.00371196f $X=-0.19 $Y=-0.245 $X2=0.98 $Y2=1.065
cc_84 VNB N_SET_B_c_1224_n 0.00210148f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB SET_B 6.21758e-19 $X=-0.19 $Y=-0.245 $X2=0.465 $Y2=2.055
cc_86 VNB N_SET_B_c_1226_n 0.0138031f $X=-0.19 $Y=-0.245 $X2=1.94 $Y2=1.975
cc_87 VNB N_SET_B_c_1227_n 0.00454843f $X=-0.19 $Y=-0.245 $X2=1.94 $Y2=1.975
cc_88 VNB N_SET_B_c_1228_n 0.0145583f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_619_368#_M1033_g 0.0274744f $X=-0.19 $Y=-0.245 $X2=1.07 $Y2=0.58
cc_90 VNB N_A_619_368#_c_1370_n 0.0166547f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=0.58
cc_91 VNB N_A_619_368#_c_1371_n 0.0316114f $X=-0.19 $Y=-0.245 $X2=0.17 $Y2=1.97
cc_92 VNB N_A_619_368#_c_1372_n 0.0104746f $X=-0.19 $Y=-0.245 $X2=0.275 $Y2=2.14
cc_93 VNB N_A_619_368#_c_1373_n 0.0184603f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_619_368#_c_1374_n 0.0235315f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_619_368#_c_1375_n 0.0186956f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_619_368#_c_1376_n 0.0222303f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_619_368#_c_1377_n 0.0127729f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_A_619_368#_c_1378_n 0.0196265f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_A_619_368#_c_1379_n 0.00936606f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_A_619_368#_c_1380_n 0.0563283f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_A_619_368#_c_1381_n 0.00824969f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_A_619_368#_c_1382_n 0.00225483f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_A_619_368#_c_1383_n 0.00368583f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_A_619_368#_c_1384_n 0.00775223f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_A_619_368#_c_1385_n 0.00164982f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_A_619_368#_c_1386_n 0.00823064f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_A_2513_258#_M1020_g 0.0355334f $X=-0.19 $Y=-0.245 $X2=0.265
+ $Y2=0.58
cc_108 VNB N_A_2513_258#_c_1646_n 0.0131618f $X=-0.19 $Y=-0.245 $X2=0.17
+ $Y2=1.97
cc_109 VNB N_A_2513_258#_c_1647_n 9.9353e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_A_2513_258#_c_1648_n 0.0163581f $X=-0.19 $Y=-0.245 $X2=0.445
+ $Y2=1.065
cc_111 VNB N_A_2513_258#_c_1649_n 0.02419f $X=-0.19 $Y=-0.245 $X2=0.98 $Y2=1.065
cc_112 VNB N_A_2513_258#_c_1650_n 0.00837366f $X=-0.19 $Y=-0.245 $X2=0.98
+ $Y2=1.065
cc_113 VNB N_A_2513_258#_c_1651_n 0.0101585f $X=-0.19 $Y=-0.245 $X2=0.465
+ $Y2=2.055
cc_114 VNB N_A_2513_258#_c_1652_n 0.00752831f $X=-0.19 $Y=-0.245 $X2=1.94
+ $Y2=1.975
cc_115 VNB N_A_2513_258#_c_1653_n 0.0155466f $X=-0.19 $Y=-0.245 $X2=1.94
+ $Y2=1.975
cc_116 VNB N_A_2067_74#_M1038_g 0.0460555f $X=-0.19 $Y=-0.245 $X2=0.17 $Y2=1.97
cc_117 VNB N_A_2067_74#_c_1749_n 0.0471136f $X=-0.19 $Y=-0.245 $X2=0.275
+ $Y2=2.465
cc_118 VNB N_A_2067_74#_M1022_g 0.0228116f $X=-0.19 $Y=-0.245 $X2=0.465
+ $Y2=2.055
cc_119 VNB N_A_2067_74#_c_1751_n 0.0122279f $X=-0.19 $Y=-0.245 $X2=1.94
+ $Y2=1.975
cc_120 VNB N_A_2067_74#_c_1752_n 0.0102776f $X=-0.19 $Y=-0.245 $X2=1.94
+ $Y2=2.055
cc_121 VNB N_A_2067_74#_M1025_g 0.0233211f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_A_2067_74#_c_1754_n 0.0136295f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB N_A_2067_74#_c_1755_n 0.058445f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_A_2067_74#_c_1756_n 0.0124376f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_A_2067_74#_M1010_g 0.0258629f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_A_2067_74#_c_1758_n 0.0103217f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_A_2067_74#_c_1759_n 0.00286548f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_A_2067_74#_c_1760_n 0.00286548f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_A_2067_74#_c_1761_n 0.00437802f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_A_2067_74#_c_1762_n 0.00783755f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_A_2067_74#_c_1763_n 0.0118908f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_A_2067_74#_c_1764_n 8.34101e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_A_2067_74#_c_1765_n 0.0137219f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_A_2067_74#_c_1766_n 0.00231564f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_A_2067_74#_c_1767_n 0.00535782f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_A_3177_368#_M1023_g 0.0228691f $X=-0.19 $Y=-0.245 $X2=2.015
+ $Y2=2.64
cc_137 VNB N_A_3177_368#_M1049_g 0.0260188f $X=-0.19 $Y=-0.245 $X2=0.275
+ $Y2=2.14
cc_138 VNB N_A_3177_368#_c_1990_n 0.0120685f $X=-0.19 $Y=-0.245 $X2=0.445
+ $Y2=1.065
cc_139 VNB N_A_3177_368#_c_1991_n 5.42215e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_A_3177_368#_c_1992_n 0.00904052f $X=-0.19 $Y=-0.245 $X2=1.94
+ $Y2=1.975
cc_141 VNB N_A_3177_368#_c_1993_n 0.00280955f $X=-0.19 $Y=-0.245 $X2=1.94
+ $Y2=2.055
cc_142 VNB N_A_3177_368#_c_1994_n 0.0752615f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_143 VNB N_VPWR_c_2057_n 0.740851f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_144 VNB N_A_304_464#_c_2257_n 0.00882071f $X=-0.19 $Y=-0.245 $X2=0.17
+ $Y2=1.97
cc_145 VNB N_A_304_464#_c_2258_n 0.0035679f $X=-0.19 $Y=-0.245 $X2=1.94
+ $Y2=2.055
cc_146 VNB N_A_304_464#_c_2259_n 0.00556247f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_147 VNB N_Q_N_c_2459_n 0.00204548f $X=-0.19 $Y=-0.245 $X2=1.07 $Y2=0.58
cc_148 VNB N_Q_N_c_2460_n 0.00257348f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_149 VNB N_Q_c_2487_n 0.00141953f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=0.58
cc_150 VNB Q 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_151 VNB Q 0.00429087f $X=-0.19 $Y=-0.245 $X2=0.17 $Y2=1.23
cc_152 VNB N_VGND_c_2517_n 0.00723643f $X=-0.19 $Y=-0.245 $X2=1.94 $Y2=2.055
cc_153 VNB N_VGND_c_2518_n 0.00970665f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_154 VNB N_VGND_c_2519_n 0.0054384f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_155 VNB N_VGND_c_2520_n 0.0152393f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_156 VNB N_VGND_c_2521_n 0.00953882f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_157 VNB N_VGND_c_2522_n 0.00396467f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_158 VNB N_VGND_c_2523_n 0.00860026f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_159 VNB N_VGND_c_2524_n 0.0144665f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_160 VNB N_VGND_c_2525_n 0.0217072f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_161 VNB N_VGND_c_2526_n 0.0146831f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_162 VNB N_VGND_c_2527_n 0.010678f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_163 VNB N_VGND_c_2528_n 0.0505285f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_164 VNB N_VGND_c_2529_n 0.0506538f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_165 VNB N_VGND_c_2530_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_166 VNB N_VGND_c_2531_n 0.0271172f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_167 VNB N_VGND_c_2532_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_168 VNB N_VGND_c_2533_n 0.0911645f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_169 VNB N_VGND_c_2534_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_170 VNB N_VGND_c_2535_n 0.0215588f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_171 VNB N_VGND_c_2536_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_172 VNB N_VGND_c_2537_n 0.0199954f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_173 VNB N_VGND_c_2538_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_174 VNB N_VGND_c_2539_n 0.0189171f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_175 VNB N_VGND_c_2540_n 0.018606f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_176 VNB N_VGND_c_2541_n 0.0671019f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_177 VNB N_VGND_c_2542_n 0.0306291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_178 VNB N_VGND_c_2543_n 0.0231281f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_179 VNB N_VGND_c_2544_n 0.0192531f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_180 VNB N_VGND_c_2545_n 0.00760052f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_181 VNB N_VGND_c_2546_n 0.00615422f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_182 VNB N_VGND_c_2547_n 0.00644364f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_183 VNB N_VGND_c_2548_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_184 VNB N_VGND_c_2549_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_185 VNB N_VGND_c_2550_n 0.99539f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_186 VNB N_A_1794_74#_c_2704_n 0.00270668f $X=-0.19 $Y=-0.245 $X2=2.015
+ $Y2=2.64
cc_187 VNB N_A_1794_74#_c_2705_n 0.00449539f $X=-0.19 $Y=-0.245 $X2=0.265
+ $Y2=0.58
cc_188 VNB N_A_1794_74#_c_2706_n 4.59673e-19 $X=-0.19 $Y=-0.245 $X2=0.28
+ $Y2=0.58
cc_189 VNB N_A_1794_74#_c_2707_n 0.00313507f $X=-0.19 $Y=-0.245 $X2=0.275
+ $Y2=2.465
cc_190 VNB N_A_1794_74#_c_2708_n 0.00251555f $X=-0.19 $Y=-0.245 $X2=0.3
+ $Y2=2.465
cc_191 VNB N_A_1794_74#_c_2709_n 0.0118588f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_192 VPB N_A_27_74#_c_379_n 0.0573013f $X=-0.19 $Y=1.66 $X2=2.015 $Y2=2.245
cc_193 VPB N_A_27_74#_c_374_n 0.0147344f $X=-0.19 $Y=1.66 $X2=0.17 $Y2=1.97
cc_194 VPB N_A_27_74#_c_381_n 0.0378239f $X=-0.19 $Y=1.66 $X2=0.3 $Y2=2.465
cc_195 VPB N_A_27_74#_c_382_n 0.0226472f $X=-0.19 $Y=1.66 $X2=1.775 $Y2=2.055
cc_196 VPB N_A_27_74#_c_383_n 0.0146808f $X=-0.19 $Y=1.66 $X2=0.275 $Y2=2.055
cc_197 VPB N_A_27_74#_c_384_n 0.00434281f $X=-0.19 $Y=1.66 $X2=1.94 $Y2=1.975
cc_198 VPB N_SCE_c_458_n 0.0231289f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_199 VPB N_SCE_c_459_n 0.0274034f $X=-0.19 $Y=1.66 $X2=1.07 $Y2=0.9
cc_200 VPB N_SCE_c_460_n 0.0179563f $X=-0.19 $Y=1.66 $X2=2.015 $Y2=2.64
cc_201 VPB N_SCE_c_461_n 0.0217424f $X=-0.19 $Y=1.66 $X2=2.015 $Y2=2.64
cc_202 VPB N_SCE_c_453_n 0.0205042f $X=-0.19 $Y=1.66 $X2=0.98 $Y2=1.065
cc_203 VPB N_D_c_535_n 0.0294353f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=2.32
cc_204 VPB N_D_c_541_n 0.0234165f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_205 VPB N_SCD_c_589_n 0.0125823f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=2.32
cc_206 VPB N_SCD_c_590_n 0.0243896f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_207 VPB N_SCD_c_591_n 0.0258796f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_208 VPB N_SCD_c_592_n 0.00933139f $X=-0.19 $Y=1.66 $X2=1.07 $Y2=0.9
cc_209 VPB N_SCD_c_585_n 0.00949905f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=0.58
cc_210 VPB N_CLK_c_635_n 0.0269913f $X=-0.19 $Y=1.66 $X2=0.135 $Y2=0.37
cc_211 VPB N_A_871_74#_c_692_n 0.012306f $X=-0.19 $Y=1.66 $X2=1.07 $Y2=0.58
cc_212 VPB N_A_871_74#_c_693_n 0.0209205f $X=-0.19 $Y=1.66 $X2=1.07 $Y2=0.58
cc_213 VPB N_A_871_74#_c_677_n 0.0285735f $X=-0.19 $Y=1.66 $X2=0.275 $Y2=2.055
cc_214 VPB N_A_871_74#_c_695_n 0.0199358f $X=-0.19 $Y=1.66 $X2=1.94 $Y2=1.975
cc_215 VPB N_A_871_74#_c_696_n 0.017836f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_216 VPB N_A_871_74#_c_697_n 0.00349515f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_217 VPB N_A_871_74#_c_698_n 0.0218722f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_218 VPB N_A_871_74#_c_699_n 0.00392415f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_219 VPB N_A_871_74#_c_681_n 0.00209765f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_220 VPB N_A_871_74#_c_682_n 0.0105641f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_221 VPB N_A_871_74#_c_683_n 0.00588447f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_222 VPB N_A_871_74#_c_703_n 0.00283177f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_223 VPB N_A_871_74#_c_704_n 0.0116178f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_224 VPB N_A_871_74#_c_705_n 0.00424862f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_225 VPB N_A_871_74#_c_706_n 0.016016f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_226 VPB N_A_871_74#_c_707_n 0.00260538f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_227 VPB N_A_871_74#_c_708_n 0.00310194f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_228 VPB N_A_871_74#_c_709_n 0.0138834f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_229 VPB N_A_871_74#_c_710_n 4.80289e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_230 VPB N_A_871_74#_c_685_n 0.0077675f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_231 VPB N_A_871_74#_c_712_n 9.20603e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_232 VPB N_A_1252_376#_c_947_n 0.0147727f $X=-0.19 $Y=1.66 $X2=1.07 $Y2=0.9
cc_233 VPB N_A_1252_376#_c_948_n 0.012809f $X=-0.19 $Y=1.66 $X2=2.015 $Y2=2.245
cc_234 VPB N_A_1252_376#_c_949_n 0.0308948f $X=-0.19 $Y=1.66 $X2=0.17 $Y2=1.23
cc_235 VPB N_A_1252_376#_c_950_n 0.0122171f $X=-0.19 $Y=1.66 $X2=0.275 $Y2=2.14
cc_236 VPB N_A_1252_376#_c_951_n 0.0357008f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_237 VPB N_A_1252_376#_c_952_n 0.00684637f $X=-0.19 $Y=1.66 $X2=0.98 $Y2=0.9
cc_238 VPB N_A_1252_376#_c_953_n 0.00243757f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_239 VPB N_A_1252_376#_c_945_n 0.00261721f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_240 VPB N_A_1069_81#_c_1032_n 0.0305354f $X=-0.19 $Y=1.66 $X2=1.07 $Y2=0.58
cc_241 VPB N_A_1069_81#_c_1053_n 0.0209064f $X=-0.19 $Y=1.66 $X2=1.07 $Y2=0.58
cc_242 VPB N_A_1069_81#_c_1035_n 0.0132763f $X=-0.19 $Y=1.66 $X2=0.275 $Y2=2.14
cc_243 VPB N_A_1069_81#_c_1055_n 0.022294f $X=-0.19 $Y=1.66 $X2=0.275 $Y2=2.465
cc_244 VPB N_A_1069_81#_c_1037_n 0.0182859f $X=-0.19 $Y=1.66 $X2=0.465 $Y2=2.055
cc_245 VPB N_A_1069_81#_c_1057_n 0.0208593f $X=-0.19 $Y=1.66 $X2=0.265 $Y2=1.065
cc_246 VPB N_A_1069_81#_c_1058_n 0.00846582f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_247 VPB N_A_1069_81#_c_1049_n 0.0108589f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_248 VPB N_SET_B_c_1229_n 0.0183162f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=2.32
cc_249 VPB N_SET_B_c_1230_n 0.0214803f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_250 VPB N_SET_B_c_1231_n 0.0219386f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=0.58
cc_251 VPB N_SET_B_c_1232_n 0.0271398f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_252 VPB N_SET_B_c_1221_n 0.0079736f $X=-0.19 $Y=1.66 $X2=0.3 $Y2=2.465
cc_253 VPB N_SET_B_c_1234_n 0.0130201f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_254 VPB N_SET_B_c_1222_n 0.0112351f $X=-0.19 $Y=1.66 $X2=0.445 $Y2=1.065
cc_255 VPB N_SET_B_c_1223_n 0.0024764f $X=-0.19 $Y=1.66 $X2=0.98 $Y2=1.065
cc_256 VPB N_SET_B_c_1224_n 0.00529978f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_257 VPB SET_B 6.00473e-19 $X=-0.19 $Y=1.66 $X2=0.465 $Y2=2.055
cc_258 VPB N_SET_B_c_1227_n 0.00391415f $X=-0.19 $Y=1.66 $X2=1.94 $Y2=1.975
cc_259 VPB N_SET_B_c_1228_n 0.0196655f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_260 VPB N_A_619_368#_c_1387_n 0.0173954f $X=-0.19 $Y=1.66 $X2=2.015 $Y2=2.64
cc_261 VPB N_A_619_368#_c_1388_n 0.0766195f $X=-0.19 $Y=1.66 $X2=0.17 $Y2=1.23
cc_262 VPB N_A_619_368#_c_1389_n 0.0602166f $X=-0.19 $Y=1.66 $X2=0.275 $Y2=2.465
cc_263 VPB N_A_619_368#_c_1390_n 0.0123948f $X=-0.19 $Y=1.66 $X2=0.3 $Y2=2.465
cc_264 VPB N_A_619_368#_c_1391_n 0.00745764f $X=-0.19 $Y=1.66 $X2=0.98 $Y2=1.065
cc_265 VPB N_A_619_368#_c_1392_n 0.0131636f $X=-0.19 $Y=1.66 $X2=0.98 $Y2=1.065
cc_266 VPB N_A_619_368#_c_1393_n 0.0176924f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_267 VPB N_A_619_368#_c_1394_n 0.2116f $X=-0.19 $Y=1.66 $X2=0.265 $Y2=1.065
cc_268 VPB N_A_619_368#_c_1395_n 0.0744302f $X=-0.19 $Y=1.66 $X2=1.94 $Y2=1.975
cc_269 VPB N_A_619_368#_c_1396_n 0.0145869f $X=-0.19 $Y=1.66 $X2=1.94 $Y2=1.975
cc_270 VPB N_A_619_368#_c_1397_n 0.014206f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_271 VPB N_A_619_368#_c_1398_n 0.0107784f $X=-0.19 $Y=1.66 $X2=0.98 $Y2=1.065
cc_272 VPB N_A_619_368#_c_1399_n 0.014619f $X=-0.19 $Y=1.66 $X2=0.98 $Y2=0.9
cc_273 VPB N_A_619_368#_c_1400_n 0.0269955f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_274 VPB N_A_619_368#_c_1401_n 0.0580487f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_275 VPB N_A_619_368#_c_1402_n 0.0712756f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_276 VPB N_A_619_368#_c_1403_n 0.0122412f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_277 VPB N_A_619_368#_c_1375_n 0.0724498f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_278 VPB N_A_619_368#_c_1377_n 0.00775791f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_279 VPB N_A_619_368#_c_1378_n 0.0119549f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_280 VPB N_A_619_368#_c_1379_n 6.04262e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_281 VPB N_A_619_368#_c_1408_n 0.0089864f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_282 VPB N_A_619_368#_c_1409_n 0.0053114f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_283 VPB N_A_619_368#_c_1382_n 7.35442e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_284 VPB N_A_619_368#_c_1411_n 0.00813764f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_285 VPB N_A_619_368#_c_1383_n 0.00170471f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_286 VPB N_A_619_368#_c_1413_n 0.0402381f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_287 VPB N_A_619_368#_c_1414_n 0.0114469f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_288 VPB N_A_619_368#_c_1386_n 0.027905f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_289 VPB N_A_619_368#_c_1416_n 0.00113419f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_290 VPB N_A_2513_258#_c_1654_n 0.022667f $X=-0.19 $Y=1.66 $X2=1.07 $Y2=0.58
cc_291 VPB N_A_2513_258#_c_1655_n 0.0225716f $X=-0.19 $Y=1.66 $X2=1.07 $Y2=0.58
cc_292 VPB N_A_2513_258#_c_1646_n 0.00827326f $X=-0.19 $Y=1.66 $X2=0.17 $Y2=1.97
cc_293 VPB N_A_2513_258#_c_1657_n 0.0153617f $X=-0.19 $Y=1.66 $X2=0.275 $Y2=2.14
cc_294 VPB N_A_2513_258#_c_1647_n 0.00137888f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_295 VPB N_A_2513_258#_c_1652_n 0.0114667f $X=-0.19 $Y=1.66 $X2=1.94 $Y2=1.975
cc_296 VPB N_A_2513_258#_c_1660_n 0.00704454f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_297 VPB N_A_2067_74#_c_1768_n 0.0147748f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_298 VPB N_A_2067_74#_c_1769_n 0.0225675f $X=-0.19 $Y=1.66 $X2=0.445 $Y2=1.065
cc_299 VPB N_A_2067_74#_c_1770_n 0.0181269f $X=-0.19 $Y=1.66 $X2=0.98 $Y2=1.065
cc_300 VPB N_A_2067_74#_c_1751_n 8.19093e-19 $X=-0.19 $Y=1.66 $X2=1.94 $Y2=1.975
cc_301 VPB N_A_2067_74#_c_1772_n 0.0228091f $X=-0.19 $Y=1.66 $X2=1.94 $Y2=1.975
cc_302 VPB N_A_2067_74#_c_1754_n 9.13218e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_303 VPB N_A_2067_74#_c_1774_n 0.0247934f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_304 VPB N_A_2067_74#_c_1756_n 9.83765e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_305 VPB N_A_2067_74#_c_1776_n 0.0255479f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_306 VPB N_A_2067_74#_c_1777_n 0.0174677f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_307 VPB N_A_2067_74#_c_1778_n 0.00960239f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_308 VPB N_A_2067_74#_c_1779_n 0.0024355f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_309 VPB N_A_2067_74#_c_1780_n 0.0152136f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_310 VPB N_A_2067_74#_c_1781_n 0.0105124f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_311 VPB N_A_2067_74#_c_1782_n 0.00884139f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_312 VPB N_A_2067_74#_c_1765_n 0.0363227f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_313 VPB N_A_2067_74#_c_1784_n 0.006122f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_314 VPB N_A_2067_74#_c_1767_n 0.00248742f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_315 VPB N_A_3177_368#_c_1995_n 0.0163465f $X=-0.19 $Y=1.66 $X2=1.07 $Y2=0.9
cc_316 VPB N_A_3177_368#_c_1996_n 0.017358f $X=-0.19 $Y=1.66 $X2=0.265 $Y2=0.58
cc_317 VPB N_A_3177_368#_c_1991_n 0.0156856f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_318 VPB N_A_3177_368#_c_1994_n 0.0169257f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_319 VPB N_VPWR_c_2058_n 0.00918275f $X=-0.19 $Y=1.66 $X2=1.94 $Y2=2.055
cc_320 VPB N_VPWR_c_2059_n 0.012364f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_321 VPB N_VPWR_c_2060_n 0.00702644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_322 VPB N_VPWR_c_2061_n 0.0313096f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_323 VPB N_VPWR_c_2062_n 0.011131f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_324 VPB N_VPWR_c_2063_n 0.00538125f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_325 VPB N_VPWR_c_2064_n 0.00982859f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_326 VPB N_VPWR_c_2065_n 0.0127416f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_327 VPB N_VPWR_c_2066_n 0.0267817f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_328 VPB N_VPWR_c_2067_n 0.0157152f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_329 VPB N_VPWR_c_2068_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_330 VPB N_VPWR_c_2069_n 0.0644986f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_331 VPB N_VPWR_c_2070_n 0.020354f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_332 VPB N_VPWR_c_2071_n 0.00460249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_333 VPB N_VPWR_c_2072_n 0.0794449f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_334 VPB N_VPWR_c_2073_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_335 VPB N_VPWR_c_2074_n 0.0380992f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_336 VPB N_VPWR_c_2075_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_337 VPB N_VPWR_c_2076_n 0.0184862f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_338 VPB N_VPWR_c_2077_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_339 VPB N_VPWR_c_2078_n 0.0193973f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_340 VPB N_VPWR_c_2079_n 0.0448083f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_341 VPB N_VPWR_c_2080_n 0.0508863f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_342 VPB N_VPWR_c_2081_n 0.0227335f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_343 VPB N_VPWR_c_2082_n 0.0203698f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_344 VPB N_VPWR_c_2083_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_345 VPB N_VPWR_c_2084_n 0.00652596f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_346 VPB N_VPWR_c_2085_n 0.0214164f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_347 VPB N_VPWR_c_2086_n 0.0224449f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_348 VPB N_VPWR_c_2087_n 0.00763133f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_349 VPB N_VPWR_c_2088_n 0.00436868f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_350 VPB N_VPWR_c_2089_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_351 VPB N_VPWR_c_2057_n 0.159462f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_352 VPB N_A_304_464#_c_2260_n 0.00846251f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=0.58
cc_353 VPB N_A_304_464#_c_2257_n 0.0147808f $X=-0.19 $Y=1.66 $X2=0.17 $Y2=1.97
cc_354 VPB N_A_304_464#_c_2262_n 0.0121196f $X=-0.19 $Y=1.66 $X2=0.275 $Y2=2.14
cc_355 VPB N_A_304_464#_c_2263_n 0.00185789f $X=-0.19 $Y=1.66 $X2=0.3 $Y2=2.465
cc_356 VPB N_A_304_464#_c_2264_n 0.00699004f $X=-0.19 $Y=1.66 $X2=0.98 $Y2=1.065
cc_357 VPB N_A_304_464#_c_2265_n 0.0103043f $X=-0.19 $Y=1.66 $X2=0.98 $Y2=0.9
cc_358 VPB N_A_304_464#_c_2259_n 0.00306764f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_359 VPB N_A_1789_424#_c_2373_n 0.00227759f $X=-0.19 $Y=1.66 $X2=0.265
+ $Y2=0.58
cc_360 VPB N_A_1789_424#_c_2374_n 0.00672758f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_361 VPB N_A_1789_424#_c_2375_n 0.00171072f $X=-0.19 $Y=1.66 $X2=0.17 $Y2=1.23
cc_362 VPB N_A_1789_424#_c_2376_n 0.00407868f $X=-0.19 $Y=1.66 $X2=0.275
+ $Y2=2.465
cc_363 VPB N_A_1789_424#_c_2377_n 0.0102485f $X=-0.19 $Y=1.66 $X2=0.445
+ $Y2=1.065
cc_364 VPB N_A_2277_455#_c_2427_n 0.00753543f $X=-0.19 $Y=1.66 $X2=1.07 $Y2=0.58
cc_365 VPB N_A_2277_455#_c_2428_n 0.0147021f $X=-0.19 $Y=1.66 $X2=2.015 $Y2=2.64
cc_366 VPB N_A_2277_455#_c_2429_n 0.00404548f $X=-0.19 $Y=1.66 $X2=2.015
+ $Y2=2.64
cc_367 VPB N_A_2277_455#_c_2430_n 0.00587602f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=0.58
cc_368 VPB N_Q_N_c_2459_n 0.00408002f $X=-0.19 $Y=1.66 $X2=1.07 $Y2=0.58
cc_369 VPB N_Q_c_2490_n 0.00257348f $X=-0.19 $Y=1.66 $X2=1.07 $Y2=0.58
cc_370 VPB N_Q_c_2491_n 0.00198321f $X=-0.19 $Y=1.66 $X2=0.265 $Y2=0.58
cc_371 VPB N_Q_c_2487_n 0.00104928f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=0.58
cc_372 N_A_27_74#_c_373_n N_SCE_M1044_g 0.011453f $X=0.28 $Y=0.58 $X2=0 $Y2=0
cc_373 N_A_27_74#_c_374_n N_SCE_M1044_g 0.00547238f $X=0.17 $Y=1.97 $X2=0 $Y2=0
cc_374 N_A_27_74#_c_375_n N_SCE_M1044_g 0.0146918f $X=0.98 $Y=1.065 $X2=0 $Y2=0
cc_375 N_A_27_74#_c_376_n N_SCE_M1044_g 0.0176381f $X=0.98 $Y=1.065 $X2=0 $Y2=0
cc_376 N_A_27_74#_c_377_n N_SCE_M1044_g 0.00812645f $X=0.265 $Y=1.065 $X2=0
+ $Y2=0
cc_377 N_A_27_74#_c_378_n N_SCE_M1044_g 0.0119253f $X=0.98 $Y=0.9 $X2=0 $Y2=0
cc_378 N_A_27_74#_c_374_n N_SCE_c_458_n 0.00413205f $X=0.17 $Y=1.97 $X2=0 $Y2=0
cc_379 N_A_27_74#_c_381_n N_SCE_c_458_n 5.33641e-19 $X=0.3 $Y=2.465 $X2=0 $Y2=0
cc_380 N_A_27_74#_c_382_n N_SCE_c_458_n 0.0131315f $X=1.775 $Y=2.055 $X2=0 $Y2=0
cc_381 N_A_27_74#_c_383_n N_SCE_c_458_n 0.00446031f $X=0.275 $Y=2.055 $X2=0
+ $Y2=0
cc_382 N_A_27_74#_c_381_n N_SCE_c_459_n 0.0137466f $X=0.3 $Y=2.465 $X2=0 $Y2=0
cc_383 N_A_27_74#_c_381_n N_SCE_c_460_n 4.83056e-19 $X=0.3 $Y=2.465 $X2=0 $Y2=0
cc_384 N_A_27_74#_c_382_n N_SCE_c_460_n 0.0162959f $X=1.775 $Y=2.055 $X2=0 $Y2=0
cc_385 N_A_27_74#_c_381_n N_SCE_c_461_n 4.6382e-19 $X=0.3 $Y=2.465 $X2=0 $Y2=0
cc_386 N_A_27_74#_c_379_n N_SCE_c_451_n 0.00140892f $X=2.015 $Y=2.245 $X2=0
+ $Y2=0
cc_387 N_A_27_74#_c_382_n N_SCE_c_451_n 0.0272489f $X=1.775 $Y=2.055 $X2=0 $Y2=0
cc_388 N_A_27_74#_c_384_n N_SCE_c_451_n 0.0194177f $X=1.94 $Y=1.975 $X2=0 $Y2=0
cc_389 N_A_27_74#_c_374_n N_SCE_c_452_n 0.0317203f $X=0.17 $Y=1.97 $X2=0 $Y2=0
cc_390 N_A_27_74#_c_375_n N_SCE_c_452_n 0.0563109f $X=0.98 $Y=1.065 $X2=0 $Y2=0
cc_391 N_A_27_74#_c_376_n N_SCE_c_452_n 0.00277723f $X=0.98 $Y=1.065 $X2=0 $Y2=0
cc_392 N_A_27_74#_c_382_n N_SCE_c_452_n 0.0460993f $X=1.775 $Y=2.055 $X2=0 $Y2=0
cc_393 N_A_27_74#_c_377_n N_SCE_c_452_n 0.00161902f $X=0.265 $Y=1.065 $X2=0
+ $Y2=0
cc_394 N_A_27_74#_c_383_n N_SCE_c_452_n 0.00328312f $X=0.275 $Y=2.055 $X2=0
+ $Y2=0
cc_395 N_A_27_74#_c_374_n N_SCE_c_453_n 0.00871649f $X=0.17 $Y=1.97 $X2=0 $Y2=0
cc_396 N_A_27_74#_c_375_n N_SCE_c_453_n 0.00180003f $X=0.98 $Y=1.065 $X2=0 $Y2=0
cc_397 N_A_27_74#_c_376_n N_SCE_c_453_n 0.0152994f $X=0.98 $Y=1.065 $X2=0 $Y2=0
cc_398 N_A_27_74#_c_382_n N_SCE_c_453_n 0.00313888f $X=1.775 $Y=2.055 $X2=0
+ $Y2=0
cc_399 N_A_27_74#_c_377_n N_SCE_c_453_n 2.0611e-19 $X=0.265 $Y=1.065 $X2=0 $Y2=0
cc_400 N_A_27_74#_c_383_n N_SCE_c_453_n 7.36532e-19 $X=0.275 $Y=2.055 $X2=0
+ $Y2=0
cc_401 N_A_27_74#_c_379_n N_SCE_c_455_n 0.00776428f $X=2.015 $Y=2.245 $X2=0
+ $Y2=0
cc_402 N_A_27_74#_c_379_n N_D_c_535_n 0.0224177f $X=2.015 $Y=2.245 $X2=0 $Y2=0
cc_403 N_A_27_74#_c_382_n N_D_c_535_n 0.0170798f $X=1.775 $Y=2.055 $X2=0 $Y2=0
cc_404 N_A_27_74#_c_384_n N_D_c_535_n 0.00116992f $X=1.94 $Y=1.975 $X2=0 $Y2=0
cc_405 N_A_27_74#_c_379_n N_D_c_541_n 0.0233104f $X=2.015 $Y=2.245 $X2=0 $Y2=0
cc_406 N_A_27_74#_c_375_n D 0.0201653f $X=0.98 $Y=1.065 $X2=0 $Y2=0
cc_407 N_A_27_74#_c_376_n D 4.18339e-19 $X=0.98 $Y=1.065 $X2=0 $Y2=0
cc_408 N_A_27_74#_c_378_n D 0.00225318f $X=0.98 $Y=0.9 $X2=0 $Y2=0
cc_409 N_A_27_74#_c_375_n N_D_c_538_n 0.00120526f $X=0.98 $Y=1.065 $X2=0 $Y2=0
cc_410 N_A_27_74#_c_376_n N_D_c_538_n 0.0255527f $X=0.98 $Y=1.065 $X2=0 $Y2=0
cc_411 N_A_27_74#_c_378_n N_D_c_539_n 0.0255527f $X=0.98 $Y=0.9 $X2=0 $Y2=0
cc_412 N_A_27_74#_c_379_n N_SCD_c_590_n 0.0383399f $X=2.015 $Y=2.245 $X2=0 $Y2=0
cc_413 N_A_27_74#_c_379_n N_SCD_c_592_n 0.0231074f $X=2.015 $Y=2.245 $X2=0 $Y2=0
cc_414 N_A_27_74#_c_384_n N_SCD_c_592_n 0.00128345f $X=1.94 $Y=1.975 $X2=0 $Y2=0
cc_415 N_A_27_74#_c_381_n N_VPWR_c_2058_n 0.0268536f $X=0.3 $Y=2.465 $X2=0 $Y2=0
cc_416 N_A_27_74#_c_382_n N_VPWR_c_2058_n 0.0275301f $X=1.775 $Y=2.055 $X2=0
+ $Y2=0
cc_417 N_A_27_74#_c_379_n N_VPWR_c_2059_n 0.00149447f $X=2.015 $Y=2.245 $X2=0
+ $Y2=0
cc_418 N_A_27_74#_c_381_n N_VPWR_c_2078_n 0.0168249f $X=0.3 $Y=2.465 $X2=0 $Y2=0
cc_419 N_A_27_74#_c_379_n N_VPWR_c_2079_n 0.00445602f $X=2.015 $Y=2.245 $X2=0
+ $Y2=0
cc_420 N_A_27_74#_c_379_n N_VPWR_c_2057_n 0.00456581f $X=2.015 $Y=2.245 $X2=0
+ $Y2=0
cc_421 N_A_27_74#_c_381_n N_VPWR_c_2057_n 0.0138933f $X=0.3 $Y=2.465 $X2=0 $Y2=0
cc_422 N_A_27_74#_c_379_n N_A_304_464#_c_2260_n 0.00939385f $X=2.015 $Y=2.245
+ $X2=0 $Y2=0
cc_423 N_A_27_74#_c_384_n N_A_304_464#_c_2260_n 0.0107144f $X=1.94 $Y=1.975
+ $X2=0 $Y2=0
cc_424 N_A_27_74#_c_379_n N_A_304_464#_c_2257_n 0.00187783f $X=2.015 $Y=2.245
+ $X2=0 $Y2=0
cc_425 N_A_27_74#_c_384_n N_A_304_464#_c_2257_n 0.0128835f $X=1.94 $Y=1.975
+ $X2=0 $Y2=0
cc_426 N_A_27_74#_c_379_n N_A_304_464#_c_2264_n 0.0213981f $X=2.015 $Y=2.245
+ $X2=0 $Y2=0
cc_427 N_A_27_74#_c_382_n N_A_304_464#_c_2264_n 0.0225954f $X=1.775 $Y=2.055
+ $X2=0 $Y2=0
cc_428 N_A_27_74#_c_384_n N_A_304_464#_c_2264_n 0.0150832f $X=1.94 $Y=1.975
+ $X2=0 $Y2=0
cc_429 N_A_27_74#_c_373_n N_VGND_c_2517_n 0.0133638f $X=0.28 $Y=0.58 $X2=0 $Y2=0
cc_430 N_A_27_74#_c_375_n N_VGND_c_2517_n 0.0255027f $X=0.98 $Y=1.065 $X2=0
+ $Y2=0
cc_431 N_A_27_74#_c_376_n N_VGND_c_2517_n 0.0038848f $X=0.98 $Y=1.065 $X2=0
+ $Y2=0
cc_432 N_A_27_74#_c_378_n N_VGND_c_2517_n 0.00981126f $X=0.98 $Y=0.9 $X2=0 $Y2=0
cc_433 N_A_27_74#_c_378_n N_VGND_c_2529_n 0.00383152f $X=0.98 $Y=0.9 $X2=0 $Y2=0
cc_434 N_A_27_74#_c_373_n N_VGND_c_2539_n 0.0159025f $X=0.28 $Y=0.58 $X2=0 $Y2=0
cc_435 N_A_27_74#_c_373_n N_VGND_c_2550_n 0.0131064f $X=0.28 $Y=0.58 $X2=0 $Y2=0
cc_436 N_A_27_74#_c_378_n N_VGND_c_2550_n 0.0075725f $X=0.98 $Y=0.9 $X2=0 $Y2=0
cc_437 N_SCE_c_451_n N_D_c_534_n 0.00445951f $X=1.965 $Y=1.485 $X2=-0.19
+ $Y2=-0.245
cc_438 N_SCE_c_453_n N_D_c_534_n 0.00828205f $X=0.92 $Y=1.635 $X2=-0.19
+ $Y2=-0.245
cc_439 N_SCE_c_451_n N_D_c_535_n 0.00429479f $X=1.965 $Y=1.485 $X2=0 $Y2=0
cc_440 N_SCE_c_453_n N_D_c_535_n 0.0172195f $X=0.92 $Y=1.635 $X2=0 $Y2=0
cc_441 N_SCE_c_454_n N_D_c_535_n 0.0014191f $X=1.085 $Y=1.6 $X2=0 $Y2=0
cc_442 N_SCE_c_460_n N_D_c_541_n 0.0172195f $X=1.025 $Y=2.155 $X2=0 $Y2=0
cc_443 N_SCE_c_461_n N_D_c_541_n 0.0370053f $X=1.025 $Y=2.245 $X2=0 $Y2=0
cc_444 N_SCE_c_451_n N_D_c_536_n 0.00572304f $X=1.965 $Y=1.485 $X2=0 $Y2=0
cc_445 N_SCE_c_455_n N_D_c_536_n 0.00964743f $X=2.13 $Y=1.065 $X2=0 $Y2=0
cc_446 N_SCE_c_456_n N_D_c_536_n 9.50384e-19 $X=2.13 $Y=1.065 $X2=0 $Y2=0
cc_447 N_SCE_c_451_n D 0.0324073f $X=1.965 $Y=1.485 $X2=0 $Y2=0
cc_448 N_SCE_c_455_n D 0.00220222f $X=2.13 $Y=1.065 $X2=0 $Y2=0
cc_449 N_SCE_c_456_n D 0.0265741f $X=2.13 $Y=1.065 $X2=0 $Y2=0
cc_450 N_SCE_c_457_n D 0.00241363f $X=2.22 $Y=0.9 $X2=0 $Y2=0
cc_451 N_SCE_c_451_n N_D_c_538_n 0.00126891f $X=1.965 $Y=1.485 $X2=0 $Y2=0
cc_452 N_SCE_c_455_n N_D_c_538_n 0.0170267f $X=2.13 $Y=1.065 $X2=0 $Y2=0
cc_453 N_SCE_c_456_n N_D_c_538_n 3.60471e-19 $X=2.13 $Y=1.065 $X2=0 $Y2=0
cc_454 N_SCE_c_455_n N_SCD_c_592_n 0.00941785f $X=2.13 $Y=1.065 $X2=0 $Y2=0
cc_455 N_SCE_c_457_n N_SCD_M1018_g 0.0341499f $X=2.22 $Y=0.9 $X2=0 $Y2=0
cc_456 N_SCE_c_455_n N_SCD_c_584_n 0.0341499f $X=2.13 $Y=1.065 $X2=0 $Y2=0
cc_457 N_SCE_c_455_n SCD 5.07628e-19 $X=2.13 $Y=1.065 $X2=0 $Y2=0
cc_458 N_SCE_c_459_n N_VPWR_c_2058_n 0.00679357f $X=0.525 $Y=2.245 $X2=0 $Y2=0
cc_459 N_SCE_c_461_n N_VPWR_c_2058_n 0.0158802f $X=1.025 $Y=2.245 $X2=0 $Y2=0
cc_460 N_SCE_c_459_n N_VPWR_c_2078_n 0.00445602f $X=0.525 $Y=2.245 $X2=0 $Y2=0
cc_461 N_SCE_c_461_n N_VPWR_c_2079_n 0.00413917f $X=1.025 $Y=2.245 $X2=0 $Y2=0
cc_462 N_SCE_c_459_n N_VPWR_c_2057_n 0.00860937f $X=0.525 $Y=2.245 $X2=0 $Y2=0
cc_463 N_SCE_c_461_n N_VPWR_c_2057_n 0.00817532f $X=1.025 $Y=2.245 $X2=0 $Y2=0
cc_464 N_SCE_c_451_n N_A_304_464#_c_2257_n 0.0129498f $X=1.965 $Y=1.485 $X2=0
+ $Y2=0
cc_465 N_SCE_c_455_n N_A_304_464#_c_2257_n 0.0142897f $X=2.13 $Y=1.065 $X2=0
+ $Y2=0
cc_466 N_SCE_c_456_n N_A_304_464#_c_2257_n 0.0356688f $X=2.13 $Y=1.065 $X2=0
+ $Y2=0
cc_467 N_SCE_c_457_n N_A_304_464#_c_2257_n 0.00470988f $X=2.22 $Y=0.9 $X2=0
+ $Y2=0
cc_468 N_SCE_c_461_n N_A_304_464#_c_2264_n 0.00192751f $X=1.025 $Y=2.245 $X2=0
+ $Y2=0
cc_469 N_SCE_c_455_n N_A_304_464#_c_2279_n 0.00233988f $X=2.13 $Y=1.065 $X2=0
+ $Y2=0
cc_470 N_SCE_c_456_n N_A_304_464#_c_2279_n 0.0260811f $X=2.13 $Y=1.065 $X2=0
+ $Y2=0
cc_471 N_SCE_c_457_n N_A_304_464#_c_2279_n 0.0150729f $X=2.22 $Y=0.9 $X2=0 $Y2=0
cc_472 N_SCE_M1044_g N_VGND_c_2517_n 0.00540268f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_473 N_SCE_c_457_n N_VGND_c_2518_n 0.00144244f $X=2.22 $Y=0.9 $X2=0 $Y2=0
cc_474 N_SCE_c_457_n N_VGND_c_2529_n 0.00314477f $X=2.22 $Y=0.9 $X2=0 $Y2=0
cc_475 N_SCE_M1044_g N_VGND_c_2539_n 0.00434272f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_476 N_SCE_M1044_g N_VGND_c_2550_n 0.00825006f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_477 N_SCE_c_457_n N_VGND_c_2550_n 0.00395526f $X=2.22 $Y=0.9 $X2=0 $Y2=0
cc_478 N_D_c_541_n N_VPWR_c_2058_n 0.00247596f $X=1.445 $Y=2.245 $X2=0 $Y2=0
cc_479 N_D_c_541_n N_VPWR_c_2079_n 0.00445602f $X=1.445 $Y=2.245 $X2=0 $Y2=0
cc_480 N_D_c_541_n N_VPWR_c_2057_n 0.00859212f $X=1.445 $Y=2.245 $X2=0 $Y2=0
cc_481 D N_A_304_464#_M1036_d 0.00795735f $X=1.595 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_482 D N_A_304_464#_c_2257_n 0.00450433f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_483 N_D_c_541_n N_A_304_464#_c_2264_n 0.0227408f $X=1.445 $Y=2.245 $X2=0
+ $Y2=0
cc_484 D N_A_304_464#_c_2279_n 0.0246293f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_485 N_D_c_539_n N_A_304_464#_c_2279_n 0.00242613f $X=1.55 $Y=0.9 $X2=0 $Y2=0
cc_486 D N_VGND_c_2517_n 0.0100693f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_487 N_D_c_539_n N_VGND_c_2517_n 0.00163952f $X=1.55 $Y=0.9 $X2=0 $Y2=0
cc_488 D N_VGND_c_2529_n 0.0118305f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_489 N_D_c_539_n N_VGND_c_2529_n 0.00304348f $X=1.55 $Y=0.9 $X2=0 $Y2=0
cc_490 D N_VGND_c_2550_n 0.0134831f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_491 N_D_c_539_n N_VGND_c_2550_n 0.00375359f $X=1.55 $Y=0.9 $X2=0 $Y2=0
cc_492 N_SCD_c_584_n N_CLK_c_635_n 0.0217622f $X=2.925 $Y=1.41 $X2=-0.19
+ $Y2=-0.245
cc_493 N_SCD_c_585_n N_CLK_c_635_n 0.00582176f $X=2.79 $Y=1.81 $X2=-0.19
+ $Y2=-0.245
cc_494 SCD N_CLK_c_635_n 0.0026011f $X=3.035 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_495 N_SCD_c_588_n N_CLK_c_636_n 0.00312834f $X=2.97 $Y=1.115 $X2=0 $Y2=0
cc_496 N_SCD_M1018_g N_A_619_368#_c_1381_n 0.00509351f $X=2.79 $Y=0.58 $X2=0
+ $Y2=0
cc_497 N_SCD_c_584_n N_A_619_368#_c_1382_n 8.82978e-19 $X=2.925 $Y=1.41 $X2=0
+ $Y2=0
cc_498 N_SCD_c_585_n N_A_619_368#_c_1382_n 0.00115574f $X=2.79 $Y=1.81 $X2=0
+ $Y2=0
cc_499 N_SCD_c_589_n N_A_619_368#_c_1414_n 9.69705e-19 $X=2.435 $Y=2.155 $X2=0
+ $Y2=0
cc_500 N_SCD_c_585_n N_A_619_368#_c_1414_n 0.00226703f $X=2.79 $Y=1.81 $X2=0
+ $Y2=0
cc_501 N_SCD_c_586_n N_A_619_368#_c_1414_n 0.0015818f $X=2.925 $Y=1.62 $X2=0
+ $Y2=0
cc_502 SCD N_A_619_368#_c_1414_n 0.011212f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_503 SCD N_A_619_368#_c_1385_n 0.0526519f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_504 N_SCD_c_588_n N_A_619_368#_c_1385_n 4.41357e-19 $X=2.97 $Y=1.115 $X2=0
+ $Y2=0
cc_505 N_SCD_c_590_n N_VPWR_c_2059_n 0.010659f $X=2.435 $Y=2.245 $X2=0 $Y2=0
cc_506 N_SCD_c_591_n N_VPWR_c_2059_n 5.29465e-19 $X=2.715 $Y=1.885 $X2=0 $Y2=0
cc_507 N_SCD_c_590_n N_VPWR_c_2079_n 0.00413917f $X=2.435 $Y=2.245 $X2=0 $Y2=0
cc_508 N_SCD_c_590_n N_VPWR_c_2057_n 0.00416516f $X=2.435 $Y=2.245 $X2=0 $Y2=0
cc_509 N_SCD_c_590_n N_A_304_464#_c_2260_n 0.0109694f $X=2.435 $Y=2.245 $X2=0
+ $Y2=0
cc_510 N_SCD_c_589_n N_A_304_464#_c_2257_n 0.0065726f $X=2.435 $Y=2.155 $X2=0
+ $Y2=0
cc_511 N_SCD_c_590_n N_A_304_464#_c_2257_n 0.00577906f $X=2.435 $Y=2.245 $X2=0
+ $Y2=0
cc_512 N_SCD_c_591_n N_A_304_464#_c_2257_n 0.00921263f $X=2.715 $Y=1.885 $X2=0
+ $Y2=0
cc_513 N_SCD_c_592_n N_A_304_464#_c_2257_n 0.00395981f $X=2.525 $Y=1.885 $X2=0
+ $Y2=0
cc_514 N_SCD_M1018_g N_A_304_464#_c_2257_n 0.0167474f $X=2.79 $Y=0.58 $X2=0
+ $Y2=0
cc_515 SCD N_A_304_464#_c_2257_n 0.0511176f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_516 N_SCD_c_591_n N_A_304_464#_c_2262_n 0.00737458f $X=2.715 $Y=1.885 $X2=0
+ $Y2=0
cc_517 N_SCD_c_586_n N_A_304_464#_c_2262_n 0.00511032f $X=2.925 $Y=1.62 $X2=0
+ $Y2=0
cc_518 N_SCD_c_590_n N_A_304_464#_c_2264_n 0.00176083f $X=2.435 $Y=2.245 $X2=0
+ $Y2=0
cc_519 N_SCD_M1018_g N_A_304_464#_c_2279_n 0.00177354f $X=2.79 $Y=0.58 $X2=0
+ $Y2=0
cc_520 N_SCD_c_590_n N_A_304_464#_c_2298_n 0.00583307f $X=2.435 $Y=2.245 $X2=0
+ $Y2=0
cc_521 N_SCD_M1018_g N_VGND_c_2518_n 0.0117409f $X=2.79 $Y=0.58 $X2=0 $Y2=0
cc_522 SCD N_VGND_c_2518_n 0.026063f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_523 N_SCD_c_588_n N_VGND_c_2518_n 0.0070747f $X=2.97 $Y=1.115 $X2=0 $Y2=0
cc_524 N_SCD_M1018_g N_VGND_c_2529_n 0.00383152f $X=2.79 $Y=0.58 $X2=0 $Y2=0
cc_525 N_SCD_M1018_g N_VGND_c_2550_n 0.0075725f $X=2.79 $Y=0.58 $X2=0 $Y2=0
cc_526 N_CLK_c_635_n N_A_619_368#_M1033_g 0.0207024f $X=3.465 $Y=1.765 $X2=0
+ $Y2=0
cc_527 N_CLK_c_636_n N_A_619_368#_M1033_g 0.0188406f $X=3.78 $Y=1.22 $X2=0 $Y2=0
cc_528 CLK N_A_619_368#_M1033_g 0.0070177f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_529 N_CLK_c_635_n N_A_619_368#_c_1387_n 0.0119921f $X=3.465 $Y=1.765 $X2=0
+ $Y2=0
cc_530 N_CLK_c_635_n N_A_619_368#_c_1377_n 0.0043393f $X=3.465 $Y=1.765 $X2=0
+ $Y2=0
cc_531 N_CLK_c_636_n N_A_619_368#_c_1381_n 6.69491e-19 $X=3.78 $Y=1.22 $X2=0
+ $Y2=0
cc_532 N_CLK_c_635_n N_A_619_368#_c_1382_n 0.0263169f $X=3.465 $Y=1.765 $X2=0
+ $Y2=0
cc_533 N_CLK_c_636_n N_A_619_368#_c_1382_n 0.00417982f $X=3.78 $Y=1.22 $X2=0
+ $Y2=0
cc_534 CLK N_A_619_368#_c_1382_n 0.0273382f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_535 N_CLK_c_635_n N_A_619_368#_c_1411_n 0.0121116f $X=3.465 $Y=1.765 $X2=0
+ $Y2=0
cc_536 CLK N_A_619_368#_c_1411_n 0.0289811f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_537 CLK N_A_619_368#_c_1383_n 0.0147056f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_538 N_CLK_c_635_n N_A_619_368#_c_1414_n 0.0140111f $X=3.465 $Y=1.765 $X2=0
+ $Y2=0
cc_539 N_CLK_c_635_n N_A_619_368#_c_1385_n 0.00438848f $X=3.465 $Y=1.765 $X2=0
+ $Y2=0
cc_540 N_CLK_c_635_n N_VPWR_c_2059_n 0.0110636f $X=3.465 $Y=1.765 $X2=0 $Y2=0
cc_541 N_CLK_c_635_n N_VPWR_c_2085_n 0.00413917f $X=3.465 $Y=1.765 $X2=0 $Y2=0
cc_542 N_CLK_c_635_n N_VPWR_c_2086_n 0.0233922f $X=3.465 $Y=1.765 $X2=0 $Y2=0
cc_543 N_CLK_c_635_n N_VPWR_c_2057_n 0.00419897f $X=3.465 $Y=1.765 $X2=0 $Y2=0
cc_544 N_CLK_c_635_n N_A_304_464#_c_2262_n 0.0142456f $X=3.465 $Y=1.765 $X2=0
+ $Y2=0
cc_545 N_CLK_c_635_n N_A_304_464#_c_2300_n 0.00453754f $X=3.465 $Y=1.765 $X2=0
+ $Y2=0
cc_546 N_CLK_c_636_n N_VGND_c_2518_n 0.00224794f $X=3.78 $Y=1.22 $X2=0 $Y2=0
cc_547 N_CLK_c_635_n N_VGND_c_2519_n 8.35753e-19 $X=3.465 $Y=1.765 $X2=0 $Y2=0
cc_548 N_CLK_c_636_n N_VGND_c_2519_n 0.0118636f $X=3.78 $Y=1.22 $X2=0 $Y2=0
cc_549 CLK N_VGND_c_2519_n 0.0254134f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_550 N_CLK_c_636_n N_VGND_c_2540_n 0.00383152f $X=3.78 $Y=1.22 $X2=0 $Y2=0
cc_551 N_CLK_c_636_n N_VGND_c_2550_n 0.00762539f $X=3.78 $Y=1.22 $X2=0 $Y2=0
cc_552 N_A_871_74#_c_703_n N_A_1252_376#_c_947_n 0.00261463f $X=6.155 $Y=2.905
+ $X2=0 $Y2=0
cc_553 N_A_871_74#_c_704_n N_A_1252_376#_c_947_n 0.00788258f $X=7.155 $Y=2.25
+ $X2=0 $Y2=0
cc_554 N_A_871_74#_c_712_n N_A_1252_376#_c_947_n 0.00252926f $X=6.187 $Y=2.25
+ $X2=0 $Y2=0
cc_555 N_A_871_74#_c_704_n N_A_1252_376#_c_948_n 0.0134562f $X=7.155 $Y=2.25
+ $X2=0 $Y2=0
cc_556 N_A_871_74#_M1027_g N_A_1252_376#_c_941_n 0.0214745f $X=6.295 $Y=0.615
+ $X2=0 $Y2=0
cc_557 N_A_871_74#_c_696_n N_A_1252_376#_c_949_n 7.74578e-19 $X=5.395 $Y=1.96
+ $X2=0 $Y2=0
cc_558 N_A_871_74#_c_683_n N_A_1252_376#_c_949_n 0.0157175f $X=6.185 $Y=1.135
+ $X2=0 $Y2=0
cc_559 N_A_871_74#_c_684_n N_A_1252_376#_c_949_n 0.00703758f $X=6.185 $Y=1.135
+ $X2=0 $Y2=0
cc_560 N_A_871_74#_c_704_n N_A_1252_376#_c_949_n 0.00686883f $X=7.155 $Y=2.25
+ $X2=0 $Y2=0
cc_561 N_A_871_74#_c_712_n N_A_1252_376#_c_949_n 0.00134941f $X=6.187 $Y=2.25
+ $X2=0 $Y2=0
cc_562 N_A_871_74#_c_683_n N_A_1252_376#_c_950_n 0.0123703f $X=6.185 $Y=1.135
+ $X2=0 $Y2=0
cc_563 N_A_871_74#_c_704_n N_A_1252_376#_c_950_n 0.053889f $X=7.155 $Y=2.25
+ $X2=0 $Y2=0
cc_564 N_A_871_74#_c_683_n N_A_1252_376#_c_951_n 0.00209505f $X=6.185 $Y=1.135
+ $X2=0 $Y2=0
cc_565 N_A_871_74#_c_706_n N_A_1252_376#_c_952_n 0.0227138f $X=7.995 $Y=2.99
+ $X2=0 $Y2=0
cc_566 N_A_871_74#_c_708_n N_A_1252_376#_c_952_n 0.0325868f $X=8.08 $Y=2.905
+ $X2=0 $Y2=0
cc_567 N_A_871_74#_c_704_n N_A_1252_376#_c_953_n 0.0128128f $X=7.155 $Y=2.25
+ $X2=0 $Y2=0
cc_568 N_A_871_74#_c_708_n N_A_1252_376#_c_953_n 0.00321202f $X=8.08 $Y=2.905
+ $X2=0 $Y2=0
cc_569 N_A_871_74#_c_710_n N_A_1252_376#_c_953_n 0.0081107f $X=8.165 $Y=2.135
+ $X2=0 $Y2=0
cc_570 N_A_871_74#_c_683_n N_A_1252_376#_c_945_n 0.00205641f $X=6.185 $Y=1.135
+ $X2=0 $Y2=0
cc_571 N_A_871_74#_c_684_n N_A_1252_376#_c_946_n 0.0337032f $X=6.185 $Y=1.135
+ $X2=0 $Y2=0
cc_572 N_A_871_74#_c_679_n N_A_1069_81#_M1019_d 4.5412e-19 $X=5.39 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_573 N_A_871_74#_c_689_n N_A_1069_81#_M1019_d 0.00650998f $X=5.395 $Y=1.29
+ $X2=-0.19 $Y2=-0.245
cc_574 N_A_871_74#_c_704_n N_A_1069_81#_c_1053_n 0.0040112f $X=7.155 $Y=2.25
+ $X2=0 $Y2=0
cc_575 N_A_871_74#_c_705_n N_A_1069_81#_c_1053_n 0.0115606f $X=7.24 $Y=2.905
+ $X2=0 $Y2=0
cc_576 N_A_871_74#_c_706_n N_A_1069_81#_c_1053_n 0.00388945f $X=7.995 $Y=2.99
+ $X2=0 $Y2=0
cc_577 N_A_871_74#_c_708_n N_A_1069_81#_c_1053_n 6.39854e-19 $X=8.08 $Y=2.905
+ $X2=0 $Y2=0
cc_578 N_A_871_74#_c_690_n N_A_1069_81#_c_1035_n 0.00918793f $X=10.38 $Y=1.365
+ $X2=0 $Y2=0
cc_579 N_A_871_74#_c_690_n N_A_1069_81#_c_1036_n 0.00550305f $X=10.38 $Y=1.365
+ $X2=0 $Y2=0
cc_580 N_A_871_74#_c_690_n N_A_1069_81#_c_1037_n 0.00827881f $X=10.38 $Y=1.365
+ $X2=0 $Y2=0
cc_581 N_A_871_74#_M1032_g N_A_1069_81#_M1009_g 0.0112306f $X=10.26 $Y=0.69
+ $X2=0 $Y2=0
cc_582 N_A_871_74#_c_687_n N_A_1069_81#_M1009_g 6.92746e-19 $X=10.545 $Y=1.365
+ $X2=0 $Y2=0
cc_583 N_A_871_74#_c_690_n N_A_1069_81#_c_1039_n 0.00404676f $X=10.38 $Y=1.365
+ $X2=0 $Y2=0
cc_584 N_A_871_74#_c_675_n N_A_1069_81#_c_1041_n 0.0180937f $X=10.835 $Y=1.41
+ $X2=0 $Y2=0
cc_585 N_A_871_74#_c_690_n N_A_1069_81#_c_1041_n 0.00373591f $X=10.38 $Y=1.365
+ $X2=0 $Y2=0
cc_586 N_A_871_74#_c_669_n N_A_1069_81#_c_1074_n 0.00361747f $X=6.02 $Y=1.365
+ $X2=0 $Y2=0
cc_587 N_A_871_74#_M1027_g N_A_1069_81#_c_1074_n 0.021861f $X=6.295 $Y=0.615
+ $X2=0 $Y2=0
cc_588 N_A_871_74#_c_683_n N_A_1069_81#_c_1074_n 0.0166876f $X=6.185 $Y=1.135
+ $X2=0 $Y2=0
cc_589 N_A_871_74#_c_684_n N_A_1069_81#_c_1074_n 0.00318891f $X=6.185 $Y=1.135
+ $X2=0 $Y2=0
cc_590 N_A_871_74#_c_689_n N_A_1069_81#_c_1078_n 0.0268483f $X=5.395 $Y=1.29
+ $X2=0 $Y2=0
cc_591 N_A_871_74#_M1027_g N_A_1069_81#_c_1042_n 0.00554569f $X=6.295 $Y=0.615
+ $X2=0 $Y2=0
cc_592 N_A_871_74#_c_683_n N_A_1069_81#_c_1042_n 0.0310926f $X=6.185 $Y=1.135
+ $X2=0 $Y2=0
cc_593 N_A_871_74#_c_683_n N_A_1069_81#_c_1044_n 0.0140103f $X=6.185 $Y=1.135
+ $X2=0 $Y2=0
cc_594 N_A_871_74#_c_684_n N_A_1069_81#_c_1044_n 0.00181486f $X=6.185 $Y=1.135
+ $X2=0 $Y2=0
cc_595 N_A_871_74#_c_704_n N_A_1069_81#_c_1044_n 0.00555233f $X=7.155 $Y=2.25
+ $X2=0 $Y2=0
cc_596 N_A_871_74#_c_686_n N_A_1069_81#_c_1046_n 0.00180199f $X=8.565 $Y=1.43
+ $X2=0 $Y2=0
cc_597 N_A_871_74#_c_686_n N_A_1069_81#_c_1047_n 0.0140773f $X=8.565 $Y=1.43
+ $X2=0 $Y2=0
cc_598 N_A_871_74#_c_690_n N_A_1069_81#_c_1047_n 0.0208175f $X=10.38 $Y=1.365
+ $X2=0 $Y2=0
cc_599 N_A_871_74#_c_686_n N_A_1069_81#_c_1048_n 8.79449e-19 $X=8.565 $Y=1.43
+ $X2=0 $Y2=0
cc_600 N_A_871_74#_c_690_n N_A_1069_81#_c_1048_n 0.0141435f $X=10.38 $Y=1.365
+ $X2=0 $Y2=0
cc_601 N_A_871_74#_c_693_n N_A_1069_81#_c_1058_n 0.00240683f $X=5.43 $Y=2.24
+ $X2=0 $Y2=0
cc_602 N_A_871_74#_c_698_n N_A_1069_81#_c_1058_n 0.0238882f $X=6.07 $Y=2.99
+ $X2=0 $Y2=0
cc_603 N_A_871_74#_c_681_n N_A_1069_81#_c_1058_n 9.31843e-19 $X=5.395 $Y=1.455
+ $X2=0 $Y2=0
cc_604 N_A_871_74#_c_703_n N_A_1069_81#_c_1058_n 0.0296994f $X=6.155 $Y=2.905
+ $X2=0 $Y2=0
cc_605 N_A_871_74#_c_692_n N_A_1069_81#_c_1049_n 0.00603316f $X=5.43 $Y=2.15
+ $X2=0 $Y2=0
cc_606 N_A_871_74#_c_693_n N_A_1069_81#_c_1049_n 4.06672e-19 $X=5.43 $Y=2.24
+ $X2=0 $Y2=0
cc_607 N_A_871_74#_c_669_n N_A_1069_81#_c_1049_n 0.0145736f $X=6.02 $Y=1.365
+ $X2=0 $Y2=0
cc_608 N_A_871_74#_M1027_g N_A_1069_81#_c_1049_n 0.00324964f $X=6.295 $Y=0.615
+ $X2=0 $Y2=0
cc_609 N_A_871_74#_c_682_n N_A_1069_81#_c_1049_n 0.00788192f $X=5.395 $Y=1.455
+ $X2=0 $Y2=0
cc_610 N_A_871_74#_c_683_n N_A_1069_81#_c_1049_n 0.0890046f $X=6.185 $Y=1.135
+ $X2=0 $Y2=0
cc_611 N_A_871_74#_c_684_n N_A_1069_81#_c_1049_n 0.00856636f $X=6.185 $Y=1.135
+ $X2=0 $Y2=0
cc_612 N_A_871_74#_c_689_n N_A_1069_81#_c_1049_n 0.0864367f $X=5.395 $Y=1.29
+ $X2=0 $Y2=0
cc_613 N_A_871_74#_c_712_n N_A_1069_81#_c_1049_n 0.0138873f $X=6.187 $Y=2.25
+ $X2=0 $Y2=0
cc_614 N_A_871_74#_c_710_n N_SET_B_c_1229_n 0.00481956f $X=8.165 $Y=2.135 $X2=0
+ $Y2=0
cc_615 N_A_871_74#_c_685_n N_SET_B_c_1229_n 0.00340414f $X=8.48 $Y=2.05 $X2=0
+ $Y2=0
cc_616 N_A_871_74#_c_706_n N_SET_B_c_1230_n 0.0024584f $X=7.995 $Y=2.99 $X2=0
+ $Y2=0
cc_617 N_A_871_74#_c_708_n N_SET_B_c_1230_n 0.0189577f $X=8.08 $Y=2.905 $X2=0
+ $Y2=0
cc_618 N_A_871_74#_c_710_n N_SET_B_c_1230_n 0.00260708f $X=8.165 $Y=2.135 $X2=0
+ $Y2=0
cc_619 N_A_871_74#_c_685_n N_SET_B_M1013_g 0.00120161f $X=8.48 $Y=2.05 $X2=0
+ $Y2=0
cc_620 N_A_871_74#_c_686_n N_SET_B_M1013_g 0.00634353f $X=8.565 $Y=1.43 $X2=0
+ $Y2=0
cc_621 N_A_871_74#_c_674_n N_SET_B_c_1222_n 0.00307898f $X=11.18 $Y=1.41 $X2=0
+ $Y2=0
cc_622 N_A_871_74#_c_675_n N_SET_B_c_1222_n 0.00454536f $X=10.835 $Y=1.41 $X2=0
+ $Y2=0
cc_623 N_A_871_74#_c_676_n N_SET_B_c_1222_n 0.0108908f $X=11.67 $Y=1.545 $X2=0
+ $Y2=0
cc_624 N_A_871_74#_c_677_n N_SET_B_c_1222_n 0.00129463f $X=11.76 $Y=2.11 $X2=0
+ $Y2=0
cc_625 N_A_871_74#_c_709_n N_SET_B_c_1222_n 0.00699781f $X=8.395 $Y=2.135 $X2=0
+ $Y2=0
cc_626 N_A_871_74#_c_710_n N_SET_B_c_1222_n 6.08327e-19 $X=8.165 $Y=2.135 $X2=0
+ $Y2=0
cc_627 N_A_871_74#_c_685_n N_SET_B_c_1222_n 0.0184668f $X=8.48 $Y=2.05 $X2=0
+ $Y2=0
cc_628 N_A_871_74#_c_687_n N_SET_B_c_1222_n 0.024823f $X=10.545 $Y=1.365 $X2=0
+ $Y2=0
cc_629 N_A_871_74#_c_690_n N_SET_B_c_1222_n 0.0532159f $X=10.38 $Y=1.365 $X2=0
+ $Y2=0
cc_630 N_A_871_74#_c_691_n N_SET_B_c_1222_n 0.00257296f $X=11.39 $Y=1.41 $X2=0
+ $Y2=0
cc_631 N_A_871_74#_c_710_n N_SET_B_c_1223_n 4.33107e-19 $X=8.165 $Y=2.135 $X2=0
+ $Y2=0
cc_632 N_A_871_74#_c_685_n N_SET_B_c_1223_n 4.56685e-19 $X=8.48 $Y=2.05 $X2=0
+ $Y2=0
cc_633 N_A_871_74#_c_709_n N_SET_B_c_1224_n 0.00418019f $X=8.395 $Y=2.135 $X2=0
+ $Y2=0
cc_634 N_A_871_74#_c_710_n N_SET_B_c_1224_n 0.0129383f $X=8.165 $Y=2.135 $X2=0
+ $Y2=0
cc_635 N_A_871_74#_c_685_n N_SET_B_c_1224_n 0.0235365f $X=8.48 $Y=2.05 $X2=0
+ $Y2=0
cc_636 N_A_871_74#_c_709_n N_SET_B_c_1228_n 0.00157943f $X=8.395 $Y=2.135 $X2=0
+ $Y2=0
cc_637 N_A_871_74#_c_710_n N_SET_B_c_1228_n 0.00245159f $X=8.165 $Y=2.135 $X2=0
+ $Y2=0
cc_638 N_A_871_74#_c_685_n N_SET_B_c_1228_n 0.00142596f $X=8.48 $Y=2.05 $X2=0
+ $Y2=0
cc_639 N_A_871_74#_c_678_n N_A_619_368#_M1033_g 0.00716152f $X=4.495 $Y=0.505
+ $X2=0 $Y2=0
cc_640 N_A_871_74#_c_680_n N_A_619_368#_M1033_g 0.00462516f $X=4.66 $Y=0.34
+ $X2=0 $Y2=0
cc_641 N_A_871_74#_c_699_n N_A_619_368#_c_1387_n 0.00143497f $X=4.72 $Y=2.99
+ $X2=0 $Y2=0
cc_642 N_A_871_74#_c_670_n N_A_619_368#_c_1370_n 0.00865427f $X=5.56 $Y=1.365
+ $X2=0 $Y2=0
cc_643 N_A_871_74#_c_681_n N_A_619_368#_c_1370_n 3.40049e-19 $X=5.395 $Y=1.455
+ $X2=0 $Y2=0
cc_644 N_A_871_74#_c_689_n N_A_619_368#_c_1370_n 7.18595e-19 $X=5.395 $Y=1.29
+ $X2=0 $Y2=0
cc_645 N_A_871_74#_c_692_n N_A_619_368#_c_1388_n 0.0073253f $X=5.43 $Y=2.15
+ $X2=0 $Y2=0
cc_646 N_A_871_74#_c_693_n N_A_619_368#_c_1388_n 0.0113006f $X=5.43 $Y=2.24
+ $X2=0 $Y2=0
cc_647 N_A_871_74#_c_696_n N_A_619_368#_c_1388_n 0.00865427f $X=5.395 $Y=1.96
+ $X2=0 $Y2=0
cc_648 N_A_871_74#_c_697_n N_A_619_368#_c_1388_n 0.00723988f $X=4.555 $Y=2.725
+ $X2=0 $Y2=0
cc_649 N_A_871_74#_c_698_n N_A_619_368#_c_1388_n 0.01157f $X=6.07 $Y=2.99 $X2=0
+ $Y2=0
cc_650 N_A_871_74#_c_670_n N_A_619_368#_c_1371_n 0.00655065f $X=5.56 $Y=1.365
+ $X2=0 $Y2=0
cc_651 N_A_871_74#_c_681_n N_A_619_368#_c_1371_n 8.57179e-19 $X=5.395 $Y=1.455
+ $X2=0 $Y2=0
cc_652 N_A_871_74#_c_684_n N_A_619_368#_c_1371_n 8.21735e-19 $X=6.185 $Y=1.135
+ $X2=0 $Y2=0
cc_653 N_A_871_74#_c_678_n N_A_619_368#_c_1372_n 0.00120198f $X=4.495 $Y=0.505
+ $X2=0 $Y2=0
cc_654 N_A_871_74#_c_679_n N_A_619_368#_c_1372_n 0.00410477f $X=5.39 $Y=0.34
+ $X2=0 $Y2=0
cc_655 N_A_871_74#_c_693_n N_A_619_368#_c_1389_n 0.00882199f $X=5.43 $Y=2.24
+ $X2=0 $Y2=0
cc_656 N_A_871_74#_c_698_n N_A_619_368#_c_1389_n 0.0147556f $X=6.07 $Y=2.99
+ $X2=0 $Y2=0
cc_657 N_A_871_74#_c_678_n N_A_619_368#_c_1373_n 0.00417367f $X=4.495 $Y=0.505
+ $X2=0 $Y2=0
cc_658 N_A_871_74#_c_679_n N_A_619_368#_c_1373_n 0.0163078f $X=5.39 $Y=0.34
+ $X2=0 $Y2=0
cc_659 N_A_871_74#_c_689_n N_A_619_368#_c_1373_n 0.013812f $X=5.395 $Y=1.29
+ $X2=0 $Y2=0
cc_660 N_A_871_74#_c_693_n N_A_619_368#_c_1391_n 0.00216849f $X=5.43 $Y=2.24
+ $X2=0 $Y2=0
cc_661 N_A_871_74#_c_703_n N_A_619_368#_c_1391_n 0.00286544f $X=6.155 $Y=2.905
+ $X2=0 $Y2=0
cc_662 N_A_871_74#_c_698_n N_A_619_368#_c_1392_n 0.0175868f $X=6.07 $Y=2.99
+ $X2=0 $Y2=0
cc_663 N_A_871_74#_c_693_n N_A_619_368#_c_1393_n 0.0125463f $X=5.43 $Y=2.24
+ $X2=0 $Y2=0
cc_664 N_A_871_74#_c_703_n N_A_619_368#_c_1393_n 0.00443587f $X=6.155 $Y=2.905
+ $X2=0 $Y2=0
cc_665 N_A_871_74#_c_712_n N_A_619_368#_c_1393_n 0.00115602f $X=6.187 $Y=2.25
+ $X2=0 $Y2=0
cc_666 N_A_871_74#_c_698_n N_A_619_368#_c_1394_n 0.00458792f $X=6.07 $Y=2.99
+ $X2=0 $Y2=0
cc_667 N_A_871_74#_c_706_n N_A_619_368#_c_1394_n 0.0149204f $X=7.995 $Y=2.99
+ $X2=0 $Y2=0
cc_668 N_A_871_74#_c_707_n N_A_619_368#_c_1394_n 0.00420304f $X=7.325 $Y=2.99
+ $X2=0 $Y2=0
cc_669 N_A_871_74#_c_708_n N_A_619_368#_c_1395_n 0.00312262f $X=8.08 $Y=2.905
+ $X2=0 $Y2=0
cc_670 N_A_871_74#_c_709_n N_A_619_368#_c_1395_n 0.00356641f $X=8.395 $Y=2.135
+ $X2=0 $Y2=0
cc_671 N_A_871_74#_c_675_n N_A_619_368#_c_1397_n 0.0147418f $X=10.835 $Y=1.41
+ $X2=0 $Y2=0
cc_672 N_A_871_74#_c_675_n N_A_619_368#_c_1398_n 0.00314037f $X=10.835 $Y=1.41
+ $X2=0 $Y2=0
cc_673 N_A_871_74#_c_677_n N_A_619_368#_c_1400_n 0.00594157f $X=11.76 $Y=2.11
+ $X2=0 $Y2=0
cc_674 N_A_871_74#_c_691_n N_A_619_368#_c_1400_n 0.0147418f $X=11.39 $Y=1.41
+ $X2=0 $Y2=0
cc_675 N_A_871_74#_c_695_n N_A_619_368#_c_1401_n 0.0180414f $X=11.76 $Y=2.2
+ $X2=0 $Y2=0
cc_676 N_A_871_74#_c_695_n N_A_619_368#_c_1402_n 0.00737233f $X=11.76 $Y=2.2
+ $X2=0 $Y2=0
cc_677 N_A_871_74#_c_676_n N_A_619_368#_c_1375_n 0.0238518f $X=11.67 $Y=1.545
+ $X2=0 $Y2=0
cc_678 N_A_871_74#_c_695_n N_A_619_368#_c_1375_n 0.0132562f $X=11.76 $Y=2.2
+ $X2=0 $Y2=0
cc_679 N_A_871_74#_c_678_n N_A_619_368#_c_1378_n 0.00155122f $X=4.495 $Y=0.505
+ $X2=0 $Y2=0
cc_680 N_A_871_74#_c_681_n N_A_619_368#_c_1379_n 3.40049e-19 $X=5.395 $Y=1.455
+ $X2=0 $Y2=0
cc_681 N_A_871_74#_c_682_n N_A_619_368#_c_1379_n 0.00865427f $X=5.395 $Y=1.455
+ $X2=0 $Y2=0
cc_682 N_A_871_74#_c_674_n N_A_619_368#_c_1409_n 0.0147418f $X=11.18 $Y=1.41
+ $X2=0 $Y2=0
cc_683 N_A_871_74#_c_676_n N_A_619_368#_c_1380_n 0.00719229f $X=11.67 $Y=1.545
+ $X2=0 $Y2=0
cc_684 N_A_871_74#_c_691_n N_A_619_368#_c_1380_n 0.00115082f $X=11.39 $Y=1.41
+ $X2=0 $Y2=0
cc_685 N_A_871_74#_M1015_d N_A_619_368#_c_1411_n 0.00379644f $X=4.37 $Y=1.84
+ $X2=0 $Y2=0
cc_686 N_A_871_74#_c_678_n N_A_619_368#_c_1383_n 0.0130668f $X=4.495 $Y=0.505
+ $X2=0 $Y2=0
cc_687 N_A_871_74#_c_675_n N_A_619_368#_c_1413_n 0.015083f $X=10.835 $Y=1.41
+ $X2=0 $Y2=0
cc_688 N_A_871_74#_c_677_n N_A_619_368#_c_1413_n 0.0122f $X=11.76 $Y=2.11 $X2=0
+ $Y2=0
cc_689 N_A_871_74#_c_687_n N_A_619_368#_c_1413_n 0.0651024f $X=10.545 $Y=1.365
+ $X2=0 $Y2=0
cc_690 N_A_871_74#_c_690_n N_A_619_368#_c_1413_n 0.0757222f $X=10.38 $Y=1.365
+ $X2=0 $Y2=0
cc_691 N_A_871_74#_c_676_n N_A_619_368#_c_1384_n 0.00963508f $X=11.67 $Y=1.545
+ $X2=0 $Y2=0
cc_692 N_A_871_74#_c_677_n N_A_619_368#_c_1384_n 0.00312843f $X=11.76 $Y=2.11
+ $X2=0 $Y2=0
cc_693 N_A_871_74#_c_688_n N_A_619_368#_c_1384_n 0.0163715f $X=11.225 $Y=1.365
+ $X2=0 $Y2=0
cc_694 N_A_871_74#_c_691_n N_A_619_368#_c_1384_n 0.0016069f $X=11.39 $Y=1.41
+ $X2=0 $Y2=0
cc_695 N_A_871_74#_c_685_n N_A_619_368#_c_1386_n 0.00575281f $X=8.48 $Y=2.05
+ $X2=0 $Y2=0
cc_696 N_A_871_74#_c_690_n N_A_619_368#_c_1386_n 0.00273126f $X=10.38 $Y=1.365
+ $X2=0 $Y2=0
cc_697 N_A_871_74#_c_685_n N_A_619_368#_c_1416_n 0.020865f $X=8.48 $Y=2.05 $X2=0
+ $Y2=0
cc_698 N_A_871_74#_c_690_n N_A_619_368#_c_1416_n 0.0204754f $X=10.38 $Y=1.365
+ $X2=0 $Y2=0
cc_699 N_A_871_74#_c_677_n N_A_2067_74#_c_1778_n 0.00412941f $X=11.76 $Y=2.11
+ $X2=0 $Y2=0
cc_700 N_A_871_74#_c_695_n N_A_2067_74#_c_1778_n 0.00690499f $X=11.76 $Y=2.2
+ $X2=0 $Y2=0
cc_701 N_A_871_74#_M1037_g N_A_2067_74#_c_1762_n 0.0108721f $X=10.76 $Y=0.69
+ $X2=0 $Y2=0
cc_702 N_A_871_74#_c_674_n N_A_2067_74#_c_1762_n 0.0127999f $X=11.18 $Y=1.41
+ $X2=0 $Y2=0
cc_703 N_A_871_74#_c_688_n N_A_2067_74#_c_1762_n 0.0484336f $X=11.225 $Y=1.365
+ $X2=0 $Y2=0
cc_704 N_A_871_74#_M1037_g N_A_2067_74#_c_1763_n 0.00325302f $X=10.76 $Y=0.69
+ $X2=0 $Y2=0
cc_705 N_A_871_74#_c_676_n N_A_2067_74#_c_1763_n 0.00296879f $X=11.67 $Y=1.545
+ $X2=0 $Y2=0
cc_706 N_A_871_74#_c_688_n N_A_2067_74#_c_1763_n 7.314e-19 $X=11.225 $Y=1.365
+ $X2=0 $Y2=0
cc_707 N_A_871_74#_c_691_n N_A_2067_74#_c_1763_n 2.19145e-19 $X=11.39 $Y=1.41
+ $X2=0 $Y2=0
cc_708 N_A_871_74#_c_695_n N_A_2067_74#_c_1779_n 0.00543714f $X=11.76 $Y=2.2
+ $X2=0 $Y2=0
cc_709 N_A_871_74#_M1032_g N_A_2067_74#_c_1766_n 0.00233014f $X=10.26 $Y=0.69
+ $X2=0 $Y2=0
cc_710 N_A_871_74#_M1037_g N_A_2067_74#_c_1766_n 0.00694931f $X=10.76 $Y=0.69
+ $X2=0 $Y2=0
cc_711 N_A_871_74#_c_675_n N_A_2067_74#_c_1766_n 0.00409869f $X=10.835 $Y=1.41
+ $X2=0 $Y2=0
cc_712 N_A_871_74#_c_687_n N_A_2067_74#_c_1766_n 0.0257498f $X=10.545 $Y=1.365
+ $X2=0 $Y2=0
cc_713 N_A_871_74#_c_677_n N_A_2067_74#_c_1784_n 0.00178103f $X=11.76 $Y=2.11
+ $X2=0 $Y2=0
cc_714 N_A_871_74#_c_695_n N_A_2067_74#_c_1784_n 0.0054952f $X=11.76 $Y=2.2
+ $X2=0 $Y2=0
cc_715 N_A_871_74#_c_676_n N_A_2067_74#_c_1767_n 4.20992e-19 $X=11.67 $Y=1.545
+ $X2=0 $Y2=0
cc_716 N_A_871_74#_c_677_n N_A_2067_74#_c_1767_n 0.00100497f $X=11.76 $Y=2.11
+ $X2=0 $Y2=0
cc_717 N_A_871_74#_c_704_n N_VPWR_M1034_d 0.0125482f $X=7.155 $Y=2.25 $X2=0
+ $Y2=0
cc_718 N_A_871_74#_c_705_n N_VPWR_M1034_d 0.0121457f $X=7.24 $Y=2.905 $X2=0
+ $Y2=0
cc_719 N_A_871_74#_c_708_n N_VPWR_M1029_d 0.00453281f $X=8.08 $Y=2.905 $X2=0
+ $Y2=0
cc_720 N_A_871_74#_c_698_n N_VPWR_c_2060_n 0.0156599f $X=6.07 $Y=2.99 $X2=0
+ $Y2=0
cc_721 N_A_871_74#_c_703_n N_VPWR_c_2060_n 0.0228376f $X=6.155 $Y=2.905 $X2=0
+ $Y2=0
cc_722 N_A_871_74#_c_704_n N_VPWR_c_2060_n 0.0419084f $X=7.155 $Y=2.25 $X2=0
+ $Y2=0
cc_723 N_A_871_74#_c_705_n N_VPWR_c_2060_n 0.0324324f $X=7.24 $Y=2.905 $X2=0
+ $Y2=0
cc_724 N_A_871_74#_c_707_n N_VPWR_c_2060_n 0.0156604f $X=7.325 $Y=2.99 $X2=0
+ $Y2=0
cc_725 N_A_871_74#_c_706_n N_VPWR_c_2061_n 0.0546768f $X=7.995 $Y=2.99 $X2=0
+ $Y2=0
cc_726 N_A_871_74#_c_707_n N_VPWR_c_2061_n 0.0115893f $X=7.325 $Y=2.99 $X2=0
+ $Y2=0
cc_727 N_A_871_74#_c_706_n N_VPWR_c_2062_n 0.0150384f $X=7.995 $Y=2.99 $X2=0
+ $Y2=0
cc_728 N_A_871_74#_c_708_n N_VPWR_c_2062_n 0.0398051f $X=8.08 $Y=2.905 $X2=0
+ $Y2=0
cc_729 N_A_871_74#_c_709_n N_VPWR_c_2062_n 0.0203752f $X=8.395 $Y=2.135 $X2=0
+ $Y2=0
cc_730 N_A_871_74#_c_698_n N_VPWR_c_2080_n 0.0975191f $X=6.07 $Y=2.99 $X2=0
+ $Y2=0
cc_731 N_A_871_74#_c_699_n N_VPWR_c_2080_n 0.0234498f $X=4.72 $Y=2.99 $X2=0
+ $Y2=0
cc_732 N_A_871_74#_c_699_n N_VPWR_c_2086_n 0.0128057f $X=4.72 $Y=2.99 $X2=0
+ $Y2=0
cc_733 N_A_871_74#_c_698_n N_VPWR_c_2057_n 0.0511446f $X=6.07 $Y=2.99 $X2=0
+ $Y2=0
cc_734 N_A_871_74#_c_699_n N_VPWR_c_2057_n 0.0127907f $X=4.72 $Y=2.99 $X2=0
+ $Y2=0
cc_735 N_A_871_74#_c_706_n N_VPWR_c_2057_n 0.028344f $X=7.995 $Y=2.99 $X2=0
+ $Y2=0
cc_736 N_A_871_74#_c_707_n N_VPWR_c_2057_n 0.00583135f $X=7.325 $Y=2.99 $X2=0
+ $Y2=0
cc_737 N_A_871_74#_c_679_n N_A_304_464#_M1019_s 0.00224741f $X=5.39 $Y=0.34
+ $X2=0 $Y2=0
cc_738 N_A_871_74#_M1015_d N_A_304_464#_c_2263_n 0.00585766f $X=4.37 $Y=1.84
+ $X2=0 $Y2=0
cc_739 N_A_871_74#_c_697_n N_A_304_464#_c_2263_n 0.0235896f $X=4.555 $Y=2.725
+ $X2=0 $Y2=0
cc_740 N_A_871_74#_c_698_n N_A_304_464#_c_2263_n 0.00442331f $X=6.07 $Y=2.99
+ $X2=0 $Y2=0
cc_741 N_A_871_74#_c_678_n N_A_304_464#_c_2258_n 0.0273357f $X=4.495 $Y=0.505
+ $X2=0 $Y2=0
cc_742 N_A_871_74#_c_679_n N_A_304_464#_c_2258_n 0.0199805f $X=5.39 $Y=0.34
+ $X2=0 $Y2=0
cc_743 N_A_871_74#_c_689_n N_A_304_464#_c_2258_n 0.0100954f $X=5.395 $Y=1.29
+ $X2=0 $Y2=0
cc_744 N_A_871_74#_c_692_n N_A_304_464#_c_2265_n 0.00101758f $X=5.43 $Y=2.15
+ $X2=0 $Y2=0
cc_745 N_A_871_74#_c_693_n N_A_304_464#_c_2265_n 0.00992949f $X=5.43 $Y=2.24
+ $X2=0 $Y2=0
cc_746 N_A_871_74#_c_696_n N_A_304_464#_c_2265_n 8.40494e-19 $X=5.395 $Y=1.96
+ $X2=0 $Y2=0
cc_747 N_A_871_74#_c_697_n N_A_304_464#_c_2265_n 0.0215555f $X=4.555 $Y=2.725
+ $X2=0 $Y2=0
cc_748 N_A_871_74#_c_698_n N_A_304_464#_c_2265_n 0.0345124f $X=6.07 $Y=2.99
+ $X2=0 $Y2=0
cc_749 N_A_871_74#_c_681_n N_A_304_464#_c_2265_n 0.012049f $X=5.395 $Y=1.455
+ $X2=0 $Y2=0
cc_750 N_A_871_74#_c_692_n N_A_304_464#_c_2259_n 0.00117754f $X=5.43 $Y=2.15
+ $X2=0 $Y2=0
cc_751 N_A_871_74#_c_670_n N_A_304_464#_c_2259_n 0.00447757f $X=5.56 $Y=1.365
+ $X2=0 $Y2=0
cc_752 N_A_871_74#_c_681_n N_A_304_464#_c_2259_n 0.0502424f $X=5.395 $Y=1.455
+ $X2=0 $Y2=0
cc_753 N_A_871_74#_c_689_n N_A_304_464#_c_2259_n 0.0181764f $X=5.395 $Y=1.29
+ $X2=0 $Y2=0
cc_754 N_A_871_74#_c_703_n A_1201_463# 0.00497225f $X=6.155 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_755 N_A_871_74#_c_709_n N_A_1789_424#_c_2377_n 0.00491328f $X=8.395 $Y=2.135
+ $X2=0 $Y2=0
cc_756 N_A_871_74#_c_695_n N_A_2277_455#_c_2427_n 0.00418069f $X=11.76 $Y=2.2
+ $X2=0 $Y2=0
cc_757 N_A_871_74#_c_695_n N_A_2277_455#_c_2428_n 0.00213109f $X=11.76 $Y=2.2
+ $X2=0 $Y2=0
cc_758 N_A_871_74#_c_680_n N_VGND_c_2519_n 0.011924f $X=4.66 $Y=0.34 $X2=0 $Y2=0
cc_759 N_A_871_74#_M1032_g N_VGND_c_2522_n 3.12362e-19 $X=10.26 $Y=0.69 $X2=0
+ $Y2=0
cc_760 N_A_871_74#_M1032_g N_VGND_c_2533_n 0.00278247f $X=10.26 $Y=0.69 $X2=0
+ $Y2=0
cc_761 N_A_871_74#_M1037_g N_VGND_c_2533_n 0.00278271f $X=10.76 $Y=0.69 $X2=0
+ $Y2=0
cc_762 N_A_871_74#_M1027_g N_VGND_c_2541_n 0.00405757f $X=6.295 $Y=0.615 $X2=0
+ $Y2=0
cc_763 N_A_871_74#_c_679_n N_VGND_c_2541_n 0.0591538f $X=5.39 $Y=0.34 $X2=0
+ $Y2=0
cc_764 N_A_871_74#_c_680_n N_VGND_c_2541_n 0.0235688f $X=4.66 $Y=0.34 $X2=0
+ $Y2=0
cc_765 N_A_871_74#_M1027_g N_VGND_c_2550_n 0.00534666f $X=6.295 $Y=0.615 $X2=0
+ $Y2=0
cc_766 N_A_871_74#_M1032_g N_VGND_c_2550_n 0.00354182f $X=10.26 $Y=0.69 $X2=0
+ $Y2=0
cc_767 N_A_871_74#_M1037_g N_VGND_c_2550_n 0.00358176f $X=10.76 $Y=0.69 $X2=0
+ $Y2=0
cc_768 N_A_871_74#_c_679_n N_VGND_c_2550_n 0.0340476f $X=5.39 $Y=0.34 $X2=0
+ $Y2=0
cc_769 N_A_871_74#_c_680_n N_VGND_c_2550_n 0.0127152f $X=4.66 $Y=0.34 $X2=0
+ $Y2=0
cc_770 N_A_871_74#_M1032_g N_A_1794_74#_c_2705_n 0.00556597f $X=10.26 $Y=0.69
+ $X2=0 $Y2=0
cc_771 N_A_871_74#_M1037_g N_A_1794_74#_c_2705_n 6.97072e-19 $X=10.76 $Y=0.69
+ $X2=0 $Y2=0
cc_772 N_A_871_74#_c_690_n N_A_1794_74#_c_2705_n 0.0650467f $X=10.38 $Y=1.365
+ $X2=0 $Y2=0
cc_773 N_A_871_74#_c_690_n N_A_1794_74#_c_2706_n 0.0189433f $X=10.38 $Y=1.365
+ $X2=0 $Y2=0
cc_774 N_A_871_74#_M1032_g N_A_1794_74#_c_2714_n 0.007555f $X=10.26 $Y=0.69
+ $X2=0 $Y2=0
cc_775 N_A_871_74#_M1037_g N_A_1794_74#_c_2714_n 6.40354e-19 $X=10.76 $Y=0.69
+ $X2=0 $Y2=0
cc_776 N_A_871_74#_M1032_g N_A_1794_74#_c_2707_n 0.0104037f $X=10.26 $Y=0.69
+ $X2=0 $Y2=0
cc_777 N_A_871_74#_M1037_g N_A_1794_74#_c_2707_n 0.0112187f $X=10.76 $Y=0.69
+ $X2=0 $Y2=0
cc_778 N_A_871_74#_M1032_g N_A_1794_74#_c_2708_n 0.00155275f $X=10.26 $Y=0.69
+ $X2=0 $Y2=0
cc_779 N_A_871_74#_M1037_g N_A_1794_74#_c_2709_n 0.00165289f $X=10.76 $Y=0.69
+ $X2=0 $Y2=0
cc_780 N_A_1252_376#_c_950_n N_A_1069_81#_c_1032_n 0.019879f $X=7.495 $Y=1.865
+ $X2=0 $Y2=0
cc_781 N_A_1252_376#_c_951_n N_A_1069_81#_c_1032_n 0.00815395f $X=6.8 $Y=1.865
+ $X2=0 $Y2=0
cc_782 N_A_1252_376#_c_953_n N_A_1069_81#_c_1032_n 0.00694514f $X=7.66 $Y=2.295
+ $X2=0 $Y2=0
cc_783 N_A_1252_376#_c_952_n N_A_1069_81#_c_1053_n 0.00515236f $X=7.66 $Y=2.515
+ $X2=0 $Y2=0
cc_784 N_A_1252_376#_c_953_n N_A_1069_81#_c_1053_n 0.00371781f $X=7.66 $Y=2.295
+ $X2=0 $Y2=0
cc_785 N_A_1252_376#_c_942_n N_A_1069_81#_M1012_g 0.0056748f $X=7.38 $Y=0.955
+ $X2=0 $Y2=0
cc_786 N_A_1252_376#_c_943_n N_A_1069_81#_M1012_g 0.0116694f $X=7.545 $Y=0.58
+ $X2=0 $Y2=0
cc_787 N_A_1252_376#_c_944_n N_A_1069_81#_M1012_g 8.40065e-19 $X=6.98 $Y=0.955
+ $X2=0 $Y2=0
cc_788 N_A_1252_376#_c_946_n N_A_1069_81#_M1012_g 0.00473478f $X=6.89 $Y=1.1
+ $X2=0 $Y2=0
cc_789 N_A_1252_376#_c_941_n N_A_1069_81#_c_1074_n 0.0113068f $X=6.685 $Y=0.935
+ $X2=0 $Y2=0
cc_790 N_A_1252_376#_c_941_n N_A_1069_81#_c_1042_n 0.00436872f $X=6.685 $Y=0.935
+ $X2=0 $Y2=0
cc_791 N_A_1252_376#_c_944_n N_A_1069_81#_c_1042_n 0.0261072f $X=6.98 $Y=0.955
+ $X2=0 $Y2=0
cc_792 N_A_1252_376#_c_946_n N_A_1069_81#_c_1042_n 0.00911922f $X=6.89 $Y=1.1
+ $X2=0 $Y2=0
cc_793 N_A_1252_376#_c_950_n N_A_1069_81#_c_1043_n 0.0532877f $X=7.495 $Y=1.865
+ $X2=0 $Y2=0
cc_794 N_A_1252_376#_c_951_n N_A_1069_81#_c_1043_n 0.00180482f $X=6.8 $Y=1.865
+ $X2=0 $Y2=0
cc_795 N_A_1252_376#_c_942_n N_A_1069_81#_c_1043_n 0.00950459f $X=7.38 $Y=0.955
+ $X2=0 $Y2=0
cc_796 N_A_1252_376#_c_944_n N_A_1069_81#_c_1043_n 0.0243532f $X=6.98 $Y=0.955
+ $X2=0 $Y2=0
cc_797 N_A_1252_376#_c_945_n N_A_1069_81#_c_1043_n 0.0113822f $X=6.8 $Y=1.7
+ $X2=0 $Y2=0
cc_798 N_A_1252_376#_c_946_n N_A_1069_81#_c_1043_n 0.00787396f $X=6.89 $Y=1.1
+ $X2=0 $Y2=0
cc_799 N_A_1252_376#_c_948_n N_A_1069_81#_c_1044_n 0.00342884f $X=6.635 $Y=1.955
+ $X2=0 $Y2=0
cc_800 N_A_1252_376#_c_950_n N_A_1069_81#_c_1044_n 8.29766e-19 $X=7.495 $Y=1.865
+ $X2=0 $Y2=0
cc_801 N_A_1252_376#_c_942_n N_A_1069_81#_c_1045_n 0.00352223f $X=7.38 $Y=0.955
+ $X2=0 $Y2=0
cc_802 N_A_1252_376#_c_942_n N_A_1069_81#_c_1046_n 0.011024f $X=7.38 $Y=0.955
+ $X2=0 $Y2=0
cc_803 N_A_1252_376#_c_949_n N_A_1069_81#_c_1049_n 0.00127968f $X=6.35 $Y=1.955
+ $X2=0 $Y2=0
cc_804 N_A_1252_376#_c_950_n N_A_1069_81#_c_1050_n 0.0251552f $X=7.495 $Y=1.865
+ $X2=0 $Y2=0
cc_805 N_A_1252_376#_c_942_n N_A_1069_81#_c_1050_n 0.0260001f $X=7.38 $Y=0.955
+ $X2=0 $Y2=0
cc_806 N_A_1252_376#_c_944_n N_A_1069_81#_c_1050_n 9.46074e-19 $X=6.98 $Y=0.955
+ $X2=0 $Y2=0
cc_807 N_A_1252_376#_c_945_n N_A_1069_81#_c_1050_n 8.62215e-19 $X=6.8 $Y=1.7
+ $X2=0 $Y2=0
cc_808 N_A_1252_376#_c_946_n N_A_1069_81#_c_1050_n 3.37949e-19 $X=6.89 $Y=1.1
+ $X2=0 $Y2=0
cc_809 N_A_1252_376#_c_950_n N_A_1069_81#_c_1051_n 0.00102424f $X=7.495 $Y=1.865
+ $X2=0 $Y2=0
cc_810 N_A_1252_376#_c_942_n N_A_1069_81#_c_1051_n 0.0090276f $X=7.38 $Y=0.955
+ $X2=0 $Y2=0
cc_811 N_A_1252_376#_c_944_n N_A_1069_81#_c_1051_n 4.25533e-19 $X=6.98 $Y=0.955
+ $X2=0 $Y2=0
cc_812 N_A_1252_376#_c_945_n N_A_1069_81#_c_1051_n 0.0170764f $X=6.8 $Y=1.7
+ $X2=0 $Y2=0
cc_813 N_A_1252_376#_c_946_n N_A_1069_81#_c_1051_n 0.0072023f $X=6.89 $Y=1.1
+ $X2=0 $Y2=0
cc_814 N_A_1252_376#_c_953_n N_SET_B_c_1229_n 0.00251983f $X=7.66 $Y=2.295 $X2=0
+ $Y2=0
cc_815 N_A_1252_376#_c_952_n N_SET_B_c_1230_n 0.00370559f $X=7.66 $Y=2.515 $X2=0
+ $Y2=0
cc_816 N_A_1252_376#_c_953_n N_SET_B_c_1230_n 4.00437e-19 $X=7.66 $Y=2.295 $X2=0
+ $Y2=0
cc_817 N_A_1252_376#_c_943_n N_SET_B_M1013_g 0.00187295f $X=7.545 $Y=0.58 $X2=0
+ $Y2=0
cc_818 N_A_1252_376#_c_950_n N_SET_B_c_1223_n 0.00142282f $X=7.495 $Y=1.865
+ $X2=0 $Y2=0
cc_819 N_A_1252_376#_c_952_n N_SET_B_c_1223_n 0.00185005f $X=7.66 $Y=2.515 $X2=0
+ $Y2=0
cc_820 N_A_1252_376#_c_950_n N_SET_B_c_1224_n 0.0122254f $X=7.495 $Y=1.865 $X2=0
+ $Y2=0
cc_821 N_A_1252_376#_c_950_n N_SET_B_c_1228_n 0.00361742f $X=7.495 $Y=1.865
+ $X2=0 $Y2=0
cc_822 N_A_1252_376#_c_947_n N_A_619_368#_c_1391_n 0.00222169f $X=6.35 $Y=2.24
+ $X2=0 $Y2=0
cc_823 N_A_1252_376#_c_947_n N_A_619_368#_c_1393_n 0.0214261f $X=6.35 $Y=2.24
+ $X2=0 $Y2=0
cc_824 N_A_1252_376#_c_949_n N_A_619_368#_c_1393_n 0.00249329f $X=6.35 $Y=1.955
+ $X2=0 $Y2=0
cc_825 N_A_1252_376#_c_947_n N_A_619_368#_c_1394_n 0.0103562f $X=6.35 $Y=2.24
+ $X2=0 $Y2=0
cc_826 N_A_1252_376#_c_947_n N_VPWR_c_2060_n 0.0120251f $X=6.35 $Y=2.24 $X2=0
+ $Y2=0
cc_827 N_A_1252_376#_c_947_n N_VPWR_c_2057_n 8.51577e-19 $X=6.35 $Y=2.24 $X2=0
+ $Y2=0
cc_828 N_A_1252_376#_c_941_n N_VGND_c_2520_n 0.00545418f $X=6.685 $Y=0.935 $X2=0
+ $Y2=0
cc_829 N_A_1252_376#_c_943_n N_VGND_c_2520_n 0.0236236f $X=7.545 $Y=0.58 $X2=0
+ $Y2=0
cc_830 N_A_1252_376#_c_944_n N_VGND_c_2520_n 0.0287015f $X=6.98 $Y=0.955 $X2=0
+ $Y2=0
cc_831 N_A_1252_376#_c_946_n N_VGND_c_2520_n 0.00217452f $X=6.89 $Y=1.1 $X2=0
+ $Y2=0
cc_832 N_A_1252_376#_c_943_n N_VGND_c_2521_n 0.0104546f $X=7.545 $Y=0.58 $X2=0
+ $Y2=0
cc_833 N_A_1252_376#_c_941_n N_VGND_c_2541_n 0.00518115f $X=6.685 $Y=0.935 $X2=0
+ $Y2=0
cc_834 N_A_1252_376#_c_943_n N_VGND_c_2542_n 0.0145794f $X=7.545 $Y=0.58 $X2=0
+ $Y2=0
cc_835 N_A_1252_376#_c_941_n N_VGND_c_2550_n 0.00534666f $X=6.685 $Y=0.935 $X2=0
+ $Y2=0
cc_836 N_A_1252_376#_c_943_n N_VGND_c_2550_n 0.0120044f $X=7.545 $Y=0.58 $X2=0
+ $Y2=0
cc_837 N_A_1069_81#_c_1032_n N_SET_B_c_1229_n 0.00668782f $X=7.435 $Y=2.15 $X2=0
+ $Y2=0
cc_838 N_A_1069_81#_c_1053_n N_SET_B_c_1230_n 0.0167374f $X=7.435 $Y=2.24 $X2=0
+ $Y2=0
cc_839 N_A_1069_81#_M1012_g N_SET_B_M1013_g 0.0537337f $X=7.76 $Y=0.58 $X2=0
+ $Y2=0
cc_840 N_A_1069_81#_c_1046_n N_SET_B_M1013_g 0.00531188f $X=8.05 $Y=1.037 $X2=0
+ $Y2=0
cc_841 N_A_1069_81#_c_1047_n N_SET_B_M1013_g 0.0172588f $X=8.695 $Y=1.065 $X2=0
+ $Y2=0
cc_842 N_A_1069_81#_c_1048_n N_SET_B_M1013_g 0.0140045f $X=8.695 $Y=1.065 $X2=0
+ $Y2=0
cc_843 N_A_1069_81#_c_1050_n N_SET_B_M1013_g 0.00108273f $X=7.51 $Y=1.295 $X2=0
+ $Y2=0
cc_844 N_A_1069_81#_c_1051_n N_SET_B_M1013_g 0.00736022f $X=7.52 $Y=1.375 $X2=0
+ $Y2=0
cc_845 N_A_1069_81#_c_1035_n N_SET_B_c_1222_n 0.00307941f $X=9.365 $Y=1.955
+ $X2=0 $Y2=0
cc_846 N_A_1069_81#_c_1037_n N_SET_B_c_1222_n 0.0037079f $X=9.815 $Y=1.955 $X2=0
+ $Y2=0
cc_847 N_A_1069_81#_c_1047_n N_SET_B_c_1222_n 0.00863597f $X=8.695 $Y=1.065
+ $X2=0 $Y2=0
cc_848 N_A_1069_81#_c_1045_n N_SET_B_c_1223_n 0.00409741f $X=7.88 $Y=1.295 $X2=0
+ $Y2=0
cc_849 N_A_1069_81#_c_1046_n N_SET_B_c_1223_n 0.00414232f $X=8.05 $Y=1.037 $X2=0
+ $Y2=0
cc_850 N_A_1069_81#_c_1047_n N_SET_B_c_1223_n 3.14556e-19 $X=8.695 $Y=1.065
+ $X2=0 $Y2=0
cc_851 N_A_1069_81#_c_1050_n N_SET_B_c_1223_n 4.88841e-19 $X=7.51 $Y=1.295 $X2=0
+ $Y2=0
cc_852 N_A_1069_81#_c_1051_n N_SET_B_c_1223_n 0.00312846f $X=7.52 $Y=1.375 $X2=0
+ $Y2=0
cc_853 N_A_1069_81#_c_1032_n N_SET_B_c_1224_n 3.68151e-19 $X=7.435 $Y=2.15 $X2=0
+ $Y2=0
cc_854 N_A_1069_81#_c_1045_n N_SET_B_c_1224_n 0.0029943f $X=7.88 $Y=1.295 $X2=0
+ $Y2=0
cc_855 N_A_1069_81#_c_1046_n N_SET_B_c_1224_n 0.0116033f $X=8.05 $Y=1.037 $X2=0
+ $Y2=0
cc_856 N_A_1069_81#_c_1047_n N_SET_B_c_1224_n 0.00565821f $X=8.695 $Y=1.065
+ $X2=0 $Y2=0
cc_857 N_A_1069_81#_c_1050_n N_SET_B_c_1224_n 9.69441e-19 $X=7.51 $Y=1.295 $X2=0
+ $Y2=0
cc_858 N_A_1069_81#_c_1051_n N_SET_B_c_1224_n 0.00262295f $X=7.52 $Y=1.375 $X2=0
+ $Y2=0
cc_859 N_A_1069_81#_c_1046_n N_SET_B_c_1228_n 0.0029438f $X=8.05 $Y=1.037 $X2=0
+ $Y2=0
cc_860 N_A_1069_81#_c_1047_n N_SET_B_c_1228_n 4.48072e-19 $X=8.695 $Y=1.065
+ $X2=0 $Y2=0
cc_861 N_A_1069_81#_c_1051_n N_SET_B_c_1228_n 0.00668782f $X=7.52 $Y=1.375 $X2=0
+ $Y2=0
cc_862 N_A_1069_81#_c_1058_n N_A_619_368#_c_1393_n 0.00627699f $X=5.705 $Y=2.515
+ $X2=0 $Y2=0
cc_863 N_A_1069_81#_c_1049_n N_A_619_368#_c_1393_n 0.00324592f $X=5.72 $Y=2.295
+ $X2=0 $Y2=0
cc_864 N_A_1069_81#_c_1053_n N_A_619_368#_c_1394_n 0.00882199f $X=7.435 $Y=2.24
+ $X2=0 $Y2=0
cc_865 N_A_1069_81#_c_1055_n N_A_619_368#_c_1395_n 0.0256685f $X=9.365 $Y=2.045
+ $X2=0 $Y2=0
cc_866 N_A_1069_81#_c_1057_n N_A_619_368#_c_1396_n 0.014266f $X=9.815 $Y=2.045
+ $X2=0 $Y2=0
cc_867 N_A_1069_81#_c_1037_n N_A_619_368#_c_1398_n 0.0089869f $X=9.815 $Y=1.955
+ $X2=0 $Y2=0
cc_868 N_A_1069_81#_c_1035_n N_A_619_368#_c_1413_n 0.0107247f $X=9.365 $Y=1.955
+ $X2=0 $Y2=0
cc_869 N_A_1069_81#_c_1036_n N_A_619_368#_c_1413_n 4.15884e-19 $X=9.725 $Y=1.31
+ $X2=0 $Y2=0
cc_870 N_A_1069_81#_c_1037_n N_A_619_368#_c_1413_n 0.0132533f $X=9.815 $Y=1.955
+ $X2=0 $Y2=0
cc_871 N_A_1069_81#_c_1035_n N_A_619_368#_c_1386_n 0.0212879f $X=9.365 $Y=1.955
+ $X2=0 $Y2=0
cc_872 N_A_1069_81#_c_1048_n N_A_619_368#_c_1386_n 0.010169f $X=8.695 $Y=1.065
+ $X2=0 $Y2=0
cc_873 N_A_1069_81#_c_1035_n N_A_619_368#_c_1416_n 7.54793e-19 $X=9.365 $Y=1.955
+ $X2=0 $Y2=0
cc_874 N_A_1069_81#_c_1057_n N_A_2067_74#_c_1804_n 2.21057e-19 $X=9.815 $Y=2.045
+ $X2=0 $Y2=0
cc_875 N_A_1069_81#_c_1057_n N_A_2067_74#_c_1805_n 3.19228e-19 $X=9.815 $Y=2.045
+ $X2=0 $Y2=0
cc_876 N_A_1069_81#_c_1055_n N_VPWR_c_2063_n 0.00975701f $X=9.365 $Y=2.045 $X2=0
+ $Y2=0
cc_877 N_A_1069_81#_c_1057_n N_VPWR_c_2063_n 0.00338591f $X=9.815 $Y=2.045 $X2=0
+ $Y2=0
cc_878 N_A_1069_81#_c_1055_n N_VPWR_c_2070_n 0.00413917f $X=9.365 $Y=2.045 $X2=0
+ $Y2=0
cc_879 N_A_1069_81#_c_1057_n N_VPWR_c_2072_n 0.0044313f $X=9.815 $Y=2.045 $X2=0
+ $Y2=0
cc_880 N_A_1069_81#_c_1055_n N_VPWR_c_2057_n 0.00818781f $X=9.365 $Y=2.045 $X2=0
+ $Y2=0
cc_881 N_A_1069_81#_c_1057_n N_VPWR_c_2057_n 0.00853445f $X=9.815 $Y=2.045 $X2=0
+ $Y2=0
cc_882 N_A_1069_81#_c_1058_n N_A_304_464#_c_2265_n 0.0182846f $X=5.705 $Y=2.515
+ $X2=0 $Y2=0
cc_883 N_A_1069_81#_c_1049_n N_A_304_464#_c_2265_n 0.0072134f $X=5.72 $Y=2.295
+ $X2=0 $Y2=0
cc_884 N_A_1069_81#_c_1049_n N_A_304_464#_c_2259_n 0.00342338f $X=5.72 $Y=2.295
+ $X2=0 $Y2=0
cc_885 N_A_1069_81#_c_1055_n N_A_1789_424#_c_2379_n 0.0155754f $X=9.365 $Y=2.045
+ $X2=0 $Y2=0
cc_886 N_A_1069_81#_c_1057_n N_A_1789_424#_c_2379_n 0.0124366f $X=9.815 $Y=2.045
+ $X2=0 $Y2=0
cc_887 N_A_1069_81#_c_1057_n N_A_1789_424#_c_2373_n 0.00167065f $X=9.815
+ $Y=2.045 $X2=0 $Y2=0
cc_888 N_A_1069_81#_c_1055_n N_A_1789_424#_c_2382_n 6.71314e-19 $X=9.365
+ $Y=2.045 $X2=0 $Y2=0
cc_889 N_A_1069_81#_c_1057_n N_A_1789_424#_c_2382_n 0.00906265f $X=9.815
+ $Y=2.045 $X2=0 $Y2=0
cc_890 N_A_1069_81#_c_1057_n N_A_1789_424#_c_2375_n 0.0032261f $X=9.815 $Y=2.045
+ $X2=0 $Y2=0
cc_891 N_A_1069_81#_c_1055_n N_A_1789_424#_c_2377_n 0.00427855f $X=9.365
+ $Y=2.045 $X2=0 $Y2=0
cc_892 N_A_1069_81#_M1012_g N_VGND_c_2520_n 0.00342558f $X=7.76 $Y=0.58 $X2=0
+ $Y2=0
cc_893 N_A_1069_81#_M1012_g N_VGND_c_2521_n 0.00149517f $X=7.76 $Y=0.58 $X2=0
+ $Y2=0
cc_894 N_A_1069_81#_c_1047_n N_VGND_c_2521_n 0.0209685f $X=8.695 $Y=1.065 $X2=0
+ $Y2=0
cc_895 N_A_1069_81#_M1009_g N_VGND_c_2522_n 0.00973428f $X=9.83 $Y=0.69 $X2=0
+ $Y2=0
cc_896 N_A_1069_81#_c_1040_n N_VGND_c_2522_n 0.0115887f $X=9.365 $Y=1.085 $X2=0
+ $Y2=0
cc_897 N_A_1069_81#_c_1040_n N_VGND_c_2531_n 0.00444681f $X=9.365 $Y=1.085 $X2=0
+ $Y2=0
cc_898 N_A_1069_81#_M1009_g N_VGND_c_2533_n 0.00383152f $X=9.83 $Y=0.69 $X2=0
+ $Y2=0
cc_899 N_A_1069_81#_c_1074_n N_VGND_c_2541_n 0.0182889f $X=6.475 $Y=0.635 $X2=0
+ $Y2=0
cc_900 N_A_1069_81#_c_1078_n N_VGND_c_2541_n 0.00491805f $X=5.9 $Y=0.635 $X2=0
+ $Y2=0
cc_901 N_A_1069_81#_M1012_g N_VGND_c_2542_n 0.00434272f $X=7.76 $Y=0.58 $X2=0
+ $Y2=0
cc_902 N_A_1069_81#_M1012_g N_VGND_c_2550_n 0.00825979f $X=7.76 $Y=0.58 $X2=0
+ $Y2=0
cc_903 N_A_1069_81#_M1009_g N_VGND_c_2550_n 0.00757637f $X=9.83 $Y=0.69 $X2=0
+ $Y2=0
cc_904 N_A_1069_81#_c_1040_n N_VGND_c_2550_n 0.00882517f $X=9.365 $Y=1.085 $X2=0
+ $Y2=0
cc_905 N_A_1069_81#_c_1074_n N_VGND_c_2550_n 0.0246945f $X=6.475 $Y=0.635 $X2=0
+ $Y2=0
cc_906 N_A_1069_81#_c_1078_n N_VGND_c_2550_n 0.00580745f $X=5.9 $Y=0.635 $X2=0
+ $Y2=0
cc_907 N_A_1069_81#_c_1074_n A_1274_81# 0.00374924f $X=6.475 $Y=0.635 $X2=-0.19
+ $Y2=-0.245
cc_908 N_A_1069_81#_c_1042_n A_1274_81# 3.0566e-19 $X=6.56 $Y=1.395 $X2=-0.19
+ $Y2=-0.245
cc_909 N_A_1069_81#_c_1040_n N_A_1794_74#_c_2704_n 4.57511e-19 $X=9.365 $Y=1.085
+ $X2=0 $Y2=0
cc_910 N_A_1069_81#_c_1047_n N_A_1794_74#_c_2704_n 0.00836125f $X=8.695 $Y=1.065
+ $X2=0 $Y2=0
cc_911 N_A_1069_81#_c_1048_n N_A_1794_74#_c_2704_n 3.95109e-19 $X=8.695 $Y=1.065
+ $X2=0 $Y2=0
cc_912 N_A_1069_81#_c_1036_n N_A_1794_74#_c_2705_n 0.00286179f $X=9.725 $Y=1.31
+ $X2=0 $Y2=0
cc_913 N_A_1069_81#_M1009_g N_A_1794_74#_c_2705_n 0.0142903f $X=9.83 $Y=0.69
+ $X2=0 $Y2=0
cc_914 N_A_1069_81#_c_1039_n N_A_1794_74#_c_2705_n 0.00494339f $X=9.365 $Y=1.16
+ $X2=0 $Y2=0
cc_915 N_A_1069_81#_c_1040_n N_A_1794_74#_c_2705_n 0.00947016f $X=9.365 $Y=1.085
+ $X2=0 $Y2=0
cc_916 N_A_1069_81#_c_1034_n N_A_1794_74#_c_2706_n 0.00940114f $X=9.275 $Y=1.16
+ $X2=0 $Y2=0
cc_917 N_A_1069_81#_c_1047_n N_A_1794_74#_c_2706_n 0.0146575f $X=8.695 $Y=1.065
+ $X2=0 $Y2=0
cc_918 N_A_1069_81#_c_1048_n N_A_1794_74#_c_2706_n 3.57917e-19 $X=8.695 $Y=1.065
+ $X2=0 $Y2=0
cc_919 N_A_1069_81#_M1009_g N_A_1794_74#_c_2708_n 9.48753e-19 $X=9.83 $Y=0.69
+ $X2=0 $Y2=0
cc_920 N_SET_B_c_1230_n N_A_619_368#_c_1394_n 0.00922046f $X=7.985 $Y=2.24 $X2=0
+ $Y2=0
cc_921 N_SET_B_c_1230_n N_A_619_368#_c_1395_n 0.0084654f $X=7.985 $Y=2.24 $X2=0
+ $Y2=0
cc_922 N_SET_B_c_1222_n N_A_619_368#_c_1374_n 0.00259421f $X=13.055 $Y=1.665
+ $X2=0 $Y2=0
cc_923 N_SET_B_c_1222_n N_A_619_368#_c_1375_n 0.00188206f $X=13.055 $Y=1.665
+ $X2=0 $Y2=0
cc_924 N_SET_B_c_1222_n N_A_619_368#_c_1380_n 0.00334987f $X=13.055 $Y=1.665
+ $X2=0 $Y2=0
cc_925 N_SET_B_c_1222_n N_A_619_368#_c_1413_n 0.0734209f $X=13.055 $Y=1.665
+ $X2=0 $Y2=0
cc_926 N_SET_B_c_1222_n N_A_619_368#_c_1384_n 0.0166357f $X=13.055 $Y=1.665
+ $X2=0 $Y2=0
cc_927 N_SET_B_c_1229_n N_A_619_368#_c_1386_n 0.00194318f $X=7.985 $Y=2.15 $X2=0
+ $Y2=0
cc_928 N_SET_B_c_1222_n N_A_619_368#_c_1386_n 0.00260077f $X=13.055 $Y=1.665
+ $X2=0 $Y2=0
cc_929 N_SET_B_c_1228_n N_A_619_368#_c_1386_n 0.00509006f $X=8.06 $Y=1.715 $X2=0
+ $Y2=0
cc_930 N_SET_B_c_1222_n N_A_619_368#_c_1416_n 0.0149981f $X=13.055 $Y=1.665
+ $X2=0 $Y2=0
cc_931 N_SET_B_c_1231_n N_A_2513_258#_c_1654_n 0.012361f $X=13.25 $Y=2.375 $X2=0
+ $Y2=0
cc_932 N_SET_B_c_1234_n N_A_2513_258#_c_1654_n 5.67665e-19 $X=13.27 $Y=1.97
+ $X2=0 $Y2=0
cc_933 N_SET_B_c_1227_n N_A_2513_258#_c_1654_n 2.00699e-19 $X=13.27 $Y=1.465
+ $X2=0 $Y2=0
cc_934 N_SET_B_c_1232_n N_A_2513_258#_c_1655_n 0.0204406f $X=13.25 $Y=2.465
+ $X2=0 $Y2=0
cc_935 N_SET_B_M1021_g N_A_2513_258#_M1020_g 0.057484f $X=13.21 $Y=0.58 $X2=0
+ $Y2=0
cc_936 N_SET_B_c_1221_n N_A_2513_258#_c_1646_n 0.0139984f $X=13.27 $Y=1.805
+ $X2=0 $Y2=0
cc_937 N_SET_B_c_1222_n N_A_2513_258#_c_1646_n 0.0013891f $X=13.055 $Y=1.665
+ $X2=0 $Y2=0
cc_938 SET_B N_A_2513_258#_c_1646_n 0.00137814f $X=13.115 $Y=1.58 $X2=0 $Y2=0
cc_939 N_SET_B_c_1234_n N_A_2513_258#_c_1657_n 0.0139984f $X=13.27 $Y=1.97 $X2=0
+ $Y2=0
cc_940 N_SET_B_M1021_g N_A_2513_258#_c_1647_n 0.00109112f $X=13.21 $Y=0.58 $X2=0
+ $Y2=0
cc_941 N_SET_B_c_1222_n N_A_2513_258#_c_1647_n 0.0304377f $X=13.055 $Y=1.665
+ $X2=0 $Y2=0
cc_942 SET_B N_A_2513_258#_c_1647_n 0.00262339f $X=13.115 $Y=1.58 $X2=0 $Y2=0
cc_943 N_SET_B_c_1226_n N_A_2513_258#_c_1647_n 8.82895e-19 $X=13.27 $Y=1.465
+ $X2=0 $Y2=0
cc_944 N_SET_B_c_1227_n N_A_2513_258#_c_1647_n 0.0453809f $X=13.27 $Y=1.465
+ $X2=0 $Y2=0
cc_945 N_SET_B_c_1226_n N_A_2513_258#_c_1648_n 0.0139984f $X=13.27 $Y=1.465
+ $X2=0 $Y2=0
cc_946 N_SET_B_c_1227_n N_A_2513_258#_c_1648_n 0.00347086f $X=13.27 $Y=1.465
+ $X2=0 $Y2=0
cc_947 N_SET_B_M1021_g N_A_2513_258#_c_1649_n 0.0144047f $X=13.21 $Y=0.58 $X2=0
+ $Y2=0
cc_948 N_SET_B_c_1222_n N_A_2513_258#_c_1649_n 0.00543614f $X=13.055 $Y=1.665
+ $X2=0 $Y2=0
cc_949 SET_B N_A_2513_258#_c_1649_n 0.00220758f $X=13.115 $Y=1.58 $X2=0 $Y2=0
cc_950 N_SET_B_c_1226_n N_A_2513_258#_c_1649_n 0.00469569f $X=13.27 $Y=1.465
+ $X2=0 $Y2=0
cc_951 N_SET_B_c_1227_n N_A_2513_258#_c_1649_n 0.0264703f $X=13.27 $Y=1.465
+ $X2=0 $Y2=0
cc_952 N_SET_B_M1021_g N_A_2513_258#_c_1651_n 9.27178e-19 $X=13.21 $Y=0.58 $X2=0
+ $Y2=0
cc_953 N_SET_B_c_1232_n N_A_2513_258#_c_1660_n 9.4089e-19 $X=13.25 $Y=2.465
+ $X2=0 $Y2=0
cc_954 N_SET_B_M1021_g N_A_2067_74#_M1038_g 0.0275785f $X=13.21 $Y=0.58 $X2=0
+ $Y2=0
cc_955 N_SET_B_c_1226_n N_A_2067_74#_c_1758_n 0.0214924f $X=13.27 $Y=1.465 $X2=0
+ $Y2=0
cc_956 N_SET_B_c_1227_n N_A_2067_74#_c_1758_n 0.00245749f $X=13.27 $Y=1.465
+ $X2=0 $Y2=0
cc_957 N_SET_B_c_1222_n N_A_2067_74#_c_1778_n 0.00657317f $X=13.055 $Y=1.665
+ $X2=0 $Y2=0
cc_958 N_SET_B_c_1222_n N_A_2067_74#_c_1805_n 0.00145175f $X=13.055 $Y=1.665
+ $X2=0 $Y2=0
cc_959 N_SET_B_c_1222_n N_A_2067_74#_c_1763_n 0.00295306f $X=13.055 $Y=1.665
+ $X2=0 $Y2=0
cc_960 N_SET_B_c_1231_n N_A_2067_74#_c_1780_n 0.0127766f $X=13.25 $Y=2.375 $X2=0
+ $Y2=0
cc_961 N_SET_B_c_1234_n N_A_2067_74#_c_1780_n 0.00143802f $X=13.27 $Y=1.97 $X2=0
+ $Y2=0
cc_962 N_SET_B_c_1222_n N_A_2067_74#_c_1780_n 0.0135949f $X=13.055 $Y=1.665
+ $X2=0 $Y2=0
cc_963 SET_B N_A_2067_74#_c_1780_n 0.00238877f $X=13.115 $Y=1.58 $X2=0 $Y2=0
cc_964 N_SET_B_c_1227_n N_A_2067_74#_c_1780_n 0.0261515f $X=13.27 $Y=1.465 $X2=0
+ $Y2=0
cc_965 N_SET_B_c_1231_n N_A_2067_74#_c_1781_n 0.00260585f $X=13.25 $Y=2.375
+ $X2=0 $Y2=0
cc_966 N_SET_B_c_1232_n N_A_2067_74#_c_1781_n 0.0121777f $X=13.25 $Y=2.465 $X2=0
+ $Y2=0
cc_967 N_SET_B_c_1231_n N_A_2067_74#_c_1782_n 0.0030803f $X=13.25 $Y=2.375 $X2=0
+ $Y2=0
cc_968 N_SET_B_c_1234_n N_A_2067_74#_c_1782_n 0.00246686f $X=13.27 $Y=1.97 $X2=0
+ $Y2=0
cc_969 N_SET_B_c_1231_n N_A_2067_74#_c_1764_n 0.00106241f $X=13.25 $Y=2.375
+ $X2=0 $Y2=0
cc_970 SET_B N_A_2067_74#_c_1764_n 0.00131157f $X=13.115 $Y=1.58 $X2=0 $Y2=0
cc_971 N_SET_B_c_1226_n N_A_2067_74#_c_1764_n 8.41851e-19 $X=13.27 $Y=1.465
+ $X2=0 $Y2=0
cc_972 N_SET_B_c_1227_n N_A_2067_74#_c_1764_n 0.0411607f $X=13.27 $Y=1.465 $X2=0
+ $Y2=0
cc_973 N_SET_B_c_1231_n N_A_2067_74#_c_1765_n 0.0146339f $X=13.25 $Y=2.375 $X2=0
+ $Y2=0
cc_974 N_SET_B_c_1221_n N_A_2067_74#_c_1765_n 0.0214924f $X=13.27 $Y=1.805 $X2=0
+ $Y2=0
cc_975 N_SET_B_c_1222_n N_A_2067_74#_c_1784_n 0.00914033f $X=13.055 $Y=1.665
+ $X2=0 $Y2=0
cc_976 N_SET_B_c_1222_n N_A_2067_74#_c_1767_n 0.0224912f $X=13.055 $Y=1.665
+ $X2=0 $Y2=0
cc_977 N_SET_B_c_1230_n N_VPWR_c_2062_n 0.00164518f $X=7.985 $Y=2.24 $X2=0 $Y2=0
cc_978 N_SET_B_c_1232_n N_VPWR_c_2064_n 0.00435973f $X=13.25 $Y=2.465 $X2=0
+ $Y2=0
cc_979 N_SET_B_c_1232_n N_VPWR_c_2074_n 0.00445602f $X=13.25 $Y=2.465 $X2=0
+ $Y2=0
cc_980 N_SET_B_c_1232_n N_VPWR_c_2057_n 0.00900303f $X=13.25 $Y=2.465 $X2=0
+ $Y2=0
cc_981 N_SET_B_c_1222_n N_A_1789_424#_c_2379_n 0.00331868f $X=13.055 $Y=1.665
+ $X2=0 $Y2=0
cc_982 N_SET_B_c_1222_n N_A_1789_424#_c_2373_n 0.00160548f $X=13.055 $Y=1.665
+ $X2=0 $Y2=0
cc_983 N_SET_B_c_1222_n N_A_1789_424#_c_2377_n 0.00197494f $X=13.055 $Y=1.665
+ $X2=0 $Y2=0
cc_984 N_SET_B_M1013_g N_VGND_c_2521_n 0.0109278f $X=8.15 $Y=0.58 $X2=0 $Y2=0
cc_985 N_SET_B_M1021_g N_VGND_c_2523_n 0.0125621f $X=13.21 $Y=0.58 $X2=0 $Y2=0
cc_986 N_SET_B_M1021_g N_VGND_c_2533_n 0.00383152f $X=13.21 $Y=0.58 $X2=0 $Y2=0
cc_987 N_SET_B_M1013_g N_VGND_c_2542_n 0.00383152f $X=8.15 $Y=0.58 $X2=0 $Y2=0
cc_988 N_SET_B_M1013_g N_VGND_c_2550_n 0.0075725f $X=8.15 $Y=0.58 $X2=0 $Y2=0
cc_989 N_SET_B_M1021_g N_VGND_c_2550_n 0.0075725f $X=13.21 $Y=0.58 $X2=0 $Y2=0
cc_990 N_A_619_368#_c_1375_n N_A_2513_258#_c_1654_n 0.0167301f $X=12.28 $Y=3.065
+ $X2=0 $Y2=0
cc_991 N_A_619_368#_c_1375_n N_A_2513_258#_c_1655_n 0.012345f $X=12.28 $Y=3.065
+ $X2=0 $Y2=0
cc_992 N_A_619_368#_c_1374_n N_A_2513_258#_M1020_g 0.00691527f $X=12.28 $Y=1.23
+ $X2=0 $Y2=0
cc_993 N_A_619_368#_c_1376_n N_A_2513_258#_M1020_g 0.0445874f $X=12.43 $Y=0.9
+ $X2=0 $Y2=0
cc_994 N_A_619_368#_c_1374_n N_A_2513_258#_c_1647_n 5.5693e-19 $X=12.28 $Y=1.23
+ $X2=0 $Y2=0
cc_995 N_A_619_368#_c_1375_n N_A_2513_258#_c_1647_n 8.7256e-19 $X=12.28 $Y=3.065
+ $X2=0 $Y2=0
cc_996 N_A_619_368#_c_1375_n N_A_2513_258#_c_1648_n 0.0424432f $X=12.28 $Y=3.065
+ $X2=0 $Y2=0
cc_997 N_A_619_368#_c_1374_n N_A_2513_258#_c_1650_n 0.00113941f $X=12.28 $Y=1.23
+ $X2=0 $Y2=0
cc_998 N_A_619_368#_c_1396_n N_A_2067_74#_c_1804_n 0.00615139f $X=10.265
+ $Y=2.045 $X2=0 $Y2=0
cc_999 N_A_619_368#_c_1399_n N_A_2067_74#_c_1804_n 0.00513213f $X=10.715
+ $Y=2.045 $X2=0 $Y2=0
cc_1000 N_A_619_368#_c_1397_n N_A_2067_74#_c_1778_n 5.44415e-19 $X=10.64 $Y=1.97
+ $X2=0 $Y2=0
cc_1001 N_A_619_368#_c_1399_n N_A_2067_74#_c_1778_n 0.0129968f $X=10.715
+ $Y=2.045 $X2=0 $Y2=0
cc_1002 N_A_619_368#_c_1400_n N_A_2067_74#_c_1778_n 0.00783144f $X=11.16 $Y=1.97
+ $X2=0 $Y2=0
cc_1003 N_A_619_368#_c_1401_n N_A_2067_74#_c_1778_n 0.0136823f $X=11.235
+ $Y=3.065 $X2=0 $Y2=0
cc_1004 N_A_619_368#_c_1409_n N_A_2067_74#_c_1778_n 0.00129623f $X=10.715
+ $Y=1.97 $X2=0 $Y2=0
cc_1005 N_A_619_368#_c_1413_n N_A_2067_74#_c_1778_n 0.0845967f $X=11.72 $Y=1.785
+ $X2=0 $Y2=0
cc_1006 N_A_619_368#_c_1396_n N_A_2067_74#_c_1805_n 0.00425563f $X=10.265
+ $Y=2.045 $X2=0 $Y2=0
cc_1007 N_A_619_368#_c_1397_n N_A_2067_74#_c_1805_n 0.00486803f $X=10.64 $Y=1.97
+ $X2=0 $Y2=0
cc_1008 N_A_619_368#_c_1398_n N_A_2067_74#_c_1805_n 2.09189e-19 $X=10.34 $Y=1.97
+ $X2=0 $Y2=0
cc_1009 N_A_619_368#_c_1413_n N_A_2067_74#_c_1805_n 0.0184869f $X=11.72 $Y=1.785
+ $X2=0 $Y2=0
cc_1010 N_A_619_368#_c_1376_n N_A_2067_74#_c_1841_n 0.00697999f $X=12.43 $Y=0.9
+ $X2=0 $Y2=0
cc_1011 N_A_619_368#_c_1380_n N_A_2067_74#_c_1841_n 0.00936164f $X=12.205
+ $Y=1.065 $X2=0 $Y2=0
cc_1012 N_A_619_368#_c_1384_n N_A_2067_74#_c_1841_n 0.0270286f $X=11.885
+ $Y=1.065 $X2=0 $Y2=0
cc_1013 N_A_619_368#_c_1380_n N_A_2067_74#_c_1763_n 0.00342686f $X=12.205
+ $Y=1.065 $X2=0 $Y2=0
cc_1014 N_A_619_368#_c_1413_n N_A_2067_74#_c_1763_n 0.00260498f $X=11.72
+ $Y=1.785 $X2=0 $Y2=0
cc_1015 N_A_619_368#_c_1384_n N_A_2067_74#_c_1763_n 0.00977037f $X=11.885
+ $Y=1.065 $X2=0 $Y2=0
cc_1016 N_A_619_368#_c_1375_n N_A_2067_74#_c_1779_n 0.0120424f $X=12.28 $Y=3.065
+ $X2=0 $Y2=0
cc_1017 N_A_619_368#_c_1375_n N_A_2067_74#_c_1780_n 5.21162e-19 $X=12.28
+ $Y=3.065 $X2=0 $Y2=0
cc_1018 N_A_619_368#_c_1401_n N_A_2067_74#_c_1784_n 8.84397e-19 $X=11.235
+ $Y=3.065 $X2=0 $Y2=0
cc_1019 N_A_619_368#_c_1375_n N_A_2067_74#_c_1784_n 0.0132729f $X=12.28 $Y=3.065
+ $X2=0 $Y2=0
cc_1020 N_A_619_368#_c_1413_n N_A_2067_74#_c_1784_n 0.0197333f $X=11.72 $Y=1.785
+ $X2=0 $Y2=0
cc_1021 N_A_619_368#_c_1374_n N_A_2067_74#_c_1767_n 0.01572f $X=12.28 $Y=1.23
+ $X2=0 $Y2=0
cc_1022 N_A_619_368#_c_1375_n N_A_2067_74#_c_1767_n 0.0183062f $X=12.28 $Y=3.065
+ $X2=0 $Y2=0
cc_1023 N_A_619_368#_c_1376_n N_A_2067_74#_c_1767_n 0.00528607f $X=12.43 $Y=0.9
+ $X2=0 $Y2=0
cc_1024 N_A_619_368#_c_1413_n N_A_2067_74#_c_1767_n 0.0133324f $X=11.72 $Y=1.785
+ $X2=0 $Y2=0
cc_1025 N_A_619_368#_c_1384_n N_A_2067_74#_c_1767_n 0.0582461f $X=11.885
+ $Y=1.065 $X2=0 $Y2=0
cc_1026 N_A_619_368#_c_1411_n N_VPWR_M1026_d 0.00859857f $X=4.39 $Y=1.875 $X2=0
+ $Y2=0
cc_1027 N_A_619_368#_c_1392_n N_VPWR_c_2060_n 8.89341e-19 $X=5.93 $Y=3.075 $X2=0
+ $Y2=0
cc_1028 N_A_619_368#_c_1394_n N_VPWR_c_2060_n 0.0392349f $X=8.72 $Y=3.15 $X2=0
+ $Y2=0
cc_1029 N_A_619_368#_c_1394_n N_VPWR_c_2061_n 0.0322942f $X=8.72 $Y=3.15 $X2=0
+ $Y2=0
cc_1030 N_A_619_368#_c_1394_n N_VPWR_c_2062_n 0.0244731f $X=8.72 $Y=3.15 $X2=0
+ $Y2=0
cc_1031 N_A_619_368#_c_1395_n N_VPWR_c_2062_n 0.0130062f $X=8.795 $Y=3.075 $X2=0
+ $Y2=0
cc_1032 N_A_619_368#_c_1394_n N_VPWR_c_2063_n 0.0020984f $X=8.72 $Y=3.15 $X2=0
+ $Y2=0
cc_1033 N_A_619_368#_c_1395_n N_VPWR_c_2063_n 6.12794e-19 $X=8.795 $Y=3.075
+ $X2=0 $Y2=0
cc_1034 N_A_619_368#_c_1375_n N_VPWR_c_2064_n 0.00189808f $X=12.28 $Y=3.065
+ $X2=0 $Y2=0
cc_1035 N_A_619_368#_c_1394_n N_VPWR_c_2070_n 0.00796123f $X=8.72 $Y=3.15 $X2=0
+ $Y2=0
cc_1036 N_A_619_368#_c_1396_n N_VPWR_c_2072_n 0.00278271f $X=10.265 $Y=2.045
+ $X2=0 $Y2=0
cc_1037 N_A_619_368#_c_1399_n N_VPWR_c_2072_n 0.00278257f $X=10.715 $Y=2.045
+ $X2=0 $Y2=0
cc_1038 N_A_619_368#_c_1403_n N_VPWR_c_2072_n 0.0286449f $X=11.31 $Y=3.14 $X2=0
+ $Y2=0
cc_1039 N_A_619_368#_c_1387_n N_VPWR_c_2080_n 0.00460063f $X=4.295 $Y=1.765
+ $X2=0 $Y2=0
cc_1040 N_A_619_368#_c_1390_n N_VPWR_c_2080_n 0.0376041f $X=4.925 $Y=3.15 $X2=0
+ $Y2=0
cc_1041 N_A_619_368#_c_1387_n N_VPWR_c_2086_n 0.00214719f $X=4.295 $Y=1.765
+ $X2=0 $Y2=0
cc_1042 N_A_619_368#_c_1390_n N_VPWR_c_2086_n 0.00232313f $X=4.925 $Y=3.15 $X2=0
+ $Y2=0
cc_1043 N_A_619_368#_c_1387_n N_VPWR_c_2057_n 0.00905135f $X=4.295 $Y=1.765
+ $X2=0 $Y2=0
cc_1044 N_A_619_368#_c_1389_n N_VPWR_c_2057_n 0.0215278f $X=5.84 $Y=3.15 $X2=0
+ $Y2=0
cc_1045 N_A_619_368#_c_1390_n N_VPWR_c_2057_n 0.00600348f $X=4.925 $Y=3.15 $X2=0
+ $Y2=0
cc_1046 N_A_619_368#_c_1394_n N_VPWR_c_2057_n 0.0676097f $X=8.72 $Y=3.15 $X2=0
+ $Y2=0
cc_1047 N_A_619_368#_c_1396_n N_VPWR_c_2057_n 0.00353907f $X=10.265 $Y=2.045
+ $X2=0 $Y2=0
cc_1048 N_A_619_368#_c_1399_n N_VPWR_c_2057_n 0.00354455f $X=10.715 $Y=2.045
+ $X2=0 $Y2=0
cc_1049 N_A_619_368#_c_1402_n N_VPWR_c_2057_n 0.0290175f $X=12.205 $Y=3.14 $X2=0
+ $Y2=0
cc_1050 N_A_619_368#_c_1403_n N_VPWR_c_2057_n 0.0114051f $X=11.31 $Y=3.14 $X2=0
+ $Y2=0
cc_1051 N_A_619_368#_c_1408_n N_VPWR_c_2057_n 0.00441524f $X=5.93 $Y=3.15 $X2=0
+ $Y2=0
cc_1052 N_A_619_368#_c_1414_n N_A_304_464#_c_2257_n 0.0143692f $X=3.545 $Y=1.965
+ $X2=0 $Y2=0
cc_1053 N_A_619_368#_M1026_s N_A_304_464#_c_2262_n 0.00840263f $X=3.095 $Y=1.84
+ $X2=0 $Y2=0
cc_1054 N_A_619_368#_c_1411_n N_A_304_464#_c_2262_n 0.00504085f $X=4.39 $Y=1.875
+ $X2=0 $Y2=0
cc_1055 N_A_619_368#_c_1414_n N_A_304_464#_c_2262_n 0.0305907f $X=3.545 $Y=1.965
+ $X2=0 $Y2=0
cc_1056 N_A_619_368#_c_1387_n N_A_304_464#_c_2263_n 0.0166148f $X=4.295 $Y=1.765
+ $X2=0 $Y2=0
cc_1057 N_A_619_368#_c_1388_n N_A_304_464#_c_2263_n 0.0132298f $X=4.85 $Y=3.075
+ $X2=0 $Y2=0
cc_1058 N_A_619_368#_c_1378_n N_A_304_464#_c_2263_n 0.00289212f $X=4.775
+ $Y=1.515 $X2=0 $Y2=0
cc_1059 N_A_619_368#_c_1411_n N_A_304_464#_c_2263_n 0.054049f $X=4.39 $Y=1.875
+ $X2=0 $Y2=0
cc_1060 N_A_619_368#_c_1387_n N_A_304_464#_c_2300_n 0.00367629f $X=4.295
+ $Y=1.765 $X2=0 $Y2=0
cc_1061 N_A_619_368#_c_1411_n N_A_304_464#_c_2300_n 0.0129609f $X=4.39 $Y=1.875
+ $X2=0 $Y2=0
cc_1062 N_A_619_368#_c_1371_n N_A_304_464#_c_2258_n 0.00547833f $X=5.195
+ $Y=0.975 $X2=0 $Y2=0
cc_1063 N_A_619_368#_c_1373_n N_A_304_464#_c_2258_n 0.00434355f $X=5.27 $Y=0.9
+ $X2=0 $Y2=0
cc_1064 N_A_619_368#_c_1387_n N_A_304_464#_c_2265_n 9.31521e-19 $X=4.295
+ $Y=1.765 $X2=0 $Y2=0
cc_1065 N_A_619_368#_c_1388_n N_A_304_464#_c_2265_n 0.0178623f $X=4.85 $Y=3.075
+ $X2=0 $Y2=0
cc_1066 N_A_619_368#_c_1393_n N_A_304_464#_c_2265_n 2.23037e-19 $X=5.93 $Y=2.81
+ $X2=0 $Y2=0
cc_1067 N_A_619_368#_M1033_g N_A_304_464#_c_2259_n 0.00150815f $X=4.28 $Y=0.74
+ $X2=0 $Y2=0
cc_1068 N_A_619_368#_c_1387_n N_A_304_464#_c_2259_n 9.26169e-19 $X=4.295
+ $Y=1.765 $X2=0 $Y2=0
cc_1069 N_A_619_368#_c_1370_n N_A_304_464#_c_2259_n 0.00891258f $X=4.85 $Y=1.35
+ $X2=0 $Y2=0
cc_1070 N_A_619_368#_c_1388_n N_A_304_464#_c_2259_n 0.0105856f $X=4.85 $Y=3.075
+ $X2=0 $Y2=0
cc_1071 N_A_619_368#_c_1371_n N_A_304_464#_c_2259_n 0.0101656f $X=5.195 $Y=0.975
+ $X2=0 $Y2=0
cc_1072 N_A_619_368#_c_1372_n N_A_304_464#_c_2259_n 0.00285843f $X=4.925
+ $Y=0.975 $X2=0 $Y2=0
cc_1073 N_A_619_368#_c_1379_n N_A_304_464#_c_2259_n 0.00807793f $X=4.85 $Y=1.515
+ $X2=0 $Y2=0
cc_1074 N_A_619_368#_c_1411_n N_A_304_464#_c_2259_n 0.0137141f $X=4.39 $Y=1.875
+ $X2=0 $Y2=0
cc_1075 N_A_619_368#_c_1383_n N_A_304_464#_c_2259_n 0.0317952f $X=4.555 $Y=1.515
+ $X2=0 $Y2=0
cc_1076 N_A_619_368#_c_1413_n N_A_1789_424#_c_2379_n 0.0252478f $X=11.72
+ $Y=1.785 $X2=0 $Y2=0
cc_1077 N_A_619_368#_c_1396_n N_A_1789_424#_c_2373_n 9.34633e-19 $X=10.265
+ $Y=2.045 $X2=0 $Y2=0
cc_1078 N_A_619_368#_c_1413_n N_A_1789_424#_c_2373_n 0.015045f $X=11.72 $Y=1.785
+ $X2=0 $Y2=0
cc_1079 N_A_619_368#_c_1396_n N_A_1789_424#_c_2382_n 0.00396311f $X=10.265
+ $Y=2.045 $X2=0 $Y2=0
cc_1080 N_A_619_368#_c_1396_n N_A_1789_424#_c_2374_n 0.0127761f $X=10.265
+ $Y=2.045 $X2=0 $Y2=0
cc_1081 N_A_619_368#_c_1399_n N_A_1789_424#_c_2374_n 0.0125787f $X=10.715
+ $Y=2.045 $X2=0 $Y2=0
cc_1082 N_A_619_368#_c_1401_n N_A_1789_424#_c_2374_n 0.00232564f $X=11.235
+ $Y=3.065 $X2=0 $Y2=0
cc_1083 N_A_619_368#_c_1396_n N_A_1789_424#_c_2376_n 7.39945e-19 $X=10.265
+ $Y=2.045 $X2=0 $Y2=0
cc_1084 N_A_619_368#_c_1399_n N_A_1789_424#_c_2376_n 0.00725376f $X=10.715
+ $Y=2.045 $X2=0 $Y2=0
cc_1085 N_A_619_368#_c_1400_n N_A_1789_424#_c_2376_n 0.00102765f $X=11.16
+ $Y=1.97 $X2=0 $Y2=0
cc_1086 N_A_619_368#_c_1401_n N_A_1789_424#_c_2376_n 0.00538716f $X=11.235
+ $Y=3.065 $X2=0 $Y2=0
cc_1087 N_A_619_368#_c_1395_n N_A_1789_424#_c_2377_n 0.0127671f $X=8.795
+ $Y=3.075 $X2=0 $Y2=0
cc_1088 N_A_619_368#_c_1413_n N_A_1789_424#_c_2377_n 0.00958835f $X=11.72
+ $Y=1.785 $X2=0 $Y2=0
cc_1089 N_A_619_368#_c_1386_n N_A_1789_424#_c_2377_n 0.00326139f $X=8.9 $Y=1.795
+ $X2=0 $Y2=0
cc_1090 N_A_619_368#_c_1416_n N_A_1789_424#_c_2377_n 0.0108129f $X=9.065
+ $Y=1.822 $X2=0 $Y2=0
cc_1091 N_A_619_368#_c_1401_n N_A_2277_455#_c_2427_n 0.00576301f $X=11.235
+ $Y=3.065 $X2=0 $Y2=0
cc_1092 N_A_619_368#_c_1375_n N_A_2277_455#_c_2427_n 0.00161392f $X=12.28
+ $Y=3.065 $X2=0 $Y2=0
cc_1093 N_A_619_368#_c_1402_n N_A_2277_455#_c_2428_n 0.00922302f $X=12.205
+ $Y=3.14 $X2=0 $Y2=0
cc_1094 N_A_619_368#_c_1375_n N_A_2277_455#_c_2428_n 0.0121403f $X=12.28
+ $Y=3.065 $X2=0 $Y2=0
cc_1095 N_A_619_368#_c_1401_n N_A_2277_455#_c_2429_n 0.00422063f $X=11.235
+ $Y=3.065 $X2=0 $Y2=0
cc_1096 N_A_619_368#_c_1402_n N_A_2277_455#_c_2429_n 0.00545232f $X=12.205
+ $Y=3.14 $X2=0 $Y2=0
cc_1097 N_A_619_368#_c_1375_n N_A_2277_455#_c_2430_n 0.00652254f $X=12.28
+ $Y=3.065 $X2=0 $Y2=0
cc_1098 N_A_619_368#_c_1381_n N_VGND_c_2518_n 0.0316927f $X=3.565 $Y=0.505 $X2=0
+ $Y2=0
cc_1099 N_A_619_368#_M1033_g N_VGND_c_2519_n 0.00470925f $X=4.28 $Y=0.74 $X2=0
+ $Y2=0
cc_1100 N_A_619_368#_c_1381_n N_VGND_c_2519_n 0.025141f $X=3.565 $Y=0.505 $X2=0
+ $Y2=0
cc_1101 N_A_619_368#_c_1376_n N_VGND_c_2533_n 0.0042336f $X=12.43 $Y=0.9 $X2=0
+ $Y2=0
cc_1102 N_A_619_368#_c_1381_n N_VGND_c_2540_n 0.0126849f $X=3.565 $Y=0.505 $X2=0
+ $Y2=0
cc_1103 N_A_619_368#_M1033_g N_VGND_c_2541_n 0.00430908f $X=4.28 $Y=0.74 $X2=0
+ $Y2=0
cc_1104 N_A_619_368#_c_1373_n N_VGND_c_2541_n 9.15902e-19 $X=5.27 $Y=0.9 $X2=0
+ $Y2=0
cc_1105 N_A_619_368#_M1033_g N_VGND_c_2550_n 0.00821169f $X=4.28 $Y=0.74 $X2=0
+ $Y2=0
cc_1106 N_A_619_368#_c_1376_n N_VGND_c_2550_n 0.0078709f $X=12.43 $Y=0.9 $X2=0
+ $Y2=0
cc_1107 N_A_619_368#_c_1381_n N_VGND_c_2550_n 0.0101411f $X=3.565 $Y=0.505 $X2=0
+ $Y2=0
cc_1108 N_A_2513_258#_c_1649_n N_A_2067_74#_M1038_g 0.0115126f $X=13.77 $Y=1.045
+ $X2=0 $Y2=0
cc_1109 N_A_2513_258#_c_1651_n N_A_2067_74#_M1038_g 0.0125515f $X=13.935 $Y=0.58
+ $X2=0 $Y2=0
cc_1110 N_A_2513_258#_c_1652_n N_A_2067_74#_M1038_g 0.00477786f $X=14.23 $Y=2.48
+ $X2=0 $Y2=0
cc_1111 N_A_2513_258#_c_1653_n N_A_2067_74#_M1038_g 0.00461905f $X=14.042
+ $Y=1.045 $X2=0 $Y2=0
cc_1112 N_A_2513_258#_c_1652_n N_A_2067_74#_c_1749_n 0.0153375f $X=14.23 $Y=2.48
+ $X2=0 $Y2=0
cc_1113 N_A_2513_258#_c_1652_n N_A_2067_74#_c_1768_n 0.00325714f $X=14.23
+ $Y=2.48 $X2=0 $Y2=0
cc_1114 N_A_2513_258#_c_1660_n N_A_2067_74#_c_1769_n 0.00897893f $X=14.23
+ $Y=2.695 $X2=0 $Y2=0
cc_1115 N_A_2513_258#_c_1652_n N_A_2067_74#_c_1770_n 0.00348266f $X=14.23
+ $Y=2.48 $X2=0 $Y2=0
cc_1116 N_A_2513_258#_c_1660_n N_A_2067_74#_c_1770_n 0.0100111f $X=14.23
+ $Y=2.695 $X2=0 $Y2=0
cc_1117 N_A_2513_258#_c_1651_n N_A_2067_74#_M1022_g 0.00441492f $X=13.935
+ $Y=0.58 $X2=0 $Y2=0
cc_1118 N_A_2513_258#_c_1652_n N_A_2067_74#_M1022_g 0.0029433f $X=14.23 $Y=2.48
+ $X2=0 $Y2=0
cc_1119 N_A_2513_258#_c_1653_n N_A_2067_74#_M1022_g 0.00323313f $X=14.042
+ $Y=1.045 $X2=0 $Y2=0
cc_1120 N_A_2513_258#_c_1652_n N_A_2067_74#_c_1751_n 0.00563716f $X=14.23
+ $Y=2.48 $X2=0 $Y2=0
cc_1121 N_A_2513_258#_c_1652_n N_A_2067_74#_c_1772_n 0.00140669f $X=14.23
+ $Y=2.48 $X2=0 $Y2=0
cc_1122 N_A_2513_258#_c_1653_n N_A_2067_74#_c_1758_n 0.0080581f $X=14.042
+ $Y=1.045 $X2=0 $Y2=0
cc_1123 N_A_2513_258#_c_1652_n N_A_2067_74#_c_1777_n 0.0090141f $X=14.23 $Y=2.48
+ $X2=0 $Y2=0
cc_1124 N_A_2513_258#_M1020_g N_A_2067_74#_c_1841_n 0.00165231f $X=12.82 $Y=0.58
+ $X2=0 $Y2=0
cc_1125 N_A_2513_258#_c_1654_n N_A_2067_74#_c_1779_n 7.26962e-19 $X=12.8
+ $Y=2.375 $X2=0 $Y2=0
cc_1126 N_A_2513_258#_c_1655_n N_A_2067_74#_c_1779_n 3.13134e-19 $X=12.8
+ $Y=2.465 $X2=0 $Y2=0
cc_1127 N_A_2513_258#_c_1654_n N_A_2067_74#_c_1780_n 0.0162892f $X=12.8 $Y=2.375
+ $X2=0 $Y2=0
cc_1128 N_A_2513_258#_c_1657_n N_A_2067_74#_c_1780_n 9.90657e-19 $X=12.73
+ $Y=1.96 $X2=0 $Y2=0
cc_1129 N_A_2513_258#_c_1647_n N_A_2067_74#_c_1780_n 0.0231756f $X=12.73
+ $Y=1.455 $X2=0 $Y2=0
cc_1130 N_A_2513_258#_c_1654_n N_A_2067_74#_c_1781_n 7.33041e-19 $X=12.8
+ $Y=2.375 $X2=0 $Y2=0
cc_1131 N_A_2513_258#_c_1655_n N_A_2067_74#_c_1781_n 3.96182e-19 $X=12.8
+ $Y=2.465 $X2=0 $Y2=0
cc_1132 N_A_2513_258#_c_1652_n N_A_2067_74#_c_1781_n 0.00614787f $X=14.23
+ $Y=2.48 $X2=0 $Y2=0
cc_1133 N_A_2513_258#_c_1660_n N_A_2067_74#_c_1781_n 0.0296215f $X=14.23
+ $Y=2.695 $X2=0 $Y2=0
cc_1134 N_A_2513_258#_c_1652_n N_A_2067_74#_c_1782_n 0.0128267f $X=14.23 $Y=2.48
+ $X2=0 $Y2=0
cc_1135 N_A_2513_258#_c_1660_n N_A_2067_74#_c_1782_n 0.00797082f $X=14.23
+ $Y=2.695 $X2=0 $Y2=0
cc_1136 N_A_2513_258#_c_1649_n N_A_2067_74#_c_1764_n 0.00941168f $X=13.77
+ $Y=1.045 $X2=0 $Y2=0
cc_1137 N_A_2513_258#_c_1652_n N_A_2067_74#_c_1764_n 0.062535f $X=14.23 $Y=2.48
+ $X2=0 $Y2=0
cc_1138 N_A_2513_258#_c_1653_n N_A_2067_74#_c_1764_n 0.0180767f $X=14.042
+ $Y=1.045 $X2=0 $Y2=0
cc_1139 N_A_2513_258#_c_1652_n N_A_2067_74#_c_1765_n 0.0118829f $X=14.23 $Y=2.48
+ $X2=0 $Y2=0
cc_1140 N_A_2513_258#_c_1654_n N_A_2067_74#_c_1767_n 0.00372173f $X=12.8
+ $Y=2.375 $X2=0 $Y2=0
cc_1141 N_A_2513_258#_M1020_g N_A_2067_74#_c_1767_n 0.00178906f $X=12.82 $Y=0.58
+ $X2=0 $Y2=0
cc_1142 N_A_2513_258#_c_1647_n N_A_2067_74#_c_1767_n 0.0605029f $X=12.73
+ $Y=1.455 $X2=0 $Y2=0
cc_1143 N_A_2513_258#_c_1648_n N_A_2067_74#_c_1767_n 0.0033491f $X=12.73
+ $Y=1.455 $X2=0 $Y2=0
cc_1144 N_A_2513_258#_c_1650_n N_A_2067_74#_c_1767_n 0.0137215f $X=12.895
+ $Y=1.045 $X2=0 $Y2=0
cc_1145 N_A_2513_258#_c_1655_n N_VPWR_c_2064_n 0.00313576f $X=12.8 $Y=2.465
+ $X2=0 $Y2=0
cc_1146 N_A_2513_258#_c_1652_n N_VPWR_c_2065_n 0.0476065f $X=14.23 $Y=2.48 $X2=0
+ $Y2=0
cc_1147 N_A_2513_258#_c_1660_n N_VPWR_c_2065_n 0.0325138f $X=14.23 $Y=2.695
+ $X2=0 $Y2=0
cc_1148 N_A_2513_258#_c_1655_n N_VPWR_c_2072_n 0.00443421f $X=12.8 $Y=2.465
+ $X2=0 $Y2=0
cc_1149 N_A_2513_258#_c_1660_n N_VPWR_c_2074_n 0.0145873f $X=14.23 $Y=2.695
+ $X2=0 $Y2=0
cc_1150 N_A_2513_258#_c_1655_n N_VPWR_c_2057_n 0.00891991f $X=12.8 $Y=2.465
+ $X2=0 $Y2=0
cc_1151 N_A_2513_258#_c_1660_n N_VPWR_c_2057_n 0.0153199f $X=14.23 $Y=2.695
+ $X2=0 $Y2=0
cc_1152 N_A_2513_258#_c_1655_n N_A_2277_455#_c_2428_n 0.00342208f $X=12.8
+ $Y=2.465 $X2=0 $Y2=0
cc_1153 N_A_2513_258#_c_1655_n N_A_2277_455#_c_2430_n 0.00483823f $X=12.8
+ $Y=2.465 $X2=0 $Y2=0
cc_1154 N_A_2513_258#_c_1652_n N_Q_N_c_2460_n 0.0210324f $X=14.23 $Y=2.48 $X2=0
+ $Y2=0
cc_1155 N_A_2513_258#_c_1653_n N_Q_N_c_2460_n 0.00612134f $X=14.042 $Y=1.045
+ $X2=0 $Y2=0
cc_1156 N_A_2513_258#_M1020_g N_VGND_c_2523_n 0.00274214f $X=12.82 $Y=0.58 $X2=0
+ $Y2=0
cc_1157 N_A_2513_258#_c_1649_n N_VGND_c_2523_n 0.0243627f $X=13.77 $Y=1.045
+ $X2=0 $Y2=0
cc_1158 N_A_2513_258#_c_1651_n N_VGND_c_2523_n 0.0165294f $X=13.935 $Y=0.58
+ $X2=0 $Y2=0
cc_1159 N_A_2513_258#_c_1651_n N_VGND_c_2524_n 0.0280059f $X=13.935 $Y=0.58
+ $X2=0 $Y2=0
cc_1160 N_A_2513_258#_M1020_g N_VGND_c_2533_n 0.00461464f $X=12.82 $Y=0.58 $X2=0
+ $Y2=0
cc_1161 N_A_2513_258#_c_1651_n N_VGND_c_2535_n 0.0145639f $X=13.935 $Y=0.58
+ $X2=0 $Y2=0
cc_1162 N_A_2513_258#_M1020_g N_VGND_c_2550_n 0.00908738f $X=12.82 $Y=0.58 $X2=0
+ $Y2=0
cc_1163 N_A_2513_258#_c_1651_n N_VGND_c_2550_n 0.0119984f $X=13.935 $Y=0.58
+ $X2=0 $Y2=0
cc_1164 N_A_2067_74#_c_1776_n N_A_3177_368#_c_1995_n 0.0144116f $X=16.255
+ $Y=1.765 $X2=0 $Y2=0
cc_1165 N_A_2067_74#_M1010_g N_A_3177_368#_M1023_g 0.0139828f $X=16.27 $Y=0.79
+ $X2=0 $Y2=0
cc_1166 N_A_2067_74#_M1025_g N_A_3177_368#_c_1990_n 0.00365834f $X=15.23 $Y=0.74
+ $X2=0 $Y2=0
cc_1167 N_A_2067_74#_M1010_g N_A_3177_368#_c_1990_n 0.016091f $X=16.27 $Y=0.79
+ $X2=0 $Y2=0
cc_1168 N_A_2067_74#_c_1754_n N_A_3177_368#_c_1991_n 0.00347777f $X=15.245
+ $Y=1.675 $X2=0 $Y2=0
cc_1169 N_A_2067_74#_c_1774_n N_A_3177_368#_c_1991_n 0.00329382f $X=15.245
+ $Y=1.765 $X2=0 $Y2=0
cc_1170 N_A_2067_74#_c_1756_n N_A_3177_368#_c_1991_n 0.00175408f $X=16.255
+ $Y=1.675 $X2=0 $Y2=0
cc_1171 N_A_2067_74#_c_1776_n N_A_3177_368#_c_1991_n 0.018379f $X=16.255
+ $Y=1.765 $X2=0 $Y2=0
cc_1172 N_A_2067_74#_c_1756_n N_A_3177_368#_c_1992_n 0.00950208f $X=16.255
+ $Y=1.675 $X2=0 $Y2=0
cc_1173 N_A_2067_74#_c_1761_n N_A_3177_368#_c_1992_n 0.0090289f $X=16.255
+ $Y=1.375 $X2=0 $Y2=0
cc_1174 N_A_2067_74#_c_1754_n N_A_3177_368#_c_1993_n 0.00515495f $X=15.245
+ $Y=1.675 $X2=0 $Y2=0
cc_1175 N_A_2067_74#_c_1755_n N_A_3177_368#_c_1993_n 0.0204535f $X=16.165
+ $Y=1.375 $X2=0 $Y2=0
cc_1176 N_A_2067_74#_c_1756_n N_A_3177_368#_c_1993_n 0.00582757f $X=16.255
+ $Y=1.675 $X2=0 $Y2=0
cc_1177 N_A_2067_74#_c_1761_n N_A_3177_368#_c_1993_n 7.76856e-19 $X=16.255
+ $Y=1.375 $X2=0 $Y2=0
cc_1178 N_A_2067_74#_c_1756_n N_A_3177_368#_c_1994_n 0.00476504f $X=16.255
+ $Y=1.675 $X2=0 $Y2=0
cc_1179 N_A_2067_74#_c_1761_n N_A_3177_368#_c_1994_n 0.0214984f $X=16.255
+ $Y=1.375 $X2=0 $Y2=0
cc_1180 N_A_2067_74#_c_1780_n N_VPWR_c_2064_n 0.0122262f $X=13.31 $Y=2.225 $X2=0
+ $Y2=0
cc_1181 N_A_2067_74#_c_1781_n N_VPWR_c_2064_n 0.0300176f $X=13.475 $Y=2.75 $X2=0
+ $Y2=0
cc_1182 N_A_2067_74#_c_1749_n N_VPWR_c_2065_n 0.00428832f $X=14.705 $Y=1.375
+ $X2=0 $Y2=0
cc_1183 N_A_2067_74#_c_1770_n N_VPWR_c_2065_n 0.00601341f $X=14.26 $Y=2.395
+ $X2=0 $Y2=0
cc_1184 N_A_2067_74#_c_1772_n N_VPWR_c_2065_n 0.0067841f $X=14.795 $Y=1.765
+ $X2=0 $Y2=0
cc_1185 N_A_2067_74#_c_1777_n N_VPWR_c_2065_n 0.0019325f $X=14.26 $Y=2.235 $X2=0
+ $Y2=0
cc_1186 N_A_2067_74#_c_1772_n N_VPWR_c_2066_n 7.29261e-19 $X=14.795 $Y=1.765
+ $X2=0 $Y2=0
cc_1187 N_A_2067_74#_c_1774_n N_VPWR_c_2066_n 0.0196894f $X=15.245 $Y=1.765
+ $X2=0 $Y2=0
cc_1188 N_A_2067_74#_c_1755_n N_VPWR_c_2066_n 0.00694774f $X=16.165 $Y=1.375
+ $X2=0 $Y2=0
cc_1189 N_A_2067_74#_c_1776_n N_VPWR_c_2066_n 0.00462006f $X=16.255 $Y=1.765
+ $X2=0 $Y2=0
cc_1190 N_A_2067_74#_c_1776_n N_VPWR_c_2067_n 0.0122251f $X=16.255 $Y=1.765
+ $X2=0 $Y2=0
cc_1191 N_A_2067_74#_c_1770_n N_VPWR_c_2074_n 0.00402251f $X=14.26 $Y=2.395
+ $X2=0 $Y2=0
cc_1192 N_A_2067_74#_c_1781_n N_VPWR_c_2074_n 0.0145781f $X=13.475 $Y=2.75 $X2=0
+ $Y2=0
cc_1193 N_A_2067_74#_c_1772_n N_VPWR_c_2076_n 0.00439937f $X=14.795 $Y=1.765
+ $X2=0 $Y2=0
cc_1194 N_A_2067_74#_c_1774_n N_VPWR_c_2076_n 0.00413917f $X=15.245 $Y=1.765
+ $X2=0 $Y2=0
cc_1195 N_A_2067_74#_c_1776_n N_VPWR_c_2081_n 0.00481995f $X=16.255 $Y=1.765
+ $X2=0 $Y2=0
cc_1196 N_A_2067_74#_c_1770_n N_VPWR_c_2057_n 0.00523671f $X=14.26 $Y=2.395
+ $X2=0 $Y2=0
cc_1197 N_A_2067_74#_c_1772_n N_VPWR_c_2057_n 0.00844048f $X=14.795 $Y=1.765
+ $X2=0 $Y2=0
cc_1198 N_A_2067_74#_c_1774_n N_VPWR_c_2057_n 0.00817726f $X=15.245 $Y=1.765
+ $X2=0 $Y2=0
cc_1199 N_A_2067_74#_c_1776_n N_VPWR_c_2057_n 0.00508379f $X=16.255 $Y=1.765
+ $X2=0 $Y2=0
cc_1200 N_A_2067_74#_c_1781_n N_VPWR_c_2057_n 0.0120405f $X=13.475 $Y=2.75 $X2=0
+ $Y2=0
cc_1201 N_A_2067_74#_c_1778_n N_A_1789_424#_M1046_d 0.00252999f $X=11.82
+ $Y=2.125 $X2=0 $Y2=0
cc_1202 N_A_2067_74#_c_1804_n N_A_1789_424#_c_2373_n 0.00639933f $X=10.49
+ $Y=2.46 $X2=0 $Y2=0
cc_1203 N_A_2067_74#_c_1805_n N_A_1789_424#_c_2373_n 0.00833572f $X=10.575
+ $Y=2.125 $X2=0 $Y2=0
cc_1204 N_A_2067_74#_c_1804_n N_A_1789_424#_c_2382_n 0.0262374f $X=10.49 $Y=2.46
+ $X2=0 $Y2=0
cc_1205 N_A_2067_74#_M1005_s N_A_1789_424#_c_2374_n 0.00238308f $X=10.34 $Y=2.12
+ $X2=0 $Y2=0
cc_1206 N_A_2067_74#_c_1804_n N_A_1789_424#_c_2374_n 0.0122792f $X=10.49 $Y=2.46
+ $X2=0 $Y2=0
cc_1207 N_A_2067_74#_c_1804_n N_A_1789_424#_c_2376_n 0.0214564f $X=10.49 $Y=2.46
+ $X2=0 $Y2=0
cc_1208 N_A_2067_74#_c_1778_n N_A_1789_424#_c_2376_n 0.0220317f $X=11.82
+ $Y=2.125 $X2=0 $Y2=0
cc_1209 N_A_2067_74#_c_1778_n N_A_2277_455#_c_2427_n 0.0204912f $X=11.82
+ $Y=2.125 $X2=0 $Y2=0
cc_1210 N_A_2067_74#_c_1779_n N_A_2277_455#_c_2427_n 0.0225147f $X=11.985
+ $Y=2.485 $X2=0 $Y2=0
cc_1211 N_A_2067_74#_c_1778_n N_A_2277_455#_c_2428_n 0.00519337f $X=11.82
+ $Y=2.125 $X2=0 $Y2=0
cc_1212 N_A_2067_74#_c_1779_n N_A_2277_455#_c_2428_n 0.0313945f $X=11.985
+ $Y=2.485 $X2=0 $Y2=0
cc_1213 N_A_2067_74#_c_1780_n N_A_2277_455#_c_2428_n 6.30153e-19 $X=13.31
+ $Y=2.225 $X2=0 $Y2=0
cc_1214 N_A_2067_74#_c_1784_n N_A_2277_455#_c_2428_n 0.0049692f $X=12.105
+ $Y=2.125 $X2=0 $Y2=0
cc_1215 N_A_2067_74#_c_1779_n N_A_2277_455#_c_2430_n 0.0143942f $X=11.985
+ $Y=2.485 $X2=0 $Y2=0
cc_1216 N_A_2067_74#_c_1780_n N_A_2277_455#_c_2430_n 0.0232278f $X=13.31
+ $Y=2.225 $X2=0 $Y2=0
cc_1217 N_A_2067_74#_c_1751_n N_Q_N_c_2459_n 0.00664874f $X=14.795 $Y=1.675
+ $X2=0 $Y2=0
cc_1218 N_A_2067_74#_c_1772_n N_Q_N_c_2459_n 0.0180168f $X=14.795 $Y=1.765 $X2=0
+ $Y2=0
cc_1219 N_A_2067_74#_c_1752_n N_Q_N_c_2459_n 0.00477651f $X=15.155 $Y=1.375
+ $X2=0 $Y2=0
cc_1220 N_A_2067_74#_c_1754_n N_Q_N_c_2459_n 0.00817929f $X=15.245 $Y=1.675
+ $X2=0 $Y2=0
cc_1221 N_A_2067_74#_c_1774_n N_Q_N_c_2459_n 0.00582203f $X=15.245 $Y=1.765
+ $X2=0 $Y2=0
cc_1222 N_A_2067_74#_c_1759_n N_Q_N_c_2459_n 0.00114549f $X=14.795 $Y=1.375
+ $X2=0 $Y2=0
cc_1223 N_A_2067_74#_M1022_g N_Q_N_c_2460_n 0.0183249f $X=14.78 $Y=0.74 $X2=0
+ $Y2=0
cc_1224 N_A_2067_74#_M1025_g N_Q_N_c_2460_n 0.0165206f $X=15.23 $Y=0.74 $X2=0
+ $Y2=0
cc_1225 N_A_2067_74#_M1022_g Q_N 0.00250547f $X=14.78 $Y=0.74 $X2=0 $Y2=0
cc_1226 N_A_2067_74#_c_1752_n Q_N 0.00824205f $X=15.155 $Y=1.375 $X2=0 $Y2=0
cc_1227 N_A_2067_74#_M1025_g Q_N 0.00308648f $X=15.23 $Y=0.74 $X2=0 $Y2=0
cc_1228 N_A_2067_74#_c_1759_n Q_N 0.0032858f $X=14.795 $Y=1.375 $X2=0 $Y2=0
cc_1229 N_A_2067_74#_c_1760_n Q_N 0.00804947f $X=15.245 $Y=1.375 $X2=0 $Y2=0
cc_1230 N_A_2067_74#_M1038_g N_VGND_c_2523_n 0.0054334f $X=13.72 $Y=0.58 $X2=0
+ $Y2=0
cc_1231 N_A_2067_74#_M1038_g N_VGND_c_2524_n 0.00358244f $X=13.72 $Y=0.58 $X2=0
+ $Y2=0
cc_1232 N_A_2067_74#_c_1749_n N_VGND_c_2524_n 0.00760021f $X=14.705 $Y=1.375
+ $X2=0 $Y2=0
cc_1233 N_A_2067_74#_M1022_g N_VGND_c_2524_n 0.00639614f $X=14.78 $Y=0.74 $X2=0
+ $Y2=0
cc_1234 N_A_2067_74#_M1025_g N_VGND_c_2525_n 0.00819758f $X=15.23 $Y=0.74 $X2=0
+ $Y2=0
cc_1235 N_A_2067_74#_c_1755_n N_VGND_c_2525_n 0.0103331f $X=16.165 $Y=1.375
+ $X2=0 $Y2=0
cc_1236 N_A_2067_74#_M1010_g N_VGND_c_2525_n 0.00377536f $X=16.27 $Y=0.79 $X2=0
+ $Y2=0
cc_1237 N_A_2067_74#_M1010_g N_VGND_c_2526_n 0.00886999f $X=16.27 $Y=0.79 $X2=0
+ $Y2=0
cc_1238 N_A_2067_74#_c_1841_n N_VGND_c_2533_n 0.0279753f $X=12.22 $Y=0.565 $X2=0
+ $Y2=0
cc_1239 N_A_2067_74#_c_1763_n N_VGND_c_2533_n 0.00610577f $X=11.55 $Y=0.565
+ $X2=0 $Y2=0
cc_1240 N_A_2067_74#_M1038_g N_VGND_c_2535_n 0.00434272f $X=13.72 $Y=0.58 $X2=0
+ $Y2=0
cc_1241 N_A_2067_74#_M1022_g N_VGND_c_2537_n 0.00456932f $X=14.78 $Y=0.74 $X2=0
+ $Y2=0
cc_1242 N_A_2067_74#_M1025_g N_VGND_c_2537_n 0.00371957f $X=15.23 $Y=0.74 $X2=0
+ $Y2=0
cc_1243 N_A_2067_74#_M1010_g N_VGND_c_2543_n 0.00485498f $X=16.27 $Y=0.79 $X2=0
+ $Y2=0
cc_1244 N_A_2067_74#_M1038_g N_VGND_c_2550_n 0.00826076f $X=13.72 $Y=0.58 $X2=0
+ $Y2=0
cc_1245 N_A_2067_74#_M1022_g N_VGND_c_2550_n 0.00894397f $X=14.78 $Y=0.74 $X2=0
+ $Y2=0
cc_1246 N_A_2067_74#_M1025_g N_VGND_c_2550_n 0.00624688f $X=15.23 $Y=0.74 $X2=0
+ $Y2=0
cc_1247 N_A_2067_74#_M1010_g N_VGND_c_2550_n 0.00514438f $X=16.27 $Y=0.79 $X2=0
+ $Y2=0
cc_1248 N_A_2067_74#_c_1762_n N_VGND_c_2550_n 0.00674927f $X=11.38 $Y=0.945
+ $X2=0 $Y2=0
cc_1249 N_A_2067_74#_c_1841_n N_VGND_c_2550_n 0.0292546f $X=12.22 $Y=0.565 $X2=0
+ $Y2=0
cc_1250 N_A_2067_74#_c_1763_n N_VGND_c_2550_n 0.00599714f $X=11.55 $Y=0.565
+ $X2=0 $Y2=0
cc_1251 N_A_2067_74#_c_1762_n N_A_1794_74#_M1037_d 0.00457257f $X=11.38 $Y=0.945
+ $X2=0 $Y2=0
cc_1252 N_A_2067_74#_c_1766_n N_A_1794_74#_c_2705_n 0.00184691f $X=10.545
+ $Y=0.81 $X2=0 $Y2=0
cc_1253 N_A_2067_74#_M1032_s N_A_1794_74#_c_2707_n 0.00250873f $X=10.335 $Y=0.37
+ $X2=0 $Y2=0
cc_1254 N_A_2067_74#_c_1762_n N_A_1794_74#_c_2707_n 0.00337267f $X=11.38
+ $Y=0.945 $X2=0 $Y2=0
cc_1255 N_A_2067_74#_c_1766_n N_A_1794_74#_c_2707_n 0.0190143f $X=10.545 $Y=0.81
+ $X2=0 $Y2=0
cc_1256 N_A_2067_74#_c_1762_n N_A_1794_74#_c_2709_n 0.02441f $X=11.38 $Y=0.945
+ $X2=0 $Y2=0
cc_1257 N_A_2067_74#_c_1763_n N_A_1794_74#_c_2709_n 0.0229927f $X=11.55 $Y=0.565
+ $X2=0 $Y2=0
cc_1258 N_A_3177_368#_c_1991_n N_VPWR_c_2066_n 0.0701154f $X=16.03 $Y=1.985
+ $X2=0 $Y2=0
cc_1259 N_A_3177_368#_c_1995_n N_VPWR_c_2067_n 0.0090241f $X=16.805 $Y=1.765
+ $X2=0 $Y2=0
cc_1260 N_A_3177_368#_c_1991_n N_VPWR_c_2067_n 0.06488f $X=16.03 $Y=1.985 $X2=0
+ $Y2=0
cc_1261 N_A_3177_368#_c_1992_n N_VPWR_c_2067_n 0.0198206f $X=16.72 $Y=1.465
+ $X2=0 $Y2=0
cc_1262 N_A_3177_368#_c_1994_n N_VPWR_c_2067_n 0.00251384f $X=17.255 $Y=1.532
+ $X2=0 $Y2=0
cc_1263 N_A_3177_368#_c_1996_n N_VPWR_c_2069_n 0.00954146f $X=17.255 $Y=1.765
+ $X2=0 $Y2=0
cc_1264 N_A_3177_368#_c_1991_n N_VPWR_c_2081_n 0.0097982f $X=16.03 $Y=1.985
+ $X2=0 $Y2=0
cc_1265 N_A_3177_368#_c_1995_n N_VPWR_c_2082_n 0.00445602f $X=16.805 $Y=1.765
+ $X2=0 $Y2=0
cc_1266 N_A_3177_368#_c_1996_n N_VPWR_c_2082_n 0.00411612f $X=17.255 $Y=1.765
+ $X2=0 $Y2=0
cc_1267 N_A_3177_368#_c_1995_n N_VPWR_c_2057_n 0.00862391f $X=16.805 $Y=1.765
+ $X2=0 $Y2=0
cc_1268 N_A_3177_368#_c_1996_n N_VPWR_c_2057_n 0.00751023f $X=17.255 $Y=1.765
+ $X2=0 $Y2=0
cc_1269 N_A_3177_368#_c_1991_n N_VPWR_c_2057_n 0.0111907f $X=16.03 $Y=1.985
+ $X2=0 $Y2=0
cc_1270 N_A_3177_368#_c_1990_n N_Q_N_c_2460_n 0.00502622f $X=16.055 $Y=0.615
+ $X2=0 $Y2=0
cc_1271 N_A_3177_368#_c_1993_n Q_N 0.00298092f $X=16.042 $Y=1.465 $X2=0 $Y2=0
cc_1272 N_A_3177_368#_c_1995_n N_Q_c_2490_n 0.0111243f $X=16.805 $Y=1.765 $X2=0
+ $Y2=0
cc_1273 N_A_3177_368#_c_1996_n N_Q_c_2490_n 0.0130738f $X=17.255 $Y=1.765 $X2=0
+ $Y2=0
cc_1274 N_A_3177_368#_c_1995_n N_Q_c_2491_n 0.00231486f $X=16.805 $Y=1.765 $X2=0
+ $Y2=0
cc_1275 N_A_3177_368#_c_1996_n N_Q_c_2491_n 0.00240464f $X=17.255 $Y=1.765 $X2=0
+ $Y2=0
cc_1276 N_A_3177_368#_c_1992_n N_Q_c_2491_n 0.00140951f $X=16.72 $Y=1.465 $X2=0
+ $Y2=0
cc_1277 N_A_3177_368#_c_1994_n N_Q_c_2491_n 0.00807114f $X=17.255 $Y=1.532 $X2=0
+ $Y2=0
cc_1278 N_A_3177_368#_M1023_g N_Q_c_2487_n 0.0025553f $X=16.835 $Y=0.74 $X2=0
+ $Y2=0
cc_1279 N_A_3177_368#_c_1996_n N_Q_c_2487_n 0.0030228f $X=17.255 $Y=1.765 $X2=0
+ $Y2=0
cc_1280 N_A_3177_368#_M1049_g N_Q_c_2487_n 0.00866774f $X=17.265 $Y=0.74 $X2=0
+ $Y2=0
cc_1281 N_A_3177_368#_c_1992_n N_Q_c_2487_n 0.0249855f $X=16.72 $Y=1.465 $X2=0
+ $Y2=0
cc_1282 N_A_3177_368#_c_1994_n N_Q_c_2487_n 0.0359592f $X=17.255 $Y=1.532 $X2=0
+ $Y2=0
cc_1283 N_A_3177_368#_M1023_g Q 0.00761048f $X=16.835 $Y=0.74 $X2=0 $Y2=0
cc_1284 N_A_3177_368#_M1049_g Q 0.0081896f $X=17.265 $Y=0.74 $X2=0 $Y2=0
cc_1285 N_A_3177_368#_M1023_g Q 0.0032018f $X=16.835 $Y=0.74 $X2=0 $Y2=0
cc_1286 N_A_3177_368#_M1049_g Q 0.00215589f $X=17.265 $Y=0.74 $X2=0 $Y2=0
cc_1287 N_A_3177_368#_c_1994_n Q 0.00244427f $X=17.255 $Y=1.532 $X2=0 $Y2=0
cc_1288 N_A_3177_368#_c_1990_n N_VGND_c_2525_n 0.048096f $X=16.055 $Y=0.615
+ $X2=0 $Y2=0
cc_1289 N_A_3177_368#_M1023_g N_VGND_c_2526_n 0.00501537f $X=16.835 $Y=0.74
+ $X2=0 $Y2=0
cc_1290 N_A_3177_368#_c_1990_n N_VGND_c_2526_n 0.0405787f $X=16.055 $Y=0.615
+ $X2=0 $Y2=0
cc_1291 N_A_3177_368#_c_1992_n N_VGND_c_2526_n 0.0213234f $X=16.72 $Y=1.465
+ $X2=0 $Y2=0
cc_1292 N_A_3177_368#_c_1994_n N_VGND_c_2526_n 0.00347105f $X=17.255 $Y=1.532
+ $X2=0 $Y2=0
cc_1293 N_A_3177_368#_M1049_g N_VGND_c_2528_n 0.00646793f $X=17.265 $Y=0.74
+ $X2=0 $Y2=0
cc_1294 N_A_3177_368#_c_1990_n N_VGND_c_2543_n 0.0111427f $X=16.055 $Y=0.615
+ $X2=0 $Y2=0
cc_1295 N_A_3177_368#_M1023_g N_VGND_c_2544_n 0.00434272f $X=16.835 $Y=0.74
+ $X2=0 $Y2=0
cc_1296 N_A_3177_368#_M1049_g N_VGND_c_2544_n 0.00422942f $X=17.265 $Y=0.74
+ $X2=0 $Y2=0
cc_1297 N_A_3177_368#_M1023_g N_VGND_c_2550_n 0.00825283f $X=16.835 $Y=0.74
+ $X2=0 $Y2=0
cc_1298 N_A_3177_368#_M1049_g N_VGND_c_2550_n 0.00787255f $X=17.265 $Y=0.74
+ $X2=0 $Y2=0
cc_1299 N_A_3177_368#_c_1990_n N_VGND_c_2550_n 0.0122012f $X=16.055 $Y=0.615
+ $X2=0 $Y2=0
cc_1300 N_VPWR_c_2057_n N_A_304_464#_c_2260_n 0.0157311f $X=17.52 $Y=3.33 $X2=0
+ $Y2=0
cc_1301 N_VPWR_M1030_d N_A_304_464#_c_2262_n 0.00308424f $X=2.51 $Y=2.32 $X2=0
+ $Y2=0
cc_1302 N_VPWR_M1026_d N_A_304_464#_c_2262_n 0.00346042f $X=3.54 $Y=1.84 $X2=0
+ $Y2=0
cc_1303 N_VPWR_c_2059_n N_A_304_464#_c_2262_n 0.0166684f $X=2.67 $Y=2.815 $X2=0
+ $Y2=0
cc_1304 N_VPWR_c_2086_n N_A_304_464#_c_2262_n 0.010424f $X=4.22 $Y=3.032 $X2=0
+ $Y2=0
cc_1305 N_VPWR_c_2057_n N_A_304_464#_c_2262_n 0.0236194f $X=17.52 $Y=3.33 $X2=0
+ $Y2=0
cc_1306 N_VPWR_M1026_d N_A_304_464#_c_2263_n 0.00888923f $X=3.54 $Y=1.84 $X2=0
+ $Y2=0
cc_1307 N_VPWR_c_2086_n N_A_304_464#_c_2263_n 0.0132442f $X=4.22 $Y=3.032 $X2=0
+ $Y2=0
cc_1308 N_VPWR_c_2058_n N_A_304_464#_c_2264_n 0.0201206f $X=0.8 $Y=2.475 $X2=0
+ $Y2=0
cc_1309 N_VPWR_c_2059_n N_A_304_464#_c_2264_n 0.0098731f $X=2.67 $Y=2.815 $X2=0
+ $Y2=0
cc_1310 N_VPWR_c_2079_n N_A_304_464#_c_2264_n 0.019885f $X=2.495 $Y=3.33 $X2=0
+ $Y2=0
cc_1311 N_VPWR_c_2057_n N_A_304_464#_c_2264_n 0.0164027f $X=17.52 $Y=3.33 $X2=0
+ $Y2=0
cc_1312 N_VPWR_M1030_d N_A_304_464#_c_2298_n 7.42828e-19 $X=2.51 $Y=2.32 $X2=0
+ $Y2=0
cc_1313 N_VPWR_c_2059_n N_A_304_464#_c_2298_n 0.00710415f $X=2.67 $Y=2.815 $X2=0
+ $Y2=0
cc_1314 N_VPWR_c_2057_n N_A_304_464#_c_2298_n 0.0014507f $X=17.52 $Y=3.33 $X2=0
+ $Y2=0
cc_1315 N_VPWR_M1026_d N_A_304_464#_c_2300_n 0.0119658f $X=3.54 $Y=1.84 $X2=0
+ $Y2=0
cc_1316 N_VPWR_c_2086_n N_A_304_464#_c_2300_n 0.0140504f $X=4.22 $Y=3.032 $X2=0
+ $Y2=0
cc_1317 N_VPWR_c_2057_n N_A_304_464#_c_2300_n 5.67209e-19 $X=17.52 $Y=3.33 $X2=0
+ $Y2=0
cc_1318 N_VPWR_M1002_s N_A_1789_424#_c_2379_n 0.00450964f $X=9.44 $Y=2.12 $X2=0
+ $Y2=0
cc_1319 N_VPWR_c_2063_n N_A_1789_424#_c_2379_n 0.0154669f $X=9.59 $Y=2.725 $X2=0
+ $Y2=0
cc_1320 N_VPWR_c_2063_n N_A_1789_424#_c_2382_n 0.0285387f $X=9.59 $Y=2.725 $X2=0
+ $Y2=0
cc_1321 N_VPWR_c_2072_n N_A_1789_424#_c_2374_n 0.0646297f $X=12.94 $Y=3.33 $X2=0
+ $Y2=0
cc_1322 N_VPWR_c_2057_n N_A_1789_424#_c_2374_n 0.0359025f $X=17.52 $Y=3.33 $X2=0
+ $Y2=0
cc_1323 N_VPWR_c_2063_n N_A_1789_424#_c_2375_n 0.012272f $X=9.59 $Y=2.725 $X2=0
+ $Y2=0
cc_1324 N_VPWR_c_2072_n N_A_1789_424#_c_2375_n 0.017869f $X=12.94 $Y=3.33 $X2=0
+ $Y2=0
cc_1325 N_VPWR_c_2057_n N_A_1789_424#_c_2375_n 0.00965079f $X=17.52 $Y=3.33
+ $X2=0 $Y2=0
cc_1326 N_VPWR_c_2062_n N_A_1789_424#_c_2377_n 0.0364847f $X=8.5 $Y=2.57 $X2=0
+ $Y2=0
cc_1327 N_VPWR_c_2063_n N_A_1789_424#_c_2377_n 0.0191298f $X=9.59 $Y=2.725 $X2=0
+ $Y2=0
cc_1328 N_VPWR_c_2070_n N_A_1789_424#_c_2377_n 0.0146357f $X=9.425 $Y=3.33 $X2=0
+ $Y2=0
cc_1329 N_VPWR_c_2057_n N_A_1789_424#_c_2377_n 0.0121141f $X=17.52 $Y=3.33 $X2=0
+ $Y2=0
cc_1330 N_VPWR_c_2064_n N_A_2277_455#_c_2428_n 0.0119055f $X=13.025 $Y=2.75
+ $X2=0 $Y2=0
cc_1331 N_VPWR_c_2072_n N_A_2277_455#_c_2428_n 0.0653329f $X=12.94 $Y=3.33 $X2=0
+ $Y2=0
cc_1332 N_VPWR_c_2057_n N_A_2277_455#_c_2428_n 0.0388334f $X=17.52 $Y=3.33 $X2=0
+ $Y2=0
cc_1333 N_VPWR_c_2072_n N_A_2277_455#_c_2429_n 0.0162012f $X=12.94 $Y=3.33 $X2=0
+ $Y2=0
cc_1334 N_VPWR_c_2057_n N_A_2277_455#_c_2429_n 0.00879606f $X=17.52 $Y=3.33
+ $X2=0 $Y2=0
cc_1335 N_VPWR_c_2064_n N_A_2277_455#_c_2430_n 0.0237693f $X=13.025 $Y=2.75
+ $X2=0 $Y2=0
cc_1336 N_VPWR_c_2065_n N_Q_N_c_2459_n 0.075588f $X=14.57 $Y=1.985 $X2=0 $Y2=0
cc_1337 N_VPWR_c_2066_n N_Q_N_c_2459_n 0.0779559f $X=15.47 $Y=1.985 $X2=0 $Y2=0
cc_1338 N_VPWR_c_2076_n N_Q_N_c_2459_n 0.0112323f $X=15.305 $Y=3.33 $X2=0 $Y2=0
cc_1339 N_VPWR_c_2057_n N_Q_N_c_2459_n 0.00925249f $X=17.52 $Y=3.33 $X2=0 $Y2=0
cc_1340 N_VPWR_c_2082_n N_Q_c_2490_n 0.0158009f $X=17.395 $Y=3.33 $X2=0 $Y2=0
cc_1341 N_VPWR_c_2057_n N_Q_c_2490_n 0.0129424f $X=17.52 $Y=3.33 $X2=0 $Y2=0
cc_1342 N_VPWR_c_2067_n N_Q_c_2491_n 0.0783173f $X=16.58 $Y=1.985 $X2=0 $Y2=0
cc_1343 N_VPWR_c_2069_n N_Q_c_2491_n 0.0887573f $X=17.48 $Y=1.985 $X2=0 $Y2=0
cc_1344 N_A_304_464#_c_2260_n A_418_464# 0.00316297f $X=2.465 $Y=2.395 $X2=-0.19
+ $Y2=-0.245
cc_1345 N_A_304_464#_c_2257_n N_VGND_c_2518_n 0.00316404f $X=2.55 $Y=2.31 $X2=0
+ $Y2=0
cc_1346 N_A_304_464#_c_2279_n N_VGND_c_2518_n 0.0172749f $X=2.155 $Y=0.565 $X2=0
+ $Y2=0
cc_1347 N_A_304_464#_c_2279_n N_VGND_c_2529_n 0.0178113f $X=2.155 $Y=0.565 $X2=0
+ $Y2=0
cc_1348 N_A_304_464#_c_2279_n N_VGND_c_2550_n 0.0216127f $X=2.155 $Y=0.565 $X2=0
+ $Y2=0
cc_1349 N_A_304_464#_c_2257_n A_495_74# 5.40786e-19 $X=2.55 $Y=2.31 $X2=-0.19
+ $Y2=-0.245
cc_1350 N_A_304_464#_c_2279_n A_495_74# 0.00326443f $X=2.155 $Y=0.565 $X2=-0.19
+ $Y2=-0.245
cc_1351 N_A_1789_424#_c_2376_n N_A_2277_455#_c_2427_n 0.0302976f $X=10.94
+ $Y=2.465 $X2=0 $Y2=0
cc_1352 N_A_1789_424#_c_2374_n N_A_2277_455#_c_2429_n 0.0104058f $X=10.775
+ $Y=2.99 $X2=0 $Y2=0
cc_1353 N_A_1789_424#_c_2376_n N_A_2277_455#_c_2429_n 0.0012809f $X=10.94
+ $Y=2.465 $X2=0 $Y2=0
cc_1354 N_Q_N_c_2460_n N_VGND_c_2524_n 0.0176944f $X=15.015 $Y=0.515 $X2=0 $Y2=0
cc_1355 N_Q_N_c_2460_n N_VGND_c_2525_n 0.0600324f $X=15.015 $Y=0.515 $X2=0 $Y2=0
cc_1356 N_Q_N_c_2460_n N_VGND_c_2537_n 0.0168417f $X=15.015 $Y=0.515 $X2=0 $Y2=0
cc_1357 N_Q_N_c_2460_n N_VGND_c_2550_n 0.0137451f $X=15.015 $Y=0.515 $X2=0 $Y2=0
cc_1358 Q N_VGND_c_2526_n 0.0295042f $X=16.955 $Y=0.47 $X2=0 $Y2=0
cc_1359 Q N_VGND_c_2528_n 0.0308798f $X=16.955 $Y=0.47 $X2=0 $Y2=0
cc_1360 Q N_VGND_c_2544_n 0.0149085f $X=16.955 $Y=0.47 $X2=0 $Y2=0
cc_1361 Q N_VGND_c_2550_n 0.0122037f $X=16.955 $Y=0.47 $X2=0 $Y2=0
cc_1362 N_VGND_c_2521_n N_A_1794_74#_c_2704_n 0.0117303f $X=8.365 $Y=0.515 $X2=0
+ $Y2=0
cc_1363 N_VGND_c_2522_n N_A_1794_74#_c_2704_n 0.0189563f $X=9.615 $Y=0.59 $X2=0
+ $Y2=0
cc_1364 N_VGND_c_2531_n N_A_1794_74#_c_2704_n 0.011066f $X=9.45 $Y=0 $X2=0 $Y2=0
cc_1365 N_VGND_c_2550_n N_A_1794_74#_c_2704_n 0.00915947f $X=17.52 $Y=0 $X2=0
+ $Y2=0
cc_1366 N_VGND_M1001_d N_A_1794_74#_c_2705_n 0.00197722f $X=9.455 $Y=0.37 $X2=0
+ $Y2=0
cc_1367 N_VGND_c_2522_n N_A_1794_74#_c_2705_n 0.0172656f $X=9.615 $Y=0.59 $X2=0
+ $Y2=0
cc_1368 N_VGND_c_2533_n N_A_1794_74#_c_2707_n 0.0423335f $X=13.26 $Y=0 $X2=0
+ $Y2=0
cc_1369 N_VGND_c_2550_n N_A_1794_74#_c_2707_n 0.0239357f $X=17.52 $Y=0 $X2=0
+ $Y2=0
cc_1370 N_VGND_c_2522_n N_A_1794_74#_c_2708_n 0.0112234f $X=9.615 $Y=0.59 $X2=0
+ $Y2=0
cc_1371 N_VGND_c_2533_n N_A_1794_74#_c_2708_n 0.0178338f $X=13.26 $Y=0 $X2=0
+ $Y2=0
cc_1372 N_VGND_c_2550_n N_A_1794_74#_c_2708_n 0.00960503f $X=17.52 $Y=0 $X2=0
+ $Y2=0
cc_1373 N_VGND_c_2533_n N_A_1794_74#_c_2709_n 0.0227418f $X=13.26 $Y=0 $X2=0
+ $Y2=0
cc_1374 N_VGND_c_2550_n N_A_1794_74#_c_2709_n 0.0126077f $X=17.52 $Y=0 $X2=0
+ $Y2=0
