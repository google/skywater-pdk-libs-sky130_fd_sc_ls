# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_ls__a21oi_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005000 1.350000 3.350000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.180000 2.755000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.447000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.435000 0.435000 1.780000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.739300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 0.350000 0.860000 0.750000 ;
        RECT 0.605000 0.750000 3.180000 0.920000 ;
        RECT 0.605000 0.920000 0.860000 1.550000 ;
        RECT 0.605000 1.550000 1.395000 1.780000 ;
        RECT 1.065000 1.780000 1.395000 2.735000 ;
        RECT 2.930000 0.920000 3.180000 1.130000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.100000  0.085000 0.430000 1.130000 ;
      RECT 0.615000  1.950000 0.895000 2.905000 ;
      RECT 0.615000  2.905000 1.845000 3.075000 ;
      RECT 1.360000  1.090000 1.775000 1.260000 ;
      RECT 1.565000  1.260000 1.775000 1.950000 ;
      RECT 1.565000  1.950000 3.690000 2.120000 ;
      RECT 1.565000  2.290000 3.705000 2.460000 ;
      RECT 1.565000  2.460000 1.845000 2.905000 ;
      RECT 2.000000  0.085000 2.330000 0.580000 ;
      RECT 2.045000  2.630000 2.305000 3.245000 ;
      RECT 2.475000  2.460000 2.805000 2.980000 ;
      RECT 2.500000  0.330000 3.690000 0.580000 ;
      RECT 3.005000  2.630000 3.175000 3.245000 ;
      RECT 3.360000  0.580000 3.690000 1.130000 ;
      RECT 3.375000  2.460000 3.705000 2.980000 ;
      RECT 3.520000  1.130000 3.690000 1.950000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_ls__a21oi_2
END LIBRARY
