* NGSPICE file created from sky130_fd_sc_ls__nor2_2.ext - technology: sky130A

.subckt sky130_fd_sc_ls__nor2_2 A B VGND VNB VPB VPWR Y
M1000 a_35_368# A VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=9.968e+11p pd=8.5e+06u as=3.36e+11p ps=2.84e+06u
M1001 Y B VGND VNB nshort w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=5.254e+11p ps=4.38e+06u
M1002 VGND A Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 Y B a_35_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=0p ps=0u
M1004 a_35_368# B Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR A a_35_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

