* File: sky130_fd_sc_ls__a2111oi_2.spice
* Created: Fri Aug 28 12:48:27 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__a2111oi_2.pex.spice"
.subckt sky130_fd_sc_ls__a2111oi_2  VNB VPB D1 C1 B1 A1 A2 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A2	A2
* A1	A1
* B1	B1
* C1	C1
* D1	D1
* VPB	VPB
* VNB	VNB
MM1009 N_Y_M1009_d N_D1_M1009_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1443 AS=0.2109 PD=1.13 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.3 A=0.111 P=1.78 MULT=1
MM1000 N_VGND_M1000_d N_C1_M1000_g N_Y_M1009_d VNB NSHORT L=0.15 W=0.74
+ AD=0.1443 AS=0.1443 PD=1.13 PS=1.13 NRD=5.664 NRS=6.48 M=1 R=4.93333
+ SA=75000.7 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1011 N_Y_M1011_d N_B1_M1011_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.74
+ AD=0.1961 AS=0.1443 PD=2.01 PS=1.13 NRD=0 NRS=12.156 M=1 R=4.93333 SA=75001.3
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1001 N_A_722_74#_M1001_d N_A1_M1001_g N_Y_M1001_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1961 AS=0.1036 PD=2.01 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.5 A=0.111 P=1.78 MULT=1
MM1014 N_A_722_74#_M1014_d N_A1_M1014_g N_Y_M1001_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1007 N_A_722_74#_M1014_d N_A2_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1073 PD=1.02 PS=1.03 NRD=0 NRS=0.804 M=1 R=4.93333 SA=75001.1
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1013 N_A_722_74#_M1013_d N_A2_M1013_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1961 AS=0.1073 PD=2.01 PS=1.03 NRD=0 NRS=0.804 M=1 R=4.93333 SA=75001.5
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1002 N_A_69_368#_M1002_d N_D1_M1002_g N_Y_M1002_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.308 AS=0.168 PD=2.79 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75001.5 A=0.168 P=2.54 MULT=1
MM1016 N_A_69_368#_M1016_d N_D1_M1016_g N_Y_M1002_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.6 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1004 N_A_69_368#_M1016_d N_C1_M1004_g N_A_334_368#_M1004_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75000.6 A=0.168 P=2.54 MULT=1
MM1008 N_A_69_368#_M1008_d N_C1_M1008_g N_A_334_368#_M1004_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.308 AS=0.168 PD=2.79 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.5 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1006 N_A_334_368#_M1006_d N_B1_M1006_g N_A_533_368#_M1006_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.308 PD=1.42 PS=2.79 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75002.4 A=0.168 P=2.54 MULT=1
MM1010 N_A_334_368#_M1006_d N_B1_M1010_g N_A_533_368#_M1010_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.6 SB=75002 A=0.168 P=2.54 MULT=1
MM1012 N_VPWR_M1012_d N_A1_M1012_g N_A_533_368#_M1010_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75001.5 A=0.168 P=2.54 MULT=1
MM1015 N_VPWR_M1012_d N_A1_M1015_g N_A_533_368#_M1015_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.5 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1003 N_VPWR_M1003_d N_A2_M1003_g N_A_533_368#_M1015_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002 SB=75000.6 A=0.168 P=2.54 MULT=1
MM1005 N_VPWR_M1003_d N_A2_M1005_g N_A_533_368#_M1005_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.308 PD=1.42 PS=2.79 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.4 SB=75000.2 A=0.168 P=2.54 MULT=1
DX17_noxref VNB VPB NWDIODE A=11.4204 P=16
*
.include "sky130_fd_sc_ls__a2111oi_2.pxi.spice"
*
.ends
*
*
