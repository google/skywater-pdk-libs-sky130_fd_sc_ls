# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_ls__a41oi_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.925000 1.300000 3.255000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.195000 1.350000 2.755000 1.780000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 1.350000 1.955000 1.780000 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005000 1.350000 1.335000 1.780000 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.300000 0.435000 1.780000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.752200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115000 0.350000 0.445000 0.960000 ;
        RECT 0.115000 0.960000 3.220000 1.130000 ;
        RECT 0.115000 1.950000 0.835000 2.120000 ;
        RECT 0.115000 2.120000 0.445000 2.980000 ;
        RECT 0.605000 1.130000 0.835000 1.950000 ;
        RECT 2.890000 0.350000 3.220000 0.960000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.615000  0.085000 1.260000 0.680000 ;
      RECT 0.615000  2.290000 1.275000 2.460000 ;
      RECT 0.615000  2.460000 0.945000 2.980000 ;
      RECT 1.105000  1.950000 3.245000 2.290000 ;
      RECT 1.115000  2.630000 1.785000 3.245000 ;
      RECT 1.445000  2.460000 1.785000 2.630000 ;
      RECT 2.405000  2.460000 2.745000 3.245000 ;
      RECT 2.915000  2.290000 3.245000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_ls__a41oi_1
END LIBRARY
