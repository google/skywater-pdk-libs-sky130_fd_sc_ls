* File: sky130_fd_sc_ls__decaphe_3.pxi.spice
* Created: Wed Sep  2 10:59:47 2020
* 
x_PM_SKY130_FD_SC_LS__DECAPHE_3%VGND N_VGND_M1000_s N_VGND_c_12_n N_VGND_M1001_g
+ VGND N_VGND_c_13_n N_VGND_c_14_n PM_SKY130_FD_SC_LS__DECAPHE_3%VGND
x_PM_SKY130_FD_SC_LS__DECAPHE_3%VPWR N_VPWR_M1001_s N_VPWR_c_21_n N_VPWR_M1000_g
+ N_VPWR_c_22_n N_VPWR_c_25_n VPWR N_VPWR_c_27_n VPWR
+ PM_SKY130_FD_SC_LS__DECAPHE_3%VPWR
cc_1 VNB N_VGND_c_12_n 0.0322953f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2.035
cc_2 VNB N_VGND_c_13_n 0.106456f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=0
cc_3 VNB N_VGND_c_14_n 0.134994f $X=-0.19 $Y=-0.245 $X2=0.26 $Y2=0.38
cc_4 VNB N_VPWR_c_21_n 0.101305f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2.035
cc_5 VNB N_VPWR_c_22_n 0.0217188f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB VPWR 0.0641695f $X=-0.19 $Y=-0.245 $X2=0.26 $Y2=0.38
cc_7 VPB N_VGND_c_12_n 0.0690098f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=2.035
cc_8 VPB N_VPWR_c_22_n 0.062346f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_9 VPB N_VPWR_c_25_n 0.0633443f $X=-0.19 $Y=1.66 $X2=0.45 $Y2=1.515
cc_10 VPB VPWR 0.0423667f $X=-0.19 $Y=1.66 $X2=0.26 $Y2=0.38
cc_11 VPB N_VPWR_c_27_n 0.0281861f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_12 N_VGND_c_12_n N_VPWR_c_21_n 0.0427369f $X=0.72 $Y=2.035 $X2=0 $Y2=0
cc_13 N_VGND_c_14_n N_VPWR_c_21_n 0.106544f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_14 N_VGND_c_12_n N_VPWR_c_22_n 0.0685154f $X=0.72 $Y=2.035 $X2=0 $Y2=0
cc_15 N_VGND_c_14_n N_VPWR_c_22_n 0.129659f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_16 N_VGND_c_12_n N_VPWR_c_25_n 0.0709167f $X=0.72 $Y=2.035 $X2=0 $Y2=0
