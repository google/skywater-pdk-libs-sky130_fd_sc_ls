* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
M1000 VGND B1_N a_62_94# VNB nshort w=640000u l=150000u
+  ad=6.474e+11p pd=6.21e+06u as=1.696e+11p ps=1.81e+06u
M1001 VPWR A1 a_241_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=9.694e+11p pd=8.27e+06u as=1.288e+12p ps=1.126e+07u
M1002 a_62_94# B1_N VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.75e+11p pd=2.55e+06u as=0p ps=0u
M1003 Y a_62_94# VGND VNB nshort w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=0p ps=0u
M1004 VGND A2 a_436_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=5.994e+11p ps=6.06e+06u
M1005 a_241_368# A2 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_241_368# A1 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND a_62_94# Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y A1 a_436_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR A2 a_241_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 Y a_62_94# a_241_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=0p ps=0u
M1011 a_436_74# A2 VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_436_74# A1 Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_241_368# a_62_94# Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
