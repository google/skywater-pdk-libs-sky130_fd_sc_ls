* File: sky130_fd_sc_ls__dfstp_4.pxi.spice
* Created: Wed Sep  2 11:01:56 2020
* 
x_PM_SKY130_FD_SC_LS__DFSTP_4%D N_D_c_270_n N_D_c_275_n N_D_M1035_g N_D_c_276_n
+ N_D_M1033_g D D N_D_c_272_n N_D_c_273_n N_D_c_278_n
+ PM_SKY130_FD_SC_LS__DFSTP_4%D
x_PM_SKY130_FD_SC_LS__DFSTP_4%CLK N_CLK_c_305_n N_CLK_M1037_g N_CLK_c_306_n
+ N_CLK_M1026_g CLK PM_SKY130_FD_SC_LS__DFSTP_4%CLK
x_PM_SKY130_FD_SC_LS__DFSTP_4%A_398_74# N_A_398_74#_M1022_d N_A_398_74#_M1034_d
+ N_A_398_74#_c_337_n N_A_398_74#_M1010_g N_A_398_74#_c_338_n
+ N_A_398_74#_M1017_g N_A_398_74#_M1003_g N_A_398_74#_c_357_n
+ N_A_398_74#_M1028_g N_A_398_74#_c_340_n N_A_398_74#_c_453_p
+ N_A_398_74#_c_341_n N_A_398_74#_c_342_n N_A_398_74#_c_358_n
+ N_A_398_74#_c_359_n N_A_398_74#_c_343_n N_A_398_74#_c_344_n
+ N_A_398_74#_c_345_n N_A_398_74#_c_363_n N_A_398_74#_c_364_n
+ N_A_398_74#_c_365_n N_A_398_74#_c_366_n N_A_398_74#_c_367_n
+ N_A_398_74#_c_368_n N_A_398_74#_c_369_n N_A_398_74#_c_370_n
+ N_A_398_74#_c_346_n N_A_398_74#_c_347_n N_A_398_74#_c_348_n
+ N_A_398_74#_c_349_n N_A_398_74#_c_372_n N_A_398_74#_c_350_n
+ N_A_398_74#_c_351_n N_A_398_74#_c_352_n N_A_398_74#_c_373_n
+ N_A_398_74#_c_353_n N_A_398_74#_c_354_n PM_SKY130_FD_SC_LS__DFSTP_4%A_398_74#
x_PM_SKY130_FD_SC_LS__DFSTP_4%A_767_402# N_A_767_402#_M1029_s
+ N_A_767_402#_M1000_d N_A_767_402#_c_604_n N_A_767_402#_M1011_g
+ N_A_767_402#_c_598_n N_A_767_402#_M1001_g N_A_767_402#_c_599_n
+ N_A_767_402#_c_600_n N_A_767_402#_c_601_n N_A_767_402#_c_606_n
+ N_A_767_402#_c_607_n N_A_767_402#_c_602_n N_A_767_402#_c_608_n
+ N_A_767_402#_c_603_n PM_SKY130_FD_SC_LS__DFSTP_4%A_767_402#
x_PM_SKY130_FD_SC_LS__DFSTP_4%A_612_74# N_A_612_74#_M1027_d N_A_612_74#_M1010_d
+ N_A_612_74#_c_684_n N_A_612_74#_c_699_n N_A_612_74#_M1000_g
+ N_A_612_74#_c_685_n N_A_612_74#_M1029_g N_A_612_74#_c_686_n
+ N_A_612_74#_M1014_g N_A_612_74#_M1031_g N_A_612_74#_c_688_n
+ N_A_612_74#_c_689_n N_A_612_74#_c_690_n N_A_612_74#_c_691_n
+ N_A_612_74#_c_701_n N_A_612_74#_c_692_n N_A_612_74#_c_693_n
+ N_A_612_74#_c_694_n N_A_612_74#_c_695_n N_A_612_74#_c_696_n
+ N_A_612_74#_c_697_n PM_SKY130_FD_SC_LS__DFSTP_4%A_612_74#
x_PM_SKY130_FD_SC_LS__DFSTP_4%SET_B N_SET_B_c_832_n N_SET_B_c_833_n
+ N_SET_B_M1007_g N_SET_B_M1020_g N_SET_B_c_822_n N_SET_B_M1005_g
+ N_SET_B_c_823_n N_SET_B_c_824_n N_SET_B_c_835_n N_SET_B_c_836_n
+ N_SET_B_M1032_g N_SET_B_c_825_n N_SET_B_c_826_n N_SET_B_c_827_n SET_B
+ N_SET_B_c_829_n N_SET_B_c_830_n N_SET_B_c_831_n
+ PM_SKY130_FD_SC_LS__DFSTP_4%SET_B
x_PM_SKY130_FD_SC_LS__DFSTP_4%A_225_74# N_A_225_74#_M1037_s N_A_225_74#_M1026_s
+ N_A_225_74#_M1022_g N_A_225_74#_c_959_n N_A_225_74#_M1034_g
+ N_A_225_74#_c_971_n N_A_225_74#_c_960_n N_A_225_74#_c_972_n
+ N_A_225_74#_c_973_n N_A_225_74#_M1027_g N_A_225_74#_c_974_n
+ N_A_225_74#_c_975_n N_A_225_74#_c_976_n N_A_225_74#_M1019_g
+ N_A_225_74#_c_977_n N_A_225_74#_M1013_g N_A_225_74#_c_962_n
+ N_A_225_74#_c_963_n N_A_225_74#_M1018_g N_A_225_74#_c_965_n
+ N_A_225_74#_c_966_n N_A_225_74#_c_983_n N_A_225_74#_c_967_n
+ N_A_225_74#_c_985_n N_A_225_74#_c_968_n N_A_225_74#_c_969_n
+ N_A_225_74#_c_987_n PM_SKY130_FD_SC_LS__DFSTP_4%A_225_74#
x_PM_SKY130_FD_SC_LS__DFSTP_4%A_1484_62# N_A_1484_62#_M1002_d
+ N_A_1484_62#_M1030_d N_A_1484_62#_M1004_g N_A_1484_62#_c_1144_n
+ N_A_1484_62#_c_1145_n N_A_1484_62#_M1024_g N_A_1484_62#_c_1138_n
+ N_A_1484_62#_c_1139_n N_A_1484_62#_c_1155_n N_A_1484_62#_c_1140_n
+ N_A_1484_62#_c_1141_n N_A_1484_62#_c_1146_n N_A_1484_62#_c_1142_n
+ N_A_1484_62#_c_1143_n PM_SKY130_FD_SC_LS__DFSTP_4%A_1484_62#
x_PM_SKY130_FD_SC_LS__DFSTP_4%A_1321_392# N_A_1321_392#_M1003_d
+ N_A_1321_392#_M1013_d N_A_1321_392#_M1032_d N_A_1321_392#_c_1227_n
+ N_A_1321_392#_M1002_g N_A_1321_392#_c_1239_n N_A_1321_392#_M1030_g
+ N_A_1321_392#_c_1229_n N_A_1321_392#_M1038_g N_A_1321_392#_c_1231_n
+ N_A_1321_392#_M1012_g N_A_1321_392#_c_1232_n N_A_1321_392#_c_1242_n
+ N_A_1321_392#_M1023_g N_A_1321_392#_c_1243_n N_A_1321_392#_c_1233_n
+ N_A_1321_392#_c_1244_n N_A_1321_392#_c_1245_n N_A_1321_392#_c_1246_n
+ N_A_1321_392#_c_1247_n N_A_1321_392#_c_1248_n N_A_1321_392#_c_1234_n
+ N_A_1321_392#_c_1235_n N_A_1321_392#_c_1236_n N_A_1321_392#_c_1237_n
+ N_A_1321_392#_c_1249_n N_A_1321_392#_c_1250_n
+ PM_SKY130_FD_SC_LS__DFSTP_4%A_1321_392#
x_PM_SKY130_FD_SC_LS__DFSTP_4%A_1940_74# N_A_1940_74#_M1038_s
+ N_A_1940_74#_M1012_d N_A_1940_74#_c_1393_n N_A_1940_74#_M1006_g
+ N_A_1940_74#_c_1394_n N_A_1940_74#_c_1395_n N_A_1940_74#_c_1396_n
+ N_A_1940_74#_M1009_g N_A_1940_74#_c_1405_n N_A_1940_74#_M1008_g
+ N_A_1940_74#_c_1406_n N_A_1940_74#_M1015_g N_A_1940_74#_c_1397_n
+ N_A_1940_74#_M1021_g N_A_1940_74#_c_1407_n N_A_1940_74#_M1016_g
+ N_A_1940_74#_c_1398_n N_A_1940_74#_M1036_g N_A_1940_74#_c_1409_n
+ N_A_1940_74#_M1025_g N_A_1940_74#_c_1400_n N_A_1940_74#_c_1401_n
+ N_A_1940_74#_c_1402_n N_A_1940_74#_c_1410_n N_A_1940_74#_c_1403_n
+ N_A_1940_74#_c_1404_n PM_SKY130_FD_SC_LS__DFSTP_4%A_1940_74#
x_PM_SKY130_FD_SC_LS__DFSTP_4%A_27_74# N_A_27_74#_M1035_s N_A_27_74#_M1027_s
+ N_A_27_74#_M1033_s N_A_27_74#_M1010_s N_A_27_74#_c_1507_n N_A_27_74#_c_1508_n
+ N_A_27_74#_c_1513_n N_A_27_74#_c_1514_n N_A_27_74#_c_1515_n
+ N_A_27_74#_c_1509_n N_A_27_74#_c_1510_n N_A_27_74#_c_1517_n
+ N_A_27_74#_c_1559_n N_A_27_74#_c_1511_n PM_SKY130_FD_SC_LS__DFSTP_4%A_27_74#
x_PM_SKY130_FD_SC_LS__DFSTP_4%VPWR N_VPWR_M1033_d N_VPWR_M1026_d N_VPWR_M1011_d
+ N_VPWR_M1007_d N_VPWR_M1024_d N_VPWR_M1030_s N_VPWR_M1012_s N_VPWR_M1023_s
+ N_VPWR_M1015_d N_VPWR_M1025_d N_VPWR_c_1577_n N_VPWR_c_1578_n N_VPWR_c_1579_n
+ N_VPWR_c_1580_n N_VPWR_c_1581_n N_VPWR_c_1582_n N_VPWR_c_1583_n
+ N_VPWR_c_1584_n N_VPWR_c_1585_n N_VPWR_c_1586_n N_VPWR_c_1587_n
+ N_VPWR_c_1588_n N_VPWR_c_1589_n N_VPWR_c_1590_n N_VPWR_c_1591_n VPWR
+ N_VPWR_c_1592_n N_VPWR_c_1593_n N_VPWR_c_1594_n N_VPWR_c_1595_n
+ N_VPWR_c_1596_n N_VPWR_c_1597_n N_VPWR_c_1598_n N_VPWR_c_1599_n
+ N_VPWR_c_1600_n N_VPWR_c_1601_n N_VPWR_c_1602_n N_VPWR_c_1603_n
+ N_VPWR_c_1604_n N_VPWR_c_1605_n N_VPWR_c_1606_n N_VPWR_c_1607_n
+ N_VPWR_c_1576_n PM_SKY130_FD_SC_LS__DFSTP_4%VPWR
x_PM_SKY130_FD_SC_LS__DFSTP_4%Q N_Q_M1006_d N_Q_M1021_d N_Q_M1008_s N_Q_M1016_s
+ N_Q_c_1758_n N_Q_c_1759_n N_Q_c_1760_n N_Q_c_1765_n N_Q_c_1766_n N_Q_c_1761_n
+ N_Q_c_1767_n N_Q_c_1762_n N_Q_c_1763_n Q Q Q N_Q_c_1770_n
+ PM_SKY130_FD_SC_LS__DFSTP_4%Q
x_PM_SKY130_FD_SC_LS__DFSTP_4%VGND N_VGND_M1035_d N_VGND_M1037_d N_VGND_M1001_d
+ N_VGND_M1020_d N_VGND_M1005_d N_VGND_M1038_d N_VGND_M1009_s N_VGND_M1036_s
+ N_VGND_c_1831_n N_VGND_c_1832_n N_VGND_c_1833_n N_VGND_c_1834_n
+ N_VGND_c_1835_n N_VGND_c_1836_n N_VGND_c_1837_n N_VGND_c_1838_n
+ N_VGND_c_1839_n N_VGND_c_1840_n N_VGND_c_1841_n VGND N_VGND_c_1842_n
+ N_VGND_c_1843_n N_VGND_c_1844_n N_VGND_c_1845_n N_VGND_c_1846_n
+ N_VGND_c_1847_n N_VGND_c_1848_n N_VGND_c_1849_n N_VGND_c_1850_n
+ N_VGND_c_1851_n N_VGND_c_1852_n N_VGND_c_1853_n N_VGND_c_1854_n
+ PM_SKY130_FD_SC_LS__DFSTP_4%VGND
cc_1 VNB N_D_c_270_n 0.0447809f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.795
cc_2 VNB N_D_M1035_g 0.0283644f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.58
cc_3 VNB N_D_c_272_n 0.025337f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.145
cc_4 VNB N_D_c_273_n 0.00250659f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.145
cc_5 VNB N_CLK_c_305_n 0.0199457f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.175
cc_6 VNB N_CLK_c_306_n 0.0394284f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.355
cc_7 VNB CLK 0.00893055f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.58
cc_8 VNB N_A_398_74#_c_337_n 0.0158101f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.58
cc_9 VNB N_A_398_74#_c_338_n 0.0227081f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.73
cc_10 VNB N_A_398_74#_M1017_g 0.0525559f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_398_74#_c_340_n 0.00169421f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.145
cc_12 VNB N_A_398_74#_c_341_n 0.0153888f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.825
cc_13 VNB N_A_398_74#_c_342_n 0.00264685f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_398_74#_c_343_n 0.00190286f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_398_74#_c_344_n 0.00125833f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_398_74#_c_345_n 0.0174283f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_398_74#_c_346_n 0.00185717f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_398_74#_c_347_n 0.00920071f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_398_74#_c_348_n 0.00225196f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_398_74#_c_349_n 0.00683192f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_398_74#_c_350_n 0.00505342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_398_74#_c_351_n 0.03212f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_398_74#_c_352_n 0.00183894f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_398_74#_c_353_n 0.0136527f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_398_74#_c_354_n 0.0192244f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_767_402#_c_598_n 0.0191692f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.73
cc_27 VNB N_A_767_402#_c_599_n 0.0117603f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_28 VNB N_A_767_402#_c_600_n 0.00887451f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_767_402#_c_601_n 0.0253986f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.145
cc_30 VNB N_A_767_402#_c_602_n 0.0141708f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_767_402#_c_603_n 0.0359736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_612_74#_c_684_n 0.0126793f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_612_74#_c_685_n 0.0192259f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_34 VNB N_A_612_74#_c_686_n 0.0341009f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_612_74#_M1031_g 0.0248687f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.825
cc_36 VNB N_A_612_74#_c_688_n 0.00472968f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.145
cc_37 VNB N_A_612_74#_c_689_n 0.0145886f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.665
cc_38 VNB N_A_612_74#_c_690_n 0.00935088f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.825
cc_39 VNB N_A_612_74#_c_691_n 0.0176834f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_612_74#_c_692_n 0.00276658f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_612_74#_c_693_n 0.00220525f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_612_74#_c_694_n 0.00959991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_612_74#_c_695_n 0.00438751f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_612_74#_c_696_n 0.00189138f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_612_74#_c_697_n 0.0434133f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_SET_B_M1020_g 0.0426396f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_SET_B_c_822_n 0.0162437f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.73
cc_48 VNB N_SET_B_c_823_n 0.0682954f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_49 VNB N_SET_B_c_824_n 0.0198191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_SET_B_c_825_n 0.00103492f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.825
cc_51 VNB N_SET_B_c_826_n 0.0123954f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.825
cc_52 VNB N_SET_B_c_827_n 0.00109498f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.825
cc_53 VNB SET_B 0.00124466f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_SET_B_c_829_n 0.00324757f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_SET_B_c_830_n 0.00628098f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_SET_B_c_831_n 0.00233764f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_225_74#_M1022_g 0.0251862f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.445
cc_58 VNB N_A_225_74#_c_959_n 0.0124352f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.73
cc_59 VNB N_A_225_74#_c_960_n 0.0336376f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.145
cc_60 VNB N_A_225_74#_M1027_g 0.0294306f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.825
cc_61 VNB N_A_225_74#_c_962_n 0.0103413f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_225_74#_c_963_n 8.10901e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_225_74#_M1018_g 0.0515873f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_225_74#_c_965_n 0.0269886f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_225_74#_c_966_n 0.0195076f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_225_74#_c_967_n 0.0115791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_225_74#_c_968_n 0.00374876f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_225_74#_c_969_n 0.013166f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_1484_62#_M1004_g 0.0336842f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.445
cc_70 VNB N_A_1484_62#_c_1138_n 0.00351864f $X=-0.19 $Y=-0.245 $X2=0.64
+ $Y2=1.145
cc_71 VNB N_A_1484_62#_c_1139_n 0.0138251f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.825
cc_72 VNB N_A_1484_62#_c_1140_n 0.00682312f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_1484_62#_c_1141_n 0.00634625f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_1484_62#_c_1142_n 0.00805698f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_1484_62#_c_1143_n 0.0430611f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_1321_392#_c_1227_n 0.00412849f $X=-0.19 $Y=-0.245 $X2=0.505
+ $Y2=2.73
cc_77 VNB N_A_1321_392#_M1002_g 0.0507006f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_1321_392#_c_1229_n 0.0753249f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.98
cc_79 VNB N_A_1321_392#_M1038_g 0.0297718f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.99
cc_80 VNB N_A_1321_392#_c_1231_n 0.0136231f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_1321_392#_c_1232_n 0.0139059f $X=-0.19 $Y=-0.245 $X2=0.64
+ $Y2=1.665
cc_82 VNB N_A_1321_392#_c_1233_n 0.00512183f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_1321_392#_c_1234_n 0.00272086f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_1321_392#_c_1235_n 0.0240576f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_1321_392#_c_1236_n 2.14136e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_1321_392#_c_1237_n 0.00243428f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_1940_74#_c_1393_n 0.0181326f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.58
cc_88 VNB N_A_1940_74#_c_1394_n 0.0145071f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.73
cc_89 VNB N_A_1940_74#_c_1395_n 0.00747839f $X=-0.19 $Y=-0.245 $X2=0.505
+ $Y2=2.73
cc_90 VNB N_A_1940_74#_c_1396_n 0.0198904f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_91 VNB N_A_1940_74#_c_1397_n 0.0203684f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.825
cc_92 VNB N_A_1940_74#_c_1398_n 0.124232f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_1940_74#_M1036_g 0.0243152f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_1940_74#_c_1400_n 0.0146895f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_1940_74#_c_1401_n 0.00151156f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_1940_74#_c_1402_n 4.11739e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_1940_74#_c_1403_n 0.00463811f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_A_1940_74#_c_1404_n 0.00402022f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_A_27_74#_c_1507_n 0.0146704f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_A_27_74#_c_1508_n 0.040185f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.145
cc_101 VNB N_A_27_74#_c_1509_n 0.00677877f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.665
cc_102 VNB N_A_27_74#_c_1510_n 0.00791533f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_A_27_74#_c_1511_n 0.0065301f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_VPWR_c_1576_n 0.541827f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_Q_c_1758_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_Q_c_1759_n 0.00542399f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.145
cc_107 VNB N_Q_c_1760_n 0.00228436f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.145
cc_108 VNB N_Q_c_1761_n 0.00280896f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_Q_c_1762_n 0.00893228f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_Q_c_1763_n 0.00372816f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB Q 0.0268803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_1831_n 0.00766994f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_1832_n 0.0223817f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_1833_n 0.00555881f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_VGND_c_1834_n 0.0166819f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_VGND_c_1835_n 0.0172166f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_VGND_c_1836_n 0.00819684f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_VGND_c_1837_n 0.0118832f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_VGND_c_1838_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_VGND_c_1839_n 0.0297496f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_VGND_c_1840_n 0.0376041f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_VGND_c_1841_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB N_VGND_c_1842_n 0.0173909f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_VGND_c_1843_n 0.0561972f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_1844_n 0.0341238f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_1845_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_VGND_c_1846_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_1847_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_1848_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_1849_n 0.00738258f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_1850_n 0.0511502f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_VGND_c_1851_n 0.0397556f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_VGND_c_1852_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_VGND_c_1853_n 0.0127911f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_VGND_c_1854_n 0.714439f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VPB N_D_c_270_n 0.0126533f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.795
cc_137 VPB N_D_c_275_n 0.0292481f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.355
cc_138 VPB N_D_c_276_n 0.0298764f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.445
cc_139 VPB N_D_c_273_n 0.00226531f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.145
cc_140 VPB N_D_c_278_n 0.0244664f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.825
cc_141 VPB N_CLK_c_306_n 0.0238122f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.355
cc_142 VPB N_A_398_74#_c_337_n 0.0598775f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.58
cc_143 VPB N_A_398_74#_c_338_n 0.0168071f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.73
cc_144 VPB N_A_398_74#_c_357_n 0.0655752f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=0.98
cc_145 VPB N_A_398_74#_c_358_n 0.0207282f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_146 VPB N_A_398_74#_c_359_n 0.00247115f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_147 VPB N_A_398_74#_c_343_n 0.00198249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_148 VPB N_A_398_74#_c_344_n 0.00593785f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_149 VPB N_A_398_74#_c_345_n 0.0189713f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_150 VPB N_A_398_74#_c_363_n 0.00277688f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_151 VPB N_A_398_74#_c_364_n 0.00885724f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_152 VPB N_A_398_74#_c_365_n 0.00435535f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_153 VPB N_A_398_74#_c_366_n 0.0169194f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_154 VPB N_A_398_74#_c_367_n 0.00322702f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_155 VPB N_A_398_74#_c_368_n 0.00244123f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_156 VPB N_A_398_74#_c_369_n 0.00795467f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_157 VPB N_A_398_74#_c_370_n 5.72606e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_158 VPB N_A_398_74#_c_346_n 0.00241745f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_159 VPB N_A_398_74#_c_372_n 0.00102708f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_160 VPB N_A_398_74#_c_373_n 8.45509e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_161 VPB N_A_398_74#_c_353_n 0.00771916f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_162 VPB N_A_767_402#_c_604_n 0.0862223f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.58
cc_163 VPB N_A_767_402#_c_601_n 0.0023708f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.145
cc_164 VPB N_A_767_402#_c_606_n 0.0132551f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.145
cc_165 VPB N_A_767_402#_c_607_n 0.00272022f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.99
cc_166 VPB N_A_767_402#_c_608_n 0.00600776f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_167 VPB N_A_612_74#_c_684_n 0.0246211f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_168 VPB N_A_612_74#_c_699_n 0.0196697f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.445
cc_169 VPB N_A_612_74#_c_686_n 0.022768f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_170 VPB N_A_612_74#_c_701_n 0.00408741f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_171 VPB N_A_612_74#_c_692_n 0.00657766f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_172 VPB N_SET_B_c_832_n 0.00995661f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.795
cc_173 VPB N_SET_B_c_833_n 0.0201009f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.99
cc_174 VPB N_SET_B_M1020_g 0.00239435f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_175 VPB N_SET_B_c_835_n 0.0328389f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.145
cc_176 VPB N_SET_B_c_836_n 0.0242498f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.145
cc_177 VPB N_SET_B_c_825_n 0.0209448f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.825
cc_178 VPB N_SET_B_c_826_n 0.0186138f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.825
cc_179 VPB N_SET_B_c_827_n 0.00156093f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.825
cc_180 VPB SET_B 0.00132511f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_181 VPB N_SET_B_c_829_n 0.00641788f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_182 VPB N_SET_B_c_830_n 0.0350478f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_183 VPB N_SET_B_c_831_n 0.00327236f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_184 VPB N_A_225_74#_c_959_n 0.0218095f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.73
cc_185 VPB N_A_225_74#_c_971_n 0.0715755f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_186 VPB N_A_225_74#_c_972_n 0.0559655f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.145
cc_187 VPB N_A_225_74#_c_973_n 0.0123764f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=0.98
cc_188 VPB N_A_225_74#_c_974_n 0.00745492f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.145
cc_189 VPB N_A_225_74#_c_975_n 0.0131636f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_190 VPB N_A_225_74#_c_976_n 0.013997f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.295
cc_191 VPB N_A_225_74#_c_977_n 0.240375f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_192 VPB N_A_225_74#_M1013_g 0.00929298f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_193 VPB N_A_225_74#_c_962_n 0.0386327f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_194 VPB N_A_225_74#_c_963_n 0.0125099f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_195 VPB N_A_225_74#_c_965_n 5.35904e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_196 VPB N_A_225_74#_c_966_n 0.0110009f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_197 VPB N_A_225_74#_c_983_n 0.0089864f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_198 VPB N_A_225_74#_c_967_n 0.00180372f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_199 VPB N_A_225_74#_c_985_n 0.0047582f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_200 VPB N_A_225_74#_c_968_n 2.33575e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_201 VPB N_A_225_74#_c_987_n 0.0138824f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_202 VPB N_A_1484_62#_c_1144_n 0.0407199f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_203 VPB N_A_1484_62#_c_1145_n 0.0203789f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_204 VPB N_A_1484_62#_c_1146_n 0.00753471f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_205 VPB N_A_1484_62#_c_1142_n 0.0182499f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_206 VPB N_A_1321_392#_c_1227_n 0.0473246f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.73
cc_207 VPB N_A_1321_392#_c_1239_n 0.0577935f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.145
cc_208 VPB N_A_1321_392#_c_1231_n 0.0224903f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_209 VPB N_A_1321_392#_c_1232_n 0.011643f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.665
cc_210 VPB N_A_1321_392#_c_1242_n 0.0157753f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.825
cc_211 VPB N_A_1321_392#_c_1243_n 0.00277544f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_212 VPB N_A_1321_392#_c_1244_n 0.00471363f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_213 VPB N_A_1321_392#_c_1245_n 0.00993643f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_214 VPB N_A_1321_392#_c_1246_n 0.00812793f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_215 VPB N_A_1321_392#_c_1247_n 0.00854122f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_216 VPB N_A_1321_392#_c_1248_n 0.0136457f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_217 VPB N_A_1321_392#_c_1249_n 0.00300538f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_218 VPB N_A_1321_392#_c_1250_n 0.00509406f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_219 VPB N_A_1940_74#_c_1405_n 0.0163145f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_220 VPB N_A_1940_74#_c_1406_n 0.0149044f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.145
cc_221 VPB N_A_1940_74#_c_1407_n 0.0148817f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.145
cc_222 VPB N_A_1940_74#_c_1398_n 0.0266595f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_223 VPB N_A_1940_74#_c_1409_n 0.0171849f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_224 VPB N_A_1940_74#_c_1410_n 0.00394633f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_225 VPB N_A_27_74#_c_1508_n 0.0275147f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.145
cc_226 VPB N_A_27_74#_c_1513_n 0.0240891f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.825
cc_227 VPB N_A_27_74#_c_1514_n 0.0258928f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.99
cc_228 VPB N_A_27_74#_c_1515_n 0.0138477f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_229 VPB N_A_27_74#_c_1509_n 0.00245721f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.665
cc_230 VPB N_A_27_74#_c_1517_n 0.0109181f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.825
cc_231 VPB N_VPWR_c_1577_n 0.0139057f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_232 VPB N_VPWR_c_1578_n 0.00396467f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_233 VPB N_VPWR_c_1579_n 0.00600137f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_234 VPB N_VPWR_c_1580_n 0.00870193f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_235 VPB N_VPWR_c_1581_n 0.00805564f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_236 VPB N_VPWR_c_1582_n 0.0123473f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_237 VPB N_VPWR_c_1583_n 0.0348994f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_238 VPB N_VPWR_c_1584_n 0.0213734f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_239 VPB N_VPWR_c_1585_n 0.0211615f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_240 VPB N_VPWR_c_1586_n 0.0026822f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_241 VPB N_VPWR_c_1587_n 0.0116916f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_242 VPB N_VPWR_c_1588_n 0.0348185f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_243 VPB N_VPWR_c_1589_n 0.00184181f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_244 VPB N_VPWR_c_1590_n 0.036062f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_245 VPB N_VPWR_c_1591_n 0.0034365f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_246 VPB N_VPWR_c_1592_n 0.0182335f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_247 VPB N_VPWR_c_1593_n 0.0214173f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_248 VPB N_VPWR_c_1594_n 0.0487365f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_249 VPB N_VPWR_c_1595_n 0.0536763f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_250 VPB N_VPWR_c_1596_n 0.020445f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_251 VPB N_VPWR_c_1597_n 0.020445f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_252 VPB N_VPWR_c_1598_n 0.0173363f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_253 VPB N_VPWR_c_1599_n 0.0159778f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_254 VPB N_VPWR_c_1600_n 0.00628551f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_255 VPB N_VPWR_c_1601_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_256 VPB N_VPWR_c_1602_n 0.00223746f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_257 VPB N_VPWR_c_1603_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_258 VPB N_VPWR_c_1604_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_259 VPB N_VPWR_c_1605_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_260 VPB N_VPWR_c_1606_n 0.00535984f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_261 VPB N_VPWR_c_1607_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_262 VPB N_VPWR_c_1576_n 0.129069f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_263 VPB N_Q_c_1765_n 0.0016237f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=0.98
cc_264 VPB N_Q_c_1766_n 0.00243101f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.825
cc_265 VPB N_Q_c_1767_n 0.00233217f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_266 VPB Q 0.00853871f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_267 VPB Q 0.0175602f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_268 VPB N_Q_c_1770_n 0.00231053f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_269 N_D_c_272_n N_CLK_c_305_n 0.00232413f $X=0.64 $Y=1.145 $X2=-0.19
+ $Y2=-0.245
cc_270 N_D_c_270_n N_CLK_c_306_n 0.0100608f $X=0.61 $Y=1.795 $X2=0 $Y2=0
cc_271 N_D_c_270_n N_A_225_74#_c_967_n 0.0035771f $X=0.61 $Y=1.795 $X2=0 $Y2=0
cc_272 N_D_M1035_g N_A_225_74#_c_969_n 0.00621603f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_273 N_D_c_272_n N_A_225_74#_c_969_n 0.0035771f $X=0.64 $Y=1.145 $X2=0 $Y2=0
cc_274 N_D_c_273_n N_A_225_74#_c_969_n 0.0557245f $X=0.64 $Y=1.145 $X2=0 $Y2=0
cc_275 N_D_c_270_n N_A_225_74#_c_987_n 0.00300389f $X=0.61 $Y=1.795 $X2=0 $Y2=0
cc_276 N_D_c_275_n N_A_225_74#_c_987_n 0.00249516f $X=0.505 $Y=2.355 $X2=0 $Y2=0
cc_277 N_D_c_273_n N_A_225_74#_c_987_n 0.02241f $X=0.64 $Y=1.145 $X2=0 $Y2=0
cc_278 N_D_M1035_g N_A_27_74#_c_1507_n 0.00146243f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_279 N_D_M1035_g N_A_27_74#_c_1508_n 0.00600966f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_280 N_D_c_272_n N_A_27_74#_c_1508_n 0.0338681f $X=0.64 $Y=1.145 $X2=0 $Y2=0
cc_281 N_D_c_273_n N_A_27_74#_c_1508_n 0.0697394f $X=0.64 $Y=1.145 $X2=0 $Y2=0
cc_282 N_D_c_276_n N_A_27_74#_c_1513_n 0.00796498f $X=0.505 $Y=2.445 $X2=0 $Y2=0
cc_283 N_D_c_275_n N_A_27_74#_c_1514_n 0.0116201f $X=0.505 $Y=2.355 $X2=0 $Y2=0
cc_284 N_D_c_276_n N_A_27_74#_c_1514_n 0.00996787f $X=0.505 $Y=2.445 $X2=0 $Y2=0
cc_285 N_D_c_273_n N_A_27_74#_c_1514_n 0.019138f $X=0.64 $Y=1.145 $X2=0 $Y2=0
cc_286 N_D_c_278_n N_A_27_74#_c_1514_n 0.00134301f $X=0.64 $Y=1.825 $X2=0 $Y2=0
cc_287 N_D_c_276_n N_VPWR_c_1577_n 0.0122026f $X=0.505 $Y=2.445 $X2=0 $Y2=0
cc_288 N_D_c_276_n N_VPWR_c_1592_n 0.00505726f $X=0.505 $Y=2.445 $X2=0 $Y2=0
cc_289 N_D_c_276_n N_VPWR_c_1576_n 0.00526498f $X=0.505 $Y=2.445 $X2=0 $Y2=0
cc_290 N_D_M1035_g N_VGND_c_1831_n 0.0137856f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_291 N_D_c_272_n N_VGND_c_1831_n 0.00175174f $X=0.64 $Y=1.145 $X2=0 $Y2=0
cc_292 N_D_c_273_n N_VGND_c_1831_n 0.0220022f $X=0.64 $Y=1.145 $X2=0 $Y2=0
cc_293 N_D_M1035_g N_VGND_c_1842_n 0.00383152f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_294 N_D_M1035_g N_VGND_c_1854_n 0.00761198f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_295 N_CLK_c_305_n N_A_225_74#_M1022_g 0.0131399f $X=1.485 $Y=1.22 $X2=0 $Y2=0
cc_296 N_CLK_c_306_n N_A_225_74#_M1022_g 0.0206752f $X=1.515 $Y=1.765 $X2=0
+ $Y2=0
cc_297 CLK N_A_225_74#_M1022_g 0.00400177f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_298 N_CLK_c_306_n N_A_225_74#_c_959_n 0.0493156f $X=1.515 $Y=1.765 $X2=0
+ $Y2=0
cc_299 N_CLK_c_305_n N_A_225_74#_c_967_n 0.00330079f $X=1.485 $Y=1.22 $X2=0
+ $Y2=0
cc_300 N_CLK_c_306_n N_A_225_74#_c_967_n 0.00653993f $X=1.515 $Y=1.765 $X2=0
+ $Y2=0
cc_301 CLK N_A_225_74#_c_967_n 0.0286813f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_302 N_CLK_c_306_n N_A_225_74#_c_985_n 0.00976072f $X=1.515 $Y=1.765 $X2=0
+ $Y2=0
cc_303 N_CLK_c_306_n N_A_225_74#_c_968_n 0.00106267f $X=1.515 $Y=1.765 $X2=0
+ $Y2=0
cc_304 CLK N_A_225_74#_c_968_n 0.0162505f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_305 N_CLK_c_305_n N_A_225_74#_c_969_n 0.00811931f $X=1.485 $Y=1.22 $X2=0
+ $Y2=0
cc_306 N_CLK_c_306_n N_A_225_74#_c_969_n 0.00114664f $X=1.515 $Y=1.765 $X2=0
+ $Y2=0
cc_307 CLK N_A_225_74#_c_969_n 0.00763035f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_308 N_CLK_c_306_n N_A_225_74#_c_987_n 0.00986362f $X=1.515 $Y=1.765 $X2=0
+ $Y2=0
cc_309 CLK N_A_225_74#_c_987_n 0.0353752f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_310 N_CLK_c_306_n N_A_27_74#_c_1514_n 0.016333f $X=1.515 $Y=1.765 $X2=0 $Y2=0
cc_311 CLK N_A_27_74#_c_1509_n 0.00460396f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_312 N_CLK_c_306_n N_VPWR_c_1577_n 0.0127382f $X=1.515 $Y=1.765 $X2=0 $Y2=0
cc_313 N_CLK_c_306_n N_VPWR_c_1578_n 0.0239849f $X=1.515 $Y=1.765 $X2=0 $Y2=0
cc_314 N_CLK_c_306_n N_VPWR_c_1593_n 0.00413917f $X=1.515 $Y=1.765 $X2=0 $Y2=0
cc_315 N_CLK_c_306_n N_VPWR_c_1576_n 0.00822528f $X=1.515 $Y=1.765 $X2=0 $Y2=0
cc_316 N_CLK_c_305_n N_VGND_c_1831_n 0.00280144f $X=1.485 $Y=1.22 $X2=0 $Y2=0
cc_317 N_CLK_c_305_n N_VGND_c_1832_n 0.00434054f $X=1.485 $Y=1.22 $X2=0 $Y2=0
cc_318 N_CLK_c_305_n N_VGND_c_1833_n 0.0027655f $X=1.485 $Y=1.22 $X2=0 $Y2=0
cc_319 CLK N_VGND_c_1833_n 0.013855f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_320 N_CLK_c_305_n N_VGND_c_1854_n 0.0082522f $X=1.485 $Y=1.22 $X2=0 $Y2=0
cc_321 N_A_398_74#_c_337_n N_A_767_402#_c_604_n 0.00106832f $X=3.005 $Y=2.24
+ $X2=0 $Y2=0
cc_322 N_A_398_74#_c_344_n N_A_767_402#_c_604_n 0.00760718f $X=3.71 $Y=1.635
+ $X2=0 $Y2=0
cc_323 N_A_398_74#_c_345_n N_A_767_402#_c_604_n 0.0088185f $X=3.71 $Y=1.635
+ $X2=0 $Y2=0
cc_324 N_A_398_74#_c_363_n N_A_767_402#_c_604_n 0.00256198f $X=3.71 $Y=2.905
+ $X2=0 $Y2=0
cc_325 N_A_398_74#_c_364_n N_A_767_402#_c_604_n 0.0325047f $X=4.515 $Y=2.25
+ $X2=0 $Y2=0
cc_326 N_A_398_74#_c_365_n N_A_767_402#_c_604_n 0.00359428f $X=4.6 $Y=2.905
+ $X2=0 $Y2=0
cc_327 N_A_398_74#_M1017_g N_A_767_402#_c_598_n 0.0422629f $X=3.585 $Y=0.58
+ $X2=0 $Y2=0
cc_328 N_A_398_74#_c_344_n N_A_767_402#_c_601_n 6.69553e-19 $X=3.71 $Y=1.635
+ $X2=0 $Y2=0
cc_329 N_A_398_74#_c_345_n N_A_767_402#_c_601_n 0.00851627f $X=3.71 $Y=1.635
+ $X2=0 $Y2=0
cc_330 N_A_398_74#_c_344_n N_A_767_402#_c_606_n 0.0123371f $X=3.71 $Y=1.635
+ $X2=0 $Y2=0
cc_331 N_A_398_74#_c_345_n N_A_767_402#_c_606_n 2.62742e-19 $X=3.71 $Y=1.635
+ $X2=0 $Y2=0
cc_332 N_A_398_74#_c_364_n N_A_767_402#_c_606_n 0.0444853f $X=4.515 $Y=2.25
+ $X2=0 $Y2=0
cc_333 N_A_398_74#_c_364_n N_A_767_402#_c_607_n 0.0104536f $X=4.515 $Y=2.25
+ $X2=0 $Y2=0
cc_334 N_A_398_74#_c_368_n N_A_767_402#_c_607_n 0.00133551f $X=5.425 $Y=2.905
+ $X2=0 $Y2=0
cc_335 N_A_398_74#_c_370_n N_A_767_402#_c_607_n 0.00848739f $X=5.51 $Y=2.18
+ $X2=0 $Y2=0
cc_336 N_A_398_74#_M1017_g N_A_767_402#_c_602_n 8.22539e-19 $X=3.585 $Y=0.58
+ $X2=0 $Y2=0
cc_337 N_A_398_74#_c_364_n N_A_767_402#_c_608_n 0.00325944f $X=4.515 $Y=2.25
+ $X2=0 $Y2=0
cc_338 N_A_398_74#_c_365_n N_A_767_402#_c_608_n 0.029467f $X=4.6 $Y=2.905 $X2=0
+ $Y2=0
cc_339 N_A_398_74#_c_366_n N_A_767_402#_c_608_n 0.0211624f $X=5.34 $Y=2.99 $X2=0
+ $Y2=0
cc_340 N_A_398_74#_c_368_n N_A_767_402#_c_608_n 0.0324793f $X=5.425 $Y=2.905
+ $X2=0 $Y2=0
cc_341 N_A_398_74#_M1017_g N_A_767_402#_c_603_n 0.00603499f $X=3.585 $Y=0.58
+ $X2=0 $Y2=0
cc_342 N_A_398_74#_c_364_n N_A_612_74#_c_699_n 0.00377878f $X=4.515 $Y=2.25
+ $X2=0 $Y2=0
cc_343 N_A_398_74#_c_365_n N_A_612_74#_c_699_n 0.0117078f $X=4.6 $Y=2.905 $X2=0
+ $Y2=0
cc_344 N_A_398_74#_c_366_n N_A_612_74#_c_699_n 0.0027223f $X=5.34 $Y=2.99 $X2=0
+ $Y2=0
cc_345 N_A_398_74#_c_368_n N_A_612_74#_c_699_n 6.03222e-19 $X=5.425 $Y=2.905
+ $X2=0 $Y2=0
cc_346 N_A_398_74#_c_368_n N_A_612_74#_c_686_n 0.00330096f $X=5.425 $Y=2.905
+ $X2=0 $Y2=0
cc_347 N_A_398_74#_c_369_n N_A_612_74#_c_686_n 0.0201389f $X=6.305 $Y=2.18 $X2=0
+ $Y2=0
cc_348 N_A_398_74#_c_346_n N_A_612_74#_c_686_n 0.00905037f $X=6.39 $Y=2.095
+ $X2=0 $Y2=0
cc_349 N_A_398_74#_c_350_n N_A_612_74#_c_686_n 0.00389788f $X=6.53 $Y=1.285
+ $X2=0 $Y2=0
cc_350 N_A_398_74#_c_351_n N_A_612_74#_c_686_n 0.0139138f $X=6.53 $Y=1.285 $X2=0
+ $Y2=0
cc_351 N_A_398_74#_c_348_n N_A_612_74#_M1031_g 0.00161751f $X=6.475 $Y=0.34
+ $X2=0 $Y2=0
cc_352 N_A_398_74#_c_351_n N_A_612_74#_M1031_g 0.00397266f $X=6.53 $Y=1.285
+ $X2=0 $Y2=0
cc_353 N_A_398_74#_c_352_n N_A_612_74#_M1031_g 0.00869284f $X=6.5 $Y=1.12 $X2=0
+ $Y2=0
cc_354 N_A_398_74#_c_354_n N_A_612_74#_M1031_g 0.0195997f $X=6.53 $Y=1.12 $X2=0
+ $Y2=0
cc_355 N_A_398_74#_M1017_g N_A_612_74#_c_688_n 0.0187196f $X=3.585 $Y=0.58 $X2=0
+ $Y2=0
cc_356 N_A_398_74#_c_341_n N_A_612_74#_c_688_n 0.00381334f $X=2.945 $Y=0.34
+ $X2=0 $Y2=0
cc_357 N_A_398_74#_c_349_n N_A_612_74#_c_688_n 0.0403355f $X=2.95 $Y=1.455 $X2=0
+ $Y2=0
cc_358 N_A_398_74#_M1017_g N_A_612_74#_c_689_n 0.0142826f $X=3.585 $Y=0.58 $X2=0
+ $Y2=0
cc_359 N_A_398_74#_c_344_n N_A_612_74#_c_689_n 0.0132987f $X=3.71 $Y=1.635 $X2=0
+ $Y2=0
cc_360 N_A_398_74#_c_345_n N_A_612_74#_c_689_n 0.0039875f $X=3.71 $Y=1.635 $X2=0
+ $Y2=0
cc_361 N_A_398_74#_c_337_n N_A_612_74#_c_701_n 0.00240563f $X=3.005 $Y=2.24
+ $X2=0 $Y2=0
cc_362 N_A_398_74#_c_338_n N_A_612_74#_c_701_n 0.00503148f $X=3.51 $Y=1.635
+ $X2=0 $Y2=0
cc_363 N_A_398_74#_c_358_n N_A_612_74#_c_701_n 0.0225127f $X=3.625 $Y=2.99 $X2=0
+ $Y2=0
cc_364 N_A_398_74#_c_337_n N_A_612_74#_c_692_n 0.0086847f $X=3.005 $Y=2.24 $X2=0
+ $Y2=0
cc_365 N_A_398_74#_c_338_n N_A_612_74#_c_692_n 0.0222601f $X=3.51 $Y=1.635 $X2=0
+ $Y2=0
cc_366 N_A_398_74#_M1017_g N_A_612_74#_c_692_n 0.00425975f $X=3.585 $Y=0.58
+ $X2=0 $Y2=0
cc_367 N_A_398_74#_c_344_n N_A_612_74#_c_692_n 0.0498141f $X=3.71 $Y=1.635 $X2=0
+ $Y2=0
cc_368 N_A_398_74#_c_349_n N_A_612_74#_c_692_n 0.0606779f $X=2.95 $Y=1.455 $X2=0
+ $Y2=0
cc_369 N_A_398_74#_c_372_n N_A_612_74#_c_692_n 0.0129296f $X=3.71 $Y=2.25 $X2=0
+ $Y2=0
cc_370 N_A_398_74#_c_338_n N_A_612_74#_c_693_n 0.00242402f $X=3.51 $Y=1.635
+ $X2=0 $Y2=0
cc_371 N_A_398_74#_M1017_g N_A_612_74#_c_693_n 0.00427915f $X=3.585 $Y=0.58
+ $X2=0 $Y2=0
cc_372 N_A_398_74#_c_349_n N_A_612_74#_c_693_n 0.0143568f $X=2.95 $Y=1.455 $X2=0
+ $Y2=0
cc_373 N_A_398_74#_M1017_g N_A_612_74#_c_694_n 0.00178188f $X=3.585 $Y=0.58
+ $X2=0 $Y2=0
cc_374 N_A_398_74#_c_344_n N_A_612_74#_c_694_n 0.00715168f $X=3.71 $Y=1.635
+ $X2=0 $Y2=0
cc_375 N_A_398_74#_c_345_n N_A_612_74#_c_694_n 9.47085e-19 $X=3.71 $Y=1.635
+ $X2=0 $Y2=0
cc_376 N_A_398_74#_c_364_n N_A_612_74#_c_694_n 0.00485285f $X=4.515 $Y=2.25
+ $X2=0 $Y2=0
cc_377 N_A_398_74#_c_369_n N_A_612_74#_c_696_n 0.00289162f $X=6.305 $Y=2.18
+ $X2=0 $Y2=0
cc_378 N_A_398_74#_c_350_n N_A_612_74#_c_696_n 0.0230196f $X=6.53 $Y=1.285 $X2=0
+ $Y2=0
cc_379 N_A_398_74#_c_351_n N_A_612_74#_c_696_n 2.80493e-19 $X=6.53 $Y=1.285
+ $X2=0 $Y2=0
cc_380 N_A_398_74#_c_370_n N_SET_B_c_832_n 0.00276362f $X=5.51 $Y=2.18 $X2=0
+ $Y2=0
cc_381 N_A_398_74#_c_366_n N_SET_B_c_833_n 0.00294574f $X=5.34 $Y=2.99 $X2=0
+ $Y2=0
cc_382 N_A_398_74#_c_368_n N_SET_B_c_833_n 0.0157239f $X=5.425 $Y=2.905 $X2=0
+ $Y2=0
cc_383 N_A_398_74#_c_370_n N_SET_B_c_833_n 0.00435079f $X=5.51 $Y=2.18 $X2=0
+ $Y2=0
cc_384 N_A_398_74#_c_357_n N_SET_B_c_826_n 0.0010485f $X=7.325 $Y=2.465 $X2=0
+ $Y2=0
cc_385 N_A_398_74#_c_369_n N_SET_B_c_826_n 0.0191764f $X=6.305 $Y=2.18 $X2=0
+ $Y2=0
cc_386 N_A_398_74#_c_346_n N_SET_B_c_826_n 0.0222258f $X=6.39 $Y=2.095 $X2=0
+ $Y2=0
cc_387 N_A_398_74#_c_350_n N_SET_B_c_826_n 0.00959624f $X=6.53 $Y=1.285 $X2=0
+ $Y2=0
cc_388 N_A_398_74#_c_373_n N_SET_B_c_826_n 0.00572674f $X=7.21 $Y=2.185 $X2=0
+ $Y2=0
cc_389 N_A_398_74#_c_353_n N_SET_B_c_826_n 0.0208316f $X=7.21 $Y=2.02 $X2=0
+ $Y2=0
cc_390 N_A_398_74#_c_369_n N_SET_B_c_827_n 0.00190675f $X=6.305 $Y=2.18 $X2=0
+ $Y2=0
cc_391 N_A_398_74#_c_370_n N_SET_B_c_827_n 8.05363e-19 $X=5.51 $Y=2.18 $X2=0
+ $Y2=0
cc_392 N_A_398_74#_c_369_n N_SET_B_c_829_n 0.00913037f $X=6.305 $Y=2.18 $X2=0
+ $Y2=0
cc_393 N_A_398_74#_c_370_n N_SET_B_c_829_n 0.0133873f $X=5.51 $Y=2.18 $X2=0
+ $Y2=0
cc_394 N_A_398_74#_c_346_n N_SET_B_c_829_n 0.00814699f $X=6.39 $Y=2.095 $X2=0
+ $Y2=0
cc_395 N_A_398_74#_c_369_n N_SET_B_c_830_n 0.00156156f $X=6.305 $Y=2.18 $X2=0
+ $Y2=0
cc_396 N_A_398_74#_c_370_n N_SET_B_c_830_n 0.00317486f $X=5.51 $Y=2.18 $X2=0
+ $Y2=0
cc_397 N_A_398_74#_c_340_n N_A_225_74#_M1022_g 0.00164183f $X=2.13 $Y=0.515
+ $X2=0 $Y2=0
cc_398 N_A_398_74#_c_342_n N_A_225_74#_M1022_g 0.00266901f $X=2.215 $Y=0.34
+ $X2=0 $Y2=0
cc_399 N_A_398_74#_c_453_p N_A_225_74#_c_959_n 0.00503544f $X=2.19 $Y=2.575
+ $X2=0 $Y2=0
cc_400 N_A_398_74#_c_359_n N_A_225_74#_c_959_n 0.00163933f $X=2.275 $Y=2.99
+ $X2=0 $Y2=0
cc_401 N_A_398_74#_c_337_n N_A_225_74#_c_971_n 0.0172835f $X=3.005 $Y=2.24 $X2=0
+ $Y2=0
cc_402 N_A_398_74#_c_453_p N_A_225_74#_c_971_n 0.00606451f $X=2.19 $Y=2.575
+ $X2=0 $Y2=0
cc_403 N_A_398_74#_c_358_n N_A_225_74#_c_971_n 0.0102166f $X=3.625 $Y=2.99 $X2=0
+ $Y2=0
cc_404 N_A_398_74#_c_343_n N_A_225_74#_c_971_n 3.80136e-19 $X=2.95 $Y=1.62 $X2=0
+ $Y2=0
cc_405 N_A_398_74#_c_337_n N_A_225_74#_c_960_n 0.0147005f $X=3.005 $Y=2.24 $X2=0
+ $Y2=0
cc_406 N_A_398_74#_c_341_n N_A_225_74#_c_960_n 0.00237694f $X=2.945 $Y=0.34
+ $X2=0 $Y2=0
cc_407 N_A_398_74#_c_343_n N_A_225_74#_c_960_n 0.00105733f $X=2.95 $Y=1.62 $X2=0
+ $Y2=0
cc_408 N_A_398_74#_c_349_n N_A_225_74#_c_960_n 0.00695648f $X=2.95 $Y=1.455
+ $X2=0 $Y2=0
cc_409 N_A_398_74#_c_337_n N_A_225_74#_c_972_n 0.00882199f $X=3.005 $Y=2.24
+ $X2=0 $Y2=0
cc_410 N_A_398_74#_c_358_n N_A_225_74#_c_972_n 0.0133466f $X=3.625 $Y=2.99 $X2=0
+ $Y2=0
cc_411 N_A_398_74#_M1017_g N_A_225_74#_M1027_g 0.0179618f $X=3.585 $Y=0.58 $X2=0
+ $Y2=0
cc_412 N_A_398_74#_c_340_n N_A_225_74#_M1027_g 0.00395905f $X=2.13 $Y=0.515
+ $X2=0 $Y2=0
cc_413 N_A_398_74#_c_341_n N_A_225_74#_M1027_g 0.010044f $X=2.945 $Y=0.34 $X2=0
+ $Y2=0
cc_414 N_A_398_74#_c_349_n N_A_225_74#_M1027_g 0.0216123f $X=2.95 $Y=1.455 $X2=0
+ $Y2=0
cc_415 N_A_398_74#_c_337_n N_A_225_74#_c_974_n 0.00215978f $X=3.005 $Y=2.24
+ $X2=0 $Y2=0
cc_416 N_A_398_74#_c_363_n N_A_225_74#_c_974_n 0.00293397f $X=3.71 $Y=2.905
+ $X2=0 $Y2=0
cc_417 N_A_398_74#_c_358_n N_A_225_74#_c_975_n 0.0181345f $X=3.625 $Y=2.99 $X2=0
+ $Y2=0
cc_418 N_A_398_74#_c_337_n N_A_225_74#_c_976_n 0.012524f $X=3.005 $Y=2.24 $X2=0
+ $Y2=0
cc_419 N_A_398_74#_c_338_n N_A_225_74#_c_976_n 0.00662218f $X=3.51 $Y=1.635
+ $X2=0 $Y2=0
cc_420 N_A_398_74#_c_363_n N_A_225_74#_c_976_n 0.00344316f $X=3.71 $Y=2.905
+ $X2=0 $Y2=0
cc_421 N_A_398_74#_c_372_n N_A_225_74#_c_976_n 0.0011228f $X=3.71 $Y=2.25 $X2=0
+ $Y2=0
cc_422 N_A_398_74#_c_357_n N_A_225_74#_c_977_n 0.00133957f $X=7.325 $Y=2.465
+ $X2=0 $Y2=0
cc_423 N_A_398_74#_c_358_n N_A_225_74#_c_977_n 0.00488406f $X=3.625 $Y=2.99
+ $X2=0 $Y2=0
cc_424 N_A_398_74#_c_366_n N_A_225_74#_c_977_n 0.0145684f $X=5.34 $Y=2.99 $X2=0
+ $Y2=0
cc_425 N_A_398_74#_c_367_n N_A_225_74#_c_977_n 0.00420304f $X=4.685 $Y=2.99
+ $X2=0 $Y2=0
cc_426 N_A_398_74#_c_357_n N_A_225_74#_M1013_g 0.00240896f $X=7.325 $Y=2.465
+ $X2=0 $Y2=0
cc_427 N_A_398_74#_c_369_n N_A_225_74#_M1013_g 0.00520345f $X=6.305 $Y=2.18
+ $X2=0 $Y2=0
cc_428 N_A_398_74#_c_346_n N_A_225_74#_M1013_g 0.00414836f $X=6.39 $Y=2.095
+ $X2=0 $Y2=0
cc_429 N_A_398_74#_c_357_n N_A_225_74#_c_962_n 0.00901519f $X=7.325 $Y=2.465
+ $X2=0 $Y2=0
cc_430 N_A_398_74#_c_373_n N_A_225_74#_c_962_n 0.00103484f $X=7.21 $Y=2.185
+ $X2=0 $Y2=0
cc_431 N_A_398_74#_c_346_n N_A_225_74#_c_963_n 0.00568179f $X=6.39 $Y=2.095
+ $X2=0 $Y2=0
cc_432 N_A_398_74#_c_350_n N_A_225_74#_c_963_n 0.00124953f $X=6.53 $Y=1.285
+ $X2=0 $Y2=0
cc_433 N_A_398_74#_c_351_n N_A_225_74#_c_963_n 0.0172051f $X=6.53 $Y=1.285 $X2=0
+ $Y2=0
cc_434 N_A_398_74#_c_346_n N_A_225_74#_M1018_g 8.38958e-19 $X=6.39 $Y=2.095
+ $X2=0 $Y2=0
cc_435 N_A_398_74#_c_347_n N_A_225_74#_M1018_g 0.0127652f $X=7.205 $Y=0.34 $X2=0
+ $Y2=0
cc_436 N_A_398_74#_c_350_n N_A_225_74#_M1018_g 3.27596e-19 $X=6.53 $Y=1.285
+ $X2=0 $Y2=0
cc_437 N_A_398_74#_c_351_n N_A_225_74#_M1018_g 0.0110658f $X=6.53 $Y=1.285 $X2=0
+ $Y2=0
cc_438 N_A_398_74#_c_353_n N_A_225_74#_M1018_g 0.00923424f $X=7.21 $Y=2.02 $X2=0
+ $Y2=0
cc_439 N_A_398_74#_c_354_n N_A_225_74#_M1018_g 0.0190732f $X=6.53 $Y=1.12 $X2=0
+ $Y2=0
cc_440 N_A_398_74#_c_337_n N_A_225_74#_c_965_n 0.0394012f $X=3.005 $Y=2.24 $X2=0
+ $Y2=0
cc_441 N_A_398_74#_c_340_n N_A_225_74#_c_965_n 5.90715e-19 $X=2.13 $Y=0.515
+ $X2=0 $Y2=0
cc_442 N_A_398_74#_c_341_n N_A_225_74#_c_965_n 9.09485e-19 $X=2.945 $Y=0.34
+ $X2=0 $Y2=0
cc_443 N_A_398_74#_c_343_n N_A_225_74#_c_965_n 3.80136e-19 $X=2.95 $Y=1.62 $X2=0
+ $Y2=0
cc_444 N_A_398_74#_c_349_n N_A_225_74#_c_965_n 8.19775e-19 $X=2.95 $Y=1.455
+ $X2=0 $Y2=0
cc_445 N_A_398_74#_c_340_n N_A_225_74#_c_966_n 0.00102731f $X=2.13 $Y=0.515
+ $X2=0 $Y2=0
cc_446 N_A_398_74#_M1034_d N_A_225_74#_c_985_n 0.00247971f $X=2.04 $Y=1.84 $X2=0
+ $Y2=0
cc_447 N_A_398_74#_c_340_n N_A_225_74#_c_968_n 0.0120964f $X=2.13 $Y=0.515 $X2=0
+ $Y2=0
cc_448 N_A_398_74#_c_347_n N_A_1484_62#_M1004_g 0.00169096f $X=7.205 $Y=0.34
+ $X2=0 $Y2=0
cc_449 N_A_398_74#_c_353_n N_A_1484_62#_M1004_g 0.00722371f $X=7.21 $Y=2.02
+ $X2=0 $Y2=0
cc_450 N_A_398_74#_c_357_n N_A_1484_62#_c_1144_n 0.0245034f $X=7.325 $Y=2.465
+ $X2=0 $Y2=0
cc_451 N_A_398_74#_c_373_n N_A_1484_62#_c_1144_n 0.00174361f $X=7.21 $Y=2.185
+ $X2=0 $Y2=0
cc_452 N_A_398_74#_c_353_n N_A_1484_62#_c_1144_n 0.00915762f $X=7.21 $Y=2.02
+ $X2=0 $Y2=0
cc_453 N_A_398_74#_c_357_n N_A_1484_62#_c_1145_n 0.0281594f $X=7.325 $Y=2.465
+ $X2=0 $Y2=0
cc_454 N_A_398_74#_c_353_n N_A_1484_62#_c_1138_n 0.0479592f $X=7.21 $Y=2.02
+ $X2=0 $Y2=0
cc_455 N_A_398_74#_c_353_n N_A_1484_62#_c_1155_n 0.0127905f $X=7.21 $Y=2.02
+ $X2=0 $Y2=0
cc_456 N_A_398_74#_c_347_n N_A_1321_392#_M1003_d 0.00205663f $X=7.205 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_457 N_A_398_74#_c_357_n N_A_1321_392#_c_1243_n 0.0056037f $X=7.325 $Y=2.465
+ $X2=0 $Y2=0
cc_458 N_A_398_74#_c_369_n N_A_1321_392#_c_1243_n 0.0120091f $X=6.305 $Y=2.18
+ $X2=0 $Y2=0
cc_459 N_A_398_74#_c_346_n N_A_1321_392#_c_1243_n 0.0193592f $X=6.39 $Y=2.095
+ $X2=0 $Y2=0
cc_460 N_A_398_74#_c_373_n N_A_1321_392#_c_1243_n 0.0185355f $X=7.21 $Y=2.185
+ $X2=0 $Y2=0
cc_461 N_A_398_74#_c_353_n N_A_1321_392#_c_1243_n 0.0100218f $X=7.21 $Y=2.02
+ $X2=0 $Y2=0
cc_462 N_A_398_74#_c_346_n N_A_1321_392#_c_1233_n 0.00689075f $X=6.39 $Y=2.095
+ $X2=0 $Y2=0
cc_463 N_A_398_74#_c_350_n N_A_1321_392#_c_1233_n 0.0251223f $X=6.53 $Y=1.285
+ $X2=0 $Y2=0
cc_464 N_A_398_74#_c_351_n N_A_1321_392#_c_1233_n 0.00226999f $X=6.53 $Y=1.285
+ $X2=0 $Y2=0
cc_465 N_A_398_74#_c_352_n N_A_1321_392#_c_1233_n 0.00627822f $X=6.5 $Y=1.12
+ $X2=0 $Y2=0
cc_466 N_A_398_74#_c_353_n N_A_1321_392#_c_1233_n 0.0496067f $X=7.21 $Y=2.02
+ $X2=0 $Y2=0
cc_467 N_A_398_74#_c_354_n N_A_1321_392#_c_1233_n 0.00150671f $X=6.53 $Y=1.12
+ $X2=0 $Y2=0
cc_468 N_A_398_74#_c_357_n N_A_1321_392#_c_1244_n 0.00962924f $X=7.325 $Y=2.465
+ $X2=0 $Y2=0
cc_469 N_A_398_74#_c_373_n N_A_1321_392#_c_1244_n 0.00826905f $X=7.21 $Y=2.185
+ $X2=0 $Y2=0
cc_470 N_A_398_74#_c_357_n N_A_1321_392#_c_1245_n 0.0147433f $X=7.325 $Y=2.465
+ $X2=0 $Y2=0
cc_471 N_A_398_74#_c_373_n N_A_1321_392#_c_1245_n 0.0181771f $X=7.21 $Y=2.185
+ $X2=0 $Y2=0
cc_472 N_A_398_74#_c_347_n N_A_1321_392#_c_1236_n 0.0218291f $X=7.205 $Y=0.34
+ $X2=0 $Y2=0
cc_473 N_A_398_74#_c_350_n N_A_1321_392#_c_1236_n 0.00246577f $X=6.53 $Y=1.285
+ $X2=0 $Y2=0
cc_474 N_A_398_74#_c_353_n N_A_1321_392#_c_1236_n 0.0150761f $X=7.21 $Y=2.02
+ $X2=0 $Y2=0
cc_475 N_A_398_74#_c_354_n N_A_1321_392#_c_1236_n 0.00408225f $X=6.53 $Y=1.12
+ $X2=0 $Y2=0
cc_476 N_A_398_74#_c_346_n N_A_1321_392#_c_1237_n 0.0101597f $X=6.39 $Y=2.095
+ $X2=0 $Y2=0
cc_477 N_A_398_74#_c_350_n N_A_1321_392#_c_1237_n 0.00157906f $X=6.53 $Y=1.285
+ $X2=0 $Y2=0
cc_478 N_A_398_74#_c_353_n N_A_1321_392#_c_1237_n 0.0119049f $X=7.21 $Y=2.02
+ $X2=0 $Y2=0
cc_479 N_A_398_74#_c_357_n N_A_1321_392#_c_1249_n 0.00385577f $X=7.325 $Y=2.465
+ $X2=0 $Y2=0
cc_480 N_A_398_74#_c_341_n N_A_27_74#_M1027_s 0.00416589f $X=2.945 $Y=0.34 $X2=0
+ $Y2=0
cc_481 N_A_398_74#_M1034_d N_A_27_74#_c_1515_n 0.00596624f $X=2.04 $Y=1.84 $X2=0
+ $Y2=0
cc_482 N_A_398_74#_c_337_n N_A_27_74#_c_1515_n 0.00882557f $X=3.005 $Y=2.24
+ $X2=0 $Y2=0
cc_483 N_A_398_74#_c_453_p N_A_27_74#_c_1515_n 0.0385621f $X=2.19 $Y=2.575 $X2=0
+ $Y2=0
cc_484 N_A_398_74#_c_358_n N_A_27_74#_c_1515_n 0.039591f $X=3.625 $Y=2.99 $X2=0
+ $Y2=0
cc_485 N_A_398_74#_c_343_n N_A_27_74#_c_1515_n 0.0182631f $X=2.95 $Y=1.62 $X2=0
+ $Y2=0
cc_486 N_A_398_74#_c_337_n N_A_27_74#_c_1509_n 0.00357538f $X=3.005 $Y=2.24
+ $X2=0 $Y2=0
cc_487 N_A_398_74#_c_340_n N_A_27_74#_c_1509_n 0.0119813f $X=2.13 $Y=0.515 $X2=0
+ $Y2=0
cc_488 N_A_398_74#_c_343_n N_A_27_74#_c_1509_n 0.0461461f $X=2.95 $Y=1.62 $X2=0
+ $Y2=0
cc_489 N_A_398_74#_c_349_n N_A_27_74#_c_1509_n 0.023467f $X=2.95 $Y=1.455 $X2=0
+ $Y2=0
cc_490 N_A_398_74#_c_340_n N_A_27_74#_c_1511_n 0.0206593f $X=2.13 $Y=0.515 $X2=0
+ $Y2=0
cc_491 N_A_398_74#_c_341_n N_A_27_74#_c_1511_n 0.0239262f $X=2.945 $Y=0.34 $X2=0
+ $Y2=0
cc_492 N_A_398_74#_c_349_n N_A_27_74#_c_1511_n 0.0244211f $X=2.95 $Y=1.455 $X2=0
+ $Y2=0
cc_493 N_A_398_74#_c_364_n N_VPWR_M1011_d 0.0102003f $X=4.515 $Y=2.25 $X2=0
+ $Y2=0
cc_494 N_A_398_74#_c_365_n N_VPWR_M1011_d 0.0115964f $X=4.6 $Y=2.905 $X2=0 $Y2=0
cc_495 N_A_398_74#_c_368_n N_VPWR_M1007_d 0.00453684f $X=5.425 $Y=2.905 $X2=0
+ $Y2=0
cc_496 N_A_398_74#_c_369_n N_VPWR_M1007_d 0.00621806f $X=6.305 $Y=2.18 $X2=0
+ $Y2=0
cc_497 N_A_398_74#_c_453_p N_VPWR_c_1578_n 0.0211373f $X=2.19 $Y=2.575 $X2=0
+ $Y2=0
cc_498 N_A_398_74#_c_359_n N_VPWR_c_1578_n 0.0125885f $X=2.275 $Y=2.99 $X2=0
+ $Y2=0
cc_499 N_A_398_74#_c_358_n N_VPWR_c_1579_n 0.0132711f $X=3.625 $Y=2.99 $X2=0
+ $Y2=0
cc_500 N_A_398_74#_c_363_n N_VPWR_c_1579_n 0.00998705f $X=3.71 $Y=2.905 $X2=0
+ $Y2=0
cc_501 N_A_398_74#_c_365_n N_VPWR_c_1579_n 0.00670109f $X=4.6 $Y=2.905 $X2=0
+ $Y2=0
cc_502 N_A_398_74#_c_367_n N_VPWR_c_1579_n 0.00852847f $X=4.685 $Y=2.99 $X2=0
+ $Y2=0
cc_503 N_A_398_74#_c_366_n N_VPWR_c_1580_n 0.0147865f $X=5.34 $Y=2.99 $X2=0
+ $Y2=0
cc_504 N_A_398_74#_c_368_n N_VPWR_c_1580_n 0.0356946f $X=5.425 $Y=2.905 $X2=0
+ $Y2=0
cc_505 N_A_398_74#_c_369_n N_VPWR_c_1580_n 0.0172533f $X=6.305 $Y=2.18 $X2=0
+ $Y2=0
cc_506 N_A_398_74#_c_363_n N_VPWR_c_1589_n 0.00929868f $X=3.71 $Y=2.905 $X2=0
+ $Y2=0
cc_507 N_A_398_74#_c_364_n N_VPWR_c_1589_n 0.0225521f $X=4.515 $Y=2.25 $X2=0
+ $Y2=0
cc_508 N_A_398_74#_c_365_n N_VPWR_c_1589_n 0.0192298f $X=4.6 $Y=2.905 $X2=0
+ $Y2=0
cc_509 N_A_398_74#_c_366_n N_VPWR_c_1590_n 0.0537108f $X=5.34 $Y=2.99 $X2=0
+ $Y2=0
cc_510 N_A_398_74#_c_367_n N_VPWR_c_1590_n 0.0115893f $X=4.685 $Y=2.99 $X2=0
+ $Y2=0
cc_511 N_A_398_74#_c_358_n N_VPWR_c_1594_n 0.0975198f $X=3.625 $Y=2.99 $X2=0
+ $Y2=0
cc_512 N_A_398_74#_c_359_n N_VPWR_c_1594_n 0.0121664f $X=2.275 $Y=2.99 $X2=0
+ $Y2=0
cc_513 N_A_398_74#_c_357_n N_VPWR_c_1595_n 0.00327026f $X=7.325 $Y=2.465 $X2=0
+ $Y2=0
cc_514 N_A_398_74#_c_357_n N_VPWR_c_1576_n 0.00420634f $X=7.325 $Y=2.465 $X2=0
+ $Y2=0
cc_515 N_A_398_74#_c_358_n N_VPWR_c_1576_n 0.0514634f $X=3.625 $Y=2.99 $X2=0
+ $Y2=0
cc_516 N_A_398_74#_c_359_n N_VPWR_c_1576_n 0.00660537f $X=2.275 $Y=2.99 $X2=0
+ $Y2=0
cc_517 N_A_398_74#_c_366_n N_VPWR_c_1576_n 0.0278398f $X=5.34 $Y=2.99 $X2=0
+ $Y2=0
cc_518 N_A_398_74#_c_367_n N_VPWR_c_1576_n 0.00583135f $X=4.685 $Y=2.99 $X2=0
+ $Y2=0
cc_519 N_A_398_74#_c_363_n A_716_463# 0.0020949f $X=3.71 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_520 N_A_398_74#_c_369_n A_1220_347# 0.0121024f $X=6.305 $Y=2.18 $X2=-0.19
+ $Y2=-0.245
cc_521 N_A_398_74#_c_346_n A_1220_347# 0.00485418f $X=6.39 $Y=2.095 $X2=-0.19
+ $Y2=-0.245
cc_522 N_A_398_74#_c_342_n N_VGND_c_1833_n 0.0109685f $X=2.215 $Y=0.34 $X2=0
+ $Y2=0
cc_523 N_A_398_74#_M1017_g N_VGND_c_1834_n 0.00126697f $X=3.585 $Y=0.58 $X2=0
+ $Y2=0
cc_524 N_A_398_74#_c_348_n N_VGND_c_1835_n 0.00917417f $X=6.475 $Y=0.34 $X2=0
+ $Y2=0
cc_525 N_A_398_74#_c_352_n N_VGND_c_1835_n 0.0285193f $X=6.5 $Y=1.12 $X2=0 $Y2=0
cc_526 N_A_398_74#_c_354_n N_VGND_c_1835_n 4.42772e-19 $X=6.53 $Y=1.12 $X2=0
+ $Y2=0
cc_527 N_A_398_74#_M1017_g N_VGND_c_1843_n 0.00434272f $X=3.585 $Y=0.58 $X2=0
+ $Y2=0
cc_528 N_A_398_74#_c_341_n N_VGND_c_1843_n 0.0586507f $X=2.945 $Y=0.34 $X2=0
+ $Y2=0
cc_529 N_A_398_74#_c_342_n N_VGND_c_1843_n 0.0121867f $X=2.215 $Y=0.34 $X2=0
+ $Y2=0
cc_530 N_A_398_74#_c_347_n N_VGND_c_1850_n 0.0587172f $X=7.205 $Y=0.34 $X2=0
+ $Y2=0
cc_531 N_A_398_74#_c_348_n N_VGND_c_1850_n 0.0121867f $X=6.475 $Y=0.34 $X2=0
+ $Y2=0
cc_532 N_A_398_74#_c_354_n N_VGND_c_1850_n 0.00278271f $X=6.53 $Y=1.12 $X2=0
+ $Y2=0
cc_533 N_A_398_74#_c_347_n N_VGND_c_1851_n 0.00636506f $X=7.205 $Y=0.34 $X2=0
+ $Y2=0
cc_534 N_A_398_74#_c_353_n N_VGND_c_1851_n 0.00405322f $X=7.21 $Y=2.02 $X2=0
+ $Y2=0
cc_535 N_A_398_74#_M1017_g N_VGND_c_1854_n 0.00822443f $X=3.585 $Y=0.58 $X2=0
+ $Y2=0
cc_536 N_A_398_74#_c_341_n N_VGND_c_1854_n 0.0333627f $X=2.945 $Y=0.34 $X2=0
+ $Y2=0
cc_537 N_A_398_74#_c_342_n N_VGND_c_1854_n 0.00660921f $X=2.215 $Y=0.34 $X2=0
+ $Y2=0
cc_538 N_A_398_74#_c_347_n N_VGND_c_1854_n 0.033365f $X=7.205 $Y=0.34 $X2=0
+ $Y2=0
cc_539 N_A_398_74#_c_348_n N_VGND_c_1854_n 0.00660921f $X=6.475 $Y=0.34 $X2=0
+ $Y2=0
cc_540 N_A_398_74#_c_354_n N_VGND_c_1854_n 0.00359494f $X=6.53 $Y=1.12 $X2=0
+ $Y2=0
cc_541 N_A_398_74#_c_348_n A_1225_74# 7.18263e-19 $X=6.475 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_542 N_A_398_74#_c_352_n A_1225_74# 0.00947773f $X=6.5 $Y=1.12 $X2=-0.19
+ $Y2=-0.245
cc_543 N_A_398_74#_c_353_n A_1436_88# 0.00181261f $X=7.21 $Y=2.02 $X2=-0.19
+ $Y2=-0.245
cc_544 N_A_767_402#_c_604_n N_A_612_74#_c_684_n 0.0185431f $X=3.925 $Y=2.24
+ $X2=0 $Y2=0
cc_545 N_A_767_402#_c_606_n N_A_612_74#_c_684_n 0.0150553f $X=4.855 $Y=1.867
+ $X2=0 $Y2=0
cc_546 N_A_767_402#_c_607_n N_A_612_74#_c_684_n 0.00439413f $X=4.94 $Y=2.295
+ $X2=0 $Y2=0
cc_547 N_A_767_402#_c_607_n N_A_612_74#_c_699_n 0.00397084f $X=4.94 $Y=2.295
+ $X2=0 $Y2=0
cc_548 N_A_767_402#_c_608_n N_A_612_74#_c_699_n 0.00775981f $X=5.085 $Y=2.515
+ $X2=0 $Y2=0
cc_549 N_A_767_402#_c_602_n N_A_612_74#_c_685_n 0.00995281f $X=4.395 $Y=1.065
+ $X2=0 $Y2=0
cc_550 N_A_767_402#_c_603_n N_A_612_74#_c_685_n 0.00382576f $X=4.395 $Y=0.975
+ $X2=0 $Y2=0
cc_551 N_A_767_402#_c_598_n N_A_612_74#_c_688_n 0.00306844f $X=3.975 $Y=0.9
+ $X2=0 $Y2=0
cc_552 N_A_767_402#_c_603_n N_A_612_74#_c_688_n 3.7427e-19 $X=4.395 $Y=0.975
+ $X2=0 $Y2=0
cc_553 N_A_767_402#_c_600_n N_A_612_74#_c_689_n 0.00297558f $X=4.05 $Y=0.975
+ $X2=0 $Y2=0
cc_554 N_A_767_402#_c_604_n N_A_612_74#_c_690_n 0.00174649f $X=3.925 $Y=2.24
+ $X2=0 $Y2=0
cc_555 N_A_767_402#_c_599_n N_A_612_74#_c_690_n 0.00182267f $X=4.23 $Y=0.975
+ $X2=0 $Y2=0
cc_556 N_A_767_402#_c_601_n N_A_612_74#_c_690_n 0.0126255f $X=4.305 $Y=1.7 $X2=0
+ $Y2=0
cc_557 N_A_767_402#_c_606_n N_A_612_74#_c_690_n 0.0475354f $X=4.855 $Y=1.867
+ $X2=0 $Y2=0
cc_558 N_A_767_402#_c_602_n N_A_612_74#_c_690_n 0.0290223f $X=4.395 $Y=1.065
+ $X2=0 $Y2=0
cc_559 N_A_767_402#_c_603_n N_A_612_74#_c_690_n 0.00105029f $X=4.395 $Y=0.975
+ $X2=0 $Y2=0
cc_560 N_A_767_402#_c_602_n N_A_612_74#_c_691_n 0.00128907f $X=4.395 $Y=1.065
+ $X2=0 $Y2=0
cc_561 N_A_767_402#_c_604_n N_A_612_74#_c_692_n 4.37211e-19 $X=3.925 $Y=2.24
+ $X2=0 $Y2=0
cc_562 N_A_767_402#_c_604_n N_A_612_74#_c_694_n 0.00308777f $X=3.925 $Y=2.24
+ $X2=0 $Y2=0
cc_563 N_A_767_402#_c_600_n N_A_612_74#_c_694_n 0.0059641f $X=4.05 $Y=0.975
+ $X2=0 $Y2=0
cc_564 N_A_767_402#_c_601_n N_A_612_74#_c_694_n 3.58867e-19 $X=4.305 $Y=1.7
+ $X2=0 $Y2=0
cc_565 N_A_767_402#_c_606_n N_A_612_74#_c_694_n 0.00151836f $X=4.855 $Y=1.867
+ $X2=0 $Y2=0
cc_566 N_A_767_402#_c_602_n N_A_612_74#_c_694_n 0.00746874f $X=4.395 $Y=1.065
+ $X2=0 $Y2=0
cc_567 N_A_767_402#_c_603_n N_A_612_74#_c_694_n 0.00363451f $X=4.395 $Y=0.975
+ $X2=0 $Y2=0
cc_568 N_A_767_402#_c_601_n N_A_612_74#_c_695_n 7.77514e-19 $X=4.305 $Y=1.7
+ $X2=0 $Y2=0
cc_569 N_A_767_402#_c_606_n N_A_612_74#_c_695_n 0.0206269f $X=4.855 $Y=1.867
+ $X2=0 $Y2=0
cc_570 N_A_767_402#_c_602_n N_A_612_74#_c_695_n 0.0261626f $X=4.395 $Y=1.065
+ $X2=0 $Y2=0
cc_571 N_A_767_402#_c_601_n N_A_612_74#_c_697_n 0.0148476f $X=4.305 $Y=1.7 $X2=0
+ $Y2=0
cc_572 N_A_767_402#_c_606_n N_A_612_74#_c_697_n 4.25161e-19 $X=4.855 $Y=1.867
+ $X2=0 $Y2=0
cc_573 N_A_767_402#_c_602_n N_A_612_74#_c_697_n 0.00234761f $X=4.395 $Y=1.065
+ $X2=0 $Y2=0
cc_574 N_A_767_402#_c_603_n N_A_612_74#_c_697_n 0.00699025f $X=4.395 $Y=0.975
+ $X2=0 $Y2=0
cc_575 N_A_767_402#_c_607_n N_SET_B_c_832_n 0.0029814f $X=4.94 $Y=2.295 $X2=0
+ $Y2=0
cc_576 N_A_767_402#_c_607_n N_SET_B_c_833_n 3.72148e-19 $X=4.94 $Y=2.295 $X2=0
+ $Y2=0
cc_577 N_A_767_402#_c_608_n N_SET_B_c_833_n 0.00158145f $X=5.085 $Y=2.515 $X2=0
+ $Y2=0
cc_578 N_A_767_402#_c_602_n N_SET_B_M1020_g 9.88858e-19 $X=4.395 $Y=1.065 $X2=0
+ $Y2=0
cc_579 N_A_767_402#_c_606_n N_SET_B_c_827_n 2.23271e-19 $X=4.855 $Y=1.867 $X2=0
+ $Y2=0
cc_580 N_A_767_402#_c_606_n N_SET_B_c_829_n 0.0156891f $X=4.855 $Y=1.867 $X2=0
+ $Y2=0
cc_581 N_A_767_402#_c_606_n N_SET_B_c_830_n 0.00255214f $X=4.855 $Y=1.867 $X2=0
+ $Y2=0
cc_582 N_A_767_402#_c_604_n N_A_225_74#_c_974_n 0.00222191f $X=3.925 $Y=2.24
+ $X2=0 $Y2=0
cc_583 N_A_767_402#_c_604_n N_A_225_74#_c_976_n 0.0239039f $X=3.925 $Y=2.24
+ $X2=0 $Y2=0
cc_584 N_A_767_402#_c_604_n N_A_225_74#_c_977_n 0.0103562f $X=3.925 $Y=2.24
+ $X2=0 $Y2=0
cc_585 N_A_767_402#_c_604_n N_VPWR_c_1579_n 0.00318511f $X=3.925 $Y=2.24 $X2=0
+ $Y2=0
cc_586 N_A_767_402#_c_604_n N_VPWR_c_1589_n 0.0030685f $X=3.925 $Y=2.24 $X2=0
+ $Y2=0
cc_587 N_A_767_402#_c_604_n N_VPWR_c_1576_n 8.51577e-19 $X=3.925 $Y=2.24 $X2=0
+ $Y2=0
cc_588 N_A_767_402#_c_602_n N_VGND_M1001_d 0.00118908f $X=4.395 $Y=1.065 $X2=0
+ $Y2=0
cc_589 N_A_767_402#_c_598_n N_VGND_c_1834_n 0.0098944f $X=3.975 $Y=0.9 $X2=0
+ $Y2=0
cc_590 N_A_767_402#_c_599_n N_VGND_c_1834_n 0.0079331f $X=4.23 $Y=0.975 $X2=0
+ $Y2=0
cc_591 N_A_767_402#_c_602_n N_VGND_c_1834_n 0.00929432f $X=4.395 $Y=1.065 $X2=0
+ $Y2=0
cc_592 N_A_767_402#_c_603_n N_VGND_c_1834_n 6.63116e-19 $X=4.395 $Y=0.975 $X2=0
+ $Y2=0
cc_593 N_A_767_402#_c_602_n N_VGND_c_1835_n 0.00958081f $X=4.395 $Y=1.065 $X2=0
+ $Y2=0
cc_594 N_A_767_402#_c_602_n N_VGND_c_1840_n 0.00824154f $X=4.395 $Y=1.065 $X2=0
+ $Y2=0
cc_595 N_A_767_402#_c_598_n N_VGND_c_1843_n 0.00383152f $X=3.975 $Y=0.9 $X2=0
+ $Y2=0
cc_596 N_A_767_402#_c_598_n N_VGND_c_1854_n 0.0075725f $X=3.975 $Y=0.9 $X2=0
+ $Y2=0
cc_597 N_A_767_402#_c_602_n N_VGND_c_1854_n 0.0209055f $X=4.395 $Y=1.065 $X2=0
+ $Y2=0
cc_598 N_A_612_74#_c_684_n N_SET_B_c_832_n 0.00538992f $X=4.86 $Y=2.15 $X2=0
+ $Y2=0
cc_599 N_A_612_74#_c_686_n N_SET_B_c_832_n 0.00523885f $X=6.025 $Y=1.66 $X2=0
+ $Y2=0
cc_600 N_A_612_74#_c_699_n N_SET_B_c_833_n 0.0141981f $X=4.86 $Y=2.24 $X2=0
+ $Y2=0
cc_601 N_A_612_74#_c_686_n N_SET_B_c_833_n 0.00677794f $X=6.025 $Y=1.66 $X2=0
+ $Y2=0
cc_602 N_A_612_74#_c_684_n N_SET_B_M1020_g 0.00427675f $X=4.86 $Y=2.15 $X2=0
+ $Y2=0
cc_603 N_A_612_74#_c_685_n N_SET_B_M1020_g 0.0531748f $X=5.1 $Y=1.12 $X2=0 $Y2=0
cc_604 N_A_612_74#_c_686_n N_SET_B_M1020_g 0.0228094f $X=6.025 $Y=1.66 $X2=0
+ $Y2=0
cc_605 N_A_612_74#_M1031_g N_SET_B_M1020_g 0.0120624f $X=6.05 $Y=0.69 $X2=0
+ $Y2=0
cc_606 N_A_612_74#_c_691_n N_SET_B_M1020_g 0.0144612f $X=5.805 $Y=1.285 $X2=0
+ $Y2=0
cc_607 N_A_612_74#_c_695_n N_SET_B_M1020_g 0.00275571f $X=4.935 $Y=1.285 $X2=0
+ $Y2=0
cc_608 N_A_612_74#_c_696_n N_SET_B_M1020_g 8.93876e-19 $X=5.97 $Y=1.285 $X2=0
+ $Y2=0
cc_609 N_A_612_74#_c_686_n N_SET_B_c_826_n 0.0110709f $X=6.025 $Y=1.66 $X2=0
+ $Y2=0
cc_610 N_A_612_74#_c_691_n N_SET_B_c_826_n 0.00599672f $X=5.805 $Y=1.285 $X2=0
+ $Y2=0
cc_611 N_A_612_74#_c_696_n N_SET_B_c_826_n 0.010239f $X=5.97 $Y=1.285 $X2=0
+ $Y2=0
cc_612 N_A_612_74#_c_686_n N_SET_B_c_827_n 0.00132786f $X=6.025 $Y=1.66 $X2=0
+ $Y2=0
cc_613 N_A_612_74#_c_691_n N_SET_B_c_827_n 0.00787805f $X=5.805 $Y=1.285 $X2=0
+ $Y2=0
cc_614 N_A_612_74#_c_684_n N_SET_B_c_829_n 0.00301198f $X=4.86 $Y=2.15 $X2=0
+ $Y2=0
cc_615 N_A_612_74#_c_686_n N_SET_B_c_829_n 0.00315116f $X=6.025 $Y=1.66 $X2=0
+ $Y2=0
cc_616 N_A_612_74#_c_691_n N_SET_B_c_829_n 0.0292376f $X=5.805 $Y=1.285 $X2=0
+ $Y2=0
cc_617 N_A_612_74#_c_695_n N_SET_B_c_829_n 0.00150495f $X=4.935 $Y=1.285 $X2=0
+ $Y2=0
cc_618 N_A_612_74#_c_684_n N_SET_B_c_830_n 0.0172323f $X=4.86 $Y=2.15 $X2=0
+ $Y2=0
cc_619 N_A_612_74#_c_686_n N_SET_B_c_830_n 0.0102234f $X=6.025 $Y=1.66 $X2=0
+ $Y2=0
cc_620 N_A_612_74#_c_691_n N_SET_B_c_830_n 0.00115614f $X=5.805 $Y=1.285 $X2=0
+ $Y2=0
cc_621 N_A_612_74#_c_693_n N_A_225_74#_c_960_n 3.27724e-19 $X=3.41 $Y=1.215
+ $X2=0 $Y2=0
cc_622 N_A_612_74#_c_688_n N_A_225_74#_M1027_g 0.00260688f $X=3.37 $Y=0.58 $X2=0
+ $Y2=0
cc_623 N_A_612_74#_c_701_n N_A_225_74#_c_976_n 0.00538483f $X=3.28 $Y=2.515
+ $X2=0 $Y2=0
cc_624 N_A_612_74#_c_692_n N_A_225_74#_c_976_n 0.00241442f $X=3.285 $Y=2.295
+ $X2=0 $Y2=0
cc_625 N_A_612_74#_c_699_n N_A_225_74#_c_977_n 0.00882199f $X=4.86 $Y=2.24 $X2=0
+ $Y2=0
cc_626 N_A_612_74#_c_686_n N_A_225_74#_c_977_n 0.0104164f $X=6.025 $Y=1.66 $X2=0
+ $Y2=0
cc_627 N_A_612_74#_c_686_n N_A_225_74#_M1013_g 0.0313943f $X=6.025 $Y=1.66 $X2=0
+ $Y2=0
cc_628 N_A_612_74#_c_686_n N_A_225_74#_c_963_n 0.00755438f $X=6.025 $Y=1.66
+ $X2=0 $Y2=0
cc_629 N_A_612_74#_c_686_n N_A_1321_392#_c_1245_n 6.56869e-19 $X=6.025 $Y=1.66
+ $X2=0 $Y2=0
cc_630 N_A_612_74#_c_701_n N_A_27_74#_c_1515_n 0.0184847f $X=3.28 $Y=2.515 $X2=0
+ $Y2=0
cc_631 N_A_612_74#_c_692_n N_A_27_74#_c_1515_n 0.00522874f $X=3.285 $Y=2.295
+ $X2=0 $Y2=0
cc_632 N_A_612_74#_c_686_n N_VPWR_c_1580_n 0.00240863f $X=6.025 $Y=1.66 $X2=0
+ $Y2=0
cc_633 N_A_612_74#_c_686_n N_VPWR_c_1576_n 9.39239e-19 $X=6.025 $Y=1.66 $X2=0
+ $Y2=0
cc_634 N_A_612_74#_c_685_n N_VGND_c_1834_n 0.00327534f $X=5.1 $Y=1.12 $X2=0
+ $Y2=0
cc_635 N_A_612_74#_c_688_n N_VGND_c_1834_n 0.00786568f $X=3.37 $Y=0.58 $X2=0
+ $Y2=0
cc_636 N_A_612_74#_c_694_n N_VGND_c_1834_n 0.00302077f $X=4.05 $Y=1.215 $X2=0
+ $Y2=0
cc_637 N_A_612_74#_c_686_n N_VGND_c_1835_n 0.00133462f $X=6.025 $Y=1.66 $X2=0
+ $Y2=0
cc_638 N_A_612_74#_M1031_g N_VGND_c_1835_n 0.0144111f $X=6.05 $Y=0.69 $X2=0
+ $Y2=0
cc_639 N_A_612_74#_c_691_n N_VGND_c_1835_n 0.010974f $X=5.805 $Y=1.285 $X2=0
+ $Y2=0
cc_640 N_A_612_74#_c_696_n N_VGND_c_1835_n 0.0156226f $X=5.97 $Y=1.285 $X2=0
+ $Y2=0
cc_641 N_A_612_74#_c_685_n N_VGND_c_1840_n 0.00417521f $X=5.1 $Y=1.12 $X2=0
+ $Y2=0
cc_642 N_A_612_74#_c_688_n N_VGND_c_1843_n 0.0109942f $X=3.37 $Y=0.58 $X2=0
+ $Y2=0
cc_643 N_A_612_74#_M1031_g N_VGND_c_1850_n 0.00383152f $X=6.05 $Y=0.69 $X2=0
+ $Y2=0
cc_644 N_A_612_74#_c_685_n N_VGND_c_1854_n 0.00479212f $X=5.1 $Y=1.12 $X2=0
+ $Y2=0
cc_645 N_A_612_74#_M1031_g N_VGND_c_1854_n 0.00758607f $X=6.05 $Y=0.69 $X2=0
+ $Y2=0
cc_646 N_A_612_74#_c_688_n N_VGND_c_1854_n 0.00904371f $X=3.37 $Y=0.58 $X2=0
+ $Y2=0
cc_647 N_SET_B_c_833_n N_A_225_74#_c_977_n 0.00909901f $X=5.31 $Y=2.24 $X2=0
+ $Y2=0
cc_648 N_SET_B_c_826_n N_A_225_74#_c_962_n 0.00400315f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_649 N_SET_B_c_826_n N_A_225_74#_c_963_n 0.00592114f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_650 N_SET_B_c_826_n N_A_225_74#_M1018_g 0.00633119f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_651 N_SET_B_c_822_n N_A_1484_62#_M1004_g 0.040286f $X=7.885 $Y=0.935 $X2=0
+ $Y2=0
cc_652 N_SET_B_c_823_n N_A_1484_62#_M1004_g 0.00387759f $X=8.31 $Y=1.385 $X2=0
+ $Y2=0
cc_653 N_SET_B_c_825_n N_A_1484_62#_c_1144_n 0.0211372f $X=8.31 $Y=1.85 $X2=0
+ $Y2=0
cc_654 N_SET_B_c_826_n N_A_1484_62#_c_1144_n 0.00374132f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_655 N_SET_B_c_831_n N_A_1484_62#_c_1144_n 0.00130941f $X=8.35 $Y=1.345 $X2=0
+ $Y2=0
cc_656 N_SET_B_c_835_n N_A_1484_62#_c_1145_n 0.0211372f $X=8.195 $Y=2.375 $X2=0
+ $Y2=0
cc_657 N_SET_B_c_836_n N_A_1484_62#_c_1145_n 0.00997743f $X=8.195 $Y=2.465 $X2=0
+ $Y2=0
cc_658 N_SET_B_c_823_n N_A_1484_62#_c_1138_n 0.0102598f $X=8.31 $Y=1.385 $X2=0
+ $Y2=0
cc_659 N_SET_B_c_826_n N_A_1484_62#_c_1138_n 0.0238932f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_660 SET_B N_A_1484_62#_c_1138_n 2.66384e-19 $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_661 N_SET_B_c_831_n N_A_1484_62#_c_1138_n 0.0214964f $X=8.35 $Y=1.345 $X2=0
+ $Y2=0
cc_662 N_SET_B_c_822_n N_A_1484_62#_c_1139_n 0.0046649f $X=7.885 $Y=0.935 $X2=0
+ $Y2=0
cc_663 N_SET_B_c_823_n N_A_1484_62#_c_1139_n 0.018828f $X=8.31 $Y=1.385 $X2=0
+ $Y2=0
cc_664 N_SET_B_c_826_n N_A_1484_62#_c_1139_n 0.00842616f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_665 SET_B N_A_1484_62#_c_1139_n 0.001949f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_666 N_SET_B_c_831_n N_A_1484_62#_c_1139_n 0.0251801f $X=8.35 $Y=1.345 $X2=0
+ $Y2=0
cc_667 N_SET_B_c_822_n N_A_1484_62#_c_1155_n 0.00326479f $X=7.885 $Y=0.935 $X2=0
+ $Y2=0
cc_668 N_SET_B_c_823_n N_A_1484_62#_c_1155_n 0.00123586f $X=8.31 $Y=1.385 $X2=0
+ $Y2=0
cc_669 N_SET_B_c_823_n N_A_1484_62#_c_1143_n 0.0230148f $X=8.31 $Y=1.385 $X2=0
+ $Y2=0
cc_670 N_SET_B_c_826_n N_A_1484_62#_c_1143_n 0.00840235f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_671 N_SET_B_c_831_n N_A_1484_62#_c_1143_n 0.00111154f $X=8.35 $Y=1.345 $X2=0
+ $Y2=0
cc_672 N_SET_B_c_824_n N_A_1321_392#_c_1227_n 0.0121016f $X=8.31 $Y=1.645 $X2=0
+ $Y2=0
cc_673 N_SET_B_c_835_n N_A_1321_392#_c_1227_n 0.00707185f $X=8.195 $Y=2.375
+ $X2=0 $Y2=0
cc_674 N_SET_B_c_823_n N_A_1321_392#_M1002_g 0.0053109f $X=8.31 $Y=1.385 $X2=0
+ $Y2=0
cc_675 N_SET_B_c_831_n N_A_1321_392#_M1002_g 0.00102865f $X=8.35 $Y=1.345 $X2=0
+ $Y2=0
cc_676 N_SET_B_c_836_n N_A_1321_392#_c_1239_n 0.00707185f $X=8.195 $Y=2.465
+ $X2=0 $Y2=0
cc_677 N_SET_B_c_826_n N_A_1321_392#_c_1243_n 0.00168835f $X=8.255 $Y=1.665
+ $X2=0 $Y2=0
cc_678 N_SET_B_c_826_n N_A_1321_392#_c_1233_n 0.0101492f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_679 N_SET_B_c_835_n N_A_1321_392#_c_1246_n 0.00510032f $X=8.195 $Y=2.375
+ $X2=0 $Y2=0
cc_680 N_SET_B_c_836_n N_A_1321_392#_c_1246_n 0.00594531f $X=8.195 $Y=2.465
+ $X2=0 $Y2=0
cc_681 N_SET_B_c_826_n N_A_1321_392#_c_1246_n 0.012116f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_682 N_SET_B_c_831_n N_A_1321_392#_c_1246_n 0.00197365f $X=8.35 $Y=1.345 $X2=0
+ $Y2=0
cc_683 N_SET_B_c_836_n N_A_1321_392#_c_1247_n 0.00859289f $X=8.195 $Y=2.465
+ $X2=0 $Y2=0
cc_684 N_SET_B_c_823_n N_A_1321_392#_c_1234_n 0.00165128f $X=8.31 $Y=1.385 $X2=0
+ $Y2=0
cc_685 N_SET_B_c_835_n N_A_1321_392#_c_1234_n 0.00252386f $X=8.195 $Y=2.375
+ $X2=0 $Y2=0
cc_686 SET_B N_A_1321_392#_c_1234_n 0.00699971f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_687 N_SET_B_c_831_n N_A_1321_392#_c_1234_n 0.0218297f $X=8.35 $Y=1.345 $X2=0
+ $Y2=0
cc_688 N_SET_B_c_823_n N_A_1321_392#_c_1235_n 0.0121016f $X=8.31 $Y=1.385 $X2=0
+ $Y2=0
cc_689 SET_B N_A_1321_392#_c_1235_n 0.00410251f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_690 N_SET_B_c_831_n N_A_1321_392#_c_1235_n 0.0022247f $X=8.35 $Y=1.345 $X2=0
+ $Y2=0
cc_691 N_SET_B_c_826_n N_A_1321_392#_c_1237_n 0.020282f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_692 N_SET_B_c_836_n N_A_1321_392#_c_1249_n 4.70987e-19 $X=8.195 $Y=2.465
+ $X2=0 $Y2=0
cc_693 N_SET_B_c_826_n N_A_1321_392#_c_1249_n 0.00323313f $X=8.255 $Y=1.665
+ $X2=0 $Y2=0
cc_694 N_SET_B_c_835_n N_A_1321_392#_c_1250_n 0.00201834f $X=8.195 $Y=2.375
+ $X2=0 $Y2=0
cc_695 N_SET_B_c_836_n N_A_1321_392#_c_1250_n 0.00307667f $X=8.195 $Y=2.465
+ $X2=0 $Y2=0
cc_696 N_SET_B_c_825_n N_A_1321_392#_c_1250_n 0.00153883f $X=8.31 $Y=1.85 $X2=0
+ $Y2=0
cc_697 SET_B N_A_1321_392#_c_1250_n 0.00301214f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_698 N_SET_B_c_831_n N_A_1321_392#_c_1250_n 0.00864852f $X=8.35 $Y=1.345 $X2=0
+ $Y2=0
cc_699 N_SET_B_c_826_n N_VPWR_M1007_d 0.00263614f $X=8.255 $Y=1.665 $X2=0 $Y2=0
cc_700 N_SET_B_c_833_n N_VPWR_c_1580_n 0.00130931f $X=5.31 $Y=2.24 $X2=0 $Y2=0
cc_701 N_SET_B_c_836_n N_VPWR_c_1581_n 0.00373065f $X=8.195 $Y=2.465 $X2=0 $Y2=0
cc_702 N_SET_B_c_836_n N_VPWR_c_1582_n 0.00327326f $X=8.195 $Y=2.465 $X2=0 $Y2=0
cc_703 N_SET_B_c_836_n N_VPWR_c_1596_n 0.00445602f $X=8.195 $Y=2.465 $X2=0 $Y2=0
cc_704 N_SET_B_c_836_n N_VPWR_c_1576_n 0.00459843f $X=8.195 $Y=2.465 $X2=0 $Y2=0
cc_705 N_SET_B_c_826_n A_1220_347# 0.00203928f $X=8.255 $Y=1.665 $X2=-0.19
+ $Y2=-0.245
cc_706 N_SET_B_M1020_g N_VGND_c_1835_n 0.0111202f $X=5.49 $Y=0.8 $X2=0 $Y2=0
cc_707 N_SET_B_c_826_n N_VGND_c_1835_n 6.575e-19 $X=8.255 $Y=1.665 $X2=0 $Y2=0
cc_708 N_SET_B_M1020_g N_VGND_c_1840_n 0.00434252f $X=5.49 $Y=0.8 $X2=0 $Y2=0
cc_709 N_SET_B_c_822_n N_VGND_c_1850_n 0.00438299f $X=7.885 $Y=0.935 $X2=0 $Y2=0
cc_710 N_SET_B_c_822_n N_VGND_c_1851_n 0.0103808f $X=7.885 $Y=0.935 $X2=0 $Y2=0
cc_711 N_SET_B_c_823_n N_VGND_c_1851_n 0.00175578f $X=8.31 $Y=1.385 $X2=0 $Y2=0
cc_712 N_SET_B_M1020_g N_VGND_c_1854_n 0.00479212f $X=5.49 $Y=0.8 $X2=0 $Y2=0
cc_713 N_SET_B_c_822_n N_VGND_c_1854_n 0.00436392f $X=7.885 $Y=0.935 $X2=0 $Y2=0
cc_714 N_A_225_74#_M1018_g N_A_1484_62#_M1004_g 0.0609879f $X=7.105 $Y=0.65
+ $X2=0 $Y2=0
cc_715 N_A_225_74#_M1018_g N_A_1484_62#_c_1144_n 0.00359614f $X=7.105 $Y=0.65
+ $X2=0 $Y2=0
cc_716 N_A_225_74#_M1013_g N_A_1321_392#_c_1243_n 0.00673155f $X=6.53 $Y=2.46
+ $X2=0 $Y2=0
cc_717 N_A_225_74#_c_962_n N_A_1321_392#_c_1243_n 0.00551206f $X=7.03 $Y=1.735
+ $X2=0 $Y2=0
cc_718 N_A_225_74#_c_963_n N_A_1321_392#_c_1243_n 0.00174454f $X=6.62 $Y=1.735
+ $X2=0 $Y2=0
cc_719 N_A_225_74#_c_962_n N_A_1321_392#_c_1233_n 0.00171411f $X=7.03 $Y=1.735
+ $X2=0 $Y2=0
cc_720 N_A_225_74#_M1018_g N_A_1321_392#_c_1233_n 0.0138144f $X=7.105 $Y=0.65
+ $X2=0 $Y2=0
cc_721 N_A_225_74#_c_977_n N_A_1321_392#_c_1245_n 3.75949e-19 $X=6.44 $Y=3.15
+ $X2=0 $Y2=0
cc_722 N_A_225_74#_M1013_g N_A_1321_392#_c_1245_n 0.00779479f $X=6.53 $Y=2.46
+ $X2=0 $Y2=0
cc_723 N_A_225_74#_c_962_n N_A_1321_392#_c_1245_n 0.00485374f $X=7.03 $Y=1.735
+ $X2=0 $Y2=0
cc_724 N_A_225_74#_M1018_g N_A_1321_392#_c_1236_n 0.00761503f $X=7.105 $Y=0.65
+ $X2=0 $Y2=0
cc_725 N_A_225_74#_c_962_n N_A_1321_392#_c_1237_n 0.0193954f $X=7.03 $Y=1.735
+ $X2=0 $Y2=0
cc_726 N_A_225_74#_M1018_g N_A_1321_392#_c_1237_n 9.78128e-19 $X=7.105 $Y=0.65
+ $X2=0 $Y2=0
cc_727 N_A_225_74#_M1026_s N_A_27_74#_c_1514_n 0.0126275f $X=1.145 $Y=1.84 $X2=0
+ $Y2=0
cc_728 N_A_225_74#_c_985_n N_A_27_74#_c_1514_n 0.00510828f $X=1.945 $Y=1.805
+ $X2=0 $Y2=0
cc_729 N_A_225_74#_c_987_n N_A_27_74#_c_1514_n 0.0327311f $X=1.455 $Y=1.895
+ $X2=0 $Y2=0
cc_730 N_A_225_74#_c_959_n N_A_27_74#_c_1515_n 0.0149286f $X=1.965 $Y=1.765
+ $X2=0 $Y2=0
cc_731 N_A_225_74#_c_971_n N_A_27_74#_c_1515_n 0.0262812f $X=2.485 $Y=3.075
+ $X2=0 $Y2=0
cc_732 N_A_225_74#_c_966_n N_A_27_74#_c_1515_n 0.00517328f $X=2.41 $Y=1.515
+ $X2=0 $Y2=0
cc_733 N_A_225_74#_c_985_n N_A_27_74#_c_1515_n 0.0265738f $X=1.945 $Y=1.805
+ $X2=0 $Y2=0
cc_734 N_A_225_74#_M1022_g N_A_27_74#_c_1509_n 9.17507e-19 $X=1.915 $Y=0.74
+ $X2=0 $Y2=0
cc_735 N_A_225_74#_c_959_n N_A_27_74#_c_1509_n 0.00117921f $X=1.965 $Y=1.765
+ $X2=0 $Y2=0
cc_736 N_A_225_74#_c_971_n N_A_27_74#_c_1509_n 0.00919077f $X=2.485 $Y=3.075
+ $X2=0 $Y2=0
cc_737 N_A_225_74#_c_960_n N_A_27_74#_c_1509_n 0.00588052f $X=2.91 $Y=1.14 $X2=0
+ $Y2=0
cc_738 N_A_225_74#_M1027_g N_A_27_74#_c_1509_n 0.00249586f $X=2.985 $Y=0.58
+ $X2=0 $Y2=0
cc_739 N_A_225_74#_c_965_n N_A_27_74#_c_1509_n 0.0199619f $X=2.485 $Y=1.14 $X2=0
+ $Y2=0
cc_740 N_A_225_74#_c_985_n N_A_27_74#_c_1509_n 0.0136281f $X=1.945 $Y=1.805
+ $X2=0 $Y2=0
cc_741 N_A_225_74#_c_968_n N_A_27_74#_c_1509_n 0.0265108f $X=2.11 $Y=1.515 $X2=0
+ $Y2=0
cc_742 N_A_225_74#_c_959_n N_A_27_74#_c_1559_n 0.0023413f $X=1.965 $Y=1.765
+ $X2=0 $Y2=0
cc_743 N_A_225_74#_c_985_n N_A_27_74#_c_1559_n 0.0108416f $X=1.945 $Y=1.805
+ $X2=0 $Y2=0
cc_744 N_A_225_74#_c_960_n N_A_27_74#_c_1511_n 0.00616968f $X=2.91 $Y=1.14 $X2=0
+ $Y2=0
cc_745 N_A_225_74#_M1027_g N_A_27_74#_c_1511_n 0.0066603f $X=2.985 $Y=0.58 $X2=0
+ $Y2=0
cc_746 N_A_225_74#_c_965_n N_A_27_74#_c_1511_n 9.04452e-19 $X=2.485 $Y=1.14
+ $X2=0 $Y2=0
cc_747 N_A_225_74#_c_985_n N_VPWR_M1026_d 0.00201531f $X=1.945 $Y=1.805 $X2=0
+ $Y2=0
cc_748 N_A_225_74#_c_959_n N_VPWR_c_1578_n 0.00784696f $X=1.965 $Y=1.765 $X2=0
+ $Y2=0
cc_749 N_A_225_74#_c_971_n N_VPWR_c_1578_n 2.02695e-19 $X=2.485 $Y=3.075 $X2=0
+ $Y2=0
cc_750 N_A_225_74#_c_973_n N_VPWR_c_1578_n 0.0024205f $X=2.56 $Y=3.15 $X2=0
+ $Y2=0
cc_751 N_A_225_74#_c_975_n N_VPWR_c_1579_n 8.25145e-19 $X=3.505 $Y=3.075 $X2=0
+ $Y2=0
cc_752 N_A_225_74#_c_977_n N_VPWR_c_1579_n 0.016318f $X=6.44 $Y=3.15 $X2=0 $Y2=0
cc_753 N_A_225_74#_c_977_n N_VPWR_c_1580_n 0.0229172f $X=6.44 $Y=3.15 $X2=0
+ $Y2=0
cc_754 N_A_225_74#_M1013_g N_VPWR_c_1580_n 0.00416432f $X=6.53 $Y=2.46 $X2=0
+ $Y2=0
cc_755 N_A_225_74#_c_977_n N_VPWR_c_1589_n 0.00416234f $X=6.44 $Y=3.15 $X2=0
+ $Y2=0
cc_756 N_A_225_74#_c_977_n N_VPWR_c_1590_n 0.0365645f $X=6.44 $Y=3.15 $X2=0
+ $Y2=0
cc_757 N_A_225_74#_c_959_n N_VPWR_c_1594_n 0.00413917f $X=1.965 $Y=1.765 $X2=0
+ $Y2=0
cc_758 N_A_225_74#_c_973_n N_VPWR_c_1594_n 0.0363678f $X=2.56 $Y=3.15 $X2=0
+ $Y2=0
cc_759 N_A_225_74#_c_977_n N_VPWR_c_1595_n 0.0241251f $X=6.44 $Y=3.15 $X2=0
+ $Y2=0
cc_760 N_A_225_74#_c_959_n N_VPWR_c_1576_n 0.0081836f $X=1.965 $Y=1.765 $X2=0
+ $Y2=0
cc_761 N_A_225_74#_c_972_n N_VPWR_c_1576_n 0.0201297f $X=3.415 $Y=3.15 $X2=0
+ $Y2=0
cc_762 N_A_225_74#_c_973_n N_VPWR_c_1576_n 0.00600062f $X=2.56 $Y=3.15 $X2=0
+ $Y2=0
cc_763 N_A_225_74#_c_977_n N_VPWR_c_1576_n 0.0938989f $X=6.44 $Y=3.15 $X2=0
+ $Y2=0
cc_764 N_A_225_74#_c_983_n N_VPWR_c_1576_n 0.00441524f $X=3.505 $Y=3.15 $X2=0
+ $Y2=0
cc_765 N_A_225_74#_c_969_n N_VGND_c_1831_n 0.0371671f $X=1.27 $Y=0.515 $X2=0
+ $Y2=0
cc_766 N_A_225_74#_c_969_n N_VGND_c_1832_n 0.0212023f $X=1.27 $Y=0.515 $X2=0
+ $Y2=0
cc_767 N_A_225_74#_M1022_g N_VGND_c_1833_n 0.0115741f $X=1.915 $Y=0.74 $X2=0
+ $Y2=0
cc_768 N_A_225_74#_c_969_n N_VGND_c_1833_n 0.0263763f $X=1.27 $Y=0.515 $X2=0
+ $Y2=0
cc_769 N_A_225_74#_M1022_g N_VGND_c_1843_n 0.00383152f $X=1.915 $Y=0.74 $X2=0
+ $Y2=0
cc_770 N_A_225_74#_M1027_g N_VGND_c_1843_n 0.00278159f $X=2.985 $Y=0.58 $X2=0
+ $Y2=0
cc_771 N_A_225_74#_M1018_g N_VGND_c_1850_n 8.27887e-19 $X=7.105 $Y=0.65 $X2=0
+ $Y2=0
cc_772 N_A_225_74#_M1022_g N_VGND_c_1854_n 0.00762539f $X=1.915 $Y=0.74 $X2=0
+ $Y2=0
cc_773 N_A_225_74#_M1027_g N_VGND_c_1854_n 0.00359882f $X=2.985 $Y=0.58 $X2=0
+ $Y2=0
cc_774 N_A_225_74#_c_969_n N_VGND_c_1854_n 0.0168959f $X=1.27 $Y=0.515 $X2=0
+ $Y2=0
cc_775 N_A_1484_62#_c_1142_n N_A_1321_392#_c_1227_n 0.0241141f $X=9.395 $Y=2.65
+ $X2=0 $Y2=0
cc_776 N_A_1484_62#_c_1139_n N_A_1321_392#_M1002_g 0.0116315f $X=9.12 $Y=0.925
+ $X2=0 $Y2=0
cc_777 N_A_1484_62#_c_1140_n N_A_1321_392#_M1002_g 0.0110008f $X=9.285 $Y=0.65
+ $X2=0 $Y2=0
cc_778 N_A_1484_62#_c_1141_n N_A_1321_392#_M1002_g 0.00495915f $X=9.285 $Y=0.925
+ $X2=0 $Y2=0
cc_779 N_A_1484_62#_c_1142_n N_A_1321_392#_M1002_g 0.0127661f $X=9.395 $Y=2.65
+ $X2=0 $Y2=0
cc_780 N_A_1484_62#_c_1146_n N_A_1321_392#_c_1239_n 0.00469259f $X=9.395
+ $Y=2.815 $X2=0 $Y2=0
cc_781 N_A_1484_62#_c_1142_n N_A_1321_392#_c_1239_n 0.00424448f $X=9.395 $Y=2.65
+ $X2=0 $Y2=0
cc_782 N_A_1484_62#_c_1142_n N_A_1321_392#_c_1229_n 0.0228841f $X=9.395 $Y=2.65
+ $X2=0 $Y2=0
cc_783 N_A_1484_62#_c_1142_n N_A_1321_392#_M1038_g 5.80505e-19 $X=9.395 $Y=2.65
+ $X2=0 $Y2=0
cc_784 N_A_1484_62#_c_1142_n N_A_1321_392#_c_1231_n 0.00645864f $X=9.395 $Y=2.65
+ $X2=0 $Y2=0
cc_785 N_A_1484_62#_c_1145_n N_A_1321_392#_c_1244_n 2.02005e-19 $X=7.745
+ $Y=2.465 $X2=0 $Y2=0
cc_786 N_A_1484_62#_c_1145_n N_A_1321_392#_c_1245_n 9.80133e-19 $X=7.745
+ $Y=2.465 $X2=0 $Y2=0
cc_787 N_A_1484_62#_c_1144_n N_A_1321_392#_c_1246_n 0.00495367f $X=7.745
+ $Y=2.375 $X2=0 $Y2=0
cc_788 N_A_1484_62#_c_1145_n N_A_1321_392#_c_1246_n 0.00529268f $X=7.745
+ $Y=2.465 $X2=0 $Y2=0
cc_789 N_A_1484_62#_c_1138_n N_A_1321_392#_c_1246_n 0.00172307f $X=7.71 $Y=1.49
+ $X2=0 $Y2=0
cc_790 N_A_1484_62#_c_1145_n N_A_1321_392#_c_1247_n 5.30429e-19 $X=7.745
+ $Y=2.465 $X2=0 $Y2=0
cc_791 N_A_1484_62#_c_1142_n N_A_1321_392#_c_1248_n 0.0135416f $X=9.395 $Y=2.65
+ $X2=0 $Y2=0
cc_792 N_A_1484_62#_c_1139_n N_A_1321_392#_c_1234_n 0.0144687f $X=9.12 $Y=0.925
+ $X2=0 $Y2=0
cc_793 N_A_1484_62#_c_1142_n N_A_1321_392#_c_1234_n 0.0696093f $X=9.395 $Y=2.65
+ $X2=0 $Y2=0
cc_794 N_A_1484_62#_c_1139_n N_A_1321_392#_c_1235_n 0.00126969f $X=9.12 $Y=0.925
+ $X2=0 $Y2=0
cc_795 N_A_1484_62#_c_1141_n N_A_1321_392#_c_1235_n 0.00163805f $X=9.285
+ $Y=0.925 $X2=0 $Y2=0
cc_796 N_A_1484_62#_c_1144_n N_A_1321_392#_c_1249_n 0.0025853f $X=7.745 $Y=2.375
+ $X2=0 $Y2=0
cc_797 N_A_1484_62#_c_1145_n N_A_1321_392#_c_1249_n 0.00708296f $X=7.745
+ $Y=2.465 $X2=0 $Y2=0
cc_798 N_A_1484_62#_c_1138_n N_A_1321_392#_c_1249_n 0.00209394f $X=7.71 $Y=1.49
+ $X2=0 $Y2=0
cc_799 N_A_1484_62#_c_1143_n N_A_1321_392#_c_1249_n 5.89701e-19 $X=7.745 $Y=1.49
+ $X2=0 $Y2=0
cc_800 N_A_1484_62#_c_1140_n N_A_1940_74#_c_1400_n 0.0282823f $X=9.285 $Y=0.65
+ $X2=0 $Y2=0
cc_801 N_A_1484_62#_c_1141_n N_A_1940_74#_c_1400_n 0.0121618f $X=9.285 $Y=0.925
+ $X2=0 $Y2=0
cc_802 N_A_1484_62#_c_1142_n N_A_1940_74#_c_1400_n 0.0198356f $X=9.395 $Y=2.65
+ $X2=0 $Y2=0
cc_803 N_A_1484_62#_c_1142_n N_A_1940_74#_c_1402_n 0.0105853f $X=9.395 $Y=2.65
+ $X2=0 $Y2=0
cc_804 N_A_1484_62#_c_1145_n N_VPWR_c_1581_n 0.00538254f $X=7.745 $Y=2.465 $X2=0
+ $Y2=0
cc_805 N_A_1484_62#_c_1146_n N_VPWR_c_1582_n 0.0221564f $X=9.395 $Y=2.815 $X2=0
+ $Y2=0
cc_806 N_A_1484_62#_c_1146_n N_VPWR_c_1583_n 0.0244397f $X=9.395 $Y=2.815 $X2=0
+ $Y2=0
cc_807 N_A_1484_62#_c_1142_n N_VPWR_c_1583_n 0.0427482f $X=9.395 $Y=2.65 $X2=0
+ $Y2=0
cc_808 N_A_1484_62#_c_1145_n N_VPWR_c_1595_n 0.00423156f $X=7.745 $Y=2.465 $X2=0
+ $Y2=0
cc_809 N_A_1484_62#_c_1146_n N_VPWR_c_1597_n 0.0142446f $X=9.395 $Y=2.815 $X2=0
+ $Y2=0
cc_810 N_A_1484_62#_c_1145_n N_VPWR_c_1576_n 0.00452425f $X=7.745 $Y=2.465 $X2=0
+ $Y2=0
cc_811 N_A_1484_62#_c_1146_n N_VPWR_c_1576_n 0.0119122f $X=9.395 $Y=2.815 $X2=0
+ $Y2=0
cc_812 N_A_1484_62#_c_1139_n N_VGND_M1005_d 0.0100699f $X=9.12 $Y=0.925 $X2=0
+ $Y2=0
cc_813 N_A_1484_62#_c_1140_n N_VGND_c_1844_n 0.0112889f $X=9.285 $Y=0.65 $X2=0
+ $Y2=0
cc_814 N_A_1484_62#_M1004_g N_VGND_c_1850_n 0.00527445f $X=7.495 $Y=0.65 $X2=0
+ $Y2=0
cc_815 N_A_1484_62#_M1004_g N_VGND_c_1851_n 0.00104583f $X=7.495 $Y=0.65 $X2=0
+ $Y2=0
cc_816 N_A_1484_62#_c_1139_n N_VGND_c_1851_n 0.0747503f $X=9.12 $Y=0.925 $X2=0
+ $Y2=0
cc_817 N_A_1484_62#_c_1140_n N_VGND_c_1851_n 0.0102732f $X=9.285 $Y=0.65 $X2=0
+ $Y2=0
cc_818 N_A_1484_62#_M1004_g N_VGND_c_1854_n 0.00523671f $X=7.495 $Y=0.65 $X2=0
+ $Y2=0
cc_819 N_A_1484_62#_c_1139_n N_VGND_c_1854_n 0.010553f $X=9.12 $Y=0.925 $X2=0
+ $Y2=0
cc_820 N_A_1484_62#_c_1155_n N_VGND_c_1854_n 0.0126596f $X=7.875 $Y=0.925 $X2=0
+ $Y2=0
cc_821 N_A_1484_62#_c_1140_n N_VGND_c_1854_n 0.0115369f $X=9.285 $Y=0.65 $X2=0
+ $Y2=0
cc_822 N_A_1484_62#_c_1155_n A_1514_88# 0.00299242f $X=7.875 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_823 N_A_1321_392#_M1038_g N_A_1940_74#_c_1393_n 0.0119421f $X=10.13 $Y=0.74
+ $X2=0 $Y2=0
cc_824 N_A_1321_392#_c_1231_n N_A_1940_74#_c_1395_n 0.0119421f $X=10.145
+ $Y=1.765 $X2=0 $Y2=0
cc_825 N_A_1321_392#_c_1232_n N_A_1940_74#_c_1395_n 0.00720145f $X=10.52 $Y=1.69
+ $X2=0 $Y2=0
cc_826 N_A_1321_392#_c_1242_n N_A_1940_74#_c_1405_n 0.014112f $X=10.595 $Y=1.765
+ $X2=0 $Y2=0
cc_827 N_A_1321_392#_c_1232_n N_A_1940_74#_c_1398_n 0.00645298f $X=10.52 $Y=1.69
+ $X2=0 $Y2=0
cc_828 N_A_1321_392#_M1002_g N_A_1940_74#_c_1400_n 0.00323395f $X=9.07 $Y=0.65
+ $X2=0 $Y2=0
cc_829 N_A_1321_392#_M1038_g N_A_1940_74#_c_1400_n 0.0230336f $X=10.13 $Y=0.74
+ $X2=0 $Y2=0
cc_830 N_A_1321_392#_c_1229_n N_A_1940_74#_c_1401_n 0.00212027f $X=10.055
+ $Y=1.492 $X2=0 $Y2=0
cc_831 N_A_1321_392#_M1038_g N_A_1940_74#_c_1401_n 0.00759579f $X=10.13 $Y=0.74
+ $X2=0 $Y2=0
cc_832 N_A_1321_392#_c_1231_n N_A_1940_74#_c_1401_n 0.00819331f $X=10.145
+ $Y=1.765 $X2=0 $Y2=0
cc_833 N_A_1321_392#_c_1229_n N_A_1940_74#_c_1402_n 0.0195173f $X=10.055
+ $Y=1.492 $X2=0 $Y2=0
cc_834 N_A_1321_392#_c_1231_n N_A_1940_74#_c_1410_n 0.0200748f $X=10.145
+ $Y=1.765 $X2=0 $Y2=0
cc_835 N_A_1321_392#_c_1232_n N_A_1940_74#_c_1410_n 0.00823448f $X=10.52 $Y=1.69
+ $X2=0 $Y2=0
cc_836 N_A_1321_392#_c_1242_n N_A_1940_74#_c_1410_n 0.0132933f $X=10.595
+ $Y=1.765 $X2=0 $Y2=0
cc_837 N_A_1321_392#_c_1232_n N_A_1940_74#_c_1403_n 0.00965439f $X=10.52 $Y=1.69
+ $X2=0 $Y2=0
cc_838 N_A_1321_392#_M1038_g N_A_1940_74#_c_1404_n 6.82259e-19 $X=10.13 $Y=0.74
+ $X2=0 $Y2=0
cc_839 N_A_1321_392#_c_1231_n N_A_1940_74#_c_1404_n 0.0145244f $X=10.145
+ $Y=1.765 $X2=0 $Y2=0
cc_840 N_A_1321_392#_c_1232_n N_A_1940_74#_c_1404_n 0.00730677f $X=10.52 $Y=1.69
+ $X2=0 $Y2=0
cc_841 N_A_1321_392#_c_1245_n N_VPWR_c_1580_n 0.0083277f $X=7.265 $Y=2.565 $X2=0
+ $Y2=0
cc_842 N_A_1321_392#_c_1245_n N_VPWR_c_1581_n 0.0092631f $X=7.265 $Y=2.565 $X2=0
+ $Y2=0
cc_843 N_A_1321_392#_c_1246_n N_VPWR_c_1581_n 0.0135931f $X=8.255 $Y=2.395 $X2=0
+ $Y2=0
cc_844 N_A_1321_392#_c_1247_n N_VPWR_c_1581_n 0.0215225f $X=8.42 $Y=2.75 $X2=0
+ $Y2=0
cc_845 N_A_1321_392#_c_1239_n N_VPWR_c_1582_n 0.00741173f $X=9.17 $Y=2.465 $X2=0
+ $Y2=0
cc_846 N_A_1321_392#_c_1247_n N_VPWR_c_1582_n 0.0244396f $X=8.42 $Y=2.75 $X2=0
+ $Y2=0
cc_847 N_A_1321_392#_c_1248_n N_VPWR_c_1582_n 0.0223194f $X=8.78 $Y=2.395 $X2=0
+ $Y2=0
cc_848 N_A_1321_392#_c_1239_n N_VPWR_c_1583_n 0.00323899f $X=9.17 $Y=2.465 $X2=0
+ $Y2=0
cc_849 N_A_1321_392#_c_1229_n N_VPWR_c_1583_n 0.00599962f $X=10.055 $Y=1.492
+ $X2=0 $Y2=0
cc_850 N_A_1321_392#_c_1231_n N_VPWR_c_1583_n 0.0112442f $X=10.145 $Y=1.765
+ $X2=0 $Y2=0
cc_851 N_A_1321_392#_c_1231_n N_VPWR_c_1584_n 0.00393873f $X=10.145 $Y=1.765
+ $X2=0 $Y2=0
cc_852 N_A_1321_392#_c_1242_n N_VPWR_c_1584_n 0.00393873f $X=10.595 $Y=1.765
+ $X2=0 $Y2=0
cc_853 N_A_1321_392#_c_1242_n N_VPWR_c_1585_n 0.00785728f $X=10.595 $Y=1.765
+ $X2=0 $Y2=0
cc_854 N_A_1321_392#_c_1244_n N_VPWR_c_1595_n 0.00387501f $X=7.545 $Y=2.565
+ $X2=0 $Y2=0
cc_855 N_A_1321_392#_c_1245_n N_VPWR_c_1595_n 0.0294395f $X=7.265 $Y=2.565 $X2=0
+ $Y2=0
cc_856 N_A_1321_392#_c_1249_n N_VPWR_c_1595_n 0.00229466f $X=7.63 $Y=2.395 $X2=0
+ $Y2=0
cc_857 N_A_1321_392#_c_1247_n N_VPWR_c_1596_n 0.0145781f $X=8.42 $Y=2.75 $X2=0
+ $Y2=0
cc_858 N_A_1321_392#_c_1239_n N_VPWR_c_1597_n 0.00445602f $X=9.17 $Y=2.465 $X2=0
+ $Y2=0
cc_859 N_A_1321_392#_c_1239_n N_VPWR_c_1576_n 0.00822944f $X=9.17 $Y=2.465 $X2=0
+ $Y2=0
cc_860 N_A_1321_392#_c_1231_n N_VPWR_c_1576_n 0.00462577f $X=10.145 $Y=1.765
+ $X2=0 $Y2=0
cc_861 N_A_1321_392#_c_1242_n N_VPWR_c_1576_n 0.00462577f $X=10.595 $Y=1.765
+ $X2=0 $Y2=0
cc_862 N_A_1321_392#_c_1244_n N_VPWR_c_1576_n 0.00704588f $X=7.545 $Y=2.565
+ $X2=0 $Y2=0
cc_863 N_A_1321_392#_c_1245_n N_VPWR_c_1576_n 0.0244971f $X=7.265 $Y=2.565 $X2=0
+ $Y2=0
cc_864 N_A_1321_392#_c_1246_n N_VPWR_c_1576_n 0.0115465f $X=8.255 $Y=2.395 $X2=0
+ $Y2=0
cc_865 N_A_1321_392#_c_1247_n N_VPWR_c_1576_n 0.0120405f $X=8.42 $Y=2.75 $X2=0
+ $Y2=0
cc_866 N_A_1321_392#_c_1248_n N_VPWR_c_1576_n 0.0105894f $X=8.78 $Y=2.395 $X2=0
+ $Y2=0
cc_867 N_A_1321_392#_c_1249_n N_VPWR_c_1576_n 0.00455301f $X=7.63 $Y=2.395 $X2=0
+ $Y2=0
cc_868 N_A_1321_392#_c_1244_n A_1480_508# 0.0018712f $X=7.545 $Y=2.565 $X2=-0.19
+ $Y2=-0.245
cc_869 N_A_1321_392#_c_1249_n A_1480_508# 0.00151742f $X=7.63 $Y=2.395 $X2=-0.19
+ $Y2=-0.245
cc_870 N_A_1321_392#_M1038_g N_VGND_c_1836_n 0.0163444f $X=10.13 $Y=0.74 $X2=0
+ $Y2=0
cc_871 N_A_1321_392#_c_1231_n N_VGND_c_1836_n 0.0012784f $X=10.145 $Y=1.765
+ $X2=0 $Y2=0
cc_872 N_A_1321_392#_M1002_g N_VGND_c_1844_n 0.00504315f $X=9.07 $Y=0.65 $X2=0
+ $Y2=0
cc_873 N_A_1321_392#_M1038_g N_VGND_c_1844_n 0.00383152f $X=10.13 $Y=0.74 $X2=0
+ $Y2=0
cc_874 N_A_1321_392#_M1002_g N_VGND_c_1851_n 0.0100857f $X=9.07 $Y=0.65 $X2=0
+ $Y2=0
cc_875 N_A_1321_392#_M1002_g N_VGND_c_1854_n 0.00523671f $X=9.07 $Y=0.65 $X2=0
+ $Y2=0
cc_876 N_A_1321_392#_M1038_g N_VGND_c_1854_n 0.00762539f $X=10.13 $Y=0.74 $X2=0
+ $Y2=0
cc_877 N_A_1940_74#_c_1402_n N_VPWR_c_1583_n 0.0134388f $X=10.01 $Y=1.405 $X2=0
+ $Y2=0
cc_878 N_A_1940_74#_c_1410_n N_VPWR_c_1583_n 0.059064f $X=10.37 $Y=1.985 $X2=0
+ $Y2=0
cc_879 N_A_1940_74#_c_1410_n N_VPWR_c_1584_n 0.00664674f $X=10.37 $Y=1.985 $X2=0
+ $Y2=0
cc_880 N_A_1940_74#_c_1394_n N_VPWR_c_1585_n 0.00111964f $X=10.985 $Y=1.3 $X2=0
+ $Y2=0
cc_881 N_A_1940_74#_c_1405_n N_VPWR_c_1585_n 0.0041061f $X=11.115 $Y=1.765 $X2=0
+ $Y2=0
cc_882 N_A_1940_74#_c_1398_n N_VPWR_c_1585_n 5.17557e-19 $X=12.395 $Y=1.32 $X2=0
+ $Y2=0
cc_883 N_A_1940_74#_c_1410_n N_VPWR_c_1585_n 0.0316306f $X=10.37 $Y=1.985 $X2=0
+ $Y2=0
cc_884 N_A_1940_74#_c_1403_n N_VPWR_c_1585_n 0.0245135f $X=11.83 $Y=1.485 $X2=0
+ $Y2=0
cc_885 N_A_1940_74#_c_1405_n N_VPWR_c_1586_n 5.50173e-19 $X=11.115 $Y=1.765
+ $X2=0 $Y2=0
cc_886 N_A_1940_74#_c_1406_n N_VPWR_c_1586_n 0.0121556f $X=11.565 $Y=1.765 $X2=0
+ $Y2=0
cc_887 N_A_1940_74#_c_1407_n N_VPWR_c_1586_n 0.0120719f $X=12.015 $Y=1.765 $X2=0
+ $Y2=0
cc_888 N_A_1940_74#_c_1409_n N_VPWR_c_1586_n 5.16933e-19 $X=12.465 $Y=1.765
+ $X2=0 $Y2=0
cc_889 N_A_1940_74#_c_1407_n N_VPWR_c_1588_n 4.98648e-19 $X=12.015 $Y=1.765
+ $X2=0 $Y2=0
cc_890 N_A_1940_74#_c_1409_n N_VPWR_c_1588_n 0.0116621f $X=12.465 $Y=1.765 $X2=0
+ $Y2=0
cc_891 N_A_1940_74#_c_1405_n N_VPWR_c_1598_n 0.00445602f $X=11.115 $Y=1.765
+ $X2=0 $Y2=0
cc_892 N_A_1940_74#_c_1406_n N_VPWR_c_1598_n 0.00413917f $X=11.565 $Y=1.765
+ $X2=0 $Y2=0
cc_893 N_A_1940_74#_c_1407_n N_VPWR_c_1599_n 0.00413917f $X=12.015 $Y=1.765
+ $X2=0 $Y2=0
cc_894 N_A_1940_74#_c_1409_n N_VPWR_c_1599_n 0.00413917f $X=12.465 $Y=1.765
+ $X2=0 $Y2=0
cc_895 N_A_1940_74#_c_1405_n N_VPWR_c_1576_n 0.00861719f $X=11.115 $Y=1.765
+ $X2=0 $Y2=0
cc_896 N_A_1940_74#_c_1406_n N_VPWR_c_1576_n 0.00817726f $X=11.565 $Y=1.765
+ $X2=0 $Y2=0
cc_897 N_A_1940_74#_c_1407_n N_VPWR_c_1576_n 0.00817726f $X=12.015 $Y=1.765
+ $X2=0 $Y2=0
cc_898 N_A_1940_74#_c_1409_n N_VPWR_c_1576_n 0.00817726f $X=12.465 $Y=1.765
+ $X2=0 $Y2=0
cc_899 N_A_1940_74#_c_1410_n N_VPWR_c_1576_n 0.00995652f $X=10.37 $Y=1.985 $X2=0
+ $Y2=0
cc_900 N_A_1940_74#_c_1393_n N_Q_c_1758_n 0.00761489f $X=10.63 $Y=1.225 $X2=0
+ $Y2=0
cc_901 N_A_1940_74#_c_1396_n N_Q_c_1758_n 0.0137392f $X=11.06 $Y=1.225 $X2=0
+ $Y2=0
cc_902 N_A_1940_74#_c_1396_n N_Q_c_1759_n 0.0127216f $X=11.06 $Y=1.225 $X2=0
+ $Y2=0
cc_903 N_A_1940_74#_c_1397_n N_Q_c_1759_n 0.0150954f $X=11.92 $Y=1.225 $X2=0
+ $Y2=0
cc_904 N_A_1940_74#_c_1398_n N_Q_c_1759_n 0.0145022f $X=12.395 $Y=1.32 $X2=0
+ $Y2=0
cc_905 N_A_1940_74#_c_1403_n N_Q_c_1759_n 0.072964f $X=11.83 $Y=1.485 $X2=0
+ $Y2=0
cc_906 N_A_1940_74#_c_1393_n N_Q_c_1760_n 0.00276819f $X=10.63 $Y=1.225 $X2=0
+ $Y2=0
cc_907 N_A_1940_74#_c_1394_n N_Q_c_1760_n 0.00224597f $X=10.985 $Y=1.3 $X2=0
+ $Y2=0
cc_908 N_A_1940_74#_c_1396_n N_Q_c_1760_n 0.00121617f $X=11.06 $Y=1.225 $X2=0
+ $Y2=0
cc_909 N_A_1940_74#_c_1400_n N_Q_c_1760_n 5.79493e-19 $X=9.845 $Y=0.515 $X2=0
+ $Y2=0
cc_910 N_A_1940_74#_c_1403_n N_Q_c_1760_n 0.0275317f $X=11.83 $Y=1.485 $X2=0
+ $Y2=0
cc_911 N_A_1940_74#_c_1405_n N_Q_c_1765_n 0.00295734f $X=11.115 $Y=1.765 $X2=0
+ $Y2=0
cc_912 N_A_1940_74#_c_1398_n N_Q_c_1765_n 0.00664878f $X=12.395 $Y=1.32 $X2=0
+ $Y2=0
cc_913 N_A_1940_74#_c_1403_n N_Q_c_1765_n 0.0235455f $X=11.83 $Y=1.485 $X2=0
+ $Y2=0
cc_914 N_A_1940_74#_c_1405_n N_Q_c_1766_n 0.00951605f $X=11.115 $Y=1.765 $X2=0
+ $Y2=0
cc_915 N_A_1940_74#_c_1406_n N_Q_c_1766_n 3.88029e-19 $X=11.565 $Y=1.765 $X2=0
+ $Y2=0
cc_916 N_A_1940_74#_c_1397_n N_Q_c_1761_n 4.78514e-19 $X=11.92 $Y=1.225 $X2=0
+ $Y2=0
cc_917 N_A_1940_74#_M1036_g N_Q_c_1761_n 0.0133757f $X=12.395 $Y=0.74 $X2=0
+ $Y2=0
cc_918 N_A_1940_74#_c_1407_n N_Q_c_1767_n 3.85296e-19 $X=12.015 $Y=1.765 $X2=0
+ $Y2=0
cc_919 N_A_1940_74#_c_1409_n N_Q_c_1767_n 3.85296e-19 $X=12.465 $Y=1.765 $X2=0
+ $Y2=0
cc_920 N_A_1940_74#_c_1398_n N_Q_c_1762_n 0.00207582f $X=12.395 $Y=1.32 $X2=0
+ $Y2=0
cc_921 N_A_1940_74#_M1036_g N_Q_c_1762_n 0.0144108f $X=12.395 $Y=0.74 $X2=0
+ $Y2=0
cc_922 N_A_1940_74#_c_1398_n N_Q_c_1763_n 0.00441672f $X=12.395 $Y=1.32 $X2=0
+ $Y2=0
cc_923 N_A_1940_74#_M1036_g N_Q_c_1763_n 0.00156147f $X=12.395 $Y=0.74 $X2=0
+ $Y2=0
cc_924 N_A_1940_74#_c_1398_n Q 0.0102248f $X=12.395 $Y=1.32 $X2=0 $Y2=0
cc_925 N_A_1940_74#_M1036_g Q 0.0121215f $X=12.395 $Y=0.74 $X2=0 $Y2=0
cc_926 N_A_1940_74#_c_1409_n Q 0.0021695f $X=12.465 $Y=1.765 $X2=0 $Y2=0
cc_927 N_A_1940_74#_c_1403_n Q 0.0100186f $X=11.83 $Y=1.485 $X2=0 $Y2=0
cc_928 N_A_1940_74#_c_1398_n Q 0.00104631f $X=12.395 $Y=1.32 $X2=0 $Y2=0
cc_929 N_A_1940_74#_c_1409_n Q 0.0219927f $X=12.465 $Y=1.765 $X2=0 $Y2=0
cc_930 N_A_1940_74#_c_1406_n N_Q_c_1770_n 0.0156734f $X=11.565 $Y=1.765 $X2=0
+ $Y2=0
cc_931 N_A_1940_74#_c_1407_n N_Q_c_1770_n 0.0170352f $X=12.015 $Y=1.765 $X2=0
+ $Y2=0
cc_932 N_A_1940_74#_c_1398_n N_Q_c_1770_n 0.0174638f $X=12.395 $Y=1.32 $X2=0
+ $Y2=0
cc_933 N_A_1940_74#_c_1403_n N_Q_c_1770_n 0.0410851f $X=11.83 $Y=1.485 $X2=0
+ $Y2=0
cc_934 N_A_1940_74#_c_1393_n N_VGND_c_1836_n 0.00590268f $X=10.63 $Y=1.225 $X2=0
+ $Y2=0
cc_935 N_A_1940_74#_c_1400_n N_VGND_c_1836_n 0.0308485f $X=9.845 $Y=0.515 $X2=0
+ $Y2=0
cc_936 N_A_1940_74#_c_1401_n N_VGND_c_1836_n 0.00164036f $X=10.205 $Y=1.405
+ $X2=0 $Y2=0
cc_937 N_A_1940_74#_c_1404_n N_VGND_c_1836_n 0.0263154f $X=10.37 $Y=1.485 $X2=0
+ $Y2=0
cc_938 N_A_1940_74#_c_1396_n N_VGND_c_1837_n 0.00322722f $X=11.06 $Y=1.225 $X2=0
+ $Y2=0
cc_939 N_A_1940_74#_c_1397_n N_VGND_c_1837_n 0.00352244f $X=11.92 $Y=1.225 $X2=0
+ $Y2=0
cc_940 N_A_1940_74#_M1036_g N_VGND_c_1839_n 0.0122304f $X=12.395 $Y=0.74 $X2=0
+ $Y2=0
cc_941 N_A_1940_74#_c_1400_n N_VGND_c_1844_n 0.0146357f $X=9.845 $Y=0.515 $X2=0
+ $Y2=0
cc_942 N_A_1940_74#_c_1393_n N_VGND_c_1845_n 0.00434272f $X=10.63 $Y=1.225 $X2=0
+ $Y2=0
cc_943 N_A_1940_74#_c_1396_n N_VGND_c_1845_n 0.00434272f $X=11.06 $Y=1.225 $X2=0
+ $Y2=0
cc_944 N_A_1940_74#_c_1397_n N_VGND_c_1846_n 0.00460063f $X=11.92 $Y=1.225 $X2=0
+ $Y2=0
cc_945 N_A_1940_74#_M1036_g N_VGND_c_1846_n 0.00434272f $X=12.395 $Y=0.74 $X2=0
+ $Y2=0
cc_946 N_A_1940_74#_c_1393_n N_VGND_c_1854_n 0.00820772f $X=10.63 $Y=1.225 $X2=0
+ $Y2=0
cc_947 N_A_1940_74#_c_1396_n N_VGND_c_1854_n 0.00823001f $X=11.06 $Y=1.225 $X2=0
+ $Y2=0
cc_948 N_A_1940_74#_c_1397_n N_VGND_c_1854_n 0.00910475f $X=11.92 $Y=1.225 $X2=0
+ $Y2=0
cc_949 N_A_1940_74#_M1036_g N_VGND_c_1854_n 0.00824368f $X=12.395 $Y=0.74 $X2=0
+ $Y2=0
cc_950 N_A_1940_74#_c_1400_n N_VGND_c_1854_n 0.0121141f $X=9.845 $Y=0.515 $X2=0
+ $Y2=0
cc_951 N_A_27_74#_c_1515_n N_VPWR_M1026_d 0.00138464f $X=2.445 $Y=2.155 $X2=0
+ $Y2=0
cc_952 N_A_27_74#_c_1559_n N_VPWR_M1026_d 0.00591605f $X=1.71 $Y=2.155 $X2=0
+ $Y2=0
cc_953 N_A_27_74#_c_1513_n N_VPWR_c_1577_n 0.0255089f $X=0.28 $Y=2.73 $X2=0
+ $Y2=0
cc_954 N_A_27_74#_c_1514_n N_VPWR_c_1577_n 0.0244079f $X=1.625 $Y=2.325 $X2=0
+ $Y2=0
cc_955 N_A_27_74#_c_1514_n N_VPWR_c_1578_n 0.00102433f $X=1.625 $Y=2.325 $X2=0
+ $Y2=0
cc_956 N_A_27_74#_c_1515_n N_VPWR_c_1578_n 0.00243978f $X=2.445 $Y=2.155 $X2=0
+ $Y2=0
cc_957 N_A_27_74#_c_1559_n N_VPWR_c_1578_n 0.0126064f $X=1.71 $Y=2.155 $X2=0
+ $Y2=0
cc_958 N_A_27_74#_c_1513_n N_VPWR_c_1592_n 0.0102563f $X=0.28 $Y=2.73 $X2=0
+ $Y2=0
cc_959 N_A_27_74#_c_1513_n N_VPWR_c_1576_n 0.0090542f $X=0.28 $Y=2.73 $X2=0
+ $Y2=0
cc_960 N_A_27_74#_c_1507_n N_VGND_c_1831_n 0.0172562f $X=0.28 $Y=0.58 $X2=0
+ $Y2=0
cc_961 N_A_27_74#_c_1507_n N_VGND_c_1842_n 0.0109681f $X=0.28 $Y=0.58 $X2=0
+ $Y2=0
cc_962 N_A_27_74#_c_1507_n N_VGND_c_1854_n 0.00912188f $X=0.28 $Y=0.58 $X2=0
+ $Y2=0
cc_963 N_VPWR_c_1585_n N_Q_c_1765_n 0.0117266f $X=10.89 $Y=1.985 $X2=0 $Y2=0
cc_964 N_VPWR_c_1585_n N_Q_c_1766_n 0.0336653f $X=10.89 $Y=1.985 $X2=0 $Y2=0
cc_965 N_VPWR_c_1586_n N_Q_c_1766_n 0.0281624f $X=11.79 $Y=2.335 $X2=0 $Y2=0
cc_966 N_VPWR_c_1598_n N_Q_c_1766_n 0.0123628f $X=11.625 $Y=3.33 $X2=0 $Y2=0
cc_967 N_VPWR_c_1576_n N_Q_c_1766_n 0.0101999f $X=12.72 $Y=3.33 $X2=0 $Y2=0
cc_968 N_VPWR_c_1586_n N_Q_c_1767_n 0.0281398f $X=11.79 $Y=2.335 $X2=0 $Y2=0
cc_969 N_VPWR_c_1588_n N_Q_c_1767_n 0.0255132f $X=12.69 $Y=2.405 $X2=0 $Y2=0
cc_970 N_VPWR_c_1599_n N_Q_c_1767_n 0.0101736f $X=12.525 $Y=3.33 $X2=0 $Y2=0
cc_971 N_VPWR_c_1576_n N_Q_c_1767_n 0.0084208f $X=12.72 $Y=3.33 $X2=0 $Y2=0
cc_972 N_VPWR_M1025_d Q 0.00426951f $X=12.54 $Y=1.84 $X2=0 $Y2=0
cc_973 N_VPWR_c_1588_n Q 0.0213356f $X=12.69 $Y=2.405 $X2=0 $Y2=0
cc_974 N_VPWR_M1015_d N_Q_c_1770_n 0.00200327f $X=11.64 $Y=1.84 $X2=0 $Y2=0
cc_975 N_VPWR_c_1586_n N_Q_c_1770_n 0.0176914f $X=11.79 $Y=2.335 $X2=0 $Y2=0
cc_976 N_Q_c_1759_n N_VGND_M1009_s 0.0089885f $X=12.015 $Y=1.065 $X2=0 $Y2=0
cc_977 N_Q_c_1762_n N_VGND_M1036_s 0.00451232f $X=12.605 $Y=1.065 $X2=0 $Y2=0
cc_978 N_Q_c_1758_n N_VGND_c_1836_n 0.0243921f $X=10.845 $Y=0.515 $X2=0 $Y2=0
cc_979 N_Q_c_1760_n N_VGND_c_1836_n 0.00711243f $X=11.01 $Y=1.065 $X2=0 $Y2=0
cc_980 N_Q_c_1758_n N_VGND_c_1837_n 0.0177638f $X=10.845 $Y=0.515 $X2=0 $Y2=0
cc_981 N_Q_c_1759_n N_VGND_c_1837_n 0.0464602f $X=12.015 $Y=1.065 $X2=0 $Y2=0
cc_982 N_Q_c_1761_n N_VGND_c_1837_n 0.0183183f $X=12.18 $Y=0.515 $X2=0 $Y2=0
cc_983 N_Q_c_1761_n N_VGND_c_1839_n 0.0180508f $X=12.18 $Y=0.515 $X2=0 $Y2=0
cc_984 N_Q_c_1762_n N_VGND_c_1839_n 0.0270821f $X=12.605 $Y=1.065 $X2=0 $Y2=0
cc_985 N_Q_c_1758_n N_VGND_c_1845_n 0.0144922f $X=10.845 $Y=0.515 $X2=0 $Y2=0
cc_986 N_Q_c_1761_n N_VGND_c_1846_n 0.0145639f $X=12.18 $Y=0.515 $X2=0 $Y2=0
cc_987 N_Q_c_1758_n N_VGND_c_1854_n 0.0118826f $X=10.845 $Y=0.515 $X2=0 $Y2=0
cc_988 N_Q_c_1761_n N_VGND_c_1854_n 0.0119984f $X=12.18 $Y=0.515 $X2=0 $Y2=0
