* NGSPICE file created from sky130_fd_sc_ls__and2b_2.ext - technology: sky130A

.subckt sky130_fd_sc_ls__and2b_2 A_N B VGND VNB VPB VPWR X
M1000 a_505_74# B VGND VNB nshort w=740000u l=150000u
+  ad=1.776e+11p pd=1.96e+06u as=8.742e+11p ps=5.41e+06u
M1001 a_198_48# a_27_74# a_505_74# VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1002 VPWR a_27_74# a_198_48# VPB phighvt w=1e+06u l=150000u
+  ad=1.53365e+12p pd=9.39e+06u as=3e+11p ps=2.6e+06u
M1003 VGND a_198_48# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.072e+11p ps=2.04e+06u
M1004 X a_198_48# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=0p ps=0u
M1005 VPWR A_N a_27_74# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=2.478e+11p ps=2.27e+06u
M1006 VPWR a_198_48# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND A_N a_27_74# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1008 X a_198_48# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_198_48# B VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

