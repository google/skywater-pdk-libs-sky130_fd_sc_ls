* File: sky130_fd_sc_ls__nor4_2.pex.spice
* Created: Fri Aug 28 13:39:56 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__NOR4_2%C 2 3 5 6 8 11 16 17 21 22 31 34 40
c72 16 0 1.10961e-19 $X=0.535 $Y=1.335
r73 32 34 0.751593 $w=2.28e-07 $l=1.5e-08 $layer=LI1_cond $X=1.68 $Y=1.65
+ $X2=1.68 $Y2=1.665
r74 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.91
+ $Y=1.485 $X2=1.91 $Y2=1.485
r75 21 31 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=1.68 $Y=1.485
+ $X2=1.91 $Y2=1.485
r76 21 32 2.85155 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=1.68 $Y=1.485
+ $X2=1.68 $Y2=1.65
r77 21 40 6.38036 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=1.68 $Y=1.485
+ $X2=1.565 $Y2=1.485
r78 21 22 16.7856 $w=2.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.68 $Y=1.7
+ $X2=1.68 $Y2=2.035
r79 21 34 1.75372 $w=2.28e-07 $l=3.5e-08 $layer=LI1_cond $X=1.68 $Y=1.7 $X2=1.68
+ $Y2=1.665
r80 17 28 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.535 $Y=1.335
+ $X2=0.535 $Y2=1.5
r81 16 19 3.14303 $w=2.73e-07 $l=7.5e-08 $layer=LI1_cond $X=0.562 $Y=1.335
+ $X2=0.562 $Y2=1.41
r82 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.535
+ $Y=1.335 $X2=0.535 $Y2=1.335
r83 14 19 3.21752 $w=1.8e-07 $l=1.38e-07 $layer=LI1_cond $X=0.7 $Y=1.41
+ $X2=0.562 $Y2=1.41
r84 14 40 53.298 $w=1.78e-07 $l=8.65e-07 $layer=LI1_cond $X=0.7 $Y=1.41
+ $X2=1.565 $Y2=1.41
r85 9 30 38.6072 $w=2.91e-07 $l=1.74714e-07 $layer=POLY_cond $X=1.93 $Y=1.32
+ $X2=1.91 $Y2=1.485
r86 9 11 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.93 $Y=1.32 $X2=1.93
+ $Y2=0.74
r87 6 30 57.6553 $w=2.91e-07 $l=2.87402e-07 $layer=POLY_cond $X=1.895 $Y=1.765
+ $X2=1.91 $Y2=1.485
r88 6 8 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.895 $Y=1.765
+ $X2=1.895 $Y2=2.4
r89 3 5 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.4
r90 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.505 $Y=1.675 $X2=0.505
+ $Y2=1.765
r91 2 28 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=0.505 $Y=1.675
+ $X2=0.505 $Y2=1.5
.ends

.subckt PM_SKY130_FD_SC_LS__NOR4_2%D 1 3 5 7 8 9 10 12 13 15 20 23
c61 23 0 6.36756e-20 $X=0.27 $Y=0.495
c62 8 0 1.10961e-19 $X=1.445 $Y=1.52
r63 20 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=0.495 $X2=0.27 $Y2=0.495
r64 16 17 1.89267 $w=3.82e-07 $l=1.5e-08 $layer=POLY_cond $X=0.97 $Y=1.475
+ $X2=0.985 $Y2=1.475
r65 13 19 24.74 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=1.46 $Y=1.185 $X2=1.46
+ $Y2=1.475
r66 13 15 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.46 $Y=1.185
+ $X2=1.46 $Y2=0.74
r67 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.445 $Y=1.765
+ $X2=1.445 $Y2=2.4
r68 9 10 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.445 $Y=1.675
+ $X2=1.445 $Y2=1.765
r69 8 19 1.89267 $w=3.82e-07 $l=1.5e-08 $layer=POLY_cond $X=1.445 $Y=1.475
+ $X2=1.46 $Y2=1.475
r70 8 17 58.0419 $w=3.82e-07 $l=4.6e-07 $layer=POLY_cond $X=1.445 $Y=1.475
+ $X2=0.985 $Y2=1.475
r71 8 9 60.25 $w=1.8e-07 $l=1.55e-07 $layer=POLY_cond $X=1.445 $Y=1.52 $X2=1.445
+ $Y2=1.675
r72 7 17 24.74 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=0.985 $Y=1.185
+ $X2=0.985 $Y2=1.475
r73 6 7 153.83 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=0.985 $Y=0.885 $X2=0.985
+ $Y2=1.185
r74 3 16 24.74 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=0.97 $Y=1.765 $X2=0.97
+ $Y2=1.475
r75 3 5 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.97 $Y=1.765
+ $X2=0.97 $Y2=2.4
r76 2 23 59.0778 $w=2.57e-07 $l=3.88844e-07 $layer=POLY_cond $X=0.435 $Y=0.81
+ $X2=0.27 $Y2=0.495
r77 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.91 $Y=0.81
+ $X2=0.985 $Y2=0.885
r78 1 2 243.564 $w=1.5e-07 $l=4.75e-07 $layer=POLY_cond $X=0.91 $Y=0.81
+ $X2=0.435 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_LS__NOR4_2%B 1 3 6 8 10 11 14 17 18 19 20 28 29 35 47
c74 6 0 7.78362e-20 $X=2.5 $Y=0.74
c75 1 0 3.55766e-19 $X=2.375 $Y=1.765
r76 35 47 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=4.05 $Y=1.71
+ $X2=4.05 $Y2=1.665
r77 33 34 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.05
+ $Y=1.465 $X2=4.05 $Y2=1.465
r78 28 29 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.05
+ $Y=0.445 $X2=4.05 $Y2=0.445
r79 26 33 10.4688 $w=4.9e-07 $l=8e-08 $layer=POLY_cond $X=3.97 $Y=1.385 $X2=3.97
+ $Y2=1.465
r80 26 28 102.638 $w=4.9e-07 $l=9.4e-07 $layer=POLY_cond $X=3.97 $Y=1.385
+ $X2=3.97 $Y2=0.445
r81 20 35 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.05 $Y=1.795 $X2=4.05
+ $Y2=1.71
r82 20 47 0.69845 $w=3.28e-07 $l=2e-08 $layer=LI1_cond $X=4.05 $Y=1.645 $X2=4.05
+ $Y2=1.665
r83 20 34 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=4.05 $Y=1.645
+ $X2=4.05 $Y2=1.465
r84 19 34 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=4.05 $Y=1.295
+ $X2=4.05 $Y2=1.465
r85 18 19 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=4.05 $Y=0.925
+ $X2=4.05 $Y2=1.295
r86 17 18 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=4.05 $Y=0.555
+ $X2=4.05 $Y2=0.925
r87 17 29 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=4.05 $Y=0.555
+ $X2=4.05 $Y2=0.445
r88 14 16 14.0074 $w=2.7e-07 $l=3.1e-07 $layer=LI1_cond $X=2.455 $Y=1.485
+ $X2=2.455 $Y2=1.795
r89 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.45
+ $Y=1.485 $X2=2.45 $Y2=1.485
r90 12 16 3.44395 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=2.625 $Y=1.795
+ $X2=2.455 $Y2=1.795
r91 11 20 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.885 $Y=1.795
+ $X2=4.05 $Y2=1.795
r92 11 12 82.2032 $w=1.68e-07 $l=1.26e-06 $layer=LI1_cond $X=3.885 $Y=1.795
+ $X2=2.625 $Y2=1.795
r93 8 33 56.3701 $w=3.79e-07 $l=3.69459e-07 $layer=POLY_cond $X=3.815 $Y=1.765
+ $X2=3.97 $Y2=1.465
r94 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.815 $Y=1.765
+ $X2=3.815 $Y2=2.4
r95 4 15 38.6072 $w=2.91e-07 $l=1.88348e-07 $layer=POLY_cond $X=2.5 $Y=1.32
+ $X2=2.45 $Y2=1.485
r96 4 6 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.5 $Y=1.32 $X2=2.5
+ $Y2=0.74
r97 1 15 57.6553 $w=2.91e-07 $l=3.15278e-07 $layer=POLY_cond $X=2.375 $Y=1.765
+ $X2=2.45 $Y2=1.485
r98 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.375 $Y=1.765
+ $X2=2.375 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__NOR4_2%A 1 3 4 6 7 9 10 15
c43 10 0 1.87727e-19 $X=3.6 $Y=1.295
r44 15 17 11.1969 $w=4.52e-07 $l=1.05e-07 $layer=POLY_cond $X=3.26 $Y=1.492
+ $X2=3.365 $Y2=1.492
r45 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.26
+ $Y=1.385 $X2=3.26 $Y2=1.385
r46 13 15 35.1903 $w=4.52e-07 $l=3.3e-07 $layer=POLY_cond $X=2.93 $Y=1.492
+ $X2=3.26 $Y2=1.492
r47 12 13 1.59956 $w=4.52e-07 $l=1.5e-08 $layer=POLY_cond $X=2.915 $Y=1.492
+ $X2=2.93 $Y2=1.492
r48 10 16 10.8842 $w=3.58e-07 $l=3.4e-07 $layer=LI1_cond $X=3.6 $Y=1.36 $X2=3.26
+ $Y2=1.36
r49 7 17 28.877 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=3.365 $Y=1.765
+ $X2=3.365 $Y2=1.492
r50 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.365 $Y=1.765
+ $X2=3.365 $Y2=2.4
r51 4 13 28.877 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=2.93 $Y=1.22 $X2=2.93
+ $Y2=1.492
r52 4 6 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.93 $Y=1.22 $X2=2.93
+ $Y2=0.74
r53 1 12 28.877 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=2.915 $Y=1.765
+ $X2=2.915 $Y2=1.492
r54 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.915 $Y=1.765
+ $X2=2.915 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__NOR4_2%A_27_368# 1 2 3 12 14 18 20 22 24 27 32
c59 32 0 1.68039e-19 $X=2.12 $Y=1.985
r60 34 35 12.4464 $w=2.48e-07 $l=2.7e-07 $layer=LI1_cond $X=2.16 $Y=2.135
+ $X2=2.16 $Y2=2.405
r61 32 34 6.91466 $w=2.48e-07 $l=1.5e-07 $layer=LI1_cond $X=2.16 $Y=1.985
+ $X2=2.16 $Y2=2.135
r62 29 30 3.67308 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=0.28 $Y=2.405
+ $X2=0.28 $Y2=2.49
r63 27 29 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=0.28 $Y=2.155
+ $X2=0.28 $Y2=2.405
r64 22 37 2.8391 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=4.072 $Y=2.22
+ $X2=4.072 $Y2=2.135
r65 22 24 25.8756 $w=2.63e-07 $l=5.95e-07 $layer=LI1_cond $X=4.072 $Y=2.22
+ $X2=4.072 $Y2=2.815
r66 21 34 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.285 $Y=2.135
+ $X2=2.16 $Y2=2.135
r67 20 37 4.40896 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=3.94 $Y=2.135
+ $X2=4.072 $Y2=2.135
r68 20 21 107.973 $w=1.68e-07 $l=1.655e-06 $layer=LI1_cond $X=3.94 $Y=2.135
+ $X2=2.285 $Y2=2.135
r69 16 35 3.91831 $w=2.48e-07 $l=8.5e-08 $layer=LI1_cond $X=2.16 $Y=2.49
+ $X2=2.16 $Y2=2.405
r70 16 18 14.9818 $w=2.48e-07 $l=3.25e-07 $layer=LI1_cond $X=2.16 $Y=2.49
+ $X2=2.16 $Y2=2.815
r71 15 29 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.445 $Y=2.405
+ $X2=0.28 $Y2=2.405
r72 14 35 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.035 $Y=2.405
+ $X2=2.16 $Y2=2.405
r73 14 15 103.733 $w=1.68e-07 $l=1.59e-06 $layer=LI1_cond $X=2.035 $Y=2.405
+ $X2=0.445 $Y2=2.405
r74 12 30 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=0.24 $Y=2.495
+ $X2=0.24 $Y2=2.49
r75 3 37 600 $w=1.7e-07 $l=3.62319e-07 $layer=licon1_PDIFF $count=1 $X=3.89
+ $Y=1.84 $X2=4.04 $Y2=2.135
r76 3 24 600 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=3.89
+ $Y=1.84 $X2=4.04 $Y2=2.815
r77 2 32 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=1.97
+ $Y=1.84 $X2=2.12 $Y2=1.985
r78 2 18 600 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.97
+ $Y=1.84 $X2=2.12 $Y2=2.815
r79 1 27 600 $w=1.7e-07 $l=3.80657e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.155
r80 1 12 300 $w=1.7e-07 $l=7.23878e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.495
.ends

.subckt PM_SKY130_FD_SC_LS__NOR4_2%A_116_368# 1 2 11
r15 8 11 33.6729 $w=3.18e-07 $l=9.35e-07 $layer=LI1_cond $X=0.735 $Y=2.82
+ $X2=1.67 $Y2=2.82
r16 2 11 600 $w=1.7e-07 $l=1.01223e-06 $layer=licon1_PDIFF $count=1 $X=1.52
+ $Y=1.84 $X2=1.67 $Y2=2.78
r17 1 8 600 $w=1.7e-07 $l=9.79439e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.84 $X2=0.735 $Y2=2.745
.ends

.subckt PM_SKY130_FD_SC_LS__NOR4_2%Y 1 2 3 11 12 13 15 18 20 24 26 31 32 36
c78 26 0 7.78362e-20 $X=1.715 $Y=0.915
r79 31 32 11.9608 $w=4.78e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.91 $X2=1.2
+ $Y2=1.91
r80 31 36 7.90124 $w=4.78e-07 $l=1.05e-07 $layer=LI1_cond $X=0.72 $Y=1.91
+ $X2=0.615 $Y2=1.91
r81 28 29 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=1.715 $Y=0.965
+ $X2=1.715 $Y2=1.065
r82 26 28 1.74613 $w=3.28e-07 $l=5e-08 $layer=LI1_cond $X=1.715 $Y=0.915
+ $X2=1.715 $Y2=0.965
r83 22 24 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=2.715 $Y=0.98
+ $X2=2.715 $Y2=0.515
r84 21 29 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.88 $Y=1.065
+ $X2=1.715 $Y2=1.065
r85 20 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.55 $Y=1.065
+ $X2=2.715 $Y2=0.98
r86 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.55 $Y=1.065
+ $X2=1.88 $Y2=1.065
r87 16 26 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=1.715 $Y=0.83
+ $X2=1.715 $Y2=0.915
r88 16 18 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=1.715 $Y=0.83
+ $X2=1.715 $Y2=0.515
r89 15 36 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=0.255 $Y=1.755
+ $X2=0.615 $Y2=1.755
r90 12 26 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.55 $Y=0.915
+ $X2=1.715 $Y2=0.915
r91 12 13 84.4866 $w=1.68e-07 $l=1.295e-06 $layer=LI1_cond $X=1.55 $Y=0.915
+ $X2=0.255 $Y2=0.915
r92 11 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.17 $Y=1.67
+ $X2=0.255 $Y2=1.755
r93 10 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.17 $Y=1
+ $X2=0.255 $Y2=0.915
r94 10 11 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.17 $Y=1 $X2=0.17
+ $Y2=1.67
r95 3 32 600 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_PDIFF $count=1 $X=1.045
+ $Y=1.84 $X2=1.205 $Y2=1.985
r96 2 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.575
+ $Y=0.37 $X2=2.715 $Y2=0.515
r97 1 28 182 $w=1.7e-07 $l=6.79062e-07 $layer=licon1_NDIFF $count=1 $X=1.535
+ $Y=0.37 $X2=1.715 $Y2=0.965
r98 1 18 182 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_NDIFF $count=1 $X=1.535
+ $Y=0.37 $X2=1.715 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__NOR4_2%A_490_368# 1 2 9 11 13 16
r28 11 18 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.63 $Y=2.56 $X2=3.63
+ $Y2=2.475
r29 11 13 12.6769 $w=2.48e-07 $l=2.75e-07 $layer=LI1_cond $X=3.63 $Y=2.56
+ $X2=3.63 $Y2=2.835
r30 10 16 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.805 $Y=2.475
+ $X2=2.64 $Y2=2.475
r31 9 18 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.505 $Y=2.475
+ $X2=3.63 $Y2=2.475
r32 9 10 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=3.505 $Y=2.475
+ $X2=2.805 $Y2=2.475
r33 2 18 600 $w=1.7e-07 $l=7.06028e-07 $layer=licon1_PDIFF $count=1 $X=3.44
+ $Y=1.84 $X2=3.59 $Y2=2.475
r34 2 13 600 $w=1.7e-07 $l=1.06737e-06 $layer=licon1_PDIFF $count=1 $X=3.44
+ $Y=1.84 $X2=3.59 $Y2=2.835
r35 1 16 300 $w=1.7e-07 $l=7.43959e-07 $layer=licon1_PDIFF $count=2 $X=2.45
+ $Y=1.84 $X2=2.64 $Y2=2.495
.ends

.subckt PM_SKY130_FD_SC_LS__NOR4_2%VPWR 1 6 8 10 20 21 24
r47 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r48 21 25 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.12 $Y2=3.33
r49 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r50 18 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.305 $Y=3.33
+ $X2=3.14 $Y2=3.33
r51 18 20 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=3.305 $Y=3.33
+ $X2=4.08 $Y2=3.33
r52 17 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r53 16 17 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r54 12 16 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=2.64 $Y2=3.33
r55 12 13 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r56 10 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.975 $Y=3.33
+ $X2=3.14 $Y2=3.33
r57 10 16 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.975 $Y=3.33
+ $X2=2.64 $Y2=3.33
r58 8 17 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r59 8 13 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=0.24 $Y2=3.33
r60 4 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.14 $Y=3.245 $X2=3.14
+ $Y2=3.33
r61 4 6 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.14 $Y=3.245 $X2=3.14
+ $Y2=2.815
r62 1 6 600 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.99
+ $Y=1.84 $X2=3.14 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_LS__NOR4_2%VGND 1 2 3 12 14 18 20 27 34 35 40 46 48 51
c52 35 0 6.36756e-20 $X=4.08 $Y=0
r53 51 52 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r54 45 46 10.7086 $w=6.83e-07 $l=1.65e-07 $layer=LI1_cond $X=1.215 $Y=0.257
+ $X2=1.38 $Y2=0.257
r55 42 45 0.261915 $w=6.83e-07 $l=1.5e-08 $layer=LI1_cond $X=1.2 $Y=0.257
+ $X2=1.215 $Y2=0.257
r56 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r57 39 43 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r58 38 42 8.38128 $w=6.83e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=0.257
+ $X2=1.2 $Y2=0.257
r59 38 40 9.83558 $w=6.83e-07 $l=1.15e-07 $layer=LI1_cond $X=0.72 $Y=0.257
+ $X2=0.605 $Y2=0.257
r60 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r61 35 52 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.12
+ $Y2=0
r62 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r63 32 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.38 $Y=0 $X2=3.215
+ $Y2=0
r64 32 34 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=3.38 $Y=0 $X2=4.08
+ $Y2=0
r65 31 43 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r66 30 46 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.68 $Y=0 $X2=1.38
+ $Y2=0
r67 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r68 27 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.05 $Y=0 $X2=2.215
+ $Y2=0
r69 27 30 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.05 $Y=0 $X2=1.68
+ $Y2=0
r70 25 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r71 24 40 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.24 $Y=0 $X2=0.605
+ $Y2=0
r72 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r73 20 52 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r74 20 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r75 20 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r76 16 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.215 $Y=0.085
+ $X2=3.215 $Y2=0
r77 16 18 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=3.215 $Y=0.085
+ $X2=3.215 $Y2=0.505
r78 15 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.38 $Y=0 $X2=2.215
+ $Y2=0
r79 14 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.05 $Y=0 $X2=3.215
+ $Y2=0
r80 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.05 $Y=0 $X2=2.38
+ $Y2=0
r81 10 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.215 $Y=0.085
+ $X2=2.215 $Y2=0
r82 10 12 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=2.215 $Y=0.085
+ $X2=2.215 $Y2=0.645
r83 3 18 91 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=2 $X=3.005
+ $Y=0.37 $X2=3.145 $Y2=0.505
r84 2 12 182 $w=1.7e-07 $l=3.65205e-07 $layer=licon1_NDIFF $count=1 $X=2.005
+ $Y=0.37 $X2=2.215 $Y2=0.645
r85 1 45 91 $w=1.7e-07 $l=6.58521e-07 $layer=licon1_NDIFF $count=2 $X=0.625
+ $Y=0.37 $X2=1.215 $Y2=0.515
.ends

