* File: sky130_fd_sc_ls__einvp_2.pex.spice
* Created: Wed Sep  2 11:07:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__EINVP_2%A 1 3 4 6 7 9 10 12 13 20
c44 10 0 1.9142e-19 $X=0.97 $Y=1.22
c45 7 0 1.88367e-19 $X=0.955 $Y=1.765
r46 20 21 1.75485 $w=4.12e-07 $l=1.5e-08 $layer=POLY_cond $X=0.955 $Y=1.492
+ $X2=0.97 $Y2=1.492
r47 19 20 48.551 $w=4.12e-07 $l=4.15e-07 $layer=POLY_cond $X=0.54 $Y=1.492
+ $X2=0.955 $Y2=1.492
r48 18 19 4.09466 $w=4.12e-07 $l=3.5e-08 $layer=POLY_cond $X=0.505 $Y=1.492
+ $X2=0.54 $Y2=1.492
r49 16 18 27.4927 $w=4.12e-07 $l=2.35e-07 $layer=POLY_cond $X=0.27 $Y=1.492
+ $X2=0.505 $Y2=1.492
r50 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.385 $X2=0.27 $Y2=1.385
r51 13 17 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.27 $Y=1.295 $X2=0.27
+ $Y2=1.385
r52 10 21 26.5862 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=0.97 $Y=1.22
+ $X2=0.97 $Y2=1.492
r53 10 12 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.97 $Y=1.22 $X2=0.97
+ $Y2=0.74
r54 7 20 26.5862 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=0.955 $Y=1.765
+ $X2=0.955 $Y2=1.492
r55 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.955 $Y=1.765
+ $X2=0.955 $Y2=2.4
r56 4 19 26.5862 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=0.54 $Y=1.22
+ $X2=0.54 $Y2=1.492
r57 4 6 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.54 $Y=1.22 $X2=0.54
+ $Y2=0.74
r58 1 18 26.5862 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=1.492
r59 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__EINVP_2%A_263_323# 1 2 7 9 10 11 12 14 17 20 21 26
+ 30
c61 11 0 6.25938e-20 $X=1.48 $Y=1.69
r62 26 28 5.95495 $w=3.83e-07 $l=1.9e-07 $layer=LI1_cond $X=2.607 $Y=0.95
+ $X2=2.607 $Y2=1.14
r63 21 30 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.58 $Y=1.72
+ $X2=2.415 $Y2=1.72
r64 20 23 26.0173 $w=3.28e-07 $l=7.45e-07 $layer=LI1_cond $X=2.58 $Y=1.72
+ $X2=2.58 $Y2=2.465
r65 20 28 20.2551 $w=3.28e-07 $l=5.8e-07 $layer=LI1_cond $X=2.58 $Y=1.72
+ $X2=2.58 $Y2=1.14
r66 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.58
+ $Y=1.72 $X2=2.58 $Y2=1.72
r67 16 17 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.93 $Y=1.69
+ $X2=1.855 $Y2=1.69
r68 16 30 248.691 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=1.93 $Y=1.69
+ $X2=2.415 $Y2=1.69
r69 12 17 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.855 $Y=1.765
+ $X2=1.855 $Y2=1.69
r70 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.855 $Y=1.765
+ $X2=1.855 $Y2=2.4
r71 10 17 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.78 $Y=1.69
+ $X2=1.855 $Y2=1.69
r72 10 11 153.83 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=1.78 $Y=1.69 $X2=1.48
+ $Y2=1.69
r73 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.405 $Y=1.765
+ $X2=1.48 $Y2=1.69
r74 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.405 $Y=1.765
+ $X2=1.405 $Y2=2.4
r75 2 23 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.49
+ $Y=2.32 $X2=2.63 $Y2=2.465
r76 1 26 182 $w=1.7e-07 $l=3.14245e-07 $layer=licon1_NDIFF $count=1 $X=2.49
+ $Y=0.7 $X2=2.635 $Y2=0.95
.ends

.subckt PM_SKY130_FD_SC_LS__EINVP_2%TE 1 3 4 5 6 8 9 12 16 17 19 21 22 25 29 31
+ 35 36
r65 35 37 36.4613 $w=2.71e-07 $l=2.05e-07 $layer=POLY_cond $X=2.645 $Y=0.425
+ $X2=2.85 $Y2=0.425
r66 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.645
+ $Y=0.425 $X2=2.645 $Y2=0.425
r67 31 36 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=2.645 $Y=0.555
+ $X2=2.645 $Y2=0.425
r68 27 29 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=2.85 $Y=1.27
+ $X2=3.06 $Y2=1.27
r69 23 25 105.117 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=2.855 $Y=2.17
+ $X2=3.06 $Y2=2.17
r70 21 25 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.06 $Y=2.095
+ $X2=3.06 $Y2=2.17
r71 20 29 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.06 $Y=1.345
+ $X2=3.06 $Y2=1.27
r72 20 21 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=3.06 $Y=1.345
+ $X2=3.06 $Y2=2.095
r73 17 23 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.855 $Y=2.245
+ $X2=2.855 $Y2=2.17
r74 17 19 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.855 $Y=2.245
+ $X2=2.855 $Y2=2.64
r75 14 27 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.85 $Y=1.195
+ $X2=2.85 $Y2=1.27
r76 14 16 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.85 $Y=1.195
+ $X2=2.85 $Y2=0.91
r77 13 37 16.5906 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.85 $Y=0.59
+ $X2=2.85 $Y2=0.425
r78 13 16 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.85 $Y=0.59
+ $X2=2.85 $Y2=0.91
r79 11 35 54.2472 $w=2.71e-07 $l=3.78616e-07 $layer=POLY_cond $X=2.34 $Y=0.59
+ $X2=2.645 $Y2=0.425
r80 11 12 305.096 $w=1.5e-07 $l=5.95e-07 $layer=POLY_cond $X=2.34 $Y=0.59
+ $X2=2.34 $Y2=1.185
r81 10 22 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.905 $Y=1.26
+ $X2=1.83 $Y2=1.26
r82 9 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.265 $Y=1.26
+ $X2=2.34 $Y2=1.185
r83 9 10 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=2.265 $Y=1.26
+ $X2=1.905 $Y2=1.26
r84 6 22 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.83 $Y=1.185
+ $X2=1.83 $Y2=1.26
r85 6 8 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.83 $Y=1.185
+ $X2=1.83 $Y2=0.74
r86 4 22 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.755 $Y=1.26
+ $X2=1.83 $Y2=1.26
r87 4 5 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.755 $Y=1.26
+ $X2=1.475 $Y2=1.26
r88 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.4 $Y=1.185
+ $X2=1.475 $Y2=1.26
r89 1 3 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.4 $Y=1.185 $X2=1.4
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__EINVP_2%A_27_368# 1 2 3 12 16 17 21 24 25 28
c50 21 0 1.40666e-19 $X=1.18 $Y=1.985
r51 28 30 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=2.04 $Y=1.985
+ $X2=2.04 $Y2=2.815
r52 26 28 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=2.04 $Y=1.65
+ $X2=2.04 $Y2=1.985
r53 24 26 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.915 $Y=1.565
+ $X2=2.04 $Y2=1.65
r54 24 25 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.915 $Y=1.565
+ $X2=1.265 $Y2=1.565
r55 21 23 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=1.18 $Y=1.985
+ $X2=1.18 $Y2=2.815
r56 19 23 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=1.18 $Y=2.905 $X2=1.18
+ $Y2=2.815
r57 18 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.18 $Y=1.65
+ $X2=1.265 $Y2=1.565
r58 18 21 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.18 $Y=1.65
+ $X2=1.18 $Y2=1.985
r59 16 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.095 $Y=2.99
+ $X2=1.18 $Y2=2.905
r60 16 17 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.095 $Y=2.99
+ $X2=0.365 $Y2=2.99
r61 12 15 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=0.24 $Y=1.985
+ $X2=0.24 $Y2=2.815
r62 10 17 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.24 $Y=2.905
+ $X2=0.365 $Y2=2.99
r63 10 15 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=0.24 $Y=2.905 $X2=0.24
+ $Y2=2.815
r64 3 30 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.93
+ $Y=1.84 $X2=2.08 $Y2=2.815
r65 3 28 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.93
+ $Y=1.84 $X2=2.08 $Y2=1.985
r66 2 23 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.03
+ $Y=1.84 $X2=1.18 $Y2=2.815
r67 2 21 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.03
+ $Y=1.84 $X2=1.18 $Y2=1.985
r68 1 15 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r69 1 12 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_LS__EINVP_2%Z 1 2 9 11 12 13 14 33
c22 11 0 6.25938e-20 $X=0.635 $Y=1.21
r23 20 33 1.53659 $w=3.13e-07 $l=4.2e-08 $layer=LI1_cond $X=0.762 $Y=1.337
+ $X2=0.762 $Y2=1.295
r24 13 14 15.3659 $w=3.13e-07 $l=4.2e-07 $layer=LI1_cond $X=0.762 $Y=1.985
+ $X2=0.762 $Y2=2.405
r25 12 13 11.7074 $w=3.13e-07 $l=3.2e-07 $layer=LI1_cond $X=0.762 $Y=1.665
+ $X2=0.762 $Y2=1.985
r26 11 33 0.804881 $w=3.13e-07 $l=2.2e-08 $layer=LI1_cond $X=0.762 $Y=1.273
+ $X2=0.762 $Y2=1.295
r27 11 31 3.92579 $w=3.13e-07 $l=9.3e-08 $layer=LI1_cond $X=0.762 $Y=1.273
+ $X2=0.762 $Y2=1.18
r28 11 12 11.2317 $w=3.13e-07 $l=3.07e-07 $layer=LI1_cond $X=0.762 $Y=1.358
+ $X2=0.762 $Y2=1.665
r29 11 20 0.768295 $w=3.13e-07 $l=2.1e-08 $layer=LI1_cond $X=0.762 $Y=1.358
+ $X2=0.762 $Y2=1.337
r30 9 31 16.5952 $w=2.48e-07 $l=3.6e-07 $layer=LI1_cond $X=0.795 $Y=0.82
+ $X2=0.795 $Y2=1.18
r31 2 13 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=0.58
+ $Y=1.84 $X2=0.73 $Y2=1.985
r32 1 9 182 $w=1.7e-07 $l=5.15267e-07 $layer=licon1_NDIFF $count=1 $X=0.615
+ $Y=0.37 $X2=0.755 $Y2=0.82
.ends

.subckt PM_SKY130_FD_SC_LS__EINVP_2%VPWR 1 2 9 13 15 17 19 27 33 37
c36 9 0 1.88367e-19 $X=1.63 $Y=1.985
r37 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r38 31 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r39 30 31 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r40 28 33 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.715 $Y=3.33
+ $X2=1.59 $Y2=3.33
r41 28 30 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=1.715 $Y=3.33
+ $X2=2.64 $Y2=3.33
r42 27 36 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=2.915 $Y=3.33
+ $X2=3.137 $Y2=3.33
r43 27 30 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.915 $Y=3.33
+ $X2=2.64 $Y2=3.33
r44 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r45 22 26 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r46 21 25 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=3.33 $X2=1.2
+ $Y2=3.33
r47 21 22 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r48 19 33 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.465 $Y=3.33
+ $X2=1.59 $Y2=3.33
r49 19 25 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.465 $Y=3.33
+ $X2=1.2 $Y2=3.33
r50 17 31 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r51 17 26 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r52 17 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r53 13 36 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=3.08 $Y=3.245
+ $X2=3.137 $Y2=3.33
r54 13 15 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=3.08 $Y=3.245
+ $X2=3.08 $Y2=2.465
r55 9 12 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=1.59 $Y=1.985
+ $X2=1.59 $Y2=2.815
r56 7 33 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.59 $Y=3.245
+ $X2=1.59 $Y2=3.33
r57 7 12 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=1.59 $Y=3.245 $X2=1.59
+ $Y2=2.815
r58 2 15 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=2.93
+ $Y=2.32 $X2=3.08 $Y2=2.465
r59 1 12 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.48
+ $Y=1.84 $X2=1.63 $Y2=2.815
r60 1 9 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.48
+ $Y=1.84 $X2=1.63 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_LS__EINVP_2%A_36_74# 1 2 3 12 14 15 19 20 21 24
r48 22 24 27.703 $w=2.58e-07 $l=6.25e-07 $layer=LI1_cond $X=2.08 $Y=1.14
+ $X2=2.08 $Y2=0.515
r49 20 22 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=1.95 $Y=1.225
+ $X2=2.08 $Y2=1.14
r50 20 21 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.95 $Y=1.225
+ $X2=1.27 $Y2=1.225
r51 17 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.185 $Y=1.14
+ $X2=1.27 $Y2=1.225
r52 17 19 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=1.185 $Y=1.14
+ $X2=1.185 $Y2=0.515
r53 16 19 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=1.185 $Y=0.425
+ $X2=1.185 $Y2=0.515
r54 14 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.1 $Y=0.34
+ $X2=1.185 $Y2=0.425
r55 14 15 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=1.1 $Y=0.34 $X2=0.49
+ $Y2=0.34
r56 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.325 $Y=0.425
+ $X2=0.49 $Y2=0.34
r57 10 12 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.325 $Y=0.425
+ $X2=0.325 $Y2=0.515
r58 3 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.905
+ $Y=0.37 $X2=2.045 $Y2=0.515
r59 2 19 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.045
+ $Y=0.37 $X2=1.185 $Y2=0.515
r60 1 12 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.18
+ $Y=0.37 $X2=0.325 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__EINVP_2%VGND 1 2 9 11 13 15 17 25 31 35
c35 9 0 1.9142e-19 $X=1.615 $Y=0.515
r36 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r37 29 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r38 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r39 26 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.78 $Y=0 $X2=1.615
+ $Y2=0
r40 26 28 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=1.78 $Y=0 $X2=2.64
+ $Y2=0
r41 25 34 4.13553 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.98 $Y=0 $X2=3.17
+ $Y2=0
r42 25 28 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.98 $Y=0 $X2=2.64
+ $Y2=0
r43 23 24 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r44 20 24 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r45 19 23 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r46 19 20 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r47 17 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.45 $Y=0 $X2=1.615
+ $Y2=0
r48 17 23 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.45 $Y=0 $X2=1.2
+ $Y2=0
r49 15 29 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r50 15 24 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r51 15 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r52 11 34 3.11253 $w=2.65e-07 $l=1.1025e-07 $layer=LI1_cond $X=3.112 $Y=0.085
+ $X2=3.17 $Y2=0
r53 11 13 33.0512 $w=2.63e-07 $l=7.6e-07 $layer=LI1_cond $X=3.112 $Y=0.085
+ $X2=3.112 $Y2=0.845
r54 7 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.615 $Y=0.085
+ $X2=1.615 $Y2=0
r55 7 9 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=1.615 $Y=0.085
+ $X2=1.615 $Y2=0.515
r56 2 13 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=2.925
+ $Y=0.7 $X2=3.07 $Y2=0.845
r57 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.475
+ $Y=0.37 $X2=1.615 $Y2=0.515
.ends

