* File: sky130_fd_sc_ls__or3_2.spice
* Created: Fri Aug 28 13:58:24 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__or3_2.pex.spice"
.subckt sky130_fd_sc_ls__or3_2  VNB VPB C B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* C	C
* VPB	VPB
* VNB	VNB
MM1008 N_VGND_M1008_d N_C_M1008_g N_A_27_74#_M1008_s VNB NSHORT L=0.15 W=0.64
+ AD=0.1616 AS=0.1824 PD=1.145 PS=1.85 NRD=20.616 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75002.6 A=0.096 P=1.58 MULT=1
MM1006 N_A_27_74#_M1006_d N_B_M1006_g N_VGND_M1008_d VNB NSHORT L=0.15 W=0.64
+ AD=0.112 AS=0.1616 PD=0.99 PS=1.145 NRD=0 NRS=21.552 M=1 R=4.26667 SA=75000.9
+ SB=75001.9 A=0.096 P=1.58 MULT=1
MM1004 N_VGND_M1004_d N_A_M1004_g N_A_27_74#_M1006_d VNB NSHORT L=0.15 W=0.64
+ AD=0.179293 AS=0.112 PD=1.21043 PS=0.99 NRD=19.68 NRS=13.116 M=1 R=4.26667
+ SA=75001.4 SB=75001.4 A=0.096 P=1.58 MULT=1
MM1005 N_X_M1005_d N_A_27_74#_M1005_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.207307 PD=1.02 PS=1.39957 NRD=0 NRS=29.184 M=1 R=4.93333
+ SA=75001.8 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1009 N_X_M1005_d N_A_27_74#_M1009_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.2627 PD=1.02 PS=2.19 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75002.3
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1003 A_150_392# N_C_M1003_g N_A_27_74#_M1003_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.295 PD=1.27 PS=2.59 NRD=15.7403 NRS=1.9503 M=1 R=6.66667 SA=75000.2
+ SB=75002.3 A=0.15 P=2.3 MULT=1
MM1002 A_234_392# N_B_M1002_g A_150_392# VPB PHIGHVT L=0.15 W=1 AD=0.21 AS=0.135
+ PD=1.42 PS=1.27 NRD=30.5153 NRS=15.7403 M=1 R=6.66667 SA=75000.6 SB=75001.9
+ A=0.15 P=2.3 MULT=1
MM1001 N_VPWR_M1001_d N_A_M1001_g A_234_392# VPB PHIGHVT L=0.15 W=1 AD=0.231981
+ AS=0.21 PD=1.49057 PS=1.42 NRD=1.9503 NRS=30.5153 M=1 R=6.66667 SA=75001.2
+ SB=75001.3 A=0.15 P=2.3 MULT=1
MM1000 N_VPWR_M1001_d N_A_27_74#_M1000_g N_X_M1000_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.259819 AS=0.168 PD=1.66943 PS=1.42 NRD=29.8849 NRS=1.7533 M=1 R=7.46667
+ SA=75001.6 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1007 N_VPWR_M1007_d N_A_27_74#_M1007_g N_X_M1000_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3864 AS=0.168 PD=2.93 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75002.1 SB=75000.3 A=0.168 P=2.54 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9564 P=11.2
*
.include "sky130_fd_sc_ls__or3_2.pxi.spice"
*
.ends
*
*
