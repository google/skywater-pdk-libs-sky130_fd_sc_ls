# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ls__fah_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ls__fah_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  13.92000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.820000 1.470000 13.490000 1.800000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.723000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.145000 1.180000 9.475000 1.550000 ;
    END
  END B
  PIN CI
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005000 1.410000 1.335000 1.780000 ;
    END
  END CI
  PIN COUT
    ANTENNADIFFAREA  0.674850 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.665000 0.730000 1.675000 0.900000 ;
        RECT 0.665000 0.900000 0.835000 1.950000 ;
        RECT 0.665000 1.950000 1.155000 2.120000 ;
        RECT 0.985000 2.120000 1.155000 2.905000 ;
        RECT 0.985000 2.905000 2.645000 3.075000 ;
        RECT 1.505000 0.400000 2.075000 0.730000 ;
        RECT 2.315000 2.875000 2.645000 2.905000 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  0.537600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.110000 0.540000 0.445000 2.980000 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 13.920000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 13.920000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 13.920000 0.085000 ;
      RECT  0.000000  3.245000 13.920000 3.415000 ;
      RECT  0.620000  0.085000  0.950000 0.560000 ;
      RECT  0.645000  2.290000  0.815000 3.245000 ;
      RECT  1.130000  1.070000  1.675000 1.240000 ;
      RECT  1.325000  1.950000  1.675000 2.535000 ;
      RECT  1.325000  2.535000  2.985000 2.625000 ;
      RECT  1.325000  2.625000  3.630000 2.705000 ;
      RECT  1.325000  2.705000  1.675000 2.735000 ;
      RECT  1.505000  1.240000  1.675000 1.950000 ;
      RECT  1.845000  0.900000  2.765000 1.070000 ;
      RECT  1.845000  1.070000  2.175000 2.195000 ;
      RECT  1.845000  2.195000  3.325000 2.285000 ;
      RECT  1.845000  2.285000  4.535000 2.365000 ;
      RECT  2.255000  0.085000  2.425000 0.730000 ;
      RECT  2.500000  1.240000  3.105000 1.410000 ;
      RECT  2.500000  1.410000  2.830000 1.635000 ;
      RECT  2.595000  0.255000  4.285000 0.425000 ;
      RECT  2.595000  0.425000  2.765000 0.900000 ;
      RECT  2.815000  2.705000  3.630000 2.795000 ;
      RECT  2.935000  0.595000  3.945000 0.765000 ;
      RECT  2.935000  0.765000  3.105000 1.240000 ;
      RECT  2.935000  2.965000  3.290000 3.245000 ;
      RECT  3.005000  1.580000  3.445000 1.855000 ;
      RECT  3.005000  1.855000  4.000000 2.025000 ;
      RECT  3.155000  2.365000  4.535000 2.455000 ;
      RECT  3.275000  0.935000  3.605000 1.185000 ;
      RECT  3.275000  1.185000  3.445000 1.580000 ;
      RECT  3.460000  2.795000  3.630000 2.905000 ;
      RECT  3.460000  2.905000  7.000000 3.075000 ;
      RECT  3.495000  2.025000  4.000000 2.115000 ;
      RECT  3.670000  1.435000  4.340000 1.595000 ;
      RECT  3.670000  1.595000  4.875000 1.685000 ;
      RECT  3.775000  0.765000  3.945000 1.095000 ;
      RECT  3.775000  1.095000  5.215000 1.265000 ;
      RECT  4.115000  0.425000  4.285000 0.755000 ;
      RECT  4.115000  0.755000  6.215000 0.765000 ;
      RECT  4.115000  0.765000  5.045000 0.925000 ;
      RECT  4.170000  1.685000  4.875000 1.765000 ;
      RECT  4.205000  2.100000  4.535000 2.285000 ;
      RECT  4.205000  2.455000  4.535000 2.735000 ;
      RECT  4.455000  0.255000  7.565000 0.425000 ;
      RECT  4.455000  0.425000  4.705000 0.585000 ;
      RECT  4.705000  1.765000  4.875000 2.730000 ;
      RECT  4.705000  2.730000  6.125000 2.905000 ;
      RECT  4.875000  0.595000  6.215000 0.755000 ;
      RECT  4.880000  1.265000  5.215000 1.425000 ;
      RECT  5.045000  1.425000  5.215000 2.320000 ;
      RECT  5.045000  2.320000  6.660000 2.490000 ;
      RECT  5.385000  0.935000  5.715000 1.035000 ;
      RECT  5.385000  1.035000  6.225000 1.205000 ;
      RECT  5.405000  1.375000  5.885000 1.705000 ;
      RECT  5.405000  1.705000  5.635000 2.150000 ;
      RECT  5.885000  0.765000  6.215000 0.865000 ;
      RECT  6.055000  1.205000  6.225000 1.950000 ;
      RECT  6.055000  1.950000  7.000000 2.120000 ;
      RECT  6.330000  2.290000  6.660000 2.320000 ;
      RECT  6.330000  2.490000  6.660000 2.640000 ;
      RECT  6.395000  0.670000  6.565000 1.550000 ;
      RECT  6.395000  1.550000  6.595000 1.780000 ;
      RECT  6.735000  0.710000  7.065000 1.380000 ;
      RECT  6.830000  2.120000  7.000000 2.905000 ;
      RECT  6.845000  1.380000  7.065000 1.550000 ;
      RECT  6.845000  1.550000  7.075000 1.780000 ;
      RECT  7.170000  1.950000  7.500000 2.925000 ;
      RECT  7.235000  0.425000  7.565000 0.620000 ;
      RECT  7.235000  0.620000 10.315000 0.790000 ;
      RECT  7.235000  0.790000  7.565000 1.130000 ;
      RECT  7.330000  1.130000  7.500000 1.950000 ;
      RECT  7.670000  1.765000  8.000000 3.245000 ;
      RECT  7.745000  0.085000  8.075000 0.450000 ;
      RECT  8.170000  0.960000  8.635000 1.210000 ;
      RECT  8.170000  1.210000  8.340000 1.880000 ;
      RECT  8.170000  1.880000  8.610000 2.905000 ;
      RECT  8.170000  2.905000 11.740000 3.075000 ;
      RECT  8.510000  1.380000  8.975000 1.710000 ;
      RECT  8.780000  1.880000  9.110000 2.565000 ;
      RECT  8.780000  2.565000 10.815000 2.735000 ;
      RECT  8.805000  0.790000  8.975000 1.380000 ;
      RECT  8.895000  0.255000 11.155000 0.425000 ;
      RECT  8.895000  0.425000  9.385000 0.450000 ;
      RECT  9.280000  1.805000 10.475000 2.395000 ;
      RECT  9.645000  0.960000  9.975000 1.805000 ;
      RECT 10.145000  0.790000 10.315000 1.220000 ;
      RECT 10.145000  1.220000 10.475000 1.550000 ;
      RECT 10.485000  0.595000 10.815000 1.050000 ;
      RECT 10.645000  1.050000 10.815000 2.565000 ;
      RECT 10.985000  0.425000 11.155000 1.550000 ;
      RECT 10.985000  1.550000 11.215000 1.780000 ;
      RECT 10.985000  1.780000 11.155000 2.735000 ;
      RECT 11.385000  1.130000 11.740000 2.905000 ;
      RECT 11.405000  0.350000 11.740000 1.130000 ;
      RECT 11.910000  0.790000 12.805000 0.960000 ;
      RECT 11.910000  0.960000 12.080000 1.720000 ;
      RECT 11.910000  1.720000 12.650000 1.940000 ;
      RECT 11.915000  0.085000 12.245000 0.620000 ;
      RECT 11.950000  2.110000 12.220000 2.330000 ;
      RECT 11.950000  2.330000 12.290000 3.245000 ;
      RECT 12.250000  1.130000 13.830000 1.300000 ;
      RECT 12.250000  1.300000 12.580000 1.550000 ;
      RECT 12.390000  1.940000 12.650000 1.970000 ;
      RECT 12.390000  1.970000 12.850000 2.160000 ;
      RECT 12.475000  0.350000 12.805000 0.790000 ;
      RECT 12.520000  2.160000 12.850000 2.980000 ;
      RECT 12.975000  0.085000 13.305000 0.960000 ;
      RECT 13.050000  1.970000 13.300000 3.245000 ;
      RECT 13.470000  1.970000 13.830000 2.980000 ;
      RECT 13.475000  0.350000 13.830000 1.130000 ;
      RECT 13.660000  1.300000 13.830000 1.970000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  1.580000  3.205000 1.750000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  1.950000  5.605000 2.120000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  1.580000  6.565000 1.750000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  1.580000  7.045000 1.750000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  8.840000  1.950000  9.010000 2.120000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT  9.885000  1.950000 10.055000 2.120000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.245000  1.950000 10.415000 2.120000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.015000  1.580000 11.185000 1.750000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.435000  1.950000 12.605000 2.120000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.245000 13.285000 3.415000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.245000 13.765000 3.415000 ;
    LAYER met1 ;
      RECT  2.975000 1.550000  3.265000 1.595000 ;
      RECT  2.975000 1.595000  6.625000 1.735000 ;
      RECT  2.975000 1.735000  3.265000 1.780000 ;
      RECT  5.375000 1.920000  5.665000 1.965000 ;
      RECT  5.375000 1.965000  9.070000 2.105000 ;
      RECT  5.375000 2.105000  5.665000 2.150000 ;
      RECT  6.335000 1.550000  6.625000 1.595000 ;
      RECT  6.335000 1.735000  6.625000 1.780000 ;
      RECT  6.815000 1.550000  7.105000 1.595000 ;
      RECT  6.815000 1.595000 11.245000 1.735000 ;
      RECT  6.815000 1.735000  7.105000 1.780000 ;
      RECT  8.780000 1.920000  9.070000 1.965000 ;
      RECT  8.780000 2.105000  9.070000 2.150000 ;
      RECT  9.825000 1.920000 10.475000 1.965000 ;
      RECT  9.825000 1.965000 12.665000 2.105000 ;
      RECT  9.825000 2.105000 10.475000 2.150000 ;
      RECT 10.955000 1.550000 11.245000 1.595000 ;
      RECT 10.955000 1.735000 11.245000 1.780000 ;
      RECT 12.375000 1.920000 12.665000 1.965000 ;
      RECT 12.375000 2.105000 12.665000 2.150000 ;
  END
END sky130_fd_sc_ls__fah_1
END LIBRARY
