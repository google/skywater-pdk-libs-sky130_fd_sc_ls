* NGSPICE file created from sky130_fd_sc_ls__and2b_4.ext - technology: sky130A

.subckt sky130_fd_sc_ls__and2b_4 A_N B VGND VNB VPB VPWR X
M1000 VGND a_218_424# X VNB nshort w=740000u l=150000u
+  ad=9.074e+11p pd=8.29e+06u as=4.218e+11p ps=4.1e+06u
M1001 VPWR a_218_424# X VPB phighvt w=1.12e+06u l=150000u
+  ad=1.7066e+12p pd=1.379e+07u as=6.72e+11p ps=5.68e+06u
M1002 a_218_424# B VPWR VPB phighvt w=840000u l=150000u
+  ad=5.04e+11p pd=4.56e+06u as=0p ps=0u
M1003 a_218_424# a_27_392# VPWR VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 X a_218_424# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_218_424# a_27_392# a_233_74# VNB nshort w=640000u l=150000u
+  ad=1.792e+11p pd=1.84e+06u as=4.16e+11p ps=3.86e+06u
M1006 VGND a_218_424# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_233_74# B VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR B a_218_424# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND A_N a_27_392# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1010 VPWR a_27_392# a_218_424# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR a_218_424# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 X a_218_424# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 X a_218_424# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_233_74# a_27_392# a_218_424# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND B a_233_74# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 X a_218_424# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR A_N a_27_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.85e+11p ps=2.57e+06u
.ends

