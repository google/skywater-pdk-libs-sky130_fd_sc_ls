* File: sky130_fd_sc_ls__sdlclkp_4.pxi.spice
* Created: Wed Sep  2 11:29:03 2020
* 
x_PM_SKY130_FD_SC_LS__SDLCLKP_4%SCE N_SCE_c_177_n N_SCE_M1009_g N_SCE_M1019_g
+ SCE N_SCE_c_179_n PM_SKY130_FD_SC_LS__SDLCLKP_4%SCE
x_PM_SKY130_FD_SC_LS__SDLCLKP_4%GATE N_GATE_c_200_n N_GATE_M1020_g
+ N_GATE_M1025_g GATE PM_SKY130_FD_SC_LS__SDLCLKP_4%GATE
x_PM_SKY130_FD_SC_LS__SDLCLKP_4%A_354_105# N_A_354_105#_M1017_d
+ N_A_354_105#_M1002_d N_A_354_105#_c_231_n N_A_354_105#_M1014_g
+ N_A_354_105#_c_232_n N_A_354_105#_M1016_g N_A_354_105#_c_234_n
+ N_A_354_105#_c_235_n N_A_354_105#_c_236_n N_A_354_105#_c_243_n
+ N_A_354_105#_c_237_n N_A_354_105#_c_238_n N_A_354_105#_c_239_n
+ PM_SKY130_FD_SC_LS__SDLCLKP_4%A_354_105#
x_PM_SKY130_FD_SC_LS__SDLCLKP_4%A_324_79# N_A_324_79#_M1011_s
+ N_A_324_79#_M1023_s N_A_324_79#_c_310_n N_A_324_79#_M1017_g
+ N_A_324_79#_c_311_n N_A_324_79#_c_312_n N_A_324_79#_c_313_n
+ N_A_324_79#_c_330_n N_A_324_79#_M1002_g N_A_324_79#_c_332_n
+ N_A_324_79#_c_333_n N_A_324_79#_c_314_n N_A_324_79#_c_315_n
+ N_A_324_79#_M1022_g N_A_324_79#_c_334_n N_A_324_79#_c_335_n
+ N_A_324_79#_c_336_n N_A_324_79#_M1012_g N_A_324_79#_c_316_n
+ N_A_324_79#_c_317_n N_A_324_79#_c_318_n N_A_324_79#_c_319_n
+ N_A_324_79#_c_320_n N_A_324_79#_c_321_n N_A_324_79#_c_322_n
+ N_A_324_79#_c_377_p N_A_324_79#_c_323_n N_A_324_79#_c_324_n
+ N_A_324_79#_c_325_n N_A_324_79#_c_365_n N_A_324_79#_c_337_n
+ N_A_324_79#_c_326_n N_A_324_79#_c_327_n N_A_324_79#_c_328_n
+ PM_SKY130_FD_SC_LS__SDLCLKP_4%A_324_79#
x_PM_SKY130_FD_SC_LS__SDLCLKP_4%A_792_48# N_A_792_48#_M1004_d
+ N_A_792_48#_M1000_d N_A_792_48#_M1005_g N_A_792_48#_c_482_n
+ N_A_792_48#_c_483_n N_A_792_48#_M1006_g N_A_792_48#_M1008_g
+ N_A_792_48#_c_476_n N_A_792_48#_M1018_g N_A_792_48#_c_485_n
+ N_A_792_48#_c_486_n N_A_792_48#_c_487_n N_A_792_48#_c_477_n
+ N_A_792_48#_c_489_n N_A_792_48#_c_490_n N_A_792_48#_c_512_n
+ N_A_792_48#_c_478_n N_A_792_48#_c_479_n N_A_792_48#_c_492_n
+ N_A_792_48#_c_493_n N_A_792_48#_c_480_n N_A_792_48#_c_481_n
+ PM_SKY130_FD_SC_LS__SDLCLKP_4%A_792_48#
x_PM_SKY130_FD_SC_LS__SDLCLKP_4%A_634_74# N_A_634_74#_M1022_d
+ N_A_634_74#_M1014_d N_A_634_74#_c_601_n N_A_634_74#_M1000_g
+ N_A_634_74#_c_602_n N_A_634_74#_M1004_g N_A_634_74#_c_603_n
+ N_A_634_74#_c_604_n N_A_634_74#_c_605_n N_A_634_74#_c_606_n
+ N_A_634_74#_c_607_n N_A_634_74#_c_608_n
+ PM_SKY130_FD_SC_LS__SDLCLKP_4%A_634_74#
x_PM_SKY130_FD_SC_LS__SDLCLKP_4%CLK N_CLK_c_680_n N_CLK_M1023_g N_CLK_c_676_n
+ N_CLK_M1011_g N_CLK_c_681_n N_CLK_M1015_g N_CLK_c_677_n N_CLK_M1007_g CLK
+ N_CLK_c_679_n PM_SKY130_FD_SC_LS__SDLCLKP_4%CLK
x_PM_SKY130_FD_SC_LS__SDLCLKP_4%A_1289_368# N_A_1289_368#_M1008_d
+ N_A_1289_368#_M1015_d N_A_1289_368#_c_740_n N_A_1289_368#_M1003_g
+ N_A_1289_368#_M1001_g N_A_1289_368#_c_741_n N_A_1289_368#_M1010_g
+ N_A_1289_368#_M1013_g N_A_1289_368#_c_742_n N_A_1289_368#_M1021_g
+ N_A_1289_368#_M1026_g N_A_1289_368#_c_743_n N_A_1289_368#_M1024_g
+ N_A_1289_368#_M1027_g N_A_1289_368#_c_744_n N_A_1289_368#_c_733_n
+ N_A_1289_368#_c_745_n N_A_1289_368#_c_746_n N_A_1289_368#_c_734_n
+ N_A_1289_368#_c_735_n N_A_1289_368#_c_736_n N_A_1289_368#_c_737_n
+ N_A_1289_368#_c_798_p N_A_1289_368#_c_738_n N_A_1289_368#_c_739_n
+ PM_SKY130_FD_SC_LS__SDLCLKP_4%A_1289_368#
x_PM_SKY130_FD_SC_LS__SDLCLKP_4%VPWR N_VPWR_M1009_s N_VPWR_M1002_s
+ N_VPWR_M1006_d N_VPWR_M1023_d N_VPWR_M1018_d N_VPWR_M1010_s N_VPWR_M1024_s
+ N_VPWR_c_853_n N_VPWR_c_854_n N_VPWR_c_855_n N_VPWR_c_856_n N_VPWR_c_857_n
+ N_VPWR_c_858_n N_VPWR_c_859_n N_VPWR_c_860_n N_VPWR_c_861_n N_VPWR_c_862_n
+ VPWR N_VPWR_c_863_n N_VPWR_c_864_n N_VPWR_c_865_n N_VPWR_c_866_n
+ N_VPWR_c_867_n N_VPWR_c_868_n N_VPWR_c_869_n N_VPWR_c_870_n N_VPWR_c_871_n
+ N_VPWR_c_852_n PM_SKY130_FD_SC_LS__SDLCLKP_4%VPWR
x_PM_SKY130_FD_SC_LS__SDLCLKP_4%A_119_143# N_A_119_143#_M1019_d
+ N_A_119_143#_M1022_s N_A_119_143#_M1020_d N_A_119_143#_M1014_s
+ N_A_119_143#_c_960_n N_A_119_143#_c_961_n N_A_119_143#_c_962_n
+ N_A_119_143#_c_963_n N_A_119_143#_c_967_n N_A_119_143#_c_968_n
+ N_A_119_143#_c_969_n N_A_119_143#_c_970_n N_A_119_143#_c_1012_n
+ N_A_119_143#_c_964_n N_A_119_143#_c_965_n
+ PM_SKY130_FD_SC_LS__SDLCLKP_4%A_119_143#
x_PM_SKY130_FD_SC_LS__SDLCLKP_4%GCLK N_GCLK_M1001_s N_GCLK_M1026_s
+ N_GCLK_M1003_d N_GCLK_M1021_d N_GCLK_c_1058_n N_GCLK_c_1053_n N_GCLK_c_1059_n
+ N_GCLK_c_1060_n N_GCLK_c_1054_n N_GCLK_c_1055_n N_GCLK_c_1061_n
+ N_GCLK_c_1056_n N_GCLK_c_1057_n N_GCLK_c_1063_n GCLK N_GCLK_c_1098_n
+ PM_SKY130_FD_SC_LS__SDLCLKP_4%GCLK
x_PM_SKY130_FD_SC_LS__SDLCLKP_4%VGND N_VGND_M1019_s N_VGND_M1025_d
+ N_VGND_M1005_d N_VGND_M1011_d N_VGND_M1001_d N_VGND_M1013_d N_VGND_M1027_d
+ N_VGND_c_1124_n N_VGND_c_1125_n N_VGND_c_1126_n N_VGND_c_1127_n
+ N_VGND_c_1128_n N_VGND_c_1129_n N_VGND_c_1130_n N_VGND_c_1131_n
+ N_VGND_c_1132_n N_VGND_c_1133_n N_VGND_c_1134_n N_VGND_c_1135_n
+ N_VGND_c_1136_n VGND N_VGND_c_1137_n N_VGND_c_1138_n N_VGND_c_1139_n
+ N_VGND_c_1140_n N_VGND_c_1141_n N_VGND_c_1142_n N_VGND_c_1143_n
+ PM_SKY130_FD_SC_LS__SDLCLKP_4%VGND
cc_1 VNB N_SCE_c_177_n 0.0230926f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.9
cc_2 VNB N_SCE_M1019_g 0.0277275f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.99
cc_3 VNB N_SCE_c_179_n 0.00872743f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.62
cc_4 VNB N_GATE_c_200_n 0.0205021f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.9
cc_5 VNB N_GATE_M1025_g 0.0240981f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.99
cc_6 VNB GATE 0.0059014f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_7 VNB N_A_354_105#_c_231_n 0.0310136f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_354_105#_c_232_n 0.0221071f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.62
cc_9 VNB N_A_354_105#_M1016_g 0.0437828f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_354_105#_c_234_n 0.00699887f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_354_105#_c_235_n 8.06639e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_354_105#_c_236_n 6.67232e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_354_105#_c_237_n 0.00206511f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_354_105#_c_238_n 0.00282247f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_354_105#_c_239_n 0.00353693f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_324_79#_c_310_n 0.0191913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_324_79#_c_311_n 0.0223453f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.62
cc_18 VNB N_A_324_79#_c_312_n 0.0128593f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.62
cc_19 VNB N_A_324_79#_c_313_n 0.0111492f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.62
cc_20 VNB N_A_324_79#_c_314_n 0.0422786f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_324_79#_c_315_n 0.0210931f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_324_79#_c_316_n 0.00491788f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_324_79#_c_317_n 0.00525298f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_324_79#_c_318_n 0.00566241f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_324_79#_c_319_n 0.00487706f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_324_79#_c_320_n 0.00149564f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_324_79#_c_321_n 0.0141001f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_324_79#_c_322_n 0.00262393f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_324_79#_c_323_n 0.0149264f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_324_79#_c_324_n 0.00222644f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_324_79#_c_325_n 0.00452749f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_324_79#_c_326_n 0.0121301f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_324_79#_c_327_n 0.0019697f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_324_79#_c_328_n 0.0569887f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_792_48#_M1005_g 0.0571831f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_792_48#_M1008_g 0.0248678f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_792_48#_c_476_n 0.0390916f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_792_48#_c_477_n 0.00941361f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_792_48#_c_478_n 0.0157893f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_792_48#_c_479_n 0.00166024f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_792_48#_c_480_n 0.00395206f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_792_48#_c_481_n 0.0115308f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_634_74#_c_601_n 0.0407121f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_634_74#_c_602_n 0.0228989f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.62
cc_45 VNB N_A_634_74#_c_603_n 0.00321093f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_634_74#_c_604_n 0.00131206f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_634_74#_c_605_n 0.0213092f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_634_74#_c_606_n 0.0035258f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_634_74#_c_607_n 0.00692367f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_634_74#_c_608_n 0.00462435f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_CLK_c_676_n 0.0200962f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.455
cc_52 VNB N_CLK_c_677_n 0.0171643f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.62
cc_53 VNB CLK 0.0075037f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.62
cc_54 VNB N_CLK_c_679_n 0.0624119f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_1289_368#_M1001_g 0.0233521f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.62
cc_56 VNB N_A_1289_368#_M1013_g 0.0209649f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_1289_368#_M1026_g 0.0202297f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_1289_368#_M1027_g 0.0260342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_1289_368#_c_733_n 0.00912363f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_1289_368#_c_734_n 0.0130086f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_1289_368#_c_735_n 0.00269775f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_1289_368#_c_736_n 0.00378119f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_1289_368#_c_737_n 2.98518e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_1289_368#_c_738_n 0.00266677f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_1289_368#_c_739_n 0.140872f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VPWR_c_852_n 0.40251f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_119_143#_c_960_n 0.00958489f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_119_143#_c_961_n 8.44192e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_119_143#_c_962_n 0.00496514f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_119_143#_c_963_n 0.00458561f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_119_143#_c_964_n 0.0096811f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_119_143#_c_965_n 0.00838916f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_GCLK_c_1053_n 0.00254365f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_GCLK_c_1054_n 0.00351355f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_GCLK_c_1055_n 0.00205014f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_GCLK_c_1056_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_GCLK_c_1057_n 5.71281e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1124_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1125_n 0.067074f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1126_n 0.0192463f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1127_n 0.00644324f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1128_n 0.00600048f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1129_n 0.0126279f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1130_n 0.00503707f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1131_n 0.010678f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1132_n 0.0505914f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1133_n 0.0643337f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1134_n 0.00617641f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1135_n 0.0380624f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1136_n 0.00615422f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_VGND_c_1137_n 0.0306291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_VGND_c_1138_n 0.0188435f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_VGND_c_1139_n 0.0193312f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_VGND_c_1140_n 0.028177f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_VGND_c_1141_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_VGND_c_1142_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_VGND_c_1143_n 0.535277f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VPB N_SCE_c_177_n 0.0444948f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.9
cc_99 VPB N_SCE_c_179_n 0.00565041f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.62
cc_100 VPB N_GATE_c_200_n 0.0388525f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.9
cc_101 VPB GATE 0.00348266f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_102 VPB N_A_354_105#_c_231_n 0.0432382f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 VPB N_A_354_105#_c_235_n 0.00167859f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB N_A_354_105#_c_236_n 0.00497365f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_105 VPB N_A_354_105#_c_243_n 0.00939143f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_A_354_105#_c_237_n 0.00371457f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB N_A_354_105#_c_238_n 6.44492e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_A_354_105#_c_239_n 0.00276779f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_109 VPB N_A_324_79#_c_313_n 0.0210657f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.62
cc_110 VPB N_A_324_79#_c_330_n 0.00701885f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_A_324_79#_M1002_g 0.0115828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_A_324_79#_c_332_n 0.125911f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_A_324_79#_c_333_n 0.0177831f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_A_324_79#_c_334_n 0.00733369f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_A_324_79#_c_335_n 0.0201791f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_A_324_79#_c_336_n 0.0198855f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_A_324_79#_c_337_n 0.00712381f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_A_324_79#_c_326_n 0.00304161f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_A_792_48#_c_482_n 0.0142562f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.62
cc_120 VPB N_A_792_48#_c_483_n 0.0237354f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.62
cc_121 VPB N_A_792_48#_c_476_n 0.0248549f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_A_792_48#_c_485_n 0.00631684f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_A_792_48#_c_486_n 0.00453835f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_A_792_48#_c_487_n 0.0140467f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_A_792_48#_c_477_n 0.00315593f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 VPB N_A_792_48#_c_489_n 0.0136815f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_127 VPB N_A_792_48#_c_490_n 0.00153807f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_A_792_48#_c_479_n 0.00816786f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_129 VPB N_A_792_48#_c_492_n 0.00440389f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_A_792_48#_c_493_n 5.03018e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_A_792_48#_c_481_n 0.0339709f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_A_634_74#_c_601_n 0.0269006f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_A_634_74#_c_604_n 0.0133562f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_CLK_c_680_n 0.0178774f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.9
cc_135 VPB N_CLK_c_681_n 0.0179379f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_CLK_c_679_n 0.0151637f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_A_1289_368#_c_740_n 0.0160835f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_A_1289_368#_c_741_n 0.016534f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_A_1289_368#_c_742_n 0.0159508f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_140 VPB N_A_1289_368#_c_743_n 0.019062f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_141 VPB N_A_1289_368#_c_744_n 0.00294323f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_142 VPB N_A_1289_368#_c_745_n 0.0040656f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_143 VPB N_A_1289_368#_c_746_n 0.00256539f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_144 VPB N_A_1289_368#_c_737_n 0.00143542f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_145 VPB N_A_1289_368#_c_739_n 0.0310227f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_146 VPB N_VPWR_c_853_n 0.0121909f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_147 VPB N_VPWR_c_854_n 0.0573835f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_148 VPB N_VPWR_c_855_n 0.0185947f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_149 VPB N_VPWR_c_856_n 0.0171686f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_150 VPB N_VPWR_c_857_n 0.00651803f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_151 VPB N_VPWR_c_858_n 0.0082016f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_152 VPB N_VPWR_c_859_n 0.0120152f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_153 VPB N_VPWR_c_860_n 0.0655155f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_154 VPB N_VPWR_c_861_n 0.023151f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_155 VPB N_VPWR_c_862_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_156 VPB N_VPWR_c_863_n 0.0330329f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_157 VPB N_VPWR_c_864_n 0.0681025f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_158 VPB N_VPWR_c_865_n 0.0387399f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_159 VPB N_VPWR_c_866_n 0.0220372f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_160 VPB N_VPWR_c_867_n 0.0185368f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_161 VPB N_VPWR_c_868_n 0.0264441f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_162 VPB N_VPWR_c_869_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_163 VPB N_VPWR_c_870_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_164 VPB N_VPWR_c_871_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_165 VPB N_VPWR_c_852_n 0.145038f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_166 VPB N_A_119_143#_c_963_n 0.00860465f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_167 VPB N_A_119_143#_c_967_n 0.0142941f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_168 VPB N_A_119_143#_c_968_n 0.00501274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_169 VPB N_A_119_143#_c_969_n 0.0120112f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_170 VPB N_A_119_143#_c_970_n 0.0226979f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_171 VPB N_GCLK_c_1058_n 0.00292742f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_172 VPB N_GCLK_c_1059_n 0.00234449f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_173 VPB N_GCLK_c_1060_n 0.00230768f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_174 VPB N_GCLK_c_1061_n 0.00289698f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_175 VPB N_GCLK_c_1057_n 0.00264854f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_176 VPB N_GCLK_c_1063_n 9.51973e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_177 N_SCE_c_177_n N_GATE_c_200_n 0.0700752f $X=0.505 $Y=1.9 $X2=-0.19
+ $Y2=-0.245
cc_178 N_SCE_c_179_n N_GATE_c_200_n 3.90315e-19 $X=0.385 $Y=1.62 $X2=-0.19
+ $Y2=-0.245
cc_179 N_SCE_M1019_g N_GATE_M1025_g 0.0177982f $X=0.52 $Y=0.99 $X2=0 $Y2=0
cc_180 N_SCE_c_177_n GATE 0.00127121f $X=0.505 $Y=1.9 $X2=0 $Y2=0
cc_181 N_SCE_c_179_n GATE 0.0171967f $X=0.385 $Y=1.62 $X2=0 $Y2=0
cc_182 N_SCE_c_177_n N_VPWR_c_854_n 0.0285041f $X=0.505 $Y=1.9 $X2=0 $Y2=0
cc_183 N_SCE_c_179_n N_VPWR_c_854_n 0.0272312f $X=0.385 $Y=1.62 $X2=0 $Y2=0
cc_184 N_SCE_c_177_n N_VPWR_c_863_n 0.00429349f $X=0.505 $Y=1.9 $X2=0 $Y2=0
cc_185 N_SCE_c_177_n N_VPWR_c_852_n 0.00454161f $X=0.505 $Y=1.9 $X2=0 $Y2=0
cc_186 N_SCE_M1019_g N_A_119_143#_c_960_n 6.33101e-19 $X=0.52 $Y=0.99 $X2=0
+ $Y2=0
cc_187 N_SCE_M1019_g N_A_119_143#_c_962_n 0.00128972f $X=0.52 $Y=0.99 $X2=0
+ $Y2=0
cc_188 N_SCE_c_177_n N_A_119_143#_c_969_n 0.00102434f $X=0.505 $Y=1.9 $X2=0
+ $Y2=0
cc_189 N_SCE_c_177_n N_A_119_143#_c_970_n 0.00150385f $X=0.505 $Y=1.9 $X2=0
+ $Y2=0
cc_190 N_SCE_c_177_n N_VGND_c_1125_n 0.00529488f $X=0.505 $Y=1.9 $X2=0 $Y2=0
cc_191 N_SCE_M1019_g N_VGND_c_1125_n 0.00746819f $X=0.52 $Y=0.99 $X2=0 $Y2=0
cc_192 N_SCE_c_179_n N_VGND_c_1125_n 0.0272945f $X=0.385 $Y=1.62 $X2=0 $Y2=0
cc_193 N_SCE_M1019_g N_VGND_c_1126_n 0.00370133f $X=0.52 $Y=0.99 $X2=0 $Y2=0
cc_194 N_SCE_M1019_g N_VGND_c_1143_n 0.00445256f $X=0.52 $Y=0.99 $X2=0 $Y2=0
cc_195 N_GATE_M1025_g N_A_324_79#_c_310_n 0.0141001f $X=0.995 $Y=0.99 $X2=0
+ $Y2=0
cc_196 N_GATE_c_200_n N_A_324_79#_c_312_n 8.07007e-19 $X=0.925 $Y=1.9 $X2=0
+ $Y2=0
cc_197 N_GATE_c_200_n N_VPWR_c_854_n 0.00307102f $X=0.925 $Y=1.9 $X2=0 $Y2=0
cc_198 N_GATE_c_200_n N_VPWR_c_863_n 0.00466857f $X=0.925 $Y=1.9 $X2=0 $Y2=0
cc_199 N_GATE_c_200_n N_VPWR_c_868_n 0.00339632f $X=0.925 $Y=1.9 $X2=0 $Y2=0
cc_200 N_GATE_c_200_n N_VPWR_c_852_n 0.00500913f $X=0.925 $Y=1.9 $X2=0 $Y2=0
cc_201 N_GATE_c_200_n N_A_119_143#_c_960_n 0.00227344f $X=0.925 $Y=1.9 $X2=0
+ $Y2=0
cc_202 N_GATE_M1025_g N_A_119_143#_c_960_n 0.0109495f $X=0.995 $Y=0.99 $X2=0
+ $Y2=0
cc_203 GATE N_A_119_143#_c_960_n 0.00907303f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_204 N_GATE_c_200_n N_A_119_143#_c_961_n 0.00126549f $X=0.925 $Y=1.9 $X2=0
+ $Y2=0
cc_205 N_GATE_M1025_g N_A_119_143#_c_961_n 0.0103937f $X=0.995 $Y=0.99 $X2=0
+ $Y2=0
cc_206 GATE N_A_119_143#_c_961_n 0.00878437f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_207 N_GATE_M1025_g N_A_119_143#_c_962_n 0.00269077f $X=0.995 $Y=0.99 $X2=0
+ $Y2=0
cc_208 N_GATE_c_200_n N_A_119_143#_c_963_n 0.00579166f $X=0.925 $Y=1.9 $X2=0
+ $Y2=0
cc_209 N_GATE_M1025_g N_A_119_143#_c_963_n 0.00678895f $X=0.995 $Y=0.99 $X2=0
+ $Y2=0
cc_210 GATE N_A_119_143#_c_963_n 0.0269205f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_211 N_GATE_c_200_n N_A_119_143#_c_969_n 0.00660871f $X=0.925 $Y=1.9 $X2=0
+ $Y2=0
cc_212 N_GATE_c_200_n N_A_119_143#_c_970_n 0.0175885f $X=0.925 $Y=1.9 $X2=0
+ $Y2=0
cc_213 GATE N_A_119_143#_c_970_n 0.0276683f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_214 N_GATE_M1025_g N_VGND_c_1126_n 0.00287494f $X=0.995 $Y=0.99 $X2=0 $Y2=0
cc_215 N_GATE_M1025_g N_VGND_c_1143_n 0.00445256f $X=0.995 $Y=0.99 $X2=0 $Y2=0
cc_216 N_A_354_105#_c_234_n N_A_324_79#_c_310_n 6.11846e-19 $X=1.91 $Y=1.12
+ $X2=0 $Y2=0
cc_217 N_A_354_105#_c_234_n N_A_324_79#_c_311_n 0.0190885f $X=1.91 $Y=1.12 $X2=0
+ $Y2=0
cc_218 N_A_354_105#_c_235_n N_A_324_79#_c_311_n 0.00248561f $X=2.365 $Y=1.65
+ $X2=0 $Y2=0
cc_219 N_A_354_105#_c_231_n N_A_324_79#_c_313_n 0.00395101f $X=3.315 $Y=1.82
+ $X2=0 $Y2=0
cc_220 N_A_354_105#_c_234_n N_A_324_79#_c_313_n 0.00306741f $X=1.91 $Y=1.12
+ $X2=0 $Y2=0
cc_221 N_A_354_105#_c_235_n N_A_324_79#_c_313_n 0.0199296f $X=2.365 $Y=1.65
+ $X2=0 $Y2=0
cc_222 N_A_354_105#_c_243_n N_A_324_79#_c_313_n 0.0132457f $X=2.53 $Y=1.975
+ $X2=0 $Y2=0
cc_223 N_A_354_105#_c_239_n N_A_324_79#_c_313_n 4.73487e-19 $X=3.09 $Y=1.57
+ $X2=0 $Y2=0
cc_224 N_A_354_105#_c_243_n N_A_324_79#_M1002_g 0.00391084f $X=2.53 $Y=1.975
+ $X2=0 $Y2=0
cc_225 N_A_354_105#_c_231_n N_A_324_79#_c_332_n 0.0103438f $X=3.315 $Y=1.82
+ $X2=0 $Y2=0
cc_226 N_A_354_105#_c_231_n N_A_324_79#_c_314_n 0.015893f $X=3.315 $Y=1.82 $X2=0
+ $Y2=0
cc_227 N_A_354_105#_c_237_n N_A_324_79#_c_314_n 0.00132308f $X=2.925 $Y=1.65
+ $X2=0 $Y2=0
cc_228 N_A_354_105#_c_238_n N_A_324_79#_c_314_n 7.91151e-19 $X=2.53 $Y=1.65
+ $X2=0 $Y2=0
cc_229 N_A_354_105#_c_239_n N_A_324_79#_c_314_n 0.00143623f $X=3.09 $Y=1.57
+ $X2=0 $Y2=0
cc_230 N_A_354_105#_M1016_g N_A_324_79#_c_315_n 0.0217463f $X=3.645 $Y=0.58
+ $X2=0 $Y2=0
cc_231 N_A_354_105#_c_231_n N_A_324_79#_c_334_n 0.00378299f $X=3.315 $Y=1.82
+ $X2=0 $Y2=0
cc_232 N_A_354_105#_c_231_n N_A_324_79#_c_336_n 0.0088366f $X=3.315 $Y=1.82
+ $X2=0 $Y2=0
cc_233 N_A_354_105#_M1016_g N_A_324_79#_c_316_n 3.16786e-19 $X=3.645 $Y=0.58
+ $X2=0 $Y2=0
cc_234 N_A_354_105#_c_237_n N_A_324_79#_c_316_n 0.0115741f $X=2.925 $Y=1.65
+ $X2=0 $Y2=0
cc_235 N_A_354_105#_c_238_n N_A_324_79#_c_316_n 0.0063017f $X=2.53 $Y=1.65 $X2=0
+ $Y2=0
cc_236 N_A_354_105#_c_239_n N_A_324_79#_c_316_n 0.00415249f $X=3.09 $Y=1.57
+ $X2=0 $Y2=0
cc_237 N_A_354_105#_M1016_g N_A_324_79#_c_318_n 0.0129965f $X=3.645 $Y=0.58
+ $X2=0 $Y2=0
cc_238 N_A_354_105#_M1016_g N_A_324_79#_c_320_n 0.00199569f $X=3.645 $Y=0.58
+ $X2=0 $Y2=0
cc_239 N_A_354_105#_M1016_g N_A_324_79#_c_322_n 0.00133148f $X=3.645 $Y=0.58
+ $X2=0 $Y2=0
cc_240 N_A_354_105#_c_234_n N_A_324_79#_c_365_n 0.0253307f $X=1.91 $Y=1.12 $X2=0
+ $Y2=0
cc_241 N_A_354_105#_c_235_n N_A_324_79#_c_365_n 0.00871007f $X=2.365 $Y=1.65
+ $X2=0 $Y2=0
cc_242 N_A_354_105#_c_238_n N_A_324_79#_c_365_n 0.0174669f $X=2.53 $Y=1.65 $X2=0
+ $Y2=0
cc_243 N_A_354_105#_c_231_n N_A_324_79#_c_328_n 0.00379557f $X=3.315 $Y=1.82
+ $X2=0 $Y2=0
cc_244 N_A_354_105#_c_234_n N_A_324_79#_c_328_n 0.00335921f $X=1.91 $Y=1.12
+ $X2=0 $Y2=0
cc_245 N_A_354_105#_c_235_n N_A_324_79#_c_328_n 0.00146387f $X=2.365 $Y=1.65
+ $X2=0 $Y2=0
cc_246 N_A_354_105#_c_238_n N_A_324_79#_c_328_n 0.00579073f $X=2.53 $Y=1.65
+ $X2=0 $Y2=0
cc_247 N_A_354_105#_c_239_n N_A_324_79#_c_328_n 6.1217e-19 $X=3.09 $Y=1.57 $X2=0
+ $Y2=0
cc_248 N_A_354_105#_c_231_n N_A_792_48#_M1005_g 0.00383961f $X=3.315 $Y=1.82
+ $X2=0 $Y2=0
cc_249 N_A_354_105#_M1016_g N_A_792_48#_M1005_g 0.0653275f $X=3.645 $Y=0.58
+ $X2=0 $Y2=0
cc_250 N_A_354_105#_c_231_n N_A_792_48#_c_481_n 0.00105613f $X=3.315 $Y=1.82
+ $X2=0 $Y2=0
cc_251 N_A_354_105#_M1016_g N_A_634_74#_c_603_n 0.00730232f $X=3.645 $Y=0.58
+ $X2=0 $Y2=0
cc_252 N_A_354_105#_c_231_n N_A_634_74#_c_604_n 0.00830893f $X=3.315 $Y=1.82
+ $X2=0 $Y2=0
cc_253 N_A_354_105#_c_232_n N_A_634_74#_c_604_n 0.0147699f $X=3.57 $Y=1.48 $X2=0
+ $Y2=0
cc_254 N_A_354_105#_c_239_n N_A_634_74#_c_604_n 0.0251391f $X=3.09 $Y=1.57 $X2=0
+ $Y2=0
cc_255 N_A_354_105#_M1016_g N_A_634_74#_c_605_n 0.00308854f $X=3.645 $Y=0.58
+ $X2=0 $Y2=0
cc_256 N_A_354_105#_c_231_n N_A_634_74#_c_606_n 0.00594497f $X=3.315 $Y=1.82
+ $X2=0 $Y2=0
cc_257 N_A_354_105#_c_232_n N_A_634_74#_c_606_n 3.55064e-19 $X=3.57 $Y=1.48
+ $X2=0 $Y2=0
cc_258 N_A_354_105#_M1016_g N_A_634_74#_c_606_n 0.00876954f $X=3.645 $Y=0.58
+ $X2=0 $Y2=0
cc_259 N_A_354_105#_c_239_n N_A_634_74#_c_606_n 0.00397264f $X=3.09 $Y=1.57
+ $X2=0 $Y2=0
cc_260 N_A_354_105#_c_232_n N_A_634_74#_c_607_n 0.00317399f $X=3.57 $Y=1.48
+ $X2=0 $Y2=0
cc_261 N_A_354_105#_M1016_g N_A_634_74#_c_607_n 0.0107752f $X=3.645 $Y=0.58
+ $X2=0 $Y2=0
cc_262 N_A_354_105#_c_231_n N_VPWR_c_852_n 9.39239e-19 $X=3.315 $Y=1.82 $X2=0
+ $Y2=0
cc_263 N_A_354_105#_c_234_n N_A_119_143#_c_963_n 0.0322212f $X=1.91 $Y=1.12
+ $X2=0 $Y2=0
cc_264 N_A_354_105#_c_236_n N_A_119_143#_c_963_n 0.0143581f $X=2.075 $Y=1.65
+ $X2=0 $Y2=0
cc_265 N_A_354_105#_M1002_d N_A_119_143#_c_967_n 0.00826344f $X=2.295 $Y=2.12
+ $X2=0 $Y2=0
cc_266 N_A_354_105#_c_231_n N_A_119_143#_c_967_n 0.00691199f $X=3.315 $Y=1.82
+ $X2=0 $Y2=0
cc_267 N_A_354_105#_c_235_n N_A_119_143#_c_967_n 0.00622309f $X=2.365 $Y=1.65
+ $X2=0 $Y2=0
cc_268 N_A_354_105#_c_236_n N_A_119_143#_c_967_n 0.00865555f $X=2.075 $Y=1.65
+ $X2=0 $Y2=0
cc_269 N_A_354_105#_c_243_n N_A_119_143#_c_967_n 0.0263817f $X=2.53 $Y=1.975
+ $X2=0 $Y2=0
cc_270 N_A_354_105#_c_237_n N_A_119_143#_c_967_n 0.00740026f $X=2.925 $Y=1.65
+ $X2=0 $Y2=0
cc_271 N_A_354_105#_c_231_n N_A_119_143#_c_968_n 0.00728875f $X=3.315 $Y=1.82
+ $X2=0 $Y2=0
cc_272 N_A_354_105#_c_243_n N_A_119_143#_c_968_n 0.0158435f $X=2.53 $Y=1.975
+ $X2=0 $Y2=0
cc_273 N_A_354_105#_c_239_n N_A_119_143#_c_968_n 0.0246052f $X=3.09 $Y=1.57
+ $X2=0 $Y2=0
cc_274 N_A_354_105#_M1017_d N_A_119_143#_c_965_n 0.00709289f $X=1.77 $Y=0.525
+ $X2=0 $Y2=0
cc_275 N_A_354_105#_c_234_n N_A_119_143#_c_965_n 0.0201545f $X=1.91 $Y=1.12
+ $X2=0 $Y2=0
cc_276 N_A_354_105#_M1016_g N_VGND_c_1127_n 3.67768e-19 $X=3.645 $Y=0.58 $X2=0
+ $Y2=0
cc_277 N_A_354_105#_M1016_g N_VGND_c_1133_n 0.00280452f $X=3.645 $Y=0.58 $X2=0
+ $Y2=0
cc_278 N_A_354_105#_M1016_g N_VGND_c_1143_n 0.00354535f $X=3.645 $Y=0.58 $X2=0
+ $Y2=0
cc_279 N_A_324_79#_c_323_n N_A_792_48#_M1004_d 0.00273752f $X=5.445 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_280 N_A_324_79#_c_318_n N_A_792_48#_M1005_g 0.00107336f $X=3.765 $Y=0.355
+ $X2=0 $Y2=0
cc_281 N_A_324_79#_c_320_n N_A_792_48#_M1005_g 0.00274065f $X=3.85 $Y=0.895
+ $X2=0 $Y2=0
cc_282 N_A_324_79#_c_321_n N_A_792_48#_M1005_g 0.0153072f $X=4.605 $Y=0.98 $X2=0
+ $Y2=0
cc_283 N_A_324_79#_c_377_p N_A_792_48#_M1005_g 0.00137341f $X=4.69 $Y=0.895
+ $X2=0 $Y2=0
cc_284 N_A_324_79#_c_324_n N_A_792_48#_M1005_g 3.77334e-19 $X=4.775 $Y=0.34
+ $X2=0 $Y2=0
cc_285 N_A_324_79#_c_334_n N_A_792_48#_c_483_n 0.00285538f $X=3.85 $Y=2.86 $X2=0
+ $Y2=0
cc_286 N_A_324_79#_c_336_n N_A_792_48#_c_483_n 0.0277971f $X=3.85 $Y=2.77 $X2=0
+ $Y2=0
cc_287 N_A_324_79#_c_337_n N_A_792_48#_c_486_n 0.013888f $X=5.605 $Y=1.985 $X2=0
+ $Y2=0
cc_288 N_A_324_79#_c_326_n N_A_792_48#_c_477_n 0.0502011f $X=5.607 $Y=1.82 $X2=0
+ $Y2=0
cc_289 N_A_324_79#_M1023_s N_A_792_48#_c_489_n 0.0129708f $X=5.46 $Y=1.84 $X2=0
+ $Y2=0
cc_290 N_A_324_79#_c_337_n N_A_792_48#_c_489_n 0.0217771f $X=5.605 $Y=1.985
+ $X2=0 $Y2=0
cc_291 N_A_324_79#_c_337_n N_A_792_48#_c_490_n 0.00416741f $X=5.605 $Y=1.985
+ $X2=0 $Y2=0
cc_292 N_A_324_79#_c_326_n N_A_792_48#_c_490_n 0.00349637f $X=5.607 $Y=1.82
+ $X2=0 $Y2=0
cc_293 N_A_324_79#_c_326_n N_A_792_48#_c_512_n 0.00220044f $X=5.607 $Y=1.82
+ $X2=0 $Y2=0
cc_294 N_A_324_79#_c_337_n N_A_792_48#_c_492_n 0.00752722f $X=5.605 $Y=1.985
+ $X2=0 $Y2=0
cc_295 N_A_324_79#_c_326_n N_A_792_48#_c_492_n 0.0074203f $X=5.607 $Y=1.82 $X2=0
+ $Y2=0
cc_296 N_A_324_79#_c_323_n N_A_792_48#_c_480_n 0.0203619f $X=5.445 $Y=0.34 $X2=0
+ $Y2=0
cc_297 N_A_324_79#_c_325_n N_A_792_48#_c_480_n 0.0397103f $X=5.67 $Y=0.515 $X2=0
+ $Y2=0
cc_298 N_A_324_79#_c_318_n N_A_634_74#_M1022_d 0.00320041f $X=3.765 $Y=0.355
+ $X2=-0.19 $Y2=-0.245
cc_299 N_A_324_79#_c_321_n N_A_634_74#_c_601_n 0.00130576f $X=4.605 $Y=0.98
+ $X2=0 $Y2=0
cc_300 N_A_324_79#_c_326_n N_A_634_74#_c_601_n 7.88608e-19 $X=5.607 $Y=1.82
+ $X2=0 $Y2=0
cc_301 N_A_324_79#_c_323_n N_A_634_74#_c_602_n 0.0156771f $X=5.445 $Y=0.34 $X2=0
+ $Y2=0
cc_302 N_A_324_79#_c_325_n N_A_634_74#_c_602_n 0.00385526f $X=5.67 $Y=0.515
+ $X2=0 $Y2=0
cc_303 N_A_324_79#_c_326_n N_A_634_74#_c_602_n 0.00125296f $X=5.607 $Y=1.82
+ $X2=0 $Y2=0
cc_304 N_A_324_79#_c_315_n N_A_634_74#_c_603_n 0.00236682f $X=3.095 $Y=1.045
+ $X2=0 $Y2=0
cc_305 N_A_324_79#_c_316_n N_A_634_74#_c_603_n 0.00641233f $X=2.805 $Y=1.15
+ $X2=0 $Y2=0
cc_306 N_A_324_79#_c_317_n N_A_634_74#_c_603_n 0.00468717f $X=2.89 $Y=1.065
+ $X2=0 $Y2=0
cc_307 N_A_324_79#_c_322_n N_A_634_74#_c_603_n 0.0100839f $X=3.935 $Y=0.98 $X2=0
+ $Y2=0
cc_308 N_A_324_79#_c_332_n N_A_634_74#_c_604_n 0.00564711f $X=3.76 $Y=3.15 $X2=0
+ $Y2=0
cc_309 N_A_324_79#_c_336_n N_A_634_74#_c_604_n 0.0165071f $X=3.85 $Y=2.77 $X2=0
+ $Y2=0
cc_310 N_A_324_79#_c_321_n N_A_634_74#_c_605_n 0.0488693f $X=4.605 $Y=0.98 $X2=0
+ $Y2=0
cc_311 N_A_324_79#_c_322_n N_A_634_74#_c_605_n 0.0143583f $X=3.935 $Y=0.98 $X2=0
+ $Y2=0
cc_312 N_A_324_79#_c_315_n N_A_634_74#_c_606_n 0.00454113f $X=3.095 $Y=1.045
+ $X2=0 $Y2=0
cc_313 N_A_324_79#_c_317_n N_A_634_74#_c_606_n 0.0136555f $X=2.89 $Y=1.065 $X2=0
+ $Y2=0
cc_314 N_A_324_79#_c_318_n N_A_634_74#_c_606_n 0.0238927f $X=3.765 $Y=0.355
+ $X2=0 $Y2=0
cc_315 N_A_324_79#_c_320_n N_A_634_74#_c_606_n 0.0151262f $X=3.85 $Y=0.895 $X2=0
+ $Y2=0
cc_316 N_A_324_79#_c_322_n N_A_634_74#_c_606_n 0.00380883f $X=3.935 $Y=0.98
+ $X2=0 $Y2=0
cc_317 N_A_324_79#_c_321_n N_A_634_74#_c_608_n 0.0135682f $X=4.605 $Y=0.98 $X2=0
+ $Y2=0
cc_318 N_A_324_79#_c_337_n N_CLK_c_680_n 0.00541719f $X=5.605 $Y=1.985 $X2=-0.19
+ $Y2=-0.245
cc_319 N_A_324_79#_c_323_n N_CLK_c_676_n 0.00462516f $X=5.445 $Y=0.34 $X2=0
+ $Y2=0
cc_320 N_A_324_79#_c_325_n N_CLK_c_676_n 0.0043874f $X=5.67 $Y=0.515 $X2=0 $Y2=0
cc_321 N_A_324_79#_c_326_n N_CLK_c_676_n 0.00343873f $X=5.607 $Y=1.82 $X2=0
+ $Y2=0
cc_322 N_A_324_79#_c_327_n N_CLK_c_676_n 0.00232496f $X=5.64 $Y=1.01 $X2=0 $Y2=0
cc_323 N_A_324_79#_c_337_n N_CLK_c_681_n 2.55992e-19 $X=5.605 $Y=1.985 $X2=0
+ $Y2=0
cc_324 N_A_324_79#_c_326_n CLK 0.0279712f $X=5.607 $Y=1.82 $X2=0 $Y2=0
cc_325 N_A_324_79#_c_327_n CLK 0.0029255f $X=5.64 $Y=1.01 $X2=0 $Y2=0
cc_326 N_A_324_79#_c_337_n N_CLK_c_679_n 7.09264e-19 $X=5.605 $Y=1.985 $X2=0
+ $Y2=0
cc_327 N_A_324_79#_c_326_n N_CLK_c_679_n 0.0147013f $X=5.607 $Y=1.82 $X2=0 $Y2=0
cc_328 N_A_324_79#_c_327_n N_CLK_c_679_n 0.00111406f $X=5.64 $Y=1.01 $X2=0 $Y2=0
cc_329 N_A_324_79#_c_334_n N_VPWR_c_855_n 0.00935475f $X=3.85 $Y=2.86 $X2=0
+ $Y2=0
cc_330 N_A_324_79#_c_333_n N_VPWR_c_864_n 0.0570707f $X=2.31 $Y=3.15 $X2=0 $Y2=0
cc_331 N_A_324_79#_M1002_g N_VPWR_c_868_n 0.0194226f $X=2.22 $Y=2.54 $X2=0 $Y2=0
cc_332 N_A_324_79#_c_333_n N_VPWR_c_868_n 0.0114039f $X=2.31 $Y=3.15 $X2=0 $Y2=0
cc_333 N_A_324_79#_c_332_n N_VPWR_c_852_n 0.0566411f $X=3.76 $Y=3.15 $X2=0 $Y2=0
cc_334 N_A_324_79#_c_333_n N_VPWR_c_852_n 0.00455307f $X=2.31 $Y=3.15 $X2=0
+ $Y2=0
cc_335 N_A_324_79#_c_317_n N_A_119_143#_M1022_s 0.00828024f $X=2.89 $Y=1.065
+ $X2=0 $Y2=0
cc_336 N_A_324_79#_c_319_n N_A_119_143#_M1022_s 9.10245e-19 $X=2.975 $Y=0.355
+ $X2=0 $Y2=0
cc_337 N_A_324_79#_c_310_n N_A_119_143#_c_960_n 4.34451e-19 $X=1.695 $Y=1.34
+ $X2=0 $Y2=0
cc_338 N_A_324_79#_c_310_n N_A_119_143#_c_963_n 0.0157986f $X=1.695 $Y=1.34
+ $X2=0 $Y2=0
cc_339 N_A_324_79#_c_312_n N_A_119_143#_c_963_n 0.005009f $X=1.77 $Y=1.415 $X2=0
+ $Y2=0
cc_340 N_A_324_79#_c_313_n N_A_119_143#_c_963_n 0.00630379f $X=2.22 $Y=1.955
+ $X2=0 $Y2=0
cc_341 N_A_324_79#_M1002_g N_A_119_143#_c_967_n 0.0243094f $X=2.22 $Y=2.54 $X2=0
+ $Y2=0
cc_342 N_A_324_79#_c_332_n N_A_119_143#_c_967_n 0.0194918f $X=3.76 $Y=3.15 $X2=0
+ $Y2=0
cc_343 N_A_324_79#_M1002_g N_A_119_143#_c_968_n 0.00404627f $X=2.22 $Y=2.54
+ $X2=0 $Y2=0
cc_344 N_A_324_79#_c_330_n N_A_119_143#_c_970_n 0.00267593f $X=2.22 $Y=2.045
+ $X2=0 $Y2=0
cc_345 N_A_324_79#_M1002_g N_A_119_143#_c_970_n 0.0076987f $X=2.22 $Y=2.54 $X2=0
+ $Y2=0
cc_346 N_A_324_79#_c_310_n N_A_119_143#_c_1012_n 0.00435069f $X=1.695 $Y=1.34
+ $X2=0 $Y2=0
cc_347 N_A_324_79#_c_310_n N_A_119_143#_c_964_n 0.00731619f $X=1.695 $Y=1.34
+ $X2=0 $Y2=0
cc_348 N_A_324_79#_c_315_n N_A_119_143#_c_964_n 0.00124433f $X=3.095 $Y=1.045
+ $X2=0 $Y2=0
cc_349 N_A_324_79#_c_316_n N_A_119_143#_c_964_n 0.00459251f $X=2.805 $Y=1.15
+ $X2=0 $Y2=0
cc_350 N_A_324_79#_c_317_n N_A_119_143#_c_964_n 0.0356041f $X=2.89 $Y=1.065
+ $X2=0 $Y2=0
cc_351 N_A_324_79#_c_319_n N_A_119_143#_c_964_n 0.00767896f $X=2.975 $Y=0.355
+ $X2=0 $Y2=0
cc_352 N_A_324_79#_c_365_n N_A_119_143#_c_964_n 0.0218607f $X=2.41 $Y=1.15 $X2=0
+ $Y2=0
cc_353 N_A_324_79#_c_328_n N_A_119_143#_c_964_n 0.00799329f $X=2.352 $Y=1.12
+ $X2=0 $Y2=0
cc_354 N_A_324_79#_c_310_n N_A_119_143#_c_965_n 0.0129997f $X=1.695 $Y=1.34
+ $X2=0 $Y2=0
cc_355 N_A_324_79#_c_311_n N_A_119_143#_c_965_n 5.7542e-19 $X=2.13 $Y=1.415
+ $X2=0 $Y2=0
cc_356 N_A_324_79#_c_365_n N_A_119_143#_c_965_n 0.00303811f $X=2.41 $Y=1.15
+ $X2=0 $Y2=0
cc_357 N_A_324_79#_c_328_n N_A_119_143#_c_965_n 0.00583436f $X=2.352 $Y=1.12
+ $X2=0 $Y2=0
cc_358 N_A_324_79#_c_321_n N_VGND_M1005_d 0.00468885f $X=4.605 $Y=0.98 $X2=0
+ $Y2=0
cc_359 N_A_324_79#_c_377_p N_VGND_M1005_d 0.00845472f $X=4.69 $Y=0.895 $X2=0
+ $Y2=0
cc_360 N_A_324_79#_c_324_n N_VGND_M1005_d 6.47853e-19 $X=4.775 $Y=0.34 $X2=0
+ $Y2=0
cc_361 N_A_324_79#_c_318_n N_VGND_c_1127_n 0.0110244f $X=3.765 $Y=0.355 $X2=0
+ $Y2=0
cc_362 N_A_324_79#_c_321_n N_VGND_c_1127_n 0.0244958f $X=4.605 $Y=0.98 $X2=0
+ $Y2=0
cc_363 N_A_324_79#_c_377_p N_VGND_c_1127_n 0.0228902f $X=4.69 $Y=0.895 $X2=0
+ $Y2=0
cc_364 N_A_324_79#_c_324_n N_VGND_c_1127_n 0.0148567f $X=4.775 $Y=0.34 $X2=0
+ $Y2=0
cc_365 N_A_324_79#_c_323_n N_VGND_c_1128_n 0.011924f $X=5.445 $Y=0.34 $X2=0
+ $Y2=0
cc_366 N_A_324_79#_c_310_n N_VGND_c_1133_n 0.00361406f $X=1.695 $Y=1.34 $X2=0
+ $Y2=0
cc_367 N_A_324_79#_c_315_n N_VGND_c_1133_n 0.00280452f $X=3.095 $Y=1.045 $X2=0
+ $Y2=0
cc_368 N_A_324_79#_c_318_n N_VGND_c_1133_n 0.056759f $X=3.765 $Y=0.355 $X2=0
+ $Y2=0
cc_369 N_A_324_79#_c_319_n N_VGND_c_1133_n 0.0111306f $X=2.975 $Y=0.355 $X2=0
+ $Y2=0
cc_370 N_A_324_79#_c_323_n N_VGND_c_1135_n 0.0705353f $X=5.445 $Y=0.34 $X2=0
+ $Y2=0
cc_371 N_A_324_79#_c_324_n N_VGND_c_1135_n 0.0121867f $X=4.775 $Y=0.34 $X2=0
+ $Y2=0
cc_372 N_A_324_79#_c_310_n N_VGND_c_1140_n 0.00218072f $X=1.695 $Y=1.34 $X2=0
+ $Y2=0
cc_373 N_A_324_79#_c_310_n N_VGND_c_1143_n 0.0049796f $X=1.695 $Y=1.34 $X2=0
+ $Y2=0
cc_374 N_A_324_79#_c_315_n N_VGND_c_1143_n 0.00359824f $X=3.095 $Y=1.045 $X2=0
+ $Y2=0
cc_375 N_A_324_79#_c_318_n N_VGND_c_1143_n 0.0346109f $X=3.765 $Y=0.355 $X2=0
+ $Y2=0
cc_376 N_A_324_79#_c_319_n N_VGND_c_1143_n 0.00656177f $X=2.975 $Y=0.355 $X2=0
+ $Y2=0
cc_377 N_A_324_79#_c_323_n N_VGND_c_1143_n 0.0395478f $X=5.445 $Y=0.34 $X2=0
+ $Y2=0
cc_378 N_A_324_79#_c_324_n N_VGND_c_1143_n 0.00660921f $X=4.775 $Y=0.34 $X2=0
+ $Y2=0
cc_379 N_A_324_79#_c_320_n A_744_74# 7.18336e-19 $X=3.85 $Y=0.895 $X2=-0.19
+ $Y2=-0.245
cc_380 N_A_792_48#_M1005_g N_A_634_74#_c_601_n 0.00800016f $X=4.035 $Y=0.58
+ $X2=0 $Y2=0
cc_381 N_A_792_48#_c_483_n N_A_634_74#_c_601_n 0.00747158f $X=4.27 $Y=2.2 $X2=0
+ $Y2=0
cc_382 N_A_792_48#_c_485_n N_A_634_74#_c_601_n 0.0136986f $X=4.88 $Y=1.82 $X2=0
+ $Y2=0
cc_383 N_A_792_48#_c_486_n N_A_634_74#_c_601_n 0.00550722f $X=5.075 $Y=2.24
+ $X2=0 $Y2=0
cc_384 N_A_792_48#_c_487_n N_A_634_74#_c_601_n 0.00612636f $X=5.045 $Y=2.73
+ $X2=0 $Y2=0
cc_385 N_A_792_48#_c_477_n N_A_634_74#_c_601_n 0.00408252f $X=5.185 $Y=1.735
+ $X2=0 $Y2=0
cc_386 N_A_792_48#_c_479_n N_A_634_74#_c_601_n 9.25858e-19 $X=4.125 $Y=1.74
+ $X2=0 $Y2=0
cc_387 N_A_792_48#_c_492_n N_A_634_74#_c_601_n 0.003104f $X=5.045 $Y=1.9 $X2=0
+ $Y2=0
cc_388 N_A_792_48#_c_493_n N_A_634_74#_c_601_n 0.00176183f $X=5.075 $Y=2.325
+ $X2=0 $Y2=0
cc_389 N_A_792_48#_c_481_n N_A_634_74#_c_601_n 0.0173674f $X=4.27 $Y=1.74 $X2=0
+ $Y2=0
cc_390 N_A_792_48#_M1005_g N_A_634_74#_c_602_n 0.0093121f $X=4.035 $Y=0.58 $X2=0
+ $Y2=0
cc_391 N_A_792_48#_c_477_n N_A_634_74#_c_602_n 0.0122125f $X=5.185 $Y=1.735
+ $X2=0 $Y2=0
cc_392 N_A_792_48#_c_480_n N_A_634_74#_c_602_n 0.00758287f $X=5.11 $Y=0.83 $X2=0
+ $Y2=0
cc_393 N_A_792_48#_M1005_g N_A_634_74#_c_603_n 9.44671e-19 $X=4.035 $Y=0.58
+ $X2=0 $Y2=0
cc_394 N_A_792_48#_M1005_g N_A_634_74#_c_604_n 0.00451039f $X=4.035 $Y=0.58
+ $X2=0 $Y2=0
cc_395 N_A_792_48#_c_482_n N_A_634_74#_c_604_n 0.00653088f $X=4.27 $Y=2.11 $X2=0
+ $Y2=0
cc_396 N_A_792_48#_c_479_n N_A_634_74#_c_604_n 0.0190551f $X=4.125 $Y=1.74 $X2=0
+ $Y2=0
cc_397 N_A_792_48#_M1005_g N_A_634_74#_c_605_n 0.0109782f $X=4.035 $Y=0.58 $X2=0
+ $Y2=0
cc_398 N_A_792_48#_c_485_n N_A_634_74#_c_605_n 0.0144756f $X=4.88 $Y=1.82 $X2=0
+ $Y2=0
cc_399 N_A_792_48#_c_479_n N_A_634_74#_c_605_n 0.0242156f $X=4.125 $Y=1.74 $X2=0
+ $Y2=0
cc_400 N_A_792_48#_c_481_n N_A_634_74#_c_605_n 0.00325243f $X=4.27 $Y=1.74 $X2=0
+ $Y2=0
cc_401 N_A_792_48#_M1005_g N_A_634_74#_c_608_n 9.69453e-19 $X=4.035 $Y=0.58
+ $X2=0 $Y2=0
cc_402 N_A_792_48#_c_485_n N_A_634_74#_c_608_n 0.0205329f $X=4.88 $Y=1.82 $X2=0
+ $Y2=0
cc_403 N_A_792_48#_c_477_n N_A_634_74#_c_608_n 0.0248004f $X=5.185 $Y=1.735
+ $X2=0 $Y2=0
cc_404 N_A_792_48#_c_492_n N_A_634_74#_c_608_n 0.00408476f $X=5.045 $Y=1.9 $X2=0
+ $Y2=0
cc_405 N_A_792_48#_c_486_n N_CLK_c_680_n 0.00325966f $X=5.075 $Y=2.24 $X2=-0.19
+ $Y2=-0.245
cc_406 N_A_792_48#_c_487_n N_CLK_c_680_n 0.0108158f $X=5.045 $Y=2.73 $X2=-0.19
+ $Y2=-0.245
cc_407 N_A_792_48#_c_489_n N_CLK_c_680_n 0.0212761f $X=6.285 $Y=2.325 $X2=-0.19
+ $Y2=-0.245
cc_408 N_A_792_48#_c_490_n N_CLK_c_680_n 0.00223446f $X=6.37 $Y=2.24 $X2=-0.19
+ $Y2=-0.245
cc_409 N_A_792_48#_c_492_n N_CLK_c_680_n 8.90288e-19 $X=5.045 $Y=1.9 $X2=-0.19
+ $Y2=-0.245
cc_410 N_A_792_48#_c_480_n N_CLK_c_676_n 5.87016e-19 $X=5.11 $Y=0.83 $X2=0 $Y2=0
cc_411 N_A_792_48#_c_476_n N_CLK_c_681_n 0.014408f $X=7.015 $Y=1.765 $X2=0 $Y2=0
cc_412 N_A_792_48#_c_489_n N_CLK_c_681_n 0.0135033f $X=6.285 $Y=2.325 $X2=0
+ $Y2=0
cc_413 N_A_792_48#_c_490_n N_CLK_c_681_n 0.0126202f $X=6.37 $Y=2.24 $X2=0 $Y2=0
cc_414 N_A_792_48#_M1008_g N_CLK_c_677_n 0.0363361f $X=6.775 $Y=0.74 $X2=0 $Y2=0
cc_415 N_A_792_48#_M1008_g CLK 2.68908e-19 $X=6.775 $Y=0.74 $X2=0 $Y2=0
cc_416 N_A_792_48#_c_512_n CLK 0.0199562f $X=6.455 $Y=1.465 $X2=0 $Y2=0
cc_417 N_A_792_48#_c_476_n N_CLK_c_679_n 0.0399896f $X=7.015 $Y=1.765 $X2=0
+ $Y2=0
cc_418 N_A_792_48#_c_489_n N_CLK_c_679_n 0.0028431f $X=6.285 $Y=2.325 $X2=0
+ $Y2=0
cc_419 N_A_792_48#_c_490_n N_CLK_c_679_n 0.00704377f $X=6.37 $Y=2.24 $X2=0 $Y2=0
cc_420 N_A_792_48#_c_512_n N_CLK_c_679_n 0.0176052f $X=6.455 $Y=1.465 $X2=0
+ $Y2=0
cc_421 N_A_792_48#_c_478_n N_CLK_c_679_n 0.00352731f $X=6.865 $Y=1.465 $X2=0
+ $Y2=0
cc_422 N_A_792_48#_c_476_n N_A_1289_368#_c_740_n 0.0279145f $X=7.015 $Y=1.765
+ $X2=0 $Y2=0
cc_423 N_A_792_48#_c_476_n N_A_1289_368#_c_744_n 0.0123006f $X=7.015 $Y=1.765
+ $X2=0 $Y2=0
cc_424 N_A_792_48#_M1008_g N_A_1289_368#_c_733_n 0.0119354f $X=6.775 $Y=0.74
+ $X2=0 $Y2=0
cc_425 N_A_792_48#_c_476_n N_A_1289_368#_c_745_n 0.0134697f $X=7.015 $Y=1.765
+ $X2=0 $Y2=0
cc_426 N_A_792_48#_c_478_n N_A_1289_368#_c_745_n 0.00532205f $X=6.865 $Y=1.465
+ $X2=0 $Y2=0
cc_427 N_A_792_48#_c_476_n N_A_1289_368#_c_746_n 0.00729244f $X=7.015 $Y=1.765
+ $X2=0 $Y2=0
cc_428 N_A_792_48#_c_490_n N_A_1289_368#_c_746_n 0.00917426f $X=6.37 $Y=2.24
+ $X2=0 $Y2=0
cc_429 N_A_792_48#_c_478_n N_A_1289_368#_c_746_n 0.0280718f $X=6.865 $Y=1.465
+ $X2=0 $Y2=0
cc_430 N_A_792_48#_M1008_g N_A_1289_368#_c_735_n 0.00395531f $X=6.775 $Y=0.74
+ $X2=0 $Y2=0
cc_431 N_A_792_48#_c_476_n N_A_1289_368#_c_735_n 0.0070975f $X=7.015 $Y=1.765
+ $X2=0 $Y2=0
cc_432 N_A_792_48#_c_478_n N_A_1289_368#_c_735_n 0.0171756f $X=6.865 $Y=1.465
+ $X2=0 $Y2=0
cc_433 N_A_792_48#_M1008_g N_A_1289_368#_c_736_n 0.00401978f $X=6.775 $Y=0.74
+ $X2=0 $Y2=0
cc_434 N_A_792_48#_c_476_n N_A_1289_368#_c_737_n 0.00319597f $X=7.015 $Y=1.765
+ $X2=0 $Y2=0
cc_435 N_A_792_48#_c_476_n N_A_1289_368#_c_738_n 0.00290882f $X=7.015 $Y=1.765
+ $X2=0 $Y2=0
cc_436 N_A_792_48#_c_478_n N_A_1289_368#_c_738_n 0.0175799f $X=6.865 $Y=1.465
+ $X2=0 $Y2=0
cc_437 N_A_792_48#_c_476_n N_A_1289_368#_c_739_n 0.0170664f $X=7.015 $Y=1.765
+ $X2=0 $Y2=0
cc_438 N_A_792_48#_c_478_n N_A_1289_368#_c_739_n 3.3999e-19 $X=6.865 $Y=1.465
+ $X2=0 $Y2=0
cc_439 N_A_792_48#_c_485_n N_VPWR_M1006_d 0.00298389f $X=4.88 $Y=1.82 $X2=0
+ $Y2=0
cc_440 N_A_792_48#_c_489_n N_VPWR_M1023_d 0.0103088f $X=6.285 $Y=2.325 $X2=0
+ $Y2=0
cc_441 N_A_792_48#_c_482_n N_VPWR_c_855_n 0.00333581f $X=4.27 $Y=2.11 $X2=0
+ $Y2=0
cc_442 N_A_792_48#_c_483_n N_VPWR_c_855_n 0.0163507f $X=4.27 $Y=2.2 $X2=0 $Y2=0
cc_443 N_A_792_48#_c_485_n N_VPWR_c_855_n 0.0202359f $X=4.88 $Y=1.82 $X2=0 $Y2=0
cc_444 N_A_792_48#_c_486_n N_VPWR_c_855_n 0.0111704f $X=5.075 $Y=2.24 $X2=0
+ $Y2=0
cc_445 N_A_792_48#_c_487_n N_VPWR_c_855_n 0.0329293f $X=5.045 $Y=2.73 $X2=0
+ $Y2=0
cc_446 N_A_792_48#_c_493_n N_VPWR_c_855_n 0.0121024f $X=5.075 $Y=2.325 $X2=0
+ $Y2=0
cc_447 N_A_792_48#_c_476_n N_VPWR_c_856_n 6.16846e-19 $X=7.015 $Y=1.765 $X2=0
+ $Y2=0
cc_448 N_A_792_48#_c_489_n N_VPWR_c_856_n 0.0220519f $X=6.285 $Y=2.325 $X2=0
+ $Y2=0
cc_449 N_A_792_48#_c_476_n N_VPWR_c_857_n 0.00766779f $X=7.015 $Y=1.765 $X2=0
+ $Y2=0
cc_450 N_A_792_48#_c_476_n N_VPWR_c_861_n 0.00445602f $X=7.015 $Y=1.765 $X2=0
+ $Y2=0
cc_451 N_A_792_48#_c_483_n N_VPWR_c_864_n 0.00410092f $X=4.27 $Y=2.2 $X2=0 $Y2=0
cc_452 N_A_792_48#_c_487_n N_VPWR_c_865_n 0.0128435f $X=5.045 $Y=2.73 $X2=0
+ $Y2=0
cc_453 N_A_792_48#_c_483_n N_VPWR_c_852_n 0.00466677f $X=4.27 $Y=2.2 $X2=0 $Y2=0
cc_454 N_A_792_48#_c_476_n N_VPWR_c_852_n 0.00858994f $X=7.015 $Y=1.765 $X2=0
+ $Y2=0
cc_455 N_A_792_48#_c_487_n N_VPWR_c_852_n 0.0135601f $X=5.045 $Y=2.73 $X2=0
+ $Y2=0
cc_456 N_A_792_48#_M1005_g N_VGND_c_1127_n 0.00667064f $X=4.035 $Y=0.58 $X2=0
+ $Y2=0
cc_457 N_A_792_48#_M1008_g N_VGND_c_1128_n 0.00242918f $X=6.775 $Y=0.74 $X2=0
+ $Y2=0
cc_458 N_A_792_48#_c_512_n N_VGND_c_1128_n 0.00198064f $X=6.455 $Y=1.465 $X2=0
+ $Y2=0
cc_459 N_A_792_48#_M1008_g N_VGND_c_1129_n 0.00353511f $X=6.775 $Y=0.74 $X2=0
+ $Y2=0
cc_460 N_A_792_48#_M1005_g N_VGND_c_1133_n 0.00444681f $X=4.035 $Y=0.58 $X2=0
+ $Y2=0
cc_461 N_A_792_48#_M1008_g N_VGND_c_1137_n 0.00434272f $X=6.775 $Y=0.74 $X2=0
+ $Y2=0
cc_462 N_A_792_48#_M1005_g N_VGND_c_1143_n 0.00877228f $X=4.035 $Y=0.58 $X2=0
+ $Y2=0
cc_463 N_A_792_48#_M1008_g N_VGND_c_1143_n 0.00825979f $X=6.775 $Y=0.74 $X2=0
+ $Y2=0
cc_464 N_A_634_74#_c_601_n N_VPWR_c_855_n 0.00818471f $X=4.82 $Y=1.68 $X2=0
+ $Y2=0
cc_465 N_A_634_74#_c_604_n N_VPWR_c_864_n 0.00640015f $X=3.54 $Y=2.07 $X2=0
+ $Y2=0
cc_466 N_A_634_74#_c_601_n N_VPWR_c_865_n 0.00504123f $X=4.82 $Y=1.68 $X2=0
+ $Y2=0
cc_467 N_A_634_74#_c_601_n N_VPWR_c_852_n 0.00519032f $X=4.82 $Y=1.68 $X2=0
+ $Y2=0
cc_468 N_A_634_74#_c_604_n N_VPWR_c_852_n 0.00771299f $X=3.54 $Y=2.07 $X2=0
+ $Y2=0
cc_469 N_A_634_74#_c_604_n N_A_119_143#_c_967_n 0.0183127f $X=3.54 $Y=2.07 $X2=0
+ $Y2=0
cc_470 N_A_634_74#_c_602_n N_VGND_c_1127_n 0.00126498f $X=4.895 $Y=1.235 $X2=0
+ $Y2=0
cc_471 N_A_634_74#_c_602_n N_VGND_c_1135_n 0.00278271f $X=4.895 $Y=1.235 $X2=0
+ $Y2=0
cc_472 N_A_634_74#_c_602_n N_VGND_c_1143_n 0.00361311f $X=4.895 $Y=1.235 $X2=0
+ $Y2=0
cc_473 N_CLK_c_681_n N_A_1289_368#_c_744_n 0.00997076f $X=6.37 $Y=1.765 $X2=0
+ $Y2=0
cc_474 N_CLK_c_677_n N_A_1289_368#_c_733_n 0.00172581f $X=6.385 $Y=1.22 $X2=0
+ $Y2=0
cc_475 N_CLK_c_681_n N_A_1289_368#_c_746_n 7.6996e-19 $X=6.37 $Y=1.765 $X2=0
+ $Y2=0
cc_476 N_CLK_c_677_n N_A_1289_368#_c_735_n 7.3019e-19 $X=6.385 $Y=1.22 $X2=0
+ $Y2=0
cc_477 N_CLK_c_680_n N_VPWR_c_856_n 0.00641581f $X=5.835 $Y=1.765 $X2=0 $Y2=0
cc_478 N_CLK_c_681_n N_VPWR_c_856_n 0.0111031f $X=6.37 $Y=1.765 $X2=0 $Y2=0
cc_479 N_CLK_c_681_n N_VPWR_c_861_n 0.00413917f $X=6.37 $Y=1.765 $X2=0 $Y2=0
cc_480 N_CLK_c_680_n N_VPWR_c_865_n 0.00402388f $X=5.835 $Y=1.765 $X2=0 $Y2=0
cc_481 N_CLK_c_680_n N_VPWR_c_852_n 0.00462577f $X=5.835 $Y=1.765 $X2=0 $Y2=0
cc_482 N_CLK_c_681_n N_VPWR_c_852_n 0.00819289f $X=6.37 $Y=1.765 $X2=0 $Y2=0
cc_483 N_CLK_c_676_n N_VGND_c_1128_n 0.00470925f $X=5.885 $Y=1.22 $X2=0 $Y2=0
cc_484 N_CLK_c_677_n N_VGND_c_1128_n 0.0156468f $X=6.385 $Y=1.22 $X2=0 $Y2=0
cc_485 CLK N_VGND_c_1128_n 0.00899f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_486 N_CLK_c_679_n N_VGND_c_1128_n 0.00507991f $X=6.37 $Y=1.492 $X2=0 $Y2=0
cc_487 N_CLK_c_676_n N_VGND_c_1135_n 0.00430908f $X=5.885 $Y=1.22 $X2=0 $Y2=0
cc_488 N_CLK_c_677_n N_VGND_c_1137_n 0.00383152f $X=6.385 $Y=1.22 $X2=0 $Y2=0
cc_489 N_CLK_c_676_n N_VGND_c_1143_n 0.00821115f $X=5.885 $Y=1.22 $X2=0 $Y2=0
cc_490 N_CLK_c_677_n N_VGND_c_1143_n 0.0075725f $X=6.385 $Y=1.22 $X2=0 $Y2=0
cc_491 N_A_1289_368#_c_745_n N_VPWR_M1018_d 0.00250594f $X=7.365 $Y=1.885 $X2=0
+ $Y2=0
cc_492 N_A_1289_368#_c_744_n N_VPWR_c_856_n 0.0193844f $X=6.79 $Y=1.985 $X2=0
+ $Y2=0
cc_493 N_A_1289_368#_c_740_n N_VPWR_c_857_n 0.0154175f $X=7.515 $Y=1.765 $X2=0
+ $Y2=0
cc_494 N_A_1289_368#_c_741_n N_VPWR_c_857_n 7.59701e-19 $X=8.095 $Y=1.765 $X2=0
+ $Y2=0
cc_495 N_A_1289_368#_c_744_n N_VPWR_c_857_n 0.0323093f $X=6.79 $Y=1.985 $X2=0
+ $Y2=0
cc_496 N_A_1289_368#_c_745_n N_VPWR_c_857_n 0.0204654f $X=7.365 $Y=1.885 $X2=0
+ $Y2=0
cc_497 N_A_1289_368#_c_741_n N_VPWR_c_858_n 0.00646055f $X=8.095 $Y=1.765 $X2=0
+ $Y2=0
cc_498 N_A_1289_368#_c_742_n N_VPWR_c_858_n 0.00620497f $X=8.595 $Y=1.765 $X2=0
+ $Y2=0
cc_499 N_A_1289_368#_c_742_n N_VPWR_c_860_n 6.43555e-19 $X=8.595 $Y=1.765 $X2=0
+ $Y2=0
cc_500 N_A_1289_368#_c_743_n N_VPWR_c_860_n 0.0174041f $X=9.09 $Y=1.765 $X2=0
+ $Y2=0
cc_501 N_A_1289_368#_c_739_n N_VPWR_c_860_n 8.22785e-19 $X=9.09 $Y=1.532 $X2=0
+ $Y2=0
cc_502 N_A_1289_368#_c_744_n N_VPWR_c_861_n 0.0145938f $X=6.79 $Y=1.985 $X2=0
+ $Y2=0
cc_503 N_A_1289_368#_c_740_n N_VPWR_c_866_n 0.00413917f $X=7.515 $Y=1.765 $X2=0
+ $Y2=0
cc_504 N_A_1289_368#_c_741_n N_VPWR_c_866_n 0.00445602f $X=8.095 $Y=1.765 $X2=0
+ $Y2=0
cc_505 N_A_1289_368#_c_742_n N_VPWR_c_867_n 0.00445602f $X=8.595 $Y=1.765 $X2=0
+ $Y2=0
cc_506 N_A_1289_368#_c_743_n N_VPWR_c_867_n 0.00429299f $X=9.09 $Y=1.765 $X2=0
+ $Y2=0
cc_507 N_A_1289_368#_c_740_n N_VPWR_c_852_n 0.00818839f $X=7.515 $Y=1.765 $X2=0
+ $Y2=0
cc_508 N_A_1289_368#_c_741_n N_VPWR_c_852_n 0.00859163f $X=8.095 $Y=1.765 $X2=0
+ $Y2=0
cc_509 N_A_1289_368#_c_742_n N_VPWR_c_852_n 0.00857795f $X=8.595 $Y=1.765 $X2=0
+ $Y2=0
cc_510 N_A_1289_368#_c_743_n N_VPWR_c_852_n 0.00848138f $X=9.09 $Y=1.765 $X2=0
+ $Y2=0
cc_511 N_A_1289_368#_c_744_n N_VPWR_c_852_n 0.0120466f $X=6.79 $Y=1.985 $X2=0
+ $Y2=0
cc_512 N_A_1289_368#_c_740_n N_GCLK_c_1058_n 0.0124709f $X=7.515 $Y=1.765 $X2=0
+ $Y2=0
cc_513 N_A_1289_368#_c_741_n N_GCLK_c_1058_n 0.0128237f $X=8.095 $Y=1.765 $X2=0
+ $Y2=0
cc_514 N_A_1289_368#_c_742_n N_GCLK_c_1058_n 7.39949e-19 $X=8.595 $Y=1.765 $X2=0
+ $Y2=0
cc_515 N_A_1289_368#_M1001_g N_GCLK_c_1053_n 4.94129e-19 $X=7.765 $Y=0.74 $X2=0
+ $Y2=0
cc_516 N_A_1289_368#_M1013_g N_GCLK_c_1053_n 4.49298e-19 $X=8.245 $Y=0.74 $X2=0
+ $Y2=0
cc_517 N_A_1289_368#_c_741_n N_GCLK_c_1059_n 0.0122806f $X=8.095 $Y=1.765 $X2=0
+ $Y2=0
cc_518 N_A_1289_368#_c_742_n N_GCLK_c_1059_n 0.014256f $X=8.595 $Y=1.765 $X2=0
+ $Y2=0
cc_519 N_A_1289_368#_c_798_p N_GCLK_c_1059_n 0.0295232f $X=8.27 $Y=1.465 $X2=0
+ $Y2=0
cc_520 N_A_1289_368#_c_739_n N_GCLK_c_1059_n 0.00941362f $X=9.09 $Y=1.532 $X2=0
+ $Y2=0
cc_521 N_A_1289_368#_c_740_n N_GCLK_c_1060_n 0.00149391f $X=7.515 $Y=1.765 $X2=0
+ $Y2=0
cc_522 N_A_1289_368#_c_741_n N_GCLK_c_1060_n 9.78171e-19 $X=8.095 $Y=1.765 $X2=0
+ $Y2=0
cc_523 N_A_1289_368#_c_745_n N_GCLK_c_1060_n 0.0149284f $X=7.365 $Y=1.885 $X2=0
+ $Y2=0
cc_524 N_A_1289_368#_c_798_p N_GCLK_c_1060_n 0.0277622f $X=8.27 $Y=1.465 $X2=0
+ $Y2=0
cc_525 N_A_1289_368#_c_739_n N_GCLK_c_1060_n 0.0083172f $X=9.09 $Y=1.532 $X2=0
+ $Y2=0
cc_526 N_A_1289_368#_M1013_g N_GCLK_c_1054_n 0.0124838f $X=8.245 $Y=0.74 $X2=0
+ $Y2=0
cc_527 N_A_1289_368#_M1026_g N_GCLK_c_1054_n 0.013917f $X=8.675 $Y=0.74 $X2=0
+ $Y2=0
cc_528 N_A_1289_368#_c_798_p N_GCLK_c_1054_n 0.0234532f $X=8.27 $Y=1.465 $X2=0
+ $Y2=0
cc_529 N_A_1289_368#_c_739_n N_GCLK_c_1054_n 0.00261961f $X=9.09 $Y=1.532 $X2=0
+ $Y2=0
cc_530 N_A_1289_368#_M1001_g N_GCLK_c_1055_n 2.44239e-19 $X=7.765 $Y=0.74 $X2=0
+ $Y2=0
cc_531 N_A_1289_368#_c_734_n N_GCLK_c_1055_n 0.0053088f $X=7.365 $Y=1.045 $X2=0
+ $Y2=0
cc_532 N_A_1289_368#_c_798_p N_GCLK_c_1055_n 0.0210853f $X=8.27 $Y=1.465 $X2=0
+ $Y2=0
cc_533 N_A_1289_368#_c_739_n N_GCLK_c_1055_n 0.00375571f $X=9.09 $Y=1.532 $X2=0
+ $Y2=0
cc_534 N_A_1289_368#_c_741_n N_GCLK_c_1061_n 6.39139e-19 $X=8.095 $Y=1.765 $X2=0
+ $Y2=0
cc_535 N_A_1289_368#_c_742_n N_GCLK_c_1061_n 0.0121198f $X=8.595 $Y=1.765 $X2=0
+ $Y2=0
cc_536 N_A_1289_368#_c_743_n N_GCLK_c_1061_n 4.36646e-19 $X=9.09 $Y=1.765 $X2=0
+ $Y2=0
cc_537 N_A_1289_368#_M1013_g N_GCLK_c_1056_n 6.74842e-19 $X=8.245 $Y=0.74 $X2=0
+ $Y2=0
cc_538 N_A_1289_368#_M1026_g N_GCLK_c_1056_n 0.00889459f $X=8.675 $Y=0.74 $X2=0
+ $Y2=0
cc_539 N_A_1289_368#_M1027_g N_GCLK_c_1056_n 0.00783249f $X=9.105 $Y=0.74 $X2=0
+ $Y2=0
cc_540 N_A_1289_368#_c_742_n N_GCLK_c_1057_n 9.08574e-19 $X=8.595 $Y=1.765 $X2=0
+ $Y2=0
cc_541 N_A_1289_368#_c_743_n N_GCLK_c_1057_n 9.38216e-19 $X=9.09 $Y=1.765 $X2=0
+ $Y2=0
cc_542 N_A_1289_368#_c_739_n N_GCLK_c_1057_n 0.0321843f $X=9.09 $Y=1.532 $X2=0
+ $Y2=0
cc_543 N_A_1289_368#_c_742_n N_GCLK_c_1063_n 0.0011248f $X=8.595 $Y=1.765 $X2=0
+ $Y2=0
cc_544 N_A_1289_368#_c_743_n N_GCLK_c_1063_n 8.54102e-19 $X=9.09 $Y=1.765 $X2=0
+ $Y2=0
cc_545 N_A_1289_368#_c_739_n N_GCLK_c_1063_n 0.00197711f $X=9.09 $Y=1.532 $X2=0
+ $Y2=0
cc_546 N_A_1289_368#_M1013_g N_GCLK_c_1098_n 9.05544e-19 $X=8.245 $Y=0.74 $X2=0
+ $Y2=0
cc_547 N_A_1289_368#_M1026_g N_GCLK_c_1098_n 0.00624222f $X=8.675 $Y=0.74 $X2=0
+ $Y2=0
cc_548 N_A_1289_368#_M1027_g N_GCLK_c_1098_n 0.0114427f $X=9.105 $Y=0.74 $X2=0
+ $Y2=0
cc_549 N_A_1289_368#_c_798_p N_GCLK_c_1098_n 0.0168342f $X=8.27 $Y=1.465 $X2=0
+ $Y2=0
cc_550 N_A_1289_368#_c_739_n N_GCLK_c_1098_n 0.0158624f $X=9.09 $Y=1.532 $X2=0
+ $Y2=0
cc_551 N_A_1289_368#_c_734_n N_VGND_M1001_d 0.00421825f $X=7.365 $Y=1.045 $X2=0
+ $Y2=0
cc_552 N_A_1289_368#_c_733_n N_VGND_c_1128_n 0.0193094f $X=6.99 $Y=0.515 $X2=0
+ $Y2=0
cc_553 N_A_1289_368#_c_735_n N_VGND_c_1128_n 0.00168579f $X=7.155 $Y=1.045 $X2=0
+ $Y2=0
cc_554 N_A_1289_368#_M1001_g N_VGND_c_1129_n 0.00416717f $X=7.765 $Y=0.74 $X2=0
+ $Y2=0
cc_555 N_A_1289_368#_c_733_n N_VGND_c_1129_n 0.0290535f $X=6.99 $Y=0.515 $X2=0
+ $Y2=0
cc_556 N_A_1289_368#_c_734_n N_VGND_c_1129_n 0.0135013f $X=7.365 $Y=1.045 $X2=0
+ $Y2=0
cc_557 N_A_1289_368#_c_798_p N_VGND_c_1129_n 0.00344427f $X=8.27 $Y=1.465 $X2=0
+ $Y2=0
cc_558 N_A_1289_368#_c_739_n N_VGND_c_1129_n 0.00242237f $X=9.09 $Y=1.532 $X2=0
+ $Y2=0
cc_559 N_A_1289_368#_M1001_g N_VGND_c_1130_n 4.61576e-19 $X=7.765 $Y=0.74 $X2=0
+ $Y2=0
cc_560 N_A_1289_368#_M1013_g N_VGND_c_1130_n 0.00903345f $X=8.245 $Y=0.74 $X2=0
+ $Y2=0
cc_561 N_A_1289_368#_M1026_g N_VGND_c_1130_n 0.00307459f $X=8.675 $Y=0.74 $X2=0
+ $Y2=0
cc_562 N_A_1289_368#_M1027_g N_VGND_c_1132_n 0.00647412f $X=9.105 $Y=0.74 $X2=0
+ $Y2=0
cc_563 N_A_1289_368#_c_733_n N_VGND_c_1137_n 0.0145639f $X=6.99 $Y=0.515 $X2=0
+ $Y2=0
cc_564 N_A_1289_368#_M1001_g N_VGND_c_1138_n 0.00461464f $X=7.765 $Y=0.74 $X2=0
+ $Y2=0
cc_565 N_A_1289_368#_M1013_g N_VGND_c_1138_n 0.00383152f $X=8.245 $Y=0.74 $X2=0
+ $Y2=0
cc_566 N_A_1289_368#_M1026_g N_VGND_c_1139_n 0.00434272f $X=8.675 $Y=0.74 $X2=0
+ $Y2=0
cc_567 N_A_1289_368#_M1027_g N_VGND_c_1139_n 0.00434272f $X=9.105 $Y=0.74 $X2=0
+ $Y2=0
cc_568 N_A_1289_368#_M1001_g N_VGND_c_1143_n 0.0091381f $X=7.765 $Y=0.74 $X2=0
+ $Y2=0
cc_569 N_A_1289_368#_M1013_g N_VGND_c_1143_n 0.00758019f $X=8.245 $Y=0.74 $X2=0
+ $Y2=0
cc_570 N_A_1289_368#_M1026_g N_VGND_c_1143_n 0.00820284f $X=8.675 $Y=0.74 $X2=0
+ $Y2=0
cc_571 N_A_1289_368#_M1027_g N_VGND_c_1143_n 0.00823942f $X=9.105 $Y=0.74 $X2=0
+ $Y2=0
cc_572 N_A_1289_368#_c_733_n N_VGND_c_1143_n 0.0119984f $X=6.99 $Y=0.515 $X2=0
+ $Y2=0
cc_573 N_VPWR_M1002_s N_A_119_143#_c_967_n 0.0189689f $X=1.565 $Y=2.12 $X2=0
+ $Y2=0
cc_574 N_VPWR_c_864_n N_A_119_143#_c_967_n 0.00755275f $X=4.43 $Y=3.33 $X2=0
+ $Y2=0
cc_575 N_VPWR_c_852_n N_A_119_143#_c_967_n 0.0319883f $X=9.36 $Y=3.33 $X2=0
+ $Y2=0
cc_576 N_VPWR_c_854_n N_A_119_143#_c_969_n 0.0103236f $X=0.28 $Y=2.12 $X2=0
+ $Y2=0
cc_577 N_VPWR_c_863_n N_A_119_143#_c_969_n 0.00874223f $X=1.545 $Y=3.33 $X2=0
+ $Y2=0
cc_578 N_VPWR_c_868_n N_A_119_143#_c_969_n 0.0130874f $X=1.99 $Y=2.775 $X2=0
+ $Y2=0
cc_579 N_VPWR_c_852_n N_A_119_143#_c_969_n 0.0107147f $X=9.36 $Y=3.33 $X2=0
+ $Y2=0
cc_580 N_VPWR_M1002_s N_A_119_143#_c_970_n 0.00618702f $X=1.565 $Y=2.12 $X2=0
+ $Y2=0
cc_581 N_VPWR_c_854_n N_A_119_143#_c_970_n 0.0161151f $X=0.28 $Y=2.12 $X2=0
+ $Y2=0
cc_582 N_VPWR_c_868_n N_A_119_143#_c_970_n 0.0448927f $X=1.99 $Y=2.775 $X2=0
+ $Y2=0
cc_583 N_VPWR_c_852_n N_A_119_143#_c_970_n 0.0108335f $X=9.36 $Y=3.33 $X2=0
+ $Y2=0
cc_584 N_VPWR_c_857_n N_GCLK_c_1058_n 0.0485394f $X=7.29 $Y=2.305 $X2=0 $Y2=0
cc_585 N_VPWR_c_858_n N_GCLK_c_1058_n 0.0563525f $X=8.32 $Y=2.305 $X2=0 $Y2=0
cc_586 N_VPWR_c_866_n N_GCLK_c_1058_n 0.0145938f $X=8.235 $Y=3.33 $X2=0 $Y2=0
cc_587 N_VPWR_c_852_n N_GCLK_c_1058_n 0.0120466f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_588 N_VPWR_M1010_s N_GCLK_c_1059_n 0.00275645f $X=8.17 $Y=1.84 $X2=0 $Y2=0
cc_589 N_VPWR_c_858_n N_GCLK_c_1059_n 0.0184684f $X=8.32 $Y=2.305 $X2=0 $Y2=0
cc_590 N_VPWR_c_858_n N_GCLK_c_1061_n 0.0322767f $X=8.32 $Y=2.305 $X2=0 $Y2=0
cc_591 N_VPWR_c_860_n N_GCLK_c_1061_n 0.0386881f $X=9.32 $Y=1.985 $X2=0 $Y2=0
cc_592 N_VPWR_c_867_n N_GCLK_c_1061_n 0.0145938f $X=9.155 $Y=3.33 $X2=0 $Y2=0
cc_593 N_VPWR_c_852_n N_GCLK_c_1061_n 0.0120466f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_594 N_VPWR_c_860_n N_GCLK_c_1063_n 0.00654084f $X=9.32 $Y=1.985 $X2=0 $Y2=0
cc_595 N_VPWR_c_854_n N_VGND_c_1125_n 3.21545e-19 $X=0.28 $Y=2.12 $X2=0 $Y2=0
cc_596 N_A_119_143#_c_961_n N_VGND_M1025_d 0.0155317f $X=1.485 $Y=0.7 $X2=0
+ $Y2=0
cc_597 N_A_119_143#_c_963_n N_VGND_M1025_d 0.00677158f $X=1.57 $Y=1.955 $X2=0
+ $Y2=0
cc_598 N_A_119_143#_c_1012_n N_VGND_M1025_d 8.26265e-19 $X=1.57 $Y=0.7 $X2=0
+ $Y2=0
cc_599 N_A_119_143#_c_960_n N_VGND_c_1125_n 0.0178065f $X=0.78 $Y=0.99 $X2=0
+ $Y2=0
cc_600 N_A_119_143#_c_962_n N_VGND_c_1125_n 0.00875128f $X=0.945 $Y=0.7 $X2=0
+ $Y2=0
cc_601 N_A_119_143#_c_961_n N_VGND_c_1126_n 0.00317977f $X=1.485 $Y=0.7 $X2=0
+ $Y2=0
cc_602 N_A_119_143#_c_962_n N_VGND_c_1126_n 0.00690349f $X=0.945 $Y=0.7 $X2=0
+ $Y2=0
cc_603 N_A_119_143#_c_1012_n N_VGND_c_1133_n 0.0012259f $X=1.57 $Y=0.7 $X2=0
+ $Y2=0
cc_604 N_A_119_143#_c_964_n N_VGND_c_1133_n 0.0144289f $X=2.525 $Y=0.62 $X2=0
+ $Y2=0
cc_605 N_A_119_143#_c_965_n N_VGND_c_1133_n 0.011464f $X=2.305 $Y=0.622 $X2=0
+ $Y2=0
cc_606 N_A_119_143#_c_961_n N_VGND_c_1140_n 0.027214f $X=1.485 $Y=0.7 $X2=0
+ $Y2=0
cc_607 N_A_119_143#_c_1012_n N_VGND_c_1140_n 0.00659988f $X=1.57 $Y=0.7 $X2=0
+ $Y2=0
cc_608 N_A_119_143#_c_961_n N_VGND_c_1143_n 0.00679534f $X=1.485 $Y=0.7 $X2=0
+ $Y2=0
cc_609 N_A_119_143#_c_962_n N_VGND_c_1143_n 0.0101259f $X=0.945 $Y=0.7 $X2=0
+ $Y2=0
cc_610 N_A_119_143#_c_1012_n N_VGND_c_1143_n 0.00319493f $X=1.57 $Y=0.7 $X2=0
+ $Y2=0
cc_611 N_A_119_143#_c_964_n N_VGND_c_1143_n 0.0120887f $X=2.525 $Y=0.62 $X2=0
+ $Y2=0
cc_612 N_A_119_143#_c_965_n N_VGND_c_1143_n 0.0187306f $X=2.305 $Y=0.622 $X2=0
+ $Y2=0
cc_613 N_GCLK_c_1054_n N_VGND_M1013_d 0.00176461f $X=8.725 $Y=1.045 $X2=0 $Y2=0
cc_614 N_GCLK_c_1053_n N_VGND_c_1129_n 0.00122648f $X=8.03 $Y=0.515 $X2=0 $Y2=0
cc_615 N_GCLK_c_1053_n N_VGND_c_1130_n 0.0158413f $X=8.03 $Y=0.515 $X2=0 $Y2=0
cc_616 N_GCLK_c_1054_n N_VGND_c_1130_n 0.0153337f $X=8.725 $Y=1.045 $X2=0 $Y2=0
cc_617 N_GCLK_c_1056_n N_VGND_c_1130_n 0.0164981f $X=8.89 $Y=0.515 $X2=0 $Y2=0
cc_618 N_GCLK_c_1056_n N_VGND_c_1132_n 0.0293763f $X=8.89 $Y=0.515 $X2=0 $Y2=0
cc_619 N_GCLK_c_1053_n N_VGND_c_1138_n 0.011066f $X=8.03 $Y=0.515 $X2=0 $Y2=0
cc_620 N_GCLK_c_1056_n N_VGND_c_1139_n 0.0144922f $X=8.89 $Y=0.515 $X2=0 $Y2=0
cc_621 N_GCLK_c_1053_n N_VGND_c_1143_n 0.00915947f $X=8.03 $Y=0.515 $X2=0 $Y2=0
cc_622 N_GCLK_c_1056_n N_VGND_c_1143_n 0.0118826f $X=8.89 $Y=0.515 $X2=0 $Y2=0
