* File: sky130_fd_sc_ls__o32a_4.spice
* Created: Wed Sep  2 11:22:54 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__o32a_4.pex.spice"
.subckt sky130_fd_sc_ls__o32a_4  VNB VPB B1 B2 A3 A2 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A2	A2
* A3	A3
* B2	B2
* B1	B1
* VPB	VPB
* VNB	VNB
MM1012 N_X_M1012_d N_A_83_256#_M1012_g N_VGND_M1012_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.2543 PD=1.02 PS=2.19 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75000.3
+ SB=75001.8 A=0.111 P=1.78 MULT=1
MM1019 N_X_M1012_d N_A_83_256#_M1019_g N_VGND_M1019_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1554 PD=1.02 PS=1.16 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75000.7
+ SB=75001.3 A=0.111 P=1.78 MULT=1
MM1024 N_X_M1024_d N_A_83_256#_M1024_g N_VGND_M1019_s VNB NSHORT L=0.15 W=0.74
+ AD=0.14985 AS=0.1554 PD=1.145 PS=1.16 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.3
+ SB=75000.8 A=0.111 P=1.78 MULT=1
MM1026 N_X_M1024_d N_A_83_256#_M1026_g N_VGND_M1026_s VNB NSHORT L=0.15 W=0.74
+ AD=0.14985 AS=0.2109 PD=1.145 PS=2.05 NRD=20.268 NRS=0 M=1 R=4.93333
+ SA=75001.8 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1008 N_A_83_256#_M1008_d N_B1_M1008_g N_A_564_74#_M1008_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.1824 PD=0.92 PS=1.85 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75004.7 A=0.096 P=1.58 MULT=1
MM1025 N_A_83_256#_M1008_d N_B1_M1025_g N_A_564_74#_M1025_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.112 PD=0.92 PS=0.99 NRD=0 NRS=13.116 M=1 R=4.26667
+ SA=75000.6 SB=75004.3 A=0.096 P=1.58 MULT=1
MM1020 N_A_564_74#_M1025_s N_B2_M1020_g N_A_83_256#_M1020_s VNB NSHORT L=0.15
+ W=0.64 AD=0.112 AS=0.112 PD=0.99 PS=0.99 NRD=0 NRS=13.116 M=1 R=4.26667
+ SA=75001.1 SB=75003.8 A=0.096 P=1.58 MULT=1
MM1021 N_A_564_74#_M1021_d N_B2_M1021_g N_A_83_256#_M1020_s VNB NSHORT L=0.15
+ W=0.64 AD=0.1216 AS=0.112 PD=1.02 PS=0.99 NRD=13.116 NRS=0 M=1 R=4.26667
+ SA=75001.6 SB=75003.3 A=0.096 P=1.58 MULT=1
MM1001 N_A_564_74#_M1021_d N_A3_M1001_g N_VGND_M1001_s VNB NSHORT L=0.15 W=0.64
+ AD=0.1216 AS=0.1184 PD=1.02 PS=1.01 NRD=5.616 NRS=7.488 M=1 R=4.26667
+ SA=75002.2 SB=75002.7 A=0.096 P=1.58 MULT=1
MM1009 N_A_564_74#_M1009_d N_A3_M1009_g N_VGND_M1001_s VNB NSHORT L=0.15 W=0.64
+ AD=0.096 AS=0.1184 PD=0.94 PS=1.01 NRD=3.744 NRS=9.372 M=1 R=4.26667
+ SA=75002.7 SB=75002.2 A=0.096 P=1.58 MULT=1
MM1003 N_A_564_74#_M1009_d N_A2_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.64
+ AD=0.096 AS=0.112 PD=0.94 PS=0.99 NRD=0 NRS=13.116 M=1 R=4.26667 SA=75003.1
+ SB=75001.8 A=0.096 P=1.58 MULT=1
MM1006 N_A_564_74#_M1006_d N_A2_M1006_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.112 PD=0.92 PS=0.99 NRD=0 NRS=0 M=1 R=4.26667 SA=75003.6
+ SB=75001.3 A=0.096 P=1.58 MULT=1
MM1004 N_VGND_M1004_d N_A1_M1004_g N_A_564_74#_M1006_d VNB NSHORT L=0.15 W=0.64
+ AD=0.152 AS=0.0896 PD=1.115 PS=0.92 NRD=17.808 NRS=0 M=1 R=4.26667 SA=75004.1
+ SB=75000.8 A=0.096 P=1.58 MULT=1
MM1011 N_VGND_M1004_d N_A1_M1011_g N_A_564_74#_M1011_s VNB NSHORT L=0.15 W=0.64
+ AD=0.152 AS=0.1824 PD=1.115 PS=1.85 NRD=18.744 NRS=0 M=1 R=4.26667 SA=75004.7
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1013 N_VPWR_M1013_d N_A_83_256#_M1013_g N_X_M1013_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75003.6 A=0.168 P=2.54 MULT=1
MM1015 N_VPWR_M1015_d N_A_83_256#_M1015_g N_X_M1013_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.196 AS=0.168 PD=1.47 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75003.2 A=0.168 P=2.54 MULT=1
MM1016 N_VPWR_M1015_d N_A_83_256#_M1016_g N_X_M1016_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.196 AS=0.2352 PD=1.47 PS=1.54 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75001.2 SB=75002.7 A=0.168 P=2.54 MULT=1
MM1022 N_VPWR_M1022_d N_A_83_256#_M1022_g N_X_M1016_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.239004 AS=0.2352 PD=1.62717 PS=1.54 NRD=1.7533 NRS=14.0658 M=1 R=7.46667
+ SA=75001.7 SB=75002.1 A=0.168 P=2.54 MULT=1
MM1000 N_VPWR_M1022_d N_B1_M1000_g N_A_534_388#_M1000_s VPB PHIGHVT L=0.15 W=1
+ AD=0.213396 AS=0.22 PD=1.45283 PS=1.44 NRD=25.5903 NRS=15.7403 M=1 R=6.66667
+ SA=75002.3 SB=75001.8 A=0.15 P=2.3 MULT=1
MM1017 N_A_83_256#_M1017_d N_B2_M1017_g N_A_534_388#_M1000_s VPB PHIGHVT L=0.15
+ W=1 AD=0.15 AS=0.22 PD=1.3 PS=1.44 NRD=1.9503 NRS=15.7403 M=1 R=6.66667
+ SA=75002.9 SB=75001.2 A=0.15 P=2.3 MULT=1
MM1023 N_A_83_256#_M1017_d N_B2_M1023_g N_A_534_388#_M1023_s VPB PHIGHVT L=0.15
+ W=1 AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75003.3 SB=75000.7 A=0.15 P=2.3 MULT=1
MM1007 N_VPWR_M1007_d N_B1_M1007_g N_A_534_388#_M1023_s VPB PHIGHVT L=0.15 W=1
+ AD=0.345 AS=0.15 PD=2.69 PS=1.3 NRD=11.8003 NRS=1.9503 M=1 R=6.66667
+ SA=75003.8 SB=75000.3 A=0.15 P=2.3 MULT=1
MM1002 N_A_83_256#_M1002_d N_A3_M1002_g N_A_961_392#_M1002_s VPB PHIGHVT L=0.15
+ W=1 AD=0.16 AS=0.295 PD=1.32 PS=2.59 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75002.7 A=0.15 P=2.3 MULT=1
MM1027 N_A_83_256#_M1002_d N_A3_M1027_g N_A_961_392#_M1027_s VPB PHIGHVT L=0.15
+ W=1 AD=0.16 AS=0.15 PD=1.32 PS=1.3 NRD=5.8903 NRS=1.9503 M=1 R=6.66667
+ SA=75000.7 SB=75002.2 A=0.15 P=2.3 MULT=1
MM1005 N_A_1234_392#_M1005_d N_A2_M1005_g N_A_961_392#_M1027_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.245 AS=0.15 PD=1.49 PS=1.3 NRD=20.685 NRS=1.9503 M=1 R=6.66667
+ SA=75001.1 SB=75001.8 A=0.15 P=2.3 MULT=1
MM1010 N_A_1234_392#_M1005_d N_A1_M1010_g N_VPWR_M1010_s VPB PHIGHVT L=0.15 W=1
+ AD=0.245 AS=0.16 PD=1.49 PS=1.32 NRD=20.685 NRS=3.9203 M=1 R=6.66667
+ SA=75001.8 SB=75001.1 A=0.15 P=2.3 MULT=1
MM1014 N_A_1234_392#_M1014_d N_A1_M1014_g N_VPWR_M1010_s VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.16 PD=1.3 PS=1.32 NRD=1.9503 NRS=3.9203 M=1 R=6.66667 SA=75002.2
+ SB=75000.7 A=0.15 P=2.3 MULT=1
MM1018 N_A_1234_392#_M1014_d N_A2_M1018_g N_A_961_392#_M1018_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.15 AS=0.295 PD=1.3 PS=2.59 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75002.7 SB=75000.2 A=0.15 P=2.3 MULT=1
DX28_noxref VNB VPB NWDIODE A=15.8844 P=20.8
*
.include "sky130_fd_sc_ls__o32a_4.pxi.spice"
*
.ends
*
*
