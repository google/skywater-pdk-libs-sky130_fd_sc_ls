* File: sky130_fd_sc_ls__decaphe_4.pex.spice
* Created: Wed Sep  2 10:59:54 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__DECAPHE_4%VGND 1 9 12 15 24 26
r14 20 22 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r15 19 26 3.14305 $w=1.475e-06 $l=3.8e-07 $layer=LI1_cond $X=0.96 $Y=0 $X2=0.96
+ $Y2=0.38
r16 19 24 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r17 19 22 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r18 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r19 16 26 9.3878 $w=1.475e-06 $l=1.31347e-06 $layer=LI1_cond $X=0.575 $Y=1.515
+ $X2=0.96 $Y2=0.38
r20 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.575
+ $Y=1.515 $X2=0.575 $Y2=1.515
r21 12 24 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=1.68
+ $Y2=0
r22 12 22 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=0.72
+ $Y2=0
r23 10 15 32.6154 $w=3.45e-07 $l=1.95e-07 $layer=POLY_cond $X=0.567 $Y=1.71
+ $X2=0.567 $Y2=1.515
r24 9 10 61.6627 $w=1.13e-06 $l=7.57e-07 $layer=POLY_cond $X=0.96 $Y=2.467
+ $X2=0.96 $Y2=1.71
r25 1 26 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=1.525
+ $Y=0.235 $X2=1.66 $Y2=0.38
r26 1 26 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=1.525
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LS__DECAPHE_4%VPWR 1 8 10 13 16 27 34
r15 28 34 0.0081048 $w=1.92e-06 $l=1.22e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=0.96 $Y2=3.208
r16 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r17 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r18 24 27 3.03205 $w=1.529e-06 $l=3.8e-07 $layer=LI1_cond $X=0.96 $Y=2.95
+ $X2=0.96 $Y2=3.33
r19 21 24 7.6998 $w=1.529e-06 $l=9.65e-07 $layer=LI1_cond $X=0.96 $Y=1.985
+ $X2=0.96 $Y2=2.95
r20 17 21 5.1864 $w=1.529e-06 $l=8.24166e-07 $layer=LI1_cond $X=1.355 $Y=1.335
+ $X2=0.96 $Y2=1.985
r21 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.355
+ $Y=1.335 $X2=1.355 $Y2=1.335
r22 13 34 6.64328e-05 $w=1.92e-06 $l=1e-09 $layer=MET1_cond $X=0.96 $Y=3.207
+ $X2=0.96 $Y2=3.208
r23 11 16 33.589 $w=3.35e-07 $l=1.95e-07 $layer=POLY_cond $X=1.357 $Y=1.14
+ $X2=1.357 $Y2=1.335
r24 10 11 29.5232 $w=3.35e-07 $l=5.18e-07 $layer=POLY_cond $X=1.357 $Y=0.622
+ $X2=1.357 $Y2=1.14
r25 8 10 19.7223 $w=1.035e-06 $l=3.97e-07 $layer=POLY_cond $X=0.96 $Y=0.622
+ $X2=1.357 $Y2=0.622
r26 1 24 400 $w=1.7e-07 $l=1.17556e-06 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.84 $X2=1.66 $Y2=2.95
r27 1 24 400 $w=1.7e-07 $l=1.17083e-06 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.84 $X2=0.26 $Y2=2.95
r28 1 21 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.84 $X2=1.66 $Y2=1.985
r29 1 21 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.84 $X2=0.26 $Y2=1.985
.ends

