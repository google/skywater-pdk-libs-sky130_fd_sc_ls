* File: sky130_fd_sc_ls__decaphe_3.pex.spice
* Created: Wed Sep  2 10:59:47 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__DECAPHE_3%VGND 1 7 9 10 19 21
r9 16 21 4.35714 $w=1.064e-06 $l=3.8e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=0.72
+ $Y2=0.38
r10 16 19 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r11 16 17 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r12 14 21 13.0141 $w=1.064e-06 $l=1.2628e-06 $layer=LI1_cond $X=0.45 $Y=1.515
+ $X2=0.72 $Y2=0.38
r13 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.45
+ $Y=1.515 $X2=0.45 $Y2=1.515
r14 10 19 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r15 10 17 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r16 7 13 41.9172 $w=6.5e-07 $l=6.40937e-07 $layer=POLY_cond $X=0.72 $Y=2.035
+ $X2=0.45 $Y2=1.515
r17 7 9 32.0345 $w=6.5e-07 $l=4.32e-07 $layer=POLY_cond $X=0.72 $Y=2.035
+ $X2=0.72 $Y2=2.467
r18 1 21 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=1.045
+ $Y=0.235 $X2=1.18 $Y2=0.38
r19 1 21 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=1.045
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LS__DECAPHE_3%VPWR 1 7 9 10 13 21 25 33
r12 26 33 0.0108064 $w=1.44e-06 $l=1.22e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.208
r13 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r14 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r15 21 33 8.85771e-05 $w=1.44e-06 $l=1e-09 $layer=MET1_cond $X=0.72 $Y=3.207
+ $X2=0.72 $Y2=3.208
r16 16 19 8.39153 $w=9.45e-07 $l=7.73305e-07 $layer=LI1_cond $X=0.99 $Y=1.335
+ $X2=0.72 $Y2=1.985
r17 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.99
+ $Y=1.335 $X2=0.99 $Y2=1.335
r18 11 25 0.920684 $w=1.438e-06 $l=8.5e-08 $layer=LI1_cond $X=0.72 $Y=3.245
+ $X2=0.72 $Y2=3.33
r19 11 13 2.83386 $w=1.268e-06 $l=2.95e-07 $layer=LI1_cond $X=0.72 $Y=3.245
+ $X2=0.72 $Y2=2.95
r20 10 19 4.85961 $w=1.27e-06 $l=4.2e-07 $layer=LI1_cond $X=0.72 $Y=2.405
+ $X2=0.72 $Y2=1.985
r21 10 13 5.23543 $w=1.268e-06 $l=5.45e-07 $layer=LI1_cond $X=0.72 $Y=2.405
+ $X2=0.72 $Y2=2.95
r22 7 17 41.9172 $w=6.5e-07 $l=6.40937e-07 $layer=POLY_cond $X=0.72 $Y=0.815
+ $X2=0.99 $Y2=1.335
r23 7 9 14.3117 $w=6.5e-07 $l=1.93e-07 $layer=POLY_cond $X=0.72 $Y=0.815
+ $X2=0.72 $Y2=0.622
r24 1 19 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.045
+ $Y=1.84 $X2=1.18 $Y2=1.985
r25 1 19 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.045
+ $Y=1.84 $X2=0.26 $Y2=1.985
r26 1 13 400 $w=1.7e-07 $l=1.17556e-06 $layer=licon1_PDIFF $count=1 $X=1.045
+ $Y=1.84 $X2=1.18 $Y2=2.95
r27 1 13 400 $w=1.7e-07 $l=1.17083e-06 $layer=licon1_PDIFF $count=1 $X=1.045
+ $Y=1.84 $X2=0.26 $Y2=2.95
.ends

