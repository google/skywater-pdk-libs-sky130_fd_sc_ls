* File: sky130_fd_sc_ls__o21ai_2.pex.spice
* Created: Fri Aug 28 13:45:18 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__O21AI_2%A1 3 5 7 10 12 14 17 20 21 23 28
c74 12 0 2.59909e-19 $X=1.955 $Y=1.765
c75 10 0 1.73347e-19 $X=1.925 $Y=0.74
c76 5 0 1.67856e-19 $X=0.505 $Y=1.765
r77 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.92
+ $Y=1.515 $X2=1.92 $Y2=1.515
r78 23 28 3.45023 $w=5.18e-07 $l=1.5e-07 $layer=LI1_cond $X=2.015 $Y=1.665
+ $X2=2.015 $Y2=1.515
r79 22 23 6.55543 $w=5.18e-07 $l=2.85e-07 $layer=LI1_cond $X=2.015 $Y=1.95
+ $X2=2.015 $Y2=1.665
r80 20 22 9.39785 $w=1.7e-07 $l=2.995e-07 $layer=LI1_cond $X=1.755 $Y=2.035
+ $X2=2.015 $Y2=1.95
r81 20 21 75.6791 $w=1.68e-07 $l=1.16e-06 $layer=LI1_cond $X=1.755 $Y=2.035
+ $X2=0.595 $Y2=2.035
r82 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.43
+ $Y=1.515 $X2=0.43 $Y2=1.515
r83 15 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.43 $Y=1.95
+ $X2=0.595 $Y2=2.035
r84 15 17 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=0.43 $Y=1.95
+ $X2=0.43 $Y2=1.515
r85 12 27 52.2586 $w=2.99e-07 $l=2.66927e-07 $layer=POLY_cond $X=1.955 $Y=1.765
+ $X2=1.92 $Y2=1.515
r86 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.955 $Y=1.765
+ $X2=1.955 $Y2=2.4
r87 8 27 38.5562 $w=2.99e-07 $l=1.67481e-07 $layer=POLY_cond $X=1.925 $Y=1.35
+ $X2=1.92 $Y2=1.515
r88 8 10 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.925 $Y=1.35
+ $X2=1.925 $Y2=0.74
r89 5 18 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.43 $Y2=1.515
r90 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.4
r91 1 18 38.5562 $w=2.99e-07 $l=1.94808e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.43 $Y2=1.515
r92 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__O21AI_2%A2 1 3 6 10 12 14 15 21 22
r57 22 23 1.97003 $w=3.67e-07 $l=1.5e-08 $layer=POLY_cond $X=1.44 $Y=1.557
+ $X2=1.455 $Y2=1.557
r58 20 22 11.8202 $w=3.67e-07 $l=9e-08 $layer=POLY_cond $X=1.35 $Y=1.557
+ $X2=1.44 $Y2=1.557
r59 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.35
+ $Y=1.515 $X2=1.35 $Y2=1.515
r60 18 20 46.624 $w=3.67e-07 $l=3.55e-07 $layer=POLY_cond $X=0.995 $Y=1.557
+ $X2=1.35 $Y2=1.557
r61 17 18 5.25341 $w=3.67e-07 $l=4e-08 $layer=POLY_cond $X=0.955 $Y=1.557
+ $X2=0.995 $Y2=1.557
r62 15 21 2.67779 $w=6.68e-07 $l=1.5e-07 $layer=LI1_cond $X=1.18 $Y=1.665
+ $X2=1.18 $Y2=1.515
r63 12 23 23.77 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.455 $Y=1.765
+ $X2=1.455 $Y2=1.557
r64 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.455 $Y=1.765
+ $X2=1.455 $Y2=2.4
r65 8 22 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.44 $Y=1.35 $X2=1.44
+ $Y2=1.557
r66 8 10 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.44 $Y=1.35 $X2=1.44
+ $Y2=0.74
r67 4 18 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.995 $Y=1.35
+ $X2=0.995 $Y2=1.557
r68 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.995 $Y=1.35
+ $X2=0.995 $Y2=0.74
r69 1 17 23.77 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.955 $Y=1.765
+ $X2=0.955 $Y2=1.557
r70 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.955 $Y=1.765
+ $X2=0.955 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__O21AI_2%B1 3 5 7 8 10 12 13 15 17
c46 17 0 1.98552e-19 $X=3.12 $Y=1.295
c47 5 0 1.86656e-19 $X=2.405 $Y=1.765
r48 20 22 14.8201 $w=3.48e-07 $l=1.07e-07 $layer=POLY_cond $X=3 $Y=1.385 $X2=3
+ $Y2=1.492
r49 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.07
+ $Y=1.385 $X2=3.07 $Y2=1.385
r50 17 21 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=3.07 $Y=1.295 $X2=3.07
+ $Y2=1.385
r51 13 20 38.7612 $w=3.48e-07 $l=2.22486e-07 $layer=POLY_cond $X=2.865 $Y=1.22
+ $X2=3 $Y2=1.385
r52 13 15 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.865 $Y=1.22
+ $X2=2.865 $Y2=0.74
r53 10 22 53.7198 $w=3.48e-07 $l=3.37808e-07 $layer=POLY_cond $X=2.855 $Y=1.765
+ $X2=3 $Y2=1.492
r54 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.855 $Y=1.765
+ $X2=2.855 $Y2=2.4
r55 8 22 11.1034 $w=2.45e-07 $l=2.35e-07 $layer=POLY_cond $X=2.765 $Y=1.492
+ $X2=3 $Y2=1.492
r56 8 9 68.4515 $w=2.45e-07 $l=2.7e-07 $layer=POLY_cond $X=2.765 $Y=1.492
+ $X2=2.495 $Y2=1.492
r57 5 9 75.954 $w=1.76e-07 $l=2.73e-07 $layer=POLY_cond $X=2.405 $Y=1.765
+ $X2=2.405 $Y2=1.492
r58 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.405 $Y=1.765
+ $X2=2.405 $Y2=2.4
r59 1 9 34.6006 $w=1.76e-07 $l=1.24475e-07 $layer=POLY_cond $X=2.4 $Y=1.37
+ $X2=2.405 $Y2=1.492
r60 1 3 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=2.4 $Y=1.37 $X2=2.4
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__O21AI_2%VPWR 1 2 3 10 12 16 18 20 24 26 31 40 44
r49 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r50 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r51 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r52 35 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r53 35 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r54 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r55 32 40 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.345 $Y=3.33
+ $X2=2.22 $Y2=3.33
r56 32 34 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.345 $Y=3.33
+ $X2=2.64 $Y2=3.33
r57 31 43 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=2.995 $Y=3.33
+ $X2=3.177 $Y2=3.33
r58 31 34 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=2.995 $Y=3.33
+ $X2=2.64 $Y2=3.33
r59 30 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r60 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r61 27 37 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.182 $Y2=3.33
r62 27 29 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.72 $Y2=3.33
r63 26 40 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.095 $Y=3.33
+ $X2=2.22 $Y2=3.33
r64 26 29 89.7059 $w=1.68e-07 $l=1.375e-06 $layer=LI1_cond $X=2.095 $Y=3.33
+ $X2=0.72 $Y2=3.33
r65 24 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r66 24 30 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r67 20 23 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=3.12 $Y=1.985
+ $X2=3.12 $Y2=2.815
r68 18 43 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=3.12 $Y=3.245
+ $X2=3.177 $Y2=3.33
r69 18 23 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=3.12 $Y=3.245
+ $X2=3.12 $Y2=2.815
r70 14 40 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.22 $Y=3.245
+ $X2=2.22 $Y2=3.33
r71 14 16 20.283 $w=2.48e-07 $l=4.4e-07 $layer=LI1_cond $X=2.22 $Y=3.245
+ $X2=2.22 $Y2=2.805
r72 10 37 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.182 $Y2=3.33
r73 10 12 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.24 $Y2=2.455
r74 3 23 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.93
+ $Y=1.84 $X2=3.08 $Y2=2.815
r75 3 20 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.93
+ $Y=1.84 $X2=3.08 $Y2=1.985
r76 2 16 600 $w=1.7e-07 $l=1.03729e-06 $layer=licon1_PDIFF $count=1 $X=2.03
+ $Y=1.84 $X2=2.18 $Y2=2.805
r77 1 12 300 $w=1.7e-07 $l=6.83667e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_LS__O21AI_2%A_116_368# 1 2 9 11 12 14
c31 14 0 1.86656e-19 $X=1.73 $Y=2.805
c32 11 0 8.35221e-20 $X=1.565 $Y=2.99
r33 14 16 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=1.73 $Y=2.805
+ $X2=1.73 $Y2=2.99
r34 11 16 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.565 $Y=2.99
+ $X2=1.73 $Y2=2.99
r35 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.565 $Y=2.99
+ $X2=0.895 $Y2=2.99
r36 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.73 $Y=2.905
+ $X2=0.895 $Y2=2.99
r37 7 9 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=0.73 $Y=2.905 $X2=0.73
+ $Y2=2.455
r38 2 14 600 $w=1.7e-07 $l=1.06029e-06 $layer=licon1_PDIFF $count=1 $X=1.53
+ $Y=1.84 $X2=1.73 $Y2=2.805
r39 1 9 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=0.58
+ $Y=1.84 $X2=0.73 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_LS__O21AI_2%Y 1 2 3 10 14 18 23 24 25 26 36 44
c42 44 0 1.76387e-19 $X=2.66 $Y=1.82
r43 32 36 1.28049 $w=2.68e-07 $l=3e-08 $layer=LI1_cond $X=2.66 $Y=1.955 $X2=2.66
+ $Y2=1.985
r44 25 33 3.46198 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.66 $Y=2.375
+ $X2=2.66 $Y2=2.29
r45 25 38 3.46198 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.66 $Y=2.375
+ $X2=2.66 $Y2=2.46
r46 25 26 12.8049 $w=2.68e-07 $l=3e-07 $layer=LI1_cond $X=2.66 $Y=2.475 $X2=2.66
+ $Y2=2.775
r47 25 38 0.640246 $w=2.68e-07 $l=1.5e-08 $layer=LI1_cond $X=2.66 $Y=2.475
+ $X2=2.66 $Y2=2.46
r48 24 32 0.128049 $w=2.68e-07 $l=3e-09 $layer=LI1_cond $X=2.66 $Y=1.952
+ $X2=2.66 $Y2=1.955
r49 24 44 6.23403 $w=2.68e-07 $l=1.32e-07 $layer=LI1_cond $X=2.66 $Y=1.952
+ $X2=2.66 $Y2=1.82
r50 24 33 10.7988 $w=2.68e-07 $l=2.53e-07 $layer=LI1_cond $X=2.66 $Y=2.037
+ $X2=2.66 $Y2=2.29
r51 24 36 2.21952 $w=2.68e-07 $l=5.2e-08 $layer=LI1_cond $X=2.66 $Y=2.037
+ $X2=2.66 $Y2=1.985
r52 23 44 36.4416 $w=2.08e-07 $l=6.9e-07 $layer=LI1_cond $X=2.63 $Y=1.13
+ $X2=2.63 $Y2=1.82
r53 18 21 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=1.23 $Y=2.375
+ $X2=1.23 $Y2=2.51
r54 12 23 6.22208 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=2.605 $Y=1 $X2=2.605
+ $Y2=1.13
r55 12 14 5.31897 $w=2.58e-07 $l=1.2e-07 $layer=LI1_cond $X=2.605 $Y=1 $X2=2.605
+ $Y2=0.88
r56 11 18 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.395 $Y=2.375
+ $X2=1.23 $Y2=2.375
r57 10 25 3.05049 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.525 $Y=2.375
+ $X2=2.66 $Y2=2.375
r58 10 11 73.7219 $w=1.68e-07 $l=1.13e-06 $layer=LI1_cond $X=2.525 $Y=2.375
+ $X2=1.395 $Y2=2.375
r59 3 25 300 $w=1.7e-07 $l=6.30555e-07 $layer=licon1_PDIFF $count=2 $X=2.48
+ $Y=1.84 $X2=2.63 $Y2=2.4
r60 3 36 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.48
+ $Y=1.84 $X2=2.63 $Y2=1.985
r61 2 21 600 $w=1.7e-07 $l=7.63479e-07 $layer=licon1_PDIFF $count=1 $X=1.03
+ $Y=1.84 $X2=1.23 $Y2=2.51
r62 1 14 182 $w=1.7e-07 $l=5.88897e-07 $layer=licon1_NDIFF $count=1 $X=2.475
+ $Y=0.37 $X2=2.645 $Y2=0.88
.ends

.subckt PM_SKY130_FD_SC_LS__O21AI_2%A_27_74# 1 2 3 4 15 17 18 21 23 25 27 31 35
c60 27 0 1.98552e-19 $X=2.915 $Y=0.435
c61 25 0 1.73347e-19 $X=2.18 $Y=0.52
c62 17 0 1.67856e-19 $X=1.125 $Y=1.095
r63 28 33 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.305 $Y=0.435
+ $X2=2.18 $Y2=0.435
r64 27 35 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.915 $Y=0.435
+ $X2=3.08 $Y2=0.435
r65 27 28 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=2.915 $Y=0.435
+ $X2=2.305 $Y2=0.435
r66 25 33 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.18 $Y=0.52 $X2=2.18
+ $Y2=0.435
r67 25 26 22.5879 $w=2.48e-07 $l=4.9e-07 $layer=LI1_cond $X=2.18 $Y=0.52
+ $X2=2.18 $Y2=1.01
r68 24 31 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.375 $Y=1.095
+ $X2=1.25 $Y2=1.095
r69 23 26 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.055 $Y=1.095
+ $X2=2.18 $Y2=1.01
r70 23 24 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.055 $Y=1.095
+ $X2=1.375 $Y2=1.095
r71 19 31 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.25 $Y=1.01
+ $X2=1.25 $Y2=1.095
r72 19 21 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=1.25 $Y=1.01
+ $X2=1.25 $Y2=0.515
r73 17 31 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.125 $Y=1.095
+ $X2=1.25 $Y2=1.095
r74 17 18 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.125 $Y=1.095
+ $X2=0.445 $Y2=1.095
r75 13 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=1.01
+ $X2=0.445 $Y2=1.095
r76 13 15 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=0.28 $Y=1.01
+ $X2=0.28 $Y2=0.515
r77 4 35 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.94
+ $Y=0.37 $X2=3.08 $Y2=0.515
r78 3 33 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2 $Y=0.37
+ $X2=2.14 $Y2=0.515
r79 2 21 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.07
+ $Y=0.37 $X2=1.21 $Y2=0.515
r80 1 15 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__O21AI_2%VGND 1 2 9 13 15 17 22 32 33 36 39
r44 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r45 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r46 30 33 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r47 29 32 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r48 29 30 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r49 27 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.875 $Y=0 $X2=1.71
+ $Y2=0
r50 27 29 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.875 $Y=0 $X2=2.16
+ $Y2=0
r51 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r52 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r53 23 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=0.78
+ $Y2=0
r54 23 25 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=1.2
+ $Y2=0
r55 22 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.545 $Y=0 $X2=1.71
+ $Y2=0
r56 22 25 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.545 $Y=0 $X2=1.2
+ $Y2=0
r57 20 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r58 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r59 17 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.78
+ $Y2=0
r60 17 19 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.24
+ $Y2=0
r61 15 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r62 15 26 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r63 15 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r64 11 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.71 $Y=0.085
+ $X2=1.71 $Y2=0
r65 11 13 20.2551 $w=3.28e-07 $l=5.8e-07 $layer=LI1_cond $X=1.71 $Y=0.085
+ $X2=1.71 $Y2=0.665
r66 7 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=0.085 $X2=0.78
+ $Y2=0
r67 7 9 20.2551 $w=3.28e-07 $l=5.8e-07 $layer=LI1_cond $X=0.78 $Y=0.085 $X2=0.78
+ $Y2=0.665
r68 2 13 182 $w=1.7e-07 $l=3.80197e-07 $layer=licon1_NDIFF $count=1 $X=1.515
+ $Y=0.37 $X2=1.71 $Y2=0.665
r69 1 9 182 $w=1.7e-07 $l=3.85973e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.78 $Y2=0.665
.ends

