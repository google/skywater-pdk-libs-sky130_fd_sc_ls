* File: sky130_fd_sc_ls__a2bb2oi_1.spice
* Created: Fri Aug 28 12:56:38 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__a2bb2oi_1.pex.spice"
.subckt sky130_fd_sc_ls__a2bb2oi_1  VNB VPB A1_N A2_N B2 B1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1	B1
* B2	B2
* A2_N	A2_N
* A1_N	A1_N
* VPB	VPB
* VNB	VNB
MM1008 N_A_126_112#_M1008_d N_A1_N_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15
+ W=0.55 AD=0.077 AS=0.14575 PD=0.83 PS=1.63 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75002.5 A=0.0825 P=1.4 MULT=1
MM1007 N_VGND_M1007_d N_A2_N_M1007_g N_A_126_112#_M1008_d VNB NSHORT L=0.15
+ W=0.55 AD=0.209064 AS=0.077 PD=1.31318 PS=0.83 NRD=70.932 NRS=0 M=1 R=3.66667
+ SA=75000.6 SB=75002 A=0.0825 P=1.4 MULT=1
MM1000 N_Y_M1000_d N_A_126_112#_M1000_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.281286 PD=1.02 PS=1.76682 NRD=0 NRS=52.716 M=1 R=4.93333
+ SA=75001.2 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1003 A_488_74# N_B2_M1003_g N_Y_M1000_d VNB NSHORT L=0.15 W=0.74 AD=0.1184
+ AS=0.1036 PD=1.06 PS=1.02 NRD=17.016 NRS=0 M=1 R=4.93333 SA=75001.6 SB=75000.7
+ A=0.111 P=1.78 MULT=1
MM1001 N_VGND_M1001_d N_B1_M1001_g A_488_74# VNB NSHORT L=0.15 W=0.74 AD=0.1961
+ AS=0.1184 PD=2.01 PS=1.06 NRD=0 NRS=17.016 M=1 R=4.93333 SA=75002.1 SB=75000.2
+ A=0.111 P=1.78 MULT=1
MM1004 A_117_392# N_A1_N_M1004_g N_VPWR_M1004_s VPB PHIGHVT L=0.15 W=1 AD=0.12
+ AS=0.275 PD=1.24 PS=2.55 NRD=12.7853 NRS=1.9503 M=1 R=6.66667 SA=75000.2
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1006 N_A_126_112#_M1006_d N_A2_N_M1006_g A_117_392# VPB PHIGHVT L=0.15 W=1
+ AD=0.275 AS=0.12 PD=2.55 PS=1.24 NRD=1.9503 NRS=12.7853 M=1 R=6.66667
+ SA=75000.6 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1005 N_A_399_368#_M1005_d N_A_126_112#_M1005_g N_Y_M1005_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.308 PD=1.42 PS=2.79 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1009 N_VPWR_M1009_d N_B2_M1009_g N_A_399_368#_M1005_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.1848 AS=0.168 PD=1.45 PS=1.42 NRD=4.3931 NRS=1.7533 M=1 R=7.46667
+ SA=75000.6 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1002 N_A_399_368#_M1002_d N_B1_M1002_g N_VPWR_M1009_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.308 AS=0.1848 PD=2.79 PS=1.45 NRD=1.7533 NRS=4.3931 M=1 R=7.46667
+ SA=75001.1 SB=75000.2 A=0.168 P=2.54 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9564 P=11.2
*
.include "sky130_fd_sc_ls__a2bb2oi_1.pxi.spice"
*
.ends
*
*
