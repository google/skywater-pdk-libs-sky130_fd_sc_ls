* NGSPICE file created from sky130_fd_sc_ls__a2bb2oi_1.ext - technology: sky130A

.subckt sky130_fd_sc_ls__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
M1000 Y a_126_112# VGND VNB nshort w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=8.322e+11p ps=6.72e+06u
M1001 VGND B1 a_488_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.368e+11p ps=2.12e+06u
M1002 a_399_368# B1 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=6.44e+11p pd=5.63e+06u as=6.446e+11p ps=5.45e+06u
M1003 a_488_74# B2 Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_117_392# A1_N VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.4e+11p pd=2.48e+06u as=0p ps=0u
M1005 a_399_368# a_126_112# Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.08e+11p ps=2.79e+06u
M1006 a_126_112# A2_N a_117_392# VPB phighvt w=1e+06u l=150000u
+  ad=2.75e+11p pd=2.55e+06u as=0p ps=0u
M1007 VGND A2_N a_126_112# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=1.54e+11p ps=1.66e+06u
M1008 a_126_112# A1_N VGND VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR B2 a_399_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

