* NGSPICE file created from sky130_fd_sc_ls__clkdlyinv5sd1_1.ext - technology: sky130A

.subckt sky130_fd_sc_ls__clkdlyinv5sd1_1 A VGND VNB VPB VPWR Y
M1000 Y a_682_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.136e+11p pd=2.8e+06u as=1.8798e+12p ps=1.011e+07u
M1001 a_549_74# a_288_74# VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=7.623e+11p ps=6.15e+06u
M1002 Y a_682_74# VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1003 VGND a_549_74# a_682_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=2.583e+11p ps=2.07e+06u
M1004 a_549_74# a_288_74# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.65e+11p pd=2.53e+06u as=0p ps=0u
M1005 VPWR a_549_74# a_682_74# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=6.1e+11p ps=3.22e+06u
M1006 VGND A a_28_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1007 VPWR A a_28_74# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1008 a_288_74# a_28_74# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.65e+11p pd=2.53e+06u as=0p ps=0u
M1009 a_288_74# a_28_74# VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
.ends

