* File: sky130_fd_sc_ls__and2_2.spice
* Created: Fri Aug 28 13:02:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__and2_2.pex.spice"
.subckt sky130_fd_sc_ls__and2_2  VNB VPB A B VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1003 A_118_74# N_A_M1003_g N_A_31_74#_M1003_s VNB NSHORT L=0.15 W=0.74
+ AD=0.0888 AS=0.2109 PD=0.98 PS=2.05 NRD=10.536 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1001 N_VGND_M1001_d N_B_M1001_g A_118_74# VNB NSHORT L=0.15 W=0.74 AD=0.1332
+ AS=0.0888 PD=1.1 PS=0.98 NRD=0 NRS=10.536 M=1 R=4.93333 SA=75000.6 SB=75001.2
+ A=0.111 P=1.78 MULT=1
MM1002 N_X_M1002_d N_A_31_74#_M1002_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1332 PD=1.02 PS=1.1 NRD=0 NRS=12.972 M=1 R=4.93333 SA=75001.1
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1007 N_X_M1002_d N_A_31_74#_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.2553 PD=1.02 PS=2.17 NRD=0 NRS=4.86 M=1 R=4.93333 SA=75001.5
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1005 N_A_31_74#_M1005_d N_A_M1005_g N_VPWR_M1005_s VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.29 PD=1.3 PS=2.58 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75000.2
+ SB=75001.6 A=0.15 P=2.3 MULT=1
MM1006 N_VPWR_M1006_d N_B_M1006_g N_A_31_74#_M1005_d VPB PHIGHVT L=0.15 W=1
+ AD=0.182453 AS=0.15 PD=1.39151 PS=1.3 NRD=11.8003 NRS=1.9503 M=1 R=6.66667
+ SA=75000.7 SB=75001.2 A=0.15 P=2.3 MULT=1
MM1000 N_VPWR_M1006_d N_A_31_74#_M1000_g N_X_M1000_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.204347 AS=0.168 PD=1.55849 PS=1.42 NRD=2.6201 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1004 N_VPWR_M1004_d N_A_31_74#_M1004_g N_X_M1000_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3192 AS=0.168 PD=2.81 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.5 SB=75000.2 A=0.168 P=2.54 MULT=1
DX8_noxref VNB VPB NWDIODE A=5.1708 P=9.28
*
.include "sky130_fd_sc_ls__and2_2.pxi.spice"
*
.ends
*
*
