* File: sky130_fd_sc_ls__a2bb2oi_1.pxi.spice
* Created: Fri Aug 28 12:56:38 2020
* 
x_PM_SKY130_FD_SC_LS__A2BB2OI_1%A1_N N_A1_N_c_61_n N_A1_N_c_66_n N_A1_N_M1004_g
+ N_A1_N_M1008_g A1_N N_A1_N_c_63_n N_A1_N_c_64_n
+ PM_SKY130_FD_SC_LS__A2BB2OI_1%A1_N
x_PM_SKY130_FD_SC_LS__A2BB2OI_1%A2_N N_A2_N_c_89_n N_A2_N_M1006_g N_A2_N_M1007_g
+ A2_N N_A2_N_c_91_n PM_SKY130_FD_SC_LS__A2BB2OI_1%A2_N
x_PM_SKY130_FD_SC_LS__A2BB2OI_1%A_126_112# N_A_126_112#_M1008_d
+ N_A_126_112#_M1006_d N_A_126_112#_c_135_n N_A_126_112#_M1005_g
+ N_A_126_112#_M1000_g N_A_126_112#_c_128_n N_A_126_112#_c_129_n
+ N_A_126_112#_c_130_n N_A_126_112#_c_131_n N_A_126_112#_c_132_n
+ N_A_126_112#_c_137_n N_A_126_112#_c_133_n N_A_126_112#_c_138_n
+ N_A_126_112#_c_134_n PM_SKY130_FD_SC_LS__A2BB2OI_1%A_126_112#
x_PM_SKY130_FD_SC_LS__A2BB2OI_1%B2 N_B2_c_198_n N_B2_M1003_g N_B2_c_199_n
+ N_B2_M1009_g N_B2_c_200_n B2 B2 PM_SKY130_FD_SC_LS__A2BB2OI_1%B2
x_PM_SKY130_FD_SC_LS__A2BB2OI_1%B1 N_B1_c_239_n N_B1_M1001_g N_B1_c_240_n
+ N_B1_M1002_g B1 PM_SKY130_FD_SC_LS__A2BB2OI_1%B1
x_PM_SKY130_FD_SC_LS__A2BB2OI_1%VPWR N_VPWR_M1004_s N_VPWR_M1009_d
+ N_VPWR_c_266_n N_VPWR_c_267_n N_VPWR_c_268_n N_VPWR_c_269_n N_VPWR_c_270_n
+ N_VPWR_c_271_n VPWR N_VPWR_c_272_n N_VPWR_c_265_n
+ PM_SKY130_FD_SC_LS__A2BB2OI_1%VPWR
x_PM_SKY130_FD_SC_LS__A2BB2OI_1%Y N_Y_M1000_d N_Y_M1005_s N_Y_c_308_n
+ N_Y_c_319_n N_Y_c_309_n Y N_Y_c_312_n PM_SKY130_FD_SC_LS__A2BB2OI_1%Y
x_PM_SKY130_FD_SC_LS__A2BB2OI_1%A_399_368# N_A_399_368#_M1005_d
+ N_A_399_368#_M1002_d N_A_399_368#_c_354_n N_A_399_368#_c_361_n
+ N_A_399_368#_c_359_n N_A_399_368#_c_355_n N_A_399_368#_c_356_n
+ N_A_399_368#_c_357_n PM_SKY130_FD_SC_LS__A2BB2OI_1%A_399_368#
x_PM_SKY130_FD_SC_LS__A2BB2OI_1%VGND N_VGND_M1008_s N_VGND_M1007_d
+ N_VGND_M1001_d N_VGND_c_382_n N_VGND_c_383_n N_VGND_c_384_n N_VGND_c_385_n
+ VGND N_VGND_c_386_n N_VGND_c_387_n N_VGND_c_388_n N_VGND_c_389_n
+ PM_SKY130_FD_SC_LS__A2BB2OI_1%VGND
cc_1 VNB N_A1_N_c_61_n 0.00441374f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.795
cc_2 VNB N_A1_N_M1008_g 0.0237325f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=0.835
cc_3 VNB N_A1_N_c_63_n 0.00807592f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.425
cc_4 VNB N_A1_N_c_64_n 0.0632721f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.425
cc_5 VNB N_A2_N_c_89_n 0.0208003f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.59
cc_6 VNB N_A2_N_M1007_g 0.0306328f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.26
cc_7 VNB N_A2_N_c_91_n 0.0040235f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.425
cc_8 VNB N_A_126_112#_c_128_n 0.0630307f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.425
cc_9 VNB N_A_126_112#_c_129_n 0.0192514f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.425
cc_10 VNB N_A_126_112#_c_130_n 0.00324684f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_126_112#_c_131_n 0.00448426f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_126_112#_c_132_n 0.00299965f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_126_112#_c_133_n 0.016101f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_126_112#_c_134_n 0.00167709f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_B2_c_198_n 0.0181973f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.59
cc_16 VNB N_B2_c_199_n 0.0378478f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.46
cc_17 VNB N_B2_c_200_n 0.012229f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB B2 0.00266487f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.425
cc_19 VNB N_B1_c_239_n 0.0214642f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.59
cc_20 VNB N_B1_c_240_n 0.0686619f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.46
cc_21 VNB B1 0.0113021f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=0.835
cc_22 VNB N_VPWR_c_265_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_Y_c_308_n 0.00408087f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_24 VNB N_Y_c_309_n 0.00214178f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.425
cc_25 VNB N_VGND_c_382_n 0.0125919f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_26 VNB N_VGND_c_383_n 0.0476835f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.425
cc_27 VNB N_VGND_c_384_n 0.0129842f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.425
cc_28 VNB N_VGND_c_385_n 0.0350088f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.425
cc_29 VNB N_VGND_c_386_n 0.0198125f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_387_n 0.029426f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_388_n 0.037158f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_389_n 0.220717f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VPB N_A1_N_c_61_n 0.00884556f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.795
cc_34 VPB N_A1_N_c_66_n 0.0274782f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.885
cc_35 VPB N_A1_N_c_63_n 0.00790246f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.425
cc_36 VPB N_A2_N_c_89_n 0.0418373f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.59
cc_37 VPB N_A2_N_c_91_n 0.0084025f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.425
cc_38 VPB N_A_126_112#_c_135_n 0.0190761f $X=-0.19 $Y=1.66 $X2=0.555 $Y2=0.835
cc_39 VPB N_A_126_112#_c_128_n 0.00725952f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.425
cc_40 VPB N_A_126_112#_c_137_n 0.0113317f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_41 VPB N_A_126_112#_c_138_n 0.0140249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_42 VPB N_A_126_112#_c_134_n 0.00592203f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_43 VPB N_B2_c_199_n 0.0228134f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=2.46
cc_44 VPB B2 0.00410131f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.425
cc_45 VPB N_B1_c_240_n 0.0310665f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=2.46
cc_46 VPB N_VPWR_c_266_n 0.0121701f $X=-0.19 $Y=1.66 $X2=0.555 $Y2=0.835
cc_47 VPB N_VPWR_c_267_n 0.0513344f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_268_n 0.0054586f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.425
cc_49 VPB N_VPWR_c_269_n 0.00150457f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_270_n 0.0561909f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_271_n 0.00307912f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_272_n 0.02286f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_265_n 0.0791058f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_Y_c_308_n 7.95989e-19 $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_55 VPB Y 0.0064256f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.665
cc_56 VPB N_Y_c_312_n 0.00789637f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_A_399_368#_c_354_n 0.00215844f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_A_399_368#_c_355_n 0.0234697f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.425
cc_59 VPB N_A_399_368#_c_356_n 0.0180958f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.665
cc_60 VPB N_A_399_368#_c_357_n 0.00717518f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 N_A1_N_c_66_n N_A2_N_c_89_n 0.0596299f $X=0.51 $Y=1.885 $X2=-0.19
+ $Y2=-0.245
cc_62 N_A1_N_c_63_n N_A2_N_c_89_n 2.2065e-19 $X=0.27 $Y=1.425 $X2=-0.19
+ $Y2=-0.245
cc_63 N_A1_N_c_64_n N_A2_N_c_89_n 0.0264272f $X=0.51 $Y=1.425 $X2=-0.19
+ $Y2=-0.245
cc_64 N_A1_N_M1008_g N_A2_N_M1007_g 0.026924f $X=0.555 $Y=0.835 $X2=0 $Y2=0
cc_65 N_A1_N_c_63_n N_A2_N_M1007_g 8.21582e-19 $X=0.27 $Y=1.425 $X2=0 $Y2=0
cc_66 N_A1_N_c_64_n N_A2_N_M1007_g 0.00166236f $X=0.51 $Y=1.425 $X2=0 $Y2=0
cc_67 N_A1_N_c_63_n N_A2_N_c_91_n 0.026906f $X=0.27 $Y=1.425 $X2=0 $Y2=0
cc_68 N_A1_N_c_64_n N_A2_N_c_91_n 0.00355419f $X=0.51 $Y=1.425 $X2=0 $Y2=0
cc_69 N_A1_N_M1008_g N_A_126_112#_c_130_n 0.00609347f $X=0.555 $Y=0.835 $X2=0
+ $Y2=0
cc_70 N_A1_N_M1008_g N_A_126_112#_c_132_n 0.00485745f $X=0.555 $Y=0.835 $X2=0
+ $Y2=0
cc_71 N_A1_N_c_66_n N_A_126_112#_c_138_n 0.00288159f $X=0.51 $Y=1.885 $X2=0
+ $Y2=0
cc_72 N_A1_N_c_66_n N_VPWR_c_267_n 0.022912f $X=0.51 $Y=1.885 $X2=0 $Y2=0
cc_73 N_A1_N_c_63_n N_VPWR_c_267_n 0.028685f $X=0.27 $Y=1.425 $X2=0 $Y2=0
cc_74 N_A1_N_c_64_n N_VPWR_c_267_n 0.00152171f $X=0.51 $Y=1.425 $X2=0 $Y2=0
cc_75 N_A1_N_c_66_n N_VPWR_c_270_n 0.00413917f $X=0.51 $Y=1.885 $X2=0 $Y2=0
cc_76 N_A1_N_c_66_n N_VPWR_c_265_n 0.00817239f $X=0.51 $Y=1.885 $X2=0 $Y2=0
cc_77 N_A1_N_M1008_g N_VGND_c_383_n 0.00759578f $X=0.555 $Y=0.835 $X2=0 $Y2=0
cc_78 N_A1_N_c_63_n N_VGND_c_383_n 0.0212796f $X=0.27 $Y=1.425 $X2=0 $Y2=0
cc_79 N_A1_N_c_64_n N_VGND_c_383_n 0.00195951f $X=0.51 $Y=1.425 $X2=0 $Y2=0
cc_80 N_A1_N_M1008_g N_VGND_c_386_n 0.0043356f $X=0.555 $Y=0.835 $X2=0 $Y2=0
cc_81 N_A1_N_M1008_g N_VGND_c_389_n 0.00487769f $X=0.555 $Y=0.835 $X2=0 $Y2=0
cc_82 N_A2_N_c_89_n N_A_126_112#_c_135_n 6.59859e-19 $X=0.9 $Y=1.885 $X2=0 $Y2=0
cc_83 N_A2_N_c_89_n N_A_126_112#_c_128_n 0.00856986f $X=0.9 $Y=1.885 $X2=0 $Y2=0
cc_84 N_A2_N_M1007_g N_A_126_112#_c_128_n 0.00790174f $X=0.985 $Y=0.835 $X2=0
+ $Y2=0
cc_85 N_A2_N_M1007_g N_A_126_112#_c_130_n 0.0115029f $X=0.985 $Y=0.835 $X2=0
+ $Y2=0
cc_86 N_A2_N_c_89_n N_A_126_112#_c_131_n 0.00310949f $X=0.9 $Y=1.885 $X2=0 $Y2=0
cc_87 N_A2_N_M1007_g N_A_126_112#_c_131_n 0.0131318f $X=0.985 $Y=0.835 $X2=0
+ $Y2=0
cc_88 N_A2_N_c_91_n N_A_126_112#_c_131_n 0.00723539f $X=1.005 $Y=1.615 $X2=0
+ $Y2=0
cc_89 N_A2_N_c_89_n N_A_126_112#_c_132_n 0.00190041f $X=0.9 $Y=1.885 $X2=0 $Y2=0
cc_90 N_A2_N_M1007_g N_A_126_112#_c_132_n 0.00204917f $X=0.985 $Y=0.835 $X2=0
+ $Y2=0
cc_91 N_A2_N_c_91_n N_A_126_112#_c_132_n 0.0179531f $X=1.005 $Y=1.615 $X2=0
+ $Y2=0
cc_92 N_A2_N_c_89_n N_A_126_112#_c_137_n 0.0144716f $X=0.9 $Y=1.885 $X2=0 $Y2=0
cc_93 N_A2_N_c_89_n N_A_126_112#_c_133_n 6.89529e-19 $X=0.9 $Y=1.885 $X2=0 $Y2=0
cc_94 N_A2_N_M1007_g N_A_126_112#_c_133_n 0.00852072f $X=0.985 $Y=0.835 $X2=0
+ $Y2=0
cc_95 N_A2_N_c_91_n N_A_126_112#_c_133_n 0.00833414f $X=1.005 $Y=1.615 $X2=0
+ $Y2=0
cc_96 N_A2_N_c_89_n N_A_126_112#_c_138_n 0.0100021f $X=0.9 $Y=1.885 $X2=0 $Y2=0
cc_97 N_A2_N_c_91_n N_A_126_112#_c_138_n 0.0116584f $X=1.005 $Y=1.615 $X2=0
+ $Y2=0
cc_98 N_A2_N_c_89_n N_A_126_112#_c_134_n 0.00782706f $X=0.9 $Y=1.885 $X2=0 $Y2=0
cc_99 N_A2_N_c_91_n N_A_126_112#_c_134_n 0.0178064f $X=1.005 $Y=1.615 $X2=0
+ $Y2=0
cc_100 N_A2_N_c_89_n N_VPWR_c_267_n 0.00343399f $X=0.9 $Y=1.885 $X2=0 $Y2=0
cc_101 N_A2_N_c_89_n N_VPWR_c_270_n 0.00445602f $X=0.9 $Y=1.885 $X2=0 $Y2=0
cc_102 N_A2_N_c_89_n N_VPWR_c_265_n 0.00862666f $X=0.9 $Y=1.885 $X2=0 $Y2=0
cc_103 N_A2_N_c_89_n Y 5.93535e-19 $X=0.9 $Y=1.885 $X2=0 $Y2=0
cc_104 N_A2_N_c_89_n N_Y_c_312_n 9.66313e-19 $X=0.9 $Y=1.885 $X2=0 $Y2=0
cc_105 N_A2_N_M1007_g N_VGND_c_386_n 0.0043356f $X=0.985 $Y=0.835 $X2=0 $Y2=0
cc_106 N_A2_N_M1007_g N_VGND_c_388_n 0.0101051f $X=0.985 $Y=0.835 $X2=0 $Y2=0
cc_107 N_A2_N_M1007_g N_VGND_c_389_n 0.00487769f $X=0.985 $Y=0.835 $X2=0 $Y2=0
cc_108 N_A_126_112#_c_129_n N_B2_c_198_n 0.0115596f $X=1.92 $Y=1.22 $X2=-0.19
+ $Y2=-0.245
cc_109 N_A_126_112#_c_135_n N_B2_c_199_n 0.0365259f $X=1.92 $Y=1.765 $X2=0 $Y2=0
cc_110 N_A_126_112#_c_128_n N_B2_c_199_n 0.0308497f $X=1.83 $Y=1.385 $X2=0 $Y2=0
cc_111 N_A_126_112#_c_128_n N_B2_c_200_n 3.62081e-19 $X=1.83 $Y=1.385 $X2=0
+ $Y2=0
cc_112 N_A_126_112#_c_138_n N_VPWR_c_267_n 0.0316462f $X=1.125 $Y=2.115 $X2=0
+ $Y2=0
cc_113 N_A_126_112#_c_135_n N_VPWR_c_268_n 5.38127e-19 $X=1.92 $Y=1.765 $X2=0
+ $Y2=0
cc_114 N_A_126_112#_c_135_n N_VPWR_c_270_n 0.00445602f $X=1.92 $Y=1.765 $X2=0
+ $Y2=0
cc_115 N_A_126_112#_c_137_n N_VPWR_c_270_n 0.0145938f $X=1.125 $Y=2.815 $X2=0
+ $Y2=0
cc_116 N_A_126_112#_c_135_n N_VPWR_c_265_n 0.00863237f $X=1.92 $Y=1.765 $X2=0
+ $Y2=0
cc_117 N_A_126_112#_c_137_n N_VPWR_c_265_n 0.0120466f $X=1.125 $Y=2.815 $X2=0
+ $Y2=0
cc_118 N_A_126_112#_c_128_n N_Y_c_308_n 0.0151646f $X=1.83 $Y=1.385 $X2=0 $Y2=0
cc_119 N_A_126_112#_c_129_n N_Y_c_308_n 0.00510828f $X=1.92 $Y=1.22 $X2=0 $Y2=0
cc_120 N_A_126_112#_c_133_n N_Y_c_308_n 0.030479f $X=1.355 $Y=1.55 $X2=0 $Y2=0
cc_121 N_A_126_112#_c_134_n N_Y_c_308_n 0.00700267f $X=1.2 $Y=1.95 $X2=0 $Y2=0
cc_122 N_A_126_112#_c_129_n N_Y_c_319_n 0.0121303f $X=1.92 $Y=1.22 $X2=0 $Y2=0
cc_123 N_A_126_112#_c_133_n N_Y_c_319_n 0.00359949f $X=1.355 $Y=1.55 $X2=0 $Y2=0
cc_124 N_A_126_112#_c_135_n Y 0.0190833f $X=1.92 $Y=1.765 $X2=0 $Y2=0
cc_125 N_A_126_112#_c_128_n Y 0.00942114f $X=1.83 $Y=1.385 $X2=0 $Y2=0
cc_126 N_A_126_112#_c_137_n Y 0.0170006f $X=1.125 $Y=2.815 $X2=0 $Y2=0
cc_127 N_A_126_112#_c_133_n Y 0.00749614f $X=1.355 $Y=1.55 $X2=0 $Y2=0
cc_128 N_A_126_112#_c_134_n Y 0.03129f $X=1.2 $Y=1.95 $X2=0 $Y2=0
cc_129 N_A_126_112#_c_135_n N_Y_c_312_n 0.00279467f $X=1.92 $Y=1.765 $X2=0 $Y2=0
cc_130 N_A_126_112#_c_137_n N_Y_c_312_n 0.0361954f $X=1.125 $Y=2.815 $X2=0 $Y2=0
cc_131 N_A_126_112#_c_135_n N_A_399_368#_c_354_n 0.00560986f $X=1.92 $Y=1.765
+ $X2=0 $Y2=0
cc_132 N_A_126_112#_c_135_n N_A_399_368#_c_359_n 0.00327885f $X=1.92 $Y=1.765
+ $X2=0 $Y2=0
cc_133 N_A_126_112#_c_131_n N_VGND_M1007_d 0.0017426f $X=1.27 $Y=1.045 $X2=0
+ $Y2=0
cc_134 N_A_126_112#_c_133_n N_VGND_M1007_d 0.00480103f $X=1.355 $Y=1.55 $X2=0
+ $Y2=0
cc_135 N_A_126_112#_c_130_n N_VGND_c_383_n 0.0157455f $X=0.77 $Y=0.835 $X2=0
+ $Y2=0
cc_136 N_A_126_112#_c_130_n N_VGND_c_386_n 0.00800702f $X=0.77 $Y=0.835 $X2=0
+ $Y2=0
cc_137 N_A_126_112#_c_129_n N_VGND_c_387_n 0.00383152f $X=1.92 $Y=1.22 $X2=0
+ $Y2=0
cc_138 N_A_126_112#_c_128_n N_VGND_c_388_n 0.00589713f $X=1.83 $Y=1.385 $X2=0
+ $Y2=0
cc_139 N_A_126_112#_c_129_n N_VGND_c_388_n 0.0120043f $X=1.92 $Y=1.22 $X2=0
+ $Y2=0
cc_140 N_A_126_112#_c_130_n N_VGND_c_388_n 0.0103109f $X=0.77 $Y=0.835 $X2=0
+ $Y2=0
cc_141 N_A_126_112#_c_131_n N_VGND_c_388_n 0.0124114f $X=1.27 $Y=1.045 $X2=0
+ $Y2=0
cc_142 N_A_126_112#_c_133_n N_VGND_c_388_n 0.0262437f $X=1.355 $Y=1.55 $X2=0
+ $Y2=0
cc_143 N_A_126_112#_c_129_n N_VGND_c_389_n 0.00753023f $X=1.92 $Y=1.22 $X2=0
+ $Y2=0
cc_144 N_A_126_112#_c_130_n N_VGND_c_389_n 0.0105477f $X=0.77 $Y=0.835 $X2=0
+ $Y2=0
cc_145 N_B2_c_198_n N_B1_c_239_n 0.036204f $X=2.365 $Y=1.22 $X2=-0.19 $Y2=-0.245
cc_146 N_B2_c_199_n N_B1_c_240_n 0.0602332f $X=2.37 $Y=1.765 $X2=0 $Y2=0
cc_147 N_B2_c_200_n N_B1_c_240_n 0.00279141f $X=2.64 $Y=1.38 $X2=0 $Y2=0
cc_148 B2 N_B1_c_240_n 0.00927274f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_149 N_B2_c_199_n B1 2.21801e-19 $X=2.37 $Y=1.765 $X2=0 $Y2=0
cc_150 N_B2_c_200_n B1 0.0262884f $X=2.64 $Y=1.38 $X2=0 $Y2=0
cc_151 B2 B1 7.69126e-19 $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_152 B2 N_VPWR_M1009_d 0.00898662f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_153 N_B2_c_199_n N_VPWR_c_268_n 0.00313506f $X=2.37 $Y=1.765 $X2=0 $Y2=0
cc_154 N_B2_c_199_n N_VPWR_c_269_n 0.00300755f $X=2.37 $Y=1.765 $X2=0 $Y2=0
cc_155 N_B2_c_199_n N_VPWR_c_270_n 0.00413917f $X=2.37 $Y=1.765 $X2=0 $Y2=0
cc_156 N_B2_c_199_n N_VPWR_c_265_n 0.00398725f $X=2.37 $Y=1.765 $X2=0 $Y2=0
cc_157 N_B2_c_198_n N_Y_c_308_n 0.00215891f $X=2.365 $Y=1.22 $X2=0 $Y2=0
cc_158 N_B2_c_199_n N_Y_c_308_n 0.00260055f $X=2.37 $Y=1.765 $X2=0 $Y2=0
cc_159 N_B2_c_200_n N_Y_c_308_n 0.0249332f $X=2.64 $Y=1.38 $X2=0 $Y2=0
cc_160 B2 N_Y_c_308_n 0.00784186f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_161 N_B2_c_198_n N_Y_c_319_n 0.00359011f $X=2.365 $Y=1.22 $X2=0 $Y2=0
cc_162 N_B2_c_199_n N_Y_c_319_n 0.00146891f $X=2.37 $Y=1.765 $X2=0 $Y2=0
cc_163 N_B2_c_200_n N_Y_c_319_n 0.00483333f $X=2.64 $Y=1.38 $X2=0 $Y2=0
cc_164 N_B2_c_198_n N_Y_c_309_n 0.0101871f $X=2.365 $Y=1.22 $X2=0 $Y2=0
cc_165 N_B2_c_199_n Y 0.00201004f $X=2.37 $Y=1.765 $X2=0 $Y2=0
cc_166 N_B2_c_200_n Y 0.001473f $X=2.64 $Y=1.38 $X2=0 $Y2=0
cc_167 B2 Y 0.00504761f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_168 N_B2_c_199_n N_A_399_368#_c_354_n 0.00492254f $X=2.37 $Y=1.765 $X2=0
+ $Y2=0
cc_169 N_B2_c_199_n N_A_399_368#_c_361_n 0.0155314f $X=2.37 $Y=1.765 $X2=0 $Y2=0
cc_170 B2 N_A_399_368#_c_361_n 0.0119897f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_171 B2 N_A_399_368#_c_355_n 0.0106226f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_172 N_B2_c_198_n N_VGND_c_385_n 0.00253877f $X=2.365 $Y=1.22 $X2=0 $Y2=0
cc_173 N_B2_c_198_n N_VGND_c_387_n 0.00434272f $X=2.365 $Y=1.22 $X2=0 $Y2=0
cc_174 N_B2_c_198_n N_VGND_c_388_n 6.57074e-19 $X=2.365 $Y=1.22 $X2=0 $Y2=0
cc_175 N_B2_c_198_n N_VGND_c_389_n 0.00821825f $X=2.365 $Y=1.22 $X2=0 $Y2=0
cc_176 N_B1_c_240_n N_VPWR_c_268_n 0.00229532f $X=2.85 $Y=1.765 $X2=0 $Y2=0
cc_177 N_B1_c_240_n N_VPWR_c_269_n 0.00325983f $X=2.85 $Y=1.765 $X2=0 $Y2=0
cc_178 N_B1_c_240_n N_VPWR_c_272_n 0.00444483f $X=2.85 $Y=1.765 $X2=0 $Y2=0
cc_179 N_B1_c_240_n N_VPWR_c_265_n 0.00442547f $X=2.85 $Y=1.765 $X2=0 $Y2=0
cc_180 N_B1_c_239_n N_Y_c_319_n 5.76856e-19 $X=2.835 $Y=1.22 $X2=0 $Y2=0
cc_181 N_B1_c_239_n N_Y_c_309_n 0.00160641f $X=2.835 $Y=1.22 $X2=0 $Y2=0
cc_182 N_B1_c_240_n N_A_399_368#_c_361_n 0.0142684f $X=2.85 $Y=1.765 $X2=0 $Y2=0
cc_183 N_B1_c_240_n N_A_399_368#_c_355_n 0.00910144f $X=2.85 $Y=1.765 $X2=0
+ $Y2=0
cc_184 B1 N_A_399_368#_c_355_n 0.0149782f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_185 N_B1_c_240_n N_A_399_368#_c_356_n 0.00533707f $X=2.85 $Y=1.765 $X2=0
+ $Y2=0
cc_186 N_B1_c_239_n N_VGND_c_385_n 0.0184513f $X=2.835 $Y=1.22 $X2=0 $Y2=0
cc_187 N_B1_c_240_n N_VGND_c_385_n 0.00192942f $X=2.85 $Y=1.765 $X2=0 $Y2=0
cc_188 B1 N_VGND_c_385_n 0.0235157f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_189 N_B1_c_239_n N_VGND_c_387_n 0.00383152f $X=2.835 $Y=1.22 $X2=0 $Y2=0
cc_190 N_B1_c_239_n N_VGND_c_389_n 0.00757998f $X=2.835 $Y=1.22 $X2=0 $Y2=0
cc_191 N_VPWR_c_270_n N_Y_c_312_n 0.0110698f $X=2.43 $Y=3.33 $X2=0 $Y2=0
cc_192 N_VPWR_c_265_n N_Y_c_312_n 0.00916093f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_193 N_VPWR_c_269_n N_A_399_368#_c_354_n 0.0168379f $X=2.61 $Y=2.815 $X2=0
+ $Y2=0
cc_194 N_VPWR_c_270_n N_A_399_368#_c_354_n 0.0109113f $X=2.43 $Y=3.33 $X2=0
+ $Y2=0
cc_195 N_VPWR_c_265_n N_A_399_368#_c_354_n 0.0090481f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_196 N_VPWR_M1009_d N_A_399_368#_c_361_n 0.00555074f $X=2.445 $Y=1.84 $X2=0
+ $Y2=0
cc_197 N_VPWR_c_269_n N_A_399_368#_c_361_n 0.0176063f $X=2.61 $Y=2.815 $X2=0
+ $Y2=0
cc_198 N_VPWR_c_265_n N_A_399_368#_c_361_n 0.0129605f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_199 N_VPWR_c_269_n N_A_399_368#_c_356_n 0.0168379f $X=2.61 $Y=2.815 $X2=0
+ $Y2=0
cc_200 N_VPWR_c_272_n N_A_399_368#_c_356_n 0.011066f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_201 N_VPWR_c_265_n N_A_399_368#_c_356_n 0.00915947f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_202 Y N_A_399_368#_M1005_d 0.0101062f $X=2.075 $Y=1.95 $X2=-0.19 $Y2=-0.245
cc_203 N_Y_c_312_n N_A_399_368#_c_354_n 0.0275831f $X=1.695 $Y=1.985 $X2=0 $Y2=0
cc_204 Y N_A_399_368#_c_361_n 5.73355e-19 $X=2.075 $Y=1.95 $X2=0 $Y2=0
cc_205 Y N_A_399_368#_c_359_n 0.0180102f $X=2.075 $Y=1.95 $X2=0 $Y2=0
cc_206 N_Y_c_312_n N_A_399_368#_c_359_n 0.0102884f $X=1.695 $Y=1.985 $X2=0 $Y2=0
cc_207 N_Y_c_319_n N_VGND_c_385_n 0.00365772f $X=2.185 $Y=0.88 $X2=0 $Y2=0
cc_208 N_Y_c_309_n N_VGND_c_385_n 0.0144183f $X=2.15 $Y=0.515 $X2=0 $Y2=0
cc_209 N_Y_c_309_n N_VGND_c_387_n 0.011237f $X=2.15 $Y=0.515 $X2=0 $Y2=0
cc_210 N_Y_c_319_n N_VGND_c_388_n 3.80876e-19 $X=2.185 $Y=0.88 $X2=0 $Y2=0
cc_211 N_Y_c_309_n N_VGND_c_388_n 0.0159304f $X=2.15 $Y=0.515 $X2=0 $Y2=0
cc_212 N_Y_c_309_n N_VGND_c_389_n 0.00933388f $X=2.15 $Y=0.515 $X2=0 $Y2=0
