* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__a222oi_2 A1 A2 B1 B2 C1 C2 VGND VNB VPB VPWR Y
X0 Y C1 a_116_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_515_392# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 Y C1 a_137_74# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X3 Y B1 a_593_74# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X4 a_116_392# B2 a_515_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_137_74# C2 VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X6 VPWR A1 a_515_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 a_116_392# C2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 VGND C2 a_137_74# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X9 a_593_74# B2 VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X10 VPWR A2 a_515_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 a_116_392# B1 a_515_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 VGND B2 a_593_74# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X13 a_593_74# B1 Y VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X14 VGND A2 a_981_74# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X15 Y C2 a_116_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 a_981_74# A1 Y VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X17 Y A1 a_981_74# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X18 a_515_392# B2 a_116_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 a_515_392# B1 a_116_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X20 a_981_74# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X21 a_137_74# C1 Y VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X22 a_116_392# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X23 a_515_392# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends
