* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__sdfrtp_4 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
M1000 a_1236_138# a_1034_392# a_415_81# VPB phighvt w=420000u l=150000u
+  ad=2.709e+11p pd=2.97e+06u as=5.047e+11p ps=5.18e+06u
M1001 a_1236_138# RESET_B VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=3.41945e+12p ps=2.648e+07u
M1002 a_415_81# D a_340_464# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1003 a_1745_74# a_1034_392# a_1367_112# VNB nshort w=640000u l=150000u
+  ad=4.33e+11p pd=3.08e+06u as=2.33e+11p ps=2.13e+06u
M1004 VPWR a_2339_74# Q VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=6.72e+11p ps=5.68e+06u
M1005 a_312_81# a_27_74# a_225_81# VNB nshort w=420000u l=150000u
+  ad=1.533e+11p pd=1.57e+06u as=2.373e+11p ps=2.81e+06u
M1006 a_415_81# D a_312_81# VNB nshort w=420000u l=150000u
+  ad=3.78e+11p pd=3.48e+06u as=0p ps=0u
M1007 VGND a_2339_74# Q VNB nshort w=740000u l=150000u
+  ad=2.36135e+12p pd=1.755e+07u as=4.144e+11p ps=4.08e+06u
M1008 a_1342_463# a_837_98# a_1236_138# VPB phighvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1009 VPWR a_1367_112# a_1342_463# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND CLK a_837_98# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.42325e+11p ps=2.38e+06u
M1011 VGND a_1745_74# a_2339_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1012 VGND RESET_B a_225_81# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_1034_392# a_837_98# VGND VNB nshort w=740000u l=150000u
+  ad=1.961e+11p pd=2.01e+06u as=0p ps=0u
M1014 a_514_464# a_27_74# a_415_81# VPB phighvt w=640000u l=150000u
+  ad=2.496e+11p pd=2.06e+06u as=0p ps=0u
M1015 a_2003_48# RESET_B VPWR VPB phighvt w=420000u l=150000u
+  ad=1.617e+11p pd=1.61e+06u as=0p ps=0u
M1016 Q a_2339_74# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 Q a_2339_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_1982_508# a_1034_392# a_1745_74# VPB phighvt w=420000u l=150000u
+  ad=1.134e+11p pd=1.38e+06u as=4.28275e+11p ps=3.57e+06u
M1019 a_1367_112# a_1236_138# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_2003_48# a_1745_74# a_2141_74# VNB nshort w=420000u l=150000u
+  ad=1.512e+11p pd=1.56e+06u as=8.82e+10p ps=1.26e+06u
M1021 VGND a_2003_48# a_1955_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1022 Q a_2339_74# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VPWR SCE a_27_74# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.888e+11p ps=1.87e+06u
M1024 VGND RESET_B a_1397_138# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1025 VPWR a_2339_74# Q VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_340_464# SCE VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_1955_74# a_837_98# a_1745_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VGND a_2339_74# Q VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPWR SCD a_514_464# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VPWR CLK a_837_98# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.95e+11p ps=2.59e+06u
M1031 a_1367_112# a_1236_138# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=3e+11p pd=2.6e+06u as=0p ps=0u
M1032 a_1236_138# a_837_98# a_415_81# VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1033 a_2339_74# a_1745_74# VPWR VPB phighvt w=840000u l=150000u
+  ad=2.52e+11p pd=2.28e+06u as=0p ps=0u
M1034 a_1034_392# a_837_98# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.95e+11p pd=2.59e+06u as=0p ps=0u
M1035 VPWR a_1745_74# a_2003_48# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 VGND SCE a_27_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1037 a_572_81# SCE a_415_81# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1038 a_2141_74# RESET_B VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 Q a_2339_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1040 a_225_81# SCD a_572_81# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1041 a_1322_138# a_1034_392# a_1236_138# VNB nshort w=420000u l=150000u
+  ad=9.45e+10p pd=1.29e+06u as=0p ps=0u
M1042 a_1745_74# a_837_98# a_1367_112# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1043 VPWR a_2003_48# a_1982_508# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1044 a_1397_138# a_1367_112# a_1322_138# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1045 a_415_81# RESET_B VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1046 VPWR a_1745_74# a_2339_74# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
