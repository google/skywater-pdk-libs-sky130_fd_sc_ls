* NGSPICE file created from sky130_fd_sc_ls__bufinv_16.ext - technology: sky130A

.subckt sky130_fd_sc_ls__bufinv_16 A VGND VNB VPB VPWR Y
M1000 VGND a_384_74# Y VNB nshort w=740000u l=150000u
+  ad=3.2079e+12p pd=2.791e+07u as=1.6576e+12p ps=1.632e+07u
M1001 Y a_384_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=2.7328e+12p pd=2.28e+07u as=4.4856e+12p ps=3.713e+07u
M1002 Y a_384_74# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_384_74# a_27_74# VGND VNB nshort w=740000u l=150000u
+  ad=6.216e+11p pd=6.12e+06u as=0p ps=0u
M1004 VPWR a_27_74# a_384_74# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=1.0304e+12p ps=8.56e+06u
M1005 VGND a_384_74# Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y a_384_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND a_27_74# a_384_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND a_27_74# a_384_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y a_384_74# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR a_384_74# Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Y a_384_74# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Y a_384_74# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR a_384_74# Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_384_74# a_27_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y a_384_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND a_27_74# a_384_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR a_384_74# Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND a_384_74# Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND a_384_74# Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 Y a_384_74# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPWR A a_27_74# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=6.664e+11p ps=5.67e+06u
M1022 a_27_74# A VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 Y a_384_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 Y a_384_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VGND A a_27_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=4.181e+11p ps=4.09e+06u
M1026 Y a_384_74# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VPWR a_27_74# a_384_74# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VPWR a_384_74# Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 Y a_384_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VGND a_384_74# Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 Y a_384_74# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 VGND a_384_74# Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VGND a_384_74# Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 VPWR A a_27_74# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 VPWR a_27_74# a_384_74# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 Y a_384_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 VPWR a_384_74# Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 VGND a_384_74# Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 VPWR a_384_74# Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1040 Y a_384_74# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1041 VGND A a_27_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1042 Y a_384_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1043 VPWR a_384_74# Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1044 a_384_74# a_27_74# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1045 a_384_74# a_27_74# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1046 a_384_74# a_27_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1047 VPWR a_384_74# Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1048 a_384_74# a_27_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1049 a_27_74# A VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

