* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__einvn_4 A TE_B VGND VNB VPB VPWR Z
M1000 a_281_74# A Z VNB nshort w=740000u l=150000u
+  ad=1.0508e+12p pd=1.024e+07u as=4.144e+11p ps=4.08e+06u
M1001 Z A a_241_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=6.72e+11p pd=5.68e+06u as=1.6688e+12p ps=1.418e+07u
M1002 a_281_74# a_114_74# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=6.253e+11p ps=6.13e+06u
M1003 VGND a_114_74# a_281_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_281_74# A Z VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_241_368# A Z VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_114_74# TE_B VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=1.0584e+12p ps=8.61e+06u
M1007 a_241_368# TE_B VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Z A a_281_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_281_74# a_114_74# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 Z A a_241_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR TE_B a_241_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR TE_B a_241_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_114_74# TE_B VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1014 a_241_368# A Z VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Z A a_281_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND a_114_74# a_281_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_241_368# TE_B VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
