* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
M1000 a_85_270# C1 a_600_392# VPB phighvt w=1e+06u l=150000u
+  ad=2.75e+11p pd=2.55e+06u as=2.7e+11p ps=2.54e+06u
M1001 a_600_392# B1 a_317_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=5.75e+11p ps=5.15e+06u
M1002 a_399_74# A2 VGND VNB nshort w=740000u l=150000u
+  ad=1.554e+11p pd=1.9e+06u as=9.731e+11p ps=7.07e+06u
M1003 VGND a_85_270# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.072e+11p ps=2.04e+06u
M1004 VPWR a_85_270# X VPB phighvt w=1.12e+06u l=150000u
+  ad=1.006e+12p pd=8.36e+06u as=3.36e+11p ps=2.84e+06u
M1005 X a_85_270# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND B1 a_85_270# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=4.847e+11p ps=4.27e+06u
M1007 VPWR A2 a_317_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_85_270# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_85_270# C1 VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_317_392# A1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_85_270# A1 a_399_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
