* File: sky130_fd_sc_ls__o41a_4.pxi.spice
* Created: Fri Aug 28 13:55:55 2020
* 
x_PM_SKY130_FD_SC_LS__O41A_4%A_110_48# N_A_110_48#_M1003_s N_A_110_48#_M1010_d
+ N_A_110_48#_M1022_s N_A_110_48#_M1006_g N_A_110_48#_c_151_n
+ N_A_110_48#_M1000_g N_A_110_48#_M1012_g N_A_110_48#_c_152_n
+ N_A_110_48#_M1004_g N_A_110_48#_M1016_g N_A_110_48#_c_153_n
+ N_A_110_48#_M1014_g N_A_110_48#_M1024_g N_A_110_48#_c_154_n
+ N_A_110_48#_M1021_g N_A_110_48#_c_147_n N_A_110_48#_c_148_n
+ N_A_110_48#_c_149_n N_A_110_48#_c_159_p N_A_110_48#_c_150_n
+ N_A_110_48#_c_156_n N_A_110_48#_c_157_n PM_SKY130_FD_SC_LS__O41A_4%A_110_48#
x_PM_SKY130_FD_SC_LS__O41A_4%B1 N_B1_c_273_n N_B1_c_279_n N_B1_M1010_g
+ N_B1_M1003_g N_B1_c_280_n N_B1_M1018_g N_B1_M1011_g B1 B1 N_B1_c_277_n
+ PM_SKY130_FD_SC_LS__O41A_4%B1
x_PM_SKY130_FD_SC_LS__O41A_4%A4 N_A4_c_335_n N_A4_M1022_g N_A4_c_331_n
+ N_A4_M1001_g N_A4_c_336_n N_A4_M1025_g N_A4_c_332_n N_A4_M1026_g A4 A4
+ N_A4_c_334_n PM_SKY130_FD_SC_LS__O41A_4%A4
x_PM_SKY130_FD_SC_LS__O41A_4%A3 N_A3_M1002_g N_A3_c_384_n N_A3_c_385_n
+ N_A3_c_393_n N_A3_M1015_g N_A3_c_386_n N_A3_c_387_n N_A3_c_388_n N_A3_M1013_g
+ N_A3_c_395_n N_A3_M1019_g A3 N_A3_c_390_n N_A3_c_391_n
+ PM_SKY130_FD_SC_LS__O41A_4%A3
x_PM_SKY130_FD_SC_LS__O41A_4%A1 N_A1_c_465_n N_A1_M1007_g N_A1_c_469_n
+ N_A1_M1008_g N_A1_c_466_n N_A1_M1009_g N_A1_c_470_n N_A1_M1027_g A1 A1
+ N_A1_c_468_n PM_SKY130_FD_SC_LS__O41A_4%A1
x_PM_SKY130_FD_SC_LS__O41A_4%A2 N_A2_M1005_g N_A2_c_519_n N_A2_c_520_n
+ N_A2_c_528_n N_A2_M1017_g N_A2_c_521_n N_A2_c_522_n N_A2_M1020_g N_A2_c_524_n
+ N_A2_c_530_n N_A2_M1023_g N_A2_c_525_n A2 PM_SKY130_FD_SC_LS__O41A_4%A2
x_PM_SKY130_FD_SC_LS__O41A_4%VPWR N_VPWR_M1000_s N_VPWR_M1004_s N_VPWR_M1021_s
+ N_VPWR_M1018_s N_VPWR_M1008_s N_VPWR_c_590_n N_VPWR_c_591_n N_VPWR_c_592_n
+ N_VPWR_c_593_n N_VPWR_c_594_n N_VPWR_c_595_n N_VPWR_c_596_n N_VPWR_c_597_n
+ N_VPWR_c_598_n N_VPWR_c_599_n N_VPWR_c_600_n N_VPWR_c_601_n N_VPWR_c_602_n
+ N_VPWR_c_603_n N_VPWR_c_604_n VPWR N_VPWR_c_605_n N_VPWR_c_589_n
+ PM_SKY130_FD_SC_LS__O41A_4%VPWR
x_PM_SKY130_FD_SC_LS__O41A_4%X N_X_M1006_d N_X_M1016_d N_X_M1000_d N_X_M1014_d
+ N_X_c_687_n N_X_c_702_n N_X_c_688_n N_X_c_692_n N_X_c_689_n N_X_c_693_n
+ N_X_c_712_n N_X_c_694_n N_X_c_690_n N_X_c_695_n N_X_c_696_n N_X_c_728_n
+ N_X_c_697_n X X X PM_SKY130_FD_SC_LS__O41A_4%X
x_PM_SKY130_FD_SC_LS__O41A_4%A_762_368# N_A_762_368#_M1015_d
+ N_A_762_368#_M1019_d N_A_762_368#_M1023_d N_A_762_368#_c_773_n
+ N_A_762_368#_c_767_n N_A_762_368#_c_783_n N_A_762_368#_c_786_n
+ N_A_762_368#_c_768_n N_A_762_368#_c_769_n N_A_762_368#_c_770_n
+ N_A_762_368#_c_771_n PM_SKY130_FD_SC_LS__O41A_4%A_762_368#
x_PM_SKY130_FD_SC_LS__O41A_4%A_851_368# N_A_851_368#_M1015_s
+ N_A_851_368#_M1025_d N_A_851_368#_c_821_n
+ PM_SKY130_FD_SC_LS__O41A_4%A_851_368#
x_PM_SKY130_FD_SC_LS__O41A_4%A_1213_368# N_A_1213_368#_M1017_s
+ N_A_1213_368#_M1027_d N_A_1213_368#_c_837_n N_A_1213_368#_c_835_n
+ N_A_1213_368#_c_836_n PM_SKY130_FD_SC_LS__O41A_4%A_1213_368#
x_PM_SKY130_FD_SC_LS__O41A_4%VGND N_VGND_M1006_s N_VGND_M1012_s N_VGND_M1024_s
+ N_VGND_M1002_s N_VGND_M1026_s N_VGND_M1005_s N_VGND_M1009_s N_VGND_c_859_n
+ N_VGND_c_860_n N_VGND_c_861_n N_VGND_c_862_n N_VGND_c_863_n N_VGND_c_864_n
+ N_VGND_c_865_n N_VGND_c_866_n N_VGND_c_867_n N_VGND_c_868_n N_VGND_c_869_n
+ N_VGND_c_870_n N_VGND_c_871_n N_VGND_c_872_n N_VGND_c_873_n VGND
+ N_VGND_c_874_n N_VGND_c_875_n N_VGND_c_876_n N_VGND_c_877_n N_VGND_c_878_n
+ N_VGND_c_879_n N_VGND_c_880_n PM_SKY130_FD_SC_LS__O41A_4%VGND
x_PM_SKY130_FD_SC_LS__O41A_4%A_523_124# N_A_523_124#_M1003_d
+ N_A_523_124#_M1011_d N_A_523_124#_M1001_d N_A_523_124#_M1013_d
+ N_A_523_124#_M1007_d N_A_523_124#_M1020_d N_A_523_124#_c_980_n
+ N_A_523_124#_c_981_n N_A_523_124#_c_982_n N_A_523_124#_c_983_n
+ N_A_523_124#_c_984_n N_A_523_124#_c_985_n N_A_523_124#_c_986_n
+ N_A_523_124#_c_987_n N_A_523_124#_c_988_n N_A_523_124#_c_989_n
+ N_A_523_124#_c_990_n N_A_523_124#_c_991_n N_A_523_124#_c_1042_n
+ N_A_523_124#_c_992_n N_A_523_124#_c_993_n N_A_523_124#_c_994_n
+ PM_SKY130_FD_SC_LS__O41A_4%A_523_124#
cc_1 VNB N_A_110_48#_M1006_g 0.021193f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=0.74
cc_2 VNB N_A_110_48#_M1012_g 0.0198267f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=0.74
cc_3 VNB N_A_110_48#_M1016_g 0.0203883f $X=-0.19 $Y=-0.245 $X2=1.555 $Y2=0.74
cc_4 VNB N_A_110_48#_M1024_g 0.0257334f $X=-0.19 $Y=-0.245 $X2=1.985 $Y2=0.74
cc_5 VNB N_A_110_48#_c_147_n 0.0185991f $X=-0.19 $Y=-0.245 $X2=2.78 $Y2=1.435
cc_6 VNB N_A_110_48#_c_148_n 0.130969f $X=-0.19 $Y=-0.245 $X2=2.11 $Y2=1.435
cc_7 VNB N_A_110_48#_c_149_n 0.00727972f $X=-0.19 $Y=-0.245 $X2=2.945 $Y2=1.6
cc_8 VNB N_A_110_48#_c_150_n 0.00170949f $X=-0.19 $Y=-0.245 $X2=3.19 $Y2=0.765
cc_9 VNB N_B1_c_273_n 0.00366516f $X=-0.19 $Y=-0.245 $X2=2.795 $Y2=1.93
cc_10 VNB N_B1_M1003_g 0.0213334f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_B1_M1011_g 0.020157f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=2.4
cc_12 VNB B1 0.00226907f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=0.74
cc_13 VNB N_B1_c_277_n 0.0427963f $X=-0.19 $Y=-0.245 $X2=1.555 $Y2=1.27
cc_14 VNB N_A4_c_331_n 0.0175218f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A4_c_332_n 0.0139587f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.27
cc_16 VNB A4 0.00518079f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=1.765
cc_17 VNB N_A4_c_334_n 0.0350844f $X=-0.19 $Y=-0.245 $X2=1.285 $Y2=2.4
cc_18 VNB N_A3_M1002_g 0.00753503f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A3_c_384_n 0.0256535f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A3_c_385_n 0.00980353f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A3_c_386_n 0.0989471f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.27
cc_22 VNB N_A3_c_387_n 0.00583879f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=0.74
cc_23 VNB N_A3_c_388_n 0.0144043f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A3_M1013_g 0.0235342f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=1.27
cc_25 VNB N_A3_c_390_n 0.0503978f $X=-0.19 $Y=-0.245 $X2=1.735 $Y2=1.765
cc_26 VNB N_A3_c_391_n 7.54705e-19 $X=-0.19 $Y=-0.245 $X2=1.985 $Y2=0.74
cc_27 VNB N_A1_c_465_n 0.0147706f $X=-0.19 $Y=-0.245 $X2=3.05 $Y2=0.62
cc_28 VNB N_A1_c_466_n 0.0146138f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB A1 0.00730714f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=1.765
cc_30 VNB N_A1_c_468_n 0.0356751f $X=-0.19 $Y=-0.245 $X2=1.285 $Y2=2.4
cc_31 VNB N_A2_M1005_g 0.0235707f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A2_c_519_n 0.00578033f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A2_c_520_n 0.0142072f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A2_c_521_n 0.137982f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.27
cc_35 VNB N_A2_c_522_n 0.00954688f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=0.74
cc_36 VNB N_A2_M1020_g 0.01277f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=2.4
cc_37 VNB N_A2_c_524_n 0.0158535f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=1.27
cc_38 VNB N_A2_c_525_n 0.0202215f $X=-0.19 $Y=-0.245 $X2=1.285 $Y2=2.4
cc_39 VNB A2 0.0401964f $X=-0.19 $Y=-0.245 $X2=1.555 $Y2=1.27
cc_40 VNB N_VPWR_c_589_n 0.342803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_X_c_687_n 0.0274757f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=1.765
cc_42 VNB N_X_c_688_n 0.00961898f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=2.4
cc_43 VNB N_X_c_689_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=1.285 $Y2=1.765
cc_44 VNB N_X_c_690_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=2.185 $Y2=1.765
cc_45 VNB N_VGND_c_859_n 0.0141307f $X=-0.19 $Y=-0.245 $X2=1.285 $Y2=2.4
cc_46 VNB N_VGND_c_860_n 0.0274339f $X=-0.19 $Y=-0.245 $X2=1.555 $Y2=1.27
cc_47 VNB N_VGND_c_861_n 0.00494723f $X=-0.19 $Y=-0.245 $X2=1.735 $Y2=1.765
cc_48 VNB N_VGND_c_862_n 0.0143472f $X=-0.19 $Y=-0.245 $X2=1.985 $Y2=0.74
cc_49 VNB N_VGND_c_863_n 0.00781633f $X=-0.19 $Y=-0.245 $X2=2.185 $Y2=2.4
cc_50 VNB N_VGND_c_864_n 0.00341672f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.435
cc_51 VNB N_VGND_c_865_n 0.00469205f $X=-0.19 $Y=-0.245 $X2=2.11 $Y2=1.435
cc_52 VNB N_VGND_c_866_n 0.0160886f $X=-0.19 $Y=-0.245 $X2=2.945 $Y2=1.6
cc_53 VNB N_VGND_c_867_n 0.0061168f $X=-0.19 $Y=-0.245 $X2=3.19 $Y2=1.1
cc_54 VNB N_VGND_c_868_n 0.0492942f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_869_n 0.00229531f $X=-0.19 $Y=-0.245 $X2=3.11 $Y2=2.035
cc_56 VNB N_VGND_c_870_n 0.0160886f $X=-0.19 $Y=-0.245 $X2=4.86 $Y2=2.035
cc_57 VNB N_VGND_c_871_n 0.00445561f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_872_n 0.0142087f $X=-0.19 $Y=-0.245 $X2=3.027 $Y2=1.435
cc_59 VNB N_VGND_c_873_n 0.00337546f $X=-0.19 $Y=-0.245 $X2=2.945 $Y2=2.035
cc_60 VNB N_VGND_c_874_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.517
cc_61 VNB N_VGND_c_875_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=1.735 $Y2=1.517
cc_62 VNB N_VGND_c_876_n 0.0272543f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_877_n 0.437198f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_878_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_879_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_880_n 0.00337546f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_523_124#_c_980_n 0.00615577f $X=-0.19 $Y=-0.245 $X2=1.285
+ $Y2=1.765
cc_68 VNB N_A_523_124#_c_981_n 0.0156685f $X=-0.19 $Y=-0.245 $X2=1.285 $Y2=2.4
cc_69 VNB N_A_523_124#_c_982_n 0.00497327f $X=-0.19 $Y=-0.245 $X2=1.555 $Y2=1.27
cc_70 VNB N_A_523_124#_c_983_n 0.00215445f $X=-0.19 $Y=-0.245 $X2=1.735
+ $Y2=1.765
cc_71 VNB N_A_523_124#_c_984_n 0.00737922f $X=-0.19 $Y=-0.245 $X2=1.735 $Y2=2.4
cc_72 VNB N_A_523_124#_c_985_n 0.00178935f $X=-0.19 $Y=-0.245 $X2=1.735 $Y2=2.4
cc_73 VNB N_A_523_124#_c_986_n 0.001978f $X=-0.19 $Y=-0.245 $X2=1.985 $Y2=0.74
cc_74 VNB N_A_523_124#_c_987_n 0.0112124f $X=-0.19 $Y=-0.245 $X2=2.185 $Y2=1.765
cc_75 VNB N_A_523_124#_c_988_n 0.00254618f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.435
cc_76 VNB N_A_523_124#_c_989_n 0.0105793f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.435
cc_77 VNB N_A_523_124#_c_990_n 0.00197771f $X=-0.19 $Y=-0.245 $X2=2.11 $Y2=1.435
cc_78 VNB N_A_523_124#_c_991_n 0.00525165f $X=-0.19 $Y=-0.245 $X2=2.945 $Y2=1.95
cc_79 VNB N_A_523_124#_c_992_n 0.00176133f $X=-0.19 $Y=-0.245 $X2=3.19 $Y2=0.765
cc_80 VNB N_A_523_124#_c_993_n 0.00322493f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_523_124#_c_994_n 0.00176197f $X=-0.19 $Y=-0.245 $X2=3.11 $Y2=2.035
cc_82 VPB N_A_110_48#_c_151_n 0.0163425f $X=-0.19 $Y=1.66 $X2=0.835 $Y2=1.765
cc_83 VPB N_A_110_48#_c_152_n 0.014923f $X=-0.19 $Y=1.66 $X2=1.285 $Y2=1.765
cc_84 VPB N_A_110_48#_c_153_n 0.014923f $X=-0.19 $Y=1.66 $X2=1.735 $Y2=1.765
cc_85 VPB N_A_110_48#_c_154_n 0.0160623f $X=-0.19 $Y=1.66 $X2=2.185 $Y2=1.765
cc_86 VPB N_A_110_48#_c_148_n 0.0273508f $X=-0.19 $Y=1.66 $X2=2.11 $Y2=1.435
cc_87 VPB N_A_110_48#_c_156_n 0.0122307f $X=-0.19 $Y=1.66 $X2=4.86 $Y2=2.035
cc_88 VPB N_A_110_48#_c_157_n 0.00348908f $X=-0.19 $Y=1.66 $X2=2.945 $Y2=2.075
cc_89 VPB N_B1_c_273_n 0.00561444f $X=-0.19 $Y=1.66 $X2=2.795 $Y2=1.93
cc_90 VPB N_B1_c_279_n 0.0216677f $X=-0.19 $Y=1.66 $X2=4.705 $Y2=1.84
cc_91 VPB N_B1_c_280_n 0.0172387f $X=-0.19 $Y=1.66 $X2=0.625 $Y2=1.27
cc_92 VPB B1 0.00822915f $X=-0.19 $Y=1.66 $X2=1.055 $Y2=0.74
cc_93 VPB N_B1_c_277_n 0.0270852f $X=-0.19 $Y=1.66 $X2=1.555 $Y2=1.27
cc_94 VPB N_A4_c_335_n 0.0158167f $X=-0.19 $Y=1.66 $X2=3.05 $Y2=0.62
cc_95 VPB N_A4_c_336_n 0.0158158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB A4 0.00642706f $X=-0.19 $Y=1.66 $X2=0.835 $Y2=1.765
cc_97 VPB N_A4_c_334_n 0.0201835f $X=-0.19 $Y=1.66 $X2=1.285 $Y2=2.4
cc_98 VPB N_A3_c_385_n 7.88789e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB N_A3_c_393_n 0.0250147f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 VPB N_A3_c_388_n 7.9375e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB N_A3_c_395_n 0.0223576f $X=-0.19 $Y=1.66 $X2=1.055 $Y2=0.74
cc_102 VPB N_A1_c_469_n 0.0160979f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 VPB N_A1_c_470_n 0.0159848f $X=-0.19 $Y=1.66 $X2=0.625 $Y2=1.27
cc_104 VPB A1 0.00704168f $X=-0.19 $Y=1.66 $X2=0.835 $Y2=1.765
cc_105 VPB N_A1_c_468_n 0.0212176f $X=-0.19 $Y=1.66 $X2=1.285 $Y2=2.4
cc_106 VPB N_A2_c_520_n 7.82949e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB N_A2_c_528_n 0.0221241f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_A2_c_524_n 0.00122646f $X=-0.19 $Y=1.66 $X2=1.055 $Y2=1.27
cc_109 VPB N_A2_c_530_n 0.0301829f $X=-0.19 $Y=1.66 $X2=1.055 $Y2=0.74
cc_110 VPB N_VPWR_c_590_n 0.0112087f $X=-0.19 $Y=1.66 $X2=1.055 $Y2=0.74
cc_111 VPB N_VPWR_c_591_n 0.00799266f $X=-0.19 $Y=1.66 $X2=1.285 $Y2=2.4
cc_112 VPB N_VPWR_c_592_n 0.0163625f $X=-0.19 $Y=1.66 $X2=1.555 $Y2=0.74
cc_113 VPB N_VPWR_c_593_n 0.0238169f $X=-0.19 $Y=1.66 $X2=1.735 $Y2=2.4
cc_114 VPB N_VPWR_c_594_n 0.00615639f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_VPWR_c_595_n 0.0173573f $X=-0.19 $Y=1.66 $X2=2.185 $Y2=2.4
cc_116 VPB N_VPWR_c_596_n 0.00324402f $X=-0.19 $Y=1.66 $X2=2.78 $Y2=1.435
cc_117 VPB N_VPWR_c_597_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0.75 $Y2=1.435
cc_118 VPB N_VPWR_c_598_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0.75 $Y2=1.435
cc_119 VPB N_VPWR_c_599_n 0.0206041f $X=-0.19 $Y=1.66 $X2=2.11 $Y2=1.435
cc_120 VPB N_VPWR_c_600_n 0.0047828f $X=-0.19 $Y=1.66 $X2=2.11 $Y2=1.435
cc_121 VPB N_VPWR_c_601_n 0.0215627f $X=-0.19 $Y=1.66 $X2=2.945 $Y2=1.6
cc_122 VPB N_VPWR_c_602_n 0.0047828f $X=-0.19 $Y=1.66 $X2=2.945 $Y2=1.95
cc_123 VPB N_VPWR_c_603_n 0.0805589f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_604_n 0.00537188f $X=-0.19 $Y=1.66 $X2=3.19 $Y2=1.1
cc_125 VPB N_VPWR_c_605_n 0.037911f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_589_n 0.131544f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_127 VPB N_X_c_687_n 0.00570873f $X=-0.19 $Y=1.66 $X2=0.835 $Y2=1.765
cc_128 VPB N_X_c_692_n 0.00897441f $X=-0.19 $Y=1.66 $X2=1.055 $Y2=1.27
cc_129 VPB N_X_c_693_n 0.00257348f $X=-0.19 $Y=1.66 $X2=1.555 $Y2=0.74
cc_130 VPB N_X_c_694_n 0.00362934f $X=-0.19 $Y=1.66 $X2=1.985 $Y2=1.27
cc_131 VPB N_X_c_695_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0.75 $Y2=1.435
cc_132 VPB N_X_c_696_n 0.00928121f $X=-0.19 $Y=1.66 $X2=2.11 $Y2=1.435
cc_133 VPB N_X_c_697_n 0.00183442f $X=-0.19 $Y=1.66 $X2=2.945 $Y2=1.6
cc_134 VPB X 0.0510143f $X=-0.19 $Y=1.66 $X2=2.945 $Y2=1.95
cc_135 VPB N_A_762_368#_c_767_n 0.00310361f $X=-0.19 $Y=1.66 $X2=0.835 $Y2=1.765
cc_136 VPB N_A_762_368#_c_768_n 0.0233531f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_A_762_368#_c_769_n 0.0357641f $X=-0.19 $Y=1.66 $X2=1.285 $Y2=2.4
cc_138 VPB N_A_762_368#_c_770_n 0.00888879f $X=-0.19 $Y=1.66 $X2=1.555 $Y2=0.74
cc_139 VPB N_A_762_368#_c_771_n 0.00180293f $X=-0.19 $Y=1.66 $X2=1.735 $Y2=2.4
cc_140 VPB N_A_851_368#_c_821_n 0.00772388f $X=-0.19 $Y=1.66 $X2=0.625 $Y2=0.74
cc_141 VPB N_A_1213_368#_c_835_n 0.00257417f $X=-0.19 $Y=1.66 $X2=0.835
+ $Y2=1.765
cc_142 VPB N_A_1213_368#_c_836_n 0.00289794f $X=-0.19 $Y=1.66 $X2=0.835 $Y2=2.4
cc_143 N_A_110_48#_c_147_n N_B1_c_273_n 0.00726507f $X=2.78 $Y=1.435 $X2=0 $Y2=0
cc_144 N_A_110_48#_c_159_p N_B1_c_273_n 0.00522018f $X=2.945 $Y=1.95 $X2=0 $Y2=0
cc_145 N_A_110_48#_c_154_n N_B1_c_279_n 0.0172138f $X=2.185 $Y=1.765 $X2=0 $Y2=0
cc_146 N_A_110_48#_c_159_p N_B1_c_279_n 0.00568468f $X=2.945 $Y=1.95 $X2=0 $Y2=0
cc_147 N_A_110_48#_c_157_n N_B1_c_279_n 0.0112303f $X=2.945 $Y=2.075 $X2=0 $Y2=0
cc_148 N_A_110_48#_c_148_n N_B1_M1003_g 0.00213441f $X=2.11 $Y=1.435 $X2=0 $Y2=0
cc_149 N_A_110_48#_c_149_n N_B1_M1003_g 0.0194369f $X=2.945 $Y=1.6 $X2=0 $Y2=0
cc_150 N_A_110_48#_c_159_p N_B1_c_280_n 0.00488611f $X=2.945 $Y=1.95 $X2=0 $Y2=0
cc_151 N_A_110_48#_c_156_n N_B1_c_280_n 0.0177821f $X=4.86 $Y=2.035 $X2=0 $Y2=0
cc_152 N_A_110_48#_c_157_n N_B1_c_280_n 0.015267f $X=2.945 $Y=2.075 $X2=0 $Y2=0
cc_153 N_A_110_48#_c_149_n N_B1_M1011_g 0.00448353f $X=2.945 $Y=1.6 $X2=0 $Y2=0
cc_154 N_A_110_48#_c_149_n B1 0.0134595f $X=2.945 $Y=1.6 $X2=0 $Y2=0
cc_155 N_A_110_48#_c_159_p B1 0.0142914f $X=2.945 $Y=1.95 $X2=0 $Y2=0
cc_156 N_A_110_48#_c_156_n B1 0.0683979f $X=4.86 $Y=2.035 $X2=0 $Y2=0
cc_157 N_A_110_48#_c_147_n N_B1_c_277_n 0.00691491f $X=2.78 $Y=1.435 $X2=0 $Y2=0
cc_158 N_A_110_48#_c_148_n N_B1_c_277_n 0.0114221f $X=2.11 $Y=1.435 $X2=0 $Y2=0
cc_159 N_A_110_48#_c_149_n N_B1_c_277_n 0.0162985f $X=2.945 $Y=1.6 $X2=0 $Y2=0
cc_160 N_A_110_48#_c_159_p N_B1_c_277_n 0.00961924f $X=2.945 $Y=1.95 $X2=0 $Y2=0
cc_161 N_A_110_48#_c_156_n N_B1_c_277_n 0.00219744f $X=4.86 $Y=2.035 $X2=0 $Y2=0
cc_162 N_A_110_48#_c_156_n N_A4_c_335_n 0.0085117f $X=4.86 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_163 N_A_110_48#_c_156_n N_A4_c_336_n 0.00353402f $X=4.86 $Y=2.035 $X2=0 $Y2=0
cc_164 N_A_110_48#_c_156_n A4 0.0385085f $X=4.86 $Y=2.035 $X2=0 $Y2=0
cc_165 N_A_110_48#_c_156_n N_A4_c_334_n 0.00136242f $X=4.86 $Y=2.035 $X2=0 $Y2=0
cc_166 N_A_110_48#_c_156_n N_A3_c_384_n 8.30342e-19 $X=4.86 $Y=2.035 $X2=0 $Y2=0
cc_167 N_A_110_48#_c_156_n N_A3_c_393_n 0.0143343f $X=4.86 $Y=2.035 $X2=0 $Y2=0
cc_168 N_A_110_48#_c_156_n N_A3_c_395_n 5.08733e-19 $X=4.86 $Y=2.035 $X2=0 $Y2=0
cc_169 N_A_110_48#_c_156_n N_VPWR_M1018_s 0.00584575f $X=4.86 $Y=2.035 $X2=0
+ $Y2=0
cc_170 N_A_110_48#_c_151_n N_VPWR_c_590_n 0.0101588f $X=0.835 $Y=1.765 $X2=0
+ $Y2=0
cc_171 N_A_110_48#_c_152_n N_VPWR_c_591_n 0.00609105f $X=1.285 $Y=1.765 $X2=0
+ $Y2=0
cc_172 N_A_110_48#_c_153_n N_VPWR_c_591_n 0.00609105f $X=1.735 $Y=1.765 $X2=0
+ $Y2=0
cc_173 N_A_110_48#_c_154_n N_VPWR_c_592_n 0.0108935f $X=2.185 $Y=1.765 $X2=0
+ $Y2=0
cc_174 N_A_110_48#_c_147_n N_VPWR_c_592_n 0.0140038f $X=2.78 $Y=1.435 $X2=0
+ $Y2=0
cc_175 N_A_110_48#_c_159_p N_VPWR_c_592_n 0.00262905f $X=2.945 $Y=1.95 $X2=0
+ $Y2=0
cc_176 N_A_110_48#_c_157_n N_VPWR_c_592_n 0.055952f $X=2.945 $Y=2.075 $X2=0
+ $Y2=0
cc_177 N_A_110_48#_c_156_n N_VPWR_c_593_n 0.0202358f $X=4.86 $Y=2.035 $X2=0
+ $Y2=0
cc_178 N_A_110_48#_c_157_n N_VPWR_c_593_n 0.0335551f $X=2.945 $Y=2.075 $X2=0
+ $Y2=0
cc_179 N_A_110_48#_c_151_n N_VPWR_c_597_n 0.00445602f $X=0.835 $Y=1.765 $X2=0
+ $Y2=0
cc_180 N_A_110_48#_c_152_n N_VPWR_c_597_n 0.00445602f $X=1.285 $Y=1.765 $X2=0
+ $Y2=0
cc_181 N_A_110_48#_c_153_n N_VPWR_c_599_n 0.00445602f $X=1.735 $Y=1.765 $X2=0
+ $Y2=0
cc_182 N_A_110_48#_c_154_n N_VPWR_c_599_n 0.00445602f $X=2.185 $Y=1.765 $X2=0
+ $Y2=0
cc_183 N_A_110_48#_c_157_n N_VPWR_c_601_n 0.00813904f $X=2.945 $Y=2.075 $X2=0
+ $Y2=0
cc_184 N_A_110_48#_c_151_n N_VPWR_c_589_n 0.00862391f $X=0.835 $Y=1.765 $X2=0
+ $Y2=0
cc_185 N_A_110_48#_c_152_n N_VPWR_c_589_n 0.00857589f $X=1.285 $Y=1.765 $X2=0
+ $Y2=0
cc_186 N_A_110_48#_c_153_n N_VPWR_c_589_n 0.00857589f $X=1.735 $Y=1.765 $X2=0
+ $Y2=0
cc_187 N_A_110_48#_c_154_n N_VPWR_c_589_n 0.00862391f $X=2.185 $Y=1.765 $X2=0
+ $Y2=0
cc_188 N_A_110_48#_c_157_n N_VPWR_c_589_n 0.0106351f $X=2.945 $Y=2.075 $X2=0
+ $Y2=0
cc_189 N_A_110_48#_M1006_g N_X_c_687_n 0.0135824f $X=0.625 $Y=0.74 $X2=0 $Y2=0
cc_190 N_A_110_48#_c_147_n N_X_c_687_n 0.0175348f $X=2.78 $Y=1.435 $X2=0 $Y2=0
cc_191 N_A_110_48#_c_148_n N_X_c_687_n 0.00429394f $X=2.11 $Y=1.435 $X2=0 $Y2=0
cc_192 N_A_110_48#_M1006_g N_X_c_702_n 0.0132299f $X=0.625 $Y=0.74 $X2=0 $Y2=0
cc_193 N_A_110_48#_c_147_n N_X_c_702_n 0.00639324f $X=2.78 $Y=1.435 $X2=0 $Y2=0
cc_194 N_A_110_48#_c_151_n N_X_c_692_n 0.01377f $X=0.835 $Y=1.765 $X2=0 $Y2=0
cc_195 N_A_110_48#_c_147_n N_X_c_692_n 0.022759f $X=2.78 $Y=1.435 $X2=0 $Y2=0
cc_196 N_A_110_48#_c_148_n N_X_c_692_n 0.00579333f $X=2.11 $Y=1.435 $X2=0 $Y2=0
cc_197 N_A_110_48#_M1006_g N_X_c_689_n 0.0121547f $X=0.625 $Y=0.74 $X2=0 $Y2=0
cc_198 N_A_110_48#_M1012_g N_X_c_689_n 2.71222e-19 $X=1.055 $Y=0.74 $X2=0 $Y2=0
cc_199 N_A_110_48#_c_151_n N_X_c_693_n 0.0135742f $X=0.835 $Y=1.765 $X2=0 $Y2=0
cc_200 N_A_110_48#_c_152_n N_X_c_693_n 0.0128074f $X=1.285 $Y=1.765 $X2=0 $Y2=0
cc_201 N_A_110_48#_c_153_n N_X_c_693_n 7.00309e-19 $X=1.735 $Y=1.765 $X2=0 $Y2=0
cc_202 N_A_110_48#_M1012_g N_X_c_712_n 0.0126527f $X=1.055 $Y=0.74 $X2=0 $Y2=0
cc_203 N_A_110_48#_M1016_g N_X_c_712_n 0.0122754f $X=1.555 $Y=0.74 $X2=0 $Y2=0
cc_204 N_A_110_48#_c_147_n N_X_c_712_n 0.061224f $X=2.78 $Y=1.435 $X2=0 $Y2=0
cc_205 N_A_110_48#_c_148_n N_X_c_712_n 0.00709665f $X=2.11 $Y=1.435 $X2=0 $Y2=0
cc_206 N_A_110_48#_c_152_n N_X_c_694_n 0.0120074f $X=1.285 $Y=1.765 $X2=0 $Y2=0
cc_207 N_A_110_48#_c_153_n N_X_c_694_n 0.0133289f $X=1.735 $Y=1.765 $X2=0 $Y2=0
cc_208 N_A_110_48#_c_154_n N_X_c_694_n 0.00410678f $X=2.185 $Y=1.765 $X2=0 $Y2=0
cc_209 N_A_110_48#_c_147_n N_X_c_694_n 0.0694546f $X=2.78 $Y=1.435 $X2=0 $Y2=0
cc_210 N_A_110_48#_c_148_n N_X_c_694_n 0.0161398f $X=2.11 $Y=1.435 $X2=0 $Y2=0
cc_211 N_A_110_48#_c_159_p N_X_c_694_n 0.00360245f $X=2.945 $Y=1.95 $X2=0 $Y2=0
cc_212 N_A_110_48#_M1012_g N_X_c_690_n 9.1509e-19 $X=1.055 $Y=0.74 $X2=0 $Y2=0
cc_213 N_A_110_48#_M1016_g N_X_c_690_n 0.00804372f $X=1.555 $Y=0.74 $X2=0 $Y2=0
cc_214 N_A_110_48#_M1024_g N_X_c_690_n 2.71222e-19 $X=1.985 $Y=0.74 $X2=0 $Y2=0
cc_215 N_A_110_48#_c_152_n N_X_c_695_n 7.00309e-19 $X=1.285 $Y=1.765 $X2=0 $Y2=0
cc_216 N_A_110_48#_c_153_n N_X_c_695_n 0.0128074f $X=1.735 $Y=1.765 $X2=0 $Y2=0
cc_217 N_A_110_48#_c_154_n N_X_c_695_n 0.0117511f $X=2.185 $Y=1.765 $X2=0 $Y2=0
cc_218 N_A_110_48#_M1006_g N_X_c_728_n 7.32094e-19 $X=0.625 $Y=0.74 $X2=0 $Y2=0
cc_219 N_A_110_48#_c_147_n N_X_c_728_n 0.0178863f $X=2.78 $Y=1.435 $X2=0 $Y2=0
cc_220 N_A_110_48#_c_148_n N_X_c_728_n 0.00272398f $X=2.11 $Y=1.435 $X2=0 $Y2=0
cc_221 N_A_110_48#_c_151_n N_X_c_697_n 0.00132156f $X=0.835 $Y=1.765 $X2=0 $Y2=0
cc_222 N_A_110_48#_c_152_n N_X_c_697_n 0.00132156f $X=1.285 $Y=1.765 $X2=0 $Y2=0
cc_223 N_A_110_48#_c_147_n N_X_c_697_n 0.0276943f $X=2.78 $Y=1.435 $X2=0 $Y2=0
cc_224 N_A_110_48#_c_148_n N_X_c_697_n 0.00835323f $X=2.11 $Y=1.435 $X2=0 $Y2=0
cc_225 N_A_110_48#_c_151_n X 0.00374056f $X=0.835 $Y=1.765 $X2=0 $Y2=0
cc_226 N_A_110_48#_c_156_n N_A_762_368#_M1015_d 0.00587962f $X=4.86 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_227 N_A_110_48#_M1022_s N_A_762_368#_c_773_n 0.00400315f $X=4.705 $Y=1.84
+ $X2=0 $Y2=0
cc_228 N_A_110_48#_c_156_n N_A_762_368#_c_773_n 0.0495398f $X=4.86 $Y=2.035
+ $X2=0 $Y2=0
cc_229 N_A_110_48#_c_156_n N_A_762_368#_c_767_n 0.00502396f $X=4.86 $Y=2.035
+ $X2=0 $Y2=0
cc_230 N_A_110_48#_c_156_n N_A_762_368#_c_770_n 0.0204259f $X=4.86 $Y=2.035
+ $X2=0 $Y2=0
cc_231 N_A_110_48#_c_156_n N_A_851_368#_M1015_s 0.0076215f $X=4.86 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_232 N_A_110_48#_M1022_s N_A_851_368#_c_821_n 0.00213554f $X=4.705 $Y=1.84
+ $X2=0 $Y2=0
cc_233 N_A_110_48#_M1006_g N_VGND_c_860_n 0.0111726f $X=0.625 $Y=0.74 $X2=0
+ $Y2=0
cc_234 N_A_110_48#_M1006_g N_VGND_c_861_n 4.80326e-19 $X=0.625 $Y=0.74 $X2=0
+ $Y2=0
cc_235 N_A_110_48#_M1012_g N_VGND_c_861_n 0.00877665f $X=1.055 $Y=0.74 $X2=0
+ $Y2=0
cc_236 N_A_110_48#_M1016_g N_VGND_c_861_n 0.00382194f $X=1.555 $Y=0.74 $X2=0
+ $Y2=0
cc_237 N_A_110_48#_M1016_g N_VGND_c_862_n 5.81525e-19 $X=1.555 $Y=0.74 $X2=0
+ $Y2=0
cc_238 N_A_110_48#_M1024_g N_VGND_c_862_n 0.0138071f $X=1.985 $Y=0.74 $X2=0
+ $Y2=0
cc_239 N_A_110_48#_c_147_n N_VGND_c_862_n 0.0248195f $X=2.78 $Y=1.435 $X2=0
+ $Y2=0
cc_240 N_A_110_48#_c_148_n N_VGND_c_862_n 0.00548538f $X=2.11 $Y=1.435 $X2=0
+ $Y2=0
cc_241 N_A_110_48#_M1006_g N_VGND_c_874_n 0.00434272f $X=0.625 $Y=0.74 $X2=0
+ $Y2=0
cc_242 N_A_110_48#_M1012_g N_VGND_c_874_n 0.00383152f $X=1.055 $Y=0.74 $X2=0
+ $Y2=0
cc_243 N_A_110_48#_M1016_g N_VGND_c_875_n 0.00434272f $X=1.555 $Y=0.74 $X2=0
+ $Y2=0
cc_244 N_A_110_48#_M1024_g N_VGND_c_875_n 0.00383152f $X=1.985 $Y=0.74 $X2=0
+ $Y2=0
cc_245 N_A_110_48#_M1006_g N_VGND_c_877_n 0.00824087f $X=0.625 $Y=0.74 $X2=0
+ $Y2=0
cc_246 N_A_110_48#_M1012_g N_VGND_c_877_n 0.0075754f $X=1.055 $Y=0.74 $X2=0
+ $Y2=0
cc_247 N_A_110_48#_M1016_g N_VGND_c_877_n 0.00820718f $X=1.555 $Y=0.74 $X2=0
+ $Y2=0
cc_248 N_A_110_48#_M1024_g N_VGND_c_877_n 0.0075754f $X=1.985 $Y=0.74 $X2=0
+ $Y2=0
cc_249 N_A_110_48#_M1024_g N_A_523_124#_c_980_n 9.31825e-19 $X=1.985 $Y=0.74
+ $X2=0 $Y2=0
cc_250 N_A_110_48#_c_147_n N_A_523_124#_c_980_n 0.00970275f $X=2.78 $Y=1.435
+ $X2=0 $Y2=0
cc_251 N_A_110_48#_c_149_n N_A_523_124#_c_980_n 0.0062953f $X=2.945 $Y=1.6 $X2=0
+ $Y2=0
cc_252 N_A_110_48#_c_150_n N_A_523_124#_c_980_n 0.0125142f $X=3.19 $Y=0.765
+ $X2=0 $Y2=0
cc_253 N_A_110_48#_c_149_n N_A_523_124#_c_981_n 0.00380631f $X=2.945 $Y=1.6
+ $X2=0 $Y2=0
cc_254 N_A_110_48#_c_150_n N_A_523_124#_c_981_n 0.0132727f $X=3.19 $Y=0.765
+ $X2=0 $Y2=0
cc_255 N_A_110_48#_M1024_g N_A_523_124#_c_982_n 5.9337e-19 $X=1.985 $Y=0.74
+ $X2=0 $Y2=0
cc_256 N_A_110_48#_c_150_n N_A_523_124#_c_983_n 0.0173112f $X=3.19 $Y=0.765
+ $X2=0 $Y2=0
cc_257 N_A_110_48#_c_149_n N_A_523_124#_c_985_n 0.00714719f $X=2.945 $Y=1.6
+ $X2=0 $Y2=0
cc_258 B1 A4 0.0224439f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_259 B1 N_A4_c_334_n 3.22268e-19 $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_260 B1 N_A3_c_384_n 0.0108947f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_261 N_B1_c_277_n N_A3_c_384_n 0.00250407f $X=3.405 $Y=1.647 $X2=0 $Y2=0
cc_262 B1 N_A3_c_385_n 0.00664537f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_263 N_B1_c_277_n N_A3_c_385_n 0.00580431f $X=3.405 $Y=1.647 $X2=0 $Y2=0
cc_264 B1 N_A3_c_393_n 0.00509853f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_265 N_B1_M1011_g N_A3_c_390_n 0.0197827f $X=3.405 $Y=0.94 $X2=0 $Y2=0
cc_266 N_B1_c_279_n N_VPWR_c_592_n 0.0107096f $X=2.72 $Y=1.855 $X2=0 $Y2=0
cc_267 N_B1_c_280_n N_VPWR_c_593_n 0.00822904f $X=3.17 $Y=1.855 $X2=0 $Y2=0
cc_268 N_B1_c_279_n N_VPWR_c_601_n 0.0044094f $X=2.72 $Y=1.855 $X2=0 $Y2=0
cc_269 N_B1_c_280_n N_VPWR_c_601_n 0.0044094f $X=3.17 $Y=1.855 $X2=0 $Y2=0
cc_270 N_B1_c_279_n N_VPWR_c_589_n 0.00487769f $X=2.72 $Y=1.855 $X2=0 $Y2=0
cc_271 N_B1_c_280_n N_VPWR_c_589_n 0.00487769f $X=3.17 $Y=1.855 $X2=0 $Y2=0
cc_272 N_B1_c_279_n N_X_c_694_n 4.41799e-19 $X=2.72 $Y=1.855 $X2=0 $Y2=0
cc_273 N_B1_M1003_g N_VGND_c_862_n 0.00500871f $X=2.975 $Y=0.94 $X2=0 $Y2=0
cc_274 N_B1_M1003_g N_VGND_c_868_n 2.27419e-19 $X=2.975 $Y=0.94 $X2=0 $Y2=0
cc_275 N_B1_M1011_g N_VGND_c_868_n 2.27419e-19 $X=3.405 $Y=0.94 $X2=0 $Y2=0
cc_276 N_B1_M1003_g N_A_523_124#_c_980_n 0.00888778f $X=2.975 $Y=0.94 $X2=0
+ $Y2=0
cc_277 N_B1_M1011_g N_A_523_124#_c_980_n 4.22299e-19 $X=3.405 $Y=0.94 $X2=0
+ $Y2=0
cc_278 N_B1_c_277_n N_A_523_124#_c_980_n 0.00125689f $X=3.405 $Y=1.647 $X2=0
+ $Y2=0
cc_279 N_B1_M1003_g N_A_523_124#_c_981_n 0.0046393f $X=2.975 $Y=0.94 $X2=0 $Y2=0
cc_280 N_B1_M1011_g N_A_523_124#_c_981_n 0.00582977f $X=3.405 $Y=0.94 $X2=0
+ $Y2=0
cc_281 N_B1_M1003_g N_A_523_124#_c_983_n 4.69875e-19 $X=2.975 $Y=0.94 $X2=0
+ $Y2=0
cc_282 N_B1_M1011_g N_A_523_124#_c_983_n 0.00880445f $X=3.405 $Y=0.94 $X2=0
+ $Y2=0
cc_283 B1 N_A_523_124#_c_984_n 0.03029f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_284 N_B1_M1011_g N_A_523_124#_c_985_n 0.00236422f $X=3.405 $Y=0.94 $X2=0
+ $Y2=0
cc_285 B1 N_A_523_124#_c_985_n 0.0213654f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_286 N_B1_c_277_n N_A_523_124#_c_985_n 0.00302844f $X=3.405 $Y=1.647 $X2=0
+ $Y2=0
cc_287 N_A4_c_331_n N_A3_M1002_g 0.00814159f $X=4.675 $Y=1.35 $X2=0 $Y2=0
cc_288 N_A4_c_331_n N_A3_c_384_n 6.90332e-19 $X=4.675 $Y=1.35 $X2=0 $Y2=0
cc_289 A4 N_A3_c_384_n 0.00282722f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_290 N_A4_c_334_n N_A3_c_384_n 0.0183984f $X=5.09 $Y=1.557 $X2=0 $Y2=0
cc_291 N_A4_c_335_n N_A3_c_393_n 0.0433698f $X=4.63 $Y=1.765 $X2=0 $Y2=0
cc_292 N_A4_c_334_n N_A3_c_393_n 0.00367105f $X=5.09 $Y=1.557 $X2=0 $Y2=0
cc_293 N_A4_c_331_n N_A3_c_386_n 0.0103098f $X=4.675 $Y=1.35 $X2=0 $Y2=0
cc_294 N_A4_c_332_n N_A3_c_386_n 0.0103186f $X=5.105 $Y=1.35 $X2=0 $Y2=0
cc_295 N_A4_c_332_n N_A3_c_387_n 0.0106756f $X=5.105 $Y=1.35 $X2=0 $Y2=0
cc_296 A4 N_A3_c_388_n 0.00215794f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_297 N_A4_c_334_n N_A3_c_388_n 0.0106756f $X=5.09 $Y=1.557 $X2=0 $Y2=0
cc_298 N_A4_c_332_n N_A3_M1013_g 0.0226172f $X=5.105 $Y=1.35 $X2=0 $Y2=0
cc_299 N_A4_c_336_n N_A3_c_395_n 0.0415254f $X=5.09 $Y=1.765 $X2=0 $Y2=0
cc_300 A4 N_A3_c_395_n 3.36673e-19 $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_301 N_A4_c_331_n N_A3_c_390_n 9.14655e-19 $X=4.675 $Y=1.35 $X2=0 $Y2=0
cc_302 N_A4_c_335_n N_VPWR_c_603_n 0.00291649f $X=4.63 $Y=1.765 $X2=0 $Y2=0
cc_303 N_A4_c_336_n N_VPWR_c_603_n 0.00291649f $X=5.09 $Y=1.765 $X2=0 $Y2=0
cc_304 N_A4_c_335_n N_VPWR_c_589_n 0.00359695f $X=4.63 $Y=1.765 $X2=0 $Y2=0
cc_305 N_A4_c_336_n N_VPWR_c_589_n 0.00359695f $X=5.09 $Y=1.765 $X2=0 $Y2=0
cc_306 N_A4_c_335_n N_A_762_368#_c_773_n 0.0107391f $X=4.63 $Y=1.765 $X2=0 $Y2=0
cc_307 N_A4_c_336_n N_A_762_368#_c_773_n 0.0122705f $X=5.09 $Y=1.765 $X2=0 $Y2=0
cc_308 A4 N_A_762_368#_c_773_n 0.00424992f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_309 N_A4_c_335_n N_A_851_368#_c_821_n 0.0132213f $X=4.63 $Y=1.765 $X2=0 $Y2=0
cc_310 N_A4_c_336_n N_A_851_368#_c_821_n 0.0132213f $X=5.09 $Y=1.765 $X2=0 $Y2=0
cc_311 N_A4_c_331_n N_VGND_c_863_n 0.00291089f $X=4.675 $Y=1.35 $X2=0 $Y2=0
cc_312 N_A4_c_331_n N_VGND_c_864_n 4.43476e-19 $X=4.675 $Y=1.35 $X2=0 $Y2=0
cc_313 N_A4_c_332_n N_VGND_c_864_n 0.0075897f $X=5.105 $Y=1.35 $X2=0 $Y2=0
cc_314 N_A4_c_331_n N_VGND_c_877_n 9.33152e-19 $X=4.675 $Y=1.35 $X2=0 $Y2=0
cc_315 N_A4_c_332_n N_VGND_c_877_n 7.83848e-19 $X=5.105 $Y=1.35 $X2=0 $Y2=0
cc_316 N_A4_c_331_n N_A_523_124#_c_984_n 0.0121471f $X=4.675 $Y=1.35 $X2=0 $Y2=0
cc_317 A4 N_A_523_124#_c_984_n 0.0209304f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_318 N_A4_c_334_n N_A_523_124#_c_984_n 0.00241504f $X=5.09 $Y=1.557 $X2=0
+ $Y2=0
cc_319 N_A4_c_331_n N_A_523_124#_c_986_n 0.0112487f $X=4.675 $Y=1.35 $X2=0 $Y2=0
cc_320 N_A4_c_332_n N_A_523_124#_c_987_n 0.0121744f $X=5.105 $Y=1.35 $X2=0 $Y2=0
cc_321 A4 N_A_523_124#_c_987_n 0.0148952f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_322 N_A4_c_331_n N_A_523_124#_c_992_n 9.00612e-19 $X=4.675 $Y=1.35 $X2=0
+ $Y2=0
cc_323 A4 N_A_523_124#_c_992_n 0.0210654f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_324 N_A4_c_334_n N_A_523_124#_c_992_n 0.00254664f $X=5.09 $Y=1.557 $X2=0
+ $Y2=0
cc_325 N_A3_M1013_g N_A2_M1005_g 0.0120828f $X=5.535 $Y=0.92 $X2=0 $Y2=0
cc_326 N_A3_c_387_n N_A2_c_519_n 0.00774643f $X=5.54 $Y=1.405 $X2=0 $Y2=0
cc_327 N_A3_c_388_n N_A2_c_520_n 0.00774643f $X=5.54 $Y=1.675 $X2=0 $Y2=0
cc_328 N_A3_c_395_n N_A2_c_528_n 0.0184213f $X=5.54 $Y=1.765 $X2=0 $Y2=0
cc_329 N_A3_c_386_n N_A2_c_522_n 0.0120828f $X=5.46 $Y=0.185 $X2=0 $Y2=0
cc_330 N_A3_c_393_n N_VPWR_c_593_n 0.00345084f $X=4.18 $Y=1.765 $X2=0 $Y2=0
cc_331 N_A3_c_393_n N_VPWR_c_603_n 0.00444483f $X=4.18 $Y=1.765 $X2=0 $Y2=0
cc_332 N_A3_c_395_n N_VPWR_c_603_n 0.00444483f $X=5.54 $Y=1.765 $X2=0 $Y2=0
cc_333 N_A3_c_393_n N_VPWR_c_589_n 0.00859578f $X=4.18 $Y=1.765 $X2=0 $Y2=0
cc_334 N_A3_c_395_n N_VPWR_c_589_n 0.0085486f $X=5.54 $Y=1.765 $X2=0 $Y2=0
cc_335 N_A3_c_393_n N_A_762_368#_c_773_n 0.0123929f $X=4.18 $Y=1.765 $X2=0 $Y2=0
cc_336 N_A3_c_395_n N_A_762_368#_c_773_n 0.0169436f $X=5.54 $Y=1.765 $X2=0 $Y2=0
cc_337 N_A3_c_395_n N_A_762_368#_c_767_n 0.0046598f $X=5.54 $Y=1.765 $X2=0 $Y2=0
cc_338 N_A3_c_395_n N_A_762_368#_c_783_n 0.00337571f $X=5.54 $Y=1.765 $X2=0
+ $Y2=0
cc_339 N_A3_c_393_n N_A_762_368#_c_770_n 0.00520662f $X=4.18 $Y=1.765 $X2=0
+ $Y2=0
cc_340 N_A3_c_395_n N_A_762_368#_c_771_n 0.0046144f $X=5.54 $Y=1.765 $X2=0 $Y2=0
cc_341 N_A3_c_393_n N_A_851_368#_c_821_n 0.00432389f $X=4.18 $Y=1.765 $X2=0
+ $Y2=0
cc_342 N_A3_c_395_n N_A_851_368#_c_821_n 0.00411781f $X=5.54 $Y=1.765 $X2=0
+ $Y2=0
cc_343 N_A3_c_391_n N_VGND_M1002_s 0.00269695f $X=4.04 $Y=0.345 $X2=0 $Y2=0
cc_344 N_A3_M1002_g N_VGND_c_863_n 0.00247081f $X=3.925 $Y=0.94 $X2=0 $Y2=0
cc_345 N_A3_c_386_n N_VGND_c_863_n 0.0160258f $X=5.46 $Y=0.185 $X2=0 $Y2=0
cc_346 N_A3_c_390_n N_VGND_c_863_n 0.0050871f $X=4.027 $Y=0.185 $X2=0 $Y2=0
cc_347 N_A3_c_391_n N_VGND_c_863_n 0.0316618f $X=4.04 $Y=0.345 $X2=0 $Y2=0
cc_348 N_A3_c_386_n N_VGND_c_864_n 0.02003f $X=5.46 $Y=0.185 $X2=0 $Y2=0
cc_349 N_A3_M1013_g N_VGND_c_864_n 0.0151923f $X=5.535 $Y=0.92 $X2=0 $Y2=0
cc_350 N_A3_c_386_n N_VGND_c_865_n 0.00157927f $X=5.46 $Y=0.185 $X2=0 $Y2=0
cc_351 N_A3_c_390_n N_VGND_c_868_n 0.0147334f $X=4.027 $Y=0.185 $X2=0 $Y2=0
cc_352 N_A3_c_391_n N_VGND_c_868_n 0.0215843f $X=4.04 $Y=0.345 $X2=0 $Y2=0
cc_353 N_A3_c_386_n N_VGND_c_870_n 0.0185349f $X=5.46 $Y=0.185 $X2=0 $Y2=0
cc_354 N_A3_c_386_n N_VGND_c_872_n 0.0048178f $X=5.46 $Y=0.185 $X2=0 $Y2=0
cc_355 N_A3_c_386_n N_VGND_c_877_n 0.0382998f $X=5.46 $Y=0.185 $X2=0 $Y2=0
cc_356 N_A3_c_390_n N_VGND_c_877_n 0.0117598f $X=4.027 $Y=0.185 $X2=0 $Y2=0
cc_357 N_A3_c_391_n N_VGND_c_877_n 0.0110944f $X=4.04 $Y=0.345 $X2=0 $Y2=0
cc_358 N_A3_c_390_n N_A_523_124#_c_981_n 0.0041408f $X=4.027 $Y=0.185 $X2=0
+ $Y2=0
cc_359 N_A3_c_391_n N_A_523_124#_c_981_n 0.0143361f $X=4.04 $Y=0.345 $X2=0 $Y2=0
cc_360 N_A3_c_390_n N_A_523_124#_c_983_n 0.0100067f $X=4.027 $Y=0.185 $X2=0
+ $Y2=0
cc_361 N_A3_c_391_n N_A_523_124#_c_983_n 0.0184329f $X=4.04 $Y=0.345 $X2=0 $Y2=0
cc_362 N_A3_M1002_g N_A_523_124#_c_984_n 0.0139445f $X=3.925 $Y=0.94 $X2=0 $Y2=0
cc_363 N_A3_c_384_n N_A_523_124#_c_984_n 0.0082136f $X=4.18 $Y=1.485 $X2=0 $Y2=0
cc_364 N_A3_c_390_n N_A_523_124#_c_984_n 7.57014e-19 $X=4.027 $Y=0.185 $X2=0
+ $Y2=0
cc_365 N_A3_c_391_n N_A_523_124#_c_984_n 0.0103418f $X=4.04 $Y=0.345 $X2=0 $Y2=0
cc_366 N_A3_M1002_g N_A_523_124#_c_985_n 3.89157e-19 $X=3.925 $Y=0.94 $X2=0
+ $Y2=0
cc_367 N_A3_c_386_n N_A_523_124#_c_986_n 0.00461056f $X=5.46 $Y=0.185 $X2=0
+ $Y2=0
cc_368 N_A3_c_387_n N_A_523_124#_c_987_n 0.00133459f $X=5.54 $Y=1.405 $X2=0
+ $Y2=0
cc_369 N_A3_M1013_g N_A_523_124#_c_987_n 0.0169534f $X=5.535 $Y=0.92 $X2=0 $Y2=0
cc_370 N_A1_c_465_n N_A2_M1005_g 0.0218812f $X=6.405 $Y=1.35 $X2=0 $Y2=0
cc_371 N_A1_c_465_n N_A2_c_519_n 0.00952883f $X=6.405 $Y=1.35 $X2=0 $Y2=0
cc_372 A1 N_A2_c_520_n 0.00167387f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_373 N_A1_c_468_n N_A2_c_520_n 0.00952883f $X=6.835 $Y=1.557 $X2=0 $Y2=0
cc_374 N_A1_c_469_n N_A2_c_528_n 0.0267621f $X=6.44 $Y=1.765 $X2=0 $Y2=0
cc_375 A1 N_A2_c_528_n 0.00247778f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_376 N_A1_c_468_n N_A2_c_528_n 0.00372657f $X=6.835 $Y=1.557 $X2=0 $Y2=0
cc_377 N_A1_c_465_n N_A2_c_521_n 0.0103098f $X=6.405 $Y=1.35 $X2=0 $Y2=0
cc_378 N_A1_c_466_n N_A2_c_521_n 0.024217f $X=6.835 $Y=1.35 $X2=0 $Y2=0
cc_379 N_A1_c_468_n N_A2_M1020_g 0.0138985f $X=6.835 $Y=1.557 $X2=0 $Y2=0
cc_380 A1 N_A2_c_524_n 0.00720243f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_381 N_A1_c_468_n N_A2_c_524_n 0.00939735f $X=6.835 $Y=1.557 $X2=0 $Y2=0
cc_382 N_A1_c_470_n N_A2_c_530_n 0.0319533f $X=6.93 $Y=1.765 $X2=0 $Y2=0
cc_383 A1 N_A2_c_530_n 3.44124e-19 $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_384 A1 N_A2_c_525_n 0.00166919f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_385 N_A1_c_469_n N_VPWR_c_594_n 0.00420441f $X=6.44 $Y=1.765 $X2=0 $Y2=0
cc_386 N_A1_c_470_n N_VPWR_c_594_n 0.00712781f $X=6.93 $Y=1.765 $X2=0 $Y2=0
cc_387 N_A1_c_469_n N_VPWR_c_603_n 0.00445602f $X=6.44 $Y=1.765 $X2=0 $Y2=0
cc_388 N_A1_c_470_n N_VPWR_c_605_n 0.00413917f $X=6.93 $Y=1.765 $X2=0 $Y2=0
cc_389 N_A1_c_469_n N_VPWR_c_589_n 0.00858046f $X=6.44 $Y=1.765 $X2=0 $Y2=0
cc_390 N_A1_c_470_n N_VPWR_c_589_n 0.00818241f $X=6.93 $Y=1.765 $X2=0 $Y2=0
cc_391 N_A1_c_469_n N_A_762_368#_c_786_n 0.0109024f $X=6.44 $Y=1.765 $X2=0 $Y2=0
cc_392 N_A1_c_470_n N_A_762_368#_c_786_n 0.0111666f $X=6.93 $Y=1.765 $X2=0 $Y2=0
cc_393 A1 N_A_762_368#_c_786_n 0.0490272f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_394 N_A1_c_468_n N_A_762_368#_c_786_n 0.00152389f $X=6.835 $Y=1.557 $X2=0
+ $Y2=0
cc_395 N_A1_c_469_n N_A_1213_368#_c_837_n 0.0120175f $X=6.44 $Y=1.765 $X2=0
+ $Y2=0
cc_396 N_A1_c_470_n N_A_1213_368#_c_837_n 0.0151166f $X=6.93 $Y=1.765 $X2=0
+ $Y2=0
cc_397 N_A1_c_469_n N_A_1213_368#_c_835_n 0.00776934f $X=6.44 $Y=1.765 $X2=0
+ $Y2=0
cc_398 N_A1_c_470_n N_A_1213_368#_c_835_n 6.13664e-19 $X=6.93 $Y=1.765 $X2=0
+ $Y2=0
cc_399 N_A1_c_470_n N_A_1213_368#_c_836_n 0.00283124f $X=6.93 $Y=1.765 $X2=0
+ $Y2=0
cc_400 N_A1_c_465_n N_VGND_c_865_n 0.00159705f $X=6.405 $Y=1.35 $X2=0 $Y2=0
cc_401 N_A1_c_465_n N_VGND_c_867_n 4.43355e-19 $X=6.405 $Y=1.35 $X2=0 $Y2=0
cc_402 N_A1_c_466_n N_VGND_c_867_n 0.00739822f $X=6.835 $Y=1.35 $X2=0 $Y2=0
cc_403 N_A1_c_465_n N_VGND_c_877_n 9.33152e-19 $X=6.405 $Y=1.35 $X2=0 $Y2=0
cc_404 N_A1_c_466_n N_VGND_c_877_n 7.83848e-19 $X=6.835 $Y=1.35 $X2=0 $Y2=0
cc_405 N_A1_c_465_n N_A_523_124#_c_989_n 0.0108924f $X=6.405 $Y=1.35 $X2=0 $Y2=0
cc_406 A1 N_A_523_124#_c_989_n 0.00895556f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_407 N_A1_c_465_n N_A_523_124#_c_990_n 0.00706136f $X=6.405 $Y=1.35 $X2=0
+ $Y2=0
cc_408 N_A1_c_466_n N_A_523_124#_c_991_n 0.0126082f $X=6.835 $Y=1.35 $X2=0 $Y2=0
cc_409 A1 N_A_523_124#_c_991_n 0.0279976f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_410 N_A1_c_468_n N_A_523_124#_c_991_n 5.80271e-19 $X=6.835 $Y=1.557 $X2=0
+ $Y2=0
cc_411 N_A1_c_466_n N_A_523_124#_c_1042_n 7.33515e-19 $X=6.835 $Y=1.35 $X2=0
+ $Y2=0
cc_412 N_A1_c_465_n N_A_523_124#_c_994_n 8.4031e-19 $X=6.405 $Y=1.35 $X2=0 $Y2=0
cc_413 A1 N_A_523_124#_c_994_n 0.0210731f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_414 N_A1_c_468_n N_A_523_124#_c_994_n 0.00253047f $X=6.835 $Y=1.557 $X2=0
+ $Y2=0
cc_415 N_A2_c_530_n N_VPWR_c_594_n 6.07762e-19 $X=7.43 $Y=1.765 $X2=0 $Y2=0
cc_416 N_A2_c_528_n N_VPWR_c_603_n 0.00445602f $X=5.99 $Y=1.765 $X2=0 $Y2=0
cc_417 N_A2_c_530_n N_VPWR_c_605_n 0.00445602f $X=7.43 $Y=1.765 $X2=0 $Y2=0
cc_418 N_A2_c_528_n N_VPWR_c_589_n 0.00858519f $X=5.99 $Y=1.765 $X2=0 $Y2=0
cc_419 N_A2_c_530_n N_VPWR_c_589_n 0.00862902f $X=7.43 $Y=1.765 $X2=0 $Y2=0
cc_420 N_A2_c_528_n N_A_762_368#_c_767_n 0.00262483f $X=5.99 $Y=1.765 $X2=0
+ $Y2=0
cc_421 N_A2_c_528_n N_A_762_368#_c_783_n 0.00337571f $X=5.99 $Y=1.765 $X2=0
+ $Y2=0
cc_422 N_A2_c_528_n N_A_762_368#_c_786_n 0.0171311f $X=5.99 $Y=1.765 $X2=0 $Y2=0
cc_423 N_A2_c_530_n N_A_762_368#_c_786_n 0.0187422f $X=7.43 $Y=1.765 $X2=0 $Y2=0
cc_424 N_A2_c_525_n N_A_762_368#_c_786_n 0.00189086f $X=7.39 $Y=1.48 $X2=0 $Y2=0
cc_425 N_A2_c_530_n N_A_762_368#_c_768_n 0.00299433f $X=7.43 $Y=1.765 $X2=0
+ $Y2=0
cc_426 N_A2_c_530_n N_A_762_368#_c_769_n 0.0169047f $X=7.43 $Y=1.765 $X2=0 $Y2=0
cc_427 N_A2_c_528_n N_A_762_368#_c_771_n 0.00183424f $X=5.99 $Y=1.765 $X2=0
+ $Y2=0
cc_428 N_A2_c_528_n N_A_1213_368#_c_835_n 0.00753224f $X=5.99 $Y=1.765 $X2=0
+ $Y2=0
cc_429 N_A2_c_530_n N_A_1213_368#_c_836_n 0.00743158f $X=7.43 $Y=1.765 $X2=0
+ $Y2=0
cc_430 N_A2_c_522_n N_VGND_c_864_n 0.00158425f $X=6.05 $Y=0.185 $X2=0 $Y2=0
cc_431 N_A2_M1005_g N_VGND_c_865_n 0.0145213f $X=5.975 $Y=0.92 $X2=0 $Y2=0
cc_432 N_A2_c_521_n N_VGND_c_865_n 0.0134054f $X=7.26 $Y=0.185 $X2=0 $Y2=0
cc_433 N_A2_c_522_n N_VGND_c_865_n 0.0024927f $X=6.05 $Y=0.185 $X2=0 $Y2=0
cc_434 N_A2_c_521_n N_VGND_c_866_n 0.0185349f $X=7.26 $Y=0.185 $X2=0 $Y2=0
cc_435 N_A2_c_521_n N_VGND_c_867_n 0.029736f $X=7.26 $Y=0.185 $X2=0 $Y2=0
cc_436 A2 N_VGND_c_867_n 0.0250425f $X=7.835 $Y=0.47 $X2=0 $Y2=0
cc_437 N_A2_c_522_n N_VGND_c_872_n 0.0048178f $X=6.05 $Y=0.185 $X2=0 $Y2=0
cc_438 N_A2_c_521_n N_VGND_c_876_n 0.0138662f $X=7.26 $Y=0.185 $X2=0 $Y2=0
cc_439 A2 N_VGND_c_876_n 0.0386817f $X=7.835 $Y=0.47 $X2=0 $Y2=0
cc_440 N_A2_c_521_n N_VGND_c_877_n 0.0400235f $X=7.26 $Y=0.185 $X2=0 $Y2=0
cc_441 N_A2_c_522_n N_VGND_c_877_n 0.00839621f $X=6.05 $Y=0.185 $X2=0 $Y2=0
cc_442 A2 N_VGND_c_877_n 0.0254788f $X=7.835 $Y=0.47 $X2=0 $Y2=0
cc_443 N_A2_M1005_g N_A_523_124#_c_989_n 0.0168696f $X=5.975 $Y=0.92 $X2=0 $Y2=0
cc_444 N_A2_c_519_n N_A_523_124#_c_989_n 0.00135482f $X=5.99 $Y=1.405 $X2=0
+ $Y2=0
cc_445 N_A2_M1005_g N_A_523_124#_c_990_n 5.60436e-19 $X=5.975 $Y=0.92 $X2=0
+ $Y2=0
cc_446 N_A2_c_521_n N_A_523_124#_c_990_n 0.00460834f $X=7.26 $Y=0.185 $X2=0
+ $Y2=0
cc_447 N_A2_M1020_g N_A_523_124#_c_991_n 0.017037f $X=7.335 $Y=0.935 $X2=0 $Y2=0
cc_448 N_A2_c_525_n N_A_523_124#_c_991_n 0.00471067f $X=7.39 $Y=1.48 $X2=0 $Y2=0
cc_449 A2 N_A_523_124#_c_991_n 0.00203938f $X=7.835 $Y=0.47 $X2=0 $Y2=0
cc_450 N_A2_c_521_n N_A_523_124#_c_1042_n 0.00157463f $X=7.26 $Y=0.185 $X2=0
+ $Y2=0
cc_451 N_A2_M1020_g N_A_523_124#_c_1042_n 0.0083412f $X=7.335 $Y=0.935 $X2=0
+ $Y2=0
cc_452 A2 N_A_523_124#_c_1042_n 0.0166591f $X=7.835 $Y=0.47 $X2=0 $Y2=0
cc_453 N_VPWR_M1000_s N_X_c_692_n 0.00508692f $X=0.465 $Y=1.84 $X2=0 $Y2=0
cc_454 N_VPWR_c_590_n N_X_c_692_n 0.0136682f $X=0.61 $Y=2.275 $X2=0 $Y2=0
cc_455 N_VPWR_c_590_n N_X_c_693_n 0.0566964f $X=0.61 $Y=2.275 $X2=0 $Y2=0
cc_456 N_VPWR_c_591_n N_X_c_693_n 0.0566964f $X=1.51 $Y=2.275 $X2=0 $Y2=0
cc_457 N_VPWR_c_597_n N_X_c_693_n 0.014552f $X=1.425 $Y=3.33 $X2=0 $Y2=0
cc_458 N_VPWR_c_589_n N_X_c_693_n 0.0119791f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_459 N_VPWR_M1004_s N_X_c_694_n 0.00247267f $X=1.36 $Y=1.84 $X2=0 $Y2=0
cc_460 N_VPWR_c_591_n N_X_c_694_n 0.0136682f $X=1.51 $Y=2.275 $X2=0 $Y2=0
cc_461 N_VPWR_c_592_n N_X_c_694_n 0.00213573f $X=2.41 $Y=2.075 $X2=0 $Y2=0
cc_462 N_VPWR_c_591_n N_X_c_695_n 0.0566964f $X=1.51 $Y=2.275 $X2=0 $Y2=0
cc_463 N_VPWR_c_592_n N_X_c_695_n 0.0697297f $X=2.41 $Y=2.075 $X2=0 $Y2=0
cc_464 N_VPWR_c_599_n N_X_c_695_n 0.014552f $X=2.325 $Y=3.33 $X2=0 $Y2=0
cc_465 N_VPWR_c_589_n N_X_c_695_n 0.0119791f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_466 N_VPWR_c_590_n X 0.0590727f $X=0.61 $Y=2.275 $X2=0 $Y2=0
cc_467 N_VPWR_c_595_n X 0.00745548f $X=0.525 $Y=3.33 $X2=0 $Y2=0
cc_468 N_VPWR_c_589_n X 0.00794958f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_469 N_VPWR_M1008_s N_A_762_368#_c_786_n 0.00437233f $X=6.515 $Y=1.84 $X2=0
+ $Y2=0
cc_470 N_VPWR_c_605_n N_A_762_368#_c_769_n 0.0146357f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_471 N_VPWR_c_589_n N_A_762_368#_c_769_n 0.0121141f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_472 N_VPWR_c_593_n N_A_762_368#_c_770_n 0.0455074f $X=3.395 $Y=2.54 $X2=0
+ $Y2=0
cc_473 N_VPWR_c_603_n N_A_762_368#_c_770_n 0.0110778f $X=6.58 $Y=3.33 $X2=0
+ $Y2=0
cc_474 N_VPWR_c_589_n N_A_762_368#_c_770_n 0.00916405f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_475 N_VPWR_c_603_n N_A_762_368#_c_771_n 0.00749631f $X=6.58 $Y=3.33 $X2=0
+ $Y2=0
cc_476 N_VPWR_c_589_n N_A_762_368#_c_771_n 0.0062048f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_477 N_VPWR_c_603_n N_A_851_368#_c_821_n 0.0516441f $X=6.58 $Y=3.33 $X2=0
+ $Y2=0
cc_478 N_VPWR_c_589_n N_A_851_368#_c_821_n 0.0431992f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_479 N_VPWR_M1008_s N_A_1213_368#_c_837_n 0.00496928f $X=6.515 $Y=1.84 $X2=0
+ $Y2=0
cc_480 N_VPWR_c_594_n N_A_1213_368#_c_837_n 0.0171845f $X=6.685 $Y=2.815 $X2=0
+ $Y2=0
cc_481 N_VPWR_c_594_n N_A_1213_368#_c_835_n 0.0224097f $X=6.685 $Y=2.815 $X2=0
+ $Y2=0
cc_482 N_VPWR_c_603_n N_A_1213_368#_c_835_n 0.0145674f $X=6.58 $Y=3.33 $X2=0
+ $Y2=0
cc_483 N_VPWR_c_589_n N_A_1213_368#_c_835_n 0.0119851f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_484 N_VPWR_c_594_n N_A_1213_368#_c_836_n 0.0129302f $X=6.685 $Y=2.815 $X2=0
+ $Y2=0
cc_485 N_VPWR_c_605_n N_A_1213_368#_c_836_n 0.0146094f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_486 N_VPWR_c_589_n N_A_1213_368#_c_836_n 0.0120527f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_487 N_X_c_702_n N_VGND_M1006_s 0.00672868f $X=0.675 $Y=1.015 $X2=-0.19
+ $Y2=-0.245
cc_488 N_X_c_688_n N_VGND_M1006_s 0.00204758f $X=0.295 $Y=1.015 $X2=-0.19
+ $Y2=-0.245
cc_489 N_X_c_712_n N_VGND_M1012_s 0.00463478f $X=1.605 $Y=1.015 $X2=0 $Y2=0
cc_490 N_X_c_702_n N_VGND_c_860_n 0.0160725f $X=0.675 $Y=1.015 $X2=0 $Y2=0
cc_491 N_X_c_688_n N_VGND_c_860_n 0.0107964f $X=0.295 $Y=1.015 $X2=0 $Y2=0
cc_492 N_X_c_689_n N_VGND_c_860_n 0.0155339f $X=0.84 $Y=0.515 $X2=0 $Y2=0
cc_493 N_X_c_689_n N_VGND_c_861_n 0.0154229f $X=0.84 $Y=0.515 $X2=0 $Y2=0
cc_494 N_X_c_712_n N_VGND_c_861_n 0.0210288f $X=1.605 $Y=1.015 $X2=0 $Y2=0
cc_495 N_X_c_690_n N_VGND_c_861_n 0.0155339f $X=1.77 $Y=0.515 $X2=0 $Y2=0
cc_496 N_X_c_690_n N_VGND_c_862_n 0.0215159f $X=1.77 $Y=0.515 $X2=0 $Y2=0
cc_497 N_X_c_689_n N_VGND_c_874_n 0.0109942f $X=0.84 $Y=0.515 $X2=0 $Y2=0
cc_498 N_X_c_690_n N_VGND_c_875_n 0.0109942f $X=1.77 $Y=0.515 $X2=0 $Y2=0
cc_499 N_X_c_689_n N_VGND_c_877_n 0.00904371f $X=0.84 $Y=0.515 $X2=0 $Y2=0
cc_500 N_X_c_690_n N_VGND_c_877_n 0.00904371f $X=1.77 $Y=0.515 $X2=0 $Y2=0
cc_501 N_A_762_368#_c_773_n N_A_851_368#_M1015_s 0.00396407f $X=5.68 $Y=2.375
+ $X2=-0.19 $Y2=1.66
cc_502 N_A_762_368#_c_773_n N_A_851_368#_M1025_d 0.00907897f $X=5.68 $Y=2.375
+ $X2=0 $Y2=0
cc_503 N_A_762_368#_c_773_n N_A_851_368#_c_821_n 0.0671352f $X=5.68 $Y=2.375
+ $X2=0 $Y2=0
cc_504 N_A_762_368#_c_770_n N_A_851_368#_c_821_n 0.0248024f $X=3.955 $Y=2.455
+ $X2=0 $Y2=0
cc_505 N_A_762_368#_c_771_n N_A_851_368#_c_821_n 0.0241317f $X=5.765 $Y=2.4
+ $X2=0 $Y2=0
cc_506 N_A_762_368#_c_786_n N_A_1213_368#_M1017_s 0.00907415f $X=7.54 $Y=2.035
+ $X2=-0.19 $Y2=1.66
cc_507 N_A_762_368#_c_786_n N_A_1213_368#_M1027_d 0.0102761f $X=7.54 $Y=2.035
+ $X2=0 $Y2=0
cc_508 N_A_762_368#_c_786_n N_A_1213_368#_c_837_n 0.0356986f $X=7.54 $Y=2.035
+ $X2=0 $Y2=0
cc_509 N_A_762_368#_c_786_n N_A_1213_368#_c_835_n 0.0173542f $X=7.54 $Y=2.035
+ $X2=0 $Y2=0
cc_510 N_A_762_368#_c_771_n N_A_1213_368#_c_835_n 0.0469254f $X=5.765 $Y=2.4
+ $X2=0 $Y2=0
cc_511 N_A_762_368#_c_786_n N_A_1213_368#_c_836_n 0.0203253f $X=7.54 $Y=2.035
+ $X2=0 $Y2=0
cc_512 N_A_762_368#_c_769_n N_A_1213_368#_c_836_n 0.0202646f $X=7.705 $Y=2.4
+ $X2=0 $Y2=0
cc_513 N_A_762_368#_c_786_n N_A_523_124#_c_991_n 0.00281217f $X=7.54 $Y=2.035
+ $X2=0 $Y2=0
cc_514 N_A_762_368#_c_768_n N_A_523_124#_c_991_n 0.00391062f $X=7.705 $Y=2.12
+ $X2=0 $Y2=0
cc_515 N_A_762_368#_c_767_n N_A_523_124#_c_993_n 0.00667642f $X=5.765 $Y=2.12
+ $X2=0 $Y2=0
cc_516 N_VGND_c_862_n N_A_523_124#_c_980_n 0.0336756f $X=2.2 $Y=0.515 $X2=0
+ $Y2=0
cc_517 N_VGND_c_868_n N_A_523_124#_c_981_n 0.0504256f $X=4.375 $Y=0 $X2=0 $Y2=0
cc_518 N_VGND_c_877_n N_A_523_124#_c_981_n 0.0295559f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_519 N_VGND_c_862_n N_A_523_124#_c_982_n 0.0121618f $X=2.2 $Y=0.515 $X2=0
+ $Y2=0
cc_520 N_VGND_c_868_n N_A_523_124#_c_982_n 0.0229068f $X=4.375 $Y=0 $X2=0 $Y2=0
cc_521 N_VGND_c_877_n N_A_523_124#_c_982_n 0.0127944f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_522 N_VGND_c_863_n N_A_523_124#_c_983_n 0.00647753f $X=4.46 $Y=0.75 $X2=0
+ $Y2=0
cc_523 N_VGND_M1002_s N_A_523_124#_c_984_n 0.0143195f $X=4 $Y=0.62 $X2=0 $Y2=0
cc_524 N_VGND_c_863_n N_A_523_124#_c_984_n 0.0135869f $X=4.46 $Y=0.75 $X2=0
+ $Y2=0
cc_525 N_VGND_c_863_n N_A_523_124#_c_986_n 0.0121933f $X=4.46 $Y=0.75 $X2=0
+ $Y2=0
cc_526 N_VGND_c_864_n N_A_523_124#_c_986_n 0.0127348f $X=5.32 $Y=0.745 $X2=0
+ $Y2=0
cc_527 N_VGND_c_870_n N_A_523_124#_c_986_n 0.00558557f $X=5.155 $Y=0 $X2=0 $Y2=0
cc_528 N_VGND_c_877_n N_A_523_124#_c_986_n 0.0068223f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_529 N_VGND_M1026_s N_A_523_124#_c_987_n 0.00176461f $X=5.18 $Y=0.6 $X2=0
+ $Y2=0
cc_530 N_VGND_c_864_n N_A_523_124#_c_987_n 0.0170777f $X=5.32 $Y=0.745 $X2=0
+ $Y2=0
cc_531 N_VGND_c_864_n N_A_523_124#_c_988_n 0.0126994f $X=5.32 $Y=0.745 $X2=0
+ $Y2=0
cc_532 N_VGND_c_865_n N_A_523_124#_c_988_n 0.0120275f $X=6.19 $Y=0.745 $X2=0
+ $Y2=0
cc_533 N_VGND_c_872_n N_A_523_124#_c_988_n 0.00405637f $X=6.025 $Y=0 $X2=0 $Y2=0
cc_534 N_VGND_c_877_n N_A_523_124#_c_988_n 0.00562174f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_535 N_VGND_M1005_s N_A_523_124#_c_989_n 0.00176461f $X=6.05 $Y=0.6 $X2=0
+ $Y2=0
cc_536 N_VGND_c_865_n N_A_523_124#_c_989_n 0.0152916f $X=6.19 $Y=0.745 $X2=0
+ $Y2=0
cc_537 N_VGND_c_865_n N_A_523_124#_c_990_n 0.0120629f $X=6.19 $Y=0.745 $X2=0
+ $Y2=0
cc_538 N_VGND_c_866_n N_A_523_124#_c_990_n 0.00558247f $X=6.885 $Y=0 $X2=0 $Y2=0
cc_539 N_VGND_c_867_n N_A_523_124#_c_990_n 0.0120629f $X=7.05 $Y=0.745 $X2=0
+ $Y2=0
cc_540 N_VGND_c_877_n N_A_523_124#_c_990_n 0.00681968f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_541 N_VGND_M1009_s N_A_523_124#_c_991_n 0.00996523f $X=6.91 $Y=0.6 $X2=0
+ $Y2=0
cc_542 N_VGND_c_867_n N_A_523_124#_c_991_n 0.015373f $X=7.05 $Y=0.745 $X2=0
+ $Y2=0
cc_543 N_VGND_c_867_n N_A_523_124#_c_1042_n 0.0130127f $X=7.05 $Y=0.745 $X2=0
+ $Y2=0
