* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__a222oi_2 A1 A2 B1 B2 C1 C2 VGND VNB VPB VPWR Y
M1000 a_137_74# C1 Y VNB nshort w=640000u l=150000u
+  ad=3.584e+11p pd=3.68e+06u as=7.232e+11p ps=7.38e+06u
M1001 a_116_392# B2 a_515_392# VPB phighvt w=1e+06u l=150000u
+  ad=1.29e+12p pd=1.058e+07u as=1.49e+12p ps=1.298e+07u
M1002 a_981_74# A1 Y VNB nshort w=640000u l=150000u
+  ad=4.032e+11p pd=3.82e+06u as=0p ps=0u
M1003 a_116_392# C1 Y VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=9.7e+11p ps=7.94e+06u
M1004 a_515_392# A2 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=6.3e+11p ps=5.26e+06u
M1005 Y A1 a_981_74# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND C2 a_137_74# VNB nshort w=640000u l=150000u
+  ad=1.01862e+12p pd=8.5e+06u as=0p ps=0u
M1007 VGND B2 a_593_74# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=3.584e+11p ps=3.68e+06u
M1008 a_137_74# C2 VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y C1 a_137_74# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 Y C2 a_116_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_515_392# B1 a_116_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR A2 a_515_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_593_74# B2 VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Y C1 a_116_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_116_392# B1 a_515_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_116_392# C2 Y VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_515_392# A1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_593_74# B1 Y VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR A1 a_515_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 Y B1 a_593_74# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_515_392# B2 a_116_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND A2 a_981_74# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_981_74# A2 VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
