* File: sky130_fd_sc_ls__o31ai_1.pex.spice
* Created: Fri Aug 28 13:53:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__O31AI_1%A1 1 3 4 6 7
c19 7 0 1.68631e-19 $X=0.24 $Y=1.295
r20 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.385 $X2=0.27 $Y2=1.385
r21 7 11 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.27 $Y=1.295 $X2=0.27
+ $Y2=1.385
r22 4 10 67.5002 $w=3.63e-07 $l=4.54247e-07 $layer=POLY_cond $X=0.52 $Y=1.765
+ $X2=0.357 $Y2=1.385
r23 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.52 $Y=1.765
+ $X2=0.52 $Y2=2.4
r24 1 10 38.952 $w=3.63e-07 $l=2.23596e-07 $layer=POLY_cond $X=0.495 $Y=1.22
+ $X2=0.357 $Y2=1.385
r25 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.495 $Y=1.22 $X2=0.495
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__O31AI_1%A2 3 5 7 8 9 10 11 18
c37 5 0 1.68631e-19 $X=0.94 $Y=1.765
r38 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.015
+ $Y=1.465 $X2=1.015 $Y2=1.465
r39 10 11 7.6965 $w=5.73e-07 $l=3.7e-07 $layer=LI1_cond $X=0.892 $Y=2.405
+ $X2=0.892 $Y2=2.775
r40 9 10 7.6965 $w=5.73e-07 $l=3.7e-07 $layer=LI1_cond $X=0.892 $Y=2.035
+ $X2=0.892 $Y2=2.405
r41 8 9 7.6965 $w=5.73e-07 $l=3.7e-07 $layer=LI1_cond $X=0.892 $Y=1.665
+ $X2=0.892 $Y2=2.035
r42 8 18 4.16027 $w=5.73e-07 $l=2e-07 $layer=LI1_cond $X=0.892 $Y=1.665
+ $X2=0.892 $Y2=1.465
r43 5 17 61.4066 $w=2.86e-07 $l=3.3541e-07 $layer=POLY_cond $X=0.94 $Y=1.765
+ $X2=1.015 $Y2=1.465
r44 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.94 $Y=1.765
+ $X2=0.94 $Y2=2.4
r45 1 17 38.6549 $w=2.86e-07 $l=2.05122e-07 $layer=POLY_cond $X=0.925 $Y=1.3
+ $X2=1.015 $Y2=1.465
r46 1 3 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.925 $Y=1.3 $X2=0.925
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__O31AI_1%A3 1 3 6 8 12
c34 12 0 1.76087e-19 $X=1.855 $Y=1.515
r35 12 14 5.27737 $w=2.74e-07 $l=3e-08 $layer=POLY_cond $X=1.855 $Y=1.557
+ $X2=1.885 $Y2=1.557
r36 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.855
+ $Y=1.515 $X2=1.855 $Y2=1.515
r37 10 12 60.6898 $w=2.74e-07 $l=3.45e-07 $layer=POLY_cond $X=1.51 $Y=1.557
+ $X2=1.855 $Y2=1.557
r38 8 13 8.1743 $w=4.28e-07 $l=3.05e-07 $layer=LI1_cond $X=2.16 $Y=1.565
+ $X2=1.855 $Y2=1.565
r39 4 14 16.847 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.885 $Y=1.35
+ $X2=1.885 $Y2=1.557
r40 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.885 $Y=1.35
+ $X2=1.885 $Y2=0.74
r41 1 10 16.847 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.51 $Y=1.765
+ $X2=1.51 $Y2=1.557
r42 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.51 $Y=1.765
+ $X2=1.51 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__O31AI_1%B1 3 5 7 8 12
c23 12 0 1.76087e-19 $X=2.61 $Y=1.465
c24 3 0 1.49438e-20 $X=2.335 $Y=0.74
r25 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.61
+ $Y=1.465 $X2=2.61 $Y2=1.465
r26 8 12 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=2.61 $Y=1.665 $X2=2.61
+ $Y2=1.465
r27 5 11 55.538 $w=4.17e-07 $l=3.74299e-07 $layer=POLY_cond $X=2.35 $Y=1.765
+ $X2=2.517 $Y2=1.465
r28 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.35 $Y=1.765
+ $X2=2.35 $Y2=2.4
r29 1 11 39.9337 $w=4.17e-07 $l=2.51305e-07 $layer=POLY_cond $X=2.335 $Y=1.3
+ $X2=2.517 $Y2=1.465
r30 1 3 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.335 $Y=1.3 $X2=2.335
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__O31AI_1%VPWR 1 2 7 9 13 15 19 21 34
r25 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r26 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r27 28 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r28 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r29 25 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r30 24 27 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.72 $Y=3.33
+ $X2=2.16 $Y2=3.33
r31 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r32 22 30 3.99177 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.38 $Y=3.33 $X2=0.19
+ $Y2=3.33
r33 22 24 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.38 $Y=3.33
+ $X2=0.72 $Y2=3.33
r34 21 33 4.67962 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=2.41 $Y=3.33
+ $X2=2.645 $Y2=3.33
r35 21 27 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.41 $Y=3.33
+ $X2=2.16 $Y2=3.33
r36 19 28 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=2.16 $Y2=3.33
r37 19 25 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=0.72 $Y2=3.33
r38 15 18 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=2.575 $Y=2.115
+ $X2=2.575 $Y2=2.815
r39 13 33 3.08656 $w=3.3e-07 $l=1.14782e-07 $layer=LI1_cond $X=2.575 $Y=3.245
+ $X2=2.645 $Y2=3.33
r40 13 18 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.575 $Y=3.245
+ $X2=2.575 $Y2=2.815
r41 9 12 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=0.255 $Y=1.985
+ $X2=0.255 $Y2=2.815
r42 7 30 3.1514 $w=2.5e-07 $l=1.12916e-07 $layer=LI1_cond $X=0.255 $Y=3.245
+ $X2=0.19 $Y2=3.33
r43 7 12 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.255 $Y=3.245
+ $X2=0.255 $Y2=2.815
r44 2 18 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.425
+ $Y=1.84 $X2=2.575 $Y2=2.815
r45 2 15 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=2.425
+ $Y=1.84 $X2=2.575 $Y2=2.115
r46 1 12 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.15
+ $Y=1.84 $X2=0.295 $Y2=2.815
r47 1 9 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.15
+ $Y=1.84 $X2=0.295 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_LS__O31AI_1%Y 1 2 9 10 13 15 16 20 21
r41 20 21 12.1537 $w=8.78e-07 $l=1.65e-07 $layer=LI1_cond $X=1.79 $Y=2.115
+ $X2=1.79 $Y2=1.95
r42 15 16 5.12955 $w=8.78e-07 $l=3.7e-07 $layer=LI1_cond $X=1.79 $Y=2.405
+ $X2=1.79 $Y2=2.775
r43 15 20 4.02045 $w=8.78e-07 $l=2.9e-07 $layer=LI1_cond $X=1.79 $Y=2.405
+ $X2=1.79 $Y2=2.115
r44 11 13 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=2.6 $Y=0.96 $X2=2.6
+ $Y2=0.515
r45 9 11 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.435 $Y=1.045
+ $X2=2.6 $Y2=0.96
r46 9 10 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=2.435 $Y=1.045
+ $X2=1.52 $Y2=1.045
r47 7 10 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.435 $Y=1.13
+ $X2=1.52 $Y2=1.045
r48 7 21 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=1.435 $Y=1.13
+ $X2=1.435 $Y2=1.95
r49 2 16 200 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=3 $X=1.585
+ $Y=1.84 $X2=1.735 $Y2=2.815
r50 2 20 200 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=3 $X=1.585
+ $Y=1.84 $X2=1.735 $Y2=2.115
r51 1 13 91 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_NDIFF $count=2 $X=2.41
+ $Y=0.37 $X2=2.6 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__O31AI_1%VGND 1 2 7 9 11 20 21 29 35
r36 33 35 7.72401 $w=5.33e-07 $l=7.5e-08 $layer=LI1_cond $X=1.68 $Y=0.182
+ $X2=1.755 $Y2=0.182
r37 33 34 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r38 31 33 2.01209 $w=5.33e-07 $l=9e-08 $layer=LI1_cond $X=1.59 $Y=0.182 $X2=1.68
+ $Y2=0.182
r39 27 31 8.71908 $w=5.33e-07 $l=3.9e-07 $layer=LI1_cond $X=1.2 $Y=0.182
+ $X2=1.59 $Y2=0.182
r40 27 29 9.28897 $w=5.33e-07 $l=1.45e-07 $layer=LI1_cond $X=1.2 $Y=0.182
+ $X2=1.055 $Y2=0.182
r41 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r42 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r43 21 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=1.68
+ $Y2=0
r44 20 35 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=2.64 $Y=0 $X2=1.755
+ $Y2=0
r45 20 21 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r46 17 28 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r47 17 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r48 16 29 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=1.055
+ $Y2=0
r49 16 17 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r50 14 24 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.222
+ $Y2=0
r51 14 16 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.72
+ $Y2=0
r52 11 34 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.68
+ $Y2=0
r53 11 28 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.2
+ $Y2=0
r54 7 24 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.222 $Y2=0
r55 7 9 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.28 $Y=0.085 $X2=0.28
+ $Y2=0.515
r56 2 31 91 $w=1.7e-07 $l=5.92495e-07 $layer=licon1_NDIFF $count=2 $X=1 $Y=0.37
+ $X2=1.59 $Y2=0.365
r57 1 9 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__O31AI_1%A_114_74# 1 2 9 12 14 16
c31 9 0 1.49438e-20 $X=1.935 $Y=0.705
r32 16 18 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=2.1 $Y=0.57 $X2=2.1
+ $Y2=0.705
r33 12 14 8.75857 $w=2.48e-07 $l=1.9e-07 $layer=LI1_cond $X=0.75 $Y=0.515
+ $X2=0.75 $Y2=0.705
r34 10 14 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.875 $Y=0.705
+ $X2=0.75 $Y2=0.705
r35 9 18 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.935 $Y=0.705
+ $X2=2.1 $Y2=0.705
r36 9 10 69.1551 $w=1.68e-07 $l=1.06e-06 $layer=LI1_cond $X=1.935 $Y=0.705
+ $X2=0.875 $Y2=0.705
r37 2 16 182 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=1 $X=1.96
+ $Y=0.37 $X2=2.1 $Y2=0.57
r38 1 12 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.515
.ends

