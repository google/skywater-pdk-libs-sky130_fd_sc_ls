* File: sky130_fd_sc_ls__nand3_1.pex.spice
* Created: Fri Aug 28 13:33:18 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__NAND3_1%C 1 3 5 6 8 9 10
r23 10 15 3.42618 $w=3.68e-07 $l=1.1e-07 $layer=LI1_cond $X=0.72 $Y=1.365
+ $X2=0.61 $Y2=1.365
r24 9 15 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=1.365
+ $X2=0.61 $Y2=1.365
r25 6 8 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.7 $Y=1.22 $X2=0.7
+ $Y2=0.74
r26 3 5 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.655 $Y=1.765
+ $X2=0.655 $Y2=2.4
r27 1 3 95.4523 $w=1.98e-07 $l=3.87427e-07 $layer=POLY_cond $X=0.67 $Y=1.385
+ $X2=0.655 $Y2=1.765
r28 1 15 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.61
+ $Y=1.385 $X2=0.61 $Y2=1.385
r29 1 6 43.1139 $w=1.98e-07 $l=1.79374e-07 $layer=POLY_cond $X=0.67 $Y=1.385
+ $X2=0.7 $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_LS__NAND3_1%B 1 3 4 6 7 8 9
c34 1 0 2.55527e-19 $X=1.09 $Y=1.22
r35 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.18
+ $Y=1.385 $X2=1.18 $Y2=1.385
r36 9 15 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=1.18 $Y=1.295 $X2=1.18
+ $Y2=1.385
r37 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.18 $Y=0.925 $X2=1.18
+ $Y2=1.295
r38 7 8 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.18 $Y=0.555 $X2=1.18
+ $Y2=0.925
r39 4 14 77.2841 $w=2.7e-07 $l=4.15812e-07 $layer=POLY_cond $X=1.105 $Y=1.765
+ $X2=1.18 $Y2=1.385
r40 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.105 $Y=1.765
+ $X2=1.105 $Y2=2.4
r41 1 14 38.9026 $w=2.7e-07 $l=2.05122e-07 $layer=POLY_cond $X=1.09 $Y=1.22
+ $X2=1.18 $Y2=1.385
r42 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.09 $Y=1.22 $X2=1.09
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__NAND3_1%A 1 3 4 6 7
c28 7 0 1.11073e-19 $X=1.68 $Y=1.295
r29 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.75
+ $Y=1.385 $X2=1.75 $Y2=1.385
r30 7 11 2.96342 $w=3.48e-07 $l=9e-08 $layer=LI1_cond $X=1.74 $Y=1.295 $X2=1.74
+ $Y2=1.385
r31 4 10 77.2841 $w=2.7e-07 $l=4.15812e-07 $layer=POLY_cond $X=1.675 $Y=1.765
+ $X2=1.75 $Y2=1.385
r32 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.675 $Y=1.765
+ $X2=1.675 $Y2=2.4
r33 1 10 38.9026 $w=2.7e-07 $l=2.05122e-07 $layer=POLY_cond $X=1.66 $Y=1.22
+ $X2=1.75 $Y2=1.385
r34 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.66 $Y=1.22 $X2=1.66
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__NAND3_1%VPWR 1 2 7 9 15 20 21 22 29 30
r29 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r30 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r31 24 33 3.93235 $w=1.7e-07 $l=2.18e-07 $layer=LI1_cond $X=0.435 $Y=3.33
+ $X2=0.217 $Y2=3.33
r32 24 26 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=0.435 $Y=3.33
+ $X2=1.2 $Y2=3.33
r33 22 30 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r34 22 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.24 $Y2=3.33
r35 22 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r36 20 26 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=1.215 $Y=3.33
+ $X2=1.2 $Y2=3.33
r37 20 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.215 $Y=3.33
+ $X2=1.38 $Y2=3.33
r38 19 29 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=1.545 $Y=3.33
+ $X2=2.16 $Y2=3.33
r39 19 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.545 $Y=3.33
+ $X2=1.38 $Y2=3.33
r40 15 18 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.38 $Y=2.145
+ $X2=1.38 $Y2=2.825
r41 13 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.38 $Y=3.245
+ $X2=1.38 $Y2=3.33
r42 13 18 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=1.38 $Y=3.245
+ $X2=1.38 $Y2=2.825
r43 9 12 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=0.31 $Y=1.985
+ $X2=0.31 $Y2=2.815
r44 7 33 3.21082 $w=2.5e-07 $l=1.28662e-07 $layer=LI1_cond $X=0.31 $Y=3.245
+ $X2=0.217 $Y2=3.33
r45 7 12 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.31 $Y=3.245 $X2=0.31
+ $Y2=2.815
r46 2 18 400 $w=1.7e-07 $l=1.08038e-06 $layer=licon1_PDIFF $count=1 $X=1.18
+ $Y=1.84 $X2=1.38 $Y2=2.825
r47 2 15 400 $w=1.7e-07 $l=3.9246e-07 $layer=licon1_PDIFF $count=1 $X=1.18
+ $Y=1.84 $X2=1.38 $Y2=2.145
r48 1 12 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.205
+ $Y=1.84 $X2=0.35 $Y2=2.815
r49 1 9 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.205
+ $Y=1.84 $X2=0.35 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_LS__NAND3_1%Y 1 2 3 10 11 14 18 23 27 29 30 31 32 37
c47 27 0 1.44454e-19 $X=2.17 $Y=0.925
r48 32 45 1.04768 $w=4.38e-07 $l=4e-08 $layer=LI1_cond $X=0.825 $Y=2.775
+ $X2=0.825 $Y2=2.815
r49 31 32 9.691 $w=4.38e-07 $l=3.7e-07 $layer=LI1_cond $X=0.825 $Y=2.405
+ $X2=0.825 $Y2=2.775
r50 30 31 9.691 $w=4.38e-07 $l=3.7e-07 $layer=LI1_cond $X=0.825 $Y=2.035
+ $X2=0.825 $Y2=2.405
r51 30 37 1.30959 $w=4.38e-07 $l=5e-08 $layer=LI1_cond $X=0.825 $Y=2.035
+ $X2=0.825 $Y2=1.985
r52 24 37 2.48823 $w=4.38e-07 $l=9.5e-08 $layer=LI1_cond $X=0.825 $Y=1.89
+ $X2=0.825 $Y2=1.985
r53 23 29 2.7724 $w=3.45e-07 $l=2.13307e-07 $layer=LI1_cond $X=2.17 $Y=1.72
+ $X2=1.995 $Y2=1.805
r54 22 27 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.17 $Y=1.01
+ $X2=2.17 $Y2=0.925
r55 22 23 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=2.17 $Y=1.01
+ $X2=2.17 $Y2=1.72
r56 18 20 19.0913 $w=5.18e-07 $l=8.3e-07 $layer=LI1_cond $X=1.995 $Y=1.985
+ $X2=1.995 $Y2=2.815
r57 16 29 2.7724 $w=3.45e-07 $l=8.5e-08 $layer=LI1_cond $X=1.995 $Y=1.89
+ $X2=1.995 $Y2=1.805
r58 16 18 2.18514 $w=5.18e-07 $l=9.5e-08 $layer=LI1_cond $X=1.995 $Y=1.89
+ $X2=1.995 $Y2=1.985
r59 12 27 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.875 $Y=0.925
+ $X2=2.17 $Y2=0.925
r60 12 14 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=1.875 $Y=0.84
+ $X2=1.875 $Y2=0.515
r61 11 24 8.71846 $w=1.7e-07 $l=2.59037e-07 $layer=LI1_cond $X=1.045 $Y=1.805
+ $X2=0.825 $Y2=1.89
r62 10 29 3.97867 $w=1.7e-07 $l=2.6e-07 $layer=LI1_cond $X=1.735 $Y=1.805
+ $X2=1.995 $Y2=1.805
r63 10 11 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.735 $Y=1.805
+ $X2=1.045 $Y2=1.805
r64 3 20 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.75
+ $Y=1.84 $X2=1.9 $Y2=2.815
r65 3 18 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.75
+ $Y=1.84 $X2=1.9 $Y2=1.985
r66 2 45 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=0.73
+ $Y=1.84 $X2=0.88 $Y2=2.815
r67 2 37 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=0.73
+ $Y=1.84 $X2=0.88 $Y2=1.985
r68 1 14 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.735
+ $Y=0.37 $X2=1.875 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__NAND3_1%VGND 1 6 9 10 11 21 22
r21 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r22 18 21 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.72 $Y=0 $X2=2.16
+ $Y2=0
r23 18 19 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r24 15 19 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r25 14 15 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r26 11 22 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r27 11 19 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r28 9 14 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=0.32 $Y=0 $X2=0.24
+ $Y2=0
r29 9 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.32 $Y=0 $X2=0.485
+ $Y2=0
r30 8 18 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=0.65 $Y=0 $X2=0.72
+ $Y2=0
r31 8 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.65 $Y=0 $X2=0.485
+ $Y2=0
r32 4 10 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.485 $Y=0.085
+ $X2=0.485 $Y2=0
r33 4 6 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.485 $Y=0.085
+ $X2=0.485 $Y2=0.515
r34 1 6 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.34
+ $Y=0.37 $X2=0.485 $Y2=0.515
.ends

