* File: sky130_fd_sc_ls__o32a_1.spice
* Created: Wed Sep  2 11:22:40 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__o32a_1.pex.spice"
.subckt sky130_fd_sc_ls__o32a_1  VNB VPB A1 A2 A3 B2 B1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* B1	B1
* B2	B2
* A3	A3
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1004 N_VGND_M1004_d N_A_83_264#_M1004_g N_X_M1004_s VNB NSHORT L=0.15 W=0.74
+ AD=0.157545 AS=0.2109 PD=1.24406 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75002.6 A=0.111 P=1.78 MULT=1
MM1009 N_A_251_74#_M1009_d N_A1_M1009_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.136255 PD=0.92 PS=1.07594 NRD=0 NRS=13.116 M=1 R=4.26667
+ SA=75000.8 SB=75002.4 A=0.096 P=1.58 MULT=1
MM1001 N_VGND_M1001_d N_A2_M1001_g N_A_251_74#_M1009_d VNB NSHORT L=0.15 W=0.64
+ AD=0.1344 AS=0.0896 PD=1.06 PS=0.92 NRD=13.116 NRS=0 M=1 R=4.26667 SA=75001.2
+ SB=75001.9 A=0.096 P=1.58 MULT=1
MM1005 N_A_251_74#_M1005_d N_A3_M1005_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.64
+ AD=0.112 AS=0.1344 PD=0.99 PS=1.06 NRD=0 NRS=13.116 M=1 R=4.26667 SA=75001.8
+ SB=75001.4 A=0.096 P=1.58 MULT=1
MM1002 N_A_83_264#_M1002_d N_B2_M1002_g N_A_251_74#_M1005_d VNB NSHORT L=0.15
+ W=0.64 AD=0.1424 AS=0.112 PD=1.085 PS=0.99 NRD=14.988 NRS=13.116 M=1 R=4.26667
+ SA=75002.3 SB=75000.9 A=0.096 P=1.58 MULT=1
MM1000 N_A_251_74#_M1000_d N_B1_M1000_g N_A_83_264#_M1002_d VNB NSHORT L=0.15
+ W=0.64 AD=0.2144 AS=0.1424 PD=1.95 PS=1.085 NRD=0 NRS=15.936 M=1 R=4.26667
+ SA=75002.9 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1007 N_VPWR_M1007_d N_A_83_264#_M1007_g N_X_M1007_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.291306 AS=0.3304 PD=1.72226 PS=2.83 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75002.7 A=0.168 P=2.54 MULT=1
MM1010 A_248_368# N_A1_M1010_g N_VPWR_M1007_d VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.260094 PD=1.27 PS=1.53774 NRD=15.7403 NRS=33.9628 M=1 R=6.66667
+ SA=75000.9 SB=75002.3 A=0.15 P=2.3 MULT=1
MM1006 A_332_368# N_A2_M1006_g A_248_368# VPB PHIGHVT L=0.15 W=1 AD=0.195
+ AS=0.135 PD=1.39 PS=1.27 NRD=27.5603 NRS=15.7403 M=1 R=6.66667 SA=75001.3
+ SB=75001.9 A=0.15 P=2.3 MULT=1
MM1011 N_A_83_264#_M1011_d N_A3_M1011_g A_332_368# VPB PHIGHVT L=0.15 W=1
+ AD=0.195 AS=0.195 PD=1.39 PS=1.39 NRD=10.8153 NRS=27.5603 M=1 R=6.66667
+ SA=75001.8 SB=75001.4 A=0.15 P=2.3 MULT=1
MM1003 A_548_368# N_B2_M1003_g N_A_83_264#_M1011_d VPB PHIGHVT L=0.15 W=1
+ AD=0.2225 AS=0.195 PD=1.445 PS=1.39 NRD=32.9778 NRS=10.8153 M=1 R=6.66667
+ SA=75002.4 SB=75000.8 A=0.15 P=2.3 MULT=1
MM1008 N_VPWR_M1008_d N_B1_M1008_g A_548_368# VPB PHIGHVT L=0.15 W=1 AD=0.295
+ AS=0.2225 PD=2.59 PS=1.445 NRD=2.9353 NRS=32.9778 M=1 R=6.66667 SA=75003
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8492 P=12.16
*
.include "sky130_fd_sc_ls__o32a_1.pxi.spice"
*
.ends
*
*
