* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__xnor2_4 A B VGND VNB VPB VPWR Y
X0 VPWR A a_950_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X1 Y a_116_368# a_511_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X2 VPWR a_116_368# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X3 a_950_368# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X4 VGND A a_511_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X5 a_511_74# B VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X6 VPWR B a_116_368# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X7 a_950_368# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X8 VGND A a_511_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X9 a_511_74# B VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X10 a_950_368# B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X11 Y a_116_368# a_511_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X12 a_511_74# A VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X13 VPWR A a_116_368# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X14 a_950_368# B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X15 Y a_116_368# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X16 a_116_368# B a_27_74# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X17 VPWR A a_950_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X18 VGND B a_511_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X19 a_511_74# a_116_368# Y VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X20 a_511_74# A VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X21 a_116_368# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X22 VGND B a_511_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X23 a_116_368# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X24 a_27_74# A VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X25 VGND A a_27_74# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X26 Y B a_950_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X27 a_27_74# B a_116_368# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X28 Y B a_950_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X29 a_511_74# a_116_368# Y VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
.ends
