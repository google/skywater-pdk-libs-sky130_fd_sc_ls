* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
M1000 a_95_306# B1 a_645_120# VNB nshort w=640000u l=150000u
+  ad=3.584e+11p pd=3.68e+06u as=3.89825e+11p ps=3.8e+06u
M1001 a_1064_123# A2 VGND VNB nshort w=640000u l=150000u
+  ad=3.584e+11p pd=3.68e+06u as=1.217e+12p ps=1.055e+07u
M1002 X a_95_306# VGND VNB nshort w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=0p ps=0u
M1003 a_95_306# A1 a_1064_123# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND a_95_306# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR A1 a_555_392# VPB phighvt w=1e+06u l=150000u
+  ad=1.767e+12p pd=1.405e+07u as=1.48e+12p ps=1.296e+07u
M1006 VPWR A2 a_555_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_95_306# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=6.72e+11p pd=5.68e+06u as=0p ps=0u
M1008 VPWR a_95_306# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_95_306# B2 a_555_392# VPB phighvt w=1e+06u l=150000u
+  ad=6e+11p pd=5.2e+06u as=0p ps=0u
M1010 a_95_306# B1 a_555_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_555_392# A1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_555_392# A2 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 X a_95_306# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_555_392# B1 a_95_306# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_555_392# B2 a_95_306# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_1064_123# A1 a_95_306# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 X a_95_306# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_645_120# B1 a_95_306# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR a_95_306# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND a_95_306# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND B2 a_645_120# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND A2 a_1064_123# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_645_120# B2 VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
