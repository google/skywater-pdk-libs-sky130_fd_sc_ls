* File: sky130_fd_sc_ls__decaphetap_2.pxi.spice
* Created: Wed Sep  2 11:00:16 2020
* 
x_PM_SKY130_FD_SC_LS__DECAPHETAP_2%VNB VNB N_VNB_R0_neg
+ PM_SKY130_FD_SC_LS__DECAPHETAP_2%VNB
x_PM_SKY130_FD_SC_LS__DECAPHETAP_2%VGND N_VGND_M1000_g N_VGND_R0_pos
+ N_VGND_c_17_n N_VGND_c_18_n N_VGND_c_19_n VGND N_VGND_c_20_n N_VGND_c_21_n
+ N_VGND_c_22_n PM_SKY130_FD_SC_LS__DECAPHETAP_2%VGND
x_PM_SKY130_FD_SC_LS__DECAPHETAP_2%VPWR N_VPWR_M1000_s N_VPWR_c_29_n VPWR
+ N_VPWR_c_31_n VPWR PM_SKY130_FD_SC_LS__DECAPHETAP_2%VPWR
cc_1 VNB N_VGND_M1000_g 0.0027366f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=2.467
cc_2 VNB N_VGND_R0_pos 0.0364474f $X=-0.19 $Y=-0.245 $X2=0.26 $Y2=0.73
cc_3 VNB N_VGND_c_17_n 0.026285f $X=-0.19 $Y=-0.245 $X2=0.172 $Y2=0.73
cc_4 VNB N_VGND_c_18_n 0.0167787f $X=-0.19 $Y=-0.245 $X2=0.277 $Y2=1.222
cc_5 VNB N_VGND_c_19_n 0.019521f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_6 VNB N_VGND_c_20_n 0.0669607f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=1.465
cc_7 VNB N_VGND_c_21_n 0.0177361f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=0
cc_8 VNB N_VGND_c_22_n 0.103334f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=0
cc_9 VNB VPWR 0.0442671f $X=-0.19 $Y=-0.245 $X2=0.277 $Y2=1.03
cc_10 VPB N_VGND_M1000_g 0.0346968f $X=-0.19 $Y=1.66 $X2=0.48 $Y2=2.467
cc_11 VPB N_VGND_c_19_n 0.00346446f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_12 VPB N_VPWR_c_29_n 0.113436f $X=-0.19 $Y=1.66 $X2=0.277 $Y2=1.222
cc_13 VPB VPWR 0.0423048f $X=-0.19 $Y=1.66 $X2=0.277 $Y2=1.03
cc_14 VPB N_VPWR_c_31_n 0.021794f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_15 N_VGND_M1000_g N_VPWR_c_29_n 0.0434328f $X=0.48 $Y=2.467 $X2=0.367
+ $Y2=0.73
cc_16 N_VGND_c_19_n N_VPWR_c_29_n 0.0320693f $X=0.27 $Y=1.465 $X2=0.367 $Y2=0.73
cc_17 N_VGND_c_20_n N_VPWR_c_29_n 0.00187508f $X=0.48 $Y=1.465 $X2=0.367
+ $Y2=0.73
