* NGSPICE file created from sky130_fd_sc_ls__dfsbp_2.ext - technology: sky130A

.subckt sky130_fd_sc_ls__dfsbp_2 CLK D SET_B VGND VNB VPB VPWR Q Q_N
M1000 a_1501_92# a_1339_74# VGND VNB nshort w=420000u l=150000u
+  ad=1.533e+11p pd=1.57e+06u as=2.28115e+12p ps=1.92e+07u
M1001 VGND a_2221_74# Q VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.072e+11p ps=2.04e+06u
M1002 a_398_74# a_225_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=2.9249e+12p ps=2.399e+07u
M1003 a_595_97# a_398_74# a_27_74# VPB phighvt w=420000u l=150000u
+  ad=1.26e+11p pd=1.44e+06u as=2.478e+11p ps=2.86e+06u
M1004 VPWR a_757_401# a_706_463# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1005 a_757_401# a_595_97# VPWR VPB phighvt w=420000u l=150000u
+  ad=1.533e+11p pd=1.57e+06u as=0p ps=0u
M1006 VGND a_1339_74# a_2221_74# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1007 VPWR a_1339_74# a_1501_92# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=2.544e+11p ps=2.27e+06u
M1008 a_1261_74# a_595_97# VGND VNB nshort w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1009 Q_N a_1339_74# VGND VNB nshort w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1010 VPWR a_1501_92# a_1521_508# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1011 Q a_2221_74# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_706_463# a_225_74# a_595_97# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_1521_508# a_398_74# a_1339_74# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=5.701e+11p ps=4.74e+06u
M1014 a_595_97# a_225_74# a_27_74# VNB nshort w=420000u l=150000u
+  ad=2.226e+11p pd=1.9e+06u as=2.394e+11p ps=2.82e+06u
M1015 a_398_74# a_225_74# VGND VNB nshort w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1016 Q a_2221_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=0p ps=0u
M1017 VPWR D a_27_74# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_1339_74# a_398_74# a_1261_74# VNB nshort w=640000u l=150000u
+  ad=2.314e+11p pd=2.12e+06u as=0p ps=0u
M1019 a_1531_118# a_1501_92# a_1453_118# VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=1.008e+11p ps=1.32e+06u
M1020 VGND a_1339_74# Q_N VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_1339_74# SET_B VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND a_757_401# a_731_97# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1023 VGND SET_B a_1001_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1024 VPWR a_1339_74# Q_N VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.36e+11p ps=2.84e+06u
M1025 VPWR a_2221_74# Q VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_1001_74# a_595_97# a_757_401# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1027 VGND D a_27_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 Q_N a_1339_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPWR CLK a_225_74# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.304e+11p ps=2.83e+06u
M1030 VPWR a_1339_74# a_2221_74# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.95e+11p ps=2.59e+06u
M1031 VGND CLK a_225_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1032 a_1258_341# a_595_97# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=3.99625e+11p pd=3.22e+06u as=0p ps=0u
M1033 a_1339_74# a_225_74# a_1258_341# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_731_97# a_398_74# a_595_97# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_1453_118# a_225_74# a_1339_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 VPWR SET_B a_757_401# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 VGND SET_B a_1531_118# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

