* File: sky130_fd_sc_ls__dlxtn_1.pex.spice
* Created: Fri Aug 28 13:20:16 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__DLXTN_1%D 1 3 5 6 8 9 14
c28 5 0 1.70828e-19 $X=0.51 $Y=1.93
c29 1 0 7.48419e-21 $X=0.495 $Y=1.235
r30 14 15 2.26646 $w=3.19e-07 $l=1.5e-08 $layer=POLY_cond $X=0.495 $Y=1.4
+ $X2=0.51 $Y2=1.4
r31 12 14 33.9969 $w=3.19e-07 $l=2.25e-07 $layer=POLY_cond $X=0.27 $Y=1.4
+ $X2=0.495 $Y2=1.4
r32 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.4 $X2=0.27 $Y2=1.4
r33 9 13 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=0.27 $Y=1.295
+ $X2=0.27 $Y2=1.4
r34 6 8 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.51 $Y=2.02 $X2=0.51
+ $Y2=2.515
r35 5 6 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.51 $Y=1.93 $X2=0.51
+ $Y2=2.02
r36 4 15 16.143 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.51 $Y=1.565
+ $X2=0.51 $Y2=1.4
r37 4 5 141.879 $w=1.8e-07 $l=3.65e-07 $layer=POLY_cond $X=0.51 $Y=1.565
+ $X2=0.51 $Y2=1.93
r38 1 14 20.418 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.235
+ $X2=0.495 $Y2=1.4
r39 1 3 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=0.495 $Y=1.235
+ $X2=0.495 $Y2=0.85
.ends

.subckt PM_SKY130_FD_SC_LS__DLXTN_1%GATE_N 1 3 6 8
c39 8 0 1.70828e-19 $X=1.2 $Y=1.665
r40 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.11
+ $Y=1.665 $X2=1.11 $Y2=1.665
r41 8 12 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=1.2 $Y=1.665 $X2=1.11
+ $Y2=1.665
r42 4 11 38.6072 $w=2.91e-07 $l=1.70895e-07 $layer=POLY_cond $X=1.085 $Y=1.5
+ $X2=1.097 $Y2=1.665
r43 4 6 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.085 $Y=1.5 $X2=1.085
+ $Y2=0.94
r44 1 11 70.0779 $w=2.91e-07 $l=3.96119e-07 $layer=POLY_cond $X=1.01 $Y=2.02
+ $X2=1.097 $Y2=1.665
r45 1 3 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.01 $Y=2.02 $X2=1.01
+ $Y2=2.515
.ends

.subckt PM_SKY130_FD_SC_LS__DLXTN_1%A_217_419# 1 2 7 9 10 12 13 15 17 19 20 22
+ 25 27 31 32 35 38 39 40 42 44 45 50 52 56 57 64
c156 56 0 1.53958e-19 $X=4.175 $Y=1.62
c157 27 0 7.48419e-21 $X=1.485 $Y=1.165
r158 66 68 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=3.805 $Y=1.62
+ $X2=3.985 $Y2=1.62
r159 57 68 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=4.175 $Y=1.62
+ $X2=3.985 $Y2=1.62
r160 56 59 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.175 $Y=1.62
+ $X2=4.175 $Y2=1.785
r161 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.175
+ $Y=1.62 $X2=4.175 $Y2=1.62
r162 53 64 45.7946 $w=5.21e-07 $l=4.95e-07 $layer=POLY_cond $X=1.72 $Y=1.535
+ $X2=2.215 $Y2=1.535
r163 53 60 13.4688 $w=3.3e-07 $l=3.5e-07 $layer=POLY_cond $X=1.72 $Y=1.535
+ $X2=1.72 $Y2=1.185
r164 52 54 8.64761 $w=3.98e-07 $l=1.65e-07 $layer=LI1_cond $X=1.685 $Y=1.605
+ $X2=1.685 $Y2=1.77
r165 52 53 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.72
+ $Y=1.605 $X2=1.72 $Y2=1.605
r166 50 60 45.4639 $w=3.3e-07 $l=2.6e-07 $layer=POLY_cond $X=1.72 $Y=0.925
+ $X2=1.72 $Y2=1.185
r167 49 50 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.72
+ $Y=0.925 $X2=1.72 $Y2=0.925
r168 45 54 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.57 $Y=2.075
+ $X2=1.57 $Y2=1.77
r169 44 46 6.81765 $w=4.98e-07 $l=2.85e-07 $layer=LI1_cond $X=1.405 $Y=2.24
+ $X2=1.405 $Y2=2.525
r170 44 45 9.51712 $w=4.98e-07 $l=1.65e-07 $layer=LI1_cond $X=1.405 $Y=2.24
+ $X2=1.405 $Y2=2.075
r171 42 59 73.0695 $w=1.68e-07 $l=1.12e-06 $layer=LI1_cond $X=4.095 $Y=2.905
+ $X2=4.095 $Y2=1.785
r172 39 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.01 $Y=2.99
+ $X2=4.095 $Y2=2.905
r173 39 40 62.9572 $w=1.68e-07 $l=9.65e-07 $layer=LI1_cond $X=4.01 $Y=2.99
+ $X2=3.045 $Y2=2.99
r174 38 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.96 $Y=2.905
+ $X2=3.045 $Y2=2.99
r175 37 38 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.96 $Y=2.61
+ $X2=2.96 $Y2=2.905
r176 36 46 7.15667 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=1.655 $Y=2.525
+ $X2=1.405 $Y2=2.525
r177 35 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.875 $Y=2.525
+ $X2=2.96 $Y2=2.61
r178 35 36 79.5936 $w=1.68e-07 $l=1.22e-06 $layer=LI1_cond $X=2.875 $Y=2.525
+ $X2=1.655 $Y2=2.525
r179 32 52 1.00839 $w=3.98e-07 $l=3.5e-08 $layer=LI1_cond $X=1.685 $Y=1.57
+ $X2=1.685 $Y2=1.605
r180 31 49 3.24963 $w=4e-07 $l=2.85e-07 $layer=LI1_cond $X=1.685 $Y=1.33
+ $X2=1.685 $Y2=1.045
r181 31 32 6.91466 $w=3.98e-07 $l=2.4e-07 $layer=LI1_cond $X=1.685 $Y=1.33
+ $X2=1.685 $Y2=1.57
r182 27 49 3.6487 $w=3.3e-07 $l=2.52982e-07 $layer=LI1_cond $X=1.485 $Y=1.165
+ $X2=1.685 $Y2=1.045
r183 27 29 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=1.485 $Y=1.165
+ $X2=1.3 $Y2=1.165
r184 23 25 110.245 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=3.59 $Y=1.185
+ $X2=3.805 $Y2=1.185
r185 20 22 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.985 $Y=2.465
+ $X2=3.985 $Y2=2.75
r186 19 20 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.985 $Y=2.375
+ $X2=3.985 $Y2=2.465
r187 18 68 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.985 $Y=1.785
+ $X2=3.985 $Y2=1.62
r188 18 19 229.339 $w=1.8e-07 $l=5.9e-07 $layer=POLY_cond $X=3.985 $Y=1.785
+ $X2=3.985 $Y2=2.375
r189 17 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.805 $Y=1.455
+ $X2=3.805 $Y2=1.62
r190 16 25 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.805 $Y=1.26
+ $X2=3.805 $Y2=1.185
r191 16 17 99.9894 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=3.805 $Y=1.26
+ $X2=3.805 $Y2=1.455
r192 13 23 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.59 $Y=1.11
+ $X2=3.59 $Y2=1.185
r193 13 15 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.59 $Y=1.11
+ $X2=3.59 $Y2=0.715
r194 10 64 12.952 $w=5.21e-07 $l=4.14126e-07 $layer=POLY_cond $X=2.355 $Y=1.185
+ $X2=2.215 $Y2=1.535
r195 10 12 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.355 $Y=1.185
+ $X2=2.355 $Y2=0.74
r196 7 64 32.4506 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=2.215 $Y=1.885
+ $X2=2.215 $Y2=1.535
r197 7 9 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.215 $Y=1.885
+ $X2=2.215 $Y2=2.38
r198 2 44 300 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=2 $X=1.085
+ $Y=2.095 $X2=1.32 $Y2=2.24
r199 1 29 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=1.16
+ $Y=0.57 $X2=1.3 $Y2=1.165
.ends

.subckt PM_SKY130_FD_SC_LS__DLXTN_1%A_27_115# 1 2 7 8 9 11 12 14 16 19 22 23 24
+ 26 27 28 30 36 41
c119 9 0 5.6227e-21 $X=2.85 $Y=1.885
c120 7 0 1.06141e-19 $X=2.85 $Y=1.555
r121 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.805
+ $Y=1.39 $X2=2.805 $Y2=1.39
r122 38 41 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=2.56 $Y=1.39
+ $X2=2.805 $Y2=1.39
r123 32 33 12.4428 $w=4.02e-07 $l=4.1e-07 $layer=LI1_cond $X=0.28 $Y=0.782
+ $X2=0.69 $Y2=0.782
r124 30 38 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.56 $Y=1.225
+ $X2=2.56 $Y2=1.39
r125 29 30 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=2.56 $Y=0.425
+ $X2=2.56 $Y2=1.225
r126 27 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.475 $Y=0.34
+ $X2=2.56 $Y2=0.425
r127 27 28 75.6791 $w=1.68e-07 $l=1.16e-06 $layer=LI1_cond $X=2.475 $Y=0.34
+ $X2=1.315 $Y2=0.34
r128 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.23 $Y=0.425
+ $X2=1.315 $Y2=0.34
r129 25 26 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=1.23 $Y=0.425
+ $X2=1.23 $Y2=0.66
r130 24 33 6.73556 $w=4.02e-07 $l=1.01833e-07 $layer=LI1_cond $X=0.775 $Y=0.745
+ $X2=0.69 $Y2=0.782
r131 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.145 $Y=0.745
+ $X2=1.23 $Y2=0.66
r132 23 24 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.145 $Y=0.745
+ $X2=0.775 $Y2=0.745
r133 22 36 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=1.735
+ $X2=0.69 $Y2=1.82
r134 21 33 5.80874 $w=1.7e-07 $l=2.28e-07 $layer=LI1_cond $X=0.69 $Y=1.01
+ $X2=0.69 $Y2=0.782
r135 21 22 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=0.69 $Y=1.01
+ $X2=0.69 $Y2=1.735
r136 17 36 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=0.285 $Y=1.82
+ $X2=0.69 $Y2=1.82
r137 17 19 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.285 $Y=1.905
+ $X2=0.285 $Y2=2.24
r138 14 16 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.2 $Y=1.11
+ $X2=3.2 $Y2=0.715
r139 13 42 34.9152 $w=2.83e-07 $l=2.75409e-07 $layer=POLY_cond $X=2.97 $Y=1.185
+ $X2=2.805 $Y2=1.39
r140 12 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.125 $Y=1.185
+ $X2=3.2 $Y2=1.11
r141 12 13 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=3.125 $Y=1.185
+ $X2=2.97 $Y2=1.185
r142 9 11 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.85 $Y=1.885
+ $X2=2.85 $Y2=2.46
r143 8 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.85 $Y=1.795 $X2=2.85
+ $Y2=1.885
r144 7 42 34.4625 $w=2.83e-07 $l=1.86145e-07 $layer=POLY_cond $X=2.85 $Y=1.555
+ $X2=2.805 $Y2=1.39
r145 7 8 93.2903 $w=1.8e-07 $l=2.4e-07 $layer=POLY_cond $X=2.85 $Y=1.555
+ $X2=2.85 $Y2=1.795
r146 2 19 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.14
+ $Y=2.095 $X2=0.285 $Y2=2.24
r147 1 32 182 $w=1.7e-07 $l=2.67862e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.28 $Y2=0.78
.ends

.subckt PM_SKY130_FD_SC_LS__DLXTN_1%A_369_392# 1 2 7 9 12 15 17 21 23 24 26 30
+ 32 38
c96 30 0 1.11763e-19 $X=3.345 $Y=1.635
c97 23 0 7.08553e-20 $X=4.19 $Y=0.42
c98 21 0 3.15497e-20 $X=3.485 $Y=0.42
r99 30 33 6.30242 $w=3.18e-07 $l=1.75e-07 $layer=LI1_cond $X=3.34 $Y=1.635
+ $X2=3.34 $Y2=1.81
r100 30 32 8.46025 $w=3.18e-07 $l=1.65e-07 $layer=LI1_cond $X=3.34 $Y=1.635
+ $X2=3.34 $Y2=1.47
r101 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.345
+ $Y=1.635 $X2=3.345 $Y2=1.635
r102 26 28 10.7754 $w=3.34e-07 $l=2.95e-07 $layer=LI1_cond $X=2.065 $Y=1.81
+ $X2=2.065 $Y2=2.105
r103 24 38 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.19 $Y=0.42
+ $X2=4.19 $Y2=0.585
r104 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.19
+ $Y=0.42 $X2=4.19 $Y2=0.42
r105 21 23 24.6204 $w=3.28e-07 $l=7.05e-07 $layer=LI1_cond $X=3.485 $Y=0.42
+ $X2=4.19 $Y2=0.42
r106 19 21 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.4 $Y=0.585
+ $X2=3.485 $Y2=0.42
r107 19 32 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=3.4 $Y=0.585
+ $X2=3.4 $Y2=1.47
r108 18 26 4.69528 $w=1.7e-07 $l=2.4e-07 $layer=LI1_cond $X=2.305 $Y=1.81
+ $X2=2.065 $Y2=1.81
r109 17 33 4.44149 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=3.18 $Y=1.81
+ $X2=3.34 $Y2=1.81
r110 17 18 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=3.18 $Y=1.81
+ $X2=2.305 $Y2=1.81
r111 13 26 3.90348 $w=3.34e-07 $l=1.51658e-07 $layer=LI1_cond $X=2.18 $Y=1.725
+ $X2=2.065 $Y2=1.81
r112 13 15 39.8745 $w=2.48e-07 $l=8.65e-07 $layer=LI1_cond $X=2.18 $Y=1.725
+ $X2=2.18 $Y2=0.86
r113 12 38 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.28 $Y=0.905
+ $X2=4.28 $Y2=0.585
r114 7 31 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=3.27 $Y=1.885
+ $X2=3.345 $Y2=1.635
r115 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.27 $Y=1.885
+ $X2=3.27 $Y2=2.46
r116 2 28 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.845
+ $Y=1.96 $X2=1.99 $Y2=2.105
r117 1 15 182 $w=1.7e-07 $l=5.57808e-07 $layer=licon1_NDIFF $count=1 $X=1.995
+ $Y=0.37 $X2=2.14 $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_LS__DLXTN_1%A_863_441# 1 2 7 9 12 14 16 19 21 22 23 30
+ 34 39 41 42 44 46
c93 39 0 1.48577e-19 $X=5.57 $Y=1.94
c94 12 0 7.08553e-20 $X=4.67 $Y=0.905
c95 7 0 1.53958e-19 $X=4.405 $Y=2.465
r96 44 47 8.64761 $w=3.98e-07 $l=1.65e-07 $layer=LI1_cond $X=5.685 $Y=1.465
+ $X2=5.685 $Y2=1.63
r97 44 46 8.64761 $w=3.98e-07 $l=1.65e-07 $layer=LI1_cond $X=5.685 $Y=1.465
+ $X2=5.685 $Y2=1.3
r98 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.72
+ $Y=1.465 $X2=5.72 $Y2=1.465
r99 42 46 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=5.57 $Y=1.135
+ $X2=5.57 $Y2=1.3
r100 39 41 5.90962 $w=2.8e-07 $l=2.56162e-07 $layer=LI1_cond $X=5.57 $Y=1.94
+ $X2=5.46 $Y2=2.147
r101 39 47 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=5.57 $Y=1.94
+ $X2=5.57 $Y2=1.63
r102 32 42 9.23056 $w=3.73e-07 $l=1.87e-07 $layer=LI1_cond $X=5.467 $Y=0.948
+ $X2=5.467 $Y2=1.135
r103 32 34 10.08 $w=3.73e-07 $l=3.28e-07 $layer=LI1_cond $X=5.467 $Y=0.948
+ $X2=5.467 $Y2=0.62
r104 28 41 5.90962 $w=2.8e-07 $l=2.08e-07 $layer=LI1_cond $X=5.46 $Y=2.355
+ $X2=5.46 $Y2=2.147
r105 28 30 13.5929 $w=3.88e-07 $l=4.6e-07 $layer=LI1_cond $X=5.46 $Y=2.355
+ $X2=5.46 $Y2=2.815
r106 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.51
+ $Y=2.19 $X2=4.51 $Y2=2.19
r107 23 41 0.758147 $w=3.3e-07 $l=2.1543e-07 $layer=LI1_cond $X=5.265 $Y=2.19
+ $X2=5.46 $Y2=2.147
r108 23 25 26.3665 $w=3.28e-07 $l=7.55e-07 $layer=LI1_cond $X=5.265 $Y=2.19
+ $X2=4.51 $Y2=2.19
r109 21 45 70.8188 $w=3.3e-07 $l=4.05e-07 $layer=POLY_cond $X=6.125 $Y=1.465
+ $X2=5.72 $Y2=1.465
r110 21 22 5.03009 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.125 $Y=1.465
+ $X2=6.125 $Y2=1.3
r111 17 22 37.0704 $w=1.5e-07 $l=9.5e-08 $layer=POLY_cond $X=6.22 $Y=1.3
+ $X2=6.125 $Y2=1.3
r112 17 19 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=6.22 $Y=1.3
+ $X2=6.22 $Y2=0.74
r113 14 22 37.0704 $w=1.5e-07 $l=5.08011e-07 $layer=POLY_cond $X=6.215 $Y=1.765
+ $X2=6.125 $Y2=1.3
r114 14 16 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.215 $Y=1.765
+ $X2=6.215 $Y2=2.4
r115 10 26 38.8445 $w=3.55e-07 $l=2.24332e-07 $layer=POLY_cond $X=4.67 $Y=2.025
+ $X2=4.53 $Y2=2.19
r116 10 12 574.298 $w=1.5e-07 $l=1.12e-06 $layer=POLY_cond $X=4.67 $Y=2.025
+ $X2=4.67 $Y2=0.905
r117 7 26 53.7797 $w=3.55e-07 $l=3.31662e-07 $layer=POLY_cond $X=4.405 $Y=2.465
+ $X2=4.53 $Y2=2.19
r118 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.405 $Y=2.465
+ $X2=4.405 $Y2=2.75
r119 2 41 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=5.28
+ $Y=1.96 $X2=5.43 $Y2=2.105
r120 2 30 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=5.28
+ $Y=1.96 $X2=5.43 $Y2=2.815
r121 1 34 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.305
+ $Y=0.475 $X2=5.445 $Y2=0.62
.ends

.subckt PM_SKY130_FD_SC_LS__DLXTN_1%A_669_392# 1 2 8 9 11 14 18 19 23 24 26 27
+ 30 31
c91 19 0 4.76483e-20 $X=3.84 $Y=0.93
c92 9 0 1.48577e-19 $X=5.205 $Y=1.885
r93 30 33 10.7882 $w=5.08e-07 $l=4.6e-07 $layer=LI1_cond $X=3.585 $Y=2.15
+ $X2=3.585 $Y2=2.61
r94 30 31 7.70264 $w=5.08e-07 $l=8.5e-08 $layer=LI1_cond $X=3.585 $Y=2.15
+ $X2=3.585 $Y2=2.065
r95 27 37 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.15 $Y=1.47
+ $X2=5.15 $Y2=1.635
r96 27 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.15 $Y=1.47
+ $X2=5.15 $Y2=1.305
r97 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.15
+ $Y=1.47 $X2=5.15 $Y2=1.47
r98 24 26 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=4.68 $Y=1.47
+ $X2=5.15 $Y2=1.47
r99 23 24 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.595 $Y=1.305
+ $X2=4.68 $Y2=1.47
r100 22 23 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=4.595 $Y=1.055
+ $X2=4.595 $Y2=1.305
r101 19 21 4.60977 $w=2.48e-07 $l=1e-07 $layer=LI1_cond $X=3.84 $Y=0.93 $X2=3.94
+ $Y2=0.93
r102 18 22 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.51 $Y=0.93
+ $X2=4.595 $Y2=1.055
r103 18 21 26.2757 $w=2.48e-07 $l=5.7e-07 $layer=LI1_cond $X=4.51 $Y=0.93
+ $X2=3.94 $Y2=0.93
r104 16 19 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.755 $Y=1.055
+ $X2=3.84 $Y2=0.93
r105 16 31 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=3.755 $Y=1.055
+ $X2=3.755 $Y2=2.065
r106 14 36 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=5.23 $Y=0.795
+ $X2=5.23 $Y2=1.305
r107 9 11 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.205 $Y=1.885
+ $X2=5.205 $Y2=2.46
r108 8 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.205 $Y=1.795
+ $X2=5.205 $Y2=1.885
r109 8 37 62.1936 $w=1.8e-07 $l=1.6e-07 $layer=POLY_cond $X=5.205 $Y=1.795
+ $X2=5.205 $Y2=1.635
r110 2 33 600 $w=1.7e-07 $l=7.60592e-07 $layer=licon1_PDIFF $count=1 $X=3.345
+ $Y=1.96 $X2=3.585 $Y2=2.61
r111 2 30 600 $w=1.7e-07 $l=3.21248e-07 $layer=licon1_PDIFF $count=1 $X=3.345
+ $Y=1.96 $X2=3.585 $Y2=2.15
r112 1 21 182 $w=1.7e-07 $l=6.17373e-07 $layer=licon1_NDIFF $count=1 $X=3.665
+ $Y=0.395 $X2=3.94 $Y2=0.89
.ends

.subckt PM_SKY130_FD_SC_LS__DLXTN_1%VPWR 1 2 3 4 15 19 23 27 32 33 34 36 41 49
+ 59 60 63 66 69
r75 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r76 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r77 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r78 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r79 57 60 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6.48 $Y2=3.33
r80 57 70 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=4.56 $Y2=3.33
r81 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r82 54 69 12.4999 $w=1.7e-07 $l=2.98e-07 $layer=LI1_cond $X=5.065 $Y=3.33
+ $X2=4.767 $Y2=3.33
r83 54 56 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=5.065 $Y=3.33
+ $X2=5.52 $Y2=3.33
r84 53 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r85 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r86 50 66 8.88104 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=2.705 $Y=3.33
+ $X2=2.532 $Y2=3.33
r87 50 52 89.7059 $w=1.68e-07 $l=1.375e-06 $layer=LI1_cond $X=2.705 $Y=3.33
+ $X2=4.08 $Y2=3.33
r88 49 69 12.4999 $w=1.7e-07 $l=2.97e-07 $layer=LI1_cond $X=4.47 $Y=3.33
+ $X2=4.767 $Y2=3.33
r89 49 52 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=4.47 $Y=3.33
+ $X2=4.08 $Y2=3.33
r90 48 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r91 47 48 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r92 45 48 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r93 45 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r94 44 47 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r95 44 45 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r96 42 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.95 $Y=3.33
+ $X2=0.785 $Y2=3.33
r97 42 44 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.95 $Y=3.33 $X2=1.2
+ $Y2=3.33
r98 41 66 8.88104 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=2.36 $Y=3.33
+ $X2=2.532 $Y2=3.33
r99 41 47 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=2.36 $Y=3.33 $X2=2.16
+ $Y2=3.33
r100 39 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r101 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r102 36 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.62 $Y=3.33
+ $X2=0.785 $Y2=3.33
r103 36 38 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=0.62 $Y=3.33
+ $X2=0.24 $Y2=3.33
r104 34 53 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=4.08 $Y2=3.33
r105 34 67 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=2.64 $Y2=3.33
r106 32 56 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.825 $Y=3.33
+ $X2=5.52 $Y2=3.33
r107 32 33 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.825 $Y=3.33
+ $X2=5.95 $Y2=3.33
r108 31 59 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=6.075 $Y=3.33
+ $X2=6.48 $Y2=3.33
r109 31 33 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.075 $Y=3.33
+ $X2=5.95 $Y2=3.33
r110 27 30 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=5.95 $Y=1.985
+ $X2=5.95 $Y2=2.815
r111 25 33 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.95 $Y=3.245
+ $X2=5.95 $Y2=3.33
r112 25 30 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=5.95 $Y=3.245
+ $X2=5.95 $Y2=2.815
r113 21 69 2.50116 $w=5.95e-07 $l=8.5e-08 $layer=LI1_cond $X=4.767 $Y=3.245
+ $X2=4.767 $Y2=3.33
r114 21 23 9.95057 $w=5.93e-07 $l=4.95e-07 $layer=LI1_cond $X=4.767 $Y=3.245
+ $X2=4.767 $Y2=2.75
r115 17 66 1.03204 $w=3.45e-07 $l=8.5e-08 $layer=LI1_cond $X=2.532 $Y=3.245
+ $X2=2.532 $Y2=3.33
r116 17 19 10.0212 $w=3.43e-07 $l=3e-07 $layer=LI1_cond $X=2.532 $Y=3.245
+ $X2=2.532 $Y2=2.945
r117 13 63 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.785 $Y=3.245
+ $X2=0.785 $Y2=3.33
r118 13 15 35.0971 $w=3.28e-07 $l=1.005e-06 $layer=LI1_cond $X=0.785 $Y=3.245
+ $X2=0.785 $Y2=2.24
r119 4 30 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=5.845
+ $Y=1.84 $X2=5.99 $Y2=2.815
r120 4 27 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=5.845
+ $Y=1.84 $X2=5.99 $Y2=1.985
r121 3 23 300 $w=1.7e-07 $l=5.95819e-07 $layer=licon1_PDIFF $count=2 $X=4.48
+ $Y=2.54 $X2=4.98 $Y2=2.75
r122 2 19 600 $w=1.7e-07 $l=1.09846e-06 $layer=licon1_PDIFF $count=1 $X=2.29
+ $Y=1.96 $X2=2.53 $Y2=2.945
r123 1 15 300 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=2.095 $X2=0.785 $Y2=2.24
.ends

.subckt PM_SKY130_FD_SC_LS__DLXTN_1%Q 1 2 7 8 9 10 11 12 13
r14 12 13 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=6.437 $Y=2.405
+ $X2=6.437 $Y2=2.775
r15 11 12 14.4485 $w=3.33e-07 $l=4.2e-07 $layer=LI1_cond $X=6.437 $Y=1.985
+ $X2=6.437 $Y2=2.405
r16 10 11 11.0084 $w=3.33e-07 $l=3.2e-07 $layer=LI1_cond $X=6.437 $Y=1.665
+ $X2=6.437 $Y2=1.985
r17 9 10 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=6.437 $Y=1.295
+ $X2=6.437 $Y2=1.665
r18 8 9 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=6.437 $Y=0.925
+ $X2=6.437 $Y2=1.295
r19 7 8 14.1045 $w=3.33e-07 $l=4.1e-07 $layer=LI1_cond $X=6.437 $Y=0.515
+ $X2=6.437 $Y2=0.925
r20 2 13 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=6.29
+ $Y=1.84 $X2=6.44 $Y2=2.815
r21 2 11 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=6.29
+ $Y=1.84 $X2=6.44 $Y2=1.985
r22 1 7 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=6.295
+ $Y=0.37 $X2=6.435 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__DLXTN_1%VGND 1 2 3 4 15 19 23 29 32 33 34 36 41 53
+ 59 60 63 66 69
r84 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r85 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r86 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r87 60 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r88 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r89 57 69 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.09 $Y=0 $X2=5.965
+ $Y2=0
r90 57 59 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=6.09 $Y=0 $X2=6.48
+ $Y2=0
r91 56 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r92 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r93 53 69 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.84 $Y=0 $X2=5.965
+ $Y2=0
r94 53 55 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=5.84 $Y=0 $X2=5.52
+ $Y2=0
r95 52 56 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.52
+ $Y2=0
r96 51 52 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r97 49 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.145 $Y=0 $X2=2.98
+ $Y2=0
r98 49 51 92.3155 $w=1.68e-07 $l=1.415e-06 $layer=LI1_cond $X=3.145 $Y=0
+ $X2=4.56 $Y2=0
r99 48 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r100 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r101 45 48 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r102 45 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r103 44 47 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r104 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r105 42 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=0.79
+ $Y2=0
r106 42 44 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=1.2
+ $Y2=0
r107 41 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.815 $Y=0 $X2=2.98
+ $Y2=0
r108 41 47 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.815 $Y=0
+ $X2=2.64 $Y2=0
r109 39 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r110 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r111 36 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.625 $Y=0 $X2=0.79
+ $Y2=0
r112 36 38 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.625 $Y=0
+ $X2=0.24 $Y2=0
r113 34 52 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=3.36 $Y=0 $X2=4.56
+ $Y2=0
r114 34 67 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.36 $Y=0
+ $X2=3.12 $Y2=0
r115 32 51 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=4.85 $Y=0 $X2=4.56
+ $Y2=0
r116 32 33 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.85 $Y=0 $X2=4.975
+ $Y2=0
r117 31 55 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=5.1 $Y=0 $X2=5.52
+ $Y2=0
r118 31 33 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.1 $Y=0 $X2=4.975
+ $Y2=0
r119 27 69 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.965 $Y=0.085
+ $X2=5.965 $Y2=0
r120 27 29 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=5.965 $Y=0.085
+ $X2=5.965 $Y2=0.515
r121 23 25 16.1342 $w=2.48e-07 $l=3.5e-07 $layer=LI1_cond $X=4.975 $Y=0.62
+ $X2=4.975 $Y2=0.97
r122 21 33 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.975 $Y=0.085
+ $X2=4.975 $Y2=0
r123 21 23 24.6623 $w=2.48e-07 $l=5.35e-07 $layer=LI1_cond $X=4.975 $Y=0.085
+ $X2=4.975 $Y2=0.62
r124 17 66 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.98 $Y=0.085
+ $X2=2.98 $Y2=0
r125 17 19 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=2.98 $Y=0.085
+ $X2=2.98 $Y2=0.54
r126 13 63 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.79 $Y=0.085
+ $X2=0.79 $Y2=0
r127 13 15 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=0.79 $Y=0.085
+ $X2=0.79 $Y2=0.325
r128 4 29 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=5.86
+ $Y=0.37 $X2=6.005 $Y2=0.515
r129 3 25 182 $w=1.7e-07 $l=3.87137e-07 $layer=licon1_NDIFF $count=1 $X=4.745
+ $Y=0.695 $X2=5.015 $Y2=0.97
r130 3 23 182 $w=1.7e-07 $l=3.05205e-07 $layer=licon1_NDIFF $count=1 $X=4.745
+ $Y=0.695 $X2=5.015 $Y2=0.62
r131 2 19 91 $w=1.7e-07 $l=6.29285e-07 $layer=licon1_NDIFF $count=2 $X=2.43
+ $Y=0.37 $X2=2.98 $Y2=0.54
r132 1 15 182 $w=1.7e-07 $l=3.42783e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.575 $X2=0.79 $Y2=0.325
.ends

