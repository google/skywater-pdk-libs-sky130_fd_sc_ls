* File: sky130_fd_sc_ls__a2bb2o_4.pxi.spice
* Created: Wed Sep  2 10:51:03 2020
* 
x_PM_SKY130_FD_SC_LS__A2BB2O_4%A_162_48# N_A_162_48#_M1015_d N_A_162_48#_M1002_s
+ N_A_162_48#_M1006_d N_A_162_48#_M1001_g N_A_162_48#_c_157_n
+ N_A_162_48#_M1003_g N_A_162_48#_M1010_g N_A_162_48#_c_158_n
+ N_A_162_48#_M1008_g N_A_162_48#_M1011_g N_A_162_48#_c_159_n
+ N_A_162_48#_M1017_g N_A_162_48#_M1019_g N_A_162_48#_c_160_n
+ N_A_162_48#_M1022_g N_A_162_48#_c_230_p N_A_162_48#_c_143_n
+ N_A_162_48#_c_144_n N_A_162_48#_c_145_n N_A_162_48#_c_146_n
+ N_A_162_48#_c_147_n N_A_162_48#_c_148_n N_A_162_48#_c_149_n
+ N_A_162_48#_c_150_n N_A_162_48#_c_151_n N_A_162_48#_c_152_n
+ N_A_162_48#_c_153_n N_A_162_48#_c_154_n N_A_162_48#_c_155_n
+ N_A_162_48#_c_156_n PM_SKY130_FD_SC_LS__A2BB2O_4%A_162_48#
x_PM_SKY130_FD_SC_LS__A2BB2O_4%A1_N N_A1_N_c_305_n N_A1_N_M1018_g N_A1_N_M1013_g
+ A1_N N_A1_N_c_307_n PM_SKY130_FD_SC_LS__A2BB2O_4%A1_N
x_PM_SKY130_FD_SC_LS__A2BB2O_4%A2_N N_A2_N_c_342_n N_A2_N_M1004_g N_A2_N_M1021_g
+ A2_N PM_SKY130_FD_SC_LS__A2BB2O_4%A2_N
x_PM_SKY130_FD_SC_LS__A2BB2O_4%A_586_94# N_A_586_94#_M1013_d N_A_586_94#_M1004_d
+ N_A_586_94#_c_374_n N_A_586_94#_M1015_g N_A_586_94#_c_384_n
+ N_A_586_94#_M1006_g N_A_586_94#_c_376_n N_A_586_94#_c_386_n
+ N_A_586_94#_M1014_g N_A_586_94#_c_377_n N_A_586_94#_c_378_n
+ N_A_586_94#_c_406_n N_A_586_94#_c_379_n N_A_586_94#_c_390_n
+ N_A_586_94#_c_391_n N_A_586_94#_c_392_n N_A_586_94#_c_380_n
+ N_A_586_94#_c_381_n N_A_586_94#_c_382_n PM_SKY130_FD_SC_LS__A2BB2O_4%A_586_94#
x_PM_SKY130_FD_SC_LS__A2BB2O_4%B2 N_B2_c_463_n N_B2_c_470_n N_B2_M1016_g
+ N_B2_M1002_g N_B2_c_465_n N_B2_c_472_n N_B2_M1020_g N_B2_M1012_g B2 B2
+ N_B2_c_468_n PM_SKY130_FD_SC_LS__A2BB2O_4%B2
x_PM_SKY130_FD_SC_LS__A2BB2O_4%B1 N_B1_c_516_n N_B1_M1007_g N_B1_c_523_n
+ N_B1_M1000_g N_B1_c_518_n N_B1_c_525_n N_B1_M1005_g N_B1_M1009_g B1 B1
+ N_B1_c_521_n PM_SKY130_FD_SC_LS__A2BB2O_4%B1
x_PM_SKY130_FD_SC_LS__A2BB2O_4%VPWR N_VPWR_M1003_s N_VPWR_M1008_s N_VPWR_M1022_s
+ N_VPWR_M1016_d N_VPWR_M1000_d N_VPWR_c_565_n N_VPWR_c_566_n N_VPWR_c_567_n
+ N_VPWR_c_568_n N_VPWR_c_569_n N_VPWR_c_570_n N_VPWR_c_571_n N_VPWR_c_572_n
+ N_VPWR_c_573_n VPWR N_VPWR_c_574_n N_VPWR_c_575_n N_VPWR_c_576_n
+ N_VPWR_c_577_n N_VPWR_c_564_n N_VPWR_c_579_n N_VPWR_c_580_n N_VPWR_c_581_n
+ PM_SKY130_FD_SC_LS__A2BB2O_4%VPWR
x_PM_SKY130_FD_SC_LS__A2BB2O_4%X N_X_M1001_s N_X_M1011_s N_X_M1003_d N_X_M1017_d
+ N_X_c_655_n N_X_c_651_n N_X_c_652_n N_X_c_657_n N_X_c_653_n N_X_c_658_n
+ N_X_c_654_n N_X_c_659_n N_X_c_660_n X X PM_SKY130_FD_SC_LS__A2BB2O_4%X
x_PM_SKY130_FD_SC_LS__A2BB2O_4%A_820_392# N_A_820_392#_M1006_s
+ N_A_820_392#_M1014_s N_A_820_392#_M1020_s N_A_820_392#_M1005_s
+ N_A_820_392#_c_721_n N_A_820_392#_c_722_n N_A_820_392#_c_723_n
+ N_A_820_392#_c_724_n N_A_820_392#_c_734_n N_A_820_392#_c_725_n
+ N_A_820_392#_c_726_n N_A_820_392#_c_727_n N_A_820_392#_c_728_n
+ N_A_820_392#_c_729_n N_A_820_392#_c_730_n
+ PM_SKY130_FD_SC_LS__A2BB2O_4%A_820_392#
x_PM_SKY130_FD_SC_LS__A2BB2O_4%VGND N_VGND_M1001_d N_VGND_M1010_d N_VGND_M1019_d
+ N_VGND_M1021_d N_VGND_M1007_s N_VGND_c_786_n N_VGND_c_787_n N_VGND_c_788_n
+ N_VGND_c_789_n N_VGND_c_790_n N_VGND_c_791_n N_VGND_c_792_n N_VGND_c_793_n
+ N_VGND_c_794_n N_VGND_c_795_n N_VGND_c_796_n N_VGND_c_797_n N_VGND_c_798_n
+ N_VGND_c_799_n VGND N_VGND_c_800_n N_VGND_c_801_n N_VGND_c_802_n
+ N_VGND_c_803_n PM_SKY130_FD_SC_LS__A2BB2O_4%VGND
x_PM_SKY130_FD_SC_LS__A2BB2O_4%A_1009_74# N_A_1009_74#_M1002_d
+ N_A_1009_74#_M1012_d N_A_1009_74#_M1009_d N_A_1009_74#_c_881_n
+ N_A_1009_74#_c_882_n N_A_1009_74#_c_883_n N_A_1009_74#_c_884_n
+ N_A_1009_74#_c_885_n PM_SKY130_FD_SC_LS__A2BB2O_4%A_1009_74#
cc_1 VNB N_A_162_48#_M1001_g 0.0237255f $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=0.74
cc_2 VNB N_A_162_48#_M1010_g 0.0203596f $X=-0.19 $Y=-0.245 $X2=1.315 $Y2=0.74
cc_3 VNB N_A_162_48#_M1011_g 0.0209199f $X=-0.19 $Y=-0.245 $X2=1.745 $Y2=0.74
cc_4 VNB N_A_162_48#_M1019_g 0.0229405f $X=-0.19 $Y=-0.245 $X2=2.175 $Y2=0.74
cc_5 VNB N_A_162_48#_c_143_n 0.00750527f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=1.095
cc_6 VNB N_A_162_48#_c_144_n 2.98445e-19 $X=-0.19 $Y=-0.245 $X2=2.73 $Y2=1.01
cc_7 VNB N_A_162_48#_c_145_n 0.0112066f $X=-0.19 $Y=-0.245 $X2=3.36 $Y2=0.34
cc_8 VNB N_A_162_48#_c_146_n 0.00241579f $X=-0.19 $Y=-0.245 $X2=2.815 $Y2=0.34
cc_9 VNB N_A_162_48#_c_147_n 7.35049e-19 $X=-0.19 $Y=-0.245 $X2=3.445 $Y2=1.01
cc_10 VNB N_A_162_48#_c_148_n 0.0132956f $X=-0.19 $Y=-0.245 $X2=4.565 $Y2=1.095
cc_11 VNB N_A_162_48#_c_149_n 0.00142487f $X=-0.19 $Y=-0.245 $X2=3.53 $Y2=1.095
cc_12 VNB N_A_162_48#_c_150_n 0.00278408f $X=-0.19 $Y=-0.245 $X2=4.69 $Y2=0.6
cc_13 VNB N_A_162_48#_c_151_n 0.0046355f $X=-0.19 $Y=-0.245 $X2=4.69 $Y2=1.01
cc_14 VNB N_A_162_48#_c_152_n 0.01106f $X=-0.19 $Y=-0.245 $X2=4.675 $Y2=2.105
cc_15 VNB N_A_162_48#_c_153_n 0.015867f $X=-0.19 $Y=-0.245 $X2=5.6 $Y2=0.515
cc_16 VNB N_A_162_48#_c_154_n 0.00148253f $X=-0.19 $Y=-0.245 $X2=2.3 $Y2=1.095
cc_17 VNB N_A_162_48#_c_155_n 0.110483f $X=-0.19 $Y=-0.245 $X2=2.22 $Y2=1.465
cc_18 VNB N_A_162_48#_c_156_n 0.00325813f $X=-0.19 $Y=-0.245 $X2=4.69 $Y2=1.095
cc_19 VNB N_A1_N_c_305_n 0.0242556f $X=-0.19 $Y=-0.245 $X2=4.51 $Y2=0.37
cc_20 VNB N_A1_N_M1013_g 0.0250245f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A1_N_c_307_n 0.00408011f $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=0.74
cc_22 VNB N_A2_N_c_342_n 0.0325434f $X=-0.19 $Y=-0.245 $X2=4.51 $Y2=0.37
cc_23 VNB N_A2_N_M1021_g 0.0298731f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB A2_N 0.00375198f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_586_94#_c_374_n 0.00596955f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_586_94#_M1015_g 0.0530923f $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=0.74
cc_27 VNB N_A_586_94#_c_376_n 0.00782844f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=2.4
cc_28 VNB N_A_586_94#_c_377_n 0.00111172f $X=-0.19 $Y=-0.245 $X2=1.4 $Y2=1.765
cc_29 VNB N_A_586_94#_c_378_n 0.0100545f $X=-0.19 $Y=-0.245 $X2=1.4 $Y2=2.4
cc_30 VNB N_A_586_94#_c_379_n 0.00576653f $X=-0.19 $Y=-0.245 $X2=1.85 $Y2=2.4
cc_31 VNB N_A_586_94#_c_380_n 0.00337719f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.465
cc_32 VNB N_A_586_94#_c_381_n 0.0217151f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.465
cc_33 VNB N_A_586_94#_c_382_n 0.00170689f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_B2_c_463_n 0.00409125f $X=-0.19 $Y=-0.245 $X2=5.46 $Y2=0.37
cc_35 VNB N_B2_M1002_g 0.0300448f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_B2_c_465_n 0.00309826f $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=0.74
cc_37 VNB N_B2_M1012_g 0.0240386f $X=-0.19 $Y=-0.245 $X2=1.315 $Y2=1.3
cc_38 VNB B2 0.00542577f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_B2_c_468_n 0.0434463f $X=-0.19 $Y=-0.245 $X2=1.85 $Y2=2.4
cc_40 VNB N_B1_c_516_n 0.00375404f $X=-0.19 $Y=-0.245 $X2=5.46 $Y2=0.37
cc_41 VNB N_B1_M1007_g 0.0245899f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_B1_c_518_n 0.00418093f $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=0.74
cc_43 VNB N_B1_M1009_g 0.0330373f $X=-0.19 $Y=-0.245 $X2=1.315 $Y2=1.3
cc_44 VNB B1 0.0210179f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_B1_c_521_n 0.0440977f $X=-0.19 $Y=-0.245 $X2=1.85 $Y2=2.4
cc_46 VNB N_VPWR_c_564_n 0.302998f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=1.532
cc_47 VNB N_X_c_651_n 0.0596433f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=1.765
cc_48 VNB N_X_c_652_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=1.315 $Y2=1.3
cc_49 VNB N_X_c_653_n 0.0046653f $X=-0.19 $Y=-0.245 $X2=1.745 $Y2=0.74
cc_50 VNB N_X_c_654_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=2.175 $Y2=1.3
cc_51 VNB N_VGND_c_786_n 0.0276293f $X=-0.19 $Y=-0.245 $X2=1.315 $Y2=0.74
cc_52 VNB N_VGND_c_787_n 0.00420208f $X=-0.19 $Y=-0.245 $X2=1.4 $Y2=2.4
cc_53 VNB N_VGND_c_788_n 0.00520439f $X=-0.19 $Y=-0.245 $X2=1.745 $Y2=0.74
cc_54 VNB N_VGND_c_789_n 0.0126152f $X=-0.19 $Y=-0.245 $X2=1.85 $Y2=2.4
cc_55 VNB N_VGND_c_790_n 0.0182134f $X=-0.19 $Y=-0.245 $X2=2.3 $Y2=2.4
cc_56 VNB N_VGND_c_791_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=2.3 $Y2=2.4
cc_57 VNB N_VGND_c_792_n 0.0172524f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.465
cc_58 VNB N_VGND_c_793_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.465
cc_59 VNB N_VGND_c_794_n 0.0172524f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_795_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=1.095
cc_61 VNB N_VGND_c_796_n 0.00114005f $X=-0.19 $Y=-0.245 $X2=2.73 $Y2=0.425
cc_62 VNB N_VGND_c_797_n 0.00500927f $X=-0.19 $Y=-0.245 $X2=2.73 $Y2=1.01
cc_63 VNB N_VGND_c_798_n 0.054636f $X=-0.19 $Y=-0.245 $X2=3.445 $Y2=0.425
cc_64 VNB N_VGND_c_799_n 0.00311272f $X=-0.19 $Y=-0.245 $X2=3.445 $Y2=1.01
cc_65 VNB N_VGND_c_800_n 0.0306025f $X=-0.19 $Y=-0.245 $X2=2.3 $Y2=1.095
cc_66 VNB N_VGND_c_801_n 0.0170727f $X=-0.19 $Y=-0.245 $X2=1.85 $Y2=1.532
cc_67 VNB N_VGND_c_802_n 0.418406f $X=-0.19 $Y=-0.245 $X2=2.175 $Y2=1.532
cc_68 VNB N_VGND_c_803_n 0.0129863f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_1009_74#_c_881_n 0.0162311f $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=1.3
cc_70 VNB N_A_1009_74#_c_882_n 0.00178301f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=2.4
cc_71 VNB N_A_1009_74#_c_883_n 0.0161319f $X=-0.19 $Y=-0.245 $X2=1.315 $Y2=0.74
cc_72 VNB N_A_1009_74#_c_884_n 0.0237116f $X=-0.19 $Y=-0.245 $X2=1.4 $Y2=2.4
cc_73 VNB N_A_1009_74#_c_885_n 0.00159638f $X=-0.19 $Y=-0.245 $X2=1.745 $Y2=0.74
cc_74 VPB N_A_162_48#_c_157_n 0.01733f $X=-0.19 $Y=1.66 $X2=0.95 $Y2=1.765
cc_75 VPB N_A_162_48#_c_158_n 0.015247f $X=-0.19 $Y=1.66 $X2=1.4 $Y2=1.765
cc_76 VPB N_A_162_48#_c_159_n 0.0152457f $X=-0.19 $Y=1.66 $X2=1.85 $Y2=1.765
cc_77 VPB N_A_162_48#_c_160_n 0.0163625f $X=-0.19 $Y=1.66 $X2=2.3 $Y2=1.765
cc_78 VPB N_A_162_48#_c_152_n 0.00269712f $X=-0.19 $Y=1.66 $X2=4.675 $Y2=2.105
cc_79 VPB N_A_162_48#_c_155_n 0.026947f $X=-0.19 $Y=1.66 $X2=2.22 $Y2=1.465
cc_80 VPB N_A1_N_c_305_n 0.0268089f $X=-0.19 $Y=1.66 $X2=4.51 $Y2=0.37
cc_81 VPB N_A1_N_c_307_n 0.00317333f $X=-0.19 $Y=1.66 $X2=0.885 $Y2=0.74
cc_82 VPB N_A2_N_c_342_n 0.0343197f $X=-0.19 $Y=1.66 $X2=4.51 $Y2=0.37
cc_83 VPB A2_N 0.00432221f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_84 VPB N_A_586_94#_c_374_n 0.00891792f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_A_586_94#_c_384_n 0.0171384f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_A_586_94#_c_376_n 0.0130408f $X=-0.19 $Y=1.66 $X2=0.95 $Y2=2.4
cc_87 VPB N_A_586_94#_c_386_n 0.0148138f $X=-0.19 $Y=1.66 $X2=1.315 $Y2=0.74
cc_88 VPB N_A_586_94#_c_377_n 0.00890359f $X=-0.19 $Y=1.66 $X2=1.4 $Y2=1.765
cc_89 VPB N_A_586_94#_c_378_n 0.0111436f $X=-0.19 $Y=1.66 $X2=1.4 $Y2=2.4
cc_90 VPB N_A_586_94#_c_379_n 0.00125525f $X=-0.19 $Y=1.66 $X2=1.85 $Y2=2.4
cc_91 VPB N_A_586_94#_c_390_n 0.0199565f $X=-0.19 $Y=1.66 $X2=2.175 $Y2=0.74
cc_92 VPB N_A_586_94#_c_391_n 0.0248332f $X=-0.19 $Y=1.66 $X2=2.3 $Y2=1.765
cc_93 VPB N_A_586_94#_c_392_n 6.41458e-19 $X=-0.19 $Y=1.66 $X2=2.3 $Y2=2.4
cc_94 VPB N_A_586_94#_c_380_n 0.00293673f $X=-0.19 $Y=1.66 $X2=1.2 $Y2=1.465
cc_95 VPB N_A_586_94#_c_381_n 0.0176996f $X=-0.19 $Y=1.66 $X2=1.2 $Y2=1.465
cc_96 VPB N_B2_c_463_n 0.00687122f $X=-0.19 $Y=1.66 $X2=5.46 $Y2=0.37
cc_97 VPB N_B2_c_470_n 0.0209621f $X=-0.19 $Y=1.66 $X2=4.525 $Y2=1.96
cc_98 VPB N_B2_c_465_n 0.00616893f $X=-0.19 $Y=1.66 $X2=0.885 $Y2=0.74
cc_99 VPB N_B2_c_472_n 0.0214822f $X=-0.19 $Y=1.66 $X2=0.885 $Y2=0.74
cc_100 VPB B2 0.00561136f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB N_B1_c_516_n 0.00729992f $X=-0.19 $Y=1.66 $X2=5.46 $Y2=0.37
cc_102 VPB N_B1_c_523_n 0.0214786f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 VPB N_B1_c_518_n 0.00847249f $X=-0.19 $Y=1.66 $X2=0.885 $Y2=0.74
cc_104 VPB N_B1_c_525_n 0.0291968f $X=-0.19 $Y=1.66 $X2=0.885 $Y2=0.74
cc_105 VPB B1 0.0110874f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_VPWR_c_565_n 0.0435331f $X=-0.19 $Y=1.66 $X2=1.315 $Y2=0.74
cc_107 VPB N_VPWR_c_566_n 0.00799266f $X=-0.19 $Y=1.66 $X2=1.4 $Y2=2.4
cc_108 VPB N_VPWR_c_567_n 0.00695663f $X=-0.19 $Y=1.66 $X2=1.745 $Y2=0.74
cc_109 VPB N_VPWR_c_568_n 0.00571271f $X=-0.19 $Y=1.66 $X2=2.175 $Y2=0.74
cc_110 VPB N_VPWR_c_569_n 0.00799266f $X=-0.19 $Y=1.66 $X2=2.3 $Y2=2.4
cc_111 VPB N_VPWR_c_570_n 0.0206041f $X=-0.19 $Y=1.66 $X2=1.2 $Y2=1.465
cc_112 VPB N_VPWR_c_571_n 0.00324402f $X=-0.19 $Y=1.66 $X2=1.2 $Y2=1.465
cc_113 VPB N_VPWR_c_572_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_VPWR_c_573_n 0.00324402f $X=-0.19 $Y=1.66 $X2=2.645 $Y2=1.095
cc_115 VPB N_VPWR_c_574_n 0.0199636f $X=-0.19 $Y=1.66 $X2=2.73 $Y2=1.01
cc_116 VPB N_VPWR_c_575_n 0.0196495f $X=-0.19 $Y=1.66 $X2=4.662 $Y2=1.18
cc_117 VPB N_VPWR_c_576_n 0.0696298f $X=-0.19 $Y=1.66 $X2=4.815 $Y2=0.475
cc_118 VPB N_VPWR_c_577_n 0.0199471f $X=-0.19 $Y=1.66 $X2=0.885 $Y2=1.532
cc_119 VPB N_VPWR_c_564_n 0.129748f $X=-0.19 $Y=1.66 $X2=0.95 $Y2=1.532
cc_120 VPB N_VPWR_c_579_n 0.0047828f $X=-0.19 $Y=1.66 $X2=1.4 $Y2=1.532
cc_121 VPB N_VPWR_c_580_n 0.00691066f $X=-0.19 $Y=1.66 $X2=2.175 $Y2=1.532
cc_122 VPB N_VPWR_c_581_n 0.00460249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_X_c_655_n 3.43452e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_X_c_651_n 0.0296822f $X=-0.19 $Y=1.66 $X2=0.95 $Y2=1.765
cc_125 VPB N_X_c_657_n 0.00257348f $X=-0.19 $Y=1.66 $X2=1.4 $Y2=1.765
cc_126 VPB N_X_c_658_n 0.00362403f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_127 VPB N_X_c_659_n 0.00257348f $X=-0.19 $Y=1.66 $X2=2.3 $Y2=1.765
cc_128 VPB N_X_c_660_n 0.00186136f $X=-0.19 $Y=1.66 $X2=1.2 $Y2=1.465
cc_129 VPB N_A_820_392#_c_721_n 0.00964539f $X=-0.19 $Y=1.66 $X2=0.95 $Y2=2.4
cc_130 VPB N_A_820_392#_c_722_n 0.00479765f $X=-0.19 $Y=1.66 $X2=1.315 $Y2=1.3
cc_131 VPB N_A_820_392#_c_723_n 0.00786769f $X=-0.19 $Y=1.66 $X2=1.315 $Y2=0.74
cc_132 VPB N_A_820_392#_c_724_n 0.00912194f $X=-0.19 $Y=1.66 $X2=1.315 $Y2=0.74
cc_133 VPB N_A_820_392#_c_725_n 0.00424615f $X=-0.19 $Y=1.66 $X2=1.4 $Y2=2.4
cc_134 VPB N_A_820_392#_c_726_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_A_820_392#_c_727_n 0.00310502f $X=-0.19 $Y=1.66 $X2=1.85 $Y2=2.4
cc_136 VPB N_A_820_392#_c_728_n 0.0105814f $X=-0.19 $Y=1.66 $X2=2.175 $Y2=1.3
cc_137 VPB N_A_820_392#_c_729_n 0.0360166f $X=-0.19 $Y=1.66 $X2=2.175 $Y2=0.74
cc_138 VPB N_A_820_392#_c_730_n 0.00419642f $X=-0.19 $Y=1.66 $X2=2.215 $Y2=1.465
cc_139 N_A_162_48#_c_160_n N_A1_N_c_305_n 0.0188843f $X=2.3 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_140 N_A_162_48#_c_143_n N_A1_N_c_305_n 0.0013817f $X=2.645 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_141 N_A_162_48#_c_154_n N_A1_N_c_305_n 3.19362e-19 $X=2.3 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_142 N_A_162_48#_c_155_n N_A1_N_c_305_n 0.0240014f $X=2.22 $Y=1.465 $X2=-0.19
+ $Y2=-0.245
cc_143 N_A_162_48#_M1019_g N_A1_N_M1013_g 0.0130514f $X=2.175 $Y=0.74 $X2=0
+ $Y2=0
cc_144 N_A_162_48#_c_143_n N_A1_N_M1013_g 0.00512257f $X=2.645 $Y=1.095 $X2=0
+ $Y2=0
cc_145 N_A_162_48#_c_144_n N_A1_N_M1013_g 0.0143856f $X=2.73 $Y=1.01 $X2=0 $Y2=0
cc_146 N_A_162_48#_c_145_n N_A1_N_M1013_g 0.00873242f $X=3.36 $Y=0.34 $X2=0
+ $Y2=0
cc_147 N_A_162_48#_c_146_n N_A1_N_M1013_g 0.00182405f $X=2.815 $Y=0.34 $X2=0
+ $Y2=0
cc_148 N_A_162_48#_c_154_n N_A1_N_M1013_g 0.00135656f $X=2.3 $Y=1.095 $X2=0
+ $Y2=0
cc_149 N_A_162_48#_c_155_n N_A1_N_M1013_g 0.00154283f $X=2.22 $Y=1.465 $X2=0
+ $Y2=0
cc_150 N_A_162_48#_c_160_n N_A1_N_c_307_n 3.53413e-19 $X=2.3 $Y=1.765 $X2=0
+ $Y2=0
cc_151 N_A_162_48#_c_143_n N_A1_N_c_307_n 0.0215242f $X=2.645 $Y=1.095 $X2=0
+ $Y2=0
cc_152 N_A_162_48#_c_154_n N_A1_N_c_307_n 0.0209458f $X=2.3 $Y=1.095 $X2=0 $Y2=0
cc_153 N_A_162_48#_c_155_n N_A1_N_c_307_n 0.00492492f $X=2.22 $Y=1.465 $X2=0
+ $Y2=0
cc_154 N_A_162_48#_c_148_n N_A2_N_c_342_n 0.00179145f $X=4.565 $Y=1.095
+ $X2=-0.19 $Y2=-0.245
cc_155 N_A_162_48#_c_149_n N_A2_N_c_342_n 0.00396026f $X=3.53 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_156 N_A_162_48#_c_144_n N_A2_N_M1021_g 6.37674e-19 $X=2.73 $Y=1.01 $X2=0
+ $Y2=0
cc_157 N_A_162_48#_c_145_n N_A2_N_M1021_g 0.0126063f $X=3.36 $Y=0.34 $X2=0 $Y2=0
cc_158 N_A_162_48#_c_147_n N_A2_N_M1021_g 0.0122699f $X=3.445 $Y=1.01 $X2=0
+ $Y2=0
cc_159 N_A_162_48#_c_149_n N_A2_N_M1021_g 0.00420304f $X=3.53 $Y=1.095 $X2=0
+ $Y2=0
cc_160 N_A_162_48#_c_148_n A2_N 0.0121728f $X=4.565 $Y=1.095 $X2=0 $Y2=0
cc_161 N_A_162_48#_c_149_n A2_N 0.0146015f $X=3.53 $Y=1.095 $X2=0 $Y2=0
cc_162 N_A_162_48#_c_148_n N_A_586_94#_c_374_n 0.00521975f $X=4.565 $Y=1.095
+ $X2=0 $Y2=0
cc_163 N_A_162_48#_c_148_n N_A_586_94#_M1015_g 0.0202752f $X=4.565 $Y=1.095
+ $X2=0 $Y2=0
cc_164 N_A_162_48#_c_150_n N_A_586_94#_M1015_g 4.60815e-19 $X=4.69 $Y=0.6 $X2=0
+ $Y2=0
cc_165 N_A_162_48#_c_152_n N_A_586_94#_M1015_g 0.0159753f $X=4.675 $Y=2.105
+ $X2=0 $Y2=0
cc_166 N_A_162_48#_c_152_n N_A_586_94#_c_384_n 0.00116514f $X=4.675 $Y=2.105
+ $X2=0 $Y2=0
cc_167 N_A_162_48#_c_152_n N_A_586_94#_c_376_n 0.0182727f $X=4.675 $Y=2.105
+ $X2=0 $Y2=0
cc_168 N_A_162_48#_c_156_n N_A_586_94#_c_376_n 0.00164342f $X=4.69 $Y=1.095
+ $X2=0 $Y2=0
cc_169 N_A_162_48#_c_152_n N_A_586_94#_c_386_n 0.00451029f $X=4.675 $Y=2.105
+ $X2=0 $Y2=0
cc_170 N_A_162_48#_c_148_n N_A_586_94#_c_377_n 0.00144804f $X=4.565 $Y=1.095
+ $X2=0 $Y2=0
cc_171 N_A_162_48#_c_152_n N_A_586_94#_c_377_n 9.5063e-19 $X=4.675 $Y=2.105
+ $X2=0 $Y2=0
cc_172 N_A_162_48#_c_152_n N_A_586_94#_c_378_n 0.00209897f $X=4.675 $Y=2.105
+ $X2=0 $Y2=0
cc_173 N_A_162_48#_c_145_n N_A_586_94#_c_406_n 0.0142089f $X=3.36 $Y=0.34 $X2=0
+ $Y2=0
cc_174 N_A_162_48#_c_143_n N_A_586_94#_c_379_n 0.00331391f $X=2.645 $Y=1.095
+ $X2=0 $Y2=0
cc_175 N_A_162_48#_c_154_n N_A_586_94#_c_379_n 0.00488541f $X=2.3 $Y=1.095 $X2=0
+ $Y2=0
cc_176 N_A_162_48#_c_152_n N_A_586_94#_c_391_n 0.00414378f $X=4.675 $Y=2.105
+ $X2=0 $Y2=0
cc_177 N_A_162_48#_c_148_n N_A_586_94#_c_380_n 0.0156104f $X=4.565 $Y=1.095
+ $X2=0 $Y2=0
cc_178 N_A_162_48#_c_152_n N_A_586_94#_c_380_n 0.0185334f $X=4.675 $Y=2.105
+ $X2=0 $Y2=0
cc_179 N_A_162_48#_c_148_n N_A_586_94#_c_381_n 0.00303502f $X=4.565 $Y=1.095
+ $X2=0 $Y2=0
cc_180 N_A_162_48#_c_143_n N_A_586_94#_c_382_n 0.00545578f $X=2.645 $Y=1.095
+ $X2=0 $Y2=0
cc_181 N_A_162_48#_c_149_n N_A_586_94#_c_382_n 0.00975088f $X=3.53 $Y=1.095
+ $X2=0 $Y2=0
cc_182 N_A_162_48#_c_152_n N_B2_c_463_n 4.18998e-19 $X=4.675 $Y=2.105 $X2=0
+ $Y2=0
cc_183 N_A_162_48#_c_151_n N_B2_M1002_g 0.00307188f $X=4.69 $Y=1.01 $X2=0 $Y2=0
cc_184 N_A_162_48#_c_152_n N_B2_M1002_g 0.00184906f $X=4.675 $Y=2.105 $X2=0
+ $Y2=0
cc_185 N_A_162_48#_c_153_n N_B2_M1002_g 0.0132302f $X=5.6 $Y=0.515 $X2=0 $Y2=0
cc_186 N_A_162_48#_c_156_n N_B2_M1002_g 0.0029913f $X=4.69 $Y=1.095 $X2=0 $Y2=0
cc_187 N_A_162_48#_c_153_n N_B2_M1012_g 0.00337267f $X=5.6 $Y=0.515 $X2=0 $Y2=0
cc_188 N_A_162_48#_c_152_n B2 0.0145622f $X=4.675 $Y=2.105 $X2=0 $Y2=0
cc_189 N_A_162_48#_c_152_n N_B2_c_468_n 0.00779214f $X=4.675 $Y=2.105 $X2=0
+ $Y2=0
cc_190 N_A_162_48#_c_157_n N_VPWR_c_565_n 0.00993564f $X=0.95 $Y=1.765 $X2=0
+ $Y2=0
cc_191 N_A_162_48#_c_158_n N_VPWR_c_566_n 0.00586501f $X=1.4 $Y=1.765 $X2=0
+ $Y2=0
cc_192 N_A_162_48#_c_159_n N_VPWR_c_566_n 0.00586501f $X=1.85 $Y=1.765 $X2=0
+ $Y2=0
cc_193 N_A_162_48#_c_160_n N_VPWR_c_567_n 0.00932553f $X=2.3 $Y=1.765 $X2=0
+ $Y2=0
cc_194 N_A_162_48#_c_157_n N_VPWR_c_570_n 0.00445602f $X=0.95 $Y=1.765 $X2=0
+ $Y2=0
cc_195 N_A_162_48#_c_158_n N_VPWR_c_570_n 0.00445602f $X=1.4 $Y=1.765 $X2=0
+ $Y2=0
cc_196 N_A_162_48#_c_159_n N_VPWR_c_575_n 0.00445602f $X=1.85 $Y=1.765 $X2=0
+ $Y2=0
cc_197 N_A_162_48#_c_160_n N_VPWR_c_575_n 0.00445602f $X=2.3 $Y=1.765 $X2=0
+ $Y2=0
cc_198 N_A_162_48#_c_157_n N_VPWR_c_564_n 0.00862391f $X=0.95 $Y=1.765 $X2=0
+ $Y2=0
cc_199 N_A_162_48#_c_158_n N_VPWR_c_564_n 0.00857589f $X=1.4 $Y=1.765 $X2=0
+ $Y2=0
cc_200 N_A_162_48#_c_159_n N_VPWR_c_564_n 0.00857589f $X=1.85 $Y=1.765 $X2=0
+ $Y2=0
cc_201 N_A_162_48#_c_160_n N_VPWR_c_564_n 0.00857749f $X=2.3 $Y=1.765 $X2=0
+ $Y2=0
cc_202 N_A_162_48#_c_157_n N_X_c_655_n 0.0149737f $X=0.95 $Y=1.765 $X2=0 $Y2=0
cc_203 N_A_162_48#_c_155_n N_X_c_655_n 0.00133221f $X=2.22 $Y=1.465 $X2=0 $Y2=0
cc_204 N_A_162_48#_M1001_g N_X_c_651_n 0.0223418f $X=0.885 $Y=0.74 $X2=0 $Y2=0
cc_205 N_A_162_48#_M1010_g N_X_c_651_n 5.75161e-19 $X=1.315 $Y=0.74 $X2=0 $Y2=0
cc_206 N_A_162_48#_c_230_p N_X_c_651_n 0.0370738f $X=2.215 $Y=1.465 $X2=0 $Y2=0
cc_207 N_A_162_48#_c_155_n N_X_c_651_n 0.0225486f $X=2.22 $Y=1.465 $X2=0 $Y2=0
cc_208 N_A_162_48#_M1001_g N_X_c_652_n 0.0128625f $X=0.885 $Y=0.74 $X2=0 $Y2=0
cc_209 N_A_162_48#_M1010_g N_X_c_652_n 3.97481e-19 $X=1.315 $Y=0.74 $X2=0 $Y2=0
cc_210 N_A_162_48#_c_157_n N_X_c_657_n 0.017229f $X=0.95 $Y=1.765 $X2=0 $Y2=0
cc_211 N_A_162_48#_c_158_n N_X_c_657_n 0.0125029f $X=1.4 $Y=1.765 $X2=0 $Y2=0
cc_212 N_A_162_48#_c_159_n N_X_c_657_n 6.9119e-19 $X=1.85 $Y=1.765 $X2=0 $Y2=0
cc_213 N_A_162_48#_M1010_g N_X_c_653_n 0.0124434f $X=1.315 $Y=0.74 $X2=0 $Y2=0
cc_214 N_A_162_48#_M1011_g N_X_c_653_n 0.0120709f $X=1.745 $Y=0.74 $X2=0 $Y2=0
cc_215 N_A_162_48#_c_230_p N_X_c_653_n 0.0657213f $X=2.215 $Y=1.465 $X2=0 $Y2=0
cc_216 N_A_162_48#_c_154_n N_X_c_653_n 0.00497192f $X=2.3 $Y=1.095 $X2=0 $Y2=0
cc_217 N_A_162_48#_c_155_n N_X_c_653_n 0.00467196f $X=2.22 $Y=1.465 $X2=0 $Y2=0
cc_218 N_A_162_48#_c_158_n N_X_c_658_n 0.0120074f $X=1.4 $Y=1.765 $X2=0 $Y2=0
cc_219 N_A_162_48#_c_159_n N_X_c_658_n 0.0129464f $X=1.85 $Y=1.765 $X2=0 $Y2=0
cc_220 N_A_162_48#_c_160_n N_X_c_658_n 0.00403157f $X=2.3 $Y=1.765 $X2=0 $Y2=0
cc_221 N_A_162_48#_c_230_p N_X_c_658_n 0.067414f $X=2.215 $Y=1.465 $X2=0 $Y2=0
cc_222 N_A_162_48#_c_154_n N_X_c_658_n 0.00205785f $X=2.3 $Y=1.095 $X2=0 $Y2=0
cc_223 N_A_162_48#_c_155_n N_X_c_658_n 0.0156879f $X=2.22 $Y=1.465 $X2=0 $Y2=0
cc_224 N_A_162_48#_M1010_g N_X_c_654_n 6.20738e-19 $X=1.315 $Y=0.74 $X2=0 $Y2=0
cc_225 N_A_162_48#_M1011_g N_X_c_654_n 0.00866629f $X=1.745 $Y=0.74 $X2=0 $Y2=0
cc_226 N_A_162_48#_M1019_g N_X_c_654_n 3.97481e-19 $X=2.175 $Y=0.74 $X2=0 $Y2=0
cc_227 N_A_162_48#_c_158_n N_X_c_659_n 6.9119e-19 $X=1.4 $Y=1.765 $X2=0 $Y2=0
cc_228 N_A_162_48#_c_159_n N_X_c_659_n 0.0125029f $X=1.85 $Y=1.765 $X2=0 $Y2=0
cc_229 N_A_162_48#_c_160_n N_X_c_659_n 0.0106924f $X=2.3 $Y=1.765 $X2=0 $Y2=0
cc_230 N_A_162_48#_c_157_n N_X_c_660_n 0.00114729f $X=0.95 $Y=1.765 $X2=0 $Y2=0
cc_231 N_A_162_48#_c_158_n N_X_c_660_n 9.27134e-19 $X=1.4 $Y=1.765 $X2=0 $Y2=0
cc_232 N_A_162_48#_c_230_p N_X_c_660_n 0.0256538f $X=2.215 $Y=1.465 $X2=0 $Y2=0
cc_233 N_A_162_48#_c_155_n N_X_c_660_n 0.00800971f $X=2.22 $Y=1.465 $X2=0 $Y2=0
cc_234 N_A_162_48#_M1006_d N_A_820_392#_c_722_n 0.00222494f $X=4.525 $Y=1.96
+ $X2=0 $Y2=0
cc_235 N_A_162_48#_c_152_n N_A_820_392#_c_722_n 0.013472f $X=4.675 $Y=2.105
+ $X2=0 $Y2=0
cc_236 N_A_162_48#_c_152_n N_A_820_392#_c_724_n 0.011904f $X=4.675 $Y=2.105
+ $X2=0 $Y2=0
cc_237 N_A_162_48#_c_152_n N_A_820_392#_c_734_n 0.0395952f $X=4.675 $Y=2.105
+ $X2=0 $Y2=0
cc_238 N_A_162_48#_c_143_n N_VGND_M1019_d 0.00860096f $X=2.645 $Y=1.095 $X2=0
+ $Y2=0
cc_239 N_A_162_48#_c_144_n N_VGND_M1019_d 0.00604133f $X=2.73 $Y=1.01 $X2=0
+ $Y2=0
cc_240 N_A_162_48#_c_154_n N_VGND_M1019_d 0.0011083f $X=2.3 $Y=1.095 $X2=0 $Y2=0
cc_241 N_A_162_48#_c_147_n N_VGND_M1021_d 0.0129017f $X=3.445 $Y=1.01 $X2=0
+ $Y2=0
cc_242 N_A_162_48#_c_148_n N_VGND_M1021_d 0.0164421f $X=4.565 $Y=1.095 $X2=0
+ $Y2=0
cc_243 N_A_162_48#_c_149_n N_VGND_M1021_d 6.25458e-19 $X=3.53 $Y=1.095 $X2=0
+ $Y2=0
cc_244 N_A_162_48#_M1001_g N_VGND_c_786_n 0.00466772f $X=0.885 $Y=0.74 $X2=0
+ $Y2=0
cc_245 N_A_162_48#_M1001_g N_VGND_c_787_n 5.05592e-19 $X=0.885 $Y=0.74 $X2=0
+ $Y2=0
cc_246 N_A_162_48#_M1010_g N_VGND_c_787_n 0.00914496f $X=1.315 $Y=0.74 $X2=0
+ $Y2=0
cc_247 N_A_162_48#_M1011_g N_VGND_c_787_n 0.00183835f $X=1.745 $Y=0.74 $X2=0
+ $Y2=0
cc_248 N_A_162_48#_M1011_g N_VGND_c_788_n 5.20618e-19 $X=1.745 $Y=0.74 $X2=0
+ $Y2=0
cc_249 N_A_162_48#_M1019_g N_VGND_c_788_n 0.0117339f $X=2.175 $Y=0.74 $X2=0
+ $Y2=0
cc_250 N_A_162_48#_c_143_n N_VGND_c_788_n 0.00724091f $X=2.645 $Y=1.095 $X2=0
+ $Y2=0
cc_251 N_A_162_48#_c_144_n N_VGND_c_788_n 0.0310611f $X=2.73 $Y=1.01 $X2=0 $Y2=0
cc_252 N_A_162_48#_c_146_n N_VGND_c_788_n 0.0146659f $X=2.815 $Y=0.34 $X2=0
+ $Y2=0
cc_253 N_A_162_48#_c_154_n N_VGND_c_788_n 0.00887034f $X=2.3 $Y=1.095 $X2=0
+ $Y2=0
cc_254 N_A_162_48#_c_155_n N_VGND_c_788_n 5.01214e-19 $X=2.22 $Y=1.465 $X2=0
+ $Y2=0
cc_255 N_A_162_48#_c_145_n N_VGND_c_789_n 0.0158668f $X=3.36 $Y=0.34 $X2=0 $Y2=0
cc_256 N_A_162_48#_c_147_n N_VGND_c_789_n 0.0337298f $X=3.445 $Y=1.01 $X2=0
+ $Y2=0
cc_257 N_A_162_48#_c_148_n N_VGND_c_789_n 0.0507639f $X=4.565 $Y=1.095 $X2=0
+ $Y2=0
cc_258 N_A_162_48#_c_150_n N_VGND_c_789_n 0.0109137f $X=4.69 $Y=0.6 $X2=0 $Y2=0
cc_259 N_A_162_48#_M1001_g N_VGND_c_792_n 0.00434272f $X=0.885 $Y=0.74 $X2=0
+ $Y2=0
cc_260 N_A_162_48#_M1010_g N_VGND_c_792_n 0.00383152f $X=1.315 $Y=0.74 $X2=0
+ $Y2=0
cc_261 N_A_162_48#_M1011_g N_VGND_c_794_n 0.00434272f $X=1.745 $Y=0.74 $X2=0
+ $Y2=0
cc_262 N_A_162_48#_M1019_g N_VGND_c_794_n 0.00383152f $X=2.175 $Y=0.74 $X2=0
+ $Y2=0
cc_263 N_A_162_48#_c_150_n N_VGND_c_798_n 0.0111552f $X=4.69 $Y=0.6 $X2=0 $Y2=0
cc_264 N_A_162_48#_c_153_n N_VGND_c_798_n 0.0388592f $X=5.6 $Y=0.515 $X2=0 $Y2=0
cc_265 N_A_162_48#_c_145_n N_VGND_c_800_n 0.0472364f $X=3.36 $Y=0.34 $X2=0 $Y2=0
cc_266 N_A_162_48#_c_146_n N_VGND_c_800_n 0.0121867f $X=2.815 $Y=0.34 $X2=0
+ $Y2=0
cc_267 N_A_162_48#_M1001_g N_VGND_c_802_n 0.00825283f $X=0.885 $Y=0.74 $X2=0
+ $Y2=0
cc_268 N_A_162_48#_M1010_g N_VGND_c_802_n 0.0075754f $X=1.315 $Y=0.74 $X2=0
+ $Y2=0
cc_269 N_A_162_48#_M1011_g N_VGND_c_802_n 0.00820284f $X=1.745 $Y=0.74 $X2=0
+ $Y2=0
cc_270 N_A_162_48#_M1019_g N_VGND_c_802_n 0.0075754f $X=2.175 $Y=0.74 $X2=0
+ $Y2=0
cc_271 N_A_162_48#_c_145_n N_VGND_c_802_n 0.027092f $X=3.36 $Y=0.34 $X2=0 $Y2=0
cc_272 N_A_162_48#_c_146_n N_VGND_c_802_n 0.00660921f $X=2.815 $Y=0.34 $X2=0
+ $Y2=0
cc_273 N_A_162_48#_c_150_n N_VGND_c_802_n 0.00923333f $X=4.69 $Y=0.6 $X2=0 $Y2=0
cc_274 N_A_162_48#_c_153_n N_VGND_c_802_n 0.033121f $X=5.6 $Y=0.515 $X2=0 $Y2=0
cc_275 N_A_162_48#_c_153_n N_A_1009_74#_M1002_d 0.00332037f $X=5.6 $Y=0.515
+ $X2=-0.19 $Y2=-0.245
cc_276 N_A_162_48#_M1002_s N_A_1009_74#_c_881_n 0.00176801f $X=5.46 $Y=0.37
+ $X2=0 $Y2=0
cc_277 N_A_162_48#_c_151_n N_A_1009_74#_c_881_n 0.0191245f $X=4.69 $Y=1.01 $X2=0
+ $Y2=0
cc_278 N_A_162_48#_c_153_n N_A_1009_74#_c_881_n 0.0438027f $X=5.6 $Y=0.515 $X2=0
+ $Y2=0
cc_279 N_A_162_48#_c_156_n N_A_1009_74#_c_881_n 0.00683847f $X=4.69 $Y=1.095
+ $X2=0 $Y2=0
cc_280 N_A_162_48#_c_153_n N_A_1009_74#_c_882_n 0.010629f $X=5.6 $Y=0.515 $X2=0
+ $Y2=0
cc_281 N_A1_N_c_305_n N_A2_N_c_342_n 0.0906855f $X=2.84 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_282 N_A1_N_c_307_n N_A2_N_c_342_n 3.74872e-19 $X=2.765 $Y=1.515 $X2=-0.19
+ $Y2=-0.245
cc_283 N_A1_N_M1013_g N_A2_N_M1021_g 0.0234549f $X=2.855 $Y=0.79 $X2=0 $Y2=0
cc_284 N_A1_N_c_305_n N_A_586_94#_c_379_n 0.00381f $X=2.84 $Y=1.765 $X2=0 $Y2=0
cc_285 N_A1_N_M1013_g N_A_586_94#_c_379_n 0.00488927f $X=2.855 $Y=0.79 $X2=0
+ $Y2=0
cc_286 N_A1_N_c_307_n N_A_586_94#_c_379_n 0.0320025f $X=2.765 $Y=1.515 $X2=0
+ $Y2=0
cc_287 N_A1_N_c_305_n N_A_586_94#_c_390_n 0.00240777f $X=2.84 $Y=1.765 $X2=0
+ $Y2=0
cc_288 N_A1_N_c_305_n N_A_586_94#_c_392_n 0.00135719f $X=2.84 $Y=1.765 $X2=0
+ $Y2=0
cc_289 N_A1_N_M1013_g N_A_586_94#_c_382_n 6.65078e-19 $X=2.855 $Y=0.79 $X2=0
+ $Y2=0
cc_290 N_A1_N_c_305_n N_VPWR_c_567_n 0.0207506f $X=2.84 $Y=1.765 $X2=0 $Y2=0
cc_291 N_A1_N_c_307_n N_VPWR_c_567_n 0.0170945f $X=2.765 $Y=1.515 $X2=0 $Y2=0
cc_292 N_A1_N_c_305_n N_VPWR_c_576_n 0.00413917f $X=2.84 $Y=1.765 $X2=0 $Y2=0
cc_293 N_A1_N_c_305_n N_VPWR_c_564_n 0.00817239f $X=2.84 $Y=1.765 $X2=0 $Y2=0
cc_294 N_A1_N_c_305_n N_X_c_658_n 6.06928e-19 $X=2.84 $Y=1.765 $X2=0 $Y2=0
cc_295 N_A1_N_c_305_n N_X_c_659_n 2.19524e-19 $X=2.84 $Y=1.765 $X2=0 $Y2=0
cc_296 N_A1_N_M1013_g N_VGND_c_788_n 0.00145351f $X=2.855 $Y=0.79 $X2=0 $Y2=0
cc_297 N_A1_N_M1013_g N_VGND_c_800_n 7.822e-19 $X=2.855 $Y=0.79 $X2=0 $Y2=0
cc_298 A2_N N_A_586_94#_M1015_g 0.00262375f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_299 N_A2_N_c_342_n N_A_586_94#_c_379_n 0.0158212f $X=3.23 $Y=1.765 $X2=0
+ $Y2=0
cc_300 A2_N N_A_586_94#_c_379_n 0.0310564f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_301 N_A2_N_c_342_n N_A_586_94#_c_390_n 0.0145288f $X=3.23 $Y=1.765 $X2=0
+ $Y2=0
cc_302 N_A2_N_c_342_n N_A_586_94#_c_392_n 0.0159494f $X=3.23 $Y=1.765 $X2=0
+ $Y2=0
cc_303 A2_N N_A_586_94#_c_392_n 0.0259161f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_304 N_A2_N_c_342_n N_A_586_94#_c_380_n 0.00228086f $X=3.23 $Y=1.765 $X2=0
+ $Y2=0
cc_305 A2_N N_A_586_94#_c_380_n 0.0243455f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_306 N_A2_N_c_342_n N_A_586_94#_c_381_n 0.0152883f $X=3.23 $Y=1.765 $X2=0
+ $Y2=0
cc_307 A2_N N_A_586_94#_c_381_n 0.0023924f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_308 N_A2_N_M1021_g N_A_586_94#_c_382_n 0.00532649f $X=3.285 $Y=0.79 $X2=0
+ $Y2=0
cc_309 N_A2_N_c_342_n N_VPWR_c_567_n 0.00310276f $X=3.23 $Y=1.765 $X2=0 $Y2=0
cc_310 N_A2_N_c_342_n N_VPWR_c_576_n 0.00445602f $X=3.23 $Y=1.765 $X2=0 $Y2=0
cc_311 N_A2_N_c_342_n N_VPWR_c_564_n 0.00862666f $X=3.23 $Y=1.765 $X2=0 $Y2=0
cc_312 N_A2_N_M1021_g N_VGND_c_789_n 4.48089e-19 $X=3.285 $Y=0.79 $X2=0 $Y2=0
cc_313 N_A2_N_M1021_g N_VGND_c_800_n 7.82463e-19 $X=3.285 $Y=0.79 $X2=0 $Y2=0
cc_314 N_A_586_94#_c_378_n N_B2_c_463_n 0.0117837f $X=4.9 $Y=1.725 $X2=0 $Y2=0
cc_315 N_A_586_94#_c_386_n N_B2_c_470_n 0.00803334f $X=4.9 $Y=1.885 $X2=0 $Y2=0
cc_316 N_A_586_94#_c_378_n B2 4.93152e-19 $X=4.9 $Y=1.725 $X2=0 $Y2=0
cc_317 N_A_586_94#_c_390_n N_VPWR_c_567_n 0.0265401f $X=3.455 $Y=2.815 $X2=0
+ $Y2=0
cc_318 N_A_586_94#_c_392_n N_VPWR_c_567_n 0.0107239f $X=3.62 $Y=2.035 $X2=0
+ $Y2=0
cc_319 N_A_586_94#_c_386_n N_VPWR_c_568_n 3.75192e-19 $X=4.9 $Y=1.885 $X2=0
+ $Y2=0
cc_320 N_A_586_94#_c_384_n N_VPWR_c_576_n 0.00278257f $X=4.45 $Y=1.885 $X2=0
+ $Y2=0
cc_321 N_A_586_94#_c_386_n N_VPWR_c_576_n 0.00278257f $X=4.9 $Y=1.885 $X2=0
+ $Y2=0
cc_322 N_A_586_94#_c_390_n N_VPWR_c_576_n 0.0145938f $X=3.455 $Y=2.815 $X2=0
+ $Y2=0
cc_323 N_A_586_94#_c_384_n N_VPWR_c_564_n 0.00358623f $X=4.45 $Y=1.885 $X2=0
+ $Y2=0
cc_324 N_A_586_94#_c_386_n N_VPWR_c_564_n 0.00353905f $X=4.9 $Y=1.885 $X2=0
+ $Y2=0
cc_325 N_A_586_94#_c_390_n N_VPWR_c_564_n 0.0120466f $X=3.455 $Y=2.815 $X2=0
+ $Y2=0
cc_326 N_A_586_94#_c_379_n A_583_368# 0.00145764f $X=3.105 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_327 N_A_586_94#_c_392_n A_583_368# 0.00481315f $X=3.62 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_328 N_A_586_94#_c_391_n N_A_820_392#_M1006_s 0.0030054f $X=3.855 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_329 N_A_586_94#_c_384_n N_A_820_392#_c_721_n 0.00789307f $X=4.45 $Y=1.885
+ $X2=0 $Y2=0
cc_330 N_A_586_94#_c_386_n N_A_820_392#_c_721_n 5.5529e-19 $X=4.9 $Y=1.885 $X2=0
+ $Y2=0
cc_331 N_A_586_94#_c_390_n N_A_820_392#_c_721_n 0.0265266f $X=3.455 $Y=2.815
+ $X2=0 $Y2=0
cc_332 N_A_586_94#_c_391_n N_A_820_392#_c_721_n 0.00813517f $X=3.855 $Y=2.035
+ $X2=0 $Y2=0
cc_333 N_A_586_94#_c_381_n N_A_820_392#_c_721_n 0.00578726f $X=3.985 $Y=1.635
+ $X2=0 $Y2=0
cc_334 N_A_586_94#_c_384_n N_A_820_392#_c_722_n 0.0107904f $X=4.45 $Y=1.885
+ $X2=0 $Y2=0
cc_335 N_A_586_94#_c_386_n N_A_820_392#_c_722_n 0.0122595f $X=4.9 $Y=1.885 $X2=0
+ $Y2=0
cc_336 N_A_586_94#_c_384_n N_A_820_392#_c_723_n 0.00262934f $X=4.45 $Y=1.885
+ $X2=0 $Y2=0
cc_337 N_A_586_94#_c_390_n N_A_820_392#_c_723_n 0.00343054f $X=3.455 $Y=2.815
+ $X2=0 $Y2=0
cc_338 N_A_586_94#_c_386_n N_A_820_392#_c_724_n 0.00254934f $X=4.9 $Y=1.885
+ $X2=0 $Y2=0
cc_339 N_A_586_94#_c_378_n N_A_820_392#_c_724_n 7.22069e-19 $X=4.9 $Y=1.725
+ $X2=0 $Y2=0
cc_340 N_A_586_94#_c_384_n N_A_820_392#_c_734_n 6.24717e-19 $X=4.45 $Y=1.885
+ $X2=0 $Y2=0
cc_341 N_A_586_94#_c_386_n N_A_820_392#_c_734_n 0.00919154f $X=4.9 $Y=1.885
+ $X2=0 $Y2=0
cc_342 N_A_586_94#_M1015_g N_VGND_c_789_n 0.016897f $X=4.435 $Y=0.74 $X2=0 $Y2=0
cc_343 N_A_586_94#_M1015_g N_VGND_c_798_n 0.00383152f $X=4.435 $Y=0.74 $X2=0
+ $Y2=0
cc_344 N_A_586_94#_M1015_g N_VGND_c_802_n 0.00762539f $X=4.435 $Y=0.74 $X2=0
+ $Y2=0
cc_345 N_B2_c_465_n N_B1_c_516_n 0.00970055f $X=5.8 $Y=1.795 $X2=0 $Y2=0
cc_346 N_B2_M1012_g N_B1_M1007_g 0.0181154f $X=5.815 $Y=0.69 $X2=0 $Y2=0
cc_347 N_B2_c_472_n N_B1_c_523_n 0.0183067f $X=5.8 $Y=1.885 $X2=0 $Y2=0
cc_348 B2 B1 0.0356352f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_349 N_B2_c_468_n B1 2.24997e-19 $X=5.815 $Y=1.425 $X2=0 $Y2=0
cc_350 B2 N_B1_c_521_n 0.00559665f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_351 N_B2_c_468_n N_B1_c_521_n 0.00970055f $X=5.815 $Y=1.425 $X2=0 $Y2=0
cc_352 N_B2_c_470_n N_VPWR_c_568_n 0.00997879f $X=5.35 $Y=1.885 $X2=0 $Y2=0
cc_353 N_B2_c_472_n N_VPWR_c_568_n 0.00526215f $X=5.8 $Y=1.885 $X2=0 $Y2=0
cc_354 N_B2_c_472_n N_VPWR_c_572_n 0.00445602f $X=5.8 $Y=1.885 $X2=0 $Y2=0
cc_355 N_B2_c_470_n N_VPWR_c_576_n 0.00413917f $X=5.35 $Y=1.885 $X2=0 $Y2=0
cc_356 N_B2_c_470_n N_VPWR_c_564_n 0.0081781f $X=5.35 $Y=1.885 $X2=0 $Y2=0
cc_357 N_B2_c_472_n N_VPWR_c_564_n 0.00857673f $X=5.8 $Y=1.885 $X2=0 $Y2=0
cc_358 N_B2_c_470_n N_A_820_392#_c_722_n 0.00125031f $X=5.35 $Y=1.885 $X2=0
+ $Y2=0
cc_359 N_B2_c_470_n N_A_820_392#_c_725_n 0.0179014f $X=5.35 $Y=1.885 $X2=0 $Y2=0
cc_360 N_B2_c_472_n N_A_820_392#_c_725_n 0.0124546f $X=5.8 $Y=1.885 $X2=0 $Y2=0
cc_361 B2 N_A_820_392#_c_725_n 0.0359957f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_362 N_B2_c_468_n N_A_820_392#_c_725_n 4.03951e-19 $X=5.815 $Y=1.425 $X2=0
+ $Y2=0
cc_363 N_B2_c_470_n N_A_820_392#_c_726_n 6.69308e-19 $X=5.35 $Y=1.885 $X2=0
+ $Y2=0
cc_364 N_B2_c_472_n N_A_820_392#_c_726_n 0.0105394f $X=5.8 $Y=1.885 $X2=0 $Y2=0
cc_365 N_B2_c_472_n N_A_820_392#_c_730_n 0.00101726f $X=5.8 $Y=1.885 $X2=0 $Y2=0
cc_366 B2 N_A_820_392#_c_730_n 0.0231165f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_367 N_B2_M1002_g N_VGND_c_798_n 0.00291649f $X=5.385 $Y=0.69 $X2=0 $Y2=0
cc_368 N_B2_M1012_g N_VGND_c_798_n 0.00433162f $X=5.815 $Y=0.69 $X2=0 $Y2=0
cc_369 N_B2_M1002_g N_VGND_c_802_n 0.0036412f $X=5.385 $Y=0.69 $X2=0 $Y2=0
cc_370 N_B2_M1012_g N_VGND_c_802_n 0.00432528f $X=5.815 $Y=0.69 $X2=0 $Y2=0
cc_371 N_B2_M1002_g N_A_1009_74#_c_881_n 0.017183f $X=5.385 $Y=0.69 $X2=0 $Y2=0
cc_372 N_B2_M1012_g N_A_1009_74#_c_881_n 0.0144965f $X=5.815 $Y=0.69 $X2=0 $Y2=0
cc_373 B2 N_A_1009_74#_c_881_n 0.0434573f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_374 N_B2_c_468_n N_A_1009_74#_c_881_n 0.00459427f $X=5.815 $Y=1.425 $X2=0
+ $Y2=0
cc_375 B2 N_A_1009_74#_c_885_n 0.015544f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_376 N_B1_c_523_n N_VPWR_c_569_n 0.00486623f $X=6.25 $Y=1.885 $X2=0 $Y2=0
cc_377 N_B1_c_525_n N_VPWR_c_569_n 0.00486623f $X=6.7 $Y=1.885 $X2=0 $Y2=0
cc_378 N_B1_c_523_n N_VPWR_c_572_n 0.00445602f $X=6.25 $Y=1.885 $X2=0 $Y2=0
cc_379 N_B1_c_525_n N_VPWR_c_577_n 0.00445602f $X=6.7 $Y=1.885 $X2=0 $Y2=0
cc_380 N_B1_c_523_n N_VPWR_c_564_n 0.00857673f $X=6.25 $Y=1.885 $X2=0 $Y2=0
cc_381 N_B1_c_525_n N_VPWR_c_564_n 0.00861067f $X=6.7 $Y=1.885 $X2=0 $Y2=0
cc_382 N_B1_c_523_n N_A_820_392#_c_726_n 0.0103374f $X=6.25 $Y=1.885 $X2=0 $Y2=0
cc_383 N_B1_c_525_n N_A_820_392#_c_726_n 6.45594e-19 $X=6.7 $Y=1.885 $X2=0 $Y2=0
cc_384 N_B1_c_523_n N_A_820_392#_c_727_n 0.016798f $X=6.25 $Y=1.885 $X2=0 $Y2=0
cc_385 N_B1_c_525_n N_A_820_392#_c_727_n 0.0124546f $X=6.7 $Y=1.885 $X2=0 $Y2=0
cc_386 B1 N_A_820_392#_c_727_n 0.0312895f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_387 N_B1_c_521_n N_A_820_392#_c_727_n 4.05102e-19 $X=6.715 $Y=1.425 $X2=0
+ $Y2=0
cc_388 N_B1_c_525_n N_A_820_392#_c_728_n 0.00108926f $X=6.7 $Y=1.885 $X2=0 $Y2=0
cc_389 B1 N_A_820_392#_c_728_n 0.0286026f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_390 N_B1_c_523_n N_A_820_392#_c_729_n 6.45594e-19 $X=6.25 $Y=1.885 $X2=0
+ $Y2=0
cc_391 N_B1_c_525_n N_A_820_392#_c_729_n 0.0104891f $X=6.7 $Y=1.885 $X2=0 $Y2=0
cc_392 N_B1_c_523_n N_A_820_392#_c_730_n 0.00192014f $X=6.25 $Y=1.885 $X2=0
+ $Y2=0
cc_393 N_B1_M1007_g N_VGND_c_796_n 0.00502457f $X=6.245 $Y=0.69 $X2=0 $Y2=0
cc_394 N_B1_M1009_g N_VGND_c_796_n 0.00503476f $X=6.715 $Y=0.69 $X2=0 $Y2=0
cc_395 N_B1_M1007_g N_VGND_c_797_n 0.00226696f $X=6.245 $Y=0.69 $X2=0 $Y2=0
cc_396 N_B1_M1009_g N_VGND_c_797_n 0.00568798f $X=6.715 $Y=0.69 $X2=0 $Y2=0
cc_397 N_B1_M1007_g N_VGND_c_798_n 0.00434272f $X=6.245 $Y=0.69 $X2=0 $Y2=0
cc_398 N_B1_M1009_g N_VGND_c_801_n 0.00383152f $X=6.715 $Y=0.69 $X2=0 $Y2=0
cc_399 N_B1_M1007_g N_VGND_c_802_n 0.00821754f $X=6.245 $Y=0.69 $X2=0 $Y2=0
cc_400 N_B1_M1009_g N_VGND_c_802_n 0.00761163f $X=6.715 $Y=0.69 $X2=0 $Y2=0
cc_401 N_B1_M1007_g N_A_1009_74#_c_883_n 0.0180055f $X=6.245 $Y=0.69 $X2=0 $Y2=0
cc_402 N_B1_M1009_g N_A_1009_74#_c_883_n 0.0140902f $X=6.715 $Y=0.69 $X2=0 $Y2=0
cc_403 B1 N_A_1009_74#_c_883_n 0.0580465f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_404 N_B1_c_521_n N_A_1009_74#_c_883_n 0.00374326f $X=6.715 $Y=1.425 $X2=0
+ $Y2=0
cc_405 N_B1_M1009_g N_A_1009_74#_c_884_n 4.43891e-19 $X=6.715 $Y=0.69 $X2=0
+ $Y2=0
cc_406 N_VPWR_M1003_s N_X_c_651_n 0.00807977f $X=0.6 $Y=1.84 $X2=0 $Y2=0
cc_407 N_VPWR_c_565_n N_X_c_651_n 0.0186335f $X=0.725 $Y=2.305 $X2=0 $Y2=0
cc_408 N_VPWR_c_565_n N_X_c_657_n 0.0563525f $X=0.725 $Y=2.305 $X2=0 $Y2=0
cc_409 N_VPWR_c_566_n N_X_c_657_n 0.0547423f $X=1.625 $Y=2.305 $X2=0 $Y2=0
cc_410 N_VPWR_c_570_n N_X_c_657_n 0.014552f $X=1.54 $Y=3.33 $X2=0 $Y2=0
cc_411 N_VPWR_c_564_n N_X_c_657_n 0.0119791f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_412 N_VPWR_M1008_s N_X_c_658_n 0.00247267f $X=1.475 $Y=1.84 $X2=0 $Y2=0
cc_413 N_VPWR_c_566_n N_X_c_658_n 0.0136682f $X=1.625 $Y=2.305 $X2=0 $Y2=0
cc_414 N_VPWR_c_566_n N_X_c_659_n 0.0547423f $X=1.625 $Y=2.305 $X2=0 $Y2=0
cc_415 N_VPWR_c_567_n N_X_c_659_n 0.0386644f $X=2.595 $Y=2.115 $X2=0 $Y2=0
cc_416 N_VPWR_c_575_n N_X_c_659_n 0.014552f $X=2.41 $Y=3.33 $X2=0 $Y2=0
cc_417 N_VPWR_c_564_n N_X_c_659_n 0.0119791f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_418 N_VPWR_c_568_n N_A_820_392#_c_722_n 0.0123543f $X=5.575 $Y=2.455 $X2=0
+ $Y2=0
cc_419 N_VPWR_c_576_n N_A_820_392#_c_722_n 0.053749f $X=5.41 $Y=3.33 $X2=0 $Y2=0
cc_420 N_VPWR_c_564_n N_A_820_392#_c_722_n 0.029846f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_421 N_VPWR_c_576_n N_A_820_392#_c_723_n 0.0236039f $X=5.41 $Y=3.33 $X2=0
+ $Y2=0
cc_422 N_VPWR_c_564_n N_A_820_392#_c_723_n 0.012761f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_423 N_VPWR_c_568_n N_A_820_392#_c_734_n 0.0403584f $X=5.575 $Y=2.455 $X2=0
+ $Y2=0
cc_424 N_VPWR_M1016_d N_A_820_392#_c_725_n 0.00222494f $X=5.425 $Y=1.96 $X2=0
+ $Y2=0
cc_425 N_VPWR_c_568_n N_A_820_392#_c_725_n 0.0154248f $X=5.575 $Y=2.455 $X2=0
+ $Y2=0
cc_426 N_VPWR_c_568_n N_A_820_392#_c_726_n 0.0462948f $X=5.575 $Y=2.455 $X2=0
+ $Y2=0
cc_427 N_VPWR_c_569_n N_A_820_392#_c_726_n 0.0449718f $X=6.475 $Y=2.455 $X2=0
+ $Y2=0
cc_428 N_VPWR_c_572_n N_A_820_392#_c_726_n 0.014552f $X=6.39 $Y=3.33 $X2=0 $Y2=0
cc_429 N_VPWR_c_564_n N_A_820_392#_c_726_n 0.0119791f $X=6.96 $Y=3.33 $X2=0
+ $Y2=0
cc_430 N_VPWR_M1000_d N_A_820_392#_c_727_n 0.00247267f $X=6.325 $Y=1.96 $X2=0
+ $Y2=0
cc_431 N_VPWR_c_569_n N_A_820_392#_c_727_n 0.0136682f $X=6.475 $Y=2.455 $X2=0
+ $Y2=0
cc_432 N_VPWR_c_569_n N_A_820_392#_c_729_n 0.0449718f $X=6.475 $Y=2.455 $X2=0
+ $Y2=0
cc_433 N_VPWR_c_577_n N_A_820_392#_c_729_n 0.0145938f $X=6.96 $Y=3.33 $X2=0
+ $Y2=0
cc_434 N_VPWR_c_564_n N_A_820_392#_c_729_n 0.0120466f $X=6.96 $Y=3.33 $X2=0
+ $Y2=0
cc_435 N_X_c_651_n N_VGND_M1001_d 0.00300749f $X=0.835 $Y=1.885 $X2=-0.19
+ $Y2=-0.245
cc_436 N_X_c_653_n N_VGND_M1010_d 0.00176461f $X=1.795 $Y=1.045 $X2=0 $Y2=0
cc_437 N_X_c_651_n N_VGND_c_786_n 0.0224079f $X=0.835 $Y=1.885 $X2=0 $Y2=0
cc_438 N_X_c_652_n N_VGND_c_786_n 0.0158413f $X=1.1 $Y=0.515 $X2=0 $Y2=0
cc_439 N_X_c_652_n N_VGND_c_787_n 0.0158413f $X=1.1 $Y=0.515 $X2=0 $Y2=0
cc_440 N_X_c_653_n N_VGND_c_787_n 0.0152916f $X=1.795 $Y=1.045 $X2=0 $Y2=0
cc_441 N_X_c_654_n N_VGND_c_787_n 0.0158413f $X=1.96 $Y=0.515 $X2=0 $Y2=0
cc_442 N_X_c_654_n N_VGND_c_788_n 0.0175587f $X=1.96 $Y=0.515 $X2=0 $Y2=0
cc_443 N_X_c_652_n N_VGND_c_792_n 0.0109942f $X=1.1 $Y=0.515 $X2=0 $Y2=0
cc_444 N_X_c_654_n N_VGND_c_794_n 0.0109942f $X=1.96 $Y=0.515 $X2=0 $Y2=0
cc_445 N_X_c_652_n N_VGND_c_802_n 0.00904371f $X=1.1 $Y=0.515 $X2=0 $Y2=0
cc_446 N_X_c_654_n N_VGND_c_802_n 0.00904371f $X=1.96 $Y=0.515 $X2=0 $Y2=0
cc_447 N_VGND_c_802_n N_A_1009_74#_c_881_n 0.00730683f $X=6.96 $Y=0 $X2=0 $Y2=0
cc_448 N_VGND_c_796_n N_A_1009_74#_c_882_n 0.0152763f $X=6.48 $Y=0.55 $X2=0
+ $Y2=0
cc_449 N_VGND_c_798_n N_A_1009_74#_c_882_n 0.00749631f $X=6.495 $Y=0 $X2=0 $Y2=0
cc_450 N_VGND_c_802_n N_A_1009_74#_c_882_n 0.0062048f $X=6.96 $Y=0 $X2=0 $Y2=0
cc_451 N_VGND_M1007_s N_A_1009_74#_c_883_n 0.00218982f $X=6.32 $Y=0.37 $X2=0
+ $Y2=0
cc_452 N_VGND_c_796_n N_A_1009_74#_c_883_n 0.019937f $X=6.48 $Y=0.55 $X2=0 $Y2=0
cc_453 N_VGND_c_796_n N_A_1009_74#_c_884_n 0.0153177f $X=6.48 $Y=0.55 $X2=0
+ $Y2=0
cc_454 N_VGND_c_801_n N_A_1009_74#_c_884_n 0.011066f $X=6.96 $Y=0 $X2=0 $Y2=0
cc_455 N_VGND_c_802_n N_A_1009_74#_c_884_n 0.00915947f $X=6.96 $Y=0 $X2=0 $Y2=0
