* File: sky130_fd_sc_ls__mux2_2.pex.spice
* Created: Wed Sep  2 11:10:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__MUX2_2%A0 1 3 4 6 7
r23 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.385 $X2=0.27 $Y2=1.385
r24 7 11 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.27 $Y=1.295 $X2=0.27
+ $Y2=1.385
r25 4 10 39.305 $w=3.85e-07 $l=2.5446e-07 $layer=POLY_cond $X=0.55 $Y=1.22
+ $X2=0.365 $Y2=1.385
r26 4 6 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.55 $Y=1.22 $X2=0.55
+ $Y2=0.74
r27 1 10 66.2218 $w=3.85e-07 $l=4.44522e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.365 $Y2=1.385
r28 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_LS__MUX2_2%A1 1 3 4 6 7 11
c30 1 0 4.93157e-20 $X=0.955 $Y=1.765
r31 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.03
+ $Y=1.385 $X2=1.03 $Y2=1.385
r32 7 11 9.6556 $w=3.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.72 $Y=1.365 $X2=1.03
+ $Y2=1.365
r33 4 10 38.9663 $w=3.64e-07 $l=2.36525e-07 $layer=POLY_cond $X=1.275 $Y=1.22
+ $X2=1.107 $Y2=1.385
r34 4 6 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.275 $Y=1.22 $X2=1.275
+ $Y2=0.74
r35 1 10 67.4361 $w=3.64e-07 $l=4.49622e-07 $layer=POLY_cond $X=0.955 $Y=1.765
+ $X2=1.107 $Y2=1.385
r36 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.955 $Y=1.765
+ $X2=0.955 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_LS__MUX2_2%S 3 5 7 9 12 14 16 17 18 20 21 22 23 29 36 39
+ 44
c97 36 0 1.85606e-19 $X=1.88 $Y=1.615
c98 14 0 1.11024e-19 $X=3.725 $Y=1.765
r99 39 44 1.92074 $w=3.28e-07 $l=5.5e-08 $layer=LI1_cond $X=2.215 $Y=1.615
+ $X2=2.16 $Y2=1.615
r100 36 38 11.073 $w=3.7e-07 $l=8.5e-08 $layer=POLY_cond $X=1.88 $Y=1.667
+ $X2=1.965 $Y2=1.667
r101 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.88
+ $Y=1.615 $X2=1.88 $Y2=1.615
r102 34 36 28.0081 $w=3.7e-07 $l=2.15e-07 $layer=POLY_cond $X=1.665 $Y=1.667
+ $X2=1.88 $Y2=1.667
r103 29 39 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.3 $Y=1.615
+ $X2=2.215 $Y2=1.615
r104 29 44 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=2.145 $Y=1.615
+ $X2=2.16 $Y2=1.615
r105 29 37 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=2.145 $Y=1.615
+ $X2=1.88 $Y2=1.615
r106 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.29
+ $Y=1.295 $X2=3.29 $Y2=1.295
r107 23 26 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=3.29 $Y=1.215 $X2=3.29
+ $Y2=1.295
r108 21 23 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.125 $Y=1.215
+ $X2=3.29 $Y2=1.215
r109 21 22 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=3.125 $Y=1.215
+ $X2=2.385 $Y2=1.215
r110 20 29 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.3 $Y=1.45 $X2=2.3
+ $Y2=1.615
r111 19 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.3 $Y=1.3
+ $X2=2.385 $Y2=1.215
r112 19 20 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=2.3 $Y=1.3 $X2=2.3
+ $Y2=1.45
r113 17 27 60.3271 $w=3.3e-07 $l=3.45e-07 $layer=POLY_cond $X=3.635 $Y=1.295
+ $X2=3.29 $Y2=1.295
r114 17 18 3.90195 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.635 $Y=1.295
+ $X2=3.725 $Y2=1.295
r115 14 16 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=3.725 $Y=1.765
+ $X2=3.725 $Y2=2.26
r116 10 18 34.7346 $w=1.65e-07 $l=1.67481e-07 $layer=POLY_cond $X=3.72 $Y=1.13
+ $X2=3.725 $Y2=1.295
r117 10 12 248.691 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=3.72 $Y=1.13
+ $X2=3.72 $Y2=0.645
r118 9 14 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.725 $Y=1.675
+ $X2=3.725 $Y2=1.765
r119 8 18 34.7346 $w=1.65e-07 $l=1.65e-07 $layer=POLY_cond $X=3.725 $Y=1.46
+ $X2=3.725 $Y2=1.295
r120 8 9 83.5726 $w=1.8e-07 $l=2.15e-07 $layer=POLY_cond $X=3.725 $Y=1.46
+ $X2=3.725 $Y2=1.675
r121 5 38 23.9667 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=1.965 $Y=1.885
+ $X2=1.965 $Y2=1.667
r122 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.965 $Y=1.885
+ $X2=1.965 $Y2=2.46
r123 1 34 23.9667 $w=1.5e-07 $l=2.17e-07 $layer=POLY_cond $X=1.665 $Y=1.45
+ $X2=1.665 $Y2=1.667
r124 1 3 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.665 $Y=1.45
+ $X2=1.665 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__MUX2_2%A_459_48# 1 2 9 11 13 14 18 23 28 29 34 36
c76 14 0 1.43329e-19 $X=3.335 $Y=1.715
r77 33 34 8.63679 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=3.567 $Y=0.77
+ $X2=3.567 $Y2=0.94
r78 29 34 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.71 $Y=1.63 $X2=3.71
+ $Y2=0.94
r79 28 31 7.93052 $w=4.58e-07 $l=3.05e-07 $layer=LI1_cond $X=3.565 $Y=1.715
+ $X2=3.565 $Y2=2.02
r80 28 29 7.19996 $w=4.58e-07 $l=8.5e-08 $layer=LI1_cond $X=3.565 $Y=1.715
+ $X2=3.565 $Y2=1.63
r81 24 36 31.269 $w=3.16e-07 $l=2.05e-07 $layer=POLY_cond $X=2.72 $Y=1.677
+ $X2=2.515 $Y2=1.677
r82 23 26 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=2.72 $Y=1.635 $X2=2.72
+ $Y2=1.715
r83 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.72
+ $Y=1.635 $X2=2.72 $Y2=1.635
r84 18 33 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=3.505 $Y=0.645
+ $X2=3.505 $Y2=0.77
r85 15 26 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.885 $Y=1.715
+ $X2=2.72 $Y2=1.715
r86 14 28 6.6364 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=3.335 $Y=1.715
+ $X2=3.565 $Y2=1.715
r87 14 15 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=3.335 $Y=1.715
+ $X2=2.885 $Y2=1.715
r88 11 36 20.1942 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.515 $Y=1.885
+ $X2=2.515 $Y2=1.677
r89 11 13 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.515 $Y=1.885
+ $X2=2.515 $Y2=2.46
r90 7 36 22.1171 $w=3.16e-07 $l=2.69933e-07 $layer=POLY_cond $X=2.37 $Y=1.47
+ $X2=2.515 $Y2=1.677
r91 7 9 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=2.37 $Y=1.47 $X2=2.37
+ $Y2=0.74
r92 2 31 600 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_PDIFF $count=1 $X=3.355
+ $Y=1.84 $X2=3.5 $Y2=2.02
r93 1 18 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=3.36
+ $Y=0.37 $X2=3.505 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_LS__MUX2_2%A_116_368# 1 2 7 9 12 16 18 20 21 26 28 30 34
+ 37 38 41 42 43 46 47 51
c105 37 0 1.6439e-20 $X=1.45 $Y=1.82
r106 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5
+ $Y=1.465 $X2=5 $Y2=1.465
r107 44 46 29.5095 $w=3.28e-07 $l=8.45e-07 $layer=LI1_cond $X=5 $Y=2.31 $X2=5
+ $Y2=1.465
r108 42 44 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.835 $Y=2.395
+ $X2=5 $Y2=2.31
r109 42 43 108.952 $w=1.68e-07 $l=1.67e-06 $layer=LI1_cond $X=4.835 $Y=2.395
+ $X2=3.165 $Y2=2.395
r110 41 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.08 $Y=2.31
+ $X2=3.165 $Y2=2.395
r111 40 41 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.08 $Y=2.14
+ $X2=3.08 $Y2=2.31
r112 39 51 3.77418 $w=2.45e-07 $l=1.16619e-07 $layer=LI1_cond $X=1.535 $Y=2.055
+ $X2=1.45 $Y2=1.98
r113 38 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.995 $Y=2.055
+ $X2=3.08 $Y2=2.14
r114 38 39 95.2513 $w=1.68e-07 $l=1.46e-06 $layer=LI1_cond $X=2.995 $Y=2.055
+ $X2=1.535 $Y2=2.055
r115 37 51 2.68609 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=1.45 $Y=1.82
+ $X2=1.45 $Y2=1.98
r116 36 37 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=1.45 $Y=1.01
+ $X2=1.45 $Y2=1.82
r117 35 50 2.90278 $w=3.2e-07 $l=1.1e-07 $layer=LI1_cond $X=0.84 $Y=1.98
+ $X2=0.73 $Y2=1.98
r118 34 51 3.77418 $w=2.45e-07 $l=8.5e-08 $layer=LI1_cond $X=1.365 $Y=1.98
+ $X2=1.45 $Y2=1.98
r119 34 35 18.9073 $w=3.18e-07 $l=5.25e-07 $layer=LI1_cond $X=1.365 $Y=1.98
+ $X2=0.84 $Y2=1.98
r120 30 36 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.365 $Y=0.845
+ $X2=1.45 $Y2=1.01
r121 30 32 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=1.365 $Y=0.845
+ $X2=0.92 $Y2=0.845
r122 26 50 4.22222 $w=2.2e-07 $l=1.6e-07 $layer=LI1_cond $X=0.73 $Y=2.14
+ $X2=0.73 $Y2=1.98
r123 26 28 22.0012 $w=2.18e-07 $l=4.2e-07 $layer=LI1_cond $X=0.73 $Y=2.14
+ $X2=0.73 $Y2=2.56
r124 24 25 0.63089 $w=3.82e-07 $l=5e-09 $layer=POLY_cond $X=4.715 $Y=1.532
+ $X2=4.72 $Y2=1.532
r125 23 24 54.2565 $w=3.82e-07 $l=4.3e-07 $layer=POLY_cond $X=4.285 $Y=1.532
+ $X2=4.715 $Y2=1.532
r126 22 23 1.89267 $w=3.82e-07 $l=1.5e-08 $layer=POLY_cond $X=4.27 $Y=1.532
+ $X2=4.285 $Y2=1.532
r127 21 47 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=4.81 $Y=1.465 $X2=5
+ $Y2=1.465
r128 21 25 12.3813 $w=3.82e-07 $l=1.1887e-07 $layer=POLY_cond $X=4.81 $Y=1.465
+ $X2=4.72 $Y2=1.532
r129 18 25 24.74 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=4.72 $Y=1.765
+ $X2=4.72 $Y2=1.532
r130 18 20 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.72 $Y=1.765
+ $X2=4.72 $Y2=2.4
r131 14 24 24.74 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=4.715 $Y=1.3
+ $X2=4.715 $Y2=1.532
r132 14 16 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.715 $Y=1.3
+ $X2=4.715 $Y2=0.74
r133 10 23 24.74 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=4.285 $Y=1.3
+ $X2=4.285 $Y2=1.532
r134 10 12 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.285 $Y=1.3
+ $X2=4.285 $Y2=0.74
r135 7 22 24.74 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=4.27 $Y=1.765
+ $X2=4.27 $Y2=1.532
r136 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.27 $Y=1.765
+ $X2=4.27 $Y2=2.4
r137 2 50 600 $w=1.7e-07 $l=2.43721e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.84 $X2=0.73 $Y2=2.02
r138 2 28 600 $w=1.7e-07 $l=7.91454e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.84 $X2=0.73 $Y2=2.56
r139 1 32 182 $w=1.7e-07 $l=6.04773e-07 $layer=licon1_NDIFF $count=1 $X=0.625
+ $Y=0.37 $X2=0.92 $Y2=0.845
.ends

.subckt PM_SKY130_FD_SC_LS__MUX2_2%A_27_368# 1 2 9 13 14 16
r29 16 18 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=1.74 $Y=2.815
+ $X2=1.74 $Y2=2.99
r30 13 18 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.575 $Y=2.99
+ $X2=1.74 $Y2=2.99
r31 13 14 73.7219 $w=1.68e-07 $l=1.13e-06 $layer=LI1_cond $X=1.575 $Y=2.99
+ $X2=0.445 $Y2=2.99
r32 9 12 24.6204 $w=3.28e-07 $l=7.05e-07 $layer=LI1_cond $X=0.28 $Y=1.99
+ $X2=0.28 $Y2=2.695
r33 7 14 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=2.905
+ $X2=0.445 $Y2=2.99
r34 7 12 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=0.28 $Y=2.905
+ $X2=0.28 $Y2=2.695
r35 2 16 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.595
+ $Y=1.96 $X2=1.74 $Y2=2.815
r36 1 12 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.695
r37 1 9 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.99
.ends

.subckt PM_SKY130_FD_SC_LS__MUX2_2%A_206_368# 1 2 7 11 17
c29 7 0 4.93157e-20 $X=2.575 $Y=2.395
r30 11 14 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=1.18 $Y=2.395
+ $X2=1.18 $Y2=2.52
r31 8 11 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.345 $Y=2.395
+ $X2=1.18 $Y2=2.395
r32 7 17 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.575 $Y=2.395
+ $X2=2.7 $Y2=2.395
r33 7 8 80.246 $w=1.68e-07 $l=1.23e-06 $layer=LI1_cond $X=2.575 $Y=2.395
+ $X2=1.345 $Y2=2.395
r34 2 17 300 $w=1.7e-07 $l=5.85214e-07 $layer=licon1_PDIFF $count=2 $X=2.59
+ $Y=1.96 $X2=2.74 $Y2=2.475
r35 1 14 600 $w=1.7e-07 $l=7.51266e-07 $layer=licon1_PDIFF $count=1 $X=1.03
+ $Y=1.84 $X2=1.18 $Y2=2.52
.ends

.subckt PM_SKY130_FD_SC_LS__MUX2_2%VPWR 1 2 3 12 16 18 20 22 24 32 40 46 49 53
r52 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r53 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r54 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r55 44 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r56 44 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r57 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r58 41 49 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=4.21 $Y=3.33 $X2=4.04
+ $Y2=3.33
r59 41 43 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=4.21 $Y=3.33
+ $X2=4.56 $Y2=3.33
r60 40 52 5.24187 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=4.78 $Y=3.33 $X2=5.03
+ $Y2=3.33
r61 40 43 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=4.78 $Y=3.33
+ $X2=4.56 $Y2=3.33
r62 39 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r63 38 39 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r64 35 38 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.64 $Y=3.33 $X2=3.6
+ $Y2=3.33
r65 33 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.405 $Y=3.33
+ $X2=2.24 $Y2=3.33
r66 33 35 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=2.405 $Y=3.33
+ $X2=2.64 $Y2=3.33
r67 32 49 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=3.87 $Y=3.33 $X2=4.04
+ $Y2=3.33
r68 32 38 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=3.87 $Y=3.33 $X2=3.6
+ $Y2=3.33
r69 31 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r70 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r71 27 31 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.68 $Y2=3.33
r72 26 30 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=1.68 $Y2=3.33
r73 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r74 24 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.075 $Y=3.33
+ $X2=2.24 $Y2=3.33
r75 24 30 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=2.075 $Y=3.33
+ $X2=1.68 $Y2=3.33
r76 22 39 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r77 22 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r78 22 35 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r79 18 52 2.99835 $w=3.85e-07 $l=1.1025e-07 $layer=LI1_cond $X=4.972 $Y=3.245
+ $X2=5.03 $Y2=3.33
r80 18 20 12.8714 $w=3.83e-07 $l=4.3e-07 $layer=LI1_cond $X=4.972 $Y=3.245
+ $X2=4.972 $Y2=2.815
r81 14 49 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=4.04 $Y=3.245
+ $X2=4.04 $Y2=3.33
r82 14 16 14.575 $w=3.38e-07 $l=4.3e-07 $layer=LI1_cond $X=4.04 $Y=3.245
+ $X2=4.04 $Y2=2.815
r83 10 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.24 $Y=3.245
+ $X2=2.24 $Y2=3.33
r84 10 12 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.24 $Y=3.245
+ $X2=2.24 $Y2=2.815
r85 3 20 600 $w=1.7e-07 $l=1.05889e-06 $layer=licon1_PDIFF $count=1 $X=4.795
+ $Y=1.84 $X2=4.97 $Y2=2.815
r86 2 16 600 $w=1.7e-07 $l=1.0884e-06 $layer=licon1_PDIFF $count=1 $X=3.8
+ $Y=1.84 $X2=4.04 $Y2=2.815
r87 1 12 600 $w=1.7e-07 $l=9.4975e-07 $layer=licon1_PDIFF $count=1 $X=2.04
+ $Y=1.96 $X2=2.24 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_LS__MUX2_2%X 1 2 7 8 9
r19 9 23 6.06583 $w=6.98e-07 $l=3.55e-07 $layer=LI1_cond $X=4.315 $Y=1.665
+ $X2=4.315 $Y2=2.02
r20 8 9 6.32213 $w=6.98e-07 $l=3.7e-07 $layer=LI1_cond $X=4.315 $Y=1.295
+ $X2=4.315 $Y2=1.665
r21 8 17 5.89496 $w=6.98e-07 $l=3.45e-07 $layer=LI1_cond $X=4.315 $Y=1.295
+ $X2=4.315 $Y2=0.95
r22 7 17 0.427171 $w=6.98e-07 $l=2.5e-08 $layer=LI1_cond $X=4.315 $Y=0.925
+ $X2=4.315 $Y2=0.95
r23 2 23 600 $w=1.7e-07 $l=2.43721e-07 $layer=licon1_PDIFF $count=1 $X=4.345
+ $Y=1.84 $X2=4.495 $Y2=2.02
r24 1 17 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=4.36
+ $Y=0.37 $X2=4.5 $Y2=0.95
.ends

.subckt PM_SKY130_FD_SC_LS__MUX2_2%A_38_74# 1 2 9 11 12 13
r29 13 16 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=2.585 $Y=0.375
+ $X2=2.585 $Y2=0.495
r30 11 13 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.42 $Y=0.375
+ $X2=2.585 $Y2=0.375
r31 11 12 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=2.42 $Y=0.375
+ $X2=0.5 $Y2=0.375
r32 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.335 $Y=0.46
+ $X2=0.5 $Y2=0.375
r33 7 9 1.92074 $w=3.28e-07 $l=5.5e-08 $layer=LI1_cond $X=0.335 $Y=0.46
+ $X2=0.335 $Y2=0.515
r34 2 16 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=2.445
+ $Y=0.37 $X2=2.585 $Y2=0.495
r35 1 9 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.19
+ $Y=0.37 $X2=0.335 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__MUX2_2%VGND 1 2 3 10 13 16 18 20 22 28 29 30 39 43
+ 49 53
c69 10 0 2.17911e-19 $X=3 $Y=0.875
r70 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r71 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r72 47 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r73 47 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r74 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r75 44 49 9.6488 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=4.23 $Y=0 $X2=4.035
+ $Y2=0
r76 44 46 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=4.23 $Y=0 $X2=4.56
+ $Y2=0
r77 43 52 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=4.835 $Y=0 $X2=5.057
+ $Y2=0
r78 43 46 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.835 $Y=0 $X2=4.56
+ $Y2=0
r79 42 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r80 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r81 39 49 9.6488 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=3.84 $Y=0 $X2=4.035
+ $Y2=0
r82 39 41 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=3.84 $Y=0 $X2=3.6
+ $Y2=0
r83 33 37 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=2.64
+ $Y2=0
r84 33 34 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r85 30 42 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r86 30 34 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=2.64 $Y=0 $X2=0.24
+ $Y2=0
r87 30 37 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r88 28 37 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=3 $Y=0 $X2=2.64
+ $Y2=0
r89 28 29 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3 $Y=0 $X2=3.085
+ $Y2=0
r90 27 41 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=3.17 $Y=0 $X2=3.6
+ $Y2=0
r91 27 29 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.17 $Y=0 $X2=3.085
+ $Y2=0
r92 22 25 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=1.88 $Y=0.875
+ $X2=1.88 $Y2=0.96
r93 18 52 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=5 $Y=0.085
+ $X2=5.057 $Y2=0
r94 18 20 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=5 $Y=0.085 $X2=5
+ $Y2=0.515
r95 14 49 1.39532 $w=3.9e-07 $l=8.5e-08 $layer=LI1_cond $X=4.035 $Y=0.085
+ $X2=4.035 $Y2=0
r96 14 16 12.7064 $w=3.88e-07 $l=4.3e-07 $layer=LI1_cond $X=4.035 $Y=0.085
+ $X2=4.035 $Y2=0.515
r97 12 29 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.085 $Y=0.085
+ $X2=3.085 $Y2=0
r98 12 13 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=3.085 $Y=0.085
+ $X2=3.085 $Y2=0.79
r99 11 22 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.045 $Y=0.875
+ $X2=1.88 $Y2=0.875
r100 10 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3 $Y=0.875
+ $X2=3.085 $Y2=0.79
r101 10 11 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=3 $Y=0.875
+ $X2=2.045 $Y2=0.875
r102 3 20 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=4.79
+ $Y=0.37 $X2=5 $Y2=0.515
r103 2 16 182 $w=1.7e-07 $l=3.03974e-07 $layer=licon1_NDIFF $count=1 $X=3.795
+ $Y=0.37 $X2=4.035 $Y2=0.515
r104 1 25 182 $w=1.7e-07 $l=6.56277e-07 $layer=licon1_NDIFF $count=1 $X=1.74
+ $Y=0.37 $X2=1.88 $Y2=0.96
.ends

