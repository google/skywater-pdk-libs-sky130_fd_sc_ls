* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__sedfxbp_2 CLK D DE SCD SCE VGND VNB VPB VPWR Q Q_N
M1000 a_691_113# a_661_87# a_1088_453# VPB phighvt w=640000u l=150000u
+  ad=5.015e+11p pd=5.17e+06u as=1.728e+11p ps=1.82e+06u
M1001 a_1586_74# a_1374_368# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=3.65505e+12p ps=2.974e+07u
M1002 VPWR a_2013_71# a_1944_508# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.512e+11p ps=1.56e+06u
M1003 a_1586_74# a_1374_368# VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=2.61097e+12p ps=2.285e+07u
M1004 a_132_464# D a_32_74# VPB phighvt w=640000u l=150000u
+  ad=1.728e+11p pd=1.82e+06u as=3.808e+11p ps=3.75e+06u
M1005 Q a_2489_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=0p ps=0u
M1006 a_32_74# a_575_87# a_527_113# VNB nshort w=420000u l=150000u
+  ad=2.835e+11p pd=3.03e+06u as=1.008e+11p ps=1.32e+06u
M1007 a_1374_368# CLK VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=0p ps=0u
M1008 a_1784_97# a_1586_74# a_691_113# VPB phighvt w=420000u l=150000u
+  ad=1.26e+11p pd=1.44e+06u as=0p ps=0u
M1009 a_2417_74# a_2013_71# VGND VNB nshort w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1010 a_691_113# a_661_87# a_32_74# VNB nshort w=420000u l=150000u
+  ad=3.885e+11p pd=4.37e+06u as=0p ps=0u
M1011 a_2489_74# a_1586_74# a_2417_74# VNB nshort w=640000u l=150000u
+  ad=2.139e+11p pd=2e+06u as=0p ps=0u
M1012 a_1088_453# SCD VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_2591_74# a_1374_368# a_2489_74# VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1014 a_575_87# a_2489_74# VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1015 a_2489_74# a_1374_368# a_2374_392# VPB phighvt w=1e+06u l=150000u
+  ad=3.328e+11p pd=2.77e+06u as=8.05e+11p ps=3.61e+06u
M1016 VPWR a_2489_74# Q VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR DE a_183_290# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.888e+11p ps=1.87e+06u
M1018 a_32_74# a_575_87# a_578_462# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.536e+11p ps=1.76e+06u
M1019 a_1944_508# a_1374_368# a_1784_97# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_575_87# a_2489_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=0p ps=0u
M1021 a_1091_125# SCD VGND VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1022 VPWR a_575_87# a_2672_508# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1023 a_2013_71# a_1784_97# VGND VNB nshort w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=0p ps=0u
M1024 a_527_113# a_183_290# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_2672_508# a_1586_74# a_2489_74# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VGND a_575_87# a_2591_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 Q_N a_575_87# VGND VNB nshort w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1028 VGND DE a_183_290# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1029 VPWR a_183_290# a_132_464# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_2013_71# a_1784_97# VPWR VPB phighvt w=840000u l=150000u
+  ad=2.478e+11p pd=2.27e+06u as=0p ps=0u
M1031 Q_N a_575_87# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=0p ps=0u
M1032 Q a_2489_74# VGND VNB nshort w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1033 a_691_113# SCE a_32_74# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 VGND a_2013_71# a_1920_97# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.953e+11p ps=1.77e+06u
M1035 a_1374_368# CLK VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1036 a_691_113# SCE a_1091_125# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_1784_97# a_1374_368# a_691_113# VNB nshort w=420000u l=150000u
+  ad=2.226e+11p pd=1.9e+06u as=0p ps=0u
M1038 VPWR a_575_87# Q_N VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 VGND SCE a_661_87# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1040 a_1920_97# a_1586_74# a_1784_97# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1041 VGND a_575_87# Q_N VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1042 VGND DE a_141_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1043 VGND a_2489_74# Q VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1044 a_578_462# DE VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1045 VPWR SCE a_661_87# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.952e+11p ps=1.89e+06u
M1046 a_2374_392# a_2013_71# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1047 a_141_74# D a_32_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
