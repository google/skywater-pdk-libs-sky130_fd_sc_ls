# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ls__nor3_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_ls__nor3_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.447000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.650000 0.310000 3.235000 0.980000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.447000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.305000 1.220000 1.635000 1.380000 ;
        RECT 1.305000 1.380000 3.255000 1.550000 ;
        RECT 2.925000 1.180000 3.255000 1.380000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.447000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.180000 0.975000 1.550000 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  0.861900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115000 0.350000 0.445000 0.840000 ;
        RECT 0.115000 0.840000 1.980000 1.010000 ;
        RECT 0.115000 1.010000 0.355000 1.720000 ;
        RECT 0.115000 1.720000 0.945000 1.890000 ;
        RECT 0.615000 1.890000 0.945000 2.735000 ;
        RECT 1.650000 0.350000 1.980000 0.840000 ;
        RECT 1.650000 1.010000 1.980000 1.050000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.115000  2.060000 0.445000 2.905000 ;
      RECT 0.115000  2.905000 1.315000 3.075000 ;
      RECT 0.615000  0.085000 1.480000 0.650000 ;
      RECT 1.145000  1.720000 3.245000 1.890000 ;
      RECT 1.145000  1.890000 1.315000 2.905000 ;
      RECT 1.515000  2.060000 2.795000 2.230000 ;
      RECT 1.515000  2.230000 1.845000 2.990000 ;
      RECT 2.015000  2.400000 2.345000 3.245000 ;
      RECT 2.150000  0.085000 2.480000 1.130000 ;
      RECT 2.515000  2.230000 2.795000 2.990000 ;
      RECT 2.965000  1.890000 3.245000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_ls__nor3_2
END LIBRARY
