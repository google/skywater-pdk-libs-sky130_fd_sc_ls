* NGSPICE file created from sky130_fd_sc_ls__o311ai_1.ext - technology: sky130A

.subckt sky130_fd_sc_ls__o311ai_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
M1000 Y C1 a_469_74# VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=2.294e+11p ps=2.1e+06u
M1001 Y A3 a_222_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=8.008e+11p pd=5.91e+06u as=4.704e+11p ps=3.08e+06u
M1002 a_128_74# A1 VGND VNB nshort w=740000u l=150000u
+  ad=4.847e+11p pd=4.27e+06u as=7.067e+11p ps=4.87e+06u
M1003 a_138_368# A1 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.024e+11p pd=2.78e+06u as=8.008e+11p ps=5.91e+06u
M1004 Y C1 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_469_74# B1 a_128_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR B1 Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND A2 a_128_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_222_368# A2 a_138_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_128_74# A3 VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

