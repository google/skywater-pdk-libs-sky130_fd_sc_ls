* File: sky130_fd_sc_ls__a41o_1.pex.spice
* Created: Fri Aug 28 13:01:10 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__A41O_1%A_83_244# 1 2 7 9 10 12 14 16 17 26 28 32 34
+ 36 37
c63 28 0 1.71268e-19 $X=1.79 $Y=1.195
c64 16 0 1.09203e-19 $X=1.095 $Y=1.385
r65 36 37 9.45624 $w=4.88e-07 $l=1.65e-07 $layer=LI1_cond $X=1.39 $Y=2.115
+ $X2=1.39 $Y2=1.95
r66 30 32 20.7789 $w=3.28e-07 $l=5.95e-07 $layer=LI1_cond $X=1.955 $Y=1.11
+ $X2=1.955 $Y2=0.515
r67 29 34 3.10218 $w=3.05e-07 $l=1.72337e-07 $layer=LI1_cond $X=1.315 $Y=1.195
+ $X2=1.23 $Y2=1.33
r68 28 30 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.79 $Y=1.195
+ $X2=1.955 $Y2=1.11
r69 28 29 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=1.79 $Y=1.195
+ $X2=1.315 $Y2=1.195
r70 24 36 1.95278 $w=4.88e-07 $l=8e-08 $layer=LI1_cond $X=1.39 $Y=2.195 $X2=1.39
+ $Y2=2.115
r71 24 26 15.1341 $w=4.88e-07 $l=6.2e-07 $layer=LI1_cond $X=1.39 $Y=2.195
+ $X2=1.39 $Y2=2.815
r72 22 34 3.51065 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=1.23 $Y=1.55 $X2=1.23
+ $Y2=1.33
r73 22 37 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=1.23 $Y=1.55 $X2=1.23
+ $Y2=1.95
r74 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.08
+ $Y=1.385 $X2=1.08 $Y2=1.385
r75 17 34 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.145 $Y=1.33
+ $X2=1.23 $Y2=1.33
r76 17 19 1.70247 $w=4.38e-07 $l=6.5e-08 $layer=LI1_cond $X=1.145 $Y=1.33
+ $X2=1.08 $Y2=1.33
r77 16 20 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.095 $Y=1.385
+ $X2=1.08 $Y2=1.385
r78 14 20 84.8077 $w=3.3e-07 $l=4.85e-07 $layer=POLY_cond $X=0.595 $Y=1.385
+ $X2=1.08 $Y2=1.385
r79 10 16 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=1.17 $Y=1.22
+ $X2=1.095 $Y2=1.385
r80 10 12 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.17 $Y=1.22 $X2=1.17
+ $Y2=0.74
r81 7 14 149.859 $w=1.8e-07 $l=3.8e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=1.385
r82 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.4
r83 2 36 400 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=1 $X=1.325
+ $Y=1.96 $X2=1.47 $Y2=2.115
r84 2 26 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.325
+ $Y=1.96 $X2=1.47 $Y2=2.815
r85 1 32 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.815
+ $Y=0.37 $X2=1.955 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__A41O_1%B1 1 3 6 8
c32 8 0 1.09203e-19 $X=1.68 $Y=1.665
r33 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.65
+ $Y=1.615 $X2=1.65 $Y2=1.615
r34 4 11 38.5916 $w=2.93e-07 $l=2.05122e-07 $layer=POLY_cond $X=1.74 $Y=1.45
+ $X2=1.65 $Y2=1.615
r35 4 6 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.74 $Y=1.45 $X2=1.74
+ $Y2=0.74
r36 1 11 55.8646 $w=2.93e-07 $l=2.91633e-07 $layer=POLY_cond $X=1.695 $Y=1.885
+ $X2=1.65 $Y2=1.615
r37 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.695 $Y=1.885
+ $X2=1.695 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_LS__A41O_1%A1 3 5 7 8
c35 8 0 1.15358e-19 $X=2.16 $Y=1.665
r36 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.19
+ $Y=1.615 $X2=2.19 $Y2=1.615
r37 5 11 55.8646 $w=2.93e-07 $l=2.72489e-07 $layer=POLY_cond $X=2.195 $Y=1.885
+ $X2=2.19 $Y2=1.615
r38 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.195 $Y=1.885
+ $X2=2.195 $Y2=2.46
r39 1 11 38.5916 $w=2.93e-07 $l=1.74714e-07 $layer=POLY_cond $X=2.17 $Y=1.45
+ $X2=2.19 $Y2=1.615
r40 1 3 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=2.17 $Y=1.45 $X2=2.17
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__A41O_1%A2 3 5 6 8 9 10 11 16 18
c41 18 0 2.09165e-19 $X=2.73 $Y=1.22
c42 16 0 1.15358e-19 $X=2.73 $Y=1.385
c43 5 0 9.71067e-20 $X=2.775 $Y=1.795
r44 16 19 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.73 $Y=1.385
+ $X2=2.73 $Y2=1.55
r45 16 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.73 $Y=1.385
+ $X2=2.73 $Y2=1.22
r46 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.73
+ $Y=1.385 $X2=2.73 $Y2=1.385
r47 11 17 2.80324 $w=3.68e-07 $l=9e-08 $layer=LI1_cond $X=2.71 $Y=1.295 $X2=2.71
+ $Y2=1.385
r48 10 11 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.71 $Y=0.925
+ $X2=2.71 $Y2=1.295
r49 9 10 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.71 $Y=0.555
+ $X2=2.71 $Y2=0.925
r50 6 8 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.775 $Y=1.885
+ $X2=2.775 $Y2=2.46
r51 5 6 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.775 $Y=1.795 $X2=2.775
+ $Y2=1.885
r52 5 19 95.2339 $w=1.8e-07 $l=2.45e-07 $layer=POLY_cond $X=2.775 $Y=1.795
+ $X2=2.775 $Y2=1.55
r53 3 18 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.64 $Y=0.74 $X2=2.64
+ $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_LS__A41O_1%A3 3 5 6 8 9 12 14
c37 9 0 3.7897e-20 $X=3.6 $Y=1.295
c38 6 0 6.00847e-21 $X=3.225 $Y=1.885
r39 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.3 $Y=1.385
+ $X2=3.3 $Y2=1.55
r40 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.3 $Y=1.385
+ $X2=3.3 $Y2=1.22
r41 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.3
+ $Y=1.385 $X2=3.3 $Y2=1.385
r42 9 13 9.34413 $w=3.68e-07 $l=3e-07 $layer=LI1_cond $X=3.6 $Y=1.365 $X2=3.3
+ $Y2=1.365
r43 6 8 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.225 $Y=1.885
+ $X2=3.225 $Y2=2.46
r44 5 6 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.225 $Y=1.795 $X2=3.225
+ $Y2=1.885
r45 5 15 95.2339 $w=1.8e-07 $l=2.45e-07 $layer=POLY_cond $X=3.225 $Y=1.795
+ $X2=3.225 $Y2=1.55
r46 3 14 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.21 $Y=0.74 $X2=3.21
+ $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_LS__A41O_1%A4 1 3 5 6 8 9 15
c28 5 0 7.12227e-20 $X=3.795 $Y=1.795
r29 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.05
+ $Y=1.385 $X2=4.05 $Y2=1.385
r30 13 15 44.5896 $w=3.3e-07 $l=2.55e-07 $layer=POLY_cond $X=3.795 $Y=1.385
+ $X2=4.05 $Y2=1.385
r31 11 13 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=3.78 $Y=1.385
+ $X2=3.795 $Y2=1.385
r32 9 16 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=4.05 $Y=1.295 $X2=4.05
+ $Y2=1.385
r33 6 8 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.795 $Y=1.885
+ $X2=3.795 $Y2=2.46
r34 5 6 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.795 $Y=1.795 $X2=3.795
+ $Y2=1.885
r35 4 13 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.795 $Y=1.55
+ $X2=3.795 $Y2=1.385
r36 4 5 95.2339 $w=1.8e-07 $l=2.45e-07 $layer=POLY_cond $X=3.795 $Y=1.55
+ $X2=3.795 $Y2=1.795
r37 1 11 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.78 $Y=1.22
+ $X2=3.78 $Y2=1.385
r38 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.78 $Y=1.22 $X2=3.78
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__A41O_1%X 1 2 7 11 13 17 19 20
r23 15 20 2.39847 $w=6.5e-07 $l=1.2e-07 $layer=LI1_cond $X=0.355 $Y=0.615
+ $X2=0.235 $Y2=0.615
r24 15 17 11.0407 $w=6.48e-07 $l=6e-07 $layer=LI1_cond $X=0.355 $Y=0.615
+ $X2=0.955 $Y2=0.615
r25 11 19 6.63994 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.28 $Y=1.985
+ $X2=0.28 $Y2=1.82
r26 11 13 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=0.28 $Y=1.985
+ $X2=0.28 $Y2=2.815
r27 7 20 6.49586 $w=2.4e-07 $l=3.25e-07 $layer=LI1_cond $X=0.235 $Y=0.94
+ $X2=0.235 $Y2=0.615
r28 7 19 42.2562 $w=2.38e-07 $l=8.8e-07 $layer=LI1_cond $X=0.235 $Y=0.94
+ $X2=0.235 $Y2=1.82
r29 2 13 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r30 2 11 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
r31 1 17 45.5 $w=1.7e-07 $l=8.8955e-07 $layer=licon1_NDIFF $count=4 $X=0.135
+ $Y=0.37 $X2=0.955 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__A41O_1%VPWR 1 2 3 14 20 24 29 30 32 33 34 47 48 51
r49 51 52 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r50 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r51 45 48 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r52 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r53 39 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r54 38 41 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r55 38 39 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r56 36 51 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=0.77 $Y2=3.33
r57 36 38 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=1.2 $Y2=3.33
r58 34 45 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r59 34 39 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.2 $Y2=3.33
r60 34 41 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r61 32 44 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=3.335 $Y=3.33
+ $X2=3.12 $Y2=3.33
r62 32 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.335 $Y=3.33
+ $X2=3.5 $Y2=3.33
r63 31 47 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=3.665 $Y=3.33
+ $X2=4.08 $Y2=3.33
r64 31 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.665 $Y=3.33
+ $X2=3.5 $Y2=3.33
r65 29 41 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=2.305 $Y=3.33
+ $X2=2.16 $Y2=3.33
r66 29 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.305 $Y=3.33
+ $X2=2.47 $Y2=3.33
r67 28 44 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=2.635 $Y=3.33
+ $X2=3.12 $Y2=3.33
r68 28 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.635 $Y=3.33
+ $X2=2.47 $Y2=3.33
r69 24 27 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=3.5 $Y=2.145 $X2=3.5
+ $Y2=2.825
r70 22 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.5 $Y=3.245 $X2=3.5
+ $Y2=3.33
r71 22 27 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=3.5 $Y=3.245 $X2=3.5
+ $Y2=2.825
r72 18 30 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.47 $Y=3.245
+ $X2=2.47 $Y2=3.33
r73 18 20 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=2.47 $Y=3.245
+ $X2=2.47 $Y2=2.455
r74 14 17 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=0.77 $Y=1.985
+ $X2=0.77 $Y2=2.815
r75 12 51 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.77 $Y=3.245
+ $X2=0.77 $Y2=3.33
r76 12 17 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.77 $Y=3.245
+ $X2=0.77 $Y2=2.815
r77 3 27 400 $w=1.7e-07 $l=9.59805e-07 $layer=licon1_PDIFF $count=1 $X=3.3
+ $Y=1.96 $X2=3.5 $Y2=2.825
r78 3 24 400 $w=1.7e-07 $l=2.77489e-07 $layer=licon1_PDIFF $count=1 $X=3.3
+ $Y=1.96 $X2=3.5 $Y2=2.145
r79 2 20 300 $w=1.7e-07 $l=5.86536e-07 $layer=licon1_PDIFF $count=2 $X=2.27
+ $Y=1.96 $X2=2.47 $Y2=2.455
r80 1 17 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.84 $X2=0.73 $Y2=2.815
r81 1 14 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.84 $X2=0.73 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_LS__A41O_1%A_354_392# 1 2 3 10 12 14 18 20 24 30
c57 30 0 7.12227e-20 $X=3 $Y=1.805
c58 20 0 9.71067e-20 $X=3.855 $Y=1.805
c59 14 0 6.00847e-21 $X=2.835 $Y=2.035
r60 32 34 2.44458 $w=3.28e-07 $l=7e-08 $layer=LI1_cond $X=3 $Y=2.035 $X2=3
+ $Y2=2.105
r61 30 32 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=3 $Y=1.805 $X2=3
+ $Y2=2.035
r62 24 26 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=4.02 $Y=2.105
+ $X2=4.02 $Y2=2.815
r63 22 24 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=4.02 $Y=1.89
+ $X2=4.02 $Y2=2.105
r64 21 30 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.165 $Y=1.805 $X2=3
+ $Y2=1.805
r65 20 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.855 $Y=1.805
+ $X2=4.02 $Y2=1.89
r66 20 21 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.855 $Y=1.805
+ $X2=3.165 $Y2=1.805
r67 16 34 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=3 $Y=2.12 $X2=3
+ $Y2=2.105
r68 16 18 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=3 $Y=2.12 $X2=3
+ $Y2=2.815
r69 15 29 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.135 $Y=2.035
+ $X2=1.97 $Y2=2.035
r70 14 32 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.835 $Y=2.035 $X2=3
+ $Y2=2.035
r71 14 15 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=2.835 $Y=2.035
+ $X2=2.135 $Y2=2.035
r72 10 29 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.97 $Y=2.12 $X2=1.97
+ $Y2=2.035
r73 10 12 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=1.97 $Y=2.12
+ $X2=1.97 $Y2=2.815
r74 3 26 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=3.87
+ $Y=1.96 $X2=4.02 $Y2=2.815
r75 3 24 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=3.87
+ $Y=1.96 $X2=4.02 $Y2=2.105
r76 2 34 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.85
+ $Y=1.96 $X2=3 $Y2=2.105
r77 2 18 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=2.85
+ $Y=1.96 $X2=3 $Y2=2.815
r78 1 29 400 $w=1.7e-07 $l=2.66458e-07 $layer=licon1_PDIFF $count=1 $X=1.77
+ $Y=1.96 $X2=1.97 $Y2=2.115
r79 1 12 400 $w=1.7e-07 $l=9.4975e-07 $layer=licon1_PDIFF $count=1 $X=1.77
+ $Y=1.96 $X2=1.97 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_LS__A41O_1%VGND 1 2 9 11 13 16 17 18 27 36
r38 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r39 33 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r40 32 33 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r41 29 32 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.68 $Y=0 $X2=3.6
+ $Y2=0
r42 29 30 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r43 27 35 4.64076 $w=1.7e-07 $l=2.45e-07 $layer=LI1_cond $X=3.83 $Y=0 $X2=4.075
+ $Y2=0
r44 27 32 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=3.83 $Y=0 $X2=3.6
+ $Y2=0
r45 26 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r46 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r47 22 26 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r48 21 25 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r49 21 22 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r50 18 33 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.6
+ $Y2=0
r51 18 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r52 16 25 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=1.29 $Y=0 $X2=1.2
+ $Y2=0
r53 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.29 $Y=0 $X2=1.455
+ $Y2=0
r54 15 29 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=1.62 $Y=0 $X2=1.68
+ $Y2=0
r55 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.62 $Y=0 $X2=1.455
+ $Y2=0
r56 11 35 3.12541 $w=3.3e-07 $l=1.18427e-07 $layer=LI1_cond $X=3.995 $Y=0.085
+ $X2=4.075 $Y2=0
r57 11 13 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.995 $Y=0.085
+ $X2=3.995 $Y2=0.515
r58 7 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.455 $Y=0.085
+ $X2=1.455 $Y2=0
r59 7 9 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=1.455 $Y=0.085
+ $X2=1.455 $Y2=0.515
r60 2 13 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.855
+ $Y=0.37 $X2=3.995 $Y2=0.515
r61 1 9 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=1.245
+ $Y=0.37 $X2=1.455 $Y2=0.515
.ends

