* File: sky130_fd_sc_ls__and3_1.pex.spice
* Created: Fri Aug 28 13:03:50 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__AND3_1%A 4 5 7 8 11 13 17 19 23
r44 19 23 3.89033 $w=4.13e-07 $l=1.15e-07 $layer=LI1_cond $X=1.2 $Y=0.462
+ $X2=1.085 $Y2=0.462
r45 16 23 17.3781 $w=3.13e-07 $l=4.75e-07 $layer=LI1_cond $X=0.61 $Y=0.412
+ $X2=1.085 $Y2=0.412
r46 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.61
+ $Y=0.405 $X2=0.61 $Y2=0.405
r47 12 13 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=0.51 $Y=1.395
+ $X2=0.51 $Y2=1.545
r48 11 12 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.53 $Y=1 $X2=0.53
+ $Y2=1.395
r49 8 17 19.6204 $w=1.5e-07 $l=2.03101e-07 $layer=POLY_cond $X=0.53 $Y=0.57
+ $X2=0.615 $Y2=0.405
r50 8 11 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=0.53 $Y=0.57 $X2=0.53
+ $Y2=1
r51 5 7 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.505 $Y=1.915
+ $X2=0.505 $Y2=2.41
r52 4 5 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.505 $Y=1.825 $X2=0.505
+ $Y2=1.915
r53 4 13 108.839 $w=1.8e-07 $l=2.8e-07 $layer=POLY_cond $X=0.505 $Y=1.825
+ $X2=0.505 $Y2=1.545
.ends

.subckt PM_SKY130_FD_SC_LS__AND3_1%B 1 3 4 6 7 8
r40 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.01
+ $Y=1.595 $X2=1.01 $Y2=1.595
r41 8 13 1.78139 $w=4.68e-07 $l=7e-08 $layer=LI1_cond $X=1.08 $Y=1.665 $X2=1.08
+ $Y2=1.595
r42 7 13 7.63454 $w=4.68e-07 $l=3e-07 $layer=LI1_cond $X=1.08 $Y=1.295 $X2=1.08
+ $Y2=1.595
r43 4 12 38.7026 $w=2.82e-07 $l=2.0106e-07 $layer=POLY_cond $X=1.09 $Y=1.43
+ $X2=1.01 $Y2=1.595
r44 4 6 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.09 $Y=1.43 $X2=1.09
+ $Y2=1
r45 1 12 65.1955 $w=2.82e-07 $l=3.4176e-07 $layer=POLY_cond $X=1.055 $Y=1.915
+ $X2=1.01 $Y2=1.595
r46 1 3 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.055 $Y=1.915
+ $X2=1.055 $Y2=2.41
.ends

.subckt PM_SKY130_FD_SC_LS__AND3_1%C 1 3 6 8
r32 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.65
+ $Y=1.615 $X2=1.65 $Y2=1.615
r33 4 11 38.6446 $w=3.36e-07 $l=1.88348e-07 $layer=POLY_cond $X=1.565 $Y=1.45
+ $X2=1.615 $Y2=1.615
r34 4 6 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.565 $Y=1.45
+ $X2=1.565 $Y2=0.92
r35 1 11 58.0107 $w=3.36e-07 $l=3.50714e-07 $layer=POLY_cond $X=1.505 $Y=1.915
+ $X2=1.615 $Y2=1.615
r36 1 3 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.505 $Y=1.915
+ $X2=1.505 $Y2=2.41
.ends

.subckt PM_SKY130_FD_SC_LS__AND3_1%A_27_398# 1 2 3 10 12 13 15 18 22 24 28 30 33
+ 34 35 37
r72 37 40 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.235 $Y=1.515
+ $X2=2.235 $Y2=1.68
r73 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.235
+ $Y=1.515 $X2=2.235 $Y2=1.515
r74 33 40 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=2.155 $Y=1.95
+ $X2=2.155 $Y2=1.68
r75 31 35 7.75133 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=1.4 $Y=2.035
+ $X2=1.257 $Y2=2.035
r76 30 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.07 $Y=2.035
+ $X2=2.155 $Y2=1.95
r77 30 31 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.07 $Y=2.035
+ $X2=1.4 $Y2=2.035
r78 26 35 0.432977 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=1.257 $Y=2.12
+ $X2=1.257 $Y2=2.035
r79 26 28 0.606549 $w=2.83e-07 $l=1.5e-08 $layer=LI1_cond $X=1.257 $Y=2.12
+ $X2=1.257 $Y2=2.135
r80 25 34 4.00616 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.48 $Y=2.035
+ $X2=0.297 $Y2=2.035
r81 24 35 7.75133 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=1.115 $Y=2.035
+ $X2=1.257 $Y2=2.035
r82 24 25 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.115 $Y=2.035
+ $X2=0.48 $Y2=2.035
r83 20 34 2.75409 $w=3.47e-07 $l=9.31128e-08 $layer=LI1_cond $X=0.28 $Y=2.12
+ $X2=0.297 $Y2=2.035
r84 20 22 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=0.28 $Y=2.12
+ $X2=0.28 $Y2=2.135
r85 16 34 2.75409 $w=3.47e-07 $l=8.5e-08 $layer=LI1_cond $X=0.297 $Y=1.95
+ $X2=0.297 $Y2=2.035
r86 16 18 31.1002 $w=3.63e-07 $l=9.85e-07 $layer=LI1_cond $X=0.297 $Y=1.95
+ $X2=0.297 $Y2=0.965
r87 13 38 50.4896 $w=3.5e-07 $l=2.99165e-07 $layer=POLY_cond $X=2.375 $Y=1.765
+ $X2=2.267 $Y2=1.515
r88 13 15 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.375 $Y=1.765
+ $X2=2.375 $Y2=2.4
r89 10 38 38.7839 $w=3.5e-07 $l=2.17612e-07 $layer=POLY_cond $X=2.145 $Y=1.35
+ $X2=2.267 $Y2=1.515
r90 10 12 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.145 $Y=1.35
+ $X2=2.145 $Y2=0.87
r91 3 28 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=1.13
+ $Y=1.99 $X2=1.28 $Y2=2.135
r92 2 22 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.99 $X2=0.28 $Y2=2.135
r93 1 18 182 $w=1.7e-07 $l=3.50071e-07 $layer=licon1_NDIFF $count=1 $X=0.17
+ $Y=0.68 $X2=0.315 $Y2=0.965
.ends

.subckt PM_SKY130_FD_SC_LS__AND3_1%VPWR 1 2 9 13 15 17 22 29 30 33 36
r38 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r39 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r40 30 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r41 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r42 27 36 14.0645 $w=1.7e-07 $l=3.7e-07 $layer=LI1_cond $X=2.31 $Y=3.33 $X2=1.94
+ $Y2=3.33
r43 27 29 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.31 $Y=3.33
+ $X2=2.64 $Y2=3.33
r44 26 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r45 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r46 23 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=0.78 $Y2=3.33
r47 23 25 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=1.2 $Y2=3.33
r48 22 36 14.0645 $w=1.7e-07 $l=3.7e-07 $layer=LI1_cond $X=1.57 $Y=3.33 $X2=1.94
+ $Y2=3.33
r49 22 25 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.57 $Y=3.33 $X2=1.2
+ $Y2=3.33
r50 20 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r51 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r52 17 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.78 $Y2=3.33
r53 17 19 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.24 $Y2=3.33
r54 15 37 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=2.16 $Y2=3.33
r55 15 26 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.2 $Y2=3.33
r56 11 36 2.97738 $w=7.4e-07 $l=8.5e-08 $layer=LI1_cond $X=1.94 $Y=3.245
+ $X2=1.94 $Y2=3.33
r57 11 13 14.062 $w=7.38e-07 $l=8.7e-07 $layer=LI1_cond $X=1.94 $Y=3.245
+ $X2=1.94 $Y2=2.375
r58 7 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=3.245 $X2=0.78
+ $Y2=3.33
r59 7 9 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=0.78 $Y=3.245 $X2=0.78
+ $Y2=2.455
r60 2 13 150 $w=1.7e-07 $l=7.32632e-07 $layer=licon1_PDIFF $count=4 $X=1.58
+ $Y=1.99 $X2=2.145 $Y2=2.375
r61 1 9 600 $w=1.7e-07 $l=5.5608e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.99 $X2=0.78 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_LS__AND3_1%X 1 2 9 15 17 18 19 27 36
r21 24 27 0.930042 $w=2.83e-07 $l=2.3e-08 $layer=LI1_cond $X=2.622 $Y=1.992
+ $X2=2.622 $Y2=2.015
r22 18 19 14.9615 $w=2.83e-07 $l=3.7e-07 $layer=LI1_cond $X=2.622 $Y=2.405
+ $X2=2.622 $Y2=2.775
r23 17 24 0.849169 $w=2.83e-07 $l=2.1e-08 $layer=LI1_cond $X=2.622 $Y=1.971
+ $X2=2.622 $Y2=1.992
r24 17 36 6.75432 $w=2.83e-07 $l=1.21e-07 $layer=LI1_cond $X=2.622 $Y=1.971
+ $X2=2.622 $Y2=1.85
r25 17 18 14.1124 $w=2.83e-07 $l=3.49e-07 $layer=LI1_cond $X=2.622 $Y=2.056
+ $X2=2.622 $Y2=2.405
r26 17 27 1.6579 $w=2.83e-07 $l=4.1e-08 $layer=LI1_cond $X=2.622 $Y=2.056
+ $X2=2.622 $Y2=2.015
r27 11 15 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.68 $Y=1.18
+ $X2=2.68 $Y2=1.095
r28 11 36 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.68 $Y=1.18
+ $X2=2.68 $Y2=1.85
r29 7 15 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2.36 $Y=1.095 $X2=2.68
+ $Y2=1.095
r30 7 9 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=2.36 $Y=1.01 $X2=2.36
+ $Y2=0.645
r31 2 19 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.45
+ $Y=1.84 $X2=2.6 $Y2=2.815
r32 2 27 400 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=1 $X=2.45
+ $Y=1.84 $X2=2.6 $Y2=2.015
r33 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.22 $Y=0.5
+ $X2=2.36 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_LS__AND3_1%VGND 1 6 11 12 13 23 24
r23 23 24 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r24 21 24 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r25 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r26 16 20 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=1.68
+ $Y2=0
r27 16 17 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r28 13 21 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.68
+ $Y2=0
r29 13 17 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.44 $Y=0 $X2=0.24
+ $Y2=0
r30 11 20 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=1.695 $Y=0 $X2=1.68
+ $Y2=0
r31 11 12 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.695 $Y=0 $X2=1.86
+ $Y2=0
r32 10 23 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=2.025 $Y=0 $X2=2.64
+ $Y2=0
r33 10 12 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.025 $Y=0 $X2=1.86
+ $Y2=0
r34 6 8 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=1.86 $Y=0.645 $X2=1.86
+ $Y2=1.065
r35 4 12 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.86 $Y=0.085 $X2=1.86
+ $Y2=0
r36 4 6 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=1.86 $Y=0.085 $X2=1.86
+ $Y2=0.645
r37 1 8 182 $w=1.7e-07 $l=5.6438e-07 $layer=licon1_NDIFF $count=1 $X=1.64 $Y=0.6
+ $X2=1.86 $Y2=1.065
r38 1 6 182 $w=1.7e-07 $l=2.41454e-07 $layer=licon1_NDIFF $count=1 $X=1.64
+ $Y=0.6 $X2=1.86 $Y2=0.645
.ends

