* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__or4b_2 A B C D_N VGND VNB VPB VPWR X
X0 X a_190_48# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X1 VPWR a_190_48# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X2 VGND C a_190_48# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X3 a_27_368# D_N VGND VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X4 VGND A a_190_48# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X5 a_27_368# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X6 a_452_392# B a_536_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 VPWR A a_452_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 X a_190_48# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X9 a_638_392# a_27_368# a_190_48# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_190_48# a_27_368# VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X11 a_536_392# C a_638_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 VGND a_190_48# X VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X13 a_190_48# B VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
.ends
