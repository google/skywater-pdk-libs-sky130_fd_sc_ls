* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__dlclkp_1 CLK GATE VGND VNB VPB VPWR GCLK
M1000 GCLK a_987_393# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=1.88295e+12p ps=1.214e+07u
M1001 a_477_124# a_309_338# a_83_260# VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=2.692e+11p ps=2.3e+06u
M1002 VGND CLK a_315_54# VNB nshort w=740000u l=150000u
+  ad=1.19302e+12p pd=9.54e+06u as=2.183e+11p ps=2.07e+06u
M1003 a_309_338# a_315_54# VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1004 VPWR CLK a_315_54# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=2.478e+11p ps=2.27e+06u
M1005 VPWR a_27_74# a_484_508# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1006 a_484_508# a_315_54# a_83_260# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=3.889e+11p ps=3.12e+06u
M1007 VPWR a_27_74# a_987_393# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=2.604e+11p ps=2.3e+06u
M1008 a_987_393# a_27_74# a_984_125# VNB nshort w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=1.536e+11p ps=1.76e+06u
M1009 a_987_393# CLK VPWR VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR a_83_260# a_27_74# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.304e+11p ps=2.83e+06u
M1011 a_984_125# CLK VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 GCLK a_987_393# VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1013 a_83_260# a_309_338# a_258_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1014 VGND a_27_74# a_477_124# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND a_83_260# a_27_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1016 a_309_338# a_315_54# VPWR VPB phighvt w=840000u l=150000u
+  ad=2.478e+11p pd=2.27e+06u as=0p ps=0u
M1017 a_258_392# GATE VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_267_80# GATE VGND VNB nshort w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1019 a_83_260# a_315_54# a_267_80# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
