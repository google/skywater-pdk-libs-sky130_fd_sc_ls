# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_ls__o311ai_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.04000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.165000 1.350000 10.435000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.765000 1.350000 7.775000 1.780000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.485000 1.430000 6.195000 1.640000 ;
        RECT 5.185000 1.640000 6.195000 1.780000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.780000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.245000 1.430000 4.195000 1.780000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.780000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.300000 1.240000 1.780000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  2.271700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545000 0.770000 1.740000 1.090000 ;
        RECT 0.545000 1.090000 6.595000 1.100000 ;
        RECT 0.740000 1.950000 6.595000 2.120000 ;
        RECT 0.740000 2.120000 1.070000 2.980000 ;
        RECT 1.410000 1.100000 6.595000 1.260000 ;
        RECT 1.740000 1.820000 2.070000 1.950000 ;
        RECT 1.740000 2.120000 2.070000 2.980000 ;
        RECT 4.685000 1.820000 5.015000 1.950000 ;
        RECT 4.685000 2.120000 5.015000 2.735000 ;
        RECT 5.685000 2.120000 6.015000 2.735000 ;
        RECT 6.365000 1.260000 6.595000 1.950000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 11.040000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 11.040000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.040000 0.085000 ;
      RECT  0.000000  3.245000 11.040000 3.415000 ;
      RECT  0.115000  0.350000  2.090000 0.600000 ;
      RECT  0.115000  0.600000  0.365000 1.130000 ;
      RECT  0.115000  1.950000  0.445000 3.245000 ;
      RECT  1.240000  2.290000  1.570000 3.245000 ;
      RECT  1.920000  0.600000  2.090000 0.750000 ;
      RECT  1.920000  0.750000  3.900000 0.920000 ;
      RECT  2.240000  2.290000  3.905000 3.245000 ;
      RECT  2.270000  0.330000  4.240000 0.580000 ;
      RECT  4.070000  0.580000  4.240000 0.750000 ;
      RECT  4.070000  0.750000  7.140000 0.920000 ;
      RECT  4.185000  2.290000  4.515000 2.905000 ;
      RECT  4.185000  2.905000  8.565000 3.075000 ;
      RECT  4.410000  0.085000  4.740000 0.580000 ;
      RECT  4.920000  0.350000  5.170000 0.750000 ;
      RECT  5.185000  2.290000  5.515000 2.905000 ;
      RECT  5.350000  0.085000  5.680000 0.580000 ;
      RECT  5.860000  0.350000  6.190000 0.750000 ;
      RECT  6.285000  2.290000  6.615000 2.905000 ;
      RECT  6.370000  0.085000  6.710000 0.580000 ;
      RECT  6.785000  1.950000 10.475000 2.120000 ;
      RECT  6.785000  2.120000  7.115000 2.735000 ;
      RECT  6.890000  0.350000  7.140000 0.750000 ;
      RECT  6.890000  0.920000  7.140000 1.010000 ;
      RECT  6.890000  1.010000  8.115000 1.180000 ;
      RECT  7.285000  2.290000  7.615000 2.905000 ;
      RECT  7.320000  0.085000  7.650000 0.825000 ;
      RECT  7.785000  2.120000 10.475000 2.150000 ;
      RECT  7.785000  2.150000  8.065000 2.735000 ;
      RECT  7.945000  0.350000  8.115000 1.010000 ;
      RECT  7.945000  1.180000  8.115000 1.300000 ;
      RECT  7.945000  1.300000  8.975000 1.470000 ;
      RECT  8.235000  2.330000  8.565000 2.905000 ;
      RECT  8.295000  0.085000  8.545000 1.130000 ;
      RECT  8.725000  0.350000  8.975000 0.960000 ;
      RECT  8.725000  0.960000 10.415000 1.130000 ;
      RECT  8.725000  1.130000  8.975000 1.300000 ;
      RECT  8.795000  2.330000  9.125000 3.245000 ;
      RECT  9.155000  0.085000  9.995000 0.790000 ;
      RECT  9.295000  2.150000  9.525000 2.980000 ;
      RECT  9.695000  2.330000 10.025000 3.245000 ;
      RECT 10.165000  0.350000 10.415000 0.960000 ;
      RECT 10.195000  2.150000 10.475000 2.980000 ;
      RECT 10.595000  0.085000 10.925000 1.130000 ;
      RECT 10.675000  1.820000 10.925000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
  END
END sky130_fd_sc_ls__o311ai_4
END LIBRARY
