* File: sky130_fd_sc_ls__dfxtp_4.pxi.spice
* Created: Fri Aug 28 13:16:55 2020
* 
x_PM_SKY130_FD_SC_LS__DFXTP_4%CLK N_CLK_M1025_g N_CLK_c_214_n N_CLK_M1015_g CLK
+ N_CLK_c_215_n PM_SKY130_FD_SC_LS__DFXTP_4%CLK
x_PM_SKY130_FD_SC_LS__DFXTP_4%A_27_74# N_A_27_74#_M1025_s N_A_27_74#_M1015_s
+ N_A_27_74#_c_246_n N_A_27_74#_M1016_g N_A_27_74#_c_247_n N_A_27_74#_M1022_g
+ N_A_27_74#_M1020_g N_A_27_74#_c_272_n N_A_27_74#_c_273_n N_A_27_74#_M1006_g
+ N_A_27_74#_c_274_n N_A_27_74#_M1018_g N_A_27_74#_c_275_n N_A_27_74#_M1028_g
+ N_A_27_74#_c_249_n N_A_27_74#_c_250_n N_A_27_74#_c_251_n N_A_27_74#_c_277_n
+ N_A_27_74#_c_278_n N_A_27_74#_c_252_n N_A_27_74#_c_253_n N_A_27_74#_c_298_n
+ N_A_27_74#_c_254_n N_A_27_74#_c_255_n N_A_27_74#_c_256_n N_A_27_74#_c_257_n
+ N_A_27_74#_c_258_n N_A_27_74#_c_259_n N_A_27_74#_c_260_n N_A_27_74#_c_261_n
+ N_A_27_74#_c_262_n N_A_27_74#_c_280_n N_A_27_74#_c_281_n N_A_27_74#_c_263_n
+ N_A_27_74#_c_264_n N_A_27_74#_c_385_p N_A_27_74#_c_386_p N_A_27_74#_c_265_n
+ N_A_27_74#_c_266_n N_A_27_74#_c_304_n N_A_27_74#_c_267_n N_A_27_74#_c_268_n
+ N_A_27_74#_c_269_n N_A_27_74#_c_270_n PM_SKY130_FD_SC_LS__DFXTP_4%A_27_74#
x_PM_SKY130_FD_SC_LS__DFXTP_4%D N_D_c_521_n N_D_M1008_g N_D_c_516_n N_D_c_517_n
+ N_D_M1019_g N_D_c_522_n N_D_c_523_n D D N_D_c_519_n D
+ PM_SKY130_FD_SC_LS__DFXTP_4%D
x_PM_SKY130_FD_SC_LS__DFXTP_4%A_206_368# N_A_206_368#_M1022_d
+ N_A_206_368#_M1016_d N_A_206_368#_c_577_n N_A_206_368#_c_578_n
+ N_A_206_368#_c_579_n N_A_206_368#_c_589_n N_A_206_368#_c_590_n
+ N_A_206_368#_c_591_n N_A_206_368#_M1010_g N_A_206_368#_M1017_g
+ N_A_206_368#_c_581_n N_A_206_368#_M1021_g N_A_206_368#_c_592_n
+ N_A_206_368#_M1001_g N_A_206_368#_c_593_n N_A_206_368#_c_582_n
+ N_A_206_368#_c_594_n N_A_206_368#_c_682_n N_A_206_368#_c_595_n
+ N_A_206_368#_c_596_n N_A_206_368#_c_643_n N_A_206_368#_c_697_p
+ N_A_206_368#_c_644_n N_A_206_368#_c_698_p N_A_206_368#_c_597_n
+ N_A_206_368#_c_598_n N_A_206_368#_c_583_n N_A_206_368#_c_584_n
+ N_A_206_368#_c_600_n N_A_206_368#_c_601_n N_A_206_368#_c_602_n
+ N_A_206_368#_c_585_n N_A_206_368#_c_604_n N_A_206_368#_c_586_n
+ N_A_206_368#_c_587_n N_A_206_368#_c_588_n N_A_206_368#_c_606_n
+ PM_SKY130_FD_SC_LS__DFXTP_4%A_206_368#
x_PM_SKY130_FD_SC_LS__DFXTP_4%A_696_458# N_A_696_458#_M1005_d
+ N_A_696_458#_M1027_d N_A_696_458#_c_826_n N_A_696_458#_M1009_g
+ N_A_696_458#_c_819_n N_A_696_458#_c_820_n N_A_696_458#_c_821_n
+ N_A_696_458#_M1011_g N_A_696_458#_c_828_n N_A_696_458#_c_822_n
+ N_A_696_458#_c_823_n N_A_696_458#_c_824_n N_A_696_458#_c_825_n
+ PM_SKY130_FD_SC_LS__DFXTP_4%A_696_458#
x_PM_SKY130_FD_SC_LS__DFXTP_4%A_544_485# N_A_544_485#_M1020_d
+ N_A_544_485#_M1010_d N_A_544_485#_c_913_n N_A_544_485#_M1027_g
+ N_A_544_485#_c_903_n N_A_544_485#_M1005_g N_A_544_485#_c_905_n
+ N_A_544_485#_c_906_n N_A_544_485#_c_907_n N_A_544_485#_c_908_n
+ N_A_544_485#_c_915_n N_A_544_485#_c_909_n N_A_544_485#_c_910_n
+ N_A_544_485#_c_917_n N_A_544_485#_c_911_n N_A_544_485#_c_912_n
+ PM_SKY130_FD_SC_LS__DFXTP_4%A_544_485#
x_PM_SKY130_FD_SC_LS__DFXTP_4%A_1226_296# N_A_1226_296#_M1024_s
+ N_A_1226_296#_M1003_s N_A_1226_296#_c_1026_n N_A_1226_296#_c_1027_n
+ N_A_1226_296#_M1023_g N_A_1226_296#_M1014_g N_A_1226_296#_M1000_g
+ N_A_1226_296#_c_1028_n N_A_1226_296#_M1002_g N_A_1226_296#_c_1029_n
+ N_A_1226_296#_M1007_g N_A_1226_296#_M1004_g N_A_1226_296#_c_1030_n
+ N_A_1226_296#_M1013_g N_A_1226_296#_M1012_g N_A_1226_296#_M1030_g
+ N_A_1226_296#_c_1031_n N_A_1226_296#_M1026_g N_A_1226_296#_c_1032_n
+ N_A_1226_296#_c_1033_n N_A_1226_296#_c_1018_n N_A_1226_296#_c_1019_n
+ N_A_1226_296#_c_1020_n N_A_1226_296#_c_1021_n N_A_1226_296#_c_1022_n
+ N_A_1226_296#_c_1023_n N_A_1226_296#_c_1024_n N_A_1226_296#_c_1025_n
+ PM_SKY130_FD_SC_LS__DFXTP_4%A_1226_296#
x_PM_SKY130_FD_SC_LS__DFXTP_4%A_1034_424# N_A_1034_424#_M1021_d
+ N_A_1034_424#_M1018_d N_A_1034_424#_c_1188_n N_A_1034_424#_M1003_g
+ N_A_1034_424#_c_1181_n N_A_1034_424#_c_1190_n N_A_1034_424#_c_1191_n
+ N_A_1034_424#_c_1192_n N_A_1034_424#_M1029_g N_A_1034_424#_c_1182_n
+ N_A_1034_424#_M1024_g N_A_1034_424#_c_1193_n N_A_1034_424#_c_1198_n
+ N_A_1034_424#_c_1194_n N_A_1034_424#_c_1195_n N_A_1034_424#_c_1183_n
+ N_A_1034_424#_c_1184_n N_A_1034_424#_c_1185_n N_A_1034_424#_c_1186_n
+ N_A_1034_424#_c_1187_n PM_SKY130_FD_SC_LS__DFXTP_4%A_1034_424#
x_PM_SKY130_FD_SC_LS__DFXTP_4%VPWR N_VPWR_M1015_d N_VPWR_M1008_s N_VPWR_M1009_d
+ N_VPWR_M1023_d N_VPWR_M1029_d N_VPWR_M1007_s N_VPWR_M1026_s N_VPWR_c_1288_n
+ N_VPWR_c_1289_n N_VPWR_c_1290_n N_VPWR_c_1291_n N_VPWR_c_1292_n
+ N_VPWR_c_1293_n N_VPWR_c_1294_n N_VPWR_c_1295_n N_VPWR_c_1296_n
+ N_VPWR_c_1297_n N_VPWR_c_1298_n VPWR N_VPWR_c_1299_n N_VPWR_c_1300_n
+ N_VPWR_c_1301_n N_VPWR_c_1302_n N_VPWR_c_1303_n N_VPWR_c_1304_n
+ N_VPWR_c_1305_n N_VPWR_c_1306_n N_VPWR_c_1287_n
+ PM_SKY130_FD_SC_LS__DFXTP_4%VPWR
x_PM_SKY130_FD_SC_LS__DFXTP_4%A_437_503# N_A_437_503#_M1019_d
+ N_A_437_503#_M1008_d N_A_437_503#_c_1417_n N_A_437_503#_c_1413_n
+ N_A_437_503#_c_1414_n N_A_437_503#_c_1415_n N_A_437_503#_c_1416_n
+ N_A_437_503#_c_1419_n PM_SKY130_FD_SC_LS__DFXTP_4%A_437_503#
x_PM_SKY130_FD_SC_LS__DFXTP_4%Q N_Q_M1000_d N_Q_M1012_d N_Q_M1002_d N_Q_M1013_d
+ N_Q_c_1474_n N_Q_c_1468_n N_Q_c_1475_n N_Q_c_1476_n N_Q_c_1469_n N_Q_c_1470_n
+ N_Q_c_1471_n N_Q_c_1472_n N_Q_c_1473_n Q Q Q Q PM_SKY130_FD_SC_LS__DFXTP_4%Q
x_PM_SKY130_FD_SC_LS__DFXTP_4%VGND N_VGND_M1025_d N_VGND_M1019_s N_VGND_M1011_d
+ N_VGND_M1014_d N_VGND_M1024_d N_VGND_M1004_s N_VGND_M1030_s N_VGND_c_1548_n
+ N_VGND_c_1549_n N_VGND_c_1550_n N_VGND_c_1551_n N_VGND_c_1552_n
+ N_VGND_c_1553_n N_VGND_c_1554_n N_VGND_c_1555_n N_VGND_c_1556_n
+ N_VGND_c_1557_n N_VGND_c_1558_n VGND N_VGND_c_1559_n N_VGND_c_1560_n
+ N_VGND_c_1561_n N_VGND_c_1562_n N_VGND_c_1563_n N_VGND_c_1564_n
+ N_VGND_c_1565_n N_VGND_c_1566_n N_VGND_c_1567_n N_VGND_c_1568_n
+ N_VGND_c_1569_n PM_SKY130_FD_SC_LS__DFXTP_4%VGND
cc_1 VNB N_CLK_M1025_g 0.0314862f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_CLK_c_214_n 0.0463134f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_3 VNB N_CLK_c_215_n 0.0163894f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=1.465
cc_4 VNB N_A_27_74#_c_246_n 0.0429298f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_5 VNB N_A_27_74#_c_247_n 0.0185497f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.465
cc_6 VNB N_A_27_74#_M1028_g 0.0383567f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_27_74#_c_249_n 0.0137015f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_27_74#_c_250_n 0.0115034f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_27_74#_c_251_n 0.02581f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_27_74#_c_252_n 0.003029f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_27_74#_c_253_n 0.00924841f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_74#_c_254_n 0.00152687f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_74#_c_255_n 0.0075881f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_74#_c_256_n 0.00137942f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_74#_c_257_n 0.00380045f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_27_74#_c_258_n 0.00734633f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_27_74#_c_259_n 0.00202332f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_27_74#_c_260_n 0.00310292f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_27_74#_c_261_n 0.0213909f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_27_74#_c_262_n 0.00177503f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_27_74#_c_263_n 0.00132271f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_27_74#_c_264_n 0.0128181f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_27_74#_c_265_n 0.00240889f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_27_74#_c_266_n 0.00509724f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_27_74#_c_267_n 0.00435855f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_27_74#_c_268_n 0.0456888f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_27_74#_c_269_n 0.0117318f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_27_74#_c_270_n 0.0261733f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_D_c_516_n 0.0287455f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_D_c_517_n 0.018154f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_31 VNB D 0.00849691f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_D_c_519_n 0.0320047f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB D 0.00141546f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_206_368#_c_577_n 0.0649996f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_35 VNB N_A_206_368#_c_578_n 0.135383f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_206_368#_c_579_n 0.0124288f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.465
cc_37 VNB N_A_206_368#_M1017_g 0.0293998f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_206_368#_c_581_n 0.0177425f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_206_368#_c_582_n 0.00196407f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_206_368#_c_583_n 0.0134612f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_206_368#_c_584_n 0.00222883f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_206_368#_c_585_n 0.00229328f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_206_368#_c_586_n 0.00506519f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_206_368#_c_587_n 0.0424638f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_206_368#_c_588_n 0.0325476f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_696_458#_c_819_n 0.0362452f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.465
cc_47 VNB N_A_696_458#_c_820_n 0.0160506f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=1.465
cc_48 VNB N_A_696_458#_c_821_n 0.0188985f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=1.465
cc_49 VNB N_A_696_458#_c_822_n 0.00675562f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_696_458#_c_823_n 0.032964f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_696_458#_c_824_n 0.00744237f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_696_458#_c_825_n 0.00785424f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_544_485#_c_903_n 0.0118371f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=1.465
cc_54 VNB N_A_544_485#_M1005_g 0.0326438f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_544_485#_c_905_n 0.0147249f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_544_485#_c_906_n 0.00170751f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_544_485#_c_907_n 0.00606768f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_544_485#_c_908_n 0.003624f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_544_485#_c_909_n 0.00355519f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_544_485#_c_910_n 0.00245988f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_544_485#_c_911_n 0.00279514f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_544_485#_c_912_n 0.0140793f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_1226_296#_M1014_g 0.0396395f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_1226_296#_M1000_g 0.0225597f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_1226_296#_M1004_g 0.0216914f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_1226_296#_M1012_g 0.0211596f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_1226_296#_M1030_g 0.0260204f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_1226_296#_c_1018_n 9.43046e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_1226_296#_c_1019_n 0.00737701f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_1226_296#_c_1020_n 0.0017939f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_1226_296#_c_1021_n 0.00343836f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_1226_296#_c_1022_n 0.00679267f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_1226_296#_c_1023_n 0.00490241f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_1226_296#_c_1024_n 0.0163456f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_1226_296#_c_1025_n 0.116715f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_1034_424#_c_1181_n 0.00737859f $X=-0.19 $Y=-0.245 $X2=0.34
+ $Y2=1.465
cc_77 VNB N_A_1034_424#_c_1182_n 0.0192903f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_1034_424#_c_1183_n 0.00110384f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_1034_424#_c_1184_n 0.00350916f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_1034_424#_c_1185_n 0.0432948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_1034_424#_c_1186_n 0.00109692f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_1034_424#_c_1187_n 0.0462154f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_VPWR_c_1287_n 0.40251f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_437_503#_c_1413_n 0.0063043f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=1.465
cc_85 VNB N_A_437_503#_c_1414_n 0.00537792f $X=-0.19 $Y=-0.245 $X2=0.315
+ $Y2=1.465
cc_86 VNB N_A_437_503#_c_1415_n 0.00352716f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_437_503#_c_1416_n 0.00186489f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_Q_c_1468_n 0.00280874f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_Q_c_1469_n 0.00237452f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_Q_c_1470_n 0.00260202f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_Q_c_1471_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_Q_c_1472_n 0.00159092f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_Q_c_1473_n 0.00181295f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_VGND_c_1548_n 0.00772186f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_VGND_c_1549_n 0.0035883f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_VGND_c_1550_n 0.00683089f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_VGND_c_1551_n 0.0185708f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_VGND_c_1552_n 0.00590547f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_VGND_c_1553_n 0.0189618f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_VGND_c_1554_n 0.00798328f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_VGND_c_1555_n 0.0114755f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_VGND_c_1556_n 0.0505702f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_VGND_c_1557_n 0.0406885f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_VGND_c_1558_n 0.00477982f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_VGND_c_1559_n 0.0194697f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_VGND_c_1560_n 0.027872f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_VGND_c_1561_n 0.0508339f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_VGND_c_1562_n 0.0188435f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_VGND_c_1563_n 0.0199286f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_1564_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_1565_n 0.0043669f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_1566_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_1567_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_1568_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_VGND_c_1569_n 0.519401f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VPB N_CLK_c_214_n 0.0289619f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_117 VPB N_CLK_c_215_n 0.0073823f $X=-0.19 $Y=1.66 $X2=0.34 $Y2=1.465
cc_118 VPB N_A_27_74#_c_246_n 0.0262962f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_119 VPB N_A_27_74#_c_272_n 0.0157713f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_A_27_74#_c_273_n 0.0204072f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_A_27_74#_c_274_n 0.0381502f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_A_27_74#_c_275_n 0.0435717f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_A_27_74#_M1028_g 0.0017983f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_A_27_74#_c_277_n 0.00758177f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_A_27_74#_c_278_n 0.035396f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 VPB N_A_27_74#_c_254_n 0.00309553f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_127 VPB N_A_27_74#_c_280_n 0.00843859f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_A_27_74#_c_281_n 0.0393075f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_129 VPB N_A_27_74#_c_264_n 5.46431e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_A_27_74#_c_270_n 0.0056647f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_D_c_521_n 0.0673339f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.3
cc_132 VPB N_D_c_522_n 0.00388284f $X=-0.19 $Y=1.66 $X2=0.34 $Y2=1.465
cc_133 VPB N_D_c_523_n 0.00469496f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_A_206_368#_c_589_n 0.0606794f $X=-0.19 $Y=1.66 $X2=0.34 $Y2=1.465
cc_135 VPB N_A_206_368#_c_590_n 0.026359f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_A_206_368#_c_591_n 0.02225f $X=-0.19 $Y=1.66 $X2=0.315 $Y2=1.665
cc_137 VPB N_A_206_368#_c_592_n 0.0624586f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_A_206_368#_c_593_n 0.00763125f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_A_206_368#_c_594_n 0.00678494f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_140 VPB N_A_206_368#_c_595_n 0.0135182f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_141 VPB N_A_206_368#_c_596_n 0.00253834f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_142 VPB N_A_206_368#_c_597_n 0.00359332f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_143 VPB N_A_206_368#_c_598_n 0.00179303f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_144 VPB N_A_206_368#_c_584_n 0.003244f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_145 VPB N_A_206_368#_c_600_n 0.00590845f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_146 VPB N_A_206_368#_c_601_n 0.00589917f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_147 VPB N_A_206_368#_c_602_n 0.0105025f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_148 VPB N_A_206_368#_c_585_n 0.00331166f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_149 VPB N_A_206_368#_c_604_n 0.00934484f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_150 VPB N_A_206_368#_c_587_n 0.0151905f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_151 VPB N_A_206_368#_c_606_n 9.0268e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_152 VPB N_A_696_458#_c_826_n 0.0168873f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_153 VPB N_A_696_458#_c_820_n 0.0310025f $X=-0.19 $Y=1.66 $X2=0.34 $Y2=1.465
cc_154 VPB N_A_696_458#_c_828_n 0.0219817f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_155 VPB N_A_696_458#_c_825_n 0.00194788f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_156 VPB N_A_544_485#_c_913_n 0.0176636f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_157 VPB N_A_544_485#_c_906_n 0.0105463f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_158 VPB N_A_544_485#_c_915_n 0.0155691f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_159 VPB N_A_544_485#_c_910_n 0.00263683f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_160 VPB N_A_544_485#_c_917_n 0.00317002f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_161 VPB N_A_544_485#_c_912_n 0.0574354f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_162 VPB N_A_1226_296#_c_1026_n 0.0375518f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_163 VPB N_A_1226_296#_c_1027_n 0.02338f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_164 VPB N_A_1226_296#_c_1028_n 0.0168783f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_165 VPB N_A_1226_296#_c_1029_n 0.0152465f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_166 VPB N_A_1226_296#_c_1030_n 0.015247f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_167 VPB N_A_1226_296#_c_1031_n 0.0174208f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_168 VPB N_A_1226_296#_c_1032_n 0.00902049f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_169 VPB N_A_1226_296#_c_1033_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_170 VPB N_A_1226_296#_c_1021_n 0.0101625f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_171 VPB N_A_1226_296#_c_1023_n 0.00492717f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_172 VPB N_A_1226_296#_c_1024_n 0.0136225f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_173 VPB N_A_1226_296#_c_1025_n 0.0303748f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_174 VPB N_A_1034_424#_c_1188_n 0.0159638f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_175 VPB N_A_1034_424#_c_1181_n 0.0139419f $X=-0.19 $Y=1.66 $X2=0.34 $Y2=1.465
cc_176 VPB N_A_1034_424#_c_1190_n 0.0192857f $X=-0.19 $Y=1.66 $X2=0.34 $Y2=1.465
cc_177 VPB N_A_1034_424#_c_1191_n 0.0123081f $X=-0.19 $Y=1.66 $X2=0.315
+ $Y2=1.465
cc_178 VPB N_A_1034_424#_c_1192_n 0.0161605f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_179 VPB N_A_1034_424#_c_1193_n 0.00823029f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_180 VPB N_A_1034_424#_c_1194_n 0.00721074f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_181 VPB N_A_1034_424#_c_1195_n 2.36146e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_182 VPB N_A_1034_424#_c_1184_n 4.86372e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_183 VPB N_VPWR_c_1288_n 0.00799266f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_184 VPB N_VPWR_c_1289_n 0.0222809f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_185 VPB N_VPWR_c_1290_n 0.00219572f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_186 VPB N_VPWR_c_1291_n 0.00750325f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_187 VPB N_VPWR_c_1292_n 0.0095345f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_188 VPB N_VPWR_c_1293_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_189 VPB N_VPWR_c_1294_n 0.00799266f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_190 VPB N_VPWR_c_1295_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_191 VPB N_VPWR_c_1296_n 0.0645754f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_192 VPB N_VPWR_c_1297_n 0.0121247f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_193 VPB N_VPWR_c_1298_n 0.0446788f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_194 VPB N_VPWR_c_1299_n 0.0543314f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_195 VPB N_VPWR_c_1300_n 0.0198086f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_196 VPB N_VPWR_c_1301_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_197 VPB N_VPWR_c_1302_n 0.0233502f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_198 VPB N_VPWR_c_1303_n 0.00324035f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_199 VPB N_VPWR_c_1304_n 0.00623744f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_200 VPB N_VPWR_c_1305_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_201 VPB N_VPWR_c_1306_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_202 VPB N_VPWR_c_1287_n 0.116556f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_203 VPB N_A_437_503#_c_1417_n 0.00567555f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_204 VPB N_A_437_503#_c_1413_n 0.00181594f $X=-0.19 $Y=1.66 $X2=0.34 $Y2=1.465
cc_205 VPB N_A_437_503#_c_1419_n 0.00519997f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_206 VPB N_Q_c_1474_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0.315 $Y2=1.665
cc_207 VPB N_Q_c_1475_n 0.00179527f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_208 VPB N_Q_c_1476_n 0.00183475f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_209 VPB N_Q_c_1472_n 8.42804e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_210 VPB Q 0.00130942f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_211 VPB Q 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_212 N_CLK_M1025_g N_A_27_74#_c_246_n 0.0040438f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_213 N_CLK_c_214_n N_A_27_74#_c_246_n 0.0455539f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_214 N_CLK_c_215_n N_A_27_74#_c_246_n 2.10754e-19 $X=0.34 $Y=1.465 $X2=0 $Y2=0
cc_215 N_CLK_M1025_g N_A_27_74#_c_247_n 0.0156678f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_216 N_CLK_M1025_g N_A_27_74#_c_251_n 0.0095711f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_217 N_CLK_c_214_n N_A_27_74#_c_277_n 0.0016558f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_218 N_CLK_c_215_n N_A_27_74#_c_277_n 0.0258609f $X=0.34 $Y=1.465 $X2=0 $Y2=0
cc_219 N_CLK_c_214_n N_A_27_74#_c_278_n 0.0104891f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_220 N_CLK_M1025_g N_A_27_74#_c_252_n 0.0128375f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_221 N_CLK_c_214_n N_A_27_74#_c_252_n 0.00100324f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_222 N_CLK_c_215_n N_A_27_74#_c_252_n 0.00433199f $X=0.34 $Y=1.465 $X2=0 $Y2=0
cc_223 N_CLK_M1025_g N_A_27_74#_c_253_n 0.00113124f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_224 N_CLK_c_214_n N_A_27_74#_c_253_n 0.0019389f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_225 N_CLK_c_215_n N_A_27_74#_c_253_n 0.0278432f $X=0.34 $Y=1.465 $X2=0 $Y2=0
cc_226 N_CLK_c_214_n N_A_27_74#_c_298_n 0.0139121f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_227 N_CLK_c_215_n N_A_27_74#_c_298_n 0.00433199f $X=0.34 $Y=1.465 $X2=0 $Y2=0
cc_228 N_CLK_c_214_n N_A_27_74#_c_254_n 0.00397589f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_229 N_CLK_M1025_g N_A_27_74#_c_266_n 0.00516055f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_230 N_CLK_c_214_n N_A_27_74#_c_266_n 0.00330504f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_231 N_CLK_c_215_n N_A_27_74#_c_266_n 0.0379192f $X=0.34 $Y=1.465 $X2=0 $Y2=0
cc_232 N_CLK_M1025_g N_A_27_74#_c_304_n 0.00177892f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_233 N_CLK_c_214_n N_A_206_368#_c_593_n 6.45668e-19 $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_234 N_CLK_c_214_n N_VPWR_c_1288_n 0.00486623f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_235 N_CLK_c_214_n N_VPWR_c_1302_n 0.00445602f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_236 N_CLK_c_214_n N_VPWR_c_1287_n 0.00861168f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_237 N_CLK_M1025_g N_VGND_c_1548_n 0.00325137f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_238 N_CLK_M1025_g N_VGND_c_1559_n 0.00434272f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_239 N_CLK_M1025_g N_VGND_c_1569_n 0.00825573f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_240 N_A_27_74#_c_250_n N_D_c_516_n 0.00789174f $X=3.145 $Y=1.24 $X2=0 $Y2=0
cc_241 N_A_27_74#_c_258_n N_D_c_516_n 8.26575e-19 $X=2.485 $Y=0.815 $X2=0 $Y2=0
cc_242 N_A_27_74#_c_270_n N_D_c_516_n 0.00133719f $X=3.287 $Y=1.75 $X2=0 $Y2=0
cc_243 N_A_27_74#_c_249_n N_D_c_517_n 0.00789174f $X=3.145 $Y=1.09 $X2=0 $Y2=0
cc_244 N_A_27_74#_c_258_n N_D_c_517_n 0.00642909f $X=2.485 $Y=0.815 $X2=0 $Y2=0
cc_245 N_A_27_74#_c_260_n N_D_c_517_n 0.00859213f $X=2.57 $Y=0.73 $X2=0 $Y2=0
cc_246 N_A_27_74#_c_261_n N_D_c_517_n 0.00155847f $X=3.705 $Y=0.34 $X2=0 $Y2=0
cc_247 N_A_27_74#_c_258_n D 0.0228259f $X=2.485 $Y=0.815 $X2=0 $Y2=0
cc_248 N_A_27_74#_c_258_n N_D_c_519_n 0.00769114f $X=2.485 $Y=0.815 $X2=0 $Y2=0
cc_249 N_A_27_74#_c_255_n N_A_206_368#_M1022_d 0.0063531f $X=1.645 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_250 N_A_27_74#_c_255_n N_A_206_368#_c_577_n 0.00779381f $X=1.645 $Y=0.34
+ $X2=0 $Y2=0
cc_251 N_A_27_74#_c_257_n N_A_206_368#_c_577_n 0.0108388f $X=1.73 $Y=0.73 $X2=0
+ $Y2=0
cc_252 N_A_27_74#_c_259_n N_A_206_368#_c_577_n 0.00938601f $X=1.815 $Y=0.815
+ $X2=0 $Y2=0
cc_253 N_A_27_74#_c_304_n N_A_206_368#_c_577_n 7.1833e-19 $X=0.905 $Y=0.96 $X2=0
+ $Y2=0
cc_254 N_A_27_74#_c_249_n N_A_206_368#_c_578_n 0.00882199f $X=3.145 $Y=1.09
+ $X2=0 $Y2=0
cc_255 N_A_27_74#_c_255_n N_A_206_368#_c_578_n 4.19731e-19 $X=1.645 $Y=0.34
+ $X2=0 $Y2=0
cc_256 N_A_27_74#_c_258_n N_A_206_368#_c_578_n 0.0061518f $X=2.485 $Y=0.815
+ $X2=0 $Y2=0
cc_257 N_A_27_74#_c_261_n N_A_206_368#_c_578_n 0.013889f $X=3.705 $Y=0.34 $X2=0
+ $Y2=0
cc_258 N_A_27_74#_c_262_n N_A_206_368#_c_578_n 0.0035998f $X=2.655 $Y=0.34 $X2=0
+ $Y2=0
cc_259 N_A_27_74#_c_247_n N_A_206_368#_c_579_n 0.0173557f $X=1.12 $Y=1.22 $X2=0
+ $Y2=0
cc_260 N_A_27_74#_c_255_n N_A_206_368#_c_579_n 0.00102791f $X=1.645 $Y=0.34
+ $X2=0 $Y2=0
cc_261 N_A_27_74#_c_270_n N_A_206_368#_c_589_n 0.00649057f $X=3.287 $Y=1.75
+ $X2=0 $Y2=0
cc_262 N_A_27_74#_c_281_n N_A_206_368#_c_590_n 0.00597913f $X=3.32 $Y=1.915
+ $X2=0 $Y2=0
cc_263 N_A_27_74#_c_272_n N_A_206_368#_c_591_n 0.00597913f $X=3.18 $Y=2.35 $X2=0
+ $Y2=0
cc_264 N_A_27_74#_c_273_n N_A_206_368#_c_591_n 0.0118532f $X=3.18 $Y=2.44 $X2=0
+ $Y2=0
cc_265 N_A_27_74#_c_249_n N_A_206_368#_M1017_g 0.00850711f $X=3.145 $Y=1.09
+ $X2=0 $Y2=0
cc_266 N_A_27_74#_c_261_n N_A_206_368#_M1017_g 0.0164125f $X=3.705 $Y=0.34 $X2=0
+ $Y2=0
cc_267 N_A_27_74#_c_280_n N_A_206_368#_M1017_g 0.00389871f $X=3.705 $Y=1.915
+ $X2=0 $Y2=0
cc_268 N_A_27_74#_c_263_n N_A_206_368#_M1017_g 0.00258579f $X=3.79 $Y=0.69 $X2=0
+ $Y2=0
cc_269 N_A_27_74#_c_264_n N_A_206_368#_M1017_g 0.00138295f $X=3.79 $Y=1.75 $X2=0
+ $Y2=0
cc_270 N_A_27_74#_M1028_g N_A_206_368#_c_581_n 0.0113184f $X=5.815 $Y=0.83 $X2=0
+ $Y2=0
cc_271 N_A_27_74#_c_267_n N_A_206_368#_c_581_n 4.97101e-19 $X=5.83 $Y=0.345
+ $X2=0 $Y2=0
cc_272 N_A_27_74#_c_268_n N_A_206_368#_c_581_n 0.00468991f $X=5.83 $Y=0.345
+ $X2=0 $Y2=0
cc_273 N_A_27_74#_c_269_n N_A_206_368#_c_581_n 0.0109765f $X=5.665 $Y=0.382
+ $X2=0 $Y2=0
cc_274 N_A_27_74#_c_274_n N_A_206_368#_c_592_n 0.0221474f $X=5.095 $Y=2.045
+ $X2=0 $Y2=0
cc_275 N_A_27_74#_c_275_n N_A_206_368#_c_592_n 0.0228077f $X=5.74 $Y=1.765 $X2=0
+ $Y2=0
cc_276 N_A_27_74#_c_246_n N_A_206_368#_c_593_n 0.00654713f $X=0.955 $Y=1.765
+ $X2=0 $Y2=0
cc_277 N_A_27_74#_c_278_n N_A_206_368#_c_593_n 0.00481788f $X=0.28 $Y=2.815
+ $X2=0 $Y2=0
cc_278 N_A_27_74#_c_247_n N_A_206_368#_c_582_n 0.00279715f $X=1.12 $Y=1.22 $X2=0
+ $Y2=0
cc_279 N_A_27_74#_c_255_n N_A_206_368#_c_582_n 0.0127042f $X=1.645 $Y=0.34 $X2=0
+ $Y2=0
cc_280 N_A_27_74#_c_257_n N_A_206_368#_c_582_n 0.00944377f $X=1.73 $Y=0.73 $X2=0
+ $Y2=0
cc_281 N_A_27_74#_c_259_n N_A_206_368#_c_582_n 0.0133618f $X=1.815 $Y=0.815
+ $X2=0 $Y2=0
cc_282 N_A_27_74#_c_304_n N_A_206_368#_c_582_n 0.0454018f $X=0.905 $Y=0.96 $X2=0
+ $Y2=0
cc_283 N_A_27_74#_c_273_n N_A_206_368#_c_595_n 0.0108338f $X=3.18 $Y=2.44 $X2=0
+ $Y2=0
cc_284 N_A_27_74#_c_273_n N_A_206_368#_c_643_n 0.00373658f $X=3.18 $Y=2.44 $X2=0
+ $Y2=0
cc_285 N_A_27_74#_c_273_n N_A_206_368#_c_644_n 0.00477971f $X=3.18 $Y=2.44 $X2=0
+ $Y2=0
cc_286 N_A_27_74#_c_274_n N_A_206_368#_c_583_n 0.00720135f $X=5.095 $Y=2.045
+ $X2=0 $Y2=0
cc_287 N_A_27_74#_M1028_g N_A_206_368#_c_583_n 7.96533e-19 $X=5.815 $Y=0.83
+ $X2=0 $Y2=0
cc_288 N_A_27_74#_c_274_n N_A_206_368#_c_584_n 0.031037f $X=5.095 $Y=2.045 $X2=0
+ $Y2=0
cc_289 N_A_27_74#_M1028_g N_A_206_368#_c_584_n 6.92466e-19 $X=5.815 $Y=0.83
+ $X2=0 $Y2=0
cc_290 N_A_27_74#_c_274_n N_A_206_368#_c_600_n 0.00926804f $X=5.095 $Y=2.045
+ $X2=0 $Y2=0
cc_291 N_A_27_74#_c_274_n N_A_206_368#_c_601_n 7.86426e-19 $X=5.095 $Y=2.045
+ $X2=0 $Y2=0
cc_292 N_A_27_74#_c_275_n N_A_206_368#_c_601_n 4.9727e-19 $X=5.74 $Y=1.765 $X2=0
+ $Y2=0
cc_293 N_A_27_74#_c_246_n N_A_206_368#_c_602_n 0.00662795f $X=0.955 $Y=1.765
+ $X2=0 $Y2=0
cc_294 N_A_27_74#_c_254_n N_A_206_368#_c_602_n 0.00584697f $X=0.76 $Y=1.95 $X2=0
+ $Y2=0
cc_295 N_A_27_74#_c_266_n N_A_206_368#_c_602_n 0.00736457f $X=0.905 $Y=1.045
+ $X2=0 $Y2=0
cc_296 N_A_27_74#_c_246_n N_A_206_368#_c_585_n 0.00268528f $X=0.955 $Y=1.765
+ $X2=0 $Y2=0
cc_297 N_A_27_74#_c_254_n N_A_206_368#_c_585_n 0.0101178f $X=0.76 $Y=1.95 $X2=0
+ $Y2=0
cc_298 N_A_27_74#_c_246_n N_A_206_368#_c_604_n 0.00572675f $X=0.955 $Y=1.765
+ $X2=0 $Y2=0
cc_299 N_A_27_74#_c_246_n N_A_206_368#_c_586_n 0.00235819f $X=0.955 $Y=1.765
+ $X2=0 $Y2=0
cc_300 N_A_27_74#_c_259_n N_A_206_368#_c_586_n 0.00573627f $X=1.815 $Y=0.815
+ $X2=0 $Y2=0
cc_301 N_A_27_74#_c_266_n N_A_206_368#_c_586_n 0.0274305f $X=0.905 $Y=1.045
+ $X2=0 $Y2=0
cc_302 N_A_27_74#_c_246_n N_A_206_368#_c_587_n 0.0211356f $X=0.955 $Y=1.765
+ $X2=0 $Y2=0
cc_303 N_A_27_74#_c_266_n N_A_206_368#_c_587_n 2.9577e-19 $X=0.905 $Y=1.045
+ $X2=0 $Y2=0
cc_304 N_A_27_74#_c_274_n N_A_206_368#_c_588_n 0.0216972f $X=5.095 $Y=2.045
+ $X2=0 $Y2=0
cc_305 N_A_27_74#_M1028_g N_A_206_368#_c_588_n 0.0201354f $X=5.815 $Y=0.83 $X2=0
+ $Y2=0
cc_306 N_A_27_74#_c_274_n N_A_206_368#_c_606_n 0.00402154f $X=5.095 $Y=2.045
+ $X2=0 $Y2=0
cc_307 N_A_27_74#_c_269_n N_A_696_458#_M1005_d 0.00205163f $X=5.665 $Y=0.382
+ $X2=-0.19 $Y2=-0.245
cc_308 N_A_27_74#_c_273_n N_A_696_458#_c_826_n 0.0324073f $X=3.18 $Y=2.44 $X2=0
+ $Y2=0
cc_309 N_A_27_74#_c_249_n N_A_696_458#_c_819_n 2.96657e-19 $X=3.145 $Y=1.09
+ $X2=0 $Y2=0
cc_310 N_A_27_74#_c_250_n N_A_696_458#_c_819_n 0.0020398f $X=3.145 $Y=1.24 $X2=0
+ $Y2=0
cc_311 N_A_27_74#_c_264_n N_A_696_458#_c_819_n 0.0119195f $X=3.79 $Y=1.75 $X2=0
+ $Y2=0
cc_312 N_A_27_74#_c_270_n N_A_696_458#_c_819_n 0.0114195f $X=3.287 $Y=1.75 $X2=0
+ $Y2=0
cc_313 N_A_27_74#_c_272_n N_A_696_458#_c_820_n 0.00698695f $X=3.18 $Y=2.35 $X2=0
+ $Y2=0
cc_314 N_A_27_74#_c_280_n N_A_696_458#_c_820_n 0.011502f $X=3.705 $Y=1.915 $X2=0
+ $Y2=0
cc_315 N_A_27_74#_c_281_n N_A_696_458#_c_820_n 0.0213588f $X=3.32 $Y=1.915 $X2=0
+ $Y2=0
cc_316 N_A_27_74#_c_264_n N_A_696_458#_c_820_n 0.0115948f $X=3.79 $Y=1.75 $X2=0
+ $Y2=0
cc_317 N_A_27_74#_c_261_n N_A_696_458#_c_821_n 3.98228e-19 $X=3.705 $Y=0.34
+ $X2=0 $Y2=0
cc_318 N_A_27_74#_c_263_n N_A_696_458#_c_821_n 0.00126253f $X=3.79 $Y=0.69 $X2=0
+ $Y2=0
cc_319 N_A_27_74#_c_264_n N_A_696_458#_c_821_n 0.00604635f $X=3.79 $Y=1.75 $X2=0
+ $Y2=0
cc_320 N_A_27_74#_c_385_p N_A_696_458#_c_821_n 0.0163588f $X=4.51 $Y=0.775 $X2=0
+ $Y2=0
cc_321 N_A_27_74#_c_386_p N_A_696_458#_c_821_n 0.00147235f $X=4.595 $Y=0.69
+ $X2=0 $Y2=0
cc_322 N_A_27_74#_c_272_n N_A_696_458#_c_828_n 0.00973828f $X=3.18 $Y=2.35 $X2=0
+ $Y2=0
cc_323 N_A_27_74#_c_280_n N_A_696_458#_c_828_n 0.00139488f $X=3.705 $Y=1.915
+ $X2=0 $Y2=0
cc_324 N_A_27_74#_c_281_n N_A_696_458#_c_828_n 3.11257e-19 $X=3.32 $Y=1.915
+ $X2=0 $Y2=0
cc_325 N_A_27_74#_c_264_n N_A_696_458#_c_822_n 0.0266789f $X=3.79 $Y=1.75 $X2=0
+ $Y2=0
cc_326 N_A_27_74#_c_385_p N_A_696_458#_c_822_n 0.0384244f $X=4.51 $Y=0.775 $X2=0
+ $Y2=0
cc_327 N_A_27_74#_c_385_p N_A_696_458#_c_823_n 0.00216189f $X=4.51 $Y=0.775
+ $X2=0 $Y2=0
cc_328 N_A_27_74#_M1028_g N_A_696_458#_c_824_n 3.19476e-19 $X=5.815 $Y=0.83
+ $X2=0 $Y2=0
cc_329 N_A_27_74#_c_385_p N_A_696_458#_c_824_n 0.00886892f $X=4.51 $Y=0.775
+ $X2=0 $Y2=0
cc_330 N_A_27_74#_c_269_n N_A_696_458#_c_824_n 0.0235144f $X=5.665 $Y=0.382
+ $X2=0 $Y2=0
cc_331 N_A_27_74#_c_274_n N_A_696_458#_c_825_n 0.0024411f $X=5.095 $Y=2.045
+ $X2=0 $Y2=0
cc_332 N_A_27_74#_c_274_n N_A_544_485#_c_913_n 0.014097f $X=5.095 $Y=2.045 $X2=0
+ $Y2=0
cc_333 N_A_27_74#_c_385_p N_A_544_485#_M1005_g 0.00231497f $X=4.51 $Y=0.775
+ $X2=0 $Y2=0
cc_334 N_A_27_74#_c_265_n N_A_544_485#_M1005_g 0.00279918f $X=4.68 $Y=0.34 $X2=0
+ $Y2=0
cc_335 N_A_27_74#_c_269_n N_A_544_485#_M1005_g 0.0104815f $X=5.665 $Y=0.382
+ $X2=0 $Y2=0
cc_336 N_A_27_74#_c_280_n N_A_544_485#_c_906_n 0.026331f $X=3.705 $Y=1.915 $X2=0
+ $Y2=0
cc_337 N_A_27_74#_c_270_n N_A_544_485#_c_906_n 0.0118712f $X=3.287 $Y=1.75 $X2=0
+ $Y2=0
cc_338 N_A_27_74#_c_250_n N_A_544_485#_c_907_n 0.00166025f $X=3.145 $Y=1.24
+ $X2=0 $Y2=0
cc_339 N_A_27_74#_c_280_n N_A_544_485#_c_907_n 0.0153093f $X=3.705 $Y=1.915
+ $X2=0 $Y2=0
cc_340 N_A_27_74#_c_281_n N_A_544_485#_c_907_n 0.00255136f $X=3.32 $Y=1.915
+ $X2=0 $Y2=0
cc_341 N_A_27_74#_c_264_n N_A_544_485#_c_907_n 0.00767638f $X=3.79 $Y=1.75 $X2=0
+ $Y2=0
cc_342 N_A_27_74#_c_270_n N_A_544_485#_c_907_n 0.0140774f $X=3.287 $Y=1.75 $X2=0
+ $Y2=0
cc_343 N_A_27_74#_c_272_n N_A_544_485#_c_915_n 0.00737544f $X=3.18 $Y=2.35 $X2=0
+ $Y2=0
cc_344 N_A_27_74#_c_273_n N_A_544_485#_c_915_n 0.0060122f $X=3.18 $Y=2.44 $X2=0
+ $Y2=0
cc_345 N_A_27_74#_c_280_n N_A_544_485#_c_915_n 0.0548044f $X=3.705 $Y=1.915
+ $X2=0 $Y2=0
cc_346 N_A_27_74#_c_281_n N_A_544_485#_c_915_n 0.00473468f $X=3.32 $Y=1.915
+ $X2=0 $Y2=0
cc_347 N_A_27_74#_c_249_n N_A_544_485#_c_909_n 0.00263846f $X=3.145 $Y=1.09
+ $X2=0 $Y2=0
cc_348 N_A_27_74#_c_250_n N_A_544_485#_c_909_n 0.00464436f $X=3.145 $Y=1.24
+ $X2=0 $Y2=0
cc_349 N_A_27_74#_c_264_n N_A_544_485#_c_909_n 0.0199406f $X=3.79 $Y=1.75 $X2=0
+ $Y2=0
cc_350 N_A_27_74#_c_270_n N_A_544_485#_c_909_n 0.00538348f $X=3.287 $Y=1.75
+ $X2=0 $Y2=0
cc_351 N_A_27_74#_c_280_n N_A_544_485#_c_910_n 0.0272824f $X=3.705 $Y=1.915
+ $X2=0 $Y2=0
cc_352 N_A_27_74#_c_264_n N_A_544_485#_c_910_n 0.00860245f $X=3.79 $Y=1.75 $X2=0
+ $Y2=0
cc_353 N_A_27_74#_c_273_n N_A_544_485#_c_917_n 0.0058613f $X=3.18 $Y=2.44 $X2=0
+ $Y2=0
cc_354 N_A_27_74#_c_249_n N_A_544_485#_c_911_n 0.00369274f $X=3.145 $Y=1.09
+ $X2=0 $Y2=0
cc_355 N_A_27_74#_c_261_n N_A_544_485#_c_911_n 0.0197592f $X=3.705 $Y=0.34 $X2=0
+ $Y2=0
cc_356 N_A_27_74#_c_264_n N_A_544_485#_c_911_n 0.00408327f $X=3.79 $Y=1.75 $X2=0
+ $Y2=0
cc_357 N_A_27_74#_c_274_n N_A_544_485#_c_912_n 0.0161801f $X=5.095 $Y=2.045
+ $X2=0 $Y2=0
cc_358 N_A_27_74#_c_280_n N_A_544_485#_c_912_n 0.00163538f $X=3.705 $Y=1.915
+ $X2=0 $Y2=0
cc_359 N_A_27_74#_c_264_n N_A_544_485#_c_912_n 7.01273e-19 $X=3.79 $Y=1.75 $X2=0
+ $Y2=0
cc_360 N_A_27_74#_c_275_n N_A_1226_296#_c_1026_n 0.00137256f $X=5.74 $Y=1.765
+ $X2=0 $Y2=0
cc_361 N_A_27_74#_M1028_g N_A_1226_296#_M1014_g 0.0373864f $X=5.815 $Y=0.83
+ $X2=0 $Y2=0
cc_362 N_A_27_74#_c_268_n N_A_1226_296#_M1014_g 0.00120024f $X=5.83 $Y=0.345
+ $X2=0 $Y2=0
cc_363 N_A_27_74#_M1028_g N_A_1226_296#_c_1023_n 0.00120248f $X=5.815 $Y=0.83
+ $X2=0 $Y2=0
cc_364 N_A_27_74#_M1028_g N_A_1226_296#_c_1024_n 0.0173687f $X=5.815 $Y=0.83
+ $X2=0 $Y2=0
cc_365 N_A_27_74#_c_274_n N_A_1034_424#_c_1193_n 0.0072886f $X=5.095 $Y=2.045
+ $X2=0 $Y2=0
cc_366 N_A_27_74#_M1028_g N_A_1034_424#_c_1198_n 0.00794457f $X=5.815 $Y=0.83
+ $X2=0 $Y2=0
cc_367 N_A_27_74#_c_267_n N_A_1034_424#_c_1198_n 0.0101797f $X=5.83 $Y=0.345
+ $X2=0 $Y2=0
cc_368 N_A_27_74#_c_268_n N_A_1034_424#_c_1198_n 5.32785e-19 $X=5.83 $Y=0.345
+ $X2=0 $Y2=0
cc_369 N_A_27_74#_c_269_n N_A_1034_424#_c_1198_n 0.0140733f $X=5.665 $Y=0.382
+ $X2=0 $Y2=0
cc_370 N_A_27_74#_c_275_n N_A_1034_424#_c_1194_n 0.0160859f $X=5.74 $Y=1.765
+ $X2=0 $Y2=0
cc_371 N_A_27_74#_c_274_n N_A_1034_424#_c_1195_n 9.55124e-19 $X=5.095 $Y=2.045
+ $X2=0 $Y2=0
cc_372 N_A_27_74#_c_275_n N_A_1034_424#_c_1195_n 0.00877163f $X=5.74 $Y=1.765
+ $X2=0 $Y2=0
cc_373 N_A_27_74#_M1028_g N_A_1034_424#_c_1183_n 0.00523836f $X=5.815 $Y=0.83
+ $X2=0 $Y2=0
cc_374 N_A_27_74#_c_275_n N_A_1034_424#_c_1184_n 0.0021257f $X=5.74 $Y=1.765
+ $X2=0 $Y2=0
cc_375 N_A_27_74#_M1028_g N_A_1034_424#_c_1184_n 0.0117463f $X=5.815 $Y=0.83
+ $X2=0 $Y2=0
cc_376 N_A_27_74#_M1028_g N_A_1034_424#_c_1185_n 0.00464647f $X=5.815 $Y=0.83
+ $X2=0 $Y2=0
cc_377 N_A_27_74#_c_267_n N_A_1034_424#_c_1185_n 0.00355696f $X=5.83 $Y=0.345
+ $X2=0 $Y2=0
cc_378 N_A_27_74#_c_268_n N_A_1034_424#_c_1185_n 0.00164778f $X=5.83 $Y=0.345
+ $X2=0 $Y2=0
cc_379 N_A_27_74#_M1028_g N_A_1034_424#_c_1186_n 0.00249192f $X=5.815 $Y=0.83
+ $X2=0 $Y2=0
cc_380 N_A_27_74#_c_298_n N_VPWR_M1015_d 0.00457874f $X=0.675 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_381 N_A_27_74#_c_254_n N_VPWR_M1015_d 0.0015936f $X=0.76 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_382 N_A_27_74#_c_246_n N_VPWR_c_1288_n 0.00486623f $X=0.955 $Y=1.765 $X2=0
+ $Y2=0
cc_383 N_A_27_74#_c_278_n N_VPWR_c_1288_n 0.0449718f $X=0.28 $Y=2.815 $X2=0
+ $Y2=0
cc_384 N_A_27_74#_c_298_n N_VPWR_c_1288_n 0.0148103f $X=0.675 $Y=2.035 $X2=0
+ $Y2=0
cc_385 N_A_27_74#_c_246_n N_VPWR_c_1289_n 0.00445602f $X=0.955 $Y=1.765 $X2=0
+ $Y2=0
cc_386 N_A_27_74#_c_246_n N_VPWR_c_1290_n 0.00246037f $X=0.955 $Y=1.765 $X2=0
+ $Y2=0
cc_387 N_A_27_74#_c_273_n N_VPWR_c_1298_n 9.63329e-19 $X=3.18 $Y=2.44 $X2=0
+ $Y2=0
cc_388 N_A_27_74#_c_274_n N_VPWR_c_1299_n 0.00278227f $X=5.095 $Y=2.045 $X2=0
+ $Y2=0
cc_389 N_A_27_74#_c_278_n N_VPWR_c_1302_n 0.0145938f $X=0.28 $Y=2.815 $X2=0
+ $Y2=0
cc_390 N_A_27_74#_c_246_n N_VPWR_c_1287_n 0.00862475f $X=0.955 $Y=1.765 $X2=0
+ $Y2=0
cc_391 N_A_27_74#_c_274_n N_VPWR_c_1287_n 0.0035639f $X=5.095 $Y=2.045 $X2=0
+ $Y2=0
cc_392 N_A_27_74#_c_278_n N_VPWR_c_1287_n 0.0120466f $X=0.28 $Y=2.815 $X2=0
+ $Y2=0
cc_393 N_A_27_74#_c_270_n N_A_437_503#_c_1413_n 0.00313016f $X=3.287 $Y=1.75
+ $X2=0 $Y2=0
cc_394 N_A_27_74#_c_249_n N_A_437_503#_c_1414_n 0.00138987f $X=3.145 $Y=1.09
+ $X2=0 $Y2=0
cc_395 N_A_27_74#_c_258_n N_A_437_503#_c_1414_n 6.4849e-19 $X=2.485 $Y=0.815
+ $X2=0 $Y2=0
cc_396 N_A_27_74#_c_261_n N_A_437_503#_c_1414_n 0.0045636f $X=3.705 $Y=0.34
+ $X2=0 $Y2=0
cc_397 N_A_27_74#_c_258_n N_A_437_503#_c_1415_n 0.0126712f $X=2.485 $Y=0.815
+ $X2=0 $Y2=0
cc_398 N_A_27_74#_c_249_n N_A_437_503#_c_1416_n 5.12891e-19 $X=3.145 $Y=1.09
+ $X2=0 $Y2=0
cc_399 N_A_27_74#_c_261_n N_A_437_503#_c_1416_n 0.0128799f $X=3.705 $Y=0.34
+ $X2=0 $Y2=0
cc_400 N_A_27_74#_c_252_n N_VGND_M1025_d 8.96075e-19 $X=0.675 $Y=1.045 $X2=-0.19
+ $Y2=-0.245
cc_401 N_A_27_74#_c_256_n N_VGND_M1025_d 5.22721e-19 $X=1.135 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_402 N_A_27_74#_c_266_n N_VGND_M1025_d 0.00979174f $X=0.905 $Y=1.045 $X2=-0.19
+ $Y2=-0.245
cc_403 N_A_27_74#_c_304_n N_VGND_M1025_d 0.00564292f $X=0.905 $Y=0.96 $X2=-0.19
+ $Y2=-0.245
cc_404 N_A_27_74#_c_258_n N_VGND_M1019_s 0.0151925f $X=2.485 $Y=0.815 $X2=0
+ $Y2=0
cc_405 N_A_27_74#_c_260_n N_VGND_M1019_s 0.0026851f $X=2.57 $Y=0.73 $X2=0 $Y2=0
cc_406 N_A_27_74#_c_385_p N_VGND_M1011_d 0.0144449f $X=4.51 $Y=0.775 $X2=0 $Y2=0
cc_407 N_A_27_74#_c_386_p N_VGND_M1011_d 0.00408409f $X=4.595 $Y=0.69 $X2=0
+ $Y2=0
cc_408 N_A_27_74#_c_265_n N_VGND_M1011_d 4.40008e-19 $X=4.68 $Y=0.34 $X2=0 $Y2=0
cc_409 N_A_27_74#_c_247_n N_VGND_c_1548_n 0.00189964f $X=1.12 $Y=1.22 $X2=0
+ $Y2=0
cc_410 N_A_27_74#_c_251_n N_VGND_c_1548_n 0.0164567f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_411 N_A_27_74#_c_252_n N_VGND_c_1548_n 0.00390521f $X=0.675 $Y=1.045 $X2=0
+ $Y2=0
cc_412 N_A_27_74#_c_256_n N_VGND_c_1548_n 0.0141863f $X=1.135 $Y=0.34 $X2=0
+ $Y2=0
cc_413 N_A_27_74#_c_266_n N_VGND_c_1548_n 0.0106391f $X=0.905 $Y=1.045 $X2=0
+ $Y2=0
cc_414 N_A_27_74#_c_304_n N_VGND_c_1548_n 0.0264745f $X=0.905 $Y=0.96 $X2=0
+ $Y2=0
cc_415 N_A_27_74#_c_255_n N_VGND_c_1549_n 0.0150375f $X=1.645 $Y=0.34 $X2=0
+ $Y2=0
cc_416 N_A_27_74#_c_257_n N_VGND_c_1549_n 0.0106642f $X=1.73 $Y=0.73 $X2=0 $Y2=0
cc_417 N_A_27_74#_c_258_n N_VGND_c_1549_n 0.025747f $X=2.485 $Y=0.815 $X2=0
+ $Y2=0
cc_418 N_A_27_74#_c_260_n N_VGND_c_1549_n 0.0104593f $X=2.57 $Y=0.73 $X2=0 $Y2=0
cc_419 N_A_27_74#_c_262_n N_VGND_c_1549_n 0.0148934f $X=2.655 $Y=0.34 $X2=0
+ $Y2=0
cc_420 N_A_27_74#_c_261_n N_VGND_c_1550_n 0.0124942f $X=3.705 $Y=0.34 $X2=0
+ $Y2=0
cc_421 N_A_27_74#_c_263_n N_VGND_c_1550_n 0.0054894f $X=3.79 $Y=0.69 $X2=0 $Y2=0
cc_422 N_A_27_74#_c_385_p N_VGND_c_1550_n 0.0191408f $X=4.51 $Y=0.775 $X2=0
+ $Y2=0
cc_423 N_A_27_74#_c_386_p N_VGND_c_1550_n 0.00706898f $X=4.595 $Y=0.69 $X2=0
+ $Y2=0
cc_424 N_A_27_74#_c_265_n N_VGND_c_1550_n 0.014421f $X=4.68 $Y=0.34 $X2=0 $Y2=0
cc_425 N_A_27_74#_c_267_n N_VGND_c_1551_n 0.0104475f $X=5.83 $Y=0.345 $X2=0
+ $Y2=0
cc_426 N_A_27_74#_c_268_n N_VGND_c_1551_n 0.00298617f $X=5.83 $Y=0.345 $X2=0
+ $Y2=0
cc_427 N_A_27_74#_c_258_n N_VGND_c_1557_n 0.00241577f $X=2.485 $Y=0.815 $X2=0
+ $Y2=0
cc_428 N_A_27_74#_c_261_n N_VGND_c_1557_n 0.0793141f $X=3.705 $Y=0.34 $X2=0
+ $Y2=0
cc_429 N_A_27_74#_c_262_n N_VGND_c_1557_n 0.0115448f $X=2.655 $Y=0.34 $X2=0
+ $Y2=0
cc_430 N_A_27_74#_c_385_p N_VGND_c_1557_n 0.00270562f $X=4.51 $Y=0.775 $X2=0
+ $Y2=0
cc_431 N_A_27_74#_c_251_n N_VGND_c_1559_n 0.0145639f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_432 N_A_27_74#_c_247_n N_VGND_c_1560_n 0.00278184f $X=1.12 $Y=1.22 $X2=0
+ $Y2=0
cc_433 N_A_27_74#_c_255_n N_VGND_c_1560_n 0.0440512f $X=1.645 $Y=0.34 $X2=0
+ $Y2=0
cc_434 N_A_27_74#_c_256_n N_VGND_c_1560_n 0.0118705f $X=1.135 $Y=0.34 $X2=0
+ $Y2=0
cc_435 N_A_27_74#_c_258_n N_VGND_c_1560_n 0.00254228f $X=2.485 $Y=0.815 $X2=0
+ $Y2=0
cc_436 N_A_27_74#_c_385_p N_VGND_c_1561_n 0.00262318f $X=4.51 $Y=0.775 $X2=0
+ $Y2=0
cc_437 N_A_27_74#_c_265_n N_VGND_c_1561_n 0.0120795f $X=4.68 $Y=0.34 $X2=0 $Y2=0
cc_438 N_A_27_74#_c_268_n N_VGND_c_1561_n 0.00653686f $X=5.83 $Y=0.345 $X2=0
+ $Y2=0
cc_439 N_A_27_74#_c_269_n N_VGND_c_1561_n 0.083814f $X=5.665 $Y=0.382 $X2=0
+ $Y2=0
cc_440 N_A_27_74#_c_247_n N_VGND_c_1569_n 0.00356305f $X=1.12 $Y=1.22 $X2=0
+ $Y2=0
cc_441 N_A_27_74#_c_251_n N_VGND_c_1569_n 0.0119984f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_442 N_A_27_74#_c_255_n N_VGND_c_1569_n 0.0245464f $X=1.645 $Y=0.34 $X2=0
+ $Y2=0
cc_443 N_A_27_74#_c_256_n N_VGND_c_1569_n 0.0061974f $X=1.135 $Y=0.34 $X2=0
+ $Y2=0
cc_444 N_A_27_74#_c_258_n N_VGND_c_1569_n 0.00901226f $X=2.485 $Y=0.815 $X2=0
+ $Y2=0
cc_445 N_A_27_74#_c_261_n N_VGND_c_1569_n 0.0418999f $X=3.705 $Y=0.34 $X2=0
+ $Y2=0
cc_446 N_A_27_74#_c_262_n N_VGND_c_1569_n 0.00582224f $X=2.655 $Y=0.34 $X2=0
+ $Y2=0
cc_447 N_A_27_74#_c_385_p N_VGND_c_1569_n 0.011451f $X=4.51 $Y=0.775 $X2=0 $Y2=0
cc_448 N_A_27_74#_c_265_n N_VGND_c_1569_n 0.00658903f $X=4.68 $Y=0.34 $X2=0
+ $Y2=0
cc_449 N_A_27_74#_c_268_n N_VGND_c_1569_n 0.0102677f $X=5.83 $Y=0.345 $X2=0
+ $Y2=0
cc_450 N_A_27_74#_c_269_n N_VGND_c_1569_n 0.0479538f $X=5.665 $Y=0.382 $X2=0
+ $Y2=0
cc_451 D N_A_206_368#_c_577_n 8.56213e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_452 N_D_c_519_n N_A_206_368#_c_577_n 0.0208842f $X=2.14 $Y=1.2 $X2=0 $Y2=0
cc_453 N_D_c_517_n N_A_206_368#_c_578_n 0.00903828f $X=2.695 $Y=1.125 $X2=0
+ $Y2=0
cc_454 N_D_c_521_n N_A_206_368#_c_589_n 0.0262574f $X=2.11 $Y=2.44 $X2=0 $Y2=0
cc_455 N_D_c_516_n N_A_206_368#_c_589_n 0.0139275f $X=2.62 $Y=1.2 $X2=0 $Y2=0
cc_456 N_D_c_522_n N_A_206_368#_c_589_n 0.00106267f $X=1.95 $Y=2.19 $X2=0 $Y2=0
cc_457 N_D_c_523_n N_A_206_368#_c_589_n 0.00402065f $X=1.95 $Y=2.025 $X2=0 $Y2=0
cc_458 N_D_c_519_n N_A_206_368#_c_589_n 0.0213315f $X=2.14 $Y=1.2 $X2=0 $Y2=0
cc_459 D N_A_206_368#_c_589_n 0.0171621f $X=2.16 $Y=1.665 $X2=0 $Y2=0
cc_460 N_D_c_521_n N_A_206_368#_c_590_n 0.0092456f $X=2.11 $Y=2.44 $X2=0 $Y2=0
cc_461 N_D_c_523_n N_A_206_368#_c_590_n 8.57545e-19 $X=1.95 $Y=2.025 $X2=0 $Y2=0
cc_462 N_D_c_521_n N_A_206_368#_c_591_n 0.0123832f $X=2.11 $Y=2.44 $X2=0 $Y2=0
cc_463 N_D_c_521_n N_A_206_368#_c_593_n 0.00442951f $X=2.11 $Y=2.44 $X2=0 $Y2=0
cc_464 D N_A_206_368#_c_582_n 0.00373037f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_465 N_D_c_521_n N_A_206_368#_c_594_n 0.0117885f $X=2.11 $Y=2.44 $X2=0 $Y2=0
cc_466 N_D_c_522_n N_A_206_368#_c_594_n 0.0233836f $X=1.95 $Y=2.19 $X2=0 $Y2=0
cc_467 N_D_c_521_n N_A_206_368#_c_682_n 0.0082193f $X=2.11 $Y=2.44 $X2=0 $Y2=0
cc_468 N_D_c_521_n N_A_206_368#_c_595_n 0.00458677f $X=2.11 $Y=2.44 $X2=0 $Y2=0
cc_469 N_D_c_521_n N_A_206_368#_c_596_n 0.00614093f $X=2.11 $Y=2.44 $X2=0 $Y2=0
cc_470 N_D_c_521_n N_A_206_368#_c_602_n 0.00725575f $X=2.11 $Y=2.44 $X2=0 $Y2=0
cc_471 N_D_c_522_n N_A_206_368#_c_602_n 0.0171484f $X=1.95 $Y=2.19 $X2=0 $Y2=0
cc_472 D N_A_206_368#_c_602_n 0.00905792f $X=2.16 $Y=1.665 $X2=0 $Y2=0
cc_473 D N_A_206_368#_c_585_n 0.00905792f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_474 N_D_c_521_n N_A_206_368#_c_604_n 0.0015521f $X=2.11 $Y=2.44 $X2=0 $Y2=0
cc_475 D N_A_206_368#_c_586_n 0.0257691f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_476 N_D_c_519_n N_A_206_368#_c_586_n 2.75227e-19 $X=2.14 $Y=1.2 $X2=0 $Y2=0
cc_477 D N_A_206_368#_c_587_n 0.00210284f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_478 N_D_c_521_n N_VPWR_c_1290_n 0.00129015f $X=2.11 $Y=2.44 $X2=0 $Y2=0
cc_479 N_D_c_521_n N_VPWR_c_1298_n 9.62598e-19 $X=2.11 $Y=2.44 $X2=0 $Y2=0
cc_480 N_D_c_521_n N_A_437_503#_c_1417_n 0.00727467f $X=2.11 $Y=2.44 $X2=0 $Y2=0
cc_481 N_D_c_522_n N_A_437_503#_c_1417_n 0.0145557f $X=1.95 $Y=2.19 $X2=0 $Y2=0
cc_482 N_D_c_516_n N_A_437_503#_c_1413_n 0.00408812f $X=2.62 $Y=1.2 $X2=0 $Y2=0
cc_483 N_D_c_523_n N_A_437_503#_c_1413_n 0.00721465f $X=1.95 $Y=2.025 $X2=0
+ $Y2=0
cc_484 D N_A_437_503#_c_1413_n 0.0410958f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_485 N_D_c_519_n N_A_437_503#_c_1413_n 0.0040357f $X=2.14 $Y=1.2 $X2=0 $Y2=0
cc_486 N_D_c_516_n N_A_437_503#_c_1414_n 0.00500174f $X=2.62 $Y=1.2 $X2=0 $Y2=0
cc_487 N_D_c_517_n N_A_437_503#_c_1414_n 0.0042308f $X=2.695 $Y=1.125 $X2=0
+ $Y2=0
cc_488 N_D_c_516_n N_A_437_503#_c_1415_n 0.00565997f $X=2.62 $Y=1.2 $X2=0 $Y2=0
cc_489 N_D_c_517_n N_A_437_503#_c_1415_n 0.00142021f $X=2.695 $Y=1.125 $X2=0
+ $Y2=0
cc_490 D N_A_437_503#_c_1415_n 0.00904419f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_491 N_D_c_517_n N_A_437_503#_c_1416_n 0.00139954f $X=2.695 $Y=1.125 $X2=0
+ $Y2=0
cc_492 N_D_c_521_n N_A_437_503#_c_1419_n 8.4471e-19 $X=2.11 $Y=2.44 $X2=0 $Y2=0
cc_493 N_D_c_523_n N_A_437_503#_c_1419_n 0.0109887f $X=1.95 $Y=2.025 $X2=0 $Y2=0
cc_494 N_D_c_517_n N_VGND_c_1549_n 5.12097e-19 $X=2.695 $Y=1.125 $X2=0 $Y2=0
cc_495 N_A_206_368#_c_597_n N_A_696_458#_M1027_d 0.00912383f $X=4.895 $Y=2.99
+ $X2=0 $Y2=0
cc_496 N_A_206_368#_c_584_n N_A_696_458#_M1027_d 0.00794144f $X=4.98 $Y=2.905
+ $X2=0 $Y2=0
cc_497 N_A_206_368#_c_595_n N_A_696_458#_c_826_n 0.00200131f $X=3.205 $Y=2.99
+ $X2=0 $Y2=0
cc_498 N_A_206_368#_c_643_n N_A_696_458#_c_826_n 0.00308339f $X=3.29 $Y=2.905
+ $X2=0 $Y2=0
cc_499 N_A_206_368#_c_697_p N_A_696_458#_c_826_n 0.0124316f $X=4.215 $Y=2.675
+ $X2=0 $Y2=0
cc_500 N_A_206_368#_c_698_p N_A_696_458#_c_826_n 0.00215988f $X=4.3 $Y=2.905
+ $X2=0 $Y2=0
cc_501 N_A_206_368#_c_598_n N_A_696_458#_c_826_n 6.88002e-19 $X=4.385 $Y=2.99
+ $X2=0 $Y2=0
cc_502 N_A_206_368#_M1017_g N_A_696_458#_c_821_n 0.036668f $X=3.6 $Y=0.72 $X2=0
+ $Y2=0
cc_503 N_A_206_368#_c_697_p N_A_696_458#_c_828_n 0.0048942f $X=4.215 $Y=2.675
+ $X2=0 $Y2=0
cc_504 N_A_206_368#_c_581_n N_A_696_458#_c_824_n 0.00883829f $X=5.23 $Y=1.15
+ $X2=0 $Y2=0
cc_505 N_A_206_368#_c_583_n N_A_696_458#_c_824_n 0.0272493f $X=4.98 $Y=1.54
+ $X2=0 $Y2=0
cc_506 N_A_206_368#_c_588_n N_A_696_458#_c_824_n 6.0283e-19 $X=5.355 $Y=1.315
+ $X2=0 $Y2=0
cc_507 N_A_206_368#_c_697_p N_A_696_458#_c_825_n 0.0113967f $X=4.215 $Y=2.675
+ $X2=0 $Y2=0
cc_508 N_A_206_368#_c_597_n N_A_696_458#_c_825_n 0.012787f $X=4.895 $Y=2.99
+ $X2=0 $Y2=0
cc_509 N_A_206_368#_c_583_n N_A_696_458#_c_825_n 0.0135469f $X=4.98 $Y=1.54
+ $X2=0 $Y2=0
cc_510 N_A_206_368#_c_584_n N_A_696_458#_c_825_n 0.086683f $X=4.98 $Y=2.905
+ $X2=0 $Y2=0
cc_511 N_A_206_368#_c_595_n N_A_544_485#_M1010_d 0.00234404f $X=3.205 $Y=2.99
+ $X2=0 $Y2=0
cc_512 N_A_206_368#_c_697_p N_A_544_485#_c_913_n 0.00634716f $X=4.215 $Y=2.675
+ $X2=0 $Y2=0
cc_513 N_A_206_368#_c_698_p N_A_544_485#_c_913_n 0.00470261f $X=4.3 $Y=2.905
+ $X2=0 $Y2=0
cc_514 N_A_206_368#_c_597_n N_A_544_485#_c_913_n 0.00981164f $X=4.895 $Y=2.99
+ $X2=0 $Y2=0
cc_515 N_A_206_368#_c_598_n N_A_544_485#_c_913_n 0.00324459f $X=4.385 $Y=2.99
+ $X2=0 $Y2=0
cc_516 N_A_206_368#_c_584_n N_A_544_485#_c_913_n 0.00225402f $X=4.98 $Y=2.905
+ $X2=0 $Y2=0
cc_517 N_A_206_368#_c_583_n N_A_544_485#_c_903_n 0.00148784f $X=4.98 $Y=1.54
+ $X2=0 $Y2=0
cc_518 N_A_206_368#_c_584_n N_A_544_485#_c_903_n 0.00530269f $X=4.98 $Y=2.905
+ $X2=0 $Y2=0
cc_519 N_A_206_368#_c_588_n N_A_544_485#_c_903_n 7.51073e-19 $X=5.355 $Y=1.315
+ $X2=0 $Y2=0
cc_520 N_A_206_368#_c_581_n N_A_544_485#_M1005_g 0.0125422f $X=5.23 $Y=1.15
+ $X2=0 $Y2=0
cc_521 N_A_206_368#_c_583_n N_A_544_485#_M1005_g 6.49327e-19 $X=4.98 $Y=1.54
+ $X2=0 $Y2=0
cc_522 N_A_206_368#_c_583_n N_A_544_485#_c_905_n 7.0138e-19 $X=4.98 $Y=1.54
+ $X2=0 $Y2=0
cc_523 N_A_206_368#_c_588_n N_A_544_485#_c_905_n 0.0125422f $X=5.355 $Y=1.315
+ $X2=0 $Y2=0
cc_524 N_A_206_368#_c_589_n N_A_544_485#_c_906_n 0.00491483f $X=2.44 $Y=1.74
+ $X2=0 $Y2=0
cc_525 N_A_206_368#_c_595_n N_A_544_485#_c_915_n 0.00429236f $X=3.205 $Y=2.99
+ $X2=0 $Y2=0
cc_526 N_A_206_368#_c_697_p N_A_544_485#_c_915_n 0.0669756f $X=4.215 $Y=2.675
+ $X2=0 $Y2=0
cc_527 N_A_206_368#_c_644_n N_A_544_485#_c_915_n 0.0108731f $X=3.375 $Y=2.675
+ $X2=0 $Y2=0
cc_528 N_A_206_368#_M1017_g N_A_544_485#_c_909_n 8.74784e-19 $X=3.6 $Y=0.72
+ $X2=0 $Y2=0
cc_529 N_A_206_368#_c_590_n N_A_544_485#_c_917_n 0.00113647f $X=2.645 $Y=2.26
+ $X2=0 $Y2=0
cc_530 N_A_206_368#_c_591_n N_A_544_485#_c_917_n 0.00467096f $X=2.645 $Y=2.35
+ $X2=0 $Y2=0
cc_531 N_A_206_368#_c_595_n N_A_544_485#_c_917_n 0.0225295f $X=3.205 $Y=2.99
+ $X2=0 $Y2=0
cc_532 N_A_206_368#_c_644_n N_A_544_485#_c_917_n 0.0120088f $X=3.375 $Y=2.675
+ $X2=0 $Y2=0
cc_533 N_A_206_368#_M1017_g N_A_544_485#_c_911_n 0.00371021f $X=3.6 $Y=0.72
+ $X2=0 $Y2=0
cc_534 N_A_206_368#_c_697_p N_A_544_485#_c_912_n 7.27956e-19 $X=4.215 $Y=2.675
+ $X2=0 $Y2=0
cc_535 N_A_206_368#_c_592_n N_A_1226_296#_c_1026_n 0.0218396f $X=5.63 $Y=2.465
+ $X2=0 $Y2=0
cc_536 N_A_206_368#_c_601_n N_A_1226_296#_c_1026_n 0.00223091f $X=5.79 $Y=2.215
+ $X2=0 $Y2=0
cc_537 N_A_206_368#_c_592_n N_A_1226_296#_c_1027_n 0.0137364f $X=5.63 $Y=2.465
+ $X2=0 $Y2=0
cc_538 N_A_206_368#_c_600_n N_A_1226_296#_c_1027_n 0.001726f $X=5.625 $Y=2.99
+ $X2=0 $Y2=0
cc_539 N_A_206_368#_c_601_n N_A_1226_296#_c_1027_n 0.00589975f $X=5.79 $Y=2.215
+ $X2=0 $Y2=0
cc_540 N_A_206_368#_c_600_n N_A_1034_424#_M1018_d 0.00579062f $X=5.625 $Y=2.99
+ $X2=0 $Y2=0
cc_541 N_A_206_368#_c_592_n N_A_1034_424#_c_1193_n 0.00555548f $X=5.63 $Y=2.465
+ $X2=0 $Y2=0
cc_542 N_A_206_368#_c_584_n N_A_1034_424#_c_1193_n 0.0602674f $X=4.98 $Y=2.905
+ $X2=0 $Y2=0
cc_543 N_A_206_368#_c_600_n N_A_1034_424#_c_1193_n 0.012787f $X=5.625 $Y=2.99
+ $X2=0 $Y2=0
cc_544 N_A_206_368#_c_601_n N_A_1034_424#_c_1193_n 0.0415397f $X=5.79 $Y=2.215
+ $X2=0 $Y2=0
cc_545 N_A_206_368#_c_583_n N_A_1034_424#_c_1198_n 0.0121339f $X=4.98 $Y=1.54
+ $X2=0 $Y2=0
cc_546 N_A_206_368#_c_588_n N_A_1034_424#_c_1198_n 0.00118963f $X=5.355 $Y=1.315
+ $X2=0 $Y2=0
cc_547 N_A_206_368#_c_592_n N_A_1034_424#_c_1194_n 0.00262346f $X=5.63 $Y=2.465
+ $X2=0 $Y2=0
cc_548 N_A_206_368#_c_583_n N_A_1034_424#_c_1194_n 0.00881428f $X=4.98 $Y=1.54
+ $X2=0 $Y2=0
cc_549 N_A_206_368#_c_601_n N_A_1034_424#_c_1194_n 0.0201862f $X=5.79 $Y=2.215
+ $X2=0 $Y2=0
cc_550 N_A_206_368#_c_583_n N_A_1034_424#_c_1195_n 0.0145175f $X=4.98 $Y=1.54
+ $X2=0 $Y2=0
cc_551 N_A_206_368#_c_584_n N_A_1034_424#_c_1195_n 0.0130363f $X=4.98 $Y=2.905
+ $X2=0 $Y2=0
cc_552 N_A_206_368#_c_581_n N_A_1034_424#_c_1183_n 0.0010414f $X=5.23 $Y=1.15
+ $X2=0 $Y2=0
cc_553 N_A_206_368#_c_583_n N_A_1034_424#_c_1184_n 0.018257f $X=4.98 $Y=1.54
+ $X2=0 $Y2=0
cc_554 N_A_206_368#_c_584_n N_A_1034_424#_c_1184_n 0.004994f $X=4.98 $Y=2.905
+ $X2=0 $Y2=0
cc_555 N_A_206_368#_c_588_n N_A_1034_424#_c_1184_n 4.99891e-19 $X=5.355 $Y=1.315
+ $X2=0 $Y2=0
cc_556 N_A_206_368#_c_583_n N_A_1034_424#_c_1186_n 0.0135592f $X=4.98 $Y=1.54
+ $X2=0 $Y2=0
cc_557 N_A_206_368#_c_588_n N_A_1034_424#_c_1186_n 6.08836e-19 $X=5.355 $Y=1.315
+ $X2=0 $Y2=0
cc_558 N_A_206_368#_c_594_n N_VPWR_M1008_s 0.01661f $X=1.995 $Y=2.61 $X2=0 $Y2=0
cc_559 N_A_206_368#_c_697_p N_VPWR_M1009_d 0.0148918f $X=4.215 $Y=2.675 $X2=0
+ $Y2=0
cc_560 N_A_206_368#_c_698_p N_VPWR_M1009_d 0.00233899f $X=4.3 $Y=2.905 $X2=0
+ $Y2=0
cc_561 N_A_206_368#_c_598_n N_VPWR_M1009_d 7.84928e-19 $X=4.385 $Y=2.99 $X2=0
+ $Y2=0
cc_562 N_A_206_368#_c_593_n N_VPWR_c_1288_n 0.0461218f $X=1.245 $Y=2.525 $X2=0
+ $Y2=0
cc_563 N_A_206_368#_c_594_n N_VPWR_c_1289_n 0.00322614f $X=1.995 $Y=2.61 $X2=0
+ $Y2=0
cc_564 N_A_206_368#_c_604_n N_VPWR_c_1289_n 0.0203945f $X=1.245 $Y=2.61 $X2=0
+ $Y2=0
cc_565 N_A_206_368#_c_594_n N_VPWR_c_1290_n 0.0128075f $X=1.995 $Y=2.61 $X2=0
+ $Y2=0
cc_566 N_A_206_368#_c_596_n N_VPWR_c_1290_n 0.0126856f $X=2.165 $Y=2.99 $X2=0
+ $Y2=0
cc_567 N_A_206_368#_c_604_n N_VPWR_c_1290_n 0.00883833f $X=1.245 $Y=2.61 $X2=0
+ $Y2=0
cc_568 N_A_206_368#_c_592_n N_VPWR_c_1291_n 5.65704e-19 $X=5.63 $Y=2.465 $X2=0
+ $Y2=0
cc_569 N_A_206_368#_c_600_n N_VPWR_c_1291_n 0.00810593f $X=5.625 $Y=2.99 $X2=0
+ $Y2=0
cc_570 N_A_206_368#_c_601_n N_VPWR_c_1291_n 0.0199785f $X=5.79 $Y=2.215 $X2=0
+ $Y2=0
cc_571 N_A_206_368#_c_595_n N_VPWR_c_1297_n 0.00788162f $X=3.205 $Y=2.99 $X2=0
+ $Y2=0
cc_572 N_A_206_368#_c_697_p N_VPWR_c_1297_n 0.0244596f $X=4.215 $Y=2.675 $X2=0
+ $Y2=0
cc_573 N_A_206_368#_c_598_n N_VPWR_c_1297_n 0.0125523f $X=4.385 $Y=2.99 $X2=0
+ $Y2=0
cc_574 N_A_206_368#_c_591_n N_VPWR_c_1298_n 7.35405e-19 $X=2.645 $Y=2.35 $X2=0
+ $Y2=0
cc_575 N_A_206_368#_c_594_n N_VPWR_c_1298_n 0.00282869f $X=1.995 $Y=2.61 $X2=0
+ $Y2=0
cc_576 N_A_206_368#_c_595_n N_VPWR_c_1298_n 0.0788186f $X=3.205 $Y=2.99 $X2=0
+ $Y2=0
cc_577 N_A_206_368#_c_596_n N_VPWR_c_1298_n 0.0119935f $X=2.165 $Y=2.99 $X2=0
+ $Y2=0
cc_578 N_A_206_368#_c_697_p N_VPWR_c_1298_n 0.00572505f $X=4.215 $Y=2.675 $X2=0
+ $Y2=0
cc_579 N_A_206_368#_c_592_n N_VPWR_c_1299_n 0.00278193f $X=5.63 $Y=2.465 $X2=0
+ $Y2=0
cc_580 N_A_206_368#_c_697_p N_VPWR_c_1299_n 0.00343944f $X=4.215 $Y=2.675 $X2=0
+ $Y2=0
cc_581 N_A_206_368#_c_597_n N_VPWR_c_1299_n 0.0324923f $X=4.895 $Y=2.99 $X2=0
+ $Y2=0
cc_582 N_A_206_368#_c_598_n N_VPWR_c_1299_n 0.0116996f $X=4.385 $Y=2.99 $X2=0
+ $Y2=0
cc_583 N_A_206_368#_c_600_n N_VPWR_c_1299_n 0.0588551f $X=5.625 $Y=2.99 $X2=0
+ $Y2=0
cc_584 N_A_206_368#_c_606_n N_VPWR_c_1299_n 0.0119597f $X=4.98 $Y=2.99 $X2=0
+ $Y2=0
cc_585 N_A_206_368#_c_592_n N_VPWR_c_1287_n 0.00356044f $X=5.63 $Y=2.465 $X2=0
+ $Y2=0
cc_586 N_A_206_368#_c_594_n N_VPWR_c_1287_n 0.0108304f $X=1.995 $Y=2.61 $X2=0
+ $Y2=0
cc_587 N_A_206_368#_c_595_n N_VPWR_c_1287_n 0.0456458f $X=3.205 $Y=2.99 $X2=0
+ $Y2=0
cc_588 N_A_206_368#_c_596_n N_VPWR_c_1287_n 0.00657291f $X=2.165 $Y=2.99 $X2=0
+ $Y2=0
cc_589 N_A_206_368#_c_697_p N_VPWR_c_1287_n 0.0169115f $X=4.215 $Y=2.675 $X2=0
+ $Y2=0
cc_590 N_A_206_368#_c_597_n N_VPWR_c_1287_n 0.0186896f $X=4.895 $Y=2.99 $X2=0
+ $Y2=0
cc_591 N_A_206_368#_c_598_n N_VPWR_c_1287_n 0.00634199f $X=4.385 $Y=2.99 $X2=0
+ $Y2=0
cc_592 N_A_206_368#_c_600_n N_VPWR_c_1287_n 0.0327104f $X=5.625 $Y=2.99 $X2=0
+ $Y2=0
cc_593 N_A_206_368#_c_604_n N_VPWR_c_1287_n 0.0168479f $X=1.245 $Y=2.61 $X2=0
+ $Y2=0
cc_594 N_A_206_368#_c_606_n N_VPWR_c_1287_n 0.00639333f $X=4.98 $Y=2.99 $X2=0
+ $Y2=0
cc_595 N_A_206_368#_c_595_n N_A_437_503#_M1008_d 0.00483859f $X=3.205 $Y=2.99
+ $X2=0 $Y2=0
cc_596 N_A_206_368#_c_590_n N_A_437_503#_c_1417_n 0.00234869f $X=2.645 $Y=2.26
+ $X2=0 $Y2=0
cc_597 N_A_206_368#_c_591_n N_A_437_503#_c_1417_n 0.00179946f $X=2.645 $Y=2.35
+ $X2=0 $Y2=0
cc_598 N_A_206_368#_c_594_n N_A_437_503#_c_1417_n 0.0133776f $X=1.995 $Y=2.61
+ $X2=0 $Y2=0
cc_599 N_A_206_368#_c_682_n N_A_437_503#_c_1417_n 0.00277431f $X=2.08 $Y=2.905
+ $X2=0 $Y2=0
cc_600 N_A_206_368#_c_595_n N_A_437_503#_c_1417_n 0.0127604f $X=3.205 $Y=2.99
+ $X2=0 $Y2=0
cc_601 N_A_206_368#_c_589_n N_A_437_503#_c_1413_n 0.0105505f $X=2.44 $Y=1.74
+ $X2=0 $Y2=0
cc_602 N_A_206_368#_c_590_n N_A_437_503#_c_1413_n 0.00357598f $X=2.645 $Y=2.26
+ $X2=0 $Y2=0
cc_603 N_A_206_368#_c_589_n N_A_437_503#_c_1414_n 5.89098e-19 $X=2.44 $Y=1.74
+ $X2=0 $Y2=0
cc_604 N_A_206_368#_c_589_n N_A_437_503#_c_1419_n 0.00557716f $X=2.44 $Y=1.74
+ $X2=0 $Y2=0
cc_605 N_A_206_368#_c_590_n N_A_437_503#_c_1419_n 0.0091371f $X=2.645 $Y=2.26
+ $X2=0 $Y2=0
cc_606 N_A_206_368#_c_595_n A_651_503# 3.89885e-19 $X=3.205 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_607 N_A_206_368#_c_643_n A_651_503# 0.0016105f $X=3.29 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_608 N_A_206_368#_c_697_p A_651_503# 0.00158555f $X=4.215 $Y=2.675 $X2=-0.19
+ $Y2=-0.245
cc_609 N_A_206_368#_c_644_n A_651_503# 6.16583e-19 $X=3.375 $Y=2.675 $X2=-0.19
+ $Y2=-0.245
cc_610 N_A_206_368#_c_600_n A_1141_508# 8.83155e-19 $X=5.625 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_611 N_A_206_368#_c_601_n A_1141_508# 0.00558111f $X=5.79 $Y=2.215 $X2=-0.19
+ $Y2=-0.245
cc_612 N_A_206_368#_c_577_n N_VGND_c_1549_n 0.00142208f $X=1.69 $Y=1.22 $X2=0
+ $Y2=0
cc_613 N_A_206_368#_c_578_n N_VGND_c_1549_n 0.0245958f $X=3.525 $Y=0.18 $X2=0
+ $Y2=0
cc_614 N_A_206_368#_c_578_n N_VGND_c_1550_n 0.00311957f $X=3.525 $Y=0.18 $X2=0
+ $Y2=0
cc_615 N_A_206_368#_M1017_g N_VGND_c_1550_n 5.84022e-19 $X=3.6 $Y=0.72 $X2=0
+ $Y2=0
cc_616 N_A_206_368#_c_578_n N_VGND_c_1557_n 0.0291559f $X=3.525 $Y=0.18 $X2=0
+ $Y2=0
cc_617 N_A_206_368#_c_579_n N_VGND_c_1560_n 0.0092256f $X=1.765 $Y=0.18 $X2=0
+ $Y2=0
cc_618 N_A_206_368#_c_581_n N_VGND_c_1561_n 7.26245e-19 $X=5.23 $Y=1.15 $X2=0
+ $Y2=0
cc_619 N_A_206_368#_c_578_n N_VGND_c_1569_n 0.0406918f $X=3.525 $Y=0.18 $X2=0
+ $Y2=0
cc_620 N_A_206_368#_c_579_n N_VGND_c_1569_n 0.00600553f $X=1.765 $Y=0.18 $X2=0
+ $Y2=0
cc_621 N_A_696_458#_c_826_n N_A_544_485#_c_913_n 0.0080054f $X=3.57 $Y=2.44
+ $X2=0 $Y2=0
cc_622 N_A_696_458#_c_820_n N_A_544_485#_c_913_n 0.00765991f $X=3.77 $Y=2.29
+ $X2=0 $Y2=0
cc_623 N_A_696_458#_c_825_n N_A_544_485#_c_913_n 0.00681984f $X=4.64 $Y=2.46
+ $X2=0 $Y2=0
cc_624 N_A_696_458#_c_825_n N_A_544_485#_c_903_n 0.00561133f $X=4.64 $Y=2.46
+ $X2=0 $Y2=0
cc_625 N_A_696_458#_c_821_n N_A_544_485#_M1005_g 0.00928538f $X=3.96 $Y=1.04
+ $X2=0 $Y2=0
cc_626 N_A_696_458#_c_823_n N_A_544_485#_M1005_g 0.0105347f $X=4.21 $Y=1.205
+ $X2=0 $Y2=0
cc_627 N_A_696_458#_c_824_n N_A_544_485#_M1005_g 0.0203393f $X=4.64 $Y=1.37
+ $X2=0 $Y2=0
cc_628 N_A_696_458#_c_819_n N_A_544_485#_c_905_n 8.00877e-19 $X=3.77 $Y=1.42
+ $X2=0 $Y2=0
cc_629 N_A_696_458#_c_823_n N_A_544_485#_c_905_n 0.00386517f $X=4.21 $Y=1.205
+ $X2=0 $Y2=0
cc_630 N_A_696_458#_c_824_n N_A_544_485#_c_905_n 0.00366748f $X=4.64 $Y=1.37
+ $X2=0 $Y2=0
cc_631 N_A_696_458#_c_825_n N_A_544_485#_c_905_n 0.00235604f $X=4.64 $Y=2.46
+ $X2=0 $Y2=0
cc_632 N_A_696_458#_c_819_n N_A_544_485#_c_907_n 0.00130712f $X=3.77 $Y=1.42
+ $X2=0 $Y2=0
cc_633 N_A_696_458#_c_820_n N_A_544_485#_c_915_n 0.00383953f $X=3.77 $Y=2.29
+ $X2=0 $Y2=0
cc_634 N_A_696_458#_c_828_n N_A_544_485#_c_915_n 0.0142234f $X=3.77 $Y=2.365
+ $X2=0 $Y2=0
cc_635 N_A_696_458#_c_825_n N_A_544_485#_c_915_n 0.0133617f $X=4.64 $Y=2.46
+ $X2=0 $Y2=0
cc_636 N_A_696_458#_c_819_n N_A_544_485#_c_909_n 0.00112127f $X=3.77 $Y=1.42
+ $X2=0 $Y2=0
cc_637 N_A_696_458#_c_820_n N_A_544_485#_c_910_n 0.00498304f $X=3.77 $Y=2.29
+ $X2=0 $Y2=0
cc_638 N_A_696_458#_c_822_n N_A_544_485#_c_910_n 0.0186936f $X=4.555 $Y=1.2
+ $X2=0 $Y2=0
cc_639 N_A_696_458#_c_823_n N_A_544_485#_c_910_n 0.00120762f $X=4.21 $Y=1.205
+ $X2=0 $Y2=0
cc_640 N_A_696_458#_c_825_n N_A_544_485#_c_910_n 0.0451133f $X=4.64 $Y=2.46
+ $X2=0 $Y2=0
cc_641 N_A_696_458#_c_820_n N_A_544_485#_c_912_n 0.0235456f $X=3.77 $Y=2.29
+ $X2=0 $Y2=0
cc_642 N_A_696_458#_c_822_n N_A_544_485#_c_912_n 0.00714445f $X=4.555 $Y=1.2
+ $X2=0 $Y2=0
cc_643 N_A_696_458#_c_823_n N_A_544_485#_c_912_n 0.0154938f $X=4.21 $Y=1.205
+ $X2=0 $Y2=0
cc_644 N_A_696_458#_c_825_n N_A_544_485#_c_912_n 0.0180063f $X=4.64 $Y=2.46
+ $X2=0 $Y2=0
cc_645 N_A_696_458#_c_824_n N_A_1034_424#_c_1183_n 0.00408737f $X=4.64 $Y=1.37
+ $X2=0 $Y2=0
cc_646 N_A_696_458#_c_824_n N_A_1034_424#_c_1186_n 3.52924e-19 $X=4.64 $Y=1.37
+ $X2=0 $Y2=0
cc_647 N_A_696_458#_c_826_n N_VPWR_c_1297_n 0.00193758f $X=3.57 $Y=2.44 $X2=0
+ $Y2=0
cc_648 N_A_696_458#_c_826_n N_VPWR_c_1298_n 0.00422085f $X=3.57 $Y=2.44 $X2=0
+ $Y2=0
cc_649 N_A_696_458#_c_826_n N_VPWR_c_1287_n 0.00537853f $X=3.57 $Y=2.44 $X2=0
+ $Y2=0
cc_650 N_A_696_458#_c_821_n N_VGND_c_1550_n 0.00165146f $X=3.96 $Y=1.04 $X2=0
+ $Y2=0
cc_651 N_A_696_458#_c_821_n N_VGND_c_1557_n 0.00374061f $X=3.96 $Y=1.04 $X2=0
+ $Y2=0
cc_652 N_A_696_458#_c_821_n N_VGND_c_1569_n 0.00502397f $X=3.96 $Y=1.04 $X2=0
+ $Y2=0
cc_653 N_A_544_485#_c_915_n N_VPWR_M1009_d 0.0031054f $X=4.055 $Y=2.335 $X2=0
+ $Y2=0
cc_654 N_A_544_485#_c_910_n N_VPWR_M1009_d 4.42249e-19 $X=4.22 $Y=1.795 $X2=0
+ $Y2=0
cc_655 N_A_544_485#_c_913_n N_VPWR_c_1297_n 9.44664e-19 $X=4.415 $Y=2.045 $X2=0
+ $Y2=0
cc_656 N_A_544_485#_c_913_n N_VPWR_c_1299_n 0.00278227f $X=4.415 $Y=2.045 $X2=0
+ $Y2=0
cc_657 N_A_544_485#_c_913_n N_VPWR_c_1287_n 0.00360398f $X=4.415 $Y=2.045 $X2=0
+ $Y2=0
cc_658 N_A_544_485#_c_906_n N_A_437_503#_c_1417_n 0.00641246f $X=2.9 $Y=2.25
+ $X2=0 $Y2=0
cc_659 N_A_544_485#_c_917_n N_A_437_503#_c_1417_n 0.0288961f $X=2.87 $Y=2.335
+ $X2=0 $Y2=0
cc_660 N_A_544_485#_c_906_n N_A_437_503#_c_1413_n 0.0268242f $X=2.9 $Y=2.25
+ $X2=0 $Y2=0
cc_661 N_A_544_485#_c_908_n N_A_437_503#_c_1413_n 0.0140664f $X=2.985 $Y=1.495
+ $X2=0 $Y2=0
cc_662 N_A_544_485#_c_909_n N_A_437_503#_c_1413_n 0.00500637f $X=3.26 $Y=1.41
+ $X2=0 $Y2=0
cc_663 N_A_544_485#_c_907_n N_A_437_503#_c_1414_n 8.03474e-19 $X=3.175 $Y=1.495
+ $X2=0 $Y2=0
cc_664 N_A_544_485#_c_908_n N_A_437_503#_c_1414_n 0.0157395f $X=2.985 $Y=1.495
+ $X2=0 $Y2=0
cc_665 N_A_544_485#_c_909_n N_A_437_503#_c_1414_n 0.0128044f $X=3.26 $Y=1.41
+ $X2=0 $Y2=0
cc_666 N_A_544_485#_c_909_n N_A_437_503#_c_1416_n 0.00579978f $X=3.26 $Y=1.41
+ $X2=0 $Y2=0
cc_667 N_A_544_485#_c_906_n N_A_437_503#_c_1419_n 0.0126271f $X=2.9 $Y=2.25
+ $X2=0 $Y2=0
cc_668 N_A_544_485#_M1005_g N_VGND_c_1550_n 8.804e-19 $X=4.755 $Y=0.655 $X2=0
+ $Y2=0
cc_669 N_A_544_485#_M1005_g N_VGND_c_1561_n 0.00390708f $X=4.755 $Y=0.655 $X2=0
+ $Y2=0
cc_670 N_A_544_485#_M1005_g N_VGND_c_1569_n 0.00542671f $X=4.755 $Y=0.655 $X2=0
+ $Y2=0
cc_671 N_A_1226_296#_c_1026_n N_A_1034_424#_c_1188_n 0.0157794f $X=6.255
+ $Y=2.375 $X2=0 $Y2=0
cc_672 N_A_1226_296#_c_1027_n N_A_1034_424#_c_1188_n 0.0127083f $X=6.255
+ $Y=2.465 $X2=0 $Y2=0
cc_673 N_A_1226_296#_c_1033_n N_A_1034_424#_c_1188_n 0.0158458f $X=6.985
+ $Y=2.265 $X2=0 $Y2=0
cc_674 N_A_1226_296#_c_1026_n N_A_1034_424#_c_1181_n 0.00192219f $X=6.255
+ $Y=2.375 $X2=0 $Y2=0
cc_675 N_A_1226_296#_c_1028_n N_A_1034_424#_c_1181_n 0.0011245f $X=7.745
+ $Y=1.765 $X2=0 $Y2=0
cc_676 N_A_1226_296#_c_1032_n N_A_1034_424#_c_1181_n 0.00392604f $X=6.82
+ $Y=1.805 $X2=0 $Y2=0
cc_677 N_A_1226_296#_c_1021_n N_A_1034_424#_c_1181_n 0.011068f $X=7.47 $Y=1.465
+ $X2=0 $Y2=0
cc_678 N_A_1226_296#_c_1023_n N_A_1034_424#_c_1181_n 0.00101768f $X=6.295
+ $Y=1.645 $X2=0 $Y2=0
cc_679 N_A_1226_296#_c_1025_n N_A_1034_424#_c_1181_n 0.00200738f $X=9.08
+ $Y=1.532 $X2=0 $Y2=0
cc_680 N_A_1226_296#_c_1028_n N_A_1034_424#_c_1190_n 0.00471449f $X=7.745
+ $Y=1.765 $X2=0 $Y2=0
cc_681 N_A_1226_296#_c_1033_n N_A_1034_424#_c_1190_n 0.00966319f $X=6.985
+ $Y=2.265 $X2=0 $Y2=0
cc_682 N_A_1226_296#_c_1021_n N_A_1034_424#_c_1190_n 0.00476867f $X=7.47
+ $Y=1.465 $X2=0 $Y2=0
cc_683 N_A_1226_296#_c_1026_n N_A_1034_424#_c_1191_n 0.00678475f $X=6.255
+ $Y=2.375 $X2=0 $Y2=0
cc_684 N_A_1226_296#_c_1032_n N_A_1034_424#_c_1191_n 0.00633358f $X=6.82
+ $Y=1.805 $X2=0 $Y2=0
cc_685 N_A_1226_296#_c_1033_n N_A_1034_424#_c_1191_n 0.00504076f $X=6.985
+ $Y=2.265 $X2=0 $Y2=0
cc_686 N_A_1226_296#_c_1028_n N_A_1034_424#_c_1192_n 0.0151007f $X=7.745
+ $Y=1.765 $X2=0 $Y2=0
cc_687 N_A_1226_296#_c_1033_n N_A_1034_424#_c_1192_n 0.0132035f $X=6.985
+ $Y=2.265 $X2=0 $Y2=0
cc_688 N_A_1226_296#_M1000_g N_A_1034_424#_c_1182_n 0.0139896f $X=7.73 $Y=0.74
+ $X2=0 $Y2=0
cc_689 N_A_1226_296#_c_1018_n N_A_1034_424#_c_1182_n 0.0119658f $X=7.015 $Y=0.88
+ $X2=0 $Y2=0
cc_690 N_A_1226_296#_c_1019_n N_A_1034_424#_c_1182_n 4.43891e-19 $X=7.055
+ $Y=0.515 $X2=0 $Y2=0
cc_691 N_A_1226_296#_c_1020_n N_A_1034_424#_c_1182_n 0.00658917f $X=7.385 $Y=1.3
+ $X2=0 $Y2=0
cc_692 N_A_1226_296#_M1014_g N_A_1034_424#_c_1198_n 9.05229e-19 $X=6.28 $Y=0.83
+ $X2=0 $Y2=0
cc_693 N_A_1226_296#_c_1026_n N_A_1034_424#_c_1194_n 9.22994e-19 $X=6.255
+ $Y=2.375 $X2=0 $Y2=0
cc_694 N_A_1226_296#_c_1023_n N_A_1034_424#_c_1194_n 0.00868849f $X=6.295
+ $Y=1.645 $X2=0 $Y2=0
cc_695 N_A_1226_296#_M1014_g N_A_1034_424#_c_1183_n 9.79059e-19 $X=6.28 $Y=0.83
+ $X2=0 $Y2=0
cc_696 N_A_1226_296#_M1014_g N_A_1034_424#_c_1184_n 9.79506e-19 $X=6.28 $Y=0.83
+ $X2=0 $Y2=0
cc_697 N_A_1226_296#_c_1023_n N_A_1034_424#_c_1184_n 0.0113414f $X=6.295
+ $Y=1.645 $X2=0 $Y2=0
cc_698 N_A_1226_296#_c_1024_n N_A_1034_424#_c_1184_n 2.81745e-19 $X=6.295
+ $Y=1.645 $X2=0 $Y2=0
cc_699 N_A_1226_296#_M1014_g N_A_1034_424#_c_1185_n 0.0186101f $X=6.28 $Y=0.83
+ $X2=0 $Y2=0
cc_700 N_A_1226_296#_c_1032_n N_A_1034_424#_c_1185_n 0.0166842f $X=6.82 $Y=1.805
+ $X2=0 $Y2=0
cc_701 N_A_1226_296#_c_1018_n N_A_1034_424#_c_1185_n 0.0182385f $X=7.015 $Y=0.88
+ $X2=0 $Y2=0
cc_702 N_A_1226_296#_c_1020_n N_A_1034_424#_c_1185_n 0.00893364f $X=7.385 $Y=1.3
+ $X2=0 $Y2=0
cc_703 N_A_1226_296#_c_1021_n N_A_1034_424#_c_1185_n 0.0467985f $X=7.47 $Y=1.465
+ $X2=0 $Y2=0
cc_704 N_A_1226_296#_c_1023_n N_A_1034_424#_c_1185_n 0.0276095f $X=6.295
+ $Y=1.645 $X2=0 $Y2=0
cc_705 N_A_1226_296#_c_1024_n N_A_1034_424#_c_1185_n 0.0013544f $X=6.295
+ $Y=1.645 $X2=0 $Y2=0
cc_706 N_A_1226_296#_M1014_g N_A_1034_424#_c_1187_n 0.0058711f $X=6.28 $Y=0.83
+ $X2=0 $Y2=0
cc_707 N_A_1226_296#_c_1018_n N_A_1034_424#_c_1187_n 0.00303145f $X=7.015
+ $Y=0.88 $X2=0 $Y2=0
cc_708 N_A_1226_296#_c_1020_n N_A_1034_424#_c_1187_n 0.00199303f $X=7.385 $Y=1.3
+ $X2=0 $Y2=0
cc_709 N_A_1226_296#_c_1021_n N_A_1034_424#_c_1187_n 0.00664738f $X=7.47
+ $Y=1.465 $X2=0 $Y2=0
cc_710 N_A_1226_296#_c_1024_n N_A_1034_424#_c_1187_n 0.0111429f $X=6.295
+ $Y=1.645 $X2=0 $Y2=0
cc_711 N_A_1226_296#_c_1025_n N_A_1034_424#_c_1187_n 0.017195f $X=9.08 $Y=1.532
+ $X2=0 $Y2=0
cc_712 N_A_1226_296#_c_1021_n N_VPWR_M1029_d 0.00189743f $X=7.47 $Y=1.465 $X2=0
+ $Y2=0
cc_713 N_A_1226_296#_c_1027_n N_VPWR_c_1291_n 0.0145978f $X=6.255 $Y=2.465 $X2=0
+ $Y2=0
cc_714 N_A_1226_296#_c_1032_n N_VPWR_c_1291_n 0.00619462f $X=6.82 $Y=1.805 $X2=0
+ $Y2=0
cc_715 N_A_1226_296#_c_1033_n N_VPWR_c_1291_n 0.0206791f $X=6.985 $Y=2.265 $X2=0
+ $Y2=0
cc_716 N_A_1226_296#_c_1023_n N_VPWR_c_1291_n 0.00531773f $X=6.295 $Y=1.645
+ $X2=0 $Y2=0
cc_717 N_A_1226_296#_c_1024_n N_VPWR_c_1291_n 6.54187e-19 $X=6.295 $Y=1.645
+ $X2=0 $Y2=0
cc_718 N_A_1226_296#_c_1028_n N_VPWR_c_1292_n 0.00727539f $X=7.745 $Y=1.765
+ $X2=0 $Y2=0
cc_719 N_A_1226_296#_c_1033_n N_VPWR_c_1292_n 0.0606477f $X=6.985 $Y=2.265 $X2=0
+ $Y2=0
cc_720 N_A_1226_296#_c_1021_n N_VPWR_c_1292_n 0.0103456f $X=7.47 $Y=1.465 $X2=0
+ $Y2=0
cc_721 N_A_1226_296#_c_1022_n N_VPWR_c_1292_n 0.00594822f $X=8.5 $Y=1.465 $X2=0
+ $Y2=0
cc_722 N_A_1226_296#_c_1028_n N_VPWR_c_1293_n 0.00445602f $X=7.745 $Y=1.765
+ $X2=0 $Y2=0
cc_723 N_A_1226_296#_c_1029_n N_VPWR_c_1293_n 0.00445602f $X=8.195 $Y=1.765
+ $X2=0 $Y2=0
cc_724 N_A_1226_296#_c_1029_n N_VPWR_c_1294_n 0.00586501f $X=8.195 $Y=1.765
+ $X2=0 $Y2=0
cc_725 N_A_1226_296#_c_1030_n N_VPWR_c_1294_n 0.00586501f $X=8.645 $Y=1.765
+ $X2=0 $Y2=0
cc_726 N_A_1226_296#_c_1031_n N_VPWR_c_1296_n 0.0100892f $X=9.095 $Y=1.765 $X2=0
+ $Y2=0
cc_727 N_A_1226_296#_c_1027_n N_VPWR_c_1299_n 0.00413917f $X=6.255 $Y=2.465
+ $X2=0 $Y2=0
cc_728 N_A_1226_296#_c_1033_n N_VPWR_c_1300_n 0.014552f $X=6.985 $Y=2.265 $X2=0
+ $Y2=0
cc_729 N_A_1226_296#_c_1030_n N_VPWR_c_1301_n 0.00445602f $X=8.645 $Y=1.765
+ $X2=0 $Y2=0
cc_730 N_A_1226_296#_c_1031_n N_VPWR_c_1301_n 0.00445602f $X=9.095 $Y=1.765
+ $X2=0 $Y2=0
cc_731 N_A_1226_296#_c_1027_n N_VPWR_c_1287_n 0.00856988f $X=6.255 $Y=2.465
+ $X2=0 $Y2=0
cc_732 N_A_1226_296#_c_1028_n N_VPWR_c_1287_n 0.00858383f $X=7.745 $Y=1.765
+ $X2=0 $Y2=0
cc_733 N_A_1226_296#_c_1029_n N_VPWR_c_1287_n 0.00857589f $X=8.195 $Y=1.765
+ $X2=0 $Y2=0
cc_734 N_A_1226_296#_c_1030_n N_VPWR_c_1287_n 0.00857589f $X=8.645 $Y=1.765
+ $X2=0 $Y2=0
cc_735 N_A_1226_296#_c_1031_n N_VPWR_c_1287_n 0.00861084f $X=9.095 $Y=1.765
+ $X2=0 $Y2=0
cc_736 N_A_1226_296#_c_1033_n N_VPWR_c_1287_n 0.0119791f $X=6.985 $Y=2.265 $X2=0
+ $Y2=0
cc_737 N_A_1226_296#_c_1028_n N_Q_c_1474_n 0.0121997f $X=7.745 $Y=1.765 $X2=0
+ $Y2=0
cc_738 N_A_1226_296#_c_1029_n N_Q_c_1474_n 0.0125029f $X=8.195 $Y=1.765 $X2=0
+ $Y2=0
cc_739 N_A_1226_296#_c_1030_n N_Q_c_1474_n 6.9119e-19 $X=8.645 $Y=1.765 $X2=0
+ $Y2=0
cc_740 N_A_1226_296#_c_1033_n N_Q_c_1474_n 0.00216738f $X=6.985 $Y=2.265 $X2=0
+ $Y2=0
cc_741 N_A_1226_296#_M1000_g N_Q_c_1468_n 4.78065e-19 $X=7.73 $Y=0.74 $X2=0
+ $Y2=0
cc_742 N_A_1226_296#_M1004_g N_Q_c_1468_n 0.00872666f $X=8.2 $Y=0.74 $X2=0 $Y2=0
cc_743 N_A_1226_296#_M1012_g N_Q_c_1468_n 6.31773e-19 $X=8.65 $Y=0.74 $X2=0
+ $Y2=0
cc_744 N_A_1226_296#_c_1029_n N_Q_c_1475_n 0.0120074f $X=8.195 $Y=1.765 $X2=0
+ $Y2=0
cc_745 N_A_1226_296#_c_1030_n N_Q_c_1475_n 0.0124686f $X=8.645 $Y=1.765 $X2=0
+ $Y2=0
cc_746 N_A_1226_296#_c_1022_n N_Q_c_1475_n 0.0389377f $X=8.5 $Y=1.465 $X2=0
+ $Y2=0
cc_747 N_A_1226_296#_c_1025_n N_Q_c_1475_n 0.00757172f $X=9.08 $Y=1.532 $X2=0
+ $Y2=0
cc_748 N_A_1226_296#_c_1028_n N_Q_c_1476_n 0.00354716f $X=7.745 $Y=1.765 $X2=0
+ $Y2=0
cc_749 N_A_1226_296#_c_1029_n N_Q_c_1476_n 9.3899e-19 $X=8.195 $Y=1.765 $X2=0
+ $Y2=0
cc_750 N_A_1226_296#_c_1033_n N_Q_c_1476_n 0.00206945f $X=6.985 $Y=2.265 $X2=0
+ $Y2=0
cc_751 N_A_1226_296#_c_1021_n N_Q_c_1476_n 0.00472878f $X=7.47 $Y=1.465 $X2=0
+ $Y2=0
cc_752 N_A_1226_296#_c_1022_n N_Q_c_1476_n 0.0276943f $X=8.5 $Y=1.465 $X2=0
+ $Y2=0
cc_753 N_A_1226_296#_c_1025_n N_Q_c_1476_n 0.00776454f $X=9.08 $Y=1.532 $X2=0
+ $Y2=0
cc_754 N_A_1226_296#_M1004_g N_Q_c_1469_n 0.01127f $X=8.2 $Y=0.74 $X2=0 $Y2=0
cc_755 N_A_1226_296#_M1012_g N_Q_c_1469_n 0.0117712f $X=8.65 $Y=0.74 $X2=0 $Y2=0
cc_756 N_A_1226_296#_c_1022_n N_Q_c_1469_n 0.0378697f $X=8.5 $Y=1.465 $X2=0
+ $Y2=0
cc_757 N_A_1226_296#_c_1025_n N_Q_c_1469_n 0.00269047f $X=9.08 $Y=1.532 $X2=0
+ $Y2=0
cc_758 N_A_1226_296#_M1000_g N_Q_c_1470_n 2.54377e-19 $X=7.73 $Y=0.74 $X2=0
+ $Y2=0
cc_759 N_A_1226_296#_M1004_g N_Q_c_1470_n 9.64852e-19 $X=8.2 $Y=0.74 $X2=0 $Y2=0
cc_760 N_A_1226_296#_c_1020_n N_Q_c_1470_n 0.00225318f $X=7.385 $Y=1.3 $X2=0
+ $Y2=0
cc_761 N_A_1226_296#_c_1022_n N_Q_c_1470_n 0.0277206f $X=8.5 $Y=1.465 $X2=0
+ $Y2=0
cc_762 N_A_1226_296#_c_1025_n N_Q_c_1470_n 0.00326139f $X=9.08 $Y=1.532 $X2=0
+ $Y2=0
cc_763 N_A_1226_296#_M1004_g N_Q_c_1471_n 6.44501e-19 $X=8.2 $Y=0.74 $X2=0 $Y2=0
cc_764 N_A_1226_296#_M1012_g N_Q_c_1471_n 0.00897582f $X=8.65 $Y=0.74 $X2=0
+ $Y2=0
cc_765 N_A_1226_296#_M1030_g N_Q_c_1471_n 0.00801138f $X=9.08 $Y=0.74 $X2=0
+ $Y2=0
cc_766 N_A_1226_296#_M1012_g N_Q_c_1472_n 0.00257108f $X=8.65 $Y=0.74 $X2=0
+ $Y2=0
cc_767 N_A_1226_296#_M1030_g N_Q_c_1472_n 0.00861468f $X=9.08 $Y=0.74 $X2=0
+ $Y2=0
cc_768 N_A_1226_296#_c_1031_n N_Q_c_1472_n 0.0019451f $X=9.095 $Y=1.765 $X2=0
+ $Y2=0
cc_769 N_A_1226_296#_c_1022_n N_Q_c_1472_n 0.022032f $X=8.5 $Y=1.465 $X2=0 $Y2=0
cc_770 N_A_1226_296#_c_1025_n N_Q_c_1472_n 0.0366525f $X=9.08 $Y=1.532 $X2=0
+ $Y2=0
cc_771 N_A_1226_296#_M1012_g N_Q_c_1473_n 0.00131511f $X=8.65 $Y=0.74 $X2=0
+ $Y2=0
cc_772 N_A_1226_296#_M1030_g N_Q_c_1473_n 0.00212711f $X=9.08 $Y=0.74 $X2=0
+ $Y2=0
cc_773 N_A_1226_296#_c_1025_n N_Q_c_1473_n 0.00148648f $X=9.08 $Y=1.532 $X2=0
+ $Y2=0
cc_774 N_A_1226_296#_c_1030_n Q 0.00114729f $X=8.645 $Y=1.765 $X2=0 $Y2=0
cc_775 N_A_1226_296#_c_1031_n Q 0.00304071f $X=9.095 $Y=1.765 $X2=0 $Y2=0
cc_776 N_A_1226_296#_c_1025_n Q 0.00466594f $X=9.08 $Y=1.532 $X2=0 $Y2=0
cc_777 N_A_1226_296#_c_1029_n Q 6.9119e-19 $X=8.195 $Y=1.765 $X2=0 $Y2=0
cc_778 N_A_1226_296#_c_1030_n Q 0.0125029f $X=8.645 $Y=1.765 $X2=0 $Y2=0
cc_779 N_A_1226_296#_c_1031_n Q 0.0118573f $X=9.095 $Y=1.765 $X2=0 $Y2=0
cc_780 N_A_1226_296#_c_1018_n N_VGND_M1024_d 0.00274889f $X=7.015 $Y=0.88 $X2=0
+ $Y2=0
cc_781 N_A_1226_296#_c_1020_n N_VGND_M1024_d 6.67814e-19 $X=7.385 $Y=1.3 $X2=0
+ $Y2=0
cc_782 N_A_1226_296#_M1014_g N_VGND_c_1551_n 0.00497913f $X=6.28 $Y=0.83 $X2=0
+ $Y2=0
cc_783 N_A_1226_296#_c_1018_n N_VGND_c_1551_n 0.00623301f $X=7.015 $Y=0.88 $X2=0
+ $Y2=0
cc_784 N_A_1226_296#_c_1019_n N_VGND_c_1551_n 0.0342287f $X=7.055 $Y=0.515 $X2=0
+ $Y2=0
cc_785 N_A_1226_296#_M1000_g N_VGND_c_1552_n 0.00336931f $X=7.73 $Y=0.74 $X2=0
+ $Y2=0
cc_786 N_A_1226_296#_c_1018_n N_VGND_c_1552_n 0.0081203f $X=7.015 $Y=0.88 $X2=0
+ $Y2=0
cc_787 N_A_1226_296#_c_1019_n N_VGND_c_1552_n 0.0136308f $X=7.055 $Y=0.515 $X2=0
+ $Y2=0
cc_788 N_A_1226_296#_c_1022_n N_VGND_c_1552_n 0.00538728f $X=8.5 $Y=1.465 $X2=0
+ $Y2=0
cc_789 N_A_1226_296#_M1000_g N_VGND_c_1553_n 0.00461464f $X=7.73 $Y=0.74 $X2=0
+ $Y2=0
cc_790 N_A_1226_296#_M1004_g N_VGND_c_1553_n 0.00434272f $X=8.2 $Y=0.74 $X2=0
+ $Y2=0
cc_791 N_A_1226_296#_M1004_g N_VGND_c_1554_n 0.00291539f $X=8.2 $Y=0.74 $X2=0
+ $Y2=0
cc_792 N_A_1226_296#_M1012_g N_VGND_c_1554_n 0.00414238f $X=8.65 $Y=0.74 $X2=0
+ $Y2=0
cc_793 N_A_1226_296#_M1030_g N_VGND_c_1556_n 0.00647072f $X=9.08 $Y=0.74 $X2=0
+ $Y2=0
cc_794 N_A_1226_296#_M1014_g N_VGND_c_1561_n 0.00417968f $X=6.28 $Y=0.83 $X2=0
+ $Y2=0
cc_795 N_A_1226_296#_c_1019_n N_VGND_c_1562_n 0.0110584f $X=7.055 $Y=0.515 $X2=0
+ $Y2=0
cc_796 N_A_1226_296#_M1012_g N_VGND_c_1563_n 0.00434272f $X=8.65 $Y=0.74 $X2=0
+ $Y2=0
cc_797 N_A_1226_296#_M1030_g N_VGND_c_1563_n 0.00428607f $X=9.08 $Y=0.74 $X2=0
+ $Y2=0
cc_798 N_A_1226_296#_M1014_g N_VGND_c_1569_n 0.00470816f $X=6.28 $Y=0.83 $X2=0
+ $Y2=0
cc_799 N_A_1226_296#_M1000_g N_VGND_c_1569_n 0.0090797f $X=7.73 $Y=0.74 $X2=0
+ $Y2=0
cc_800 N_A_1226_296#_M1004_g N_VGND_c_1569_n 0.00820868f $X=8.2 $Y=0.74 $X2=0
+ $Y2=0
cc_801 N_A_1226_296#_M1012_g N_VGND_c_1569_n 0.00820929f $X=8.65 $Y=0.74 $X2=0
+ $Y2=0
cc_802 N_A_1226_296#_M1030_g N_VGND_c_1569_n 0.00805681f $X=9.08 $Y=0.74 $X2=0
+ $Y2=0
cc_803 N_A_1226_296#_c_1019_n N_VGND_c_1569_n 0.00915653f $X=7.055 $Y=0.515
+ $X2=0 $Y2=0
cc_804 N_A_1034_424#_c_1188_n N_VPWR_c_1291_n 0.00606538f $X=6.76 $Y=2.045 $X2=0
+ $Y2=0
cc_805 N_A_1034_424#_c_1192_n N_VPWR_c_1292_n 0.0110424f $X=7.21 $Y=2.045 $X2=0
+ $Y2=0
cc_806 N_A_1034_424#_c_1188_n N_VPWR_c_1300_n 0.00445602f $X=6.76 $Y=2.045 $X2=0
+ $Y2=0
cc_807 N_A_1034_424#_c_1192_n N_VPWR_c_1300_n 0.00445602f $X=7.21 $Y=2.045 $X2=0
+ $Y2=0
cc_808 N_A_1034_424#_c_1188_n N_VPWR_c_1287_n 0.00857473f $X=6.76 $Y=2.045 $X2=0
+ $Y2=0
cc_809 N_A_1034_424#_c_1192_n N_VPWR_c_1287_n 0.00858495f $X=7.21 $Y=2.045 $X2=0
+ $Y2=0
cc_810 N_A_1034_424#_c_1190_n N_Q_c_1474_n 2.97544e-19 $X=7.135 $Y=1.97 $X2=0
+ $Y2=0
cc_811 N_A_1034_424#_c_1192_n N_Q_c_1474_n 2.69808e-19 $X=7.21 $Y=2.045 $X2=0
+ $Y2=0
cc_812 N_A_1034_424#_c_1190_n N_Q_c_1476_n 2.97674e-19 $X=7.135 $Y=1.97 $X2=0
+ $Y2=0
cc_813 N_A_1034_424#_c_1182_n N_VGND_c_1551_n 0.00255519f $X=7.27 $Y=1.22 $X2=0
+ $Y2=0
cc_814 N_A_1034_424#_c_1185_n N_VGND_c_1551_n 0.0205361f $X=6.63 $Y=1.225 $X2=0
+ $Y2=0
cc_815 N_A_1034_424#_c_1182_n N_VGND_c_1552_n 0.00860377f $X=7.27 $Y=1.22 $X2=0
+ $Y2=0
cc_816 N_A_1034_424#_c_1182_n N_VGND_c_1562_n 0.00383152f $X=7.27 $Y=1.22 $X2=0
+ $Y2=0
cc_817 N_A_1034_424#_c_1182_n N_VGND_c_1569_n 0.00762539f $X=7.27 $Y=1.22 $X2=0
+ $Y2=0
cc_818 N_VPWR_c_1292_n N_Q_c_1474_n 0.0617165f $X=7.52 $Y=2.225 $X2=0 $Y2=0
cc_819 N_VPWR_c_1293_n N_Q_c_1474_n 0.014552f $X=8.335 $Y=3.33 $X2=0 $Y2=0
cc_820 N_VPWR_c_1294_n N_Q_c_1474_n 0.0547423f $X=8.42 $Y=2.305 $X2=0 $Y2=0
cc_821 N_VPWR_c_1287_n N_Q_c_1474_n 0.0119791f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_822 N_VPWR_M1007_s N_Q_c_1475_n 0.00247267f $X=8.27 $Y=1.84 $X2=0 $Y2=0
cc_823 N_VPWR_c_1294_n N_Q_c_1475_n 0.0136682f $X=8.42 $Y=2.305 $X2=0 $Y2=0
cc_824 N_VPWR_c_1296_n Q 0.0107081f $X=9.32 $Y=1.985 $X2=0 $Y2=0
cc_825 N_VPWR_c_1294_n Q 0.0547423f $X=8.42 $Y=2.305 $X2=0 $Y2=0
cc_826 N_VPWR_c_1296_n Q 0.0677182f $X=9.32 $Y=1.985 $X2=0 $Y2=0
cc_827 N_VPWR_c_1301_n Q 0.014552f $X=9.235 $Y=3.33 $X2=0 $Y2=0
cc_828 N_VPWR_c_1287_n Q 0.0119791f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_829 N_Q_c_1469_n N_VGND_M1004_s 0.0025002f $X=8.7 $Y=1.045 $X2=0 $Y2=0
cc_830 N_Q_c_1468_n N_VGND_c_1552_n 0.00158095f $X=7.985 $Y=0.515 $X2=0 $Y2=0
cc_831 N_Q_c_1468_n N_VGND_c_1553_n 0.0145639f $X=7.985 $Y=0.515 $X2=0 $Y2=0
cc_832 N_Q_c_1468_n N_VGND_c_1554_n 0.0164567f $X=7.985 $Y=0.515 $X2=0 $Y2=0
cc_833 N_Q_c_1469_n N_VGND_c_1554_n 0.0135869f $X=8.7 $Y=1.045 $X2=0 $Y2=0
cc_834 N_Q_c_1471_n N_VGND_c_1554_n 0.028721f $X=8.865 $Y=0.515 $X2=0 $Y2=0
cc_835 N_Q_c_1471_n N_VGND_c_1556_n 0.0231198f $X=8.865 $Y=0.515 $X2=0 $Y2=0
cc_836 N_Q_c_1473_n N_VGND_c_1556_n 0.00774108f $X=8.867 $Y=1.045 $X2=0 $Y2=0
cc_837 N_Q_c_1471_n N_VGND_c_1563_n 0.0147003f $X=8.865 $Y=0.515 $X2=0 $Y2=0
cc_838 N_Q_c_1468_n N_VGND_c_1569_n 0.0119984f $X=7.985 $Y=0.515 $X2=0 $Y2=0
cc_839 N_Q_c_1471_n N_VGND_c_1569_n 0.0120432f $X=8.865 $Y=0.515 $X2=0 $Y2=0
