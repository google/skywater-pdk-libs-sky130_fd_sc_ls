* File: sky130_fd_sc_ls__a21oi_4.pex.spice
* Created: Wed Sep  2 10:49:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__A21OI_4%A2 1 3 6 8 10 13 15 17 20 22 24 27 29 30 31
+ 47
c86 31 0 1.12387e-19 $X=2.16 $Y=1.665
c87 27 0 7.99896e-20 $X=2.05 $Y=0.74
r88 47 48 0.651351 $w=3.7e-07 $l=5e-09 $layer=POLY_cond $X=2.045 $Y=1.557
+ $X2=2.05 $Y2=1.557
r89 45 47 9.77027 $w=3.7e-07 $l=7.5e-08 $layer=POLY_cond $X=1.97 $Y=1.557
+ $X2=2.045 $Y2=1.557
r90 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.97
+ $Y=1.515 $X2=1.97 $Y2=1.515
r91 43 45 45.5946 $w=3.7e-07 $l=3.5e-07 $layer=POLY_cond $X=1.62 $Y=1.557
+ $X2=1.97 $Y2=1.557
r92 42 43 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=1.595 $Y=1.557
+ $X2=1.62 $Y2=1.557
r93 41 42 52.7595 $w=3.7e-07 $l=4.05e-07 $layer=POLY_cond $X=1.19 $Y=1.557
+ $X2=1.595 $Y2=1.557
r94 40 41 5.86216 $w=3.7e-07 $l=4.5e-08 $layer=POLY_cond $X=1.145 $Y=1.557
+ $X2=1.19 $Y2=1.557
r95 38 40 25.4027 $w=3.7e-07 $l=1.95e-07 $layer=POLY_cond $X=0.95 $Y=1.557
+ $X2=1.145 $Y2=1.557
r96 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.95
+ $Y=1.515 $X2=0.95 $Y2=1.515
r97 36 38 24.7514 $w=3.7e-07 $l=1.9e-07 $layer=POLY_cond $X=0.76 $Y=1.557
+ $X2=0.95 $Y2=1.557
r98 35 36 8.46757 $w=3.7e-07 $l=6.5e-08 $layer=POLY_cond $X=0.695 $Y=1.557
+ $X2=0.76 $Y2=1.557
r99 31 46 5.09219 $w=4.28e-07 $l=1.9e-07 $layer=LI1_cond $X=2.16 $Y=1.565
+ $X2=1.97 $Y2=1.565
r100 30 46 7.77229 $w=4.28e-07 $l=2.9e-07 $layer=LI1_cond $X=1.68 $Y=1.565
+ $X2=1.97 $Y2=1.565
r101 29 30 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.565
+ $X2=1.68 $Y2=1.565
r102 29 39 6.70025 $w=4.28e-07 $l=2.5e-07 $layer=LI1_cond $X=1.2 $Y=1.565
+ $X2=0.95 $Y2=1.565
r103 25 48 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.05 $Y=1.35
+ $X2=2.05 $Y2=1.557
r104 25 27 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.05 $Y=1.35
+ $X2=2.05 $Y2=0.74
r105 22 47 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.045 $Y=1.765
+ $X2=2.045 $Y2=1.557
r106 22 24 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.045 $Y=1.765
+ $X2=2.045 $Y2=2.4
r107 18 43 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.62 $Y=1.35
+ $X2=1.62 $Y2=1.557
r108 18 20 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.62 $Y=1.35
+ $X2=1.62 $Y2=0.74
r109 15 42 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.595 $Y=1.765
+ $X2=1.595 $Y2=1.557
r110 15 17 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.595 $Y=1.765
+ $X2=1.595 $Y2=2.4
r111 11 41 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.19 $Y=1.35
+ $X2=1.19 $Y2=1.557
r112 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.19 $Y=1.35
+ $X2=1.19 $Y2=0.74
r113 8 40 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.145 $Y=1.765
+ $X2=1.145 $Y2=1.557
r114 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.145 $Y=1.765
+ $X2=1.145 $Y2=2.4
r115 4 36 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.76 $Y=1.35
+ $X2=0.76 $Y2=1.557
r116 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.76 $Y=1.35 $X2=0.76
+ $Y2=0.74
r117 1 35 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.695 $Y=1.765
+ $X2=0.695 $Y2=1.557
r118 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.695 $Y=1.765
+ $X2=0.695 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__A21OI_4%A1 3 5 7 10 12 14 17 19 21 24 26 28 29 30 43
+ 44
c87 44 0 9.44733e-20 $X=3.77 $Y=1.515
c88 26 0 1.59665e-20 $X=3.845 $Y=1.765
c89 17 0 6.95413e-20 $X=3.34 $Y=0.74
c90 10 0 6.95443e-20 $X=2.91 $Y=0.74
c91 5 0 1.12387e-19 $X=2.495 $Y=1.765
c92 3 0 1.9142e-19 $X=2.48 $Y=0.74
r93 43 45 9.77027 $w=3.7e-07 $l=7.5e-08 $layer=POLY_cond $X=3.77 $Y=1.557
+ $X2=3.845 $Y2=1.557
r94 43 44 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.77
+ $Y=1.515 $X2=3.77 $Y2=1.515
r95 41 43 48.8514 $w=3.7e-07 $l=3.75e-07 $layer=POLY_cond $X=3.395 $Y=1.557
+ $X2=3.77 $Y2=1.557
r96 40 41 7.16487 $w=3.7e-07 $l=5.5e-08 $layer=POLY_cond $X=3.34 $Y=1.557
+ $X2=3.395 $Y2=1.557
r97 38 40 32.5676 $w=3.7e-07 $l=2.5e-07 $layer=POLY_cond $X=3.09 $Y=1.557
+ $X2=3.34 $Y2=1.557
r98 38 39 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.09
+ $Y=1.515 $X2=3.09 $Y2=1.515
r99 36 38 18.8892 $w=3.7e-07 $l=1.45e-07 $layer=POLY_cond $X=2.945 $Y=1.557
+ $X2=3.09 $Y2=1.557
r100 35 36 4.55946 $w=3.7e-07 $l=3.5e-08 $layer=POLY_cond $X=2.91 $Y=1.557
+ $X2=2.945 $Y2=1.557
r101 34 35 54.0622 $w=3.7e-07 $l=4.15e-07 $layer=POLY_cond $X=2.495 $Y=1.557
+ $X2=2.91 $Y2=1.557
r102 33 34 1.95405 $w=3.7e-07 $l=1.5e-08 $layer=POLY_cond $X=2.48 $Y=1.557
+ $X2=2.495 $Y2=1.557
r103 30 44 4.55617 $w=4.28e-07 $l=1.7e-07 $layer=LI1_cond $X=3.6 $Y=1.565
+ $X2=3.77 $Y2=1.565
r104 29 30 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=3.12 $Y=1.565
+ $X2=3.6 $Y2=1.565
r105 29 39 0.80403 $w=4.28e-07 $l=3e-08 $layer=LI1_cond $X=3.12 $Y=1.565
+ $X2=3.09 $Y2=1.565
r106 26 45 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.845 $Y=1.765
+ $X2=3.845 $Y2=1.557
r107 26 28 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.845 $Y=1.765
+ $X2=3.845 $Y2=2.4
r108 22 43 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.77 $Y=1.35
+ $X2=3.77 $Y2=1.557
r109 22 24 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.77 $Y=1.35
+ $X2=3.77 $Y2=0.74
r110 19 41 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.395 $Y=1.765
+ $X2=3.395 $Y2=1.557
r111 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.395 $Y=1.765
+ $X2=3.395 $Y2=2.4
r112 15 40 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.34 $Y=1.35
+ $X2=3.34 $Y2=1.557
r113 15 17 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.34 $Y=1.35
+ $X2=3.34 $Y2=0.74
r114 12 36 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.945 $Y=1.765
+ $X2=2.945 $Y2=1.557
r115 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.945 $Y=1.765
+ $X2=2.945 $Y2=2.4
r116 8 35 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.91 $Y=1.35
+ $X2=2.91 $Y2=1.557
r117 8 10 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.91 $Y=1.35
+ $X2=2.91 $Y2=0.74
r118 5 34 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.495 $Y=1.765
+ $X2=2.495 $Y2=1.557
r119 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.495 $Y=1.765
+ $X2=2.495 $Y2=2.4
r120 1 33 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.48 $Y=1.35
+ $X2=2.48 $Y2=1.557
r121 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.48 $Y=1.35 $X2=2.48
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__A21OI_4%B1 1 3 4 6 9 11 13 16 18 19 20 22 23 25 26
+ 37
c65 37 0 1.59665e-20 $X=5.08 $Y=1.515
c66 1 0 9.44733e-20 $X=4.295 $Y=1.765
r67 38 39 1.97003 $w=3.67e-07 $l=1.5e-08 $layer=POLY_cond $X=5.195 $Y=1.557
+ $X2=5.21 $Y2=1.557
r68 36 38 15.1035 $w=3.67e-07 $l=1.15e-07 $layer=POLY_cond $X=5.08 $Y=1.557
+ $X2=5.195 $Y2=1.557
r69 36 37 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=5.08
+ $Y=1.515 $X2=5.08 $Y2=1.515
r70 34 36 39.4005 $w=3.67e-07 $l=3e-07 $layer=POLY_cond $X=4.78 $Y=1.557
+ $X2=5.08 $Y2=1.557
r71 33 34 4.59673 $w=3.67e-07 $l=3.5e-08 $layer=POLY_cond $X=4.745 $Y=1.557
+ $X2=4.78 $Y2=1.557
r72 31 33 45.3106 $w=3.67e-07 $l=3.45e-07 $layer=POLY_cond $X=4.4 $Y=1.557
+ $X2=4.745 $Y2=1.557
r73 31 32 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=4.4
+ $Y=1.515 $X2=4.4 $Y2=1.515
r74 29 31 13.7902 $w=3.67e-07 $l=1.05e-07 $layer=POLY_cond $X=4.295 $Y=1.557
+ $X2=4.4 $Y2=1.557
r75 26 37 1.07204 $w=4.28e-07 $l=4e-08 $layer=LI1_cond $X=5.04 $Y=1.565 $X2=5.08
+ $Y2=1.565
r76 25 26 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=4.56 $Y=1.565
+ $X2=5.04 $Y2=1.565
r77 25 32 4.28816 $w=4.28e-07 $l=1.6e-07 $layer=LI1_cond $X=4.56 $Y=1.565
+ $X2=4.4 $Y2=1.565
r78 20 23 64.3434 $w=1.8e-07 $l=1.6e-07 $layer=POLY_cond $X=5.645 $Y=1.765
+ $X2=5.645 $Y2=1.605
r79 20 22 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.645 $Y=1.765
+ $X2=5.645 $Y2=2.4
r80 19 39 27.1901 $w=3.67e-07 $l=9.60469e-08 $layer=POLY_cond $X=5.285 $Y=1.605
+ $X2=5.21 $Y2=1.557
r81 18 23 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=5.555 $Y=1.605
+ $X2=5.645 $Y2=1.605
r82 18 19 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=5.555 $Y=1.605
+ $X2=5.285 $Y2=1.605
r83 14 39 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.21 $Y=1.35 $X2=5.21
+ $Y2=1.557
r84 14 16 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.21 $Y=1.35
+ $X2=5.21 $Y2=0.74
r85 11 38 23.77 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=5.195 $Y=1.765
+ $X2=5.195 $Y2=1.557
r86 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.195 $Y=1.765
+ $X2=5.195 $Y2=2.4
r87 7 34 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.78 $Y=1.35 $X2=4.78
+ $Y2=1.557
r88 7 9 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.78 $Y=1.35 $X2=4.78
+ $Y2=0.74
r89 4 33 23.77 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=4.745 $Y=1.765
+ $X2=4.745 $Y2=1.557
r90 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.745 $Y=1.765
+ $X2=4.745 $Y2=2.4
r91 1 29 23.77 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=4.295 $Y=1.765
+ $X2=4.295 $Y2=1.557
r92 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.295 $Y=1.765
+ $X2=4.295 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__A21OI_4%A_69_368# 1 2 3 4 5 6 7 22 24 26 30 32 34 35
+ 38 40 44 46 47 48 49 52 54 58 65 68 70 73
r107 58 61 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=5.91 $Y=1.985
+ $X2=5.91 $Y2=2.815
r108 56 61 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=5.91 $Y=2.905
+ $X2=5.91 $Y2=2.815
r109 55 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.055 $Y=2.99
+ $X2=4.97 $Y2=2.99
r110 54 56 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.785 $Y=2.99
+ $X2=5.91 $Y2=2.905
r111 54 55 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=5.785 $Y=2.99
+ $X2=5.055 $Y2=2.99
r112 50 73 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.97 $Y=2.905
+ $X2=4.97 $Y2=2.99
r113 50 52 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=4.97 $Y=2.905
+ $X2=4.97 $Y2=2.455
r114 48 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.885 $Y=2.99
+ $X2=4.97 $Y2=2.99
r115 48 49 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=4.885 $Y=2.99
+ $X2=4.155 $Y2=2.99
r116 47 49 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.03 $Y=2.905
+ $X2=4.155 $Y2=2.99
r117 46 72 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.03 $Y=2.46
+ $X2=4.03 $Y2=2.375
r118 46 47 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=4.03 $Y=2.46
+ $X2=4.03 $Y2=2.905
r119 45 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.335 $Y=2.375
+ $X2=3.17 $Y2=2.375
r120 44 72 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.905 $Y=2.375
+ $X2=4.03 $Y2=2.375
r121 44 45 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=3.905 $Y=2.375
+ $X2=3.335 $Y2=2.375
r122 41 68 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.355 $Y=2.375
+ $X2=2.23 $Y2=2.375
r123 40 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.005 $Y=2.375
+ $X2=3.17 $Y2=2.375
r124 40 41 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=3.005 $Y=2.375
+ $X2=2.355 $Y2=2.375
r125 36 68 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.23 $Y=2.46
+ $X2=2.23 $Y2=2.375
r126 36 38 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=2.23 $Y=2.46
+ $X2=2.23 $Y2=2.465
r127 35 68 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.23 $Y=2.29
+ $X2=2.23 $Y2=2.375
r128 34 67 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.23 $Y=2.12
+ $X2=2.23 $Y2=2.035
r129 34 35 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=2.23 $Y=2.12
+ $X2=2.23 $Y2=2.29
r130 33 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.535 $Y=2.035
+ $X2=1.37 $Y2=2.035
r131 32 67 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.105 $Y=2.035
+ $X2=2.23 $Y2=2.035
r132 32 33 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=2.105 $Y=2.035
+ $X2=1.535 $Y2=2.035
r133 28 65 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.37 $Y=2.12
+ $X2=1.37 $Y2=2.035
r134 28 30 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=1.37 $Y=2.12
+ $X2=1.37 $Y2=2.815
r135 27 63 3.99177 $w=1.7e-07 $l=1.5411e-07 $layer=LI1_cond $X=0.555 $Y=2.035
+ $X2=0.43 $Y2=1.97
r136 26 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.205 $Y=2.035
+ $X2=1.37 $Y2=2.035
r137 26 27 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.205 $Y=2.035
+ $X2=0.555 $Y2=2.035
r138 22 63 3.1514 $w=2.5e-07 $l=1.5e-07 $layer=LI1_cond $X=0.43 $Y=2.12 $X2=0.43
+ $Y2=1.97
r139 22 24 12.9074 $w=2.48e-07 $l=2.8e-07 $layer=LI1_cond $X=0.43 $Y=2.12
+ $X2=0.43 $Y2=2.4
r140 7 61 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=5.72
+ $Y=1.84 $X2=5.87 $Y2=2.815
r141 7 58 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=5.72
+ $Y=1.84 $X2=5.87 $Y2=1.985
r142 6 52 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=4.82
+ $Y=1.84 $X2=4.97 $Y2=2.455
r143 5 72 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=3.92
+ $Y=1.84 $X2=4.07 $Y2=2.455
r144 4 70 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=3.02
+ $Y=1.84 $X2=3.17 $Y2=2.455
r145 3 67 600 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=2.12
+ $Y=1.84 $X2=2.27 $Y2=2.115
r146 3 38 300 $w=1.7e-07 $l=6.95971e-07 $layer=licon1_PDIFF $count=2 $X=2.12
+ $Y=1.84 $X2=2.27 $Y2=2.465
r147 2 65 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=1.22
+ $Y=1.84 $X2=1.37 $Y2=2.115
r148 2 30 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.22
+ $Y=1.84 $X2=1.37 $Y2=2.815
r149 1 63 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.345
+ $Y=1.84 $X2=0.47 $Y2=1.985
r150 1 24 300 $w=1.7e-07 $l=6.19354e-07 $layer=licon1_PDIFF $count=2 $X=0.345
+ $Y=1.84 $X2=0.47 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__A21OI_4%VPWR 1 2 3 4 15 19 23 25 29 32 33 35 36 37
+ 46 55 56 59 62
r86 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r87 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r88 55 56 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r89 53 56 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.08 $Y=3.33 $X2=6
+ $Y2=3.33
r90 53 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r91 52 55 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.08 $Y=3.33 $X2=6
+ $Y2=3.33
r92 52 53 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r93 50 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.705 $Y=3.33
+ $X2=3.62 $Y2=3.33
r94 50 52 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=3.705 $Y=3.33
+ $X2=4.08 $Y2=3.33
r95 49 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r96 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r97 46 59 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.555 $Y=3.33
+ $X2=2.68 $Y2=3.33
r98 46 48 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=2.555 $Y=3.33
+ $X2=2.16 $Y2=3.33
r99 45 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r100 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r101 41 45 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r102 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r103 37 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r104 37 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r105 35 44 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=1.735 $Y=3.33
+ $X2=1.68 $Y2=3.33
r106 35 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.735 $Y=3.33
+ $X2=1.82 $Y2=3.33
r107 34 48 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.905 $Y=3.33
+ $X2=2.16 $Y2=3.33
r108 34 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.905 $Y=3.33
+ $X2=1.82 $Y2=3.33
r109 32 40 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=0.755 $Y=3.33
+ $X2=0.72 $Y2=3.33
r110 32 33 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.755 $Y=3.33
+ $X2=0.88 $Y2=3.33
r111 31 44 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=1.005 $Y=3.33
+ $X2=1.68 $Y2=3.33
r112 31 33 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.005 $Y=3.33
+ $X2=0.88 $Y2=3.33
r113 27 62 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.62 $Y=3.245
+ $X2=3.62 $Y2=3.33
r114 27 29 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=3.62 $Y=3.245
+ $X2=3.62 $Y2=2.805
r115 26 59 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.805 $Y=3.33
+ $X2=2.68 $Y2=3.33
r116 25 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.535 $Y=3.33
+ $X2=3.62 $Y2=3.33
r117 25 26 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=3.535 $Y=3.33
+ $X2=2.805 $Y2=3.33
r118 21 59 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.68 $Y=3.245
+ $X2=2.68 $Y2=3.33
r119 21 23 20.283 $w=2.48e-07 $l=4.4e-07 $layer=LI1_cond $X=2.68 $Y=3.245
+ $X2=2.68 $Y2=2.805
r120 17 36 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.82 $Y=3.245
+ $X2=1.82 $Y2=3.33
r121 17 19 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=1.82 $Y=3.245
+ $X2=1.82 $Y2=2.455
r122 13 33 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.88 $Y=3.245
+ $X2=0.88 $Y2=3.33
r123 13 15 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=0.88 $Y=3.245
+ $X2=0.88 $Y2=2.455
r124 4 29 600 $w=1.7e-07 $l=1.03729e-06 $layer=licon1_PDIFF $count=1 $X=3.47
+ $Y=1.84 $X2=3.62 $Y2=2.805
r125 3 23 600 $w=1.7e-07 $l=1.03729e-06 $layer=licon1_PDIFF $count=1 $X=2.57
+ $Y=1.84 $X2=2.72 $Y2=2.805
r126 2 19 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=1.67
+ $Y=1.84 $X2=1.82 $Y2=2.455
r127 1 15 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=0.77
+ $Y=1.84 $X2=0.92 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_LS__A21OI_4%Y 1 2 3 4 5 6 19 20 21 29 31 33 39 43 44 46
+ 47 48 49 54
c101 47 0 7.99896e-20 $X=2.64 $Y=0.925
r102 48 49 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.64 $Y=1.295
+ $X2=2.64 $Y2=1.665
r103 48 57 5.76222 $w=2.28e-07 $l=1.15e-07 $layer=LI1_cond $X=2.64 $Y=1.295
+ $X2=2.64 $Y2=1.18
r104 47 54 6.14322 $w=2.42e-07 $l=1.5e-07 $layer=LI1_cond $X=2.652 $Y=1.03
+ $X2=2.652 $Y2=0.88
r105 47 57 6.14322 $w=2.42e-07 $l=1.55885e-07 $layer=LI1_cond $X=2.652 $Y=1.03
+ $X2=2.64 $Y2=1.18
r106 47 54 0.956863 $w=2.55e-07 $l=2e-08 $layer=LI1_cond $X=2.652 $Y=0.86
+ $X2=2.652 $Y2=0.88
r107 41 49 14.2803 $w=2.28e-07 $l=2.85e-07 $layer=LI1_cond $X=2.64 $Y=1.95
+ $X2=2.64 $Y2=1.665
r108 37 39 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=5.465 $Y=1.01
+ $X2=5.465 $Y2=0.515
r109 34 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.685 $Y=2.035
+ $X2=4.52 $Y2=2.035
r110 33 46 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.255 $Y=2.035
+ $X2=5.42 $Y2=2.035
r111 33 34 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=5.255 $Y=2.035
+ $X2=4.685 $Y2=2.035
r112 32 44 5.43733 $w=2.35e-07 $l=1.5411e-07 $layer=LI1_cond $X=4.65 $Y=1.095
+ $X2=4.525 $Y2=1.03
r113 31 37 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.34 $Y=1.095
+ $X2=5.465 $Y2=1.01
r114 31 32 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.34 $Y=1.095
+ $X2=4.65 $Y2=1.095
r115 27 44 1.12072 $w=2.5e-07 $l=1.5e-07 $layer=LI1_cond $X=4.525 $Y=0.88
+ $X2=4.525 $Y2=1.03
r116 27 29 16.8257 $w=2.48e-07 $l=3.65e-07 $layer=LI1_cond $X=4.525 $Y=0.88
+ $X2=4.525 $Y2=0.515
r117 22 47 0.588783 $w=3e-07 $l=1.28e-07 $layer=LI1_cond $X=2.78 $Y=1.03
+ $X2=2.652 $Y2=1.03
r118 22 24 29.7714 $w=2.98e-07 $l=7.75e-07 $layer=LI1_cond $X=2.78 $Y=1.03
+ $X2=3.555 $Y2=1.03
r119 21 44 5.43733 $w=2.35e-07 $l=1.25e-07 $layer=LI1_cond $X=4.4 $Y=1.03
+ $X2=4.525 $Y2=1.03
r120 21 24 32.4605 $w=2.98e-07 $l=8.45e-07 $layer=LI1_cond $X=4.4 $Y=1.03
+ $X2=3.555 $Y2=1.03
r121 20 41 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=2.755 $Y=2.035
+ $X2=2.64 $Y2=1.95
r122 19 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.355 $Y=2.035
+ $X2=4.52 $Y2=2.035
r123 19 20 104.385 $w=1.68e-07 $l=1.6e-06 $layer=LI1_cond $X=4.355 $Y=2.035
+ $X2=2.755 $Y2=2.035
r124 6 46 300 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=2 $X=5.27
+ $Y=1.84 $X2=5.42 $Y2=2.115
r125 5 43 300 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=2 $X=4.37
+ $Y=1.84 $X2=4.52 $Y2=2.115
r126 4 39 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.285
+ $Y=0.37 $X2=5.425 $Y2=0.515
r127 3 29 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=4.44
+ $Y=0.37 $X2=4.565 $Y2=0.515
r128 2 24 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=3.415
+ $Y=0.37 $X2=3.555 $Y2=0.965
r129 1 47 182 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_NDIFF $count=1 $X=2.555
+ $Y=0.37 $X2=2.695 $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_LS__A21OI_4%A_84_74# 1 2 3 4 5 18 20 21 24 26 32 33 34
+ 36 37 42
c72 34 0 6.95443e-20 $X=3.82 $Y=0.34
c73 32 0 6.95413e-20 $X=2.96 $Y=0.34
r74 42 45 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=3.985 $Y=0.34
+ $X2=3.985 $Y2=0.53
r75 37 40 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=3.125 $Y=0.34
+ $X2=3.125 $Y2=0.53
r76 35 37 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.29 $Y=0.34
+ $X2=3.125 $Y2=0.34
r77 34 42 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.82 $Y=0.34
+ $X2=3.985 $Y2=0.34
r78 34 35 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.82 $Y=0.34
+ $X2=3.29 $Y2=0.34
r79 32 37 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.96 $Y=0.34
+ $X2=3.125 $Y2=0.34
r80 32 33 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=2.96 $Y=0.34
+ $X2=2.35 $Y2=0.34
r81 29 31 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=2.265 $Y=1.01
+ $X2=2.265 $Y2=0.515
r82 28 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.265 $Y=0.425
+ $X2=2.35 $Y2=0.34
r83 28 31 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=2.265 $Y=0.425
+ $X2=2.265 $Y2=0.515
r84 27 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.49 $Y=1.095
+ $X2=1.405 $Y2=1.095
r85 26 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.18 $Y=1.095
+ $X2=2.265 $Y2=1.01
r86 26 27 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.18 $Y=1.095
+ $X2=1.49 $Y2=1.095
r87 22 36 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.405 $Y=1.01
+ $X2=1.405 $Y2=1.095
r88 22 24 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=1.405 $Y=1.01
+ $X2=1.405 $Y2=0.515
r89 20 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.32 $Y=1.095
+ $X2=1.405 $Y2=1.095
r90 20 21 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.32 $Y=1.095
+ $X2=0.63 $Y2=1.095
r91 16 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.505 $Y=1.01
+ $X2=0.63 $Y2=1.095
r92 16 18 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=0.505 $Y=1.01
+ $X2=0.505 $Y2=0.515
r93 5 45 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=3.845
+ $Y=0.37 $X2=3.985 $Y2=0.53
r94 4 40 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=2.985
+ $Y=0.37 $X2=3.125 $Y2=0.53
r95 3 31 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.125
+ $Y=0.37 $X2=2.265 $Y2=0.515
r96 2 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.265
+ $Y=0.37 $X2=1.405 $Y2=0.515
r97 1 18 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.42
+ $Y=0.37 $X2=0.545 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__A21OI_4%VGND 1 2 3 12 14 18 22 24 25 26 32 42 43 46
+ 49
c69 18 0 1.9142e-19 $X=1.835 $Y=0.595
r70 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r71 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r72 43 50 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.04
+ $Y2=0
r73 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6 $Y2=0
r74 40 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.16 $Y=0 $X2=4.995
+ $Y2=0
r75 40 42 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=5.16 $Y=0 $X2=6
+ $Y2=0
r76 39 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r77 38 39 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r78 36 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r79 35 38 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=2.16 $Y=0 $X2=4.56
+ $Y2=0
r80 35 36 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r81 33 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2 $Y=0 $X2=1.835
+ $Y2=0
r82 33 35 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=2 $Y=0 $X2=2.16
+ $Y2=0
r83 32 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.83 $Y=0 $X2=4.995
+ $Y2=0
r84 32 38 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=4.83 $Y=0 $X2=4.56
+ $Y2=0
r85 30 47 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r86 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r87 26 39 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=3.12 $Y=0 $X2=4.56
+ $Y2=0
r88 26 36 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.16
+ $Y2=0
r89 24 29 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=0.81 $Y=0 $X2=0.72
+ $Y2=0
r90 24 25 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.81 $Y=0 $X2=0.975
+ $Y2=0
r91 20 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.995 $Y=0.085
+ $X2=4.995 $Y2=0
r92 20 22 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=4.995 $Y=0.085
+ $X2=4.995 $Y2=0.595
r93 16 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.835 $Y=0.085
+ $X2=1.835 $Y2=0
r94 16 18 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=1.835 $Y=0.085
+ $X2=1.835 $Y2=0.595
r95 15 25 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.14 $Y=0 $X2=0.975
+ $Y2=0
r96 14 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.67 $Y=0 $X2=1.835
+ $Y2=0
r97 14 15 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.67 $Y=0 $X2=1.14
+ $Y2=0
r98 10 25 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.975 $Y=0.085
+ $X2=0.975 $Y2=0
r99 10 12 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=0.975 $Y=0.085
+ $X2=0.975 $Y2=0.595
r100 3 22 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=4.855
+ $Y=0.37 $X2=4.995 $Y2=0.595
r101 2 18 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=1.695
+ $Y=0.37 $X2=1.835 $Y2=0.595
r102 1 12 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=0.835
+ $Y=0.37 $X2=0.975 $Y2=0.595
.ends

