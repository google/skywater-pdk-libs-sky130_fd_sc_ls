* File: sky130_fd_sc_ls__and4bb_2.pxi.spice
* Created: Wed Sep  2 10:56:10 2020
* 
x_PM_SKY130_FD_SC_LS__AND4BB_2%A_N N_A_N_M1015_g N_A_N_c_97_n N_A_N_M1000_g A_N
+ N_A_N_c_98_n PM_SKY130_FD_SC_LS__AND4BB_2%A_N
x_PM_SKY130_FD_SC_LS__AND4BB_2%A_27_74# N_A_27_74#_M1015_s N_A_27_74#_M1000_s
+ N_A_27_74#_c_133_n N_A_27_74#_M1014_g N_A_27_74#_M1002_g N_A_27_74#_c_128_n
+ N_A_27_74#_c_129_n N_A_27_74#_c_130_n N_A_27_74#_c_134_n N_A_27_74#_c_131_n
+ N_A_27_74#_c_136_n N_A_27_74#_c_137_n N_A_27_74#_c_132_n
+ PM_SKY130_FD_SC_LS__AND4BB_2%A_27_74#
x_PM_SKY130_FD_SC_LS__AND4BB_2%A_354_252# N_A_354_252#_M1005_d
+ N_A_354_252#_M1004_d N_A_354_252#_M1003_g N_A_354_252#_c_194_n
+ N_A_354_252#_c_203_n N_A_354_252#_M1009_g N_A_354_252#_c_195_n
+ N_A_354_252#_c_196_n N_A_354_252#_c_197_n N_A_354_252#_c_247_p
+ N_A_354_252#_c_228_p N_A_354_252#_c_232_p N_A_354_252#_c_284_p
+ N_A_354_252#_c_198_n N_A_354_252#_c_199_n N_A_354_252#_c_205_n
+ N_A_354_252#_c_206_n N_A_354_252#_c_207_n N_A_354_252#_c_288_p
+ N_A_354_252#_c_200_n N_A_354_252#_c_201_n
+ PM_SKY130_FD_SC_LS__AND4BB_2%A_354_252#
x_PM_SKY130_FD_SC_LS__AND4BB_2%C N_C_M1010_g N_C_c_310_n N_C_M1006_g C
+ PM_SKY130_FD_SC_LS__AND4BB_2%C
x_PM_SKY130_FD_SC_LS__AND4BB_2%D N_D_M1013_g N_D_c_344_n N_D_M1011_g D
+ PM_SKY130_FD_SC_LS__AND4BB_2%D
x_PM_SKY130_FD_SC_LS__AND4BB_2%A_225_82# N_A_225_82#_M1002_s N_A_225_82#_M1014_d
+ N_A_225_82#_M1006_d N_A_225_82#_M1001_g N_A_225_82#_c_385_n
+ N_A_225_82#_M1007_g N_A_225_82#_M1008_g N_A_225_82#_c_386_n
+ N_A_225_82#_M1012_g N_A_225_82#_c_380_n N_A_225_82#_c_381_n
+ N_A_225_82#_c_388_n N_A_225_82#_c_389_n N_A_225_82#_c_390_n
+ N_A_225_82#_c_391_n N_A_225_82#_c_392_n N_A_225_82#_c_382_n
+ N_A_225_82#_c_393_n N_A_225_82#_c_394_n N_A_225_82#_c_383_n
+ N_A_225_82#_c_384_n PM_SKY130_FD_SC_LS__AND4BB_2%A_225_82#
x_PM_SKY130_FD_SC_LS__AND4BB_2%B_N N_B_N_c_503_n N_B_N_M1004_g N_B_N_c_504_n
+ N_B_N_M1005_g B_N PM_SKY130_FD_SC_LS__AND4BB_2%B_N
x_PM_SKY130_FD_SC_LS__AND4BB_2%VPWR N_VPWR_M1000_d N_VPWR_M1009_d N_VPWR_M1011_d
+ N_VPWR_M1012_s N_VPWR_c_530_n N_VPWR_c_531_n N_VPWR_c_532_n N_VPWR_c_533_n
+ N_VPWR_c_534_n N_VPWR_c_535_n N_VPWR_c_536_n N_VPWR_c_537_n N_VPWR_c_538_n
+ N_VPWR_c_539_n VPWR N_VPWR_c_540_n N_VPWR_c_541_n N_VPWR_c_529_n
+ N_VPWR_c_543_n PM_SKY130_FD_SC_LS__AND4BB_2%VPWR
x_PM_SKY130_FD_SC_LS__AND4BB_2%X N_X_M1001_d N_X_M1007_d N_X_c_599_n X X X X
+ N_X_c_600_n PM_SKY130_FD_SC_LS__AND4BB_2%X
x_PM_SKY130_FD_SC_LS__AND4BB_2%VGND N_VGND_M1015_d N_VGND_M1013_d N_VGND_M1008_s
+ N_VGND_c_634_n N_VGND_c_635_n VGND N_VGND_c_636_n N_VGND_c_637_n
+ N_VGND_c_638_n N_VGND_c_639_n N_VGND_c_640_n N_VGND_c_641_n N_VGND_c_642_n
+ N_VGND_c_643_n PM_SKY130_FD_SC_LS__AND4BB_2%VGND
cc_1 VNB N_A_N_M1015_g 0.0555342f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.645
cc_2 VNB N_A_N_c_97_n 0.026968f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.885
cc_3 VNB N_A_N_c_98_n 0.00891974f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_4 VNB N_A_27_74#_M1002_g 0.0222037f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_5 VNB N_A_27_74#_c_128_n 0.0327895f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_6 VNB N_A_27_74#_c_129_n 0.00630734f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_27_74#_c_130_n 0.00985767f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_27_74#_c_131_n 0.0182802f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_27_74#_c_132_n 0.0501833f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_354_252#_c_194_n 0.00461139f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.615
cc_11 VNB N_A_354_252#_c_195_n 0.00340503f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_354_252#_c_196_n 0.0330202f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_354_252#_c_197_n 0.0244392f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_354_252#_c_198_n 0.00968485f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_354_252#_c_199_n 8.10761e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_354_252#_c_200_n 0.0205529f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_354_252#_c_201_n 0.0161531f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_C_M1010_g 0.0271198f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.645
cc_19 VNB N_C_c_310_n 0.0185033f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.885
cc_20 VNB C 0.00463605f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_21 VNB N_D_M1013_g 0.0299553f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.645
cc_22 VNB N_D_c_344_n 0.0261406f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.885
cc_23 VNB D 0.00272145f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_24 VNB N_A_225_82#_M1001_g 0.0243113f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_25 VNB N_A_225_82#_M1008_g 0.0210013f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_225_82#_c_380_n 0.00817637f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_225_82#_c_381_n 0.00423086f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_225_82#_c_382_n 0.00611436f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_225_82#_c_383_n 0.00307202f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_225_82#_c_384_n 0.0469531f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_B_N_c_503_n 0.066553f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.45
cc_32 VNB N_B_N_c_504_n 0.0234298f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB B_N 0.00853765f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=2.38
cc_34 VNB N_VPWR_c_529_n 0.223389f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_X_c_599_n 0.00239705f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_36 VNB N_X_c_600_n 0.00191711f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_634_n 0.0158429f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_38 VNB N_VGND_c_635_n 0.00992069f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_39 VNB N_VGND_c_636_n 0.0173909f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_637_n 0.063202f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_638_n 0.0282128f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_639_n 0.019529f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_640_n 0.35573f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_641_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_642_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_643_n 0.0208183f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VPB N_A_N_c_97_n 0.0503769f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.885
cc_48 VPB N_A_N_c_98_n 0.00783763f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.615
cc_49 VPB N_A_27_74#_c_133_n 0.019325f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=2.38
cc_50 VPB N_A_27_74#_c_134_n 0.00147287f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_51 VPB N_A_27_74#_c_131_n 0.00251227f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_A_27_74#_c_136_n 0.00494613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_A_27_74#_c_137_n 0.0391303f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_A_27_74#_c_132_n 0.0209288f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_A_354_252#_c_194_n 0.00916667f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.615
cc_56 VPB N_A_354_252#_c_203_n 0.0263296f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.615
cc_57 VPB N_A_354_252#_c_198_n 0.00192121f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_A_354_252#_c_205_n 0.0142544f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_A_354_252#_c_206_n 8.17396e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_A_354_252#_c_207_n 0.0337804f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_C_c_310_n 0.0361288f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.885
cc_62 VPB C 0.00464027f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_63 VPB N_D_c_344_n 0.0412215f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.885
cc_64 VPB D 0.00175937f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_65 VPB N_A_225_82#_c_385_n 0.0176323f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_A_225_82#_c_386_n 0.0161104f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_A_225_82#_c_381_n 0.00675668f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_A_225_82#_c_388_n 0.00334339f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_A_225_82#_c_389_n 0.010143f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_A_225_82#_c_390_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_A_225_82#_c_391_n 0.00735735f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_A_225_82#_c_392_n 0.00283301f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_A_225_82#_c_393_n 0.00694775f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_A_225_82#_c_394_n 0.00589681f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_A_225_82#_c_384_n 0.0264158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_B_N_c_503_n 0.0298923f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.45
cc_77 VPB N_VPWR_c_530_n 0.0125615f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_531_n 0.00990292f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_532_n 0.00998098f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_533_n 0.0190281f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_534_n 0.025094f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_535_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_536_n 0.0229908f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_537_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_538_n 0.0237111f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_539_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_540_n 0.0276061f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_541_n 0.0217627f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_529_n 0.10744f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_543_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB X 0.00105619f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_92 VPB X 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_X_c_600_n 0.00131273f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 N_A_N_c_97_n N_A_27_74#_c_133_n 0.0156621f $X=0.6 $Y=1.885 $X2=0 $Y2=0
cc_95 N_A_N_M1015_g N_A_27_74#_c_128_n 0.0108396f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_96 N_A_N_M1015_g N_A_27_74#_c_129_n 0.017498f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_97 N_A_N_c_97_n N_A_27_74#_c_129_n 0.00436366f $X=0.6 $Y=1.885 $X2=0 $Y2=0
cc_98 N_A_N_c_98_n N_A_27_74#_c_129_n 0.0133796f $X=0.385 $Y=1.615 $X2=0 $Y2=0
cc_99 N_A_N_c_97_n N_A_27_74#_c_130_n 0.00337787f $X=0.6 $Y=1.885 $X2=0 $Y2=0
cc_100 N_A_N_c_98_n N_A_27_74#_c_130_n 0.0206322f $X=0.385 $Y=1.615 $X2=0 $Y2=0
cc_101 N_A_N_c_97_n N_A_27_74#_c_134_n 0.0135008f $X=0.6 $Y=1.885 $X2=0 $Y2=0
cc_102 N_A_N_c_98_n N_A_27_74#_c_134_n 6.80235e-19 $X=0.385 $Y=1.615 $X2=0 $Y2=0
cc_103 N_A_N_M1015_g N_A_27_74#_c_131_n 0.0048164f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_104 N_A_N_c_97_n N_A_27_74#_c_131_n 0.00192367f $X=0.6 $Y=1.885 $X2=0 $Y2=0
cc_105 N_A_N_c_98_n N_A_27_74#_c_131_n 0.0154119f $X=0.385 $Y=1.615 $X2=0 $Y2=0
cc_106 N_A_N_c_97_n N_A_27_74#_c_136_n 0.00523982f $X=0.6 $Y=1.885 $X2=0 $Y2=0
cc_107 N_A_N_c_98_n N_A_27_74#_c_136_n 0.0069965f $X=0.385 $Y=1.615 $X2=0 $Y2=0
cc_108 N_A_N_c_97_n N_A_27_74#_c_137_n 0.0211541f $X=0.6 $Y=1.885 $X2=0 $Y2=0
cc_109 N_A_N_c_98_n N_A_27_74#_c_137_n 0.0278035f $X=0.385 $Y=1.615 $X2=0 $Y2=0
cc_110 N_A_N_M1015_g N_A_27_74#_c_132_n 0.00318303f $X=0.495 $Y=0.645 $X2=0
+ $Y2=0
cc_111 N_A_N_c_97_n N_A_27_74#_c_132_n 0.0146002f $X=0.6 $Y=1.885 $X2=0 $Y2=0
cc_112 N_A_N_M1015_g N_A_225_82#_c_380_n 0.00139595f $X=0.495 $Y=0.645 $X2=0
+ $Y2=0
cc_113 N_A_N_M1015_g N_A_225_82#_c_382_n 0.00476143f $X=0.495 $Y=0.645 $X2=0
+ $Y2=0
cc_114 N_A_N_c_97_n N_VPWR_c_530_n 0.00794677f $X=0.6 $Y=1.885 $X2=0 $Y2=0
cc_115 N_A_N_c_97_n N_VPWR_c_534_n 0.00458031f $X=0.6 $Y=1.885 $X2=0 $Y2=0
cc_116 N_A_N_c_97_n N_VPWR_c_529_n 0.0049649f $X=0.6 $Y=1.885 $X2=0 $Y2=0
cc_117 N_A_N_M1015_g N_VGND_c_634_n 0.018223f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_118 N_A_N_M1015_g N_VGND_c_636_n 0.00383152f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_119 N_A_N_M1015_g N_VGND_c_640_n 0.00761198f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_120 N_A_27_74#_c_132_n N_A_354_252#_c_194_n 0.00416622f $X=1.17 $Y=1.612
+ $X2=0 $Y2=0
cc_121 N_A_27_74#_c_133_n N_A_354_252#_c_203_n 0.0162053f $X=1.17 $Y=1.885 $X2=0
+ $Y2=0
cc_122 N_A_27_74#_M1002_g N_A_354_252#_c_195_n 5.41695e-19 $X=1.485 $Y=0.78
+ $X2=0 $Y2=0
cc_123 N_A_27_74#_M1002_g N_A_354_252#_c_196_n 0.0143574f $X=1.485 $Y=0.78 $X2=0
+ $Y2=0
cc_124 N_A_27_74#_c_132_n N_A_354_252#_c_196_n 0.00175421f $X=1.17 $Y=1.612
+ $X2=0 $Y2=0
cc_125 N_A_27_74#_M1002_g N_A_354_252#_c_201_n 0.0510069f $X=1.485 $Y=0.78 $X2=0
+ $Y2=0
cc_126 N_A_27_74#_M1002_g N_A_225_82#_c_380_n 0.0124106f $X=1.485 $Y=0.78 $X2=0
+ $Y2=0
cc_127 N_A_27_74#_c_133_n N_A_225_82#_c_381_n 6.15178e-19 $X=1.17 $Y=1.885 $X2=0
+ $Y2=0
cc_128 N_A_27_74#_M1002_g N_A_225_82#_c_381_n 0.00481006f $X=1.485 $Y=0.78 $X2=0
+ $Y2=0
cc_129 N_A_27_74#_c_131_n N_A_225_82#_c_381_n 0.0310645f $X=0.85 $Y=1.67 $X2=0
+ $Y2=0
cc_130 N_A_27_74#_c_136_n N_A_225_82#_c_381_n 0.00959708f $X=0.85 $Y=1.95 $X2=0
+ $Y2=0
cc_131 N_A_27_74#_c_132_n N_A_225_82#_c_381_n 0.0106853f $X=1.17 $Y=1.612 $X2=0
+ $Y2=0
cc_132 N_A_27_74#_c_133_n N_A_225_82#_c_388_n 0.011494f $X=1.17 $Y=1.885 $X2=0
+ $Y2=0
cc_133 N_A_27_74#_M1002_g N_A_225_82#_c_382_n 0.00559356f $X=1.485 $Y=0.78 $X2=0
+ $Y2=0
cc_134 N_A_27_74#_c_131_n N_A_225_82#_c_382_n 0.0185168f $X=0.85 $Y=1.67 $X2=0
+ $Y2=0
cc_135 N_A_27_74#_c_132_n N_A_225_82#_c_382_n 0.00737103f $X=1.17 $Y=1.612 $X2=0
+ $Y2=0
cc_136 N_A_27_74#_c_133_n N_A_225_82#_c_393_n 0.00242489f $X=1.17 $Y=1.885 $X2=0
+ $Y2=0
cc_137 N_A_27_74#_c_134_n N_A_225_82#_c_393_n 0.00692332f $X=0.765 $Y=2.035
+ $X2=0 $Y2=0
cc_138 N_A_27_74#_c_136_n N_A_225_82#_c_393_n 3.58645e-19 $X=0.85 $Y=1.95 $X2=0
+ $Y2=0
cc_139 N_A_27_74#_c_134_n N_VPWR_M1000_d 0.00652706f $X=0.765 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_140 N_A_27_74#_c_133_n N_VPWR_c_530_n 0.0181079f $X=1.17 $Y=1.885 $X2=0 $Y2=0
cc_141 N_A_27_74#_c_134_n N_VPWR_c_530_n 0.0138849f $X=0.765 $Y=2.035 $X2=0
+ $Y2=0
cc_142 N_A_27_74#_c_131_n N_VPWR_c_530_n 0.00417773f $X=0.85 $Y=1.67 $X2=0 $Y2=0
cc_143 N_A_27_74#_c_137_n N_VPWR_c_530_n 0.0316073f $X=0.375 $Y=2.115 $X2=0
+ $Y2=0
cc_144 N_A_27_74#_c_132_n N_VPWR_c_530_n 7.23795e-19 $X=1.17 $Y=1.612 $X2=0
+ $Y2=0
cc_145 N_A_27_74#_c_137_n N_VPWR_c_534_n 0.00880551f $X=0.375 $Y=2.115 $X2=0
+ $Y2=0
cc_146 N_A_27_74#_c_133_n N_VPWR_c_540_n 0.00413917f $X=1.17 $Y=1.885 $X2=0
+ $Y2=0
cc_147 N_A_27_74#_c_133_n N_VPWR_c_529_n 0.00819732f $X=1.17 $Y=1.885 $X2=0
+ $Y2=0
cc_148 N_A_27_74#_c_137_n N_VPWR_c_529_n 0.0108814f $X=0.375 $Y=2.115 $X2=0
+ $Y2=0
cc_149 N_A_27_74#_M1002_g N_VGND_c_634_n 0.00391641f $X=1.485 $Y=0.78 $X2=0
+ $Y2=0
cc_150 N_A_27_74#_c_128_n N_VGND_c_634_n 0.0226023f $X=0.28 $Y=0.645 $X2=0 $Y2=0
cc_151 N_A_27_74#_c_129_n N_VGND_c_634_n 0.0182601f $X=0.765 $Y=1.195 $X2=0
+ $Y2=0
cc_152 N_A_27_74#_c_131_n N_VGND_c_634_n 0.010213f $X=0.85 $Y=1.67 $X2=0 $Y2=0
cc_153 N_A_27_74#_c_128_n N_VGND_c_636_n 0.011066f $X=0.28 $Y=0.645 $X2=0 $Y2=0
cc_154 N_A_27_74#_M1002_g N_VGND_c_637_n 0.00393863f $X=1.485 $Y=0.78 $X2=0
+ $Y2=0
cc_155 N_A_27_74#_M1002_g N_VGND_c_640_n 0.00533081f $X=1.485 $Y=0.78 $X2=0
+ $Y2=0
cc_156 N_A_27_74#_c_128_n N_VGND_c_640_n 0.00915947f $X=0.28 $Y=0.645 $X2=0
+ $Y2=0
cc_157 N_A_354_252#_c_195_n N_C_M1010_g 0.0030537f $X=1.935 $Y=1.425 $X2=0 $Y2=0
cc_158 N_A_354_252#_c_196_n N_C_M1010_g 0.00891742f $X=1.935 $Y=1.425 $X2=0
+ $Y2=0
cc_159 N_A_354_252#_c_197_n N_C_M1010_g 0.0164446f $X=3.475 $Y=1.085 $X2=0 $Y2=0
cc_160 N_A_354_252#_c_201_n N_C_M1010_g 0.0343132f $X=1.935 $Y=1.26 $X2=0 $Y2=0
cc_161 N_A_354_252#_c_194_n N_C_c_310_n 0.00940882f $X=1.89 $Y=1.795 $X2=0 $Y2=0
cc_162 N_A_354_252#_c_203_n N_C_c_310_n 0.0205338f $X=1.89 $Y=1.885 $X2=0 $Y2=0
cc_163 N_A_354_252#_c_195_n N_C_c_310_n 2.13462e-19 $X=1.935 $Y=1.425 $X2=0
+ $Y2=0
cc_164 N_A_354_252#_c_196_n N_C_c_310_n 0.0107049f $X=1.935 $Y=1.425 $X2=0 $Y2=0
cc_165 N_A_354_252#_c_197_n N_C_c_310_n 0.00433303f $X=3.475 $Y=1.085 $X2=0
+ $Y2=0
cc_166 N_A_354_252#_c_194_n C 0.00163055f $X=1.89 $Y=1.795 $X2=0 $Y2=0
cc_167 N_A_354_252#_c_195_n C 0.0110064f $X=1.935 $Y=1.425 $X2=0 $Y2=0
cc_168 N_A_354_252#_c_196_n C 5.88671e-19 $X=1.935 $Y=1.425 $X2=0 $Y2=0
cc_169 N_A_354_252#_c_197_n C 0.0251515f $X=3.475 $Y=1.085 $X2=0 $Y2=0
cc_170 N_A_354_252#_c_197_n N_D_M1013_g 0.0185539f $X=3.475 $Y=1.085 $X2=0 $Y2=0
cc_171 N_A_354_252#_c_228_p N_D_M1013_g 0.00271323f $X=3.56 $Y=1 $X2=0 $Y2=0
cc_172 N_A_354_252#_c_197_n N_D_c_344_n 0.00164497f $X=3.475 $Y=1.085 $X2=0
+ $Y2=0
cc_173 N_A_354_252#_c_197_n D 0.0183765f $X=3.475 $Y=1.085 $X2=0 $Y2=0
cc_174 N_A_354_252#_c_197_n N_A_225_82#_M1001_g 0.00161928f $X=3.475 $Y=1.085
+ $X2=0 $Y2=0
cc_175 N_A_354_252#_c_232_p N_A_225_82#_M1001_g 0.0135356f $X=4.365 $Y=0.665
+ $X2=0 $Y2=0
cc_176 N_A_354_252#_c_232_p N_A_225_82#_M1008_g 0.014255f $X=4.365 $Y=0.665
+ $X2=0 $Y2=0
cc_177 N_A_354_252#_c_198_n N_A_225_82#_M1008_g 0.00761203f $X=4.45 $Y=1.76
+ $X2=0 $Y2=0
cc_178 N_A_354_252#_c_206_n N_A_225_82#_c_386_n 0.00151518f $X=4.535 $Y=1.845
+ $X2=0 $Y2=0
cc_179 N_A_354_252#_c_207_n N_A_225_82#_c_386_n 5.96295e-19 $X=4.99 $Y=1.985
+ $X2=0 $Y2=0
cc_180 N_A_354_252#_c_201_n N_A_225_82#_c_380_n 0.00207976f $X=1.935 $Y=1.26
+ $X2=0 $Y2=0
cc_181 N_A_354_252#_c_194_n N_A_225_82#_c_381_n 0.00664175f $X=1.89 $Y=1.795
+ $X2=0 $Y2=0
cc_182 N_A_354_252#_c_203_n N_A_225_82#_c_381_n 0.00119554f $X=1.89 $Y=1.885
+ $X2=0 $Y2=0
cc_183 N_A_354_252#_c_195_n N_A_225_82#_c_381_n 0.0318557f $X=1.935 $Y=1.425
+ $X2=0 $Y2=0
cc_184 N_A_354_252#_c_196_n N_A_225_82#_c_381_n 0.00210056f $X=1.935 $Y=1.425
+ $X2=0 $Y2=0
cc_185 N_A_354_252#_c_203_n N_A_225_82#_c_388_n 0.0066357f $X=1.89 $Y=1.885
+ $X2=0 $Y2=0
cc_186 N_A_354_252#_c_203_n N_A_225_82#_c_389_n 0.0188406f $X=1.89 $Y=1.885
+ $X2=0 $Y2=0
cc_187 N_A_354_252#_c_195_n N_A_225_82#_c_389_n 0.0141669f $X=1.935 $Y=1.425
+ $X2=0 $Y2=0
cc_188 N_A_354_252#_c_196_n N_A_225_82#_c_389_n 8.86618e-19 $X=1.935 $Y=1.425
+ $X2=0 $Y2=0
cc_189 N_A_354_252#_c_203_n N_A_225_82#_c_390_n 8.61223e-19 $X=1.89 $Y=1.885
+ $X2=0 $Y2=0
cc_190 N_A_354_252#_c_247_p N_A_225_82#_c_382_n 0.00173038f $X=2.1 $Y=1.085
+ $X2=0 $Y2=0
cc_191 N_A_354_252#_c_201_n N_A_225_82#_c_382_n 4.31478e-19 $X=1.935 $Y=1.26
+ $X2=0 $Y2=0
cc_192 N_A_354_252#_c_203_n N_A_225_82#_c_393_n 3.05651e-19 $X=1.89 $Y=1.885
+ $X2=0 $Y2=0
cc_193 N_A_354_252#_c_197_n N_A_225_82#_c_383_n 0.0126261f $X=3.475 $Y=1.085
+ $X2=0 $Y2=0
cc_194 N_A_354_252#_c_232_p N_A_225_82#_c_383_n 0.0037988f $X=4.365 $Y=0.665
+ $X2=0 $Y2=0
cc_195 N_A_354_252#_c_197_n N_A_225_82#_c_384_n 0.00277924f $X=3.475 $Y=1.085
+ $X2=0 $Y2=0
cc_196 N_A_354_252#_c_198_n N_A_225_82#_c_384_n 0.00413158f $X=4.45 $Y=1.76
+ $X2=0 $Y2=0
cc_197 N_A_354_252#_c_198_n N_B_N_c_503_n 0.00703202f $X=4.45 $Y=1.76 $X2=-0.19
+ $Y2=-0.245
cc_198 N_A_354_252#_c_205_n N_B_N_c_503_n 0.0221723f $X=4.82 $Y=1.845 $X2=-0.19
+ $Y2=-0.245
cc_199 N_A_354_252#_c_207_n N_B_N_c_503_n 0.0133575f $X=4.99 $Y=1.985 $X2=-0.19
+ $Y2=-0.245
cc_200 N_A_354_252#_c_200_n N_B_N_c_503_n 0.0016773f $X=5 $Y=0.665 $X2=-0.19
+ $Y2=-0.245
cc_201 N_A_354_252#_c_198_n N_B_N_c_504_n 0.00664614f $X=4.45 $Y=1.76 $X2=0
+ $Y2=0
cc_202 N_A_354_252#_c_199_n N_B_N_c_504_n 0.0124991f $X=4.835 $Y=0.665 $X2=0
+ $Y2=0
cc_203 N_A_354_252#_c_200_n N_B_N_c_504_n 0.00587758f $X=5 $Y=0.665 $X2=0 $Y2=0
cc_204 N_A_354_252#_c_198_n B_N 0.0206499f $X=4.45 $Y=1.76 $X2=0 $Y2=0
cc_205 N_A_354_252#_c_199_n B_N 3.09683e-19 $X=4.835 $Y=0.665 $X2=0 $Y2=0
cc_206 N_A_354_252#_c_205_n B_N 0.0281059f $X=4.82 $Y=1.845 $X2=0 $Y2=0
cc_207 N_A_354_252#_c_200_n B_N 0.0246489f $X=5 $Y=0.665 $X2=0 $Y2=0
cc_208 N_A_354_252#_c_205_n N_VPWR_M1012_s 0.00136333f $X=4.82 $Y=1.845 $X2=0
+ $Y2=0
cc_209 N_A_354_252#_c_206_n N_VPWR_M1012_s 0.00321156f $X=4.535 $Y=1.845 $X2=0
+ $Y2=0
cc_210 N_A_354_252#_c_203_n N_VPWR_c_531_n 0.0109035f $X=1.89 $Y=1.885 $X2=0
+ $Y2=0
cc_211 N_A_354_252#_c_205_n N_VPWR_c_533_n 0.00639085f $X=4.82 $Y=1.845 $X2=0
+ $Y2=0
cc_212 N_A_354_252#_c_206_n N_VPWR_c_533_n 0.0152373f $X=4.535 $Y=1.845 $X2=0
+ $Y2=0
cc_213 N_A_354_252#_c_207_n N_VPWR_c_533_n 0.0396375f $X=4.99 $Y=1.985 $X2=0
+ $Y2=0
cc_214 N_A_354_252#_c_203_n N_VPWR_c_540_n 0.00461464f $X=1.89 $Y=1.885 $X2=0
+ $Y2=0
cc_215 N_A_354_252#_c_207_n N_VPWR_c_541_n 0.00698636f $X=4.99 $Y=1.985 $X2=0
+ $Y2=0
cc_216 N_A_354_252#_c_203_n N_VPWR_c_529_n 0.00913375f $X=1.89 $Y=1.885 $X2=0
+ $Y2=0
cc_217 N_A_354_252#_c_207_n N_VPWR_c_529_n 0.0104303f $X=4.99 $Y=1.985 $X2=0
+ $Y2=0
cc_218 N_A_354_252#_c_232_p N_X_M1001_d 0.00438182f $X=4.365 $Y=0.665 $X2=-0.19
+ $Y2=-0.245
cc_219 N_A_354_252#_c_197_n N_X_c_599_n 0.0073895f $X=3.475 $Y=1.085 $X2=0 $Y2=0
cc_220 N_A_354_252#_c_232_p N_X_c_599_n 0.0193287f $X=4.365 $Y=0.665 $X2=0 $Y2=0
cc_221 N_A_354_252#_c_198_n N_X_c_599_n 0.018632f $X=4.45 $Y=1.76 $X2=0 $Y2=0
cc_222 N_A_354_252#_c_207_n X 0.00434494f $X=4.99 $Y=1.985 $X2=0 $Y2=0
cc_223 N_A_354_252#_c_198_n N_X_c_600_n 0.0421223f $X=4.45 $Y=1.76 $X2=0 $Y2=0
cc_224 N_A_354_252#_c_206_n N_X_c_600_n 0.0138633f $X=4.535 $Y=1.845 $X2=0 $Y2=0
cc_225 N_A_354_252#_c_197_n N_VGND_M1013_d 0.0128486f $X=3.475 $Y=1.085 $X2=0
+ $Y2=0
cc_226 N_A_354_252#_c_228_p N_VGND_M1013_d 0.00423184f $X=3.56 $Y=1 $X2=0 $Y2=0
cc_227 N_A_354_252#_c_284_p N_VGND_M1013_d 0.0046727f $X=3.645 $Y=0.665 $X2=0
+ $Y2=0
cc_228 N_A_354_252#_c_232_p N_VGND_M1008_s 0.00178542f $X=4.365 $Y=0.665 $X2=0
+ $Y2=0
cc_229 N_A_354_252#_c_198_n N_VGND_M1008_s 0.0104856f $X=4.45 $Y=1.76 $X2=0
+ $Y2=0
cc_230 N_A_354_252#_c_199_n N_VGND_M1008_s 0.005464f $X=4.835 $Y=0.665 $X2=0
+ $Y2=0
cc_231 N_A_354_252#_c_288_p N_VGND_M1008_s 0.00253983f $X=4.45 $Y=0.665 $X2=0
+ $Y2=0
cc_232 N_A_354_252#_c_197_n N_VGND_c_635_n 0.0218816f $X=3.475 $Y=1.085 $X2=0
+ $Y2=0
cc_233 N_A_354_252#_c_228_p N_VGND_c_635_n 0.00607742f $X=3.56 $Y=1 $X2=0 $Y2=0
cc_234 N_A_354_252#_c_284_p N_VGND_c_635_n 0.0144778f $X=3.645 $Y=0.665 $X2=0
+ $Y2=0
cc_235 N_A_354_252#_c_201_n N_VGND_c_637_n 0.00548708f $X=1.935 $Y=1.26 $X2=0
+ $Y2=0
cc_236 N_A_354_252#_c_232_p N_VGND_c_638_n 0.0113015f $X=4.365 $Y=0.665 $X2=0
+ $Y2=0
cc_237 N_A_354_252#_c_284_p N_VGND_c_638_n 0.00354771f $X=3.645 $Y=0.665 $X2=0
+ $Y2=0
cc_238 N_A_354_252#_c_199_n N_VGND_c_639_n 0.00346124f $X=4.835 $Y=0.665 $X2=0
+ $Y2=0
cc_239 N_A_354_252#_c_200_n N_VGND_c_639_n 0.00717525f $X=5 $Y=0.665 $X2=0 $Y2=0
cc_240 N_A_354_252#_c_232_p N_VGND_c_640_n 0.0201945f $X=4.365 $Y=0.665 $X2=0
+ $Y2=0
cc_241 N_A_354_252#_c_284_p N_VGND_c_640_n 0.00533675f $X=3.645 $Y=0.665 $X2=0
+ $Y2=0
cc_242 N_A_354_252#_c_199_n N_VGND_c_640_n 0.00587114f $X=4.835 $Y=0.665 $X2=0
+ $Y2=0
cc_243 N_A_354_252#_c_288_p N_VGND_c_640_n 9.58892e-19 $X=4.45 $Y=0.665 $X2=0
+ $Y2=0
cc_244 N_A_354_252#_c_200_n N_VGND_c_640_n 0.0101296f $X=5 $Y=0.665 $X2=0 $Y2=0
cc_245 N_A_354_252#_c_201_n N_VGND_c_640_n 0.00533081f $X=1.935 $Y=1.26 $X2=0
+ $Y2=0
cc_246 N_A_354_252#_c_232_p N_VGND_c_643_n 0.00285472f $X=4.365 $Y=0.665 $X2=0
+ $Y2=0
cc_247 N_A_354_252#_c_199_n N_VGND_c_643_n 0.00892769f $X=4.835 $Y=0.665 $X2=0
+ $Y2=0
cc_248 N_A_354_252#_c_288_p N_VGND_c_643_n 0.0140478f $X=4.45 $Y=0.665 $X2=0
+ $Y2=0
cc_249 N_A_354_252#_c_197_n A_390_82# 0.00707549f $X=3.475 $Y=1.085 $X2=-0.19
+ $Y2=-0.245
cc_250 N_A_354_252#_c_247_p A_390_82# 0.0040802f $X=2.1 $Y=1.085 $X2=-0.19
+ $Y2=-0.245
cc_251 N_A_354_252#_c_197_n A_498_82# 0.00938627f $X=3.475 $Y=1.085 $X2=-0.19
+ $Y2=-0.245
cc_252 N_C_M1010_g N_D_M1013_g 0.0418504f $X=2.415 $Y=0.78 $X2=0 $Y2=0
cc_253 N_C_c_310_n N_D_c_344_n 0.0363929f $X=2.55 $Y=1.885 $X2=0 $Y2=0
cc_254 C N_D_c_344_n 0.00246628f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_255 N_C_c_310_n D 3.20914e-19 $X=2.55 $Y=1.885 $X2=0 $Y2=0
cc_256 C D 0.0291574f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_257 N_C_c_310_n N_A_225_82#_c_389_n 0.0142752f $X=2.55 $Y=1.885 $X2=0 $Y2=0
cc_258 C N_A_225_82#_c_389_n 0.022783f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_259 N_C_c_310_n N_A_225_82#_c_390_n 0.0113926f $X=2.55 $Y=1.885 $X2=0 $Y2=0
cc_260 N_C_c_310_n N_A_225_82#_c_394_n 9.78637e-19 $X=2.55 $Y=1.885 $X2=0 $Y2=0
cc_261 C N_A_225_82#_c_394_n 0.0127141f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_262 N_C_c_310_n N_VPWR_c_531_n 0.0103491f $X=2.55 $Y=1.885 $X2=0 $Y2=0
cc_263 N_C_c_310_n N_VPWR_c_536_n 0.00445602f $X=2.55 $Y=1.885 $X2=0 $Y2=0
cc_264 N_C_c_310_n N_VPWR_c_529_n 0.00859665f $X=2.55 $Y=1.885 $X2=0 $Y2=0
cc_265 N_C_M1010_g N_VGND_c_635_n 0.00258673f $X=2.415 $Y=0.78 $X2=0 $Y2=0
cc_266 N_C_M1010_g N_VGND_c_637_n 0.00548708f $X=2.415 $Y=0.78 $X2=0 $Y2=0
cc_267 N_C_M1010_g N_VGND_c_640_n 0.00533081f $X=2.415 $Y=0.78 $X2=0 $Y2=0
cc_268 N_D_M1013_g N_A_225_82#_M1001_g 0.0104375f $X=2.925 $Y=0.78 $X2=0 $Y2=0
cc_269 N_D_c_344_n N_A_225_82#_c_385_n 0.0163641f $X=3 $Y=1.885 $X2=0 $Y2=0
cc_270 N_D_c_344_n N_A_225_82#_c_390_n 0.0160543f $X=3 $Y=1.885 $X2=0 $Y2=0
cc_271 N_D_c_344_n N_A_225_82#_c_391_n 0.0145817f $X=3 $Y=1.885 $X2=0 $Y2=0
cc_272 D N_A_225_82#_c_391_n 0.024017f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_273 N_D_c_344_n N_A_225_82#_c_392_n 0.00373014f $X=3 $Y=1.885 $X2=0 $Y2=0
cc_274 D N_A_225_82#_c_392_n 0.00651523f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_275 N_D_c_344_n N_A_225_82#_c_394_n 0.0041631f $X=3 $Y=1.885 $X2=0 $Y2=0
cc_276 D N_A_225_82#_c_394_n 0.00113045f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_277 N_D_M1013_g N_A_225_82#_c_383_n 0.00141277f $X=2.925 $Y=0.78 $X2=0 $Y2=0
cc_278 N_D_c_344_n N_A_225_82#_c_383_n 0.00166013f $X=3 $Y=1.885 $X2=0 $Y2=0
cc_279 D N_A_225_82#_c_383_n 0.0154006f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_280 N_D_M1013_g N_A_225_82#_c_384_n 0.00141849f $X=2.925 $Y=0.78 $X2=0 $Y2=0
cc_281 N_D_c_344_n N_A_225_82#_c_384_n 0.0135551f $X=3 $Y=1.885 $X2=0 $Y2=0
cc_282 D N_A_225_82#_c_384_n 3.00649e-19 $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_283 N_D_c_344_n N_VPWR_c_532_n 0.010844f $X=3 $Y=1.885 $X2=0 $Y2=0
cc_284 N_D_c_344_n N_VPWR_c_536_n 0.00445602f $X=3 $Y=1.885 $X2=0 $Y2=0
cc_285 N_D_c_344_n N_VPWR_c_529_n 0.00860729f $X=3 $Y=1.885 $X2=0 $Y2=0
cc_286 N_D_M1013_g N_VGND_c_635_n 0.0147594f $X=2.925 $Y=0.78 $X2=0 $Y2=0
cc_287 N_D_M1013_g N_VGND_c_637_n 0.00455951f $X=2.925 $Y=0.78 $X2=0 $Y2=0
cc_288 N_D_M1013_g N_VGND_c_640_n 0.00447788f $X=2.925 $Y=0.78 $X2=0 $Y2=0
cc_289 N_A_225_82#_M1008_g N_B_N_c_503_n 0.00182278f $X=4.195 $Y=0.78 $X2=-0.19
+ $Y2=-0.245
cc_290 N_A_225_82#_c_386_n N_B_N_c_503_n 0.0179666f $X=4.225 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_291 N_A_225_82#_c_384_n N_B_N_c_503_n 0.0124013f $X=4.195 $Y=1.552 $X2=-0.19
+ $Y2=-0.245
cc_292 N_A_225_82#_M1008_g N_B_N_c_504_n 0.0170269f $X=4.195 $Y=0.78 $X2=0 $Y2=0
cc_293 N_A_225_82#_c_389_n N_VPWR_M1009_d 0.00740139f $X=2.61 $Y=2.035 $X2=0
+ $Y2=0
cc_294 N_A_225_82#_c_391_n N_VPWR_M1011_d 0.0167791f $X=3.495 $Y=2.035 $X2=0
+ $Y2=0
cc_295 N_A_225_82#_c_392_n N_VPWR_M1011_d 0.0023678f $X=3.58 $Y=1.95 $X2=0 $Y2=0
cc_296 N_A_225_82#_c_388_n N_VPWR_c_530_n 0.0330122f $X=1.595 $Y=2.815 $X2=0
+ $Y2=0
cc_297 N_A_225_82#_c_388_n N_VPWR_c_531_n 0.0185533f $X=1.595 $Y=2.815 $X2=0
+ $Y2=0
cc_298 N_A_225_82#_c_389_n N_VPWR_c_531_n 0.0266856f $X=2.61 $Y=2.035 $X2=0
+ $Y2=0
cc_299 N_A_225_82#_c_390_n N_VPWR_c_531_n 0.0447456f $X=2.775 $Y=2.815 $X2=0
+ $Y2=0
cc_300 N_A_225_82#_c_385_n N_VPWR_c_532_n 0.0104271f $X=3.775 $Y=1.765 $X2=0
+ $Y2=0
cc_301 N_A_225_82#_c_390_n N_VPWR_c_532_n 0.0387012f $X=2.775 $Y=2.815 $X2=0
+ $Y2=0
cc_302 N_A_225_82#_c_391_n N_VPWR_c_532_n 0.026815f $X=3.495 $Y=2.035 $X2=0
+ $Y2=0
cc_303 N_A_225_82#_c_386_n N_VPWR_c_533_n 0.00825088f $X=4.225 $Y=1.765 $X2=0
+ $Y2=0
cc_304 N_A_225_82#_c_390_n N_VPWR_c_536_n 0.014552f $X=2.775 $Y=2.815 $X2=0
+ $Y2=0
cc_305 N_A_225_82#_c_385_n N_VPWR_c_538_n 0.00445602f $X=3.775 $Y=1.765 $X2=0
+ $Y2=0
cc_306 N_A_225_82#_c_386_n N_VPWR_c_538_n 0.00411612f $X=4.225 $Y=1.765 $X2=0
+ $Y2=0
cc_307 N_A_225_82#_c_388_n N_VPWR_c_540_n 0.0146357f $X=1.595 $Y=2.815 $X2=0
+ $Y2=0
cc_308 N_A_225_82#_c_385_n N_VPWR_c_529_n 0.00860645f $X=3.775 $Y=1.765 $X2=0
+ $Y2=0
cc_309 N_A_225_82#_c_386_n N_VPWR_c_529_n 0.00752331f $X=4.225 $Y=1.765 $X2=0
+ $Y2=0
cc_310 N_A_225_82#_c_388_n N_VPWR_c_529_n 0.0121141f $X=1.595 $Y=2.815 $X2=0
+ $Y2=0
cc_311 N_A_225_82#_c_390_n N_VPWR_c_529_n 0.0119791f $X=2.775 $Y=2.815 $X2=0
+ $Y2=0
cc_312 N_A_225_82#_M1001_g N_X_c_599_n 0.00349132f $X=3.765 $Y=0.78 $X2=0 $Y2=0
cc_313 N_A_225_82#_M1008_g N_X_c_599_n 0.00488473f $X=4.195 $Y=0.78 $X2=0 $Y2=0
cc_314 N_A_225_82#_c_383_n N_X_c_599_n 0.0029987f $X=3.69 $Y=1.505 $X2=0 $Y2=0
cc_315 N_A_225_82#_c_384_n N_X_c_599_n 0.00269894f $X=4.195 $Y=1.552 $X2=0 $Y2=0
cc_316 N_A_225_82#_c_385_n X 0.00198005f $X=3.775 $Y=1.765 $X2=0 $Y2=0
cc_317 N_A_225_82#_c_386_n X 0.00291296f $X=4.225 $Y=1.765 $X2=0 $Y2=0
cc_318 N_A_225_82#_c_383_n X 0.00126392f $X=3.69 $Y=1.505 $X2=0 $Y2=0
cc_319 N_A_225_82#_c_384_n X 0.00466761f $X=4.195 $Y=1.552 $X2=0 $Y2=0
cc_320 N_A_225_82#_c_385_n X 0.0183391f $X=3.775 $Y=1.765 $X2=0 $Y2=0
cc_321 N_A_225_82#_c_386_n X 0.0130018f $X=4.225 $Y=1.765 $X2=0 $Y2=0
cc_322 N_A_225_82#_M1001_g N_X_c_600_n 0.00344857f $X=3.765 $Y=0.78 $X2=0 $Y2=0
cc_323 N_A_225_82#_c_385_n N_X_c_600_n 5.7161e-19 $X=3.775 $Y=1.765 $X2=0 $Y2=0
cc_324 N_A_225_82#_M1008_g N_X_c_600_n 0.00356046f $X=4.195 $Y=0.78 $X2=0 $Y2=0
cc_325 N_A_225_82#_c_386_n N_X_c_600_n 0.00138061f $X=4.225 $Y=1.765 $X2=0 $Y2=0
cc_326 N_A_225_82#_c_392_n N_X_c_600_n 0.00754692f $X=3.58 $Y=1.95 $X2=0 $Y2=0
cc_327 N_A_225_82#_c_383_n N_X_c_600_n 0.023711f $X=3.69 $Y=1.505 $X2=0 $Y2=0
cc_328 N_A_225_82#_c_384_n N_X_c_600_n 0.0178955f $X=4.195 $Y=1.552 $X2=0 $Y2=0
cc_329 N_A_225_82#_c_380_n N_VGND_c_634_n 0.0382158f $X=1.27 $Y=0.555 $X2=0
+ $Y2=0
cc_330 N_A_225_82#_M1001_g N_VGND_c_635_n 0.00689129f $X=3.765 $Y=0.78 $X2=0
+ $Y2=0
cc_331 N_A_225_82#_c_380_n N_VGND_c_637_n 0.018524f $X=1.27 $Y=0.555 $X2=0 $Y2=0
cc_332 N_A_225_82#_M1001_g N_VGND_c_638_n 0.00414982f $X=3.765 $Y=0.78 $X2=0
+ $Y2=0
cc_333 N_A_225_82#_M1008_g N_VGND_c_638_n 0.00414982f $X=4.195 $Y=0.78 $X2=0
+ $Y2=0
cc_334 N_A_225_82#_M1001_g N_VGND_c_640_n 0.00533081f $X=3.765 $Y=0.78 $X2=0
+ $Y2=0
cc_335 N_A_225_82#_M1008_g N_VGND_c_640_n 0.00533081f $X=4.195 $Y=0.78 $X2=0
+ $Y2=0
cc_336 N_A_225_82#_c_380_n N_VGND_c_640_n 0.0176287f $X=1.27 $Y=0.555 $X2=0
+ $Y2=0
cc_337 N_A_225_82#_M1008_g N_VGND_c_643_n 0.00546687f $X=4.195 $Y=0.78 $X2=0
+ $Y2=0
cc_338 N_B_N_c_503_n N_VPWR_c_533_n 0.00823143f $X=4.76 $Y=1.765 $X2=0 $Y2=0
cc_339 N_B_N_c_503_n N_VPWR_c_541_n 0.00393873f $X=4.76 $Y=1.765 $X2=0 $Y2=0
cc_340 N_B_N_c_503_n N_VPWR_c_529_n 0.00462577f $X=4.76 $Y=1.765 $X2=0 $Y2=0
cc_341 N_B_N_c_503_n X 7.09034e-19 $X=4.76 $Y=1.765 $X2=0 $Y2=0
cc_342 N_B_N_c_503_n N_X_c_600_n 2.38613e-19 $X=4.76 $Y=1.765 $X2=0 $Y2=0
cc_343 N_B_N_c_504_n N_VGND_c_639_n 0.0032796f $X=4.785 $Y=1.26 $X2=0 $Y2=0
cc_344 N_B_N_c_504_n N_VGND_c_640_n 0.00476395f $X=4.785 $Y=1.26 $X2=0 $Y2=0
cc_345 N_VPWR_c_532_n X 0.0344701f $X=3.365 $Y=2.405 $X2=0 $Y2=0
cc_346 N_VPWR_c_533_n X 0.0673472f $X=4.45 $Y=2.265 $X2=0 $Y2=0
cc_347 N_VPWR_c_538_n X 0.0158009f $X=4.365 $Y=3.33 $X2=0 $Y2=0
cc_348 N_VPWR_c_529_n X 0.0129424f $X=5.04 $Y=3.33 $X2=0 $Y2=0
