* NGSPICE file created from sky130_fd_sc_ls__a2111oi_1.ext - technology: sky130A

.subckt sky130_fd_sc_ls__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
M1000 a_234_368# C1 a_156_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=4.368e+11p pd=3.02e+06u as=2.688e+11p ps=2.72e+06u
M1001 VGND A2 a_461_74# VNB nshort w=740000u l=150000u
+  ad=7.77e+11p pd=6.54e+06u as=2.368e+11p ps=2.12e+06u
M1002 a_461_74# A1 Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=4.144e+11p ps=4.08e+06u
M1003 Y D1 VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_342_368# A2 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=7.448e+11p pd=5.81e+06u as=4.368e+11p ps=3.02e+06u
M1005 a_342_368# B1 a_234_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND C1 Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_156_368# D1 Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.08e+11p ps=2.79e+06u
M1008 Y B1 VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR A1 a_342_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

