* File: sky130_fd_sc_ls__dfstp_1.pex.spice
* Created: Wed Sep  2 11:01:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__DFSTP_1%D 2 4 7 9 11 12 13 17 18 21
c35 18 0 7.5678e-20 $X=0.64 $Y=1.145
r36 21 23 39.9775 $w=4e-07 $l=1.65e-07 $layer=POLY_cond $X=0.605 $Y=1.825
+ $X2=0.605 $Y2=1.99
r37 21 22 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.64
+ $Y=1.825 $X2=0.64 $Y2=1.825
r38 17 19 45.6753 $w=4e-07 $l=1.65e-07 $layer=POLY_cond $X=0.605 $Y=1.145
+ $X2=0.605 $Y2=0.98
r39 17 18 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.64
+ $Y=1.145 $X2=0.64 $Y2=1.145
r40 13 22 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=0.64 $Y=1.665
+ $X2=0.64 $Y2=1.825
r41 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.64 $Y=1.295
+ $X2=0.64 $Y2=1.665
r42 12 18 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=0.64 $Y=1.295
+ $X2=0.64 $Y2=1.145
r43 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.495 $Y=2.465
+ $X2=0.495 $Y2=2.75
r44 7 19 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=0.495 $Y=0.58 $X2=0.495
+ $Y2=0.98
r45 4 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.495 $Y=2.375 $X2=0.495
+ $Y2=2.465
r46 4 23 149.653 $w=1.8e-07 $l=3.85e-07 $layer=POLY_cond $X=0.495 $Y=2.375
+ $X2=0.495 $Y2=1.99
r47 2 21 4.86635 $w=4e-07 $l=3.5e-08 $layer=POLY_cond $X=0.605 $Y=1.79 $X2=0.605
+ $Y2=1.825
r48 1 17 4.86635 $w=4e-07 $l=3.5e-08 $layer=POLY_cond $X=0.605 $Y=1.18 $X2=0.605
+ $Y2=1.145
r49 1 2 84.8135 $w=4e-07 $l=6.1e-07 $layer=POLY_cond $X=0.605 $Y=1.18 $X2=0.605
+ $Y2=1.79
.ends

.subckt PM_SKY130_FD_SC_LS__DFSTP_1%CLK 1 3 4 6 7
c33 1 0 1.72487e-19 $X=1.48 $Y=1.675
r34 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.465
+ $Y=1.385 $X2=1.465 $Y2=1.385
r35 7 11 6.69663 $w=3.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.68 $Y=1.365
+ $X2=1.465 $Y2=1.365
r36 4 10 38.6342 $w=2.88e-07 $l=1.74714e-07 $layer=POLY_cond $X=1.485 $Y=1.22
+ $X2=1.465 $Y2=1.385
r37 4 6 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.485 $Y=1.22 $X2=1.485
+ $Y2=0.74
r38 1 10 59.5544 $w=2.88e-07 $l=2.97405e-07 $layer=POLY_cond $X=1.48 $Y=1.675
+ $X2=1.465 $Y2=1.385
r39 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.48 $Y=1.675
+ $X2=1.48 $Y2=2.31
.ends

.subckt PM_SKY130_FD_SC_LS__DFSTP_1%A_398_74# 1 2 7 9 10 11 14 18 19 21 23 26 30
+ 32 33 34 35 36 38 39 45 49 50 53 54 55 57 58 59 61 62 63 67 68 69 71 72 73 75
+ 76 77 80 84 89
c282 76 0 2.26502e-20 $X=6.48 $Y=1.285
c283 75 0 8.25365e-20 $X=6.48 $Y=1.285
c284 67 0 1.10875e-19 $X=6.32 $Y=1.715
c285 59 0 5.18726e-20 $X=5.365 $Y=2.405
c286 50 0 1.73639e-19 $X=4.4 $Y=2.17
c287 14 0 8.43983e-20 $X=3.625 $Y=0.58
r288 84 85 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=3.67 $Y=1.51
+ $X2=3.67 $Y2=1.435
r289 80 82 5.14244 $w=3.44e-07 $l=1.45e-07 $layer=LI1_cond $X=7.095 $Y=2.162
+ $X2=7.24 $Y2=2.162
r290 80 81 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.095
+ $Y=2.185 $X2=7.095 $Y2=2.185
r291 76 89 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.48 $Y=1.285
+ $X2=6.48 $Y2=1.12
r292 75 78 8.69073 $w=4.08e-07 $l=1.65e-07 $layer=LI1_cond $X=6.44 $Y=1.285
+ $X2=6.44 $Y2=1.45
r293 75 77 8.69073 $w=4.08e-07 $l=1.65e-07 $layer=LI1_cond $X=6.44 $Y=1.285
+ $X2=6.44 $Y2=1.12
r294 75 76 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.48
+ $Y=1.285 $X2=6.48 $Y2=1.285
r295 71 82 4.87082 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=7.24 $Y=1.97
+ $X2=7.24 $Y2=2.162
r296 70 71 100.797 $w=1.68e-07 $l=1.545e-06 $layer=LI1_cond $X=7.24 $Y=0.425
+ $X2=7.24 $Y2=1.97
r297 68 70 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.155 $Y=0.34
+ $X2=7.24 $Y2=0.425
r298 68 69 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=7.155 $Y=0.34
+ $X2=6.405 $Y2=0.34
r299 67 78 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=6.32 $Y=1.715
+ $X2=6.32 $Y2=1.45
r300 64 69 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.32 $Y=0.425
+ $X2=6.405 $Y2=0.34
r301 64 77 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=6.32 $Y=0.425
+ $X2=6.32 $Y2=1.12
r302 62 67 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.235 $Y=1.8
+ $X2=6.32 $Y2=1.715
r303 62 63 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=6.235 $Y=1.8
+ $X2=5.975 $Y2=1.8
r304 60 63 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.89 $Y=1.885
+ $X2=5.975 $Y2=1.8
r305 60 61 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=5.89 $Y=1.885
+ $X2=5.89 $Y2=2.32
r306 58 61 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.805 $Y=2.405
+ $X2=5.89 $Y2=2.32
r307 58 59 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=5.805 $Y=2.405
+ $X2=5.365 $Y2=2.405
r308 56 59 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.28 $Y=2.49
+ $X2=5.365 $Y2=2.405
r309 56 57 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=5.28 $Y=2.49
+ $X2=5.28 $Y2=2.905
r310 54 57 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.195 $Y=2.99
+ $X2=5.28 $Y2=2.905
r311 54 55 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=5.195 $Y=2.99
+ $X2=4.57 $Y2=2.99
r312 53 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.485 $Y=2.905
+ $X2=4.57 $Y2=2.99
r313 52 53 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=4.485 $Y=2.255
+ $X2=4.485 $Y2=2.905
r314 51 73 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.755 $Y=2.17
+ $X2=3.67 $Y2=2.17
r315 50 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.4 $Y=2.17
+ $X2=4.485 $Y2=2.255
r316 50 51 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=4.4 $Y=2.17
+ $X2=3.755 $Y2=2.17
r317 48 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.67 $Y=2.255
+ $X2=3.67 $Y2=2.17
r318 48 49 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=3.67 $Y=2.255
+ $X2=3.67 $Y2=2.905
r319 46 84 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.67 $Y=1.6 $X2=3.67
+ $Y2=1.51
r320 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.67
+ $Y=1.6 $X2=3.67 $Y2=1.6
r321 43 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.67 $Y=2.085
+ $X2=3.67 $Y2=2.17
r322 43 45 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=3.67 $Y=2.085
+ $X2=3.67 $Y2=1.6
r323 41 72 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=2.99 $Y=0.425
+ $X2=2.99 $Y2=1.435
r324 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.95
+ $Y=1.6 $X2=2.95 $Y2=1.6
r325 36 72 6.82988 $w=2.43e-07 $l=1.22e-07 $layer=LI1_cond $X=2.952 $Y=1.557
+ $X2=2.952 $Y2=1.435
r326 36 38 2.02266 $w=2.43e-07 $l=4.3e-08 $layer=LI1_cond $X=2.952 $Y=1.557
+ $X2=2.952 $Y2=1.6
r327 34 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.585 $Y=2.99
+ $X2=3.67 $Y2=2.905
r328 34 35 82.5294 $w=1.68e-07 $l=1.265e-06 $layer=LI1_cond $X=3.585 $Y=2.99
+ $X2=2.32 $Y2=2.99
r329 32 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.905 $Y=0.34
+ $X2=2.99 $Y2=0.425
r330 32 33 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=2.905 $Y=0.34
+ $X2=2.295 $Y2=0.34
r331 28 35 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.195 $Y=2.905
+ $X2=2.32 $Y2=2.99
r332 28 30 11.9854 $w=2.48e-07 $l=2.6e-07 $layer=LI1_cond $X=2.195 $Y=2.905
+ $X2=2.195 $Y2=2.645
r333 24 33 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.13 $Y=0.425
+ $X2=2.295 $Y2=0.34
r334 24 26 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=2.13 $Y=0.425
+ $X2=2.13 $Y2=0.515
r335 23 39 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.95 $Y=1.94
+ $X2=2.95 $Y2=1.6
r336 22 39 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=2.95 $Y=1.585
+ $X2=2.95 $Y2=1.6
r337 19 81 55.8714 $w=3.2e-07 $l=3.24037e-07 $layer=POLY_cond $X=7.21 $Y=2.465
+ $X2=7.115 $Y2=2.185
r338 19 21 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.21 $Y=2.465
+ $X2=7.21 $Y2=2.75
r339 18 89 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=6.525 $Y=0.69
+ $X2=6.525 $Y2=1.12
r340 14 85 438.415 $w=1.5e-07 $l=8.55e-07 $layer=POLY_cond $X=3.625 $Y=0.58
+ $X2=3.625 $Y2=1.435
r341 11 22 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=3.115 $Y=1.51
+ $X2=2.95 $Y2=1.585
r342 10 84 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.505 $Y=1.51
+ $X2=3.67 $Y2=1.51
r343 10 11 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=3.505 $Y=1.51
+ $X2=3.115 $Y2=1.51
r344 7 23 55.1908 $w=2.62e-07 $l=3.09839e-07 $layer=POLY_cond $X=2.97 $Y=2.24
+ $X2=2.95 $Y2=1.94
r345 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.97 $Y=2.24 $X2=2.97
+ $Y2=2.525
r346 2 30 600 $w=1.7e-07 $l=9.67096e-07 $layer=licon1_PDIFF $count=1 $X=2.005
+ $Y=1.75 $X2=2.155 $Y2=2.645
r347 1 26 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.99
+ $Y=0.37 $X2=2.13 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__DFSTP_1%A_760_395# 1 2 7 9 10 12 14 15 23 25 30 31
+ 35
c82 35 0 9.9779e-20 $X=4.31 $Y=1.065
c83 25 0 8.43983e-20 $X=4.43 $Y=1.065
r84 30 31 10.151 $w=2.83e-07 $l=2.05e-07 $layer=LI1_cond $X=4.882 $Y=2.525
+ $X2=4.882 $Y2=2.32
r85 26 35 23.3226 $w=2.48e-07 $l=1.2e-07 $layer=POLY_cond $X=4.43 $Y=1.065
+ $X2=4.31 $Y2=1.065
r86 25 28 13.0154 $w=3.89e-07 $l=4.15e-07 $layer=LI1_cond $X=4.43 $Y=0.872
+ $X2=4.845 $Y2=0.872
r87 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.43
+ $Y=1.065 $X2=4.43 $Y2=1.065
r88 20 23 9.07524 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.22 $Y=1.8
+ $X2=4.385 $Y2=1.8
r89 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.22
+ $Y=1.8 $X2=4.22 $Y2=1.8
r90 17 31 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=4.825 $Y=1.915
+ $X2=4.825 $Y2=2.32
r91 15 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.74 $Y=1.83
+ $X2=4.825 $Y2=1.915
r92 15 23 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=4.74 $Y=1.83
+ $X2=4.385 $Y2=1.83
r93 14 21 45.364 $w=3.18e-07 $l=3.05457e-07 $layer=POLY_cond $X=4.31 $Y=1.59
+ $X2=4.092 $Y2=1.8
r94 13 35 14.534 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.31 $Y=1.23
+ $X2=4.31 $Y2=1.065
r95 13 14 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=4.31 $Y=1.23
+ $X2=4.31 $Y2=1.59
r96 10 35 57.3347 $w=2.48e-07 $l=3.68375e-07 $layer=POLY_cond $X=4.015 $Y=0.9
+ $X2=4.31 $Y2=1.065
r97 10 12 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.015 $Y=0.9
+ $X2=4.015 $Y2=0.58
r98 7 21 80.2256 $w=3.18e-07 $l=5.31488e-07 $layer=POLY_cond $X=3.89 $Y=2.24
+ $X2=4.092 $Y2=1.8
r99 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.89 $Y=2.24 $X2=3.89
+ $Y2=2.525
r100 2 30 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=4.79
+ $Y=2.315 $X2=4.94 $Y2=2.525
r101 1 28 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.705
+ $Y=0.59 $X2=4.845 $Y2=0.8
.ends

.subckt PM_SKY130_FD_SC_LS__DFSTP_1%A_604_74# 1 2 8 9 11 14 16 18 21 25 29 32 34
+ 37 38 40 44 45 47 48
c143 37 0 9.9779e-20 $X=4.97 $Y=1.38
c144 16 0 6.04515e-20 $X=5.91 $Y=1.63
c145 9 0 2.25511e-19 $X=4.715 $Y=2.24
r146 44 45 10.3582 $w=3.33e-07 $l=2.2e-07 $layer=LI1_cond $X=3.247 $Y=2.515
+ $X2=3.247 $Y2=2.295
r147 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.9
+ $Y=1.38 $X2=5.9 $Y2=1.38
r148 38 51 13.6415 $w=3.18e-07 $l=9e-08 $layer=POLY_cond $X=4.97 $Y=1.447
+ $X2=5.06 $Y2=1.447
r149 38 49 38.6509 $w=3.18e-07 $l=2.55e-07 $layer=POLY_cond $X=4.97 $Y=1.447
+ $X2=4.715 $Y2=1.447
r150 37 48 7.72582 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.97 $Y=1.38
+ $X2=4.805 $Y2=1.38
r151 37 40 32.4779 $w=3.28e-07 $l=9.3e-07 $layer=LI1_cond $X=4.97 $Y=1.38
+ $X2=5.9 $Y2=1.38
r152 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.97
+ $Y=1.38 $X2=4.97 $Y2=1.38
r153 34 48 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=4.095 $Y=1.43
+ $X2=4.805 $Y2=1.43
r154 32 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.01 $Y=1.345
+ $X2=4.095 $Y2=1.43
r155 31 32 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=4.01 $Y=1.02
+ $X2=4.01 $Y2=1.345
r156 30 47 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.575 $Y=0.935
+ $X2=3.41 $Y2=0.935
r157 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.925 $Y=0.935
+ $X2=4.01 $Y2=1.02
r158 29 30 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=3.925 $Y=0.935
+ $X2=3.575 $Y2=0.935
r159 27 47 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=3.33 $Y=1.02
+ $X2=3.41 $Y2=0.935
r160 27 45 83.1818 $w=1.68e-07 $l=1.275e-06 $layer=LI1_cond $X=3.33 $Y=1.02
+ $X2=3.33 $Y2=2.295
r161 23 47 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.41 $Y=0.85
+ $X2=3.41 $Y2=0.935
r162 23 25 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=3.41 $Y=0.85
+ $X2=3.41 $Y2=0.58
r163 19 41 38.5336 $w=3.07e-07 $l=2.07123e-07 $layer=POLY_cond $X=6 $Y=1.215
+ $X2=5.905 $Y2=1.38
r164 19 21 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=6 $Y=1.215 $X2=6
+ $Y2=0.69
r165 16 41 51.8789 $w=3.07e-07 $l=2.52488e-07 $layer=POLY_cond $X=5.91 $Y=1.63
+ $X2=5.905 $Y2=1.38
r166 16 18 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.91 $Y=1.63
+ $X2=5.91 $Y2=2.205
r167 12 51 20.3436 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=5.06 $Y=1.215
+ $X2=5.06 $Y2=1.447
r168 12 14 212.798 $w=1.5e-07 $l=4.15e-07 $layer=POLY_cond $X=5.06 $Y=1.215
+ $X2=5.06 $Y2=0.8
r169 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.715 $Y=2.24
+ $X2=4.715 $Y2=2.525
r170 8 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=4.715 $Y=2.15 $X2=4.715
+ $Y2=2.24
r171 7 49 16.0701 $w=1.8e-07 $l=2.33e-07 $layer=POLY_cond $X=4.715 $Y=1.68
+ $X2=4.715 $Y2=1.447
r172 7 8 182.694 $w=1.8e-07 $l=4.7e-07 $layer=POLY_cond $X=4.715 $Y=1.68
+ $X2=4.715 $Y2=2.15
r173 2 44 600 $w=1.7e-07 $l=2.82843e-07 $layer=licon1_PDIFF $count=1 $X=3.045
+ $Y=2.315 $X2=3.245 $Y2=2.515
r174 1 25 182 $w=1.7e-07 $l=4.83735e-07 $layer=licon1_NDIFF $count=1 $X=3.02
+ $Y=0.37 $X2=3.41 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_LS__DFSTP_1%SET_B 1 3 6 8 10 11 12 13 15 16 17 18 19 22
+ 24 32
c129 32 0 7.26887e-20 $X=8.35 $Y=1.295
r130 34 35 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=8.35
+ $Y=1.975 $X2=8.35 $Y2=1.975
r131 32 35 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=8.35 $Y=1.295
+ $X2=8.35 $Y2=1.975
r132 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.245
+ $Y=1.985 $X2=5.245 $Y2=1.985
r133 24 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=2.035
+ $X2=8.4 $Y2=2.035
r134 22 28 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=5.52 $Y=1.985
+ $X2=5.245 $Y2=1.985
r135 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=2.035
+ $X2=5.52 $Y2=2.035
r136 19 21 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.665 $Y=2.035
+ $X2=5.52 $Y2=2.035
r137 18 24 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.255 $Y=2.035
+ $X2=8.4 $Y2=2.035
r138 18 19 3.20544 $w=1.4e-07 $l=2.59e-06 $layer=MET1_cond $X=8.255 $Y=2.035
+ $X2=5.665 $Y2=2.035
r139 17 34 9.54844 $w=4.95e-07 $l=8.91852e-08 $layer=POLY_cond $X=8.267 $Y=1.893
+ $X2=8.252 $Y2=1.975
r140 16 32 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=8.35
+ $Y=1.295 $X2=8.35 $Y2=1.295
r141 16 17 55.7728 $w=4.95e-07 $l=5.16e-07 $layer=POLY_cond $X=8.267 $Y=1.377
+ $X2=8.267 $Y2=1.893
r142 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=8.08 $Y=2.465
+ $X2=8.08 $Y2=2.75
r143 12 13 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=8.08 $Y=2.375
+ $X2=8.08 $Y2=2.465
r144 11 34 45.3963 $w=4.1e-07 $l=3.29977e-07 $layer=POLY_cond $X=8.08 $Y=2.23
+ $X2=8.252 $Y2=1.975
r145 11 12 56.3629 $w=1.8e-07 $l=1.45e-07 $layer=POLY_cond $X=8.08 $Y=2.23
+ $X2=8.08 $Y2=2.375
r146 8 16 82.838 $w=2.63e-07 $l=7.02544e-07 $layer=POLY_cond $X=7.815 $Y=0.865
+ $X2=8.267 $Y2=1.377
r147 8 10 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.815 $Y=0.865
+ $X2=7.815 $Y2=0.58
r148 4 27 39.0253 $w=3.68e-07 $l=2.22486e-07 $layer=POLY_cond $X=5.42 $Y=1.82
+ $X2=5.285 $Y2=1.985
r149 4 6 523.021 $w=1.5e-07 $l=1.02e-06 $layer=POLY_cond $X=5.42 $Y=1.82
+ $X2=5.42 $Y2=0.8
r150 1 27 50.8133 $w=3.68e-07 $l=3.09233e-07 $layer=POLY_cond $X=5.165 $Y=2.24
+ $X2=5.285 $Y2=1.985
r151 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=5.165 $Y=2.24
+ $X2=5.165 $Y2=2.525
.ends

.subckt PM_SKY130_FD_SC_LS__DFSTP_1%A_224_350# 1 2 9 11 13 15 16 18 19 22 24 25
+ 26 28 29 34 35 36 39 42 43 44 45 47 48 52 56 63
c192 42 0 6.14252e-20 $X=1.93 $Y=1.467
c193 35 0 8.25365e-20 $X=6.96 $Y=1.735
c194 26 0 1.22961e-19 $X=3.47 $Y=2.81
r195 62 63 8.47192 $w=3.38e-07 $l=1.65e-07 $layer=LI1_cond $X=1.255 $Y=1.89
+ $X2=1.42 $Y2=1.89
r196 59 62 6.6096 $w=3.38e-07 $l=1.95e-07 $layer=LI1_cond $X=1.06 $Y=1.89
+ $X2=1.255 $Y2=1.89
r197 56 58 17.8607 $w=4.58e-07 $l=4.95e-07 $layer=LI1_cond $X=1.205 $Y=0.515
+ $X2=1.205 $Y2=1.01
r198 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.15
+ $Y=1.425 $X2=2.15 $Y2=1.425
r199 50 52 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.15 $Y=1.72
+ $X2=2.15 $Y2=1.425
r200 48 50 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.985 $Y=1.805
+ $X2=2.15 $Y2=1.72
r201 48 63 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=1.985 $Y=1.805
+ $X2=1.42 $Y2=1.805
r202 47 59 4.80115 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=1.06 $Y=1.72
+ $X2=1.06 $Y2=1.89
r203 47 58 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=1.06 $Y=1.72
+ $X2=1.06 $Y2=1.01
r204 43 53 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=2.375 $Y=1.425
+ $X2=2.15 $Y2=1.425
r205 43 44 13.5877 $w=2.4e-07 $l=1.40584e-07 $layer=POLY_cond $X=2.375 $Y=1.425
+ $X2=2.45 $Y2=1.317
r206 41 53 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=2.02 $Y=1.425
+ $X2=2.15 $Y2=1.425
r207 41 42 5.03009 $w=3.3e-07 $l=1.08995e-07 $layer=POLY_cond $X=2.02 $Y=1.425
+ $X2=1.93 $Y2=1.467
r208 37 39 553.787 $w=1.5e-07 $l=1.08e-06 $layer=POLY_cond $X=7.035 $Y=1.66
+ $X2=7.035 $Y2=0.58
r209 35 37 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.96 $Y=1.735
+ $X2=7.035 $Y2=1.66
r210 35 36 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=6.96 $Y=1.735
+ $X2=6.505 $Y2=1.735
r211 32 34 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.415 $Y=3.035
+ $X2=6.415 $Y2=2.46
r212 31 36 26.9307 $w=1.5e-07 $l=1.89737e-07 $layer=POLY_cond $X=6.415 $Y=1.885
+ $X2=6.505 $Y2=1.735
r213 31 34 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.415 $Y=1.885
+ $X2=6.415 $Y2=2.46
r214 30 45 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.56 $Y=3.15 $X2=3.47
+ $Y2=3.15
r215 29 32 26.9307 $w=1.5e-07 $l=1.53542e-07 $layer=POLY_cond $X=6.325 $Y=3.15
+ $X2=6.415 $Y2=3.035
r216 29 30 1417.8 $w=1.5e-07 $l=2.765e-06 $layer=POLY_cond $X=6.325 $Y=3.15
+ $X2=3.56 $Y2=3.15
r217 26 28 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.47 $Y=2.81
+ $X2=3.47 $Y2=2.525
r218 25 45 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=3.47 $Y=3.075
+ $X2=3.47 $Y2=3.15
r219 24 26 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.47 $Y=2.9 $X2=3.47
+ $Y2=2.81
r220 24 25 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=3.47 $Y=2.9
+ $X2=3.47 $Y2=3.075
r221 20 22 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.945 $Y=1.045
+ $X2=2.945 $Y2=0.58
r222 18 45 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.38 $Y=3.15 $X2=3.47
+ $Y2=3.15
r223 18 19 438.415 $w=1.5e-07 $l=8.55e-07 $layer=POLY_cond $X=3.38 $Y=3.15
+ $X2=2.525 $Y2=3.15
r224 17 44 13.5877 $w=2.4e-07 $l=2.31482e-07 $layer=POLY_cond $X=2.525 $Y=1.12
+ $X2=2.45 $Y2=1.317
r225 16 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.87 $Y=1.12
+ $X2=2.945 $Y2=1.045
r226 16 17 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=2.87 $Y=1.12
+ $X2=2.525 $Y2=1.12
r227 15 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.45 $Y=3.075
+ $X2=2.525 $Y2=3.15
r228 14 44 12.1617 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=2.45 $Y=1.59
+ $X2=2.45 $Y2=1.317
r229 14 15 761.457 $w=1.5e-07 $l=1.485e-06 $layer=POLY_cond $X=2.45 $Y=1.59
+ $X2=2.45 $Y2=3.075
r230 11 42 37.0704 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.93 $Y=1.675
+ $X2=1.93 $Y2=1.467
r231 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.93 $Y=1.675
+ $X2=1.93 $Y2=2.31
r232 7 42 37.0704 $w=1.5e-07 $l=2.14369e-07 $layer=POLY_cond $X=1.915 $Y=1.26
+ $X2=1.93 $Y2=1.467
r233 7 9 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=1.915 $Y=1.26
+ $X2=1.915 $Y2=0.74
r234 2 62 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.12
+ $Y=1.75 $X2=1.255 $Y2=1.895
r235 1 56 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=1.125
+ $Y=0.37 $X2=1.27 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__DFSTP_1%A_1470_48# 1 2 9 12 13 15 18 21 22 23 25 32
+ 33 38
c90 21 0 1.66339e-19 $X=8.93 $Y=0.875
c91 9 0 7.26887e-20 $X=7.425 $Y=0.58
r92 32 33 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=9.28 $Y=2.815
+ $X2=9.28 $Y2=2.65
r93 27 33 94.5989 $w=1.68e-07 $l=1.45e-06 $layer=LI1_cond $X=9.36 $Y=1.2
+ $X2=9.36 $Y2=2.65
r94 23 27 12.9839 $w=2.49e-07 $l=3.52916e-07 $layer=LI1_cond $X=9.095 $Y=0.995
+ $X2=9.36 $Y2=1.2
r95 23 25 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=9.095 $Y=0.79
+ $X2=9.095 $Y2=0.58
r96 21 23 9.32073 $w=2.49e-07 $l=2.16852e-07 $layer=LI1_cond $X=8.93 $Y=0.875
+ $X2=9.095 $Y2=0.995
r97 21 22 78.2888 $w=1.68e-07 $l=1.2e-06 $layer=LI1_cond $X=8.93 $Y=0.875
+ $X2=7.73 $Y2=0.875
r98 19 38 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=7.615 $Y=1.39
+ $X2=7.63 $Y2=1.39
r99 19 35 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=7.615 $Y=1.39
+ $X2=7.425 $Y2=1.39
r100 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.615
+ $Y=1.39 $X2=7.615 $Y2=1.39
r101 16 22 7.04737 $w=1.7e-07 $l=1.54771e-07 $layer=LI1_cond $X=7.612 $Y=0.96
+ $X2=7.73 $Y2=0.875
r102 16 18 21.0873 $w=2.33e-07 $l=4.3e-07 $layer=LI1_cond $X=7.612 $Y=0.96
+ $X2=7.612 $Y2=1.39
r103 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.63 $Y=2.465
+ $X2=7.63 $Y2=2.75
r104 12 13 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=7.63 $Y=2.375
+ $X2=7.63 $Y2=2.465
r105 11 38 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.63 $Y=1.555
+ $X2=7.63 $Y2=1.39
r106 11 12 318.742 $w=1.8e-07 $l=8.2e-07 $layer=POLY_cond $X=7.63 $Y=1.555
+ $X2=7.63 $Y2=2.375
r107 7 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.425 $Y=1.225
+ $X2=7.425 $Y2=1.39
r108 7 9 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=7.425 $Y=1.225
+ $X2=7.425 $Y2=0.58
r109 2 32 600 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=9.13
+ $Y=2.54 $X2=9.28 $Y2=2.815
r110 1 25 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=8.955
+ $Y=0.37 $X2=9.095 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_LS__DFSTP_1%A_1298_392# 1 2 3 11 14 16 18 19 23 25 27 29
+ 30 32 35 38 39 43 45 46 47 50 52 56 57 61 63 64 68 72 74
c184 72 0 5.52031e-20 $X=6.9 $Y=1.715
c185 64 0 5.24842e-21 $X=6.642 $Y=2.05
c186 63 0 2.26502e-20 $X=6.645 $Y=2.155
c187 57 0 1.66339e-19 $X=8.94 $Y=1.535
r188 66 68 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=6.74 $Y=0.76 $X2=6.9
+ $Y2=0.76
r189 63 64 4.6525 $w=3.33e-07 $l=1.05e-07 $layer=LI1_cond $X=6.642 $Y=2.155
+ $X2=6.642 $Y2=2.05
r190 60 61 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=8.94
+ $Y=2.215 $X2=8.94 $Y2=2.215
r191 57 77 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=8.945 $Y=1.535
+ $X2=8.945 $Y2=1.37
r192 56 60 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=8.94 $Y=1.535
+ $X2=8.94 $Y2=2.215
r193 56 57 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=8.94
+ $Y=1.535 $X2=8.94 $Y2=1.535
r194 54 60 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=8.94 $Y=2.31
+ $X2=8.94 $Y2=2.215
r195 53 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.47 $Y=2.395
+ $X2=8.305 $Y2=2.395
r196 52 54 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.775 $Y=2.395
+ $X2=8.94 $Y2=2.31
r197 52 53 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=8.775 $Y=2.395
+ $X2=8.47 $Y2=2.395
r198 48 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.305 $Y=2.48
+ $X2=8.305 $Y2=2.395
r199 48 50 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=8.305 $Y=2.48
+ $X2=8.305 $Y2=2.765
r200 46 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.14 $Y=2.395
+ $X2=8.305 $Y2=2.395
r201 46 47 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=8.14 $Y=2.395
+ $X2=7.6 $Y2=2.395
r202 44 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.515 $Y=2.48
+ $X2=7.6 $Y2=2.395
r203 44 45 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=7.515 $Y=2.48
+ $X2=7.515 $Y2=2.625
r204 43 72 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.9 $Y=1.63 $X2=6.9
+ $Y2=1.715
r205 42 68 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.9 $Y=0.925
+ $X2=6.9 $Y2=0.76
r206 42 43 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=6.9 $Y=0.925
+ $X2=6.9 $Y2=1.63
r207 39 41 5.68106 $w=3.53e-07 $l=1.75e-07 $layer=LI1_cond $X=6.81 $Y=2.802
+ $X2=6.985 $Y2=2.802
r208 38 45 7.97992 $w=3.55e-07 $l=2.15346e-07 $layer=LI1_cond $X=7.43 $Y=2.802
+ $X2=7.515 $Y2=2.625
r209 38 41 14.4461 $w=3.53e-07 $l=4.45e-07 $layer=LI1_cond $X=7.43 $Y=2.802
+ $X2=6.985 $Y2=2.802
r210 36 72 13.5701 $w=1.68e-07 $l=2.08e-07 $layer=LI1_cond $X=6.692 $Y=1.715
+ $X2=6.9 $Y2=1.715
r211 36 64 12.26 $w=2.33e-07 $l=2.5e-07 $layer=LI1_cond $X=6.692 $Y=1.8
+ $X2=6.692 $Y2=2.05
r212 35 39 6.82394 $w=3.55e-07 $l=2.47113e-07 $layer=LI1_cond $X=6.642 $Y=2.625
+ $X2=6.81 $Y2=2.802
r213 34 63 2.13288 $w=3.33e-07 $l=6.2e-08 $layer=LI1_cond $X=6.642 $Y=2.217
+ $X2=6.642 $Y2=2.155
r214 34 35 14.0357 $w=3.33e-07 $l=4.08e-07 $layer=LI1_cond $X=6.642 $Y=2.217
+ $X2=6.642 $Y2=2.625
r215 31 32 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=9.87 $Y=1.865
+ $X2=10.025 $Y2=1.865
r216 30 61 2.54577 $w=3.4e-07 $l=1.5e-08 $layer=POLY_cond $X=8.945 $Y=2.23
+ $X2=8.945 $Y2=2.215
r217 28 61 46.6725 $w=3.4e-07 $l=2.75e-07 $layer=POLY_cond $X=8.945 $Y=1.94
+ $X2=8.945 $Y2=2.215
r218 28 29 9.89174 $w=3.4e-07 $l=7.5e-08 $layer=POLY_cond $X=8.945 $Y=1.94
+ $X2=8.945 $Y2=1.865
r219 25 32 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.025 $Y=1.94
+ $X2=10.025 $Y2=1.865
r220 25 27 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=10.025 $Y=1.94
+ $X2=10.025 $Y2=2.435
r221 21 31 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.87 $Y=1.79
+ $X2=9.87 $Y2=1.865
r222 21 23 587.117 $w=1.5e-07 $l=1.145e-06 $layer=POLY_cond $X=9.87 $Y=1.79
+ $X2=9.87 $Y2=0.645
r223 20 29 17.3855 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=9.115 $Y=1.865
+ $X2=8.945 $Y2=1.865
r224 19 31 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.795 $Y=1.865
+ $X2=9.87 $Y2=1.865
r225 19 20 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=9.795 $Y=1.865
+ $X2=9.115 $Y2=1.865
r226 16 30 37.6312 $w=3.01e-07 $l=2.84737e-07 $layer=POLY_cond $X=9.055 $Y=2.465
+ $X2=8.945 $Y2=2.23
r227 16 18 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=9.055 $Y=2.465
+ $X2=9.055 $Y2=2.75
r228 14 77 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=8.88 $Y=0.58
+ $X2=8.88 $Y2=1.37
r229 11 29 9.89174 $w=3.4e-07 $l=7.5e-08 $layer=POLY_cond $X=8.945 $Y=1.79
+ $X2=8.945 $Y2=1.865
r230 10 57 0.848592 $w=3.4e-07 $l=5e-09 $layer=POLY_cond $X=8.945 $Y=1.54
+ $X2=8.945 $Y2=1.535
r231 10 11 42.4296 $w=3.4e-07 $l=2.5e-07 $layer=POLY_cond $X=8.945 $Y=1.54
+ $X2=8.945 $Y2=1.79
r232 3 50 600 $w=1.7e-07 $l=2.90474e-07 $layer=licon1_PDIFF $count=1 $X=8.155
+ $Y=2.54 $X2=8.305 $Y2=2.765
r233 2 63 300 $w=1.7e-07 $l=2.61247e-07 $layer=licon1_PDIFF $count=2 $X=6.49
+ $Y=1.96 $X2=6.645 $Y2=2.155
r234 2 41 300 $w=1.7e-07 $l=1.09487e-06 $layer=licon1_PDIFF $count=2 $X=6.49
+ $Y=1.96 $X2=6.985 $Y2=2.835
r235 1 66 182 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_NDIFF $count=1 $X=6.6
+ $Y=0.37 $X2=6.74 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_LS__DFSTP_1%A_1902_74# 1 2 7 9 10 12 15 18 21 25 28 29
r55 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.35
+ $Y=1.385 $X2=10.35 $Y2=1.385
r56 23 29 0.466467 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=9.965 $Y=1.385
+ $X2=9.8 $Y2=1.385
r57 23 25 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=9.965 $Y=1.385
+ $X2=10.35 $Y2=1.385
r58 19 29 6.31733 $w=2.57e-07 $l=1.65e-07 $layer=LI1_cond $X=9.8 $Y=1.55 $X2=9.8
+ $Y2=1.385
r59 19 21 21.3027 $w=3.28e-07 $l=6.1e-07 $layer=LI1_cond $X=9.8 $Y=1.55 $X2=9.8
+ $Y2=2.16
r60 18 29 6.31733 $w=2.57e-07 $l=1.98167e-07 $layer=LI1_cond $X=9.727 $Y=1.22
+ $X2=9.8 $Y2=1.385
r61 18 28 21.5823 $w=1.83e-07 $l=3.6e-07 $layer=LI1_cond $X=9.727 $Y=1.22
+ $X2=9.727 $Y2=0.86
r62 13 28 7.96936 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=9.655 $Y=0.695
+ $X2=9.655 $Y2=0.86
r63 13 15 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=9.655 $Y=0.695
+ $X2=9.655 $Y2=0.605
r64 10 26 68.9212 $w=3.43e-07 $l=4.4238e-07 $layer=POLY_cond $X=10.545 $Y=1.765
+ $X2=10.41 $Y2=1.385
r65 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=10.545 $Y=1.765
+ $X2=10.545 $Y2=2.4
r66 7 26 38.7084 $w=3.43e-07 $l=1.83916e-07 $layer=POLY_cond $X=10.45 $Y=1.22
+ $X2=10.41 $Y2=1.385
r67 7 9 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=10.45 $Y=1.22 $X2=10.45
+ $Y2=0.74
r68 2 21 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=9.675
+ $Y=2.015 $X2=9.8 $Y2=2.16
r69 1 15 182 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_NDIFF $count=1 $X=9.51
+ $Y=0.37 $X2=9.655 $Y2=0.605
.ends

.subckt PM_SKY130_FD_SC_LS__DFSTP_1%A_27_74# 1 2 3 4 15 18 21 23 25 28 29 30 31
+ 36
c68 28 0 6.14252e-20 $X=2.572 $Y=2.06
c69 25 0 1.22961e-19 $X=2.485 $Y=2.145
r70 36 38 8.65635 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=2.61 $Y=0.76
+ $X2=2.61 $Y2=0.925
r71 31 33 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.675 $Y=2.145
+ $X2=1.675 $Y2=2.315
r72 28 38 71.9325 $w=1.73e-07 $l=1.135e-06 $layer=LI1_cond $X=2.572 $Y=2.06
+ $X2=2.572 $Y2=0.925
r73 26 31 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.76 $Y=2.145
+ $X2=1.675 $Y2=2.145
r74 25 41 13.515 $w=3.34e-07 $l=4.64047e-07 $layer=LI1_cond $X=2.485 $Y=2.145
+ $X2=2.697 $Y2=2.515
r75 25 28 5.85659 $w=3.34e-07 $l=1.22327e-07 $layer=LI1_cond $X=2.485 $Y=2.145
+ $X2=2.572 $Y2=2.06
r76 25 26 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=2.485 $Y=2.145
+ $X2=1.76 $Y2=2.145
r77 24 30 2.11342 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.355 $Y=2.315
+ $X2=0.23 $Y2=2.315
r78 23 33 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.59 $Y=2.315
+ $X2=1.675 $Y2=2.315
r79 23 24 80.5722 $w=1.68e-07 $l=1.235e-06 $layer=LI1_cond $X=1.59 $Y=2.315
+ $X2=0.355 $Y2=2.315
r80 19 30 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.23 $Y=2.4 $X2=0.23
+ $Y2=2.315
r81 19 21 16.1342 $w=2.48e-07 $l=3.5e-07 $layer=LI1_cond $X=0.23 $Y=2.4 $X2=0.23
+ $Y2=2.75
r82 18 30 4.3182 $w=2.1e-07 $l=1.03078e-07 $layer=LI1_cond $X=0.19 $Y=2.23
+ $X2=0.23 $Y2=2.315
r83 18 29 92.6417 $w=1.68e-07 $l=1.42e-06 $layer=LI1_cond $X=0.19 $Y=2.23
+ $X2=0.19 $Y2=0.81
r84 13 29 7.14225 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=0.235 $Y=0.68
+ $X2=0.235 $Y2=0.81
r85 13 15 4.43247 $w=2.58e-07 $l=1e-07 $layer=LI1_cond $X=0.235 $Y=0.68
+ $X2=0.235 $Y2=0.58
r86 4 41 600 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=1 $X=2.6
+ $Y=2.315 $X2=2.745 $Y2=2.515
r87 3 21 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.54 $X2=0.27 $Y2=2.75
r88 2 36 182 $w=1.7e-07 $l=4.48163e-07 $layer=licon1_NDIFF $count=1 $X=2.525
+ $Y=0.37 $X2=2.65 $Y2=0.76
r89 1 15 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_LS__DFSTP_1%VPWR 1 2 3 4 5 6 7 24 28 32 36 40 44 48 55
+ 56 58 59 60 62 67 72 93 97 104 105 108 111 114 117 120
r131 120 121 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r132 117 118 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r133 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r134 111 112 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r135 108 109 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r136 105 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=10.32 $Y2=3.33
r137 104 105 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r138 102 120 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.485 $Y=3.33
+ $X2=10.32 $Y2=3.33
r139 102 104 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=10.485 $Y=3.33
+ $X2=10.8 $Y2=3.33
r140 101 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=10.32 $Y2=3.33
r141 101 118 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=8.88 $Y2=3.33
r142 100 101 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r143 98 117 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.915 $Y=3.33
+ $X2=8.79 $Y2=3.33
r144 98 100 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=8.915 $Y=3.33
+ $X2=9.84 $Y2=3.33
r145 97 120 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.155 $Y=3.33
+ $X2=10.32 $Y2=3.33
r146 97 100 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=10.155 $Y=3.33
+ $X2=9.84 $Y2=3.33
r147 96 118 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=8.88 $Y2=3.33
r148 95 96 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r149 93 117 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.665 $Y=3.33
+ $X2=8.79 $Y2=3.33
r150 93 95 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=8.665 $Y=3.33
+ $X2=8.4 $Y2=3.33
r151 92 96 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=8.4 $Y2=3.33
r152 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r153 89 92 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=7.44 $Y2=3.33
r154 88 91 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=6 $Y=3.33 $X2=7.44
+ $Y2=3.33
r155 88 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r156 83 115 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r157 82 85 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r158 82 83 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r159 80 114 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=4.23 $Y=3.33
+ $X2=4.09 $Y2=3.33
r160 80 82 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=4.23 $Y=3.33
+ $X2=4.56 $Y2=3.33
r161 79 115 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r162 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r163 76 79 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.6 $Y2=3.33
r164 76 112 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r165 75 78 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=3.6 $Y2=3.33
r166 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r167 73 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.87 $Y=3.33
+ $X2=1.705 $Y2=3.33
r168 73 75 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.87 $Y=3.33
+ $X2=2.16 $Y2=3.33
r169 72 114 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=3.95 $Y=3.33
+ $X2=4.09 $Y2=3.33
r170 72 78 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=3.95 $Y=3.33
+ $X2=3.6 $Y2=3.33
r171 71 112 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r172 71 109 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r173 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r174 68 108 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.885 $Y=3.33
+ $X2=0.72 $Y2=3.33
r175 68 70 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.885 $Y=3.33
+ $X2=1.2 $Y2=3.33
r176 67 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.54 $Y=3.33
+ $X2=1.705 $Y2=3.33
r177 67 70 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.54 $Y=3.33
+ $X2=1.2 $Y2=3.33
r178 65 109 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r179 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r180 62 108 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.555 $Y=3.33
+ $X2=0.72 $Y2=3.33
r181 62 64 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.555 $Y=3.33
+ $X2=0.24 $Y2=3.33
r182 60 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33 $X2=6
+ $Y2=3.33
r183 60 83 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=4.56 $Y2=3.33
r184 60 85 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r185 58 91 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=7.77 $Y=3.33
+ $X2=7.44 $Y2=3.33
r186 58 59 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.77 $Y=3.33
+ $X2=7.855 $Y2=3.33
r187 57 95 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=7.94 $Y=3.33
+ $X2=8.4 $Y2=3.33
r188 57 59 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.94 $Y=3.33
+ $X2=7.855 $Y2=3.33
r189 55 85 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=5.535 $Y=3.33
+ $X2=5.52 $Y2=3.33
r190 55 56 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.535 $Y=3.33
+ $X2=5.66 $Y2=3.33
r191 54 88 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=5.785 $Y=3.33
+ $X2=6 $Y2=3.33
r192 54 56 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.785 $Y=3.33
+ $X2=5.66 $Y2=3.33
r193 51 53 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=10.32 $Y=2.4
+ $X2=10.32 $Y2=2.815
r194 48 51 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=10.32 $Y=1.985
+ $X2=10.32 $Y2=2.4
r195 46 120 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.32 $Y=3.245
+ $X2=10.32 $Y2=3.33
r196 46 53 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=10.32 $Y=3.245
+ $X2=10.32 $Y2=2.815
r197 42 117 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.79 $Y=3.245
+ $X2=8.79 $Y2=3.33
r198 42 44 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=8.79 $Y=3.245
+ $X2=8.79 $Y2=2.815
r199 38 59 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.855 $Y=3.245
+ $X2=7.855 $Y2=3.33
r200 38 40 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=7.855 $Y=3.245
+ $X2=7.855 $Y2=2.815
r201 34 56 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.66 $Y=3.245
+ $X2=5.66 $Y2=3.33
r202 34 36 19.361 $w=2.48e-07 $l=4.2e-07 $layer=LI1_cond $X=5.66 $Y=3.245
+ $X2=5.66 $Y2=2.825
r203 30 114 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=4.09 $Y=3.245
+ $X2=4.09 $Y2=3.33
r204 30 32 26.9589 $w=2.78e-07 $l=6.55e-07 $layer=LI1_cond $X=4.09 $Y=3.245
+ $X2=4.09 $Y2=2.59
r205 26 111 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.705 $Y=3.245
+ $X2=1.705 $Y2=3.33
r206 26 28 19.382 $w=3.28e-07 $l=5.55e-07 $layer=LI1_cond $X=1.705 $Y=3.245
+ $X2=1.705 $Y2=2.69
r207 22 108 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.72 $Y=3.245
+ $X2=0.72 $Y2=3.33
r208 22 24 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=0.72 $Y=3.245
+ $X2=0.72 $Y2=2.775
r209 7 53 600 $w=1.7e-07 $l=9.03327e-07 $layer=licon1_PDIFF $count=1 $X=10.1
+ $Y=2.015 $X2=10.32 $Y2=2.815
r210 7 51 600 $w=1.7e-07 $l=4.82623e-07 $layer=licon1_PDIFF $count=1 $X=10.1
+ $Y=2.015 $X2=10.32 $Y2=2.4
r211 7 48 600 $w=1.7e-07 $l=2.34521e-07 $layer=licon1_PDIFF $count=1 $X=10.1
+ $Y=2.015 $X2=10.32 $Y2=1.985
r212 6 44 600 $w=1.7e-07 $l=3.33729e-07 $layer=licon1_PDIFF $count=1 $X=8.7
+ $Y=2.54 $X2=8.83 $Y2=2.815
r213 5 40 600 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=7.705
+ $Y=2.54 $X2=7.855 $Y2=2.815
r214 4 36 600 $w=1.7e-07 $l=6.73721e-07 $layer=licon1_PDIFF $count=1 $X=5.24
+ $Y=2.315 $X2=5.62 $Y2=2.825
r215 3 32 600 $w=1.7e-07 $l=3.47851e-07 $layer=licon1_PDIFF $count=1 $X=3.965
+ $Y=2.315 $X2=4.13 $Y2=2.59
r216 2 28 600 $w=1.7e-07 $l=1.01223e-06 $layer=licon1_PDIFF $count=1 $X=1.555
+ $Y=1.75 $X2=1.705 $Y2=2.69
r217 1 24 600 $w=1.7e-07 $l=3.00791e-07 $layer=licon1_PDIFF $count=1 $X=0.57
+ $Y=2.54 $X2=0.72 $Y2=2.775
.ends

.subckt PM_SKY130_FD_SC_LS__DFSTP_1%Q 1 2 7 8 9 10 11 12 13 23
r18 12 13 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=10.81 $Y=2.405
+ $X2=10.81 $Y2=2.775
r19 11 12 19.361 $w=2.48e-07 $l=4.2e-07 $layer=LI1_cond $X=10.81 $Y=1.985
+ $X2=10.81 $Y2=2.405
r20 10 11 14.7513 $w=2.48e-07 $l=3.2e-07 $layer=LI1_cond $X=10.81 $Y=1.665
+ $X2=10.81 $Y2=1.985
r21 9 10 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=10.81 $Y=1.295
+ $X2=10.81 $Y2=1.665
r22 9 43 11.2939 $w=2.48e-07 $l=2.45e-07 $layer=LI1_cond $X=10.81 $Y=1.295
+ $X2=10.81 $Y2=1.05
r23 8 43 5.37855 $w=4.33e-07 $l=1.25e-07 $layer=LI1_cond $X=10.717 $Y=0.925
+ $X2=10.717 $Y2=1.05
r24 8 21 2.43735 $w=4.33e-07 $l=9.2e-08 $layer=LI1_cond $X=10.717 $Y=0.925
+ $X2=10.717 $Y2=0.833
r25 7 21 7.36504 $w=4.33e-07 $l=2.78e-07 $layer=LI1_cond $X=10.717 $Y=0.555
+ $X2=10.717 $Y2=0.833
r26 7 23 1.05972 $w=4.33e-07 $l=4e-08 $layer=LI1_cond $X=10.717 $Y=0.555
+ $X2=10.717 $Y2=0.515
r27 2 13 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=10.62
+ $Y=1.84 $X2=10.77 $Y2=2.815
r28 2 11 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=10.62
+ $Y=1.84 $X2=10.77 $Y2=1.985
r29 1 23 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.525
+ $Y=0.37 $X2=10.665 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__DFSTP_1%VGND 1 2 3 4 5 6 21 23 27 31 35 39 44 45 47
+ 48 49 51 56 80 81 84 87 90 95 101
c116 27 0 9.68091e-20 $X=1.7 $Y=0.495
r117 100 101 10.7086 $w=6.83e-07 $l=1.65e-07 $layer=LI1_cond $X=8.595 $Y=0.257
+ $X2=8.76 $Y2=0.257
r118 97 100 3.40489 $w=6.83e-07 $l=1.95e-07 $layer=LI1_cond $X=8.4 $Y=0.257
+ $X2=8.595 $Y2=0.257
r119 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r120 94 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.4
+ $Y2=0
r121 93 97 8.38128 $w=6.83e-07 $l=4.8e-07 $layer=LI1_cond $X=7.92 $Y=0.257
+ $X2=8.4 $Y2=0.257
r122 93 95 8.70061 $w=6.83e-07 $l=5e-08 $layer=LI1_cond $X=7.92 $Y=0.257
+ $X2=7.87 $Y2=0.257
r123 93 94 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r124 90 91 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r125 87 88 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r126 85 88 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r127 84 85 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r128 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.8 $Y=0 $X2=10.8
+ $Y2=0
r129 78 81 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.84 $Y=0 $X2=10.8
+ $Y2=0
r130 77 78 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r131 75 78 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=9.84
+ $Y2=0
r132 75 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=8.4
+ $Y2=0
r133 74 77 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=8.88 $Y=0 $X2=9.84
+ $Y2=0
r134 74 101 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=8.88 $Y=0 $X2=8.76
+ $Y2=0
r135 74 75 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r136 71 94 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6 $Y=0 $X2=7.92
+ $Y2=0
r137 70 95 122 $w=1.68e-07 $l=1.87e-06 $layer=LI1_cond $X=6 $Y=0 $X2=7.87 $Y2=0
r138 70 71 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6
+ $Y2=0
r139 64 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r140 63 66 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.56 $Y=0 $X2=5.52
+ $Y2=0
r141 63 64 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r142 61 90 9.6488 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=4.455 $Y=0 $X2=4.26
+ $Y2=0
r143 61 63 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=4.455 $Y=0
+ $X2=4.56 $Y2=0
r144 60 91 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=4.08 $Y2=0
r145 60 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r146 59 60 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r147 57 87 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.785 $Y=0 $X2=1.7
+ $Y2=0
r148 57 59 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.785 $Y=0
+ $X2=2.16 $Y2=0
r149 56 90 9.6488 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=4.065 $Y=0 $X2=4.26
+ $Y2=0
r150 56 59 124.283 $w=1.68e-07 $l=1.905e-06 $layer=LI1_cond $X=4.065 $Y=0
+ $X2=2.16 $Y2=0
r151 54 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r152 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r153 51 84 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.67
+ $Y2=0
r154 51 53 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0
+ $X2=0.24 $Y2=0
r155 49 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r156 49 64 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=4.56
+ $Y2=0
r157 49 66 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r158 47 77 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=10 $Y=0 $X2=9.84
+ $Y2=0
r159 47 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10 $Y=0 $X2=10.165
+ $Y2=0
r160 46 80 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=10.33 $Y=0 $X2=10.8
+ $Y2=0
r161 46 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.33 $Y=0
+ $X2=10.165 $Y2=0
r162 44 66 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=5.62 $Y=0 $X2=5.52
+ $Y2=0
r163 44 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.62 $Y=0 $X2=5.785
+ $Y2=0
r164 43 70 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=5.95 $Y=0 $X2=6 $Y2=0
r165 43 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.95 $Y=0 $X2=5.785
+ $Y2=0
r166 39 41 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=10.165 $Y=0.495
+ $X2=10.165 $Y2=0.93
r167 37 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.165 $Y=0.085
+ $X2=10.165 $Y2=0
r168 37 39 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=10.165 $Y=0.085
+ $X2=10.165 $Y2=0.495
r169 33 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.785 $Y=0.085
+ $X2=5.785 $Y2=0
r170 33 35 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=5.785 $Y=0.085
+ $X2=5.785 $Y2=0.515
r171 29 90 1.39532 $w=3.9e-07 $l=8.5e-08 $layer=LI1_cond $X=4.26 $Y=0.085
+ $X2=4.26 $Y2=0
r172 29 31 12.7064 $w=3.88e-07 $l=4.3e-07 $layer=LI1_cond $X=4.26 $Y=0.085
+ $X2=4.26 $Y2=0.515
r173 25 87 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.7 $Y=0.085 $X2=1.7
+ $Y2=0
r174 25 27 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=1.7 $Y=0.085
+ $X2=1.7 $Y2=0.495
r175 24 84 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.795 $Y=0 $X2=0.67
+ $Y2=0
r176 23 87 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.615 $Y=0 $X2=1.7
+ $Y2=0
r177 23 24 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=1.615 $Y=0
+ $X2=0.795 $Y2=0
r178 19 84 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.67 $Y=0.085
+ $X2=0.67 $Y2=0
r179 19 21 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=0.67 $Y=0.085
+ $X2=0.67 $Y2=0.58
r180 6 41 182 $w=1.7e-07 $l=6.60908e-07 $layer=licon1_NDIFF $count=1 $X=9.945
+ $Y=0.37 $X2=10.165 $Y2=0.93
r181 6 39 182 $w=1.7e-07 $l=2.755e-07 $layer=licon1_NDIFF $count=1 $X=9.945
+ $Y=0.37 $X2=10.165 $Y2=0.495
r182 5 100 91 $w=1.7e-07 $l=7.74112e-07 $layer=licon1_NDIFF $count=2 $X=7.89
+ $Y=0.37 $X2=8.595 $Y2=0.515
r183 4 35 91 $w=1.7e-07 $l=3.25346e-07 $layer=licon1_NDIFF $count=2 $X=5.495
+ $Y=0.59 $X2=5.785 $Y2=0.515
r184 3 31 182 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_NDIFF $count=1 $X=4.09
+ $Y=0.37 $X2=4.26 $Y2=0.515
r185 2 27 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.56
+ $Y=0.37 $X2=1.7 $Y2=0.495
r186 1 21 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.58
.ends

