* File: sky130_fd_sc_ls__o2111ai_1.spice
* Created: Wed Sep  2 11:16:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__o2111ai_1.pex.spice"
.subckt sky130_fd_sc_ls__o2111ai_1  VNB VPB D1 C1 B1 A2 A1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A1	A1
* A2	A2
* B1	B1
* C1	C1
* D1	D1
* VPB	VPB
* VNB	VNB
MM1006 A_182_74# N_D1_M1006_g N_Y_M1006_s VNB NSHORT L=0.15 W=0.74 AD=0.0888
+ AS=0.4625 PD=0.98 PS=2.73 NRD=10.536 NRS=0 M=1 R=4.93333 SA=75000.6 SB=75002.2
+ A=0.111 P=1.78 MULT=1
MM1007 A_260_74# N_C1_M1007_g A_182_74# VNB NSHORT L=0.15 W=0.74 AD=0.1443
+ AS=0.0888 PD=1.13 PS=0.98 NRD=22.692 NRS=10.536 M=1 R=4.93333 SA=75000.9
+ SB=75001.8 A=0.111 P=1.78 MULT=1
MM1001 N_A_368_74#_M1001_d N_B1_M1001_g A_260_74# VNB NSHORT L=0.15 W=0.74
+ AD=0.1332 AS=0.1443 PD=1.1 PS=1.13 NRD=1.62 NRS=22.692 M=1 R=4.93333
+ SA=75001.5 SB=75001.3 A=0.111 P=1.78 MULT=1
MM1002 N_VGND_M1002_d N_A2_M1002_g N_A_368_74#_M1001_d VNB NSHORT L=0.15 W=0.74
+ AD=0.1628 AS=0.1332 PD=1.18 PS=1.1 NRD=7.296 NRS=11.34 M=1 R=4.93333 SA=75002
+ SB=75000.8 A=0.111 P=1.78 MULT=1
MM1004 N_A_368_74#_M1004_d N_A1_M1004_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.1628 PD=2.05 PS=1.18 NRD=0 NRS=18.648 M=1 R=4.93333 SA=75002.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1003 N_Y_M1003_d N_D1_M1003_g N_VPWR_M1003_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.3864 PD=1.42 PS=2.93 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75000.3 SB=75002.2 A=0.168 P=2.54 MULT=1
MM1005 N_VPWR_M1005_d N_C1_M1005_g N_Y_M1003_d VPB PHIGHVT L=0.15 W=1.12
+ AD=0.2688 AS=0.168 PD=1.6 PS=1.42 NRD=29.0181 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75001.8 A=0.168 P=2.54 MULT=1
MM1000 N_Y_M1000_d N_B1_M1000_g N_VPWR_M1005_d VPB PHIGHVT L=0.15 W=1.12
+ AD=0.182 AS=0.2688 PD=1.445 PS=1.6 NRD=6.1464 NRS=6.1464 M=1 R=7.46667
+ SA=75001.3 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1008 A_490_368# N_A2_M1008_g N_Y_M1000_d VPB PHIGHVT L=0.15 W=1.12 AD=0.1708
+ AS=0.182 PD=1.425 PS=1.445 NRD=17.139 NRS=1.7533 M=1 R=7.46667 SA=75001.8
+ SB=75000.7 A=0.168 P=2.54 MULT=1
MM1009 N_VPWR_M1009_d N_A1_M1009_g A_490_368# VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.1708 PD=2.83 PS=1.425 NRD=1.7533 NRS=17.139 M=1 R=7.46667
+ SA=75002.3 SB=75000.2 A=0.168 P=2.54 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9564 P=11.2
*
.include "sky130_fd_sc_ls__o2111ai_1.pxi.spice"
*
.ends
*
*
