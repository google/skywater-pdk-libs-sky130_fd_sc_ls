* File: sky130_fd_sc_ls__sdfrtn_1.pex.spice
* Created: Wed Sep  2 11:27:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__SDFRTN_1%SCE 3 6 7 9 12 15 22 23 25 26 27 33 35
c68 22 0 8.65763e-20 $X=0.7 $Y=1.575
r69 32 35 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=2.385 $Y=1.12
+ $X2=2.615 $Y2=1.12
r70 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.385
+ $Y=1.12 $X2=2.385 $Y2=1.12
r71 27 33 5.91467 $w=4.53e-07 $l=2.25e-07 $layer=LI1_cond $X=2.16 $Y=1.182
+ $X2=2.385 $Y2=1.182
r72 26 27 3.02306 $w=4.53e-07 $l=1.15e-07 $layer=LI1_cond $X=2.045 $Y=1.182
+ $X2=2.16 $Y2=1.182
r73 25 26 9.38335 $w=4.53e-07 $l=1.7e-07 $layer=LI1_cond $X=1.875 $Y=1.267
+ $X2=2.045 $Y2=1.267
r74 23 30 46.8028 $w=4.45e-07 $l=1.65e-07 $layer=POLY_cond $X=0.642 $Y=1.575
+ $X2=0.642 $Y2=1.41
r75 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.7
+ $Y=1.575 $X2=0.7 $Y2=1.575
r76 20 22 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.865 $Y=1.495
+ $X2=0.7 $Y2=1.495
r77 20 25 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=0.865 $Y=1.495
+ $X2=1.875 $Y2=1.495
r78 13 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.615 $Y=0.955
+ $X2=2.615 $Y2=1.12
r79 13 15 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=2.615 $Y=0.955
+ $X2=2.615 $Y2=0.615
r80 7 12 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.955 $Y=2.245
+ $X2=0.955 $Y2=2.64
r81 7 9 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.505 $Y=2.245
+ $X2=0.505 $Y2=2.64
r82 6 7 31.2407 $w=4.86e-07 $l=4.4477e-07 $layer=POLY_cond $X=0.642 $Y=1.93
+ $X2=0.955 $Y2=2.245
r83 5 23 7.12377 $w=4.45e-07 $l=5.7e-08 $layer=POLY_cond $X=0.642 $Y=1.632
+ $X2=0.642 $Y2=1.575
r84 5 6 37.2436 $w=4.45e-07 $l=2.98e-07 $layer=POLY_cond $X=0.642 $Y=1.632
+ $X2=0.642 $Y2=1.93
r85 3 30 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=0.495 $Y=0.65
+ $X2=0.495 $Y2=1.41
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTN_1%A_27_88# 1 2 9 11 12 14 17 20 23 25 31 32
+ 34 35 37 38 39 42
c92 11 0 1.86156e-19 $X=2.28 $Y=2.155
r93 38 42 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.455 $Y=1.1
+ $X2=1.455 $Y2=0.935
r94 37 39 7.86356 $w=3.03e-07 $l=1.65e-07 $layer=LI1_cond $X=1.455 $Y=1.087
+ $X2=1.29 $Y2=1.087
r95 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.455
+ $Y=1.1 $X2=1.455 $Y2=1.1
r96 32 44 17.4861 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=2.38 $Y=1.72 $X2=2.28
+ $Y2=1.72
r97 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.38
+ $Y=1.72 $X2=2.38 $Y2=1.72
r98 29 31 19.9058 $w=3.28e-07 $l=5.7e-07 $layer=LI1_cond $X=2.38 $Y=2.29
+ $X2=2.38 $Y2=1.72
r99 28 34 2.90107 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=0.445 $Y=1.145
+ $X2=0.28 $Y2=1.145
r100 28 39 49.3254 $w=1.88e-07 $l=8.45e-07 $layer=LI1_cond $X=0.445 $Y=1.145
+ $X2=1.29 $Y2=1.145
r101 26 35 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.365 $Y=2.375
+ $X2=0.24 $Y2=2.375
r102 25 29 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.215 $Y=2.375
+ $X2=2.38 $Y2=2.29
r103 25 26 120.695 $w=1.68e-07 $l=1.85e-06 $layer=LI1_cond $X=2.215 $Y=2.375
+ $X2=0.365 $Y2=2.375
r104 21 35 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.24 $Y=2.46
+ $X2=0.24 $Y2=2.375
r105 21 23 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=0.24 $Y=2.46
+ $X2=0.24 $Y2=2.465
r106 20 35 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.24 $Y=2.29
+ $X2=0.24 $Y2=2.375
r107 19 34 3.58697 $w=2.9e-07 $l=1.13248e-07 $layer=LI1_cond $X=0.24 $Y=1.24
+ $X2=0.28 $Y2=1.145
r108 19 20 48.4026 $w=2.48e-07 $l=1.05e-06 $layer=LI1_cond $X=0.24 $Y=1.24
+ $X2=0.24 $Y2=2.29
r109 15 34 3.58697 $w=2.9e-07 $l=9.5e-08 $layer=LI1_cond $X=0.28 $Y=1.05
+ $X2=0.28 $Y2=1.145
r110 15 17 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=0.28 $Y=1.05 $X2=0.28
+ $Y2=0.65
r111 12 14 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.28 $Y=2.245
+ $X2=2.28 $Y2=2.64
r112 11 12 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.28 $Y=2.155
+ $X2=2.28 $Y2=2.245
r113 10 44 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.28 $Y=1.885
+ $X2=2.28 $Y2=1.72
r114 10 11 104.952 $w=1.8e-07 $l=2.7e-07 $layer=POLY_cond $X=2.28 $Y=1.885
+ $X2=2.28 $Y2=2.155
r115 9 42 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.545 $Y=0.615
+ $X2=1.545 $Y2=0.935
r116 2 23 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.32 $X2=0.28 $Y2=2.465
r117 1 17 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.44 $X2=0.28 $Y2=0.65
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTN_1%D 1 3 4 8 10 12 13 17 18
c40 18 0 1.86156e-19 $X=1.815 $Y=1.945
c41 10 0 8.65763e-20 $X=1.345 $Y=2.035
r42 17 20 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.815 $Y=1.945
+ $X2=1.815 $Y2=2.035
r43 17 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.815 $Y=1.945
+ $X2=1.815 $Y2=1.78
r44 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.815
+ $Y=1.945 $X2=1.815 $Y2=1.945
r45 13 18 4.57588 $w=3.38e-07 $l=1.35e-07 $layer=LI1_cond $X=1.68 $Y=1.95
+ $X2=1.815 $Y2=1.95
r46 12 13 16.2698 $w=3.38e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.95 $X2=1.68
+ $Y2=1.95
r47 8 19 597.372 $w=1.5e-07 $l=1.165e-06 $layer=POLY_cond $X=1.905 $Y=0.615
+ $X2=1.905 $Y2=1.78
r48 5 10 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=1.435 $Y=2.035 $X2=1.345
+ $Y2=2.035
r49 4 20 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.65 $Y=2.035
+ $X2=1.815 $Y2=2.035
r50 4 5 110.245 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=1.65 $Y=2.035
+ $X2=1.435 $Y2=2.035
r51 1 10 83.7788 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=1.345 $Y=2.245
+ $X2=1.345 $Y2=2.035
r52 1 3 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.345 $Y=2.245
+ $X2=1.345 $Y2=2.64
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTN_1%SCD 1 3 5 8 12 14 15 19
c51 5 0 1.38402e-19 $X=2.875 $Y=2.095
r52 19 22 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.965 $Y=1.69
+ $X2=2.965 $Y2=1.855
r53 19 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.965 $Y=1.69
+ $X2=2.965 $Y2=1.525
r54 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.965
+ $Y=1.69 $X2=2.965 $Y2=1.69
r55 15 20 9.14007 $w=4.33e-07 $l=3.45e-07 $layer=LI1_cond $X=3.017 $Y=2.035
+ $X2=3.017 $Y2=1.69
r56 14 20 0.662324 $w=4.33e-07 $l=2.5e-08 $layer=LI1_cond $X=3.017 $Y=1.665
+ $X2=3.017 $Y2=1.69
r57 10 12 105.117 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=2.67 $Y=2.17
+ $X2=2.875 $Y2=2.17
r58 8 21 466.617 $w=1.5e-07 $l=9.1e-07 $layer=POLY_cond $X=3.005 $Y=0.615
+ $X2=3.005 $Y2=1.525
r59 5 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.875 $Y=2.095
+ $X2=2.875 $Y2=2.17
r60 5 22 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=2.875 $Y=2.095
+ $X2=2.875 $Y2=1.855
r61 1 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.67 $Y=2.245
+ $X2=2.67 $Y2=2.17
r62 1 3 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.67 $Y=2.245
+ $X2=2.67 $Y2=2.64
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTN_1%CLK_N 1 3 6 8 9 10
c39 10 0 6.18507e-21 $X=4.56 $Y=1.295
c40 6 0 2.04547e-19 $X=4.72 $Y=2.235
r41 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.44
+ $Y=1.385 $X2=4.44 $Y2=1.385
r42 10 14 4.06745 $w=3.38e-07 $l=1.2e-07 $layer=LI1_cond $X=4.56 $Y=1.38
+ $X2=4.44 $Y2=1.38
r43 9 13 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=4.645 $Y=1.385
+ $X2=4.44 $Y2=1.385
r44 8 13 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=4.27 $Y=1.385
+ $X2=4.44 $Y2=1.385
r45 4 9 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=4.72 $Y=1.55
+ $X2=4.645 $Y2=1.385
r46 4 6 351.245 $w=1.5e-07 $l=6.85e-07 $layer=POLY_cond $X=4.72 $Y=1.55 $X2=4.72
+ $Y2=2.235
r47 1 8 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=4.195 $Y=1.22
+ $X2=4.27 $Y2=1.385
r48 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.195 $Y=1.22 $X2=4.195
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTN_1%A_1049_347# 1 2 7 9 12 15 16 18 19 21 23 25
+ 27 28 32 33 34 37 38 39 43 46 49 51 52 53 55 67
c183 27 0 1.4087e-19 $X=5.55 $Y=1.735
c184 12 0 1.13453e-19 $X=6.63 $Y=2.525
c185 7 0 1.7914e-19 $X=6.285 $Y=0.505
r186 59 70 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.66 $Y=1.065
+ $X2=9.66 $Y2=1.23
r187 59 67 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=9.66 $Y=1.065
+ $X2=9.66 $Y2=0.94
r188 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.66
+ $Y=1.065 $X2=9.66 $Y2=1.065
r189 55 58 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=9.66 $Y=0.875
+ $X2=9.66 $Y2=1.065
r190 51 53 5.33982 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=6.63 $Y=1.9
+ $X2=6.495 $Y2=1.9
r191 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.63
+ $Y=1.9 $X2=6.63 $Y2=1.9
r192 49 61 34.7923 $w=3.4e-07 $l=2.05e-07 $layer=POLY_cond $X=6.49 $Y=0.335
+ $X2=6.285 $Y2=0.335
r193 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.49
+ $Y=0.34 $X2=6.49 $Y2=0.34
r194 43 45 4.02231 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=5.51 $Y=0.99
+ $X2=5.51 $Y2=1.085
r195 38 55 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.495 $Y=0.875
+ $X2=9.66 $Y2=0.875
r196 38 39 115.802 $w=1.68e-07 $l=1.775e-06 $layer=LI1_cond $X=9.495 $Y=0.875
+ $X2=7.72 $Y2=0.875
r197 37 39 6.9898 $w=1.7e-07 $l=1.49579e-07 $layer=LI1_cond $X=7.607 $Y=0.79
+ $X2=7.72 $Y2=0.875
r198 36 37 12.5488 $w=2.23e-07 $l=2.45e-07 $layer=LI1_cond $X=7.607 $Y=0.545
+ $X2=7.607 $Y2=0.79
r199 35 48 2.74877 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.495 $Y=0.4
+ $X2=6.41 $Y2=0.4
r200 34 36 6.95868 $w=2.9e-07 $l=1.93041e-07 $layer=LI1_cond $X=7.495 $Y=0.4
+ $X2=7.607 $Y2=0.545
r201 34 35 39.7394 $w=2.88e-07 $l=1e-06 $layer=LI1_cond $X=7.495 $Y=0.4
+ $X2=6.495 $Y2=0.4
r202 32 48 4.68908 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=6.41 $Y=0.545
+ $X2=6.41 $Y2=0.4
r203 32 33 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=6.41 $Y=0.545
+ $X2=6.41 $Y2=1.265
r204 31 41 3.39346 $w=2.55e-07 $l=2.23e-07 $layer=LI1_cond $X=5.675 $Y=1.862
+ $X2=5.452 $Y2=1.862
r205 31 53 37.059 $w=2.53e-07 $l=8.2e-07 $layer=LI1_cond $X=5.675 $Y=1.862
+ $X2=6.495 $Y2=1.862
r206 29 46 2.15711 $w=2e-07 $l=1.25e-07 $layer=LI1_cond $X=5.675 $Y=1.365
+ $X2=5.55 $Y2=1.365
r207 28 33 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=6.325 $Y=1.365
+ $X2=6.41 $Y2=1.265
r208 28 29 36.0455 $w=1.98e-07 $l=6.5e-07 $layer=LI1_cond $X=6.325 $Y=1.365
+ $X2=5.675 $Y2=1.365
r209 27 41 3.4239 $w=2.5e-07 $l=1.69041e-07 $layer=LI1_cond $X=5.55 $Y=1.735
+ $X2=5.452 $Y2=1.862
r210 26 46 4.27425 $w=2.5e-07 $l=1e-07 $layer=LI1_cond $X=5.55 $Y=1.465 $X2=5.55
+ $Y2=1.365
r211 26 27 12.4464 $w=2.48e-07 $l=2.7e-07 $layer=LI1_cond $X=5.55 $Y=1.465
+ $X2=5.55 $Y2=1.735
r212 25 46 4.27425 $w=2.5e-07 $l=1e-07 $layer=LI1_cond $X=5.55 $Y=1.265 $X2=5.55
+ $Y2=1.365
r213 25 45 8.29759 $w=2.48e-07 $l=1.8e-07 $layer=LI1_cond $X=5.55 $Y=1.265
+ $X2=5.55 $Y2=1.085
r214 21 23 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=10.29 $Y=0.865
+ $X2=10.29 $Y2=0.58
r215 20 67 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.825 $Y=0.94
+ $X2=9.66 $Y2=0.94
r216 19 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.215 $Y=0.94
+ $X2=10.29 $Y2=0.865
r217 19 20 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=10.215 $Y=0.94
+ $X2=9.825 $Y2=0.94
r218 16 18 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=9.62 $Y=1.885
+ $X2=9.62 $Y2=2.46
r219 15 16 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=9.62 $Y=1.795
+ $X2=9.62 $Y2=1.885
r220 15 70 219.621 $w=1.8e-07 $l=5.65e-07 $layer=POLY_cond $X=9.62 $Y=1.795
+ $X2=9.62 $Y2=1.23
r221 10 52 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.63 $Y=2.065
+ $X2=6.63 $Y2=1.9
r222 10 12 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=6.63 $Y=2.065
+ $X2=6.63 $Y2=2.525
r223 7 61 21.9347 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=6.285 $Y=0.505
+ $X2=6.285 $Y2=0.335
r224 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.285 $Y=0.505
+ $X2=6.285 $Y2=0.825
r225 2 41 600 $w=1.7e-07 $l=2.33238e-07 $layer=licon1_PDIFF $count=1 $X=5.245
+ $Y=1.735 $X2=5.395 $Y2=1.905
r226 1 43 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=5.37
+ $Y=0.395 $X2=5.51 $Y2=0.99
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTN_1%A_1402_308# 1 2 9 13 17 20 21 22 26 31 32
+ 37
c96 37 0 1.50769e-20 $X=7.37 $Y=1.705
c97 31 0 1.69146e-19 $X=8.96 $Y=2.135
c98 17 0 1.5858e-20 $X=7.31 $Y=1.705
c99 13 0 8.36181e-20 $X=7.37 $Y=0.825
r100 31 33 0.276272 $w=8.73e-07 $l=5e-09 $layer=LI1_cond $X=9.127 $Y=2.135
+ $X2=9.127 $Y2=2.14
r101 31 32 12.1237 $w=8.73e-07 $l=1.65e-07 $layer=LI1_cond $X=9.127 $Y=2.135
+ $X2=9.127 $Y2=1.97
r102 26 33 10.4851 $w=7.68e-07 $l=6.75e-07 $layer=LI1_cond $X=9.18 $Y=2.815
+ $X2=9.18 $Y2=2.14
r103 22 29 3.40825 $w=1.7e-07 $l=1.16619e-07 $layer=LI1_cond $X=8.775 $Y=1.3
+ $X2=8.85 $Y2=1.215
r104 22 32 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.775 $Y=1.3
+ $X2=8.775 $Y2=1.97
r105 20 29 3.40825 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=8.69 $Y=1.215
+ $X2=8.85 $Y2=1.215
r106 20 21 79.2674 $w=1.68e-07 $l=1.215e-06 $layer=LI1_cond $X=8.69 $Y=1.215
+ $X2=7.475 $Y2=1.215
r107 18 37 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=7.31 $Y=1.705
+ $X2=7.37 $Y2=1.705
r108 18 34 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=7.31 $Y=1.705
+ $X2=7.085 $Y2=1.705
r109 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.31
+ $Y=1.705 $X2=7.31 $Y2=1.705
r110 15 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=7.35 $Y=1.3
+ $X2=7.475 $Y2=1.215
r111 15 17 18.6696 $w=2.48e-07 $l=4.05e-07 $layer=LI1_cond $X=7.35 $Y=1.3
+ $X2=7.35 $Y2=1.705
r112 11 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.37 $Y=1.54
+ $X2=7.37 $Y2=1.705
r113 11 13 366.628 $w=1.5e-07 $l=7.15e-07 $layer=POLY_cond $X=7.37 $Y=1.54
+ $X2=7.37 $Y2=0.825
r114 7 34 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.085 $Y=1.87
+ $X2=7.085 $Y2=1.705
r115 7 9 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=7.085 $Y=1.87
+ $X2=7.085 $Y2=2.525
r116 2 31 200 $w=1.7e-07 $l=2.73861e-07 $layer=licon1_PDIFF $count=3 $X=8.76
+ $Y=1.96 $X2=8.96 $Y2=2.135
r117 2 26 200 $w=1.7e-07 $l=9.4975e-07 $layer=licon1_PDIFF $count=3 $X=8.76
+ $Y=1.96 $X2=8.96 $Y2=2.815
r118 1 29 182 $w=1.7e-07 $l=6.19375e-07 $layer=licon1_NDIFF $count=1 $X=8.425
+ $Y=0.72 $X2=8.705 $Y2=1.215
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTN_1%RESET_B 4 5 6 9 12 16 19 22 25 28 29 31 34
+ 36 38 39 40 41 46 49 52 53 56 57 61 62
c243 61 0 1.97052e-19 $X=11.16 $Y=1.375
c244 57 0 8.36181e-20 $X=7.85 $Y=1.635
c245 53 0 1.38402e-19 $X=3.57 $Y=1.52
c246 36 0 2.78046e-19 $X=11.25 $Y=2.375
c247 34 0 1.5858e-20 $X=7.76 $Y=2.16
r248 61 64 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=11.16 $Y=1.375
+ $X2=11.16 $Y2=1.54
r249 61 63 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=11.16 $Y=1.375
+ $X2=11.16 $Y2=1.21
r250 61 62 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.16
+ $Y=1.375 $X2=11.16 $Y2=1.375
r251 56 59 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.85 $Y=1.635
+ $X2=7.85 $Y2=1.8
r252 56 58 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.85 $Y=1.635
+ $X2=7.85 $Y2=1.47
r253 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.85
+ $Y=1.635 $X2=7.85 $Y2=1.635
r254 52 54 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=3.552 $Y=1.52
+ $X2=3.552 $Y2=1.355
r255 52 53 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.57
+ $Y=1.52 $X2=3.57 $Y2=1.52
r256 49 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=1.665
+ $X2=3.6 $Y2=1.665
r257 47 62 11.2317 $w=3.15e-07 $l=2.9e-07 $layer=LI1_cond $X=11.195 $Y=1.665
+ $X2=11.195 $Y2=1.375
r258 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=1.665
+ $X2=11.28 $Y2=1.665
r259 43 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=1.665
+ $X2=7.92 $Y2=1.665
r260 41 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.065 $Y=1.665
+ $X2=7.92 $Y2=1.665
r261 40 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=11.135 $Y=1.665
+ $X2=11.28 $Y2=1.665
r262 40 41 3.7995 $w=1.4e-07 $l=3.07e-06 $layer=MET1_cond $X=11.135 $Y=1.665
+ $X2=8.065 $Y2=1.665
r263 39 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.745 $Y=1.665
+ $X2=3.6 $Y2=1.665
r264 38 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.775 $Y=1.665
+ $X2=7.92 $Y2=1.665
r265 38 39 4.98761 $w=1.4e-07 $l=4.03e-06 $layer=MET1_cond $X=7.775 $Y=1.665
+ $X2=3.745 $Y2=1.665
r266 36 37 19.6163 $w=1.72e-07 $l=7e-08 $layer=POLY_cond $X=11.25 $Y=2.375
+ $X2=11.32 $Y2=2.375
r267 32 34 104.279 $w=1.6e-07 $l=2.25e-07 $layer=POLY_cond $X=7.535 $Y=2.16
+ $X2=7.76 $Y2=2.16
r268 29 37 6.07713 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=11.32 $Y=2.465
+ $X2=11.32 $Y2=2.375
r269 29 31 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=11.32 $Y=2.465
+ $X2=11.32 $Y2=2.75
r270 28 36 6.07713 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=11.25 $Y=2.285
+ $X2=11.25 $Y2=2.375
r271 28 64 382.011 $w=1.5e-07 $l=7.45e-07 $layer=POLY_cond $X=11.25 $Y=2.285
+ $X2=11.25 $Y2=1.54
r272 25 63 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=11.25 $Y=0.58
+ $X2=11.25 $Y2=1.21
r273 22 34 4.37345 $w=1.5e-07 $l=8e-08 $layer=POLY_cond $X=7.76 $Y=2.08 $X2=7.76
+ $Y2=2.16
r274 22 59 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=7.76 $Y=2.08
+ $X2=7.76 $Y2=1.8
r275 19 58 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=7.76 $Y=0.825
+ $X2=7.76 $Y2=1.47
r276 14 16 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=7.535 $Y=3.075
+ $X2=7.535 $Y2=2.525
r277 13 32 4.37345 $w=1.5e-07 $l=8e-08 $layer=POLY_cond $X=7.535 $Y=2.24
+ $X2=7.535 $Y2=2.16
r278 13 16 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.535 $Y=2.24
+ $X2=7.535 $Y2=2.525
r279 11 52 2.68759 $w=3.65e-07 $l=1.7e-08 $layer=POLY_cond $X=3.552 $Y=1.537
+ $X2=3.552 $Y2=1.52
r280 11 12 48.3767 $w=3.65e-07 $l=3.06e-07 $layer=POLY_cond $X=3.552 $Y=1.537
+ $X2=3.552 $Y2=1.843
r281 9 54 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=3.445 $Y=0.615
+ $X2=3.445 $Y2=1.355
r282 5 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.46 $Y=3.15
+ $X2=7.535 $Y2=3.075
r283 5 6 2099.78 $w=1.5e-07 $l=4.095e-06 $layer=POLY_cond $X=7.46 $Y=3.15
+ $X2=3.365 $Y2=3.15
r284 2 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.29 $Y=3.075
+ $X2=3.365 $Y2=3.15
r285 2 4 223.053 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.29 $Y=3.075
+ $X2=3.29 $Y2=2.64
r286 1 12 62.5045 $w=3.1e-07 $l=5.16651e-07 $layer=POLY_cond $X=3.29 $Y=2.245
+ $X2=3.552 $Y2=1.843
r287 1 4 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.29 $Y=2.245
+ $X2=3.29 $Y2=2.64
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTN_1%A_1251_463# 1 2 3 10 12 13 15 18 20 21 23
+ 24 28 30 34 35 40 42 45
c128 40 0 1.76356e-19 $X=6.97 $Y=0.91
c129 34 0 7.49297e-20 $X=8.39 $Y=1.635
c130 23 0 1.7914e-19 $X=6.97 $Y=2.04
r131 38 40 6.69663 $w=3.68e-07 $l=2.15e-07 $layer=LI1_cond $X=6.755 $Y=0.91
+ $X2=6.97 $Y2=0.91
r132 35 48 39.8291 $w=3.57e-07 $l=2.95e-07 $layer=POLY_cond $X=8.39 $Y=1.677
+ $X2=8.685 $Y2=1.677
r133 35 46 5.40056 $w=3.57e-07 $l=4e-08 $layer=POLY_cond $X=8.39 $Y=1.677
+ $X2=8.35 $Y2=1.677
r134 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.39
+ $Y=1.635 $X2=8.39 $Y2=1.635
r135 32 34 13.0871 $w=2.93e-07 $l=3.35e-07 $layer=LI1_cond $X=8.372 $Y=1.97
+ $X2=8.372 $Y2=1.635
r136 31 45 9.39981 $w=1.7e-07 $l=3.82426e-07 $layer=LI1_cond $X=7.95 $Y=2.055
+ $X2=7.575 $Y2=2.04
r137 30 32 7.47753 $w=1.7e-07 $l=1.84673e-07 $layer=LI1_cond $X=8.225 $Y=2.055
+ $X2=8.372 $Y2=1.97
r138 30 31 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=8.225 $Y=2.055
+ $X2=7.95 $Y2=2.055
r139 26 45 1.28102 $w=3.75e-07 $l=2.58378e-07 $layer=LI1_cond $X=7.762 $Y=2.21
+ $X2=7.575 $Y2=2.04
r140 26 28 10.2952 $w=3.73e-07 $l=3.35e-07 $layer=LI1_cond $X=7.762 $Y=2.21
+ $X2=7.762 $Y2=2.545
r141 25 42 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.055 $Y=2.125
+ $X2=6.97 $Y2=2.125
r142 24 45 9.39981 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.575 $Y=2.125
+ $X2=7.575 $Y2=2.04
r143 24 25 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=7.575 $Y=2.125
+ $X2=7.055 $Y2=2.125
r144 23 42 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=6.97 $Y=2.04
+ $X2=6.97 $Y2=2.125
r145 22 40 5.30706 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=6.97 $Y=1.095
+ $X2=6.97 $Y2=0.91
r146 22 23 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=6.97 $Y=1.095
+ $X2=6.97 $Y2=2.04
r147 20 42 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=6.97 $Y=2.34
+ $X2=6.97 $Y2=2.125
r148 20 21 16.6364 $w=2.08e-07 $l=3.15e-07 $layer=LI1_cond $X=6.885 $Y=2.34
+ $X2=6.57 $Y2=2.34
r149 16 21 7.02201 $w=2.1e-07 $l=1.88319e-07 $layer=LI1_cond $X=6.427 $Y=2.445
+ $X2=6.57 $Y2=2.34
r150 16 18 4.04366 $w=2.83e-07 $l=1e-07 $layer=LI1_cond $X=6.427 $Y=2.445
+ $X2=6.427 $Y2=2.545
r151 13 48 23.1043 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=8.685 $Y=1.885
+ $X2=8.685 $Y2=1.677
r152 13 15 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=8.685 $Y=1.885
+ $X2=8.685 $Y2=2.46
r153 10 46 23.1043 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=8.35 $Y=1.47
+ $X2=8.35 $Y2=1.677
r154 10 12 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=8.35 $Y=1.47
+ $X2=8.35 $Y2=1.04
r155 3 28 600 $w=1.7e-07 $l=2.95635e-07 $layer=licon1_PDIFF $count=1 $X=7.61
+ $Y=2.315 $X2=7.76 $Y2=2.545
r156 2 18 600 $w=1.7e-07 $l=2.95635e-07 $layer=licon1_PDIFF $count=1 $X=6.255
+ $Y=2.315 $X2=6.405 $Y2=2.545
r157 1 38 182 $w=1.7e-07 $l=5.14441e-07 $layer=licon1_NDIFF $count=1 $X=6.36
+ $Y=0.615 $X2=6.755 $Y2=0.89
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTN_1%A_854_74# 1 2 7 9 11 13 14 18 20 22 27 28
+ 29 33 35 36 38 39 40 44 48 53 59 61 63 65 68 70 71 72
c207 35 0 1.69146e-19 $X=10.135 $Y=2.375
c208 22 0 1.61279e-19 $X=6.905 $Y=1.225
c209 11 0 6.18507e-21 $X=5.295 $Y=1.245
r210 71 80 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=10.23 $Y=1.39
+ $X2=10.135 $Y2=1.39
r211 70 72 8.46257 $w=3.13e-07 $l=1.65e-07 $layer=LI1_cond $X=10.23 $Y=1.382
+ $X2=10.065 $Y2=1.382
r212 70 71 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.23
+ $Y=1.39 $X2=10.23 $Y2=1.39
r213 68 76 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=9.155 $Y=1.635
+ $X2=9.06 $Y2=1.635
r214 67 68 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.155
+ $Y=1.635 $X2=9.155 $Y2=1.635
r215 65 67 7.70526 $w=2.85e-07 $l=1.8e-07 $layer=LI1_cond $X=9.19 $Y=1.455
+ $X2=9.19 $Y2=1.635
r216 62 75 5.37047 $w=3.59e-07 $l=4e-08 $layer=POLY_cond $X=5.187 $Y=1.41
+ $X2=5.187 $Y2=1.45
r217 61 64 8.99425 $w=4.08e-07 $l=1.95e-07 $layer=LI1_cond $X=5.05 $Y=1.41
+ $X2=5.05 $Y2=1.605
r218 61 63 5.5054 $w=4.08e-07 $l=1.75e-07 $layer=LI1_cond $X=5.05 $Y=1.41
+ $X2=5.05 $Y2=1.235
r219 61 62 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.17
+ $Y=1.41 $X2=5.17 $Y2=1.41
r220 57 59 6.51648 $w=1.78e-07 $l=1.05e-07 $layer=LI1_cond $X=4.495 $Y=1.91
+ $X2=4.6 $Y2=1.91
r221 55 65 3.76007 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=9.35 $Y=1.455
+ $X2=9.19 $Y2=1.455
r222 55 72 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=9.35 $Y=1.455
+ $X2=10.065 $Y2=1.455
r223 53 64 12.8894 $w=1.83e-07 $l=2.15e-07 $layer=LI1_cond $X=4.937 $Y=1.82
+ $X2=4.937 $Y2=1.605
r224 50 63 7.0227 $w=3.18e-07 $l=1.95e-07 $layer=LI1_cond $X=5.005 $Y=1.04
+ $X2=5.005 $Y2=1.235
r225 48 53 6.83233 $w=1.7e-07 $l=1.27609e-07 $layer=LI1_cond $X=4.845 $Y=1.905
+ $X2=4.937 $Y2=1.82
r226 48 59 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=4.845 $Y=1.905
+ $X2=4.6 $Y2=1.905
r227 44 50 7.68211 $w=1.7e-07 $l=1.9799e-07 $layer=LI1_cond $X=4.845 $Y=0.955
+ $X2=5.005 $Y2=1.04
r228 44 46 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=4.845 $Y=0.955
+ $X2=4.41 $Y2=0.955
r229 40 42 115.372 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=6.675 $Y=1.225
+ $X2=6.675 $Y2=1.45
r230 36 38 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=10.135 $Y=2.465
+ $X2=10.135 $Y2=2.75
r231 35 36 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=10.135 $Y=2.375
+ $X2=10.135 $Y2=2.465
r232 34 80 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=10.135 $Y=1.555
+ $X2=10.135 $Y2=1.39
r233 34 35 318.742 $w=1.8e-07 $l=8.2e-07 $layer=POLY_cond $X=10.135 $Y=1.555
+ $X2=10.135 $Y2=2.375
r234 31 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.06 $Y=1.47
+ $X2=9.06 $Y2=1.635
r235 31 33 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=9.06 $Y=1.47
+ $X2=9.06 $Y2=1.04
r236 30 33 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=9.06 $Y=0.275
+ $X2=9.06 $Y2=1.04
r237 28 30 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.985 $Y=0.2
+ $X2=9.06 $Y2=0.275
r238 28 29 989.638 $w=1.5e-07 $l=1.93e-06 $layer=POLY_cond $X=8.985 $Y=0.2
+ $X2=7.055 $Y2=0.2
r239 25 27 166.649 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=6.98 $Y=1.15
+ $X2=6.98 $Y2=0.825
r240 24 29 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.98 $Y=0.275
+ $X2=7.055 $Y2=0.2
r241 24 27 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=6.98 $Y=0.275
+ $X2=6.98 $Y2=0.825
r242 23 40 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.75 $Y=1.225
+ $X2=6.675 $Y2=1.225
r243 22 25 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.905 $Y=1.225
+ $X2=6.98 $Y2=1.15
r244 22 23 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=6.905 $Y=1.225
+ $X2=6.75 $Y2=1.225
r245 21 39 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.255 $Y=1.45
+ $X2=6.18 $Y2=1.45
r246 20 42 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.6 $Y=1.45
+ $X2=6.675 $Y2=1.45
r247 20 21 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=6.6 $Y=1.45
+ $X2=6.255 $Y2=1.45
r248 16 39 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.18 $Y=1.525
+ $X2=6.18 $Y2=1.45
r249 16 18 512.766 $w=1.5e-07 $l=1e-06 $layer=POLY_cond $X=6.18 $Y=1.525
+ $X2=6.18 $Y2=2.525
r250 15 75 23.2387 $w=1.5e-07 $l=1.83e-07 $layer=POLY_cond $X=5.37 $Y=1.45
+ $X2=5.187 $Y2=1.45
r251 14 39 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.105 $Y=1.45
+ $X2=6.18 $Y2=1.45
r252 14 15 376.883 $w=1.5e-07 $l=7.35e-07 $layer=POLY_cond $X=6.105 $Y=1.45
+ $X2=5.37 $Y2=1.45
r253 11 62 38.8967 $w=3.59e-07 $l=2.12238e-07 $layer=POLY_cond $X=5.295 $Y=1.245
+ $X2=5.187 $Y2=1.41
r254 11 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.295 $Y=1.245
+ $X2=5.295 $Y2=0.765
r255 7 75 33.5262 $w=3.59e-07 $l=1.33229e-07 $layer=POLY_cond $X=5.17 $Y=1.575
+ $X2=5.187 $Y2=1.45
r256 7 9 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.17 $Y=1.575
+ $X2=5.17 $Y2=2.235
r257 2 57 600 $w=1.7e-07 $l=2.56271e-07 $layer=licon1_PDIFF $count=1 $X=4.31
+ $Y=1.735 $X2=4.495 $Y2=1.905
r258 1 46 182 $w=1.7e-07 $l=6.51249e-07 $layer=licon1_NDIFF $count=1 $X=4.27
+ $Y=0.37 $X2=4.41 $Y2=0.955
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTN_1%A_2087_410# 1 2 7 9 12 14 18 20 24 27 29 34
c91 29 0 9.65573e-20 $X=10.6 $Y=2.215
c92 12 0 1.91401e-20 $X=10.69 $Y=0.58
r93 29 32 7.37564 $w=2.48e-07 $l=1.6e-07 $layer=LI1_cond $X=10.56 $Y=2.215
+ $X2=10.56 $Y2=2.375
r94 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.6
+ $Y=2.215 $X2=10.6 $Y2=2.215
r95 26 27 103.733 $w=1.68e-07 $l=1.59e-06 $layer=LI1_cond $X=12.15 $Y=0.7
+ $X2=12.15 $Y2=2.29
r96 25 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.71 $Y=2.375
+ $X2=11.545 $Y2=2.375
r97 24 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=12.065 $Y=2.375
+ $X2=12.15 $Y2=2.29
r98 24 25 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=12.065 $Y=2.375
+ $X2=11.71 $Y2=2.375
r99 20 26 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=12.065 $Y=0.575
+ $X2=12.15 $Y2=0.7
r100 20 22 4.84026 $w=2.48e-07 $l=1.05e-07 $layer=LI1_cond $X=12.065 $Y=0.575
+ $X2=11.96 $Y2=0.575
r101 16 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.545 $Y=2.46
+ $X2=11.545 $Y2=2.375
r102 16 18 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=11.545 $Y=2.46
+ $X2=11.545 $Y2=2.75
r103 15 32 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.685 $Y=2.375
+ $X2=10.56 $Y2=2.375
r104 14 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.38 $Y=2.375
+ $X2=11.545 $Y2=2.375
r105 14 15 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=11.38 $Y=2.375
+ $X2=10.685 $Y2=2.375
r106 10 30 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=10.69 $Y=2.05
+ $X2=10.6 $Y2=2.215
r107 10 12 753.766 $w=1.5e-07 $l=1.47e-06 $layer=POLY_cond $X=10.69 $Y=2.05
+ $X2=10.69 $Y2=0.58
r108 7 30 52.2586 $w=2.99e-07 $l=2.76134e-07 $layer=POLY_cond $X=10.545 $Y=2.465
+ $X2=10.6 $Y2=2.215
r109 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=10.545 $Y=2.465
+ $X2=10.545 $Y2=2.75
r110 2 18 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=11.395
+ $Y=2.54 $X2=11.545 $Y2=2.75
r111 1 22 182 $w=1.7e-07 $l=3.46482e-07 $layer=licon1_NDIFF $count=1 $X=11.715
+ $Y=0.37 $X2=11.96 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTN_1%A_1827_144# 1 2 7 9 11 13 15 16 18 19 21 23
+ 25 26 28 29 30 35 39 40 41 42 43 44 45 50 51 53 54
c159 54 0 1.97052e-19 $X=10.94 $Y=1.795
c160 40 0 1.91401e-20 $X=10.08 $Y=0.87
c161 21 0 1.07922e-19 $X=12.77 $Y=1.07
c162 19 0 1.07922e-19 $X=12.755 $Y=1.97
r163 54 56 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=10.94 $Y=1.795
+ $X2=10.94 $Y2=2.035
r164 50 51 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=11.73
+ $Y=1.065 $X2=11.73 $Y2=1.065
r165 48 50 30.9064 $w=3.28e-07 $l=8.85e-07 $layer=LI1_cond $X=11.73 $Y=1.95
+ $X2=11.73 $Y2=1.065
r166 47 50 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=11.73 $Y=1.04
+ $X2=11.73 $Y2=1.065
r167 46 56 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.025 $Y=2.035
+ $X2=10.94 $Y2=2.035
r168 45 48 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=11.565 $Y=2.035
+ $X2=11.73 $Y2=1.95
r169 45 46 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=11.565 $Y=2.035
+ $X2=11.025 $Y2=2.035
r170 43 47 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=11.565 $Y=0.955
+ $X2=11.73 $Y2=1.04
r171 43 44 91.3369 $w=1.68e-07 $l=1.4e-06 $layer=LI1_cond $X=11.565 $Y=0.955
+ $X2=10.165 $Y2=0.955
r172 41 54 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.855 $Y=1.795
+ $X2=10.94 $Y2=1.795
r173 41 42 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=10.855 $Y=1.795
+ $X2=10.065 $Y2=1.795
r174 40 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.08 $Y=0.87
+ $X2=10.165 $Y2=0.955
r175 39 53 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.08 $Y=0.62
+ $X2=10.08 $Y2=0.455
r176 39 40 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=10.08 $Y=0.62
+ $X2=10.08 $Y2=0.87
r177 35 37 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=9.9 $Y=2.135
+ $X2=9.9 $Y2=2.815
r178 33 42 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.9 $Y=1.88
+ $X2=10.065 $Y2=1.795
r179 33 35 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=9.9 $Y=1.88
+ $X2=9.9 $Y2=2.135
r180 26 28 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=12.845 $Y=0.995
+ $X2=12.845 $Y2=0.645
r181 23 25 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=12.83 $Y=2.045
+ $X2=12.83 $Y2=2.54
r182 22 51 12.1617 $w=1.5e-07 $l=1.8747e-07 $layer=POLY_cond $X=11.895 $Y=1.07
+ $X2=11.73 $Y2=1.022
r183 21 26 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=12.77 $Y=1.07
+ $X2=12.845 $Y2=0.995
r184 21 22 448.67 $w=1.5e-07 $l=8.75e-07 $layer=POLY_cond $X=12.77 $Y=1.07
+ $X2=11.895 $Y2=1.07
r185 20 30 6.66866 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=11.86 $Y=1.97
+ $X2=11.77 $Y2=1.97
r186 19 23 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=12.755 $Y=1.97
+ $X2=12.83 $Y2=2.045
r187 19 20 458.926 $w=1.5e-07 $l=8.95e-07 $layer=POLY_cond $X=12.755 $Y=1.97
+ $X2=11.86 $Y2=1.97
r188 16 18 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=11.77 $Y=2.465
+ $X2=11.77 $Y2=2.75
r189 15 16 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=11.77 $Y=2.375
+ $X2=11.77 $Y2=2.465
r190 14 30 18.8402 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=11.77 $Y=2.045
+ $X2=11.77 $Y2=1.97
r191 14 15 128.274 $w=1.8e-07 $l=3.3e-07 $layer=POLY_cond $X=11.77 $Y=2.045
+ $X2=11.77 $Y2=2.375
r192 13 30 18.8402 $w=1.65e-07 $l=8.21584e-08 $layer=POLY_cond $X=11.755
+ $Y=1.895 $X2=11.77 $Y2=1.97
r193 13 29 166.649 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=11.755 $Y=1.895
+ $X2=11.755 $Y2=1.57
r194 11 29 38.9318 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=11.73 $Y=1.405
+ $X2=11.73 $Y2=1.57
r195 10 51 13.5877 $w=2.4e-07 $l=1.23e-07 $layer=POLY_cond $X=11.73 $Y=1.145
+ $X2=11.73 $Y2=1.022
r196 10 11 45.4639 $w=3.3e-07 $l=2.6e-07 $layer=POLY_cond $X=11.73 $Y=1.145
+ $X2=11.73 $Y2=1.405
r197 7 51 13.5877 $w=2.4e-07 $l=1.60823e-07 $layer=POLY_cond $X=11.64 $Y=0.9
+ $X2=11.73 $Y2=1.022
r198 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=11.64 $Y=0.9
+ $X2=11.64 $Y2=0.58
r199 2 37 600 $w=1.7e-07 $l=9.51998e-07 $layer=licon1_PDIFF $count=1 $X=9.695
+ $Y=1.96 $X2=9.9 $Y2=2.815
r200 2 35 300 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=2 $X=9.695
+ $Y=1.96 $X2=9.845 $Y2=2.135
r201 1 53 91 $w=1.7e-07 $l=9.83616e-07 $layer=licon1_NDIFF $count=2 $X=9.135
+ $Y=0.72 $X2=9.995 $Y2=0.455
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTN_1%A_2492_424# 1 2 7 9 12 14 15 18 22 25
c45 25 0 2.15844e-19 $X=12.645 $Y=1.52
r46 25 28 5.13927 $w=3.68e-07 $l=1.65e-07 $layer=LI1_cond $X=12.625 $Y=1.52
+ $X2=12.625 $Y2=1.685
r47 25 27 5.13927 $w=3.68e-07 $l=1.65e-07 $layer=LI1_cond $X=12.625 $Y=1.52
+ $X2=12.625 $Y2=1.355
r48 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.645
+ $Y=1.52 $X2=12.645 $Y2=1.52
r49 22 28 18.8286 $w=3.53e-07 $l=5.8e-07 $layer=LI1_cond $X=12.617 $Y=2.265
+ $X2=12.617 $Y2=1.685
r50 18 27 23.0489 $w=3.53e-07 $l=7.1e-07 $layer=LI1_cond $X=12.617 $Y=0.645
+ $X2=12.617 $Y2=1.355
r51 14 26 118.031 $w=3.3e-07 $l=6.75e-07 $layer=POLY_cond $X=13.32 $Y=1.52
+ $X2=12.645 $Y2=1.52
r52 14 15 5.03009 $w=3.3e-07 $l=1.08167e-07 $layer=POLY_cond $X=13.32 $Y=1.52
+ $X2=13.41 $Y2=1.56
r53 10 15 37.0704 $w=1.5e-07 $l=2.12368e-07 $layer=POLY_cond $X=13.425 $Y=1.355
+ $X2=13.41 $Y2=1.56
r54 10 12 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=13.425 $Y=1.355
+ $X2=13.425 $Y2=0.74
r55 7 15 37.0704 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=13.41 $Y=1.765
+ $X2=13.41 $Y2=1.56
r56 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=13.41 $Y=1.765
+ $X2=13.41 $Y2=2.4
r57 2 22 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=12.46
+ $Y=2.12 $X2=12.605 $Y2=2.265
r58 1 18 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=12.485
+ $Y=0.37 $X2=12.63 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTN_1%VPWR 1 2 3 4 5 6 7 8 27 31 35 39 43 47 52
+ 53 55 56 57 59 64 72 81 85 97 103 104 107 110 117 120 123 130
c139 123 0 1.81488e-19 $X=10.905 $Y=2.815
c140 5 0 7.49297e-20 $X=8.325 $Y=1.96
r141 130 131 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=3.33
+ $X2=13.2 $Y2=3.33
r142 120 121 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r143 117 118 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r144 113 114 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r145 110 113 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.98 $Y=3.055
+ $X2=2.98 $Y2=3.33
r146 107 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r147 104 131 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=3.33
+ $X2=13.2 $Y2=3.33
r148 103 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=3.33
+ $X2=13.68 $Y2=3.33
r149 101 130 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.305 $Y=3.33
+ $X2=13.14 $Y2=3.33
r150 101 103 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=13.305 $Y=3.33
+ $X2=13.68 $Y2=3.33
r151 100 131 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=13.2 $Y2=3.33
r152 99 100 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r153 97 130 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.975 $Y=3.33
+ $X2=13.14 $Y2=3.33
r154 97 99 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=12.975 $Y=3.33
+ $X2=12.72 $Y2=3.33
r155 96 100 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=12.72 $Y2=3.33
r156 96 127 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=10.8 $Y2=3.33
r157 95 96 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r158 93 95 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=11.21 $Y=3.33
+ $X2=11.76 $Y2=3.33
r159 92 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=10.8 $Y2=3.33
r160 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r161 89 92 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=10.32 $Y2=3.33
r162 89 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=8.4 $Y2=3.33
r163 88 91 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=8.88 $Y=3.33
+ $X2=10.32 $Y2=3.33
r164 88 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r165 86 120 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.625 $Y=3.33
+ $X2=8.46 $Y2=3.33
r166 86 88 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=8.625 $Y=3.33
+ $X2=8.88 $Y2=3.33
r167 85 93 8.37032 $w=1.7e-07 $l=3.03e-07 $layer=LI1_cond $X=10.907 $Y=3.33
+ $X2=11.21 $Y2=3.33
r168 85 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r169 85 123 10.1815 $w=6.03e-07 $l=5.15e-07 $layer=LI1_cond $X=10.907 $Y=3.33
+ $X2=10.907 $Y2=2.815
r170 85 91 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=10.605 $Y=3.33
+ $X2=10.32 $Y2=3.33
r171 84 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r172 83 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r173 81 120 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.295 $Y=3.33
+ $X2=8.46 $Y2=3.33
r174 81 83 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=8.295 $Y=3.33
+ $X2=7.92 $Y2=3.33
r175 77 117 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.11 $Y=3.33
+ $X2=4.945 $Y2=3.33
r176 77 79 120.695 $w=1.68e-07 $l=1.85e-06 $layer=LI1_cond $X=5.11 $Y=3.33
+ $X2=6.96 $Y2=3.33
r177 76 118 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r178 76 114 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=3.12 $Y2=3.33
r179 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r180 73 113 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.145 $Y=3.33
+ $X2=2.98 $Y2=3.33
r181 73 75 92.3155 $w=1.68e-07 $l=1.415e-06 $layer=LI1_cond $X=3.145 $Y=3.33
+ $X2=4.56 $Y2=3.33
r182 72 117 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.78 $Y=3.33
+ $X2=4.945 $Y2=3.33
r183 72 75 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=4.78 $Y=3.33
+ $X2=4.56 $Y2=3.33
r184 71 114 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r185 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r186 68 71 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r187 68 108 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r188 67 70 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r189 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r190 65 107 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=0.73 $Y2=3.33
r191 65 67 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=1.2 $Y2=3.33
r192 64 113 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.815 $Y=3.33
+ $X2=2.98 $Y2=3.33
r193 64 70 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.815 $Y=3.33
+ $X2=2.64 $Y2=3.33
r194 62 108 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r195 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r196 59 107 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.73 $Y2=3.33
r197 59 61 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.24 $Y2=3.33
r198 57 84 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.92 $Y2=3.33
r199 57 118 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=5.04 $Y2=3.33
r200 57 79 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r201 55 95 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=11.88 $Y=3.33
+ $X2=11.76 $Y2=3.33
r202 55 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.88 $Y=3.33
+ $X2=12.045 $Y2=3.33
r203 54 99 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=12.21 $Y=3.33
+ $X2=12.72 $Y2=3.33
r204 54 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.21 $Y=3.33
+ $X2=12.045 $Y2=3.33
r205 52 79 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=7.225 $Y=3.33
+ $X2=6.96 $Y2=3.33
r206 52 53 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.225 $Y=3.33
+ $X2=7.31 $Y2=3.33
r207 51 83 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=7.395 $Y=3.33
+ $X2=7.92 $Y2=3.33
r208 51 53 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.395 $Y=3.33
+ $X2=7.31 $Y2=3.33
r209 47 50 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=13.14 $Y=1.985
+ $X2=13.14 $Y2=2.4
r210 45 130 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.14 $Y=3.245
+ $X2=13.14 $Y2=3.33
r211 45 50 29.5095 $w=3.28e-07 $l=8.45e-07 $layer=LI1_cond $X=13.14 $Y=3.245
+ $X2=13.14 $Y2=2.4
r212 41 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.045 $Y=3.245
+ $X2=12.045 $Y2=3.33
r213 41 43 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=12.045 $Y=3.245
+ $X2=12.045 $Y2=2.805
r214 37 120 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.46 $Y=3.245
+ $X2=8.46 $Y2=3.33
r215 37 39 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=8.46 $Y=3.245
+ $X2=8.46 $Y2=2.475
r216 33 53 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.31 $Y=3.245
+ $X2=7.31 $Y2=3.33
r217 33 35 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=7.31 $Y=3.245
+ $X2=7.31 $Y2=2.545
r218 29 117 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.945 $Y=3.245
+ $X2=4.945 $Y2=3.33
r219 29 31 23.0489 $w=3.28e-07 $l=6.6e-07 $layer=LI1_cond $X=4.945 $Y=3.245
+ $X2=4.945 $Y2=2.585
r220 25 107 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=3.33
r221 25 27 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=2.805
r222 8 50 300 $w=1.7e-07 $l=3.79737e-07 $layer=licon1_PDIFF $count=2 $X=12.905
+ $Y=2.12 $X2=13.14 $Y2=2.4
r223 8 47 600 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_PDIFF $count=1 $X=12.905
+ $Y=2.12 $X2=13.14 $Y2=1.985
r224 7 43 600 $w=1.7e-07 $l=3.51034e-07 $layer=licon1_PDIFF $count=1 $X=11.845
+ $Y=2.54 $X2=12.045 $Y2=2.805
r225 6 123 600 $w=1.7e-07 $l=3.995e-07 $layer=licon1_PDIFF $count=1 $X=10.62
+ $Y=2.54 $X2=10.905 $Y2=2.815
r226 5 39 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=8.325
+ $Y=1.96 $X2=8.46 $Y2=2.475
r227 4 35 600 $w=1.7e-07 $l=2.95635e-07 $layer=licon1_PDIFF $count=1 $X=7.16
+ $Y=2.315 $X2=7.31 $Y2=2.545
r228 3 31 600 $w=1.7e-07 $l=9.21954e-07 $layer=licon1_PDIFF $count=1 $X=4.795
+ $Y=1.735 $X2=4.945 $Y2=2.585
r229 2 110 600 $w=1.7e-07 $l=8.44364e-07 $layer=licon1_PDIFF $count=1 $X=2.745
+ $Y=2.32 $X2=2.98 $Y2=3.055
r230 1 27 600 $w=1.7e-07 $l=5.54955e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=2.32 $X2=0.73 $Y2=2.805
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTN_1%A_284_464# 1 2 3 4 5 18 22 25 26 27 29 31
+ 32 33 35 37 38 39 40 42 46 50 53 54 57 58
c158 46 0 1.13453e-19 $X=5.955 $Y=2.545
r159 53 54 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.055 $Y=2.795
+ $X2=2.22 $Y2=2.795
r160 48 50 7.60612 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=6.03 $Y=0.7
+ $X2=6.03 $Y2=0.865
r161 44 46 9.52982 $w=2.58e-07 $l=2.15e-07 $layer=LI1_cond $X=5.985 $Y=2.33
+ $X2=5.985 $Y2=2.545
r162 42 44 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=5.855 $Y=2.245
+ $X2=5.985 $Y2=2.33
r163 42 43 74.0481 $w=1.68e-07 $l=1.135e-06 $layer=LI1_cond $X=5.855 $Y=2.245
+ $X2=4.72 $Y2=2.245
r164 41 58 4.27425 $w=2.12e-07 $l=8.5e-08 $layer=LI1_cond $X=4.075 $Y=2.282
+ $X2=3.99 $Y2=2.282
r165 40 43 10.9158 $w=2.09e-07 $l=2.04666e-07 $layer=LI1_cond $X=4.533 $Y=2.282
+ $X2=4.72 $Y2=2.245
r166 40 41 23.4586 $w=2.23e-07 $l=4.58e-07 $layer=LI1_cond $X=4.533 $Y=2.282
+ $X2=4.075 $Y2=2.282
r167 38 48 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.905 $Y=0.615
+ $X2=6.03 $Y2=0.7
r168 38 39 119.39 $w=1.68e-07 $l=1.83e-06 $layer=LI1_cond $X=5.905 $Y=0.615
+ $X2=4.075 $Y2=0.615
r169 37 58 2.15711 $w=1.7e-07 $l=1.12e-07 $layer=LI1_cond $X=3.99 $Y=2.17
+ $X2=3.99 $Y2=2.282
r170 36 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.99 $Y=1.185
+ $X2=3.99 $Y2=1.1
r171 36 37 64.262 $w=1.68e-07 $l=9.85e-07 $layer=LI1_cond $X=3.99 $Y=1.185
+ $X2=3.99 $Y2=2.17
r172 35 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.99 $Y=1.015
+ $X2=3.99 $Y2=1.1
r173 34 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.99 $Y=0.7
+ $X2=4.075 $Y2=0.615
r174 34 35 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=3.99 $Y=0.7
+ $X2=3.99 $Y2=1.015
r175 32 58 4.27425 $w=2.12e-07 $l=9.12688e-08 $layer=LI1_cond $X=3.905 $Y=2.295
+ $X2=3.99 $Y2=2.282
r176 32 33 12.4773 $w=1.98e-07 $l=2.25e-07 $layer=LI1_cond $X=3.905 $Y=2.295
+ $X2=3.68 $Y2=2.295
r177 29 56 3.20527 $w=2.5e-07 $l=1.75e-07 $layer=LI1_cond $X=3.555 $Y=2.63
+ $X2=3.555 $Y2=2.805
r178 29 31 7.60612 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=3.555 $Y=2.63
+ $X2=3.555 $Y2=2.465
r179 28 33 6.92652 $w=2e-07 $l=1.67705e-07 $layer=LI1_cond $X=3.555 $Y=2.395
+ $X2=3.68 $Y2=2.295
r180 28 31 3.22684 $w=2.48e-07 $l=7e-08 $layer=LI1_cond $X=3.555 $Y=2.395
+ $X2=3.555 $Y2=2.465
r181 26 57 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.905 $Y=1.1
+ $X2=3.99 $Y2=1.1
r182 26 27 66.2193 $w=1.68e-07 $l=1.015e-06 $layer=LI1_cond $X=3.905 $Y=1.1
+ $X2=2.89 $Y2=1.1
r183 25 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.805 $Y=1.015
+ $X2=2.89 $Y2=1.1
r184 24 25 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.805 $Y=0.765
+ $X2=2.805 $Y2=1.015
r185 22 56 3.9379 $w=1.7e-07 $l=1.63936e-07 $layer=LI1_cond $X=3.43 $Y=2.715
+ $X2=3.555 $Y2=2.805
r186 22 54 78.9412 $w=1.68e-07 $l=1.21e-06 $layer=LI1_cond $X=3.43 $Y=2.715
+ $X2=2.22 $Y2=2.715
r187 18 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.72 $Y=0.68
+ $X2=2.805 $Y2=0.765
r188 18 20 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=2.72 $Y=0.68
+ $X2=2.26 $Y2=0.68
r189 5 46 600 $w=1.7e-07 $l=2.93684e-07 $layer=licon1_PDIFF $count=1 $X=5.81
+ $Y=2.315 $X2=5.955 $Y2=2.545
r190 4 56 600 $w=1.7e-07 $l=5.65044e-07 $layer=licon1_PDIFF $count=1 $X=3.365
+ $Y=2.32 $X2=3.515 $Y2=2.815
r191 4 31 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=3.365
+ $Y=2.32 $X2=3.515 $Y2=2.465
r192 3 53 300 $w=1.7e-07 $l=8.39553e-07 $layer=licon1_PDIFF $count=2 $X=1.42
+ $Y=2.32 $X2=2.055 $Y2=2.795
r193 2 50 182 $w=1.7e-07 $l=3.14245e-07 $layer=licon1_NDIFF $count=1 $X=5.925
+ $Y=0.615 $X2=6.07 $Y2=0.865
r194 1 20 182 $w=1.7e-07 $l=3.94208e-07 $layer=licon1_NDIFF $count=1 $X=1.98
+ $Y=0.405 $X2=2.26 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTN_1%Q 1 2 7 8 9 10 11 12 13
r13 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=13.64 $Y=2.405
+ $X2=13.64 $Y2=2.775
r14 11 12 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=13.64 $Y=1.985
+ $X2=13.64 $Y2=2.405
r15 10 11 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=13.64 $Y=1.665
+ $X2=13.64 $Y2=1.985
r16 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=13.64 $Y=1.295
+ $X2=13.64 $Y2=1.665
r17 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=13.64 $Y=0.925
+ $X2=13.64 $Y2=1.295
r18 7 8 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=13.64 $Y=0.515
+ $X2=13.64 $Y2=0.925
r19 2 13 400 $w=1.7e-07 $l=1.04964e-06 $layer=licon1_PDIFF $count=1 $X=13.485
+ $Y=1.84 $X2=13.64 $Y2=2.815
r20 2 11 400 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=1 $X=13.485
+ $Y=1.84 $X2=13.64 $Y2=1.985
r21 1 7 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=13.5
+ $Y=0.37 $X2=13.64 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTN_1%VGND 1 2 3 4 5 6 21 25 29 33 37 39 49 54 59
+ 64 74 75 78 83 86 89 95 98 101
r117 101 102 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=0
+ $X2=13.2 $Y2=0
r118 98 99 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=10.8 $Y=0 $X2=10.8
+ $Y2=0
r119 95 96 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r120 89 92 8.80338 $w=3.58e-07 $l=2.75e-07 $layer=LI1_cond $X=4.985 $Y=0
+ $X2=4.985 $Y2=0.275
r121 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r122 85 86 10.9331 $w=4.43e-07 $l=2.45e-07 $layer=LI1_cond $X=3.82 $Y=0.137
+ $X2=4.065 $Y2=0.137
r123 81 85 5.69747 $w=4.43e-07 $l=2.2e-07 $layer=LI1_cond $X=3.6 $Y=0.137
+ $X2=3.82 $Y2=0.137
r124 81 83 5.23558 $w=4.43e-07 $l=2.5e-08 $layer=LI1_cond $X=3.6 $Y=0.137
+ $X2=3.575 $Y2=0.137
r125 81 82 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r126 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r127 75 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=0
+ $X2=13.2 $Y2=0
r128 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=0
+ $X2=13.68 $Y2=0
r129 72 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.305 $Y=0
+ $X2=13.14 $Y2=0
r130 72 74 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=13.305 $Y=0
+ $X2=13.68 $Y2=0
r131 71 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=0
+ $X2=13.2 $Y2=0
r132 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r133 68 71 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=12.72 $Y2=0
r134 68 99 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=10.8 $Y2=0
r135 67 70 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=11.28 $Y=0
+ $X2=12.72 $Y2=0
r136 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r137 65 98 10.873 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=11.2 $Y=0 $X2=10.965
+ $Y2=0
r138 65 67 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=11.2 $Y=0 $X2=11.28
+ $Y2=0
r139 64 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.975 $Y=0
+ $X2=13.14 $Y2=0
r140 64 70 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=12.975 $Y=0
+ $X2=12.72 $Y2=0
r141 63 99 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=8.4 $Y=0 $X2=10.8
+ $Y2=0
r142 63 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=7.92
+ $Y2=0
r143 62 63 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r144 60 95 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.22 $Y=0 $X2=8.055
+ $Y2=0
r145 60 62 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=8.22 $Y=0 $X2=8.4
+ $Y2=0
r146 59 98 10.873 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=10.73 $Y=0
+ $X2=10.965 $Y2=0
r147 59 62 152.011 $w=1.68e-07 $l=2.33e-06 $layer=LI1_cond $X=10.73 $Y=0 $X2=8.4
+ $Y2=0
r148 58 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r149 57 58 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r150 55 89 5.14255 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=5.165 $Y=0 $X2=4.985
+ $Y2=0
r151 55 57 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=5.165 $Y=0
+ $X2=5.52 $Y2=0
r152 54 95 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.89 $Y=0 $X2=8.055
+ $Y2=0
r153 54 57 154.62 $w=1.68e-07 $l=2.37e-06 $layer=LI1_cond $X=7.89 $Y=0 $X2=5.52
+ $Y2=0
r154 53 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r155 53 82 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=3.6
+ $Y2=0
r156 52 86 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=4.56 $Y=0
+ $X2=4.065 $Y2=0
r157 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r158 49 89 5.14255 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=4.805 $Y=0 $X2=4.985
+ $Y2=0
r159 49 52 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=4.805 $Y=0 $X2=4.56
+ $Y2=0
r160 48 82 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=3.6
+ $Y2=0
r161 48 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r162 47 83 154.947 $w=1.68e-07 $l=2.375e-06 $layer=LI1_cond $X=1.2 $Y=0
+ $X2=3.575 $Y2=0
r163 47 48 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r164 45 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=0.78
+ $Y2=0
r165 45 47 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=1.2
+ $Y2=0
r166 42 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r167 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r168 39 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.78
+ $Y2=0
r169 39 41 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=0
+ $X2=0.24 $Y2=0
r170 37 96 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.92
+ $Y2=0
r171 37 58 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=6.96 $Y=0
+ $X2=5.52 $Y2=0
r172 33 35 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=13.14 $Y=0.555
+ $X2=13.14 $Y2=0.965
r173 31 101 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.14 $Y=0.085
+ $X2=13.14 $Y2=0
r174 31 33 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=13.14 $Y=0.085
+ $X2=13.14 $Y2=0.555
r175 27 98 1.91284 $w=4.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.965 $Y=0.085
+ $X2=10.965 $Y2=0
r176 27 29 10.9428 $w=4.68e-07 $l=4.3e-07 $layer=LI1_cond $X=10.965 $Y=0.085
+ $X2=10.965 $Y2=0.515
r177 23 95 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.055 $Y=0.085
+ $X2=8.055 $Y2=0
r178 23 25 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=8.055 $Y=0.085
+ $X2=8.055 $Y2=0.535
r179 19 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=0.085
+ $X2=0.78 $Y2=0
r180 19 21 19.7312 $w=3.28e-07 $l=5.65e-07 $layer=LI1_cond $X=0.78 $Y=0.085
+ $X2=0.78 $Y2=0.65
r181 6 35 182 $w=1.7e-07 $l=7.25655e-07 $layer=licon1_NDIFF $count=1 $X=12.92
+ $Y=0.37 $X2=13.21 $Y2=0.965
r182 6 33 182 $w=1.7e-07 $l=2.98496e-07 $layer=licon1_NDIFF $count=1 $X=12.92
+ $Y=0.37 $X2=13.14 $Y2=0.555
r183 5 29 182 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_NDIFF $count=1 $X=10.765
+ $Y=0.37 $X2=10.965 $Y2=0.515
r184 4 25 182 $w=1.7e-07 $l=2.56905e-07 $layer=licon1_NDIFF $count=1 $X=7.835
+ $Y=0.615 $X2=8.055 $Y2=0.535
r185 3 92 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=4.825
+ $Y=0.135 $X2=4.985 $Y2=0.275
r186 2 85 182 $w=1.7e-07 $l=3.59166e-07 $layer=licon1_NDIFF $count=1 $X=3.52
+ $Y=0.405 $X2=3.82 $Y2=0.275
r187 1 21 182 $w=1.7e-07 $l=2.96985e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.44 $X2=0.78 $Y2=0.65
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTN_1%noxref_24 1 2 9 11 12 15
r37 13 15 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=3.225 $Y=0.425
+ $X2=3.225 $Y2=0.615
r38 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.06 $Y=0.34
+ $X2=3.225 $Y2=0.425
r39 11 12 102.102 $w=1.68e-07 $l=1.565e-06 $layer=LI1_cond $X=3.06 $Y=0.34
+ $X2=1.495 $Y2=0.34
r40 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.33 $Y=0.425
+ $X2=1.495 $Y2=0.34
r41 7 9 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.33 $Y=0.425 $X2=1.33
+ $Y2=0.575
r42 2 15 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=3.08
+ $Y=0.405 $X2=3.225 $Y2=0.615
r43 1 9 182 $w=1.7e-07 $l=2.27706e-07 $layer=licon1_NDIFF $count=1 $X=1.195
+ $Y=0.405 $X2=1.33 $Y2=0.575
.ends

