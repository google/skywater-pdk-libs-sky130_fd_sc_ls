* File: sky130_fd_sc_ls__a41oi_1.spice
* Created: Wed Sep  2 10:53:46 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__a41oi_1.pex.spice"
.subckt sky130_fd_sc_ls__a41oi_1  VNB VPB B1 A4 A3 A2 A1 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A1	A1
* A2	A2
* A3	A3
* A4	A4
* B1	B1
* VPB	VPB
* VNB	VNB
MM1008 N_VGND_M1008_d N_B1_M1008_g N_Y_M1008_s VNB NSHORT L=0.15 W=0.74
+ AD=0.24605 AS=0.2109 PD=1.405 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75002.6 A=0.111 P=1.78 MULT=1
MM1002 A_277_74# N_A4_M1002_g N_VGND_M1008_d VNB NSHORT L=0.15 W=0.74 AD=0.0888
+ AS=0.24605 PD=0.98 PS=1.405 NRD=10.536 NRS=0 M=1 R=4.93333 SA=75001 SB=75001.7
+ A=0.111 P=1.78 MULT=1
MM1003 A_355_74# N_A3_M1003_g A_277_74# VNB NSHORT L=0.15 W=0.74 AD=0.1554
+ AS=0.0888 PD=1.16 PS=0.98 NRD=25.128 NRS=10.536 M=1 R=4.93333 SA=75001.4
+ SB=75001.4 A=0.111 P=1.78 MULT=1
MM1009 A_469_74# N_A2_M1009_g A_355_74# VNB NSHORT L=0.15 W=0.74 AD=0.1554
+ AS=0.1554 PD=1.16 PS=1.16 NRD=25.128 NRS=25.128 M=1 R=4.93333 SA=75002
+ SB=75000.8 A=0.111 P=1.78 MULT=1
MM1000 N_Y_M1000_d N_A1_M1000_g A_469_74# VNB NSHORT L=0.15 W=0.74 AD=0.2109
+ AS=0.1554 PD=2.05 PS=1.16 NRD=0 NRS=25.128 M=1 R=4.93333 SA=75002.6 SB=75000.2
+ A=0.111 P=1.78 MULT=1
MM1007 N_A_116_368#_M1007_d N_B1_M1007_g N_Y_M1007_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.196 AS=0.3304 PD=1.47 PS=2.83 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75002.6 A=0.168 P=2.54 MULT=1
MM1006 N_VPWR_M1006_d N_A4_M1006_g N_A_116_368#_M1007_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.3864 AS=0.196 PD=1.81 PS=1.47 NRD=51.0033 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75002.1 A=0.168 P=2.54 MULT=1
MM1001 N_A_116_368#_M1001_d N_A3_M1001_g N_VPWR_M1006_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.3864 PD=1.42 PS=1.81 NRD=1.7533 NRS=51.0033 M=1 R=7.46667
+ SA=75001.6 SB=75001.2 A=0.168 P=2.54 MULT=1
MM1004 N_VPWR_M1004_d N_A2_M1004_g N_A_116_368#_M1001_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.2296 AS=0.168 PD=1.53 PS=1.42 NRD=11.426 NRS=1.7533 M=1 R=7.46667
+ SA=75002 SB=75000.8 A=0.168 P=2.54 MULT=1
MM1005 N_A_116_368#_M1005_d N_A1_M1005_g N_VPWR_M1004_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.3304 AS=0.2296 PD=2.83 PS=1.53 NRD=1.7533 NRS=11.426 M=1 R=7.46667
+ SA=75002.6 SB=75000.2 A=0.168 P=2.54 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9564 P=11.2
*
.include "sky130_fd_sc_ls__a41oi_1.pxi.spice"
*
.ends
*
*
