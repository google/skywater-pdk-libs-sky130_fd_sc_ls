* File: sky130_fd_sc_ls__nand4bb_1.pex.spice
* Created: Fri Aug 28 13:35:54 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__NAND4BB_1%A_N 1 2 3 5 9 11 15 17
r30 14 17 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=0.315 $Y=0.42
+ $X2=0.52 $Y2=0.42
r31 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.315
+ $Y=0.42 $X2=0.315 $Y2=0.42
r32 11 15 4.38253 $w=3.53e-07 $l=1.35e-07 $layer=LI1_cond $X=0.302 $Y=0.555
+ $X2=0.302 $Y2=0.42
r33 9 10 207.67 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=0.52 $Y=0.97 $X2=0.52
+ $Y2=1.375
r34 6 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.52 $Y=0.585
+ $X2=0.52 $Y2=0.42
r35 6 9 197.415 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=0.52 $Y=0.585
+ $X2=0.52 $Y2=0.97
r36 3 5 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.505 $Y=1.915
+ $X2=0.505 $Y2=2.41
r37 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.505 $Y=1.825 $X2=0.505
+ $Y2=1.915
r38 1 10 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.505 $Y=1.465
+ $X2=0.505 $Y2=1.375
r39 1 2 139.935 $w=1.8e-07 $l=3.6e-07 $layer=POLY_cond $X=0.505 $Y=1.465
+ $X2=0.505 $Y2=1.825
.ends

.subckt PM_SKY130_FD_SC_LS__NAND4BB_1%B_N 1 3 6 8 9
c30 1 0 8.08011e-20 $X=1.055 $Y=1.915
r31 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.01
+ $Y=1.635 $X2=1.01 $Y2=1.635
r32 9 14 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=1.2 $Y=1.635 $X2=1.01
+ $Y2=1.635
r33 8 14 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=0.72 $Y=1.635
+ $X2=1.01 $Y2=1.635
r34 4 13 38.6072 $w=2.91e-07 $l=2.05122e-07 $layer=POLY_cond $X=1.1 $Y=1.47
+ $X2=1.01 $Y2=1.635
r35 4 6 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=1.1 $Y=1.47 $X2=1.1
+ $Y2=0.925
r36 1 13 57.6553 $w=2.91e-07 $l=3.01662e-07 $layer=POLY_cond $X=1.055 $Y=1.915
+ $X2=1.01 $Y2=1.635
r37 1 3 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.055 $Y=1.915
+ $X2=1.055 $Y2=2.41
.ends

.subckt PM_SKY130_FD_SC_LS__NAND4BB_1%A_27_398# 1 2 7 9 10 12 17 19 25 26 27
c61 27 0 8.08011e-20 $X=1.85 $Y=1.215
c62 7 0 3.99753e-20 $X=2.065 $Y=1.765
r63 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.85
+ $Y=1.385 $X2=1.85 $Y2=1.385
r64 27 30 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=1.85 $Y=1.215
+ $X2=1.85 $Y2=1.385
r65 24 25 9.2801 $w=4.58e-07 $l=1.65e-07 $layer=LI1_cond $X=0.305 $Y=1.07
+ $X2=0.47 $Y2=1.07
r66 21 24 2.73018 $w=4.58e-07 $l=1.05e-07 $layer=LI1_cond $X=0.2 $Y=1.07
+ $X2=0.305 $Y2=1.07
r67 19 27 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.685 $Y=1.215
+ $X2=1.85 $Y2=1.215
r68 19 25 79.2674 $w=1.68e-07 $l=1.215e-06 $layer=LI1_cond $X=1.685 $Y=1.215
+ $X2=0.47 $Y2=1.215
r69 17 26 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.28 $Y=2.135
+ $X2=0.28 $Y2=1.97
r70 13 21 6.6364 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=0.2 $Y=1.3 $X2=0.2
+ $Y2=1.07
r71 13 26 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.2 $Y=1.3 $X2=0.2
+ $Y2=1.97
r72 10 31 39.0103 $w=3.67e-07 $l=2.38642e-07 $layer=POLY_cond $X=2.1 $Y=1.22
+ $X2=1.93 $Y2=1.385
r73 10 12 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.1 $Y=1.22 $X2=2.1
+ $Y2=0.74
r74 7 31 67.2473 $w=3.67e-07 $l=4.4238e-07 $layer=POLY_cond $X=2.065 $Y=1.765
+ $X2=1.93 $Y2=1.385
r75 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.065 $Y=1.765
+ $X2=2.065 $Y2=2.4
r76 2 17 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.99 $X2=0.28 $Y2=2.135
r77 1 24 182 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_NDIFF $count=1 $X=0.16
+ $Y=0.86 $X2=0.305 $Y2=1.05
.ends

.subckt PM_SKY130_FD_SC_LS__NAND4BB_1%A_226_398# 1 2 7 9 10 12 15 17 20 22 24 28
+ 32
c71 10 0 1.04695e-19 $X=2.655 $Y=1.765
r72 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.58
+ $Y=1.385 $X2=2.58 $Y2=1.385
r73 29 32 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=2.27 $Y=1.385
+ $X2=2.58 $Y2=1.385
r74 26 28 8.63679 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=1.32 $Y=0.795
+ $X2=1.49 $Y2=0.795
r75 21 29 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.27 $Y=1.55
+ $X2=2.27 $Y2=1.385
r76 21 22 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=2.27 $Y=1.55
+ $X2=2.27 $Y2=1.97
r77 20 29 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.27 $Y=1.22
+ $X2=2.27 $Y2=1.385
r78 19 20 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=2.27 $Y=0.96
+ $X2=2.27 $Y2=1.22
r79 17 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.185 $Y=0.875
+ $X2=2.27 $Y2=0.96
r80 17 28 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=2.185 $Y=0.875
+ $X2=1.49 $Y2=0.875
r81 16 24 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.445 $Y=2.055
+ $X2=1.28 $Y2=2.055
r82 15 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.185 $Y=2.055
+ $X2=2.27 $Y2=1.97
r83 15 16 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=2.185 $Y=2.055
+ $X2=1.445 $Y2=2.055
r84 10 33 77.2841 $w=2.7e-07 $l=4.15812e-07 $layer=POLY_cond $X=2.655 $Y=1.765
+ $X2=2.58 $Y2=1.385
r85 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.655 $Y=1.765
+ $X2=2.655 $Y2=2.4
r86 7 33 38.9026 $w=2.7e-07 $l=2.05122e-07 $layer=POLY_cond $X=2.49 $Y=1.22
+ $X2=2.58 $Y2=1.385
r87 7 9 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.49 $Y=1.22 $X2=2.49
+ $Y2=0.74
r88 2 24 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=1.13
+ $Y=1.99 $X2=1.28 $Y2=2.135
r89 1 26 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=1.175
+ $Y=0.65 $X2=1.32 $Y2=0.795
.ends

.subckt PM_SKY130_FD_SC_LS__NAND4BB_1%C 1 3 4 6 7 8
r39 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.15
+ $Y=1.385 $X2=3.15 $Y2=1.385
r40 8 13 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=3.15 $Y=1.295 $X2=3.15
+ $Y2=1.385
r41 7 8 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.15 $Y=0.925 $X2=3.15
+ $Y2=1.295
r42 4 12 77.2841 $w=2.7e-07 $l=3.82492e-07 $layer=POLY_cond $X=3.155 $Y=1.765
+ $X2=3.15 $Y2=1.385
r43 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.155 $Y=1.765
+ $X2=3.155 $Y2=2.4
r44 1 12 38.9026 $w=2.7e-07 $l=2.05122e-07 $layer=POLY_cond $X=3.06 $Y=1.22
+ $X2=3.15 $Y2=1.385
r45 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.06 $Y=1.22 $X2=3.06
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__NAND4BB_1%D 3 5 7 8 12
r34 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.72
+ $Y=1.515 $X2=3.72 $Y2=1.515
r35 8 12 4.32166 $w=3.98e-07 $l=1.5e-07 $layer=LI1_cond $X=3.685 $Y=1.665
+ $X2=3.685 $Y2=1.515
r36 5 11 52.2586 $w=2.99e-07 $l=2.57391e-07 $layer=POLY_cond $X=3.705 $Y=1.765
+ $X2=3.72 $Y2=1.515
r37 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.705 $Y=1.765
+ $X2=3.705 $Y2=2.4
r38 1 11 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=3.63 $Y=1.35
+ $X2=3.72 $Y2=1.515
r39 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.63 $Y=1.35 $X2=3.63
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__NAND4BB_1%VPWR 1 2 3 12 16 20 23 24 26 27 28 30 46
+ 47 50
r57 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r58 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r59 44 47 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r60 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r61 38 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r62 37 40 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r63 37 38 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r64 35 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=0.78 $Y2=3.33
r65 35 37 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=1.2 $Y2=3.33
r66 33 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r67 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r68 30 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.78 $Y2=3.33
r69 30 32 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.24 $Y2=3.33
r70 28 44 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r71 28 38 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.2 $Y2=3.33
r72 28 40 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r73 26 43 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=3.265 $Y=3.33
+ $X2=3.12 $Y2=3.33
r74 26 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.265 $Y=3.33
+ $X2=3.43 $Y2=3.33
r75 25 46 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=3.595 $Y=3.33
+ $X2=4.08 $Y2=3.33
r76 25 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.595 $Y=3.33
+ $X2=3.43 $Y2=3.33
r77 23 40 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=2.175 $Y=3.33
+ $X2=2.16 $Y2=3.33
r78 23 24 10.1275 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=2.175 $Y=3.33
+ $X2=2.385 $Y2=3.33
r79 22 43 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=2.595 $Y=3.33
+ $X2=3.12 $Y2=3.33
r80 22 24 10.1275 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=2.595 $Y=3.33
+ $X2=2.385 $Y2=3.33
r81 18 27 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.43 $Y=3.245
+ $X2=3.43 $Y2=3.33
r82 18 20 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=3.43 $Y=3.245
+ $X2=3.43 $Y2=2.455
r83 14 24 1.60615 $w=4.2e-07 $l=8.5e-08 $layer=LI1_cond $X=2.385 $Y=3.245
+ $X2=2.385 $Y2=3.33
r84 14 16 11.7988 $w=4.18e-07 $l=4.3e-07 $layer=LI1_cond $X=2.385 $Y=3.245
+ $X2=2.385 $Y2=2.815
r85 10 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=3.245
+ $X2=0.78 $Y2=3.33
r86 10 12 38.764 $w=3.28e-07 $l=1.11e-06 $layer=LI1_cond $X=0.78 $Y=3.245
+ $X2=0.78 $Y2=2.135
r87 3 20 300 $w=1.7e-07 $l=7.07972e-07 $layer=licon1_PDIFF $count=2 $X=3.23
+ $Y=1.84 $X2=3.43 $Y2=2.455
r88 2 16 600 $w=1.7e-07 $l=1.09064e-06 $layer=licon1_PDIFF $count=1 $X=2.14
+ $Y=1.84 $X2=2.385 $Y2=2.815
r89 1 12 300 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=2 $X=0.58
+ $Y=1.99 $X2=0.78 $Y2=2.135
.ends

.subckt PM_SKY130_FD_SC_LS__NAND4BB_1%Y 1 2 3 4 15 19 23 26 27 28 31 34 36 38 39
+ 42 48
c86 42 0 3.99753e-20 $X=2.93 $Y=1.985
c87 23 0 1.04695e-19 $X=3.765 $Y=2.035
r88 46 48 0.104919 $w=5.68e-07 $l=5e-09 $layer=LI1_cond $X=2.81 $Y=2.395
+ $X2=2.81 $Y2=2.4
r89 39 46 7.55418 $w=5.68e-07 $l=3.6e-07 $layer=LI1_cond $X=2.81 $Y=2.035
+ $X2=2.81 $Y2=2.395
r90 39 42 1.04919 $w=5.68e-07 $l=5e-08 $layer=LI1_cond $X=2.81 $Y=2.035 $X2=2.81
+ $Y2=1.985
r91 34 38 3.01263 $w=3.15e-07 $l=1.8262e-07 $layer=LI1_cond $X=4.14 $Y=1.95
+ $X2=3.995 $Y2=2.035
r92 33 34 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=4.14 $Y=1.18
+ $X2=4.14 $Y2=1.95
r93 29 38 3.01263 $w=3.15e-07 $l=8.5e-08 $layer=LI1_cond $X=3.995 $Y=2.12
+ $X2=3.995 $Y2=2.035
r94 29 31 18.0712 $w=4.58e-07 $l=6.95e-07 $layer=LI1_cond $X=3.995 $Y=2.12
+ $X2=3.995 $Y2=2.815
r95 27 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.055 $Y=1.095
+ $X2=4.14 $Y2=1.18
r96 27 28 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=4.055 $Y=1.095
+ $X2=3.655 $Y2=1.095
r97 26 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.57 $Y=1.01
+ $X2=3.655 $Y2=1.095
r98 25 26 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=3.57 $Y=0.62
+ $X2=3.57 $Y2=1.01
r99 24 39 7.98728 $w=1.7e-07 $l=2.85e-07 $layer=LI1_cond $X=3.095 $Y=2.035
+ $X2=2.81 $Y2=2.035
r100 23 38 3.63293 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=3.765 $Y=2.035
+ $X2=3.995 $Y2=2.035
r101 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.765 $Y=2.035
+ $X2=3.095 $Y2=2.035
r102 20 36 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.005 $Y=2.395
+ $X2=1.84 $Y2=2.395
r103 19 46 7.98728 $w=1.7e-07 $l=2.85e-07 $layer=LI1_cond $X=2.525 $Y=2.395
+ $X2=2.81 $Y2=2.395
r104 19 20 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.525 $Y=2.395
+ $X2=2.005 $Y2=2.395
r105 15 25 7.28469 $w=2.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=3.485 $Y=0.485
+ $X2=3.57 $Y2=0.62
r106 15 17 68.2929 $w=2.68e-07 $l=1.6e-06 $layer=LI1_cond $X=3.485 $Y=0.485
+ $X2=1.885 $Y2=0.485
r107 4 38 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=3.78
+ $Y=1.84 $X2=3.93 $Y2=2.115
r108 4 31 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=3.78
+ $Y=1.84 $X2=3.93 $Y2=2.815
r109 3 48 300 $w=1.7e-07 $l=6.5238e-07 $layer=licon1_PDIFF $count=2 $X=2.73
+ $Y=1.84 $X2=2.93 $Y2=2.4
r110 3 42 600 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=1 $X=2.73
+ $Y=1.84 $X2=2.93 $Y2=1.985
r111 2 36 300 $w=1.7e-07 $l=7.03776e-07 $layer=licon1_PDIFF $count=2 $X=1.695
+ $Y=1.84 $X2=1.84 $Y2=2.475
r112 1 17 182 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=1 $X=1.74
+ $Y=0.37 $X2=1.885 $Y2=0.525
.ends

.subckt PM_SKY130_FD_SC_LS__NAND4BB_1%VGND 1 2 11 13 15 17 19 28 32
r37 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r38 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r39 26 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r40 25 26 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r41 23 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r42 22 25 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=3.6
+ $Y2=0
r43 22 23 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r44 20 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.98 $Y=0 $X2=0.815
+ $Y2=0
r45 20 22 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.98 $Y=0 $X2=1.2
+ $Y2=0
r46 19 31 4.63344 $w=1.7e-07 $l=2.47e-07 $layer=LI1_cond $X=3.825 $Y=0 $X2=4.072
+ $Y2=0
r47 19 25 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=3.825 $Y=0 $X2=3.6
+ $Y2=0
r48 17 26 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.6
+ $Y2=0
r49 17 23 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.2
+ $Y2=0
r50 13 31 3.13273 $w=3.3e-07 $l=1.19143e-07 $layer=LI1_cond $X=3.99 $Y=0.085
+ $X2=4.072 $Y2=0
r51 13 15 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=3.99 $Y=0.085
+ $X2=3.99 $Y2=0.595
r52 9 28 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=0.085
+ $X2=0.815 $Y2=0
r53 9 11 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.815 $Y=0.085
+ $X2=0.815 $Y2=0.795
r54 2 15 182 $w=1.7e-07 $l=3.81248e-07 $layer=licon1_NDIFF $count=1 $X=3.705
+ $Y=0.37 $X2=3.99 $Y2=0.595
r55 1 11 182 $w=1.7e-07 $l=2.6533e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.695 $X2=0.815 $Y2=0.795
.ends

