* NGSPICE file created from sky130_fd_sc_ls__a32oi_1.ext - technology: sky130A

.subckt sky130_fd_sc_ls__a32oi_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
M1000 VGND A3 a_469_74# VNB nshort w=740000u l=150000u
+  ad=4.403e+11p pd=4.15e+06u as=3.108e+11p ps=2.32e+06u
M1001 a_27_368# A2 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=1.1816e+12p pd=8.83e+06u as=1.0472e+12p ps=6.35e+06u
M1002 a_119_74# B2 VGND VNB nshort w=740000u l=150000u
+  ad=1.776e+11p pd=1.96e+06u as=0p ps=0u
M1003 VPWR A3 a_27_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_27_368# B1 Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.92e+11p ps=2.94e+06u
M1005 a_391_74# A1 Y VNB nshort w=740000u l=150000u
+  ad=1.776e+11p pd=1.96e+06u as=6.068e+11p ps=3.12e+06u
M1006 Y B2 a_27_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_469_74# A2 a_391_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y B1 a_119_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR A1 a_27_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

