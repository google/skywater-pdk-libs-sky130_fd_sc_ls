* NGSPICE file created from sky130_fd_sc_ls__clkbuf_4.ext - technology: sky130A

.subckt sky130_fd_sc_ls__clkbuf_4 A VGND VNB VPB VPWR X
M1000 VPWR a_83_270# X VPB phighvt w=1.12e+06u l=150000u
+  ad=1.0584e+12p pd=8.61e+06u as=6.72e+11p ps=5.68e+06u
M1001 VGND a_83_270# X VNB nshort w=420000u l=150000u
+  ad=3.969e+11p pd=4.41e+06u as=2.52e+11p ps=2.88e+06u
M1002 a_83_270# A VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=0p ps=0u
M1003 a_83_270# A VGND VNB nshort w=420000u l=150000u
+  ad=1.26e+11p pd=1.44e+06u as=0p ps=0u
M1004 X a_83_270# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 X a_83_270# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR a_83_270# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_83_270# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_83_270# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND a_83_270# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

