* File: sky130_fd_sc_ls__nor2_8.spice
* Created: Fri Aug 28 13:37:18 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__nor2_8.pex.spice"
.subckt sky130_fd_sc_ls__nor2_8  VNB VPB A B VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1004 N_VGND_M1004_d N_A_M1004_g N_Y_M1004_s VNB NSHORT L=0.15 W=0.74 AD=0.7881
+ AS=0.1295 PD=3.61 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75001 SB=75004.8
+ A=0.111 P=1.78 MULT=1
MM1007 N_VGND_M1007_d N_A_M1007_g N_Y_M1004_s VNB NSHORT L=0.15 W=0.74 AD=0.2775
+ AS=0.1295 PD=1.49 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.5 SB=75004.3
+ A=0.111 P=1.78 MULT=1
MM1012 N_VGND_M1007_d N_A_M1012_g N_Y_M1012_s VNB NSHORT L=0.15 W=0.74 AD=0.2775
+ AS=0.1295 PD=1.49 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.4 SB=75003.4
+ A=0.111 P=1.78 MULT=1
MM1015 N_VGND_M1015_d N_A_M1015_g N_Y_M1012_s VNB NSHORT L=0.15 W=0.74 AD=0.1295
+ AS=0.1295 PD=1.09 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75002.9 SB=75002.9
+ A=0.111 P=1.78 MULT=1
MM1003 N_VGND_M1015_d N_B_M1003_g N_Y_M1003_s VNB NSHORT L=0.15 W=0.74 AD=0.1295
+ AS=0.35705 PD=1.09 PS=1.705 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75003.4
+ SB=75002.4 A=0.111 P=1.78 MULT=1
MM1009 N_VGND_M1009_d N_B_M1009_g N_Y_M1003_s VNB NSHORT L=0.15 W=0.74 AD=0.1554
+ AS=0.35705 PD=1.16 PS=1.705 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75004.5
+ SB=75001.3 A=0.111 P=1.78 MULT=1
MM1010 N_VGND_M1009_d N_B_M1010_g N_Y_M1010_s VNB NSHORT L=0.15 W=0.74 AD=0.1554
+ AS=0.1036 PD=1.16 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75005.1 SB=75000.7
+ A=0.111 P=1.78 MULT=1
MM1020 N_VGND_M1020_d N_B_M1020_g N_Y_M1010_s VNB NSHORT L=0.15 W=0.74 AD=0.2627
+ AS=0.1036 PD=2.19 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75005.5 SB=75000.3
+ A=0.111 P=1.78 MULT=1
MM1000 N_A_27_368#_M1000_d N_A_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.196 PD=2.83 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75000.2 SB=75007.4 A=0.168 P=2.54 MULT=1
MM1005 N_A_27_368#_M1005_d N_A_M1005_g N_VPWR_M1000_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75006.9 A=0.168 P=2.54 MULT=1
MM1013 N_A_27_368#_M1005_d N_A_M1013_g N_VPWR_M1013_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.2 SB=75006.4 A=0.168 P=2.54 MULT=1
MM1016 N_A_27_368#_M1016_d N_A_M1016_g N_VPWR_M1013_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.6 SB=75006 A=0.168 P=2.54 MULT=1
MM1017 N_A_27_368#_M1016_d N_A_M1017_g N_VPWR_M1017_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75002.1 SB=75005.5 A=0.168 P=2.54 MULT=1
MM1019 N_A_27_368#_M1019_d N_A_M1019_g N_VPWR_M1017_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.6 SB=75005 A=0.168 P=2.54 MULT=1
MM1021 N_A_27_368#_M1019_d N_A_M1021_g N_VPWR_M1021_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.224 PD=1.42 PS=1.52 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75003 SB=75004.6 A=0.168 P=2.54 MULT=1
MM1023 N_A_27_368#_M1023_d N_A_M1023_g N_VPWR_M1021_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.224 PD=1.42 PS=1.52 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75003.6 SB=75004 A=0.168 P=2.54 MULT=1
MM1001 N_A_27_368#_M1023_d N_B_M1001_g N_Y_M1001_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75004 SB=75003.6 A=0.168 P=2.54 MULT=1
MM1002 N_A_27_368#_M1002_d N_B_M1002_g N_Y_M1001_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.196 AS=0.196 PD=1.47 PS=1.47 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75004.5 SB=75003.1 A=0.168 P=2.54 MULT=1
MM1006 N_A_27_368#_M1002_d N_B_M1006_g N_Y_M1006_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.196 AS=0.168 PD=1.47 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75005
+ SB=75002.6 A=0.168 P=2.54 MULT=1
MM1008 N_A_27_368#_M1008_d N_B_M1008_g N_Y_M1006_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75005.5 SB=75002.1 A=0.168 P=2.54 MULT=1
MM1011 N_A_27_368#_M1008_d N_B_M1011_g N_Y_M1011_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75005.9 SB=75001.7 A=0.168 P=2.54 MULT=1
MM1014 N_A_27_368#_M1014_d N_B_M1014_g N_Y_M1011_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.196 AS=0.168 PD=1.47 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75006.4 SB=75001.2 A=0.168 P=2.54 MULT=1
MM1018 N_A_27_368#_M1014_d N_B_M1018_g N_Y_M1018_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.196 AS=0.168 PD=1.47 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75006.9 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1022 N_A_27_368#_M1022_d N_B_M1022_g N_Y_M1018_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3864 AS=0.168 PD=2.93 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75007.3 SB=75000.3 A=0.168 P=2.54 MULT=1
DX24_noxref VNB VPB NWDIODE A=15.8844 P=20.8
*
.include "sky130_fd_sc_ls__nor2_8.pxi.spice"
*
.ends
*
*
