* File: sky130_fd_sc_ls__and2_2.pex.spice
* Created: Wed Sep  2 10:54:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__AND2_2%A 2 3 5 8 10 14 17
c29 14 0 1.00841e-19 $X=0.27 $Y=1.465
r30 16 17 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.5 $Y=1.465
+ $X2=0.515 $Y2=1.465
r31 13 16 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=0.27 $Y=1.465
+ $X2=0.5 $Y2=1.465
r32 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.465 $X2=0.27 $Y2=1.465
r33 10 14 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=0.27 $Y=1.665 $X2=0.27
+ $Y2=1.465
r34 6 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.515 $Y=1.3
+ $X2=0.515 $Y2=1.465
r35 6 8 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.515 $Y=1.3 $X2=0.515
+ $Y2=0.74
r36 3 5 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.5 $Y=1.885 $X2=0.5
+ $Y2=2.46
r37 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.5 $Y=1.795 $X2=0.5
+ $Y2=1.885
r38 1 16 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.5 $Y=1.63 $X2=0.5
+ $Y2=1.465
r39 1 2 64.1371 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.5 $Y=1.63 $X2=0.5
+ $Y2=1.795
.ends

.subckt PM_SKY130_FD_SC_LS__AND2_2%B 3 6 7 9 10 13 14
c45 14 0 4.02182e-20 $X=0.965 $Y=1.465
c46 6 0 1.00841e-19 $X=0.95 $Y=1.795
c47 3 0 1.29733e-19 $X=0.905 $Y=0.74
r48 13 16 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.965 $Y=1.465
+ $X2=0.965 $Y2=1.63
r49 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.965 $Y=1.465
+ $X2=0.965 $Y2=1.3
r50 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.965
+ $Y=1.465 $X2=0.965 $Y2=1.465
r51 10 14 6.10498 $w=4.78e-07 $l=2.45e-07 $layer=LI1_cond $X=0.72 $Y=1.54
+ $X2=0.965 $Y2=1.54
r52 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.95 $Y=1.885
+ $X2=0.95 $Y2=2.46
r53 6 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.95 $Y=1.795 $X2=0.95
+ $Y2=1.885
r54 6 16 64.1371 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.95 $Y=1.795
+ $X2=0.95 $Y2=1.63
r55 3 15 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.905 $Y=0.74
+ $X2=0.905 $Y2=1.3
.ends

.subckt PM_SKY130_FD_SC_LS__AND2_2%A_31_74# 1 2 7 9 10 12 13 15 16 18 21 23 24
+ 25 27 29 31 32 42
c93 42 0 6.76218e-20 $X=1.845 $Y=1.492
c94 10 0 4.02182e-20 $X=1.455 $Y=1.765
r95 42 43 6.45536 $w=4.48e-07 $l=6e-08 $layer=POLY_cond $X=1.845 $Y=1.492
+ $X2=1.905 $Y2=1.492
r96 39 40 4.30357 $w=4.48e-07 $l=4e-08 $layer=POLY_cond $X=1.415 $Y=1.492
+ $X2=1.455 $Y2=1.492
r97 38 42 36.5804 $w=4.48e-07 $l=3.4e-07 $layer=POLY_cond $X=1.505 $Y=1.492
+ $X2=1.845 $Y2=1.492
r98 38 40 5.37946 $w=4.48e-07 $l=5e-08 $layer=POLY_cond $X=1.505 $Y=1.492
+ $X2=1.455 $Y2=1.492
r99 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.505
+ $Y=1.385 $X2=1.505 $Y2=1.385
r100 31 37 8.96794 $w=3.07e-07 $l=2.17612e-07 $layer=LI1_cond $X=1.34 $Y=1.55
+ $X2=1.462 $Y2=1.385
r101 31 32 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=1.34 $Y=1.55 $X2=1.34
+ $Y2=1.95
r102 30 34 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.89 $Y=2.035
+ $X2=0.765 $Y2=2.035
r103 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.255 $Y=2.035
+ $X2=1.34 $Y2=1.95
r104 29 30 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.255 $Y=2.035
+ $X2=0.89 $Y2=2.035
r105 25 34 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.765 $Y=2.12
+ $X2=0.765 $Y2=2.035
r106 25 27 32.0379 $w=2.48e-07 $l=6.95e-07 $layer=LI1_cond $X=0.765 $Y=2.12
+ $X2=0.765 $Y2=2.815
r107 23 37 13.5114 $w=3.07e-07 $l=4.31254e-07 $layer=LI1_cond $X=1.255 $Y=1.045
+ $X2=1.462 $Y2=1.385
r108 23 24 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=1.255 $Y=1.045
+ $X2=0.465 $Y2=1.045
r109 19 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.3 $Y=0.96
+ $X2=0.465 $Y2=1.045
r110 19 21 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=0.3 $Y=0.96
+ $X2=0.3 $Y2=0.515
r111 16 43 28.6558 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=1.905 $Y=1.765
+ $X2=1.905 $Y2=1.492
r112 16 18 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.905 $Y=1.765
+ $X2=1.905 $Y2=2.4
r113 13 42 28.6558 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=1.845 $Y=1.22
+ $X2=1.845 $Y2=1.492
r114 13 15 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.845 $Y=1.22
+ $X2=1.845 $Y2=0.74
r115 10 40 28.6558 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=1.455 $Y=1.765
+ $X2=1.455 $Y2=1.492
r116 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.455 $Y=1.765
+ $X2=1.455 $Y2=2.4
r117 7 39 28.6558 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=1.415 $Y=1.22
+ $X2=1.415 $Y2=1.492
r118 7 9 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.415 $Y=1.22
+ $X2=1.415 $Y2=0.74
r119 2 34 400 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=1 $X=0.575
+ $Y=1.96 $X2=0.725 $Y2=2.115
r120 2 27 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=0.575
+ $Y=1.96 $X2=0.725 $Y2=2.815
r121 1 21 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.155
+ $Y=0.37 $X2=0.3 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__AND2_2%VPWR 1 2 3 10 12 18 20 22 24 26 31 40 44
r38 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r39 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r40 35 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r41 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r42 32 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.39 $Y=3.33
+ $X2=1.225 $Y2=3.33
r43 32 34 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.39 $Y=3.33
+ $X2=1.68 $Y2=3.33
r44 31 43 4.02656 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=2.045 $Y=3.33
+ $X2=2.222 $Y2=3.33
r45 31 34 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.045 $Y=3.33
+ $X2=1.68 $Y2=3.33
r46 30 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r47 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r48 27 37 4.746 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=0.44 $Y=3.33 $X2=0.22
+ $Y2=3.33
r49 27 29 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.44 $Y=3.33
+ $X2=0.72 $Y2=3.33
r50 26 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.06 $Y=3.33
+ $X2=1.225 $Y2=3.33
r51 26 29 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.06 $Y=3.33
+ $X2=0.72 $Y2=3.33
r52 24 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r53 24 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r54 24 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r55 20 43 3.1166 $w=2.5e-07 $l=1.07912e-07 $layer=LI1_cond $X=2.17 $Y=3.245
+ $X2=2.222 $Y2=3.33
r56 20 22 47.0197 $w=2.48e-07 $l=1.02e-06 $layer=LI1_cond $X=2.17 $Y=3.245
+ $X2=2.17 $Y2=2.225
r57 16 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.225 $Y=3.245
+ $X2=1.225 $Y2=3.33
r58 16 18 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=1.225 $Y=3.245
+ $X2=1.225 $Y2=2.455
r59 12 15 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=0.275 $Y=2.115
+ $X2=0.275 $Y2=2.815
r60 10 37 3.02018 $w=3.3e-07 $l=1.09087e-07 $layer=LI1_cond $X=0.275 $Y=3.245
+ $X2=0.22 $Y2=3.33
r61 10 15 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.275 $Y=3.245
+ $X2=0.275 $Y2=2.815
r62 3 22 300 $w=1.7e-07 $l=4.53845e-07 $layer=licon1_PDIFF $count=2 $X=1.98
+ $Y=1.84 $X2=2.13 $Y2=2.225
r63 2 18 300 $w=1.7e-07 $l=5.86536e-07 $layer=licon1_PDIFF $count=2 $X=1.025
+ $Y=1.96 $X2=1.225 $Y2=2.455
r64 1 15 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.275 $Y2=2.815
r65 1 12 400 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.275 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_LS__AND2_2%X 1 2 7 8 14 16 17 18
c33 7 0 1.29733e-19 $X=1.925 $Y=1.02
r34 17 18 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=1.72 $Y=2.405
+ $X2=1.72 $Y2=2.775
r35 16 17 19.361 $w=2.48e-07 $l=4.2e-07 $layer=LI1_cond $X=1.72 $Y=1.985
+ $X2=1.72 $Y2=2.405
r36 12 16 4.37928 $w=2.48e-07 $l=9.5e-08 $layer=LI1_cond $X=1.72 $Y=1.89
+ $X2=1.72 $Y2=1.985
r37 12 14 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.72 $Y=1.805
+ $X2=1.925 $Y2=1.805
r38 8 14 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.925 $Y=1.72
+ $X2=1.925 $Y2=1.805
r39 7 10 19.526 $w=3.29e-07 $l=5.35817e-07 $layer=LI1_cond $X=1.925 $Y=1.02
+ $X2=1.737 $Y2=0.57
r40 7 8 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.925 $Y=1.02 $X2=1.925
+ $Y2=1.72
r41 2 18 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.53
+ $Y=1.84 $X2=1.68 $Y2=2.815
r42 2 16 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.53
+ $Y=1.84 $X2=1.68 $Y2=1.985
r43 1 10 182 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=1 $X=1.49
+ $Y=0.37 $X2=1.63 $Y2=0.57
.ends

.subckt PM_SKY130_FD_SC_LS__AND2_2%VGND 1 2 9 11 13 15 17 22 28 32
c32 13 0 6.76218e-20 $X=2.09 $Y=0.515
r33 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r34 26 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r35 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r36 23 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.285 $Y=0 $X2=1.12
+ $Y2=0
r37 23 25 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.285 $Y=0 $X2=1.68
+ $Y2=0
r38 22 31 4.55093 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=1.975 $Y=0 $X2=2.187
+ $Y2=0
r39 22 25 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.975 $Y=0 $X2=1.68
+ $Y2=0
r40 19 20 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r41 17 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=1.12
+ $Y2=0
r42 17 19 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=0.72
+ $Y2=0
r43 15 26 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r44 15 20 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r45 15 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r46 11 31 3.04826 $w=3.1e-07 $l=1.09864e-07 $layer=LI1_cond $X=2.13 $Y=0.085
+ $X2=2.187 $Y2=0
r47 11 13 15.9855 $w=3.08e-07 $l=4.3e-07 $layer=LI1_cond $X=2.13 $Y=0.085
+ $X2=2.13 $Y2=0.515
r48 7 28 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=0.085 $X2=1.12
+ $Y2=0
r49 7 9 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=1.12 $Y=0.085
+ $X2=1.12 $Y2=0.57
r50 2 13 182 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_NDIFF $count=1 $X=1.92
+ $Y=0.37 $X2=2.09 $Y2=0.515
r51 1 9 182 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=1 $X=0.98
+ $Y=0.37 $X2=1.12 $Y2=0.57
.ends

