* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__sdfrbp_1 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q Q_N
M1000 a_1320_119# a_1034_392# a_1234_119# VNB nshort w=420000u l=150000u
+  ad=9.87e+10p pd=1.31e+06u as=1.176e+11p ps=1.4e+06u
M1001 VGND a_1747_74# a_2513_424# VNB nshort w=550000u l=150000u
+  ad=1.77802e+12p pd=1.475e+07u as=1.4575e+11p ps=1.63e+06u
M1002 Q_N a_1747_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=2.27322e+12p ps=1.901e+07u
M1003 VGND a_2008_48# a_1966_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1004 a_1234_119# RESET_B VPWR VPB phighvt w=420000u l=150000u
+  ad=2.499e+11p pd=2.87e+06u as=0p ps=0u
M1005 a_2124_74# RESET_B VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1006 Q_N a_1747_74# VGND VNB nshort w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1007 a_2008_48# a_1747_74# a_2124_74# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1008 a_312_81# a_27_74# a_225_81# VNB nshort w=420000u l=150000u
+  ad=1.407e+11p pd=1.51e+06u as=2.499e+11p ps=2.87e+06u
M1009 a_1966_74# a_835_98# a_1747_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=4.519e+11p ps=3.17e+06u
M1010 a_1332_457# a_835_98# a_1234_119# VPB phighvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1011 VGND RESET_B a_1397_119# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1012 a_409_81# D a_312_81# VNB nshort w=420000u l=150000u
+  ad=3.339e+11p pd=3.27e+06u as=0p ps=0u
M1013 a_1747_74# a_835_98# a_1367_93# VPB phighvt w=1e+06u l=150000u
+  ad=4.1485e+11p pd=3.51e+06u as=3e+11p ps=2.6e+06u
M1014 a_409_81# D a_338_464# VPB phighvt w=640000u l=150000u
+  ad=5.047e+11p pd=5.18e+06u as=1.728e+11p ps=1.82e+06u
M1015 a_1969_489# a_1034_392# a_1747_74# VPB phighvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1016 a_225_81# SCD a_545_81# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1017 VPWR a_2008_48# a_1969_489# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 Q a_2513_424# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.08e+11p pd=2.79e+06u as=0p ps=0u
M1019 a_512_464# a_27_74# a_409_81# VPB phighvt w=640000u l=150000u
+  ad=2.56e+11p pd=2.08e+06u as=0p ps=0u
M1020 a_1747_74# a_1034_392# a_1367_93# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=1.856e+11p ps=1.86e+06u
M1021 a_1397_119# a_1367_93# a_1320_119# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_545_81# SCE a_409_81# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VPWR SCD a_512_464# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VPWR CLK a_835_98# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.95e+11p ps=2.59e+06u
M1025 VGND CLK a_835_98# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.619e+11p ps=2.38e+06u
M1026 VPWR SCE a_27_74# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=5.792e+11p ps=3.09e+06u
M1027 a_2008_48# RESET_B VPWR VPB phighvt w=420000u l=150000u
+  ad=1.26e+11p pd=1.44e+06u as=0p ps=0u
M1028 a_1034_392# a_835_98# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.95e+11p pd=2.59e+06u as=0p ps=0u
M1029 VPWR a_1747_74# a_2513_424# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=2.31e+11p ps=2.23e+06u
M1030 a_1367_93# a_1234_119# VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 Q a_2513_424# VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1032 VGND SCE a_27_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1033 a_1034_392# a_835_98# VGND VNB nshort w=740000u l=150000u
+  ad=1.961e+11p pd=2.01e+06u as=0p ps=0u
M1034 VPWR a_1367_93# a_1332_457# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_1234_119# a_835_98# a_409_81# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 VGND RESET_B a_225_81# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_338_464# SCE VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 a_409_81# RESET_B VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_1234_119# a_1034_392# a_409_81# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1040 a_1367_93# a_1234_119# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1041 VPWR a_1747_74# a_2008_48# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
