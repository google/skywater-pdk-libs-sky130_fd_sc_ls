* File: sky130_fd_sc_ls__a22oi_4.pxi.spice
* Created: Wed Sep  2 10:50:44 2020
* 
x_PM_SKY130_FD_SC_LS__A22OI_4%B2 N_B2_c_125_n N_B2_M1005_g N_B2_M1007_g
+ N_B2_M1013_g N_B2_c_126_n N_B2_M1010_g N_B2_M1017_g N_B2_c_127_n N_B2_M1011_g
+ N_B2_M1028_g N_B2_c_128_n N_B2_M1020_g B2 B2 B2 N_B2_c_129_n N_B2_c_124_n
+ PM_SKY130_FD_SC_LS__A22OI_4%B2
x_PM_SKY130_FD_SC_LS__A22OI_4%B1 N_B1_M1004_g N_B1_c_209_n N_B1_M1000_g
+ N_B1_M1006_g N_B1_c_210_n N_B1_M1008_g N_B1_M1023_g N_B1_c_211_n N_B1_M1016_g
+ N_B1_M1024_g N_B1_c_212_n N_B1_M1025_g B1 B1 N_B1_c_208_n
+ PM_SKY130_FD_SC_LS__A22OI_4%B1
x_PM_SKY130_FD_SC_LS__A22OI_4%A1 N_A1_c_308_n N_A1_M1001_g N_A1_c_300_n
+ N_A1_M1012_g N_A1_c_309_n N_A1_M1021_g N_A1_M1019_g N_A1_c_310_n N_A1_M1022_g
+ N_A1_M1026_g N_A1_c_311_n N_A1_M1031_g N_A1_M1030_g N_A1_c_305_n A1 A1 A1
+ N_A1_c_307_n PM_SKY130_FD_SC_LS__A22OI_4%A1
x_PM_SKY130_FD_SC_LS__A22OI_4%A2 N_A2_c_396_n N_A2_M1002_g N_A2_M1014_g
+ N_A2_c_397_n N_A2_M1003_g N_A2_M1015_g N_A2_c_398_n N_A2_M1009_g N_A2_M1018_g
+ N_A2_M1029_g N_A2_c_399_n N_A2_M1027_g A2 A2 A2 N_A2_c_394_n N_A2_c_395_n
+ PM_SKY130_FD_SC_LS__A22OI_4%A2
x_PM_SKY130_FD_SC_LS__A22OI_4%A_45_368# N_A_45_368#_M1005_d N_A_45_368#_M1010_d
+ N_A_45_368#_M1020_d N_A_45_368#_M1008_d N_A_45_368#_M1025_d
+ N_A_45_368#_M1021_s N_A_45_368#_M1031_s N_A_45_368#_M1003_d
+ N_A_45_368#_M1027_d N_A_45_368#_c_468_n N_A_45_368#_c_469_n
+ N_A_45_368#_c_470_n N_A_45_368#_c_486_n N_A_45_368#_c_471_n
+ N_A_45_368#_c_492_n N_A_45_368#_c_472_n N_A_45_368#_c_501_n
+ N_A_45_368#_c_473_n N_A_45_368#_c_474_n N_A_45_368#_c_509_n
+ N_A_45_368#_c_517_n N_A_45_368#_c_475_n N_A_45_368#_c_524_n
+ N_A_45_368#_c_476_n N_A_45_368#_c_535_n N_A_45_368#_c_477_n
+ N_A_45_368#_c_541_n N_A_45_368#_c_478_n N_A_45_368#_c_479_n
+ N_A_45_368#_c_480_n N_A_45_368#_c_481_n N_A_45_368#_c_482_n
+ N_A_45_368#_c_530_n N_A_45_368#_c_533_n N_A_45_368#_c_548_n
+ PM_SKY130_FD_SC_LS__A22OI_4%A_45_368#
x_PM_SKY130_FD_SC_LS__A22OI_4%Y N_Y_M1004_s N_Y_M1023_s N_Y_M1012_s N_Y_M1026_s
+ N_Y_M1005_s N_Y_M1011_s N_Y_M1000_s N_Y_M1016_s N_Y_c_624_n N_Y_c_627_n
+ N_Y_c_629_n N_Y_c_633_n N_Y_c_635_n N_Y_c_642_n N_Y_c_645_n N_Y_c_618_n
+ N_Y_c_619_n N_Y_c_655_n N_Y_c_623_n N_Y_c_620_n N_Y_c_637_n N_Y_c_668_n
+ N_Y_c_670_n N_Y_c_621_n N_Y_c_622_n Y Y PM_SKY130_FD_SC_LS__A22OI_4%Y
x_PM_SKY130_FD_SC_LS__A22OI_4%VPWR N_VPWR_M1001_d N_VPWR_M1022_d N_VPWR_M1002_s
+ N_VPWR_M1009_s N_VPWR_c_733_n N_VPWR_c_734_n N_VPWR_c_735_n N_VPWR_c_736_n
+ N_VPWR_c_737_n N_VPWR_c_738_n N_VPWR_c_739_n N_VPWR_c_740_n VPWR
+ N_VPWR_c_741_n N_VPWR_c_742_n N_VPWR_c_743_n N_VPWR_c_732_n N_VPWR_c_745_n
+ N_VPWR_c_746_n PM_SKY130_FD_SC_LS__A22OI_4%VPWR
x_PM_SKY130_FD_SC_LS__A22OI_4%A_48_74# N_A_48_74#_M1007_s N_A_48_74#_M1013_s
+ N_A_48_74#_M1028_s N_A_48_74#_M1006_d N_A_48_74#_M1024_d N_A_48_74#_c_833_n
+ N_A_48_74#_c_834_n N_A_48_74#_c_835_n N_A_48_74#_c_836_n N_A_48_74#_c_837_n
+ N_A_48_74#_c_838_n N_A_48_74#_c_839_n N_A_48_74#_c_840_n N_A_48_74#_c_841_n
+ N_A_48_74#_c_842_n PM_SKY130_FD_SC_LS__A22OI_4%A_48_74#
x_PM_SKY130_FD_SC_LS__A22OI_4%VGND N_VGND_M1007_d N_VGND_M1017_d N_VGND_M1014_d
+ N_VGND_M1018_d N_VGND_c_899_n N_VGND_c_900_n N_VGND_c_901_n N_VGND_c_902_n
+ N_VGND_c_903_n N_VGND_c_904_n N_VGND_c_905_n N_VGND_c_906_n VGND
+ N_VGND_c_907_n N_VGND_c_908_n N_VGND_c_909_n N_VGND_c_910_n N_VGND_c_911_n
+ N_VGND_c_912_n PM_SKY130_FD_SC_LS__A22OI_4%VGND
x_PM_SKY130_FD_SC_LS__A22OI_4%A_840_74# N_A_840_74#_M1012_d N_A_840_74#_M1019_d
+ N_A_840_74#_M1030_d N_A_840_74#_M1015_s N_A_840_74#_M1029_s
+ N_A_840_74#_c_993_n N_A_840_74#_c_994_n N_A_840_74#_c_995_n
+ N_A_840_74#_c_996_n N_A_840_74#_c_997_n N_A_840_74#_c_998_n
+ N_A_840_74#_c_999_n N_A_840_74#_c_1000_n N_A_840_74#_c_1001_n
+ PM_SKY130_FD_SC_LS__A22OI_4%A_840_74#
cc_1 VNB N_B2_M1007_g 0.0318708f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=0.74
cc_2 VNB N_B2_M1013_g 0.0230578f $X=-0.19 $Y=-0.245 $X2=1.01 $Y2=0.74
cc_3 VNB N_B2_M1017_g 0.0224931f $X=-0.19 $Y=-0.245 $X2=1.44 $Y2=0.74
cc_4 VNB N_B2_M1028_g 0.0229726f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=0.74
cc_5 VNB N_B2_c_124_n 0.08144f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=1.557
cc_6 VNB N_B1_M1004_g 0.0213573f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=2.4
cc_7 VNB N_B1_M1006_g 0.0206638f $X=-0.19 $Y=-0.245 $X2=1.01 $Y2=0.74
cc_8 VNB N_B1_M1023_g 0.0206542f $X=-0.19 $Y=-0.245 $X2=1.44 $Y2=0.74
cc_9 VNB N_B1_M1024_g 0.0248723f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=0.74
cc_10 VNB B1 0.0014908f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_11 VNB N_B1_c_208_n 0.0814765f $X=-0.19 $Y=-0.245 $X2=1.79 $Y2=1.515
cc_12 VNB N_A1_c_300_n 0.013191f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.35
cc_13 VNB N_A1_M1012_g 0.0269428f $X=-0.19 $Y=-0.245 $X2=1.01 $Y2=1.35
cc_14 VNB N_A1_M1019_g 0.0234062f $X=-0.19 $Y=-0.245 $X2=1.44 $Y2=1.35
cc_15 VNB N_A1_M1026_g 0.0234234f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=1.35
cc_16 VNB N_A1_M1030_g 0.0240886f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_17 VNB N_A1_c_305_n 0.0114234f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_18 VNB A1 0.00163664f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=1.557
cc_19 VNB N_A1_c_307_n 0.063517f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A2_M1014_g 0.0230056f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=0.74
cc_21 VNB N_A2_M1015_g 0.0230578f $X=-0.19 $Y=-0.245 $X2=1.025 $Y2=2.4
cc_22 VNB N_A2_M1018_g 0.0224931f $X=-0.19 $Y=-0.245 $X2=1.475 $Y2=2.4
cc_23 VNB N_A2_M1029_g 0.0326336f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=0.74
cc_24 VNB N_A2_c_394_n 0.00356131f $X=-0.19 $Y=-0.245 $X2=1.79 $Y2=1.515
cc_25 VNB N_A2_c_395_n 0.0801686f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=1.557
cc_26 VNB N_Y_c_618_n 0.00224682f $X=-0.19 $Y=-0.245 $X2=1.79 $Y2=1.515
cc_27 VNB N_Y_c_619_n 0.00229069f $X=-0.19 $Y=-0.245 $X2=1.79 $Y2=1.515
cc_28 VNB N_Y_c_620_n 0.0229782f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_Y_c_621_n 0.00510981f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_Y_c_622_n 0.00826357f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VPWR_c_732_n 0.342803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_48_74#_c_833_n 0.0270834f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_48_74#_c_834_n 0.00400183f $X=-0.19 $Y=-0.245 $X2=1.475 $Y2=2.4
cc_34 VNB N_A_48_74#_c_835_n 0.0120073f $X=-0.19 $Y=-0.245 $X2=1.475 $Y2=2.4
cc_35 VNB N_A_48_74#_c_836_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=0.74
cc_36 VNB N_A_48_74#_c_837_n 0.0102323f $X=-0.19 $Y=-0.245 $X2=1.925 $Y2=1.765
cc_37 VNB N_A_48_74#_c_838_n 0.00299433f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_48_74#_c_839_n 0.00211517f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_48_74#_c_840_n 0.00938494f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.557
cc_40 VNB N_A_48_74#_c_841_n 0.00178779f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=1.515
cc_41 VNB N_A_48_74#_c_842_n 0.00164253f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=1.515
cc_42 VNB N_VGND_c_899_n 0.00481913f $X=-0.19 $Y=-0.245 $X2=1.44 $Y2=1.35
cc_43 VNB N_VGND_c_900_n 0.00334323f $X=-0.19 $Y=-0.245 $X2=1.475 $Y2=1.765
cc_44 VNB N_VGND_c_901_n 0.00481913f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=0.74
cc_45 VNB N_VGND_c_902_n 0.00497771f $X=-0.19 $Y=-0.245 $X2=1.925 $Y2=2.4
cc_46 VNB N_VGND_c_903_n 0.108097f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_47 VNB N_VGND_c_904_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_48 VNB N_VGND_c_905_n 0.0172524f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_906_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_907_n 0.0200958f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=1.557
cc_51 VNB N_VGND_c_908_n 0.0172524f $X=-0.19 $Y=-0.245 $X2=1.44 $Y2=1.557
cc_52 VNB N_VGND_c_909_n 0.0231293f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_910_n 0.445534f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_911_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_912_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_840_74#_c_993_n 0.00754101f $X=-0.19 $Y=-0.245 $X2=1.44 $Y2=0.74
cc_57 VNB N_A_840_74#_c_994_n 0.0016059f $X=-0.19 $Y=-0.245 $X2=1.475 $Y2=2.4
cc_58 VNB N_A_840_74#_c_995_n 0.00257879f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=0.74
cc_59 VNB N_A_840_74#_c_996_n 0.00230622f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_840_74#_c_997_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=1.925 $Y2=2.4
cc_61 VNB N_A_840_74#_c_998_n 0.0166385f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_62 VNB N_A_840_74#_c_999_n 0.0281813f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_840_74#_c_1000_n 0.00646965f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=1.515
cc_64 VNB N_A_840_74#_c_1001_n 0.00178779f $X=-0.19 $Y=-0.245 $X2=1.44 $Y2=1.557
cc_65 VPB N_B2_c_125_n 0.0183915f $X=-0.19 $Y=1.66 $X2=0.575 $Y2=1.765
cc_66 VPB N_B2_c_126_n 0.014659f $X=-0.19 $Y=1.66 $X2=1.025 $Y2=1.765
cc_67 VPB N_B2_c_127_n 0.0146598f $X=-0.19 $Y=1.66 $X2=1.475 $Y2=1.765
cc_68 VPB N_B2_c_128_n 0.0148576f $X=-0.19 $Y=1.66 $X2=1.925 $Y2=1.765
cc_69 VPB N_B2_c_129_n 0.00839387f $X=-0.19 $Y=1.66 $X2=1.79 $Y2=1.515
cc_70 VPB N_B2_c_124_n 0.0494747f $X=-0.19 $Y=1.66 $X2=1.87 $Y2=1.557
cc_71 VPB N_B1_c_209_n 0.0147854f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=0.74
cc_72 VPB N_B1_c_210_n 0.0146577f $X=-0.19 $Y=1.66 $X2=1.025 $Y2=1.765
cc_73 VPB N_B1_c_211_n 0.0146889f $X=-0.19 $Y=1.66 $X2=1.475 $Y2=1.765
cc_74 VPB N_B1_c_212_n 0.0147551f $X=-0.19 $Y=1.66 $X2=1.925 $Y2=1.765
cc_75 VPB B1 0.00685912f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_76 VPB N_B1_c_208_n 0.0481133f $X=-0.19 $Y=1.66 $X2=1.79 $Y2=1.515
cc_77 VPB N_A1_c_308_n 0.0153891f $X=-0.19 $Y=1.66 $X2=0.575 $Y2=1.765
cc_78 VPB N_A1_c_309_n 0.0149981f $X=-0.19 $Y=1.66 $X2=1.01 $Y2=0.74
cc_79 VPB N_A1_c_310_n 0.0170119f $X=-0.19 $Y=1.66 $X2=1.44 $Y2=0.74
cc_80 VPB N_A1_c_311_n 0.0174109f $X=-0.19 $Y=1.66 $X2=1.87 $Y2=0.74
cc_81 VPB N_A1_c_305_n 0.00646634f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.58
cc_82 VPB A1 0.010329f $X=-0.19 $Y=1.66 $X2=0.575 $Y2=1.557
cc_83 VPB N_A1_c_307_n 0.0429772f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_84 VPB N_A2_c_396_n 0.0153053f $X=-0.19 $Y=1.66 $X2=0.575 $Y2=1.765
cc_85 VPB N_A2_c_397_n 0.0149968f $X=-0.19 $Y=1.66 $X2=1.01 $Y2=1.35
cc_86 VPB N_A2_c_398_n 0.014996f $X=-0.19 $Y=1.66 $X2=1.44 $Y2=1.35
cc_87 VPB N_A2_c_399_n 0.0199141f $X=-0.19 $Y=1.66 $X2=1.925 $Y2=1.765
cc_88 VPB N_A2_c_394_n 0.0113536f $X=-0.19 $Y=1.66 $X2=1.79 $Y2=1.515
cc_89 VPB N_A2_c_395_n 0.0492591f $X=-0.19 $Y=1.66 $X2=1.87 $Y2=1.557
cc_90 VPB N_A_45_368#_c_468_n 0.0454805f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_91 VPB N_A_45_368#_c_469_n 0.00259172f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_92 VPB N_A_45_368#_c_470_n 0.00939918f $X=-0.19 $Y=1.66 $X2=0.575 $Y2=1.557
cc_93 VPB N_A_45_368#_c_471_n 0.00213603f $X=-0.19 $Y=1.66 $X2=1.01 $Y2=1.557
cc_94 VPB N_A_45_368#_c_472_n 0.00213603f $X=-0.19 $Y=1.66 $X2=1.79 $Y2=1.515
cc_95 VPB N_A_45_368#_c_473_n 0.00479765f $X=-0.19 $Y=1.66 $X2=0.77 $Y2=1.565
cc_96 VPB N_A_45_368#_c_474_n 0.00287037f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_A_45_368#_c_475_n 0.00216998f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_A_45_368#_c_476_n 0.00216998f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB N_A_45_368#_c_477_n 0.00180921f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 VPB N_A_45_368#_c_478_n 0.0169052f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB N_A_45_368#_c_479_n 0.0345863f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_102 VPB N_A_45_368#_c_480_n 0.0021839f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 VPB N_A_45_368#_c_481_n 0.0021839f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB N_A_45_368#_c_482_n 0.0021839f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_105 VPB N_Y_c_623_n 0.00251102f $X=-0.19 $Y=1.66 $X2=0.77 $Y2=1.565
cc_106 VPB N_VPWR_c_733_n 0.00335558f $X=-0.19 $Y=1.66 $X2=1.44 $Y2=1.35
cc_107 VPB N_VPWR_c_734_n 0.00948205f $X=-0.19 $Y=1.66 $X2=1.475 $Y2=1.765
cc_108 VPB N_VPWR_c_735_n 0.0026822f $X=-0.19 $Y=1.66 $X2=1.87 $Y2=0.74
cc_109 VPB N_VPWR_c_736_n 0.00329129f $X=-0.19 $Y=1.66 $X2=1.925 $Y2=2.4
cc_110 VPB N_VPWR_c_737_n 0.0994019f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_111 VPB N_VPWR_c_738_n 0.00601644f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.58
cc_112 VPB N_VPWR_c_739_n 0.0164465f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_VPWR_c_740_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_VPWR_c_741_n 0.0175706f $X=-0.19 $Y=1.66 $X2=1.79 $Y2=1.557
cc_115 VPB N_VPWR_c_742_n 0.0175706f $X=-0.19 $Y=1.66 $X2=1.925 $Y2=1.557
cc_116 VPB N_VPWR_c_743_n 0.0212096f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_732_n 0.0973001f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_745_n 0.0088221f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_746_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 N_B2_M1028_g N_B1_M1004_g 0.0189918f $X=1.87 $Y=0.74 $X2=0 $Y2=0
cc_121 N_B2_c_128_n N_B1_c_209_n 0.0255159f $X=1.925 $Y=1.765 $X2=0 $Y2=0
cc_122 N_B2_c_129_n B1 0.0227446f $X=1.79 $Y=1.515 $X2=0 $Y2=0
cc_123 N_B2_c_124_n B1 0.00203324f $X=1.87 $Y=1.557 $X2=0 $Y2=0
cc_124 N_B2_c_129_n N_B1_c_208_n 7.84039e-19 $X=1.79 $Y=1.515 $X2=0 $Y2=0
cc_125 N_B2_c_124_n N_B1_c_208_n 0.0234647f $X=1.87 $Y=1.557 $X2=0 $Y2=0
cc_126 N_B2_c_125_n N_A_45_368#_c_468_n 0.00835508f $X=0.575 $Y=1.765 $X2=0
+ $Y2=0
cc_127 N_B2_c_125_n N_A_45_368#_c_469_n 0.0137046f $X=0.575 $Y=1.765 $X2=0 $Y2=0
cc_128 N_B2_c_126_n N_A_45_368#_c_469_n 0.0108414f $X=1.025 $Y=1.765 $X2=0 $Y2=0
cc_129 N_B2_c_125_n N_A_45_368#_c_486_n 6.2388e-19 $X=0.575 $Y=1.765 $X2=0 $Y2=0
cc_130 N_B2_c_126_n N_A_45_368#_c_486_n 0.00850468f $X=1.025 $Y=1.765 $X2=0
+ $Y2=0
cc_131 N_B2_c_127_n N_A_45_368#_c_486_n 0.00830261f $X=1.475 $Y=1.765 $X2=0
+ $Y2=0
cc_132 N_B2_c_128_n N_A_45_368#_c_486_n 5.7112e-19 $X=1.925 $Y=1.765 $X2=0 $Y2=0
cc_133 N_B2_c_127_n N_A_45_368#_c_471_n 0.0108414f $X=1.475 $Y=1.765 $X2=0 $Y2=0
cc_134 N_B2_c_128_n N_A_45_368#_c_471_n 0.0108414f $X=1.925 $Y=1.765 $X2=0 $Y2=0
cc_135 N_B2_c_127_n N_A_45_368#_c_492_n 5.7112e-19 $X=1.475 $Y=1.765 $X2=0 $Y2=0
cc_136 N_B2_c_128_n N_A_45_368#_c_492_n 0.00828741f $X=1.925 $Y=1.765 $X2=0
+ $Y2=0
cc_137 N_B2_c_126_n N_A_45_368#_c_480_n 0.00175197f $X=1.025 $Y=1.765 $X2=0
+ $Y2=0
cc_138 N_B2_c_127_n N_A_45_368#_c_480_n 0.00175197f $X=1.475 $Y=1.765 $X2=0
+ $Y2=0
cc_139 N_B2_c_128_n N_A_45_368#_c_481_n 0.00171731f $X=1.925 $Y=1.765 $X2=0
+ $Y2=0
cc_140 N_B2_c_125_n N_Y_c_624_n 0.00203651f $X=0.575 $Y=1.765 $X2=0 $Y2=0
cc_141 N_B2_c_129_n N_Y_c_624_n 0.0193936f $X=1.79 $Y=1.515 $X2=0 $Y2=0
cc_142 N_B2_c_124_n N_Y_c_624_n 0.00124229f $X=1.87 $Y=1.557 $X2=0 $Y2=0
cc_143 N_B2_c_125_n N_Y_c_627_n 0.0082032f $X=0.575 $Y=1.765 $X2=0 $Y2=0
cc_144 N_B2_c_126_n N_Y_c_627_n 0.00576017f $X=1.025 $Y=1.765 $X2=0 $Y2=0
cc_145 N_B2_c_126_n N_Y_c_629_n 0.0126853f $X=1.025 $Y=1.765 $X2=0 $Y2=0
cc_146 N_B2_c_127_n N_Y_c_629_n 0.0126853f $X=1.475 $Y=1.765 $X2=0 $Y2=0
cc_147 N_B2_c_129_n N_Y_c_629_n 0.0477183f $X=1.79 $Y=1.515 $X2=0 $Y2=0
cc_148 N_B2_c_124_n N_Y_c_629_n 0.00169221f $X=1.87 $Y=1.557 $X2=0 $Y2=0
cc_149 N_B2_c_127_n N_Y_c_633_n 0.00532448f $X=1.475 $Y=1.765 $X2=0 $Y2=0
cc_150 N_B2_c_128_n N_Y_c_633_n 0.00532448f $X=1.925 $Y=1.765 $X2=0 $Y2=0
cc_151 N_B2_c_128_n N_Y_c_635_n 0.0139291f $X=1.925 $Y=1.765 $X2=0 $Y2=0
cc_152 N_B2_c_129_n N_Y_c_635_n 0.0106982f $X=1.79 $Y=1.515 $X2=0 $Y2=0
cc_153 N_B2_c_129_n N_Y_c_637_n 0.0150275f $X=1.79 $Y=1.515 $X2=0 $Y2=0
cc_154 N_B2_c_124_n N_Y_c_637_n 0.00104225f $X=1.87 $Y=1.557 $X2=0 $Y2=0
cc_155 N_B2_c_125_n N_VPWR_c_737_n 0.00278271f $X=0.575 $Y=1.765 $X2=0 $Y2=0
cc_156 N_B2_c_126_n N_VPWR_c_737_n 0.00278257f $X=1.025 $Y=1.765 $X2=0 $Y2=0
cc_157 N_B2_c_127_n N_VPWR_c_737_n 0.00278257f $X=1.475 $Y=1.765 $X2=0 $Y2=0
cc_158 N_B2_c_128_n N_VPWR_c_737_n 0.00278257f $X=1.925 $Y=1.765 $X2=0 $Y2=0
cc_159 N_B2_c_125_n N_VPWR_c_732_n 0.00357527f $X=0.575 $Y=1.765 $X2=0 $Y2=0
cc_160 N_B2_c_126_n N_VPWR_c_732_n 0.00353822f $X=1.025 $Y=1.765 $X2=0 $Y2=0
cc_161 N_B2_c_127_n N_VPWR_c_732_n 0.00353822f $X=1.475 $Y=1.765 $X2=0 $Y2=0
cc_162 N_B2_c_128_n N_VPWR_c_732_n 0.00353905f $X=1.925 $Y=1.765 $X2=0 $Y2=0
cc_163 N_B2_M1007_g N_A_48_74#_c_833_n 0.00159319f $X=0.58 $Y=0.74 $X2=0 $Y2=0
cc_164 N_B2_M1007_g N_A_48_74#_c_834_n 0.0167076f $X=0.58 $Y=0.74 $X2=0 $Y2=0
cc_165 N_B2_M1013_g N_A_48_74#_c_834_n 0.01115f $X=1.01 $Y=0.74 $X2=0 $Y2=0
cc_166 N_B2_c_129_n N_A_48_74#_c_834_n 0.0342156f $X=1.79 $Y=1.515 $X2=0 $Y2=0
cc_167 N_B2_c_124_n N_A_48_74#_c_834_n 0.00238888f $X=1.87 $Y=1.557 $X2=0 $Y2=0
cc_168 N_B2_M1007_g N_A_48_74#_c_836_n 6.58468e-19 $X=0.58 $Y=0.74 $X2=0 $Y2=0
cc_169 N_B2_M1013_g N_A_48_74#_c_836_n 0.00918302f $X=1.01 $Y=0.74 $X2=0 $Y2=0
cc_170 N_B2_M1017_g N_A_48_74#_c_836_n 3.97481e-19 $X=1.44 $Y=0.74 $X2=0 $Y2=0
cc_171 N_B2_M1017_g N_A_48_74#_c_837_n 0.0130453f $X=1.44 $Y=0.74 $X2=0 $Y2=0
cc_172 N_B2_M1028_g N_A_48_74#_c_837_n 0.0128967f $X=1.87 $Y=0.74 $X2=0 $Y2=0
cc_173 N_B2_c_129_n N_A_48_74#_c_837_n 0.0483191f $X=1.79 $Y=1.515 $X2=0 $Y2=0
cc_174 N_B2_c_124_n N_A_48_74#_c_837_n 0.00503902f $X=1.87 $Y=1.557 $X2=0 $Y2=0
cc_175 N_B2_M1028_g N_A_48_74#_c_839_n 9.48753e-19 $X=1.87 $Y=0.74 $X2=0 $Y2=0
cc_176 N_B2_M1013_g N_A_48_74#_c_841_n 0.00157732f $X=1.01 $Y=0.74 $X2=0 $Y2=0
cc_177 N_B2_c_129_n N_A_48_74#_c_841_n 0.0213626f $X=1.79 $Y=1.515 $X2=0 $Y2=0
cc_178 N_B2_c_124_n N_A_48_74#_c_841_n 0.00232957f $X=1.87 $Y=1.557 $X2=0 $Y2=0
cc_179 N_B2_M1007_g N_VGND_c_899_n 0.0128874f $X=0.58 $Y=0.74 $X2=0 $Y2=0
cc_180 N_B2_M1013_g N_VGND_c_899_n 0.00204878f $X=1.01 $Y=0.74 $X2=0 $Y2=0
cc_181 N_B2_M1013_g N_VGND_c_900_n 5.19194e-19 $X=1.01 $Y=0.74 $X2=0 $Y2=0
cc_182 N_B2_M1017_g N_VGND_c_900_n 0.0108127f $X=1.44 $Y=0.74 $X2=0 $Y2=0
cc_183 N_B2_M1028_g N_VGND_c_900_n 0.0100301f $X=1.87 $Y=0.74 $X2=0 $Y2=0
cc_184 N_B2_M1028_g N_VGND_c_903_n 0.00383152f $X=1.87 $Y=0.74 $X2=0 $Y2=0
cc_185 N_B2_M1007_g N_VGND_c_907_n 0.00383152f $X=0.58 $Y=0.74 $X2=0 $Y2=0
cc_186 N_B2_M1013_g N_VGND_c_908_n 0.00434272f $X=1.01 $Y=0.74 $X2=0 $Y2=0
cc_187 N_B2_M1017_g N_VGND_c_908_n 0.00383152f $X=1.44 $Y=0.74 $X2=0 $Y2=0
cc_188 N_B2_M1007_g N_VGND_c_910_n 0.00761455f $X=0.58 $Y=0.74 $X2=0 $Y2=0
cc_189 N_B2_M1013_g N_VGND_c_910_n 0.00820284f $X=1.01 $Y=0.74 $X2=0 $Y2=0
cc_190 N_B2_M1017_g N_VGND_c_910_n 0.0075754f $X=1.44 $Y=0.74 $X2=0 $Y2=0
cc_191 N_B2_M1028_g N_VGND_c_910_n 0.00757637f $X=1.87 $Y=0.74 $X2=0 $Y2=0
cc_192 N_B1_c_212_n N_A1_c_308_n 0.00968263f $X=3.725 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_193 N_B1_c_208_n N_A1_M1012_g 0.0020658f $X=3.59 $Y=1.542 $X2=0 $Y2=0
cc_194 N_B1_c_208_n N_A1_c_305_n 0.0138384f $X=3.59 $Y=1.542 $X2=0 $Y2=0
cc_195 N_B1_c_208_n A1 8.7484e-19 $X=3.59 $Y=1.542 $X2=0 $Y2=0
cc_196 N_B1_c_209_n N_A_45_368#_c_492_n 0.00828741f $X=2.375 $Y=1.765 $X2=0
+ $Y2=0
cc_197 N_B1_c_210_n N_A_45_368#_c_492_n 5.7112e-19 $X=2.825 $Y=1.765 $X2=0 $Y2=0
cc_198 N_B1_c_209_n N_A_45_368#_c_472_n 0.0108414f $X=2.375 $Y=1.765 $X2=0 $Y2=0
cc_199 N_B1_c_210_n N_A_45_368#_c_472_n 0.0108414f $X=2.825 $Y=1.765 $X2=0 $Y2=0
cc_200 N_B1_c_209_n N_A_45_368#_c_501_n 5.7112e-19 $X=2.375 $Y=1.765 $X2=0 $Y2=0
cc_201 N_B1_c_210_n N_A_45_368#_c_501_n 0.00830261f $X=2.825 $Y=1.765 $X2=0
+ $Y2=0
cc_202 N_B1_c_211_n N_A_45_368#_c_501_n 0.00830261f $X=3.275 $Y=1.765 $X2=0
+ $Y2=0
cc_203 N_B1_c_212_n N_A_45_368#_c_501_n 5.7112e-19 $X=3.725 $Y=1.765 $X2=0 $Y2=0
cc_204 N_B1_c_211_n N_A_45_368#_c_473_n 0.0107904f $X=3.275 $Y=1.765 $X2=0 $Y2=0
cc_205 N_B1_c_212_n N_A_45_368#_c_473_n 0.0122595f $X=3.725 $Y=1.765 $X2=0 $Y2=0
cc_206 N_B1_c_212_n N_A_45_368#_c_474_n 0.00331158f $X=3.725 $Y=1.765 $X2=0
+ $Y2=0
cc_207 N_B1_c_208_n N_A_45_368#_c_474_n 4.64745e-19 $X=3.59 $Y=1.542 $X2=0 $Y2=0
cc_208 N_B1_c_211_n N_A_45_368#_c_509_n 5.98281e-19 $X=3.275 $Y=1.765 $X2=0
+ $Y2=0
cc_209 N_B1_c_212_n N_A_45_368#_c_509_n 0.00925416f $X=3.725 $Y=1.765 $X2=0
+ $Y2=0
cc_210 N_B1_c_209_n N_A_45_368#_c_481_n 0.00171731f $X=2.375 $Y=1.765 $X2=0
+ $Y2=0
cc_211 N_B1_c_210_n N_A_45_368#_c_482_n 0.00175197f $X=2.825 $Y=1.765 $X2=0
+ $Y2=0
cc_212 N_B1_c_211_n N_A_45_368#_c_482_n 0.00175197f $X=3.275 $Y=1.765 $X2=0
+ $Y2=0
cc_213 N_B1_c_209_n N_Y_c_635_n 0.0126342f $X=2.375 $Y=1.765 $X2=0 $Y2=0
cc_214 B1 N_Y_c_635_n 0.0154983f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_215 N_B1_c_208_n N_Y_c_635_n 0.0011179f $X=3.59 $Y=1.542 $X2=0 $Y2=0
cc_216 N_B1_M1004_g N_Y_c_642_n 0.00525476f $X=2.3 $Y=0.74 $X2=0 $Y2=0
cc_217 N_B1_M1006_g N_Y_c_642_n 0.00642147f $X=2.73 $Y=0.74 $X2=0 $Y2=0
cc_218 N_B1_M1023_g N_Y_c_642_n 5.71377e-19 $X=3.16 $Y=0.74 $X2=0 $Y2=0
cc_219 N_B1_c_209_n N_Y_c_645_n 0.00532448f $X=2.375 $Y=1.765 $X2=0 $Y2=0
cc_220 N_B1_c_210_n N_Y_c_645_n 0.00532448f $X=2.825 $Y=1.765 $X2=0 $Y2=0
cc_221 N_B1_M1006_g N_Y_c_618_n 0.00900535f $X=2.73 $Y=0.74 $X2=0 $Y2=0
cc_222 N_B1_M1023_g N_Y_c_618_n 0.00841735f $X=3.16 $Y=0.74 $X2=0 $Y2=0
cc_223 B1 N_Y_c_618_n 0.0396537f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_224 N_B1_c_208_n N_Y_c_618_n 0.00239847f $X=3.59 $Y=1.542 $X2=0 $Y2=0
cc_225 N_B1_M1004_g N_Y_c_619_n 0.00413664f $X=2.3 $Y=0.74 $X2=0 $Y2=0
cc_226 N_B1_M1006_g N_Y_c_619_n 0.00277633f $X=2.73 $Y=0.74 $X2=0 $Y2=0
cc_227 B1 N_Y_c_619_n 0.027784f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_228 N_B1_c_208_n N_Y_c_619_n 0.00244236f $X=3.59 $Y=1.542 $X2=0 $Y2=0
cc_229 N_B1_c_210_n N_Y_c_655_n 0.0126342f $X=2.825 $Y=1.765 $X2=0 $Y2=0
cc_230 N_B1_c_211_n N_Y_c_655_n 0.0149075f $X=3.275 $Y=1.765 $X2=0 $Y2=0
cc_231 B1 N_Y_c_655_n 0.039209f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_232 N_B1_c_208_n N_Y_c_655_n 0.00253386f $X=3.59 $Y=1.542 $X2=0 $Y2=0
cc_233 N_B1_c_211_n N_Y_c_623_n 0.00386833f $X=3.275 $Y=1.765 $X2=0 $Y2=0
cc_234 N_B1_c_212_n N_Y_c_623_n 0.00187771f $X=3.725 $Y=1.765 $X2=0 $Y2=0
cc_235 B1 N_Y_c_623_n 0.0200227f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_236 N_B1_c_208_n N_Y_c_623_n 0.014168f $X=3.59 $Y=1.542 $X2=0 $Y2=0
cc_237 N_B1_M1006_g N_Y_c_620_n 5.1907e-19 $X=2.73 $Y=0.74 $X2=0 $Y2=0
cc_238 N_B1_M1023_g N_Y_c_620_n 0.0093565f $X=3.16 $Y=0.74 $X2=0 $Y2=0
cc_239 N_B1_M1024_g N_Y_c_620_n 0.0241822f $X=3.59 $Y=0.74 $X2=0 $Y2=0
cc_240 B1 N_Y_c_620_n 0.0195623f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_241 N_B1_c_208_n N_Y_c_620_n 0.0314039f $X=3.59 $Y=1.542 $X2=0 $Y2=0
cc_242 B1 N_Y_c_668_n 0.0150275f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_243 N_B1_c_208_n N_Y_c_668_n 0.00103903f $X=3.59 $Y=1.542 $X2=0 $Y2=0
cc_244 N_B1_c_211_n N_Y_c_670_n 0.00515316f $X=3.275 $Y=1.765 $X2=0 $Y2=0
cc_245 N_B1_c_208_n N_Y_c_670_n 0.00127229f $X=3.59 $Y=1.542 $X2=0 $Y2=0
cc_246 N_B1_c_212_n N_VPWR_c_733_n 3.85248e-19 $X=3.725 $Y=1.765 $X2=0 $Y2=0
cc_247 N_B1_c_209_n N_VPWR_c_737_n 0.00278257f $X=2.375 $Y=1.765 $X2=0 $Y2=0
cc_248 N_B1_c_210_n N_VPWR_c_737_n 0.00278257f $X=2.825 $Y=1.765 $X2=0 $Y2=0
cc_249 N_B1_c_211_n N_VPWR_c_737_n 0.00278257f $X=3.275 $Y=1.765 $X2=0 $Y2=0
cc_250 N_B1_c_212_n N_VPWR_c_737_n 0.00278257f $X=3.725 $Y=1.765 $X2=0 $Y2=0
cc_251 N_B1_c_209_n N_VPWR_c_732_n 0.00353905f $X=2.375 $Y=1.765 $X2=0 $Y2=0
cc_252 N_B1_c_210_n N_VPWR_c_732_n 0.00353822f $X=2.825 $Y=1.765 $X2=0 $Y2=0
cc_253 N_B1_c_211_n N_VPWR_c_732_n 0.00353822f $X=3.275 $Y=1.765 $X2=0 $Y2=0
cc_254 N_B1_c_212_n N_VPWR_c_732_n 0.00353905f $X=3.725 $Y=1.765 $X2=0 $Y2=0
cc_255 N_B1_M1004_g N_A_48_74#_c_837_n 5.7448e-19 $X=2.3 $Y=0.74 $X2=0 $Y2=0
cc_256 N_B1_M1004_g N_A_48_74#_c_838_n 0.0119575f $X=2.3 $Y=0.74 $X2=0 $Y2=0
cc_257 N_B1_M1006_g N_A_48_74#_c_838_n 0.00942802f $X=2.73 $Y=0.74 $X2=0 $Y2=0
cc_258 N_B1_M1023_g N_A_48_74#_c_840_n 0.0135458f $X=3.16 $Y=0.74 $X2=0 $Y2=0
cc_259 N_B1_M1024_g N_A_48_74#_c_840_n 0.013953f $X=3.59 $Y=0.74 $X2=0 $Y2=0
cc_260 N_B1_M1006_g N_A_48_74#_c_842_n 2.84754e-19 $X=2.73 $Y=0.74 $X2=0 $Y2=0
cc_261 N_B1_M1023_g N_A_48_74#_c_842_n 2.84754e-19 $X=3.16 $Y=0.74 $X2=0 $Y2=0
cc_262 N_B1_M1004_g N_VGND_c_903_n 0.00278271f $X=2.3 $Y=0.74 $X2=0 $Y2=0
cc_263 N_B1_M1006_g N_VGND_c_903_n 0.00278271f $X=2.73 $Y=0.74 $X2=0 $Y2=0
cc_264 N_B1_M1023_g N_VGND_c_903_n 0.00278271f $X=3.16 $Y=0.74 $X2=0 $Y2=0
cc_265 N_B1_M1024_g N_VGND_c_903_n 0.00278271f $X=3.59 $Y=0.74 $X2=0 $Y2=0
cc_266 N_B1_M1004_g N_VGND_c_910_n 0.00353526f $X=2.3 $Y=0.74 $X2=0 $Y2=0
cc_267 N_B1_M1006_g N_VGND_c_910_n 0.00353428f $X=2.73 $Y=0.74 $X2=0 $Y2=0
cc_268 N_B1_M1023_g N_VGND_c_910_n 0.00353428f $X=3.16 $Y=0.74 $X2=0 $Y2=0
cc_269 N_B1_M1024_g N_VGND_c_910_n 0.00358427f $X=3.59 $Y=0.74 $X2=0 $Y2=0
cc_270 N_B1_M1024_g N_A_840_74#_c_1000_n 5.02354e-19 $X=3.59 $Y=0.74 $X2=0 $Y2=0
cc_271 N_A1_c_311_n N_A2_c_396_n 0.00978533f $X=5.755 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_272 N_A1_M1030_g N_A2_M1014_g 0.019323f $X=5.83 $Y=0.74 $X2=0 $Y2=0
cc_273 A1 N_A2_c_394_n 0.0274602f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_274 N_A1_c_307_n N_A2_c_394_n 0.0116557f $X=5.755 $Y=1.557 $X2=0 $Y2=0
cc_275 N_A1_c_307_n N_A2_c_395_n 0.0252148f $X=5.755 $Y=1.557 $X2=0 $Y2=0
cc_276 N_A1_c_308_n N_A_45_368#_c_473_n 0.00125031f $X=4.175 $Y=1.765 $X2=0
+ $Y2=0
cc_277 N_A1_c_308_n N_A_45_368#_c_474_n 0.00285814f $X=4.175 $Y=1.765 $X2=0
+ $Y2=0
cc_278 N_A1_c_308_n N_A_45_368#_c_509_n 0.00592667f $X=4.175 $Y=1.765 $X2=0
+ $Y2=0
cc_279 N_A1_c_308_n N_A_45_368#_c_517_n 0.0150614f $X=4.175 $Y=1.765 $X2=0 $Y2=0
cc_280 N_A1_c_300_n N_A_45_368#_c_517_n 0.0050955f $X=4.465 $Y=1.575 $X2=0 $Y2=0
cc_281 N_A1_c_309_n N_A_45_368#_c_517_n 0.0126853f $X=4.625 $Y=1.765 $X2=0 $Y2=0
cc_282 A1 N_A_45_368#_c_517_n 0.0202749f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_283 N_A1_c_309_n N_A_45_368#_c_475_n 0.00610108f $X=4.625 $Y=1.765 $X2=0
+ $Y2=0
cc_284 N_A1_c_310_n N_A_45_368#_c_475_n 0.0106335f $X=5.075 $Y=1.765 $X2=0 $Y2=0
cc_285 N_A1_c_311_n N_A_45_368#_c_475_n 8.2412e-19 $X=5.755 $Y=1.765 $X2=0 $Y2=0
cc_286 N_A1_c_310_n N_A_45_368#_c_524_n 0.0130095f $X=5.075 $Y=1.765 $X2=0 $Y2=0
cc_287 N_A1_c_311_n N_A_45_368#_c_524_n 0.017102f $X=5.755 $Y=1.765 $X2=0 $Y2=0
cc_288 A1 N_A_45_368#_c_524_n 0.0459409f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_289 N_A1_c_307_n N_A_45_368#_c_524_n 0.00244209f $X=5.755 $Y=1.557 $X2=0
+ $Y2=0
cc_290 N_A1_c_310_n N_A_45_368#_c_476_n 8.2412e-19 $X=5.075 $Y=1.765 $X2=0 $Y2=0
cc_291 N_A1_c_311_n N_A_45_368#_c_476_n 0.0109276f $X=5.755 $Y=1.765 $X2=0 $Y2=0
cc_292 N_A1_c_310_n N_A_45_368#_c_530_n 4.27055e-19 $X=5.075 $Y=1.765 $X2=0
+ $Y2=0
cc_293 A1 N_A_45_368#_c_530_n 0.0193936f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_294 N_A1_c_307_n N_A_45_368#_c_530_n 0.00123805f $X=5.755 $Y=1.557 $X2=0
+ $Y2=0
cc_295 N_A1_c_311_n N_A_45_368#_c_533_n 9.50925e-19 $X=5.755 $Y=1.765 $X2=0
+ $Y2=0
cc_296 N_A1_c_305_n N_Y_c_623_n 7.94101e-19 $X=4.175 $Y=1.575 $X2=0 $Y2=0
cc_297 N_A1_M1012_g N_Y_c_620_n 0.0102495f $X=4.54 $Y=0.74 $X2=0 $Y2=0
cc_298 N_A1_c_305_n N_Y_c_620_n 0.00595089f $X=4.175 $Y=1.575 $X2=0 $Y2=0
cc_299 A1 N_Y_c_620_n 0.0118787f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_300 N_A1_c_307_n N_Y_c_620_n 7.30532e-19 $X=5.755 $Y=1.557 $X2=0 $Y2=0
cc_301 N_A1_M1019_g N_Y_c_621_n 3.85913e-19 $X=4.97 $Y=0.74 $X2=0 $Y2=0
cc_302 N_A1_M1026_g N_Y_c_621_n 0.00304036f $X=5.4 $Y=0.74 $X2=0 $Y2=0
cc_303 N_A1_M1030_g N_Y_c_621_n 0.0054657f $X=5.83 $Y=0.74 $X2=0 $Y2=0
cc_304 N_A1_c_307_n N_Y_c_621_n 0.00271214f $X=5.755 $Y=1.557 $X2=0 $Y2=0
cc_305 N_A1_M1012_g N_Y_c_622_n 0.0156902f $X=4.54 $Y=0.74 $X2=0 $Y2=0
cc_306 N_A1_M1019_g N_Y_c_622_n 0.0123927f $X=4.97 $Y=0.74 $X2=0 $Y2=0
cc_307 N_A1_M1026_g N_Y_c_622_n 0.0106768f $X=5.4 $Y=0.74 $X2=0 $Y2=0
cc_308 N_A1_c_305_n N_Y_c_622_n 0.00767097f $X=4.175 $Y=1.575 $X2=0 $Y2=0
cc_309 A1 N_Y_c_622_n 0.0766192f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_310 N_A1_c_307_n N_Y_c_622_n 0.00448048f $X=5.755 $Y=1.557 $X2=0 $Y2=0
cc_311 N_A1_c_308_n N_VPWR_c_733_n 0.011002f $X=4.175 $Y=1.765 $X2=0 $Y2=0
cc_312 N_A1_c_309_n N_VPWR_c_733_n 0.011748f $X=4.625 $Y=1.765 $X2=0 $Y2=0
cc_313 N_A1_c_310_n N_VPWR_c_733_n 5.5582e-19 $X=5.075 $Y=1.765 $X2=0 $Y2=0
cc_314 N_A1_c_310_n N_VPWR_c_734_n 0.00722304f $X=5.075 $Y=1.765 $X2=0 $Y2=0
cc_315 N_A1_c_311_n N_VPWR_c_734_n 0.00722304f $X=5.755 $Y=1.765 $X2=0 $Y2=0
cc_316 N_A1_c_311_n N_VPWR_c_735_n 5.51351e-19 $X=5.755 $Y=1.765 $X2=0 $Y2=0
cc_317 N_A1_c_308_n N_VPWR_c_737_n 0.00413917f $X=4.175 $Y=1.765 $X2=0 $Y2=0
cc_318 N_A1_c_309_n N_VPWR_c_741_n 0.00413917f $X=4.625 $Y=1.765 $X2=0 $Y2=0
cc_319 N_A1_c_310_n N_VPWR_c_741_n 0.00445602f $X=5.075 $Y=1.765 $X2=0 $Y2=0
cc_320 N_A1_c_311_n N_VPWR_c_742_n 0.00445602f $X=5.755 $Y=1.765 $X2=0 $Y2=0
cc_321 N_A1_c_308_n N_VPWR_c_732_n 0.0081781f $X=4.175 $Y=1.765 $X2=0 $Y2=0
cc_322 N_A1_c_309_n N_VPWR_c_732_n 0.00817726f $X=4.625 $Y=1.765 $X2=0 $Y2=0
cc_323 N_A1_c_310_n N_VPWR_c_732_n 0.00858715f $X=5.075 $Y=1.765 $X2=0 $Y2=0
cc_324 N_A1_c_311_n N_VPWR_c_732_n 0.00858799f $X=5.755 $Y=1.765 $X2=0 $Y2=0
cc_325 N_A1_M1012_g N_A_48_74#_c_840_n 0.0032792f $X=4.54 $Y=0.74 $X2=0 $Y2=0
cc_326 N_A1_M1030_g N_VGND_c_901_n 6.37019e-19 $X=5.83 $Y=0.74 $X2=0 $Y2=0
cc_327 N_A1_M1012_g N_VGND_c_903_n 0.00291649f $X=4.54 $Y=0.74 $X2=0 $Y2=0
cc_328 N_A1_M1019_g N_VGND_c_903_n 0.00291649f $X=4.97 $Y=0.74 $X2=0 $Y2=0
cc_329 N_A1_M1026_g N_VGND_c_903_n 0.00291649f $X=5.4 $Y=0.74 $X2=0 $Y2=0
cc_330 N_A1_M1030_g N_VGND_c_903_n 0.00291649f $X=5.83 $Y=0.74 $X2=0 $Y2=0
cc_331 N_A1_M1012_g N_VGND_c_910_n 0.0036412f $X=4.54 $Y=0.74 $X2=0 $Y2=0
cc_332 N_A1_M1019_g N_VGND_c_910_n 0.00359121f $X=4.97 $Y=0.74 $X2=0 $Y2=0
cc_333 N_A1_M1026_g N_VGND_c_910_n 0.00359121f $X=5.4 $Y=0.74 $X2=0 $Y2=0
cc_334 N_A1_M1030_g N_VGND_c_910_n 0.00359219f $X=5.83 $Y=0.74 $X2=0 $Y2=0
cc_335 N_A1_M1012_g N_A_840_74#_c_993_n 0.00920696f $X=4.54 $Y=0.74 $X2=0 $Y2=0
cc_336 N_A1_M1019_g N_A_840_74#_c_993_n 0.0106927f $X=4.97 $Y=0.74 $X2=0 $Y2=0
cc_337 N_A1_M1026_g N_A_840_74#_c_993_n 0.0105443f $X=5.4 $Y=0.74 $X2=0 $Y2=0
cc_338 N_A1_M1030_g N_A_840_74#_c_993_n 0.014175f $X=5.83 $Y=0.74 $X2=0 $Y2=0
cc_339 N_A1_M1030_g N_A_840_74#_c_996_n 0.0017668f $X=5.83 $Y=0.74 $X2=0 $Y2=0
cc_340 N_A1_M1012_g N_A_840_74#_c_1000_n 0.00296395f $X=4.54 $Y=0.74 $X2=0 $Y2=0
cc_341 N_A1_M1019_g N_A_840_74#_c_1000_n 3.85913e-19 $X=4.97 $Y=0.74 $X2=0 $Y2=0
cc_342 N_A2_c_396_n N_A_45_368#_c_476_n 0.00623248f $X=6.205 $Y=1.765 $X2=0
+ $Y2=0
cc_343 N_A2_c_396_n N_A_45_368#_c_535_n 0.0126853f $X=6.205 $Y=1.765 $X2=0 $Y2=0
cc_344 N_A2_c_397_n N_A_45_368#_c_535_n 0.0126853f $X=6.655 $Y=1.765 $X2=0 $Y2=0
cc_345 N_A2_c_394_n N_A_45_368#_c_535_n 0.0477183f $X=7.3 $Y=1.515 $X2=0 $Y2=0
cc_346 N_A2_c_395_n N_A_45_368#_c_535_n 0.00150005f $X=7.55 $Y=1.557 $X2=0 $Y2=0
cc_347 N_A2_c_397_n N_A_45_368#_c_477_n 0.00572499f $X=6.655 $Y=1.765 $X2=0
+ $Y2=0
cc_348 N_A2_c_398_n N_A_45_368#_c_477_n 0.00572499f $X=7.105 $Y=1.765 $X2=0
+ $Y2=0
cc_349 N_A2_c_398_n N_A_45_368#_c_541_n 0.0126853f $X=7.105 $Y=1.765 $X2=0 $Y2=0
cc_350 N_A2_c_399_n N_A_45_368#_c_541_n 0.017059f $X=7.555 $Y=1.765 $X2=0 $Y2=0
cc_351 N_A2_c_394_n N_A_45_368#_c_541_n 0.0330867f $X=7.3 $Y=1.515 $X2=0 $Y2=0
cc_352 N_A2_c_395_n N_A_45_368#_c_541_n 0.00150005f $X=7.55 $Y=1.557 $X2=0 $Y2=0
cc_353 N_A2_c_399_n N_A_45_368#_c_478_n 0.00314968f $X=7.555 $Y=1.765 $X2=0
+ $Y2=0
cc_354 N_A2_c_399_n N_A_45_368#_c_479_n 0.00729586f $X=7.555 $Y=1.765 $X2=0
+ $Y2=0
cc_355 N_A2_c_394_n N_A_45_368#_c_533_n 0.0158218f $X=7.3 $Y=1.515 $X2=0 $Y2=0
cc_356 N_A2_c_394_n N_A_45_368#_c_548_n 0.0150275f $X=7.3 $Y=1.515 $X2=0 $Y2=0
cc_357 N_A2_c_395_n N_A_45_368#_c_548_n 0.00104296f $X=7.55 $Y=1.557 $X2=0 $Y2=0
cc_358 N_A2_c_396_n N_VPWR_c_735_n 0.011748f $X=6.205 $Y=1.765 $X2=0 $Y2=0
cc_359 N_A2_c_397_n N_VPWR_c_735_n 0.0116643f $X=6.655 $Y=1.765 $X2=0 $Y2=0
cc_360 N_A2_c_398_n N_VPWR_c_735_n 5.35985e-19 $X=7.105 $Y=1.765 $X2=0 $Y2=0
cc_361 N_A2_c_397_n N_VPWR_c_736_n 5.35985e-19 $X=6.655 $Y=1.765 $X2=0 $Y2=0
cc_362 N_A2_c_398_n N_VPWR_c_736_n 0.0116643f $X=7.105 $Y=1.765 $X2=0 $Y2=0
cc_363 N_A2_c_399_n N_VPWR_c_736_n 0.0147395f $X=7.555 $Y=1.765 $X2=0 $Y2=0
cc_364 N_A2_c_397_n N_VPWR_c_739_n 0.00413917f $X=6.655 $Y=1.765 $X2=0 $Y2=0
cc_365 N_A2_c_398_n N_VPWR_c_739_n 0.00413917f $X=7.105 $Y=1.765 $X2=0 $Y2=0
cc_366 N_A2_c_396_n N_VPWR_c_742_n 0.00413917f $X=6.205 $Y=1.765 $X2=0 $Y2=0
cc_367 N_A2_c_399_n N_VPWR_c_743_n 0.00413917f $X=7.555 $Y=1.765 $X2=0 $Y2=0
cc_368 N_A2_c_396_n N_VPWR_c_732_n 0.0081781f $X=6.205 $Y=1.765 $X2=0 $Y2=0
cc_369 N_A2_c_397_n N_VPWR_c_732_n 0.00817726f $X=6.655 $Y=1.765 $X2=0 $Y2=0
cc_370 N_A2_c_398_n N_VPWR_c_732_n 0.00817726f $X=7.105 $Y=1.765 $X2=0 $Y2=0
cc_371 N_A2_c_399_n N_VPWR_c_732_n 0.00821508f $X=7.555 $Y=1.765 $X2=0 $Y2=0
cc_372 N_A2_M1014_g N_VGND_c_901_n 0.00977449f $X=6.26 $Y=0.74 $X2=0 $Y2=0
cc_373 N_A2_M1015_g N_VGND_c_901_n 0.00192252f $X=6.69 $Y=0.74 $X2=0 $Y2=0
cc_374 N_A2_M1015_g N_VGND_c_902_n 5.20618e-19 $X=6.69 $Y=0.74 $X2=0 $Y2=0
cc_375 N_A2_M1018_g N_VGND_c_902_n 0.00985915f $X=7.12 $Y=0.74 $X2=0 $Y2=0
cc_376 N_A2_M1029_g N_VGND_c_902_n 0.00328502f $X=7.55 $Y=0.74 $X2=0 $Y2=0
cc_377 N_A2_M1014_g N_VGND_c_903_n 0.00383152f $X=6.26 $Y=0.74 $X2=0 $Y2=0
cc_378 N_A2_M1015_g N_VGND_c_905_n 0.00434272f $X=6.69 $Y=0.74 $X2=0 $Y2=0
cc_379 N_A2_M1018_g N_VGND_c_905_n 0.00383152f $X=7.12 $Y=0.74 $X2=0 $Y2=0
cc_380 N_A2_M1029_g N_VGND_c_909_n 0.00434272f $X=7.55 $Y=0.74 $X2=0 $Y2=0
cc_381 N_A2_M1014_g N_VGND_c_910_n 0.00757637f $X=6.26 $Y=0.74 $X2=0 $Y2=0
cc_382 N_A2_M1015_g N_VGND_c_910_n 0.00820284f $X=6.69 $Y=0.74 $X2=0 $Y2=0
cc_383 N_A2_M1018_g N_VGND_c_910_n 0.0075754f $X=7.12 $Y=0.74 $X2=0 $Y2=0
cc_384 N_A2_M1029_g N_VGND_c_910_n 0.00824275f $X=7.55 $Y=0.74 $X2=0 $Y2=0
cc_385 N_A2_M1014_g N_A_840_74#_c_995_n 0.0128967f $X=6.26 $Y=0.74 $X2=0 $Y2=0
cc_386 N_A2_M1015_g N_A_840_74#_c_995_n 0.0111034f $X=6.69 $Y=0.74 $X2=0 $Y2=0
cc_387 N_A2_c_394_n N_A_840_74#_c_995_n 0.0456932f $X=7.3 $Y=1.515 $X2=0 $Y2=0
cc_388 N_A2_c_395_n N_A_840_74#_c_995_n 0.00368969f $X=7.55 $Y=1.557 $X2=0 $Y2=0
cc_389 N_A2_c_394_n N_A_840_74#_c_996_n 0.0152645f $X=7.3 $Y=1.515 $X2=0 $Y2=0
cc_390 N_A2_c_395_n N_A_840_74#_c_996_n 3.65737e-19 $X=7.55 $Y=1.557 $X2=0 $Y2=0
cc_391 N_A2_M1014_g N_A_840_74#_c_997_n 7.09663e-19 $X=6.26 $Y=0.74 $X2=0 $Y2=0
cc_392 N_A2_M1015_g N_A_840_74#_c_997_n 0.00918302f $X=6.69 $Y=0.74 $X2=0 $Y2=0
cc_393 N_A2_M1018_g N_A_840_74#_c_997_n 3.97481e-19 $X=7.12 $Y=0.74 $X2=0 $Y2=0
cc_394 N_A2_M1018_g N_A_840_74#_c_998_n 0.0130918f $X=7.12 $Y=0.74 $X2=0 $Y2=0
cc_395 N_A2_M1029_g N_A_840_74#_c_998_n 0.0180105f $X=7.55 $Y=0.74 $X2=0 $Y2=0
cc_396 N_A2_c_394_n N_A_840_74#_c_998_n 0.0358403f $X=7.3 $Y=1.515 $X2=0 $Y2=0
cc_397 N_A2_c_395_n N_A_840_74#_c_998_n 0.0031669f $X=7.55 $Y=1.557 $X2=0 $Y2=0
cc_398 N_A2_M1018_g N_A_840_74#_c_999_n 7.07591e-19 $X=7.12 $Y=0.74 $X2=0 $Y2=0
cc_399 N_A2_M1029_g N_A_840_74#_c_999_n 0.0100626f $X=7.55 $Y=0.74 $X2=0 $Y2=0
cc_400 N_A2_M1015_g N_A_840_74#_c_1001_n 0.00157732f $X=6.69 $Y=0.74 $X2=0 $Y2=0
cc_401 N_A2_c_394_n N_A_840_74#_c_1001_n 0.0213626f $X=7.3 $Y=1.515 $X2=0 $Y2=0
cc_402 N_A2_c_395_n N_A_840_74#_c_1001_n 0.00232957f $X=7.55 $Y=1.557 $X2=0
+ $Y2=0
cc_403 N_A_45_368#_c_469_n N_Y_M1005_s 0.00222494f $X=1.085 $Y=2.99 $X2=0 $Y2=0
cc_404 N_A_45_368#_c_471_n N_Y_M1011_s 0.00247267f $X=1.985 $Y=2.99 $X2=0 $Y2=0
cc_405 N_A_45_368#_c_472_n N_Y_M1000_s 0.00247267f $X=2.885 $Y=2.99 $X2=0 $Y2=0
cc_406 N_A_45_368#_c_473_n N_Y_M1016_s 0.00222494f $X=3.785 $Y=2.99 $X2=0 $Y2=0
cc_407 N_A_45_368#_c_468_n N_Y_c_624_n 0.0121024f $X=0.35 $Y=1.985 $X2=0 $Y2=0
cc_408 N_A_45_368#_c_468_n N_Y_c_627_n 0.0403609f $X=0.35 $Y=1.985 $X2=0 $Y2=0
cc_409 N_A_45_368#_c_469_n N_Y_c_627_n 0.0144323f $X=1.085 $Y=2.99 $X2=0 $Y2=0
cc_410 N_A_45_368#_c_486_n N_Y_c_627_n 0.0298377f $X=1.25 $Y=2.375 $X2=0 $Y2=0
cc_411 N_A_45_368#_M1010_d N_Y_c_629_n 0.00359365f $X=1.1 $Y=1.84 $X2=0 $Y2=0
cc_412 N_A_45_368#_c_486_n N_Y_c_629_n 0.0171813f $X=1.25 $Y=2.375 $X2=0 $Y2=0
cc_413 N_A_45_368#_c_486_n N_Y_c_633_n 0.0289859f $X=1.25 $Y=2.375 $X2=0 $Y2=0
cc_414 N_A_45_368#_c_471_n N_Y_c_633_n 0.012787f $X=1.985 $Y=2.99 $X2=0 $Y2=0
cc_415 N_A_45_368#_c_492_n N_Y_c_633_n 0.0289859f $X=2.15 $Y=2.375 $X2=0 $Y2=0
cc_416 N_A_45_368#_M1020_d N_Y_c_635_n 0.00865978f $X=2 $Y=1.84 $X2=0 $Y2=0
cc_417 N_A_45_368#_c_492_n N_Y_c_635_n 0.0171814f $X=2.15 $Y=2.375 $X2=0 $Y2=0
cc_418 N_A_45_368#_c_492_n N_Y_c_645_n 0.0289859f $X=2.15 $Y=2.375 $X2=0 $Y2=0
cc_419 N_A_45_368#_c_472_n N_Y_c_645_n 0.012787f $X=2.885 $Y=2.99 $X2=0 $Y2=0
cc_420 N_A_45_368#_c_501_n N_Y_c_645_n 0.0289859f $X=3.05 $Y=2.375 $X2=0 $Y2=0
cc_421 N_A_45_368#_M1008_d N_Y_c_655_n 0.00359365f $X=2.9 $Y=1.84 $X2=0 $Y2=0
cc_422 N_A_45_368#_c_501_n N_Y_c_655_n 0.0171813f $X=3.05 $Y=2.375 $X2=0 $Y2=0
cc_423 N_A_45_368#_c_474_n N_Y_c_623_n 0.0054205f $X=3.91 $Y=2.12 $X2=0 $Y2=0
cc_424 N_A_45_368#_c_474_n N_Y_c_620_n 0.0155233f $X=3.91 $Y=2.12 $X2=0 $Y2=0
cc_425 N_A_45_368#_c_517_n N_Y_c_620_n 0.00503654f $X=4.765 $Y=2.035 $X2=0 $Y2=0
cc_426 N_A_45_368#_c_501_n N_Y_c_670_n 0.0293393f $X=3.05 $Y=2.375 $X2=0 $Y2=0
cc_427 N_A_45_368#_c_473_n N_Y_c_670_n 0.013472f $X=3.785 $Y=2.99 $X2=0 $Y2=0
cc_428 N_A_45_368#_c_517_n N_VPWR_M1001_d 0.0041741f $X=4.765 $Y=2.035 $X2=-0.19
+ $Y2=1.66
cc_429 N_A_45_368#_c_524_n N_VPWR_M1022_d 0.00961821f $X=5.815 $Y=2.035 $X2=0
+ $Y2=0
cc_430 N_A_45_368#_c_535_n N_VPWR_M1002_s 0.00359365f $X=6.795 $Y=2.035 $X2=0
+ $Y2=0
cc_431 N_A_45_368#_c_541_n N_VPWR_M1009_s 0.00359365f $X=7.695 $Y=2.035 $X2=0
+ $Y2=0
cc_432 N_A_45_368#_c_473_n N_VPWR_c_733_n 0.0125885f $X=3.785 $Y=2.99 $X2=0
+ $Y2=0
cc_433 N_A_45_368#_c_509_n N_VPWR_c_733_n 0.0412023f $X=3.95 $Y=2.4 $X2=0 $Y2=0
cc_434 N_A_45_368#_c_517_n N_VPWR_c_733_n 0.0171814f $X=4.765 $Y=2.035 $X2=0
+ $Y2=0
cc_435 N_A_45_368#_c_475_n N_VPWR_c_733_n 0.0462948f $X=4.85 $Y=2.415 $X2=0
+ $Y2=0
cc_436 N_A_45_368#_c_475_n N_VPWR_c_734_n 0.0256432f $X=4.85 $Y=2.415 $X2=0
+ $Y2=0
cc_437 N_A_45_368#_c_524_n N_VPWR_c_734_n 0.0338452f $X=5.815 $Y=2.035 $X2=0
+ $Y2=0
cc_438 N_A_45_368#_c_476_n N_VPWR_c_734_n 0.0256432f $X=5.98 $Y=2.465 $X2=0
+ $Y2=0
cc_439 N_A_45_368#_c_476_n N_VPWR_c_735_n 0.0462948f $X=5.98 $Y=2.465 $X2=0
+ $Y2=0
cc_440 N_A_45_368#_c_535_n N_VPWR_c_735_n 0.0171813f $X=6.795 $Y=2.035 $X2=0
+ $Y2=0
cc_441 N_A_45_368#_c_477_n N_VPWR_c_735_n 0.0449718f $X=6.88 $Y=2.465 $X2=0
+ $Y2=0
cc_442 N_A_45_368#_c_477_n N_VPWR_c_736_n 0.0449718f $X=6.88 $Y=2.465 $X2=0
+ $Y2=0
cc_443 N_A_45_368#_c_541_n N_VPWR_c_736_n 0.0171813f $X=7.695 $Y=2.035 $X2=0
+ $Y2=0
cc_444 N_A_45_368#_c_479_n N_VPWR_c_736_n 0.0462948f $X=7.78 $Y=2.4 $X2=0 $Y2=0
cc_445 N_A_45_368#_c_469_n N_VPWR_c_737_n 0.0409869f $X=1.085 $Y=2.99 $X2=0
+ $Y2=0
cc_446 N_A_45_368#_c_470_n N_VPWR_c_737_n 0.0179217f $X=0.435 $Y=2.99 $X2=0
+ $Y2=0
cc_447 N_A_45_368#_c_471_n N_VPWR_c_737_n 0.03588f $X=1.985 $Y=2.99 $X2=0 $Y2=0
cc_448 N_A_45_368#_c_472_n N_VPWR_c_737_n 0.03588f $X=2.885 $Y=2.99 $X2=0 $Y2=0
cc_449 N_A_45_368#_c_473_n N_VPWR_c_737_n 0.053749f $X=3.785 $Y=2.99 $X2=0 $Y2=0
cc_450 N_A_45_368#_c_480_n N_VPWR_c_737_n 0.0235512f $X=1.25 $Y=2.99 $X2=0 $Y2=0
cc_451 N_A_45_368#_c_481_n N_VPWR_c_737_n 0.0235512f $X=2.15 $Y=2.99 $X2=0 $Y2=0
cc_452 N_A_45_368#_c_482_n N_VPWR_c_737_n 0.0235512f $X=3.05 $Y=2.99 $X2=0 $Y2=0
cc_453 N_A_45_368#_c_477_n N_VPWR_c_739_n 0.00749631f $X=6.88 $Y=2.465 $X2=0
+ $Y2=0
cc_454 N_A_45_368#_c_475_n N_VPWR_c_741_n 0.0110241f $X=4.85 $Y=2.415 $X2=0
+ $Y2=0
cc_455 N_A_45_368#_c_476_n N_VPWR_c_742_n 0.0110241f $X=5.98 $Y=2.465 $X2=0
+ $Y2=0
cc_456 N_A_45_368#_c_479_n N_VPWR_c_743_n 0.011066f $X=7.78 $Y=2.4 $X2=0 $Y2=0
cc_457 N_A_45_368#_c_469_n N_VPWR_c_732_n 0.0231342f $X=1.085 $Y=2.99 $X2=0
+ $Y2=0
cc_458 N_A_45_368#_c_470_n N_VPWR_c_732_n 0.00971942f $X=0.435 $Y=2.99 $X2=0
+ $Y2=0
cc_459 N_A_45_368#_c_471_n N_VPWR_c_732_n 0.0201952f $X=1.985 $Y=2.99 $X2=0
+ $Y2=0
cc_460 N_A_45_368#_c_472_n N_VPWR_c_732_n 0.0201952f $X=2.885 $Y=2.99 $X2=0
+ $Y2=0
cc_461 N_A_45_368#_c_473_n N_VPWR_c_732_n 0.029846f $X=3.785 $Y=2.99 $X2=0 $Y2=0
cc_462 N_A_45_368#_c_475_n N_VPWR_c_732_n 0.00909194f $X=4.85 $Y=2.415 $X2=0
+ $Y2=0
cc_463 N_A_45_368#_c_476_n N_VPWR_c_732_n 0.00909194f $X=5.98 $Y=2.465 $X2=0
+ $Y2=0
cc_464 N_A_45_368#_c_477_n N_VPWR_c_732_n 0.0062048f $X=6.88 $Y=2.465 $X2=0
+ $Y2=0
cc_465 N_A_45_368#_c_479_n N_VPWR_c_732_n 0.00915947f $X=7.78 $Y=2.4 $X2=0 $Y2=0
cc_466 N_A_45_368#_c_480_n N_VPWR_c_732_n 0.0126924f $X=1.25 $Y=2.99 $X2=0 $Y2=0
cc_467 N_A_45_368#_c_481_n N_VPWR_c_732_n 0.0126924f $X=2.15 $Y=2.99 $X2=0 $Y2=0
cc_468 N_A_45_368#_c_482_n N_VPWR_c_732_n 0.0126924f $X=3.05 $Y=2.99 $X2=0 $Y2=0
cc_469 N_A_45_368#_c_468_n N_A_48_74#_c_835_n 0.00864987f $X=0.35 $Y=1.985 $X2=0
+ $Y2=0
cc_470 N_A_45_368#_c_478_n N_A_840_74#_c_998_n 0.00868683f $X=7.82 $Y=2.12 $X2=0
+ $Y2=0
cc_471 N_Y_c_618_n N_A_48_74#_M1006_d 0.00176461f $X=3.21 $Y=1.095 $X2=0 $Y2=0
cc_472 N_Y_c_620_n N_A_48_74#_M1024_d 0.00386132f $X=4.195 $Y=0.99 $X2=0 $Y2=0
cc_473 N_Y_c_619_n N_A_48_74#_c_837_n 0.00997012f $X=2.68 $Y=1.095 $X2=0 $Y2=0
cc_474 N_Y_M1004_s N_A_48_74#_c_838_n 0.00176461f $X=2.375 $Y=0.37 $X2=0 $Y2=0
cc_475 N_Y_c_642_n N_A_48_74#_c_838_n 0.0157965f $X=2.515 $Y=0.76 $X2=0 $Y2=0
cc_476 N_Y_c_618_n N_A_48_74#_c_838_n 0.0030313f $X=3.21 $Y=1.095 $X2=0 $Y2=0
cc_477 N_Y_M1023_s N_A_48_74#_c_840_n 0.00180346f $X=3.235 $Y=0.37 $X2=0 $Y2=0
cc_478 N_Y_c_618_n N_A_48_74#_c_840_n 0.00436902f $X=3.21 $Y=1.095 $X2=0 $Y2=0
cc_479 N_Y_c_620_n N_A_48_74#_c_840_n 0.0472031f $X=4.195 $Y=0.99 $X2=0 $Y2=0
cc_480 N_Y_c_618_n N_A_48_74#_c_842_n 0.0133411f $X=3.21 $Y=1.095 $X2=0 $Y2=0
cc_481 N_Y_c_620_n N_VGND_c_910_n 0.00898375f $X=4.195 $Y=0.99 $X2=0 $Y2=0
cc_482 N_Y_c_622_n N_A_840_74#_M1012_d 0.00344035f $X=5.45 $Y=0.95 $X2=-0.19
+ $Y2=-0.245
cc_483 N_Y_c_622_n N_A_840_74#_M1019_d 0.00209854f $X=5.45 $Y=0.95 $X2=0 $Y2=0
cc_484 N_Y_M1012_s N_A_840_74#_c_993_n 0.00212678f $X=4.615 $Y=0.37 $X2=0 $Y2=0
cc_485 N_Y_M1026_s N_A_840_74#_c_993_n 0.00179007f $X=5.475 $Y=0.37 $X2=0 $Y2=0
cc_486 N_Y_c_621_n N_A_840_74#_c_993_n 0.016201f $X=5.615 $Y=0.95 $X2=0 $Y2=0
cc_487 N_Y_c_622_n N_A_840_74#_c_993_n 0.0379865f $X=5.45 $Y=0.95 $X2=0 $Y2=0
cc_488 N_Y_c_621_n N_A_840_74#_c_996_n 0.00561736f $X=5.615 $Y=0.95 $X2=0 $Y2=0
cc_489 N_Y_c_620_n N_A_840_74#_c_1000_n 0.0030156f $X=4.195 $Y=0.99 $X2=0 $Y2=0
cc_490 N_Y_c_622_n N_A_840_74#_c_1000_n 0.0182263f $X=5.45 $Y=0.95 $X2=0 $Y2=0
cc_491 N_A_48_74#_c_834_n N_VGND_M1007_d 0.00176461f $X=1.06 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_492 N_A_48_74#_c_837_n N_VGND_M1017_d 0.00176461f $X=2 $Y=1.095 $X2=0 $Y2=0
cc_493 N_A_48_74#_c_833_n N_VGND_c_899_n 0.0175587f $X=0.365 $Y=0.515 $X2=0
+ $Y2=0
cc_494 N_A_48_74#_c_834_n N_VGND_c_899_n 0.0152916f $X=1.06 $Y=1.095 $X2=0 $Y2=0
cc_495 N_A_48_74#_c_836_n N_VGND_c_899_n 0.0175587f $X=1.225 $Y=0.515 $X2=0
+ $Y2=0
cc_496 N_A_48_74#_c_836_n N_VGND_c_900_n 0.0182902f $X=1.225 $Y=0.515 $X2=0
+ $Y2=0
cc_497 N_A_48_74#_c_837_n N_VGND_c_900_n 0.0170777f $X=2 $Y=1.095 $X2=0 $Y2=0
cc_498 N_A_48_74#_c_839_n N_VGND_c_900_n 0.0112234f $X=2.17 $Y=0.34 $X2=0 $Y2=0
cc_499 N_A_48_74#_c_838_n N_VGND_c_903_n 0.0435462f $X=2.86 $Y=0.34 $X2=0 $Y2=0
cc_500 N_A_48_74#_c_839_n N_VGND_c_903_n 0.0121867f $X=2.17 $Y=0.34 $X2=0 $Y2=0
cc_501 N_A_48_74#_c_840_n N_VGND_c_903_n 0.0626962f $X=3.805 $Y=0.515 $X2=0
+ $Y2=0
cc_502 N_A_48_74#_c_842_n N_VGND_c_903_n 0.0119073f $X=2.945 $Y=0.34 $X2=0 $Y2=0
cc_503 N_A_48_74#_c_833_n N_VGND_c_907_n 0.011066f $X=0.365 $Y=0.515 $X2=0 $Y2=0
cc_504 N_A_48_74#_c_836_n N_VGND_c_908_n 0.0109942f $X=1.225 $Y=0.515 $X2=0
+ $Y2=0
cc_505 N_A_48_74#_c_833_n N_VGND_c_910_n 0.00915947f $X=0.365 $Y=0.515 $X2=0
+ $Y2=0
cc_506 N_A_48_74#_c_836_n N_VGND_c_910_n 0.00904371f $X=1.225 $Y=0.515 $X2=0
+ $Y2=0
cc_507 N_A_48_74#_c_838_n N_VGND_c_910_n 0.0245733f $X=2.86 $Y=0.34 $X2=0 $Y2=0
cc_508 N_A_48_74#_c_839_n N_VGND_c_910_n 0.00660921f $X=2.17 $Y=0.34 $X2=0 $Y2=0
cc_509 N_A_48_74#_c_840_n N_VGND_c_910_n 0.0345365f $X=3.805 $Y=0.515 $X2=0
+ $Y2=0
cc_510 N_A_48_74#_c_842_n N_VGND_c_910_n 0.00650586f $X=2.945 $Y=0.34 $X2=0
+ $Y2=0
cc_511 N_A_48_74#_c_840_n N_A_840_74#_c_1000_n 0.0214676f $X=3.805 $Y=0.515
+ $X2=0 $Y2=0
cc_512 N_VGND_c_901_n N_A_840_74#_c_994_n 0.00947603f $X=6.475 $Y=0.595 $X2=0
+ $Y2=0
cc_513 N_VGND_c_903_n N_A_840_74#_c_994_n 0.00758556f $X=6.31 $Y=0 $X2=0 $Y2=0
cc_514 N_VGND_c_910_n N_A_840_74#_c_994_n 0.00627867f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_515 N_VGND_M1014_d N_A_840_74#_c_995_n 0.00176461f $X=6.335 $Y=0.37 $X2=0
+ $Y2=0
cc_516 N_VGND_c_901_n N_A_840_74#_c_995_n 0.0153337f $X=6.475 $Y=0.595 $X2=0
+ $Y2=0
cc_517 N_VGND_c_901_n N_A_840_74#_c_997_n 0.0175587f $X=6.475 $Y=0.595 $X2=0
+ $Y2=0
cc_518 N_VGND_c_902_n N_A_840_74#_c_997_n 0.0175587f $X=7.335 $Y=0.595 $X2=0
+ $Y2=0
cc_519 N_VGND_c_905_n N_A_840_74#_c_997_n 0.0109942f $X=7.17 $Y=0 $X2=0 $Y2=0
cc_520 N_VGND_c_910_n N_A_840_74#_c_997_n 0.00904371f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_521 N_VGND_M1018_d N_A_840_74#_c_998_n 0.00176461f $X=7.195 $Y=0.37 $X2=0
+ $Y2=0
cc_522 N_VGND_c_902_n N_A_840_74#_c_998_n 0.0153337f $X=7.335 $Y=0.595 $X2=0
+ $Y2=0
cc_523 N_VGND_c_902_n N_A_840_74#_c_999_n 0.0182902f $X=7.335 $Y=0.595 $X2=0
+ $Y2=0
cc_524 N_VGND_c_909_n N_A_840_74#_c_999_n 0.0145639f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_525 N_VGND_c_910_n N_A_840_74#_c_999_n 0.0119984f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_526 N_VGND_c_903_n N_A_840_74#_c_1000_n 0.0731929f $X=6.31 $Y=0 $X2=0 $Y2=0
cc_527 N_VGND_c_910_n N_A_840_74#_c_1000_n 0.0615691f $X=7.92 $Y=0 $X2=0 $Y2=0
