* NGSPICE file created from sky130_fd_sc_ls__fa_2.ext - technology: sky130A

.subckt sky130_fd_sc_ls__fa_2 A B CIN VGND VNB VPB VPWR COUT SUM
M1000 a_1205_79# B a_1119_79# VNB nshort w=740000u l=150000u
+  ad=1.776e+11p pd=1.96e+06u as=2.072e+11p ps=2.04e+06u
M1001 VGND A a_1205_79# VNB nshort w=740000u l=150000u
+  ad=2.36723e+12p pd=1.592e+07u as=0p ps=0u
M1002 COUT a_336_347# VGND VNB nshort w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1003 a_27_79# B VGND VNB nshort w=740000u l=150000u
+  ad=6.327e+11p pd=4.67e+06u as=0p ps=0u
M1004 SUM a_992_347# VGND VNB nshort w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1005 a_27_378# B VPWR VPB phighvt w=1e+06u l=150000u
+  ad=5.95e+11p pd=5.19e+06u as=2.80985e+12p ps=1.858e+07u
M1006 a_683_347# CIN VPWR VPB phighvt w=1e+06u l=150000u
+  ad=6.82125e+11p pd=5.62e+06u as=0p ps=0u
M1007 VPWR A a_27_378# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND a_336_347# COUT VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 COUT a_336_347# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=4.424e+11p pd=3.03e+06u as=0p ps=0u
M1010 VGND a_992_347# SUM VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND B a_701_79# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=5.18e+11p ps=4.36e+06u
M1012 a_336_347# CIN a_27_378# VPB phighvt w=1e+06u l=150000u
+  ad=5.9e+11p pd=3.18e+06u as=0p ps=0u
M1013 a_701_79# A VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 SUM a_992_347# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=0p ps=0u
M1015 VGND A a_27_79# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR A a_484_347# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1017 a_1119_79# CIN a_992_347# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.59e+11p ps=2.18e+06u
M1018 a_683_347# A VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND A a_487_79# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=1.776e+11p ps=1.96e+06u
M1020 VPWR A a_1202_368# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1021 a_487_79# B a_336_347# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.59e+11p ps=2.18e+06u
M1022 a_484_347# B a_336_347# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VPWR B a_683_347# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VPWR a_992_347# SUM VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_1094_347# CIN a_992_347# VPB phighvt w=1e+06u l=150000u
+  ad=4.047e+11p pd=2.99e+06u as=3.6e+11p ps=2.72e+06u
M1026 a_1202_368# B a_1094_347# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VPWR a_336_347# COUT VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_336_347# CIN a_27_79# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_701_79# CIN VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_992_347# a_336_347# a_683_347# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_992_347# a_336_347# a_701_79# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

