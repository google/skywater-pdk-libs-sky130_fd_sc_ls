* File: sky130_fd_sc_ls__nor4_4.spice
* Created: Fri Aug 28 13:40:06 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__nor4_4.pex.spice"
.subckt sky130_fd_sc_ls__nor4_4  VNB VPB D C B A Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A	A
* B	B
* C	C
* D	D
* VPB	VPB
* VNB	VNB
MM1002 N_VGND_M1002_d N_D_M1002_g N_Y_M1002_s VNB NSHORT L=0.15 W=0.74 AD=0.2442
+ AS=0.4329 PD=2.14 PS=1.91 NRD=7.296 NRS=0 M=1 R=4.93333 SA=75000.3 SB=75007.6
+ A=0.111 P=1.78 MULT=1
MM1020 N_VGND_M1020_d N_D_M1020_g N_Y_M1002_s VNB NSHORT L=0.15 W=0.74 AD=0.1295
+ AS=0.4329 PD=1.09 PS=1.91 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.6 SB=75006.3
+ A=0.111 P=1.78 MULT=1
MM1008 N_VGND_M1020_d N_C_M1008_g N_Y_M1008_s VNB NSHORT L=0.15 W=0.74 AD=0.1295
+ AS=0.444 PD=1.09 PS=1.94 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75002.1 SB=75005.8
+ A=0.111 P=1.78 MULT=1
MM1022 N_VGND_M1022_d N_C_M1022_g N_Y_M1008_s VNB NSHORT L=0.15 W=0.74 AD=0.1295
+ AS=0.444 PD=1.09 PS=1.94 NRD=0 NRS=0 M=1 R=4.93333 SA=75003.4 SB=75004.5
+ A=0.111 P=1.78 MULT=1
MM1007 N_Y_M1007_d N_B_M1007_g N_VGND_M1022_d VNB NSHORT L=0.15 W=0.74 AD=0.1036
+ AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75003.9 SB=75004
+ A=0.111 P=1.78 MULT=1
MM1015 N_Y_M1007_d N_B_M1015_g N_VGND_M1015_s VNB NSHORT L=0.15 W=0.74 AD=0.1036
+ AS=0.8621 PD=1.02 PS=3.07 NRD=0 NRS=0 M=1 R=4.93333 SA=75004.4 SB=75003.5
+ A=0.111 P=1.78 MULT=1
MM1010 N_Y_M1010_d N_A_M1010_g N_VGND_M1015_s VNB NSHORT L=0.15 W=0.74 AD=0.2627
+ AS=0.8621 PD=1.45 PS=3.07 NRD=48.648 NRS=0 M=1 R=4.93333 SA=75006.8 SB=75001.1
+ A=0.111 P=1.78 MULT=1
MM1017 N_Y_M1010_d N_A_M1017_g N_VGND_M1017_s VNB NSHORT L=0.15 W=0.74 AD=0.2627
+ AS=0.2109 PD=1.45 PS=2.05 NRD=48.648 NRS=0 M=1 R=4.93333 SA=75007.7 SB=75000.2
+ A=0.111 P=1.78 MULT=1
MM1000 N_A_27_368#_M1000_d N_D_M1000_g N_Y_M1000_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3864 AS=0.168 PD=2.93 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75000.3 SB=75003.4 A=0.168 P=2.54 MULT=1
MM1012 N_A_27_368#_M1012_d N_D_M1012_g N_Y_M1000_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75003 A=0.168 P=2.54 MULT=1
MM1013 N_A_27_368#_M1012_d N_D_M1013_g N_Y_M1013_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75001.2 SB=75002.5 A=0.168 P=2.54 MULT=1
MM1018 N_A_27_368#_M1018_d N_D_M1018_g N_Y_M1013_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.7 SB=75002 A=0.168 P=2.54 MULT=1
MM1005 N_A_496_368#_M1005_d N_C_M1005_g N_A_27_368#_M1018_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.1 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1011 N_A_496_368#_M1005_d N_C_M1011_g N_A_27_368#_M1011_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.6 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1016 N_A_496_368#_M1016_d N_C_M1016_g N_A_27_368#_M1011_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75003 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1021 N_A_496_368#_M1016_d N_C_M1021_g N_A_27_368#_M1021_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75003.5 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1003 N_A_496_368#_M1003_d N_B_M1003_g N_A_879_368#_M1003_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75003.6 A=0.168 P=2.54 MULT=1
MM1004 N_A_496_368#_M1003_d N_B_M1004_g N_A_879_368#_M1004_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.1792 PD=1.42 PS=1.44 NRD=1.7533 NRS=3.5066 M=1 R=7.46667
+ SA=75000.7 SB=75003.1 A=0.168 P=2.54 MULT=1
MM1006 N_A_496_368#_M1006_d N_B_M1006_g N_A_879_368#_M1004_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.1792 PD=1.42 PS=1.44 NRD=1.7533 NRS=3.5066 M=1 R=7.46667
+ SA=75001.1 SB=75002.7 A=0.168 P=2.54 MULT=1
MM1023 N_A_496_368#_M1006_d N_B_M1023_g N_A_879_368#_M1023_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.6 SB=75002.2 A=0.168 P=2.54 MULT=1
MM1001 N_A_879_368#_M1023_s N_A_M1001_g N_VPWR_M1001_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.224 PD=1.42 PS=1.52 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75002 SB=75001.8 A=0.168 P=2.54 MULT=1
MM1009 N_A_879_368#_M1009_d N_A_M1009_g N_VPWR_M1001_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.224 PD=1.42 PS=1.52 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75002.6 SB=75001.2 A=0.168 P=2.54 MULT=1
MM1014 N_A_879_368#_M1009_d N_A_M1014_g N_VPWR_M1014_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.224 PD=1.42 PS=1.52 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75003 SB=75000.8 A=0.168 P=2.54 MULT=1
MM1019 N_A_879_368#_M1019_d N_A_M1019_g N_VPWR_M1014_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.224 PD=2.83 PS=1.52 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75003.6 SB=75000.2 A=0.168 P=2.54 MULT=1
DX24_noxref VNB VPB NWDIODE A=16.7772 P=21.76
*
.include "sky130_fd_sc_ls__nor4_4.pxi.spice"
*
.ends
*
*
