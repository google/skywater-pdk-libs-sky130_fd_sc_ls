* File: sky130_fd_sc_ls__nand4bb_2.pxi.spice
* Created: Wed Sep  2 11:13:36 2020
* 
x_PM_SKY130_FD_SC_LS__NAND4BB_2%A_N N_A_N_c_111_n N_A_N_M1011_g N_A_N_M1018_g
+ A_N N_A_N_c_113_n PM_SKY130_FD_SC_LS__NAND4BB_2%A_N
x_PM_SKY130_FD_SC_LS__NAND4BB_2%B_N N_B_N_M1002_g N_B_N_c_148_n N_B_N_c_152_n
+ N_B_N_M1010_g B_N N_B_N_c_150_n PM_SKY130_FD_SC_LS__NAND4BB_2%B_N
x_PM_SKY130_FD_SC_LS__NAND4BB_2%A_27_368# N_A_27_368#_M1018_s
+ N_A_27_368#_M1011_s N_A_27_368#_c_186_n N_A_27_368#_M1008_g
+ N_A_27_368#_c_194_n N_A_27_368#_M1012_g N_A_27_368#_c_187_n
+ N_A_27_368#_M1016_g N_A_27_368#_c_195_n N_A_27_368#_M1017_g
+ N_A_27_368#_c_188_n N_A_27_368#_c_189_n N_A_27_368#_c_190_n
+ N_A_27_368#_c_198_n N_A_27_368#_c_199_n N_A_27_368#_c_191_n
+ N_A_27_368#_c_192_n N_A_27_368#_c_201_n N_A_27_368#_c_193_n
+ PM_SKY130_FD_SC_LS__NAND4BB_2%A_27_368#
x_PM_SKY130_FD_SC_LS__NAND4BB_2%A_231_74# N_A_231_74#_M1002_d
+ N_A_231_74#_M1010_d N_A_231_74#_c_291_n N_A_231_74#_M1001_g
+ N_A_231_74#_M1000_g N_A_231_74#_c_292_n N_A_231_74#_M1007_g
+ N_A_231_74#_M1014_g N_A_231_74#_c_293_n N_A_231_74#_c_285_n
+ N_A_231_74#_c_286_n N_A_231_74#_c_287_n N_A_231_74#_c_323_n
+ N_A_231_74#_c_325_n N_A_231_74#_c_288_n N_A_231_74#_c_357_p
+ N_A_231_74#_c_289_n N_A_231_74#_c_290_n
+ PM_SKY130_FD_SC_LS__NAND4BB_2%A_231_74#
x_PM_SKY130_FD_SC_LS__NAND4BB_2%C N_C_c_390_n N_C_M1004_g N_C_M1013_g
+ N_C_c_391_n N_C_M1006_g N_C_M1019_g C C N_C_c_388_n N_C_c_389_n
+ PM_SKY130_FD_SC_LS__NAND4BB_2%C
x_PM_SKY130_FD_SC_LS__NAND4BB_2%D N_D_c_448_n N_D_M1009_g N_D_M1003_g
+ N_D_c_449_n N_D_M1015_g N_D_M1005_g D N_D_c_446_n N_D_c_447_n
+ PM_SKY130_FD_SC_LS__NAND4BB_2%D
x_PM_SKY130_FD_SC_LS__NAND4BB_2%VPWR N_VPWR_M1011_d N_VPWR_M1012_s
+ N_VPWR_M1017_s N_VPWR_M1007_s N_VPWR_M1006_s N_VPWR_M1015_s N_VPWR_c_495_n
+ N_VPWR_c_496_n N_VPWR_c_497_n N_VPWR_c_498_n N_VPWR_c_499_n N_VPWR_c_500_n
+ N_VPWR_c_501_n N_VPWR_c_502_n N_VPWR_c_503_n N_VPWR_c_504_n N_VPWR_c_505_n
+ VPWR N_VPWR_c_506_n N_VPWR_c_507_n N_VPWR_c_508_n N_VPWR_c_509_n
+ N_VPWR_c_510_n N_VPWR_c_511_n N_VPWR_c_494_n
+ PM_SKY130_FD_SC_LS__NAND4BB_2%VPWR
x_PM_SKY130_FD_SC_LS__NAND4BB_2%Y N_Y_M1008_s N_Y_M1012_d N_Y_M1001_d
+ N_Y_M1004_d N_Y_M1009_d N_Y_c_592_n N_Y_c_586_n N_Y_c_587_n N_Y_c_600_n
+ N_Y_c_601_n N_Y_c_582_n N_Y_c_583_n N_Y_c_588_n N_Y_c_627_n N_Y_c_637_n
+ N_Y_c_589_n N_Y_c_641_n N_Y_c_644_n N_Y_c_590_n N_Y_c_606_n N_Y_c_646_n
+ N_Y_c_647_n Y N_Y_c_584_n Y PM_SKY130_FD_SC_LS__NAND4BB_2%Y
x_PM_SKY130_FD_SC_LS__NAND4BB_2%VGND N_VGND_M1018_d N_VGND_M1003_s
+ N_VGND_c_703_n N_VGND_c_704_n VGND N_VGND_c_705_n N_VGND_c_706_n
+ N_VGND_c_707_n N_VGND_c_708_n N_VGND_c_709_n N_VGND_c_710_n
+ PM_SKY130_FD_SC_LS__NAND4BB_2%VGND
x_PM_SKY130_FD_SC_LS__NAND4BB_2%A_373_74# N_A_373_74#_M1008_d
+ N_A_373_74#_M1016_d N_A_373_74#_M1014_d N_A_373_74#_c_762_n
+ N_A_373_74#_c_763_n N_A_373_74#_c_764_n N_A_373_74#_c_769_n
+ N_A_373_74#_c_770_n N_A_373_74#_c_765_n
+ PM_SKY130_FD_SC_LS__NAND4BB_2%A_373_74#
x_PM_SKY130_FD_SC_LS__NAND4BB_2%A_678_74# N_A_678_74#_M1000_s
+ N_A_678_74#_M1013_s N_A_678_74#_c_800_n N_A_678_74#_c_808_n
+ N_A_678_74#_c_801_n PM_SKY130_FD_SC_LS__NAND4BB_2%A_678_74#
x_PM_SKY130_FD_SC_LS__NAND4BB_2%A_886_74# N_A_886_74#_M1013_d
+ N_A_886_74#_M1019_d N_A_886_74#_M1005_d N_A_886_74#_c_828_n
+ N_A_886_74#_c_829_n N_A_886_74#_c_830_n N_A_886_74#_c_831_n
+ N_A_886_74#_c_832_n N_A_886_74#_c_833_n N_A_886_74#_c_834_n
+ PM_SKY130_FD_SC_LS__NAND4BB_2%A_886_74#
cc_1 VNB N_A_N_c_111_n 0.0365336f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_2 VNB N_A_N_M1018_g 0.03514f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.69
cc_3 VNB N_A_N_c_113_n 0.00693888f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.465
cc_4 VNB N_B_N_M1002_g 0.026521f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.34
cc_5 VNB N_B_N_c_148_n 0.0101242f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.69
cc_6 VNB B_N 0.00413281f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.465
cc_7 VNB N_B_N_c_150_n 0.0359383f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.465
cc_8 VNB N_A_27_368#_c_186_n 0.0187505f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_27_368#_c_187_n 0.0160904f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.465
cc_10 VNB N_A_27_368#_c_188_n 0.0301512f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_27_368#_c_189_n 0.0575891f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_368#_c_190_n 0.0227309f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_368#_c_191_n 0.00308008f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_368#_c_192_n 0.0136634f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_368#_c_193_n 0.0298922f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_231_74#_M1000_g 0.0242412f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.465
cc_17 VNB N_A_231_74#_M1014_g 0.02636f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_231_74#_c_285_n 0.0273422f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_231_74#_c_286_n 0.00999249f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_231_74#_c_287_n 0.0158903f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_231_74#_c_288_n 7.56474e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_231_74#_c_289_n 0.0059109f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_231_74#_c_290_n 0.0410517f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_C_M1013_g 0.0283133f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.69
cc_25 VNB N_C_M1019_g 0.0242061f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.465
cc_26 VNB N_C_c_388_n 0.0444016f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_C_c_389_n 0.00659658f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_D_M1003_g 0.0245196f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.69
cc_29 VNB N_D_M1005_g 0.0328675f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.465
cc_30 VNB D 0.016099f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_D_c_446_n 0.0390496f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_D_c_447_n 0.00283578f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VPWR_c_494_n 0.283096f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_Y_c_582_n 0.00765485f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_Y_c_583_n 2.81032e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_Y_c_584_n 0.00350986f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB Y 0.00973795f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_703_n 0.0160994f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_704_n 0.00635889f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.465
cc_40 VNB N_VGND_c_705_n 0.0193554f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_706_n 0.119321f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_707_n 0.01755f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_708_n 0.376185f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_709_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_710_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_373_74#_c_762_n 0.0030355f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.465
cc_47 VNB N_A_373_74#_c_763_n 0.00374022f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_373_74#_c_764_n 0.0045977f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.665
cc_49 VNB N_A_373_74#_c_765_n 0.00190736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_678_74#_c_800_n 0.0197769f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_678_74#_c_801_n 0.00201273f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.465
cc_52 VNB N_A_886_74#_c_828_n 0.00516762f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.465
cc_53 VNB N_A_886_74#_c_829_n 0.00396309f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_886_74#_c_830_n 0.00600345f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.665
cc_55 VNB N_A_886_74#_c_831_n 0.00206647f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_886_74#_c_832_n 0.0129966f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_886_74#_c_833_n 0.0266107f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_886_74#_c_834_n 0.00847193f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VPB N_A_N_c_111_n 0.0269721f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_60 VPB N_A_N_c_113_n 0.00484126f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.465
cc_61 VPB N_B_N_c_148_n 0.00101326f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=0.69
cc_62 VPB N_B_N_c_152_n 0.0254031f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_A_27_368#_c_194_n 0.0162433f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.465
cc_64 VPB N_A_27_368#_c_195_n 0.0165146f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_A_27_368#_c_188_n 0.0117307f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_A_27_368#_c_189_n 0.0136612f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_A_27_368#_c_198_n 0.0210799f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_A_27_368#_c_199_n 0.0169352f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_A_27_368#_c_191_n 0.00740183f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_A_27_368#_c_201_n 0.0179311f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_A_27_368#_c_193_n 0.0127393f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_A_231_74#_c_291_n 0.0166133f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_A_231_74#_c_292_n 0.0164104f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_A_231_74#_c_293_n 0.0106388f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_A_231_74#_c_286_n 0.00375326f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_A_231_74#_c_288_n 2.3955e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_A_231_74#_c_290_n 0.0222647f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_C_c_390_n 0.0167476f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_79 VPB N_C_c_391_n 0.0164867f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_80 VPB N_C_c_388_n 0.0248223f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_C_c_389_n 0.00834289f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 VPB N_D_c_448_n 0.0169259f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_83 VPB N_D_c_449_n 0.0190394f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_84 VPB D 0.00795763f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_D_c_446_n 0.0223745f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_D_c_447_n 8.96742e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_495_n 0.0195293f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_496_n 0.0187976f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_497_n 0.00830446f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_498_n 0.0128241f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_499_n 0.00830446f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_500_n 0.0120198f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_501_n 0.0484608f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_502_n 0.0274624f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_503_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_504_n 0.0186948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_505_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_506_n 0.0186948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_507_n 0.0186948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_508_n 0.0185368f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_509_n 0.0270017f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_102 VPB N_VPWR_c_510_n 0.0145925f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 VPB N_VPWR_c_511_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB N_VPWR_c_494_n 0.105548f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_105 VPB N_Y_c_586_n 0.00201649f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_Y_c_587_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB N_Y_c_588_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_Y_c_589_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_109 VPB N_Y_c_590_n 0.00289674f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_110 VPB Y 0.00475965f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 N_A_N_M1018_g N_B_N_M1002_g 0.0242833f $X=0.51 $Y=0.69 $X2=0 $Y2=0
cc_112 N_A_N_c_111_n N_B_N_c_148_n 0.00811074f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_113 N_A_N_c_113_n N_B_N_c_148_n 0.00312372f $X=0.6 $Y=1.465 $X2=0 $Y2=0
cc_114 N_A_N_c_111_n N_B_N_c_152_n 0.0266926f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_115 N_A_N_c_111_n B_N 2.32259e-19 $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_116 N_A_N_M1018_g B_N 6.76537e-19 $X=0.51 $Y=0.69 $X2=0 $Y2=0
cc_117 N_A_N_c_113_n B_N 0.0168772f $X=0.6 $Y=1.465 $X2=0 $Y2=0
cc_118 N_A_N_c_111_n N_B_N_c_150_n 0.0110681f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_119 N_A_N_c_113_n N_B_N_c_150_n 0.00129152f $X=0.6 $Y=1.465 $X2=0 $Y2=0
cc_120 N_A_N_M1018_g N_A_27_368#_c_190_n 0.00575762f $X=0.51 $Y=0.69 $X2=0 $Y2=0
cc_121 N_A_N_c_111_n N_A_27_368#_c_198_n 0.00698933f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_122 N_A_N_c_111_n N_A_27_368#_c_199_n 0.0150373f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_123 N_A_N_c_113_n N_A_27_368#_c_199_n 0.0135156f $X=0.6 $Y=1.465 $X2=0 $Y2=0
cc_124 N_A_N_c_111_n N_A_27_368#_c_192_n 8.32806e-19 $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_125 N_A_N_M1018_g N_A_27_368#_c_192_n 0.0029049f $X=0.51 $Y=0.69 $X2=0 $Y2=0
cc_126 N_A_N_c_113_n N_A_27_368#_c_192_n 0.00130596f $X=0.6 $Y=1.465 $X2=0 $Y2=0
cc_127 N_A_N_c_111_n N_A_27_368#_c_201_n 0.0068122f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_128 N_A_N_c_113_n N_A_27_368#_c_201_n 6.59727e-19 $X=0.6 $Y=1.465 $X2=0 $Y2=0
cc_129 N_A_N_c_111_n N_A_27_368#_c_193_n 0.0137873f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_130 N_A_N_M1018_g N_A_27_368#_c_193_n 0.00751517f $X=0.51 $Y=0.69 $X2=0 $Y2=0
cc_131 N_A_N_c_113_n N_A_27_368#_c_193_n 0.0365737f $X=0.6 $Y=1.465 $X2=0 $Y2=0
cc_132 N_A_N_c_111_n N_A_231_74#_c_293_n 0.00108102f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_133 N_A_N_c_113_n N_A_231_74#_c_286_n 0.0082347f $X=0.6 $Y=1.465 $X2=0 $Y2=0
cc_134 N_A_N_c_111_n N_VPWR_c_495_n 0.00598876f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_135 N_A_N_c_111_n N_VPWR_c_509_n 0.00481995f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_136 N_A_N_c_111_n N_VPWR_c_494_n 0.00508379f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_137 N_A_N_c_111_n N_VGND_c_703_n 9.50251e-19 $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_138 N_A_N_M1018_g N_VGND_c_703_n 0.0072585f $X=0.51 $Y=0.69 $X2=0 $Y2=0
cc_139 N_A_N_c_113_n N_VGND_c_703_n 0.0114275f $X=0.6 $Y=1.465 $X2=0 $Y2=0
cc_140 N_A_N_M1018_g N_VGND_c_705_n 0.00434272f $X=0.51 $Y=0.69 $X2=0 $Y2=0
cc_141 N_A_N_M1018_g N_VGND_c_708_n 0.0082502f $X=0.51 $Y=0.69 $X2=0 $Y2=0
cc_142 N_B_N_c_148_n N_A_27_368#_c_188_n 0.0020421f $X=1.125 $Y=1.675 $X2=0
+ $Y2=0
cc_143 N_B_N_c_150_n N_A_27_368#_c_188_n 0.00278569f $X=1.17 $Y=1.345 $X2=0
+ $Y2=0
cc_144 N_B_N_M1002_g N_A_27_368#_c_190_n 2.21897e-19 $X=1.08 $Y=0.69 $X2=0 $Y2=0
cc_145 N_B_N_c_152_n N_A_27_368#_c_199_n 0.021774f $X=1.125 $Y=1.765 $X2=0 $Y2=0
cc_146 N_B_N_c_152_n N_A_27_368#_c_191_n 0.00465428f $X=1.125 $Y=1.765 $X2=0
+ $Y2=0
cc_147 N_B_N_c_152_n N_A_27_368#_c_201_n 0.00214904f $X=1.125 $Y=1.765 $X2=0
+ $Y2=0
cc_148 N_B_N_c_152_n N_A_231_74#_c_293_n 0.0118192f $X=1.125 $Y=1.765 $X2=0
+ $Y2=0
cc_149 B_N N_A_231_74#_c_293_n 0.00733608f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_150 N_B_N_c_150_n N_A_231_74#_c_293_n 7.70522e-19 $X=1.17 $Y=1.345 $X2=0
+ $Y2=0
cc_151 N_B_N_M1002_g N_A_231_74#_c_285_n 0.0136048f $X=1.08 $Y=0.69 $X2=0 $Y2=0
cc_152 B_N N_A_231_74#_c_285_n 0.0142214f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_153 N_B_N_c_150_n N_A_231_74#_c_285_n 0.00123144f $X=1.17 $Y=1.345 $X2=0
+ $Y2=0
cc_154 N_B_N_c_148_n N_A_231_74#_c_286_n 0.00371505f $X=1.125 $Y=1.675 $X2=0
+ $Y2=0
cc_155 N_B_N_c_152_n N_A_231_74#_c_286_n 0.00145939f $X=1.125 $Y=1.765 $X2=0
+ $Y2=0
cc_156 B_N N_A_231_74#_c_286_n 0.0247641f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_157 N_B_N_c_150_n N_A_231_74#_c_286_n 0.00522964f $X=1.17 $Y=1.345 $X2=0
+ $Y2=0
cc_158 N_B_N_c_152_n N_VPWR_c_495_n 0.0112541f $X=1.125 $Y=1.765 $X2=0 $Y2=0
cc_159 N_B_N_c_152_n N_VPWR_c_496_n 0.00885633f $X=1.125 $Y=1.765 $X2=0 $Y2=0
cc_160 N_B_N_c_152_n N_VPWR_c_502_n 0.0049405f $X=1.125 $Y=1.765 $X2=0 $Y2=0
cc_161 N_B_N_c_152_n N_VPWR_c_494_n 0.00508379f $X=1.125 $Y=1.765 $X2=0 $Y2=0
cc_162 N_B_N_M1002_g N_VGND_c_703_n 0.00725816f $X=1.08 $Y=0.69 $X2=0 $Y2=0
cc_163 N_B_N_M1002_g N_VGND_c_706_n 0.00433139f $X=1.08 $Y=0.69 $X2=0 $Y2=0
cc_164 N_B_N_M1002_g N_VGND_c_708_n 0.00822643f $X=1.08 $Y=0.69 $X2=0 $Y2=0
cc_165 N_B_N_M1002_g N_A_373_74#_c_764_n 6.96305e-19 $X=1.08 $Y=0.69 $X2=0 $Y2=0
cc_166 N_A_27_368#_c_199_n N_A_231_74#_M1010_d 0.0184953f $X=1.845 $Y=2.325
+ $X2=0 $Y2=0
cc_167 N_A_27_368#_c_195_n N_A_231_74#_c_291_n 0.030654f $X=2.735 $Y=1.765 $X2=0
+ $Y2=0
cc_168 N_A_27_368#_c_187_n N_A_231_74#_M1000_g 0.0210727f $X=2.725 $Y=1.185
+ $X2=0 $Y2=0
cc_169 N_A_27_368#_c_189_n N_A_231_74#_M1000_g 0.00555143f $X=2.725 $Y=1.475
+ $X2=0 $Y2=0
cc_170 N_A_27_368#_c_199_n N_A_231_74#_c_293_n 0.0335903f $X=1.845 $Y=2.325
+ $X2=0 $Y2=0
cc_171 N_A_27_368#_c_191_n N_A_231_74#_c_293_n 0.021559f $X=2.01 $Y=1.515 $X2=0
+ $Y2=0
cc_172 N_A_27_368#_c_186_n N_A_231_74#_c_285_n 0.00551647f $X=2.27 $Y=1.185
+ $X2=0 $Y2=0
cc_173 N_A_27_368#_c_186_n N_A_231_74#_c_286_n 0.00338988f $X=2.27 $Y=1.185
+ $X2=0 $Y2=0
cc_174 N_A_27_368#_c_188_n N_A_231_74#_c_286_n 0.00356856f $X=2.195 $Y=1.515
+ $X2=0 $Y2=0
cc_175 N_A_27_368#_c_191_n N_A_231_74#_c_286_n 0.0358639f $X=2.01 $Y=1.515 $X2=0
+ $Y2=0
cc_176 N_A_27_368#_c_186_n N_A_231_74#_c_287_n 0.018062f $X=2.27 $Y=1.185 $X2=0
+ $Y2=0
cc_177 N_A_27_368#_c_187_n N_A_231_74#_c_287_n 0.00121168f $X=2.725 $Y=1.185
+ $X2=0 $Y2=0
cc_178 N_A_27_368#_c_188_n N_A_231_74#_c_287_n 0.00308089f $X=2.195 $Y=1.515
+ $X2=0 $Y2=0
cc_179 N_A_27_368#_c_191_n N_A_231_74#_c_287_n 0.0262124f $X=2.01 $Y=1.515 $X2=0
+ $Y2=0
cc_180 N_A_27_368#_c_189_n N_A_231_74#_c_323_n 0.0158912f $X=2.725 $Y=1.475
+ $X2=0 $Y2=0
cc_181 N_A_27_368#_c_191_n N_A_231_74#_c_323_n 0.00567911f $X=2.01 $Y=1.515
+ $X2=0 $Y2=0
cc_182 N_A_27_368#_c_189_n N_A_231_74#_c_325_n 0.00650229f $X=2.725 $Y=1.475
+ $X2=0 $Y2=0
cc_183 N_A_27_368#_c_191_n N_A_231_74#_c_325_n 0.0135702f $X=2.01 $Y=1.515 $X2=0
+ $Y2=0
cc_184 N_A_27_368#_c_189_n N_A_231_74#_c_288_n 5.14709e-19 $X=2.725 $Y=1.475
+ $X2=0 $Y2=0
cc_185 N_A_27_368#_c_189_n N_A_231_74#_c_289_n 0.0169413f $X=2.725 $Y=1.475
+ $X2=0 $Y2=0
cc_186 N_A_27_368#_c_189_n N_A_231_74#_c_290_n 0.0182673f $X=2.725 $Y=1.475
+ $X2=0 $Y2=0
cc_187 N_A_27_368#_c_199_n N_VPWR_M1011_d 0.0147844f $X=1.845 $Y=2.325 $X2=-0.19
+ $Y2=-0.245
cc_188 N_A_27_368#_c_199_n N_VPWR_M1012_s 0.00589703f $X=1.845 $Y=2.325 $X2=0
+ $Y2=0
cc_189 N_A_27_368#_c_191_n N_VPWR_M1012_s 0.0060416f $X=2.01 $Y=1.515 $X2=0
+ $Y2=0
cc_190 N_A_27_368#_c_198_n N_VPWR_c_495_n 0.0189321f $X=0.28 $Y=2.715 $X2=0
+ $Y2=0
cc_191 N_A_27_368#_c_199_n N_VPWR_c_495_n 0.0266856f $X=1.845 $Y=2.325 $X2=0
+ $Y2=0
cc_192 N_A_27_368#_c_194_n N_VPWR_c_496_n 0.0112021f $X=2.285 $Y=1.765 $X2=0
+ $Y2=0
cc_193 N_A_27_368#_c_199_n N_VPWR_c_496_n 0.0277468f $X=1.845 $Y=2.325 $X2=0
+ $Y2=0
cc_194 N_A_27_368#_c_195_n N_VPWR_c_497_n 0.00658161f $X=2.735 $Y=1.765 $X2=0
+ $Y2=0
cc_195 N_A_27_368#_c_194_n N_VPWR_c_504_n 0.00445602f $X=2.285 $Y=1.765 $X2=0
+ $Y2=0
cc_196 N_A_27_368#_c_195_n N_VPWR_c_504_n 0.00445602f $X=2.735 $Y=1.765 $X2=0
+ $Y2=0
cc_197 N_A_27_368#_c_198_n N_VPWR_c_509_n 0.0103978f $X=0.28 $Y=2.715 $X2=0
+ $Y2=0
cc_198 N_A_27_368#_c_194_n N_VPWR_c_494_n 0.00861719f $X=2.285 $Y=1.765 $X2=0
+ $Y2=0
cc_199 N_A_27_368#_c_195_n N_VPWR_c_494_n 0.00857825f $X=2.735 $Y=1.765 $X2=0
+ $Y2=0
cc_200 N_A_27_368#_c_198_n N_VPWR_c_494_n 0.0118739f $X=0.28 $Y=2.715 $X2=0
+ $Y2=0
cc_201 N_A_27_368#_c_187_n N_Y_c_592_n 0.00669329f $X=2.725 $Y=1.185 $X2=0 $Y2=0
cc_202 N_A_27_368#_c_189_n N_Y_c_592_n 0.00140079f $X=2.725 $Y=1.475 $X2=0 $Y2=0
cc_203 N_A_27_368#_c_194_n N_Y_c_586_n 0.00249249f $X=2.285 $Y=1.765 $X2=0 $Y2=0
cc_204 N_A_27_368#_c_195_n N_Y_c_586_n 0.00129805f $X=2.735 $Y=1.765 $X2=0 $Y2=0
cc_205 N_A_27_368#_c_189_n N_Y_c_586_n 0.00795655f $X=2.725 $Y=1.475 $X2=0 $Y2=0
cc_206 N_A_27_368#_c_191_n N_Y_c_586_n 0.00908697f $X=2.01 $Y=1.515 $X2=0 $Y2=0
cc_207 N_A_27_368#_c_194_n N_Y_c_587_n 0.0161044f $X=2.285 $Y=1.765 $X2=0 $Y2=0
cc_208 N_A_27_368#_c_195_n N_Y_c_587_n 0.0119101f $X=2.735 $Y=1.765 $X2=0 $Y2=0
cc_209 N_A_27_368#_c_195_n N_Y_c_600_n 0.0128707f $X=2.735 $Y=1.765 $X2=0 $Y2=0
cc_210 N_A_27_368#_c_186_n N_Y_c_601_n 7.63784e-19 $X=2.27 $Y=1.185 $X2=0 $Y2=0
cc_211 N_A_27_368#_c_187_n N_Y_c_601_n 0.00734808f $X=2.725 $Y=1.185 $X2=0 $Y2=0
cc_212 N_A_27_368#_c_187_n N_Y_c_583_n 0.00302705f $X=2.725 $Y=1.185 $X2=0 $Y2=0
cc_213 N_A_27_368#_c_189_n N_Y_c_583_n 0.00586261f $X=2.725 $Y=1.475 $X2=0 $Y2=0
cc_214 N_A_27_368#_c_195_n N_Y_c_588_n 3.75838e-19 $X=2.735 $Y=1.765 $X2=0 $Y2=0
cc_215 N_A_27_368#_c_195_n N_Y_c_606_n 3.07173e-19 $X=2.735 $Y=1.765 $X2=0 $Y2=0
cc_216 N_A_27_368#_c_190_n N_VGND_c_703_n 0.0259022f $X=0.295 $Y=0.515 $X2=0
+ $Y2=0
cc_217 N_A_27_368#_c_190_n N_VGND_c_705_n 0.0161257f $X=0.295 $Y=0.515 $X2=0
+ $Y2=0
cc_218 N_A_27_368#_c_186_n N_VGND_c_706_n 0.00288916f $X=2.27 $Y=1.185 $X2=0
+ $Y2=0
cc_219 N_A_27_368#_c_187_n N_VGND_c_706_n 0.00288916f $X=2.725 $Y=1.185 $X2=0
+ $Y2=0
cc_220 N_A_27_368#_c_186_n N_VGND_c_708_n 0.00362434f $X=2.27 $Y=1.185 $X2=0
+ $Y2=0
cc_221 N_A_27_368#_c_187_n N_VGND_c_708_n 0.0035883f $X=2.725 $Y=1.185 $X2=0
+ $Y2=0
cc_222 N_A_27_368#_c_190_n N_VGND_c_708_n 0.013291f $X=0.295 $Y=0.515 $X2=0
+ $Y2=0
cc_223 N_A_27_368#_c_186_n N_A_373_74#_c_763_n 0.0110252f $X=2.27 $Y=1.185 $X2=0
+ $Y2=0
cc_224 N_A_27_368#_c_187_n N_A_373_74#_c_763_n 0.0104231f $X=2.725 $Y=1.185
+ $X2=0 $Y2=0
cc_225 N_A_27_368#_c_187_n N_A_373_74#_c_769_n 0.00376849f $X=2.725 $Y=1.185
+ $X2=0 $Y2=0
cc_226 N_A_27_368#_c_187_n N_A_373_74#_c_770_n 6.66863e-19 $X=2.725 $Y=1.185
+ $X2=0 $Y2=0
cc_227 N_A_27_368#_c_187_n N_A_678_74#_c_801_n 4.68114e-19 $X=2.725 $Y=1.185
+ $X2=0 $Y2=0
cc_228 N_A_231_74#_c_291_n N_VPWR_c_497_n 0.00658161f $X=3.285 $Y=1.765 $X2=0
+ $Y2=0
cc_229 N_A_231_74#_c_292_n N_VPWR_c_498_n 0.00399808f $X=3.735 $Y=1.765 $X2=0
+ $Y2=0
cc_230 N_A_231_74#_c_291_n N_VPWR_c_506_n 0.00445602f $X=3.285 $Y=1.765 $X2=0
+ $Y2=0
cc_231 N_A_231_74#_c_292_n N_VPWR_c_506_n 0.00445602f $X=3.735 $Y=1.765 $X2=0
+ $Y2=0
cc_232 N_A_231_74#_c_291_n N_VPWR_c_494_n 0.00857825f $X=3.285 $Y=1.765 $X2=0
+ $Y2=0
cc_233 N_A_231_74#_c_292_n N_VPWR_c_494_n 0.00861719f $X=3.735 $Y=1.765 $X2=0
+ $Y2=0
cc_234 N_A_231_74#_c_287_n N_Y_M1008_s 0.00210949f $X=2.345 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_235 N_A_231_74#_c_287_n N_Y_c_592_n 0.00908783f $X=2.345 $Y=1.095 $X2=0 $Y2=0
cc_236 N_A_231_74#_c_289_n N_Y_c_592_n 0.003567f $X=3.125 $Y=1.555 $X2=0 $Y2=0
cc_237 N_A_231_74#_c_325_n N_Y_c_586_n 0.0122119f $X=2.515 $Y=1.515 $X2=0 $Y2=0
cc_238 N_A_231_74#_c_289_n N_Y_c_586_n 0.0105528f $X=3.125 $Y=1.555 $X2=0 $Y2=0
cc_239 N_A_231_74#_c_291_n N_Y_c_587_n 6.8381e-19 $X=3.285 $Y=1.765 $X2=0 $Y2=0
cc_240 N_A_231_74#_c_291_n N_Y_c_600_n 0.0124513f $X=3.285 $Y=1.765 $X2=0 $Y2=0
cc_241 N_A_231_74#_c_288_n N_Y_c_600_n 0.0134692f $X=3.375 $Y=1.555 $X2=0 $Y2=0
cc_242 N_A_231_74#_c_289_n N_Y_c_600_n 0.0227293f $X=3.125 $Y=1.555 $X2=0 $Y2=0
cc_243 N_A_231_74#_c_290_n N_Y_c_600_n 0.0014773f $X=3.735 $Y=1.557 $X2=0 $Y2=0
cc_244 N_A_231_74#_c_287_n N_Y_c_601_n 0.0062804f $X=2.345 $Y=1.095 $X2=0 $Y2=0
cc_245 N_A_231_74#_M1000_g N_Y_c_582_n 0.0111766f $X=3.315 $Y=0.74 $X2=0 $Y2=0
cc_246 N_A_231_74#_M1014_g N_Y_c_582_n 0.0123305f $X=3.745 $Y=0.74 $X2=0 $Y2=0
cc_247 N_A_231_74#_c_289_n N_Y_c_582_n 0.0684994f $X=3.125 $Y=1.555 $X2=0 $Y2=0
cc_248 N_A_231_74#_c_290_n N_Y_c_582_n 0.00559961f $X=3.735 $Y=1.557 $X2=0 $Y2=0
cc_249 N_A_231_74#_c_287_n N_Y_c_583_n 0.00798859f $X=2.345 $Y=1.095 $X2=0 $Y2=0
cc_250 N_A_231_74#_c_323_n N_Y_c_583_n 0.00603279f $X=2.43 $Y=1.43 $X2=0 $Y2=0
cc_251 N_A_231_74#_c_289_n N_Y_c_583_n 0.0130428f $X=3.125 $Y=1.555 $X2=0 $Y2=0
cc_252 N_A_231_74#_c_291_n N_Y_c_588_n 0.00957133f $X=3.285 $Y=1.765 $X2=0 $Y2=0
cc_253 N_A_231_74#_c_292_n N_Y_c_588_n 0.0146973f $X=3.735 $Y=1.765 $X2=0 $Y2=0
cc_254 N_A_231_74#_c_292_n N_Y_c_627_n 0.0178738f $X=3.735 $Y=1.765 $X2=0 $Y2=0
cc_255 N_A_231_74#_c_357_p N_Y_c_627_n 0.00864511f $X=3.63 $Y=1.515 $X2=0 $Y2=0
cc_256 N_A_231_74#_c_291_n N_Y_c_606_n 0.00239007f $X=3.285 $Y=1.765 $X2=0 $Y2=0
cc_257 N_A_231_74#_c_292_n N_Y_c_606_n 5.58885e-19 $X=3.735 $Y=1.765 $X2=0 $Y2=0
cc_258 N_A_231_74#_c_288_n N_Y_c_606_n 0.021414f $X=3.375 $Y=1.555 $X2=0 $Y2=0
cc_259 N_A_231_74#_c_290_n N_Y_c_606_n 0.00670438f $X=3.735 $Y=1.557 $X2=0 $Y2=0
cc_260 N_A_231_74#_c_292_n Y 0.00302973f $X=3.735 $Y=1.765 $X2=0 $Y2=0
cc_261 N_A_231_74#_M1014_g Y 0.00324507f $X=3.745 $Y=0.74 $X2=0 $Y2=0
cc_262 N_A_231_74#_c_357_p Y 0.0202512f $X=3.63 $Y=1.515 $X2=0 $Y2=0
cc_263 N_A_231_74#_c_290_n Y 0.0135557f $X=3.735 $Y=1.557 $X2=0 $Y2=0
cc_264 N_A_231_74#_c_285_n N_VGND_c_703_n 0.0276751f $X=1.59 $Y=1.18 $X2=0 $Y2=0
cc_265 N_A_231_74#_M1000_g N_VGND_c_706_n 0.00328473f $X=3.315 $Y=0.74 $X2=0
+ $Y2=0
cc_266 N_A_231_74#_M1014_g N_VGND_c_706_n 0.00278646f $X=3.745 $Y=0.74 $X2=0
+ $Y2=0
cc_267 N_A_231_74#_c_285_n N_VGND_c_706_n 0.0242075f $X=1.59 $Y=1.18 $X2=0 $Y2=0
cc_268 N_A_231_74#_M1000_g N_VGND_c_708_n 0.00429295f $X=3.315 $Y=0.74 $X2=0
+ $Y2=0
cc_269 N_A_231_74#_M1014_g N_VGND_c_708_n 0.00357517f $X=3.745 $Y=0.74 $X2=0
+ $Y2=0
cc_270 N_A_231_74#_c_285_n N_VGND_c_708_n 0.019994f $X=1.59 $Y=1.18 $X2=0 $Y2=0
cc_271 N_A_231_74#_c_287_n N_A_373_74#_M1008_d 0.00372399f $X=2.345 $Y=1.095
+ $X2=-0.19 $Y2=-0.245
cc_272 N_A_231_74#_c_285_n N_A_373_74#_c_762_n 0.0295158f $X=1.59 $Y=1.18 $X2=0
+ $Y2=0
cc_273 N_A_231_74#_c_287_n N_A_373_74#_c_762_n 0.0232663f $X=2.345 $Y=1.095
+ $X2=0 $Y2=0
cc_274 N_A_231_74#_M1000_g N_A_373_74#_c_763_n 0.00122855f $X=3.315 $Y=0.74
+ $X2=0 $Y2=0
cc_275 N_A_231_74#_c_287_n N_A_373_74#_c_763_n 0.0041185f $X=2.345 $Y=1.095
+ $X2=0 $Y2=0
cc_276 N_A_231_74#_c_285_n N_A_373_74#_c_764_n 0.0138246f $X=1.59 $Y=1.18 $X2=0
+ $Y2=0
cc_277 N_A_231_74#_M1000_g N_A_373_74#_c_765_n 0.011936f $X=3.315 $Y=0.74 $X2=0
+ $Y2=0
cc_278 N_A_231_74#_M1014_g N_A_373_74#_c_765_n 0.0090691f $X=3.745 $Y=0.74 $X2=0
+ $Y2=0
cc_279 N_A_231_74#_M1014_g N_A_678_74#_c_800_n 0.0100577f $X=3.745 $Y=0.74 $X2=0
+ $Y2=0
cc_280 N_A_231_74#_M1000_g N_A_678_74#_c_801_n 0.00591536f $X=3.315 $Y=0.74
+ $X2=0 $Y2=0
cc_281 N_A_231_74#_M1014_g N_A_678_74#_c_801_n 0.00947051f $X=3.745 $Y=0.74
+ $X2=0 $Y2=0
cc_282 N_A_231_74#_M1014_g N_A_886_74#_c_828_n 0.00192867f $X=3.745 $Y=0.74
+ $X2=0 $Y2=0
cc_283 N_A_231_74#_M1014_g N_A_886_74#_c_830_n 0.00225492f $X=3.745 $Y=0.74
+ $X2=0 $Y2=0
cc_284 N_C_c_391_n N_D_c_448_n 0.0317819f $X=5.165 $Y=1.765 $X2=-0.19 $Y2=-0.245
cc_285 N_C_c_389_n N_D_c_448_n 3.59818e-19 $X=5.22 $Y=1.515 $X2=-0.19 $Y2=-0.245
cc_286 N_C_M1019_g N_D_M1003_g 0.0195547f $X=5.29 $Y=0.74 $X2=0 $Y2=0
cc_287 N_C_c_388_n N_D_c_446_n 0.0207293f $X=5.22 $Y=1.515 $X2=0 $Y2=0
cc_288 N_C_c_389_n N_D_c_446_n 0.00265154f $X=5.22 $Y=1.515 $X2=0 $Y2=0
cc_289 N_C_c_388_n N_D_c_447_n 4.12009e-19 $X=5.22 $Y=1.515 $X2=0 $Y2=0
cc_290 N_C_c_389_n N_D_c_447_n 0.0210188f $X=5.22 $Y=1.515 $X2=0 $Y2=0
cc_291 N_C_c_390_n N_VPWR_c_498_n 0.00399808f $X=4.715 $Y=1.765 $X2=0 $Y2=0
cc_292 N_C_c_391_n N_VPWR_c_499_n 0.00598632f $X=5.165 $Y=1.765 $X2=0 $Y2=0
cc_293 N_C_c_390_n N_VPWR_c_507_n 0.00445602f $X=4.715 $Y=1.765 $X2=0 $Y2=0
cc_294 N_C_c_391_n N_VPWR_c_507_n 0.00445602f $X=5.165 $Y=1.765 $X2=0 $Y2=0
cc_295 N_C_c_390_n N_VPWR_c_494_n 0.00861719f $X=4.715 $Y=1.765 $X2=0 $Y2=0
cc_296 N_C_c_391_n N_VPWR_c_494_n 0.00857825f $X=5.165 $Y=1.765 $X2=0 $Y2=0
cc_297 N_C_c_390_n N_Y_c_637_n 0.0139279f $X=4.715 $Y=1.765 $X2=0 $Y2=0
cc_298 N_C_c_389_n N_Y_c_637_n 0.0232781f $X=5.22 $Y=1.515 $X2=0 $Y2=0
cc_299 N_C_c_390_n N_Y_c_589_n 0.0144423f $X=4.715 $Y=1.765 $X2=0 $Y2=0
cc_300 N_C_c_391_n N_Y_c_589_n 0.0103138f $X=5.165 $Y=1.765 $X2=0 $Y2=0
cc_301 N_C_c_391_n N_Y_c_641_n 0.0124513f $X=5.165 $Y=1.765 $X2=0 $Y2=0
cc_302 N_C_c_388_n N_Y_c_641_n 6.25269e-19 $X=5.22 $Y=1.515 $X2=0 $Y2=0
cc_303 N_C_c_389_n N_Y_c_641_n 0.0192955f $X=5.22 $Y=1.515 $X2=0 $Y2=0
cc_304 N_C_c_391_n N_Y_c_644_n 4.54145e-19 $X=5.165 $Y=1.765 $X2=0 $Y2=0
cc_305 N_C_c_391_n N_Y_c_590_n 6.63528e-19 $X=5.165 $Y=1.765 $X2=0 $Y2=0
cc_306 N_C_c_390_n N_Y_c_646_n 0.00307612f $X=4.715 $Y=1.765 $X2=0 $Y2=0
cc_307 N_C_c_390_n N_Y_c_647_n 4.27055e-19 $X=4.715 $Y=1.765 $X2=0 $Y2=0
cc_308 N_C_c_391_n N_Y_c_647_n 4.27055e-19 $X=5.165 $Y=1.765 $X2=0 $Y2=0
cc_309 N_C_c_388_n N_Y_c_647_n 0.00144303f $X=5.22 $Y=1.515 $X2=0 $Y2=0
cc_310 N_C_c_389_n N_Y_c_647_n 0.0237598f $X=5.22 $Y=1.515 $X2=0 $Y2=0
cc_311 N_C_M1013_g N_Y_c_584_n 0.00266115f $X=4.79 $Y=0.74 $X2=0 $Y2=0
cc_312 N_C_c_390_n Y 0.00193306f $X=4.715 $Y=1.765 $X2=0 $Y2=0
cc_313 N_C_M1013_g Y 0.00218978f $X=4.79 $Y=0.74 $X2=0 $Y2=0
cc_314 N_C_c_388_n Y 0.0019102f $X=5.22 $Y=1.515 $X2=0 $Y2=0
cc_315 N_C_c_389_n Y 0.0281718f $X=5.22 $Y=1.515 $X2=0 $Y2=0
cc_316 N_C_M1013_g N_VGND_c_706_n 0.00278271f $X=4.79 $Y=0.74 $X2=0 $Y2=0
cc_317 N_C_M1019_g N_VGND_c_706_n 0.00430908f $X=5.29 $Y=0.74 $X2=0 $Y2=0
cc_318 N_C_M1013_g N_VGND_c_708_n 0.00359085f $X=4.79 $Y=0.74 $X2=0 $Y2=0
cc_319 N_C_M1019_g N_VGND_c_708_n 0.00817424f $X=5.29 $Y=0.74 $X2=0 $Y2=0
cc_320 N_C_M1013_g N_A_678_74#_c_800_n 0.0132866f $X=4.79 $Y=0.74 $X2=0 $Y2=0
cc_321 N_C_M1019_g N_A_678_74#_c_800_n 0.0051084f $X=5.29 $Y=0.74 $X2=0 $Y2=0
cc_322 N_C_M1019_g N_A_678_74#_c_808_n 0.00472624f $X=5.29 $Y=0.74 $X2=0 $Y2=0
cc_323 N_C_M1013_g N_A_886_74#_c_828_n 0.00667517f $X=4.79 $Y=0.74 $X2=0 $Y2=0
cc_324 N_C_M1019_g N_A_886_74#_c_828_n 8.48828e-19 $X=5.29 $Y=0.74 $X2=0 $Y2=0
cc_325 N_C_M1013_g N_A_886_74#_c_829_n 0.0093986f $X=4.79 $Y=0.74 $X2=0 $Y2=0
cc_326 N_C_M1019_g N_A_886_74#_c_829_n 0.0134906f $X=5.29 $Y=0.74 $X2=0 $Y2=0
cc_327 N_C_c_388_n N_A_886_74#_c_829_n 0.00441409f $X=5.22 $Y=1.515 $X2=0 $Y2=0
cc_328 N_C_c_389_n N_A_886_74#_c_829_n 0.0484156f $X=5.22 $Y=1.515 $X2=0 $Y2=0
cc_329 N_C_M1013_g N_A_886_74#_c_830_n 0.00417978f $X=4.79 $Y=0.74 $X2=0 $Y2=0
cc_330 N_C_c_388_n N_A_886_74#_c_830_n 0.00239344f $X=5.22 $Y=1.515 $X2=0 $Y2=0
cc_331 N_C_c_389_n N_A_886_74#_c_830_n 0.0256033f $X=5.22 $Y=1.515 $X2=0 $Y2=0
cc_332 N_C_M1019_g N_A_886_74#_c_831_n 3.97173e-19 $X=5.29 $Y=0.74 $X2=0 $Y2=0
cc_333 N_D_c_448_n N_VPWR_c_499_n 0.00598632f $X=5.715 $Y=1.765 $X2=0 $Y2=0
cc_334 N_D_c_448_n N_VPWR_c_501_n 5.87829e-19 $X=5.715 $Y=1.765 $X2=0 $Y2=0
cc_335 N_D_c_449_n N_VPWR_c_501_n 0.0137469f $X=6.205 $Y=1.765 $X2=0 $Y2=0
cc_336 D N_VPWR_c_501_n 0.0203491f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_337 N_D_c_447_n N_VPWR_c_501_n 0.00356189f $X=6.365 $Y=1.565 $X2=0 $Y2=0
cc_338 N_D_c_448_n N_VPWR_c_508_n 0.00445602f $X=5.715 $Y=1.765 $X2=0 $Y2=0
cc_339 N_D_c_449_n N_VPWR_c_508_n 0.00444681f $X=6.205 $Y=1.765 $X2=0 $Y2=0
cc_340 N_D_c_448_n N_VPWR_c_494_n 0.00858197f $X=5.715 $Y=1.765 $X2=0 $Y2=0
cc_341 N_D_c_449_n N_VPWR_c_494_n 0.00878088f $X=6.205 $Y=1.765 $X2=0 $Y2=0
cc_342 N_D_c_448_n N_Y_c_589_n 6.63528e-19 $X=5.715 $Y=1.765 $X2=0 $Y2=0
cc_343 N_D_c_448_n N_Y_c_641_n 0.012969f $X=5.715 $Y=1.765 $X2=0 $Y2=0
cc_344 N_D_c_447_n N_Y_c_641_n 0.00702711f $X=6.365 $Y=1.565 $X2=0 $Y2=0
cc_345 N_D_c_448_n N_Y_c_644_n 0.00236769f $X=5.715 $Y=1.765 $X2=0 $Y2=0
cc_346 N_D_c_446_n N_Y_c_644_n 0.00727595f $X=6.205 $Y=1.557 $X2=0 $Y2=0
cc_347 N_D_c_447_n N_Y_c_644_n 0.0231738f $X=6.365 $Y=1.565 $X2=0 $Y2=0
cc_348 N_D_c_448_n N_Y_c_590_n 0.0105414f $X=5.715 $Y=1.765 $X2=0 $Y2=0
cc_349 N_D_c_449_n N_Y_c_590_n 2.77576e-19 $X=6.205 $Y=1.765 $X2=0 $Y2=0
cc_350 N_D_M1003_g N_VGND_c_704_n 0.00429635f $X=5.72 $Y=0.74 $X2=0 $Y2=0
cc_351 N_D_M1005_g N_VGND_c_704_n 0.0131831f $X=6.22 $Y=0.74 $X2=0 $Y2=0
cc_352 N_D_M1003_g N_VGND_c_706_n 0.00434272f $X=5.72 $Y=0.74 $X2=0 $Y2=0
cc_353 N_D_M1005_g N_VGND_c_707_n 0.00383152f $X=6.22 $Y=0.74 $X2=0 $Y2=0
cc_354 N_D_M1003_g N_VGND_c_708_n 0.00820816f $X=5.72 $Y=0.74 $X2=0 $Y2=0
cc_355 N_D_M1005_g N_VGND_c_708_n 0.00761215f $X=6.22 $Y=0.74 $X2=0 $Y2=0
cc_356 N_D_M1003_g N_A_678_74#_c_800_n 3.17554e-19 $X=5.72 $Y=0.74 $X2=0 $Y2=0
cc_357 N_D_M1003_g N_A_886_74#_c_831_n 0.00934902f $X=5.72 $Y=0.74 $X2=0 $Y2=0
cc_358 N_D_M1005_g N_A_886_74#_c_831_n 0.00101123f $X=6.22 $Y=0.74 $X2=0 $Y2=0
cc_359 N_D_M1003_g N_A_886_74#_c_832_n 0.0115433f $X=5.72 $Y=0.74 $X2=0 $Y2=0
cc_360 N_D_M1005_g N_A_886_74#_c_832_n 0.0140711f $X=6.22 $Y=0.74 $X2=0 $Y2=0
cc_361 N_D_c_446_n N_A_886_74#_c_832_n 0.00381149f $X=6.205 $Y=1.557 $X2=0 $Y2=0
cc_362 N_D_c_447_n N_A_886_74#_c_832_n 0.0722592f $X=6.365 $Y=1.565 $X2=0 $Y2=0
cc_363 N_D_M1005_g N_A_886_74#_c_833_n 0.00159319f $X=6.22 $Y=0.74 $X2=0 $Y2=0
cc_364 N_D_M1003_g N_A_886_74#_c_834_n 0.00155819f $X=5.72 $Y=0.74 $X2=0 $Y2=0
cc_365 N_D_c_446_n N_A_886_74#_c_834_n 5.01936e-19 $X=6.205 $Y=1.557 $X2=0 $Y2=0
cc_366 N_D_c_447_n N_A_886_74#_c_834_n 0.00368228f $X=6.365 $Y=1.565 $X2=0 $Y2=0
cc_367 N_VPWR_c_496_n N_Y_c_587_n 0.0157994f $X=2.01 $Y=2.78 $X2=0 $Y2=0
cc_368 N_VPWR_c_497_n N_Y_c_587_n 0.0304332f $X=3.01 $Y=2.355 $X2=0 $Y2=0
cc_369 N_VPWR_c_504_n N_Y_c_587_n 0.014552f $X=2.845 $Y=3.33 $X2=0 $Y2=0
cc_370 N_VPWR_c_494_n N_Y_c_587_n 0.0119791f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_371 N_VPWR_M1017_s N_Y_c_600_n 0.00689416f $X=2.81 $Y=1.84 $X2=0 $Y2=0
cc_372 N_VPWR_c_497_n N_Y_c_600_n 0.0232685f $X=3.01 $Y=2.355 $X2=0 $Y2=0
cc_373 N_VPWR_c_497_n N_Y_c_588_n 0.0304332f $X=3.01 $Y=2.355 $X2=0 $Y2=0
cc_374 N_VPWR_c_498_n N_Y_c_588_n 0.0267725f $X=4.49 $Y=2.455 $X2=0 $Y2=0
cc_375 N_VPWR_c_506_n N_Y_c_588_n 0.014552f $X=3.845 $Y=3.33 $X2=0 $Y2=0
cc_376 N_VPWR_c_494_n N_Y_c_588_n 0.0119791f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_377 N_VPWR_M1007_s N_Y_c_627_n 0.00284152f $X=3.81 $Y=1.84 $X2=0 $Y2=0
cc_378 N_VPWR_c_498_n N_Y_c_627_n 0.00819043f $X=4.49 $Y=2.455 $X2=0 $Y2=0
cc_379 N_VPWR_M1007_s N_Y_c_637_n 0.0175401f $X=3.81 $Y=1.84 $X2=0 $Y2=0
cc_380 N_VPWR_c_498_n N_Y_c_637_n 0.0315306f $X=4.49 $Y=2.455 $X2=0 $Y2=0
cc_381 N_VPWR_c_498_n N_Y_c_589_n 0.0267725f $X=4.49 $Y=2.455 $X2=0 $Y2=0
cc_382 N_VPWR_c_499_n N_Y_c_589_n 0.0266809f $X=5.44 $Y=2.455 $X2=0 $Y2=0
cc_383 N_VPWR_c_507_n N_Y_c_589_n 0.014552f $X=5.275 $Y=3.33 $X2=0 $Y2=0
cc_384 N_VPWR_c_494_n N_Y_c_589_n 0.0119791f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_385 N_VPWR_M1006_s N_Y_c_641_n 0.0117318f $X=5.24 $Y=1.84 $X2=0 $Y2=0
cc_386 N_VPWR_c_499_n N_Y_c_641_n 0.0232685f $X=5.44 $Y=2.455 $X2=0 $Y2=0
cc_387 N_VPWR_c_499_n N_Y_c_590_n 0.0266809f $X=5.44 $Y=2.455 $X2=0 $Y2=0
cc_388 N_VPWR_c_501_n N_Y_c_590_n 0.0330597f $X=6.44 $Y=2.115 $X2=0 $Y2=0
cc_389 N_VPWR_c_508_n N_Y_c_590_n 0.0145938f $X=6.275 $Y=3.33 $X2=0 $Y2=0
cc_390 N_VPWR_c_494_n N_Y_c_590_n 0.0120466f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_391 N_VPWR_M1007_s N_Y_c_646_n 0.00731928f $X=3.81 $Y=1.84 $X2=0 $Y2=0
cc_392 N_VPWR_c_498_n N_Y_c_646_n 0.020647f $X=4.49 $Y=2.455 $X2=0 $Y2=0
cc_393 N_VPWR_M1007_s Y 3.45784e-19 $X=3.81 $Y=1.84 $X2=0 $Y2=0
cc_394 N_Y_c_582_n N_A_373_74#_M1016_d 0.00505217f $X=3.965 $Y=1.175 $X2=0 $Y2=0
cc_395 N_Y_c_582_n N_A_373_74#_M1014_d 9.27081e-19 $X=3.965 $Y=1.175 $X2=0 $Y2=0
cc_396 N_Y_c_584_n N_A_373_74#_M1014_d 0.00234035f $X=4.08 $Y=1.26 $X2=0 $Y2=0
cc_397 N_Y_M1008_s N_A_373_74#_c_763_n 0.00193522f $X=2.345 $Y=0.37 $X2=0 $Y2=0
cc_398 N_Y_c_592_n N_A_373_74#_c_763_n 0.023659f $X=2.685 $Y=0.755 $X2=0 $Y2=0
cc_399 N_Y_c_582_n N_A_373_74#_c_763_n 0.00480411f $X=3.965 $Y=1.175 $X2=0 $Y2=0
cc_400 N_Y_c_582_n N_A_373_74#_c_770_n 0.0127069f $X=3.965 $Y=1.175 $X2=0 $Y2=0
cc_401 N_Y_c_582_n N_A_373_74#_c_765_n 0.0387128f $X=3.965 $Y=1.175 $X2=0 $Y2=0
cc_402 N_Y_c_584_n N_A_373_74#_c_765_n 0.0175541f $X=4.08 $Y=1.26 $X2=0 $Y2=0
cc_403 N_Y_c_582_n N_A_678_74#_M1000_s 0.00176891f $X=3.965 $Y=1.175 $X2=-0.19
+ $Y2=-0.245
cc_404 N_Y_c_584_n N_A_678_74#_c_800_n 4.87282e-19 $X=4.08 $Y=1.26 $X2=0 $Y2=0
cc_405 N_Y_c_584_n N_A_886_74#_c_830_n 0.00714078f $X=4.08 $Y=1.26 $X2=0 $Y2=0
cc_406 N_VGND_c_706_n N_A_373_74#_c_763_n 0.0442921f $X=5.84 $Y=0 $X2=0 $Y2=0
cc_407 N_VGND_c_708_n N_A_373_74#_c_763_n 0.0353647f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_408 N_VGND_c_706_n N_A_373_74#_c_764_n 0.0156771f $X=5.84 $Y=0 $X2=0 $Y2=0
cc_409 N_VGND_c_708_n N_A_373_74#_c_764_n 0.0122201f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_410 N_VGND_c_706_n N_A_373_74#_c_765_n 0.00193679f $X=5.84 $Y=0 $X2=0 $Y2=0
cc_411 N_VGND_c_708_n N_A_373_74#_c_765_n 0.00572201f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_412 N_VGND_c_704_n N_A_678_74#_c_800_n 0.00302522f $X=6.005 $Y=0.65 $X2=0
+ $Y2=0
cc_413 N_VGND_c_706_n N_A_678_74#_c_800_n 0.100668f $X=5.84 $Y=0 $X2=0 $Y2=0
cc_414 N_VGND_c_708_n N_A_678_74#_c_800_n 0.057077f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_415 N_VGND_c_706_n N_A_678_74#_c_801_n 0.0221127f $X=5.84 $Y=0 $X2=0 $Y2=0
cc_416 N_VGND_c_708_n N_A_678_74#_c_801_n 0.012301f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_417 N_VGND_c_704_n N_A_886_74#_c_831_n 0.0175116f $X=6.005 $Y=0.65 $X2=0
+ $Y2=0
cc_418 N_VGND_c_706_n N_A_886_74#_c_831_n 0.0109942f $X=5.84 $Y=0 $X2=0 $Y2=0
cc_419 N_VGND_c_708_n N_A_886_74#_c_831_n 0.00904371f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_420 N_VGND_M1003_s N_A_886_74#_c_832_n 0.00266f $X=5.795 $Y=0.37 $X2=0 $Y2=0
cc_421 N_VGND_c_704_n N_A_886_74#_c_832_n 0.018932f $X=6.005 $Y=0.65 $X2=0 $Y2=0
cc_422 N_VGND_c_704_n N_A_886_74#_c_833_n 0.0173942f $X=6.005 $Y=0.65 $X2=0
+ $Y2=0
cc_423 N_VGND_c_707_n N_A_886_74#_c_833_n 0.011066f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_424 N_VGND_c_708_n N_A_886_74#_c_833_n 0.00915947f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_425 N_A_373_74#_c_765_n N_A_678_74#_M1000_s 0.0033542f $X=3.985 $Y=0.835
+ $X2=-0.19 $Y2=-0.245
cc_426 N_A_373_74#_M1014_d N_A_678_74#_c_800_n 0.0045553f $X=3.82 $Y=0.37 $X2=0
+ $Y2=0
cc_427 N_A_373_74#_c_765_n N_A_678_74#_c_800_n 0.0164472f $X=3.985 $Y=0.835
+ $X2=0 $Y2=0
cc_428 N_A_373_74#_c_763_n N_A_678_74#_c_801_n 0.00822726f $X=3.025 $Y=0.415
+ $X2=0 $Y2=0
cc_429 N_A_373_74#_c_765_n N_A_678_74#_c_801_n 0.0155728f $X=3.985 $Y=0.835
+ $X2=0 $Y2=0
cc_430 N_A_373_74#_c_765_n N_A_886_74#_c_828_n 0.0120186f $X=3.985 $Y=0.835
+ $X2=0 $Y2=0
cc_431 N_A_678_74#_c_800_n N_A_886_74#_M1013_d 0.00288367f $X=4.91 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_432 N_A_678_74#_c_800_n N_A_886_74#_c_828_n 0.0179715f $X=4.91 $Y=0.34 $X2=0
+ $Y2=0
cc_433 N_A_678_74#_M1013_s N_A_886_74#_c_829_n 0.00266f $X=4.865 $Y=0.37 $X2=0
+ $Y2=0
cc_434 N_A_678_74#_c_800_n N_A_886_74#_c_829_n 0.00304353f $X=4.91 $Y=0.34 $X2=0
+ $Y2=0
cc_435 N_A_678_74#_c_808_n N_A_886_74#_c_829_n 0.0186354f $X=5.075 $Y=0.65 $X2=0
+ $Y2=0
cc_436 N_A_678_74#_c_800_n N_A_886_74#_c_831_n 0.00374778f $X=4.91 $Y=0.34 $X2=0
+ $Y2=0
