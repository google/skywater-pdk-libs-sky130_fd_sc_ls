* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__or3b_4 A B C_N VGND VNB VPB VPWR X
X0 a_307_392# B a_217_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_409_392# a_27_392# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X2 X a_409_392# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X3 a_217_392# B a_307_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 a_217_392# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 VGND a_409_392# X VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X6 VPWR a_409_392# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X7 VPWR a_409_392# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X8 X a_409_392# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X9 a_409_392# a_27_392# a_307_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_27_392# C_N VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X11 a_27_392# C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 a_307_392# a_27_392# a_409_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 X a_409_392# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X14 VPWR A a_217_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 VGND B a_409_392# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X16 a_409_392# A VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X17 X a_409_392# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X18 VGND a_409_392# X VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
.ends
