* NGSPICE file created from sky130_fd_sc_ls__nor2b_1.ext - technology: sky130A

.subckt sky130_fd_sc_ls__nor2b_1 A B_N VGND VNB VPB VPWR Y
M1000 Y a_27_112# a_278_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=4.2e+11p pd=2.99e+06u as=3.024e+11p ps=2.78e+06u
M1001 VGND a_27_112# Y VNB nshort w=740000u l=150000u
+  ad=5.6985e+11p pd=4.59e+06u as=2.627e+11p ps=2.19e+06u
M1002 a_278_368# A VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=4.69e+11p ps=3.16e+06u
M1003 VPWR B_N a_27_112# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=2.478e+11p ps=2.27e+06u
M1004 VGND B_N a_27_112# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=2.805e+11p ps=2.12e+06u
M1005 Y A VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

