# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ls__o2111ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_ls__o2111ai_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.08000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.285000 1.350000 7.635000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.805000 1.350000 9.490000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.780000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445000 1.350000 6.115000 1.780000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.780000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.210000 1.300000 4.195000 1.630000 ;
        RECT 3.965000 1.630000 4.195000 1.780000 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.780000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.350000 1.350000 1.780000 ;
    END
  END D1
  PIN Y
    ANTENNADIFFAREA  3.411800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115000 1.950000 9.515000 1.970000 ;
        RECT 0.115000 1.970000 2.200000 2.120000 ;
        RECT 0.115000 2.120000 1.200000 2.980000 ;
        RECT 0.615000 0.770000 1.805000 1.130000 ;
        RECT 1.565000 1.130000 1.805000 1.550000 ;
        RECT 1.565000 1.550000 2.040000 1.780000 ;
        RECT 1.870000 1.780000 2.040000 1.800000 ;
        RECT 1.870000 1.800000 3.520000 1.950000 ;
        RECT 1.870000 2.120000 2.200000 2.980000 ;
        RECT 3.190000 1.970000 9.515000 2.120000 ;
        RECT 3.190000 2.120000 3.520000 2.980000 ;
        RECT 4.190000 2.120000 4.520000 2.980000 ;
        RECT 8.185000 2.120000 8.515000 2.735000 ;
        RECT 9.185000 2.120000 9.515000 2.735000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.080000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 10.080000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.080000 0.085000 ;
      RECT 0.000000  3.245000 10.080000 3.415000 ;
      RECT 0.115000  0.350000  2.155000 0.600000 ;
      RECT 0.115000  0.600000  0.445000 1.130000 ;
      RECT 1.370000  2.290000  1.700000 3.245000 ;
      RECT 1.985000  0.600000  2.155000 0.815000 ;
      RECT 1.985000  0.815000  3.955000 1.130000 ;
      RECT 2.335000  0.350000  5.805000 0.645000 ;
      RECT 2.370000  2.140000  3.020000 3.245000 ;
      RECT 3.690000  2.290000  4.020000 3.245000 ;
      RECT 4.185000  0.815000  4.515000 0.850000 ;
      RECT 4.185000  0.850000  6.305000 1.010000 ;
      RECT 4.185000  1.010000  9.965000 1.130000 ;
      RECT 4.750000  2.290000  8.015000 2.460000 ;
      RECT 4.750000  2.460000  6.165000 2.980000 ;
      RECT 5.045000  1.130000  9.965000 1.180000 ;
      RECT 5.475000  0.645000  5.805000 0.680000 ;
      RECT 5.975000  0.350000  6.305000 0.850000 ;
      RECT 6.335000  2.630000  6.585000 3.245000 ;
      RECT 6.475000  0.085000  6.805000 0.820000 ;
      RECT 6.785000  2.460000  7.115000 2.980000 ;
      RECT 6.985000  0.350000  7.155000 1.010000 ;
      RECT 7.315000  2.630000  7.485000 3.245000 ;
      RECT 7.335000  0.085000  7.665000 0.820000 ;
      RECT 7.685000  2.460000  8.015000 2.905000 ;
      RECT 7.685000  2.905000  9.965000 3.075000 ;
      RECT 7.845000  0.350000  8.095000 1.010000 ;
      RECT 8.265000  0.085000  8.595000 0.820000 ;
      RECT 8.685000  2.290000  9.015000 2.905000 ;
      RECT 8.775000  0.350000  9.025000 1.010000 ;
      RECT 9.205000  0.085000  9.535000 0.820000 ;
      RECT 9.715000  0.350000  9.965000 1.010000 ;
      RECT 9.715000  1.820000  9.965000 2.905000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
      RECT 9.275000 -0.085000 9.445000 0.085000 ;
      RECT 9.275000  3.245000 9.445000 3.415000 ;
      RECT 9.755000 -0.085000 9.925000 0.085000 ;
      RECT 9.755000  3.245000 9.925000 3.415000 ;
  END
END sky130_fd_sc_ls__o2111ai_4
END LIBRARY
