* File: sky130_fd_sc_ls__or3_2.pxi.spice
* Created: Wed Sep  2 11:24:52 2020
* 
x_PM_SKY130_FD_SC_LS__OR3_2%C N_C_M1008_g N_C_c_61_n N_C_c_66_n N_C_M1003_g C C
+ N_C_c_62_n N_C_c_63_n N_C_c_64_n PM_SKY130_FD_SC_LS__OR3_2%C
x_PM_SKY130_FD_SC_LS__OR3_2%B N_B_c_103_n N_B_M1002_g N_B_M1006_g N_B_c_99_n
+ N_B_c_100_n B B B N_B_c_101_n N_B_c_102_n PM_SKY130_FD_SC_LS__OR3_2%B
x_PM_SKY130_FD_SC_LS__OR3_2%A N_A_M1004_g N_A_c_147_n N_A_c_151_n N_A_M1001_g A
+ N_A_c_149_n PM_SKY130_FD_SC_LS__OR3_2%A
x_PM_SKY130_FD_SC_LS__OR3_2%A_27_74# N_A_27_74#_M1008_s N_A_27_74#_M1006_d
+ N_A_27_74#_M1003_s N_A_27_74#_c_199_n N_A_27_74#_M1000_g N_A_27_74#_M1005_g
+ N_A_27_74#_c_200_n N_A_27_74#_M1007_g N_A_27_74#_M1009_g N_A_27_74#_c_191_n
+ N_A_27_74#_c_192_n N_A_27_74#_c_202_n N_A_27_74#_c_211_n N_A_27_74#_c_193_n
+ N_A_27_74#_c_234_n N_A_27_74#_c_194_n N_A_27_74#_c_195_n N_A_27_74#_c_196_n
+ N_A_27_74#_c_197_n N_A_27_74#_c_203_n N_A_27_74#_c_226_n N_A_27_74#_c_198_n
+ PM_SKY130_FD_SC_LS__OR3_2%A_27_74#
x_PM_SKY130_FD_SC_LS__OR3_2%VPWR N_VPWR_M1001_d N_VPWR_M1007_d N_VPWR_c_298_n
+ N_VPWR_c_299_n N_VPWR_c_300_n N_VPWR_c_301_n N_VPWR_c_302_n VPWR
+ N_VPWR_c_303_n N_VPWR_c_297_n PM_SKY130_FD_SC_LS__OR3_2%VPWR
x_PM_SKY130_FD_SC_LS__OR3_2%X N_X_M1005_d N_X_M1000_s N_X_c_337_n N_X_c_333_n
+ N_X_c_338_n N_X_c_339_n N_X_c_334_n N_X_c_335_n X X
+ PM_SKY130_FD_SC_LS__OR3_2%X
x_PM_SKY130_FD_SC_LS__OR3_2%VGND N_VGND_M1008_d N_VGND_M1004_d N_VGND_M1009_s
+ N_VGND_c_379_n N_VGND_c_380_n N_VGND_c_381_n VGND N_VGND_c_382_n
+ N_VGND_c_383_n N_VGND_c_384_n N_VGND_c_385_n N_VGND_c_386_n
+ PM_SKY130_FD_SC_LS__OR3_2%VGND
cc_1 VNB N_C_c_61_n 0.0264575f $X=-0.19 $Y=-0.245 $X2=0.592 $Y2=1.618
cc_2 VNB N_C_c_62_n 0.0180279f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.285
cc_3 VNB N_C_c_63_n 0.00582239f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.285
cc_4 VNB N_C_c_64_n 0.0231661f $X=-0.19 $Y=-0.245 $X2=0.592 $Y2=1.12
cc_5 VNB N_B_c_99_n 0.0207084f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=2.46
cc_6 VNB N_B_c_100_n 0.0256663f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_7 VNB N_B_c_101_n 0.016747f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.285
cc_8 VNB N_B_c_102_n 0.00168225f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_M1004_g 0.0253763f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.69
cc_10 VNB N_A_c_147_n 0.00654081f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=1.885
cc_11 VNB A 0.00702351f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_12 VNB N_A_c_149_n 0.0310448f $X=-0.19 $Y=-0.245 $X2=0.592 $Y2=1.285
cc_13 VNB N_A_27_74#_M1005_g 0.023704f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.285
cc_14 VNB N_A_27_74#_M1009_g 0.0225458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_74#_c_191_n 0.0195766f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_27_74#_c_192_n 0.0324859f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_27_74#_c_193_n 0.00279936f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_27_74#_c_194_n 0.00321738f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_27_74#_c_195_n 0.00704396f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_27_74#_c_196_n 0.00174694f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_27_74#_c_197_n 0.00717518f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_27_74#_c_198_n 0.0585368f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VPWR_c_297_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_X_c_333_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.285
cc_25 VNB N_X_c_334_n 0.00924703f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.295
cc_26 VNB N_X_c_335_n 0.00230427f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB X 0.0270256f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_379_n 0.00993412f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_380_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.285
cc_30 VNB N_VGND_c_381_n 0.0289902f $X=-0.19 $Y=-0.245 $X2=0.592 $Y2=1.12
cc_31 VNB N_VGND_c_382_n 0.0189953f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_383_n 0.0362797f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_384_n 0.0187266f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_385_n 0.00795684f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_386_n 0.200397f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VPB N_C_c_61_n 0.0211471f $X=-0.19 $Y=1.66 $X2=0.592 $Y2=1.618
cc_37 VPB N_C_c_66_n 0.0196207f $X=-0.19 $Y=1.66 $X2=0.675 $Y2=1.885
cc_38 VPB N_C_c_63_n 0.0049966f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.285
cc_39 VPB N_B_c_103_n 0.0161098f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.12
cc_40 VPB N_B_c_100_n 0.0195927f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_41 VPB N_B_c_102_n 0.00253786f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_42 VPB N_A_c_147_n 0.00820914f $X=-0.19 $Y=1.66 $X2=0.675 $Y2=1.885
cc_43 VPB N_A_c_151_n 0.0244819f $X=-0.19 $Y=1.66 $X2=0.675 $Y2=2.46
cc_44 VPB N_A_27_74#_c_199_n 0.0167734f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_45 VPB N_A_27_74#_c_200_n 0.0164424f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.285
cc_46 VPB N_A_27_74#_c_192_n 0.0151944f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB N_A_27_74#_c_202_n 0.0351085f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 VPB N_A_27_74#_c_203_n 0.0163805f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 VPB N_A_27_74#_c_198_n 0.0144913f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_298_n 0.00943661f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_51 VPB N_VPWR_c_299_n 0.0147428f $X=-0.19 $Y=1.66 $X2=0.592 $Y2=1.285
cc_52 VPB N_VPWR_c_300_n 0.0445933f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.285
cc_53 VPB N_VPWR_c_301_n 0.0521687f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_302_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.295
cc_55 VPB N_VPWR_c_303_n 0.0221952f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_297_n 0.089671f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_X_c_337_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_58 VPB N_X_c_338_n 0.0134285f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.285
cc_59 VPB N_X_c_339_n 0.00183475f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB X 0.00753623f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 N_C_c_66_n N_B_c_103_n 0.0535209f $X=0.675 $Y=1.885 $X2=-0.19 $Y2=-0.245
cc_62 N_C_c_62_n N_B_c_99_n 3.44629e-19 $X=0.6 $Y=1.285 $X2=0 $Y2=0
cc_63 N_C_c_63_n N_B_c_99_n 2.2459e-19 $X=0.6 $Y=1.285 $X2=0 $Y2=0
cc_64 N_C_c_64_n N_B_c_99_n 0.0169682f $X=0.592 $Y=1.12 $X2=0 $Y2=0
cc_65 N_C_c_61_n N_B_c_100_n 0.0199009f $X=0.592 $Y=1.618 $X2=0 $Y2=0
cc_66 N_C_c_62_n N_B_c_101_n 0.0199009f $X=0.6 $Y=1.285 $X2=0 $Y2=0
cc_67 N_C_c_63_n N_B_c_101_n 0.00405211f $X=0.6 $Y=1.285 $X2=0 $Y2=0
cc_68 N_C_c_61_n N_B_c_102_n 6.25805e-19 $X=0.592 $Y=1.618 $X2=0 $Y2=0
cc_69 N_C_c_66_n N_B_c_102_n 0.00412162f $X=0.675 $Y=1.885 $X2=0 $Y2=0
cc_70 N_C_c_62_n N_B_c_102_n 7.27895e-19 $X=0.6 $Y=1.285 $X2=0 $Y2=0
cc_71 N_C_c_63_n N_B_c_102_n 0.0529675f $X=0.6 $Y=1.285 $X2=0 $Y2=0
cc_72 N_C_c_64_n N_A_27_74#_c_191_n 0.00889707f $X=0.592 $Y=1.12 $X2=0 $Y2=0
cc_73 N_C_c_61_n N_A_27_74#_c_192_n 0.00282974f $X=0.592 $Y=1.618 $X2=0 $Y2=0
cc_74 N_C_c_66_n N_A_27_74#_c_192_n 0.00212559f $X=0.675 $Y=1.885 $X2=0 $Y2=0
cc_75 N_C_c_63_n N_A_27_74#_c_192_n 0.0510277f $X=0.6 $Y=1.285 $X2=0 $Y2=0
cc_76 N_C_c_64_n N_A_27_74#_c_192_n 0.0212678f $X=0.592 $Y=1.12 $X2=0 $Y2=0
cc_77 N_C_c_66_n N_A_27_74#_c_202_n 0.0129179f $X=0.675 $Y=1.885 $X2=0 $Y2=0
cc_78 N_C_c_62_n N_A_27_74#_c_211_n 0.00123205f $X=0.6 $Y=1.285 $X2=0 $Y2=0
cc_79 N_C_c_63_n N_A_27_74#_c_211_n 0.028434f $X=0.6 $Y=1.285 $X2=0 $Y2=0
cc_80 N_C_c_64_n N_A_27_74#_c_211_n 0.0093151f $X=0.592 $Y=1.12 $X2=0 $Y2=0
cc_81 N_C_c_64_n N_A_27_74#_c_193_n 8.22913e-19 $X=0.592 $Y=1.12 $X2=0 $Y2=0
cc_82 N_C_c_63_n N_A_27_74#_c_197_n 7.54612e-19 $X=0.6 $Y=1.285 $X2=0 $Y2=0
cc_83 N_C_c_64_n N_A_27_74#_c_197_n 0.00348058f $X=0.592 $Y=1.12 $X2=0 $Y2=0
cc_84 N_C_c_61_n N_A_27_74#_c_203_n 0.00160893f $X=0.592 $Y=1.618 $X2=0 $Y2=0
cc_85 N_C_c_66_n N_A_27_74#_c_203_n 0.00262461f $X=0.675 $Y=1.885 $X2=0 $Y2=0
cc_86 N_C_c_63_n N_A_27_74#_c_203_n 0.0119028f $X=0.6 $Y=1.285 $X2=0 $Y2=0
cc_87 N_C_c_66_n N_VPWR_c_301_n 0.00445602f $X=0.675 $Y=1.885 $X2=0 $Y2=0
cc_88 N_C_c_66_n N_VPWR_c_297_n 0.00862094f $X=0.675 $Y=1.885 $X2=0 $Y2=0
cc_89 N_C_c_64_n N_VGND_c_379_n 0.00525591f $X=0.592 $Y=1.12 $X2=0 $Y2=0
cc_90 N_C_c_64_n N_VGND_c_382_n 0.00434272f $X=0.592 $Y=1.12 $X2=0 $Y2=0
cc_91 N_C_c_64_n N_VGND_c_386_n 0.00437823f $X=0.592 $Y=1.12 $X2=0 $Y2=0
cc_92 N_B_c_99_n N_A_M1004_g 0.0226312f $X=1.17 $Y=1.13 $X2=0 $Y2=0
cc_93 N_B_c_101_n N_A_M1004_g 0.0182474f $X=1.17 $Y=1.295 $X2=0 $Y2=0
cc_94 N_B_c_102_n N_A_M1004_g 7.88302e-19 $X=1.17 $Y=1.295 $X2=0 $Y2=0
cc_95 N_B_c_100_n N_A_c_147_n 0.0182474f $X=1.17 $Y=1.635 $X2=0 $Y2=0
cc_96 N_B_c_102_n N_A_c_147_n 0.00163762f $X=1.17 $Y=1.295 $X2=0 $Y2=0
cc_97 N_B_c_103_n N_A_c_151_n 0.0293813f $X=1.095 $Y=1.885 $X2=0 $Y2=0
cc_98 N_B_c_100_n N_A_c_151_n 0.00223184f $X=1.17 $Y=1.635 $X2=0 $Y2=0
cc_99 N_B_c_102_n N_A_c_151_n 0.0113634f $X=1.17 $Y=1.295 $X2=0 $Y2=0
cc_100 N_B_c_101_n A 0.00225967f $X=1.17 $Y=1.295 $X2=0 $Y2=0
cc_101 N_B_c_102_n A 0.0233956f $X=1.17 $Y=1.295 $X2=0 $Y2=0
cc_102 N_B_c_99_n N_A_27_74#_c_191_n 8.22365e-19 $X=1.17 $Y=1.13 $X2=0 $Y2=0
cc_103 N_B_c_103_n N_A_27_74#_c_202_n 0.00122402f $X=1.095 $Y=1.885 $X2=0 $Y2=0
cc_104 N_B_c_99_n N_A_27_74#_c_211_n 0.00936587f $X=1.17 $Y=1.13 $X2=0 $Y2=0
cc_105 N_B_c_101_n N_A_27_74#_c_211_n 3.45553e-19 $X=1.17 $Y=1.295 $X2=0 $Y2=0
cc_106 N_B_c_102_n N_A_27_74#_c_211_n 0.0122553f $X=1.17 $Y=1.295 $X2=0 $Y2=0
cc_107 N_B_c_99_n N_A_27_74#_c_193_n 0.00804273f $X=1.17 $Y=1.13 $X2=0 $Y2=0
cc_108 N_B_c_99_n N_A_27_74#_c_226_n 0.0025058f $X=1.17 $Y=1.13 $X2=0 $Y2=0
cc_109 N_B_c_101_n N_A_27_74#_c_226_n 6.74766e-19 $X=1.17 $Y=1.295 $X2=0 $Y2=0
cc_110 N_B_c_102_n N_A_27_74#_c_226_n 0.00901973f $X=1.17 $Y=1.295 $X2=0 $Y2=0
cc_111 N_B_c_102_n A_234_392# 0.0131191f $X=1.17 $Y=1.295 $X2=-0.19 $Y2=-0.245
cc_112 N_B_c_103_n N_VPWR_c_298_n 0.00173122f $X=1.095 $Y=1.885 $X2=0 $Y2=0
cc_113 N_B_c_102_n N_VPWR_c_298_n 0.0389709f $X=1.17 $Y=1.295 $X2=0 $Y2=0
cc_114 N_B_c_103_n N_VPWR_c_301_n 0.00303293f $X=1.095 $Y=1.885 $X2=0 $Y2=0
cc_115 N_B_c_102_n N_VPWR_c_301_n 0.00909385f $X=1.17 $Y=1.295 $X2=0 $Y2=0
cc_116 N_B_c_103_n N_VPWR_c_297_n 0.00372936f $X=1.095 $Y=1.885 $X2=0 $Y2=0
cc_117 N_B_c_102_n N_VPWR_c_297_n 0.0106888f $X=1.17 $Y=1.295 $X2=0 $Y2=0
cc_118 N_B_c_99_n N_VGND_c_379_n 0.00380067f $X=1.17 $Y=1.13 $X2=0 $Y2=0
cc_119 N_B_c_99_n N_VGND_c_383_n 0.00479783f $X=1.17 $Y=1.13 $X2=0 $Y2=0
cc_120 N_B_c_99_n N_VGND_c_386_n 0.00434877f $X=1.17 $Y=1.13 $X2=0 $Y2=0
cc_121 N_A_c_147_n N_A_27_74#_c_199_n 0.00359537f $X=1.665 $Y=1.795 $X2=0 $Y2=0
cc_122 N_A_c_151_n N_A_27_74#_c_199_n 0.0129424f $X=1.665 $Y=1.885 $X2=0 $Y2=0
cc_123 N_A_M1004_g N_A_27_74#_M1005_g 0.0147473f $X=1.65 $Y=0.69 $X2=0 $Y2=0
cc_124 N_A_c_149_n N_A_27_74#_M1005_g 0.00187922f $X=1.74 $Y=1.385 $X2=0 $Y2=0
cc_125 N_A_M1004_g N_A_27_74#_c_193_n 0.00230442f $X=1.65 $Y=0.69 $X2=0 $Y2=0
cc_126 N_A_M1004_g N_A_27_74#_c_234_n 0.0131982f $X=1.65 $Y=0.69 $X2=0 $Y2=0
cc_127 A N_A_27_74#_c_234_n 0.0191834f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_128 N_A_c_149_n N_A_27_74#_c_234_n 9.50988e-19 $X=1.74 $Y=1.385 $X2=0 $Y2=0
cc_129 N_A_M1004_g N_A_27_74#_c_194_n 0.00420198f $X=1.65 $Y=0.69 $X2=0 $Y2=0
cc_130 A N_A_27_74#_c_194_n 0.00916736f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_131 N_A_c_149_n N_A_27_74#_c_194_n 5.96051e-19 $X=1.74 $Y=1.385 $X2=0 $Y2=0
cc_132 N_A_c_147_n N_A_27_74#_c_195_n 0.00192809f $X=1.665 $Y=1.795 $X2=0 $Y2=0
cc_133 A N_A_27_74#_c_195_n 0.0211265f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_134 N_A_c_149_n N_A_27_74#_c_195_n 0.00163329f $X=1.74 $Y=1.385 $X2=0 $Y2=0
cc_135 N_A_c_147_n N_A_27_74#_c_198_n 0.00692915f $X=1.665 $Y=1.795 $X2=0 $Y2=0
cc_136 A N_A_27_74#_c_198_n 2.73033e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_137 N_A_c_149_n N_A_27_74#_c_198_n 0.0132233f $X=1.74 $Y=1.385 $X2=0 $Y2=0
cc_138 N_A_c_151_n N_VPWR_c_298_n 0.0211204f $X=1.665 $Y=1.885 $X2=0 $Y2=0
cc_139 A N_VPWR_c_298_n 0.00810648f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_140 N_A_c_149_n N_VPWR_c_298_n 0.00105498f $X=1.74 $Y=1.385 $X2=0 $Y2=0
cc_141 N_A_c_151_n N_VPWR_c_301_n 0.00413917f $X=1.665 $Y=1.885 $X2=0 $Y2=0
cc_142 N_A_c_151_n N_VPWR_c_297_n 0.00818781f $X=1.665 $Y=1.885 $X2=0 $Y2=0
cc_143 N_A_c_151_n N_X_c_337_n 2.93406e-19 $X=1.665 $Y=1.885 $X2=0 $Y2=0
cc_144 N_A_M1004_g N_X_c_333_n 0.0010435f $X=1.65 $Y=0.69 $X2=0 $Y2=0
cc_145 N_A_c_151_n N_X_c_339_n 6.37522e-19 $X=1.665 $Y=1.885 $X2=0 $Y2=0
cc_146 N_A_M1004_g N_VGND_c_383_n 0.0159537f $X=1.65 $Y=0.69 $X2=0 $Y2=0
cc_147 N_A_M1004_g N_VGND_c_386_n 0.00374187f $X=1.65 $Y=0.69 $X2=0 $Y2=0
cc_148 N_A_27_74#_c_199_n N_VPWR_c_298_n 0.0128259f $X=2.275 $Y=1.765 $X2=0
+ $Y2=0
cc_149 N_A_27_74#_c_200_n N_VPWR_c_300_n 0.0212063f $X=2.725 $Y=1.765 $X2=0
+ $Y2=0
cc_150 N_A_27_74#_c_202_n N_VPWR_c_301_n 0.0145938f $X=0.45 $Y=2.815 $X2=0 $Y2=0
cc_151 N_A_27_74#_c_199_n N_VPWR_c_303_n 0.00445602f $X=2.275 $Y=1.765 $X2=0
+ $Y2=0
cc_152 N_A_27_74#_c_200_n N_VPWR_c_303_n 0.00445602f $X=2.725 $Y=1.765 $X2=0
+ $Y2=0
cc_153 N_A_27_74#_c_199_n N_VPWR_c_297_n 0.00859686f $X=2.275 $Y=1.765 $X2=0
+ $Y2=0
cc_154 N_A_27_74#_c_200_n N_VPWR_c_297_n 0.00860769f $X=2.725 $Y=1.765 $X2=0
+ $Y2=0
cc_155 N_A_27_74#_c_202_n N_VPWR_c_297_n 0.0120466f $X=0.45 $Y=2.815 $X2=0 $Y2=0
cc_156 N_A_27_74#_c_199_n N_X_c_337_n 0.0134506f $X=2.275 $Y=1.765 $X2=0 $Y2=0
cc_157 N_A_27_74#_c_200_n N_X_c_337_n 0.0165744f $X=2.725 $Y=1.765 $X2=0 $Y2=0
cc_158 N_A_27_74#_M1005_g N_X_c_333_n 0.00983911f $X=2.365 $Y=0.74 $X2=0 $Y2=0
cc_159 N_A_27_74#_M1009_g N_X_c_333_n 0.0131993f $X=2.795 $Y=0.74 $X2=0 $Y2=0
cc_160 N_A_27_74#_c_200_n N_X_c_338_n 0.0135579f $X=2.725 $Y=1.765 $X2=0 $Y2=0
cc_161 N_A_27_74#_c_196_n N_X_c_338_n 0.010734f $X=2.65 $Y=1.465 $X2=0 $Y2=0
cc_162 N_A_27_74#_c_198_n N_X_c_338_n 0.00184626f $X=2.725 $Y=1.532 $X2=0 $Y2=0
cc_163 N_A_27_74#_c_199_n N_X_c_339_n 0.00414322f $X=2.275 $Y=1.765 $X2=0 $Y2=0
cc_164 N_A_27_74#_c_200_n N_X_c_339_n 9.3899e-19 $X=2.725 $Y=1.765 $X2=0 $Y2=0
cc_165 N_A_27_74#_c_196_n N_X_c_339_n 0.0276943f $X=2.65 $Y=1.465 $X2=0 $Y2=0
cc_166 N_A_27_74#_c_198_n N_X_c_339_n 0.00792231f $X=2.725 $Y=1.532 $X2=0 $Y2=0
cc_167 N_A_27_74#_M1009_g N_X_c_334_n 0.0132378f $X=2.795 $Y=0.74 $X2=0 $Y2=0
cc_168 N_A_27_74#_c_196_n N_X_c_334_n 0.00496499f $X=2.65 $Y=1.465 $X2=0 $Y2=0
cc_169 N_A_27_74#_M1005_g N_X_c_335_n 0.00237641f $X=2.365 $Y=0.74 $X2=0 $Y2=0
cc_170 N_A_27_74#_M1009_g N_X_c_335_n 9.7541e-19 $X=2.795 $Y=0.74 $X2=0 $Y2=0
cc_171 N_A_27_74#_c_194_n N_X_c_335_n 0.00787895f $X=2.16 $Y=1.3 $X2=0 $Y2=0
cc_172 N_A_27_74#_c_196_n N_X_c_335_n 0.0276081f $X=2.65 $Y=1.465 $X2=0 $Y2=0
cc_173 N_A_27_74#_c_198_n N_X_c_335_n 0.00232957f $X=2.725 $Y=1.532 $X2=0 $Y2=0
cc_174 N_A_27_74#_c_200_n X 0.00116193f $X=2.725 $Y=1.765 $X2=0 $Y2=0
cc_175 N_A_27_74#_M1009_g X 0.0104281f $X=2.795 $Y=0.74 $X2=0 $Y2=0
cc_176 N_A_27_74#_c_196_n X 0.0246264f $X=2.65 $Y=1.465 $X2=0 $Y2=0
cc_177 N_A_27_74#_c_198_n X 0.00607246f $X=2.725 $Y=1.532 $X2=0 $Y2=0
cc_178 N_A_27_74#_c_211_n N_VGND_M1008_d 0.0140026f $X=1.2 $Y=0.865 $X2=-0.19
+ $Y2=-0.245
cc_179 N_A_27_74#_c_234_n N_VGND_M1004_d 0.0157029f $X=2.075 $Y=0.875 $X2=0
+ $Y2=0
cc_180 N_A_27_74#_c_194_n N_VGND_M1004_d 0.00326802f $X=2.16 $Y=1.3 $X2=0 $Y2=0
cc_181 N_A_27_74#_c_191_n N_VGND_c_379_n 0.0102838f $X=0.28 $Y=0.65 $X2=0 $Y2=0
cc_182 N_A_27_74#_c_211_n N_VGND_c_379_n 0.0295211f $X=1.2 $Y=0.865 $X2=0 $Y2=0
cc_183 N_A_27_74#_c_193_n N_VGND_c_379_n 0.010199f $X=1.365 $Y=0.78 $X2=0 $Y2=0
cc_184 N_A_27_74#_M1009_g N_VGND_c_381_n 0.0118431f $X=2.795 $Y=0.74 $X2=0 $Y2=0
cc_185 N_A_27_74#_c_191_n N_VGND_c_382_n 0.0153852f $X=0.28 $Y=0.65 $X2=0 $Y2=0
cc_186 N_A_27_74#_M1005_g N_VGND_c_383_n 0.00411273f $X=2.365 $Y=0.74 $X2=0
+ $Y2=0
cc_187 N_A_27_74#_c_193_n N_VGND_c_383_n 0.0253687f $X=1.365 $Y=0.78 $X2=0 $Y2=0
cc_188 N_A_27_74#_c_234_n N_VGND_c_383_n 0.0353491f $X=2.075 $Y=0.875 $X2=0
+ $Y2=0
cc_189 N_A_27_74#_c_198_n N_VGND_c_383_n 2.76634e-19 $X=2.725 $Y=1.532 $X2=0
+ $Y2=0
cc_190 N_A_27_74#_M1005_g N_VGND_c_384_n 0.00434272f $X=2.365 $Y=0.74 $X2=0
+ $Y2=0
cc_191 N_A_27_74#_M1009_g N_VGND_c_384_n 0.00434272f $X=2.795 $Y=0.74 $X2=0
+ $Y2=0
cc_192 N_A_27_74#_M1005_g N_VGND_c_386_n 0.00822235f $X=2.365 $Y=0.74 $X2=0
+ $Y2=0
cc_193 N_A_27_74#_M1009_g N_VGND_c_386_n 0.00823934f $X=2.795 $Y=0.74 $X2=0
+ $Y2=0
cc_194 N_A_27_74#_c_191_n N_VGND_c_386_n 0.0127091f $X=0.28 $Y=0.65 $X2=0 $Y2=0
cc_195 N_A_27_74#_c_211_n N_VGND_c_386_n 0.0121035f $X=1.2 $Y=0.865 $X2=0 $Y2=0
cc_196 N_A_27_74#_c_193_n N_VGND_c_386_n 0.0119539f $X=1.365 $Y=0.78 $X2=0 $Y2=0
cc_197 N_A_27_74#_c_234_n N_VGND_c_386_n 0.00729135f $X=2.075 $Y=0.875 $X2=0
+ $Y2=0
cc_198 N_VPWR_c_298_n N_X_c_337_n 0.0534912f $X=1.89 $Y=2.105 $X2=0 $Y2=0
cc_199 N_VPWR_c_300_n N_X_c_337_n 0.0323093f $X=3 $Y=2.225 $X2=0 $Y2=0
cc_200 N_VPWR_c_303_n N_X_c_337_n 0.014552f $X=2.835 $Y=3.33 $X2=0 $Y2=0
cc_201 N_VPWR_c_297_n N_X_c_337_n 0.0119791f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_202 N_VPWR_M1007_d N_X_c_338_n 0.00429065f $X=2.8 $Y=1.84 $X2=0 $Y2=0
cc_203 N_VPWR_c_300_n N_X_c_338_n 0.0264075f $X=3 $Y=2.225 $X2=0 $Y2=0
cc_204 N_VPWR_c_298_n N_X_c_339_n 0.00168189f $X=1.89 $Y=2.105 $X2=0 $Y2=0
cc_205 N_X_c_334_n N_VGND_M1009_s 0.00470604f $X=3.005 $Y=1.045 $X2=0 $Y2=0
cc_206 N_X_c_333_n N_VGND_c_381_n 0.0173003f $X=2.58 $Y=0.515 $X2=0 $Y2=0
cc_207 N_X_c_334_n N_VGND_c_381_n 0.0270821f $X=3.005 $Y=1.045 $X2=0 $Y2=0
cc_208 N_X_c_333_n N_VGND_c_383_n 0.0102333f $X=2.58 $Y=0.515 $X2=0 $Y2=0
cc_209 N_X_c_333_n N_VGND_c_384_n 0.0144922f $X=2.58 $Y=0.515 $X2=0 $Y2=0
cc_210 N_X_c_333_n N_VGND_c_386_n 0.0118826f $X=2.58 $Y=0.515 $X2=0 $Y2=0
