# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_ls__nand4_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.800000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.885000 1.350000 4.215000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.680000 1.350000 3.715000 1.780000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.430000 1.350000 2.440000 1.780000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.350000 1.090000 1.780000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  1.633200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.635000 1.950000 4.675000 2.120000 ;
        RECT 0.635000 2.120000 0.900000 2.980000 ;
        RECT 1.570000 2.120000 1.900000 2.980000 ;
        RECT 2.830000 2.120000 3.160000 2.980000 ;
        RECT 3.840000 2.120000 4.675000 2.150000 ;
        RECT 3.840000 2.150000 4.125000 2.980000 ;
        RECT 3.845000 0.645000 4.175000 1.010000 ;
        RECT 3.845000 1.010000 4.675000 1.180000 ;
        RECT 4.445000 1.180000 4.675000 1.950000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.800000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.800000 0.085000 ;
      RECT 0.000000  3.245000 4.800000 3.415000 ;
      RECT 0.115000  0.350000 0.445000 1.010000 ;
      RECT 0.115000  1.010000 1.315000 1.180000 ;
      RECT 0.115000  1.950000 0.450000 3.245000 ;
      RECT 0.615000  0.085000 0.945000 0.840000 ;
      RECT 1.070000  2.290000 1.400000 3.245000 ;
      RECT 1.145000  0.255000 2.325000 0.425000 ;
      RECT 1.145000  0.425000 1.315000 1.010000 ;
      RECT 1.495000  0.595000 1.825000 1.010000 ;
      RECT 1.495000  1.010000 3.315000 1.180000 ;
      RECT 1.995000  0.425000 2.325000 0.840000 ;
      RECT 2.080000  2.290000 2.650000 3.245000 ;
      RECT 2.555000  0.255000 4.675000 0.425000 ;
      RECT 2.555000  0.425000 2.815000 0.840000 ;
      RECT 2.985000  0.645000 3.315000 1.010000 ;
      RECT 3.330000  2.290000 3.660000 3.245000 ;
      RECT 3.485000  0.425000 3.675000 1.130000 ;
      RECT 4.295000  2.320000 4.625000 3.245000 ;
      RECT 4.345000  0.425000 4.675000 0.840000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
  END
END sky130_fd_sc_ls__nand4_2
