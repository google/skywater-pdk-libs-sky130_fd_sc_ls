* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__dfxtp_1 CLK D VGND VNB VPB VPWR Q
X0 VPWR a_561_463# a_713_458# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X1 VPWR a_1210_314# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X2 a_713_458# a_206_368# a_1011_424# VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X3 a_561_463# a_27_74# a_668_503# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 a_1168_124# a_1210_314# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_713_458# a_27_74# a_1011_424# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X6 a_561_463# a_206_368# a_731_101# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_1011_424# a_27_74# a_1168_124# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_27_74# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X9 a_454_503# a_206_368# a_561_463# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X10 VGND D a_454_503# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 a_1118_508# a_1210_314# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X12 a_454_503# a_27_74# a_561_463# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 VGND a_561_463# a_713_458# VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X14 a_731_101# a_713_458# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 a_1210_314# a_1011_424# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X16 VPWR a_27_74# a_206_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X17 a_27_74# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X18 VGND a_27_74# a_206_368# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X19 a_1011_424# a_206_368# a_1118_508# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X20 VPWR D a_454_503# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X21 a_668_503# a_713_458# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X22 VGND a_1210_314# Q VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X23 a_1210_314# a_1011_424# VGND VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
.ends
