* NGSPICE file created from sky130_fd_sc_ls__sdlclkp_1.ext - technology: sky130A

.subckt sky130_fd_sc_ls__sdlclkp_1 CLK GATE SCE VGND VNB VPB VPWR GCLK
M1000 a_318_74# a_288_48# VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=1.3368e+12p ps=1.136e+07u
M1001 VPWR a_709_54# a_722_492# VPB phighvt w=420000u l=150000u
+  ad=1.92175e+12p pd=1.454e+07u as=1.008e+11p ps=1.32e+06u
M1002 VGND CLK a_288_48# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.072e+11p ps=2.04e+06u
M1003 a_1166_94# CLK VGND VNB nshort w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1004 a_318_74# a_288_48# VPWR VPB phighvt w=840000u l=150000u
+  ad=2.478e+11p pd=2.27e+06u as=0p ps=0u
M1005 a_1238_94# a_709_54# a_1166_94# VNB nshort w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=0p ps=0u
M1006 a_566_74# a_318_74# a_114_112# VPB phighvt w=840000u l=150000u
+  ad=3.10975e+11p pd=2.74e+06u as=4.956e+11p ps=4.54e+06u
M1007 a_709_54# a_566_74# VGND VNB nshort w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1008 VGND GATE a_114_112# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=4.4825e+11p ps=3.83e+06u
M1009 a_114_112# SCE VGND VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_1238_94# CLK VPWR VPB phighvt w=840000u l=150000u
+  ad=2.52e+11p pd=2.28e+06u as=0p ps=0u
M1011 GCLK a_1238_94# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=4.256e+11p pd=3e+06u as=0p ps=0u
M1012 a_667_80# a_318_74# a_566_74# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.846e+11p ps=1.81e+06u
M1013 VGND a_709_54# a_667_80# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_116_424# SCE VPWR VPB phighvt w=840000u l=150000u
+  ad=2.016e+11p pd=2.16e+06u as=0p ps=0u
M1015 a_566_74# a_288_48# a_114_112# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_709_54# a_566_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=0p ps=0u
M1017 VPWR a_709_54# a_1238_94# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 GCLK a_1238_94# VGND VNB nshort w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1019 a_114_112# GATE a_116_424# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_722_492# a_288_48# a_566_74# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPWR CLK a_288_48# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=2.478e+11p ps=2.27e+06u
.ends

