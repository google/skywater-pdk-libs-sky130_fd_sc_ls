* File: sky130_fd_sc_ls__nand4bb_4.pex.spice
* Created: Wed Sep  2 11:13:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__NAND4BB_4%A_N 3 6 7 9 10 12 16 18 21
c49 21 0 1.99278e-19 $X=0.605 $Y=1.615
c50 10 0 3.39396e-20 $X=0.955 $Y=2.045
r51 21 23 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.595 $Y=1.615
+ $X2=0.595 $Y2=1.45
r52 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.605
+ $Y=1.615 $X2=0.605 $Y2=1.615
r53 18 22 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=0.72 $Y=1.615
+ $X2=0.605 $Y2=1.615
r54 10 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.955 $Y=2.045
+ $X2=0.955 $Y2=1.97
r55 10 12 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.955 $Y=2.045
+ $X2=0.955 $Y2=2.54
r56 7 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.505 $Y=2.045
+ $X2=0.505 $Y2=1.97
r57 7 9 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.505 $Y=2.045
+ $X2=0.505 $Y2=2.54
r58 6 16 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=0.595 $Y=1.97
+ $X2=0.955 $Y2=1.97
r59 6 13 46.1489 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=0.595 $Y=1.97 $X2=0.505
+ $Y2=1.97
r60 5 21 1.64869 $w=3.5e-07 $l=1e-08 $layer=POLY_cond $X=0.595 $Y=1.625
+ $X2=0.595 $Y2=1.615
r61 5 6 44.5147 $w=3.5e-07 $l=2.7e-07 $layer=POLY_cond $X=0.595 $Y=1.625
+ $X2=0.595 $Y2=1.895
r62 3 23 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=0.495 $Y=0.94
+ $X2=0.495 $Y2=1.45
.ends

.subckt PM_SKY130_FD_SC_LS__NAND4BB_4%B_N 3 5 6 7 9 10 12 13 17
c58 10 0 1.98429e-19 $X=1.855 $Y=2.045
c59 7 0 5.52958e-20 $X=1.405 $Y=2.045
r60 15 17 25.0462 $w=4.33e-07 $l=2.25e-07 $layer=POLY_cond $X=1.405 $Y=1.775
+ $X2=1.63 $Y2=1.775
r61 13 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.63
+ $Y=1.715 $X2=1.63 $Y2=1.715
r62 10 17 25.0462 $w=4.33e-07 $l=3.65582e-07 $layer=POLY_cond $X=1.855 $Y=2.045
+ $X2=1.63 $Y2=1.775
r63 10 12 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.855 $Y=2.045
+ $X2=1.855 $Y2=2.54
r64 7 15 27.8114 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=1.405 $Y=2.045
+ $X2=1.405 $Y2=1.775
r65 7 9 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.405 $Y=2.045
+ $X2=1.405 $Y2=2.54
r66 5 15 31.9371 $w=4.33e-07 $l=2.35743e-07 $layer=POLY_cond $X=1.315 $Y=1.58
+ $X2=1.405 $Y2=1.775
r67 5 6 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=1.315 $Y=1.58
+ $X2=1.16 $Y2=1.58
r68 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.085 $Y=1.505
+ $X2=1.16 $Y2=1.58
r69 1 3 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=1.085 $Y=1.505
+ $X2=1.085 $Y2=0.94
.ends

.subckt PM_SKY130_FD_SC_LS__NAND4BB_4%A_27_114# 1 2 7 9 10 12 13 15 16 18 19 21
+ 22 24 27 29 30 31 33 34 35 37 38 39 40 44 47 49 50 55 60 61
c159 31 0 1.90572e-19 $X=3.975 $Y=1.765
c160 27 0 1.79504e-19 $X=3.635 $Y=0.74
c161 19 0 7.06753e-20 $X=3.205 $Y=1.22
c162 13 0 7.06753e-20 $X=2.765 $Y=1.22
r163 68 69 31.5419 $w=4.89e-07 $l=3.2e-07 $layer=POLY_cond $X=3.205 $Y=1.492
+ $X2=3.525 $Y2=1.492
r164 67 68 12.8139 $w=4.89e-07 $l=1.3e-07 $layer=POLY_cond $X=3.075 $Y=1.492
+ $X2=3.205 $Y2=1.492
r165 62 63 34.0061 $w=4.89e-07 $l=3.45e-07 $layer=POLY_cond $X=2.23 $Y=1.492
+ $X2=2.575 $Y2=1.492
r166 56 67 7.39264 $w=4.89e-07 $l=7.5e-08 $layer=POLY_cond $X=3 $Y=1.492
+ $X2=3.075 $Y2=1.492
r167 56 65 23.1636 $w=4.89e-07 $l=2.35e-07 $layer=POLY_cond $X=3 $Y=1.492
+ $X2=2.765 $Y2=1.492
r168 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3
+ $Y=1.385 $X2=3 $Y2=1.385
r169 53 65 10.3497 $w=4.89e-07 $l=1.05e-07 $layer=POLY_cond $X=2.66 $Y=1.492
+ $X2=2.765 $Y2=1.492
r170 53 63 8.37832 $w=4.89e-07 $l=8.5e-08 $layer=POLY_cond $X=2.66 $Y=1.492
+ $X2=2.575 $Y2=1.492
r171 52 55 11.5244 $w=3.38e-07 $l=3.4e-07 $layer=LI1_cond $X=2.66 $Y=1.38 $X2=3
+ $Y2=1.38
r172 52 53 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.66
+ $Y=1.385 $X2=2.66 $Y2=1.385
r173 50 61 14.4036 $w=3.38e-07 $l=3.4e-07 $layer=LI1_cond $X=2.495 $Y=1.38
+ $X2=2.155 $Y2=1.38
r174 50 52 5.59274 $w=3.38e-07 $l=1.65e-07 $layer=LI1_cond $X=2.495 $Y=1.38
+ $X2=2.66 $Y2=1.38
r175 49 61 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.76 $Y=1.295
+ $X2=2.155 $Y2=1.295
r176 47 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.675 $Y=1.21
+ $X2=1.76 $Y2=1.295
r177 46 47 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=1.675 $Y=0.83
+ $X2=1.675 $Y2=1.21
r178 42 44 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=0.73 $Y=2.12
+ $X2=0.73 $Y2=2.265
r179 41 59 4.8908 $w=1.7e-07 $l=1.98605e-07 $layer=LI1_cond $X=0.445 $Y=0.745
+ $X2=0.272 $Y2=0.69
r180 40 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.59 $Y=0.745
+ $X2=1.675 $Y2=0.83
r181 40 41 74.7005 $w=1.68e-07 $l=1.145e-06 $layer=LI1_cond $X=1.59 $Y=0.745
+ $X2=0.445 $Y2=0.745
r182 38 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.645 $Y=2.035
+ $X2=0.73 $Y2=2.12
r183 38 39 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.645 $Y=2.035
+ $X2=0.27 $Y2=2.035
r184 37 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.185 $Y=1.95
+ $X2=0.27 $Y2=2.035
r185 37 60 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.185 $Y=1.95
+ $X2=0.185 $Y2=1.28
r186 35 60 8.71323 $w=3.43e-07 $l=1.72e-07 $layer=LI1_cond $X=0.272 $Y=1.108
+ $X2=0.272 $Y2=1.28
r187 34 59 3.00312 $w=3.45e-07 $l=1.4e-07 $layer=LI1_cond $X=0.272 $Y=0.83
+ $X2=0.272 $Y2=0.69
r188 34 35 9.28635 $w=3.43e-07 $l=2.78e-07 $layer=LI1_cond $X=0.272 $Y=0.83
+ $X2=0.272 $Y2=1.108
r189 31 33 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.975 $Y=1.765
+ $X2=3.975 $Y2=2.4
r190 29 31 26.9307 $w=1.5e-07 $l=1.53542e-07 $layer=POLY_cond $X=3.885 $Y=1.65
+ $X2=3.975 $Y2=1.765
r191 29 30 89.734 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=3.885 $Y=1.65
+ $X2=3.71 $Y2=1.65
r192 25 30 32.7723 $w=4.89e-07 $l=1.9187e-07 $layer=POLY_cond $X=3.635 $Y=1.492
+ $X2=3.71 $Y2=1.65
r193 25 69 10.8425 $w=4.89e-07 $l=1.1e-07 $layer=POLY_cond $X=3.635 $Y=1.492
+ $X2=3.525 $Y2=1.492
r194 25 27 299.968 $w=1.5e-07 $l=5.85e-07 $layer=POLY_cond $X=3.635 $Y=1.325
+ $X2=3.635 $Y2=0.74
r195 22 69 30.8469 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=3.525 $Y=1.765
+ $X2=3.525 $Y2=1.492
r196 22 24 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.525 $Y=1.765
+ $X2=3.525 $Y2=2.4
r197 19 68 30.8469 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=3.205 $Y=1.22
+ $X2=3.205 $Y2=1.492
r198 19 21 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.205 $Y=1.22
+ $X2=3.205 $Y2=0.74
r199 16 67 30.8469 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=3.075 $Y=1.765
+ $X2=3.075 $Y2=1.492
r200 16 18 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.075 $Y=1.765
+ $X2=3.075 $Y2=2.4
r201 13 65 30.8469 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=2.765 $Y=1.22
+ $X2=2.765 $Y2=1.492
r202 13 15 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.765 $Y=1.22
+ $X2=2.765 $Y2=0.74
r203 10 63 30.8469 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=2.575 $Y=1.765
+ $X2=2.575 $Y2=1.492
r204 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.575 $Y=1.765
+ $X2=2.575 $Y2=2.4
r205 7 62 30.8469 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=2.23 $Y=1.22
+ $X2=2.23 $Y2=1.492
r206 7 9 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.23 $Y=1.22 $X2=2.23
+ $Y2=0.74
r207 2 44 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=0.58
+ $Y=2.12 $X2=0.73 $Y2=2.265
r208 1 59 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.57 $X2=0.28 $Y2=0.715
.ends

.subckt PM_SKY130_FD_SC_LS__NAND4BB_4%A_232_114# 1 2 7 9 10 11 12 14 15 17 18 20
+ 21 23 24 26 27 29 30 32 34 35 36 39 42 43 44 45 50 56 59 72
c177 45 0 1.90572e-19 $X=4.315 $Y=1.555
c178 34 0 2.88513e-19 $X=1.21 $Y=2.05
c179 18 0 6.63463e-21 $X=4.875 $Y=1.765
r180 71 72 14.6061 $w=4.62e-07 $l=1.4e-07 $layer=POLY_cond $X=5.375 $Y=1.475
+ $X2=5.515 $Y2=1.475
r181 68 69 5.21645 $w=4.62e-07 $l=5e-08 $layer=POLY_cond $X=4.875 $Y=1.475
+ $X2=4.925 $Y2=1.475
r182 65 66 7.30303 $w=4.62e-07 $l=7e-08 $layer=POLY_cond $X=4.425 $Y=1.475
+ $X2=4.495 $Y2=1.475
r183 53 56 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=1.21 $Y=1.165
+ $X2=1.315 $Y2=1.165
r184 51 71 20.3442 $w=4.62e-07 $l=1.95e-07 $layer=POLY_cond $X=5.18 $Y=1.475
+ $X2=5.375 $Y2=1.475
r185 51 69 26.6039 $w=4.62e-07 $l=2.55e-07 $layer=POLY_cond $X=5.18 $Y=1.475
+ $X2=4.925 $Y2=1.475
r186 50 51 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=5.18
+ $Y=1.515 $X2=5.18 $Y2=1.515
r187 48 68 39.1234 $w=4.62e-07 $l=3.75e-07 $layer=POLY_cond $X=4.5 $Y=1.475
+ $X2=4.875 $Y2=1.475
r188 48 66 0.521645 $w=4.62e-07 $l=5e-09 $layer=POLY_cond $X=4.5 $Y=1.475
+ $X2=4.495 $Y2=1.475
r189 47 50 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=4.5 $Y=1.555
+ $X2=5.18 $Y2=1.555
r190 47 48 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=4.5
+ $Y=1.515 $X2=4.5 $Y2=1.515
r191 45 63 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=4.23 $Y=1.555
+ $X2=4.23 $Y2=1.805
r192 45 47 8.52808 $w=2.48e-07 $l=1.85e-07 $layer=LI1_cond $X=4.315 $Y=1.555
+ $X2=4.5 $Y2=1.555
r193 43 63 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.145 $Y=1.805
+ $X2=4.23 $Y2=1.805
r194 43 44 131.134 $w=1.68e-07 $l=2.01e-06 $layer=LI1_cond $X=4.145 $Y=1.805
+ $X2=2.135 $Y2=1.805
r195 42 59 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.05 $Y=2.05
+ $X2=2.05 $Y2=2.135
r196 41 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.05 $Y=1.89
+ $X2=2.135 $Y2=1.805
r197 41 42 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=2.05 $Y=1.89
+ $X2=2.05 $Y2=2.05
r198 37 59 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.655 $Y=2.135
+ $X2=2.05 $Y2=2.135
r199 37 39 1.85214 $w=2.78e-07 $l=4.5e-08 $layer=LI1_cond $X=1.655 $Y=2.22
+ $X2=1.655 $Y2=2.265
r200 35 37 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=1.515 $Y=2.135
+ $X2=1.655 $Y2=2.135
r201 35 36 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=1.515 $Y=2.135
+ $X2=1.295 $Y2=2.135
r202 34 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.21 $Y=2.05
+ $X2=1.295 $Y2=2.135
r203 33 53 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.21 $Y=1.33
+ $X2=1.21 $Y2=1.165
r204 33 34 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=1.21 $Y=1.33
+ $X2=1.21 $Y2=2.05
r205 30 72 32.342 $w=4.62e-07 $l=4.31277e-07 $layer=POLY_cond $X=5.825 $Y=1.765
+ $X2=5.515 $Y2=1.475
r206 30 32 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.825 $Y=1.765
+ $X2=5.825 $Y2=2.4
r207 27 72 29.4226 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=5.515 $Y=1.185
+ $X2=5.515 $Y2=1.475
r208 27 29 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=5.515 $Y=1.185
+ $X2=5.515 $Y2=0.74
r209 24 71 29.4226 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=5.375 $Y=1.765
+ $X2=5.375 $Y2=1.475
r210 24 26 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.375 $Y=1.765
+ $X2=5.375 $Y2=2.4
r211 21 69 29.4226 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=4.925 $Y=1.185
+ $X2=4.925 $Y2=1.475
r212 21 23 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=4.925 $Y=1.185
+ $X2=4.925 $Y2=0.74
r213 18 68 29.4226 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=4.875 $Y=1.765
+ $X2=4.875 $Y2=1.475
r214 18 20 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.875 $Y=1.765
+ $X2=4.875 $Y2=2.4
r215 15 66 29.4226 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=4.495 $Y=1.185
+ $X2=4.495 $Y2=1.475
r216 15 17 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=4.495 $Y=1.185
+ $X2=4.495 $Y2=0.74
r217 12 65 29.4226 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=4.425 $Y=1.765
+ $X2=4.425 $Y2=1.475
r218 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.425 $Y=1.765
+ $X2=4.425 $Y2=2.4
r219 10 65 33.1446 $w=4.62e-07 $l=2.56076e-07 $layer=POLY_cond $X=4.335 $Y=1.26
+ $X2=4.425 $Y2=1.475
r220 10 11 99.9894 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=4.335 $Y=1.26
+ $X2=4.14 $Y2=1.26
r221 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.065 $Y=1.185
+ $X2=4.14 $Y2=1.26
r222 7 9 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=4.065 $Y=1.185
+ $X2=4.065 $Y2=0.74
r223 2 39 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=1.48
+ $Y=2.12 $X2=1.63 $Y2=2.265
r224 1 56 182 $w=1.7e-07 $l=6.68019e-07 $layer=licon1_NDIFF $count=1 $X=1.16
+ $Y=0.57 $X2=1.315 $Y2=1.165
.ends

.subckt PM_SKY130_FD_SC_LS__NAND4BB_4%C 1 3 6 8 10 13 15 17 20 22 24 27 36 39 49
+ 52 54
c97 54 0 1.90128e-19 $X=7.075 $Y=1.55
c98 22 0 6.20142e-20 $X=7.725 $Y=1.765
c99 8 0 1.227e-20 $X=6.725 $Y=1.765
r100 49 50 9.04558 $w=3.73e-07 $l=7e-08 $layer=POLY_cond $X=7.725 $Y=1.542
+ $X2=7.795 $Y2=1.542
r101 46 47 11.63 $w=3.73e-07 $l=9e-08 $layer=POLY_cond $X=7.275 $Y=1.542
+ $X2=7.365 $Y2=1.542
r102 45 46 43.9357 $w=3.73e-07 $l=3.4e-07 $layer=POLY_cond $X=6.935 $Y=1.542
+ $X2=7.275 $Y2=1.542
r103 44 45 27.1367 $w=3.73e-07 $l=2.1e-07 $layer=POLY_cond $X=6.725 $Y=1.542
+ $X2=6.935 $Y2=1.542
r104 43 44 28.429 $w=3.73e-07 $l=2.2e-07 $layer=POLY_cond $X=6.505 $Y=1.542
+ $X2=6.725 $Y2=1.542
r105 39 54 3.96409 $w=4.58e-07 $l=1.15e-07 $layer=LI1_cond $X=6.96 $Y=1.55
+ $X2=7.075 $Y2=1.55
r106 39 52 3.96409 $w=4.58e-07 $l=1.15e-07 $layer=LI1_cond $X=6.96 $Y=1.55
+ $X2=6.845 $Y2=1.55
r107 37 49 36.1823 $w=3.73e-07 $l=2.8e-07 $layer=POLY_cond $X=7.445 $Y=1.542
+ $X2=7.725 $Y2=1.542
r108 37 47 10.3378 $w=3.73e-07 $l=8e-08 $layer=POLY_cond $X=7.445 $Y=1.542
+ $X2=7.365 $Y2=1.542
r109 36 54 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=7.445 $Y=1.485
+ $X2=7.075 $Y2=1.485
r110 36 37 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.445
+ $Y=1.485 $X2=7.445 $Y2=1.485
r111 32 43 10.3378 $w=3.73e-07 $l=8e-08 $layer=POLY_cond $X=6.425 $Y=1.542
+ $X2=6.505 $Y2=1.542
r112 32 41 19.3834 $w=3.73e-07 $l=1.5e-07 $layer=POLY_cond $X=6.425 $Y=1.542
+ $X2=6.275 $Y2=1.542
r113 31 52 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=6.425 $Y=1.485
+ $X2=6.845 $Y2=1.485
r114 31 32 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.425
+ $Y=1.485 $X2=6.425 $Y2=1.485
r115 25 50 24.162 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=7.795 $Y=1.32
+ $X2=7.795 $Y2=1.542
r116 25 27 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=7.795 $Y=1.32
+ $X2=7.795 $Y2=0.74
r117 22 49 24.162 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=7.725 $Y=1.765
+ $X2=7.725 $Y2=1.542
r118 22 24 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.725 $Y=1.765
+ $X2=7.725 $Y2=2.4
r119 18 47 24.162 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=7.365 $Y=1.32
+ $X2=7.365 $Y2=1.542
r120 18 20 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=7.365 $Y=1.32
+ $X2=7.365 $Y2=0.74
r121 15 46 24.162 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=7.275 $Y=1.765
+ $X2=7.275 $Y2=1.542
r122 15 17 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.275 $Y=1.765
+ $X2=7.275 $Y2=2.4
r123 11 45 24.162 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=6.935 $Y=1.32
+ $X2=6.935 $Y2=1.542
r124 11 13 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.935 $Y=1.32
+ $X2=6.935 $Y2=0.74
r125 8 44 24.162 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=6.725 $Y=1.765
+ $X2=6.725 $Y2=1.542
r126 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.725 $Y=1.765
+ $X2=6.725 $Y2=2.4
r127 4 43 24.162 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=6.505 $Y=1.32
+ $X2=6.505 $Y2=1.542
r128 4 6 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.505 $Y=1.32
+ $X2=6.505 $Y2=0.74
r129 1 41 24.162 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=6.275 $Y=1.765
+ $X2=6.275 $Y2=1.542
r130 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.275 $Y=1.765
+ $X2=6.275 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__NAND4BB_4%D 3 5 7 10 12 14 17 19 21 22 24 27 29 30
+ 31 32 46
c86 32 0 6.20142e-20 $X=9.84 $Y=1.665
r87 48 49 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=9.765
+ $Y=1.465 $X2=9.765 $Y2=1.465
r88 46 48 22.712 $w=3.82e-07 $l=1.8e-07 $layer=POLY_cond $X=9.585 $Y=1.532
+ $X2=9.765 $Y2=1.532
r89 45 46 1.26178 $w=3.82e-07 $l=1e-08 $layer=POLY_cond $X=9.575 $Y=1.532
+ $X2=9.585 $Y2=1.532
r90 44 45 56.7801 $w=3.82e-07 $l=4.5e-07 $layer=POLY_cond $X=9.125 $Y=1.532
+ $X2=9.575 $Y2=1.532
r91 43 44 5.04712 $w=3.82e-07 $l=4e-08 $layer=POLY_cond $X=9.085 $Y=1.532
+ $X2=9.125 $Y2=1.532
r92 42 43 51.733 $w=3.82e-07 $l=4.1e-07 $layer=POLY_cond $X=8.675 $Y=1.532
+ $X2=9.085 $Y2=1.532
r93 41 42 2.52356 $w=3.82e-07 $l=2e-08 $layer=POLY_cond $X=8.655 $Y=1.532
+ $X2=8.675 $Y2=1.532
r94 39 41 31.5445 $w=3.82e-07 $l=2.5e-07 $layer=POLY_cond $X=8.405 $Y=1.532
+ $X2=8.655 $Y2=1.532
r95 39 40 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=8.405
+ $Y=1.465 $X2=8.405 $Y2=1.465
r96 37 39 22.712 $w=3.82e-07 $l=1.8e-07 $layer=POLY_cond $X=8.225 $Y=1.532
+ $X2=8.405 $Y2=1.532
r97 32 49 1.86887 $w=4.78e-07 $l=7.5e-08 $layer=LI1_cond $X=9.84 $Y=1.54
+ $X2=9.765 $Y2=1.54
r98 31 49 10.0919 $w=4.78e-07 $l=4.05e-07 $layer=LI1_cond $X=9.36 $Y=1.54
+ $X2=9.765 $Y2=1.54
r99 30 31 11.9608 $w=4.78e-07 $l=4.8e-07 $layer=LI1_cond $X=8.88 $Y=1.54
+ $X2=9.36 $Y2=1.54
r100 30 40 11.8362 $w=4.78e-07 $l=4.75e-07 $layer=LI1_cond $X=8.88 $Y=1.54
+ $X2=8.405 $Y2=1.54
r101 29 40 0.124591 $w=4.78e-07 $l=5e-09 $layer=LI1_cond $X=8.4 $Y=1.54
+ $X2=8.405 $Y2=1.54
r102 25 46 24.74 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=9.585 $Y=1.3
+ $X2=9.585 $Y2=1.532
r103 25 27 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=9.585 $Y=1.3
+ $X2=9.585 $Y2=0.74
r104 22 45 24.74 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=9.575 $Y=1.765
+ $X2=9.575 $Y2=1.532
r105 22 24 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=9.575 $Y=1.765
+ $X2=9.575 $Y2=2.4
r106 19 44 24.74 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=9.125 $Y=1.765
+ $X2=9.125 $Y2=1.532
r107 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=9.125 $Y=1.765
+ $X2=9.125 $Y2=2.4
r108 15 43 24.74 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=9.085 $Y=1.3
+ $X2=9.085 $Y2=1.532
r109 15 17 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=9.085 $Y=1.3
+ $X2=9.085 $Y2=0.74
r110 12 42 24.74 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=8.675 $Y=1.765
+ $X2=8.675 $Y2=1.532
r111 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.675 $Y=1.765
+ $X2=8.675 $Y2=2.4
r112 8 41 24.74 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=8.655 $Y=1.3
+ $X2=8.655 $Y2=1.532
r113 8 10 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=8.655 $Y=1.3
+ $X2=8.655 $Y2=0.74
r114 5 37 24.74 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=8.225 $Y=1.765
+ $X2=8.225 $Y2=1.532
r115 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.225 $Y=1.765
+ $X2=8.225 $Y2=2.4
r116 1 37 24.74 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=8.225 $Y=1.3
+ $X2=8.225 $Y2=1.532
r117 1 3 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=8.225 $Y=1.3
+ $X2=8.225 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__NAND4BB_4%VPWR 1 2 3 4 5 6 7 8 9 10 11 34 36 40 44
+ 48 50 54 56 60 64 68 70 74 76 80 82 84 88 89 90 92 97 106 111 116 125 128 131
+ 134 137 140 143 146 150
r174 149 150 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r175 146 147 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r176 144 147 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.88 $Y2=3.33
r177 143 144 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r178 141 144 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.92 $Y2=3.33
r179 140 141 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r180 137 138 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r181 131 132 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r182 128 129 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r183 125 126 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r184 122 123 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r185 120 150 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=9.84 $Y2=3.33
r186 120 147 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=8.88 $Y2=3.33
r187 119 120 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r188 117 146 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.985 $Y=3.33
+ $X2=8.9 $Y2=3.33
r189 117 119 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=8.985 $Y=3.33
+ $X2=9.36 $Y2=3.33
r190 116 149 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=9.715 $Y=3.33
+ $X2=9.897 $Y2=3.33
r191 116 119 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=9.715 $Y=3.33
+ $X2=9.36 $Y2=3.33
r192 115 141 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6.96 $Y2=3.33
r193 115 138 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6 $Y2=3.33
r194 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r195 112 137 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.135 $Y=3.33
+ $X2=6.01 $Y2=3.33
r196 112 114 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=6.135 $Y=3.33
+ $X2=6.48 $Y2=3.33
r197 111 140 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.835 $Y=3.33
+ $X2=7 $Y2=3.33
r198 111 114 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=6.835 $Y=3.33
+ $X2=6.48 $Y2=3.33
r199 110 138 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6 $Y2=3.33
r200 109 110 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r201 107 134 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.315 $Y=3.33
+ $X2=5.15 $Y2=3.33
r202 107 109 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=5.315 $Y=3.33
+ $X2=5.52 $Y2=3.33
r203 106 137 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.885 $Y=3.33
+ $X2=6.01 $Y2=3.33
r204 106 109 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=5.885 $Y=3.33
+ $X2=5.52 $Y2=3.33
r205 105 132 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r206 105 129 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.16 $Y2=3.33
r207 104 105 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r208 102 128 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.335 $Y=3.33
+ $X2=2.17 $Y2=3.33
r209 102 104 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=2.335 $Y=3.33
+ $X2=3.12 $Y2=3.33
r210 101 129 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r211 101 126 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r212 100 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r213 98 125 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.345 $Y=3.33
+ $X2=1.18 $Y2=3.33
r214 98 100 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.345 $Y=3.33
+ $X2=1.68 $Y2=3.33
r215 97 128 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.005 $Y=3.33
+ $X2=2.17 $Y2=3.33
r216 97 100 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.005 $Y=3.33
+ $X2=1.68 $Y2=3.33
r217 96 126 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r218 96 123 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r219 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r220 93 122 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.222 $Y2=3.33
r221 93 95 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.72 $Y2=3.33
r222 92 125 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.015 $Y=3.33
+ $X2=1.18 $Y2=3.33
r223 92 95 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.015 $Y=3.33
+ $X2=0.72 $Y2=3.33
r224 90 110 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r225 90 132 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.08 $Y2=3.33
r226 90 134 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r227 88 104 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=3.135 $Y=3.33
+ $X2=3.12 $Y2=3.33
r228 88 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.135 $Y=3.33
+ $X2=3.3 $Y2=3.33
r229 84 87 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=9.84 $Y=2.115
+ $X2=9.84 $Y2=2.815
r230 82 149 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=9.84 $Y=3.245
+ $X2=9.897 $Y2=3.33
r231 82 87 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=9.84 $Y=3.245
+ $X2=9.84 $Y2=2.815
r232 78 146 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.9 $Y=3.245
+ $X2=8.9 $Y2=3.33
r233 78 80 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=8.9 $Y=3.245
+ $X2=8.9 $Y2=2.455
r234 77 143 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.115 $Y=3.33
+ $X2=7.99 $Y2=3.33
r235 76 146 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.815 $Y=3.33
+ $X2=8.9 $Y2=3.33
r236 76 77 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=8.815 $Y=3.33
+ $X2=8.115 $Y2=3.33
r237 72 143 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.99 $Y=3.245
+ $X2=7.99 $Y2=3.33
r238 72 74 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=7.99 $Y=3.245
+ $X2=7.99 $Y2=2.455
r239 71 140 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.165 $Y=3.33
+ $X2=7 $Y2=3.33
r240 70 143 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.865 $Y=3.33
+ $X2=7.99 $Y2=3.33
r241 70 71 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=7.865 $Y=3.33
+ $X2=7.165 $Y2=3.33
r242 66 140 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7 $Y=3.245 $X2=7
+ $Y2=3.33
r243 66 68 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=7 $Y=3.245 $X2=7
+ $Y2=2.455
r244 62 137 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.01 $Y=3.245
+ $X2=6.01 $Y2=3.33
r245 62 64 42.4099 $w=2.48e-07 $l=9.2e-07 $layer=LI1_cond $X=6.01 $Y=3.245
+ $X2=6.01 $Y2=2.325
r246 58 134 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.15 $Y=3.245
+ $X2=5.15 $Y2=3.33
r247 58 60 31.081 $w=3.28e-07 $l=8.9e-07 $layer=LI1_cond $X=5.15 $Y=3.245
+ $X2=5.15 $Y2=2.355
r248 57 131 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.365 $Y=3.33
+ $X2=4.2 $Y2=3.33
r249 56 134 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.985 $Y=3.33
+ $X2=5.15 $Y2=3.33
r250 56 57 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=4.985 $Y=3.33
+ $X2=4.365 $Y2=3.33
r251 52 131 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.2 $Y=3.245
+ $X2=4.2 $Y2=3.33
r252 52 54 26.1919 $w=3.28e-07 $l=7.5e-07 $layer=LI1_cond $X=4.2 $Y=3.245
+ $X2=4.2 $Y2=2.495
r253 51 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.465 $Y=3.33
+ $X2=3.3 $Y2=3.33
r254 50 131 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.035 $Y=3.33
+ $X2=4.2 $Y2=3.33
r255 50 51 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=4.035 $Y=3.33
+ $X2=3.465 $Y2=3.33
r256 46 89 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.3 $Y=3.245 $X2=3.3
+ $Y2=3.33
r257 46 48 26.1919 $w=3.28e-07 $l=7.5e-07 $layer=LI1_cond $X=3.3 $Y=3.245
+ $X2=3.3 $Y2=2.495
r258 42 128 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.17 $Y=3.245
+ $X2=2.17 $Y2=3.33
r259 42 44 26.1919 $w=3.28e-07 $l=7.5e-07 $layer=LI1_cond $X=2.17 $Y=3.245
+ $X2=2.17 $Y2=2.495
r260 38 125 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.18 $Y=3.245
+ $X2=1.18 $Y2=3.33
r261 38 40 26.1919 $w=3.28e-07 $l=7.5e-07 $layer=LI1_cond $X=1.18 $Y=3.245
+ $X2=1.18 $Y2=2.495
r262 34 122 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.222 $Y2=3.33
r263 34 36 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.28 $Y2=2.455
r264 11 87 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=9.65
+ $Y=1.84 $X2=9.8 $Y2=2.815
r265 11 84 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=9.65
+ $Y=1.84 $X2=9.8 $Y2=2.115
r266 10 80 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=8.75
+ $Y=1.84 $X2=8.9 $Y2=2.455
r267 9 74 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=7.8
+ $Y=1.84 $X2=7.95 $Y2=2.455
r268 8 68 300 $w=1.7e-07 $l=7.07972e-07 $layer=licon1_PDIFF $count=2 $X=6.8
+ $Y=1.84 $X2=7 $Y2=2.455
r269 7 64 300 $w=1.7e-07 $l=5.54955e-07 $layer=licon1_PDIFF $count=2 $X=5.9
+ $Y=1.84 $X2=6.05 $Y2=2.325
r270 6 60 300 $w=1.7e-07 $l=6.06815e-07 $layer=licon1_PDIFF $count=2 $X=4.95
+ $Y=1.84 $X2=5.15 $Y2=2.355
r271 5 54 300 $w=1.7e-07 $l=7.26137e-07 $layer=licon1_PDIFF $count=2 $X=4.05
+ $Y=1.84 $X2=4.2 $Y2=2.495
r272 4 48 300 $w=1.7e-07 $l=7.26137e-07 $layer=licon1_PDIFF $count=2 $X=3.15
+ $Y=1.84 $X2=3.3 $Y2=2.495
r273 3 44 300 $w=1.7e-07 $l=4.80234e-07 $layer=licon1_PDIFF $count=2 $X=1.93
+ $Y=2.12 $X2=2.17 $Y2=2.495
r274 2 40 300 $w=1.7e-07 $l=4.43706e-07 $layer=licon1_PDIFF $count=2 $X=1.03
+ $Y=2.12 $X2=1.18 $Y2=2.495
r275 1 36 300 $w=1.7e-07 $l=4.00999e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.12 $X2=0.28 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_LS__NAND4BB_4%Y 1 2 3 4 5 6 7 8 9 10 31 33 35 38 42 44
+ 48 50 53 56 58 62 64 68 70 74 76 78 80 83 87 90 94 95 102 103 109 111 114 115
c202 87 0 1.98429e-19 $X=2.745 $Y=2.23
c203 58 0 1.227e-20 $X=6.335 $Y=1.905
c204 44 0 6.63463e-21 $X=4.485 $Y=2.145
c205 38 0 2.42988e-20 $X=5.515 $Y=1.175
r206 115 121 7.59565 $w=4.38e-07 $l=2.9e-07 $layer=LI1_cond $X=2.745 $Y=2.775
+ $X2=2.745 $Y2=2.485
r207 114 121 2.09535 $w=4.38e-07 $l=8e-08 $layer=LI1_cond $X=2.745 $Y=2.405
+ $X2=2.745 $Y2=2.485
r208 106 107 1.74613 $w=3.28e-07 $l=5e-08 $layer=LI1_cond $X=6.5 $Y=1.985
+ $X2=6.5 $Y2=2.035
r209 103 106 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=6.5 $Y=1.905 $X2=6.5
+ $Y2=1.985
r210 99 100 3.26614 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=4.65 $Y=2.145
+ $X2=4.65 $Y2=2.23
r211 98 99 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=4.65 $Y=2.015
+ $X2=4.65 $Y2=2.145
r212 95 98 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=4.65 $Y=1.935 $X2=4.65
+ $Y2=2.015
r213 90 91 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=3.42 $Y=0.955
+ $X2=3.42 $Y2=1.175
r214 87 114 4.58358 $w=4.38e-07 $l=1.75e-07 $layer=LI1_cond $X=2.745 $Y=2.23
+ $X2=2.745 $Y2=2.405
r215 87 89 2.42973 $w=4.4e-07 $l=8.5e-08 $layer=LI1_cond $X=2.745 $Y=2.23
+ $X2=2.745 $Y2=2.145
r216 83 85 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=2.485 $Y=0.815
+ $X2=2.485 $Y2=0.955
r217 78 113 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.35 $Y=2.12
+ $X2=9.35 $Y2=2.035
r218 78 80 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=9.35 $Y=2.12
+ $X2=9.35 $Y2=2.815
r219 77 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.615 $Y=2.035
+ $X2=8.45 $Y2=2.035
r220 76 113 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.185 $Y=2.035
+ $X2=9.35 $Y2=2.035
r221 76 77 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=9.185 $Y=2.035
+ $X2=8.615 $Y2=2.035
r222 72 111 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.45 $Y=2.12
+ $X2=8.45 $Y2=2.035
r223 72 74 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=8.45 $Y=2.12
+ $X2=8.45 $Y2=2.815
r224 71 109 8.61065 $w=1.7e-07 $l=1.94808e-07 $layer=LI1_cond $X=7.665 $Y=2.035
+ $X2=7.5 $Y2=1.97
r225 70 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.285 $Y=2.035
+ $X2=8.45 $Y2=2.035
r226 70 71 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=8.285 $Y=2.035
+ $X2=7.665 $Y2=2.035
r227 66 109 0.89609 $w=3.3e-07 $l=1.5e-07 $layer=LI1_cond $X=7.5 $Y=2.12 $X2=7.5
+ $Y2=1.97
r228 66 68 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=7.5 $Y=2.12
+ $X2=7.5 $Y2=2.815
r229 65 107 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.665 $Y=2.035
+ $X2=6.5 $Y2=2.035
r230 64 109 8.61065 $w=1.7e-07 $l=1.94808e-07 $layer=LI1_cond $X=7.335 $Y=2.035
+ $X2=7.5 $Y2=1.97
r231 64 65 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.335 $Y=2.035
+ $X2=6.665 $Y2=2.035
r232 60 107 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=6.5 $Y=2.12
+ $X2=6.5 $Y2=2.035
r233 60 62 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=6.5 $Y=2.12
+ $X2=6.5 $Y2=2.815
r234 59 102 3.05 $w=1.7e-07 $l=9.21954e-08 $layer=LI1_cond $X=5.685 $Y=1.905
+ $X2=5.6 $Y2=1.92
r235 58 103 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.335 $Y=1.905
+ $X2=6.5 $Y2=1.905
r236 58 59 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=6.335 $Y=1.905
+ $X2=5.685 $Y2=1.905
r237 54 102 3.05 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=5.6 $Y=2.02 $X2=5.6
+ $Y2=1.92
r238 54 56 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=5.6 $Y=2.02
+ $X2=5.6 $Y2=2.815
r239 53 102 3.05 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=5.6 $Y=1.82 $X2=5.6
+ $Y2=1.92
r240 52 53 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=5.6 $Y=1.26 $X2=5.6
+ $Y2=1.82
r241 51 95 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.815 $Y=1.935
+ $X2=4.65 $Y2=1.935
r242 50 102 3.05 $w=1.7e-07 $l=9.21954e-08 $layer=LI1_cond $X=5.515 $Y=1.935
+ $X2=5.6 $Y2=1.92
r243 50 51 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=5.515 $Y=1.935
+ $X2=4.815 $Y2=1.935
r244 48 100 7.61436 $w=2.78e-07 $l=1.85e-07 $layer=LI1_cond $X=4.675 $Y=2.415
+ $X2=4.675 $Y2=2.23
r245 45 94 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=3.865 $Y=2.145
+ $X2=3.75 $Y2=2.145
r246 44 99 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.485 $Y=2.145
+ $X2=4.65 $Y2=2.145
r247 44 45 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=4.485 $Y=2.145
+ $X2=3.865 $Y2=2.145
r248 40 94 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.75 $Y=2.23
+ $X2=3.75 $Y2=2.145
r249 40 42 12.7771 $w=2.28e-07 $l=2.55e-07 $layer=LI1_cond $X=3.75 $Y=2.23
+ $X2=3.75 $Y2=2.485
r250 39 91 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.505 $Y=1.175
+ $X2=3.42 $Y2=1.175
r251 38 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.515 $Y=1.175
+ $X2=5.6 $Y2=1.26
r252 38 39 131.134 $w=1.68e-07 $l=2.01e-06 $layer=LI1_cond $X=5.515 $Y=1.175
+ $X2=3.505 $Y2=1.175
r253 35 90 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.42 $Y=0.87
+ $X2=3.42 $Y2=0.955
r254 35 37 0.717647 $w=1.7e-07 $l=1e-08 $layer=LI1_cond $X=3.42 $Y=0.87 $X2=3.42
+ $Y2=0.86
r255 34 89 6.28872 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=2.965 $Y=2.145
+ $X2=2.745 $Y2=2.145
r256 33 94 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=3.635 $Y=2.145
+ $X2=3.75 $Y2=2.145
r257 33 34 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.635 $Y=2.145
+ $X2=2.965 $Y2=2.145
r258 32 85 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.65 $Y=0.955
+ $X2=2.485 $Y2=0.955
r259 31 90 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.335 $Y=0.955
+ $X2=3.42 $Y2=0.955
r260 31 32 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=3.335 $Y=0.955
+ $X2=2.65 $Y2=0.955
r261 10 113 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=9.2
+ $Y=1.84 $X2=9.35 $Y2=2.115
r262 10 80 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=9.2
+ $Y=1.84 $X2=9.35 $Y2=2.815
r263 9 111 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=8.3
+ $Y=1.84 $X2=8.45 $Y2=2.115
r264 9 74 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=8.3
+ $Y=1.84 $X2=8.45 $Y2=2.815
r265 8 109 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=7.35
+ $Y=1.84 $X2=7.5 $Y2=1.985
r266 8 68 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=7.35
+ $Y=1.84 $X2=7.5 $Y2=2.815
r267 7 106 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=6.35
+ $Y=1.84 $X2=6.5 $Y2=1.985
r268 7 62 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=6.35
+ $Y=1.84 $X2=6.5 $Y2=2.815
r269 6 102 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=5.45
+ $Y=1.84 $X2=5.6 $Y2=1.985
r270 6 56 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=5.45
+ $Y=1.84 $X2=5.6 $Y2=2.815
r271 5 98 600 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=1 $X=4.5
+ $Y=1.84 $X2=4.65 $Y2=2.015
r272 5 48 300 $w=1.7e-07 $l=6.45659e-07 $layer=licon1_PDIFF $count=2 $X=4.5
+ $Y=1.84 $X2=4.65 $Y2=2.415
r273 4 94 600 $w=1.7e-07 $l=3.72525e-07 $layer=licon1_PDIFF $count=1 $X=3.6
+ $Y=1.84 $X2=3.75 $Y2=2.145
r274 4 42 300 $w=1.7e-07 $l=7.16083e-07 $layer=licon1_PDIFF $count=2 $X=3.6
+ $Y=1.84 $X2=3.75 $Y2=2.485
r275 3 121 300 $w=1.7e-07 $l=7.16083e-07 $layer=licon1_PDIFF $count=2 $X=2.65
+ $Y=1.84 $X2=2.8 $Y2=2.485
r276 3 89 600 $w=1.7e-07 $l=3.72525e-07 $layer=licon1_PDIFF $count=1 $X=2.65
+ $Y=1.84 $X2=2.8 $Y2=2.145
r277 2 37 182 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_NDIFF $count=1 $X=3.28
+ $Y=0.37 $X2=3.42 $Y2=0.86
r278 1 83 182 $w=1.7e-07 $l=5.27376e-07 $layer=licon1_NDIFF $count=1 $X=2.305
+ $Y=0.37 $X2=2.485 $Y2=0.815
.ends

.subckt PM_SKY130_FD_SC_LS__NAND4BB_4%VGND 1 2 3 12 16 20 22 24 29 37 44 45 48
+ 51 54
r94 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r95 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r96 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r97 45 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0 $X2=9.36
+ $Y2=0
r98 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r99 42 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.465 $Y=0 $X2=9.3
+ $Y2=0
r100 42 44 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=9.465 $Y=0
+ $X2=9.84 $Y2=0
r101 41 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=9.36
+ $Y2=0
r102 41 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=8.4
+ $Y2=0
r103 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r104 38 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.605 $Y=0 $X2=8.44
+ $Y2=0
r105 38 40 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=8.605 $Y=0
+ $X2=8.88 $Y2=0
r106 37 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.135 $Y=0 $X2=9.3
+ $Y2=0
r107 37 40 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=9.135 $Y=0
+ $X2=8.88 $Y2=0
r108 36 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.4
+ $Y2=0
r109 35 36 1.24 $w=1.7e-07 $l=1.275e-06 $layer=mcon $count=7 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r110 33 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r111 32 35 438.417 $w=1.68e-07 $l=6.72e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=7.92
+ $Y2=0
r112 32 33 1.24 $w=1.7e-07 $l=1.275e-06 $layer=mcon $count=7 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r113 30 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=0.79
+ $Y2=0
r114 30 32 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=1.2
+ $Y2=0
r115 29 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.275 $Y=0 $X2=8.44
+ $Y2=0
r116 29 35 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=8.275 $Y=0
+ $X2=7.92 $Y2=0
r117 27 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r118 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r119 24 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.625 $Y=0 $X2=0.79
+ $Y2=0
r120 24 26 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.625 $Y=0
+ $X2=0.24 $Y2=0
r121 22 36 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=7.92 $Y2=0
r122 22 33 1.07034 $w=4.9e-07 $l=3.84e-06 $layer=MET1_cond $X=5.04 $Y=0 $X2=1.2
+ $Y2=0
r123 18 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.3 $Y=0.085 $X2=9.3
+ $Y2=0
r124 18 20 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=9.3 $Y=0.085
+ $X2=9.3 $Y2=0.57
r125 14 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.44 $Y=0.085
+ $X2=8.44 $Y2=0
r126 14 16 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=8.44 $Y=0.085
+ $X2=8.44 $Y2=0.57
r127 10 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.79 $Y=0.085
+ $X2=0.79 $Y2=0
r128 10 12 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=0.79 $Y=0.085
+ $X2=0.79 $Y2=0.325
r129 3 20 182 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=1 $X=9.16
+ $Y=0.37 $X2=9.3 $Y2=0.57
r130 2 16 182 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=1 $X=8.3
+ $Y=0.37 $X2=8.44 $Y2=0.57
r131 1 12 182 $w=1.7e-07 $l=3.37528e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.57 $X2=0.79 $Y2=0.325
.ends

.subckt PM_SKY130_FD_SC_LS__NAND4BB_4%A_374_74# 1 2 3 4 5 18 20 21 22 27 28 29
+ 32 38
c63 22 0 7.06753e-20 $X=3.685 $Y=0.34
c64 20 0 7.06753e-20 $X=2.82 $Y=0.34
r65 38 40 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=5.73 $Y=0.715
+ $X2=5.73 $Y2=0.835
r66 32 35 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=2.985 $Y=0.34
+ $X2=2.985 $Y2=0.525
r67 29 31 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=3.935 $Y=0.835
+ $X2=4.71 $Y2=0.835
r68 28 40 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.565 $Y=0.835
+ $X2=5.73 $Y2=0.835
r69 28 31 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=5.565 $Y=0.835
+ $X2=4.71 $Y2=0.835
r70 25 29 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.81 $Y=0.75
+ $X2=3.935 $Y2=0.835
r71 25 27 5.30124 $w=2.48e-07 $l=1.15e-07 $layer=LI1_cond $X=3.81 $Y=0.75
+ $X2=3.81 $Y2=0.635
r72 24 27 9.68052 $w=2.48e-07 $l=2.1e-07 $layer=LI1_cond $X=3.81 $Y=0.425
+ $X2=3.81 $Y2=0.635
r73 23 32 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.15 $Y=0.34
+ $X2=2.985 $Y2=0.34
r74 22 24 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.685 $Y=0.34
+ $X2=3.81 $Y2=0.425
r75 22 23 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=3.685 $Y=0.34
+ $X2=3.15 $Y2=0.34
r76 20 32 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.82 $Y=0.34
+ $X2=2.985 $Y2=0.34
r77 20 21 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=2.82 $Y=0.34 $X2=2.1
+ $Y2=0.34
r78 16 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.015 $Y=0.425
+ $X2=2.1 $Y2=0.34
r79 16 18 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=2.015 $Y=0.425
+ $X2=2.015 $Y2=0.515
r80 5 38 182 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_NDIFF $count=1 $X=5.59
+ $Y=0.37 $X2=5.73 $Y2=0.715
r81 4 31 182 $w=1.7e-07 $l=5.30401e-07 $layer=licon1_NDIFF $count=1 $X=4.57
+ $Y=0.37 $X2=4.71 $Y2=0.835
r82 3 27 182 $w=1.7e-07 $l=3.27605e-07 $layer=licon1_NDIFF $count=1 $X=3.71
+ $Y=0.37 $X2=3.85 $Y2=0.635
r83 2 35 182 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=1 $X=2.84
+ $Y=0.37 $X2=2.985 $Y2=0.525
r84 1 18 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=1.87
+ $Y=0.37 $X2=2.015 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__NAND4BB_4%A_828_74# 1 2 3 4 13 19 23 25 29 31 32
c51 19 0 2.42988e-20 $X=6.555 $Y=0.34
c52 13 0 1.79504e-19 $X=5.223 $Y=0.417
r53 27 29 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=7.58 $Y=0.425
+ $X2=7.58 $Y2=0.58
r54 26 32 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.885 $Y=0.34
+ $X2=6.72 $Y2=0.34
r55 25 27 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.415 $Y=0.34
+ $X2=7.58 $Y2=0.425
r56 25 26 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=7.415 $Y=0.34
+ $X2=6.885 $Y2=0.34
r57 21 32 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.72 $Y=0.425
+ $X2=6.72 $Y2=0.34
r58 21 23 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=6.72 $Y=0.425
+ $X2=6.72 $Y2=0.58
r59 19 32 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.555 $Y=0.34
+ $X2=6.72 $Y2=0.34
r60 19 31 76.3316 $w=1.68e-07 $l=1.17e-06 $layer=LI1_cond $X=6.555 $Y=0.34
+ $X2=5.385 $Y2=0.34
r61 15 18 33.3322 $w=3.23e-07 $l=9.4e-07 $layer=LI1_cond $X=4.28 $Y=0.417
+ $X2=5.22 $Y2=0.417
r62 13 31 8.35379 $w=3.23e-07 $l=1.62e-07 $layer=LI1_cond $X=5.223 $Y=0.417
+ $X2=5.385 $Y2=0.417
r63 13 18 0.106379 $w=3.23e-07 $l=3e-09 $layer=LI1_cond $X=5.223 $Y=0.417
+ $X2=5.22 $Y2=0.417
r64 4 29 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=7.44
+ $Y=0.37 $X2=7.58 $Y2=0.58
r65 3 23 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=6.58
+ $Y=0.37 $X2=6.72 $Y2=0.58
r66 2 18 182 $w=1.7e-07 $l=2.755e-07 $layer=licon1_NDIFF $count=1 $X=5 $Y=0.37
+ $X2=5.22 $Y2=0.495
r67 1 15 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=4.14
+ $Y=0.37 $X2=4.28 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LS__NAND4BB_4%A_1229_74# 1 2 3 4 5 18 20 21 24 26 30 32
+ 36 38 42 44 45 46
r73 40 42 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=9.8 $Y=0.96 $X2=9.8
+ $Y2=0.515
r74 39 46 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.955 $Y=1.045
+ $X2=8.87 $Y2=1.045
r75 38 40 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.635 $Y=1.045
+ $X2=9.8 $Y2=0.96
r76 38 39 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=9.635 $Y=1.045
+ $X2=8.955 $Y2=1.045
r77 34 46 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.87 $Y=0.96 $X2=8.87
+ $Y2=1.045
r78 34 36 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=8.87 $Y=0.96
+ $X2=8.87 $Y2=0.515
r79 33 45 5.16603 $w=1.7e-07 $l=8.9861e-08 $layer=LI1_cond $X=8.095 $Y=1.045
+ $X2=8.01 $Y2=1.055
r80 32 46 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.785 $Y=1.045
+ $X2=8.87 $Y2=1.045
r81 32 33 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=8.785 $Y=1.045
+ $X2=8.095 $Y2=1.045
r82 28 45 1.34256 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=8.01 $Y=0.96 $X2=8.01
+ $Y2=1.055
r83 28 30 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=8.01 $Y=0.96
+ $X2=8.01 $Y2=0.515
r84 27 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.235 $Y=1.065
+ $X2=7.15 $Y2=1.065
r85 26 45 5.16603 $w=1.7e-07 $l=8.9861e-08 $layer=LI1_cond $X=7.925 $Y=1.065
+ $X2=8.01 $Y2=1.055
r86 26 27 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=7.925 $Y=1.065
+ $X2=7.235 $Y2=1.065
r87 22 44 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.15 $Y=0.98 $X2=7.15
+ $Y2=1.065
r88 22 24 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=7.15 $Y=0.98
+ $X2=7.15 $Y2=0.86
r89 20 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.065 $Y=1.065
+ $X2=7.15 $Y2=1.065
r90 20 21 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=7.065 $Y=1.065
+ $X2=6.375 $Y2=1.065
r91 16 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.25 $Y=0.98
+ $X2=6.375 $Y2=1.065
r92 16 18 5.53173 $w=2.48e-07 $l=1.2e-07 $layer=LI1_cond $X=6.25 $Y=0.98
+ $X2=6.25 $Y2=0.86
r93 5 42 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.66
+ $Y=0.37 $X2=9.8 $Y2=0.515
r94 4 36 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.73
+ $Y=0.37 $X2=8.87 $Y2=0.515
r95 3 30 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.87
+ $Y=0.37 $X2=8.01 $Y2=0.515
r96 2 24 182 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_NDIFF $count=1 $X=7.01
+ $Y=0.37 $X2=7.15 $Y2=0.86
r97 1 18 182 $w=1.7e-07 $l=5.57808e-07 $layer=licon1_NDIFF $count=1 $X=6.145
+ $Y=0.37 $X2=6.29 $Y2=0.86
.ends

