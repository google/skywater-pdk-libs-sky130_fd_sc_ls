* File: sky130_fd_sc_ls__decaphe_18.pxi.spice
* Created: Fri Aug 28 13:11:52 2020
* 
x_PM_SKY130_FD_SC_LS__DECAPHE_18%VPWR N_VPWR_M1001_s N_VPWR_c_15_n
+ N_VPWR_M1000_g N_VPWR_c_16_n VPWR N_VPWR_c_17_n N_VPWR_c_18_n N_VPWR_c_19_n
+ N_VPWR_c_20_n N_VPWR_c_21_n N_VPWR_c_22_n VPWR
+ PM_SKY130_FD_SC_LS__DECAPHE_18%VPWR
x_PM_SKY130_FD_SC_LS__DECAPHE_18%VGND N_VGND_M1000_s VGND N_VGND_M1001_g
+ N_VGND_c_39_n N_VGND_c_40_n N_VGND_c_41_n VGND
+ PM_SKY130_FD_SC_LS__DECAPHE_18%VGND
cc_1 VNB N_VPWR_c_15_n 0.158308f $X=-0.19 $Y=-0.245 $X2=2.005 $Y2=0.622
cc_2 VNB N_VPWR_c_16_n 0.235581f $X=-0.19 $Y=-0.245 $X2=6.615 $Y2=0.622
cc_3 VNB N_VPWR_c_17_n 0.0757653f $X=-0.19 $Y=-0.245 $X2=3.095 $Y2=0.802
cc_4 VNB N_VPWR_c_18_n 0.084437f $X=-0.19 $Y=-0.245 $X2=3.765 $Y2=0.802
cc_5 VNB N_VPWR_c_19_n 0.0757653f $X=-0.19 $Y=-0.245 $X2=4.855 $Y2=0.802
cc_6 VNB N_VPWR_c_20_n 0.084437f $X=-0.19 $Y=-0.245 $X2=5.525 $Y2=0.802
cc_7 VNB N_VPWR_c_21_n 0.0268417f $X=-0.19 $Y=-0.245 $X2=8.38 $Y2=1.985
cc_8 VNB N_VPWR_c_22_n 0.362705f $X=-0.19 $Y=-0.245 $X2=8.4 $Y2=3.33
cc_9 VNB N_VGND_c_39_n 0.218881f $X=-0.19 $Y=-0.245 $X2=3.6 $Y2=1.335
cc_10 VNB N_VGND_c_40_n 0.286178f $X=-0.19 $Y=-0.245 $X2=3.6 $Y2=2.332
cc_11 VNB N_VGND_c_41_n 0.40592f $X=-0.19 $Y=-0.245 $X2=8.38 $Y2=2.332
cc_12 VPB N_VPWR_c_21_n 0.252637f $X=-0.19 $Y=1.66 $X2=8.38 $Y2=1.985
cc_13 VPB N_VPWR_c_22_n 0.0432146f $X=-0.19 $Y=1.66 $X2=8.4 $Y2=3.33
cc_14 VPB N_VGND_c_39_n 0.550081f $X=-0.19 $Y=1.66 $X2=3.6 $Y2=1.335
cc_15 N_VPWR_c_15_n N_VGND_c_39_n 0.113678f $X=2.005 $Y=0.622 $X2=0 $Y2=0
cc_16 N_VPWR_c_16_n N_VGND_c_39_n 0.160088f $X=6.615 $Y=0.622 $X2=0 $Y2=0
cc_17 N_VPWR_c_17_n N_VGND_c_39_n 0.045102f $X=3.095 $Y=0.802 $X2=0 $Y2=0
cc_18 N_VPWR_c_18_n N_VGND_c_39_n 0.0634323f $X=3.765 $Y=0.802 $X2=0 $Y2=0
cc_19 N_VPWR_c_19_n N_VGND_c_39_n 0.045102f $X=4.855 $Y=0.802 $X2=0 $Y2=0
cc_20 N_VPWR_c_20_n N_VGND_c_39_n 0.0634323f $X=5.525 $Y=0.802 $X2=0 $Y2=0
cc_21 N_VPWR_c_21_n N_VGND_c_39_n 1.43347f $X=8.38 $Y=1.985 $X2=0 $Y2=0
cc_22 N_VPWR_c_15_n N_VGND_c_40_n 0.224087f $X=2.005 $Y=0.622 $X2=0 $Y2=0
cc_23 N_VPWR_c_16_n N_VGND_c_40_n 0.371271f $X=6.615 $Y=0.622 $X2=0 $Y2=0
cc_24 N_VPWR_c_17_n N_VGND_c_40_n 0.144464f $X=3.095 $Y=0.802 $X2=0 $Y2=0
cc_25 N_VPWR_c_18_n N_VGND_c_40_n 0.0959058f $X=3.765 $Y=0.802 $X2=0 $Y2=0
cc_26 N_VPWR_c_19_n N_VGND_c_40_n 0.144464f $X=4.855 $Y=0.802 $X2=0 $Y2=0
cc_27 N_VPWR_c_20_n N_VGND_c_40_n 0.0959058f $X=5.525 $Y=0.802 $X2=0 $Y2=0
cc_28 N_VPWR_c_21_n N_VGND_c_40_n 0.841455f $X=8.38 $Y=1.985 $X2=0 $Y2=0
