* File: sky130_fd_sc_ls__a22o_1.pex.spice
* Created: Wed Sep  2 10:50:11 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__A22O_1%A2 1 2 3 5 9 11 17
r31 14 17 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=0.395 $Y=0.34
+ $X2=0.6 $Y2=0.34
r32 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.395
+ $Y=0.34 $X2=0.395 $Y2=0.34
r33 11 15 7.43059 $w=3.53e-07 $l=2.15e-07 $layer=LI1_cond $X=0.342 $Y=0.555
+ $X2=0.342 $Y2=0.34
r34 9 10 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.6 $Y=0.935 $X2=0.6
+ $Y2=1.33
r35 6 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.6 $Y=0.505 $X2=0.6
+ $Y2=0.34
r36 6 9 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=0.6 $Y=0.505 $X2=0.6
+ $Y2=0.935
r37 3 5 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.585 $Y=1.885
+ $X2=0.585 $Y2=2.46
r38 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.585 $Y=1.795 $X2=0.585
+ $Y2=1.885
r39 1 10 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.585 $Y=1.42 $X2=0.585
+ $Y2=1.33
r40 1 2 145.766 $w=1.8e-07 $l=3.75e-07 $layer=POLY_cond $X=0.585 $Y=1.42
+ $X2=0.585 $Y2=1.795
.ends

.subckt PM_SKY130_FD_SC_LS__A22O_1%B2 1 3 6 8 9 14
r35 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.05
+ $Y=1.635 $X2=1.05 $Y2=1.635
r36 9 14 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=0.72 $Y=1.635
+ $X2=1.05 $Y2=1.635
r37 8 9 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.24 $Y=1.635 $X2=0.72
+ $Y2=1.635
r38 4 13 38.5562 $w=2.99e-07 $l=1.77059e-07 $layer=POLY_cond $X=1.075 $Y=1.47
+ $X2=1.05 $Y2=1.635
r39 4 6 387.138 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=1.075 $Y=1.47
+ $X2=1.075 $Y2=0.715
r40 1 13 52.2586 $w=2.99e-07 $l=2.57391e-07 $layer=POLY_cond $X=1.035 $Y=1.885
+ $X2=1.05 $Y2=1.635
r41 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.035 $Y=1.885
+ $X2=1.035 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_LS__A22O_1%B1 3 5 6 8 9 10 11
c36 10 0 2.0037e-19 $X=1.467 $Y=1.26
c37 9 0 4.51155e-20 $X=1.467 $Y=1.11
r38 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.59
+ $Y=1.635 $X2=1.59 $Y2=1.635
r39 11 15 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=1.68 $Y=1.635 $X2=1.59
+ $Y2=1.635
r40 9 10 44.7709 $w=2.15e-07 $l=1.5e-07 $layer=POLY_cond $X=1.467 $Y=1.11
+ $X2=1.467 $Y2=1.26
r41 6 14 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=1.515 $Y=1.885
+ $X2=1.59 $Y2=1.635
r42 6 8 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.515 $Y=1.885
+ $X2=1.515 $Y2=2.46
r43 5 14 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=1.5 $Y=1.47
+ $X2=1.59 $Y2=1.635
r44 5 10 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=1.5 $Y=1.47 $X2=1.5
+ $Y2=1.26
r45 3 9 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.435 $Y=0.715
+ $X2=1.435 $Y2=1.11
.ends

.subckt PM_SKY130_FD_SC_LS__A22O_1%A1 1 3 4 6 7 11
r35 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.13
+ $Y=1.515 $X2=2.13 $Y2=1.515
r36 7 11 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=2.13 $Y=1.665
+ $X2=2.13 $Y2=1.515
r37 4 10 75.8144 $w=2.68e-07 $l=3.76444e-07 $layer=POLY_cond $X=2.055 $Y=1.885
+ $X2=2.042 $Y2=1.515
r38 4 6 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.055 $Y=1.885
+ $X2=2.055 $Y2=2.46
r39 1 10 82.1092 $w=2.68e-07 $l=4.855e-07 $layer=POLY_cond $X=1.865 $Y=1.11
+ $X2=2.042 $Y2=1.515
r40 1 3 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.865 $Y=1.11
+ $X2=1.865 $Y2=0.715
.ends

.subckt PM_SKY130_FD_SC_LS__A22O_1%A_222_392# 1 2 7 9 12 16 18 23 26 28
c57 18 0 8.56871e-20 $X=2.505 $Y=1.095
r58 28 30 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=1.65 $Y=0.885
+ $X2=1.65 $Y2=1.095
r59 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.67
+ $Y=1.465 $X2=2.67 $Y2=1.465
r60 21 23 23.2793 $w=2.48e-07 $l=5.05e-07 $layer=LI1_cond $X=2.63 $Y=1.97
+ $X2=2.63 $Y2=1.465
r61 20 23 13.1378 $w=2.48e-07 $l=2.85e-07 $layer=LI1_cond $X=2.63 $Y=1.18
+ $X2=2.63 $Y2=1.465
r62 19 30 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.815 $Y=1.095
+ $X2=1.65 $Y2=1.095
r63 18 20 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.505 $Y=1.095
+ $X2=2.63 $Y2=1.18
r64 18 19 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.505 $Y=1.095
+ $X2=1.815 $Y2=1.095
r65 17 26 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.425 $Y=2.055
+ $X2=1.26 $Y2=2.055
r66 16 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.505 $Y=2.055
+ $X2=2.63 $Y2=1.97
r67 16 17 70.4599 $w=1.68e-07 $l=1.08e-06 $layer=LI1_cond $X=2.505 $Y=2.055
+ $X2=1.425 $Y2=2.055
r68 10 24 38.6704 $w=3.39e-07 $l=2.27255e-07 $layer=POLY_cond $X=2.875 $Y=1.3
+ $X2=2.727 $Y2=1.465
r69 10 12 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.875 $Y=1.3
+ $X2=2.875 $Y2=0.74
r70 7 24 57.8651 $w=3.39e-07 $l=3.27719e-07 $layer=POLY_cond $X=2.785 $Y=1.765
+ $X2=2.727 $Y2=1.465
r71 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.785 $Y=1.765
+ $X2=2.785 $Y2=2.4
r72 2 26 300 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=2 $X=1.11
+ $Y=1.96 $X2=1.26 $Y2=2.135
r73 1 28 182 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_NDIFF $count=1 $X=1.51
+ $Y=0.395 $X2=1.65 $Y2=0.885
.ends

.subckt PM_SKY130_FD_SC_LS__A22O_1%VPWR 1 2 7 9 15 17 19 29 30 36
r35 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r36 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r37 30 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r38 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r39 27 36 12.0744 $w=1.7e-07 $l=2.8e-07 $layer=LI1_cond $X=2.725 $Y=3.33
+ $X2=2.445 $Y2=3.33
r40 27 29 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=2.725 $Y=3.33
+ $X2=3.12 $Y2=3.33
r41 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r42 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r43 23 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r44 22 25 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.72 $Y=3.33
+ $X2=2.16 $Y2=3.33
r45 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r46 20 33 3.92346 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.222 $Y2=3.33
r47 20 22 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.72 $Y2=3.33
r48 19 36 12.0744 $w=1.7e-07 $l=2.8e-07 $layer=LI1_cond $X=2.165 $Y=3.33
+ $X2=2.445 $Y2=3.33
r49 19 25 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=2.165 $Y=3.33
+ $X2=2.16 $Y2=3.33
r50 17 26 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r51 17 23 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r52 13 36 2.35715 $w=5.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.445 $Y=3.245
+ $X2=2.445 $Y2=3.33
r53 13 15 17.4072 $w=5.58e-07 $l=8.15e-07 $layer=LI1_cond $X=2.445 $Y=3.245
+ $X2=2.445 $Y2=2.43
r54 9 12 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=0.32 $Y=2.135
+ $X2=0.32 $Y2=2.815
r55 7 33 3.2197 $w=2.5e-07 $l=1.33918e-07 $layer=LI1_cond $X=0.32 $Y=3.245
+ $X2=0.222 $Y2=3.33
r56 7 12 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.32 $Y=3.245 $X2=0.32
+ $Y2=2.815
r57 2 15 300 $w=1.7e-07 $l=6.50385e-07 $layer=licon1_PDIFF $count=2 $X=2.13
+ $Y=1.96 $X2=2.56 $Y2=2.43
r58 1 12 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.235
+ $Y=1.96 $X2=0.36 $Y2=2.815
r59 1 9 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.235
+ $Y=1.96 $X2=0.36 $Y2=2.135
.ends

.subckt PM_SKY130_FD_SC_LS__A22O_1%A_132_392# 1 2 9 13 14 17
r22 15 17 12.3888 $w=3.98e-07 $l=4.3e-07 $layer=LI1_cond $X=1.795 $Y=2.905
+ $X2=1.795 $Y2=2.475
r23 13 15 8.37092 $w=1.7e-07 $l=2.38747e-07 $layer=LI1_cond $X=1.595 $Y=2.99
+ $X2=1.795 $Y2=2.905
r24 13 14 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.595 $Y=2.99
+ $X2=0.895 $Y2=2.99
r25 9 12 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=0.77 $Y=2.135
+ $X2=0.77 $Y2=2.815
r26 7 14 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.77 $Y=2.905
+ $X2=0.895 $Y2=2.99
r27 7 12 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=0.77 $Y=2.905 $X2=0.77
+ $Y2=2.815
r28 2 17 300 $w=1.7e-07 $l=6.08933e-07 $layer=licon1_PDIFF $count=2 $X=1.59
+ $Y=1.96 $X2=1.795 $Y2=2.475
r29 1 12 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=0.66
+ $Y=1.96 $X2=0.81 $Y2=2.815
r30 1 9 400 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=1 $X=0.66
+ $Y=1.96 $X2=0.81 $Y2=2.135
.ends

.subckt PM_SKY130_FD_SC_LS__A22O_1%X 1 2 7 8 9 10 11 12 13
r13 13 40 1.3969 $w=3.28e-07 $l=4e-08 $layer=LI1_cond $X=3.09 $Y=2.775 $X2=3.09
+ $Y2=2.815
r14 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.09 $Y=2.405
+ $X2=3.09 $Y2=2.775
r15 11 12 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.09 $Y=2.035
+ $X2=3.09 $Y2=2.405
r16 11 32 1.74613 $w=3.28e-07 $l=5e-08 $layer=LI1_cond $X=3.09 $Y=2.035 $X2=3.09
+ $Y2=1.985
r17 10 32 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=3.09 $Y=1.665
+ $X2=3.09 $Y2=1.985
r18 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.09 $Y=1.295
+ $X2=3.09 $Y2=1.665
r19 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.09 $Y=0.925 $X2=3.09
+ $Y2=1.295
r20 7 8 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=3.09 $Y=0.515 $X2=3.09
+ $Y2=0.925
r21 2 40 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.86
+ $Y=1.84 $X2=3.01 $Y2=2.815
r22 2 32 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.86
+ $Y=1.84 $X2=3.01 $Y2=1.985
r23 1 7 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.95
+ $Y=0.37 $X2=3.09 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__A22O_1%A_52_123# 1 2 7 10 11 13 16
c43 13 0 1.59798e-19 $X=2.08 $Y=0.54
r44 16 18 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=0.385 $Y=1.055
+ $X2=0.385 $Y2=1.215
r45 11 13 36.6477 $w=2.48e-07 $l=7.95e-07 $layer=LI1_cond $X=1.285 $Y=0.5
+ $X2=2.08 $Y2=0.5
r46 9 11 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.2 $Y=0.625
+ $X2=1.285 $Y2=0.5
r47 9 10 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=1.2 $Y=0.625 $X2=1.2
+ $Y2=1.13
r48 8 18 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.55 $Y=1.215
+ $X2=0.385 $Y2=1.215
r49 7 10 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.115 $Y=1.215
+ $X2=1.2 $Y2=1.13
r50 7 8 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=1.115 $Y=1.215
+ $X2=0.55 $Y2=1.215
r51 2 13 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1.94
+ $Y=0.395 $X2=2.08 $Y2=0.54
r52 1 16 182 $w=1.7e-07 $l=4.98598e-07 $layer=licon1_NDIFF $count=1 $X=0.26
+ $Y=0.615 $X2=0.385 $Y2=1.055
.ends

.subckt PM_SKY130_FD_SC_LS__A22O_1%VGND 1 2 9 13 16 17 18 24 33 34 37
r39 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r40 34 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r41 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r42 31 37 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.745 $Y=0 $X2=2.62
+ $Y2=0
r43 31 33 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=2.745 $Y=0 $X2=3.12
+ $Y2=0
r44 30 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r45 29 30 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r46 26 29 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r47 26 27 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r48 24 37 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.495 $Y=0 $X2=2.62
+ $Y2=0
r49 24 29 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.495 $Y=0 $X2=2.16
+ $Y2=0
r50 22 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r51 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r52 18 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r53 18 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r54 16 21 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=0.73 $Y=0 $X2=0.72
+ $Y2=0
r55 16 17 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=0.73 $Y=0 $X2=0.837
+ $Y2=0
r56 15 26 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=1.2
+ $Y2=0
r57 15 17 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=0.837
+ $Y2=0
r58 11 37 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.62 $Y=0.085
+ $X2=2.62 $Y2=0
r59 11 13 27.1977 $w=2.48e-07 $l=5.9e-07 $layer=LI1_cond $X=2.62 $Y=0.085
+ $X2=2.62 $Y2=0.675
r60 7 17 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=0.837 $Y=0.085
+ $X2=0.837 $Y2=0
r61 7 9 36.9854 $w=2.13e-07 $l=6.9e-07 $layer=LI1_cond $X=0.837 $Y=0.085
+ $X2=0.837 $Y2=0.775
r62 2 13 182 $w=1.7e-07 $l=3.62146e-07 $layer=licon1_NDIFF $count=1 $X=2.535
+ $Y=0.37 $X2=2.66 $Y2=0.675
r63 1 9 182 $w=1.7e-07 $l=2.26274e-07 $layer=licon1_NDIFF $count=1 $X=0.675
+ $Y=0.615 $X2=0.835 $Y2=0.775
.ends

