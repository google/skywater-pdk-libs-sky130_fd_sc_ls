* File: sky130_fd_sc_ls__and2b_1.spice
* Created: Wed Sep  2 10:54:24 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__and2b_1.pex.spice"
.subckt sky130_fd_sc_ls__and2b_1  VNB VPB A_N B VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B	B
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1006 N_VGND_M1006_d N_A_N_M1006_g N_A_27_74#_M1006_s VNB NSHORT L=0.15 W=0.55
+ AD=0.19525 AS=0.15675 PD=1.81 PS=1.67 NRD=15.264 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75000.3 A=0.0825 P=1.4 MULT=1
MM1000 A_353_98# N_A_27_74#_M1000_g N_A_266_98#_M1000_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0768 AS=0.1824 PD=0.88 PS=1.85 NRD=12.18 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75001.4 A=0.096 P=1.58 MULT=1
MM1001 N_VGND_M1001_d N_B_M1001_g A_353_98# VNB NSHORT L=0.15 W=0.64 AD=0.20007
+ AS=0.0768 PD=1.27536 PS=0.88 NRD=0 NRS=12.18 M=1 R=4.26667 SA=75000.6 SB=75001
+ A=0.096 P=1.58 MULT=1
MM1002 N_X_M1002_d N_A_266_98#_M1002_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.23133 PD=2.05 PS=1.47464 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1003 N_VPWR_M1003_d N_A_N_M1003_g N_A_27_74#_M1003_s VPB PHIGHVT L=0.15 W=0.84
+ AD=0.126 AS=0.8526 PD=1.14 PS=3.71 NRD=2.3443 NRS=2.3443 M=1 R=5.6 SA=75000.9
+ SB=75001.7 A=0.126 P=1.98 MULT=1
MM1005 N_A_266_98#_M1005_d N_A_27_74#_M1005_g N_VPWR_M1003_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.126 AS=0.126 PD=1.14 PS=1.14 NRD=2.3443 NRS=2.3443 M=1 R=5.6
+ SA=75001.4 SB=75001.3 A=0.126 P=1.98 MULT=1
MM1007 N_VPWR_M1007_d N_B_M1007_g N_A_266_98#_M1005_d VPB PHIGHVT L=0.15 W=0.84
+ AD=0.198 AS=0.126 PD=1.33286 PS=1.14 NRD=22.261 NRS=2.3443 M=1 R=5.6
+ SA=75001.8 SB=75000.8 A=0.126 P=1.98 MULT=1
MM1004 N_X_M1004_d N_A_266_98#_M1004_g N_VPWR_M1007_d VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.264 PD=2.83 PS=1.77714 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75001.9 SB=75000.2 A=0.168 P=2.54 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.9564 P=11.2
*
.include "sky130_fd_sc_ls__and2b_1.pxi.spice"
*
.ends
*
*
