* File: sky130_fd_sc_ls__clkbuf_2.spice
* Created: Wed Sep  2 10:57:37 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__clkbuf_2.pex.spice"
.subckt sky130_fd_sc_ls__clkbuf_2  VNB VPB A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1004 N_X_M1004_d N_A_43_192#_M1004_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75001.1
+ A=0.063 P=1.14 MULT=1
MM1005 N_X_M1004_d N_A_43_192#_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0735 PD=0.7 PS=0.77 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75000.7
+ A=0.063 P=1.14 MULT=1
MM1001 N_A_43_192#_M1001_d N_A_M1001_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0735 PD=1.41 PS=0.77 NRD=0 NRS=19.992 M=1 R=2.8 SA=75001.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1002 N_X_M1002_d N_A_43_192#_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.3192 PD=1.42 PS=2.81 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1003 N_X_M1002_d N_A_43_192#_M1003_g N_VPWR_M1003_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1000 N_A_43_192#_M1000_d N_A_M1000_g N_VPWR_M1003_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3528 AS=0.168 PD=2.87 PS=1.42 NRD=3.5066 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75000.2 A=0.168 P=2.54 MULT=1
DX6_noxref VNB VPB NWDIODE A=4.278 P=8.32
*
.include "sky130_fd_sc_ls__clkbuf_2.pxi.spice"
*
.ends
*
*
