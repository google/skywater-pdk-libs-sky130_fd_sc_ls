* File: sky130_fd_sc_ls__sedfxbp_2.pex.spice
* Created: Fri Aug 28 14:07:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__SEDFXBP_2%D 2 3 5 8 12 13 18 19 21 23
c43 23 0 2.19166e-19 $X=0.54 $Y=1.99
c44 18 0 8.95046e-20 $X=0.54 $Y=1.145
r45 21 23 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.54 $Y=1.825
+ $X2=0.54 $Y2=1.99
r46 21 22 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.54
+ $Y=1.825 $X2=0.54 $Y2=1.825
r47 18 21 118.906 $w=3.3e-07 $l=6.8e-07 $layer=POLY_cond $X=0.54 $Y=1.145
+ $X2=0.54 $Y2=1.825
r48 18 19 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.54
+ $Y=1.145 $X2=0.54 $Y2=1.145
r49 13 22 4.49734 $w=4.08e-07 $l=1.6e-07 $layer=LI1_cond $X=0.63 $Y=1.665
+ $X2=0.63 $Y2=1.825
r50 12 13 10.4001 $w=4.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.63 $Y=1.295
+ $X2=0.63 $Y2=1.665
r51 12 19 4.21625 $w=4.08e-07 $l=1.5e-07 $layer=LI1_cond $X=0.63 $Y=1.295
+ $X2=0.63 $Y2=1.145
r52 11 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.54 $Y=0.98
+ $X2=0.54 $Y2=1.145
r53 8 11 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=0.63 $Y=0.58 $X2=0.63
+ $Y2=0.98
r54 3 5 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.585 $Y=2.245
+ $X2=0.585 $Y2=2.64
r55 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.585 $Y=2.155 $X2=0.585
+ $Y2=2.245
r56 2 23 64.1371 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.585 $Y=2.155
+ $X2=0.585 $Y2=1.99
.ends

.subckt PM_SKY130_FD_SC_LS__SEDFXBP_2%A_183_290# 1 2 7 9 12 14 18 19 20 21 22 23
+ 26 30 32 36 37 39
c113 23 0 3.35759e-20 $X=1.335 $Y=2.035
c114 21 0 8.95046e-20 $X=1.335 $Y=1.195
r115 37 43 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.47 $Y=1.68
+ $X2=2.47 $Y2=1.515
r116 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.47
+ $Y=1.68 $X2=2.47 $Y2=1.68
r117 34 36 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=2.47 $Y=1.95
+ $X2=2.47 $Y2=1.68
r118 33 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.995 $Y=2.035
+ $X2=1.91 $Y2=2.035
r119 32 34 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.305 $Y=2.035
+ $X2=2.47 $Y2=1.95
r120 32 33 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=2.305 $Y=2.035
+ $X2=1.995 $Y2=2.035
r121 28 39 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.91 $Y=2.12
+ $X2=1.91 $Y2=2.035
r122 28 30 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=1.91 $Y=2.12
+ $X2=1.91 $Y2=2.51
r123 24 26 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.845 $Y=1.11
+ $X2=1.845 $Y2=0.775
r124 22 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.825 $Y=2.035
+ $X2=1.91 $Y2=2.035
r125 22 23 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=1.825 $Y=2.035
+ $X2=1.335 $Y2=2.035
r126 20 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.68 $Y=1.195
+ $X2=1.845 $Y2=1.11
r127 20 21 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.68 $Y=1.195
+ $X2=1.335 $Y2=1.195
r128 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.17
+ $Y=1.615 $X2=1.17 $Y2=1.615
r129 16 23 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.17 $Y=1.95
+ $X2=1.335 $Y2=2.035
r130 16 18 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.17 $Y=1.95
+ $X2=1.17 $Y2=1.615
r131 15 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.17 $Y=1.28
+ $X2=1.335 $Y2=1.195
r132 15 18 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.17 $Y=1.28
+ $X2=1.17 $Y2=1.615
r133 14 19 39.0632 $w=4.2e-07 $l=2.95e-07 $layer=POLY_cond $X=1.125 $Y=1.91
+ $X2=1.125 $Y2=1.615
r134 12 43 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=2.56 $Y=0.775
+ $X2=2.56 $Y2=1.515
r135 7 14 48.9303 $w=3.3e-07 $l=3.90416e-07 $layer=POLY_cond $X=1.005 $Y=2.245
+ $X2=1.125 $Y2=1.91
r136 7 9 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.005 $Y=2.245
+ $X2=1.005 $Y2=2.64
r137 2 30 600 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=1 $X=1.765
+ $Y=2.31 $X2=1.91 $Y2=2.51
r138 1 26 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=1.7
+ $Y=0.565 $X2=1.845 $Y2=0.775
.ends

.subckt PM_SKY130_FD_SC_LS__SEDFXBP_2%DE 3 5 6 9 12 13 14 15 17 18 20 21 23 25
+ 26 27 28 31 33
c95 21 0 1.25679e-19 $X=2.74 $Y=2.16
r96 31 34 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.74 $Y=1.615
+ $X2=1.74 $Y2=1.78
r97 31 33 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.74 $Y=1.615
+ $X2=1.74 $Y2=1.45
r98 28 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.74
+ $Y=1.615 $X2=1.74 $Y2=1.615
r99 23 25 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.815 $Y=2.235
+ $X2=2.815 $Y2=2.63
r100 22 27 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.21 $Y=2.16
+ $X2=2.135 $Y2=2.16
r101 21 23 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.74 $Y=2.16
+ $X2=2.815 $Y2=2.235
r102 21 22 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.74 $Y=2.16
+ $X2=2.21 $Y2=2.16
r103 18 27 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.135 $Y=2.235
+ $X2=2.135 $Y2=2.16
r104 18 20 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.135 $Y=2.235
+ $X2=2.135 $Y2=2.63
r105 15 17 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.06 $Y=1.06
+ $X2=2.06 $Y2=0.775
r106 13 27 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.06 $Y=2.16
+ $X2=2.135 $Y2=2.16
r107 13 14 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=2.06 $Y=2.16
+ $X2=1.905 $Y2=2.16
r108 12 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.83 $Y=2.085
+ $X2=1.905 $Y2=2.16
r109 12 34 156.394 $w=1.5e-07 $l=3.05e-07 $layer=POLY_cond $X=1.83 $Y=2.085
+ $X2=1.83 $Y2=1.78
r110 10 26 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.725 $Y=1.135
+ $X2=1.65 $Y2=1.135
r111 9 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.985 $Y=1.135
+ $X2=2.06 $Y2=1.06
r112 9 10 133.319 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=1.985 $Y=1.135
+ $X2=1.725 $Y2=1.135
r113 7 26 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.65 $Y=1.21
+ $X2=1.65 $Y2=1.135
r114 7 33 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=1.65 $Y=1.21
+ $X2=1.65 $Y2=1.45
r115 5 26 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.575 $Y=1.135
+ $X2=1.65 $Y2=1.135
r116 5 6 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.575 $Y=1.135
+ $X2=1.095 $Y2=1.135
r117 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.02 $Y=1.06
+ $X2=1.095 $Y2=1.135
r118 1 3 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.02 $Y=1.06 $X2=1.02
+ $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_LS__SEDFXBP_2%A_575_87# 1 2 9 12 13 15 16 18 19 20 21 23
+ 25 28 30 32 35 37 39 40 45 47 51 54 55 58 59 63 66 67 73 80 81 87
c290 80 0 1.25679e-19 $X=3.04 $Y=1.68
c291 73 0 1.80649e-19 $X=15.12 $Y=1.665
c292 66 0 8.32079e-20 $X=14.975 $Y=1.665
c293 30 0 1.4807e-19 $X=16.325 $Y=1.765
c294 20 0 4.92549e-20 $X=13.345 $Y=0.94
c295 13 0 1.69943e-19 $X=3.205 $Y=2.235
r296 95 96 3.23498 $w=7.09e-07 $l=1.88e-07 $layer=LI1_cond $X=14.855 $Y=2.217
+ $X2=14.855 $Y2=2.405
r297 94 95 3.9921 $w=7.09e-07 $l=2.32e-07 $layer=LI1_cond $X=14.855 $Y=1.985
+ $X2=14.855 $Y2=2.217
r298 87 88 4.74877 $w=4.06e-07 $l=4e-08 $layer=POLY_cond $X=16.735 $Y=1.532
+ $X2=16.775 $Y2=1.532
r299 84 85 2.37438 $w=4.06e-07 $l=2e-08 $layer=POLY_cond $X=16.305 $Y=1.532
+ $X2=16.325 $Y2=1.532
r300 79 81 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.04 $Y=1.68
+ $X2=3.205 $Y2=1.68
r301 79 80 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.04
+ $Y=1.68 $X2=3.04 $Y2=1.68
r302 76 79 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.95 $Y=1.68 $X2=3.04
+ $Y2=1.68
r303 74 94 5.50635 $w=7.09e-07 $l=3.2e-07 $layer=LI1_cond $X=14.855 $Y=1.665
+ $X2=14.855 $Y2=1.985
r304 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.12 $Y=1.665
+ $X2=15.12 $Y2=1.665
r305 69 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=1.665
+ $X2=3.12 $Y2=1.665
r306 67 69 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.265 $Y=1.665
+ $X2=3.12 $Y2=1.665
r307 66 73 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=14.975 $Y=1.665
+ $X2=15.12 $Y2=1.665
r308 66 67 14.4925 $w=1.4e-07 $l=1.171e-05 $layer=MET1_cond $X=14.975 $Y=1.665
+ $X2=3.265 $Y2=1.665
r309 64 87 40.3645 $w=4.06e-07 $l=3.4e-07 $layer=POLY_cond $X=16.395 $Y=1.532
+ $X2=16.735 $Y2=1.532
r310 64 85 8.31034 $w=4.06e-07 $l=7e-08 $layer=POLY_cond $X=16.395 $Y=1.532
+ $X2=16.325 $Y2=1.532
r311 63 64 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=16.395
+ $Y=1.465 $X2=16.395 $Y2=1.465
r312 60 63 10.4924 $w=3.33e-07 $l=3.05e-07 $layer=LI1_cond $X=16.09 $Y=1.467
+ $X2=16.395 $Y2=1.467
r313 57 60 4.05585 $w=1.9e-07 $l=1.68e-07 $layer=LI1_cond $X=16.09 $Y=1.635
+ $X2=16.09 $Y2=1.467
r314 57 58 39.9856 $w=1.88e-07 $l=6.85e-07 $layer=LI1_cond $X=16.09 $Y=1.635
+ $X2=16.09 $Y2=2.32
r315 56 96 9.40575 $w=1.7e-07 $l=3.8e-07 $layer=LI1_cond $X=15.235 $Y=2.405
+ $X2=14.855 $Y2=2.405
r316 55 58 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=15.995 $Y=2.405
+ $X2=16.09 $Y2=2.32
r317 55 56 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=15.995 $Y=2.405
+ $X2=15.235 $Y2=2.405
r318 54 74 10.2197 $w=7.09e-07 $l=1.5906e-07 $layer=LI1_cond $X=14.75 $Y=1.55
+ $X2=14.855 $Y2=1.665
r319 54 59 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=14.75 $Y=1.55
+ $X2=14.75 $Y2=1.13
r320 49 59 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=14.67 $Y=0.965
+ $X2=14.67 $Y2=1.13
r321 49 51 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=14.67 $Y=0.965
+ $X2=14.67 $Y2=0.515
r322 45 96 4.4124 $w=7.09e-07 $l=2.38747e-07 $layer=LI1_cond $X=14.655 $Y=2.49
+ $X2=14.855 $Y2=2.405
r323 45 47 10.404 $w=3.58e-07 $l=3.25e-07 $layer=LI1_cond $X=14.655 $Y=2.49
+ $X2=14.655 $Y2=2.815
r324 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.75
+ $Y=2.215 $X2=13.75 $Y2=2.215
r325 40 95 5.32966 $w=3.25e-07 $l=3.8e-07 $layer=LI1_cond $X=14.475 $Y=2.217
+ $X2=14.855 $Y2=2.217
r326 40 42 25.7083 $w=3.23e-07 $l=7.25e-07 $layer=LI1_cond $X=14.475 $Y=2.217
+ $X2=13.75 $Y2=2.217
r327 37 88 26.2263 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=16.775 $Y=1.765
+ $X2=16.775 $Y2=1.532
r328 37 39 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=16.775 $Y=1.765
+ $X2=16.775 $Y2=2.4
r329 33 87 26.2263 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=16.735 $Y=1.3
+ $X2=16.735 $Y2=1.532
r330 33 35 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=16.735 $Y=1.3
+ $X2=16.735 $Y2=0.74
r331 30 85 26.2263 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=16.325 $Y=1.765
+ $X2=16.325 $Y2=1.532
r332 30 32 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=16.325 $Y=1.765
+ $X2=16.325 $Y2=2.4
r333 26 84 26.2263 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=16.305 $Y=1.3
+ $X2=16.305 $Y2=1.532
r334 26 28 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=16.305 $Y=1.3
+ $X2=16.305 $Y2=0.74
r335 25 43 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=13.84 $Y=2.05
+ $X2=13.75 $Y2=2.215
r336 24 25 530.713 $w=1.5e-07 $l=1.035e-06 $layer=POLY_cond $X=13.84 $Y=1.015
+ $X2=13.84 $Y2=2.05
r337 21 43 52.2586 $w=2.99e-07 $l=2.7157e-07 $layer=POLY_cond $X=13.705 $Y=2.465
+ $X2=13.75 $Y2=2.215
r338 21 23 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=13.705 $Y=2.465
+ $X2=13.705 $Y2=2.75
r339 19 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=13.765 $Y=0.94
+ $X2=13.84 $Y2=1.015
r340 19 20 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=13.765 $Y=0.94
+ $X2=13.345 $Y2=0.94
r341 16 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=13.27 $Y=0.865
+ $X2=13.345 $Y2=0.94
r342 16 18 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=13.27 $Y=0.865
+ $X2=13.27 $Y2=0.58
r343 13 15 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.205 $Y=2.235
+ $X2=3.205 $Y2=2.63
r344 12 13 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.205 $Y=2.145
+ $X2=3.205 $Y2=2.235
r345 11 81 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.205 $Y=1.845
+ $X2=3.205 $Y2=1.68
r346 11 12 116.613 $w=1.8e-07 $l=3e-07 $layer=POLY_cond $X=3.205 $Y=1.845
+ $X2=3.205 $Y2=2.145
r347 7 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.95 $Y=1.515
+ $X2=2.95 $Y2=1.68
r348 7 9 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=2.95 $Y=1.515
+ $X2=2.95 $Y2=0.775
r349 2 94 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=14.49
+ $Y=1.84 $X2=14.64 $Y2=1.985
r350 2 47 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=14.49
+ $Y=1.84 $X2=14.64 $Y2=2.815
r351 1 51 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=14.53
+ $Y=0.37 $X2=14.67 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__SEDFXBP_2%A_661_87# 1 2 7 9 10 11 12 14 17 18 19 22
+ 25 28 30 34 35 38 43 46 47
c111 46 0 1.27569e-19 $X=5.97 $Y=1.58
r112 46 49 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=5.97 $Y=1.58
+ $X2=5.97 $Y2=1.765
r113 46 47 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.97
+ $Y=1.58 $X2=5.97 $Y2=1.58
r114 40 43 5.37015 $w=4.88e-07 $l=2.2e-07 $layer=LI1_cond $X=4.22 $Y=2.49
+ $X2=4.44 $Y2=2.49
r115 37 39 8.79328 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=4.18 $Y=1.89
+ $X2=4.18 $Y2=2.055
r116 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.18
+ $Y=1.89 $X2=4.18 $Y2=1.89
r117 35 37 5.76222 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=4.18 $Y=1.765
+ $X2=4.18 $Y2=1.89
r118 33 34 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.18
+ $Y=0.53 $X2=4.18 $Y2=0.53
r119 31 35 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.305 $Y=1.765
+ $X2=4.18 $Y2=1.765
r120 30 49 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.805 $Y=1.765
+ $X2=5.97 $Y2=1.765
r121 30 31 97.861 $w=1.68e-07 $l=1.5e-06 $layer=LI1_cond $X=5.805 $Y=1.765
+ $X2=4.305 $Y2=1.765
r122 26 33 3.15958 $w=4.05e-07 $l=1.75e-07 $layer=LI1_cond $X=4.305 $Y=0.807
+ $X2=4.18 $Y2=0.687
r123 26 28 9.10572 $w=4.03e-07 $l=3.2e-07 $layer=LI1_cond $X=4.305 $Y=0.807
+ $X2=4.625 $Y2=0.807
r124 25 40 7.03003 $w=1.7e-07 $l=2.45e-07 $layer=LI1_cond $X=4.22 $Y=2.245
+ $X2=4.22 $Y2=2.49
r125 25 39 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=4.22 $Y=2.245
+ $X2=4.22 $Y2=2.055
r126 23 38 118.906 $w=3.3e-07 $l=6.8e-07 $layer=POLY_cond $X=4.18 $Y=1.21
+ $X2=4.18 $Y2=1.89
r127 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.18
+ $Y=1.21 $X2=4.18 $Y2=1.21
r128 20 35 3.91831 $w=2.48e-07 $l=8.5e-08 $layer=LI1_cond $X=4.18 $Y=1.68
+ $X2=4.18 $Y2=1.765
r129 20 22 21.6659 $w=2.48e-07 $l=4.7e-07 $layer=LI1_cond $X=4.18 $Y=1.68
+ $X2=4.18 $Y2=1.21
r130 19 33 4.16548 $w=2.5e-07 $l=3.23e-07 $layer=LI1_cond $X=4.18 $Y=1.01
+ $X2=4.18 $Y2=0.687
r131 19 22 9.21954 $w=2.48e-07 $l=2e-07 $layer=LI1_cond $X=4.18 $Y=1.01 $X2=4.18
+ $Y2=1.21
r132 18 47 36.0236 $w=4.4e-07 $l=2.85e-07 $layer=POLY_cond $X=5.915 $Y=1.865
+ $X2=5.915 $Y2=1.58
r133 17 23 10.1687 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.18 $Y=1.135
+ $X2=4.18 $Y2=1.21
r134 15 34 92.6765 $w=3.3e-07 $l=5.3e-07 $layer=POLY_cond $X=4.18 $Y=1.06
+ $X2=4.18 $Y2=0.53
r135 15 17 10.1687 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.18 $Y=1.06
+ $X2=4.18 $Y2=1.135
r136 12 18 44.0028 $w=3.56e-07 $l=3.84545e-07 $layer=POLY_cond $X=5.785 $Y=2.19
+ $X2=5.915 $Y2=1.865
r137 12 14 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=5.785 $Y=2.19
+ $X2=5.785 $Y2=2.585
r138 10 17 16.9349 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.015 $Y=1.135
+ $X2=4.18 $Y2=1.135
r139 10 11 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.015 $Y=1.135
+ $X2=3.455 $Y2=1.135
r140 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.38 $Y=1.06
+ $X2=3.455 $Y2=1.135
r141 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.38 $Y=1.06 $X2=3.38
+ $Y2=0.775
r142 2 43 600 $w=1.7e-07 $l=2.88531e-07 $layer=licon1_PDIFF $count=1 $X=4.295
+ $Y=2.265 $X2=4.44 $Y2=2.49
r143 1 28 182 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_NDIFF $count=1 $X=4.48
+ $Y=0.625 $X2=4.625 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LS__SEDFXBP_2%SCD 2 3 5 8 10 13
r46 13 16 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.29 $Y=1.345
+ $X2=5.29 $Y2=1.51
r47 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.29 $Y=1.345
+ $X2=5.29 $Y2=1.18
r48 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.29
+ $Y=1.345 $X2=5.29 $Y2=1.345
r49 10 14 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=5.52 $Y=1.345
+ $X2=5.29 $Y2=1.345
r50 8 15 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=5.38 $Y=0.835
+ $X2=5.38 $Y2=1.18
r51 3 5 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=5.365 $Y=2.19
+ $X2=5.365 $Y2=2.585
r52 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.365 $Y=2.1 $X2=5.365
+ $Y2=2.19
r53 2 16 229.339 $w=1.8e-07 $l=5.9e-07 $layer=POLY_cond $X=5.365 $Y=2.1
+ $X2=5.365 $Y2=1.51
.ends

.subckt PM_SKY130_FD_SC_LS__SEDFXBP_2%SCE 1 3 4 5 7 8 11 15 16 17 20 22 25 26
c83 20 0 1.27569e-19 $X=5.77 $Y=0.835
c84 1 0 3.24615e-19 $X=3.655 $Y=3.025
r85 25 28 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.75 $Y=1.345
+ $X2=4.75 $Y2=1.51
r86 25 27 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.75 $Y=1.345
+ $X2=4.75 $Y2=1.18
r87 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.75
+ $Y=1.345 $X2=4.75 $Y2=1.345
r88 22 26 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=4.56 $Y=1.345
+ $X2=4.75 $Y2=1.345
r89 18 20 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=5.77 $Y=0.255
+ $X2=5.77 $Y2=0.835
r90 16 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.695 $Y=0.18
+ $X2=5.77 $Y2=0.255
r91 16 17 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=5.695 $Y=0.18
+ $X2=4.915 $Y2=0.18
r92 15 27 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=4.84 $Y=0.835
+ $X2=4.84 $Y2=1.18
r93 12 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.84 $Y=0.255
+ $X2=4.915 $Y2=0.18
r94 12 15 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=4.84 $Y=0.255
+ $X2=4.84 $Y2=0.835
r95 9 11 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=4.675 $Y=2.98
+ $X2=4.675 $Y2=2.585
r96 8 11 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=4.675 $Y=2.19
+ $X2=4.675 $Y2=2.585
r97 7 8 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=4.675 $Y=2.1 $X2=4.675
+ $Y2=2.19
r98 7 28 229.339 $w=1.8e-07 $l=5.9e-07 $layer=POLY_cond $X=4.675 $Y=2.1
+ $X2=4.675 $Y2=1.51
r99 4 9 26.9307 $w=1.5e-07 $l=1.58745e-07 $layer=POLY_cond $X=4.585 $Y=3.1
+ $X2=4.675 $Y2=2.98
r100 4 5 438.415 $w=1.5e-07 $l=8.55e-07 $layer=POLY_cond $X=4.585 $Y=3.1
+ $X2=3.73 $Y2=3.1
r101 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.655 $Y=3.025
+ $X2=3.73 $Y2=3.1
r102 1 3 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.655 $Y=3.025
+ $X2=3.655 $Y2=2.63
.ends

.subckt PM_SKY130_FD_SC_LS__SEDFXBP_2%CLK 1 3 4 6 7
r36 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.87
+ $Y=1.385 $X2=6.87 $Y2=1.385
r37 7 11 3.05058 $w=3.38e-07 $l=9e-08 $layer=LI1_cond $X=6.875 $Y=1.295
+ $X2=6.875 $Y2=1.385
r38 4 10 38.9026 $w=2.7e-07 $l=1.67481e-07 $layer=POLY_cond $X=6.865 $Y=1.22
+ $X2=6.87 $Y2=1.385
r39 4 6 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=6.865 $Y=1.22 $X2=6.865
+ $Y2=0.74
r40 1 10 77.2841 $w=2.7e-07 $l=4.15812e-07 $layer=POLY_cond $X=6.795 $Y=1.765
+ $X2=6.87 $Y2=1.385
r41 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.795 $Y=1.765
+ $X2=6.795 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__SEDFXBP_2%A_1586_74# 1 2 7 9 10 12 15 18 19 21 24 26
+ 27 28 34 37 40 41 43 46 47 48 50 51 52 53 55 58 60 61 64 66 67 70 74 84
c239 84 0 5.95143e-20 $X=12.37 $Y=1.635
c240 70 0 9.34686e-20 $X=13.36 $Y=1.215
c241 64 0 1.97544e-19 $X=8.89 $Y=2.14
c242 60 0 1.82067e-19 $X=8.89 $Y=1.98
c243 37 0 1.94394e-19 $X=9.65 $Y=0.85
c244 19 0 1.60159e-19 $X=13.285 $Y=2.465
c245 18 0 1.09438e-19 $X=13.285 $Y=2.375
r246 74 88 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=13.36 $Y=1.39
+ $X2=13.36 $Y2=1.555
r247 73 74 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.36
+ $Y=1.39 $X2=13.36 $Y2=1.39
r248 70 73 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=13.36 $Y=1.215
+ $X2=13.36 $Y2=1.39
r249 68 69 15.5982 $w=2.19e-07 $l=2.8e-07 $layer=LI1_cond $X=12.23 $Y=0.935
+ $X2=12.23 $Y2=1.215
r250 64 77 47.886 $w=3.07e-07 $l=3.05e-07 $layer=POLY_cond $X=8.89 $Y=2.22
+ $X2=9.195 $Y2=2.22
r251 63 64 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.89
+ $Y=2.14 $X2=8.89 $Y2=2.14
r252 60 63 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=8.89 $Y=1.98
+ $X2=8.89 $Y2=2.14
r253 60 61 8.28756 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=8.89 $Y=1.98
+ $X2=8.89 $Y2=1.82
r254 59 69 2.22295 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=12.38 $Y=1.215
+ $X2=12.23 $Y2=1.215
r255 58 70 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.195 $Y=1.215
+ $X2=13.36 $Y2=1.215
r256 58 59 53.1711 $w=1.68e-07 $l=8.15e-07 $layer=LI1_cond $X=13.195 $Y=1.215
+ $X2=12.38 $Y2=1.215
r257 56 84 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=12.26 $Y=1.635
+ $X2=12.37 $Y2=1.635
r258 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.26
+ $Y=1.635 $X2=12.26 $Y2=1.635
r259 53 69 4.36852 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.23 $Y=1.3 $X2=12.23
+ $Y2=1.215
r260 53 55 12.8689 $w=2.98e-07 $l=3.35e-07 $layer=LI1_cond $X=12.23 $Y=1.3
+ $X2=12.23 $Y2=1.635
r261 51 68 2.22295 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=12.08 $Y=0.935
+ $X2=12.23 $Y2=0.935
r262 51 52 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=12.08 $Y=0.935
+ $X2=11.54 $Y2=0.935
r263 50 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.455 $Y=0.85
+ $X2=11.54 $Y2=0.935
r264 49 50 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=11.455 $Y=0.425
+ $X2=11.455 $Y2=0.85
r265 47 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.37 $Y=0.34
+ $X2=11.455 $Y2=0.425
r266 47 48 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=11.37 $Y=0.34
+ $X2=10.86 $Y2=0.34
r267 45 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.775 $Y=0.425
+ $X2=10.86 $Y2=0.34
r268 45 46 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=10.775 $Y=0.425
+ $X2=10.775 $Y2=0.85
r269 44 67 2.45049 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=9.855 $Y=0.935
+ $X2=9.71 $Y2=0.935
r270 43 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.69 $Y=0.935
+ $X2=10.775 $Y2=0.85
r271 43 44 54.4759 $w=1.68e-07 $l=8.35e-07 $layer=LI1_cond $X=10.69 $Y=0.935
+ $X2=9.855 $Y2=0.935
r272 41 78 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.69 $Y=1.18
+ $X2=9.525 $Y2=1.18
r273 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.69
+ $Y=1.18 $X2=9.69 $Y2=1.18
r274 38 67 3.98977 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.71 $Y=1.02
+ $X2=9.71 $Y2=0.935
r275 38 40 6.35831 $w=2.88e-07 $l=1.6e-07 $layer=LI1_cond $X=9.71 $Y=1.02
+ $X2=9.71 $Y2=1.18
r276 37 67 3.98977 $w=2.3e-07 $l=1.11018e-07 $layer=LI1_cond $X=9.65 $Y=0.85
+ $X2=9.71 $Y2=0.935
r277 36 37 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=9.65 $Y=0.425
+ $X2=9.65 $Y2=0.85
r278 35 66 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.055 $Y=0.34
+ $X2=8.97 $Y2=0.34
r279 34 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.565 $Y=0.34
+ $X2=9.65 $Y2=0.425
r280 34 35 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=9.565 $Y=0.34
+ $X2=9.055 $Y2=0.34
r281 32 66 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.97 $Y=0.425
+ $X2=8.97 $Y2=0.34
r282 32 61 91.0107 $w=1.68e-07 $l=1.395e-06 $layer=LI1_cond $X=8.97 $Y=0.425
+ $X2=8.97 $Y2=1.82
r283 28 60 0.903439 $w=3.2e-07 $l=1.65e-07 $layer=LI1_cond $X=8.725 $Y=1.98
+ $X2=8.89 $Y2=1.98
r284 28 30 11.3444 $w=3.18e-07 $l=3.15e-07 $layer=LI1_cond $X=8.725 $Y=1.98
+ $X2=8.41 $Y2=1.98
r285 26 66 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.885 $Y=0.34
+ $X2=8.97 $Y2=0.34
r286 26 27 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=8.885 $Y=0.34
+ $X2=8.235 $Y2=0.34
r287 22 27 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.07 $Y=0.425
+ $X2=8.235 $Y2=0.34
r288 22 24 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=8.07 $Y=0.425
+ $X2=8.07 $Y2=0.515
r289 19 21 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=13.285 $Y=2.465
+ $X2=13.285 $Y2=2.75
r290 18 19 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=13.285 $Y=2.375
+ $X2=13.285 $Y2=2.465
r291 18 88 318.742 $w=1.8e-07 $l=8.2e-07 $layer=POLY_cond $X=13.285 $Y=2.375
+ $X2=13.285 $Y2=1.555
r292 13 84 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=12.37 $Y=1.47
+ $X2=12.37 $Y2=1.635
r293 13 15 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=12.37 $Y=1.47
+ $X2=12.37 $Y2=0.69
r294 10 78 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.525 $Y=1.015
+ $X2=9.525 $Y2=1.18
r295 10 12 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=9.525 $Y=1.015
+ $X2=9.525 $Y2=0.695
r296 7 77 19.5117 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=9.195 $Y=2.465
+ $X2=9.195 $Y2=2.22
r297 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=9.195 $Y=2.465
+ $X2=9.195 $Y2=2.75
r298 2 30 600 $w=1.7e-07 $l=2.43721e-07 $layer=licon1_PDIFF $count=1 $X=8.26
+ $Y=1.84 $X2=8.41 $Y2=2.02
r299 1 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.93
+ $Y=0.37 $X2=8.07 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__SEDFXBP_2%A_1374_368# 1 2 11 13 15 17 18 22 24 27 28
+ 30 31 33 36 38 39 40 46 49 51 55 56 57 61 67 73
c190 67 0 1.09438e-19 $X=12.82 $Y=1.635
c191 61 0 1.97544e-19 $X=9.69 $Y=2.195
c192 46 0 1.60159e-19 $X=12.55 $Y=2.475
c193 31 0 9.34686e-20 $X=12.75 $Y=1.885
c194 27 0 1.82067e-19 $X=9.6 $Y=2.03
c195 22 0 1.94394e-19 $X=8.845 $Y=0.695
c196 13 0 5.76754e-20 $X=8.095 $Y=1.66
r197 67 68 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.82
+ $Y=1.635 $X2=12.82 $Y2=1.635
r198 64 67 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=12.635 $Y=1.635
+ $X2=12.82 $Y2=1.635
r199 61 62 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.69
+ $Y=2.195 $X2=9.69 $Y2=2.195
r200 55 58 9.0362 $w=4.38e-07 $l=3.45e-07 $layer=LI1_cond $X=7.435 $Y=1.635
+ $X2=7.435 $Y2=1.98
r201 55 57 8.83531 $w=4.38e-07 $l=1.65e-07 $layer=LI1_cond $X=7.435 $Y=1.635
+ $X2=7.435 $Y2=1.47
r202 55 56 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.49
+ $Y=1.635 $X2=7.49 $Y2=1.635
r203 53 57 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=7.3 $Y=1.01 $X2=7.3
+ $Y2=1.47
r204 51 53 17.7356 $w=4.68e-07 $l=4.95e-07 $layer=LI1_cond $X=7.15 $Y=0.515
+ $X2=7.15 $Y2=1.01
r205 48 64 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.635 $Y=1.8
+ $X2=12.635 $Y2=1.635
r206 48 49 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=12.635 $Y=1.8
+ $X2=12.635 $Y2=2.39
r207 47 61 11.8611 $w=2.88e-07 $l=3.58887e-07 $layer=LI1_cond $X=9.925 $Y=2.475
+ $X2=9.745 $Y2=2.195
r208 46 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=12.55 $Y=2.475
+ $X2=12.635 $Y2=2.39
r209 46 47 171.257 $w=1.68e-07 $l=2.625e-06 $layer=LI1_cond $X=12.55 $Y=2.475
+ $X2=9.925 $Y2=2.475
r210 40 58 2.60351 $w=3.2e-07 $l=2.2e-07 $layer=LI1_cond $X=7.215 $Y=1.98
+ $X2=7.435 $Y2=1.98
r211 40 42 7.0227 $w=3.18e-07 $l=1.95e-07 $layer=LI1_cond $X=7.215 $Y=1.98
+ $X2=7.02 $Y2=1.98
r212 34 68 38.5562 $w=2.99e-07 $l=1.92678e-07 $layer=POLY_cond $X=12.88 $Y=1.47
+ $X2=12.82 $Y2=1.635
r213 34 36 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=12.88 $Y=1.47
+ $X2=12.88 $Y2=0.58
r214 31 68 52.2586 $w=2.99e-07 $l=2.82843e-07 $layer=POLY_cond $X=12.75 $Y=1.885
+ $X2=12.82 $Y2=1.635
r215 31 33 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=12.75 $Y=1.885
+ $X2=12.75 $Y2=2.46
r216 28 62 55.8646 $w=2.93e-07 $l=2.91633e-07 $layer=POLY_cond $X=9.645 $Y=2.465
+ $X2=9.69 $Y2=2.195
r217 28 30 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=9.645 $Y=2.465
+ $X2=9.645 $Y2=2.75
r218 27 62 38.5916 $w=2.93e-07 $l=2.05122e-07 $layer=POLY_cond $X=9.6 $Y=2.03
+ $X2=9.69 $Y2=2.195
r219 26 27 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=9.6 $Y=1.735
+ $X2=9.6 $Y2=2.03
r220 25 39 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.92 $Y=1.66
+ $X2=8.845 $Y2=1.66
r221 24 26 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.525 $Y=1.66
+ $X2=9.6 $Y2=1.735
r222 24 25 310.223 $w=1.5e-07 $l=6.05e-07 $layer=POLY_cond $X=9.525 $Y=1.66
+ $X2=8.92 $Y2=1.66
r223 20 39 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.845 $Y=1.585
+ $X2=8.845 $Y2=1.66
r224 20 22 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=8.845 $Y=1.585
+ $X2=8.845 $Y2=0.695
r225 19 38 20.4101 $w=1.5e-07 $l=9.72111e-08 $layer=POLY_cond $X=8.275 $Y=1.66
+ $X2=8.185 $Y2=1.675
r226 18 39 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.77 $Y=1.66
+ $X2=8.845 $Y2=1.66
r227 18 19 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=8.77 $Y=1.66
+ $X2=8.275 $Y2=1.66
r228 15 38 5.30422 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=8.185 $Y=1.765
+ $X2=8.185 $Y2=1.675
r229 15 17 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.185 $Y=1.765
+ $X2=8.185 $Y2=2.4
r230 13 38 20.4101 $w=1.5e-07 $l=9.72111e-08 $layer=POLY_cond $X=8.095 $Y=1.66
+ $X2=8.185 $Y2=1.675
r231 13 73 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.095 $Y=1.66
+ $X2=7.93 $Y2=1.66
r232 9 73 28.1815 $w=2.65e-07 $l=7.5e-08 $layer=POLY_cond $X=7.855 $Y=1.602
+ $X2=7.93 $Y2=1.602
r233 9 56 82.6235 $w=2.65e-07 $l=3.65e-07 $layer=POLY_cond $X=7.855 $Y=1.602
+ $X2=7.49 $Y2=1.602
r234 9 11 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=7.855 $Y=1.47
+ $X2=7.855 $Y2=0.74
r235 2 42 600 $w=1.7e-07 $l=2.43721e-07 $layer=licon1_PDIFF $count=1 $X=6.87
+ $Y=1.84 $X2=7.02 $Y2=2.02
r236 1 51 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.94
+ $Y=0.37 $X2=7.08 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__SEDFXBP_2%A_2013_71# 1 2 9 12 13 15 18 19 20 22 23
+ 25 26 28 34 37 38 40 41 43 47
c114 47 0 2.55325e-20 $X=10.23 $Y=1.355
c115 43 0 1.43495e-19 $X=10.23 $Y=1.275
c116 40 0 5.95143e-20 $X=11.72 $Y=1.355
r117 49 50 9.1748 $w=2.46e-07 $l=1.85e-07 $layer=LI1_cond $X=11.115 $Y=1.355
+ $X2=11.3 $Y2=1.355
r118 47 53 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.23 $Y=1.355
+ $X2=10.23 $Y2=1.52
r119 47 52 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.23 $Y=1.355
+ $X2=10.23 $Y2=1.19
r120 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.23
+ $Y=1.355 $X2=10.23 $Y2=1.355
r121 43 46 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=10.23 $Y=1.275
+ $X2=10.23 $Y2=1.355
r122 40 41 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=11.72
+ $Y=1.355 $X2=11.72 $Y2=1.355
r123 38 50 3.95924 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.385 $Y=1.355
+ $X2=11.3 $Y2=1.355
r124 38 40 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=11.385 $Y=1.355
+ $X2=11.72 $Y2=1.355
r125 36 50 2.90119 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.3 $Y=1.52
+ $X2=11.3 $Y2=1.355
r126 36 37 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=11.3 $Y=1.52
+ $X2=11.3 $Y2=2.05
r127 32 49 2.90119 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.115 $Y=1.19
+ $X2=11.115 $Y2=1.355
r128 32 34 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=11.115 $Y=1.19
+ $X2=11.115 $Y2=0.805
r129 28 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.215 $Y=2.135
+ $X2=11.3 $Y2=2.05
r130 28 30 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=11.215 $Y=2.135
+ $X2=10.925 $Y2=2.135
r131 27 43 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.395 $Y=1.275
+ $X2=10.23 $Y2=1.275
r132 26 49 5.39088 $w=2.46e-07 $l=1.18427e-07 $layer=LI1_cond $X=11.03 $Y=1.275
+ $X2=11.115 $Y2=1.355
r133 26 27 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=11.03 $Y=1.275
+ $X2=10.395 $Y2=1.275
r134 23 25 134.96 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=12.01 $Y=1.11
+ $X2=12.01 $Y2=0.69
r135 20 22 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=11.795 $Y=1.885
+ $X2=11.795 $Y2=2.46
r136 19 20 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=11.795 $Y=1.795
+ $X2=11.795 $Y2=1.885
r137 18 23 37.9597 $w=2.73e-07 $l=3.7229e-07 $layer=POLY_cond $X=11.795 $Y=1.39
+ $X2=12.01 $Y2=1.11
r138 18 41 13.2418 $w=2.73e-07 $l=7.5e-08 $layer=POLY_cond $X=11.795 $Y=1.39
+ $X2=11.72 $Y2=1.39
r139 18 19 106.895 $w=1.8e-07 $l=2.75e-07 $layer=POLY_cond $X=11.795 $Y=1.52
+ $X2=11.795 $Y2=1.795
r140 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=10.155 $Y=2.465
+ $X2=10.155 $Y2=2.75
r141 12 13 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=10.155 $Y=2.375
+ $X2=10.155 $Y2=2.465
r142 12 53 332.347 $w=1.8e-07 $l=8.55e-07 $layer=POLY_cond $X=10.155 $Y=2.375
+ $X2=10.155 $Y2=1.52
r143 9 52 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=10.14 $Y=0.695
+ $X2=10.14 $Y2=1.19
r144 2 30 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=10.775
+ $Y=1.99 $X2=10.925 $Y2=2.135
r145 1 34 182 $w=1.7e-07 $l=5.00125e-07 $layer=licon1_NDIFF $count=1 $X=10.975
+ $Y=0.37 $X2=11.115 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LS__SEDFXBP_2%A_1784_97# 1 2 7 9 12 16 20 22 24 25 28
c85 7 0 1.43495e-19 $X=10.7 $Y=1.915
r86 28 31 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=10.775 $Y=1.665
+ $X2=10.775 $Y2=1.775
r87 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.775
+ $Y=1.665 $X2=10.775 $Y2=1.665
r88 24 25 10.4318 $w=3.58e-07 $l=2.25e-07 $layer=LI1_cond $X=9.405 $Y=2.755
+ $X2=9.405 $Y2=2.53
r89 21 22 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.395 $Y=1.775
+ $X2=9.31 $Y2=1.775
r90 20 31 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.61 $Y=1.775
+ $X2=10.775 $Y2=1.775
r91 20 21 79.2674 $w=1.68e-07 $l=1.215e-06 $layer=LI1_cond $X=10.61 $Y=1.775
+ $X2=9.395 $Y2=1.775
r92 18 22 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.31 $Y=1.86 $X2=9.31
+ $Y2=1.775
r93 18 25 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.31 $Y=1.86
+ $X2=9.31 $Y2=2.53
r94 14 22 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.31 $Y=1.69 $X2=9.31
+ $Y2=1.775
r95 14 16 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=9.31 $Y=1.69
+ $X2=9.31 $Y2=0.76
r96 10 29 38.5818 $w=3.27e-07 $l=2.12238e-07 $layer=POLY_cond $X=10.9 $Y=1.5
+ $X2=10.792 $Y2=1.665
r97 10 12 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=10.9 $Y=1.5 $X2=10.9
+ $Y2=0.69
r98 7 29 51.1109 $w=3.27e-07 $l=2.92404e-07 $layer=POLY_cond $X=10.7 $Y=1.915
+ $X2=10.792 $Y2=1.665
r99 7 9 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=10.7 $Y=1.915 $X2=10.7
+ $Y2=2.41
r100 2 24 600 $w=1.7e-07 $l=2.80134e-07 $layer=licon1_PDIFF $count=1 $X=9.27
+ $Y=2.54 $X2=9.42 $Y2=2.755
r101 1 16 182 $w=1.7e-07 $l=5.09264e-07 $layer=licon1_NDIFF $count=1 $X=8.92
+ $Y=0.485 $X2=9.31 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_LS__SEDFXBP_2%A_2489_74# 1 2 7 9 12 14 15 16 18 21 25 27
+ 29 32 33 35 37 40 41 42 44 45 47 55
c155 47 0 1.80649e-19 $X=14.33 $Y=1.465
c156 42 0 4.92549e-20 $X=13.325 $Y=1.8
c157 33 0 1.45871e-19 $X=12.585 $Y=0.77
r158 61 62 4.86869 $w=3.96e-07 $l=4e-08 $layer=POLY_cond $X=14.415 $Y=1.532
+ $X2=14.455 $Y2=1.532
r159 53 55 6.89045 $w=4.58e-07 $l=2.65e-07 $layer=LI1_cond $X=12.975 $Y=2.75
+ $X2=13.24 $Y2=2.75
r160 48 61 10.346 $w=3.96e-07 $l=8.5e-08 $layer=POLY_cond $X=14.33 $Y=1.532
+ $X2=14.415 $Y2=1.532
r161 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=14.33
+ $Y=1.465 $X2=14.33 $Y2=1.465
r162 45 58 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=13.78 $Y=1.465
+ $X2=13.78 $Y2=1.8
r163 45 47 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=13.865 $Y=1.465
+ $X2=14.33 $Y2=1.465
r164 44 45 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=13.78 $Y=1.3
+ $X2=13.78 $Y2=1.465
r165 43 44 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=13.78 $Y=0.94
+ $X2=13.78 $Y2=1.3
r166 41 58 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.695 $Y=1.8
+ $X2=13.78 $Y2=1.8
r167 41 42 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=13.695 $Y=1.8
+ $X2=13.325 $Y2=1.8
r168 40 55 6.6364 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=13.24 $Y=2.52
+ $X2=13.24 $Y2=2.75
r169 39 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=13.24 $Y=1.885
+ $X2=13.325 $Y2=1.8
r170 39 40 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=13.24 $Y=1.885
+ $X2=13.24 $Y2=2.52
r171 38 51 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.75 $Y=0.855
+ $X2=12.585 $Y2=0.855
r172 37 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=13.695 $Y=0.855
+ $X2=13.78 $Y2=0.94
r173 37 38 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=13.695 $Y=0.855
+ $X2=12.75 $Y2=0.855
r174 33 51 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.585 $Y=0.77
+ $X2=12.585 $Y2=0.855
r175 33 35 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=12.585 $Y=0.77
+ $X2=12.585 $Y2=0.515
r176 31 32 50.9238 $w=4.07e-07 $l=4.3e-07 $layer=POLY_cond $X=15.445 $Y=1.532
+ $X2=15.875 $Y2=1.532
r177 30 31 2.36855 $w=4.07e-07 $l=2e-08 $layer=POLY_cond $X=15.425 $Y=1.532
+ $X2=15.445 $Y2=1.532
r178 27 32 26.2866 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=15.875 $Y=1.765
+ $X2=15.875 $Y2=1.532
r179 27 29 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=15.875 $Y=1.765
+ $X2=15.875 $Y2=2.4
r180 23 32 26.2866 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=15.875 $Y=1.3
+ $X2=15.875 $Y2=1.532
r181 23 25 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=15.875 $Y=1.3
+ $X2=15.875 $Y2=0.74
r182 19 31 26.2866 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=15.445 $Y=1.3
+ $X2=15.445 $Y2=1.532
r183 19 21 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=15.445 $Y=1.3
+ $X2=15.445 $Y2=0.74
r184 16 30 26.2866 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=15.425 $Y=1.765
+ $X2=15.425 $Y2=1.532
r185 16 18 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=15.425 $Y=1.765
+ $X2=15.425 $Y2=2.4
r186 15 62 10.6098 $w=3.96e-07 $l=1.03199e-07 $layer=POLY_cond $X=14.53 $Y=1.465
+ $X2=14.455 $Y2=1.532
r187 14 30 12.5251 $w=4.07e-07 $l=1.1887e-07 $layer=POLY_cond $X=15.335 $Y=1.465
+ $X2=15.425 $Y2=1.532
r188 14 15 140.763 $w=3.3e-07 $l=8.05e-07 $layer=POLY_cond $X=15.335 $Y=1.465
+ $X2=14.53 $Y2=1.465
r189 10 62 25.6164 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=14.455 $Y=1.3
+ $X2=14.455 $Y2=1.532
r190 10 12 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=14.455 $Y=1.3
+ $X2=14.455 $Y2=0.74
r191 7 61 25.6164 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=14.415 $Y=1.765
+ $X2=14.415 $Y2=1.532
r192 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=14.415 $Y=1.765
+ $X2=14.415 $Y2=2.4
r193 2 53 600 $w=1.7e-07 $l=8.61742e-07 $layer=licon1_PDIFF $count=1 $X=12.825
+ $Y=1.96 $X2=12.975 $Y2=2.75
r194 1 51 182 $w=1.7e-07 $l=5.50568e-07 $layer=licon1_NDIFF $count=1 $X=12.445
+ $Y=0.37 $X2=12.585 $Y2=0.855
r195 1 35 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=12.445
+ $Y=0.37 $X2=12.585 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__SEDFXBP_2%A_32_74# 1 2 3 4 14 17 19 22 23 24 26 27
+ 28 31 36 40 42 45 48
c119 48 0 3.24615e-19 $X=3.43 $Y=2.455
c120 19 0 1.8559e-19 $X=1.485 $Y=2.375
r121 37 40 9.10802 $w=3.08e-07 $l=2.45e-07 $layer=LI1_cond $X=0.17 $Y=0.575
+ $X2=0.415 $Y2=0.575
r122 36 48 4.06715 $w=2.25e-07 $l=1.09087e-07 $layer=LI1_cond $X=3.46 $Y=2.29
+ $X2=3.405 $Y2=2.375
r123 35 45 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.46 $Y=1.345
+ $X2=3.46 $Y2=1.26
r124 35 36 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=3.46 $Y=1.345
+ $X2=3.46 $Y2=2.29
r125 29 45 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.165 $Y=1.26
+ $X2=3.46 $Y2=1.26
r126 29 31 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=3.165 $Y=1.175
+ $X2=3.165 $Y2=0.775
r127 27 48 2.36881 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=3.265 $Y=2.375
+ $X2=3.405 $Y2=2.375
r128 27 28 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=3.265 $Y=2.375
+ $X2=2.335 $Y2=2.375
r129 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.25 $Y=2.46
+ $X2=2.335 $Y2=2.375
r130 25 26 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=2.25 $Y=2.46
+ $X2=2.25 $Y2=2.905
r131 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.165 $Y=2.99
+ $X2=2.25 $Y2=2.905
r132 23 24 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=2.165 $Y=2.99
+ $X2=1.655 $Y2=2.99
r133 22 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.57 $Y=2.905
+ $X2=1.655 $Y2=2.99
r134 21 22 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=1.57 $Y=2.46
+ $X2=1.57 $Y2=2.905
r135 20 42 3.51065 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=0.525 $Y=2.375
+ $X2=0.305 $Y2=2.375
r136 19 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.485 $Y=2.375
+ $X2=1.57 $Y2=2.46
r137 19 20 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.485 $Y=2.375
+ $X2=0.525 $Y2=2.375
r138 15 42 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.305 $Y=2.46
+ $X2=0.305 $Y2=2.375
r139 15 17 0.130959 $w=4.38e-07 $l=5e-09 $layer=LI1_cond $X=0.305 $Y=2.46
+ $X2=0.305 $Y2=2.465
r140 14 42 3.10218 $w=3.05e-07 $l=1.72337e-07 $layer=LI1_cond $X=0.17 $Y=2.29
+ $X2=0.305 $Y2=2.375
r141 13 37 4.25403 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=0.17 $Y=0.73
+ $X2=0.17 $Y2=0.575
r142 13 14 101.775 $w=1.68e-07 $l=1.56e-06 $layer=LI1_cond $X=0.17 $Y=0.73
+ $X2=0.17 $Y2=2.29
r143 4 48 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=3.28
+ $Y=2.31 $X2=3.43 $Y2=2.455
r144 3 17 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.215
+ $Y=2.32 $X2=0.36 $Y2=2.465
r145 2 31 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.025
+ $Y=0.565 $X2=3.165 $Y2=0.775
r146 1 40 182 $w=1.7e-07 $l=3.46194e-07 $layer=licon1_NDIFF $count=1 $X=0.16
+ $Y=0.37 $X2=0.415 $Y2=0.585
.ends

.subckt PM_SKY130_FD_SC_LS__SEDFXBP_2%VPWR 1 2 3 4 5 6 7 8 9 10 11 36 40 44 48
+ 52 56 60 64 68 72 74 76 79 80 82 83 84 86 91 96 108 112 124 131 136 141 147
+ 150 153 156 159 162 165 168 172
r199 171 172 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=17.04 $Y=3.33
+ $X2=17.04 $Y2=3.33
r200 168 169 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=16.08 $Y=3.33
+ $X2=16.08 $Y2=3.33
r201 165 166 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.12 $Y=3.33
+ $X2=15.12 $Y2=3.33
r202 162 163 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.16 $Y=3.33
+ $X2=14.16 $Y2=3.33
r203 159 160 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r204 156 157 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r205 153 154 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r206 150 151 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r207 147 148 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r208 145 172 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=16.56 $Y=3.33
+ $X2=17.04 $Y2=3.33
r209 145 169 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=16.56 $Y=3.33
+ $X2=16.08 $Y2=3.33
r210 144 145 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=16.56 $Y=3.33
+ $X2=16.56 $Y2=3.33
r211 142 168 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=16.265 $Y=3.33
+ $X2=16.1 $Y2=3.33
r212 142 144 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=16.265 $Y=3.33
+ $X2=16.56 $Y2=3.33
r213 141 171 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=16.835 $Y=3.33
+ $X2=17.057 $Y2=3.33
r214 141 144 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=16.835 $Y=3.33
+ $X2=16.56 $Y2=3.33
r215 140 169 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=15.6 $Y=3.33
+ $X2=16.08 $Y2=3.33
r216 140 166 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=15.6 $Y=3.33
+ $X2=15.12 $Y2=3.33
r217 139 140 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.6 $Y=3.33
+ $X2=15.6 $Y2=3.33
r218 137 165 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=15.365 $Y=3.33
+ $X2=15.2 $Y2=3.33
r219 137 139 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=15.365 $Y=3.33
+ $X2=15.6 $Y2=3.33
r220 136 168 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=15.935 $Y=3.33
+ $X2=16.1 $Y2=3.33
r221 136 139 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=15.935 $Y=3.33
+ $X2=15.6 $Y2=3.33
r222 135 166 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.64 $Y=3.33
+ $X2=15.12 $Y2=3.33
r223 135 163 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.64 $Y=3.33
+ $X2=14.16 $Y2=3.33
r224 134 135 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.64 $Y=3.33
+ $X2=14.64 $Y2=3.33
r225 132 162 11.8214 $w=1.7e-07 $l=2.7e-07 $layer=LI1_cond $X=14.305 $Y=3.33
+ $X2=14.035 $Y2=3.33
r226 132 134 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=14.305 $Y=3.33
+ $X2=14.64 $Y2=3.33
r227 131 165 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=15.035 $Y=3.33
+ $X2=15.2 $Y2=3.33
r228 131 134 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=15.035 $Y=3.33
+ $X2=14.64 $Y2=3.33
r229 130 163 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=3.33
+ $X2=14.16 $Y2=3.33
r230 129 130 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=13.68 $Y=3.33
+ $X2=13.68 $Y2=3.33
r231 127 130 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=13.68 $Y2=3.33
r232 126 129 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=11.76 $Y=3.33
+ $X2=13.68 $Y2=3.33
r233 126 127 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r234 124 162 11.8214 $w=1.7e-07 $l=2.7e-07 $layer=LI1_cond $X=13.765 $Y=3.33
+ $X2=14.035 $Y2=3.33
r235 124 129 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=13.765 $Y=3.33
+ $X2=13.68 $Y2=3.33
r236 123 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=11.76 $Y2=3.33
r237 123 160 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=10.32 $Y2=3.33
r238 122 123 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r239 120 159 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.555 $Y=3.33
+ $X2=10.39 $Y2=3.33
r240 120 122 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=10.555 $Y=3.33
+ $X2=11.28 $Y2=3.33
r241 119 160 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=10.32 $Y2=3.33
r242 118 119 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r243 116 157 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=7.92 $Y2=3.33
r244 115 118 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=8.4 $Y=3.33
+ $X2=9.84 $Y2=3.33
r245 115 116 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r246 113 156 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.125 $Y=3.33
+ $X2=7.96 $Y2=3.33
r247 113 115 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=8.125 $Y=3.33
+ $X2=8.4 $Y2=3.33
r248 112 159 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.225 $Y=3.33
+ $X2=10.39 $Y2=3.33
r249 112 118 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=10.225 $Y=3.33
+ $X2=9.84 $Y2=3.33
r250 111 157 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r251 110 111 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r252 108 156 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.795 $Y=3.33
+ $X2=7.96 $Y2=3.33
r253 108 110 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=7.795 $Y=3.33
+ $X2=7.44 $Y2=3.33
r254 107 111 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=7.44 $Y2=3.33
r255 106 107 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r256 104 107 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6.48 $Y2=3.33
r257 104 154 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=5.04 $Y2=3.33
r258 103 106 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=5.52 $Y=3.33
+ $X2=6.48 $Y2=3.33
r259 103 104 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r260 101 153 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.305 $Y=3.33
+ $X2=5.17 $Y2=3.33
r261 101 103 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=5.305 $Y=3.33
+ $X2=5.52 $Y2=3.33
r262 100 154 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=5.04 $Y2=3.33
r263 100 151 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r264 99 100 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r265 97 150 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.755 $Y=3.33
+ $X2=2.63 $Y2=3.33
r266 97 99 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.755 $Y=3.33
+ $X2=3.12 $Y2=3.33
r267 96 153 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.035 $Y=3.33
+ $X2=5.17 $Y2=3.33
r268 96 99 124.936 $w=1.68e-07 $l=1.915e-06 $layer=LI1_cond $X=5.035 $Y=3.33
+ $X2=3.12 $Y2=3.33
r269 95 151 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r270 95 148 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.2 $Y2=3.33
r271 94 95 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r272 92 147 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.315 $Y=3.33
+ $X2=1.19 $Y2=3.33
r273 92 94 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=1.315 $Y=3.33
+ $X2=2.16 $Y2=3.33
r274 91 150 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.505 $Y=3.33
+ $X2=2.63 $Y2=3.33
r275 91 94 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.505 $Y=3.33
+ $X2=2.16 $Y2=3.33
r276 89 148 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r277 88 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r278 86 147 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.065 $Y=3.33
+ $X2=1.19 $Y2=3.33
r279 86 88 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.065 $Y=3.33
+ $X2=0.72 $Y2=3.33
r280 84 119 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=8.64 $Y=3.33
+ $X2=9.84 $Y2=3.33
r281 84 116 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=8.64 $Y=3.33
+ $X2=8.4 $Y2=3.33
r282 82 122 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=11.32 $Y=3.33
+ $X2=11.28 $Y2=3.33
r283 82 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.32 $Y=3.33
+ $X2=11.485 $Y2=3.33
r284 81 126 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=11.65 $Y=3.33
+ $X2=11.76 $Y2=3.33
r285 81 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.65 $Y=3.33
+ $X2=11.485 $Y2=3.33
r286 79 106 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=6.485 $Y=3.33
+ $X2=6.48 $Y2=3.33
r287 79 80 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.485 $Y=3.33
+ $X2=6.61 $Y2=3.33
r288 78 110 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=6.735 $Y=3.33
+ $X2=7.44 $Y2=3.33
r289 78 80 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.735 $Y=3.33
+ $X2=6.61 $Y2=3.33
r290 74 171 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=17 $Y=3.245
+ $X2=17.057 $Y2=3.33
r291 74 76 34.7479 $w=3.28e-07 $l=9.95e-07 $layer=LI1_cond $X=17 $Y=3.245 $X2=17
+ $Y2=2.25
r292 70 168 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=16.1 $Y=3.245
+ $X2=16.1 $Y2=3.33
r293 70 72 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=16.1 $Y=3.245
+ $X2=16.1 $Y2=2.78
r294 66 165 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=15.2 $Y=3.245
+ $X2=15.2 $Y2=3.33
r295 66 68 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=15.2 $Y=3.245
+ $X2=15.2 $Y2=2.78
r296 62 162 2.26835 $w=5.4e-07 $l=8.5e-08 $layer=LI1_cond $X=14.035 $Y=3.245
+ $X2=14.035 $Y2=3.33
r297 62 64 9.52433 $w=5.38e-07 $l=4.3e-07 $layer=LI1_cond $X=14.035 $Y=3.245
+ $X2=14.035 $Y2=2.815
r298 58 83 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.485 $Y=3.245
+ $X2=11.485 $Y2=3.33
r299 58 60 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=11.485 $Y=3.245
+ $X2=11.485 $Y2=2.895
r300 54 159 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.39 $Y=3.245
+ $X2=10.39 $Y2=3.33
r301 54 56 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=10.39 $Y=3.245
+ $X2=10.39 $Y2=2.815
r302 50 156 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.96 $Y=3.245
+ $X2=7.96 $Y2=3.33
r303 50 52 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=7.96 $Y=3.245
+ $X2=7.96 $Y2=2.815
r304 46 80 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.61 $Y=3.245
+ $X2=6.61 $Y2=3.33
r305 46 48 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=6.61 $Y=3.245
+ $X2=6.61 $Y2=2.815
r306 42 153 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.17 $Y=3.245
+ $X2=5.17 $Y2=3.33
r307 42 44 20.7013 $w=2.68e-07 $l=4.85e-07 $layer=LI1_cond $X=5.17 $Y=3.245
+ $X2=5.17 $Y2=2.76
r308 38 150 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.63 $Y=3.245
+ $X2=2.63 $Y2=3.33
r309 38 40 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=2.63 $Y=3.245
+ $X2=2.63 $Y2=2.8
r310 34 147 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.19 $Y=3.245
+ $X2=1.19 $Y2=3.33
r311 34 36 20.283 $w=2.48e-07 $l=4.4e-07 $layer=LI1_cond $X=1.19 $Y=3.245
+ $X2=1.19 $Y2=2.805
r312 11 76 300 $w=1.7e-07 $l=4.79166e-07 $layer=licon1_PDIFF $count=2 $X=16.85
+ $Y=1.84 $X2=17 $Y2=2.25
r313 10 72 600 $w=1.7e-07 $l=1.01223e-06 $layer=licon1_PDIFF $count=1 $X=15.95
+ $Y=1.84 $X2=16.1 $Y2=2.78
r314 9 68 600 $w=1.7e-07 $l=1.0099e-06 $layer=licon1_PDIFF $count=1 $X=15.055
+ $Y=1.84 $X2=15.2 $Y2=2.78
r315 8 64 600 $w=1.7e-07 $l=3.81772e-07 $layer=licon1_PDIFF $count=1 $X=13.78
+ $Y=2.54 $X2=14.035 $Y2=2.815
r316 7 60 600 $w=1.7e-07 $l=1.00489e-06 $layer=licon1_PDIFF $count=1 $X=11.34
+ $Y=1.96 $X2=11.485 $Y2=2.895
r317 6 56 600 $w=1.7e-07 $l=3.45868e-07 $layer=licon1_PDIFF $count=1 $X=10.23
+ $Y=2.54 $X2=10.39 $Y2=2.815
r318 5 52 600 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=7.815
+ $Y=1.84 $X2=7.96 $Y2=2.815
r319 4 48 600 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=6.425
+ $Y=1.84 $X2=6.57 $Y2=2.815
r320 3 44 600 $w=1.7e-07 $l=6.58122e-07 $layer=licon1_PDIFF $count=1 $X=4.75
+ $Y=2.265 $X2=5.13 $Y2=2.76
r321 2 40 600 $w=1.7e-07 $l=6.52917e-07 $layer=licon1_PDIFF $count=1 $X=2.21
+ $Y=2.31 $X2=2.59 $Y2=2.8
r322 1 36 600 $w=1.7e-07 $l=5.54955e-07 $layer=licon1_PDIFF $count=1 $X=1.08
+ $Y=2.32 $X2=1.23 $Y2=2.805
.ends

.subckt PM_SKY130_FD_SC_LS__SEDFXBP_2%A_691_113# 1 2 3 4 5 6 21 24 25 26 28 29
+ 30 33 36 37 38 40 41 42 43 47 49 53 56 59 62 67 68
c186 21 0 1.69943e-19 $X=3.84 $Y=2.415
r187 68 70 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=8.38 $Y=2.395
+ $X2=8.38 $Y2=2.565
r188 58 59 83.8342 $w=1.68e-07 $l=1.285e-06 $layer=LI1_cond $X=3.8 $Y=1.005
+ $X2=3.8 $Y2=2.29
r189 56 58 10.5346 $w=3.83e-07 $l=2.3e-07 $layer=LI1_cond $X=3.692 $Y=0.775
+ $X2=3.692 $Y2=1.005
r190 51 53 4.60977 $w=2.48e-07 $l=1e-07 $layer=LI1_cond $X=8.93 $Y=2.65 $X2=8.93
+ $Y2=2.75
r191 50 70 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.465 $Y=2.565
+ $X2=8.38 $Y2=2.565
r192 49 51 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=8.805 $Y=2.565
+ $X2=8.93 $Y2=2.65
r193 49 50 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=8.805 $Y=2.565
+ $X2=8.465 $Y2=2.565
r194 45 47 33.1904 $w=2.48e-07 $l=7.2e-07 $layer=LI1_cond $X=8.59 $Y=1.48
+ $X2=8.59 $Y2=0.76
r195 44 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.075 $Y=2.395
+ $X2=7.99 $Y2=2.395
r196 43 68 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.295 $Y=2.395
+ $X2=8.38 $Y2=2.395
r197 43 44 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=8.295 $Y=2.395
+ $X2=8.075 $Y2=2.395
r198 41 45 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=8.465 $Y=1.565
+ $X2=8.59 $Y2=1.48
r199 41 42 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=8.465 $Y=1.565
+ $X2=8.075 $Y2=1.565
r200 40 67 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.99 $Y=2.31
+ $X2=7.99 $Y2=2.395
r201 39 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.99 $Y=1.65
+ $X2=8.075 $Y2=1.565
r202 39 40 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=7.99 $Y=1.65
+ $X2=7.99 $Y2=2.31
r203 37 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.905 $Y=2.395
+ $X2=7.99 $Y2=2.395
r204 37 38 93.2941 $w=1.68e-07 $l=1.43e-06 $layer=LI1_cond $X=7.905 $Y=2.395
+ $X2=6.475 $Y2=2.395
r205 36 38 8.2443 $w=5.49e-07 $l=1.77482e-07 $layer=LI1_cond $X=6.39 $Y=2.255
+ $X2=6.475 $Y2=2.395
r206 36 65 8.44444 $w=5.49e-07 $l=5.21248e-07 $layer=LI1_cond $X=6.39 $Y=2.255
+ $X2=6.01 $Y2=2.59
r207 35 62 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.39 $Y=1.26
+ $X2=6.39 $Y2=1.175
r208 35 36 64.9144 $w=1.68e-07 $l=9.95e-07 $layer=LI1_cond $X=6.39 $Y=1.26
+ $X2=6.39 $Y2=2.255
r209 31 62 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=5.985 $Y=1.175
+ $X2=6.39 $Y2=1.175
r210 31 33 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=5.985 $Y=1.09
+ $X2=5.985 $Y2=0.835
r211 29 65 10.0221 $w=5.49e-07 $l=3.22102e-07 $layer=LI1_cond $X=5.845 $Y=2.34
+ $X2=6.01 $Y2=2.59
r212 29 30 63.9358 $w=1.68e-07 $l=9.8e-07 $layer=LI1_cond $X=5.845 $Y=2.34
+ $X2=4.865 $Y2=2.34
r213 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.78 $Y=2.425
+ $X2=4.865 $Y2=2.34
r214 27 28 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=4.78 $Y=2.425
+ $X2=4.78 $Y2=2.905
r215 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.695 $Y=2.99
+ $X2=4.78 $Y2=2.905
r216 25 26 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=4.695 $Y=2.99
+ $X2=3.965 $Y2=2.99
r217 22 26 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.84 $Y=2.905
+ $X2=3.965 $Y2=2.99
r218 22 24 20.744 $w=2.48e-07 $l=4.5e-07 $layer=LI1_cond $X=3.84 $Y=2.905
+ $X2=3.84 $Y2=2.455
r219 21 59 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=3.84 $Y=2.415
+ $X2=3.84 $Y2=2.29
r220 21 24 1.84391 $w=2.48e-07 $l=4e-08 $layer=LI1_cond $X=3.84 $Y=2.415
+ $X2=3.84 $Y2=2.455
r221 6 53 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=8.825
+ $Y=2.54 $X2=8.97 $Y2=2.75
r222 5 65 300 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=2 $X=5.86
+ $Y=2.265 $X2=6.01 $Y2=2.42
r223 4 24 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=3.73
+ $Y=2.31 $X2=3.88 $Y2=2.455
r224 3 47 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=8.485
+ $Y=0.485 $X2=8.63 $Y2=0.76
r225 2 33 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=5.845
+ $Y=0.625 $X2=5.985 $Y2=0.835
r226 1 56 182 $w=1.7e-07 $l=2.96985e-07 $layer=licon1_NDIFF $count=1 $X=3.455
+ $Y=0.565 $X2=3.665 $Y2=0.775
.ends

.subckt PM_SKY130_FD_SC_LS__SEDFXBP_2%Q 1 2 7 8 9 10 11
r19 10 11 10.8465 $w=3.38e-07 $l=3.2e-07 $layer=LI1_cond $X=15.655 $Y=1.665
+ $X2=15.655 $Y2=1.985
r20 9 10 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=15.655 $Y=1.295
+ $X2=15.655 $Y2=1.665
r21 8 9 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=15.655 $Y=0.925
+ $X2=15.655 $Y2=1.295
r22 7 8 13.8971 $w=3.38e-07 $l=4.1e-07 $layer=LI1_cond $X=15.655 $Y=0.515
+ $X2=15.655 $Y2=0.925
r23 2 11 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=15.5
+ $Y=1.84 $X2=15.65 $Y2=1.985
r24 1 7 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=15.52
+ $Y=0.37 $X2=15.66 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__SEDFXBP_2%Q_N 1 2 7 8 9 10 11 12 13 28 32
c33 8 0 1.4807e-19 $X=16.932 $Y=1.805
r34 29 32 0.501062 $w=2.28e-07 $l=1e-08 $layer=LI1_cond $X=16.55 $Y=1.975
+ $X2=16.55 $Y2=1.985
r35 21 28 1.22229 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=16.52 $Y=0.96
+ $X2=16.52 $Y2=0.925
r36 12 13 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=16.55 $Y=2.405
+ $X2=16.55 $Y2=2.775
r37 11 29 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=16.56 $Y=1.89
+ $X2=16.55 $Y2=1.89
r38 11 12 17.938 $w=2.28e-07 $l=3.58e-07 $layer=LI1_cond $X=16.55 $Y=2.047
+ $X2=16.55 $Y2=2.405
r39 11 32 3.10659 $w=2.28e-07 $l=6.2e-08 $layer=LI1_cond $X=16.55 $Y=2.047
+ $X2=16.55 $Y2=1.985
r40 10 21 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=16.56 $Y=1.045
+ $X2=16.52 $Y2=1.045
r41 10 28 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=16.52 $Y=0.9
+ $X2=16.52 $Y2=0.925
r42 9 10 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=16.52 $Y=0.515
+ $X2=16.52 $Y2=0.9
r43 8 11 24.2695 $w=1.68e-07 $l=3.72e-07 $layer=LI1_cond $X=16.932 $Y=1.89
+ $X2=16.56 $Y2=1.89
r44 7 10 24.2695 $w=1.68e-07 $l=3.72e-07 $layer=LI1_cond $X=16.932 $Y=1.045
+ $X2=16.56 $Y2=1.045
r45 7 8 17.3624 $w=4.63e-07 $l=6.75e-07 $layer=LI1_cond $X=16.932 $Y=1.13
+ $X2=16.932 $Y2=1.805
r46 2 32 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=16.4
+ $Y=1.84 $X2=16.55 $Y2=1.985
r47 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=16.38
+ $Y=0.37 $X2=16.52 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__SEDFXBP_2%VGND 1 2 3 4 5 6 7 8 9 10 11 36 40 44 48
+ 52 56 60 62 63 68 70 74 76 80 82 84 87 88 90 91 93 94 96 105 109 118 122 134
+ 140 143 146 149 152 155 159 162 166
r220 165 166 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=17.04 $Y=0
+ $X2=17.04 $Y2=0
r221 162 163 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=16.08 $Y=0
+ $X2=16.08 $Y2=0
r222 160 163 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=15.12 $Y=0
+ $X2=16.08 $Y2=0
r223 159 160 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=15.12 $Y=0
+ $X2=15.12 $Y2=0
r224 156 160 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=14.16 $Y=0
+ $X2=15.12 $Y2=0
r225 155 156 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=14.16 $Y=0
+ $X2=14.16 $Y2=0
r226 152 153 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r227 149 150 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r228 146 147 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r229 143 144 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r230 140 141 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r231 138 166 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=16.56 $Y=0
+ $X2=17.04 $Y2=0
r232 138 163 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=16.56 $Y=0
+ $X2=16.08 $Y2=0
r233 137 138 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=16.56 $Y=0
+ $X2=16.56 $Y2=0
r234 135 162 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=16.175 $Y=0
+ $X2=16.09 $Y2=0
r235 135 137 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=16.175 $Y=0
+ $X2=16.56 $Y2=0
r236 134 165 4.03428 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=16.855 $Y=0
+ $X2=17.067 $Y2=0
r237 134 137 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=16.855 $Y=0
+ $X2=16.56 $Y2=0
r238 133 156 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=13.2 $Y=0
+ $X2=14.16 $Y2=0
r239 132 133 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=13.2 $Y=0
+ $X2=13.2 $Y2=0
r240 130 133 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=13.2 $Y2=0
r241 130 153 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=11.76 $Y2=0
r242 129 132 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=12.24 $Y=0
+ $X2=13.2 $Y2=0
r243 129 130 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r244 127 152 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.96 $Y=0
+ $X2=11.835 $Y2=0
r245 127 129 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=11.96 $Y=0
+ $X2=12.24 $Y2=0
r246 126 153 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=11.76 $Y2=0
r247 126 150 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=10.32 $Y2=0
r248 125 126 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.8 $Y=0
+ $X2=10.8 $Y2=0
r249 123 149 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.52 $Y=0
+ $X2=10.395 $Y2=0
r250 123 125 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=10.52 $Y=0
+ $X2=10.8 $Y2=0
r251 122 152 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.71 $Y=0
+ $X2=11.835 $Y2=0
r252 122 125 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=11.71 $Y=0
+ $X2=10.8 $Y2=0
r253 120 121 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r254 118 149 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.27 $Y=0
+ $X2=10.395 $Y2=0
r255 118 120 153.316 $w=1.68e-07 $l=2.35e-06 $layer=LI1_cond $X=10.27 $Y=0
+ $X2=7.92 $Y2=0
r256 117 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=7.92 $Y2=0
r257 117 147 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=6.48 $Y2=0
r258 116 117 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r259 114 146 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.745 $Y=0
+ $X2=6.58 $Y2=0
r260 114 116 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=6.745 $Y=0
+ $X2=7.44 $Y2=0
r261 113 147 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0
+ $X2=6.48 $Y2=0
r262 113 144 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0
+ $X2=5.04 $Y2=0
r263 112 113 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r264 110 143 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.29 $Y=0
+ $X2=5.125 $Y2=0
r265 110 112 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=5.29 $Y=0
+ $X2=5.52 $Y2=0
r266 109 146 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.415 $Y=0
+ $X2=6.58 $Y2=0
r267 109 112 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=6.415 $Y=0
+ $X2=5.52 $Y2=0
r268 108 144 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=5.04 $Y2=0
r269 107 108 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r270 105 143 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.96 $Y=0
+ $X2=5.125 $Y2=0
r271 105 107 151.358 $w=1.68e-07 $l=2.32e-06 $layer=LI1_cond $X=4.96 $Y=0
+ $X2=2.64 $Y2=0
r272 104 108 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=2.64 $Y2=0
r273 104 141 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=1.2 $Y2=0
r274 103 104 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r275 101 140 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.4 $Y=0
+ $X2=1.235 $Y2=0
r276 101 103 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=1.4 $Y=0 $X2=2.16
+ $Y2=0
r277 99 141 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r278 98 99 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r279 96 140 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.07 $Y=0
+ $X2=1.235 $Y2=0
r280 96 98 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.07 $Y=0 $X2=0.72
+ $Y2=0
r281 94 150 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=8.64 $Y=0
+ $X2=10.32 $Y2=0
r282 94 121 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=8.64 $Y=0
+ $X2=7.92 $Y2=0
r283 93 132 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=13.32 $Y=0
+ $X2=13.2 $Y2=0
r284 90 116 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=7.555 $Y=0
+ $X2=7.44 $Y2=0
r285 90 91 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.555 $Y=0 $X2=7.64
+ $Y2=0
r286 89 120 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=7.725 $Y=0
+ $X2=7.92 $Y2=0
r287 89 91 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.725 $Y=0 $X2=7.64
+ $Y2=0
r288 87 103 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=2.18 $Y=0 $X2=2.16
+ $Y2=0
r289 87 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.18 $Y=0 $X2=2.345
+ $Y2=0
r290 86 107 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=2.51 $Y=0 $X2=2.64
+ $Y2=0
r291 86 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.51 $Y=0 $X2=2.345
+ $Y2=0
r292 82 165 3.17794 $w=2.6e-07 $l=1.19143e-07 $layer=LI1_cond $X=16.985 $Y=0.085
+ $X2=17.067 $Y2=0
r293 82 84 23.9354 $w=2.58e-07 $l=5.4e-07 $layer=LI1_cond $X=16.985 $Y=0.085
+ $X2=16.985 $Y2=0.625
r294 78 162 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=16.09 $Y=0.085
+ $X2=16.09 $Y2=0
r295 78 80 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=16.09 $Y=0.085
+ $X2=16.09 $Y2=0.515
r296 77 159 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=15.315 $Y=0
+ $X2=15.19 $Y2=0
r297 76 162 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=16.005 $Y=0
+ $X2=16.09 $Y2=0
r298 76 77 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=16.005 $Y=0
+ $X2=15.315 $Y2=0
r299 72 159 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=15.19 $Y=0.085
+ $X2=15.19 $Y2=0
r300 72 74 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=15.19 $Y=0.085
+ $X2=15.19 $Y2=0.515
r301 71 155 3.47156 $w=4.27e-07 $l=3.17402e-07 $layer=LI1_cond $X=14.335 $Y=0
+ $X2=14.2 $Y2=0.257
r302 70 159 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=15.065 $Y=0
+ $X2=15.19 $Y2=0
r303 70 71 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=15.065 $Y=0
+ $X2=14.335 $Y2=0
r304 66 155 3.03886 $w=2.7e-07 $l=3.43e-07 $layer=LI1_cond $X=14.2 $Y=0.6
+ $X2=14.2 $Y2=0.257
r305 66 68 15.1525 $w=2.68e-07 $l=3.55e-07 $layer=LI1_cond $X=14.2 $Y=0.6
+ $X2=14.2 $Y2=0.955
r306 63 93 13.7992 $w=6.83e-07 $l=3.42e-07 $layer=LI1_cond $X=13.662 $Y=0.257
+ $X2=13.32 $Y2=0.257
r307 63 65 3.19536 $w=6.83e-07 $l=1.83e-07 $layer=LI1_cond $X=13.662 $Y=0.257
+ $X2=13.845 $Y2=0.257
r308 62 155 3.47156 $w=4.27e-07 $l=1.35e-07 $layer=LI1_cond $X=14.065 $Y=0.257
+ $X2=14.2 $Y2=0.257
r309 62 65 3.84142 $w=6.83e-07 $l=2.2e-07 $layer=LI1_cond $X=14.065 $Y=0.257
+ $X2=13.845 $Y2=0.257
r310 58 152 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=11.835 $Y=0.085
+ $X2=11.835 $Y2=0
r311 58 60 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=11.835 $Y=0.085
+ $X2=11.835 $Y2=0.515
r312 54 149 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=10.395 $Y=0.085
+ $X2=10.395 $Y2=0
r313 54 56 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=10.395 $Y=0.085
+ $X2=10.395 $Y2=0.515
r314 50 91 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.64 $Y=0.085
+ $X2=7.64 $Y2=0
r315 50 52 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=7.64 $Y=0.085
+ $X2=7.64 $Y2=0.515
r316 46 146 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.58 $Y=0.085
+ $X2=6.58 $Y2=0
r317 46 48 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=6.58 $Y=0.085
+ $X2=6.58 $Y2=0.495
r318 42 143 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.125 $Y=0.085
+ $X2=5.125 $Y2=0
r319 42 44 25.1442 $w=3.28e-07 $l=7.2e-07 $layer=LI1_cond $X=5.125 $Y=0.085
+ $X2=5.125 $Y2=0.805
r320 38 88 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.345 $Y=0.085
+ $X2=2.345 $Y2=0
r321 38 40 24.0965 $w=3.28e-07 $l=6.9e-07 $layer=LI1_cond $X=2.345 $Y=0.085
+ $X2=2.345 $Y2=0.775
r322 34 140 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.235 $Y=0.085
+ $X2=1.235 $Y2=0
r323 34 36 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=1.235 $Y=0.085
+ $X2=1.235 $Y2=0.58
r324 11 84 182 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=1 $X=16.81
+ $Y=0.37 $X2=16.95 $Y2=0.625
r325 10 80 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=15.95
+ $Y=0.37 $X2=16.09 $Y2=0.515
r326 9 74 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=15.085
+ $Y=0.37 $X2=15.23 $Y2=0.515
r327 8 155 182 $w=1.7e-07 $l=9.6478e-07 $layer=licon1_NDIFF $count=1 $X=13.345
+ $Y=0.37 $X2=14.24 $Y2=0.515
r328 8 68 182 $w=1.7e-07 $l=1.15091e-06 $layer=licon1_NDIFF $count=1 $X=13.345
+ $Y=0.37 $X2=14.24 $Y2=0.955
r329 8 65 91 $w=1.7e-07 $l=5.67891e-07 $layer=licon1_NDIFF $count=2 $X=13.345
+ $Y=0.37 $X2=13.845 $Y2=0.515
r330 7 60 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=11.65
+ $Y=0.37 $X2=11.795 $Y2=0.515
r331 6 56 182 $w=1.7e-07 $l=2.34521e-07 $layer=licon1_NDIFF $count=1 $X=10.215
+ $Y=0.485 $X2=10.435 $Y2=0.515
r332 5 52 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=7.495
+ $Y=0.37 $X2=7.64 $Y2=0.515
r333 4 48 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=6.435
+ $Y=0.37 $X2=6.58 $Y2=0.495
r334 3 44 182 $w=1.7e-07 $l=2.86182e-07 $layer=licon1_NDIFF $count=1 $X=4.915
+ $Y=0.625 $X2=5.125 $Y2=0.805
r335 2 40 182 $w=1.7e-07 $l=2.96985e-07 $layer=licon1_NDIFF $count=1 $X=2.135
+ $Y=0.565 $X2=2.345 $Y2=0.775
r336 1 36 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.095
+ $Y=0.37 $X2=1.235 $Y2=0.58
.ends

