* File: sky130_fd_sc_ls__or3_4.spice
* Created: Wed Sep  2 11:24:59 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__or3_4.pex.spice"
.subckt sky130_fd_sc_ls__or3_4  VNB VPB A B C VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* C	C
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1008 N_VGND_M1008_d N_C_M1008_g N_A_302_388#_M1008_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1332 AS=0.2109 PD=1.1 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75003.1 A=0.111 P=1.78 MULT=1
MM1012 N_A_302_388#_M1012_d N_B_M1012_g N_VGND_M1008_d VNB NSHORT L=0.15 W=0.74
+ AD=0.1258 AS=0.1332 PD=1.08 PS=1.1 NRD=9.72 NRS=1.62 M=1 R=4.93333 SA=75000.7
+ SB=75002.6 A=0.111 P=1.78 MULT=1
MM1004 N_VGND_M1004_d N_A_M1004_g N_A_302_388#_M1012_d VNB NSHORT L=0.15 W=0.74
+ AD=0.1295 AS=0.1258 PD=1.09 PS=1.08 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75001.2
+ SB=75002.1 A=0.111 P=1.78 MULT=1
MM1001 N_X_M1001_d N_A_302_388#_M1001_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.74
+ AD=0.10545 AS=0.1295 PD=1.025 PS=1.09 NRD=0.804 NRS=0 M=1 R=4.93333 SA=75001.7
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1007 N_X_M1001_d N_A_302_388#_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.74
+ AD=0.10545 AS=0.1258 PD=1.025 PS=1.08 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.1
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1009 N_X_M1009_d N_A_302_388#_M1009_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1258 PD=1.02 PS=1.08 NRD=0 NRS=9.72 M=1 R=4.93333 SA=75002.6
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1015 N_X_M1009_d N_A_302_388#_M1015_g N_VGND_M1015_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75003.1
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1002 N_A_116_388#_M1002_d N_A_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.295 PD=1.3 PS=2.59 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75000.2
+ SB=75004.5 A=0.15 P=2.3 MULT=1
MM1000 N_A_116_388#_M1002_d N_B_M1000_g N_A_206_388#_M1000_s VPB PHIGHVT L=0.15
+ W=1 AD=0.15 AS=0.165 PD=1.3 PS=1.33 NRD=1.9503 NRS=4.9053 M=1 R=6.66667
+ SA=75000.7 SB=75004 A=0.15 P=2.3 MULT=1
MM1013 N_A_302_388#_M1013_d N_C_M1013_g N_A_206_388#_M1000_s VPB PHIGHVT L=0.15
+ W=1 AD=0.15 AS=0.165 PD=1.3 PS=1.33 NRD=1.9503 NRS=4.9053 M=1 R=6.66667
+ SA=75001.1 SB=75003.6 A=0.15 P=2.3 MULT=1
MM1016 N_A_302_388#_M1013_d N_C_M1016_g N_A_206_388#_M1016_s VPB PHIGHVT L=0.15
+ W=1 AD=0.15 AS=0.1775 PD=1.3 PS=1.355 NRD=1.9503 NRS=6.8753 M=1 R=6.66667
+ SA=75001.6 SB=75003.1 A=0.15 P=2.3 MULT=1
MM1003 N_A_116_388#_M1003_d N_B_M1003_g N_A_206_388#_M1016_s VPB PHIGHVT L=0.15
+ W=1 AD=0.175 AS=0.1775 PD=1.35 PS=1.355 NRD=11.8003 NRS=7.8603 M=1 R=6.66667
+ SA=75002.1 SB=75002.6 A=0.15 P=2.3 MULT=1
MM1006 N_A_116_388#_M1003_d N_A_M1006_g N_VPWR_M1006_s VPB PHIGHVT L=0.15 W=1
+ AD=0.175 AS=0.196887 PD=1.35 PS=1.41981 NRD=1.9503 NRS=18.715 M=1 R=6.66667
+ SA=75002.6 SB=75002.1 A=0.15 P=2.3 MULT=1
MM1005 N_X_M1005_d N_A_302_388#_M1005_g N_VPWR_M1006_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.220513 PD=1.42 PS=1.59019 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.8 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1010 N_X_M1005_d N_A_302_388#_M1010_g N_VPWR_M1010_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75003.3 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1011 N_X_M1011_d N_A_302_388#_M1011_g N_VPWR_M1010_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75003.7 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1014 N_X_M1011_d N_A_302_388#_M1014_g N_VPWR_M1014_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75004.2 SB=75000.2 A=0.168 P=2.54 MULT=1
DX17_noxref VNB VPB NWDIODE A=10.5276 P=15.04
*
.include "sky130_fd_sc_ls__or3_4.pxi.spice"
*
.ends
*
*
