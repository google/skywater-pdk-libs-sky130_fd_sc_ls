* File: sky130_fd_sc_ls__o211ai_2.pxi.spice
* Created: Fri Aug 28 13:43:52 2020
* 
x_PM_SKY130_FD_SC_LS__O211AI_2%C1 N_C1_M1002_g N_C1_c_88_n N_C1_M1014_g
+ N_C1_M1003_g N_C1_c_89_n N_C1_M1015_g C1 N_C1_c_86_n N_C1_c_87_n
+ PM_SKY130_FD_SC_LS__O211AI_2%C1
x_PM_SKY130_FD_SC_LS__O211AI_2%B1 N_B1_c_135_n N_B1_M1005_g N_B1_M1000_g
+ N_B1_c_136_n N_B1_M1008_g N_B1_M1013_g B1 B1 N_B1_c_133_n N_B1_c_134_n
+ PM_SKY130_FD_SC_LS__O211AI_2%B1
x_PM_SKY130_FD_SC_LS__O211AI_2%A2 N_A2_c_188_n N_A2_M1011_g N_A2_M1004_g
+ N_A2_c_189_n N_A2_M1012_g N_A2_M1009_g A2 A2 N_A2_c_185_n N_A2_c_186_n
+ N_A2_c_187_n PM_SKY130_FD_SC_LS__O211AI_2%A2
x_PM_SKY130_FD_SC_LS__O211AI_2%A1 N_A1_c_245_n N_A1_M1001_g N_A1_M1006_g
+ N_A1_M1010_g N_A1_c_246_n N_A1_M1007_g A1 N_A1_c_243_n N_A1_c_244_n
+ PM_SKY130_FD_SC_LS__O211AI_2%A1
x_PM_SKY130_FD_SC_LS__O211AI_2%VPWR N_VPWR_M1014_s N_VPWR_M1015_s N_VPWR_M1008_s
+ N_VPWR_M1001_d N_VPWR_c_290_n N_VPWR_c_291_n N_VPWR_c_292_n N_VPWR_c_293_n
+ N_VPWR_c_294_n N_VPWR_c_295_n VPWR N_VPWR_c_296_n N_VPWR_c_297_n
+ N_VPWR_c_298_n N_VPWR_c_289_n N_VPWR_c_300_n N_VPWR_c_301_n N_VPWR_c_302_n
+ PM_SKY130_FD_SC_LS__O211AI_2%VPWR
x_PM_SKY130_FD_SC_LS__O211AI_2%Y N_Y_M1002_d N_Y_M1014_d N_Y_M1005_d N_Y_M1011_d
+ N_Y_c_360_n N_Y_c_354_n N_Y_c_368_n N_Y_c_357_n N_Y_c_358_n N_Y_c_355_n
+ N_Y_c_373_n N_Y_c_386_n N_Y_c_394_n Y Y PM_SKY130_FD_SC_LS__O211AI_2%Y
x_PM_SKY130_FD_SC_LS__O211AI_2%A_505_368# N_A_505_368#_M1011_s
+ N_A_505_368#_M1012_s N_A_505_368#_M1007_s N_A_505_368#_c_423_n
+ N_A_505_368#_c_424_n N_A_505_368#_c_425_n N_A_505_368#_c_426_n
+ N_A_505_368#_c_433_n N_A_505_368#_c_427_n N_A_505_368#_c_428_n
+ N_A_505_368#_c_429_n PM_SKY130_FD_SC_LS__O211AI_2%A_505_368#
x_PM_SKY130_FD_SC_LS__O211AI_2%A_30_84# N_A_30_84#_M1002_s N_A_30_84#_M1003_s
+ N_A_30_84#_M1013_s N_A_30_84#_c_467_n N_A_30_84#_c_468_n N_A_30_84#_c_469_n
+ N_A_30_84#_c_470_n N_A_30_84#_c_471_n PM_SKY130_FD_SC_LS__O211AI_2%A_30_84#
x_PM_SKY130_FD_SC_LS__O211AI_2%A_303_84# N_A_303_84#_M1000_d N_A_303_84#_M1004_s
+ N_A_303_84#_M1006_d N_A_303_84#_c_505_n N_A_303_84#_c_506_n
+ N_A_303_84#_c_507_n N_A_303_84#_c_508_n N_A_303_84#_c_509_n
+ N_A_303_84#_c_510_n PM_SKY130_FD_SC_LS__O211AI_2%A_303_84#
x_PM_SKY130_FD_SC_LS__O211AI_2%VGND N_VGND_M1004_d N_VGND_M1009_d N_VGND_M1010_s
+ N_VGND_c_552_n N_VGND_c_553_n N_VGND_c_554_n N_VGND_c_555_n VGND
+ N_VGND_c_556_n N_VGND_c_557_n N_VGND_c_558_n N_VGND_c_559_n N_VGND_c_560_n
+ N_VGND_c_561_n PM_SKY130_FD_SC_LS__O211AI_2%VGND
cc_1 VNB N_C1_M1002_g 0.0263047f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.79
cc_2 VNB N_C1_M1003_g 0.0196764f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=0.79
cc_3 VNB N_C1_c_86_n 0.0165723f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.515
cc_4 VNB N_C1_c_87_n 0.0622332f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=1.557
cc_5 VNB N_B1_M1000_g 0.0212084f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=2.4
cc_6 VNB N_B1_M1013_g 0.0270227f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=2.4
cc_7 VNB N_B1_c_133_n 0.00829772f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=1.557
cc_8 VNB N_B1_c_134_n 0.0363355f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.515
cc_9 VNB N_A2_M1004_g 0.0288139f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=2.4
cc_10 VNB N_A2_M1009_g 0.0215493f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=2.4
cc_11 VNB A2 0.00397139f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A2_c_185_n 0.0383468f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.515
cc_13 VNB N_A2_c_186_n 0.0397412f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A2_c_187_n 0.00344733f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A1_M1006_g 0.0211184f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=2.4
cc_16 VNB N_A1_M1010_g 0.0256402f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=0.79
cc_17 VNB A1 0.0263416f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.557
cc_18 VNB N_A1_c_243_n 0.084182f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.665
cc_19 VNB N_A1_c_244_n 0.00232983f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_VPWR_c_289_n 0.203486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_Y_c_354_n 0.00148201f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.515
cc_22 VNB N_Y_c_355_n 0.00410134f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_30_84#_c_467_n 0.0296889f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=1.765
cc_24 VNB N_A_30_84#_c_468_n 0.00482743f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=2.4
cc_25 VNB N_A_30_84#_c_469_n 0.00951014f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_26 VNB N_A_30_84#_c_470_n 0.0119635f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.557
cc_27 VNB N_A_30_84#_c_471_n 0.00572319f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=1.557
cc_28 VNB N_A_303_84#_c_505_n 0.0174175f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=0.79
cc_29 VNB N_A_303_84#_c_506_n 0.00178908f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=2.4
cc_30 VNB N_A_303_84#_c_507_n 0.00814736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_303_84#_c_508_n 0.00229554f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.557
cc_32 VNB N_A_303_84#_c_509_n 0.00243322f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_303_84#_c_510_n 0.00126893f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.665
cc_34 VNB N_VGND_c_552_n 0.0103499f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=1.765
cc_35 VNB N_VGND_c_553_n 0.00257504f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_554_n 0.0125081f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.515
cc_37 VNB N_VGND_c_555_n 0.0342758f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.557
cc_38 VNB N_VGND_c_556_n 0.0629405f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.515
cc_39 VNB N_VGND_c_557_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_558_n 0.016335f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_559_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_560_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_561_n 0.289293f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VPB N_C1_c_88_n 0.0179926f $X=-0.19 $Y=1.66 $X2=0.535 $Y2=1.765
cc_45 VPB N_C1_c_89_n 0.0159125f $X=-0.19 $Y=1.66 $X2=0.985 $Y2=1.765
cc_46 VPB N_C1_c_86_n 0.0102315f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.515
cc_47 VPB N_C1_c_87_n 0.0209876f $X=-0.19 $Y=1.66 $X2=0.94 $Y2=1.557
cc_48 VPB N_B1_c_135_n 0.0158124f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.35
cc_49 VPB N_B1_c_136_n 0.0179811f $X=-0.19 $Y=1.66 $X2=0.94 $Y2=1.35
cc_50 VPB N_B1_c_133_n 0.00856079f $X=-0.19 $Y=1.66 $X2=0.985 $Y2=1.557
cc_51 VPB N_B1_c_134_n 0.0217863f $X=-0.19 $Y=1.66 $X2=0.337 $Y2=1.515
cc_52 VPB N_A2_c_188_n 0.0184685f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.35
cc_53 VPB N_A2_c_189_n 0.0149065f $X=-0.19 $Y=1.66 $X2=0.94 $Y2=1.35
cc_54 VPB A2 0.00342544f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_A2_c_186_n 0.014191f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_A2_c_187_n 0.00510321f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_A1_c_245_n 0.0155495f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.35
cc_58 VPB N_A1_c_246_n 0.0210231f $X=-0.19 $Y=1.66 $X2=0.985 $Y2=1.765
cc_59 VPB N_A1_c_243_n 0.0164986f $X=-0.19 $Y=1.66 $X2=0.337 $Y2=1.665
cc_60 VPB N_VPWR_c_290_n 0.0116091f $X=-0.19 $Y=1.66 $X2=0.985 $Y2=2.4
cc_61 VPB N_VPWR_c_291_n 0.049587f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_62 VPB N_VPWR_c_292_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.515
cc_63 VPB N_VPWR_c_293_n 0.00799266f $X=-0.19 $Y=1.66 $X2=0.985 $Y2=1.557
cc_64 VPB N_VPWR_c_294_n 0.0149773f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_295_n 0.00651803f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_296_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_297_n 0.0389676f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_298_n 0.0191515f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_289_n 0.083841f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_300_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_301_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_302_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_Y_c_354_n 0.00251262f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.515
cc_74 VPB N_Y_c_357_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0.985 $Y2=1.557
cc_75 VPB N_Y_c_358_n 0.0167585f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB Y 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_A_505_368#_c_423_n 0.0055788f $X=-0.19 $Y=1.66 $X2=0.985 $Y2=1.765
cc_78 VPB N_A_505_368#_c_424_n 0.00523584f $X=-0.19 $Y=1.66 $X2=0.985 $Y2=2.4
cc_79 VPB N_A_505_368#_c_425_n 0.00384138f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_80 VPB N_A_505_368#_c_426_n 0.00318541f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_A_505_368#_c_427_n 0.00279022f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.557
cc_82 VPB N_A_505_368#_c_428_n 0.00907732f $X=-0.19 $Y=1.66 $X2=0.94 $Y2=1.557
cc_83 VPB N_A_505_368#_c_429_n 0.0403323f $X=-0.19 $Y=1.66 $X2=0.337 $Y2=1.515
cc_84 N_C1_c_89_n N_B1_c_135_n 0.0242681f $X=0.985 $Y=1.765 $X2=-0.19 $Y2=-0.245
cc_85 N_C1_M1003_g N_B1_M1000_g 0.0214079f $X=0.94 $Y=0.79 $X2=0 $Y2=0
cc_86 N_C1_c_87_n N_B1_c_133_n 0.00441801f $X=0.94 $Y=1.557 $X2=0 $Y2=0
cc_87 N_C1_c_87_n N_B1_c_134_n 0.0189721f $X=0.94 $Y=1.557 $X2=0 $Y2=0
cc_88 N_C1_c_88_n N_VPWR_c_291_n 0.00831454f $X=0.535 $Y=1.765 $X2=0 $Y2=0
cc_89 N_C1_c_86_n N_VPWR_c_291_n 0.0220584f $X=0.385 $Y=1.515 $X2=0 $Y2=0
cc_90 N_C1_c_87_n N_VPWR_c_291_n 0.00107017f $X=0.94 $Y=1.557 $X2=0 $Y2=0
cc_91 N_C1_c_88_n N_VPWR_c_292_n 0.00445602f $X=0.535 $Y=1.765 $X2=0 $Y2=0
cc_92 N_C1_c_89_n N_VPWR_c_292_n 0.00445602f $X=0.985 $Y=1.765 $X2=0 $Y2=0
cc_93 N_C1_c_89_n N_VPWR_c_293_n 0.00486623f $X=0.985 $Y=1.765 $X2=0 $Y2=0
cc_94 N_C1_c_88_n N_VPWR_c_289_n 0.00861179f $X=0.535 $Y=1.765 $X2=0 $Y2=0
cc_95 N_C1_c_89_n N_VPWR_c_289_n 0.00857673f $X=0.985 $Y=1.765 $X2=0 $Y2=0
cc_96 N_C1_M1002_g N_Y_c_360_n 0.00489796f $X=0.51 $Y=0.79 $X2=0 $Y2=0
cc_97 N_C1_M1003_g N_Y_c_360_n 0.00460661f $X=0.94 $Y=0.79 $X2=0 $Y2=0
cc_98 N_C1_M1002_g N_Y_c_354_n 0.002587f $X=0.51 $Y=0.79 $X2=0 $Y2=0
cc_99 N_C1_c_88_n N_Y_c_354_n 0.00279375f $X=0.535 $Y=1.765 $X2=0 $Y2=0
cc_100 N_C1_M1003_g N_Y_c_354_n 0.00463156f $X=0.94 $Y=0.79 $X2=0 $Y2=0
cc_101 N_C1_c_89_n N_Y_c_354_n 0.00201369f $X=0.985 $Y=1.765 $X2=0 $Y2=0
cc_102 N_C1_c_86_n N_Y_c_354_n 0.0318657f $X=0.385 $Y=1.515 $X2=0 $Y2=0
cc_103 N_C1_c_87_n N_Y_c_354_n 0.0185648f $X=0.94 $Y=1.557 $X2=0 $Y2=0
cc_104 N_C1_c_89_n N_Y_c_368_n 0.0159694f $X=0.985 $Y=1.765 $X2=0 $Y2=0
cc_105 N_C1_c_89_n N_Y_c_357_n 6.45594e-19 $X=0.985 $Y=1.765 $X2=0 $Y2=0
cc_106 N_C1_M1002_g N_Y_c_355_n 0.00325382f $X=0.51 $Y=0.79 $X2=0 $Y2=0
cc_107 N_C1_M1003_g N_Y_c_355_n 0.00190678f $X=0.94 $Y=0.79 $X2=0 $Y2=0
cc_108 N_C1_c_87_n N_Y_c_355_n 0.00191597f $X=0.94 $Y=1.557 $X2=0 $Y2=0
cc_109 N_C1_c_88_n N_Y_c_373_n 0.00256038f $X=0.535 $Y=1.765 $X2=0 $Y2=0
cc_110 N_C1_c_89_n N_Y_c_373_n 9.50925e-19 $X=0.985 $Y=1.765 $X2=0 $Y2=0
cc_111 N_C1_c_87_n N_Y_c_373_n 0.0028713f $X=0.94 $Y=1.557 $X2=0 $Y2=0
cc_112 N_C1_c_88_n Y 0.00960826f $X=0.535 $Y=1.765 $X2=0 $Y2=0
cc_113 N_C1_c_89_n Y 0.0103431f $X=0.985 $Y=1.765 $X2=0 $Y2=0
cc_114 N_C1_M1002_g N_A_30_84#_c_467_n 0.00159319f $X=0.51 $Y=0.79 $X2=0 $Y2=0
cc_115 N_C1_c_86_n N_A_30_84#_c_467_n 0.0217837f $X=0.385 $Y=1.515 $X2=0 $Y2=0
cc_116 N_C1_c_87_n N_A_30_84#_c_467_n 0.00125844f $X=0.94 $Y=1.557 $X2=0 $Y2=0
cc_117 N_C1_M1002_g N_A_30_84#_c_468_n 0.0141481f $X=0.51 $Y=0.79 $X2=0 $Y2=0
cc_118 N_C1_M1003_g N_A_30_84#_c_468_n 0.0134522f $X=0.94 $Y=0.79 $X2=0 $Y2=0
cc_119 N_C1_M1003_g N_A_30_84#_c_471_n 0.00240868f $X=0.94 $Y=0.79 $X2=0 $Y2=0
cc_120 N_C1_c_87_n N_A_30_84#_c_471_n 6.37393e-19 $X=0.94 $Y=1.557 $X2=0 $Y2=0
cc_121 N_C1_M1002_g N_VGND_c_556_n 8.76084e-19 $X=0.51 $Y=0.79 $X2=0 $Y2=0
cc_122 N_C1_M1003_g N_VGND_c_556_n 8.76084e-19 $X=0.94 $Y=0.79 $X2=0 $Y2=0
cc_123 N_B1_M1013_g N_A2_c_185_n 0.00856729f $X=1.94 $Y=0.79 $X2=0 $Y2=0
cc_124 N_B1_c_133_n N_A2_c_185_n 3.61578e-19 $X=1.85 $Y=1.515 $X2=0 $Y2=0
cc_125 N_B1_c_133_n N_A2_c_187_n 0.0184224f $X=1.85 $Y=1.515 $X2=0 $Y2=0
cc_126 N_B1_c_134_n N_A2_c_187_n 0.00112552f $X=1.885 $Y=1.557 $X2=0 $Y2=0
cc_127 N_B1_c_135_n N_VPWR_c_293_n 0.00486623f $X=1.435 $Y=1.765 $X2=0 $Y2=0
cc_128 N_B1_c_136_n N_VPWR_c_294_n 0.00714506f $X=1.885 $Y=1.765 $X2=0 $Y2=0
cc_129 N_B1_c_135_n N_VPWR_c_296_n 0.00445602f $X=1.435 $Y=1.765 $X2=0 $Y2=0
cc_130 N_B1_c_136_n N_VPWR_c_296_n 0.00445602f $X=1.885 $Y=1.765 $X2=0 $Y2=0
cc_131 N_B1_c_135_n N_VPWR_c_289_n 0.00857673f $X=1.435 $Y=1.765 $X2=0 $Y2=0
cc_132 N_B1_c_136_n N_VPWR_c_289_n 0.00862391f $X=1.885 $Y=1.765 $X2=0 $Y2=0
cc_133 N_B1_M1000_g N_Y_c_354_n 7.9877e-19 $X=1.44 $Y=0.79 $X2=0 $Y2=0
cc_134 N_B1_c_133_n N_Y_c_354_n 0.0317179f $X=1.85 $Y=1.515 $X2=0 $Y2=0
cc_135 N_B1_c_135_n N_Y_c_368_n 0.0119563f $X=1.435 $Y=1.765 $X2=0 $Y2=0
cc_136 N_B1_c_133_n N_Y_c_368_n 0.0284881f $X=1.85 $Y=1.515 $X2=0 $Y2=0
cc_137 N_B1_c_135_n N_Y_c_357_n 0.0103431f $X=1.435 $Y=1.765 $X2=0 $Y2=0
cc_138 N_B1_c_136_n N_Y_c_357_n 0.01498f $X=1.885 $Y=1.765 $X2=0 $Y2=0
cc_139 N_B1_c_136_n N_Y_c_358_n 0.0139279f $X=1.885 $Y=1.765 $X2=0 $Y2=0
cc_140 N_B1_c_133_n N_Y_c_358_n 0.0121995f $X=1.85 $Y=1.515 $X2=0 $Y2=0
cc_141 N_B1_c_135_n N_Y_c_386_n 4.27055e-19 $X=1.435 $Y=1.765 $X2=0 $Y2=0
cc_142 N_B1_c_136_n N_Y_c_386_n 4.27055e-19 $X=1.885 $Y=1.765 $X2=0 $Y2=0
cc_143 N_B1_c_133_n N_Y_c_386_n 0.0237598f $X=1.85 $Y=1.515 $X2=0 $Y2=0
cc_144 N_B1_c_134_n N_Y_c_386_n 0.00144657f $X=1.885 $Y=1.557 $X2=0 $Y2=0
cc_145 N_B1_c_135_n Y 6.45594e-19 $X=1.435 $Y=1.765 $X2=0 $Y2=0
cc_146 N_B1_M1000_g N_A_30_84#_c_470_n 0.0168204f $X=1.44 $Y=0.79 $X2=0 $Y2=0
cc_147 N_B1_M1013_g N_A_30_84#_c_470_n 0.0198009f $X=1.94 $Y=0.79 $X2=0 $Y2=0
cc_148 N_B1_c_133_n N_A_30_84#_c_470_n 0.00395247f $X=1.85 $Y=1.515 $X2=0 $Y2=0
cc_149 N_B1_M1000_g N_A_30_84#_c_471_n 0.0105901f $X=1.44 $Y=0.79 $X2=0 $Y2=0
cc_150 N_B1_M1013_g N_A_30_84#_c_471_n 6.5477e-19 $X=1.94 $Y=0.79 $X2=0 $Y2=0
cc_151 N_B1_c_133_n N_A_30_84#_c_471_n 0.0271148f $X=1.85 $Y=1.515 $X2=0 $Y2=0
cc_152 N_B1_c_134_n N_A_30_84#_c_471_n 5.01936e-19 $X=1.885 $Y=1.557 $X2=0 $Y2=0
cc_153 N_B1_M1013_g N_A_303_84#_c_505_n 0.00994167f $X=1.94 $Y=0.79 $X2=0 $Y2=0
cc_154 N_B1_c_133_n N_A_303_84#_c_505_n 0.00797813f $X=1.85 $Y=1.515 $X2=0 $Y2=0
cc_155 N_B1_M1000_g N_A_303_84#_c_509_n 0.0015116f $X=1.44 $Y=0.79 $X2=0 $Y2=0
cc_156 N_B1_M1013_g N_A_303_84#_c_509_n 0.00598046f $X=1.94 $Y=0.79 $X2=0 $Y2=0
cc_157 N_B1_c_133_n N_A_303_84#_c_509_n 0.0261926f $X=1.85 $Y=1.515 $X2=0 $Y2=0
cc_158 N_B1_c_134_n N_A_303_84#_c_509_n 0.0038569f $X=1.885 $Y=1.557 $X2=0 $Y2=0
cc_159 N_B1_M1013_g N_VGND_c_552_n 0.0023272f $X=1.94 $Y=0.79 $X2=0 $Y2=0
cc_160 N_B1_M1000_g N_VGND_c_556_n 8.94875e-19 $X=1.44 $Y=0.79 $X2=0 $Y2=0
cc_161 N_B1_M1013_g N_VGND_c_556_n 8.76084e-19 $X=1.94 $Y=0.79 $X2=0 $Y2=0
cc_162 N_A2_c_189_n N_A1_c_245_n 0.00967787f $X=3.345 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_163 N_A2_M1009_g N_A1_M1006_g 0.0299183f $X=3.37 $Y=0.74 $X2=0 $Y2=0
cc_164 N_A2_M1009_g N_A1_c_243_n 0.0196111f $X=3.37 $Y=0.74 $X2=0 $Y2=0
cc_165 A2 N_A1_c_243_n 4.12017e-19 $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_166 N_A2_c_186_n N_A1_c_243_n 0.00568023f $X=3.345 $Y=1.542 $X2=0 $Y2=0
cc_167 A2 N_A1_c_244_n 0.0210188f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_168 N_A2_c_186_n N_A1_c_244_n 4.12009e-19 $X=3.345 $Y=1.542 $X2=0 $Y2=0
cc_169 N_A2_c_188_n N_VPWR_c_294_n 8.40374e-19 $X=2.895 $Y=1.765 $X2=0 $Y2=0
cc_170 N_A2_c_188_n N_VPWR_c_297_n 0.00278271f $X=2.895 $Y=1.765 $X2=0 $Y2=0
cc_171 N_A2_c_189_n N_VPWR_c_297_n 0.00278271f $X=3.345 $Y=1.765 $X2=0 $Y2=0
cc_172 N_A2_c_188_n N_VPWR_c_289_n 0.00358624f $X=2.895 $Y=1.765 $X2=0 $Y2=0
cc_173 N_A2_c_189_n N_VPWR_c_289_n 0.00353907f $X=3.345 $Y=1.765 $X2=0 $Y2=0
cc_174 N_A2_c_188_n N_Y_c_358_n 0.0139279f $X=2.895 $Y=1.765 $X2=0 $Y2=0
cc_175 N_A2_c_185_n N_Y_c_358_n 0.00181184f $X=2.805 $Y=1.485 $X2=0 $Y2=0
cc_176 N_A2_c_187_n N_Y_c_358_n 0.0387567f $X=3.005 $Y=1.55 $X2=0 $Y2=0
cc_177 N_A2_c_188_n N_Y_c_394_n 0.0134092f $X=2.895 $Y=1.765 $X2=0 $Y2=0
cc_178 N_A2_c_189_n N_Y_c_394_n 0.00924457f $X=3.345 $Y=1.765 $X2=0 $Y2=0
cc_179 A2 N_Y_c_394_n 0.0201187f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_180 N_A2_c_186_n N_Y_c_394_n 0.00129651f $X=3.345 $Y=1.542 $X2=0 $Y2=0
cc_181 N_A2_c_187_n N_Y_c_394_n 0.0026794f $X=3.005 $Y=1.55 $X2=0 $Y2=0
cc_182 N_A2_c_188_n N_A_505_368#_c_424_n 0.0136535f $X=2.895 $Y=1.765 $X2=0
+ $Y2=0
cc_183 N_A2_c_189_n N_A_505_368#_c_424_n 0.012504f $X=3.345 $Y=1.765 $X2=0 $Y2=0
cc_184 N_A2_c_189_n N_A_505_368#_c_426_n 0.00378881f $X=3.345 $Y=1.765 $X2=0
+ $Y2=0
cc_185 N_A2_c_189_n N_A_505_368#_c_433_n 0.00584968f $X=3.345 $Y=1.765 $X2=0
+ $Y2=0
cc_186 N_A2_M1004_g N_A_30_84#_c_470_n 0.00137242f $X=2.94 $Y=0.74 $X2=0 $Y2=0
cc_187 N_A2_M1004_g N_A_303_84#_c_505_n 0.0147855f $X=2.94 $Y=0.74 $X2=0 $Y2=0
cc_188 A2 N_A_303_84#_c_505_n 0.00496209f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_189 N_A2_c_185_n N_A_303_84#_c_505_n 0.00981932f $X=2.805 $Y=1.485 $X2=0
+ $Y2=0
cc_190 N_A2_c_187_n N_A_303_84#_c_505_n 0.0433508f $X=3.005 $Y=1.55 $X2=0 $Y2=0
cc_191 N_A2_M1004_g N_A_303_84#_c_506_n 3.92313e-19 $X=2.94 $Y=0.74 $X2=0 $Y2=0
cc_192 N_A2_M1009_g N_A_303_84#_c_506_n 3.92313e-19 $X=3.37 $Y=0.74 $X2=0 $Y2=0
cc_193 N_A2_M1009_g N_A_303_84#_c_507_n 0.0127084f $X=3.37 $Y=0.74 $X2=0 $Y2=0
cc_194 A2 N_A_303_84#_c_507_n 0.0148851f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_195 A2 N_A_303_84#_c_510_n 0.0147323f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_196 N_A2_c_186_n N_A_303_84#_c_510_n 7.91474e-19 $X=3.345 $Y=1.542 $X2=0
+ $Y2=0
cc_197 N_A2_M1004_g N_VGND_c_552_n 0.0112914f $X=2.94 $Y=0.74 $X2=0 $Y2=0
cc_198 N_A2_M1009_g N_VGND_c_552_n 4.58208e-19 $X=3.37 $Y=0.74 $X2=0 $Y2=0
cc_199 N_A2_M1004_g N_VGND_c_553_n 4.58208e-19 $X=2.94 $Y=0.74 $X2=0 $Y2=0
cc_200 N_A2_M1009_g N_VGND_c_553_n 0.0096639f $X=3.37 $Y=0.74 $X2=0 $Y2=0
cc_201 N_A2_M1004_g N_VGND_c_557_n 0.00383152f $X=2.94 $Y=0.74 $X2=0 $Y2=0
cc_202 N_A2_M1009_g N_VGND_c_557_n 0.00383152f $X=3.37 $Y=0.74 $X2=0 $Y2=0
cc_203 N_A2_M1004_g N_VGND_c_561_n 0.0075754f $X=2.94 $Y=0.74 $X2=0 $Y2=0
cc_204 N_A2_M1009_g N_VGND_c_561_n 0.0075754f $X=3.37 $Y=0.74 $X2=0 $Y2=0
cc_205 N_A1_c_245_n N_VPWR_c_295_n 0.0128268f $X=3.795 $Y=1.765 $X2=0 $Y2=0
cc_206 N_A1_c_246_n N_VPWR_c_295_n 0.00756136f $X=4.295 $Y=1.765 $X2=0 $Y2=0
cc_207 N_A1_c_245_n N_VPWR_c_297_n 0.00413917f $X=3.795 $Y=1.765 $X2=0 $Y2=0
cc_208 N_A1_c_246_n N_VPWR_c_298_n 0.00445602f $X=4.295 $Y=1.765 $X2=0 $Y2=0
cc_209 N_A1_c_245_n N_VPWR_c_289_n 0.0081781f $X=3.795 $Y=1.765 $X2=0 $Y2=0
cc_210 N_A1_c_246_n N_VPWR_c_289_n 0.00860873f $X=4.295 $Y=1.765 $X2=0 $Y2=0
cc_211 N_A1_c_245_n N_A_505_368#_c_424_n 0.00125031f $X=3.795 $Y=1.765 $X2=0
+ $Y2=0
cc_212 N_A1_c_245_n N_A_505_368#_c_433_n 0.00585153f $X=3.795 $Y=1.765 $X2=0
+ $Y2=0
cc_213 N_A1_c_245_n N_A_505_368#_c_427_n 0.0131491f $X=3.795 $Y=1.765 $X2=0
+ $Y2=0
cc_214 N_A1_c_246_n N_A_505_368#_c_427_n 0.0122806f $X=4.295 $Y=1.765 $X2=0
+ $Y2=0
cc_215 N_A1_c_243_n N_A_505_368#_c_427_n 0.00967642f $X=4.295 $Y=1.532 $X2=0
+ $Y2=0
cc_216 N_A1_c_244_n N_A_505_368#_c_427_n 0.0492535f $X=4.365 $Y=1.415 $X2=0
+ $Y2=0
cc_217 N_A1_c_246_n N_A_505_368#_c_428_n 8.3017e-19 $X=4.295 $Y=1.765 $X2=0
+ $Y2=0
cc_218 N_A1_c_243_n N_A_505_368#_c_428_n 0.00268037f $X=4.295 $Y=1.532 $X2=0
+ $Y2=0
cc_219 N_A1_c_244_n N_A_505_368#_c_428_n 0.0296882f $X=4.365 $Y=1.415 $X2=0
+ $Y2=0
cc_220 N_A1_c_245_n N_A_505_368#_c_429_n 9.60989e-19 $X=3.795 $Y=1.765 $X2=0
+ $Y2=0
cc_221 N_A1_c_246_n N_A_505_368#_c_429_n 0.0125008f $X=4.295 $Y=1.765 $X2=0
+ $Y2=0
cc_222 N_A1_M1006_g N_A_303_84#_c_507_n 0.0128457f $X=3.805 $Y=0.74 $X2=0 $Y2=0
cc_223 N_A1_M1010_g N_A_303_84#_c_507_n 0.00127757f $X=4.28 $Y=0.74 $X2=0 $Y2=0
cc_224 N_A1_c_243_n N_A_303_84#_c_507_n 0.0046047f $X=4.295 $Y=1.532 $X2=0 $Y2=0
cc_225 N_A1_c_244_n N_A_303_84#_c_507_n 0.0371669f $X=4.365 $Y=1.415 $X2=0 $Y2=0
cc_226 N_A1_M1006_g N_A_303_84#_c_508_n 4.44262e-19 $X=3.805 $Y=0.74 $X2=0 $Y2=0
cc_227 N_A1_M1010_g N_A_303_84#_c_508_n 4.4892e-19 $X=4.28 $Y=0.74 $X2=0 $Y2=0
cc_228 N_A1_M1006_g N_VGND_c_553_n 0.00949565f $X=3.805 $Y=0.74 $X2=0 $Y2=0
cc_229 N_A1_M1010_g N_VGND_c_553_n 4.51649e-19 $X=4.28 $Y=0.74 $X2=0 $Y2=0
cc_230 N_A1_M1006_g N_VGND_c_555_n 4.93565e-19 $X=3.805 $Y=0.74 $X2=0 $Y2=0
cc_231 N_A1_M1010_g N_VGND_c_555_n 0.0124427f $X=4.28 $Y=0.74 $X2=0 $Y2=0
cc_232 A1 N_VGND_c_555_n 0.0263105f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_233 N_A1_c_243_n N_VGND_c_555_n 0.0017669f $X=4.295 $Y=1.532 $X2=0 $Y2=0
cc_234 N_A1_c_244_n N_VGND_c_555_n 0.00136555f $X=4.365 $Y=1.415 $X2=0 $Y2=0
cc_235 N_A1_M1006_g N_VGND_c_558_n 0.00398535f $X=3.805 $Y=0.74 $X2=0 $Y2=0
cc_236 N_A1_M1010_g N_VGND_c_558_n 0.00383152f $X=4.28 $Y=0.74 $X2=0 $Y2=0
cc_237 N_A1_M1006_g N_VGND_c_561_n 0.00787968f $X=3.805 $Y=0.74 $X2=0 $Y2=0
cc_238 N_A1_M1010_g N_VGND_c_561_n 0.00757973f $X=4.28 $Y=0.74 $X2=0 $Y2=0
cc_239 N_VPWR_M1015_s N_Y_c_368_n 0.00445471f $X=1.06 $Y=1.84 $X2=0 $Y2=0
cc_240 N_VPWR_c_293_n N_Y_c_368_n 0.0136682f $X=1.21 $Y=2.455 $X2=0 $Y2=0
cc_241 N_VPWR_c_293_n N_Y_c_357_n 0.0449718f $X=1.21 $Y=2.455 $X2=0 $Y2=0
cc_242 N_VPWR_c_294_n N_Y_c_357_n 0.0462948f $X=2.11 $Y=2.455 $X2=0 $Y2=0
cc_243 N_VPWR_c_296_n N_Y_c_357_n 0.014552f $X=2.025 $Y=3.33 $X2=0 $Y2=0
cc_244 N_VPWR_c_289_n N_Y_c_357_n 0.0119791f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_245 N_VPWR_M1008_s N_Y_c_358_n 0.0129281f $X=1.96 $Y=1.84 $X2=0 $Y2=0
cc_246 N_VPWR_c_294_n N_Y_c_358_n 0.0202359f $X=2.11 $Y=2.455 $X2=0 $Y2=0
cc_247 N_VPWR_c_291_n N_Y_c_373_n 0.0121024f $X=0.31 $Y=2.115 $X2=0 $Y2=0
cc_248 N_VPWR_c_291_n Y 0.0576605f $X=0.31 $Y=2.115 $X2=0 $Y2=0
cc_249 N_VPWR_c_292_n Y 0.014552f $X=1.125 $Y=3.33 $X2=0 $Y2=0
cc_250 N_VPWR_c_293_n Y 0.0449718f $X=1.21 $Y=2.455 $X2=0 $Y2=0
cc_251 N_VPWR_c_289_n Y 0.0119791f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_252 N_VPWR_c_294_n N_A_505_368#_c_423_n 0.0397233f $X=2.11 $Y=2.455 $X2=0
+ $Y2=0
cc_253 N_VPWR_c_295_n N_A_505_368#_c_424_n 0.0125885f $X=4.02 $Y=2.325 $X2=0
+ $Y2=0
cc_254 N_VPWR_c_297_n N_A_505_368#_c_424_n 0.0582805f $X=3.855 $Y=3.33 $X2=0
+ $Y2=0
cc_255 N_VPWR_c_289_n N_A_505_368#_c_424_n 0.0326824f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_256 N_VPWR_c_294_n N_A_505_368#_c_425_n 0.0119251f $X=2.11 $Y=2.455 $X2=0
+ $Y2=0
cc_257 N_VPWR_c_297_n N_A_505_368#_c_425_n 0.0179217f $X=3.855 $Y=3.33 $X2=0
+ $Y2=0
cc_258 N_VPWR_c_289_n N_A_505_368#_c_425_n 0.00971942f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_259 N_VPWR_c_295_n N_A_505_368#_c_433_n 0.0484948f $X=4.02 $Y=2.325 $X2=0
+ $Y2=0
cc_260 N_VPWR_M1001_d N_A_505_368#_c_427_n 0.00250873f $X=3.87 $Y=1.84 $X2=0
+ $Y2=0
cc_261 N_VPWR_c_295_n N_A_505_368#_c_427_n 0.0202249f $X=4.02 $Y=2.325 $X2=0
+ $Y2=0
cc_262 N_VPWR_c_295_n N_A_505_368#_c_429_n 0.0315588f $X=4.02 $Y=2.325 $X2=0
+ $Y2=0
cc_263 N_VPWR_c_298_n N_A_505_368#_c_429_n 0.0145938f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_264 N_VPWR_c_289_n N_A_505_368#_c_429_n 0.0120466f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_265 N_Y_c_358_n N_A_505_368#_M1011_s 0.00594057f $X=2.955 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_266 N_Y_c_358_n N_A_505_368#_c_423_n 0.0202359f $X=2.955 $Y=2.035 $X2=0 $Y2=0
cc_267 N_Y_c_394_n N_A_505_368#_c_423_n 0.0298377f $X=3.12 $Y=2.115 $X2=0 $Y2=0
cc_268 N_Y_M1011_d N_A_505_368#_c_424_n 0.00197722f $X=2.97 $Y=1.84 $X2=0 $Y2=0
cc_269 N_Y_c_394_n N_A_505_368#_c_424_n 0.0160777f $X=3.12 $Y=2.115 $X2=0 $Y2=0
cc_270 N_Y_c_394_n N_A_505_368#_c_426_n 0.00308048f $X=3.12 $Y=2.115 $X2=0 $Y2=0
cc_271 N_Y_c_394_n N_A_505_368#_c_433_n 0.0489989f $X=3.12 $Y=2.115 $X2=0 $Y2=0
cc_272 N_Y_c_360_n N_A_30_84#_c_467_n 0.0216593f $X=0.725 $Y=0.68 $X2=0 $Y2=0
cc_273 N_Y_M1002_d N_A_30_84#_c_468_n 0.00176461f $X=0.585 $Y=0.42 $X2=0 $Y2=0
cc_274 N_Y_c_360_n N_A_30_84#_c_468_n 0.0158928f $X=0.725 $Y=0.68 $X2=0 $Y2=0
cc_275 N_Y_c_360_n N_A_30_84#_c_471_n 0.017638f $X=0.725 $Y=0.68 $X2=0 $Y2=0
cc_276 N_A_505_368#_c_426_n N_A_303_84#_c_507_n 0.00549175f $X=3.57 $Y=1.99
+ $X2=0 $Y2=0
cc_277 N_A_505_368#_c_427_n N_A_303_84#_c_507_n 8.52231e-19 $X=4.355 $Y=1.905
+ $X2=0 $Y2=0
cc_278 N_A_30_84#_c_470_n N_A_303_84#_M1000_d 0.00244396f $X=2.16 $Y=0.565
+ $X2=-0.19 $Y2=-0.245
cc_279 N_A_30_84#_M1013_s N_A_303_84#_c_505_n 0.0131383f $X=2.015 $Y=0.42 $X2=0
+ $Y2=0
cc_280 N_A_30_84#_c_470_n N_A_303_84#_c_505_n 0.0220402f $X=2.16 $Y=0.565 $X2=0
+ $Y2=0
cc_281 N_A_30_84#_c_470_n N_A_303_84#_c_509_n 0.0210984f $X=2.16 $Y=0.565 $X2=0
+ $Y2=0
cc_282 N_A_30_84#_c_471_n N_A_303_84#_c_509_n 0.0112335f $X=1.225 $Y=0.565 $X2=0
+ $Y2=0
cc_283 N_A_30_84#_c_470_n N_VGND_c_552_n 0.0338381f $X=2.16 $Y=0.565 $X2=0 $Y2=0
cc_284 N_A_30_84#_c_468_n N_VGND_c_556_n 0.0437462f $X=1.06 $Y=0.34 $X2=0 $Y2=0
cc_285 N_A_30_84#_c_469_n N_VGND_c_556_n 0.0179217f $X=0.38 $Y=0.34 $X2=0 $Y2=0
cc_286 N_A_30_84#_c_470_n N_VGND_c_556_n 0.065133f $X=2.16 $Y=0.565 $X2=0 $Y2=0
cc_287 N_A_30_84#_c_471_n N_VGND_c_556_n 0.0236566f $X=1.225 $Y=0.565 $X2=0
+ $Y2=0
cc_288 N_A_30_84#_c_468_n N_VGND_c_561_n 0.0255585f $X=1.06 $Y=0.34 $X2=0 $Y2=0
cc_289 N_A_30_84#_c_469_n N_VGND_c_561_n 0.00971942f $X=0.38 $Y=0.34 $X2=0 $Y2=0
cc_290 N_A_30_84#_c_470_n N_VGND_c_561_n 0.0361835f $X=2.16 $Y=0.565 $X2=0 $Y2=0
cc_291 N_A_30_84#_c_471_n N_VGND_c_561_n 0.0128296f $X=1.225 $Y=0.565 $X2=0
+ $Y2=0
cc_292 N_A_303_84#_c_505_n N_VGND_M1004_d 0.00326148f $X=3.07 $Y=1.065 $X2=-0.19
+ $Y2=-0.245
cc_293 N_A_303_84#_c_507_n N_VGND_M1009_d 0.00188382f $X=3.935 $Y=1.065 $X2=0
+ $Y2=0
cc_294 N_A_303_84#_c_505_n N_VGND_c_552_n 0.0205937f $X=3.07 $Y=1.065 $X2=0
+ $Y2=0
cc_295 N_A_303_84#_c_506_n N_VGND_c_552_n 0.016636f $X=3.155 $Y=0.515 $X2=0
+ $Y2=0
cc_296 N_A_303_84#_c_506_n N_VGND_c_553_n 0.016636f $X=3.155 $Y=0.515 $X2=0
+ $Y2=0
cc_297 N_A_303_84#_c_507_n N_VGND_c_553_n 0.0160414f $X=3.935 $Y=1.065 $X2=0
+ $Y2=0
cc_298 N_A_303_84#_c_508_n N_VGND_c_553_n 0.0163061f $X=4.02 $Y=0.515 $X2=0
+ $Y2=0
cc_299 N_A_303_84#_c_508_n N_VGND_c_555_n 0.0246508f $X=4.02 $Y=0.515 $X2=0
+ $Y2=0
cc_300 N_A_303_84#_c_506_n N_VGND_c_557_n 0.00749631f $X=3.155 $Y=0.515 $X2=0
+ $Y2=0
cc_301 N_A_303_84#_c_508_n N_VGND_c_558_n 0.00995046f $X=4.02 $Y=0.515 $X2=0
+ $Y2=0
cc_302 N_A_303_84#_c_506_n N_VGND_c_561_n 0.0062048f $X=3.155 $Y=0.515 $X2=0
+ $Y2=0
cc_303 N_A_303_84#_c_508_n N_VGND_c_561_n 0.00823613f $X=4.02 $Y=0.515 $X2=0
+ $Y2=0
