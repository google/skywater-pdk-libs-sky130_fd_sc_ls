# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_ls__a221oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_ls__a221oi_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.56000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445000 1.430000 6.115000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.430000 4.265000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.365000 1.430000 8.095000 1.780000 ;
        RECT 6.730000 1.350000 8.095000 1.430000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.285000 1.350000 9.955000 1.780000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.525000 1.350000 1.875000 1.780000 ;
    END
  END C1
  PIN VNB
    PORT
      LAYER pwell ;
        RECT 0.000000 0.000000 10.560000 0.245000 ;
    END
  END VNB
  PIN VPB
    PORT
      LAYER nwell ;
        RECT -0.190000 1.660000 10.750000 3.520000 ;
    END
  END VPB
  PIN Y
    ANTENNADIFFAREA  2.380200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 0.350000 0.495000 1.010000 ;
        RECT 0.105000 1.010000 2.295000 1.090000 ;
        RECT 0.105000 1.090000 8.210000 1.180000 ;
        RECT 0.105000 1.180000 0.355000 2.905000 ;
        RECT 0.105000 2.905000 2.235000 3.075000 ;
        RECT 1.005000 2.290000 1.335000 2.905000 ;
        RECT 1.185000 0.350000 1.355000 1.010000 ;
        RECT 1.905000 2.290000 2.235000 2.905000 ;
        RECT 2.045000 0.350000 2.295000 1.010000 ;
        RECT 2.045000 1.180000 6.530000 1.260000 ;
        RECT 4.850000 0.640000 5.040000 1.090000 ;
        RECT 5.710000 0.640000 5.900000 1.090000 ;
        RECT 6.360000 0.850000 8.210000 1.090000 ;
        RECT 7.915000 0.770000 8.210000 0.850000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.560000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 10.560000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 10.560000 0.085000 ;
      RECT  0.000000  3.245000 10.560000 3.415000 ;
      RECT  0.555000  1.950000  9.925000 2.120000 ;
      RECT  0.555000  2.120000  0.835000 2.735000 ;
      RECT  0.675000  0.085000  1.005000 0.840000 ;
      RECT  1.505000  2.120000  1.735000 2.735000 ;
      RECT  1.535000  0.085000  1.865000 0.840000 ;
      RECT  2.615000  2.290000  6.725000 2.460000 ;
      RECT  2.615000  2.460000  2.945000 2.980000 ;
      RECT  2.630000  0.350000  2.880000 0.750000 ;
      RECT  2.630000  0.750000  4.680000 0.920000 ;
      RECT  3.060000  0.085000  3.390000 0.580000 ;
      RECT  3.145000  2.630000  3.315000 3.245000 ;
      RECT  3.515000  2.460000  3.845000 2.980000 ;
      RECT  3.570000  0.350000  3.740000 0.750000 ;
      RECT  3.920000  0.085000  4.250000 0.580000 ;
      RECT  4.045000  2.630000  4.215000 3.245000 ;
      RECT  4.415000  2.460000  4.745000 2.980000 ;
      RECT  4.430000  0.300000  6.400000 0.470000 ;
      RECT  4.430000  0.470000  4.680000 0.750000 ;
      RECT  4.945000  2.630000  5.115000 3.245000 ;
      RECT  5.210000  0.470000  5.540000 0.920000 ;
      RECT  5.315000  2.460000  5.645000 2.980000 ;
      RECT  5.815000  2.630000  6.275000 3.245000 ;
      RECT  6.070000  0.470000  6.400000 0.680000 ;
      RECT  6.445000  2.460000  6.725000 2.905000 ;
      RECT  6.445000  2.905000 10.375000 3.075000 ;
      RECT  6.590000  0.350000  8.560000 0.600000 ;
      RECT  6.590000  0.600000  6.920000 0.680000 ;
      RECT  6.895000  2.120000  7.225000 2.735000 ;
      RECT  7.395000  2.290000  7.625000 2.905000 ;
      RECT  7.450000  0.600000  7.745000 0.680000 ;
      RECT  7.795000  2.120000  8.125000 2.735000 ;
      RECT  8.295000  2.290000  8.525000 2.905000 ;
      RECT  8.390000  0.600000  8.560000 1.010000 ;
      RECT  8.390000  1.010000 10.360000 1.180000 ;
      RECT  8.695000  2.120000  9.025000 2.735000 ;
      RECT  8.740000  0.085000  9.070000 0.840000 ;
      RECT  9.195000  2.290000  9.425000 2.905000 ;
      RECT  9.250000  0.350000  9.420000 1.010000 ;
      RECT  9.595000  2.120000  9.925000 2.735000 ;
      RECT  9.600000  0.085000  9.930000 0.840000 ;
      RECT 10.110000  0.350000 10.360000 1.010000 ;
      RECT 10.125000  1.820000 10.375000 2.905000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
  END
END sky130_fd_sc_ls__a221oi_4
END LIBRARY
