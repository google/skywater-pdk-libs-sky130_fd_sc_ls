* File: sky130_fd_sc_ls__sedfxbp_2.pxi.spice
* Created: Fri Aug 28 14:07:12 2020
* 
x_PM_SKY130_FD_SC_LS__SEDFXBP_2%D N_D_c_350_n N_D_c_351_n N_D_M1004_g
+ N_D_M1047_g D D N_D_c_347_n N_D_c_348_n N_D_c_349_n N_D_c_354_n
+ PM_SKY130_FD_SC_LS__SEDFXBP_2%D
x_PM_SKY130_FD_SC_LS__SEDFXBP_2%A_183_290# N_A_183_290#_M1028_s
+ N_A_183_290#_M1017_s N_A_183_290#_c_397_n N_A_183_290#_M1029_g
+ N_A_183_290#_M1024_g N_A_183_290#_c_398_n N_A_183_290#_c_390_n
+ N_A_183_290#_c_391_n N_A_183_290#_c_392_n N_A_183_290#_c_393_n
+ N_A_183_290#_c_400_n N_A_183_290#_c_401_n N_A_183_290#_c_394_n
+ N_A_183_290#_c_402_n N_A_183_290#_c_403_n N_A_183_290#_c_395_n
+ N_A_183_290#_c_396_n N_A_183_290#_c_406_n
+ PM_SKY130_FD_SC_LS__SEDFXBP_2%A_183_290#
x_PM_SKY130_FD_SC_LS__SEDFXBP_2%DE N_DE_M1042_g N_DE_c_503_n N_DE_c_504_n
+ N_DE_c_505_n N_DE_c_511_n N_DE_c_512_n N_DE_c_513_n N_DE_c_506_n N_DE_M1028_g
+ N_DE_c_514_n N_DE_M1017_g N_DE_c_515_n N_DE_c_516_n N_DE_M1044_g N_DE_c_507_n
+ N_DE_c_517_n DE N_DE_c_509_n N_DE_c_510_n PM_SKY130_FD_SC_LS__SEDFXBP_2%DE
x_PM_SKY130_FD_SC_LS__SEDFXBP_2%A_575_87# N_A_575_87#_M1014_d
+ N_A_575_87#_M1020_d N_A_575_87#_M1006_g N_A_575_87#_c_615_n
+ N_A_575_87#_c_616_n N_A_575_87#_M1018_g N_A_575_87#_c_598_n
+ N_A_575_87#_M1026_g N_A_575_87#_c_599_n N_A_575_87#_c_600_n
+ N_A_575_87#_c_617_n N_A_575_87#_M1022_g N_A_575_87#_c_601_n
+ N_A_575_87#_M1027_g N_A_575_87#_c_619_n N_A_575_87#_M1031_g
+ N_A_575_87#_M1041_g N_A_575_87#_c_620_n N_A_575_87#_M1038_g
+ N_A_575_87#_c_621_n N_A_575_87#_c_604_n N_A_575_87#_c_623_n
+ N_A_575_87#_c_605_n N_A_575_87#_c_606_n N_A_575_87#_c_727_p
+ N_A_575_87#_c_607_n N_A_575_87#_c_608_n N_A_575_87#_c_609_n
+ N_A_575_87#_c_610_n N_A_575_87#_c_633_n N_A_575_87#_c_611_n
+ N_A_575_87#_c_612_n N_A_575_87#_c_613_n N_A_575_87#_c_614_n
+ PM_SKY130_FD_SC_LS__SEDFXBP_2%A_575_87#
x_PM_SKY130_FD_SC_LS__SEDFXBP_2%A_661_87# N_A_661_87#_M1039_s
+ N_A_661_87#_M1045_s N_A_661_87#_c_887_n N_A_661_87#_M1010_g
+ N_A_661_87#_c_888_n N_A_661_87#_c_889_n N_A_661_87#_c_896_n
+ N_A_661_87#_M1000_g N_A_661_87#_c_890_n N_A_661_87#_c_897_n
+ N_A_661_87#_c_891_n N_A_661_87#_c_907_n N_A_661_87#_c_898_n
+ N_A_661_87#_c_892_n N_A_661_87#_c_899_n N_A_661_87#_c_893_n
+ N_A_661_87#_c_900_n N_A_661_87#_c_894_n N_A_661_87#_c_902_n
+ N_A_661_87#_c_903_n N_A_661_87#_c_895_n
+ PM_SKY130_FD_SC_LS__SEDFXBP_2%A_661_87#
x_PM_SKY130_FD_SC_LS__SEDFXBP_2%SCD N_SCD_c_998_n N_SCD_c_1003_n N_SCD_M1012_g
+ N_SCD_M1021_g SCD N_SCD_c_1001_n PM_SKY130_FD_SC_LS__SEDFXBP_2%SCD
x_PM_SKY130_FD_SC_LS__SEDFXBP_2%SCE N_SCE_c_1051_n N_SCE_M1033_g N_SCE_c_1052_n
+ N_SCE_c_1053_n N_SCE_c_1044_n N_SCE_c_1055_n N_SCE_M1045_g N_SCE_M1039_g
+ N_SCE_c_1046_n N_SCE_c_1047_n N_SCE_M1036_g SCE N_SCE_c_1049_n N_SCE_c_1050_n
+ PM_SKY130_FD_SC_LS__SEDFXBP_2%SCE
x_PM_SKY130_FD_SC_LS__SEDFXBP_2%CLK N_CLK_c_1127_n N_CLK_M1007_g N_CLK_c_1128_n
+ N_CLK_M1035_g CLK PM_SKY130_FD_SC_LS__SEDFXBP_2%CLK
x_PM_SKY130_FD_SC_LS__SEDFXBP_2%A_1586_74# N_A_1586_74#_M1003_d
+ N_A_1586_74#_M1001_d N_A_1586_74#_c_1187_n N_A_1586_74#_M1008_g
+ N_A_1586_74#_c_1163_n N_A_1586_74#_M1040_g N_A_1586_74#_M1011_g
+ N_A_1586_74#_c_1165_n N_A_1586_74#_c_1189_n N_A_1586_74#_M1025_g
+ N_A_1586_74#_c_1166_n N_A_1586_74#_c_1167_n N_A_1586_74#_c_1168_n
+ N_A_1586_74#_c_1190_n N_A_1586_74#_c_1169_n N_A_1586_74#_c_1170_n
+ N_A_1586_74#_c_1171_n N_A_1586_74#_c_1172_n N_A_1586_74#_c_1173_n
+ N_A_1586_74#_c_1273_p N_A_1586_74#_c_1174_n N_A_1586_74#_c_1175_n
+ N_A_1586_74#_c_1176_n N_A_1586_74#_c_1177_n N_A_1586_74#_c_1178_n
+ N_A_1586_74#_c_1179_n N_A_1586_74#_c_1180_n N_A_1586_74#_c_1181_n
+ N_A_1586_74#_c_1192_n N_A_1586_74#_c_1182_n N_A_1586_74#_c_1194_n
+ N_A_1586_74#_c_1183_n N_A_1586_74#_c_1311_p N_A_1586_74#_c_1184_n
+ N_A_1586_74#_c_1185_n N_A_1586_74#_c_1186_n
+ PM_SKY130_FD_SC_LS__SEDFXBP_2%A_1586_74#
x_PM_SKY130_FD_SC_LS__SEDFXBP_2%A_1374_368# N_A_1374_368#_M1035_d
+ N_A_1374_368#_M1007_d N_A_1374_368#_M1003_g N_A_1374_368#_c_1403_n
+ N_A_1374_368#_c_1417_n N_A_1374_368#_M1001_g N_A_1374_368#_c_1404_n
+ N_A_1374_368#_M1037_g N_A_1374_368#_c_1406_n N_A_1374_368#_c_1420_n
+ N_A_1374_368#_c_1421_n N_A_1374_368#_M1019_g N_A_1374_368#_c_1407_n
+ N_A_1374_368#_M1015_g N_A_1374_368#_M1013_g N_A_1374_368#_c_1409_n
+ N_A_1374_368#_c_1410_n N_A_1374_368#_c_1425_n N_A_1374_368#_c_1426_n
+ N_A_1374_368#_c_1427_n N_A_1374_368#_c_1411_n N_A_1374_368#_c_1412_n
+ N_A_1374_368#_c_1429_n N_A_1374_368#_c_1413_n N_A_1374_368#_c_1430_n
+ N_A_1374_368#_c_1414_n N_A_1374_368#_c_1415_n
+ PM_SKY130_FD_SC_LS__SEDFXBP_2%A_1374_368#
x_PM_SKY130_FD_SC_LS__SEDFXBP_2%A_2013_71# N_A_2013_71#_M1023_d
+ N_A_2013_71#_M1030_d N_A_2013_71#_M1034_g N_A_2013_71#_c_1593_n
+ N_A_2013_71#_c_1606_n N_A_2013_71#_M1002_g N_A_2013_71#_c_1594_n
+ N_A_2013_71#_c_1595_n N_A_2013_71#_c_1608_n N_A_2013_71#_M1046_g
+ N_A_2013_71#_c_1596_n N_A_2013_71#_M1009_g N_A_2013_71#_c_1597_n
+ N_A_2013_71#_c_1609_n N_A_2013_71#_c_1598_n N_A_2013_71#_c_1599_n
+ N_A_2013_71#_c_1600_n N_A_2013_71#_c_1601_n N_A_2013_71#_c_1602_n
+ N_A_2013_71#_c_1603_n N_A_2013_71#_c_1604_n
+ PM_SKY130_FD_SC_LS__SEDFXBP_2%A_2013_71#
x_PM_SKY130_FD_SC_LS__SEDFXBP_2%A_1784_97# N_A_1784_97#_M1037_d
+ N_A_1784_97#_M1008_d N_A_1784_97#_c_1706_n N_A_1784_97#_M1030_g
+ N_A_1784_97#_M1023_g N_A_1784_97#_c_1708_n N_A_1784_97#_c_1710_n
+ N_A_1784_97#_c_1711_n N_A_1784_97#_c_1712_n N_A_1784_97#_c_1713_n
+ N_A_1784_97#_c_1714_n PM_SKY130_FD_SC_LS__SEDFXBP_2%A_1784_97#
x_PM_SKY130_FD_SC_LS__SEDFXBP_2%A_2489_74# N_A_2489_74#_M1011_d
+ N_A_2489_74#_M1015_d N_A_2489_74#_c_1802_n N_A_2489_74#_M1020_g
+ N_A_2489_74#_M1014_g N_A_2489_74#_c_1792_n N_A_2489_74#_c_1793_n
+ N_A_2489_74#_c_1804_n N_A_2489_74#_M1005_g N_A_2489_74#_M1032_g
+ N_A_2489_74#_M1043_g N_A_2489_74#_c_1805_n N_A_2489_74#_M1016_g
+ N_A_2489_74#_c_1796_n N_A_2489_74#_c_1871_n N_A_2489_74#_c_1797_n
+ N_A_2489_74#_c_1798_n N_A_2489_74#_c_1807_n N_A_2489_74#_c_1808_n
+ N_A_2489_74#_c_1809_n N_A_2489_74#_c_1799_n N_A_2489_74#_c_1800_n
+ N_A_2489_74#_c_1801_n N_A_2489_74#_c_1811_n
+ PM_SKY130_FD_SC_LS__SEDFXBP_2%A_2489_74#
x_PM_SKY130_FD_SC_LS__SEDFXBP_2%A_32_74# N_A_32_74#_M1047_s N_A_32_74#_M1006_d
+ N_A_32_74#_M1004_s N_A_32_74#_M1018_d N_A_32_74#_c_1946_n N_A_32_74#_c_1952_n
+ N_A_32_74#_c_1953_n N_A_32_74#_c_1954_n N_A_32_74#_c_1955_n
+ N_A_32_74#_c_1956_n N_A_32_74#_c_1987_n N_A_32_74#_c_1957_n
+ N_A_32_74#_c_1958_n N_A_32_74#_c_1947_n N_A_32_74#_c_1948_n
+ N_A_32_74#_c_1949_n N_A_32_74#_c_1960_n N_A_32_74#_c_1950_n
+ N_A_32_74#_c_1961_n PM_SKY130_FD_SC_LS__SEDFXBP_2%A_32_74#
x_PM_SKY130_FD_SC_LS__SEDFXBP_2%VPWR N_VPWR_M1029_d N_VPWR_M1017_d
+ N_VPWR_M1045_d N_VPWR_M1007_s N_VPWR_M1001_s N_VPWR_M1002_d N_VPWR_M1046_s
+ N_VPWR_M1022_d N_VPWR_M1005_s N_VPWR_M1016_s N_VPWR_M1038_s N_VPWR_c_2067_n
+ N_VPWR_c_2068_n N_VPWR_c_2069_n N_VPWR_c_2070_n N_VPWR_c_2071_n
+ N_VPWR_c_2072_n N_VPWR_c_2073_n N_VPWR_c_2074_n N_VPWR_c_2075_n
+ N_VPWR_c_2076_n N_VPWR_c_2077_n N_VPWR_c_2078_n N_VPWR_c_2079_n
+ N_VPWR_c_2080_n N_VPWR_c_2081_n N_VPWR_c_2082_n VPWR N_VPWR_c_2083_n
+ N_VPWR_c_2084_n N_VPWR_c_2085_n N_VPWR_c_2086_n N_VPWR_c_2087_n
+ N_VPWR_c_2088_n N_VPWR_c_2089_n N_VPWR_c_2090_n N_VPWR_c_2091_n
+ N_VPWR_c_2092_n N_VPWR_c_2093_n N_VPWR_c_2094_n N_VPWR_c_2095_n
+ N_VPWR_c_2096_n N_VPWR_c_2097_n N_VPWR_c_2098_n N_VPWR_c_2099_n
+ N_VPWR_c_2066_n PM_SKY130_FD_SC_LS__SEDFXBP_2%VPWR
x_PM_SKY130_FD_SC_LS__SEDFXBP_2%A_691_113# N_A_691_113#_M1010_d
+ N_A_691_113#_M1036_d N_A_691_113#_M1037_s N_A_691_113#_M1033_d
+ N_A_691_113#_M1000_d N_A_691_113#_M1008_s N_A_691_113#_c_2274_n
+ N_A_691_113#_c_2339_n N_A_691_113#_c_2275_n N_A_691_113#_c_2286_n
+ N_A_691_113#_c_2302_n N_A_691_113#_c_2276_n N_A_691_113#_c_2277_n
+ N_A_691_113#_c_2266_n N_A_691_113#_c_2267_n N_A_691_113#_c_2279_n
+ N_A_691_113#_c_2280_n N_A_691_113#_c_2281_n N_A_691_113#_c_2268_n
+ N_A_691_113#_c_2269_n N_A_691_113#_c_2295_n N_A_691_113#_c_2270_n
+ N_A_691_113#_c_2282_n N_A_691_113#_c_2283_n N_A_691_113#_c_2271_n
+ N_A_691_113#_c_2272_n N_A_691_113#_c_2273_n N_A_691_113#_c_2438_n
+ N_A_691_113#_c_2375_n PM_SKY130_FD_SC_LS__SEDFXBP_2%A_691_113#
x_PM_SKY130_FD_SC_LS__SEDFXBP_2%Q N_Q_M1032_d N_Q_M1005_d Q Q Q Q Q
+ PM_SKY130_FD_SC_LS__SEDFXBP_2%Q
x_PM_SKY130_FD_SC_LS__SEDFXBP_2%Q_N N_Q_N_M1027_d N_Q_N_M1031_d N_Q_N_c_2476_n
+ N_Q_N_c_2477_n Q_N Q_N Q_N Q_N Q_N Q_N Q_N PM_SKY130_FD_SC_LS__SEDFXBP_2%Q_N
x_PM_SKY130_FD_SC_LS__SEDFXBP_2%VGND N_VGND_M1042_d N_VGND_M1028_d
+ N_VGND_M1039_d N_VGND_M1035_s N_VGND_M1003_s N_VGND_M1034_d N_VGND_M1009_s
+ N_VGND_M1026_d N_VGND_M1032_s N_VGND_M1043_s N_VGND_M1041_s N_VGND_c_2509_n
+ N_VGND_c_2510_n N_VGND_c_2511_n N_VGND_c_2512_n N_VGND_c_2513_n
+ N_VGND_c_2514_n N_VGND_c_2515_n N_VGND_c_2516_n N_VGND_c_2517_n
+ N_VGND_c_2518_n N_VGND_c_2519_n N_VGND_c_2520_n N_VGND_c_2521_n
+ N_VGND_c_2522_n N_VGND_c_2523_n N_VGND_c_2524_n N_VGND_c_2525_n
+ N_VGND_c_2526_n N_VGND_c_2527_n N_VGND_c_2528_n N_VGND_c_2529_n VGND
+ N_VGND_c_2530_n N_VGND_c_2531_n N_VGND_c_2532_n N_VGND_c_2533_n
+ N_VGND_c_2534_n N_VGND_c_2535_n N_VGND_c_2536_n N_VGND_c_2537_n
+ N_VGND_c_2538_n N_VGND_c_2539_n N_VGND_c_2540_n N_VGND_c_2541_n
+ N_VGND_c_2542_n N_VGND_c_2543_n N_VGND_c_2544_n
+ PM_SKY130_FD_SC_LS__SEDFXBP_2%VGND
cc_1 VNB N_D_M1047_g 0.0264128f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.58
cc_2 VNB N_D_c_347_n 0.0166671f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.145
cc_3 VNB N_D_c_348_n 0.0120671f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.145
cc_4 VNB N_D_c_349_n 0.0398527f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.825
cc_5 VNB N_A_183_290#_M1024_g 0.0449705f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_6 VNB N_A_183_290#_c_390_n 0.00295485f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.145
cc_7 VNB N_A_183_290#_c_391_n 0.0231869f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.145
cc_8 VNB N_A_183_290#_c_392_n 0.0073121f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.825
cc_9 VNB N_A_183_290#_c_393_n 4.59932e-19 $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.825
cc_10 VNB N_A_183_290#_c_394_n 0.00999719f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.295
cc_11 VNB N_A_183_290#_c_395_n 0.00268811f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_183_290#_c_396_n 0.0162115f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_DE_M1042_g 0.0299417f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=2.245
cc_14 VNB N_DE_c_503_n 0.0304597f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=2.64
cc_15 VNB N_DE_c_504_n 0.00725655f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.98
cc_16 VNB N_DE_c_505_n 0.0266857f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_DE_c_506_n 0.0179672f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_DE_c_507_n 0.00950241f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.295
cc_19 VNB DE 0.0038178f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.665
cc_20 VNB N_DE_c_509_n 0.0165295f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_DE_c_510_n 0.0196098f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_575_87#_M1006_g 0.0399729f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_575_87#_c_598_n 0.0170882f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.825
cc_24 VNB N_A_575_87#_c_599_n 0.0400986f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.145
cc_25 VNB N_A_575_87#_c_600_n 0.00716283f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.825
cc_26 VNB N_A_575_87#_c_601_n 0.0335071f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_575_87#_M1027_g 0.0215195f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.665
cc_28 VNB N_A_575_87#_M1041_g 0.023699f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_575_87#_c_604_n 5.3143e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_575_87#_c_605_n 0.00811762f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_575_87#_c_606_n 0.00364338f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_575_87#_c_607_n 9.39012e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_575_87#_c_608_n 0.00301273f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_575_87#_c_609_n 0.01027f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_575_87#_c_610_n 0.0465057f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_575_87#_c_611_n 2.4907e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_575_87#_c_612_n 0.00101108f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_575_87#_c_613_n 0.01914f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_575_87#_c_614_n 0.0506567f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_661_87#_c_887_n 0.0164494f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.58
cc_41 VNB N_A_661_87#_c_888_n 0.0374808f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.145
cc_42 VNB N_A_661_87#_c_889_n 0.00865069f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=0.98
cc_43 VNB N_A_661_87#_c_890_n 0.00880625f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.145
cc_44 VNB N_A_661_87#_c_891_n 0.00219983f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.145
cc_45 VNB N_A_661_87#_c_892_n 0.00716145f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.665
cc_46 VNB N_A_661_87#_c_893_n 0.0680445f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_661_87#_c_894_n 0.0346451f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_661_87#_c_895_n 0.032224f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_SCD_c_998_n 0.00875717f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=2.155
cc_50 VNB N_SCD_M1021_g 0.0175076f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.58
cc_51 VNB SCD 0.0142331f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.145
cc_52 VNB N_SCD_c_1001_n 0.0311734f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_53 VNB N_SCE_c_1044_n 0.00875383f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.58
cc_54 VNB N_SCE_M1039_g 0.0334855f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_SCE_c_1046_n 0.0681329f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.825
cc_56 VNB N_SCE_c_1047_n 0.012806f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.145
cc_57 VNB N_SCE_M1036_g 0.0359126f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.825
cc_58 VNB N_SCE_c_1049_n 0.027336f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_SCE_c_1050_n 0.0059654f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.295
cc_60 VNB N_CLK_c_1127_n 0.0450332f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.99
cc_61 VNB N_CLK_c_1128_n 0.0212689f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=2.64
cc_62 VNB CLK 0.00807833f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.58
cc_63 VNB N_A_1586_74#_c_1163_n 0.0185214f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.145
cc_64 VNB N_A_1586_74#_M1011_g 0.035432f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_1586_74#_c_1165_n 0.00537699f $X=-0.19 $Y=-0.245 $X2=0.54
+ $Y2=1.145
cc_66 VNB N_A_1586_74#_c_1166_n 0.00958186f $X=-0.19 $Y=-0.245 $X2=0.63
+ $Y2=1.145
cc_67 VNB N_A_1586_74#_c_1167_n 0.0189124f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.295
cc_68 VNB N_A_1586_74#_c_1168_n 0.00279267f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_1586_74#_c_1169_n 0.017477f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_1586_74#_c_1170_n 5.87492e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_1586_74#_c_1171_n 0.0022144f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_1586_74#_c_1172_n 0.0434353f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_1586_74#_c_1173_n 0.0082121f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_1586_74#_c_1174_n 0.00904398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_1586_74#_c_1175_n 0.00203028f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_1586_74#_c_1176_n 0.00953978f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_1586_74#_c_1177_n 0.00466954f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_1586_74#_c_1178_n 0.00313816f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_1586_74#_c_1179_n 0.00318285f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_1586_74#_c_1180_n 0.00302573f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_1586_74#_c_1181_n 0.0116019f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_1586_74#_c_1182_n 0.00571213f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_1586_74#_c_1183_n 0.00123754f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_1586_74#_c_1184_n 0.00280784f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_1586_74#_c_1185_n 0.0296806f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_1586_74#_c_1186_n 0.0174662f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_1374_368#_M1003_g 0.0392551f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=0.98
cc_88 VNB N_A_1374_368#_c_1403_n 0.00338809f $X=-0.19 $Y=-0.245 $X2=0.635
+ $Y2=1.58
cc_89 VNB N_A_1374_368#_c_1404_n 0.0154657f $X=-0.19 $Y=-0.245 $X2=0.54
+ $Y2=1.145
cc_90 VNB N_A_1374_368#_M1037_g 0.053968f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.825
cc_91 VNB N_A_1374_368#_c_1406_n 0.030791f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.145
cc_92 VNB N_A_1374_368#_c_1407_n 0.0151197f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_1374_368#_M1013_g 0.0511607f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_1374_368#_c_1409_n 0.00657241f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_1374_368#_c_1410_n 0.00119395f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_1374_368#_c_1411_n 0.0123224f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_1374_368#_c_1412_n 0.010047f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_A_1374_368#_c_1413_n 0.00894163f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_A_1374_368#_c_1414_n 0.00381838f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_A_1374_368#_c_1415_n 0.0326992f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_A_2013_71#_M1034_g 0.030024f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_A_2013_71#_c_1593_n 0.00884039f $X=-0.19 $Y=-0.245 $X2=0.635
+ $Y2=1.21
cc_103 VNB N_A_2013_71#_c_1594_n 0.0300468f $X=-0.19 $Y=-0.245 $X2=0.54
+ $Y2=1.145
cc_104 VNB N_A_2013_71#_c_1595_n 0.0086274f $X=-0.19 $Y=-0.245 $X2=0.54
+ $Y2=1.145
cc_105 VNB N_A_2013_71#_c_1596_n 0.0198235f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.99
cc_106 VNB N_A_2013_71#_c_1597_n 0.00999316f $X=-0.19 $Y=-0.245 $X2=0.63
+ $Y2=1.295
cc_107 VNB N_A_2013_71#_c_1598_n 0.00548308f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_A_2013_71#_c_1599_n 0.00253632f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_A_2013_71#_c_1600_n 0.00496828f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_A_2013_71#_c_1601_n 0.00184523f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_A_2013_71#_c_1602_n 0.0564399f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_A_2013_71#_c_1603_n 0.00274233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_A_2013_71#_c_1604_n 0.0364327f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_A_1784_97#_c_1706_n 0.0192526f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.58
cc_115 VNB N_A_1784_97#_M1023_g 0.0420339f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_116 VNB N_A_1784_97#_c_1708_n 0.013135f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.825
cc_117 VNB N_A_2489_74#_M1014_g 0.0257653f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_118 VNB N_A_2489_74#_c_1792_n 0.0754252f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_A_2489_74#_c_1793_n 0.0317828f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_A_2489_74#_M1032_g 0.022963f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.825
cc_121 VNB N_A_2489_74#_M1043_g 0.0208419f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_A_2489_74#_c_1796_n 0.0427532f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB N_A_2489_74#_c_1797_n 0.00286498f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_A_2489_74#_c_1798_n 0.00321929f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_A_2489_74#_c_1799_n 0.00525878f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_A_2489_74#_c_1800_n 0.00283454f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_A_2489_74#_c_1801_n 0.0083479f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_A_32_74#_c_1946_n 0.0434942f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_A_32_74#_c_1947_n 0.00382371f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_A_32_74#_c_1948_n 0.00641878f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_A_32_74#_c_1949_n 0.0138478f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_A_32_74#_c_1950_n 0.00433514f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_VPWR_c_2066_n 0.720949f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_A_691_113#_c_2266_n 0.0105451f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_A_691_113#_c_2267_n 0.0100696f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_A_691_113#_c_2268_n 0.0104521f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_A_691_113#_c_2269_n 0.00181722f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB N_A_691_113#_c_2270_n 0.0173316f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VNB N_A_691_113#_c_2271_n 0.00973194f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_A_691_113#_c_2272_n 0.00794098f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_141 VNB N_A_691_113#_c_2273_n 0.0192996f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_142 VNB Q 0.00240191f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.58
cc_143 VNB N_Q_N_c_2476_n 0.0132008f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.58
cc_144 VNB N_Q_N_c_2477_n 0.0239423f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.58
cc_145 VNB Q_N 0.00239713f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_146 VNB N_VGND_c_2509_n 0.0193314f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_147 VNB N_VGND_c_2510_n 0.0301467f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_148 VNB N_VGND_c_2511_n 0.0105113f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_149 VNB N_VGND_c_2512_n 0.0172622f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_150 VNB N_VGND_c_2513_n 0.00978559f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_151 VNB N_VGND_c_2514_n 0.0106328f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_152 VNB N_VGND_c_2515_n 0.00590394f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_153 VNB N_VGND_c_2516_n 0.0119255f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_154 VNB N_VGND_c_2517_n 0.00982717f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_155 VNB N_VGND_c_2518_n 0.00206318f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_156 VNB N_VGND_c_2519_n 0.0206041f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_157 VNB N_VGND_c_2520_n 0.0192796f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_158 VNB N_VGND_c_2521_n 0.0192531f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_159 VNB N_VGND_c_2522_n 0.00984545f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_160 VNB N_VGND_c_2523_n 0.0124653f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_161 VNB N_VGND_c_2524_n 0.0280494f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_162 VNB N_VGND_c_2525_n 0.023012f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_163 VNB N_VGND_c_2526_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_164 VNB N_VGND_c_2527_n 0.0220562f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_165 VNB N_VGND_c_2528_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_166 VNB N_VGND_c_2529_n 0.0403351f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_167 VNB N_VGND_c_2530_n 0.032665f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_168 VNB N_VGND_c_2531_n 0.0688863f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_169 VNB N_VGND_c_2532_n 0.0331395f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_170 VNB N_VGND_c_2533_n 0.0636008f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_171 VNB N_VGND_c_2534_n 0.0296519f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_172 VNB N_VGND_c_2535_n 0.019013f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_173 VNB N_VGND_c_2536_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_174 VNB N_VGND_c_2537_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_175 VNB N_VGND_c_2538_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_176 VNB N_VGND_c_2539_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_177 VNB N_VGND_c_2540_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_178 VNB N_VGND_c_2541_n 0.0112842f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_179 VNB N_VGND_c_2542_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_180 VNB N_VGND_c_2543_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_181 VNB N_VGND_c_2544_n 0.938824f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_182 VPB N_D_c_350_n 0.00985685f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=2.155
cc_183 VPB N_D_c_351_n 0.0256671f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=2.245
cc_184 VPB N_D_c_348_n 0.00461728f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.145
cc_185 VPB N_D_c_349_n 0.0112765f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.825
cc_186 VPB N_D_c_354_n 0.0156268f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.99
cc_187 VPB N_A_183_290#_c_397_n 0.0184393f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=0.58
cc_188 VPB N_A_183_290#_c_398_n 0.03334f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_189 VPB N_A_183_290#_c_391_n 0.020582f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.145
cc_190 VPB N_A_183_290#_c_400_n 0.0113728f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.825
cc_191 VPB N_A_183_290#_c_401_n 0.00224433f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.99
cc_192 VPB N_A_183_290#_c_402_n 0.00268948f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.825
cc_193 VPB N_A_183_290#_c_403_n 0.0123271f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_194 VPB N_A_183_290#_c_395_n 0.00274132f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_195 VPB N_A_183_290#_c_396_n 0.0179737f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_196 VPB N_A_183_290#_c_406_n 0.00136575f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_197 VPB N_DE_c_511_n 0.0193526f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_198 VPB N_DE_c_512_n 0.011356f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_199 VPB N_DE_c_513_n 0.0115848f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_200 VPB N_DE_c_514_n 0.0170592f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.145
cc_201 VPB N_DE_c_515_n 0.0413577f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.825
cc_202 VPB N_DE_c_516_n 0.0151132f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.99
cc_203 VPB N_DE_c_517_n 0.00666874f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_204 VPB DE 0.0020259f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.665
cc_205 VPB N_DE_c_509_n 0.0123229f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_206 VPB N_A_575_87#_c_615_n 0.0216256f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_207 VPB N_A_575_87#_c_616_n 0.0201112f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_208 VPB N_A_575_87#_c_617_n 0.0537867f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.825
cc_209 VPB N_A_575_87#_c_601_n 0.0227764f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_210 VPB N_A_575_87#_c_619_n 0.015159f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.825
cc_211 VPB N_A_575_87#_c_620_n 0.0175065f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_212 VPB N_A_575_87#_c_621_n 0.0059015f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_213 VPB N_A_575_87#_c_604_n 0.0151067f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_214 VPB N_A_575_87#_c_623_n 0.00879621f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_215 VPB N_A_575_87#_c_607_n 0.0029429f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_216 VPB N_A_575_87#_c_610_n 0.0575069f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_217 VPB N_A_575_87#_c_611_n 0.00131138f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_218 VPB N_A_575_87#_c_612_n 0.00129194f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_219 VPB N_A_575_87#_c_613_n 0.0226993f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_220 VPB N_A_575_87#_c_614_n 0.0149891f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_221 VPB N_A_661_87#_c_896_n 0.016921f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_222 VPB N_A_661_87#_c_897_n 0.0354087f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.145
cc_223 VPB N_A_661_87#_c_898_n 0.00434515f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_224 VPB N_A_661_87#_c_899_n 0.0208166f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.825
cc_225 VPB N_A_661_87#_c_900_n 0.00321747f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_226 VPB N_A_661_87#_c_894_n 0.0418704f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_227 VPB N_A_661_87#_c_902_n 0.00985185f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_228 VPB N_A_661_87#_c_903_n 0.00242577f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_229 VPB N_A_661_87#_c_895_n 0.0173634f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_230 VPB N_SCD_c_998_n 0.0256075f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=2.155
cc_231 VPB N_SCD_c_1003_n 0.0221674f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=2.245
cc_232 VPB N_SCE_c_1051_n 0.0189243f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.99
cc_233 VPB N_SCE_c_1052_n 0.0844158f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=2.64
cc_234 VPB N_SCE_c_1053_n 0.0133945f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=2.64
cc_235 VPB N_SCE_c_1044_n 0.0258986f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=0.58
cc_236 VPB N_SCE_c_1055_n 0.00754596f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=0.58
cc_237 VPB N_SCE_M1045_g 0.00964732f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=0.98
cc_238 VPB N_CLK_c_1127_n 0.0293371f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.99
cc_239 VPB N_A_1586_74#_c_1187_n 0.01905f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=0.58
cc_240 VPB N_A_1586_74#_c_1165_n 0.0376285f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.145
cc_241 VPB N_A_1586_74#_c_1189_n 0.0219712f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.145
cc_242 VPB N_A_1586_74#_c_1190_n 0.00468789f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.665
cc_243 VPB N_A_1586_74#_c_1180_n 0.00648383f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_244 VPB N_A_1586_74#_c_1192_n 0.00503963f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_245 VPB N_A_1586_74#_c_1182_n 0.00178697f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_246 VPB N_A_1586_74#_c_1194_n 0.061127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_247 VPB N_A_1586_74#_c_1186_n 0.0189353f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_248 VPB N_A_1374_368#_c_1403_n 0.0060259f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_249 VPB N_A_1374_368#_c_1417_n 0.0215025f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_250 VPB N_A_1374_368#_c_1404_n 0.0195938f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.145
cc_251 VPB N_A_1374_368#_c_1406_n 0.0199367f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.145
cc_252 VPB N_A_1374_368#_c_1420_n 0.0180856f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_253 VPB N_A_1374_368#_c_1421_n 0.0538565f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.665
cc_254 VPB N_A_1374_368#_c_1407_n 0.0440014f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_255 VPB N_A_1374_368#_c_1409_n 0.00438246f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_256 VPB N_A_1374_368#_c_1410_n 0.00298346f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_257 VPB N_A_1374_368#_c_1425_n 0.0040461f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_258 VPB N_A_1374_368#_c_1426_n 0.0121562f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_259 VPB N_A_1374_368#_c_1427_n 0.00261599f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_260 VPB N_A_1374_368#_c_1412_n 0.00682253f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_261 VPB N_A_1374_368#_c_1429_n 0.0406368f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_262 VPB N_A_1374_368#_c_1430_n 0.00756028f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_263 VPB N_A_1374_368#_c_1414_n 0.00210725f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_264 VPB N_A_1374_368#_c_1415_n 0.0153862f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_265 VPB N_A_2013_71#_c_1593_n 0.0417122f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_266 VPB N_A_2013_71#_c_1606_n 0.0228032f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_267 VPB N_A_2013_71#_c_1595_n 0.00835609f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.145
cc_268 VPB N_A_2013_71#_c_1608_n 0.0291381f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.825
cc_269 VPB N_A_2013_71#_c_1609_n 0.00602683f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.665
cc_270 VPB N_A_2013_71#_c_1599_n 0.00903944f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_271 VPB N_A_1784_97#_c_1706_n 0.0440232f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=0.58
cc_272 VPB N_A_1784_97#_c_1710_n 0.0162618f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.825
cc_273 VPB N_A_1784_97#_c_1711_n 0.00117381f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.825
cc_274 VPB N_A_1784_97#_c_1712_n 0.00492079f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.145
cc_275 VPB N_A_1784_97#_c_1713_n 0.00721525f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_276 VPB N_A_1784_97#_c_1714_n 0.0017703f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.665
cc_277 VPB N_A_2489_74#_c_1802_n 0.0192283f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=0.58
cc_278 VPB N_A_2489_74#_c_1793_n 0.00809164f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_279 VPB N_A_2489_74#_c_1804_n 0.0169125f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.825
cc_280 VPB N_A_2489_74#_c_1805_n 0.0148841f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_281 VPB N_A_2489_74#_c_1796_n 0.0128322f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_282 VPB N_A_2489_74#_c_1807_n 0.00595698f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_283 VPB N_A_2489_74#_c_1808_n 0.0110034f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_284 VPB N_A_2489_74#_c_1809_n 0.0015169f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_285 VPB N_A_2489_74#_c_1800_n 0.0014512f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_286 VPB N_A_2489_74#_c_1811_n 0.00455915f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_287 VPB N_A_32_74#_c_1946_n 0.0303411f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_288 VPB N_A_32_74#_c_1952_n 0.026226f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.145
cc_289 VPB N_A_32_74#_c_1953_n 0.015704f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.145
cc_290 VPB N_A_32_74#_c_1954_n 0.00998336f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.825
cc_291 VPB N_A_32_74#_c_1955_n 0.00941149f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.99
cc_292 VPB N_A_32_74#_c_1956_n 0.00349119f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.145
cc_293 VPB N_A_32_74#_c_1957_n 0.00718892f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_294 VPB N_A_32_74#_c_1958_n 0.00104602f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.665
cc_295 VPB N_A_32_74#_c_1948_n 0.0123413f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_296 VPB N_A_32_74#_c_1960_n 0.0140676f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_297 VPB N_A_32_74#_c_1961_n 0.00428149f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_298 VPB N_VPWR_c_2067_n 0.00600898f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_299 VPB N_VPWR_c_2068_n 0.00589284f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_300 VPB N_VPWR_c_2069_n 0.00823648f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_301 VPB N_VPWR_c_2070_n 0.00751218f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_302 VPB N_VPWR_c_2071_n 0.0220447f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_303 VPB N_VPWR_c_2072_n 0.0115779f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_304 VPB N_VPWR_c_2073_n 0.0162479f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_305 VPB N_VPWR_c_2074_n 0.00880467f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_306 VPB N_VPWR_c_2075_n 0.00916914f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_307 VPB N_VPWR_c_2076_n 0.00261791f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_308 VPB N_VPWR_c_2077_n 0.0120106f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_309 VPB N_VPWR_c_2078_n 0.0405468f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_310 VPB N_VPWR_c_2079_n 0.0342477f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_311 VPB N_VPWR_c_2080_n 0.00460249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_312 VPB N_VPWR_c_2081_n 0.0242802f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_313 VPB N_VPWR_c_2082_n 0.00632182f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_314 VPB N_VPWR_c_2083_n 0.0324541f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_315 VPB N_VPWR_c_2084_n 0.0296515f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_316 VPB N_VPWR_c_2085_n 0.0590043f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_317 VPB N_VPWR_c_2086_n 0.0335097f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_318 VPB N_VPWR_c_2087_n 0.059622f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_319 VPB N_VPWR_c_2088_n 0.0636904f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_320 VPB N_VPWR_c_2089_n 0.0203698f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_321 VPB N_VPWR_c_2090_n 0.0177589f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_322 VPB N_VPWR_c_2091_n 0.01587f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_323 VPB N_VPWR_c_2092_n 0.00460249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_324 VPB N_VPWR_c_2093_n 0.00467461f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_325 VPB N_VPWR_c_2094_n 0.00516749f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_326 VPB N_VPWR_c_2095_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_327 VPB N_VPWR_c_2096_n 0.00615076f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_328 VPB N_VPWR_c_2097_n 0.0101806f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_329 VPB N_VPWR_c_2098_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_330 VPB N_VPWR_c_2099_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_331 VPB N_VPWR_c_2066_n 0.211753f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_332 VPB N_A_691_113#_c_2274_n 0.00174855f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.825
cc_333 VPB N_A_691_113#_c_2275_n 0.0119484f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_334 VPB N_A_691_113#_c_2276_n 0.00810814f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_335 VPB N_A_691_113#_c_2277_n 0.001333f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.825
cc_336 VPB N_A_691_113#_c_2267_n 0.00915521f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_337 VPB N_A_691_113#_c_2279_n 0.0192891f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_338 VPB N_A_691_113#_c_2280_n 0.0204232f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_339 VPB N_A_691_113#_c_2281_n 0.00161618f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_340 VPB N_A_691_113#_c_2282_n 0.00986275f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_341 VPB N_A_691_113#_c_2283_n 0.00723316f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_342 VPB N_A_691_113#_c_2272_n 0.0099146f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_343 VPB N_Q_N_c_2477_n 0.017779f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=0.58
cc_344 VPB Q_N 0.00281782f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_345 N_D_c_351_n N_A_183_290#_c_397_n 0.0383559f $X=0.585 $Y=2.245 $X2=0 $Y2=0
cc_346 N_D_c_350_n N_A_183_290#_c_398_n 0.0143845f $X=0.585 $Y=2.155 $X2=0 $Y2=0
cc_347 N_D_c_354_n N_A_183_290#_c_398_n 0.0169614f $X=0.54 $Y=1.99 $X2=0 $Y2=0
cc_348 N_D_c_348_n N_A_183_290#_c_390_n 0.0545333f $X=0.54 $Y=1.145 $X2=0 $Y2=0
cc_349 N_D_c_349_n N_A_183_290#_c_390_n 0.00133474f $X=0.54 $Y=1.825 $X2=0 $Y2=0
cc_350 N_D_c_348_n N_A_183_290#_c_391_n 0.00384651f $X=0.54 $Y=1.145 $X2=0 $Y2=0
cc_351 N_D_c_349_n N_A_183_290#_c_391_n 0.0169614f $X=0.54 $Y=1.825 $X2=0 $Y2=0
cc_352 N_D_c_348_n N_A_183_290#_c_393_n 0.0148197f $X=0.54 $Y=1.145 $X2=0 $Y2=0
cc_353 N_D_c_349_n N_A_183_290#_c_393_n 4.03978e-19 $X=0.54 $Y=1.825 $X2=0 $Y2=0
cc_354 N_D_c_350_n N_A_183_290#_c_401_n 6.9419e-19 $X=0.585 $Y=2.155 $X2=0 $Y2=0
cc_355 N_D_c_348_n N_A_183_290#_c_401_n 0.00341199f $X=0.54 $Y=1.145 $X2=0 $Y2=0
cc_356 N_D_M1047_g N_DE_M1042_g 0.025244f $X=0.63 $Y=0.58 $X2=0 $Y2=0
cc_357 N_D_c_348_n N_DE_M1042_g 0.00420913f $X=0.54 $Y=1.145 $X2=0 $Y2=0
cc_358 N_D_c_347_n N_DE_c_504_n 0.025244f $X=0.54 $Y=1.145 $X2=0 $Y2=0
cc_359 N_D_c_350_n N_A_32_74#_c_1946_n 0.00823508f $X=0.585 $Y=2.155 $X2=0 $Y2=0
cc_360 N_D_c_351_n N_A_32_74#_c_1946_n 0.00137514f $X=0.585 $Y=2.245 $X2=0 $Y2=0
cc_361 N_D_M1047_g N_A_32_74#_c_1946_n 0.00669921f $X=0.63 $Y=0.58 $X2=0 $Y2=0
cc_362 N_D_c_347_n N_A_32_74#_c_1946_n 0.0239763f $X=0.54 $Y=1.145 $X2=0 $Y2=0
cc_363 N_D_c_348_n N_A_32_74#_c_1946_n 0.0771054f $X=0.54 $Y=1.145 $X2=0 $Y2=0
cc_364 N_D_c_351_n N_A_32_74#_c_1952_n 0.00949192f $X=0.585 $Y=2.245 $X2=0 $Y2=0
cc_365 N_D_c_351_n N_A_32_74#_c_1953_n 0.0127112f $X=0.585 $Y=2.245 $X2=0 $Y2=0
cc_366 N_D_c_348_n N_A_32_74#_c_1953_n 0.0161746f $X=0.54 $Y=1.145 $X2=0 $Y2=0
cc_367 N_D_M1047_g N_A_32_74#_c_1949_n 0.0058515f $X=0.63 $Y=0.58 $X2=0 $Y2=0
cc_368 N_D_c_347_n N_A_32_74#_c_1949_n 0.00276862f $X=0.54 $Y=1.145 $X2=0 $Y2=0
cc_369 N_D_c_348_n N_A_32_74#_c_1949_n 0.00757623f $X=0.54 $Y=1.145 $X2=0 $Y2=0
cc_370 N_D_c_351_n N_A_32_74#_c_1960_n 0.00164796f $X=0.585 $Y=2.245 $X2=0 $Y2=0
cc_371 N_D_c_348_n N_A_32_74#_c_1960_n 0.00569905f $X=0.54 $Y=1.145 $X2=0 $Y2=0
cc_372 N_D_c_354_n N_A_32_74#_c_1960_n 0.00263932f $X=0.54 $Y=1.99 $X2=0 $Y2=0
cc_373 N_D_c_351_n N_VPWR_c_2067_n 0.001556f $X=0.585 $Y=2.245 $X2=0 $Y2=0
cc_374 N_D_c_351_n N_VPWR_c_2083_n 0.00445602f $X=0.585 $Y=2.245 $X2=0 $Y2=0
cc_375 N_D_c_351_n N_VPWR_c_2066_n 0.00861888f $X=0.585 $Y=2.245 $X2=0 $Y2=0
cc_376 N_D_M1047_g N_VGND_c_2509_n 0.00218592f $X=0.63 $Y=0.58 $X2=0 $Y2=0
cc_377 N_D_M1047_g N_VGND_c_2530_n 0.004347f $X=0.63 $Y=0.58 $X2=0 $Y2=0
cc_378 N_D_M1047_g N_VGND_c_2544_n 0.00822933f $X=0.63 $Y=0.58 $X2=0 $Y2=0
cc_379 N_A_183_290#_c_394_n N_DE_M1042_g 0.00659112f $X=1.845 $Y=0.775 $X2=0
+ $Y2=0
cc_380 N_A_183_290#_c_392_n N_DE_c_503_n 0.0130203f $X=1.68 $Y=1.195 $X2=0 $Y2=0
cc_381 N_A_183_290#_c_393_n N_DE_c_503_n 0.00791665f $X=1.335 $Y=1.195 $X2=0
+ $Y2=0
cc_382 N_A_183_290#_c_391_n N_DE_c_504_n 0.0226593f $X=1.17 $Y=1.615 $X2=0 $Y2=0
cc_383 N_A_183_290#_c_393_n N_DE_c_504_n 0.00629125f $X=1.335 $Y=1.195 $X2=0
+ $Y2=0
cc_384 N_A_183_290#_c_392_n N_DE_c_505_n 0.00690186f $X=1.68 $Y=1.195 $X2=0
+ $Y2=0
cc_385 N_A_183_290#_c_394_n N_DE_c_505_n 0.00596863f $X=1.845 $Y=0.775 $X2=0
+ $Y2=0
cc_386 N_A_183_290#_c_390_n N_DE_c_511_n 9.54411e-19 $X=1.17 $Y=1.615 $X2=0
+ $Y2=0
cc_387 N_A_183_290#_c_391_n N_DE_c_511_n 0.00491474f $X=1.17 $Y=1.615 $X2=0
+ $Y2=0
cc_388 N_A_183_290#_c_400_n N_DE_c_511_n 0.00391046f $X=1.825 $Y=2.035 $X2=0
+ $Y2=0
cc_389 N_A_183_290#_c_395_n N_DE_c_511_n 0.00303743f $X=2.47 $Y=1.68 $X2=0 $Y2=0
cc_390 N_A_183_290#_c_406_n N_DE_c_511_n 0.00539719f $X=1.91 $Y=2.035 $X2=0
+ $Y2=0
cc_391 N_A_183_290#_c_402_n N_DE_c_512_n 0.00796868f $X=1.91 $Y=2.51 $X2=0 $Y2=0
cc_392 N_A_183_290#_c_403_n N_DE_c_512_n 0.00366629f $X=2.305 $Y=2.035 $X2=0
+ $Y2=0
cc_393 N_A_183_290#_c_406_n N_DE_c_512_n 0.00180964f $X=1.91 $Y=2.035 $X2=0
+ $Y2=0
cc_394 N_A_183_290#_c_398_n N_DE_c_513_n 0.00794913f $X=1.125 $Y=1.91 $X2=0
+ $Y2=0
cc_395 N_A_183_290#_c_400_n N_DE_c_513_n 0.00339243f $X=1.825 $Y=2.035 $X2=0
+ $Y2=0
cc_396 N_A_183_290#_c_402_n N_DE_c_513_n 0.00689062f $X=1.91 $Y=2.51 $X2=0 $Y2=0
cc_397 N_A_183_290#_c_406_n N_DE_c_513_n 2.6366e-19 $X=1.91 $Y=2.035 $X2=0 $Y2=0
cc_398 N_A_183_290#_M1024_g N_DE_c_506_n 0.0184318f $X=2.56 $Y=0.775 $X2=0 $Y2=0
cc_399 N_A_183_290#_c_394_n N_DE_c_506_n 0.00860606f $X=1.845 $Y=0.775 $X2=0
+ $Y2=0
cc_400 N_A_183_290#_c_402_n N_DE_c_514_n 0.00434248f $X=1.91 $Y=2.51 $X2=0 $Y2=0
cc_401 N_A_183_290#_c_403_n N_DE_c_515_n 0.0108361f $X=2.305 $Y=2.035 $X2=0
+ $Y2=0
cc_402 N_A_183_290#_c_396_n N_DE_c_515_n 0.0181259f $X=2.47 $Y=1.68 $X2=0 $Y2=0
cc_403 N_A_183_290#_c_392_n N_DE_c_507_n 0.00525481f $X=1.68 $Y=1.195 $X2=0
+ $Y2=0
cc_404 N_A_183_290#_c_394_n N_DE_c_507_n 0.00353956f $X=1.845 $Y=0.775 $X2=0
+ $Y2=0
cc_405 N_A_183_290#_c_403_n N_DE_c_517_n 0.00829073f $X=2.305 $Y=2.035 $X2=0
+ $Y2=0
cc_406 N_A_183_290#_M1024_g DE 3.21021e-19 $X=2.56 $Y=0.775 $X2=0 $Y2=0
cc_407 N_A_183_290#_c_390_n DE 0.020843f $X=1.17 $Y=1.615 $X2=0 $Y2=0
cc_408 N_A_183_290#_c_391_n DE 0.00206473f $X=1.17 $Y=1.615 $X2=0 $Y2=0
cc_409 N_A_183_290#_c_392_n DE 0.0270293f $X=1.68 $Y=1.195 $X2=0 $Y2=0
cc_410 N_A_183_290#_c_400_n DE 0.019286f $X=1.825 $Y=2.035 $X2=0 $Y2=0
cc_411 N_A_183_290#_c_395_n DE 0.00999033f $X=2.47 $Y=1.68 $X2=0 $Y2=0
cc_412 N_A_183_290#_c_396_n DE 0.00111448f $X=2.47 $Y=1.68 $X2=0 $Y2=0
cc_413 N_A_183_290#_c_406_n DE 0.00638598f $X=1.91 $Y=2.035 $X2=0 $Y2=0
cc_414 N_A_183_290#_M1024_g N_DE_c_509_n 9.94929e-19 $X=2.56 $Y=0.775 $X2=0
+ $Y2=0
cc_415 N_A_183_290#_c_390_n N_DE_c_509_n 4.11485e-19 $X=1.17 $Y=1.615 $X2=0
+ $Y2=0
cc_416 N_A_183_290#_c_391_n N_DE_c_509_n 0.0179198f $X=1.17 $Y=1.615 $X2=0 $Y2=0
cc_417 N_A_183_290#_c_392_n N_DE_c_509_n 0.00127783f $X=1.68 $Y=1.195 $X2=0
+ $Y2=0
cc_418 N_A_183_290#_c_400_n N_DE_c_509_n 0.00462669f $X=1.825 $Y=2.035 $X2=0
+ $Y2=0
cc_419 N_A_183_290#_c_395_n N_DE_c_509_n 7.04955e-19 $X=2.47 $Y=1.68 $X2=0 $Y2=0
cc_420 N_A_183_290#_c_396_n N_DE_c_509_n 0.00950624f $X=2.47 $Y=1.68 $X2=0 $Y2=0
cc_421 N_A_183_290#_c_390_n N_DE_c_510_n 0.00581511f $X=1.17 $Y=1.615 $X2=0
+ $Y2=0
cc_422 N_A_183_290#_c_392_n N_DE_c_510_n 0.00597544f $X=1.68 $Y=1.195 $X2=0
+ $Y2=0
cc_423 N_A_183_290#_M1024_g N_A_575_87#_M1006_g 0.0369397f $X=2.56 $Y=0.775
+ $X2=0 $Y2=0
cc_424 N_A_183_290#_c_403_n N_A_575_87#_c_615_n 0.00421101f $X=2.305 $Y=2.035
+ $X2=0 $Y2=0
cc_425 N_A_183_290#_c_395_n N_A_575_87#_c_615_n 0.00283945f $X=2.47 $Y=1.68
+ $X2=0 $Y2=0
cc_426 N_A_183_290#_c_395_n N_A_575_87#_c_633_n 0.00127953f $X=2.47 $Y=1.68
+ $X2=0 $Y2=0
cc_427 N_A_183_290#_c_395_n N_A_575_87#_c_612_n 0.0172952f $X=2.47 $Y=1.68 $X2=0
+ $Y2=0
cc_428 N_A_183_290#_c_396_n N_A_575_87#_c_612_n 0.00120934f $X=2.47 $Y=1.68
+ $X2=0 $Y2=0
cc_429 N_A_183_290#_c_395_n N_A_575_87#_c_613_n 4.18224e-19 $X=2.47 $Y=1.68
+ $X2=0 $Y2=0
cc_430 N_A_183_290#_c_396_n N_A_575_87#_c_613_n 0.0369397f $X=2.47 $Y=1.68 $X2=0
+ $Y2=0
cc_431 N_A_183_290#_c_397_n N_A_32_74#_c_1952_n 0.00181882f $X=1.005 $Y=2.245
+ $X2=0 $Y2=0
cc_432 N_A_183_290#_c_397_n N_A_32_74#_c_1953_n 0.0184872f $X=1.005 $Y=2.245
+ $X2=0 $Y2=0
cc_433 N_A_183_290#_c_398_n N_A_32_74#_c_1953_n 0.00284279f $X=1.125 $Y=1.91
+ $X2=0 $Y2=0
cc_434 N_A_183_290#_c_400_n N_A_32_74#_c_1953_n 0.0255781f $X=1.825 $Y=2.035
+ $X2=0 $Y2=0
cc_435 N_A_183_290#_c_401_n N_A_32_74#_c_1953_n 0.0260073f $X=1.335 $Y=2.035
+ $X2=0 $Y2=0
cc_436 N_A_183_290#_c_402_n N_A_32_74#_c_1953_n 0.0141582f $X=1.91 $Y=2.51 $X2=0
+ $Y2=0
cc_437 N_A_183_290#_c_397_n N_A_32_74#_c_1954_n 0.00426176f $X=1.005 $Y=2.245
+ $X2=0 $Y2=0
cc_438 N_A_183_290#_c_402_n N_A_32_74#_c_1954_n 0.0203028f $X=1.91 $Y=2.51 $X2=0
+ $Y2=0
cc_439 N_A_183_290#_M1017_s N_A_32_74#_c_1955_n 0.0031801f $X=1.765 $Y=2.31
+ $X2=0 $Y2=0
cc_440 N_A_183_290#_c_402_n N_A_32_74#_c_1955_n 0.012787f $X=1.91 $Y=2.51 $X2=0
+ $Y2=0
cc_441 N_A_183_290#_c_397_n N_A_32_74#_c_1956_n 6.5162e-19 $X=1.005 $Y=2.245
+ $X2=0 $Y2=0
cc_442 N_A_183_290#_c_402_n N_A_32_74#_c_1987_n 0.0192722f $X=1.91 $Y=2.51 $X2=0
+ $Y2=0
cc_443 N_A_183_290#_c_403_n N_A_32_74#_c_1957_n 0.0237119f $X=2.305 $Y=2.035
+ $X2=0 $Y2=0
cc_444 N_A_183_290#_c_402_n N_A_32_74#_c_1958_n 0.0133878f $X=1.91 $Y=2.51 $X2=0
+ $Y2=0
cc_445 N_A_183_290#_c_403_n N_A_32_74#_c_1958_n 0.0136791f $X=2.305 $Y=2.035
+ $X2=0 $Y2=0
cc_446 N_A_183_290#_M1024_g N_A_32_74#_c_1947_n 0.00214472f $X=2.56 $Y=0.775
+ $X2=0 $Y2=0
cc_447 N_A_183_290#_M1024_g N_A_32_74#_c_1950_n 8.2814e-19 $X=2.56 $Y=0.775
+ $X2=0 $Y2=0
cc_448 N_A_183_290#_c_397_n N_VPWR_c_2067_n 0.0107235f $X=1.005 $Y=2.245 $X2=0
+ $Y2=0
cc_449 N_A_183_290#_c_397_n N_VPWR_c_2083_n 0.00413917f $X=1.005 $Y=2.245 $X2=0
+ $Y2=0
cc_450 N_A_183_290#_c_397_n N_VPWR_c_2066_n 0.00817532f $X=1.005 $Y=2.245 $X2=0
+ $Y2=0
cc_451 N_A_183_290#_c_391_n N_VGND_c_2509_n 2.63289e-19 $X=1.17 $Y=1.615 $X2=0
+ $Y2=0
cc_452 N_A_183_290#_c_392_n N_VGND_c_2509_n 0.00336712f $X=1.68 $Y=1.195 $X2=0
+ $Y2=0
cc_453 N_A_183_290#_c_393_n N_VGND_c_2509_n 0.0152311f $X=1.335 $Y=1.195 $X2=0
+ $Y2=0
cc_454 N_A_183_290#_c_394_n N_VGND_c_2509_n 0.0156036f $X=1.845 $Y=0.775 $X2=0
+ $Y2=0
cc_455 N_A_183_290#_M1024_g N_VGND_c_2510_n 0.0129344f $X=2.56 $Y=0.775 $X2=0
+ $Y2=0
cc_456 N_A_183_290#_c_394_n N_VGND_c_2510_n 0.0188413f $X=1.845 $Y=0.775 $X2=0
+ $Y2=0
cc_457 N_A_183_290#_c_395_n N_VGND_c_2510_n 0.00772803f $X=2.47 $Y=1.68 $X2=0
+ $Y2=0
cc_458 N_A_183_290#_c_396_n N_VGND_c_2510_n 0.0011905f $X=2.47 $Y=1.68 $X2=0
+ $Y2=0
cc_459 N_A_183_290#_c_394_n N_VGND_c_2525_n 0.00805126f $X=1.845 $Y=0.775 $X2=0
+ $Y2=0
cc_460 N_A_183_290#_M1024_g N_VGND_c_2531_n 0.00372658f $X=2.56 $Y=0.775 $X2=0
+ $Y2=0
cc_461 N_A_183_290#_M1024_g N_VGND_c_2544_n 0.00408518f $X=2.56 $Y=0.775 $X2=0
+ $Y2=0
cc_462 N_A_183_290#_c_394_n N_VGND_c_2544_n 0.0106012f $X=1.845 $Y=0.775 $X2=0
+ $Y2=0
cc_463 N_DE_c_515_n N_A_575_87#_c_615_n 0.0105652f $X=2.74 $Y=2.16 $X2=0 $Y2=0
cc_464 N_DE_c_516_n N_A_575_87#_c_616_n 0.043765f $X=2.815 $Y=2.235 $X2=0 $Y2=0
cc_465 N_DE_c_515_n N_A_575_87#_c_613_n 0.00173282f $X=2.74 $Y=2.16 $X2=0 $Y2=0
cc_466 N_DE_c_514_n N_A_32_74#_c_1954_n 0.00326422f $X=2.135 $Y=2.235 $X2=0
+ $Y2=0
cc_467 N_DE_c_512_n N_A_32_74#_c_1955_n 7.49315e-19 $X=2.06 $Y=2.16 $X2=0 $Y2=0
cc_468 N_DE_c_513_n N_A_32_74#_c_1955_n 0.00219966f $X=1.905 $Y=2.16 $X2=0 $Y2=0
cc_469 N_DE_c_514_n N_A_32_74#_c_1955_n 0.0134726f $X=2.135 $Y=2.235 $X2=0 $Y2=0
cc_470 N_DE_c_516_n N_A_32_74#_c_1955_n 4.32305e-19 $X=2.815 $Y=2.235 $X2=0
+ $Y2=0
cc_471 N_DE_c_514_n N_A_32_74#_c_1987_n 0.0118088f $X=2.135 $Y=2.235 $X2=0 $Y2=0
cc_472 N_DE_c_516_n N_A_32_74#_c_1987_n 0.00283455f $X=2.815 $Y=2.235 $X2=0
+ $Y2=0
cc_473 N_DE_c_515_n N_A_32_74#_c_1957_n 0.00753877f $X=2.74 $Y=2.16 $X2=0 $Y2=0
cc_474 N_DE_c_516_n N_A_32_74#_c_1957_n 0.0187002f $X=2.815 $Y=2.235 $X2=0 $Y2=0
cc_475 N_DE_c_514_n N_A_32_74#_c_1958_n 0.00588346f $X=2.135 $Y=2.235 $X2=0
+ $Y2=0
cc_476 N_DE_c_515_n N_A_32_74#_c_1958_n 8.05635e-19 $X=2.74 $Y=2.16 $X2=0 $Y2=0
cc_477 N_DE_M1042_g N_A_32_74#_c_1949_n 8.70603e-19 $X=1.02 $Y=0.58 $X2=0 $Y2=0
cc_478 N_DE_c_516_n N_A_32_74#_c_1961_n 0.00177861f $X=2.815 $Y=2.235 $X2=0
+ $Y2=0
cc_479 N_DE_c_514_n N_VPWR_c_2068_n 0.00142894f $X=2.135 $Y=2.235 $X2=0 $Y2=0
cc_480 N_DE_c_516_n N_VPWR_c_2068_n 0.00959893f $X=2.815 $Y=2.235 $X2=0 $Y2=0
cc_481 N_DE_c_514_n N_VPWR_c_2084_n 0.00390665f $X=2.135 $Y=2.235 $X2=0 $Y2=0
cc_482 N_DE_c_516_n N_VPWR_c_2085_n 0.00512473f $X=2.815 $Y=2.235 $X2=0 $Y2=0
cc_483 N_DE_c_514_n N_VPWR_c_2066_n 0.00542671f $X=2.135 $Y=2.235 $X2=0 $Y2=0
cc_484 N_DE_c_516_n N_VPWR_c_2066_n 0.00492022f $X=2.815 $Y=2.235 $X2=0 $Y2=0
cc_485 N_DE_M1042_g N_VGND_c_2509_n 0.0143553f $X=1.02 $Y=0.58 $X2=0 $Y2=0
cc_486 N_DE_c_503_n N_VGND_c_2509_n 0.00425745f $X=1.575 $Y=1.135 $X2=0 $Y2=0
cc_487 N_DE_c_506_n N_VGND_c_2509_n 0.00322863f $X=2.06 $Y=1.06 $X2=0 $Y2=0
cc_488 N_DE_c_506_n N_VGND_c_2510_n 0.00564371f $X=2.06 $Y=1.06 $X2=0 $Y2=0
cc_489 N_DE_c_506_n N_VGND_c_2525_n 0.00430863f $X=2.06 $Y=1.06 $X2=0 $Y2=0
cc_490 N_DE_M1042_g N_VGND_c_2530_n 0.00383152f $X=1.02 $Y=0.58 $X2=0 $Y2=0
cc_491 N_DE_M1042_g N_VGND_c_2544_n 0.0075725f $X=1.02 $Y=0.58 $X2=0 $Y2=0
cc_492 N_DE_c_506_n N_VGND_c_2544_n 0.00486331f $X=2.06 $Y=1.06 $X2=0 $Y2=0
cc_493 N_A_575_87#_M1006_g N_A_661_87#_c_887_n 0.0180128f $X=2.95 $Y=0.775 $X2=0
+ $Y2=0
cc_494 N_A_575_87#_c_610_n N_A_661_87#_c_888_n 0.00616126f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_495 N_A_575_87#_c_610_n N_A_661_87#_c_907_n 0.0186276f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_496 N_A_575_87#_c_610_n N_A_661_87#_c_892_n 0.00389277f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_497 N_A_575_87#_c_610_n N_A_661_87#_c_899_n 0.0516509f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_498 N_A_575_87#_c_610_n N_A_661_87#_c_900_n 0.00884701f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_499 N_A_575_87#_c_610_n N_A_661_87#_c_894_n 0.00594097f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_500 N_A_575_87#_c_613_n N_A_661_87#_c_894_n 0.00551319f $X=3.205 $Y=1.68
+ $X2=0 $Y2=0
cc_501 N_A_575_87#_c_610_n N_A_661_87#_c_902_n 0.00183705f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_502 N_A_575_87#_c_610_n N_A_661_87#_c_903_n 0.0192345f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_503 N_A_575_87#_c_610_n N_A_661_87#_c_895_n 0.00382946f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_504 N_A_575_87#_c_610_n N_SCD_c_998_n 0.00279625f $X=14.975 $Y=1.665 $X2=0
+ $Y2=0
cc_505 N_A_575_87#_c_610_n SCD 0.0135615f $X=14.975 $Y=1.665 $X2=0 $Y2=0
cc_506 N_A_575_87#_c_610_n N_SCD_c_1001_n 0.00380723f $X=14.975 $Y=1.665 $X2=0
+ $Y2=0
cc_507 N_A_575_87#_c_616_n N_SCE_c_1051_n 0.00740543f $X=3.205 $Y=2.235
+ $X2=-0.19 $Y2=-0.245
cc_508 N_A_575_87#_c_610_n N_SCE_c_1051_n 0.00322369f $X=14.975 $Y=1.665
+ $X2=-0.19 $Y2=-0.245
cc_509 N_A_575_87#_c_616_n N_SCE_c_1053_n 0.00286907f $X=3.205 $Y=2.235 $X2=0
+ $Y2=0
cc_510 N_A_575_87#_c_610_n N_SCE_c_1044_n 0.00267168f $X=14.975 $Y=1.665 $X2=0
+ $Y2=0
cc_511 N_A_575_87#_c_610_n N_SCE_M1036_g 5.5049e-19 $X=14.975 $Y=1.665 $X2=0
+ $Y2=0
cc_512 N_A_575_87#_c_610_n N_SCE_c_1049_n 0.0043941f $X=14.975 $Y=1.665 $X2=0
+ $Y2=0
cc_513 N_A_575_87#_c_610_n N_SCE_c_1050_n 0.0115832f $X=14.975 $Y=1.665 $X2=0
+ $Y2=0
cc_514 N_A_575_87#_c_610_n N_CLK_c_1127_n 0.00760554f $X=14.975 $Y=1.665
+ $X2=-0.19 $Y2=-0.245
cc_515 N_A_575_87#_c_610_n CLK 0.012981f $X=14.975 $Y=1.665 $X2=0 $Y2=0
cc_516 N_A_575_87#_c_617_n N_A_1586_74#_c_1165_n 0.0198888f $X=13.705 $Y=2.465
+ $X2=0 $Y2=0
cc_517 N_A_575_87#_c_601_n N_A_1586_74#_c_1165_n 0.0151002f $X=13.84 $Y=2.05
+ $X2=0 $Y2=0
cc_518 N_A_575_87#_c_621_n N_A_1586_74#_c_1165_n 0.00104433f $X=14.475 $Y=2.217
+ $X2=0 $Y2=0
cc_519 N_A_575_87#_c_610_n N_A_1586_74#_c_1165_n 0.00305397f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_520 N_A_575_87#_c_617_n N_A_1586_74#_c_1189_n 0.0320696f $X=13.705 $Y=2.465
+ $X2=0 $Y2=0
cc_521 N_A_575_87#_c_610_n N_A_1586_74#_c_1166_n 0.00221507f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_522 N_A_575_87#_c_610_n N_A_1586_74#_c_1190_n 0.0119703f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_523 N_A_575_87#_c_610_n N_A_1586_74#_c_1171_n 0.0070403f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_524 N_A_575_87#_c_610_n N_A_1586_74#_c_1172_n 7.16649e-19 $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_525 N_A_575_87#_c_610_n N_A_1586_74#_c_1173_n 0.00501141f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_526 N_A_575_87#_c_610_n N_A_1586_74#_c_1177_n 0.00603531f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_527 N_A_575_87#_c_610_n N_A_1586_74#_c_1178_n 3.66988e-19 $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_528 N_A_575_87#_c_610_n N_A_1586_74#_c_1180_n 0.0387409f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_529 N_A_575_87#_c_610_n N_A_1586_74#_c_1181_n 0.0165713f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_530 N_A_575_87#_c_610_n N_A_1586_74#_c_1192_n 0.00818568f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_531 N_A_575_87#_c_610_n N_A_1586_74#_c_1182_n 0.0201078f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_532 N_A_575_87#_c_610_n N_A_1586_74#_c_1194_n 0.0010178f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_533 N_A_575_87#_c_600_n N_A_1586_74#_c_1184_n 0.00221728f $X=13.345 $Y=0.94
+ $X2=0 $Y2=0
cc_534 N_A_575_87#_c_601_n N_A_1586_74#_c_1184_n 9.53696e-19 $X=13.84 $Y=2.05
+ $X2=0 $Y2=0
cc_535 N_A_575_87#_c_610_n N_A_1586_74#_c_1184_n 0.00886866f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_536 N_A_575_87#_c_600_n N_A_1586_74#_c_1185_n 0.0204808f $X=13.345 $Y=0.94
+ $X2=0 $Y2=0
cc_537 N_A_575_87#_c_601_n N_A_1586_74#_c_1185_n 0.0173096f $X=13.84 $Y=2.05
+ $X2=0 $Y2=0
cc_538 N_A_575_87#_c_610_n N_A_1586_74#_c_1185_n 0.00391026f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_539 N_A_575_87#_c_610_n N_A_1586_74#_c_1186_n 0.00371475f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_540 N_A_575_87#_c_610_n N_A_1374_368#_c_1404_n 0.00307977f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_541 N_A_575_87#_c_610_n N_A_1374_368#_c_1406_n 0.0122449f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_542 N_A_575_87#_c_610_n N_A_1374_368#_c_1407_n 6.94548e-19 $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_543 N_A_575_87#_c_598_n N_A_1374_368#_M1013_g 0.0417021f $X=13.27 $Y=0.865
+ $X2=0 $Y2=0
cc_544 N_A_575_87#_c_610_n N_A_1374_368#_c_1409_n 0.00236152f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_545 N_A_575_87#_c_610_n N_A_1374_368#_c_1410_n 0.00496775f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_546 N_A_575_87#_c_610_n N_A_1374_368#_c_1425_n 0.0146295f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_547 N_A_575_87#_c_610_n N_A_1374_368#_c_1427_n 0.0015259f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_548 N_A_575_87#_c_610_n N_A_1374_368#_c_1411_n 0.00629485f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_549 N_A_575_87#_c_610_n N_A_1374_368#_c_1412_n 0.0400993f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_550 N_A_575_87#_c_610_n N_A_1374_368#_c_1430_n 0.00208407f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_551 N_A_575_87#_c_610_n N_A_1374_368#_c_1414_n 0.030391f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_552 N_A_575_87#_c_610_n N_A_1374_368#_c_1415_n 0.00899734f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_553 N_A_575_87#_c_610_n N_A_2013_71#_c_1593_n 0.00298149f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_554 N_A_575_87#_c_610_n N_A_2013_71#_c_1594_n 0.00463613f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_555 N_A_575_87#_c_610_n N_A_2013_71#_c_1595_n 0.0126745f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_556 N_A_575_87#_c_610_n N_A_2013_71#_c_1597_n 0.0112107f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_557 N_A_575_87#_c_610_n N_A_2013_71#_c_1609_n 0.0117248f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_558 N_A_575_87#_c_610_n N_A_2013_71#_c_1599_n 0.0215524f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_559 N_A_575_87#_c_610_n N_A_2013_71#_c_1600_n 0.00903406f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_560 N_A_575_87#_c_610_n N_A_2013_71#_c_1601_n 0.0240966f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_561 N_A_575_87#_c_610_n N_A_2013_71#_c_1602_n 0.00849763f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_562 N_A_575_87#_c_610_n N_A_2013_71#_c_1603_n 0.00853542f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_563 N_A_575_87#_c_610_n N_A_1784_97#_c_1706_n 0.00373529f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_564 N_A_575_87#_c_610_n N_A_1784_97#_c_1708_n 0.0141202f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_565 N_A_575_87#_c_610_n N_A_1784_97#_c_1710_n 0.0600244f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_566 N_A_575_87#_c_610_n N_A_1784_97#_c_1711_n 0.00882231f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_567 N_A_575_87#_c_610_n N_A_1784_97#_c_1714_n 0.0224528f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_568 N_A_575_87#_c_617_n N_A_2489_74#_c_1802_n 0.0121797f $X=13.705 $Y=2.465
+ $X2=0 $Y2=0
cc_569 N_A_575_87#_c_601_n N_A_2489_74#_c_1802_n 0.0163791f $X=13.84 $Y=2.05
+ $X2=0 $Y2=0
cc_570 N_A_575_87#_c_621_n N_A_2489_74#_c_1802_n 0.0185932f $X=14.475 $Y=2.217
+ $X2=0 $Y2=0
cc_571 N_A_575_87#_c_604_n N_A_2489_74#_c_1802_n 0.0113716f $X=14.655 $Y=2.49
+ $X2=0 $Y2=0
cc_572 N_A_575_87#_c_623_n N_A_2489_74#_c_1802_n 0.00776817f $X=14.64 $Y=2.815
+ $X2=0 $Y2=0
cc_573 N_A_575_87#_c_599_n N_A_2489_74#_M1014_g 0.00727204f $X=13.765 $Y=0.94
+ $X2=0 $Y2=0
cc_574 N_A_575_87#_c_605_n N_A_2489_74#_M1014_g 0.00834476f $X=14.67 $Y=0.515
+ $X2=0 $Y2=0
cc_575 N_A_575_87#_c_606_n N_A_2489_74#_M1014_g 0.00600966f $X=14.75 $Y=1.55
+ $X2=0 $Y2=0
cc_576 N_A_575_87#_c_608_n N_A_2489_74#_M1014_g 0.00278814f $X=14.67 $Y=1.13
+ $X2=0 $Y2=0
cc_577 N_A_575_87#_c_604_n N_A_2489_74#_c_1792_n 0.0305492f $X=14.655 $Y=2.49
+ $X2=0 $Y2=0
cc_578 N_A_575_87#_c_606_n N_A_2489_74#_c_1792_n 0.0185398f $X=14.75 $Y=1.55
+ $X2=0 $Y2=0
cc_579 N_A_575_87#_c_727_p N_A_2489_74#_c_1792_n 0.00169922f $X=15.995 $Y=2.405
+ $X2=0 $Y2=0
cc_580 N_A_575_87#_c_608_n N_A_2489_74#_c_1792_n 0.00135743f $X=14.67 $Y=1.13
+ $X2=0 $Y2=0
cc_581 N_A_575_87#_c_610_n N_A_2489_74#_c_1792_n 0.00296264f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_582 N_A_575_87#_c_611_n N_A_2489_74#_c_1792_n 0.00679929f $X=15.12 $Y=1.665
+ $X2=0 $Y2=0
cc_583 N_A_575_87#_c_601_n N_A_2489_74#_c_1793_n 0.0216215f $X=13.84 $Y=2.05
+ $X2=0 $Y2=0
cc_584 N_A_575_87#_c_621_n N_A_2489_74#_c_1793_n 0.00194123f $X=14.475 $Y=2.217
+ $X2=0 $Y2=0
cc_585 N_A_575_87#_c_604_n N_A_2489_74#_c_1793_n 0.00925467f $X=14.655 $Y=2.49
+ $X2=0 $Y2=0
cc_586 N_A_575_87#_c_610_n N_A_2489_74#_c_1793_n 0.00702919f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_587 N_A_575_87#_c_604_n N_A_2489_74#_c_1804_n 0.0161488f $X=14.655 $Y=2.49
+ $X2=0 $Y2=0
cc_588 N_A_575_87#_c_623_n N_A_2489_74#_c_1804_n 0.00410525f $X=14.64 $Y=2.815
+ $X2=0 $Y2=0
cc_589 N_A_575_87#_c_727_p N_A_2489_74#_c_1804_n 0.0180339f $X=15.995 $Y=2.405
+ $X2=0 $Y2=0
cc_590 N_A_575_87#_c_611_n N_A_2489_74#_c_1804_n 3.64599e-19 $X=15.12 $Y=1.665
+ $X2=0 $Y2=0
cc_591 N_A_575_87#_c_605_n N_A_2489_74#_M1032_g 0.00393219f $X=14.67 $Y=0.515
+ $X2=0 $Y2=0
cc_592 N_A_575_87#_M1027_g N_A_2489_74#_M1043_g 0.0151259f $X=16.305 $Y=0.74
+ $X2=0 $Y2=0
cc_593 N_A_575_87#_c_619_n N_A_2489_74#_c_1805_n 0.0331706f $X=16.325 $Y=1.765
+ $X2=0 $Y2=0
cc_594 N_A_575_87#_c_727_p N_A_2489_74#_c_1805_n 0.0153666f $X=15.995 $Y=2.405
+ $X2=0 $Y2=0
cc_595 N_A_575_87#_c_607_n N_A_2489_74#_c_1805_n 0.00274426f $X=16.09 $Y=2.32
+ $X2=0 $Y2=0
cc_596 N_A_575_87#_c_604_n N_A_2489_74#_c_1796_n 0.00303238f $X=14.655 $Y=2.49
+ $X2=0 $Y2=0
cc_597 N_A_575_87#_c_727_p N_A_2489_74#_c_1796_n 6.08229e-19 $X=15.995 $Y=2.405
+ $X2=0 $Y2=0
cc_598 N_A_575_87#_c_607_n N_A_2489_74#_c_1796_n 9.72868e-19 $X=16.09 $Y=2.32
+ $X2=0 $Y2=0
cc_599 N_A_575_87#_c_609_n N_A_2489_74#_c_1796_n 0.00326544f $X=16.395 $Y=1.465
+ $X2=0 $Y2=0
cc_600 N_A_575_87#_c_611_n N_A_2489_74#_c_1796_n 0.00397573f $X=15.12 $Y=1.665
+ $X2=0 $Y2=0
cc_601 N_A_575_87#_c_614_n N_A_2489_74#_c_1796_n 0.0211137f $X=16.735 $Y=1.532
+ $X2=0 $Y2=0
cc_602 N_A_575_87#_c_598_n N_A_2489_74#_c_1798_n 0.00739677f $X=13.27 $Y=0.865
+ $X2=0 $Y2=0
cc_603 N_A_575_87#_c_599_n N_A_2489_74#_c_1798_n 0.0200523f $X=13.765 $Y=0.94
+ $X2=0 $Y2=0
cc_604 N_A_575_87#_c_600_n N_A_2489_74#_c_1798_n 0.00284537f $X=13.345 $Y=0.94
+ $X2=0 $Y2=0
cc_605 N_A_575_87#_c_617_n N_A_2489_74#_c_1807_n 0.0012434f $X=13.705 $Y=2.465
+ $X2=0 $Y2=0
cc_606 N_A_575_87#_c_601_n N_A_2489_74#_c_1807_n 8.72783e-19 $X=13.84 $Y=2.05
+ $X2=0 $Y2=0
cc_607 N_A_575_87#_c_621_n N_A_2489_74#_c_1807_n 0.0174688f $X=14.475 $Y=2.217
+ $X2=0 $Y2=0
cc_608 N_A_575_87#_c_617_n N_A_2489_74#_c_1808_n 0.00275459f $X=13.705 $Y=2.465
+ $X2=0 $Y2=0
cc_609 N_A_575_87#_c_601_n N_A_2489_74#_c_1808_n 3.91756e-19 $X=13.84 $Y=2.05
+ $X2=0 $Y2=0
cc_610 N_A_575_87#_c_621_n N_A_2489_74#_c_1808_n 0.00772483f $X=14.475 $Y=2.217
+ $X2=0 $Y2=0
cc_611 N_A_575_87#_c_610_n N_A_2489_74#_c_1808_n 0.0191403f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_612 N_A_575_87#_c_610_n N_A_2489_74#_c_1809_n 0.0108527f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_613 N_A_575_87#_c_599_n N_A_2489_74#_c_1799_n 0.00639798f $X=13.765 $Y=0.94
+ $X2=0 $Y2=0
cc_614 N_A_575_87#_c_601_n N_A_2489_74#_c_1799_n 0.00974521f $X=13.84 $Y=2.05
+ $X2=0 $Y2=0
cc_615 N_A_575_87#_c_608_n N_A_2489_74#_c_1799_n 2.36907e-19 $X=14.67 $Y=1.13
+ $X2=0 $Y2=0
cc_616 N_A_575_87#_c_617_n N_A_2489_74#_c_1800_n 0.00189071f $X=13.705 $Y=2.465
+ $X2=0 $Y2=0
cc_617 N_A_575_87#_c_601_n N_A_2489_74#_c_1800_n 0.0154484f $X=13.84 $Y=2.05
+ $X2=0 $Y2=0
cc_618 N_A_575_87#_c_621_n N_A_2489_74#_c_1800_n 0.0128991f $X=14.475 $Y=2.217
+ $X2=0 $Y2=0
cc_619 N_A_575_87#_c_604_n N_A_2489_74#_c_1800_n 0.00223915f $X=14.655 $Y=2.49
+ $X2=0 $Y2=0
cc_620 N_A_575_87#_c_610_n N_A_2489_74#_c_1800_n 0.0191046f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_621 N_A_575_87#_c_601_n N_A_2489_74#_c_1801_n 0.00891743f $X=13.84 $Y=2.05
+ $X2=0 $Y2=0
cc_622 N_A_575_87#_c_621_n N_A_2489_74#_c_1801_n 0.0134213f $X=14.475 $Y=2.217
+ $X2=0 $Y2=0
cc_623 N_A_575_87#_c_604_n N_A_2489_74#_c_1801_n 0.00718983f $X=14.655 $Y=2.49
+ $X2=0 $Y2=0
cc_624 N_A_575_87#_c_606_n N_A_2489_74#_c_1801_n 0.0188124f $X=14.75 $Y=1.55
+ $X2=0 $Y2=0
cc_625 N_A_575_87#_c_610_n N_A_2489_74#_c_1801_n 0.0309319f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_626 N_A_575_87#_c_617_n N_A_2489_74#_c_1811_n 0.00186889f $X=13.705 $Y=2.465
+ $X2=0 $Y2=0
cc_627 N_A_575_87#_c_616_n N_A_32_74#_c_1957_n 0.0130721f $X=3.205 $Y=2.235
+ $X2=0 $Y2=0
cc_628 N_A_575_87#_c_633_n N_A_32_74#_c_1957_n 0.00295921f $X=3.265 $Y=1.665
+ $X2=0 $Y2=0
cc_629 N_A_575_87#_c_612_n N_A_32_74#_c_1957_n 0.0102375f $X=3.04 $Y=1.68 $X2=0
+ $Y2=0
cc_630 N_A_575_87#_c_613_n N_A_32_74#_c_1957_n 0.00427623f $X=3.205 $Y=1.68
+ $X2=0 $Y2=0
cc_631 N_A_575_87#_M1006_g N_A_32_74#_c_1947_n 0.0139535f $X=2.95 $Y=0.775 $X2=0
+ $Y2=0
cc_632 N_A_575_87#_M1006_g N_A_32_74#_c_1948_n 0.00479218f $X=2.95 $Y=0.775
+ $X2=0 $Y2=0
cc_633 N_A_575_87#_c_616_n N_A_32_74#_c_1948_n 0.0012384f $X=3.205 $Y=2.235
+ $X2=0 $Y2=0
cc_634 N_A_575_87#_c_610_n N_A_32_74#_c_1948_n 0.0165546f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_635 N_A_575_87#_c_633_n N_A_32_74#_c_1948_n 0.00240104f $X=3.265 $Y=1.665
+ $X2=0 $Y2=0
cc_636 N_A_575_87#_c_612_n N_A_32_74#_c_1948_n 0.0226176f $X=3.04 $Y=1.68 $X2=0
+ $Y2=0
cc_637 N_A_575_87#_c_613_n N_A_32_74#_c_1948_n 0.0160465f $X=3.205 $Y=1.68 $X2=0
+ $Y2=0
cc_638 N_A_575_87#_M1006_g N_A_32_74#_c_1950_n 0.00700496f $X=2.95 $Y=0.775
+ $X2=0 $Y2=0
cc_639 N_A_575_87#_c_610_n N_A_32_74#_c_1950_n 0.00516988f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_640 N_A_575_87#_c_633_n N_A_32_74#_c_1950_n 0.00394327f $X=3.265 $Y=1.665
+ $X2=0 $Y2=0
cc_641 N_A_575_87#_c_612_n N_A_32_74#_c_1950_n 0.0139741f $X=3.04 $Y=1.68 $X2=0
+ $Y2=0
cc_642 N_A_575_87#_c_613_n N_A_32_74#_c_1950_n 0.00812585f $X=3.205 $Y=1.68
+ $X2=0 $Y2=0
cc_643 N_A_575_87#_c_616_n N_A_32_74#_c_1961_n 0.0102922f $X=3.205 $Y=2.235
+ $X2=0 $Y2=0
cc_644 N_A_575_87#_c_610_n N_A_32_74#_c_1961_n 0.00385085f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_645 N_A_575_87#_c_621_n N_VPWR_M1022_d 0.00684327f $X=14.475 $Y=2.217 $X2=0
+ $Y2=0
cc_646 N_A_575_87#_c_604_n N_VPWR_M1005_s 0.0125424f $X=14.655 $Y=2.49 $X2=0
+ $Y2=0
cc_647 N_A_575_87#_c_727_p N_VPWR_M1005_s 0.00136304f $X=15.995 $Y=2.405 $X2=0
+ $Y2=0
cc_648 N_A_575_87#_c_727_p N_VPWR_M1016_s 0.00410137f $X=15.995 $Y=2.405 $X2=0
+ $Y2=0
cc_649 N_A_575_87#_c_607_n N_VPWR_M1016_s 0.00803013f $X=16.09 $Y=2.32 $X2=0
+ $Y2=0
cc_650 N_A_575_87#_c_616_n N_VPWR_c_2068_n 0.00149083f $X=3.205 $Y=2.235 $X2=0
+ $Y2=0
cc_651 N_A_575_87#_c_617_n N_VPWR_c_2074_n 0.0184408f $X=13.705 $Y=2.465 $X2=0
+ $Y2=0
cc_652 N_A_575_87#_c_621_n N_VPWR_c_2074_n 0.0292563f $X=14.475 $Y=2.217 $X2=0
+ $Y2=0
cc_653 N_A_575_87#_c_623_n N_VPWR_c_2074_n 0.0133999f $X=14.64 $Y=2.815 $X2=0
+ $Y2=0
cc_654 N_A_575_87#_c_604_n N_VPWR_c_2075_n 0.0175754f $X=14.655 $Y=2.49 $X2=0
+ $Y2=0
cc_655 N_A_575_87#_c_623_n N_VPWR_c_2075_n 0.0239305f $X=14.64 $Y=2.815 $X2=0
+ $Y2=0
cc_656 N_A_575_87#_c_727_p N_VPWR_c_2075_n 0.00558175f $X=15.995 $Y=2.405 $X2=0
+ $Y2=0
cc_657 N_A_575_87#_c_619_n N_VPWR_c_2076_n 0.00725426f $X=16.325 $Y=1.765 $X2=0
+ $Y2=0
cc_658 N_A_575_87#_c_620_n N_VPWR_c_2076_n 3.29061e-19 $X=16.775 $Y=1.765 $X2=0
+ $Y2=0
cc_659 N_A_575_87#_c_727_p N_VPWR_c_2076_n 0.0166202f $X=15.995 $Y=2.405 $X2=0
+ $Y2=0
cc_660 N_A_575_87#_c_619_n N_VPWR_c_2078_n 4.63588e-19 $X=16.325 $Y=1.765 $X2=0
+ $Y2=0
cc_661 N_A_575_87#_c_620_n N_VPWR_c_2078_n 0.0155262f $X=16.775 $Y=1.765 $X2=0
+ $Y2=0
cc_662 N_A_575_87#_c_616_n N_VPWR_c_2085_n 0.0055545f $X=3.205 $Y=2.235 $X2=0
+ $Y2=0
cc_663 N_A_575_87#_c_617_n N_VPWR_c_2088_n 0.00413917f $X=13.705 $Y=2.465 $X2=0
+ $Y2=0
cc_664 N_A_575_87#_c_623_n N_VPWR_c_2089_n 0.0159324f $X=14.64 $Y=2.815 $X2=0
+ $Y2=0
cc_665 N_A_575_87#_c_619_n N_VPWR_c_2091_n 0.00413917f $X=16.325 $Y=1.765 $X2=0
+ $Y2=0
cc_666 N_A_575_87#_c_620_n N_VPWR_c_2091_n 0.00413917f $X=16.775 $Y=1.765 $X2=0
+ $Y2=0
cc_667 N_A_575_87#_c_616_n N_VPWR_c_2066_n 0.00542671f $X=3.205 $Y=2.235 $X2=0
+ $Y2=0
cc_668 N_A_575_87#_c_617_n N_VPWR_c_2066_n 0.00852225f $X=13.705 $Y=2.465 $X2=0
+ $Y2=0
cc_669 N_A_575_87#_c_619_n N_VPWR_c_2066_n 0.00817726f $X=16.325 $Y=1.765 $X2=0
+ $Y2=0
cc_670 N_A_575_87#_c_620_n N_VPWR_c_2066_n 0.00817726f $X=16.775 $Y=1.765 $X2=0
+ $Y2=0
cc_671 N_A_575_87#_c_604_n N_VPWR_c_2066_n 0.00864971f $X=14.655 $Y=2.49 $X2=0
+ $Y2=0
cc_672 N_A_575_87#_c_623_n N_VPWR_c_2066_n 0.0131546f $X=14.64 $Y=2.815 $X2=0
+ $Y2=0
cc_673 N_A_575_87#_c_727_p N_VPWR_c_2066_n 0.0190963f $X=15.995 $Y=2.405 $X2=0
+ $Y2=0
cc_674 N_A_575_87#_c_610_n N_A_691_113#_c_2274_n 0.00288899f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_675 N_A_575_87#_c_616_n N_A_691_113#_c_2286_n 5.12161e-19 $X=3.205 $Y=2.235
+ $X2=0 $Y2=0
cc_676 N_A_575_87#_c_610_n N_A_691_113#_c_2276_n 0.00532122f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_677 N_A_575_87#_c_610_n N_A_691_113#_c_2277_n 0.00111174f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_678 N_A_575_87#_c_610_n N_A_691_113#_c_2267_n 0.0202067f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_679 N_A_575_87#_c_610_n N_A_691_113#_c_2279_n 0.0197782f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_680 N_A_575_87#_c_610_n N_A_691_113#_c_2280_n 0.0076514f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_681 N_A_575_87#_c_610_n N_A_691_113#_c_2281_n 0.013888f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_682 N_A_575_87#_c_610_n N_A_691_113#_c_2268_n 0.0347249f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_683 N_A_575_87#_c_610_n N_A_691_113#_c_2269_n 0.00439964f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_684 N_A_575_87#_c_610_n N_A_691_113#_c_2295_n 0.00276274f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_685 N_A_575_87#_c_610_n N_A_691_113#_c_2271_n 0.00579027f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_686 N_A_575_87#_M1006_g N_A_691_113#_c_2272_n 5.8879e-19 $X=2.95 $Y=0.775
+ $X2=0 $Y2=0
cc_687 N_A_575_87#_c_610_n N_A_691_113#_c_2272_n 0.0186936f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_688 N_A_575_87#_c_610_n N_A_691_113#_c_2273_n 0.00878755f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_689 N_A_575_87#_c_727_p N_Q_M1005_d 0.00558496f $X=15.995 $Y=2.405 $X2=0
+ $Y2=0
cc_690 N_A_575_87#_M1027_g Q 0.0010619f $X=16.305 $Y=0.74 $X2=0 $Y2=0
cc_691 N_A_575_87#_c_604_n Q 0.0328167f $X=14.655 $Y=2.49 $X2=0 $Y2=0
cc_692 N_A_575_87#_c_606_n Q 0.0104168f $X=14.75 $Y=1.55 $X2=0 $Y2=0
cc_693 N_A_575_87#_c_727_p Q 0.0179431f $X=15.995 $Y=2.405 $X2=0 $Y2=0
cc_694 N_A_575_87#_c_607_n Q 0.0271809f $X=16.09 $Y=2.32 $X2=0 $Y2=0
cc_695 N_A_575_87#_c_609_n Q 0.0275006f $X=16.395 $Y=1.465 $X2=0 $Y2=0
cc_696 N_A_575_87#_c_611_n Q 0.00675851f $X=15.12 $Y=1.665 $X2=0 $Y2=0
cc_697 N_A_575_87#_c_614_n Q 2.32349e-19 $X=16.735 $Y=1.532 $X2=0 $Y2=0
cc_698 N_A_575_87#_M1027_g N_Q_N_c_2476_n 0.00237533f $X=16.305 $Y=0.74 $X2=0
+ $Y2=0
cc_699 N_A_575_87#_M1041_g N_Q_N_c_2476_n 0.0131327f $X=16.735 $Y=0.74 $X2=0
+ $Y2=0
cc_700 N_A_575_87#_c_609_n N_Q_N_c_2476_n 0.0115705f $X=16.395 $Y=1.465 $X2=0
+ $Y2=0
cc_701 N_A_575_87#_c_614_n N_Q_N_c_2476_n 0.002804f $X=16.735 $Y=1.532 $X2=0
+ $Y2=0
cc_702 N_A_575_87#_M1027_g N_Q_N_c_2477_n 9.68429e-19 $X=16.305 $Y=0.74 $X2=0
+ $Y2=0
cc_703 N_A_575_87#_c_619_n N_Q_N_c_2477_n 3.4717e-19 $X=16.325 $Y=1.765 $X2=0
+ $Y2=0
cc_704 N_A_575_87#_M1041_g N_Q_N_c_2477_n 0.00816363f $X=16.735 $Y=0.74 $X2=0
+ $Y2=0
cc_705 N_A_575_87#_c_620_n N_Q_N_c_2477_n 0.0150088f $X=16.775 $Y=1.765 $X2=0
+ $Y2=0
cc_706 N_A_575_87#_c_607_n N_Q_N_c_2477_n 0.0115912f $X=16.09 $Y=2.32 $X2=0
+ $Y2=0
cc_707 N_A_575_87#_c_609_n N_Q_N_c_2477_n 0.0303602f $X=16.395 $Y=1.465 $X2=0
+ $Y2=0
cc_708 N_A_575_87#_c_614_n N_Q_N_c_2477_n 0.0311749f $X=16.735 $Y=1.532 $X2=0
+ $Y2=0
cc_709 N_A_575_87#_M1027_g Q_N 0.00756419f $X=16.305 $Y=0.74 $X2=0 $Y2=0
cc_710 N_A_575_87#_M1041_g Q_N 0.013384f $X=16.735 $Y=0.74 $X2=0 $Y2=0
cc_711 N_A_575_87#_c_619_n Q_N 0.00402046f $X=16.325 $Y=1.765 $X2=0 $Y2=0
cc_712 N_A_575_87#_c_620_n Q_N 0.00402046f $X=16.775 $Y=1.765 $X2=0 $Y2=0
cc_713 N_A_575_87#_M1006_g N_VGND_c_2510_n 0.0018473f $X=2.95 $Y=0.775 $X2=0
+ $Y2=0
cc_714 N_A_575_87#_c_610_n N_VGND_c_2511_n 0.00383642f $X=14.975 $Y=1.665 $X2=0
+ $Y2=0
cc_715 N_A_575_87#_c_610_n N_VGND_c_2513_n 0.00319228f $X=14.975 $Y=1.665 $X2=0
+ $Y2=0
cc_716 N_A_575_87#_c_599_n N_VGND_c_2516_n 0.00216966f $X=13.765 $Y=0.94 $X2=0
+ $Y2=0
cc_717 N_A_575_87#_c_598_n N_VGND_c_2517_n 0.0105517f $X=13.27 $Y=0.865 $X2=0
+ $Y2=0
cc_718 N_A_575_87#_c_599_n N_VGND_c_2517_n 0.00310568f $X=13.765 $Y=0.94 $X2=0
+ $Y2=0
cc_719 N_A_575_87#_c_599_n N_VGND_c_2518_n 0.00246324f $X=13.765 $Y=0.94 $X2=0
+ $Y2=0
cc_720 N_A_575_87#_c_605_n N_VGND_c_2518_n 0.0198374f $X=14.67 $Y=0.515 $X2=0
+ $Y2=0
cc_721 N_A_575_87#_c_610_n N_VGND_c_2518_n 0.00126635f $X=14.975 $Y=1.665 $X2=0
+ $Y2=0
cc_722 N_A_575_87#_c_605_n N_VGND_c_2519_n 0.0145639f $X=14.67 $Y=0.515 $X2=0
+ $Y2=0
cc_723 N_A_575_87#_c_604_n N_VGND_c_2520_n 0.00440301f $X=14.655 $Y=2.49 $X2=0
+ $Y2=0
cc_724 N_A_575_87#_c_605_n N_VGND_c_2520_n 0.0514703f $X=14.67 $Y=0.515 $X2=0
+ $Y2=0
cc_725 N_A_575_87#_c_611_n N_VGND_c_2520_n 0.00254943f $X=15.12 $Y=1.665 $X2=0
+ $Y2=0
cc_726 N_A_575_87#_M1027_g N_VGND_c_2522_n 0.00315608f $X=16.305 $Y=0.74 $X2=0
+ $Y2=0
cc_727 N_A_575_87#_c_609_n N_VGND_c_2522_n 0.0148775f $X=16.395 $Y=1.465 $X2=0
+ $Y2=0
cc_728 N_A_575_87#_M1041_g N_VGND_c_2524_n 0.00611725f $X=16.735 $Y=0.74 $X2=0
+ $Y2=0
cc_729 N_A_575_87#_c_598_n N_VGND_c_2529_n 0.00383152f $X=13.27 $Y=0.865 $X2=0
+ $Y2=0
cc_730 N_A_575_87#_M1006_g N_VGND_c_2531_n 0.00430863f $X=2.95 $Y=0.775 $X2=0
+ $Y2=0
cc_731 N_A_575_87#_M1027_g N_VGND_c_2535_n 0.00434272f $X=16.305 $Y=0.74 $X2=0
+ $Y2=0
cc_732 N_A_575_87#_M1041_g N_VGND_c_2535_n 0.00434272f $X=16.735 $Y=0.74 $X2=0
+ $Y2=0
cc_733 N_A_575_87#_c_605_n N_VGND_c_2541_n 0.0103109f $X=14.67 $Y=0.515 $X2=0
+ $Y2=0
cc_734 N_A_575_87#_M1006_g N_VGND_c_2544_n 0.00486331f $X=2.95 $Y=0.775 $X2=0
+ $Y2=0
cc_735 N_A_575_87#_c_598_n N_VGND_c_2544_n 0.00367447f $X=13.27 $Y=0.865 $X2=0
+ $Y2=0
cc_736 N_A_575_87#_M1027_g N_VGND_c_2544_n 0.00820382f $X=16.305 $Y=0.74 $X2=0
+ $Y2=0
cc_737 N_A_575_87#_M1041_g N_VGND_c_2544_n 0.00823877f $X=16.735 $Y=0.74 $X2=0
+ $Y2=0
cc_738 N_A_575_87#_c_605_n N_VGND_c_2544_n 0.0119984f $X=14.67 $Y=0.515 $X2=0
+ $Y2=0
cc_739 N_A_661_87#_c_897_n N_SCD_c_998_n 0.0223471f $X=5.915 $Y=1.865 $X2=0
+ $Y2=0
cc_740 N_A_661_87#_c_899_n N_SCD_c_998_n 0.0127814f $X=5.805 $Y=1.765 $X2=0
+ $Y2=0
cc_741 N_A_661_87#_c_903_n N_SCD_c_998_n 0.00130006f $X=5.97 $Y=1.58 $X2=0 $Y2=0
cc_742 N_A_661_87#_c_896_n N_SCD_c_1003_n 0.0386525f $X=5.785 $Y=2.19 $X2=0
+ $Y2=0
cc_743 N_A_661_87#_c_899_n SCD 0.0330694f $X=5.805 $Y=1.765 $X2=0 $Y2=0
cc_744 N_A_661_87#_c_903_n SCD 0.00650547f $X=5.97 $Y=1.58 $X2=0 $Y2=0
cc_745 N_A_661_87#_c_895_n SCD 8.85081e-19 $X=5.97 $Y=1.58 $X2=0 $Y2=0
cc_746 N_A_661_87#_c_899_n N_SCD_c_1001_n 0.00329296f $X=5.805 $Y=1.765 $X2=0
+ $Y2=0
cc_747 N_A_661_87#_c_903_n N_SCD_c_1001_n 0.00122864f $X=5.97 $Y=1.58 $X2=0
+ $Y2=0
cc_748 N_A_661_87#_c_895_n N_SCD_c_1001_n 0.0223471f $X=5.97 $Y=1.58 $X2=0 $Y2=0
cc_749 N_A_661_87#_c_898_n N_SCE_c_1051_n 3.10849e-19 $X=4.22 $Y=2.245 $X2=-0.19
+ $Y2=-0.245
cc_750 N_A_661_87#_c_902_n N_SCE_c_1051_n 0.00105023f $X=4.44 $Y=2.49 $X2=-0.19
+ $Y2=-0.245
cc_751 N_A_661_87#_c_902_n N_SCE_c_1052_n 0.00224682f $X=4.44 $Y=2.49 $X2=0
+ $Y2=0
cc_752 N_A_661_87#_c_898_n N_SCE_c_1044_n 0.00416364f $X=4.22 $Y=2.245 $X2=0
+ $Y2=0
cc_753 N_A_661_87#_c_899_n N_SCE_c_1044_n 0.0152143f $X=5.805 $Y=1.765 $X2=0
+ $Y2=0
cc_754 N_A_661_87#_c_900_n N_SCE_c_1044_n 0.00200108f $X=4.18 $Y=1.765 $X2=0
+ $Y2=0
cc_755 N_A_661_87#_c_894_n N_SCE_c_1044_n 0.0241622f $X=4.18 $Y=1.89 $X2=0 $Y2=0
cc_756 N_A_661_87#_c_898_n N_SCE_M1045_g 0.00163272f $X=4.22 $Y=2.245 $X2=0
+ $Y2=0
cc_757 N_A_661_87#_c_902_n N_SCE_M1045_g 0.00358656f $X=4.44 $Y=2.49 $X2=0 $Y2=0
cc_758 N_A_661_87#_c_891_n N_SCE_M1039_g 8.75597e-19 $X=4.18 $Y=1.01 $X2=0 $Y2=0
cc_759 N_A_661_87#_c_907_n N_SCE_M1039_g 8.91698e-19 $X=4.18 $Y=1.21 $X2=0 $Y2=0
cc_760 N_A_661_87#_c_892_n N_SCE_M1039_g 0.00549146f $X=4.625 $Y=0.805 $X2=0
+ $Y2=0
cc_761 N_A_661_87#_c_893_n N_SCE_M1039_g 0.0176733f $X=4.18 $Y=0.53 $X2=0 $Y2=0
cc_762 N_A_661_87#_c_899_n N_SCE_M1036_g 7.90301e-19 $X=5.805 $Y=1.765 $X2=0
+ $Y2=0
cc_763 N_A_661_87#_c_895_n N_SCE_M1036_g 0.0100355f $X=5.97 $Y=1.58 $X2=0 $Y2=0
cc_764 N_A_661_87#_c_890_n N_SCE_c_1049_n 0.0241622f $X=4.18 $Y=1.135 $X2=0
+ $Y2=0
cc_765 N_A_661_87#_c_907_n N_SCE_c_1049_n 9.78573e-19 $X=4.18 $Y=1.21 $X2=0
+ $Y2=0
cc_766 N_A_661_87#_c_892_n N_SCE_c_1049_n 0.00467945f $X=4.625 $Y=0.805 $X2=0
+ $Y2=0
cc_767 N_A_661_87#_c_899_n N_SCE_c_1049_n 0.00388395f $X=5.805 $Y=1.765 $X2=0
+ $Y2=0
cc_768 N_A_661_87#_c_890_n N_SCE_c_1050_n 0.00222389f $X=4.18 $Y=1.135 $X2=0
+ $Y2=0
cc_769 N_A_661_87#_c_907_n N_SCE_c_1050_n 0.0261395f $X=4.18 $Y=1.21 $X2=0 $Y2=0
cc_770 N_A_661_87#_c_892_n N_SCE_c_1050_n 0.0223339f $X=4.625 $Y=0.805 $X2=0
+ $Y2=0
cc_771 N_A_661_87#_c_899_n N_SCE_c_1050_n 0.0283146f $X=5.805 $Y=1.765 $X2=0
+ $Y2=0
cc_772 N_A_661_87#_c_895_n N_CLK_c_1127_n 0.0100232f $X=5.97 $Y=1.58 $X2=-0.19
+ $Y2=-0.245
cc_773 N_A_661_87#_c_887_n N_A_32_74#_c_1947_n 0.00745701f $X=3.38 $Y=1.06 $X2=0
+ $Y2=0
cc_774 N_A_661_87#_c_889_n N_A_32_74#_c_1947_n 0.00424876f $X=3.455 $Y=1.135
+ $X2=0 $Y2=0
cc_775 N_A_661_87#_c_889_n N_A_32_74#_c_1948_n 9.15581e-19 $X=3.455 $Y=1.135
+ $X2=0 $Y2=0
cc_776 N_A_661_87#_c_888_n N_A_32_74#_c_1950_n 0.00486125f $X=4.015 $Y=1.135
+ $X2=0 $Y2=0
cc_777 N_A_661_87#_c_889_n N_A_32_74#_c_1950_n 0.00908768f $X=3.455 $Y=1.135
+ $X2=0 $Y2=0
cc_778 N_A_661_87#_c_896_n N_VPWR_c_2069_n 0.00148326f $X=5.785 $Y=2.19 $X2=0
+ $Y2=0
cc_779 N_A_661_87#_c_896_n N_VPWR_c_2070_n 0.00280498f $X=5.785 $Y=2.19 $X2=0
+ $Y2=0
cc_780 N_A_661_87#_c_896_n N_VPWR_c_2079_n 0.00522998f $X=5.785 $Y=2.19 $X2=0
+ $Y2=0
cc_781 N_A_661_87#_c_896_n N_VPWR_c_2066_n 0.00528353f $X=5.785 $Y=2.19 $X2=0
+ $Y2=0
cc_782 N_A_661_87#_c_902_n N_A_691_113#_c_2274_n 0.0362007f $X=4.44 $Y=2.49
+ $X2=0 $Y2=0
cc_783 N_A_661_87#_c_902_n N_A_691_113#_c_2275_n 0.0295498f $X=4.44 $Y=2.49
+ $X2=0 $Y2=0
cc_784 N_A_661_87#_c_902_n N_A_691_113#_c_2302_n 0.0232577f $X=4.44 $Y=2.49
+ $X2=0 $Y2=0
cc_785 N_A_661_87#_c_896_n N_A_691_113#_c_2276_n 0.0122978f $X=5.785 $Y=2.19
+ $X2=0 $Y2=0
cc_786 N_A_661_87#_c_897_n N_A_691_113#_c_2276_n 4.93938e-19 $X=5.915 $Y=1.865
+ $X2=0 $Y2=0
cc_787 N_A_661_87#_c_899_n N_A_691_113#_c_2276_n 0.0309344f $X=5.805 $Y=1.765
+ $X2=0 $Y2=0
cc_788 N_A_661_87#_c_903_n N_A_691_113#_c_2276_n 0.00284364f $X=5.97 $Y=1.58
+ $X2=0 $Y2=0
cc_789 N_A_661_87#_c_899_n N_A_691_113#_c_2277_n 0.00604348f $X=5.805 $Y=1.765
+ $X2=0 $Y2=0
cc_790 N_A_661_87#_c_902_n N_A_691_113#_c_2277_n 0.0142675f $X=4.44 $Y=2.49
+ $X2=0 $Y2=0
cc_791 N_A_661_87#_c_896_n N_A_691_113#_c_2267_n 0.00163973f $X=5.785 $Y=2.19
+ $X2=0 $Y2=0
cc_792 N_A_661_87#_c_897_n N_A_691_113#_c_2267_n 0.00278924f $X=5.915 $Y=1.865
+ $X2=0 $Y2=0
cc_793 N_A_661_87#_c_903_n N_A_691_113#_c_2267_n 0.0481738f $X=5.97 $Y=1.58
+ $X2=0 $Y2=0
cc_794 N_A_661_87#_c_895_n N_A_691_113#_c_2267_n 0.00643452f $X=5.97 $Y=1.58
+ $X2=0 $Y2=0
cc_795 N_A_661_87#_c_896_n N_A_691_113#_c_2280_n 0.0099462f $X=5.785 $Y=2.19
+ $X2=0 $Y2=0
cc_796 N_A_661_87#_c_897_n N_A_691_113#_c_2280_n 0.00247726f $X=5.915 $Y=1.865
+ $X2=0 $Y2=0
cc_797 N_A_661_87#_c_903_n N_A_691_113#_c_2280_n 0.0247389f $X=5.97 $Y=1.58
+ $X2=0 $Y2=0
cc_798 N_A_661_87#_c_887_n N_A_691_113#_c_2271_n 0.00364479f $X=3.38 $Y=1.06
+ $X2=0 $Y2=0
cc_799 N_A_661_87#_c_888_n N_A_691_113#_c_2271_n 0.00746942f $X=4.015 $Y=1.135
+ $X2=0 $Y2=0
cc_800 N_A_661_87#_c_891_n N_A_691_113#_c_2271_n 0.0390571f $X=4.18 $Y=1.01
+ $X2=0 $Y2=0
cc_801 N_A_661_87#_c_893_n N_A_691_113#_c_2271_n 0.00543315f $X=4.18 $Y=0.53
+ $X2=0 $Y2=0
cc_802 N_A_661_87#_c_887_n N_A_691_113#_c_2272_n 4.83295e-19 $X=3.38 $Y=1.06
+ $X2=0 $Y2=0
cc_803 N_A_661_87#_c_888_n N_A_691_113#_c_2272_n 0.0150982f $X=4.015 $Y=1.135
+ $X2=0 $Y2=0
cc_804 N_A_661_87#_c_907_n N_A_691_113#_c_2272_n 0.0753924f $X=4.18 $Y=1.21
+ $X2=0 $Y2=0
cc_805 N_A_661_87#_c_898_n N_A_691_113#_c_2272_n 0.0109073f $X=4.22 $Y=2.245
+ $X2=0 $Y2=0
cc_806 N_A_661_87#_c_894_n N_A_691_113#_c_2272_n 0.013121f $X=4.18 $Y=1.89 $X2=0
+ $Y2=0
cc_807 N_A_661_87#_c_902_n N_A_691_113#_c_2272_n 0.00268195f $X=4.44 $Y=2.49
+ $X2=0 $Y2=0
cc_808 N_A_661_87#_c_903_n N_A_691_113#_c_2273_n 0.0235691f $X=5.97 $Y=1.58
+ $X2=0 $Y2=0
cc_809 N_A_661_87#_c_895_n N_A_691_113#_c_2273_n 0.00784966f $X=5.97 $Y=1.58
+ $X2=0 $Y2=0
cc_810 N_A_661_87#_c_891_n N_VGND_c_2511_n 0.00663031f $X=4.18 $Y=1.01 $X2=0
+ $Y2=0
cc_811 N_A_661_87#_c_892_n N_VGND_c_2511_n 0.0177281f $X=4.625 $Y=0.805 $X2=0
+ $Y2=0
cc_812 N_A_661_87#_c_899_n N_VGND_c_2511_n 0.00247704f $X=5.805 $Y=1.765 $X2=0
+ $Y2=0
cc_813 N_A_661_87#_c_887_n N_VGND_c_2531_n 0.00430863f $X=3.38 $Y=1.06 $X2=0
+ $Y2=0
cc_814 N_A_661_87#_c_891_n N_VGND_c_2531_n 0.00979148f $X=4.18 $Y=1.01 $X2=0
+ $Y2=0
cc_815 N_A_661_87#_c_892_n N_VGND_c_2531_n 0.00989191f $X=4.625 $Y=0.805 $X2=0
+ $Y2=0
cc_816 N_A_661_87#_c_893_n N_VGND_c_2531_n 0.0036882f $X=4.18 $Y=0.53 $X2=0
+ $Y2=0
cc_817 N_A_661_87#_c_887_n N_VGND_c_2544_n 0.00486331f $X=3.38 $Y=1.06 $X2=0
+ $Y2=0
cc_818 N_A_661_87#_c_891_n N_VGND_c_2544_n 0.00893856f $X=4.18 $Y=1.01 $X2=0
+ $Y2=0
cc_819 N_A_661_87#_c_892_n N_VGND_c_2544_n 0.0145109f $X=4.625 $Y=0.805 $X2=0
+ $Y2=0
cc_820 N_A_661_87#_c_893_n N_VGND_c_2544_n 0.00270334f $X=4.18 $Y=0.53 $X2=0
+ $Y2=0
cc_821 N_SCD_c_1003_n N_SCE_c_1052_n 9.69788e-19 $X=5.365 $Y=2.19 $X2=0 $Y2=0
cc_822 N_SCD_c_998_n N_SCE_c_1044_n 0.00902607f $X=5.365 $Y=2.1 $X2=0 $Y2=0
cc_823 N_SCD_c_1003_n N_SCE_c_1055_n 0.00902607f $X=5.365 $Y=2.19 $X2=0 $Y2=0
cc_824 N_SCD_c_1003_n N_SCE_M1045_g 0.0109972f $X=5.365 $Y=2.19 $X2=0 $Y2=0
cc_825 N_SCD_M1021_g N_SCE_M1039_g 0.013329f $X=5.38 $Y=0.835 $X2=0 $Y2=0
cc_826 N_SCD_M1021_g N_SCE_c_1046_n 0.00907339f $X=5.38 $Y=0.835 $X2=0 $Y2=0
cc_827 N_SCD_M1021_g N_SCE_M1036_g 0.0345301f $X=5.38 $Y=0.835 $X2=0 $Y2=0
cc_828 SCD N_SCE_c_1049_n 4.12687e-19 $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_829 N_SCD_c_1001_n N_SCE_c_1049_n 0.0214313f $X=5.29 $Y=1.345 $X2=0 $Y2=0
cc_830 SCD N_SCE_c_1050_n 0.0221522f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_831 N_SCD_c_1001_n N_SCE_c_1050_n 4.13447e-19 $X=5.29 $Y=1.345 $X2=0 $Y2=0
cc_832 N_SCD_c_1003_n N_VPWR_c_2069_n 0.00976838f $X=5.365 $Y=2.19 $X2=0 $Y2=0
cc_833 N_SCD_c_1003_n N_VPWR_c_2079_n 0.0048289f $X=5.365 $Y=2.19 $X2=0 $Y2=0
cc_834 N_SCD_c_1003_n N_VPWR_c_2066_n 0.0047904f $X=5.365 $Y=2.19 $X2=0 $Y2=0
cc_835 N_SCD_c_1003_n N_A_691_113#_c_2275_n 3.44487e-19 $X=5.365 $Y=2.19 $X2=0
+ $Y2=0
cc_836 N_SCD_c_1003_n N_A_691_113#_c_2302_n 0.00275933f $X=5.365 $Y=2.19 $X2=0
+ $Y2=0
cc_837 N_SCD_c_1003_n N_A_691_113#_c_2276_n 0.0175715f $X=5.365 $Y=2.19 $X2=0
+ $Y2=0
cc_838 N_SCD_M1021_g N_A_691_113#_c_2266_n 0.00156538f $X=5.38 $Y=0.835 $X2=0
+ $Y2=0
cc_839 SCD N_A_691_113#_c_2267_n 0.00535427f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_840 N_SCD_c_1003_n N_A_691_113#_c_2280_n 0.00176441f $X=5.365 $Y=2.19 $X2=0
+ $Y2=0
cc_841 N_SCD_M1021_g N_A_691_113#_c_2273_n 5.99886e-19 $X=5.38 $Y=0.835 $X2=0
+ $Y2=0
cc_842 SCD N_A_691_113#_c_2273_n 0.00671568f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_843 N_SCD_c_1001_n N_A_691_113#_c_2273_n 4.02826e-19 $X=5.29 $Y=1.345 $X2=0
+ $Y2=0
cc_844 N_SCD_M1021_g N_VGND_c_2511_n 0.0036597f $X=5.38 $Y=0.835 $X2=0 $Y2=0
cc_845 SCD N_VGND_c_2511_n 0.0114218f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_846 N_SCD_c_1001_n N_VGND_c_2511_n 0.00375077f $X=5.29 $Y=1.345 $X2=0 $Y2=0
cc_847 N_SCD_M1021_g N_VGND_c_2544_n 9.49986e-19 $X=5.38 $Y=0.835 $X2=0 $Y2=0
cc_848 N_SCE_c_1051_n N_A_32_74#_c_1948_n 8.17475e-19 $X=3.655 $Y=3.025 $X2=0
+ $Y2=0
cc_849 N_SCE_c_1052_n N_VPWR_c_2069_n 0.00310851f $X=4.585 $Y=3.1 $X2=0 $Y2=0
cc_850 N_SCE_M1045_g N_VPWR_c_2069_n 0.00119166f $X=4.675 $Y=2.585 $X2=0 $Y2=0
cc_851 N_SCE_c_1053_n N_VPWR_c_2085_n 0.0250818f $X=3.73 $Y=3.1 $X2=0 $Y2=0
cc_852 N_SCE_c_1052_n N_VPWR_c_2066_n 0.0262386f $X=4.585 $Y=3.1 $X2=0 $Y2=0
cc_853 N_SCE_c_1053_n N_VPWR_c_2066_n 0.0111009f $X=3.73 $Y=3.1 $X2=0 $Y2=0
cc_854 N_SCE_c_1051_n N_A_691_113#_c_2274_n 0.00154181f $X=3.655 $Y=3.025 $X2=0
+ $Y2=0
cc_855 N_SCE_M1045_g N_A_691_113#_c_2274_n 0.00423625f $X=4.675 $Y=2.585 $X2=0
+ $Y2=0
cc_856 N_SCE_c_1051_n N_A_691_113#_c_2339_n 0.00461132f $X=3.655 $Y=3.025 $X2=0
+ $Y2=0
cc_857 N_SCE_c_1052_n N_A_691_113#_c_2275_n 0.0235692f $X=4.585 $Y=3.1 $X2=0
+ $Y2=0
cc_858 N_SCE_M1045_g N_A_691_113#_c_2275_n 0.0077662f $X=4.675 $Y=2.585 $X2=0
+ $Y2=0
cc_859 N_SCE_c_1051_n N_A_691_113#_c_2286_n 0.00342836f $X=3.655 $Y=3.025 $X2=0
+ $Y2=0
cc_860 N_SCE_c_1052_n N_A_691_113#_c_2286_n 0.00845974f $X=4.585 $Y=3.1 $X2=0
+ $Y2=0
cc_861 N_SCE_c_1053_n N_A_691_113#_c_2286_n 0.00108712f $X=3.73 $Y=3.1 $X2=0
+ $Y2=0
cc_862 N_SCE_M1045_g N_A_691_113#_c_2302_n 0.0165657f $X=4.675 $Y=2.585 $X2=0
+ $Y2=0
cc_863 N_SCE_c_1055_n N_A_691_113#_c_2277_n 5.28827e-19 $X=4.675 $Y=2.19 $X2=0
+ $Y2=0
cc_864 N_SCE_M1045_g N_A_691_113#_c_2277_n 0.00655934f $X=4.675 $Y=2.585 $X2=0
+ $Y2=0
cc_865 N_SCE_M1036_g N_A_691_113#_c_2266_n 0.0109232f $X=5.77 $Y=0.835 $X2=0
+ $Y2=0
cc_866 N_SCE_c_1051_n N_A_691_113#_c_2272_n 0.00327539f $X=3.655 $Y=3.025 $X2=0
+ $Y2=0
cc_867 N_SCE_M1036_g N_A_691_113#_c_2273_n 0.00377254f $X=5.77 $Y=0.835 $X2=0
+ $Y2=0
cc_868 N_SCE_M1039_g N_VGND_c_2511_n 0.0126683f $X=4.84 $Y=0.835 $X2=0 $Y2=0
cc_869 N_SCE_c_1046_n N_VGND_c_2511_n 0.0244098f $X=5.695 $Y=0.18 $X2=0 $Y2=0
cc_870 N_SCE_M1036_g N_VGND_c_2511_n 0.00789535f $X=5.77 $Y=0.835 $X2=0 $Y2=0
cc_871 N_SCE_c_1046_n N_VGND_c_2512_n 0.0109961f $X=5.695 $Y=0.18 $X2=0 $Y2=0
cc_872 N_SCE_M1036_g N_VGND_c_2512_n 6.60132e-19 $X=5.77 $Y=0.835 $X2=0 $Y2=0
cc_873 N_SCE_c_1047_n N_VGND_c_2531_n 0.00729633f $X=4.915 $Y=0.18 $X2=0 $Y2=0
cc_874 N_SCE_c_1046_n N_VGND_c_2532_n 0.0201823f $X=5.695 $Y=0.18 $X2=0 $Y2=0
cc_875 N_SCE_c_1046_n N_VGND_c_2544_n 0.0326416f $X=5.695 $Y=0.18 $X2=0 $Y2=0
cc_876 N_SCE_c_1047_n N_VGND_c_2544_n 0.0106185f $X=4.915 $Y=0.18 $X2=0 $Y2=0
cc_877 N_CLK_c_1127_n N_A_1374_368#_c_1425_n 0.00710614f $X=6.795 $Y=1.765 $X2=0
+ $Y2=0
cc_878 CLK N_A_1374_368#_c_1425_n 0.00659815f $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_879 N_CLK_c_1127_n N_A_1374_368#_c_1411_n 5.12853e-19 $X=6.795 $Y=1.765 $X2=0
+ $Y2=0
cc_880 N_CLK_c_1128_n N_A_1374_368#_c_1411_n 0.0115578f $X=6.865 $Y=1.22 $X2=0
+ $Y2=0
cc_881 CLK N_A_1374_368#_c_1411_n 0.00829649f $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_882 N_CLK_c_1127_n N_A_1374_368#_c_1412_n 0.00487523f $X=6.795 $Y=1.765 $X2=0
+ $Y2=0
cc_883 N_CLK_c_1127_n N_A_1374_368#_c_1429_n 0.00502083f $X=6.795 $Y=1.765 $X2=0
+ $Y2=0
cc_884 N_CLK_c_1127_n N_A_1374_368#_c_1413_n 0.00200244f $X=6.795 $Y=1.765 $X2=0
+ $Y2=0
cc_885 N_CLK_c_1128_n N_A_1374_368#_c_1413_n 0.00389062f $X=6.865 $Y=1.22 $X2=0
+ $Y2=0
cc_886 CLK N_A_1374_368#_c_1413_n 0.0298284f $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_887 N_CLK_c_1127_n N_A_1374_368#_c_1415_n 0.00895263f $X=6.795 $Y=1.765 $X2=0
+ $Y2=0
cc_888 CLK N_A_1374_368#_c_1415_n 2.18476e-19 $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_889 N_CLK_c_1127_n N_VPWR_c_2070_n 0.0209712f $X=6.795 $Y=1.765 $X2=0 $Y2=0
cc_890 N_CLK_c_1127_n N_VPWR_c_2086_n 0.00413917f $X=6.795 $Y=1.765 $X2=0 $Y2=0
cc_891 N_CLK_c_1127_n N_VPWR_c_2066_n 0.00421563f $X=6.795 $Y=1.765 $X2=0 $Y2=0
cc_892 N_CLK_c_1128_n N_A_691_113#_c_2266_n 0.00440404f $X=6.865 $Y=1.22 $X2=0
+ $Y2=0
cc_893 N_CLK_c_1127_n N_A_691_113#_c_2267_n 0.0168923f $X=6.795 $Y=1.765 $X2=0
+ $Y2=0
cc_894 CLK N_A_691_113#_c_2267_n 0.0174202f $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_895 N_CLK_c_1127_n N_A_691_113#_c_2279_n 0.0172284f $X=6.795 $Y=1.765 $X2=0
+ $Y2=0
cc_896 N_CLK_c_1127_n N_A_691_113#_c_2280_n 0.00677945f $X=6.795 $Y=1.765 $X2=0
+ $Y2=0
cc_897 N_CLK_c_1127_n N_A_691_113#_c_2273_n 8.76987e-19 $X=6.795 $Y=1.765 $X2=0
+ $Y2=0
cc_898 N_CLK_c_1128_n N_A_691_113#_c_2273_n 0.00334486f $X=6.865 $Y=1.22 $X2=0
+ $Y2=0
cc_899 CLK N_A_691_113#_c_2273_n 0.0054797f $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_900 N_CLK_c_1127_n N_VGND_c_2512_n 2.21461e-19 $X=6.795 $Y=1.765 $X2=0 $Y2=0
cc_901 N_CLK_c_1128_n N_VGND_c_2512_n 0.0157427f $X=6.865 $Y=1.22 $X2=0 $Y2=0
cc_902 CLK N_VGND_c_2512_n 0.00209233f $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_903 N_CLK_c_1128_n N_VGND_c_2513_n 0.00305448f $X=6.865 $Y=1.22 $X2=0 $Y2=0
cc_904 N_CLK_c_1128_n N_VGND_c_2527_n 0.00434272f $X=6.865 $Y=1.22 $X2=0 $Y2=0
cc_905 N_CLK_c_1128_n N_VGND_c_2544_n 0.00830058f $X=6.865 $Y=1.22 $X2=0 $Y2=0
cc_906 N_A_1586_74#_c_1166_n N_A_1374_368#_M1003_g 0.00979223f $X=8.07 $Y=0.515
+ $X2=0 $Y2=0
cc_907 N_A_1586_74#_c_1168_n N_A_1374_368#_M1003_g 0.00474255f $X=8.235 $Y=0.34
+ $X2=0 $Y2=0
cc_908 N_A_1586_74#_c_1166_n N_A_1374_368#_c_1403_n 0.0012801f $X=8.07 $Y=0.515
+ $X2=0 $Y2=0
cc_909 N_A_1586_74#_c_1190_n N_A_1374_368#_c_1417_n 0.0038875f $X=8.725 $Y=1.98
+ $X2=0 $Y2=0
cc_910 N_A_1586_74#_c_1192_n N_A_1374_368#_c_1417_n 4.56175e-19 $X=8.89 $Y=1.98
+ $X2=0 $Y2=0
cc_911 N_A_1586_74#_c_1182_n N_A_1374_368#_c_1417_n 0.00115424f $X=8.89 $Y=1.82
+ $X2=0 $Y2=0
cc_912 N_A_1586_74#_c_1194_n N_A_1374_368#_c_1417_n 0.00503455f $X=8.89 $Y=2.14
+ $X2=0 $Y2=0
cc_913 N_A_1586_74#_c_1190_n N_A_1374_368#_c_1404_n 0.00871102f $X=8.725 $Y=1.98
+ $X2=0 $Y2=0
cc_914 N_A_1586_74#_c_1192_n N_A_1374_368#_c_1404_n 0.00441444f $X=8.89 $Y=1.98
+ $X2=0 $Y2=0
cc_915 N_A_1586_74#_c_1194_n N_A_1374_368#_c_1404_n 0.0186888f $X=8.89 $Y=2.14
+ $X2=0 $Y2=0
cc_916 N_A_1586_74#_c_1163_n N_A_1374_368#_M1037_g 0.013497f $X=9.525 $Y=1.015
+ $X2=0 $Y2=0
cc_917 N_A_1586_74#_c_1166_n N_A_1374_368#_M1037_g 0.00327787f $X=8.07 $Y=0.515
+ $X2=0 $Y2=0
cc_918 N_A_1586_74#_c_1167_n N_A_1374_368#_M1037_g 0.00929412f $X=8.885 $Y=0.34
+ $X2=0 $Y2=0
cc_919 N_A_1586_74#_c_1182_n N_A_1374_368#_M1037_g 0.0298706f $X=8.89 $Y=1.82
+ $X2=0 $Y2=0
cc_920 N_A_1586_74#_c_1183_n N_A_1374_368#_M1037_g 0.00206916f $X=8.97 $Y=0.34
+ $X2=0 $Y2=0
cc_921 N_A_1586_74#_c_1171_n N_A_1374_368#_c_1406_n 4.9149e-19 $X=9.69 $Y=1.18
+ $X2=0 $Y2=0
cc_922 N_A_1586_74#_c_1172_n N_A_1374_368#_c_1406_n 0.0133907f $X=9.69 $Y=1.18
+ $X2=0 $Y2=0
cc_923 N_A_1586_74#_c_1182_n N_A_1374_368#_c_1406_n 0.0076216f $X=8.89 $Y=1.82
+ $X2=0 $Y2=0
cc_924 N_A_1586_74#_c_1194_n N_A_1374_368#_c_1406_n 0.00712942f $X=8.89 $Y=2.14
+ $X2=0 $Y2=0
cc_925 N_A_1586_74#_c_1182_n N_A_1374_368#_c_1420_n 4.63241e-19 $X=8.89 $Y=1.82
+ $X2=0 $Y2=0
cc_926 N_A_1586_74#_c_1194_n N_A_1374_368#_c_1420_n 0.00326764f $X=8.89 $Y=2.14
+ $X2=0 $Y2=0
cc_927 N_A_1586_74#_c_1187_n N_A_1374_368#_c_1421_n 0.0100863f $X=9.195 $Y=2.465
+ $X2=0 $Y2=0
cc_928 N_A_1586_74#_c_1172_n N_A_1374_368#_c_1421_n 0.00184435f $X=9.69 $Y=1.18
+ $X2=0 $Y2=0
cc_929 N_A_1586_74#_c_1194_n N_A_1374_368#_c_1421_n 0.0152709f $X=8.89 $Y=2.14
+ $X2=0 $Y2=0
cc_930 N_A_1586_74#_c_1165_n N_A_1374_368#_c_1407_n 0.0192432f $X=13.285
+ $Y=2.375 $X2=0 $Y2=0
cc_931 N_A_1586_74#_c_1189_n N_A_1374_368#_c_1407_n 0.0131701f $X=13.285
+ $Y=2.465 $X2=0 $Y2=0
cc_932 N_A_1586_74#_c_1180_n N_A_1374_368#_c_1407_n 3.6914e-19 $X=12.26 $Y=1.635
+ $X2=0 $Y2=0
cc_933 N_A_1586_74#_c_1181_n N_A_1374_368#_c_1407_n 0.00456417f $X=13.195
+ $Y=1.215 $X2=0 $Y2=0
cc_934 N_A_1586_74#_c_1185_n N_A_1374_368#_c_1407_n 0.0213123f $X=13.36 $Y=1.39
+ $X2=0 $Y2=0
cc_935 N_A_1586_74#_c_1186_n N_A_1374_368#_c_1407_n 0.021367f $X=12.37 $Y=1.635
+ $X2=0 $Y2=0
cc_936 N_A_1586_74#_M1011_g N_A_1374_368#_M1013_g 0.0293304f $X=12.37 $Y=0.69
+ $X2=0 $Y2=0
cc_937 N_A_1586_74#_c_1180_n N_A_1374_368#_M1013_g 8.82425e-19 $X=12.26 $Y=1.635
+ $X2=0 $Y2=0
cc_938 N_A_1586_74#_c_1181_n N_A_1374_368#_M1013_g 0.0114972f $X=13.195 $Y=1.215
+ $X2=0 $Y2=0
cc_939 N_A_1586_74#_c_1184_n N_A_1374_368#_M1013_g 0.00153298f $X=13.36 $Y=1.215
+ $X2=0 $Y2=0
cc_940 N_A_1586_74#_c_1185_n N_A_1374_368#_M1013_g 0.0135859f $X=13.36 $Y=1.39
+ $X2=0 $Y2=0
cc_941 N_A_1586_74#_c_1190_n N_A_1374_368#_c_1409_n 3.47737e-19 $X=8.725 $Y=1.98
+ $X2=0 $Y2=0
cc_942 N_A_1586_74#_c_1182_n N_A_1374_368#_c_1409_n 6.6446e-19 $X=8.89 $Y=1.82
+ $X2=0 $Y2=0
cc_943 N_A_1586_74#_c_1182_n N_A_1374_368#_c_1410_n 0.00342855f $X=8.89 $Y=1.82
+ $X2=0 $Y2=0
cc_944 N_A_1586_74#_c_1180_n N_A_1374_368#_c_1426_n 0.00881567f $X=12.26
+ $Y=1.635 $X2=0 $Y2=0
cc_945 N_A_1586_74#_c_1186_n N_A_1374_368#_c_1426_n 0.00321743f $X=12.37
+ $Y=1.635 $X2=0 $Y2=0
cc_946 N_A_1586_74#_c_1165_n N_A_1374_368#_c_1427_n 6.17953e-19 $X=13.285
+ $Y=2.375 $X2=0 $Y2=0
cc_947 N_A_1586_74#_c_1180_n N_A_1374_368#_c_1414_n 0.0248923f $X=12.26 $Y=1.635
+ $X2=0 $Y2=0
cc_948 N_A_1586_74#_c_1181_n N_A_1374_368#_c_1414_n 0.0303637f $X=13.195
+ $Y=1.215 $X2=0 $Y2=0
cc_949 N_A_1586_74#_c_1184_n N_A_1374_368#_c_1414_n 0.00481086f $X=13.36
+ $Y=1.215 $X2=0 $Y2=0
cc_950 N_A_1586_74#_c_1185_n N_A_1374_368#_c_1414_n 0.00193886f $X=13.36 $Y=1.39
+ $X2=0 $Y2=0
cc_951 N_A_1586_74#_c_1186_n N_A_1374_368#_c_1414_n 0.00195577f $X=12.37
+ $Y=1.635 $X2=0 $Y2=0
cc_952 N_A_1586_74#_c_1174_n N_A_2013_71#_M1023_d 0.00350583f $X=11.37 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_953 N_A_1586_74#_c_1163_n N_A_2013_71#_M1034_g 0.013612f $X=9.525 $Y=1.015
+ $X2=0 $Y2=0
cc_954 N_A_1586_74#_c_1169_n N_A_2013_71#_M1034_g 7.07453e-19 $X=9.565 $Y=0.34
+ $X2=0 $Y2=0
cc_955 N_A_1586_74#_c_1170_n N_A_2013_71#_M1034_g 0.00524926f $X=9.65 $Y=0.85
+ $X2=0 $Y2=0
cc_956 N_A_1586_74#_c_1171_n N_A_2013_71#_M1034_g 0.00166923f $X=9.69 $Y=1.18
+ $X2=0 $Y2=0
cc_957 N_A_1586_74#_c_1172_n N_A_2013_71#_M1034_g 0.0210021f $X=9.69 $Y=1.18
+ $X2=0 $Y2=0
cc_958 N_A_1586_74#_c_1173_n N_A_2013_71#_M1034_g 0.0138659f $X=10.69 $Y=0.935
+ $X2=0 $Y2=0
cc_959 N_A_1586_74#_c_1273_p N_A_2013_71#_M1034_g 0.00308709f $X=10.775 $Y=0.85
+ $X2=0 $Y2=0
cc_960 N_A_1586_74#_M1011_g N_A_2013_71#_c_1594_n 0.0056233f $X=12.37 $Y=0.69
+ $X2=0 $Y2=0
cc_961 N_A_1586_74#_c_1179_n N_A_2013_71#_c_1594_n 0.00681315f $X=12.23 $Y=1.3
+ $X2=0 $Y2=0
cc_962 N_A_1586_74#_c_1180_n N_A_2013_71#_c_1594_n 0.00612418f $X=12.26 $Y=1.635
+ $X2=0 $Y2=0
cc_963 N_A_1586_74#_c_1186_n N_A_2013_71#_c_1594_n 0.0210373f $X=12.37 $Y=1.635
+ $X2=0 $Y2=0
cc_964 N_A_1586_74#_M1011_g N_A_2013_71#_c_1596_n 0.0605761f $X=12.37 $Y=0.69
+ $X2=0 $Y2=0
cc_965 N_A_1586_74#_c_1174_n N_A_2013_71#_c_1596_n 6.63977e-19 $X=11.37 $Y=0.34
+ $X2=0 $Y2=0
cc_966 N_A_1586_74#_c_1176_n N_A_2013_71#_c_1596_n 0.004173f $X=11.455 $Y=0.85
+ $X2=0 $Y2=0
cc_967 N_A_1586_74#_c_1177_n N_A_2013_71#_c_1596_n 0.0123107f $X=12.08 $Y=0.935
+ $X2=0 $Y2=0
cc_968 N_A_1586_74#_c_1179_n N_A_2013_71#_c_1596_n 0.0052319f $X=12.23 $Y=1.3
+ $X2=0 $Y2=0
cc_969 N_A_1586_74#_c_1173_n N_A_2013_71#_c_1597_n 0.035239f $X=10.69 $Y=0.935
+ $X2=0 $Y2=0
cc_970 N_A_1586_74#_c_1173_n N_A_2013_71#_c_1598_n 0.00750114f $X=10.69 $Y=0.935
+ $X2=0 $Y2=0
cc_971 N_A_1586_74#_c_1174_n N_A_2013_71#_c_1598_n 0.0127109f $X=11.37 $Y=0.34
+ $X2=0 $Y2=0
cc_972 N_A_1586_74#_c_1176_n N_A_2013_71#_c_1598_n 0.0188234f $X=11.455 $Y=0.85
+ $X2=0 $Y2=0
cc_973 N_A_1586_74#_c_1178_n N_A_2013_71#_c_1598_n 0.0141448f $X=11.54 $Y=0.935
+ $X2=0 $Y2=0
cc_974 N_A_1586_74#_c_1178_n N_A_2013_71#_c_1600_n 0.00130064f $X=11.54 $Y=0.935
+ $X2=0 $Y2=0
cc_975 N_A_1586_74#_M1011_g N_A_2013_71#_c_1601_n 2.44748e-19 $X=12.37 $Y=0.69
+ $X2=0 $Y2=0
cc_976 N_A_1586_74#_c_1177_n N_A_2013_71#_c_1601_n 0.0251569f $X=12.08 $Y=0.935
+ $X2=0 $Y2=0
cc_977 N_A_1586_74#_c_1178_n N_A_2013_71#_c_1601_n 0.01265f $X=11.54 $Y=0.935
+ $X2=0 $Y2=0
cc_978 N_A_1586_74#_c_1179_n N_A_2013_71#_c_1601_n 0.00844044f $X=12.23 $Y=1.3
+ $X2=0 $Y2=0
cc_979 N_A_1586_74#_c_1180_n N_A_2013_71#_c_1601_n 0.0163961f $X=12.26 $Y=1.635
+ $X2=0 $Y2=0
cc_980 N_A_1586_74#_c_1174_n N_A_2013_71#_c_1602_n 0.00351137f $X=11.37 $Y=0.34
+ $X2=0 $Y2=0
cc_981 N_A_1586_74#_c_1177_n N_A_2013_71#_c_1602_n 0.0113034f $X=12.08 $Y=0.935
+ $X2=0 $Y2=0
cc_982 N_A_1586_74#_c_1178_n N_A_2013_71#_c_1602_n 0.00455524f $X=11.54 $Y=0.935
+ $X2=0 $Y2=0
cc_983 N_A_1586_74#_c_1171_n N_A_2013_71#_c_1603_n 0.00972664f $X=9.69 $Y=1.18
+ $X2=0 $Y2=0
cc_984 N_A_1586_74#_c_1172_n N_A_2013_71#_c_1603_n 5.60957e-19 $X=9.69 $Y=1.18
+ $X2=0 $Y2=0
cc_985 N_A_1586_74#_c_1173_n N_A_2013_71#_c_1603_n 0.0235913f $X=10.69 $Y=0.935
+ $X2=0 $Y2=0
cc_986 N_A_1586_74#_c_1173_n N_A_2013_71#_c_1604_n 0.00125903f $X=10.69 $Y=0.935
+ $X2=0 $Y2=0
cc_987 N_A_1586_74#_c_1182_n N_A_1784_97#_M1037_d 0.0043242f $X=8.89 $Y=1.82
+ $X2=-0.19 $Y2=-0.245
cc_988 N_A_1586_74#_c_1173_n N_A_1784_97#_M1023_g 0.00576525f $X=10.69 $Y=0.935
+ $X2=0 $Y2=0
cc_989 N_A_1586_74#_c_1273_p N_A_1784_97#_M1023_g 0.0116034f $X=10.775 $Y=0.85
+ $X2=0 $Y2=0
cc_990 N_A_1586_74#_c_1174_n N_A_1784_97#_M1023_g 0.0112842f $X=11.37 $Y=0.34
+ $X2=0 $Y2=0
cc_991 N_A_1586_74#_c_1175_n N_A_1784_97#_M1023_g 0.00332344f $X=10.86 $Y=0.34
+ $X2=0 $Y2=0
cc_992 N_A_1586_74#_c_1176_n N_A_1784_97#_M1023_g 0.00327684f $X=11.455 $Y=0.85
+ $X2=0 $Y2=0
cc_993 N_A_1586_74#_c_1163_n N_A_1784_97#_c_1708_n 0.00497183f $X=9.525 $Y=1.015
+ $X2=0 $Y2=0
cc_994 N_A_1586_74#_c_1169_n N_A_1784_97#_c_1708_n 0.012971f $X=9.565 $Y=0.34
+ $X2=0 $Y2=0
cc_995 N_A_1586_74#_c_1171_n N_A_1784_97#_c_1708_n 0.0241468f $X=9.69 $Y=1.18
+ $X2=0 $Y2=0
cc_996 N_A_1586_74#_c_1182_n N_A_1784_97#_c_1708_n 0.0805264f $X=8.89 $Y=1.82
+ $X2=0 $Y2=0
cc_997 N_A_1586_74#_c_1311_p N_A_1784_97#_c_1708_n 0.0114261f $X=9.71 $Y=0.935
+ $X2=0 $Y2=0
cc_998 N_A_1586_74#_c_1171_n N_A_1784_97#_c_1710_n 0.0087019f $X=9.69 $Y=1.18
+ $X2=0 $Y2=0
cc_999 N_A_1586_74#_c_1172_n N_A_1784_97#_c_1710_n 0.00188502f $X=9.69 $Y=1.18
+ $X2=0 $Y2=0
cc_1000 N_A_1586_74#_c_1173_n N_A_1784_97#_c_1710_n 0.00312506f $X=10.69
+ $Y=0.935 $X2=0 $Y2=0
cc_1001 N_A_1586_74#_c_1182_n N_A_1784_97#_c_1711_n 0.0136362f $X=8.89 $Y=1.82
+ $X2=0 $Y2=0
cc_1002 N_A_1586_74#_c_1187_n N_A_1784_97#_c_1712_n 0.00658301f $X=9.195
+ $Y=2.465 $X2=0 $Y2=0
cc_1003 N_A_1586_74#_c_1187_n N_A_1784_97#_c_1713_n 0.00163453f $X=9.195
+ $Y=2.465 $X2=0 $Y2=0
cc_1004 N_A_1586_74#_c_1192_n N_A_1784_97#_c_1713_n 0.0333201f $X=8.89 $Y=1.98
+ $X2=0 $Y2=0
cc_1005 N_A_1586_74#_c_1194_n N_A_1784_97#_c_1713_n 0.01442f $X=8.89 $Y=2.14
+ $X2=0 $Y2=0
cc_1006 N_A_1586_74#_M1011_g N_A_2489_74#_c_1871_n 0.00274767f $X=12.37 $Y=0.69
+ $X2=0 $Y2=0
cc_1007 N_A_1586_74#_c_1181_n N_A_2489_74#_c_1871_n 0.0224089f $X=13.195
+ $Y=1.215 $X2=0 $Y2=0
cc_1008 N_A_1586_74#_M1011_g N_A_2489_74#_c_1797_n 0.00726238f $X=12.37 $Y=0.69
+ $X2=0 $Y2=0
cc_1009 N_A_1586_74#_c_1181_n N_A_2489_74#_c_1798_n 0.0298078f $X=13.195
+ $Y=1.215 $X2=0 $Y2=0
cc_1010 N_A_1586_74#_c_1184_n N_A_2489_74#_c_1798_n 0.0233024f $X=13.36 $Y=1.215
+ $X2=0 $Y2=0
cc_1011 N_A_1586_74#_c_1185_n N_A_2489_74#_c_1798_n 3.05108e-19 $X=13.36 $Y=1.39
+ $X2=0 $Y2=0
cc_1012 N_A_1586_74#_c_1165_n N_A_2489_74#_c_1807_n 0.0139101f $X=13.285
+ $Y=2.375 $X2=0 $Y2=0
cc_1013 N_A_1586_74#_c_1189_n N_A_2489_74#_c_1807_n 0.00535595f $X=13.285
+ $Y=2.465 $X2=0 $Y2=0
cc_1014 N_A_1586_74#_c_1165_n N_A_2489_74#_c_1808_n 0.00547079f $X=13.285
+ $Y=2.375 $X2=0 $Y2=0
cc_1015 N_A_1586_74#_c_1184_n N_A_2489_74#_c_1808_n 0.0129484f $X=13.36 $Y=1.215
+ $X2=0 $Y2=0
cc_1016 N_A_1586_74#_c_1185_n N_A_2489_74#_c_1808_n 0.00334366f $X=13.36 $Y=1.39
+ $X2=0 $Y2=0
cc_1017 N_A_1586_74#_c_1165_n N_A_2489_74#_c_1809_n 0.00374558f $X=13.285
+ $Y=2.375 $X2=0 $Y2=0
cc_1018 N_A_1586_74#_c_1181_n N_A_2489_74#_c_1809_n 0.00104657f $X=13.195
+ $Y=1.215 $X2=0 $Y2=0
cc_1019 N_A_1586_74#_c_1184_n N_A_2489_74#_c_1809_n 0.00824827f $X=13.36
+ $Y=1.215 $X2=0 $Y2=0
cc_1020 N_A_1586_74#_c_1184_n N_A_2489_74#_c_1799_n 0.0315436f $X=13.36 $Y=1.215
+ $X2=0 $Y2=0
cc_1021 N_A_1586_74#_c_1185_n N_A_2489_74#_c_1799_n 0.00202138f $X=13.36 $Y=1.39
+ $X2=0 $Y2=0
cc_1022 N_A_1586_74#_c_1165_n N_A_2489_74#_c_1800_n 0.00242749f $X=13.285
+ $Y=2.375 $X2=0 $Y2=0
cc_1023 N_A_1586_74#_c_1189_n N_A_2489_74#_c_1811_n 0.0180456f $X=13.285
+ $Y=2.465 $X2=0 $Y2=0
cc_1024 N_A_1586_74#_c_1189_n N_VPWR_c_2074_n 0.00145008f $X=13.285 $Y=2.465
+ $X2=0 $Y2=0
cc_1025 N_A_1586_74#_c_1187_n N_VPWR_c_2087_n 0.00411612f $X=9.195 $Y=2.465
+ $X2=0 $Y2=0
cc_1026 N_A_1586_74#_c_1189_n N_VPWR_c_2088_n 0.00331272f $X=13.285 $Y=2.465
+ $X2=0 $Y2=0
cc_1027 N_A_1586_74#_c_1187_n N_VPWR_c_2066_n 0.00753176f $X=9.195 $Y=2.465
+ $X2=0 $Y2=0
cc_1028 N_A_1586_74#_c_1189_n N_VPWR_c_2066_n 0.00525375f $X=13.285 $Y=2.465
+ $X2=0 $Y2=0
cc_1029 N_A_1586_74#_c_1194_n N_VPWR_c_2066_n 3.3237e-19 $X=8.89 $Y=2.14 $X2=0
+ $Y2=0
cc_1030 N_A_1586_74#_c_1190_n N_A_691_113#_c_2281_n 0.013384f $X=8.725 $Y=1.98
+ $X2=0 $Y2=0
cc_1031 N_A_1586_74#_c_1192_n N_A_691_113#_c_2281_n 0.0020663f $X=8.89 $Y=1.98
+ $X2=0 $Y2=0
cc_1032 N_A_1586_74#_c_1166_n N_A_691_113#_c_2268_n 0.00680159f $X=8.07 $Y=0.515
+ $X2=0 $Y2=0
cc_1033 N_A_1586_74#_c_1190_n N_A_691_113#_c_2268_n 0.0306411f $X=8.725 $Y=1.98
+ $X2=0 $Y2=0
cc_1034 N_A_1586_74#_c_1182_n N_A_691_113#_c_2268_n 0.0128117f $X=8.89 $Y=1.82
+ $X2=0 $Y2=0
cc_1035 N_A_1586_74#_c_1166_n N_A_691_113#_c_2269_n 0.00798758f $X=8.07 $Y=0.515
+ $X2=0 $Y2=0
cc_1036 N_A_1586_74#_c_1190_n N_A_691_113#_c_2295_n 0.00100393f $X=8.725 $Y=1.98
+ $X2=0 $Y2=0
cc_1037 N_A_1586_74#_c_1166_n N_A_691_113#_c_2270_n 0.0353265f $X=8.07 $Y=0.515
+ $X2=0 $Y2=0
cc_1038 N_A_1586_74#_c_1167_n N_A_691_113#_c_2270_n 0.0191962f $X=8.885 $Y=0.34
+ $X2=0 $Y2=0
cc_1039 N_A_1586_74#_c_1182_n N_A_691_113#_c_2270_n 0.0528515f $X=8.89 $Y=1.82
+ $X2=0 $Y2=0
cc_1040 N_A_1586_74#_M1001_d N_A_691_113#_c_2282_n 0.00421995f $X=8.26 $Y=1.84
+ $X2=0 $Y2=0
cc_1041 N_A_1586_74#_c_1187_n N_A_691_113#_c_2282_n 0.00203673f $X=9.195
+ $Y=2.465 $X2=0 $Y2=0
cc_1042 N_A_1586_74#_c_1190_n N_A_691_113#_c_2282_n 0.0124469f $X=8.725 $Y=1.98
+ $X2=0 $Y2=0
cc_1043 N_A_1586_74#_c_1192_n N_A_691_113#_c_2282_n 0.0270109f $X=8.89 $Y=1.98
+ $X2=0 $Y2=0
cc_1044 N_A_1586_74#_c_1194_n N_A_691_113#_c_2282_n 0.00245339f $X=8.89 $Y=2.14
+ $X2=0 $Y2=0
cc_1045 N_A_1586_74#_c_1187_n N_A_691_113#_c_2283_n 0.00164129f $X=9.195
+ $Y=2.465 $X2=0 $Y2=0
cc_1046 N_A_1586_74#_M1001_d N_A_691_113#_c_2375_n 0.00806736f $X=8.26 $Y=1.84
+ $X2=0 $Y2=0
cc_1047 N_A_1586_74#_c_1187_n N_A_691_113#_c_2375_n 3.23029e-19 $X=9.195
+ $Y=2.465 $X2=0 $Y2=0
cc_1048 N_A_1586_74#_c_1190_n N_A_691_113#_c_2375_n 0.0115323f $X=8.725 $Y=1.98
+ $X2=0 $Y2=0
cc_1049 N_A_1586_74#_c_1194_n N_A_691_113#_c_2375_n 0.00333296f $X=8.89 $Y=2.14
+ $X2=0 $Y2=0
cc_1050 N_A_1586_74#_c_1173_n N_VGND_M1034_d 0.00719284f $X=10.69 $Y=0.935 $X2=0
+ $Y2=0
cc_1051 N_A_1586_74#_c_1273_p N_VGND_M1034_d 0.00493253f $X=10.775 $Y=0.85 $X2=0
+ $Y2=0
cc_1052 N_A_1586_74#_c_1175_n N_VGND_M1034_d 5.37788e-19 $X=10.86 $Y=0.34 $X2=0
+ $Y2=0
cc_1053 N_A_1586_74#_c_1177_n N_VGND_M1009_s 0.00391333f $X=12.08 $Y=0.935 $X2=0
+ $Y2=0
cc_1054 N_A_1586_74#_c_1166_n N_VGND_c_2513_n 0.0259189f $X=8.07 $Y=0.515 $X2=0
+ $Y2=0
cc_1055 N_A_1586_74#_c_1168_n N_VGND_c_2513_n 0.010974f $X=8.235 $Y=0.34 $X2=0
+ $Y2=0
cc_1056 N_A_1586_74#_c_1169_n N_VGND_c_2514_n 0.00662337f $X=9.565 $Y=0.34 $X2=0
+ $Y2=0
cc_1057 N_A_1586_74#_c_1170_n N_VGND_c_2514_n 0.00506803f $X=9.65 $Y=0.85 $X2=0
+ $Y2=0
cc_1058 N_A_1586_74#_c_1173_n N_VGND_c_2514_n 0.0196718f $X=10.69 $Y=0.935 $X2=0
+ $Y2=0
cc_1059 N_A_1586_74#_c_1273_p N_VGND_c_2514_n 0.0190358f $X=10.775 $Y=0.85 $X2=0
+ $Y2=0
cc_1060 N_A_1586_74#_c_1175_n N_VGND_c_2514_n 0.0145685f $X=10.86 $Y=0.34 $X2=0
+ $Y2=0
cc_1061 N_A_1586_74#_M1011_g N_VGND_c_2515_n 0.00147043f $X=12.37 $Y=0.69 $X2=0
+ $Y2=0
cc_1062 N_A_1586_74#_c_1174_n N_VGND_c_2515_n 0.0146661f $X=11.37 $Y=0.34 $X2=0
+ $Y2=0
cc_1063 N_A_1586_74#_c_1176_n N_VGND_c_2515_n 0.0193741f $X=11.455 $Y=0.85 $X2=0
+ $Y2=0
cc_1064 N_A_1586_74#_c_1177_n N_VGND_c_2515_n 0.015048f $X=12.08 $Y=0.935 $X2=0
+ $Y2=0
cc_1065 N_A_1586_74#_M1011_g N_VGND_c_2529_n 0.00434272f $X=12.37 $Y=0.69 $X2=0
+ $Y2=0
cc_1066 N_A_1586_74#_c_1163_n N_VGND_c_2533_n 7.53287e-19 $X=9.525 $Y=1.015
+ $X2=0 $Y2=0
cc_1067 N_A_1586_74#_c_1167_n N_VGND_c_2533_n 0.0418136f $X=8.885 $Y=0.34 $X2=0
+ $Y2=0
cc_1068 N_A_1586_74#_c_1168_n N_VGND_c_2533_n 0.0235688f $X=8.235 $Y=0.34 $X2=0
+ $Y2=0
cc_1069 N_A_1586_74#_c_1169_n N_VGND_c_2533_n 0.0449818f $X=9.565 $Y=0.34 $X2=0
+ $Y2=0
cc_1070 N_A_1586_74#_c_1183_n N_VGND_c_2533_n 0.0121867f $X=8.97 $Y=0.34 $X2=0
+ $Y2=0
cc_1071 N_A_1586_74#_c_1174_n N_VGND_c_2534_n 0.0446499f $X=11.37 $Y=0.34 $X2=0
+ $Y2=0
cc_1072 N_A_1586_74#_c_1175_n N_VGND_c_2534_n 0.0120637f $X=10.86 $Y=0.34 $X2=0
+ $Y2=0
cc_1073 N_A_1586_74#_M1011_g N_VGND_c_2544_n 0.00821463f $X=12.37 $Y=0.69 $X2=0
+ $Y2=0
cc_1074 N_A_1586_74#_c_1167_n N_VGND_c_2544_n 0.0244305f $X=8.885 $Y=0.34 $X2=0
+ $Y2=0
cc_1075 N_A_1586_74#_c_1168_n N_VGND_c_2544_n 0.0127152f $X=8.235 $Y=0.34 $X2=0
+ $Y2=0
cc_1076 N_A_1586_74#_c_1169_n N_VGND_c_2544_n 0.025776f $X=9.565 $Y=0.34 $X2=0
+ $Y2=0
cc_1077 N_A_1586_74#_c_1173_n N_VGND_c_2544_n 0.0203559f $X=10.69 $Y=0.935 $X2=0
+ $Y2=0
cc_1078 N_A_1586_74#_c_1174_n N_VGND_c_2544_n 0.0252533f $X=11.37 $Y=0.34 $X2=0
+ $Y2=0
cc_1079 N_A_1586_74#_c_1175_n N_VGND_c_2544_n 0.00644906f $X=10.86 $Y=0.34 $X2=0
+ $Y2=0
cc_1080 N_A_1586_74#_c_1177_n N_VGND_c_2544_n 0.00988673f $X=12.08 $Y=0.935
+ $X2=0 $Y2=0
cc_1081 N_A_1586_74#_c_1179_n N_VGND_c_2544_n 0.00660638f $X=12.23 $Y=1.3 $X2=0
+ $Y2=0
cc_1082 N_A_1586_74#_c_1183_n N_VGND_c_2544_n 0.00660921f $X=8.97 $Y=0.34 $X2=0
+ $Y2=0
cc_1083 N_A_1586_74#_c_1311_p N_VGND_c_2544_n 0.00454674f $X=9.71 $Y=0.935 $X2=0
+ $Y2=0
cc_1084 N_A_1586_74#_c_1170_n A_1920_97# 0.00506914f $X=9.65 $Y=0.85 $X2=-0.19
+ $Y2=-0.245
cc_1085 N_A_1586_74#_c_1173_n A_1920_97# 0.00308187f $X=10.69 $Y=0.935 $X2=-0.19
+ $Y2=-0.245
cc_1086 N_A_1586_74#_c_1311_p A_1920_97# 0.00274383f $X=9.71 $Y=0.935 $X2=-0.19
+ $Y2=-0.245
cc_1087 N_A_1586_74#_c_1179_n A_2417_74# 0.00229931f $X=12.23 $Y=1.3 $X2=-0.19
+ $Y2=-0.245
cc_1088 N_A_1374_368#_c_1426_n N_A_2013_71#_M1030_d 0.0079555f $X=12.55 $Y=2.475
+ $X2=0 $Y2=0
cc_1089 N_A_1374_368#_c_1406_n N_A_2013_71#_c_1593_n 0.014422f $X=9.525 $Y=1.66
+ $X2=0 $Y2=0
cc_1090 N_A_1374_368#_c_1421_n N_A_2013_71#_c_1593_n 0.0229417f $X=9.645
+ $Y=2.465 $X2=0 $Y2=0
cc_1091 N_A_1374_368#_c_1430_n N_A_2013_71#_c_1593_n 0.00864601f $X=9.69
+ $Y=2.195 $X2=0 $Y2=0
cc_1092 N_A_1374_368#_c_1421_n N_A_2013_71#_c_1606_n 0.0201335f $X=9.645
+ $Y=2.465 $X2=0 $Y2=0
cc_1093 N_A_1374_368#_c_1426_n N_A_2013_71#_c_1606_n 0.0153246f $X=12.55
+ $Y=2.475 $X2=0 $Y2=0
cc_1094 N_A_1374_368#_c_1426_n N_A_2013_71#_c_1608_n 0.0203243f $X=12.55
+ $Y=2.475 $X2=0 $Y2=0
cc_1095 N_A_1374_368#_c_1427_n N_A_2013_71#_c_1608_n 0.0119913f $X=12.635
+ $Y=2.39 $X2=0 $Y2=0
cc_1096 N_A_1374_368#_c_1426_n N_A_2013_71#_c_1609_n 0.0432777f $X=12.55
+ $Y=2.475 $X2=0 $Y2=0
cc_1097 N_A_1374_368#_c_1426_n N_A_1784_97#_c_1706_n 0.0157356f $X=12.55
+ $Y=2.475 $X2=0 $Y2=0
cc_1098 N_A_1374_368#_M1037_g N_A_1784_97#_c_1708_n 0.00328193f $X=8.845
+ $Y=0.695 $X2=0 $Y2=0
cc_1099 N_A_1374_368#_c_1406_n N_A_1784_97#_c_1708_n 0.00874168f $X=9.525
+ $Y=1.66 $X2=0 $Y2=0
cc_1100 N_A_1374_368#_c_1406_n N_A_1784_97#_c_1710_n 0.00795059f $X=9.525
+ $Y=1.66 $X2=0 $Y2=0
cc_1101 N_A_1374_368#_c_1420_n N_A_1784_97#_c_1710_n 0.0086077f $X=9.6 $Y=2.03
+ $X2=0 $Y2=0
cc_1102 N_A_1374_368#_c_1421_n N_A_1784_97#_c_1710_n 7.55709e-19 $X=9.645
+ $Y=2.465 $X2=0 $Y2=0
cc_1103 N_A_1374_368#_c_1426_n N_A_1784_97#_c_1710_n 0.0210569f $X=12.55
+ $Y=2.475 $X2=0 $Y2=0
cc_1104 N_A_1374_368#_c_1430_n N_A_1784_97#_c_1710_n 0.025582f $X=9.69 $Y=2.195
+ $X2=0 $Y2=0
cc_1105 N_A_1374_368#_c_1406_n N_A_1784_97#_c_1711_n 0.00465441f $X=9.525
+ $Y=1.66 $X2=0 $Y2=0
cc_1106 N_A_1374_368#_c_1421_n N_A_1784_97#_c_1712_n 0.0108277f $X=9.645
+ $Y=2.465 $X2=0 $Y2=0
cc_1107 N_A_1374_368#_c_1430_n N_A_1784_97#_c_1712_n 0.00306263f $X=9.69
+ $Y=2.195 $X2=0 $Y2=0
cc_1108 N_A_1374_368#_c_1420_n N_A_1784_97#_c_1713_n 0.00778971f $X=9.6 $Y=2.03
+ $X2=0 $Y2=0
cc_1109 N_A_1374_368#_c_1421_n N_A_1784_97#_c_1713_n 0.0013164f $X=9.645
+ $Y=2.465 $X2=0 $Y2=0
cc_1110 N_A_1374_368#_c_1430_n N_A_1784_97#_c_1713_n 0.0334058f $X=9.69 $Y=2.195
+ $X2=0 $Y2=0
cc_1111 N_A_1374_368#_c_1426_n N_A_1784_97#_c_1714_n 0.00401604f $X=12.55
+ $Y=2.475 $X2=0 $Y2=0
cc_1112 N_A_1374_368#_M1013_g N_A_2489_74#_c_1797_n 0.00236994f $X=12.88 $Y=0.58
+ $X2=0 $Y2=0
cc_1113 N_A_1374_368#_M1013_g N_A_2489_74#_c_1798_n 0.0118688f $X=12.88 $Y=0.58
+ $X2=0 $Y2=0
cc_1114 N_A_1374_368#_c_1407_n N_A_2489_74#_c_1807_n 0.00439856f $X=12.75
+ $Y=1.885 $X2=0 $Y2=0
cc_1115 N_A_1374_368#_c_1426_n N_A_2489_74#_c_1807_n 0.00511041f $X=12.55
+ $Y=2.475 $X2=0 $Y2=0
cc_1116 N_A_1374_368#_c_1427_n N_A_2489_74#_c_1807_n 0.0178676f $X=12.635
+ $Y=2.39 $X2=0 $Y2=0
cc_1117 N_A_1374_368#_c_1407_n N_A_2489_74#_c_1809_n 9.91152e-19 $X=12.75
+ $Y=1.885 $X2=0 $Y2=0
cc_1118 N_A_1374_368#_c_1427_n N_A_2489_74#_c_1809_n 0.00334249f $X=12.635
+ $Y=2.39 $X2=0 $Y2=0
cc_1119 N_A_1374_368#_c_1414_n N_A_2489_74#_c_1809_n 0.00682912f $X=12.82
+ $Y=1.635 $X2=0 $Y2=0
cc_1120 N_A_1374_368#_c_1407_n N_A_2489_74#_c_1811_n 0.010632f $X=12.75 $Y=1.885
+ $X2=0 $Y2=0
cc_1121 N_A_1374_368#_c_1426_n N_A_2489_74#_c_1811_n 0.00329601f $X=12.55
+ $Y=2.475 $X2=0 $Y2=0
cc_1122 N_A_1374_368#_c_1426_n N_VPWR_M1002_d 0.00710844f $X=12.55 $Y=2.475
+ $X2=0 $Y2=0
cc_1123 N_A_1374_368#_c_1426_n N_VPWR_M1046_s 0.0164191f $X=12.55 $Y=2.475 $X2=0
+ $Y2=0
cc_1124 N_A_1374_368#_c_1417_n N_VPWR_c_2071_n 0.0217145f $X=8.185 $Y=1.765
+ $X2=0 $Y2=0
cc_1125 N_A_1374_368#_c_1421_n N_VPWR_c_2072_n 0.00126038f $X=9.645 $Y=2.465
+ $X2=0 $Y2=0
cc_1126 N_A_1374_368#_c_1426_n N_VPWR_c_2072_n 0.0213705f $X=12.55 $Y=2.475
+ $X2=0 $Y2=0
cc_1127 N_A_1374_368#_c_1426_n N_VPWR_c_2073_n 0.0259982f $X=12.55 $Y=2.475
+ $X2=0 $Y2=0
cc_1128 N_A_1374_368#_c_1417_n N_VPWR_c_2087_n 0.00413917f $X=8.185 $Y=1.765
+ $X2=0 $Y2=0
cc_1129 N_A_1374_368#_c_1421_n N_VPWR_c_2087_n 0.00445602f $X=9.645 $Y=2.465
+ $X2=0 $Y2=0
cc_1130 N_A_1374_368#_c_1407_n N_VPWR_c_2088_n 0.00461464f $X=12.75 $Y=1.885
+ $X2=0 $Y2=0
cc_1131 N_A_1374_368#_c_1417_n N_VPWR_c_2066_n 0.00421563f $X=8.185 $Y=1.765
+ $X2=0 $Y2=0
cc_1132 N_A_1374_368#_c_1421_n N_VPWR_c_2066_n 0.00893971f $X=9.645 $Y=2.465
+ $X2=0 $Y2=0
cc_1133 N_A_1374_368#_c_1407_n N_VPWR_c_2066_n 0.00776565f $X=12.75 $Y=1.885
+ $X2=0 $Y2=0
cc_1134 N_A_1374_368#_c_1426_n N_VPWR_c_2066_n 0.078766f $X=12.55 $Y=2.475 $X2=0
+ $Y2=0
cc_1135 N_A_1374_368#_c_1430_n N_VPWR_c_2066_n 0.00695798f $X=9.69 $Y=2.195
+ $X2=0 $Y2=0
cc_1136 N_A_1374_368#_c_1425_n N_A_691_113#_c_2267_n 0.0127791f $X=7.215 $Y=1.98
+ $X2=0 $Y2=0
cc_1137 N_A_1374_368#_M1007_d N_A_691_113#_c_2279_n 0.00838267f $X=6.87 $Y=1.84
+ $X2=0 $Y2=0
cc_1138 N_A_1374_368#_c_1425_n N_A_691_113#_c_2279_n 0.0225386f $X=7.215 $Y=1.98
+ $X2=0 $Y2=0
cc_1139 N_A_1374_368#_c_1412_n N_A_691_113#_c_2279_n 0.0346f $X=7.49 $Y=1.635
+ $X2=0 $Y2=0
cc_1140 N_A_1374_368#_c_1429_n N_A_691_113#_c_2279_n 0.00229113f $X=7.49
+ $Y=1.635 $X2=0 $Y2=0
cc_1141 N_A_1374_368#_c_1415_n N_A_691_113#_c_2279_n 0.0047155f $X=7.93 $Y=1.602
+ $X2=0 $Y2=0
cc_1142 N_A_1374_368#_c_1403_n N_A_691_113#_c_2281_n 0.0066893f $X=8.095 $Y=1.66
+ $X2=0 $Y2=0
cc_1143 N_A_1374_368#_c_1417_n N_A_691_113#_c_2281_n 0.00696918f $X=8.185
+ $Y=1.765 $X2=0 $Y2=0
cc_1144 N_A_1374_368#_c_1409_n N_A_691_113#_c_2281_n 8.20479e-19 $X=8.185
+ $Y=1.675 $X2=0 $Y2=0
cc_1145 N_A_1374_368#_c_1412_n N_A_691_113#_c_2281_n 0.0264305f $X=7.49 $Y=1.635
+ $X2=0 $Y2=0
cc_1146 N_A_1374_368#_c_1429_n N_A_691_113#_c_2281_n 0.00319604f $X=7.49
+ $Y=1.635 $X2=0 $Y2=0
cc_1147 N_A_1374_368#_c_1415_n N_A_691_113#_c_2281_n 0.00171162f $X=7.93
+ $Y=1.602 $X2=0 $Y2=0
cc_1148 N_A_1374_368#_c_1403_n N_A_691_113#_c_2268_n 6.16439e-19 $X=8.095
+ $Y=1.66 $X2=0 $Y2=0
cc_1149 N_A_1374_368#_c_1404_n N_A_691_113#_c_2268_n 0.0129394f $X=8.77 $Y=1.66
+ $X2=0 $Y2=0
cc_1150 N_A_1374_368#_M1037_g N_A_691_113#_c_2268_n 0.00239961f $X=8.845
+ $Y=0.695 $X2=0 $Y2=0
cc_1151 N_A_1374_368#_c_1409_n N_A_691_113#_c_2268_n 0.00709359f $X=8.185
+ $Y=1.675 $X2=0 $Y2=0
cc_1152 N_A_1374_368#_c_1403_n N_A_691_113#_c_2269_n 0.00178115f $X=8.095
+ $Y=1.66 $X2=0 $Y2=0
cc_1153 N_A_1374_368#_c_1412_n N_A_691_113#_c_2269_n 0.00922738f $X=7.49
+ $Y=1.635 $X2=0 $Y2=0
cc_1154 N_A_1374_368#_c_1415_n N_A_691_113#_c_2269_n 0.00619128f $X=7.93
+ $Y=1.602 $X2=0 $Y2=0
cc_1155 N_A_1374_368#_c_1417_n N_A_691_113#_c_2295_n 0.0161605f $X=8.185
+ $Y=1.765 $X2=0 $Y2=0
cc_1156 N_A_1374_368#_M1003_g N_A_691_113#_c_2270_n 0.00963337f $X=7.855 $Y=0.74
+ $X2=0 $Y2=0
cc_1157 N_A_1374_368#_M1037_g N_A_691_113#_c_2270_n 0.0127542f $X=8.845 $Y=0.695
+ $X2=0 $Y2=0
cc_1158 N_A_1374_368#_c_1417_n N_A_691_113#_c_2283_n 0.00798501f $X=8.185
+ $Y=1.765 $X2=0 $Y2=0
cc_1159 N_A_1374_368#_c_1426_n A_1944_508# 0.00183207f $X=12.55 $Y=2.475
+ $X2=-0.19 $Y2=-0.245
cc_1160 N_A_1374_368#_c_1430_n A_1944_508# 0.00332423f $X=9.69 $Y=2.195
+ $X2=-0.19 $Y2=-0.245
cc_1161 N_A_1374_368#_c_1426_n A_2374_392# 0.0334166f $X=12.55 $Y=2.475
+ $X2=-0.19 $Y2=-0.245
cc_1162 N_A_1374_368#_c_1427_n A_2374_392# 0.00765757f $X=12.635 $Y=2.39
+ $X2=-0.19 $Y2=-0.245
cc_1163 N_A_1374_368#_c_1411_n N_VGND_c_2512_n 0.023367f $X=7.08 $Y=0.515 $X2=0
+ $Y2=0
cc_1164 N_A_1374_368#_M1003_g N_VGND_c_2513_n 0.00467695f $X=7.855 $Y=0.74 $X2=0
+ $Y2=0
cc_1165 N_A_1374_368#_c_1411_n N_VGND_c_2513_n 0.0618465f $X=7.08 $Y=0.515 $X2=0
+ $Y2=0
cc_1166 N_A_1374_368#_c_1412_n N_VGND_c_2513_n 0.00440058f $X=7.49 $Y=1.635
+ $X2=0 $Y2=0
cc_1167 N_A_1374_368#_c_1415_n N_VGND_c_2513_n 0.00324689f $X=7.93 $Y=1.602
+ $X2=0 $Y2=0
cc_1168 N_A_1374_368#_M1013_g N_VGND_c_2517_n 0.00128745f $X=12.88 $Y=0.58 $X2=0
+ $Y2=0
cc_1169 N_A_1374_368#_c_1411_n N_VGND_c_2527_n 0.0207821f $X=7.08 $Y=0.515 $X2=0
+ $Y2=0
cc_1170 N_A_1374_368#_M1013_g N_VGND_c_2529_n 0.00461464f $X=12.88 $Y=0.58 $X2=0
+ $Y2=0
cc_1171 N_A_1374_368#_M1003_g N_VGND_c_2533_n 0.00430908f $X=7.855 $Y=0.74 $X2=0
+ $Y2=0
cc_1172 N_A_1374_368#_M1037_g N_VGND_c_2533_n 7.53287e-19 $X=8.845 $Y=0.695
+ $X2=0 $Y2=0
cc_1173 N_A_1374_368#_M1003_g N_VGND_c_2544_n 0.0082568f $X=7.855 $Y=0.74 $X2=0
+ $Y2=0
cc_1174 N_A_1374_368#_M1013_g N_VGND_c_2544_n 0.00447595f $X=12.88 $Y=0.58 $X2=0
+ $Y2=0
cc_1175 N_A_1374_368#_c_1411_n N_VGND_c_2544_n 0.0171578f $X=7.08 $Y=0.515 $X2=0
+ $Y2=0
cc_1176 N_A_2013_71#_c_1593_n N_A_1784_97#_c_1706_n 0.0326265f $X=10.155
+ $Y=2.375 $X2=0 $Y2=0
cc_1177 N_A_2013_71#_c_1606_n N_A_1784_97#_c_1706_n 0.00936349f $X=10.155
+ $Y=2.465 $X2=0 $Y2=0
cc_1178 N_A_2013_71#_c_1597_n N_A_1784_97#_c_1706_n 0.00565038f $X=11.03
+ $Y=1.275 $X2=0 $Y2=0
cc_1179 N_A_2013_71#_c_1609_n N_A_1784_97#_c_1706_n 0.00609197f $X=11.215
+ $Y=2.135 $X2=0 $Y2=0
cc_1180 N_A_2013_71#_c_1599_n N_A_1784_97#_c_1706_n 0.0103522f $X=11.3 $Y=2.05
+ $X2=0 $Y2=0
cc_1181 N_A_2013_71#_c_1604_n N_A_1784_97#_c_1706_n 0.00132858f $X=10.23
+ $Y=1.355 $X2=0 $Y2=0
cc_1182 N_A_2013_71#_M1034_g N_A_1784_97#_M1023_g 0.0125129f $X=10.14 $Y=0.695
+ $X2=0 $Y2=0
cc_1183 N_A_2013_71#_c_1597_n N_A_1784_97#_M1023_g 0.0144178f $X=11.03 $Y=1.275
+ $X2=0 $Y2=0
cc_1184 N_A_2013_71#_c_1598_n N_A_1784_97#_M1023_g 0.00603479f $X=11.115
+ $Y=0.805 $X2=0 $Y2=0
cc_1185 N_A_2013_71#_c_1600_n N_A_1784_97#_M1023_g 0.0010369f $X=11.385 $Y=1.355
+ $X2=0 $Y2=0
cc_1186 N_A_2013_71#_c_1602_n N_A_1784_97#_M1023_g 0.0214312f $X=11.72 $Y=1.355
+ $X2=0 $Y2=0
cc_1187 N_A_2013_71#_c_1603_n N_A_1784_97#_M1023_g 8.94976e-19 $X=10.23 $Y=1.275
+ $X2=0 $Y2=0
cc_1188 N_A_2013_71#_c_1604_n N_A_1784_97#_M1023_g 0.00852329f $X=10.23 $Y=1.355
+ $X2=0 $Y2=0
cc_1189 N_A_2013_71#_M1034_g N_A_1784_97#_c_1708_n 0.00400396f $X=10.14 $Y=0.695
+ $X2=0 $Y2=0
cc_1190 N_A_2013_71#_c_1593_n N_A_1784_97#_c_1708_n 4.86365e-19 $X=10.155
+ $Y=2.375 $X2=0 $Y2=0
cc_1191 N_A_2013_71#_c_1603_n N_A_1784_97#_c_1708_n 0.00461219f $X=10.23
+ $Y=1.275 $X2=0 $Y2=0
cc_1192 N_A_2013_71#_c_1593_n N_A_1784_97#_c_1710_n 0.0137448f $X=10.155
+ $Y=2.375 $X2=0 $Y2=0
cc_1193 N_A_2013_71#_c_1597_n N_A_1784_97#_c_1710_n 0.00704001f $X=11.03
+ $Y=1.275 $X2=0 $Y2=0
cc_1194 N_A_2013_71#_c_1603_n N_A_1784_97#_c_1710_n 0.0208348f $X=10.23 $Y=1.275
+ $X2=0 $Y2=0
cc_1195 N_A_2013_71#_c_1604_n N_A_1784_97#_c_1710_n 9.81093e-19 $X=10.23
+ $Y=1.355 $X2=0 $Y2=0
cc_1196 N_A_2013_71#_c_1606_n N_A_1784_97#_c_1712_n 0.00157058f $X=10.155
+ $Y=2.465 $X2=0 $Y2=0
cc_1197 N_A_2013_71#_c_1593_n N_A_1784_97#_c_1714_n 0.001345f $X=10.155 $Y=2.375
+ $X2=0 $Y2=0
cc_1198 N_A_2013_71#_c_1597_n N_A_1784_97#_c_1714_n 0.0224081f $X=11.03 $Y=1.275
+ $X2=0 $Y2=0
cc_1199 N_A_2013_71#_c_1609_n N_A_1784_97#_c_1714_n 0.0101788f $X=11.215
+ $Y=2.135 $X2=0 $Y2=0
cc_1200 N_A_2013_71#_c_1599_n N_A_1784_97#_c_1714_n 0.0158264f $X=11.3 $Y=2.05
+ $X2=0 $Y2=0
cc_1201 N_A_2013_71#_c_1596_n N_A_2489_74#_c_1871_n 4.65641e-19 $X=12.01 $Y=1.11
+ $X2=0 $Y2=0
cc_1202 N_A_2013_71#_c_1596_n N_A_2489_74#_c_1797_n 0.00134647f $X=12.01 $Y=1.11
+ $X2=0 $Y2=0
cc_1203 N_A_2013_71#_c_1609_n N_VPWR_M1046_s 0.00351827f $X=11.215 $Y=2.135
+ $X2=0 $Y2=0
cc_1204 N_A_2013_71#_c_1599_n N_VPWR_M1046_s 0.00139771f $X=11.3 $Y=2.05 $X2=0
+ $Y2=0
cc_1205 N_A_2013_71#_c_1606_n N_VPWR_c_2072_n 0.00920075f $X=10.155 $Y=2.465
+ $X2=0 $Y2=0
cc_1206 N_A_2013_71#_c_1608_n N_VPWR_c_2073_n 0.0148532f $X=11.795 $Y=1.885
+ $X2=0 $Y2=0
cc_1207 N_A_2013_71#_c_1606_n N_VPWR_c_2087_n 0.00444681f $X=10.155 $Y=2.465
+ $X2=0 $Y2=0
cc_1208 N_A_2013_71#_c_1608_n N_VPWR_c_2088_n 0.00461464f $X=11.795 $Y=1.885
+ $X2=0 $Y2=0
cc_1209 N_A_2013_71#_c_1606_n N_VPWR_c_2066_n 0.00428411f $X=10.155 $Y=2.465
+ $X2=0 $Y2=0
cc_1210 N_A_2013_71#_c_1608_n N_VPWR_c_2066_n 0.0045644f $X=11.795 $Y=1.885
+ $X2=0 $Y2=0
cc_1211 N_A_2013_71#_M1034_g N_VGND_c_2514_n 0.00364778f $X=10.14 $Y=0.695 $X2=0
+ $Y2=0
cc_1212 N_A_2013_71#_c_1596_n N_VGND_c_2515_n 0.010393f $X=12.01 $Y=1.11 $X2=0
+ $Y2=0
cc_1213 N_A_2013_71#_c_1596_n N_VGND_c_2529_n 0.00383152f $X=12.01 $Y=1.11 $X2=0
+ $Y2=0
cc_1214 N_A_2013_71#_M1034_g N_VGND_c_2533_n 0.00497279f $X=10.14 $Y=0.695 $X2=0
+ $Y2=0
cc_1215 N_A_2013_71#_M1034_g N_VGND_c_2544_n 0.00509887f $X=10.14 $Y=0.695 $X2=0
+ $Y2=0
cc_1216 N_A_2013_71#_c_1596_n N_VGND_c_2544_n 0.0038545f $X=12.01 $Y=1.11 $X2=0
+ $Y2=0
cc_1217 N_A_1784_97#_c_1706_n N_VPWR_c_2072_n 0.00644269f $X=10.7 $Y=1.915 $X2=0
+ $Y2=0
cc_1218 N_A_1784_97#_c_1712_n N_VPWR_c_2072_n 0.00626449f $X=9.42 $Y=2.755 $X2=0
+ $Y2=0
cc_1219 N_A_1784_97#_c_1706_n N_VPWR_c_2073_n 0.0057683f $X=10.7 $Y=1.915 $X2=0
+ $Y2=0
cc_1220 N_A_1784_97#_c_1706_n N_VPWR_c_2081_n 0.00487664f $X=10.7 $Y=1.915 $X2=0
+ $Y2=0
cc_1221 N_A_1784_97#_c_1712_n N_VPWR_c_2087_n 0.0155564f $X=9.42 $Y=2.755 $X2=0
+ $Y2=0
cc_1222 N_A_1784_97#_c_1706_n N_VPWR_c_2066_n 0.00505379f $X=10.7 $Y=1.915 $X2=0
+ $Y2=0
cc_1223 N_A_1784_97#_c_1712_n N_VPWR_c_2066_n 0.0128478f $X=9.42 $Y=2.755 $X2=0
+ $Y2=0
cc_1224 N_A_1784_97#_c_1713_n N_A_691_113#_c_2282_n 0.0138271f $X=9.405 $Y=2.53
+ $X2=0 $Y2=0
cc_1225 N_A_1784_97#_c_1712_n N_A_691_113#_c_2283_n 0.0252345f $X=9.42 $Y=2.755
+ $X2=0 $Y2=0
cc_1226 N_A_1784_97#_M1023_g N_VGND_c_2514_n 0.00193352f $X=10.9 $Y=0.69 $X2=0
+ $Y2=0
cc_1227 N_A_1784_97#_M1023_g N_VGND_c_2534_n 0.00278237f $X=10.9 $Y=0.69 $X2=0
+ $Y2=0
cc_1228 N_A_1784_97#_M1023_g N_VGND_c_2544_n 0.00363424f $X=10.9 $Y=0.69 $X2=0
+ $Y2=0
cc_1229 N_A_2489_74#_c_1802_n N_VPWR_c_2074_n 0.00634677f $X=14.415 $Y=1.765
+ $X2=0 $Y2=0
cc_1230 N_A_2489_74#_c_1811_n N_VPWR_c_2074_n 0.0121555f $X=13.24 $Y=2.75 $X2=0
+ $Y2=0
cc_1231 N_A_2489_74#_c_1802_n N_VPWR_c_2075_n 0.00322903f $X=14.415 $Y=1.765
+ $X2=0 $Y2=0
cc_1232 N_A_2489_74#_c_1804_n N_VPWR_c_2075_n 0.0106215f $X=15.425 $Y=1.765
+ $X2=0 $Y2=0
cc_1233 N_A_2489_74#_c_1805_n N_VPWR_c_2075_n 0.00127141f $X=15.875 $Y=1.765
+ $X2=0 $Y2=0
cc_1234 N_A_2489_74#_c_1804_n N_VPWR_c_2076_n 0.00127141f $X=15.425 $Y=1.765
+ $X2=0 $Y2=0
cc_1235 N_A_2489_74#_c_1805_n N_VPWR_c_2076_n 0.00959143f $X=15.875 $Y=1.765
+ $X2=0 $Y2=0
cc_1236 N_A_2489_74#_c_1811_n N_VPWR_c_2088_n 0.0184478f $X=13.24 $Y=2.75 $X2=0
+ $Y2=0
cc_1237 N_A_2489_74#_c_1802_n N_VPWR_c_2089_n 0.00445602f $X=14.415 $Y=1.765
+ $X2=0 $Y2=0
cc_1238 N_A_2489_74#_c_1804_n N_VPWR_c_2090_n 0.00413917f $X=15.425 $Y=1.765
+ $X2=0 $Y2=0
cc_1239 N_A_2489_74#_c_1805_n N_VPWR_c_2090_n 0.00413917f $X=15.875 $Y=1.765
+ $X2=0 $Y2=0
cc_1240 N_A_2489_74#_c_1802_n N_VPWR_c_2066_n 0.00863669f $X=14.415 $Y=1.765
+ $X2=0 $Y2=0
cc_1241 N_A_2489_74#_c_1804_n N_VPWR_c_2066_n 0.00414505f $X=15.425 $Y=1.765
+ $X2=0 $Y2=0
cc_1242 N_A_2489_74#_c_1805_n N_VPWR_c_2066_n 0.00414505f $X=15.875 $Y=1.765
+ $X2=0 $Y2=0
cc_1243 N_A_2489_74#_c_1811_n N_VPWR_c_2066_n 0.0152882f $X=13.24 $Y=2.75 $X2=0
+ $Y2=0
cc_1244 N_A_2489_74#_c_1804_n Q 0.00572978f $X=15.425 $Y=1.765 $X2=0 $Y2=0
cc_1245 N_A_2489_74#_M1032_g Q 0.016221f $X=15.445 $Y=0.74 $X2=0 $Y2=0
cc_1246 N_A_2489_74#_M1043_g Q 0.0145925f $X=15.875 $Y=0.74 $X2=0 $Y2=0
cc_1247 N_A_2489_74#_c_1805_n Q 0.00514983f $X=15.875 $Y=1.765 $X2=0 $Y2=0
cc_1248 N_A_2489_74#_c_1796_n Q 0.037668f $X=15.875 $Y=1.532 $X2=0 $Y2=0
cc_1249 N_A_2489_74#_c_1798_n N_VGND_M1026_d 0.00511003f $X=13.695 $Y=0.855
+ $X2=0 $Y2=0
cc_1250 N_A_2489_74#_c_1797_n N_VGND_c_2515_n 0.010811f $X=12.585 $Y=0.515 $X2=0
+ $Y2=0
cc_1251 N_A_2489_74#_c_1798_n N_VGND_c_2516_n 0.0147778f $X=13.695 $Y=0.855
+ $X2=0 $Y2=0
cc_1252 N_A_2489_74#_c_1797_n N_VGND_c_2517_n 0.00419512f $X=12.585 $Y=0.515
+ $X2=0 $Y2=0
cc_1253 N_A_2489_74#_c_1798_n N_VGND_c_2517_n 0.024775f $X=13.695 $Y=0.855 $X2=0
+ $Y2=0
cc_1254 N_A_2489_74#_M1014_g N_VGND_c_2518_n 0.00106276f $X=14.455 $Y=0.74 $X2=0
+ $Y2=0
cc_1255 N_A_2489_74#_c_1793_n N_VGND_c_2518_n 0.00393223f $X=14.53 $Y=1.465
+ $X2=0 $Y2=0
cc_1256 N_A_2489_74#_c_1798_n N_VGND_c_2518_n 0.0125741f $X=13.695 $Y=0.855
+ $X2=0 $Y2=0
cc_1257 N_A_2489_74#_c_1799_n N_VGND_c_2518_n 0.011522f $X=13.78 $Y=1.3 $X2=0
+ $Y2=0
cc_1258 N_A_2489_74#_c_1801_n N_VGND_c_2518_n 0.0210027f $X=14.33 $Y=1.465 $X2=0
+ $Y2=0
cc_1259 N_A_2489_74#_M1014_g N_VGND_c_2519_n 0.00434272f $X=14.455 $Y=0.74 $X2=0
+ $Y2=0
cc_1260 N_A_2489_74#_M1014_g N_VGND_c_2520_n 0.00413259f $X=14.455 $Y=0.74 $X2=0
+ $Y2=0
cc_1261 N_A_2489_74#_c_1792_n N_VGND_c_2520_n 0.00657295f $X=15.335 $Y=1.465
+ $X2=0 $Y2=0
cc_1262 N_A_2489_74#_M1032_g N_VGND_c_2520_n 0.00646793f $X=15.445 $Y=0.74 $X2=0
+ $Y2=0
cc_1263 N_A_2489_74#_M1032_g N_VGND_c_2521_n 0.00422942f $X=15.445 $Y=0.74 $X2=0
+ $Y2=0
cc_1264 N_A_2489_74#_M1043_g N_VGND_c_2521_n 0.00434272f $X=15.875 $Y=0.74 $X2=0
+ $Y2=0
cc_1265 N_A_2489_74#_M1043_g N_VGND_c_2522_n 0.00313962f $X=15.875 $Y=0.74 $X2=0
+ $Y2=0
cc_1266 N_A_2489_74#_c_1797_n N_VGND_c_2529_n 0.014415f $X=12.585 $Y=0.515 $X2=0
+ $Y2=0
cc_1267 N_A_2489_74#_M1014_g N_VGND_c_2541_n 0.005596f $X=14.455 $Y=0.74 $X2=0
+ $Y2=0
cc_1268 N_A_2489_74#_M1014_g N_VGND_c_2544_n 0.00830035f $X=14.455 $Y=0.74 $X2=0
+ $Y2=0
cc_1269 N_A_2489_74#_M1032_g N_VGND_c_2544_n 0.00788596f $X=15.445 $Y=0.74 $X2=0
+ $Y2=0
cc_1270 N_A_2489_74#_M1043_g N_VGND_c_2544_n 0.00820382f $X=15.875 $Y=0.74 $X2=0
+ $Y2=0
cc_1271 N_A_2489_74#_c_1797_n N_VGND_c_2544_n 0.0119404f $X=12.585 $Y=0.515
+ $X2=0 $Y2=0
cc_1272 N_A_2489_74#_c_1798_n N_VGND_c_2544_n 0.0209551f $X=13.695 $Y=0.855
+ $X2=0 $Y2=0
cc_1273 N_A_2489_74#_c_1798_n A_2591_74# 0.0023798f $X=13.695 $Y=0.855 $X2=-0.19
+ $Y2=-0.245
cc_1274 N_A_32_74#_c_1953_n A_132_464# 0.00595227f $X=1.485 $Y=2.375 $X2=-0.19
+ $Y2=-0.245
cc_1275 N_A_32_74#_c_1953_n N_VPWR_M1029_d 0.00509381f $X=1.485 $Y=2.375
+ $X2=-0.19 $Y2=-0.245
cc_1276 N_A_32_74#_c_1955_n N_VPWR_M1017_d 4.29284e-19 $X=2.165 $Y=2.99 $X2=0
+ $Y2=0
cc_1277 N_A_32_74#_c_1987_n N_VPWR_M1017_d 0.00490162f $X=2.25 $Y=2.905 $X2=0
+ $Y2=0
cc_1278 N_A_32_74#_c_1957_n N_VPWR_M1017_d 0.00977001f $X=3.265 $Y=2.375 $X2=0
+ $Y2=0
cc_1279 N_A_32_74#_c_1952_n N_VPWR_c_2067_n 0.0101952f $X=0.36 $Y=2.465 $X2=0
+ $Y2=0
cc_1280 N_A_32_74#_c_1953_n N_VPWR_c_2067_n 0.0154248f $X=1.485 $Y=2.375 $X2=0
+ $Y2=0
cc_1281 N_A_32_74#_c_1954_n N_VPWR_c_2067_n 0.0208967f $X=1.57 $Y=2.905 $X2=0
+ $Y2=0
cc_1282 N_A_32_74#_c_1956_n N_VPWR_c_2067_n 0.0146662f $X=1.655 $Y=2.99 $X2=0
+ $Y2=0
cc_1283 N_A_32_74#_c_1955_n N_VPWR_c_2068_n 0.0146002f $X=2.165 $Y=2.99 $X2=0
+ $Y2=0
cc_1284 N_A_32_74#_c_1987_n N_VPWR_c_2068_n 0.0205316f $X=2.25 $Y=2.905 $X2=0
+ $Y2=0
cc_1285 N_A_32_74#_c_1957_n N_VPWR_c_2068_n 0.0154248f $X=3.265 $Y=2.375 $X2=0
+ $Y2=0
cc_1286 N_A_32_74#_c_1961_n N_VPWR_c_2068_n 0.0100549f $X=3.43 $Y=2.455 $X2=0
+ $Y2=0
cc_1287 N_A_32_74#_c_1952_n N_VPWR_c_2083_n 0.0195149f $X=0.36 $Y=2.465 $X2=0
+ $Y2=0
cc_1288 N_A_32_74#_c_1955_n N_VPWR_c_2084_n 0.0445209f $X=2.165 $Y=2.99 $X2=0
+ $Y2=0
cc_1289 N_A_32_74#_c_1956_n N_VPWR_c_2084_n 0.0121867f $X=1.655 $Y=2.99 $X2=0
+ $Y2=0
cc_1290 N_A_32_74#_c_1961_n N_VPWR_c_2085_n 0.0118846f $X=3.43 $Y=2.455 $X2=0
+ $Y2=0
cc_1291 N_A_32_74#_c_1952_n N_VPWR_c_2066_n 0.0161142f $X=0.36 $Y=2.465 $X2=0
+ $Y2=0
cc_1292 N_A_32_74#_c_1955_n N_VPWR_c_2066_n 0.0256906f $X=2.165 $Y=2.99 $X2=0
+ $Y2=0
cc_1293 N_A_32_74#_c_1956_n N_VPWR_c_2066_n 0.00660921f $X=1.655 $Y=2.99 $X2=0
+ $Y2=0
cc_1294 N_A_32_74#_c_1961_n N_VPWR_c_2066_n 0.0101938f $X=3.43 $Y=2.455 $X2=0
+ $Y2=0
cc_1295 N_A_32_74#_c_1957_n A_578_462# 0.0048076f $X=3.265 $Y=2.375 $X2=-0.19
+ $Y2=-0.245
cc_1296 N_A_32_74#_c_1961_n N_A_691_113#_c_2274_n 0.00699177f $X=3.43 $Y=2.455
+ $X2=0 $Y2=0
cc_1297 N_A_32_74#_c_1961_n N_A_691_113#_c_2286_n 0.00351237f $X=3.43 $Y=2.455
+ $X2=0 $Y2=0
cc_1298 N_A_32_74#_c_1947_n N_A_691_113#_c_2271_n 0.0188786f $X=3.165 $Y=0.775
+ $X2=0 $Y2=0
cc_1299 N_A_32_74#_c_1950_n N_A_691_113#_c_2271_n 0.00333703f $X=3.46 $Y=1.26
+ $X2=0 $Y2=0
cc_1300 N_A_32_74#_c_1947_n N_A_691_113#_c_2272_n 0.00645754f $X=3.165 $Y=0.775
+ $X2=0 $Y2=0
cc_1301 N_A_32_74#_c_1948_n N_A_691_113#_c_2272_n 0.0697173f $X=3.46 $Y=2.29
+ $X2=0 $Y2=0
cc_1302 N_A_32_74#_c_1950_n N_A_691_113#_c_2272_n 0.0136555f $X=3.46 $Y=1.26
+ $X2=0 $Y2=0
cc_1303 N_A_32_74#_c_1949_n N_VGND_c_2509_n 0.0100909f $X=0.415 $Y=0.585 $X2=0
+ $Y2=0
cc_1304 N_A_32_74#_c_1947_n N_VGND_c_2510_n 0.0145731f $X=3.165 $Y=0.775 $X2=0
+ $Y2=0
cc_1305 N_A_32_74#_c_1949_n N_VGND_c_2530_n 0.0149954f $X=0.415 $Y=0.585 $X2=0
+ $Y2=0
cc_1306 N_A_32_74#_c_1947_n N_VGND_c_2531_n 0.00794834f $X=3.165 $Y=0.775 $X2=0
+ $Y2=0
cc_1307 N_A_32_74#_c_1947_n N_VGND_c_2544_n 0.0105391f $X=3.165 $Y=0.775 $X2=0
+ $Y2=0
cc_1308 N_A_32_74#_c_1949_n N_VGND_c_2544_n 0.0168506f $X=0.415 $Y=0.585 $X2=0
+ $Y2=0
cc_1309 N_VPWR_c_2069_n N_A_691_113#_c_2275_n 0.0148243f $X=5.13 $Y=2.76 $X2=0
+ $Y2=0
cc_1310 N_VPWR_c_2085_n N_A_691_113#_c_2275_n 0.0567624f $X=5.035 $Y=3.33 $X2=0
+ $Y2=0
cc_1311 N_VPWR_c_2066_n N_A_691_113#_c_2275_n 0.0303734f $X=17.04 $Y=3.33 $X2=0
+ $Y2=0
cc_1312 N_VPWR_c_2085_n N_A_691_113#_c_2286_n 0.0170104f $X=5.035 $Y=3.33 $X2=0
+ $Y2=0
cc_1313 N_VPWR_c_2066_n N_A_691_113#_c_2286_n 0.00854122f $X=17.04 $Y=3.33 $X2=0
+ $Y2=0
cc_1314 N_VPWR_M1045_d N_A_691_113#_c_2302_n 0.00528719f $X=4.75 $Y=2.265 $X2=0
+ $Y2=0
cc_1315 N_VPWR_c_2069_n N_A_691_113#_c_2302_n 0.0232873f $X=5.13 $Y=2.76 $X2=0
+ $Y2=0
cc_1316 N_VPWR_M1045_d N_A_691_113#_c_2276_n 0.0101647f $X=4.75 $Y=2.265 $X2=0
+ $Y2=0
cc_1317 N_VPWR_c_2069_n N_A_691_113#_c_2276_n 0.017052f $X=5.13 $Y=2.76 $X2=0
+ $Y2=0
cc_1318 N_VPWR_M1007_s N_A_691_113#_c_2267_n 0.00613089f $X=6.425 $Y=1.84 $X2=0
+ $Y2=0
cc_1319 N_VPWR_M1007_s N_A_691_113#_c_2279_n 0.00635059f $X=6.425 $Y=1.84 $X2=0
+ $Y2=0
cc_1320 N_VPWR_M1001_s N_A_691_113#_c_2279_n 0.00250916f $X=7.815 $Y=1.84 $X2=0
+ $Y2=0
cc_1321 N_VPWR_c_2070_n N_A_691_113#_c_2279_n 0.0150987f $X=6.57 $Y=2.815 $X2=0
+ $Y2=0
cc_1322 N_VPWR_c_2071_n N_A_691_113#_c_2279_n 0.00870407f $X=7.96 $Y=2.815 $X2=0
+ $Y2=0
cc_1323 N_VPWR_c_2066_n N_A_691_113#_c_2279_n 0.0368914f $X=17.04 $Y=3.33 $X2=0
+ $Y2=0
cc_1324 N_VPWR_M1007_s N_A_691_113#_c_2280_n 0.00259343f $X=6.425 $Y=1.84 $X2=0
+ $Y2=0
cc_1325 N_VPWR_c_2069_n N_A_691_113#_c_2280_n 0.00972078f $X=5.13 $Y=2.76 $X2=0
+ $Y2=0
cc_1326 N_VPWR_c_2070_n N_A_691_113#_c_2280_n 0.0217988f $X=6.57 $Y=2.815 $X2=0
+ $Y2=0
cc_1327 N_VPWR_c_2079_n N_A_691_113#_c_2280_n 0.0167396f $X=6.485 $Y=3.33 $X2=0
+ $Y2=0
cc_1328 N_VPWR_c_2066_n N_A_691_113#_c_2280_n 0.0229958f $X=17.04 $Y=3.33 $X2=0
+ $Y2=0
cc_1329 N_VPWR_M1001_s N_A_691_113#_c_2281_n 0.0114611f $X=7.815 $Y=1.84 $X2=0
+ $Y2=0
cc_1330 N_VPWR_c_2071_n N_A_691_113#_c_2295_n 0.00100191f $X=7.96 $Y=2.815 $X2=0
+ $Y2=0
cc_1331 N_VPWR_c_2066_n N_A_691_113#_c_2295_n 0.00503485f $X=17.04 $Y=3.33 $X2=0
+ $Y2=0
cc_1332 N_VPWR_c_2087_n N_A_691_113#_c_2282_n 0.00557176f $X=10.225 $Y=3.33
+ $X2=0 $Y2=0
cc_1333 N_VPWR_c_2066_n N_A_691_113#_c_2282_n 0.00937585f $X=17.04 $Y=3.33 $X2=0
+ $Y2=0
cc_1334 N_VPWR_c_2087_n N_A_691_113#_c_2283_n 0.0108228f $X=10.225 $Y=3.33 $X2=0
+ $Y2=0
cc_1335 N_VPWR_c_2066_n N_A_691_113#_c_2283_n 0.00906589f $X=17.04 $Y=3.33 $X2=0
+ $Y2=0
cc_1336 N_VPWR_M1001_s N_A_691_113#_c_2438_n 0.00184106f $X=7.815 $Y=1.84 $X2=0
+ $Y2=0
cc_1337 N_VPWR_c_2071_n N_A_691_113#_c_2438_n 0.0129915f $X=7.96 $Y=2.815 $X2=0
+ $Y2=0
cc_1338 N_VPWR_c_2066_n N_A_691_113#_c_2438_n 6.0606e-19 $X=17.04 $Y=3.33 $X2=0
+ $Y2=0
cc_1339 N_VPWR_c_2087_n N_A_691_113#_c_2375_n 0.00263412f $X=10.225 $Y=3.33
+ $X2=0 $Y2=0
cc_1340 N_VPWR_c_2066_n N_A_691_113#_c_2375_n 0.00477661f $X=17.04 $Y=3.33 $X2=0
+ $Y2=0
cc_1341 N_VPWR_M1038_s N_Q_N_c_2477_n 0.00329576f $X=16.85 $Y=1.84 $X2=0 $Y2=0
cc_1342 N_VPWR_c_2078_n N_Q_N_c_2477_n 0.0219924f $X=17 $Y=2.25 $X2=0 $Y2=0
cc_1343 N_VPWR_c_2076_n Q_N 0.015063f $X=16.1 $Y=2.78 $X2=0 $Y2=0
cc_1344 N_VPWR_c_2078_n Q_N 0.034387f $X=17 $Y=2.25 $X2=0 $Y2=0
cc_1345 N_VPWR_c_2091_n Q_N 0.0115612f $X=16.835 $Y=3.33 $X2=0 $Y2=0
cc_1346 N_VPWR_c_2066_n Q_N 0.00856962f $X=17.04 $Y=3.33 $X2=0 $Y2=0
cc_1347 N_A_691_113#_c_2276_n A_1088_453# 0.00595227f $X=5.845 $Y=2.34 $X2=-0.19
+ $Y2=-0.245
cc_1348 N_A_691_113#_c_2273_n N_VGND_M1035_s 7.58458e-19 $X=6.39 $Y=1.175 $X2=0
+ $Y2=0
cc_1349 N_A_691_113#_c_2266_n N_VGND_c_2511_n 0.00634222f $X=5.985 $Y=0.835
+ $X2=0 $Y2=0
cc_1350 N_A_691_113#_c_2266_n N_VGND_c_2512_n 0.0192622f $X=5.985 $Y=0.835 $X2=0
+ $Y2=0
cc_1351 N_A_691_113#_c_2273_n N_VGND_c_2512_n 0.00485909f $X=6.39 $Y=1.175 $X2=0
+ $Y2=0
cc_1352 N_A_691_113#_c_2271_n N_VGND_c_2531_n 0.00932016f $X=3.665 $Y=0.775
+ $X2=0 $Y2=0
cc_1353 N_A_691_113#_c_2266_n N_VGND_c_2532_n 0.00684598f $X=5.985 $Y=0.835
+ $X2=0 $Y2=0
cc_1354 N_A_691_113#_c_2266_n N_VGND_c_2544_n 0.00989908f $X=5.985 $Y=0.835
+ $X2=0 $Y2=0
cc_1355 N_A_691_113#_c_2271_n N_VGND_c_2544_n 0.0122951f $X=3.665 $Y=0.775 $X2=0
+ $Y2=0
cc_1356 Q N_VGND_c_2520_n 0.0309174f $X=15.515 $Y=0.47 $X2=0 $Y2=0
cc_1357 Q N_VGND_c_2521_n 0.0149085f $X=15.515 $Y=0.47 $X2=0 $Y2=0
cc_1358 Q N_VGND_c_2522_n 0.0294574f $X=15.515 $Y=0.47 $X2=0 $Y2=0
cc_1359 Q N_VGND_c_2544_n 0.0122037f $X=15.515 $Y=0.47 $X2=0 $Y2=0
cc_1360 N_Q_N_c_2476_n N_VGND_M1041_s 0.00328964f $X=16.932 $Y=1.13 $X2=0 $Y2=0
cc_1361 N_Q_N_c_2476_n N_VGND_c_2522_n 0.00741094f $X=16.932 $Y=1.13 $X2=0 $Y2=0
cc_1362 Q_N N_VGND_c_2522_n 0.0225498f $X=16.475 $Y=0.47 $X2=0 $Y2=0
cc_1363 N_Q_N_c_2476_n N_VGND_c_2524_n 0.0201545f $X=16.932 $Y=1.13 $X2=0 $Y2=0
cc_1364 Q_N N_VGND_c_2524_n 0.0172723f $X=16.475 $Y=0.47 $X2=0 $Y2=0
cc_1365 Q_N N_VGND_c_2535_n 0.014379f $X=16.475 $Y=0.47 $X2=0 $Y2=0
cc_1366 Q_N N_VGND_c_2544_n 0.0118382f $X=16.475 $Y=0.47 $X2=0 $Y2=0
