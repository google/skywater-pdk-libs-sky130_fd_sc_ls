* File: sky130_fd_sc_ls__sdlclkp_4.spice
* Created: Wed Sep  2 11:29:03 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__sdlclkp_4.pex.spice"
.subckt sky130_fd_sc_ls__sdlclkp_4  VNB VPB SCE GATE CLK VPWR GCLK VGND
* 
* VGND	VGND
* GCLK	GCLK
* VPWR	VPWR
* CLK	CLK
* GATE	GATE
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1019 N_A_119_143#_M1019_d N_SCE_M1019_g N_VGND_M1019_s VNB NSHORT L=0.15
+ W=0.55 AD=0.089375 AS=0.1705 PD=0.875 PS=1.72 NRD=9.816 NRS=5.448 M=1
+ R=3.66667 SA=75000.2 SB=75001.4 A=0.0825 P=1.4 MULT=1
MM1025 N_VGND_M1025_d N_GATE_M1025_g N_A_119_143#_M1019_d VNB NSHORT L=0.15
+ W=0.55 AD=0.233963 AS=0.089375 PD=1.43256 PS=0.875 NRD=80.808 NRS=0 M=1
+ R=3.66667 SA=75000.7 SB=75000.9 A=0.0825 P=1.4 MULT=1
MM1017 N_A_354_105#_M1017_d N_A_324_79#_M1017_g N_VGND_M1025_d VNB NSHORT L=0.15
+ W=0.74 AD=0.2109 AS=0.314787 PD=2.05 PS=1.92744 NRD=0 NRS=60.06 M=1 R=4.93333
+ SA=75001.2 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1022 N_A_634_74#_M1022_d N_A_324_79#_M1022_g N_A_119_143#_M1022_s VNB NSHORT
+ L=0.15 W=0.55 AD=0.119214 AS=0.38225 PD=1.07732 PS=2.49 NRD=4.356 NRS=77.448
+ M=1 R=3.66667 SA=75000.6 SB=75001.6 A=0.0825 P=1.4 MULT=1
MM1016 A_744_74# N_A_354_105#_M1016_g N_A_634_74#_M1022_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.0910361 PD=0.66 PS=0.82268 NRD=18.564 NRS=30 M=1 R=2.8
+ SA=75001.2 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1005_d N_A_792_48#_M1005_g A_744_74# VNB NSHORT L=0.15 W=0.42
+ AD=0.136934 AS=0.0504 PD=1.05 PS=0.66 NRD=5.712 NRS=18.564 M=1 R=2.8
+ SA=75001.6 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1004 N_A_792_48#_M1004_d N_A_634_74#_M1004_g N_VGND_M1005_d VNB NSHORT L=0.15
+ W=0.74 AD=0.2109 AS=0.241266 PD=2.05 PS=1.85 NRD=0 NRS=66.48 M=1 R=4.93333
+ SA=75001.4 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1011 N_VGND_M1011_d N_CLK_M1011_g N_A_324_79#_M1011_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1295 AS=0.2109 PD=1.09 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1007 A_1292_74# N_CLK_M1007_g N_VGND_M1011_d VNB NSHORT L=0.15 W=0.74
+ AD=0.0888 AS=0.1295 PD=0.98 PS=1.09 NRD=10.536 NRS=0 M=1 R=4.93333 SA=75000.7
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1008 N_A_1289_368#_M1008_d N_A_792_48#_M1008_g A_1292_74# VNB NSHORT L=0.15
+ W=0.74 AD=0.2109 AS=0.0888 PD=2.05 PS=0.98 NRD=0 NRS=10.536 M=1 R=4.93333
+ SA=75001.1 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1001 N_VGND_M1001_d N_A_1289_368#_M1001_g N_GCLK_M1001_s VNB NSHORT L=0.15
+ W=0.74 AD=0.2109 AS=0.1221 PD=2.05 PS=1.07 NRD=0 NRS=8.1 M=1 R=4.93333
+ SA=75000.2 SB=75001.6 A=0.111 P=1.78 MULT=1
MM1013 N_VGND_M1013_d N_A_1289_368#_M1013_g N_GCLK_M1001_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1221 PD=1.02 PS=1.07 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.7 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1026 N_VGND_M1013_d N_A_1289_368#_M1026_g N_GCLK_M1026_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.1 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1027 N_VGND_M1027_d N_A_1289_368#_M1027_g N_GCLK_M1026_s VNB NSHORT L=0.15
+ W=0.74 AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1009 A_116_395# N_SCE_M1009_g N_VPWR_M1009_s VPB PHIGHVT L=0.15 W=0.84
+ AD=0.1134 AS=0.2478 PD=1.11 PS=2.27 NRD=18.7544 NRS=2.3443 M=1 R=5.6
+ SA=75000.2 SB=75000.6 A=0.126 P=1.98 MULT=1
MM1020 N_A_119_143#_M1020_d N_GATE_M1020_g A_116_395# VPB PHIGHVT L=0.15 W=0.84
+ AD=0.2478 AS=0.1134 PD=2.27 PS=1.11 NRD=2.3443 NRS=18.7544 M=1 R=5.6
+ SA=75000.6 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1002 N_A_354_105#_M1002_d N_A_324_79#_M1002_g N_VPWR_M1002_s VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.4033 AS=0.4872 PD=3.02 PS=2.84 NRD=99.682 NRS=3.5066 M=1
+ R=5.6 SA=75000.5 SB=75000.3 A=0.126 P=1.98 MULT=1
MM1014 N_A_634_74#_M1014_d N_A_354_105#_M1014_g N_A_119_143#_M1014_s VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.1904 AS=0.2478 PD=1.63333 PS=2.27 NRD=2.3443 NRS=2.3443 M=1
+ R=5.6 SA=75000.2 SB=75001 A=0.126 P=1.98 MULT=1
MM1012 A_785_455# N_A_324_79#_M1012_g N_A_634_74#_M1014_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0567 AS=0.0952 PD=0.69 PS=0.816667 NRD=37.5088 NRS=44.5417 M=1
+ R=2.8 SA=75000.8 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1006 N_VPWR_M1006_d N_A_792_48#_M1006_g A_785_455# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.102136 AS=0.0567 PD=0.829091 PS=0.69 NRD=53.9386 NRS=37.5088 M=1 R=2.8
+ SA=75001.2 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1000 N_A_792_48#_M1000_d N_A_634_74#_M1000_g N_VPWR_M1006_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.3304 AS=0.272364 PD=2.83 PS=2.21091 NRD=1.7533 NRS=1.7533 M=1
+ R=7.46667 SA=75000.8 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1023 N_VPWR_M1023_d N_CLK_M1023_g N_A_324_79#_M1023_s VPB PHIGHVT L=0.15
+ W=0.84 AD=0.174 AS=0.252 PD=1.29 PS=2.28 NRD=35.6767 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75003.5 A=0.126 P=1.98 MULT=1
MM1015 N_A_1289_368#_M1015_d N_CLK_M1015_g N_VPWR_M1023_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.2772 AS=0.232 PD=1.615 PS=1.72 NRD=36.051 NRS=1.7533 M=1 R=7.46667
+ SA=75000.6 SB=75002.9 A=0.168 P=2.54 MULT=1
MM1018 N_VPWR_M1018_d N_A_792_48#_M1018_g N_A_1289_368#_M1015_d VPB PHIGHVT
+ L=0.15 W=1.12 AD=0.196 AS=0.2772 PD=1.47 PS=1.615 NRD=10.5395 NRS=1.7533 M=1
+ R=7.46667 SA=75001.3 SB=75002.3 A=0.168 P=2.54 MULT=1
MM1003 N_GCLK_M1003_d N_A_1289_368#_M1003_g N_VPWR_M1018_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.2408 AS=0.196 PD=1.55 PS=1.47 NRD=24.6053 NRS=1.7533 M=1 R=7.46667
+ SA=75001.8 SB=75001.8 A=0.168 P=2.54 MULT=1
MM1010 N_GCLK_M1003_d N_A_1289_368#_M1010_g N_VPWR_M1010_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.2408 AS=0.196 PD=1.55 PS=1.47 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.3 SB=75001.2 A=0.168 P=2.54 MULT=1
MM1021 N_GCLK_M1021_d N_A_1289_368#_M1021_g N_VPWR_M1010_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.1932 AS=0.196 PD=1.465 PS=1.47 NRD=1.7533 NRS=10.5395 M=1
+ R=7.46667 SA=75002.8 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1024 N_GCLK_M1021_d N_A_1289_368#_M1024_g N_VPWR_M1024_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.1932 AS=0.336 PD=1.465 PS=2.84 NRD=9.6727 NRS=2.6201 M=1 R=7.46667
+ SA=75003.3 SB=75000.2 A=0.168 P=2.54 MULT=1
DX28_noxref VNB VPB NWDIODE A=18.6851 P=23.85
*
.include "sky130_fd_sc_ls__sdlclkp_4.pxi.spice"
*
.ends
*
*
