* File: sky130_fd_sc_ls__mux4_4.spice
* Created: Fri Aug 28 13:31:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__mux4_4.pex.spice"
.subckt sky130_fd_sc_ls__mux4_4  VNB VPB A1 A0 S0 A2 A3 S1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* S1	S1
* A3	A3
* A2	A2
* S0	S0
* A0	A0
* A1	A1
* VPB	VPB
* VNB	VNB
MM1025 N_VGND_M1025_d N_A1_M1025_g N_A_114_126#_M1025_s VNB NSHORT L=0.15 W=0.64
+ AD=0.1824 AS=0.0896 PD=1.85 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75001.6 A=0.096 P=1.58 MULT=1
MM1028 N_VGND_M1028_d N_A1_M1028_g N_A_114_126#_M1025_s VNB NSHORT L=0.15 W=0.64
+ AD=0.1104 AS=0.0896 PD=0.985 PS=0.92 NRD=5.616 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75001.2 A=0.096 P=1.58 MULT=1
MM1021 N_A_299_126#_M1021_d N_A0_M1021_g N_VGND_M1028_d VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.1104 PD=0.92 PS=0.985 NRD=0 NRS=6.552 M=1 R=4.26667 SA=75001.1
+ SB=75000.7 A=0.096 P=1.58 MULT=1
MM1022 N_A_299_126#_M1021_d N_A0_M1022_g N_VGND_M1022_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.3525 PD=0.92 PS=2.83 NRD=0 NRS=92.952 M=1 R=4.26667 SA=75001.6
+ SB=75000.3 A=0.096 P=1.58 MULT=1
MM1004 N_A_509_392#_M1004_d N_S0_M1004_g N_A_114_126#_M1004_s VNB NSHORT L=0.15
+ W=0.64 AD=0.31625 AS=0.104 PD=2.58 PS=0.965 NRD=82.332 NRS=0 M=1 R=4.26667
+ SA=75000.3 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1047 N_A_509_392#_M1047_d N_S0_M1047_g N_A_114_126#_M1004_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.104 PD=0.92 PS=0.965 NRD=0 NRS=8.436 M=1 R=4.26667
+ SA=75000.8 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1036 N_A_299_126#_M1036_d N_A_758_306#_M1036_g N_A_509_392#_M1047_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.2 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1042 N_A_299_126#_M1036_d N_A_758_306#_M1042_g N_A_509_392#_M1042_s VNB NSHORT
+ L=0.15 W=0.64 AD=0.0896 AS=0.1824 PD=0.92 PS=1.85 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.6 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1012 N_VGND_M1012_d N_S0_M1012_g N_A_758_306#_M1012_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.2109 PD=2.05 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1002 N_A_1191_121#_M1002_d N_A_758_306#_M1002_g N_A_1278_121#_M1002_s VNB
+ NSHORT L=0.15 W=0.64 AD=0.1824 AS=0.0896 PD=1.85 PS=0.92 NRD=0 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1051 N_A_1191_121#_M1051_d N_A_758_306#_M1051_g N_A_1278_121#_M1002_s VNB
+ NSHORT L=0.15 W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1
+ R=4.26667 SA=75000.6 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1006 N_A_1450_121#_M1006_d N_S0_M1006_g N_A_1191_121#_M1051_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.1 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1040 N_A_1450_121#_M1006_d N_S0_M1040_g N_A_1191_121#_M1040_s VNB NSHORT
+ L=0.15 W=0.64 AD=0.0896 AS=0.2336 PD=0.92 PS=2.01 NRD=0 NRS=14.988 M=1
+ R=4.26667 SA=75001.5 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1018 N_A_1278_121#_M1018_d N_A2_M1018_g N_VGND_M1018_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.2887 PD=0.92 PS=2.39 NRD=0 NRS=74.256 M=1 R=4.26667
+ SA=75000.3 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1038 N_A_1278_121#_M1018_d N_A2_M1038_g N_VGND_M1038_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.7 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1014 N_A_1450_121#_M1014_d N_A3_M1014_g N_VGND_M1038_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.1 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1027 N_A_1450_121#_M1014_d N_A3_M1027_g N_VGND_M1027_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.1824 PD=0.92 PS=1.85 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.6 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1013 N_A_1191_121#_M1013_d N_S1_M1013_g N_A_2199_74#_M1013_s VNB NSHORT L=0.15
+ W=0.64 AD=0.166175 AS=0.1824 PD=1.255 PS=1.85 NRD=38.364 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75002.1 A=0.096 P=1.58 MULT=1
MM1015 N_A_1191_121#_M1013_d N_S1_M1015_g N_A_2199_74#_M1015_s VNB NSHORT L=0.15
+ W=0.64 AD=0.166175 AS=0.224 PD=1.255 PS=1.34 NRD=38.364 NRS=0 M=1 R=4.26667
+ SA=75000.8 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1009 N_A_2199_74#_M1015_s N_A_2489_347#_M1009_g N_A_509_392#_M1009_s VNB
+ NSHORT L=0.15 W=0.64 AD=0.224 AS=0.0896 PD=1.34 PS=0.92 NRD=13.116 NRS=0 M=1
+ R=4.26667 SA=75001.6 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1048 N_A_2199_74#_M1048_d N_A_2489_347#_M1048_g N_A_509_392#_M1009_s VNB
+ NSHORT L=0.15 W=0.64 AD=0.2272 AS=0.0896 PD=1.99 PS=0.92 NRD=6.552 NRS=0 M=1
+ R=4.26667 SA=75002.1 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1010 N_VGND_M1010_d N_S1_M1010_g N_A_2489_347#_M1010_s VNB NSHORT L=0.15
+ W=0.74 AD=0.2146 AS=0.2109 PD=1.32 PS=2.05 NRD=48.648 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75002.2 A=0.111 P=1.78 MULT=1
MM1016 N_X_M1016_d N_A_2199_74#_M1016_g N_VGND_M1010_d VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.2146 PD=1.02 PS=1.32 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.9
+ SB=75001.5 A=0.111 P=1.78 MULT=1
MM1026 N_X_M1016_d N_A_2199_74#_M1026_g N_VGND_M1026_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.4
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1029 N_X_M1029_d N_A_2199_74#_M1029_g N_VGND_M1026_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.8
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1050 N_X_M1029_d N_A_2199_74#_M1050_g N_VGND_M1050_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1039 N_VPWR_M1039_d N_A1_M1039_g N_A_116_392#_M1039_s VPB PHIGHVT L=0.15 W=1
+ AD=0.295 AS=0.15 PD=2.59 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75000.2
+ SB=75001.6 A=0.15 P=2.3 MULT=1
MM1041 N_VPWR_M1041_d N_A1_M1041_g N_A_116_392#_M1039_s VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75000.7
+ SB=75001.2 A=0.15 P=2.3 MULT=1
MM1000 N_A_296_392#_M1000_d N_A0_M1000_g N_VPWR_M1041_d VPB PHIGHVT L=0.15 W=1
+ AD=0.175 AS=0.15 PD=1.35 PS=1.3 NRD=11.8003 NRS=1.9503 M=1 R=6.66667
+ SA=75001.1 SB=75000.7 A=0.15 P=2.3 MULT=1
MM1008 N_A_296_392#_M1000_d N_A0_M1008_g N_VPWR_M1008_s VPB PHIGHVT L=0.15 W=1
+ AD=0.175 AS=0.295 PD=1.35 PS=2.59 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75001.6 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1003 N_A_296_392#_M1003_d N_S0_M1003_g N_A_509_392#_M1003_s VPB PHIGHVT L=0.15
+ W=1 AD=0.1625 AS=0.31 PD=1.325 PS=2.62 NRD=1.9503 NRS=3.9203 M=1 R=6.66667
+ SA=75000.2 SB=75001.6 A=0.15 P=2.3 MULT=1
MM1043 N_A_296_392#_M1003_d N_S0_M1043_g N_A_509_392#_M1043_s VPB PHIGHVT L=0.15
+ W=1 AD=0.1625 AS=0.1625 PD=1.325 PS=1.325 NRD=6.8753 NRS=6.8753 M=1 R=6.66667
+ SA=75000.7 SB=75001.1 A=0.15 P=2.3 MULT=1
MM1023 N_A_116_392#_M1023_d N_A_758_306#_M1023_g N_A_509_392#_M1043_s VPB
+ PHIGHVT L=0.15 W=1 AD=0.15 AS=0.1625 PD=1.3 PS=1.325 NRD=1.9503 NRS=1.9503 M=1
+ R=6.66667 SA=75001.2 SB=75000.7 A=0.15 P=2.3 MULT=1
MM1035 N_A_116_392#_M1023_d N_A_758_306#_M1035_g N_A_509_392#_M1035_s VPB
+ PHIGHVT L=0.15 W=1 AD=0.15 AS=0.295 PD=1.3 PS=2.59 NRD=1.9503 NRS=1.9503 M=1
+ R=6.66667 SA=75001.6 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1030 N_VPWR_M1030_d N_S0_M1030_g N_A_758_306#_M1030_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.3304 AS=0.3304 PD=2.83 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1019 N_A_1285_377#_M1019_d N_A_758_306#_M1019_g N_A_1191_121#_M1019_s VPB
+ PHIGHVT L=0.15 W=1 AD=0.15 AS=0.295 PD=1.3 PS=2.59 NRD=1.9503 NRS=1.9503 M=1
+ R=6.66667 SA=75000.2 SB=75001.6 A=0.15 P=2.3 MULT=1
MM1031 N_A_1285_377#_M1019_d N_A_758_306#_M1031_g N_A_1191_121#_M1031_s VPB
+ PHIGHVT L=0.15 W=1 AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1
+ R=6.66667 SA=75000.7 SB=75001.1 A=0.15 P=2.3 MULT=1
MM1005 N_A_1191_121#_M1031_s N_S0_M1005_g N_A_1465_377#_M1005_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75001.1 SB=75000.7 A=0.15 P=2.3 MULT=1
MM1045 N_A_1191_121#_M1045_d N_S0_M1045_g N_A_1465_377#_M1005_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.295 AS=0.15 PD=2.59 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75001.6 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1007 N_A_1465_377#_M1007_d N_A2_M1007_g N_VPWR_M1007_s VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.44815 PD=1.3 PS=3.23 NRD=1.9503 NRS=77.4407 M=1 R=6.66667
+ SA=75000.3 SB=75001.7 A=0.15 P=2.3 MULT=1
MM1017 N_A_1465_377#_M1007_d N_A2_M1017_g N_VPWR_M1017_s VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.27525 PD=1.3 PS=1.715 NRD=1.9503 NRS=43.3794 M=1 R=6.66667
+ SA=75000.8 SB=75001.3 A=0.15 P=2.3 MULT=1
MM1033 N_VPWR_M1017_s N_A3_M1033_g N_A_1285_377#_M1033_s VPB PHIGHVT L=0.15 W=1
+ AD=0.27525 AS=0.15 PD=1.715 PS=1.3 NRD=43.3794 NRS=1.9503 M=1 R=6.66667
+ SA=75001.4 SB=75000.7 A=0.15 P=2.3 MULT=1
MM1046 N_VPWR_M1046_d N_A3_M1046_g N_A_1285_377#_M1033_s VPB PHIGHVT L=0.15 W=1
+ AD=0.295 AS=0.15 PD=2.59 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75001.8
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1001 N_A_2199_74#_M1001_d N_S1_M1001_g N_A_509_392#_M1001_s VPB PHIGHVT L=0.15
+ W=1 AD=0.295 AS=0.175 PD=2.59 PS=1.35 NRD=1.9503 NRS=11.8003 M=1 R=6.66667
+ SA=75000.2 SB=75001.8 A=0.15 P=2.3 MULT=1
MM1044 N_A_2199_74#_M1044_d N_S1_M1044_g N_A_509_392#_M1001_s VPB PHIGHVT L=0.15
+ W=1 AD=0.175 AS=0.175 PD=1.35 PS=1.35 NRD=11.8003 NRS=1.9503 M=1 R=6.66667
+ SA=75000.7 SB=75001.3 A=0.15 P=2.3 MULT=1
MM1011 N_A_1191_121#_M1011_d N_A_2489_347#_M1011_g N_A_2199_74#_M1044_d VPB
+ PHIGHVT L=0.15 W=1 AD=0.175 AS=0.175 PD=1.35 PS=1.35 NRD=11.8003 NRS=1.9503
+ M=1 R=6.66667 SA=75001.2 SB=75000.8 A=0.15 P=2.3 MULT=1
MM1020 N_A_1191_121#_M1011_d N_A_2489_347#_M1020_g N_A_2199_74#_M1020_s VPB
+ PHIGHVT L=0.15 W=1 AD=0.175 AS=0.345 PD=1.35 PS=2.69 NRD=1.9503 NRS=11.8003
+ M=1 R=6.66667 SA=75001.7 SB=75000.3 A=0.15 P=2.3 MULT=1
MM1037 N_VPWR_M1037_d N_S1_M1037_g N_A_2489_347#_M1037_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.2044 AS=0.3696 PD=1.485 PS=2.9 NRD=4.3931 NRS=7.8997 M=1 R=7.46667
+ SA=75000.3 SB=75002.2 A=0.168 P=2.54 MULT=1
MM1024 N_VPWR_M1037_d N_A_2199_74#_M1024_g N_X_M1024_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.2044 AS=0.168 PD=1.485 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75000.8 SB=75001.7 A=0.168 P=2.54 MULT=1
MM1032 N_VPWR_M1032_d N_A_2199_74#_M1032_g N_X_M1024_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.196 AS=0.168 PD=1.47 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.2 SB=75001.2 A=0.168 P=2.54 MULT=1
MM1034 N_VPWR_M1032_d N_A_2199_74#_M1034_g N_X_M1034_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.196 AS=0.168 PD=1.47 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75001.7 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1049 N_VPWR_M1049_d N_A_2199_74#_M1049_g N_X_M1034_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3864 AS=0.168 PD=2.93 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75002.2 SB=75000.3 A=0.168 P=2.54 MULT=1
DX52_noxref VNB VPB NWDIODE A=31.9548 P=38.08
*
.include "sky130_fd_sc_ls__mux4_4.pxi.spice"
*
.ends
*
*
