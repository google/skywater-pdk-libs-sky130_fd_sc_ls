* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__dlxbp_1 D GATE VGND VNB VPB VPWR Q Q_N
X0 a_589_80# a_373_82# a_664_392# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X1 Q a_863_98# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X2 VPWR a_1347_424# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X3 a_27_413# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X4 a_815_124# a_863_98# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 VPWR a_27_413# a_586_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 Q a_863_98# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X7 a_373_82# a_231_74# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X8 VGND a_27_413# a_589_80# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X9 VPWR GATE a_231_74# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X10 a_770_508# a_863_98# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X11 a_27_413# D VGND VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X12 a_373_82# a_231_74# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X13 VPWR a_664_392# a_863_98# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X14 VGND GATE a_231_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X15 a_586_392# a_231_74# a_664_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 VPWR a_863_98# a_1347_424# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X17 VGND a_664_392# a_863_98# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X18 VGND a_863_98# a_1347_424# VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X19 a_664_392# a_373_82# a_770_508# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X20 VGND a_1347_424# Q_N VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X21 a_664_392# a_231_74# a_815_124# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
