* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__sdfsbp_2 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q Q_N
M1000 Q_N a_2067_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=3.668e+12p ps=2.764e+07u
M1001 VGND a_1069_81# a_1794_74# VNB nshort w=640000u l=150000u
+  ad=2.2419e+12p pd=2.069e+07u as=6.208e+11p ps=5.78e+06u
M1002 a_1789_424# a_1069_81# VPWR VPB phighvt w=840000u l=150000u
+  ad=7.896e+11p pd=6.92e+06u as=0p ps=0u
M1003 VPWR a_2513_258# a_2277_455# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=2.499e+11p ps=2.87e+06u
M1004 VPWR a_2067_74# a_3177_368# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.95e+11p ps=2.59e+06u
M1005 a_1789_424# a_619_368# a_2067_74# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=4.998e+11p ps=5.14e+06u
M1006 a_220_464# SCE VPWR VPB phighvt w=640000u l=150000u
+  ad=1.728e+11p pd=1.82e+06u as=0p ps=0u
M1007 a_2501_74# a_619_368# a_2067_74# VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=5.999e+11p ps=4.61e+06u
M1008 VPWR SCE a_27_74# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.888e+11p ps=1.87e+06u
M1009 a_1794_74# a_1069_81# VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND a_2067_74# a_3177_368# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1011 Q a_3177_368# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=0p ps=0u
M1012 a_1567_74# a_1069_81# a_1252_376# VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=1.197e+11p ps=1.41e+06u
M1013 VGND SET_B a_1567_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_2067_74# SET_B VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_871_74# a_619_368# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.696e+11p pd=2.9e+06u as=0p ps=0u
M1016 a_1252_376# a_1069_81# VPWR VPB phighvt w=420000u l=150000u
+  ad=1.68e+11p pd=1.64e+06u as=0p ps=0u
M1017 a_495_74# SCE a_304_464# VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=4.515e+11p ps=3.83e+06u
M1018 VGND SCD a_495_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_1069_81# a_619_368# a_304_464# VNB nshort w=420000u l=150000u
+  ad=3.675e+11p pd=2.59e+06u as=0p ps=0u
M1020 a_2579_74# a_2513_258# a_2501_74# VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1021 VGND SET_B a_2579_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 Q_N a_2067_74# VGND VNB nshort w=740000u l=150000u
+  ad=2.22e+11p pd=2.08e+06u as=0p ps=0u
M1023 Q a_3177_368# VGND VNB nshort w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1024 VGND a_1252_376# a_1274_81# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1025 VGND a_2067_74# Q_N VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VPWR CLK a_619_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.304e+11p ps=2.83e+06u
M1027 a_1274_81# a_871_74# a_1069_81# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VPWR a_3177_368# Q VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPWR SET_B a_1252_376# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VPWR SCD a_418_464# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1031 a_1069_81# a_871_74# a_304_464# VPB phighvt w=420000u l=150000u
+  ad=1.47e+11p pd=1.54e+06u as=3.927e+11p ps=3.55e+06u
M1032 a_1794_74# a_871_74# a_2067_74# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_871_74# a_619_368# VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1034 VPWR a_1252_376# a_1201_463# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1035 a_229_74# a_27_74# VGND VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1036 a_304_464# D a_229_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_2067_74# a_871_74# a_1794_74# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 a_2513_258# a_2067_74# VGND VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1039 VGND CLK a_619_368# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1040 a_1201_463# a_619_368# a_1069_81# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1041 VPWR a_2067_74# a_2513_258# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.239e+11p ps=1.43e+06u
M1042 a_418_464# a_27_74# a_304_464# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1043 VPWR a_1069_81# a_1789_424# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1044 VGND SCE a_27_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1045 VPWR a_2067_74# Q_N VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1046 a_2067_74# a_619_368# a_1789_424# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1047 a_2067_74# a_871_74# a_2277_455# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1048 a_304_464# D a_220_464# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1049 VGND a_3177_368# Q VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
