* File: sky130_fd_sc_ls__a21oi_4.spice
* Created: Fri Aug 28 12:52:22 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__a21oi_4.pex.spice"
.subckt sky130_fd_sc_ls__a21oi_4  VNB VPB A2 A1 B1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1	B1
* A1	A1
* A2	A2
* VPB	VPB
* VNB	VNB
MM1001 N_A_84_74#_M1001_d N_A2_M1001_g N_VGND_M1001_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1961 AS=0.1036 PD=2.01 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75003.2 A=0.111 P=1.78 MULT=1
MM1013 N_A_84_74#_M1013_d N_A2_M1013_g N_VGND_M1001_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75002.8 A=0.111 P=1.78 MULT=1
MM1014 N_A_84_74#_M1013_d N_A2_M1014_g N_VGND_M1014_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75002.4 A=0.111 P=1.78 MULT=1
MM1015 N_A_84_74#_M1015_d N_A2_M1015_g N_VGND_M1014_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75001.9 A=0.111 P=1.78 MULT=1
MM1009 N_A_84_74#_M1015_d N_A1_M1009_g N_Y_M1009_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.9
+ SB=75001.5 A=0.111 P=1.78 MULT=1
MM1012 N_A_84_74#_M1012_d N_A1_M1012_g N_Y_M1009_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.3
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1020 N_A_84_74#_M1012_d N_A1_M1020_g N_Y_M1020_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.8
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1021 N_A_84_74#_M1021_d N_A1_M1021_g N_Y_M1020_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75003.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1008 N_VGND_M1008_d N_B1_M1008_g N_Y_M1008_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1961 PD=1.02 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1019 N_VGND_M1008_d N_B1_M1019_g N_Y_M1019_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1961 PD=1.02 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1002 N_A_69_368#_M1002_d N_A2_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.308 AS=0.168 PD=2.79 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75005.1 A=0.168 P=2.54 MULT=1
MM1003 N_A_69_368#_M1003_d N_A2_M1003_g N_VPWR_M1002_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.6 SB=75004.7 A=0.168 P=2.54 MULT=1
MM1005 N_A_69_368#_M1003_d N_A2_M1005_g N_VPWR_M1005_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75004.2 A=0.168 P=2.54 MULT=1
MM1018 N_A_69_368#_M1018_d N_A2_M1018_g N_VPWR_M1005_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.5 SB=75003.8 A=0.168 P=2.54 MULT=1
MM1000 N_A_69_368#_M1018_d N_A1_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75002
+ SB=75003.3 A=0.168 P=2.54 MULT=1
MM1006 N_A_69_368#_M1006_d N_A1_M1006_g N_VPWR_M1000_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.4 SB=75002.9 A=0.168 P=2.54 MULT=1
MM1010 N_A_69_368#_M1006_d N_A1_M1010_g N_VPWR_M1010_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.9 SB=75002.4 A=0.168 P=2.54 MULT=1
MM1016 N_A_69_368#_M1016_d N_A1_M1016_g N_VPWR_M1010_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75003.3 SB=75002 A=0.168 P=2.54 MULT=1
MM1004 N_Y_M1004_d N_B1_M1004_g N_A_69_368#_M1016_d VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75003.8 SB=75001.5 A=0.168 P=2.54 MULT=1
MM1007 N_Y_M1004_d N_B1_M1007_g N_A_69_368#_M1007_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75004.2 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1011 N_Y_M1011_d N_B1_M1011_g N_A_69_368#_M1007_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75004.7 SB=75000.6 A=0.168 P=2.54 MULT=1
MM1017 N_Y_M1011_d N_B1_M1017_g N_A_69_368#_M1017_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.308 PD=1.42 PS=2.79 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75005.1 SB=75000.2 A=0.168 P=2.54 MULT=1
DX22_noxref VNB VPB NWDIODE A=12.3132 P=16.96
*
.include "sky130_fd_sc_ls__a21oi_4.pxi.spice"
*
.ends
*
*
