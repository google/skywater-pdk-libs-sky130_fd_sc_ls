* File: sky130_fd_sc_ls__o31ai_1.pxi.spice
* Created: Fri Aug 28 13:53:17 2020
* 
x_PM_SKY130_FD_SC_LS__O31AI_1%A1 N_A1_c_43_n N_A1_M1005_g N_A1_c_44_n
+ N_A1_M1001_g A1 PM_SKY130_FD_SC_LS__O31AI_1%A1
x_PM_SKY130_FD_SC_LS__O31AI_1%A2 N_A2_M1006_g N_A2_c_63_n N_A2_M1007_g A2 A2 A2
+ A2 N_A2_c_64_n PM_SKY130_FD_SC_LS__O31AI_1%A2
x_PM_SKY130_FD_SC_LS__O31AI_1%A3 N_A3_c_102_n N_A3_M1004_g N_A3_M1000_g A3
+ N_A3_c_101_n PM_SKY130_FD_SC_LS__O31AI_1%A3
x_PM_SKY130_FD_SC_LS__O31AI_1%B1 N_B1_M1003_g N_B1_c_134_n N_B1_M1002_g B1
+ N_B1_c_135_n PM_SKY130_FD_SC_LS__O31AI_1%B1
x_PM_SKY130_FD_SC_LS__O31AI_1%VPWR N_VPWR_M1001_s N_VPWR_M1002_d N_VPWR_c_157_n
+ N_VPWR_c_158_n N_VPWR_c_159_n N_VPWR_c_160_n VPWR N_VPWR_c_161_n
+ N_VPWR_c_156_n PM_SKY130_FD_SC_LS__O31AI_1%VPWR
x_PM_SKY130_FD_SC_LS__O31AI_1%Y N_Y_M1003_d N_Y_M1004_d N_Y_c_185_n N_Y_c_186_n
+ N_Y_c_187_n Y Y N_Y_c_189_n N_Y_c_188_n PM_SKY130_FD_SC_LS__O31AI_1%Y
x_PM_SKY130_FD_SC_LS__O31AI_1%VGND N_VGND_M1005_s N_VGND_M1006_d N_VGND_c_226_n
+ N_VGND_c_227_n VGND N_VGND_c_228_n N_VGND_c_229_n N_VGND_c_230_n
+ N_VGND_c_231_n PM_SKY130_FD_SC_LS__O31AI_1%VGND
x_PM_SKY130_FD_SC_LS__O31AI_1%A_114_74# N_A_114_74#_M1005_d N_A_114_74#_M1000_d
+ N_A_114_74#_c_266_n N_A_114_74#_c_262_n N_A_114_74#_c_263_n
+ N_A_114_74#_c_264_n PM_SKY130_FD_SC_LS__O31AI_1%A_114_74#
cc_1 VNB N_A1_c_43_n 0.0213825f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.22
cc_2 VNB N_A1_c_44_n 0.0685421f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.765
cc_3 VNB A1 0.0103026f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_A2_M1006_g 0.0235915f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_5 VNB N_A2_c_63_n 0.0343495f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=2.4
cc_6 VNB N_A2_c_64_n 0.00639141f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A3_M1000_g 0.026895f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=2.4
cc_8 VNB A3 0.0037708f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A3_c_101_n 0.0355833f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.295
cc_10 VNB N_B1_M1003_g 0.0302921f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_11 VNB N_B1_c_134_n 0.0613222f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=2.4
cc_12 VNB N_B1_c_135_n 0.00461578f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.295
cc_13 VNB N_VPWR_c_156_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_Y_c_185_n 0.0150819f $X=-0.19 $Y=-0.245 $X2=0.357 $Y2=1.385
cc_15 VNB N_Y_c_186_n 3.20099e-19 $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_16 VNB N_Y_c_187_n 0.0262708f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_Y_c_188_n 0.00868892f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_VGND_c_226_n 0.0120272f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_19 VNB N_VGND_c_227_n 0.0337878f $X=-0.19 $Y=-0.245 $X2=0.357 $Y2=1.385
cc_20 VNB N_VGND_c_228_n 0.0319663f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_229_n 0.179964f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_230_n 0.0164203f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_231_n 0.0228461f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_114_74#_c_262_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.295
cc_25 VNB N_A_114_74#_c_263_n 0.00231275f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_114_74#_c_264_n 0.002553f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VPB N_A1_c_44_n 0.0275936f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.765
cc_28 VPB N_A2_c_63_n 0.0220077f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=2.4
cc_29 VPB N_A2_c_64_n 0.00184546f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_30 VPB N_A3_c_102_n 0.0187717f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.22
cc_31 VPB A3 0.00738154f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_32 VPB N_A3_c_101_n 0.0197506f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.295
cc_33 VPB N_B1_c_134_n 0.0285488f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=2.4
cc_34 VPB N_B1_c_135_n 0.00926038f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.295
cc_35 VPB N_VPWR_c_157_n 0.0111306f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_36 VPB N_VPWR_c_158_n 0.0564169f $X=-0.19 $Y=1.66 $X2=0.357 $Y2=1.385
cc_37 VPB N_VPWR_c_159_n 0.012808f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_38 VPB N_VPWR_c_160_n 0.0485722f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_39 VPB N_VPWR_c_161_n 0.0537671f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_40 VPB N_VPWR_c_156_n 0.0678121f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_41 VPB N_Y_c_189_n 0.00696328f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_42 VPB N_Y_c_188_n 0.00117474f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_43 N_A1_c_43_n N_A2_M1006_g 0.0106343f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_44 A1 N_A2_M1006_g 5.69588e-19 $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_45 N_A1_c_44_n N_A2_c_63_n 0.0874177f $X=0.52 $Y=1.765 $X2=0 $Y2=0
cc_46 N_A1_c_44_n N_A2_c_64_n 0.0232306f $X=0.52 $Y=1.765 $X2=0 $Y2=0
cc_47 A1 N_A2_c_64_n 0.0200321f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_48 N_A1_c_44_n N_VPWR_c_158_n 0.0139619f $X=0.52 $Y=1.765 $X2=0 $Y2=0
cc_49 A1 N_VPWR_c_158_n 0.0149782f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_50 N_A1_c_44_n N_VPWR_c_161_n 0.00461464f $X=0.52 $Y=1.765 $X2=0 $Y2=0
cc_51 N_A1_c_44_n N_VPWR_c_156_n 0.009123f $X=0.52 $Y=1.765 $X2=0 $Y2=0
cc_52 N_A1_c_43_n N_VGND_c_227_n 0.0130745f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_53 N_A1_c_44_n N_VGND_c_227_n 0.00199898f $X=0.52 $Y=1.765 $X2=0 $Y2=0
cc_54 A1 N_VGND_c_227_n 0.025255f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_55 N_A1_c_43_n N_VGND_c_229_n 0.00757637f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_56 N_A1_c_43_n N_VGND_c_230_n 0.00383152f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_57 N_A1_c_43_n N_A_114_74#_c_262_n 8.89831e-19 $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_58 N_A2_c_63_n N_A3_c_102_n 0.0348431f $X=0.94 $Y=1.765 $X2=-0.19 $Y2=-0.245
cc_59 N_A2_c_64_n N_A3_c_102_n 0.0039107f $X=1.015 $Y=1.465 $X2=-0.19 $Y2=-0.245
cc_60 N_A2_c_63_n N_A3_M1000_g 5.59819e-19 $X=0.94 $Y=1.765 $X2=0 $Y2=0
cc_61 N_A2_c_63_n N_A3_c_101_n 0.0123445f $X=0.94 $Y=1.765 $X2=0 $Y2=0
cc_62 N_A2_c_64_n N_A3_c_101_n 5.84032e-19 $X=1.015 $Y=1.465 $X2=0 $Y2=0
cc_63 N_A2_c_64_n N_VPWR_c_158_n 0.0341984f $X=1.015 $Y=1.465 $X2=0 $Y2=0
cc_64 N_A2_c_63_n N_VPWR_c_161_n 0.00303293f $X=0.94 $Y=1.765 $X2=0 $Y2=0
cc_65 N_A2_c_64_n N_VPWR_c_161_n 0.0155345f $X=1.015 $Y=1.465 $X2=0 $Y2=0
cc_66 N_A2_c_63_n N_VPWR_c_156_n 0.00372936f $X=0.94 $Y=1.765 $X2=0 $Y2=0
cc_67 N_A2_c_64_n N_VPWR_c_156_n 0.0192311f $X=1.015 $Y=1.465 $X2=0 $Y2=0
cc_68 N_A2_c_64_n A_119_368# 0.00389278f $X=1.015 $Y=1.465 $X2=-0.19 $Y2=-0.245
cc_69 N_A2_c_64_n A_203_368# 0.0109027f $X=1.015 $Y=1.465 $X2=-0.19 $Y2=-0.245
cc_70 N_A2_M1006_g N_Y_c_186_n 0.00330111f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_71 N_A2_c_63_n N_Y_c_189_n 0.00214029f $X=0.94 $Y=1.765 $X2=0 $Y2=0
cc_72 N_A2_M1006_g N_Y_c_188_n 0.00477786f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_73 N_A2_c_63_n N_Y_c_188_n 0.00627607f $X=0.94 $Y=1.765 $X2=0 $Y2=0
cc_74 N_A2_c_64_n N_Y_c_188_n 0.135015f $X=1.015 $Y=1.465 $X2=0 $Y2=0
cc_75 N_A2_M1006_g N_VGND_c_227_n 5.69788e-19 $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_76 N_A2_M1006_g N_VGND_c_229_n 0.00404728f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_77 N_A2_M1006_g N_VGND_c_230_n 0.00320194f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_78 N_A2_M1006_g N_VGND_c_231_n 0.00531017f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_79 N_A2_M1006_g N_A_114_74#_c_266_n 0.0122762f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_80 N_A2_c_63_n N_A_114_74#_c_266_n 7.85764e-19 $X=0.94 $Y=1.765 $X2=0 $Y2=0
cc_81 N_A2_c_64_n N_A_114_74#_c_266_n 0.008902f $X=1.015 $Y=1.465 $X2=0 $Y2=0
cc_82 N_A2_M1006_g N_A_114_74#_c_262_n 0.010161f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_83 N_A2_M1006_g N_A_114_74#_c_263_n 0.0107236f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_84 N_A2_c_64_n N_A_114_74#_c_263_n 0.0230199f $X=1.015 $Y=1.465 $X2=0 $Y2=0
cc_85 N_A3_M1000_g N_B1_M1003_g 0.0316207f $X=1.885 $Y=0.74 $X2=0 $Y2=0
cc_86 N_A3_c_102_n N_B1_c_134_n 0.0057915f $X=1.51 $Y=1.765 $X2=0 $Y2=0
cc_87 A3 N_B1_c_134_n 0.0115059f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_88 N_A3_c_101_n N_B1_c_134_n 0.0190819f $X=1.855 $Y=1.515 $X2=0 $Y2=0
cc_89 N_A3_M1000_g N_B1_c_135_n 2.15196e-19 $X=1.885 $Y=0.74 $X2=0 $Y2=0
cc_90 A3 N_B1_c_135_n 0.0343232f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_91 N_A3_c_102_n N_VPWR_c_161_n 0.00291513f $X=1.51 $Y=1.765 $X2=0 $Y2=0
cc_92 N_A3_c_102_n N_VPWR_c_156_n 0.00363065f $X=1.51 $Y=1.765 $X2=0 $Y2=0
cc_93 N_A3_M1000_g N_Y_c_185_n 0.0125598f $X=1.885 $Y=0.74 $X2=0 $Y2=0
cc_94 A3 N_Y_c_185_n 0.0374035f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_95 N_A3_c_101_n N_Y_c_185_n 0.00884428f $X=1.855 $Y=1.515 $X2=0 $Y2=0
cc_96 N_A3_c_102_n N_Y_c_189_n 0.0281338f $X=1.51 $Y=1.765 $X2=0 $Y2=0
cc_97 A3 N_Y_c_189_n 0.0471524f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_98 N_A3_c_101_n N_Y_c_189_n 0.00443454f $X=1.855 $Y=1.515 $X2=0 $Y2=0
cc_99 N_A3_c_102_n N_Y_c_188_n 0.00943478f $X=1.51 $Y=1.765 $X2=0 $Y2=0
cc_100 N_A3_M1000_g N_Y_c_188_n 0.00612746f $X=1.885 $Y=0.74 $X2=0 $Y2=0
cc_101 A3 N_Y_c_188_n 0.033267f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_102 N_A3_c_101_n N_Y_c_188_n 0.00961308f $X=1.855 $Y=1.515 $X2=0 $Y2=0
cc_103 N_A3_M1000_g N_VGND_c_228_n 0.00320194f $X=1.885 $Y=0.74 $X2=0 $Y2=0
cc_104 N_A3_M1000_g N_VGND_c_229_n 0.00404912f $X=1.885 $Y=0.74 $X2=0 $Y2=0
cc_105 N_A3_M1000_g N_VGND_c_231_n 0.00703231f $X=1.885 $Y=0.74 $X2=0 $Y2=0
cc_106 N_A3_M1000_g N_A_114_74#_c_266_n 0.0108636f $X=1.885 $Y=0.74 $X2=0 $Y2=0
cc_107 N_A3_M1000_g N_A_114_74#_c_264_n 0.0106282f $X=1.885 $Y=0.74 $X2=0 $Y2=0
cc_108 N_B1_c_134_n N_VPWR_c_160_n 0.0202043f $X=2.35 $Y=1.765 $X2=0 $Y2=0
cc_109 N_B1_c_135_n N_VPWR_c_160_n 0.0246455f $X=2.61 $Y=1.465 $X2=0 $Y2=0
cc_110 N_B1_c_134_n N_VPWR_c_161_n 0.00413917f $X=2.35 $Y=1.765 $X2=0 $Y2=0
cc_111 N_B1_c_134_n N_VPWR_c_156_n 0.00820326f $X=2.35 $Y=1.765 $X2=0 $Y2=0
cc_112 N_B1_M1003_g N_Y_c_185_n 0.0174305f $X=2.335 $Y=0.74 $X2=0 $Y2=0
cc_113 N_B1_c_134_n N_Y_c_185_n 0.00401927f $X=2.35 $Y=1.765 $X2=0 $Y2=0
cc_114 N_B1_c_135_n N_Y_c_185_n 0.0277433f $X=2.61 $Y=1.465 $X2=0 $Y2=0
cc_115 N_B1_M1003_g N_Y_c_187_n 0.00164953f $X=2.335 $Y=0.74 $X2=0 $Y2=0
cc_116 N_B1_c_134_n N_Y_c_189_n 2.57779e-19 $X=2.35 $Y=1.765 $X2=0 $Y2=0
cc_117 N_B1_M1003_g N_VGND_c_228_n 0.00456932f $X=2.335 $Y=0.74 $X2=0 $Y2=0
cc_118 N_B1_M1003_g N_VGND_c_229_n 0.00894956f $X=2.335 $Y=0.74 $X2=0 $Y2=0
cc_119 N_B1_M1003_g N_A_114_74#_c_264_n 0.004688f $X=2.335 $Y=0.74 $X2=0 $Y2=0
cc_120 N_VPWR_c_160_n N_Y_c_189_n 0.0377637f $X=2.575 $Y=2.115 $X2=0 $Y2=0
cc_121 N_VPWR_c_161_n N_Y_c_189_n 0.0387288f $X=2.41 $Y=3.33 $X2=0 $Y2=0
cc_122 N_VPWR_c_156_n N_Y_c_189_n 0.031704f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_123 A_203_368# N_Y_c_189_n 0.00984915f $X=1.015 $Y=1.84 $X2=0 $Y2=0
cc_124 A_203_368# N_Y_c_188_n 9.72352e-19 $X=1.015 $Y=1.84 $X2=0.892 $Y2=1.665
cc_125 N_Y_c_185_n N_VGND_M1006_d 0.00337116f $X=2.435 $Y=1.045 $X2=0 $Y2=0
cc_126 N_Y_c_186_n N_VGND_M1006_d 0.00548721f $X=1.52 $Y=1.045 $X2=0 $Y2=0
cc_127 N_Y_c_187_n N_VGND_c_228_n 0.0146357f $X=2.6 $Y=0.515 $X2=0 $Y2=0
cc_128 N_Y_c_187_n N_VGND_c_229_n 0.0121141f $X=2.6 $Y=0.515 $X2=0 $Y2=0
cc_129 N_Y_c_185_n N_A_114_74#_M1000_d 0.00197722f $X=2.435 $Y=1.045 $X2=0 $Y2=0
cc_130 N_Y_c_185_n N_A_114_74#_c_266_n 0.0253598f $X=2.435 $Y=1.045 $X2=0 $Y2=0
cc_131 N_Y_c_186_n N_A_114_74#_c_266_n 0.013831f $X=1.52 $Y=1.045 $X2=0 $Y2=0
cc_132 N_Y_c_186_n N_A_114_74#_c_263_n 0.0062517f $X=1.52 $Y=1.045 $X2=0 $Y2=0
cc_133 N_Y_c_185_n N_A_114_74#_c_264_n 0.016668f $X=2.435 $Y=1.045 $X2=0 $Y2=0
cc_134 N_Y_c_187_n N_A_114_74#_c_264_n 0.0173003f $X=2.6 $Y=0.515 $X2=0 $Y2=0
cc_135 N_VGND_M1006_d N_A_114_74#_c_266_n 0.023923f $X=1 $Y=0.37 $X2=0 $Y2=0
cc_136 N_VGND_c_228_n N_A_114_74#_c_266_n 0.00266409f $X=2.64 $Y=0 $X2=0 $Y2=0
cc_137 N_VGND_c_229_n N_A_114_74#_c_266_n 0.0123863f $X=2.64 $Y=0 $X2=0 $Y2=0
cc_138 N_VGND_c_230_n N_A_114_74#_c_266_n 0.00266409f $X=1.055 $Y=0.182 $X2=0
+ $Y2=0
cc_139 N_VGND_c_231_n N_A_114_74#_c_266_n 0.0525207f $X=1.755 $Y=0.182 $X2=0
+ $Y2=0
cc_140 N_VGND_c_227_n N_A_114_74#_c_262_n 0.0243832f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_141 N_VGND_c_229_n N_A_114_74#_c_262_n 0.00904371f $X=2.64 $Y=0 $X2=0 $Y2=0
cc_142 N_VGND_c_230_n N_A_114_74#_c_262_n 0.0109942f $X=1.055 $Y=0.182 $X2=0
+ $Y2=0
cc_143 N_VGND_c_231_n N_A_114_74#_c_262_n 0.00426994f $X=1.755 $Y=0.182 $X2=0
+ $Y2=0
cc_144 N_VGND_c_228_n N_A_114_74#_c_264_n 0.0141059f $X=2.64 $Y=0 $X2=0 $Y2=0
cc_145 N_VGND_c_229_n N_A_114_74#_c_264_n 0.0118064f $X=2.64 $Y=0 $X2=0 $Y2=0
cc_146 N_VGND_c_231_n N_A_114_74#_c_264_n 0.00441839f $X=1.755 $Y=0.182 $X2=0
+ $Y2=0
