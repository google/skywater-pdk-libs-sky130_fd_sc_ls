* File: sky130_fd_sc_ls__maj3_2.spice
* Created: Wed Sep  2 11:09:55 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__maj3_2.pex.spice"
.subckt sky130_fd_sc_ls__maj3_2  VNB VPB B C A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* C	C
* B	B
* VPB	VPB
* VNB	VNB
MM1010 N_VGND_M1010_d N_A_87_264#_M1010_g N_X_M1010_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75004 A=0.111 P=1.78 MULT=1
MM1013 N_VGND_M1013_d N_A_87_264#_M1013_g N_X_M1010_s VNB NSHORT L=0.15 W=0.74
+ AD=0.33115 AS=0.1036 PD=1.635 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75003.5 A=0.111 P=1.78 MULT=1
MM1008 A_413_74# N_A_M1008_g N_VGND_M1013_d VNB NSHORT L=0.15 W=0.74 AD=0.0888
+ AS=0.33115 PD=0.98 PS=1.635 NRD=10.536 NRS=10.536 M=1 R=4.93333 SA=75001.7
+ SB=75002.5 A=0.111 P=1.78 MULT=1
MM1009 N_A_87_264#_M1009_d N_B_M1009_g A_413_74# VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.0888 PD=1.02 PS=0.98 NRD=0 NRS=10.536 M=1 R=4.93333 SA=75002.1
+ SB=75002.1 A=0.111 P=1.78 MULT=1
MM1001 A_577_74# N_B_M1001_g N_A_87_264#_M1009_d VNB NSHORT L=0.15 W=0.74
+ AD=0.1221 AS=0.1036 PD=1.07 PS=1.02 NRD=17.832 NRS=0 M=1 R=4.93333 SA=75002.5
+ SB=75001.7 A=0.111 P=1.78 MULT=1
MM1004 N_VGND_M1004_d N_C_M1004_g A_577_74# VNB NSHORT L=0.15 W=0.74 AD=0.1665
+ AS=0.1221 PD=1.19 PS=1.07 NRD=13.776 NRS=17.832 M=1 R=4.93333 SA=75003
+ SB=75001.2 A=0.111 P=1.78 MULT=1
MM1011 A_793_74# N_A_M1011_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.74 AD=0.0888
+ AS=0.1665 PD=0.98 PS=1.19 NRD=10.536 NRS=13.776 M=1 R=4.93333 SA=75003.6
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1012 N_A_87_264#_M1012_d N_C_M1012_g A_793_74# VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.0888 PD=2.05 PS=0.98 NRD=0 NRS=10.536 M=1 R=4.93333 SA=75004
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1002 N_X_M1002_d N_A_87_264#_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75003.4 A=0.168 P=2.54 MULT=1
MM1003 N_X_M1002_d N_A_87_264#_M1003_g N_VPWR_M1003_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.426023 PD=1.42 PS=1.9917 NRD=1.7533 NRS=2.6201 M=1 R=7.46667
+ SA=75000.7 SB=75003 A=0.168 P=2.54 MULT=1
MM1006 A_393_368# N_A_M1006_g N_VPWR_M1003_s VPB PHIGHVT L=0.15 W=1 AD=0.186687
+ AS=0.380377 PD=1.46 PS=1.7783 NRD=25.9252 NRS=2.9353 M=1 R=6.66667 SA=75001.6
+ SB=75002.4 A=0.15 P=2.3 MULT=1
MM1014 N_A_87_264#_M1014_d N_B_M1014_g A_393_368# VPB PHIGHVT L=0.15 W=1 AD=0.15
+ AS=0.186687 PD=1.3 PS=1.46 NRD=1.9503 NRS=25.9252 M=1 R=6.66667 SA=75001.9
+ SB=75002 A=0.15 P=2.3 MULT=1
MM1015 A_584_347# N_B_M1015_g N_A_87_264#_M1014_d VPB PHIGHVT L=0.15 W=1
+ AD=0.155 AS=0.15 PD=1.31 PS=1.3 NRD=19.6803 NRS=1.9503 M=1 R=6.66667
+ SA=75002.3 SB=75001.6 A=0.15 P=2.3 MULT=1
MM1000 N_VPWR_M1000_d N_C_M1000_g A_584_347# VPB PHIGHVT L=0.15 W=1 AD=0.2184
+ AS=0.155 PD=1.525 PS=1.31 NRD=26.1025 NRS=19.6803 M=1 R=6.66667 SA=75002.8
+ SB=75001.1 A=0.15 P=2.3 MULT=1
MM1007 A_790_368# N_A_M1007_g N_VPWR_M1000_d VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.2184 PD=1.27 PS=1.525 NRD=15.7403 NRS=1.9503 M=1 R=6.66667 SA=75003.2
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1005 N_A_87_264#_M1005_d N_C_M1005_g A_790_368# VPB PHIGHVT L=0.15 W=1
+ AD=0.295 AS=0.135 PD=2.59 PS=1.27 NRD=1.9503 NRS=15.7403 M=1 R=6.66667
+ SA=75003.6 SB=75000.2 A=0.15 P=2.3 MULT=1
DX16_noxref VNB VPB NWDIODE A=9.83955 P=14.29
*
.include "sky130_fd_sc_ls__maj3_2.pxi.spice"
*
.ends
*
*
