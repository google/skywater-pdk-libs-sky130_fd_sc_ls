* File: sky130_fd_sc_ls__xnor3_4.pex.spice
* Created: Wed Sep  2 11:30:46 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__XNOR3_4%A_75_227# 1 2 3 4 14 15 17 20 22 23 25 26 27
+ 30 34 35 36 38 39 43 48 49 52 57
c134 34 0 1.89638e-19 $X=1.26 $Y=0.53
r135 52 54 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=3.515 $Y=2.795
+ $X2=3.515 $Y2=2.99
r136 48 49 9.77977 $w=1.88e-07 $l=1.65e-07 $layer=LI1_cond $X=3.365 $Y=0.35
+ $X2=3.2 $Y2=0.35
r137 43 58 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.54 $Y=1.3
+ $X2=0.54 $Y2=1.465
r138 43 57 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.54 $Y=1.3
+ $X2=0.54 $Y2=1.135
r139 42 44 8.79328 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=0.58 $Y=1.3
+ $X2=0.58 $Y2=1.465
r140 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.54
+ $Y=1.3 $X2=0.54 $Y2=1.3
r141 39 42 8.29759 $w=2.48e-07 $l=1.8e-07 $layer=LI1_cond $X=0.58 $Y=1.12
+ $X2=0.58 $Y2=1.3
r142 38 49 115.802 $w=1.68e-07 $l=1.775e-06 $layer=LI1_cond $X=1.425 $Y=0.34
+ $X2=3.2 $Y2=0.34
r143 35 54 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.35 $Y=2.99
+ $X2=3.515 $Y2=2.99
r144 35 36 127.545 $w=1.68e-07 $l=1.955e-06 $layer=LI1_cond $X=3.35 $Y=2.99
+ $X2=1.395 $Y2=2.99
r145 32 34 23.2793 $w=2.48e-07 $l=5.05e-07 $layer=LI1_cond $X=1.3 $Y=1.035
+ $X2=1.3 $Y2=0.53
r146 31 38 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.3 $Y=0.425
+ $X2=1.425 $Y2=0.34
r147 31 34 4.84026 $w=2.48e-07 $l=1.05e-07 $layer=LI1_cond $X=1.3 $Y=0.425
+ $X2=1.3 $Y2=0.53
r148 28 36 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.23 $Y=2.905
+ $X2=1.395 $Y2=2.99
r149 28 30 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=1.23 $Y=2.905
+ $X2=1.23 $Y2=2.72
r150 27 46 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.23 $Y=2.12 $X2=1.23
+ $Y2=2.035
r151 27 30 20.9535 $w=3.28e-07 $l=6e-07 $layer=LI1_cond $X=1.23 $Y=2.12 $X2=1.23
+ $Y2=2.72
r152 25 46 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.065 $Y=2.035
+ $X2=1.23 $Y2=2.035
r153 25 26 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=1.065 $Y=2.035
+ $X2=0.705 $Y2=2.035
r154 24 39 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.705 $Y=1.12
+ $X2=0.58 $Y2=1.12
r155 23 32 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.175 $Y=1.12
+ $X2=1.3 $Y2=1.035
r156 23 24 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=1.175 $Y=1.12
+ $X2=0.705 $Y2=1.12
r157 22 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.62 $Y=1.95
+ $X2=0.705 $Y2=2.035
r158 22 44 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=0.62 $Y=1.95
+ $X2=0.62 $Y2=1.465
r159 20 57 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=0.545 $Y=0.705
+ $X2=0.545 $Y2=1.135
r160 15 17 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.505 $Y=1.79
+ $X2=0.505 $Y2=2.365
r161 14 15 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.505 $Y=1.7
+ $X2=0.505 $Y2=1.79
r162 14 58 91.3468 $w=1.8e-07 $l=2.35e-07 $layer=POLY_cond $X=0.505 $Y=1.7
+ $X2=0.505 $Y2=1.465
r163 4 52 600 $w=1.7e-07 $l=1.04089e-06 $layer=licon1_PDIFF $count=1 $X=3.28
+ $Y=1.865 $X2=3.515 $Y2=2.795
r164 3 46 300 $w=1.7e-07 $l=2.33238e-07 $layer=licon1_PDIFF $count=2 $X=1.08
+ $Y=1.865 $X2=1.23 $Y2=2.035
r165 3 30 600 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=1.08
+ $Y=1.865 $X2=1.23 $Y2=2.72
r166 2 48 182 $w=1.7e-07 $l=3.37528e-07 $layer=licon1_NDIFF $count=1 $X=3.145
+ $Y=0.605 $X2=3.365 $Y2=0.36
r167 1 34 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.12
+ $Y=0.385 $X2=1.26 $Y2=0.53
.ends

.subckt PM_SKY130_FD_SC_LS__XNOR3_4%A 1 3 6 8 12
c44 6 0 1.6832e-19 $X=1.045 $Y=0.705
c45 1 0 9.56919e-20 $X=1.005 $Y=1.79
r46 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.08
+ $Y=1.54 $X2=1.08 $Y2=1.54
r47 8 12 3.60138 $w=3.98e-07 $l=1.25e-07 $layer=LI1_cond $X=1.115 $Y=1.665
+ $X2=1.115 $Y2=1.54
r48 4 11 38.5562 $w=2.99e-07 $l=1.81659e-07 $layer=POLY_cond $X=1.045 $Y=1.375
+ $X2=1.08 $Y2=1.54
r49 4 6 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=1.045 $Y=1.375
+ $X2=1.045 $Y2=0.705
r50 1 11 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=1.005 $Y=1.79
+ $X2=1.08 $Y2=1.54
r51 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.005 $Y=1.79
+ $X2=1.005 $Y2=2.365
.ends

.subckt PM_SKY130_FD_SC_LS__XNOR3_4%A_386_23# 1 2 10 11 12 13 14 15 17 21 22 24
+ 29 35 37 38 40 42 44 46
c128 37 0 4.27592e-20 $X=3.685 $Y=1.95
c129 22 0 1.9098e-19 $X=3.205 $Y=1.79
c130 14 0 8.8275e-20 $X=2.245 $Y=1.7
c131 11 0 1.46697e-19 $X=2.995 $Y=0.19
c132 10 0 7.08805e-20 $X=2.005 $Y=0.815
r133 42 44 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=3.77 $Y=2.075
+ $X2=4.105 $Y2=2.075
r134 38 40 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=3.77 $Y=1.04
+ $X2=3.925 $Y2=1.04
r135 37 42 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.685 $Y=1.95
+ $X2=3.77 $Y2=2.075
r136 36 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.685 $Y=1.705
+ $X2=3.685 $Y2=1.54
r137 36 37 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=3.685 $Y=1.705
+ $X2=3.685 $Y2=1.95
r138 35 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.685 $Y=1.375
+ $X2=3.685 $Y2=1.54
r139 34 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.685 $Y=1.125
+ $X2=3.77 $Y2=1.04
r140 34 35 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.685 $Y=1.125
+ $X2=3.685 $Y2=1.375
r141 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.16
+ $Y=1.54 $X2=3.16 $Y2=1.54
r142 29 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.6 $Y=1.54
+ $X2=3.685 $Y2=1.54
r143 29 31 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=3.6 $Y=1.54
+ $X2=3.16 $Y2=1.54
r144 22 32 52.2586 $w=2.99e-07 $l=2.7157e-07 $layer=POLY_cond $X=3.205 $Y=1.79
+ $X2=3.16 $Y2=1.54
r145 22 24 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=3.205 $Y=1.79
+ $X2=3.205 $Y2=2.285
r146 19 32 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=3.07 $Y=1.375
+ $X2=3.16 $Y2=1.54
r147 19 21 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=3.07 $Y=1.375
+ $X2=3.07 $Y2=0.925
r148 18 21 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.07 $Y=0.265
+ $X2=3.07 $Y2=0.925
r149 15 17 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.245 $Y=1.79
+ $X2=2.245 $Y2=2.185
r150 14 15 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.245 $Y=1.7
+ $X2=2.245 $Y2=1.79
r151 13 25 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=2.245 $Y=1.395
+ $X2=2.005 $Y2=1.395
r152 13 14 89.4032 $w=1.8e-07 $l=2.3e-07 $layer=POLY_cond $X=2.245 $Y=1.47
+ $X2=2.245 $Y2=1.7
r153 11 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.995 $Y=0.19
+ $X2=3.07 $Y2=0.265
r154 11 12 469.181 $w=1.5e-07 $l=9.15e-07 $layer=POLY_cond $X=2.995 $Y=0.19
+ $X2=2.08 $Y2=0.19
r155 8 25 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.005 $Y=1.32
+ $X2=2.005 $Y2=1.395
r156 8 10 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=2.005 $Y=1.32
+ $X2=2.005 $Y2=0.815
r157 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.005 $Y=0.265
+ $X2=2.08 $Y2=0.19
r158 7 10 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.005 $Y=0.265
+ $X2=2.005 $Y2=0.815
r159 2 44 600 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=3.96
+ $Y=1.84 $X2=4.105 $Y2=2.115
r160 1 40 182 $w=1.7e-07 $l=6.63551e-07 $layer=licon1_NDIFF $count=1 $X=3.78
+ $Y=0.445 $X2=3.925 $Y2=1.04
.ends

.subckt PM_SKY130_FD_SC_LS__XNOR3_4%B 3 5 6 7 10 11 12 15 17 18 22 23 26 29 31
+ 33 37 39 40 45 46
c153 46 0 4.27592e-20 $X=4.14 $Y=1.557
c154 45 0 1.9098e-19 $X=4.105 $Y=1.515
c155 26 0 2.21365e-20 $X=3.81 $Y=3.075
c156 22 0 8.1711e-21 $X=2.695 $Y=2.185
c157 7 0 1.19763e-19 $X=1.545 $Y=1.79
c158 3 0 1.70469e-19 $X=1.53 $Y=0.705
r159 46 47 30.7315 $w=2.98e-07 $l=1.9e-07 $layer=POLY_cond $X=4.14 $Y=1.557
+ $X2=4.33 $Y2=1.557
r160 44 46 5.66107 $w=2.98e-07 $l=3.5e-08 $layer=POLY_cond $X=4.105 $Y=1.557
+ $X2=4.14 $Y2=1.557
r161 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.105
+ $Y=1.515 $X2=4.105 $Y2=1.515
r162 40 45 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=4.105 $Y=1.665
+ $X2=4.105 $Y2=1.515
r163 35 37 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.62 $Y=1.715
+ $X2=2.695 $Y2=1.715
r164 31 47 18.8112 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=4.33 $Y=1.765
+ $X2=4.33 $Y2=1.557
r165 31 33 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.33 $Y=1.765
+ $X2=4.33 $Y2=2.4
r166 27 46 18.8112 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.14 $Y=1.35
+ $X2=4.14 $Y2=1.557
r167 27 29 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=4.14 $Y=1.35
+ $X2=4.14 $Y2=0.815
r168 25 44 47.7148 $w=2.98e-07 $l=2.95e-07 $layer=POLY_cond $X=3.81 $Y=1.557
+ $X2=4.105 $Y2=1.557
r169 25 26 715.309 $w=1.5e-07 $l=1.395e-06 $layer=POLY_cond $X=3.81 $Y=1.68
+ $X2=3.81 $Y2=3.075
r170 24 39 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.785 $Y=3.15
+ $X2=2.695 $Y2=3.15
r171 23 26 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.735 $Y=3.15
+ $X2=3.81 $Y2=3.075
r172 23 24 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=3.735 $Y=3.15
+ $X2=2.785 $Y2=3.15
r173 20 22 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.695 $Y=2.58
+ $X2=2.695 $Y2=2.185
r174 19 37 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.695 $Y=1.79
+ $X2=2.695 $Y2=1.715
r175 19 22 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.695 $Y=1.79
+ $X2=2.695 $Y2=2.185
r176 18 39 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=2.695 $Y=3.075
+ $X2=2.695 $Y2=3.15
r177 17 20 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.695 $Y=2.67
+ $X2=2.695 $Y2=2.58
r178 17 18 157.427 $w=1.8e-07 $l=4.05e-07 $layer=POLY_cond $X=2.695 $Y=2.67
+ $X2=2.695 $Y2=3.075
r179 13 35 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.62 $Y=1.64
+ $X2=2.62 $Y2=1.715
r180 13 15 366.628 $w=1.5e-07 $l=7.15e-07 $layer=POLY_cond $X=2.62 $Y=1.64
+ $X2=2.62 $Y2=0.925
r181 11 39 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.605 $Y=3.15
+ $X2=2.695 $Y2=3.15
r182 11 12 497.383 $w=1.5e-07 $l=9.7e-07 $layer=POLY_cond $X=2.605 $Y=3.15
+ $X2=1.635 $Y2=3.15
r183 8 10 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.545 $Y=2.78
+ $X2=1.545 $Y2=2.285
r184 7 34 58.3064 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=1.545 $Y=1.79
+ $X2=1.545 $Y2=1.64
r185 7 10 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.545 $Y=1.79
+ $X2=1.545 $Y2=2.285
r186 6 12 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=1.545 $Y=3.075
+ $X2=1.635 $Y2=3.15
r187 5 8 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.545 $Y=2.87 $X2=1.545
+ $Y2=2.78
r188 5 6 79.6855 $w=1.8e-07 $l=2.05e-07 $layer=POLY_cond $X=1.545 $Y=2.87
+ $X2=1.545 $Y2=3.075
r189 3 34 479.436 $w=1.5e-07 $l=9.35e-07 $layer=POLY_cond $X=1.53 $Y=0.705
+ $X2=1.53 $Y2=1.64
.ends

.subckt PM_SKY130_FD_SC_LS__XNOR3_4%A_1024_300# 1 2 9 11 13 14 17 19 24 26 29 33
r82 30 33 6.33218 $w=5.08e-07 $l=2.7e-07 $layer=LI1_cond $X=6.525 $Y=2.245
+ $X2=6.795 $Y2=2.245
r83 26 28 4.25191 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=6.555 $Y=1.085
+ $X2=6.555 $Y2=1.17
r84 21 24 9.07524 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=5.285 $Y=1.665
+ $X2=5.45 $Y2=1.665
r85 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.285
+ $Y=1.665 $X2=5.285 $Y2=1.665
r86 19 30 7.28118 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=6.525 $Y=1.99
+ $X2=6.525 $Y2=2.245
r87 18 29 4.60183 $w=1.95e-07 $l=9.66954e-08 $layer=LI1_cond $X=6.525 $Y=1.72
+ $X2=6.5 $Y2=1.635
r88 18 19 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=6.525 $Y=1.72
+ $X2=6.525 $Y2=1.99
r89 17 29 4.60183 $w=1.95e-07 $l=8.5e-08 $layer=LI1_cond $X=6.5 $Y=1.55 $X2=6.5
+ $Y2=1.635
r90 17 28 19.9058 $w=2.18e-07 $l=3.8e-07 $layer=LI1_cond $X=6.5 $Y=1.55 $X2=6.5
+ $Y2=1.17
r91 14 29 1.84097 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=6.39 $Y=1.635 $X2=6.5
+ $Y2=1.635
r92 14 24 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=6.39 $Y=1.635
+ $X2=5.45 $Y2=1.635
r93 11 22 52.2586 $w=2.99e-07 $l=2.76134e-07 $layer=POLY_cond $X=5.34 $Y=1.915
+ $X2=5.285 $Y2=1.665
r94 11 13 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=5.34 $Y=1.915
+ $X2=5.34 $Y2=2.41
r95 7 22 38.5562 $w=2.99e-07 $l=1.98997e-07 $layer=POLY_cond $X=5.21 $Y=1.5
+ $X2=5.285 $Y2=1.665
r96 7 9 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=5.21 $Y=1.5 $X2=5.21
+ $Y2=0.69
r97 2 33 600 $w=1.7e-07 $l=4.61844e-07 $layer=licon1_PDIFF $count=1 $X=6.65
+ $Y=1.84 $X2=6.795 $Y2=2.235
r98 1 26 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=6.41
+ $Y=0.81 $X2=6.555 $Y2=1.085
.ends

.subckt PM_SKY130_FD_SC_LS__XNOR3_4%C 3 6 7 9 10 11 12 14 15 17 21 26
c75 12 0 2.47917e-19 $X=6.77 $Y=1.35
r76 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.945
+ $Y=1.515 $X2=6.945 $Y2=1.515
r77 23 25 11.8525 $w=3.66e-07 $l=9e-08 $layer=POLY_cond $X=6.902 $Y=1.425
+ $X2=6.902 $Y2=1.515
r78 21 26 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=6.945 $Y=1.665
+ $X2=6.945 $Y2=1.515
r79 15 25 50.1894 $w=3.66e-07 $l=3.03315e-07 $layer=POLY_cond $X=7.02 $Y=1.765
+ $X2=6.902 $Y2=1.515
r80 15 17 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=7.02 $Y=1.765
+ $X2=7.02 $Y2=2.16
r81 12 23 27.143 $w=3.66e-07 $l=1.653e-07 $layer=POLY_cond $X=6.77 $Y=1.35
+ $X2=6.902 $Y2=1.425
r82 12 14 106.04 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=6.77 $Y=1.35 $X2=6.77
+ $Y2=1.02
r83 10 23 23.7042 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.695 $Y=1.425
+ $X2=6.902 $Y2=1.425
r84 10 11 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=6.695 $Y=1.425
+ $X2=6.05 $Y2=1.425
r85 7 9 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=5.96 $Y=1.915 $X2=5.96
+ $Y2=2.41
r86 6 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.96 $Y=1.825 $X2=5.96
+ $Y2=1.915
r87 5 11 46.1489 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=5.96 $Y=1.425 $X2=6.05
+ $Y2=1.425
r88 5 18 99.9894 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=5.96 $Y=1.425
+ $X2=5.765 $Y2=1.425
r89 5 6 126.331 $w=1.8e-07 $l=3.25e-07 $layer=POLY_cond $X=5.96 $Y=1.5 $X2=5.96
+ $Y2=1.825
r90 1 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.765 $Y=1.35
+ $X2=5.765 $Y2=1.425
r91 1 3 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.765 $Y=1.35
+ $X2=5.765 $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_LS__XNOR3_4%A_1057_74# 1 2 7 9 10 12 13 15 16 18 19 21
+ 22 24 25 27 28 30 33 35 36 37 40 41 42 44 45 46 48 50 52 55 59 65 68 70 80
c159 70 0 1.96868e-19 $X=8.13 $Y=1.505
c160 68 0 1.17951e-19 $X=7.485 $Y=1.505
r161 80 81 1.93834 $w=3.73e-07 $l=1.5e-08 $layer=POLY_cond $X=9.57 $Y=1.552
+ $X2=9.585 $Y2=1.552
r162 79 80 53.6273 $w=3.73e-07 $l=4.15e-07 $layer=POLY_cond $X=9.155 $Y=1.552
+ $X2=9.57 $Y2=1.552
r163 78 79 4.52279 $w=3.73e-07 $l=3.5e-08 $layer=POLY_cond $X=9.12 $Y=1.552
+ $X2=9.155 $Y2=1.552
r164 77 78 51.0429 $w=3.73e-07 $l=3.95e-07 $layer=POLY_cond $X=8.725 $Y=1.552
+ $X2=9.12 $Y2=1.552
r165 76 77 7.10724 $w=3.73e-07 $l=5.5e-08 $layer=POLY_cond $X=8.67 $Y=1.552
+ $X2=8.725 $Y2=1.552
r166 75 76 48.4584 $w=3.73e-07 $l=3.75e-07 $layer=POLY_cond $X=8.295 $Y=1.552
+ $X2=8.67 $Y2=1.552
r167 74 75 9.69169 $w=3.73e-07 $l=7.5e-08 $layer=POLY_cond $X=8.22 $Y=1.552
+ $X2=8.295 $Y2=1.552
r168 69 70 112.786 $w=3.3e-07 $l=6.45e-07 $layer=POLY_cond $X=7.485 $Y=1.505
+ $X2=8.13 $Y2=1.505
r169 68 69 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=7.485
+ $Y=1.505 $X2=7.485 $Y2=1.505
r170 63 65 11.939 $w=1.68e-07 $l=1.83e-07 $layer=LI1_cond $X=7.222 $Y=2.035
+ $X2=7.405 $Y2=2.035
r171 59 61 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=5.65 $Y=2.895
+ $X2=5.65 $Y2=2.99
r172 56 74 7.10724 $w=3.73e-07 $l=5.5e-08 $layer=POLY_cond $X=8.165 $Y=1.552
+ $X2=8.22 $Y2=1.552
r173 56 70 5.28177 $w=3.73e-07 $l=6.20806e-08 $layer=POLY_cond $X=8.165 $Y=1.552
+ $X2=8.13 $Y2=1.505
r174 55 56 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=8.165
+ $Y=1.505 $X2=8.165 $Y2=1.505
r175 53 68 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.49 $Y=1.505
+ $X2=7.405 $Y2=1.505
r176 53 55 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=7.49 $Y=1.505
+ $X2=8.165 $Y2=1.505
r177 52 65 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.405 $Y=1.95
+ $X2=7.405 $Y2=2.035
r178 51 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.405 $Y=1.67
+ $X2=7.405 $Y2=1.505
r179 51 52 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=7.405 $Y=1.67
+ $X2=7.405 $Y2=1.95
r180 50 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.405 $Y=1.34
+ $X2=7.405 $Y2=1.505
r181 49 50 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=7.405 $Y=1.18
+ $X2=7.405 $Y2=1.34
r182 47 63 0.22998 $w=1.85e-07 $l=8.5e-08 $layer=LI1_cond $X=7.222 $Y=2.12
+ $X2=7.222 $Y2=2.035
r183 47 48 47.0614 $w=1.83e-07 $l=7.85e-07 $layer=LI1_cond $X=7.222 $Y=2.12
+ $X2=7.222 $Y2=2.905
r184 45 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.32 $Y=1.095
+ $X2=7.405 $Y2=1.18
r185 45 46 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=7.32 $Y=1.095
+ $X2=7.06 $Y2=1.095
r186 44 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.975 $Y=1.01
+ $X2=7.06 $Y2=1.095
r187 43 44 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=6.975 $Y=0.83
+ $X2=6.975 $Y2=1.01
r188 41 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.89 $Y=0.745
+ $X2=6.975 $Y2=0.83
r189 41 42 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=6.89 $Y=0.745
+ $X2=6.5 $Y2=0.745
r190 40 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.415 $Y=0.66
+ $X2=6.5 $Y2=0.745
r191 39 40 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=6.415 $Y=0.425
+ $X2=6.415 $Y2=0.66
r192 38 61 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.815 $Y=2.99
+ $X2=5.65 $Y2=2.99
r193 37 48 6.83233 $w=1.7e-07 $l=1.27609e-07 $layer=LI1_cond $X=7.13 $Y=2.99
+ $X2=7.222 $Y2=2.905
r194 37 38 85.7914 $w=1.68e-07 $l=1.315e-06 $layer=LI1_cond $X=7.13 $Y=2.99
+ $X2=5.815 $Y2=2.99
r195 35 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.33 $Y=0.34
+ $X2=6.415 $Y2=0.425
r196 35 36 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.33 $Y=0.34
+ $X2=5.66 $Y2=0.34
r197 31 36 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.495 $Y=0.425
+ $X2=5.66 $Y2=0.34
r198 31 33 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=5.495 $Y=0.425
+ $X2=5.495 $Y2=0.515
r199 28 81 24.162 $w=1.5e-07 $l=2.12e-07 $layer=POLY_cond $X=9.585 $Y=1.34
+ $X2=9.585 $Y2=1.552
r200 28 30 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=9.585 $Y=1.34
+ $X2=9.585 $Y2=0.86
r201 25 80 24.162 $w=1.5e-07 $l=2.13e-07 $layer=POLY_cond $X=9.57 $Y=1.765
+ $X2=9.57 $Y2=1.552
r202 25 27 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=9.57 $Y=1.765
+ $X2=9.57 $Y2=2.4
r203 22 79 24.162 $w=1.5e-07 $l=2.12e-07 $layer=POLY_cond $X=9.155 $Y=1.34
+ $X2=9.155 $Y2=1.552
r204 22 24 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=9.155 $Y=1.34
+ $X2=9.155 $Y2=0.86
r205 19 78 24.162 $w=1.5e-07 $l=2.13e-07 $layer=POLY_cond $X=9.12 $Y=1.765
+ $X2=9.12 $Y2=1.552
r206 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=9.12 $Y=1.765
+ $X2=9.12 $Y2=2.4
r207 16 77 24.162 $w=1.5e-07 $l=2.12e-07 $layer=POLY_cond $X=8.725 $Y=1.34
+ $X2=8.725 $Y2=1.552
r208 16 18 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=8.725 $Y=1.34
+ $X2=8.725 $Y2=0.86
r209 13 76 24.162 $w=1.5e-07 $l=2.13e-07 $layer=POLY_cond $X=8.67 $Y=1.765
+ $X2=8.67 $Y2=1.552
r210 13 15 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.67 $Y=1.765
+ $X2=8.67 $Y2=2.4
r211 10 75 24.162 $w=1.5e-07 $l=2.12e-07 $layer=POLY_cond $X=8.295 $Y=1.34
+ $X2=8.295 $Y2=1.552
r212 10 12 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=8.295 $Y=1.34
+ $X2=8.295 $Y2=0.86
r213 7 74 24.162 $w=1.5e-07 $l=2.13e-07 $layer=POLY_cond $X=8.22 $Y=1.765
+ $X2=8.22 $Y2=1.552
r214 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.22 $Y=1.765
+ $X2=8.22 $Y2=2.4
r215 2 59 600 $w=1.7e-07 $l=1.01573e-06 $layer=licon1_PDIFF $count=1 $X=5.415
+ $Y=1.99 $X2=5.65 $Y2=2.895
r216 1 33 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=5.285
+ $Y=0.37 $X2=5.495 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__XNOR3_4%A_27_373# 1 2 3 4 15 17 18 20 23 24 25 29 34
+ 38 39 45 46 49
c112 29 0 6.75216e-20 $X=2.3 $Y=1.1
c113 25 0 1.83967e-19 $X=1.665 $Y=1.475
c114 20 0 1.6832e-19 $X=0.33 $Y=0.615
c115 17 0 8.1711e-21 $X=2.305 $Y=2.65
r116 49 51 29.2227 $w=2.78e-07 $l=7.1e-07 $layer=LI1_cond $X=0.225 $Y=2.01
+ $X2=0.225 $Y2=2.72
r117 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=2.035
+ $X2=1.68 $Y2=2.035
r118 41 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=2.035
+ $X2=0.24 $Y2=2.035
r119 39 41 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.385 $Y=2.035
+ $X2=0.24 $Y2=2.035
r120 38 45 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.535 $Y=2.035
+ $X2=1.68 $Y2=2.035
r121 38 39 1.42326 $w=1.4e-07 $l=1.15e-06 $layer=MET1_cond $X=1.535 $Y=2.035
+ $X2=0.385 $Y2=2.035
r122 34 36 7.40856 $w=4.18e-07 $l=2.7e-07 $layer=LI1_cond $X=2.515 $Y=2.38
+ $X2=2.515 $Y2=2.65
r123 29 31 6.91466 $w=2.48e-07 $l=1.5e-07 $layer=LI1_cond $X=2.26 $Y=1.1
+ $X2=2.26 $Y2=1.25
r124 27 46 29.3909 $w=1.98e-07 $l=5.3e-07 $layer=LI1_cond $X=1.665 $Y=2.565
+ $X2=1.665 $Y2=2.035
r125 25 46 31.0545 $w=1.98e-07 $l=5.6e-07 $layer=LI1_cond $X=1.665 $Y=1.475
+ $X2=1.665 $Y2=2.035
r126 25 26 13.8873 $w=2e-07 $l=2.25e-07 $layer=LI1_cond $X=1.665 $Y=1.475
+ $X2=1.665 $Y2=1.25
r127 23 49 1.02897 $w=2.78e-07 $l=2.5e-08 $layer=LI1_cond $X=0.225 $Y=1.985
+ $X2=0.225 $Y2=2.01
r128 23 24 6.72007 $w=2.78e-07 $l=1.4e-07 $layer=LI1_cond $X=0.225 $Y=1.985
+ $X2=0.225 $Y2=1.845
r129 22 24 54.3455 $w=1.98e-07 $l=9.8e-07 $layer=LI1_cond $X=0.185 $Y=0.865
+ $X2=0.185 $Y2=1.845
r130 20 22 10.0564 $w=4.08e-07 $l=2.5e-07 $layer=LI1_cond $X=0.29 $Y=0.615
+ $X2=0.29 $Y2=0.865
r131 18 27 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=1.765 $Y=2.65
+ $X2=1.665 $Y2=2.565
r132 17 36 6.07598 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=2.305 $Y=2.65
+ $X2=2.515 $Y2=2.65
r133 17 18 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=2.305 $Y=2.65
+ $X2=1.765 $Y2=2.65
r134 16 26 1.02909 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=1.765 $Y=1.25
+ $X2=1.665 $Y2=1.25
r135 15 31 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.135 $Y=1.25
+ $X2=2.26 $Y2=1.25
r136 15 16 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.135 $Y=1.25
+ $X2=1.765 $Y2=1.25
r137 4 34 600 $w=1.7e-07 $l=5.85214e-07 $layer=licon1_PDIFF $count=1 $X=2.32
+ $Y=1.865 $X2=2.47 $Y2=2.38
r138 3 51 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.865 $X2=0.28 $Y2=2.72
r139 3 49 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.865 $X2=0.28 $Y2=2.01
r140 2 29 182 $w=1.7e-07 $l=5.94916e-07 $layer=licon1_NDIFF $count=1 $X=2.08
+ $Y=0.605 $X2=2.3 $Y2=1.1
r141 1 20 182 $w=1.7e-07 $l=2.93684e-07 $layer=licon1_NDIFF $count=1 $X=0.185
+ $Y=0.385 $X2=0.33 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_LS__XNOR3_4%VPWR 1 2 3 4 5 18 22 25 28 30 34 38 40 45 47
+ 49 54 62 70 76 79 82 85 89
r107 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r108 85 86 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r109 83 86 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.88 $Y2=3.33
r110 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r111 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r112 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r113 74 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=9.84 $Y2=3.33
r114 74 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=8.88 $Y2=3.33
r115 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r116 71 85 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.98 $Y=3.33
+ $X2=8.895 $Y2=3.33
r117 71 73 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=8.98 $Y=3.33
+ $X2=9.36 $Y2=3.33
r118 70 88 4.0045 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=9.71 $Y=3.33
+ $X2=9.895 $Y2=3.33
r119 70 73 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=9.71 $Y=3.33
+ $X2=9.36 $Y2=3.33
r120 69 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r121 68 69 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r122 65 68 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=5.04 $Y=3.33
+ $X2=7.44 $Y2=3.33
r123 63 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.72 $Y=3.33
+ $X2=4.555 $Y2=3.33
r124 63 65 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=4.72 $Y=3.33
+ $X2=5.04 $Y2=3.33
r125 62 82 12.8484 $w=1.7e-07 $l=3.12e-07 $layer=LI1_cond $X=7.485 $Y=3.33
+ $X2=7.797 $Y2=3.33
r126 62 68 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=7.485 $Y=3.33
+ $X2=7.44 $Y2=3.33
r127 61 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r128 60 61 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r129 58 61 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=4.08 $Y2=3.33
r130 58 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r131 57 60 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=4.08 $Y2=3.33
r132 57 58 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r133 55 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=0.73 $Y2=3.33
r134 55 57 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=1.2 $Y2=3.33
r135 54 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.39 $Y=3.33
+ $X2=4.555 $Y2=3.33
r136 54 60 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=4.39 $Y=3.33
+ $X2=4.08 $Y2=3.33
r137 52 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r138 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r139 49 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.73 $Y2=3.33
r140 49 51 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.24 $Y2=3.33
r141 47 69 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=7.44 $Y2=3.33
r142 47 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r143 47 65 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r144 45 46 3.52857 $w=6.23e-07 $l=1.2e-07 $layer=LI1_cond $X=7.797 $Y=2.41
+ $X2=7.797 $Y2=2.29
r145 40 43 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=9.835 $Y=1.985
+ $X2=9.835 $Y2=2.815
r146 38 88 3.13866 $w=2.5e-07 $l=1.11018e-07 $layer=LI1_cond $X=9.835 $Y=3.245
+ $X2=9.895 $Y2=3.33
r147 38 43 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=9.835 $Y=3.245
+ $X2=9.835 $Y2=2.815
r148 34 37 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=8.895 $Y=1.985
+ $X2=8.895 $Y2=2.815
r149 32 85 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.895 $Y=3.245
+ $X2=8.895 $Y2=3.33
r150 32 37 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=8.895 $Y=3.245
+ $X2=8.895 $Y2=2.815
r151 31 82 12.8484 $w=1.7e-07 $l=3.13e-07 $layer=LI1_cond $X=8.11 $Y=3.33
+ $X2=7.797 $Y2=3.33
r152 30 85 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.81 $Y=3.33
+ $X2=8.895 $Y2=3.33
r153 30 31 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=8.81 $Y=3.33 $X2=8.11
+ $Y2=3.33
r154 28 46 7.72815 $w=4.23e-07 $l=2.85e-07 $layer=LI1_cond $X=7.897 $Y=2.005
+ $X2=7.897 $Y2=2.29
r155 25 82 2.61429 $w=6.25e-07 $l=8.5e-08 $layer=LI1_cond $X=7.797 $Y=3.245
+ $X2=7.797 $Y2=3.33
r156 24 45 3.67435 $w=6.23e-07 $l=1.92e-07 $layer=LI1_cond $X=7.797 $Y=2.602
+ $X2=7.797 $Y2=2.41
r157 24 25 12.3053 $w=6.23e-07 $l=6.43e-07 $layer=LI1_cond $X=7.797 $Y=2.602
+ $X2=7.797 $Y2=3.245
r158 20 79 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.555 $Y=3.245
+ $X2=4.555 $Y2=3.33
r159 20 22 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=4.555 $Y=3.245
+ $X2=4.555 $Y2=2.815
r160 16 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=3.33
r161 16 18 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=2.375
r162 5 43 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=9.645
+ $Y=1.84 $X2=9.795 $Y2=2.815
r163 5 40 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=9.645
+ $Y=1.84 $X2=9.795 $Y2=1.985
r164 4 37 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=8.745
+ $Y=1.84 $X2=8.895 $Y2=2.815
r165 4 34 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=8.745
+ $Y=1.84 $X2=8.895 $Y2=1.985
r166 3 45 150 $w=1.7e-07 $l=1.15022e-06 $layer=licon1_PDIFF $count=4 $X=7.095
+ $Y=1.84 $X2=7.995 $Y2=2.41
r167 3 28 600 $w=1.7e-07 $l=7.52994e-07 $layer=licon1_PDIFF $count=1 $X=7.095
+ $Y=1.84 $X2=7.77 $Y2=2.005
r168 2 22 600 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=4.405
+ $Y=1.84 $X2=4.555 $Y2=2.815
r169 1 18 300 $w=1.7e-07 $l=5.80172e-07 $layer=licon1_PDIFF $count=2 $X=0.58
+ $Y=1.865 $X2=0.73 $Y2=2.375
.ends

.subckt PM_SKY130_FD_SC_LS__XNOR3_4%A_324_373# 1 2 3 4 14 15 16 18 20 22 23 25
+ 30 33 35 36 42 43 46
c128 16 0 2.40512e-19 $X=2.245 $Y=1.59
r129 43 47 7.46954 $w=2.68e-07 $l=1.75e-07 $layer=LI1_cond $X=5.04 $Y=2.085
+ $X2=4.865 $Y2=2.085
r130 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=2.035
+ $X2=5.04 $Y2=2.035
r131 38 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=2.035
+ $X2=2.16 $Y2=2.035
r132 36 38 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.305 $Y=2.035
+ $X2=2.16 $Y2=2.035
r133 35 42 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.895 $Y=2.035
+ $X2=5.04 $Y2=2.035
r134 35 36 3.20544 $w=1.4e-07 $l=2.59e-06 $layer=MET1_cond $X=4.895 $Y=2.035
+ $X2=2.305 $Y2=2.035
r135 27 30 8.75857 $w=2.48e-07 $l=1.9e-07 $layer=LI1_cond $X=2.655 $Y=1.08
+ $X2=2.845 $Y2=1.08
r136 23 33 32.9995 $w=1.98e-07 $l=5.9e-07 $layer=LI1_cond $X=5.995 $Y=1.28
+ $X2=5.405 $Y2=1.28
r137 23 25 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=5.995 $Y=1.18
+ $X2=5.995 $Y2=0.81
r138 22 33 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=4.95 $Y=1.295
+ $X2=5.405 $Y2=1.295
r139 20 47 3.44395 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.865 $Y=1.95
+ $X2=4.865 $Y2=2.085
r140 19 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.865 $Y=1.38
+ $X2=4.95 $Y2=1.295
r141 19 20 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=4.865 $Y=1.38
+ $X2=4.865 $Y2=1.95
r142 17 27 2.04652 $w=2e-07 $l=1.25e-07 $layer=LI1_cond $X=2.655 $Y=1.205
+ $X2=2.655 $Y2=1.08
r143 17 18 16.6364 $w=1.98e-07 $l=3e-07 $layer=LI1_cond $X=2.655 $Y=1.205
+ $X2=2.655 $Y2=1.505
r144 15 18 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=2.555 $Y=1.59
+ $X2=2.655 $Y2=1.505
r145 15 16 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=2.555 $Y=1.59
+ $X2=2.245 $Y2=1.59
r146 14 46 1.05747 $w=3.1e-07 $l=2.5e-08 $layer=LI1_cond $X=2.09 $Y=1.965
+ $X2=2.09 $Y2=1.99
r147 13 16 7.59919 $w=1.7e-07 $l=1.92873e-07 $layer=LI1_cond $X=2.09 $Y=1.675
+ $X2=2.245 $Y2=1.59
r148 13 14 10.7809 $w=3.08e-07 $l=2.9e-07 $layer=LI1_cond $X=2.09 $Y=1.675
+ $X2=2.09 $Y2=1.965
r149 4 43 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=4.97
+ $Y=1.99 $X2=5.115 $Y2=2.135
r150 3 46 600 $w=1.7e-07 $l=4.58258e-07 $layer=licon1_PDIFF $count=1 $X=1.62
+ $Y=1.865 $X2=2.02 $Y2=1.99
r151 2 25 182 $w=1.7e-07 $l=5.11664e-07 $layer=licon1_NDIFF $count=1 $X=5.84
+ $Y=0.37 $X2=5.995 $Y2=0.81
r152 1 30 182 $w=1.7e-07 $l=5.04455e-07 $layer=licon1_NDIFF $count=1 $X=2.695
+ $Y=0.605 $X2=2.845 $Y2=1.04
.ends

.subckt PM_SKY130_FD_SC_LS__XNOR3_4%A_321_77# 1 2 3 4 15 19 21 22 24 25 29 31 36
+ 37 38 41
c131 37 0 2.17577e-19 $X=2.725 $Y=0.69
c132 22 0 2.21365e-20 $X=3.145 $Y=2.455
r133 38 40 10.6978 $w=5.36e-07 $l=4.7e-07 $layer=LI1_cond $X=4.525 $Y=0.69
+ $X2=4.995 $Y2=0.69
r134 36 37 9.92344 $w=1.88e-07 $l=1.7e-07 $layer=LI1_cond $X=2.555 $Y=0.69
+ $X2=2.725 $Y2=0.69
r135 31 34 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=1.79 $Y=0.68
+ $X2=1.79 $Y2=0.795
r136 27 29 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=6.145 $Y=2.39
+ $X2=6.145 $Y2=2.135
r137 26 41 5.16603 $w=1.7e-07 $l=8.9861e-08 $layer=LI1_cond $X=4.61 $Y=2.475
+ $X2=4.525 $Y2=2.465
r138 25 27 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.02 $Y=2.475
+ $X2=6.145 $Y2=2.39
r139 25 26 91.9893 $w=1.68e-07 $l=1.41e-06 $layer=LI1_cond $X=6.02 $Y=2.475
+ $X2=4.61 $Y2=2.475
r140 24 41 1.34256 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.525 $Y=2.37
+ $X2=4.525 $Y2=2.465
r141 23 38 7.59541 $w=1.7e-07 $l=3.4e-07 $layer=LI1_cond $X=4.525 $Y=1.03
+ $X2=4.525 $Y2=0.69
r142 23 24 87.4225 $w=1.68e-07 $l=1.34e-06 $layer=LI1_cond $X=4.525 $Y=1.03
+ $X2=4.525 $Y2=2.37
r143 21 41 5.16603 $w=1.7e-07 $l=8.9861e-08 $layer=LI1_cond $X=4.44 $Y=2.455
+ $X2=4.525 $Y2=2.465
r144 21 22 84.4866 $w=1.68e-07 $l=1.295e-06 $layer=LI1_cond $X=4.44 $Y=2.455
+ $X2=3.145 $Y2=2.455
r145 17 22 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.02 $Y=2.37
+ $X2=3.145 $Y2=2.455
r146 17 19 15.2122 $w=2.48e-07 $l=3.3e-07 $layer=LI1_cond $X=3.02 $Y=2.37
+ $X2=3.02 $Y2=2.04
r147 15 38 8.11642 $w=5.36e-07 $l=8.9861e-08 $layer=LI1_cond $X=4.44 $Y=0.7
+ $X2=4.525 $Y2=0.69
r148 15 37 111.888 $w=1.68e-07 $l=1.715e-06 $layer=LI1_cond $X=4.44 $Y=0.7
+ $X2=2.725 $Y2=0.7
r149 14 31 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.955 $Y=0.68
+ $X2=1.79 $Y2=0.68
r150 14 36 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=1.955 $Y=0.68
+ $X2=2.555 $Y2=0.68
r151 4 29 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=6.035
+ $Y=1.99 $X2=6.185 $Y2=2.135
r152 3 19 300 $w=1.7e-07 $l=2.84341e-07 $layer=licon1_PDIFF $count=2 $X=2.77
+ $Y=1.865 $X2=2.98 $Y2=2.04
r153 2 40 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=4.85
+ $Y=0.37 $X2=4.995 $Y2=0.515
r154 1 34 182 $w=1.7e-07 $l=4.93913e-07 $layer=licon1_NDIFF $count=1 $X=1.605
+ $Y=0.385 $X2=1.79 $Y2=0.795
.ends

.subckt PM_SKY130_FD_SC_LS__XNOR3_4%X 1 2 3 4 15 19 22 25 28 29 30 31 32 33 34
+ 35 36 37 38 58
r58 56 58 1.29853 $w=3.53e-07 $l=4e-08 $layer=LI1_cond $X=9.357 $Y=1.625
+ $X2=9.357 $Y2=1.665
r59 37 38 12.0114 $w=3.53e-07 $l=3.7e-07 $layer=LI1_cond $X=9.357 $Y=2.405
+ $X2=9.357 $Y2=2.775
r60 36 37 13.6345 $w=3.53e-07 $l=4.2e-07 $layer=LI1_cond $X=9.357 $Y=1.985
+ $X2=9.357 $Y2=2.405
r61 35 47 3.3083 $w=3.42e-07 $l=1.08305e-07 $layer=LI1_cond $X=9.357 $Y=1.522
+ $X2=9.37 $Y2=1.42
r62 35 56 3.3083 $w=3.42e-07 $l=1.03e-07 $layer=LI1_cond $X=9.357 $Y=1.522
+ $X2=9.357 $Y2=1.625
r63 35 36 9.67403 $w=3.53e-07 $l=2.98e-07 $layer=LI1_cond $X=9.357 $Y=1.687
+ $X2=9.357 $Y2=1.985
r64 35 58 0.71419 $w=3.53e-07 $l=2.2e-08 $layer=LI1_cond $X=9.357 $Y=1.687
+ $X2=9.357 $Y2=1.665
r65 34 47 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=9.37 $Y=1.295
+ $X2=9.37 $Y2=1.42
r66 33 34 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=9.37 $Y=0.925
+ $X2=9.37 $Y2=1.295
r67 32 33 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=9.37 $Y=0.555
+ $X2=9.37 $Y2=0.925
r68 28 29 8.51103 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=8.46 $Y=2.005
+ $X2=8.46 $Y2=1.84
r69 26 31 1.0233 $w=2.05e-07 $l=1.03e-07 $layer=LI1_cond $X=8.675 $Y=1.522
+ $X2=8.572 $Y2=1.522
r70 25 35 3.24129 $w=2.05e-07 $l=1.77e-07 $layer=LI1_cond $X=9.18 $Y=1.522
+ $X2=9.357 $Y2=1.522
r71 25 26 27.3215 $w=2.03e-07 $l=5.05e-07 $layer=LI1_cond $X=9.18 $Y=1.522
+ $X2=8.675 $Y2=1.522
r72 23 31 5.56063 $w=1.87e-07 $l=1.11176e-07 $layer=LI1_cond $X=8.555 $Y=1.625
+ $X2=8.572 $Y2=1.522
r73 23 29 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=8.555 $Y=1.625
+ $X2=8.555 $Y2=1.84
r74 22 31 5.56063 $w=1.87e-07 $l=1.02e-07 $layer=LI1_cond $X=8.572 $Y=1.42
+ $X2=8.572 $Y2=1.522
r75 22 30 13.5255 $w=2.03e-07 $l=2.5e-07 $layer=LI1_cond $X=8.572 $Y=1.42
+ $X2=8.572 $Y2=1.17
r76 17 30 7.40596 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=8.51 $Y=1.005
+ $X2=8.51 $Y2=1.17
r77 17 19 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=8.51 $Y=1.005
+ $X2=8.51 $Y2=0.635
r78 13 28 0.480185 $w=3.58e-07 $l=1.5e-08 $layer=LI1_cond $X=8.46 $Y=2.02
+ $X2=8.46 $Y2=2.005
r79 13 15 25.4498 $w=3.58e-07 $l=7.95e-07 $layer=LI1_cond $X=8.46 $Y=2.02
+ $X2=8.46 $Y2=2.815
r80 4 38 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=9.195
+ $Y=1.84 $X2=9.345 $Y2=2.815
r81 4 36 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=9.195
+ $Y=1.84 $X2=9.345 $Y2=1.985
r82 3 28 400 $w=1.7e-07 $l=2.2798e-07 $layer=licon1_PDIFF $count=1 $X=8.295
+ $Y=1.84 $X2=8.445 $Y2=2.005
r83 3 15 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=8.295
+ $Y=1.84 $X2=8.445 $Y2=2.815
r84 2 32 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.23
+ $Y=0.49 $X2=9.37 $Y2=0.635
r85 1 19 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.37
+ $Y=0.49 $X2=8.51 $Y2=0.635
.ends

.subckt PM_SKY130_FD_SC_LS__XNOR3_4%VGND 1 2 3 4 5 20 24 26 30 32 33 36 38 40 42
+ 44 52 58 61 77 81
c100 20 0 1.02947e-19 $X=0.83 $Y=0.615
r101 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r102 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r103 74 75 0.585834 $w=8.33e-07 $l=4e-08 $layer=LI1_cond $X=8 $Y=0.377 $X2=8.04
+ $Y2=0.377
r104 72 78 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.88
+ $Y2=0
r105 71 74 1.17167 $w=8.33e-07 $l=8e-08 $layer=LI1_cond $X=7.92 $Y=0.377 $X2=8
+ $Y2=0.377
r106 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r107 69 71 5.71188 $w=8.33e-07 $l=3.9e-07 $layer=LI1_cond $X=7.53 $Y=0.377
+ $X2=7.92 $Y2=0.377
r108 67 69 6.81032 $w=8.33e-07 $l=4.65e-07 $layer=LI1_cond $X=7.065 $Y=0.377
+ $X2=7.53 $Y2=0.377
r109 65 72 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.92
+ $Y2=0
r110 64 67 1.53782 $w=8.33e-07 $l=1.05e-07 $layer=LI1_cond $X=6.96 $Y=0.377
+ $X2=7.065 $Y2=0.377
r111 64 65 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r112 61 62 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r113 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r114 56 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0 $X2=9.84
+ $Y2=0
r115 56 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0 $X2=8.88
+ $Y2=0
r116 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r117 53 77 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.025 $Y=0 $X2=8.94
+ $Y2=0
r118 53 55 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=9.025 $Y=0
+ $X2=9.36 $Y2=0
r119 52 80 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=9.715 $Y=0
+ $X2=9.897 $Y2=0
r120 52 55 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=9.715 $Y=0
+ $X2=9.36 $Y2=0
r121 51 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r122 50 51 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r123 48 51 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=4.08
+ $Y2=0
r124 48 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r125 47 50 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=4.08
+ $Y2=0
r126 47 48 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=1.2 $Y=0
+ $X2=1.2 $Y2=0
r127 45 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.995 $Y=0 $X2=0.83
+ $Y2=0
r128 45 47 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=0.995 $Y=0 $X2=1.2
+ $Y2=0
r129 44 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.27 $Y=0 $X2=4.435
+ $Y2=0
r130 44 50 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=4.27 $Y=0 $X2=4.08
+ $Y2=0
r131 42 65 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=6.96 $Y2=0
r132 42 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.56
+ $Y2=0
r133 38 80 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=9.84 $Y=0.085
+ $X2=9.897 $Y2=0
r134 38 40 25.3537 $w=2.48e-07 $l=5.5e-07 $layer=LI1_cond $X=9.84 $Y=0.085
+ $X2=9.84 $Y2=0.635
r135 34 77 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.94 $Y=0.085
+ $X2=8.94 $Y2=0
r136 34 36 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=8.94 $Y=0.085
+ $X2=8.94 $Y2=0.635
r137 33 75 11.282 $w=8.33e-07 $l=4.35033e-07 $layer=LI1_cond $X=8.165 $Y=0
+ $X2=8.04 $Y2=0.377
r138 32 77 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.855 $Y=0 $X2=8.94
+ $Y2=0
r139 32 33 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=8.855 $Y=0 $X2=8.165
+ $Y2=0
r140 28 75 7.9472 $w=2.5e-07 $l=4.63e-07 $layer=LI1_cond $X=8.04 $Y=0.84
+ $X2=8.04 $Y2=0.377
r141 28 30 7.60612 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=8.04 $Y=0.84
+ $X2=8.04 $Y2=1.005
r142 27 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.6 $Y=0 $X2=4.435
+ $Y2=0
r143 26 64 10.33 $w=8.33e-07 $l=4.05893e-07 $layer=LI1_cond $X=6.9 $Y=0 $X2=6.96
+ $Y2=0.377
r144 26 27 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=6.9 $Y=0 $X2=4.6
+ $Y2=0
r145 22 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.435 $Y=0.085
+ $X2=4.435 $Y2=0
r146 22 24 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=4.435 $Y=0.085
+ $X2=4.435 $Y2=0.36
r147 18 58 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.83 $Y=0.085
+ $X2=0.83 $Y2=0
r148 18 20 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=0.83 $Y=0.085
+ $X2=0.83 $Y2=0.615
r149 5 40 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.66
+ $Y=0.49 $X2=9.8 $Y2=0.635
r150 4 36 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.8
+ $Y=0.49 $X2=8.94 $Y2=0.635
r151 3 74 91 $w=1.7e-07 $l=1.3763e-06 $layer=licon1_NDIFF $count=2 $X=6.845
+ $Y=0.81 $X2=8 $Y2=0.325
r152 3 69 91 $w=1.7e-07 $l=8.95237e-07 $layer=licon1_NDIFF $count=2 $X=6.845
+ $Y=0.81 $X2=7.53 $Y2=0.325
r153 3 67 91 $w=1.7e-07 $l=5.84744e-07 $layer=licon1_NDIFF $count=2 $X=6.845
+ $Y=0.81 $X2=7.065 $Y2=0.325
r154 3 30 182 $w=1.7e-07 $l=1.32893e-06 $layer=licon1_NDIFF $count=1 $X=6.845
+ $Y=0.81 $X2=8.08 $Y2=1.005
r155 2 24 182 $w=1.7e-07 $l=2.59037e-07 $layer=licon1_NDIFF $count=1 $X=4.215
+ $Y=0.445 $X2=4.435 $Y2=0.36
r156 1 20 182 $w=1.7e-07 $l=3.18119e-07 $layer=licon1_NDIFF $count=1 $X=0.62
+ $Y=0.385 $X2=0.83 $Y2=0.615
.ends

