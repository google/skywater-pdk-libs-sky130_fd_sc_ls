* File: sky130_fd_sc_ls__o311a_1.pxi.spice
* Created: Fri Aug 28 13:51:20 2020
* 
x_PM_SKY130_FD_SC_LS__O311A_1%C1 N_C1_c_79_n N_C1_c_84_n N_C1_M1006_g
+ N_C1_M1002_g C1 N_C1_c_82_n PM_SKY130_FD_SC_LS__O311A_1%C1
x_PM_SKY130_FD_SC_LS__O311A_1%B1 N_B1_M1001_g N_B1_c_110_n N_B1_c_114_n
+ N_B1_M1009_g B1 N_B1_c_112_n PM_SKY130_FD_SC_LS__O311A_1%B1
x_PM_SKY130_FD_SC_LS__O311A_1%A2 N_A2_M1005_g N_A2_c_149_n N_A2_M1010_g
+ N_A2_c_150_n N_A2_c_165_p N_A2_c_195_p N_A2_c_151_n A2 N_A2_c_152_n
+ N_A2_c_153_n PM_SKY130_FD_SC_LS__O311A_1%A2
x_PM_SKY130_FD_SC_LS__O311A_1%A3 N_A3_c_221_n N_A3_M1008_g N_A3_c_222_n
+ N_A3_c_223_n N_A3_c_217_n N_A3_M1003_g A3 A3 A3 N_A3_c_219_n N_A3_c_220_n
+ PM_SKY130_FD_SC_LS__O311A_1%A3
x_PM_SKY130_FD_SC_LS__O311A_1%A1 N_A1_c_262_n N_A1_c_267_n N_A1_M1007_g
+ N_A1_M1011_g A1 N_A1_c_263_n N_A1_c_264_n N_A1_c_265_n
+ PM_SKY130_FD_SC_LS__O311A_1%A1
x_PM_SKY130_FD_SC_LS__O311A_1%A_31_387# N_A_31_387#_M1002_s N_A_31_387#_M1006_s
+ N_A_31_387#_M1009_d N_A_31_387#_c_304_n N_A_31_387#_M1000_g
+ N_A_31_387#_M1004_g N_A_31_387#_c_315_n N_A_31_387#_c_306_n
+ N_A_31_387#_c_307_n N_A_31_387#_c_308_n N_A_31_387#_c_309_n
+ N_A_31_387#_c_318_n N_A_31_387#_c_334_n N_A_31_387#_c_319_n
+ N_A_31_387#_c_320_n N_A_31_387#_c_310_n N_A_31_387#_c_311_n
+ N_A_31_387#_c_312_n N_A_31_387#_c_313_n PM_SKY130_FD_SC_LS__O311A_1%A_31_387#
x_PM_SKY130_FD_SC_LS__O311A_1%VPWR N_VPWR_M1006_d N_VPWR_M1007_d N_VPWR_c_428_n
+ N_VPWR_c_429_n VPWR N_VPWR_c_430_n N_VPWR_c_431_n N_VPWR_c_432_n
+ N_VPWR_c_427_n N_VPWR_c_434_n N_VPWR_c_435_n PM_SKY130_FD_SC_LS__O311A_1%VPWR
x_PM_SKY130_FD_SC_LS__O311A_1%X N_X_M1004_d N_X_M1000_d N_X_c_480_n N_X_c_481_n
+ N_X_c_477_n X X X PM_SKY130_FD_SC_LS__O311A_1%X
x_PM_SKY130_FD_SC_LS__O311A_1%A_209_74# N_A_209_74#_M1001_d N_A_209_74#_M1003_d
+ N_A_209_74#_c_503_n N_A_209_74#_c_506_n N_A_209_74#_c_504_n
+ PM_SKY130_FD_SC_LS__O311A_1%A_209_74#
x_PM_SKY130_FD_SC_LS__O311A_1%VGND N_VGND_M1005_d N_VGND_M1011_d N_VGND_c_531_n
+ N_VGND_c_522_n VGND N_VGND_c_523_n N_VGND_c_524_n N_VGND_c_525_n
+ N_VGND_c_526_n PM_SKY130_FD_SC_LS__O311A_1%VGND
cc_1 VNB N_C1_c_79_n 0.0154393f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.77
cc_2 VNB N_C1_M1002_g 0.02469f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=0.69
cc_3 VNB C1 0.0121164f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_C1_c_82_n 0.0546617f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.305
cc_5 VNB N_B1_M1001_g 0.0196196f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.86
cc_6 VNB N_B1_c_110_n 0.0130036f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.14
cc_7 VNB B1 0.00308495f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_8 VNB N_B1_c_112_n 0.0295848f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.305
cc_9 VNB N_A2_M1005_g 0.0210444f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.86
cc_10 VNB N_A2_c_149_n 0.0257012f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=2.435
cc_11 VNB N_A2_c_150_n 0.00351602f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A2_c_151_n 0.00486902f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.305
cc_13 VNB N_A2_c_152_n 0.0298977f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A2_c_153_n 0.00245544f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A3_c_217_n 0.0114682f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=0.69
cc_16 VNB A3 0.00138988f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A3_c_219_n 0.0473444f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A3_c_220_n 0.0213502f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A1_c_262_n 0.011579f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.77
cc_20 VNB N_A1_c_263_n 0.0340747f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.305
cc_21 VNB N_A1_c_264_n 0.0166185f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.305
cc_22 VNB N_A1_c_265_n 0.0221309f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.305
cc_23 VNB N_A_31_387#_c_304_n 0.0291516f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_24 VNB N_A_31_387#_M1004_g 0.0312993f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_31_387#_c_306_n 0.019793f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_31_387#_c_307_n 0.00527983f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_31_387#_c_308_n 0.0106214f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_31_387#_c_309_n 0.00304476f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_31_387#_c_310_n 0.00424542f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_31_387#_c_311_n 7.98615e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_31_387#_c_312_n 0.00695823f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_31_387#_c_313_n 0.00336822f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VPWR_c_427_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_X_c_477_n 0.0250799f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB X 0.0267037f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.305
cc_36 VNB X 0.013364f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.305
cc_37 VNB N_A_209_74#_c_503_n 0.00406087f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=0.69
cc_38 VNB N_A_209_74#_c_504_n 0.0147102f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.305
cc_39 VNB N_VGND_c_522_n 0.00647919f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.305
cc_40 VNB N_VGND_c_523_n 0.0873829f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.305
cc_41 VNB N_VGND_c_524_n 0.0193554f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_525_n 0.261122f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_526_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VPB N_C1_c_79_n 0.00701719f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=1.77
cc_45 VPB N_C1_c_84_n 0.0269814f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=1.86
cc_46 VPB N_B1_c_110_n 0.00609143f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=1.14
cc_47 VPB N_B1_c_114_n 0.021265f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=0.69
cc_48 VPB N_A2_c_149_n 0.03817f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=2.435
cc_49 VPB N_A2_c_150_n 0.0017688f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_A2_c_151_n 0.00175132f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.305
cc_51 VPB N_A3_c_221_n 0.0179776f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=1.47
cc_52 VPB N_A3_c_222_n 0.03749f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=2.435
cc_53 VPB N_A3_c_223_n 0.00778788f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=2.435
cc_54 VPB N_A3_c_217_n 0.00271961f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=0.69
cc_55 VPB A3 0.00233286f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_A1_c_262_n 0.0052455f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=1.77
cc_57 VPB N_A1_c_267_n 0.0232475f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=1.86
cc_58 VPB N_A_31_387#_c_304_n 0.0328318f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_59 VPB N_A_31_387#_c_315_n 0.047466f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_A_31_387#_c_308_n 0.00309737f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_A_31_387#_c_309_n 0.00935005f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_A_31_387#_c_318_n 0.00268475f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_A_31_387#_c_319_n 0.0122419f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_A_31_387#_c_320_n 9.40627e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_A_31_387#_c_310_n 0.00552421f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_A_31_387#_c_311_n 7.96937e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_A_31_387#_c_313_n 0.00368195f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_428_n 0.0115862f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_429_n 0.0105324f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_430_n 0.0198977f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_431_n 0.0607653f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_432_n 0.0193973f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_427_n 0.0836881f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_434_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_435_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_X_c_480_n 0.0367571f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_X_c_481_n 0.00768928f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.305
cc_78 VPB N_X_c_477_n 0.0132189f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 N_C1_M1002_g N_B1_M1001_g 0.0311169f $X=0.58 $Y=0.69 $X2=0 $Y2=0
cc_80 N_C1_c_79_n N_B1_c_110_n 0.00578733f $X=0.525 $Y=1.77 $X2=0 $Y2=0
cc_81 N_C1_c_84_n N_B1_c_114_n 0.0311397f $X=0.525 $Y=1.86 $X2=0 $Y2=0
cc_82 N_C1_c_82_n B1 3.30694e-19 $X=0.58 $Y=1.305 $X2=0 $Y2=0
cc_83 N_C1_c_82_n N_B1_c_112_n 0.0311169f $X=0.58 $Y=1.305 $X2=0 $Y2=0
cc_84 N_C1_c_84_n N_A_31_387#_c_315_n 0.0163444f $X=0.525 $Y=1.86 $X2=0 $Y2=0
cc_85 N_C1_M1002_g N_A_31_387#_c_306_n 0.00844889f $X=0.58 $Y=0.69 $X2=0 $Y2=0
cc_86 N_C1_c_79_n N_A_31_387#_c_307_n 0.00868484f $X=0.525 $Y=1.77 $X2=0 $Y2=0
cc_87 N_C1_M1002_g N_A_31_387#_c_307_n 0.00858018f $X=0.58 $Y=0.69 $X2=0 $Y2=0
cc_88 C1 N_A_31_387#_c_307_n 0.0233985f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_89 N_C1_c_82_n N_A_31_387#_c_307_n 0.00911304f $X=0.58 $Y=1.305 $X2=0 $Y2=0
cc_90 N_C1_c_79_n N_A_31_387#_c_309_n 0.0106881f $X=0.525 $Y=1.77 $X2=0 $Y2=0
cc_91 N_C1_c_84_n N_A_31_387#_c_309_n 0.00867655f $X=0.525 $Y=1.86 $X2=0 $Y2=0
cc_92 C1 N_A_31_387#_c_309_n 0.0206681f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_93 N_C1_c_82_n N_A_31_387#_c_309_n 0.00704075f $X=0.58 $Y=1.305 $X2=0 $Y2=0
cc_94 N_C1_c_84_n N_A_31_387#_c_334_n 6.84479e-19 $X=0.525 $Y=1.86 $X2=0 $Y2=0
cc_95 N_C1_M1002_g N_A_31_387#_c_312_n 0.00848905f $X=0.58 $Y=0.69 $X2=0 $Y2=0
cc_96 C1 N_A_31_387#_c_312_n 0.0155323f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_97 N_C1_c_82_n N_A_31_387#_c_312_n 0.00717614f $X=0.58 $Y=1.305 $X2=0 $Y2=0
cc_98 N_C1_c_84_n N_VPWR_c_428_n 0.00909794f $X=0.525 $Y=1.86 $X2=0 $Y2=0
cc_99 N_C1_c_84_n N_VPWR_c_430_n 0.00544739f $X=0.525 $Y=1.86 $X2=0 $Y2=0
cc_100 N_C1_c_84_n N_VPWR_c_427_n 0.00537853f $X=0.525 $Y=1.86 $X2=0 $Y2=0
cc_101 N_C1_M1002_g N_VGND_c_523_n 0.00434272f $X=0.58 $Y=0.69 $X2=0 $Y2=0
cc_102 N_C1_M1002_g N_VGND_c_525_n 0.00442932f $X=0.58 $Y=0.69 $X2=0 $Y2=0
cc_103 N_B1_M1001_g N_A2_M1005_g 0.0159664f $X=0.97 $Y=0.69 $X2=0 $Y2=0
cc_104 N_B1_c_110_n N_A2_c_150_n 0.00467281f $X=1.075 $Y=1.77 $X2=0 $Y2=0
cc_105 B1 N_A2_c_152_n 0.00193925f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_106 N_B1_c_112_n N_A2_c_152_n 0.020587f $X=1.06 $Y=1.305 $X2=0 $Y2=0
cc_107 B1 N_A2_c_153_n 0.0265356f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_108 N_B1_c_112_n N_A2_c_153_n 3.50521e-19 $X=1.06 $Y=1.305 $X2=0 $Y2=0
cc_109 N_B1_c_114_n N_A3_c_221_n 0.00860888f $X=1.075 $Y=1.86 $X2=-0.19
+ $Y2=-0.245
cc_110 N_B1_c_110_n N_A3_c_223_n 0.00711621f $X=1.075 $Y=1.77 $X2=0 $Y2=0
cc_111 N_B1_c_114_n N_A_31_387#_c_315_n 7.20022e-19 $X=1.075 $Y=1.86 $X2=0 $Y2=0
cc_112 N_B1_M1001_g N_A_31_387#_c_306_n 0.00129834f $X=0.97 $Y=0.69 $X2=0 $Y2=0
cc_113 N_B1_M1001_g N_A_31_387#_c_307_n 0.00553928f $X=0.97 $Y=0.69 $X2=0 $Y2=0
cc_114 N_B1_c_110_n N_A_31_387#_c_307_n 0.00341339f $X=1.075 $Y=1.77 $X2=0 $Y2=0
cc_115 B1 N_A_31_387#_c_307_n 0.0249634f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_116 N_B1_c_110_n N_A_31_387#_c_308_n 0.00857366f $X=1.075 $Y=1.77 $X2=0 $Y2=0
cc_117 N_B1_c_114_n N_A_31_387#_c_308_n 0.00816456f $X=1.075 $Y=1.86 $X2=0 $Y2=0
cc_118 B1 N_A_31_387#_c_308_n 0.0283256f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_119 N_B1_c_112_n N_A_31_387#_c_308_n 0.00414882f $X=1.06 $Y=1.305 $X2=0 $Y2=0
cc_120 N_B1_c_114_n N_A_31_387#_c_318_n 0.0020229f $X=1.075 $Y=1.86 $X2=0 $Y2=0
cc_121 N_B1_c_114_n N_A_31_387#_c_334_n 0.0129347f $X=1.075 $Y=1.86 $X2=0 $Y2=0
cc_122 N_B1_M1001_g N_A_31_387#_c_312_n 0.00138573f $X=0.97 $Y=0.69 $X2=0 $Y2=0
cc_123 N_B1_c_114_n N_VPWR_c_428_n 0.00909759f $X=1.075 $Y=1.86 $X2=0 $Y2=0
cc_124 N_B1_c_114_n N_VPWR_c_431_n 0.0054367f $X=1.075 $Y=1.86 $X2=0 $Y2=0
cc_125 N_B1_c_114_n N_VPWR_c_427_n 0.00537853f $X=1.075 $Y=1.86 $X2=0 $Y2=0
cc_126 N_B1_M1001_g N_A_209_74#_c_503_n 0.00276611f $X=0.97 $Y=0.69 $X2=0 $Y2=0
cc_127 B1 N_A_209_74#_c_506_n 0.0169224f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_128 N_B1_c_112_n N_A_209_74#_c_506_n 0.00410213f $X=1.06 $Y=1.305 $X2=0 $Y2=0
cc_129 N_B1_M1001_g N_VGND_c_523_n 0.00461464f $X=0.97 $Y=0.69 $X2=0 $Y2=0
cc_130 N_B1_M1001_g N_VGND_c_525_n 0.00910057f $X=0.97 $Y=0.69 $X2=0 $Y2=0
cc_131 N_A2_c_150_n N_A3_c_221_n 0.00920271f $X=1.72 $Y=2.32 $X2=-0.19
+ $Y2=-0.245
cc_132 N_A2_c_150_n N_A3_c_222_n 0.0123672f $X=1.72 $Y=2.32 $X2=0 $Y2=0
cc_133 N_A2_c_165_p N_A3_c_222_n 0.00484151f $X=2.515 $Y=2.405 $X2=0 $Y2=0
cc_134 N_A2_c_153_n N_A3_c_222_n 2.41637e-19 $X=1.72 $Y=1.305 $X2=0 $Y2=0
cc_135 N_A2_c_152_n N_A3_c_223_n 0.0195985f $X=1.6 $Y=1.305 $X2=0 $Y2=0
cc_136 N_A2_c_153_n N_A3_c_223_n 0.00126382f $X=1.72 $Y=1.305 $X2=0 $Y2=0
cc_137 N_A2_c_149_n N_A3_c_217_n 0.0110399f $X=2.605 $Y=1.86 $X2=0 $Y2=0
cc_138 N_A2_c_150_n N_A3_c_217_n 0.00456493f $X=1.72 $Y=2.32 $X2=0 $Y2=0
cc_139 N_A2_c_151_n N_A3_c_217_n 4.03153e-19 $X=2.68 $Y=1.61 $X2=0 $Y2=0
cc_140 N_A2_c_149_n A3 0.00518787f $X=2.605 $Y=1.86 $X2=0 $Y2=0
cc_141 N_A2_c_150_n A3 0.0510888f $X=1.72 $Y=2.32 $X2=0 $Y2=0
cc_142 N_A2_c_165_p A3 0.0266856f $X=2.515 $Y=2.405 $X2=0 $Y2=0
cc_143 N_A2_c_151_n A3 0.0407438f $X=2.68 $Y=1.61 $X2=0 $Y2=0
cc_144 N_A2_c_152_n A3 3.76918e-19 $X=1.6 $Y=1.305 $X2=0 $Y2=0
cc_145 N_A2_c_153_n A3 0.02617f $X=1.72 $Y=1.305 $X2=0 $Y2=0
cc_146 N_A2_M1005_g N_A3_c_219_n 0.00206579f $X=1.51 $Y=0.69 $X2=0 $Y2=0
cc_147 N_A2_c_149_n N_A3_c_219_n 3.04703e-19 $X=2.605 $Y=1.86 $X2=0 $Y2=0
cc_148 N_A2_c_152_n N_A3_c_219_n 0.0205549f $X=1.6 $Y=1.305 $X2=0 $Y2=0
cc_149 N_A2_c_153_n N_A3_c_219_n 0.00184761f $X=1.72 $Y=1.305 $X2=0 $Y2=0
cc_150 N_A2_M1005_g N_A3_c_220_n 0.0166563f $X=1.51 $Y=0.69 $X2=0 $Y2=0
cc_151 N_A2_c_149_n N_A1_c_262_n 0.0176963f $X=2.605 $Y=1.86 $X2=0 $Y2=0
cc_152 N_A2_c_151_n N_A1_c_262_n 0.00128926f $X=2.68 $Y=1.61 $X2=0 $Y2=0
cc_153 N_A2_c_149_n N_A1_c_267_n 0.0333879f $X=2.605 $Y=1.86 $X2=0 $Y2=0
cc_154 N_A2_c_165_p N_A1_c_267_n 6.12011e-19 $X=2.515 $Y=2.405 $X2=0 $Y2=0
cc_155 N_A2_c_151_n N_A1_c_267_n 0.00173704f $X=2.68 $Y=1.61 $X2=0 $Y2=0
cc_156 N_A2_c_149_n N_A1_c_263_n 3.52691e-19 $X=2.605 $Y=1.86 $X2=0 $Y2=0
cc_157 N_A2_c_150_n N_A_31_387#_c_308_n 0.0135297f $X=1.72 $Y=2.32 $X2=0 $Y2=0
cc_158 N_A2_c_152_n N_A_31_387#_c_308_n 6.39279e-19 $X=1.6 $Y=1.305 $X2=0 $Y2=0
cc_159 N_A2_c_153_n N_A_31_387#_c_308_n 8.43332e-19 $X=1.72 $Y=1.305 $X2=0 $Y2=0
cc_160 N_A2_c_150_n N_A_31_387#_c_334_n 0.02354f $X=1.72 $Y=2.32 $X2=0 $Y2=0
cc_161 N_A2_c_149_n N_A_31_387#_c_319_n 0.0134116f $X=2.605 $Y=1.86 $X2=0 $Y2=0
cc_162 N_A2_c_165_p N_A_31_387#_c_319_n 0.0413727f $X=2.515 $Y=2.405 $X2=0 $Y2=0
cc_163 N_A2_c_195_p N_A_31_387#_c_319_n 0.0072142f $X=1.805 $Y=2.405 $X2=0 $Y2=0
cc_164 N_A2_c_149_n N_A_31_387#_c_320_n 0.00698595f $X=2.605 $Y=1.86 $X2=0 $Y2=0
cc_165 N_A2_c_165_p N_A_31_387#_c_320_n 0.0138308f $X=2.515 $Y=2.405 $X2=0 $Y2=0
cc_166 N_A2_c_151_n N_A_31_387#_c_320_n 0.0408386f $X=2.68 $Y=1.61 $X2=0 $Y2=0
cc_167 N_A2_c_149_n N_A_31_387#_c_311_n 0.00103439f $X=2.605 $Y=1.86 $X2=0 $Y2=0
cc_168 N_A2_c_151_n N_A_31_387#_c_311_n 0.0142132f $X=2.68 $Y=1.61 $X2=0 $Y2=0
cc_169 N_A2_c_149_n N_VPWR_c_431_n 0.00399513f $X=2.605 $Y=1.86 $X2=0 $Y2=0
cc_170 N_A2_c_149_n N_VPWR_c_427_n 0.00537853f $X=2.605 $Y=1.86 $X2=0 $Y2=0
cc_171 N_A2_c_150_n A_320_387# 0.0110094f $X=1.72 $Y=2.32 $X2=-0.19 $Y2=-0.245
cc_172 N_A2_c_165_p A_320_387# 0.0262931f $X=2.515 $Y=2.405 $X2=-0.19 $Y2=-0.245
cc_173 N_A2_c_195_p A_320_387# 0.00345505f $X=1.805 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_174 N_A2_c_165_p A_536_387# 0.00302979f $X=2.515 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_175 N_A2_c_151_n A_536_387# 0.00338565f $X=2.68 $Y=1.61 $X2=-0.19 $Y2=-0.245
cc_176 N_A2_M1005_g N_A_209_74#_c_504_n 0.0203628f $X=1.51 $Y=0.69 $X2=0 $Y2=0
cc_177 N_A2_c_153_n N_A_209_74#_c_504_n 0.00310605f $X=1.72 $Y=1.305 $X2=0 $Y2=0
cc_178 N_A2_M1005_g N_VGND_c_531_n 0.0056177f $X=1.51 $Y=0.69 $X2=0 $Y2=0
cc_179 N_A2_c_149_n N_VGND_c_531_n 0.0017834f $X=2.605 $Y=1.86 $X2=0 $Y2=0
cc_180 N_A2_c_151_n N_VGND_c_531_n 0.0111729f $X=2.68 $Y=1.61 $X2=0 $Y2=0
cc_181 N_A2_c_152_n N_VGND_c_531_n 0.00385043f $X=1.6 $Y=1.305 $X2=0 $Y2=0
cc_182 N_A2_c_153_n N_VGND_c_531_n 0.0148018f $X=1.72 $Y=1.305 $X2=0 $Y2=0
cc_183 N_A2_M1005_g N_VGND_c_523_n 0.00281891f $X=1.51 $Y=0.69 $X2=0 $Y2=0
cc_184 N_A2_M1005_g N_VGND_c_525_n 0.00357277f $X=1.51 $Y=0.69 $X2=0 $Y2=0
cc_185 N_A3_c_223_n N_A_31_387#_c_308_n 0.00301767f $X=1.6 $Y=1.785 $X2=0 $Y2=0
cc_186 N_A3_c_221_n N_A_31_387#_c_318_n 6.07096e-19 $X=1.525 $Y=1.86 $X2=0 $Y2=0
cc_187 N_A3_c_221_n N_A_31_387#_c_334_n 0.0196746f $X=1.525 $Y=1.86 $X2=0 $Y2=0
cc_188 N_A3_c_223_n N_A_31_387#_c_334_n 0.00175313f $X=1.6 $Y=1.785 $X2=0 $Y2=0
cc_189 N_A3_c_221_n N_A_31_387#_c_319_n 0.0135012f $X=1.525 $Y=1.86 $X2=0 $Y2=0
cc_190 N_A3_c_221_n N_VPWR_c_431_n 0.00399501f $X=1.525 $Y=1.86 $X2=0 $Y2=0
cc_191 N_A3_c_221_n N_VPWR_c_427_n 0.00537853f $X=1.525 $Y=1.86 $X2=0 $Y2=0
cc_192 A3 A_320_387# 0.00965894f $X=2.075 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_193 N_A3_c_220_n N_A_209_74#_c_504_n 0.0159594f $X=2.14 $Y=1.085 $X2=0 $Y2=0
cc_194 A3 N_VGND_c_531_n 0.0233403f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_195 N_A3_c_219_n N_VGND_c_531_n 0.00471366f $X=2.14 $Y=1.285 $X2=0 $Y2=0
cc_196 N_A3_c_220_n N_VGND_c_531_n 0.0136627f $X=2.14 $Y=1.085 $X2=0 $Y2=0
cc_197 N_A3_c_220_n N_VGND_c_523_n 0.00281891f $X=2.14 $Y=1.085 $X2=0 $Y2=0
cc_198 N_A3_c_220_n N_VGND_c_525_n 0.00361247f $X=2.14 $Y=1.085 $X2=0 $Y2=0
cc_199 N_A1_c_262_n N_A_31_387#_c_304_n 0.0136207f $X=3.175 $Y=1.77 $X2=0 $Y2=0
cc_200 N_A1_c_267_n N_A_31_387#_c_304_n 0.0202664f $X=3.175 $Y=1.86 $X2=0 $Y2=0
cc_201 N_A1_c_263_n N_A_31_387#_c_304_n 0.0063017f $X=3.22 $Y=1.285 $X2=0 $Y2=0
cc_202 N_A1_c_264_n N_A_31_387#_c_304_n 3.45132e-19 $X=3.22 $Y=1.285 $X2=0 $Y2=0
cc_203 N_A1_c_264_n N_A_31_387#_M1004_g 0.00133094f $X=3.22 $Y=1.285 $X2=0 $Y2=0
cc_204 N_A1_c_265_n N_A_31_387#_M1004_g 0.022713f $X=3.22 $Y=1.12 $X2=0 $Y2=0
cc_205 N_A1_c_267_n N_A_31_387#_c_319_n 0.00603074f $X=3.175 $Y=1.86 $X2=0 $Y2=0
cc_206 N_A1_c_267_n N_A_31_387#_c_320_n 0.0248218f $X=3.175 $Y=1.86 $X2=0 $Y2=0
cc_207 N_A1_c_262_n N_A_31_387#_c_310_n 0.00416531f $X=3.175 $Y=1.77 $X2=0 $Y2=0
cc_208 N_A1_c_267_n N_A_31_387#_c_310_n 0.00380473f $X=3.175 $Y=1.86 $X2=0 $Y2=0
cc_209 N_A1_c_263_n N_A_31_387#_c_310_n 0.00316326f $X=3.22 $Y=1.285 $X2=0 $Y2=0
cc_210 N_A1_c_264_n N_A_31_387#_c_310_n 0.0146979f $X=3.22 $Y=1.285 $X2=0 $Y2=0
cc_211 N_A1_c_262_n N_A_31_387#_c_311_n 0.00348446f $X=3.175 $Y=1.77 $X2=0 $Y2=0
cc_212 N_A1_c_267_n N_A_31_387#_c_311_n 3.22226e-19 $X=3.175 $Y=1.86 $X2=0 $Y2=0
cc_213 N_A1_c_263_n N_A_31_387#_c_311_n 6.9887e-19 $X=3.22 $Y=1.285 $X2=0 $Y2=0
cc_214 N_A1_c_264_n N_A_31_387#_c_311_n 0.0140509f $X=3.22 $Y=1.285 $X2=0 $Y2=0
cc_215 N_A1_c_262_n N_A_31_387#_c_313_n 0.00118121f $X=3.175 $Y=1.77 $X2=0 $Y2=0
cc_216 N_A1_c_264_n N_A_31_387#_c_313_n 0.00631056f $X=3.22 $Y=1.285 $X2=0 $Y2=0
cc_217 N_A1_c_267_n N_VPWR_c_429_n 0.0118174f $X=3.175 $Y=1.86 $X2=0 $Y2=0
cc_218 N_A1_c_267_n N_VPWR_c_431_n 0.00468858f $X=3.175 $Y=1.86 $X2=0 $Y2=0
cc_219 N_A1_c_267_n N_VPWR_c_427_n 0.00537853f $X=3.175 $Y=1.86 $X2=0 $Y2=0
cc_220 N_A1_c_264_n X 2.93139e-19 $X=3.22 $Y=1.285 $X2=0 $Y2=0
cc_221 N_A1_c_265_n X 6.59557e-19 $X=3.22 $Y=1.12 $X2=0 $Y2=0
cc_222 N_A1_c_265_n N_A_209_74#_c_504_n 0.00664776f $X=3.22 $Y=1.12 $X2=0 $Y2=0
cc_223 N_A1_c_263_n N_VGND_c_531_n 0.00450164f $X=3.22 $Y=1.285 $X2=0 $Y2=0
cc_224 N_A1_c_264_n N_VGND_c_531_n 0.0251429f $X=3.22 $Y=1.285 $X2=0 $Y2=0
cc_225 N_A1_c_265_n N_VGND_c_531_n 0.0111167f $X=3.22 $Y=1.12 $X2=0 $Y2=0
cc_226 N_A1_c_265_n N_VGND_c_522_n 0.0146844f $X=3.22 $Y=1.12 $X2=0 $Y2=0
cc_227 N_A1_c_265_n N_VGND_c_523_n 0.00383152f $X=3.22 $Y=1.12 $X2=0 $Y2=0
cc_228 N_A1_c_265_n N_VGND_c_525_n 0.00374822f $X=3.22 $Y=1.12 $X2=0 $Y2=0
cc_229 N_A_31_387#_c_315_n N_VPWR_c_428_n 0.0373748f $X=0.3 $Y=2.08 $X2=0 $Y2=0
cc_230 N_A_31_387#_c_309_n N_VPWR_c_428_n 0.0251994f $X=0.75 $Y=1.725 $X2=0
+ $Y2=0
cc_231 N_A_31_387#_c_318_n N_VPWR_c_428_n 0.00795491f $X=1.3 $Y=2.785 $X2=0
+ $Y2=0
cc_232 N_A_31_387#_c_304_n N_VPWR_c_429_n 0.0110742f $X=3.795 $Y=1.765 $X2=0
+ $Y2=0
cc_233 N_A_31_387#_c_319_n N_VPWR_c_429_n 0.0140387f $X=3.015 $Y=2.87 $X2=0
+ $Y2=0
cc_234 N_A_31_387#_c_320_n N_VPWR_c_429_n 0.0610102f $X=3.1 $Y=2.785 $X2=0 $Y2=0
cc_235 N_A_31_387#_c_310_n N_VPWR_c_429_n 0.0197628f $X=3.595 $Y=1.705 $X2=0
+ $Y2=0
cc_236 N_A_31_387#_c_313_n N_VPWR_c_429_n 0.00688187f $X=3.76 $Y=1.515 $X2=0
+ $Y2=0
cc_237 N_A_31_387#_c_315_n N_VPWR_c_430_n 0.0132586f $X=0.3 $Y=2.08 $X2=0 $Y2=0
cc_238 N_A_31_387#_c_318_n N_VPWR_c_431_n 0.0132602f $X=1.3 $Y=2.785 $X2=0 $Y2=0
cc_239 N_A_31_387#_c_319_n N_VPWR_c_431_n 0.0628064f $X=3.015 $Y=2.87 $X2=0
+ $Y2=0
cc_240 N_A_31_387#_c_304_n N_VPWR_c_432_n 0.00445602f $X=3.795 $Y=1.765 $X2=0
+ $Y2=0
cc_241 N_A_31_387#_c_304_n N_VPWR_c_427_n 0.00865278f $X=3.795 $Y=1.765 $X2=0
+ $Y2=0
cc_242 N_A_31_387#_c_315_n N_VPWR_c_427_n 0.0119178f $X=0.3 $Y=2.08 $X2=0 $Y2=0
cc_243 N_A_31_387#_c_318_n N_VPWR_c_427_n 0.0119651f $X=1.3 $Y=2.785 $X2=0 $Y2=0
cc_244 N_A_31_387#_c_319_n N_VPWR_c_427_n 0.0597297f $X=3.015 $Y=2.87 $X2=0
+ $Y2=0
cc_245 N_A_31_387#_c_319_n A_320_387# 0.0158797f $X=3.015 $Y=2.87 $X2=-0.19
+ $Y2=-0.245
cc_246 N_A_31_387#_c_319_n A_536_387# 0.00840874f $X=3.015 $Y=2.87 $X2=-0.19
+ $Y2=-0.245
cc_247 N_A_31_387#_c_320_n A_536_387# 0.00884873f $X=3.1 $Y=2.785 $X2=-0.19
+ $Y2=-0.245
cc_248 N_A_31_387#_c_304_n N_X_c_480_n 0.0085677f $X=3.795 $Y=1.765 $X2=0 $Y2=0
cc_249 N_A_31_387#_c_304_n N_X_c_481_n 0.00202785f $X=3.795 $Y=1.765 $X2=0 $Y2=0
cc_250 N_A_31_387#_c_313_n N_X_c_481_n 0.00215794f $X=3.76 $Y=1.515 $X2=0 $Y2=0
cc_251 N_A_31_387#_c_304_n N_X_c_477_n 0.0124144f $X=3.795 $Y=1.765 $X2=0 $Y2=0
cc_252 N_A_31_387#_M1004_g N_X_c_477_n 0.00580334f $X=3.82 $Y=0.74 $X2=0 $Y2=0
cc_253 N_A_31_387#_c_313_n N_X_c_477_n 0.0332755f $X=3.76 $Y=1.515 $X2=0 $Y2=0
cc_254 N_A_31_387#_M1004_g X 0.00812529f $X=3.82 $Y=0.74 $X2=0 $Y2=0
cc_255 N_A_31_387#_c_304_n X 0.0012634f $X=3.795 $Y=1.765 $X2=0 $Y2=0
cc_256 N_A_31_387#_M1004_g X 0.0042952f $X=3.82 $Y=0.74 $X2=0 $Y2=0
cc_257 N_A_31_387#_c_313_n X 0.00153012f $X=3.76 $Y=1.515 $X2=0 $Y2=0
cc_258 N_A_31_387#_c_307_n A_131_74# 5.66122e-19 $X=0.665 $Y=1.64 $X2=-0.19
+ $Y2=-0.245
cc_259 N_A_31_387#_c_312_n A_131_74# 0.00269364f $X=0.665 $Y=0.885 $X2=-0.19
+ $Y2=-0.245
cc_260 N_A_31_387#_c_306_n N_A_209_74#_c_503_n 0.00424699f $X=0.365 $Y=0.515
+ $X2=0 $Y2=0
cc_261 N_A_31_387#_c_308_n N_A_209_74#_c_506_n 0.00334383f $X=1.135 $Y=1.725
+ $X2=0 $Y2=0
cc_262 N_A_31_387#_c_304_n N_VGND_c_531_n 6.53733e-19 $X=3.795 $Y=1.765 $X2=0
+ $Y2=0
cc_263 N_A_31_387#_c_310_n N_VGND_c_531_n 0.00547315f $X=3.595 $Y=1.705 $X2=0
+ $Y2=0
cc_264 N_A_31_387#_c_313_n N_VGND_c_531_n 0.00405649f $X=3.76 $Y=1.515 $X2=0
+ $Y2=0
cc_265 N_A_31_387#_M1004_g N_VGND_c_522_n 0.00538108f $X=3.82 $Y=0.74 $X2=0
+ $Y2=0
cc_266 N_A_31_387#_c_306_n N_VGND_c_523_n 0.0141395f $X=0.365 $Y=0.515 $X2=0
+ $Y2=0
cc_267 N_A_31_387#_M1004_g N_VGND_c_524_n 0.00434272f $X=3.82 $Y=0.74 $X2=0
+ $Y2=0
cc_268 N_A_31_387#_M1004_g N_VGND_c_525_n 0.00824752f $X=3.82 $Y=0.74 $X2=0
+ $Y2=0
cc_269 N_A_31_387#_c_306_n N_VGND_c_525_n 0.0118342f $X=0.365 $Y=0.515 $X2=0
+ $Y2=0
cc_270 N_A_31_387#_c_312_n N_VGND_c_525_n 0.00703783f $X=0.665 $Y=0.885 $X2=0
+ $Y2=0
cc_271 N_VPWR_c_432_n N_X_c_480_n 0.0168249f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_272 N_VPWR_c_427_n N_X_c_480_n 0.0138933f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_273 N_VPWR_c_429_n N_X_c_481_n 0.0398603f $X=3.52 $Y=2.125 $X2=0 $Y2=0
cc_274 X N_VGND_c_522_n 0.0164106f $X=3.995 $Y=0.47 $X2=0 $Y2=0
cc_275 X N_VGND_c_524_n 0.0161257f $X=3.995 $Y=0.47 $X2=0 $Y2=0
cc_276 X N_VGND_c_525_n 0.013291f $X=3.995 $Y=0.47 $X2=0 $Y2=0
cc_277 N_A_209_74#_c_504_n N_VGND_M1005_d 0.00743158f $X=3.015 $Y=0.525
+ $X2=-0.19 $Y2=-0.245
cc_278 N_A_209_74#_M1003_d N_VGND_c_531_n 0.0325693f $X=2.305 $Y=0.37 $X2=0
+ $Y2=0
cc_279 N_A_209_74#_c_504_n N_VGND_c_531_n 0.106422f $X=3.015 $Y=0.525 $X2=0
+ $Y2=0
cc_280 N_A_209_74#_c_504_n N_VGND_c_522_n 0.0157478f $X=3.015 $Y=0.525 $X2=0
+ $Y2=0
cc_281 N_A_209_74#_c_503_n N_VGND_c_523_n 0.0204446f $X=1.225 $Y=0.61 $X2=0
+ $Y2=0
cc_282 N_A_209_74#_c_504_n N_VGND_c_523_n 0.103511f $X=3.015 $Y=0.525 $X2=0
+ $Y2=0
cc_283 N_A_209_74#_c_503_n N_VGND_c_525_n 0.0126791f $X=1.225 $Y=0.61 $X2=0
+ $Y2=0
cc_284 N_A_209_74#_c_504_n N_VGND_c_525_n 0.0659666f $X=3.015 $Y=0.525 $X2=0
+ $Y2=0
