* File: sky130_fd_sc_ls__einvn_8.pxi.spice
* Created: Wed Sep  2 11:06:57 2020
* 
x_PM_SKY130_FD_SC_LS__EINVN_8%A_126_74# N_A_126_74#_M1032_d N_A_126_74#_M1020_d
+ N_A_126_74#_c_173_n N_A_126_74#_c_174_n N_A_126_74#_c_175_n
+ N_A_126_74#_M1003_g N_A_126_74#_c_176_n N_A_126_74#_c_177_n
+ N_A_126_74#_M1005_g N_A_126_74#_c_178_n N_A_126_74#_c_179_n
+ N_A_126_74#_M1015_g N_A_126_74#_c_180_n N_A_126_74#_c_181_n
+ N_A_126_74#_M1016_g N_A_126_74#_c_182_n N_A_126_74#_c_183_n
+ N_A_126_74#_M1019_g N_A_126_74#_c_184_n N_A_126_74#_c_185_n
+ N_A_126_74#_M1026_g N_A_126_74#_c_186_n N_A_126_74#_c_187_n
+ N_A_126_74#_M1030_g N_A_126_74#_c_188_n N_A_126_74#_c_189_n
+ N_A_126_74#_M1033_g N_A_126_74#_c_190_n N_A_126_74#_c_191_n
+ N_A_126_74#_c_192_n N_A_126_74#_c_193_n N_A_126_74#_c_194_n
+ N_A_126_74#_c_195_n N_A_126_74#_c_196_n N_A_126_74#_c_197_n
+ N_A_126_74#_c_198_n N_A_126_74#_c_199_n N_A_126_74#_c_200_n
+ PM_SKY130_FD_SC_LS__EINVN_8%A_126_74#
x_PM_SKY130_FD_SC_LS__EINVN_8%TE_B N_TE_B_M1032_g N_TE_B_c_326_n N_TE_B_M1020_g
+ N_TE_B_c_327_n N_TE_B_c_345_n N_TE_B_M1000_g N_TE_B_c_328_n N_TE_B_c_347_n
+ N_TE_B_M1002_g N_TE_B_c_329_n N_TE_B_c_349_n N_TE_B_M1008_g N_TE_B_c_330_n
+ N_TE_B_c_351_n N_TE_B_M1012_g N_TE_B_c_331_n N_TE_B_c_353_n N_TE_B_M1018_g
+ N_TE_B_c_332_n N_TE_B_c_355_n N_TE_B_M1023_g N_TE_B_c_333_n N_TE_B_c_357_n
+ N_TE_B_M1027_g N_TE_B_c_334_n N_TE_B_c_359_n N_TE_B_M1031_g N_TE_B_c_335_n
+ N_TE_B_c_336_n N_TE_B_c_337_n N_TE_B_c_338_n N_TE_B_c_339_n N_TE_B_c_340_n
+ N_TE_B_c_341_n TE_B PM_SKY130_FD_SC_LS__EINVN_8%TE_B
x_PM_SKY130_FD_SC_LS__EINVN_8%A N_A_M1004_g N_A_c_503_n N_A_M1001_g N_A_M1007_g
+ N_A_c_504_n N_A_M1006_g N_A_M1010_g N_A_c_505_n N_A_M1009_g N_A_M1013_g
+ N_A_c_506_n N_A_M1011_g N_A_M1017_g N_A_c_507_n N_A_M1014_g N_A_M1022_g
+ N_A_c_508_n N_A_M1021_g N_A_M1024_g N_A_c_509_n N_A_M1025_g N_A_c_510_n
+ N_A_M1028_g N_A_M1029_g A A A A A N_A_c_502_n PM_SKY130_FD_SC_LS__EINVN_8%A
x_PM_SKY130_FD_SC_LS__EINVN_8%VPWR N_VPWR_M1020_s N_VPWR_M1000_d N_VPWR_M1008_d
+ N_VPWR_M1018_d N_VPWR_M1027_d N_VPWR_c_653_n N_VPWR_c_654_n N_VPWR_c_655_n
+ N_VPWR_c_656_n N_VPWR_c_657_n N_VPWR_c_658_n N_VPWR_c_659_n N_VPWR_c_660_n
+ N_VPWR_c_661_n VPWR N_VPWR_c_662_n N_VPWR_c_663_n N_VPWR_c_652_n
+ N_VPWR_c_665_n N_VPWR_c_666_n N_VPWR_c_667_n N_VPWR_c_668_n
+ PM_SKY130_FD_SC_LS__EINVN_8%VPWR
x_PM_SKY130_FD_SC_LS__EINVN_8%A_239_368# N_A_239_368#_M1000_s
+ N_A_239_368#_M1002_s N_A_239_368#_M1012_s N_A_239_368#_M1023_s
+ N_A_239_368#_M1031_s N_A_239_368#_M1006_s N_A_239_368#_M1011_s
+ N_A_239_368#_M1021_s N_A_239_368#_M1028_s N_A_239_368#_c_758_n
+ N_A_239_368#_c_759_n N_A_239_368#_c_760_n N_A_239_368#_c_761_n
+ N_A_239_368#_c_762_n N_A_239_368#_c_763_n N_A_239_368#_c_764_n
+ N_A_239_368#_c_765_n N_A_239_368#_c_817_n N_A_239_368#_c_819_n
+ N_A_239_368#_c_820_n N_A_239_368#_c_766_n N_A_239_368#_c_767_n
+ N_A_239_368#_c_842_n N_A_239_368#_c_768_n N_A_239_368#_c_902_p
+ N_A_239_368#_c_769_n N_A_239_368#_c_906_p N_A_239_368#_c_770_n
+ N_A_239_368#_c_771_n N_A_239_368#_c_783_n N_A_239_368#_c_784_n
+ N_A_239_368#_c_772_n N_A_239_368#_c_773_n N_A_239_368#_c_774_n
+ N_A_239_368#_c_775_n PM_SKY130_FD_SC_LS__EINVN_8%A_239_368#
x_PM_SKY130_FD_SC_LS__EINVN_8%Z N_Z_M1004_d N_Z_M1010_d N_Z_M1017_d N_Z_M1024_d
+ N_Z_M1001_d N_Z_M1009_d N_Z_M1014_d N_Z_M1025_d N_Z_c_944_n N_Z_c_931_n
+ N_Z_c_938_n N_Z_c_951_n N_Z_c_953_n N_Z_c_957_n N_Z_c_932_n N_Z_c_962_n
+ N_Z_c_1044_p N_Z_c_933_n N_Z_c_971_n N_Z_c_1049_p N_Z_c_934_n N_Z_c_940_n
+ N_Z_c_1023_n N_Z_c_935_n N_Z_c_936_n N_Z_c_989_n N_Z_c_937_n N_Z_c_994_n
+ N_Z_c_1000_n Z PM_SKY130_FD_SC_LS__EINVN_8%Z
x_PM_SKY130_FD_SC_LS__EINVN_8%VGND N_VGND_M1032_s N_VGND_M1003_d N_VGND_M1015_d
+ N_VGND_M1019_d N_VGND_M1030_d N_VGND_c_1052_n N_VGND_c_1053_n N_VGND_c_1054_n
+ N_VGND_c_1055_n N_VGND_c_1056_n N_VGND_c_1057_n N_VGND_c_1058_n
+ N_VGND_c_1059_n N_VGND_c_1060_n N_VGND_c_1061_n N_VGND_c_1062_n
+ N_VGND_c_1063_n N_VGND_c_1064_n N_VGND_c_1065_n VGND N_VGND_c_1066_n
+ N_VGND_c_1067_n PM_SKY130_FD_SC_LS__EINVN_8%VGND
x_PM_SKY130_FD_SC_LS__EINVN_8%A_293_74# N_A_293_74#_M1003_s N_A_293_74#_M1005_s
+ N_A_293_74#_M1016_s N_A_293_74#_M1026_s N_A_293_74#_M1033_s
+ N_A_293_74#_M1007_s N_A_293_74#_M1013_s N_A_293_74#_M1022_s
+ N_A_293_74#_M1029_s N_A_293_74#_c_1160_n N_A_293_74#_c_1161_n
+ N_A_293_74#_c_1162_n N_A_293_74#_c_1163_n N_A_293_74#_c_1164_n
+ N_A_293_74#_c_1165_n N_A_293_74#_c_1166_n N_A_293_74#_c_1167_n
+ N_A_293_74#_c_1168_n N_A_293_74#_c_1169_n N_A_293_74#_c_1170_n
+ N_A_293_74#_c_1171_n N_A_293_74#_c_1172_n N_A_293_74#_c_1243_n
+ N_A_293_74#_c_1173_n N_A_293_74#_c_1174_n N_A_293_74#_c_1175_n
+ N_A_293_74#_c_1176_n N_A_293_74#_c_1177_n N_A_293_74#_c_1178_n
+ N_A_293_74#_c_1179_n PM_SKY130_FD_SC_LS__EINVN_8%A_293_74#
cc_1 VNB N_A_126_74#_c_173_n 0.0195256f $X=-0.19 $Y=-0.245 $X2=1.75 $Y2=1.26
cc_2 VNB N_A_126_74#_c_174_n 0.0116503f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=1.26
cc_3 VNB N_A_126_74#_c_175_n 0.0175595f $X=-0.19 $Y=-0.245 $X2=1.825 $Y2=1.185
cc_4 VNB N_A_126_74#_c_176_n 0.009775f $X=-0.19 $Y=-0.245 $X2=2.18 $Y2=1.26
cc_5 VNB N_A_126_74#_c_177_n 0.0149561f $X=-0.19 $Y=-0.245 $X2=2.255 $Y2=1.185
cc_6 VNB N_A_126_74#_c_178_n 0.0105004f $X=-0.19 $Y=-0.245 $X2=2.61 $Y2=1.26
cc_7 VNB N_A_126_74#_c_179_n 0.0151386f $X=-0.19 $Y=-0.245 $X2=2.685 $Y2=1.185
cc_8 VNB N_A_126_74#_c_180_n 0.013192f $X=-0.19 $Y=-0.245 $X2=3.11 $Y2=1.26
cc_9 VNB N_A_126_74#_c_181_n 0.0154922f $X=-0.19 $Y=-0.245 $X2=3.185 $Y2=1.185
cc_10 VNB N_A_126_74#_c_182_n 0.0105004f $X=-0.19 $Y=-0.245 $X2=3.54 $Y2=1.26
cc_11 VNB N_A_126_74#_c_183_n 0.0151383f $X=-0.19 $Y=-0.245 $X2=3.615 $Y2=1.185
cc_12 VNB N_A_126_74#_c_184_n 0.0131804f $X=-0.19 $Y=-0.245 $X2=4.04 $Y2=1.26
cc_13 VNB N_A_126_74#_c_185_n 0.0154922f $X=-0.19 $Y=-0.245 $X2=4.115 $Y2=1.185
cc_14 VNB N_A_126_74#_c_186_n 0.0105004f $X=-0.19 $Y=-0.245 $X2=4.47 $Y2=1.26
cc_15 VNB N_A_126_74#_c_187_n 0.0146944f $X=-0.19 $Y=-0.245 $X2=4.545 $Y2=1.185
cc_16 VNB N_A_126_74#_c_188_n 0.016112f $X=-0.19 $Y=-0.245 $X2=4.9 $Y2=1.26
cc_17 VNB N_A_126_74#_c_189_n 0.0150038f $X=-0.19 $Y=-0.245 $X2=4.975 $Y2=1.185
cc_18 VNB N_A_126_74#_c_190_n 0.00412378f $X=-0.19 $Y=-0.245 $X2=1.825 $Y2=1.26
cc_19 VNB N_A_126_74#_c_191_n 0.00411221f $X=-0.19 $Y=-0.245 $X2=2.255 $Y2=1.26
cc_20 VNB N_A_126_74#_c_192_n 0.00412378f $X=-0.19 $Y=-0.245 $X2=2.685 $Y2=1.26
cc_21 VNB N_A_126_74#_c_193_n 0.00411221f $X=-0.19 $Y=-0.245 $X2=3.185 $Y2=1.26
cc_22 VNB N_A_126_74#_c_194_n 0.00412378f $X=-0.19 $Y=-0.245 $X2=3.615 $Y2=1.26
cc_23 VNB N_A_126_74#_c_195_n 0.00411221f $X=-0.19 $Y=-0.245 $X2=4.115 $Y2=1.26
cc_24 VNB N_A_126_74#_c_196_n 0.00411221f $X=-0.19 $Y=-0.245 $X2=4.545 $Y2=1.26
cc_25 VNB N_A_126_74#_c_197_n 0.00607853f $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=1.985
cc_26 VNB N_A_126_74#_c_198_n 0.00623379f $X=-0.19 $Y=-0.245 $X2=1.19 $Y2=0.49
cc_27 VNB N_A_126_74#_c_199_n 0.0727067f $X=-0.19 $Y=-0.245 $X2=1.19 $Y2=0.49
cc_28 VNB N_A_126_74#_c_200_n 0.00657985f $X=-0.19 $Y=-0.245 $X2=1.19 $Y2=1.17
cc_29 VNB N_TE_B_M1032_g 0.0278801f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_TE_B_c_326_n 0.0585644f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_TE_B_c_327_n 0.0257209f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=1.26
cc_32 VNB N_TE_B_c_328_n 0.00838936f $X=-0.19 $Y=-0.245 $X2=1.9 $Y2=1.26
cc_33 VNB N_TE_B_c_329_n 0.00707023f $X=-0.19 $Y=-0.245 $X2=2.33 $Y2=1.26
cc_34 VNB N_TE_B_c_330_n 0.00838938f $X=-0.19 $Y=-0.245 $X2=2.76 $Y2=1.26
cc_35 VNB N_TE_B_c_331_n 0.00707022f $X=-0.19 $Y=-0.245 $X2=3.26 $Y2=1.26
cc_36 VNB N_TE_B_c_332_n 0.00838938f $X=-0.19 $Y=-0.245 $X2=3.69 $Y2=1.26
cc_37 VNB N_TE_B_c_333_n 0.00707021f $X=-0.19 $Y=-0.245 $X2=4.19 $Y2=1.26
cc_38 VNB N_TE_B_c_334_n 0.014922f $X=-0.19 $Y=-0.245 $X2=4.62 $Y2=1.26
cc_39 VNB N_TE_B_c_335_n 0.004883f $X=-0.19 $Y=-0.245 $X2=1.825 $Y2=1.26
cc_40 VNB N_TE_B_c_336_n 0.0048708f $X=-0.19 $Y=-0.245 $X2=2.255 $Y2=1.26
cc_41 VNB N_TE_B_c_337_n 0.00487072f $X=-0.19 $Y=-0.245 $X2=2.685 $Y2=1.26
cc_42 VNB N_TE_B_c_338_n 0.0048708f $X=-0.19 $Y=-0.245 $X2=3.185 $Y2=1.26
cc_43 VNB N_TE_B_c_339_n 0.00487074f $X=-0.19 $Y=-0.245 $X2=3.615 $Y2=1.26
cc_44 VNB N_TE_B_c_340_n 0.0048708f $X=-0.19 $Y=-0.245 $X2=4.115 $Y2=1.26
cc_45 VNB N_TE_B_c_341_n 0.00487632f $X=-0.19 $Y=-0.245 $X2=4.545 $Y2=1.26
cc_46 VNB TE_B 0.0103923f $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=1.335
cc_47 VNB N_A_M1004_g 0.0221898f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_M1007_g 0.0225221f $X=-0.19 $Y=-0.245 $X2=1.825 $Y2=0.74
cc_49 VNB N_A_M1010_g 0.0223938f $X=-0.19 $Y=-0.245 $X2=2.61 $Y2=1.26
cc_50 VNB N_A_M1013_g 0.023211f $X=-0.19 $Y=-0.245 $X2=3.185 $Y2=1.185
cc_51 VNB N_A_M1017_g 0.0231908f $X=-0.19 $Y=-0.245 $X2=3.615 $Y2=0.74
cc_52 VNB N_A_M1022_g 0.0222089f $X=-0.19 $Y=-0.245 $X2=4.19 $Y2=1.26
cc_53 VNB N_A_M1024_g 0.0240746f $X=-0.19 $Y=-0.245 $X2=4.975 $Y2=0.74
cc_54 VNB N_A_M1029_g 0.0335013f $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=1.335
cc_55 VNB A 0.0168057f $X=-0.19 $Y=-0.245 $X2=1.02 $Y2=1.13
cc_56 VNB N_A_c_502_n 0.155021f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_VPWR_c_652_n 0.382608f $X=-0.19 $Y=-0.245 $X2=1.19 $Y2=0.49
cc_58 VNB N_Z_c_931_n 0.00202243f $X=-0.19 $Y=-0.245 $X2=3.185 $Y2=0.74
cc_59 VNB N_Z_c_932_n 0.00317099f $X=-0.19 $Y=-0.245 $X2=4.545 $Y2=0.74
cc_60 VNB N_Z_c_933_n 0.00651605f $X=-0.19 $Y=-0.245 $X2=3.185 $Y2=1.26
cc_61 VNB N_Z_c_934_n 0.0056064f $X=-0.19 $Y=-0.245 $X2=1.19 $Y2=0.49
cc_62 VNB N_Z_c_935_n 0.00612864f $X=-0.19 $Y=-0.245 $X2=1.19 $Y2=1.17
cc_63 VNB N_Z_c_936_n 0.00228886f $X=-0.19 $Y=-0.245 $X2=1.19 $Y2=1.17
cc_64 VNB N_Z_c_937_n 0.00124857f $X=-0.19 $Y=-0.245 $X2=1.19 $Y2=0.49
cc_65 VNB N_VGND_c_1052_n 0.0139411f $X=-0.19 $Y=-0.245 $X2=2.255 $Y2=0.74
cc_66 VNB N_VGND_c_1053_n 0.0336621f $X=-0.19 $Y=-0.245 $X2=2.33 $Y2=1.26
cc_67 VNB N_VGND_c_1054_n 0.00642423f $X=-0.19 $Y=-0.245 $X2=3.11 $Y2=1.26
cc_68 VNB N_VGND_c_1055_n 0.00707795f $X=-0.19 $Y=-0.245 $X2=3.185 $Y2=0.74
cc_69 VNB N_VGND_c_1056_n 0.00706502f $X=-0.19 $Y=-0.245 $X2=3.615 $Y2=0.74
cc_70 VNB N_VGND_c_1057_n 0.00333063f $X=-0.19 $Y=-0.245 $X2=4.115 $Y2=1.185
cc_71 VNB N_VGND_c_1058_n 0.0364238f $X=-0.19 $Y=-0.245 $X2=4.47 $Y2=1.26
cc_72 VNB N_VGND_c_1059_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=4.19 $Y2=1.26
cc_73 VNB N_VGND_c_1060_n 0.0172524f $X=-0.19 $Y=-0.245 $X2=4.545 $Y2=0.74
cc_74 VNB N_VGND_c_1061_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=4.545 $Y2=0.74
cc_75 VNB N_VGND_c_1062_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=4.62 $Y2=1.26
cc_76 VNB N_VGND_c_1063_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=4.975 $Y2=1.185
cc_77 VNB N_VGND_c_1064_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=4.975 $Y2=0.74
cc_78 VNB N_VGND_c_1065_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=1.19 $Y2=1.185
cc_79 VNB N_VGND_c_1066_n 0.0976923f $X=-0.19 $Y=-0.245 $X2=1.19 $Y2=1.17
cc_80 VNB N_VGND_c_1067_n 0.488671f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=1.13
cc_81 VNB N_A_293_74#_c_1160_n 0.00280512f $X=-0.19 $Y=-0.245 $X2=3.615 $Y2=0.74
cc_82 VNB N_A_293_74#_c_1161_n 0.00371275f $X=-0.19 $Y=-0.245 $X2=4.04 $Y2=1.26
cc_83 VNB N_A_293_74#_c_1162_n 0.00323505f $X=-0.19 $Y=-0.245 $X2=3.69 $Y2=1.26
cc_84 VNB N_A_293_74#_c_1163_n 0.00270303f $X=-0.19 $Y=-0.245 $X2=4.115 $Y2=0.74
cc_85 VNB N_A_293_74#_c_1164_n 0.0041406f $X=-0.19 $Y=-0.245 $X2=4.19 $Y2=1.26
cc_86 VNB N_A_293_74#_c_1165_n 0.00270303f $X=-0.19 $Y=-0.245 $X2=4.9 $Y2=1.26
cc_87 VNB N_A_293_74#_c_1166_n 0.0041347f $X=-0.19 $Y=-0.245 $X2=4.975 $Y2=1.185
cc_88 VNB N_A_293_74#_c_1167_n 0.00277134f $X=-0.19 $Y=-0.245 $X2=1.825 $Y2=1.26
cc_89 VNB N_A_293_74#_c_1168_n 0.0105983f $X=-0.19 $Y=-0.245 $X2=2.685 $Y2=1.26
cc_90 VNB N_A_293_74#_c_1169_n 0.00211517f $X=-0.19 $Y=-0.245 $X2=3.615 $Y2=1.26
cc_91 VNB N_A_293_74#_c_1170_n 0.00162202f $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=1.335
cc_92 VNB N_A_293_74#_c_1171_n 0.00700214f $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=1.985
cc_93 VNB N_A_293_74#_c_1172_n 0.00199363f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_293_74#_c_1173_n 0.0129598f $X=-0.19 $Y=-0.245 $X2=1.02 $Y2=0.515
cc_95 VNB N_A_293_74#_c_1174_n 0.0301984f $X=-0.19 $Y=-0.245 $X2=1.19 $Y2=1.17
cc_96 VNB N_A_293_74#_c_1175_n 0.0015613f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=1.335
cc_97 VNB N_A_293_74#_c_1176_n 0.0015611f $X=-0.19 $Y=-0.245 $X2=1.19 $Y2=0.49
cc_98 VNB N_A_293_74#_c_1177_n 0.00522494f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_A_293_74#_c_1178_n 0.00241737f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_A_293_74#_c_1179_n 0.00203217f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VPB N_A_126_74#_c_197_n 0.013792f $X=-0.19 $Y=1.66 $X2=0.78 $Y2=1.985
cc_102 VPB N_TE_B_c_326_n 0.0436579f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 VPB N_TE_B_c_327_n 0.0336578f $X=-0.19 $Y=1.66 $X2=1.355 $Y2=1.26
cc_104 VPB N_TE_B_c_345_n 0.0190765f $X=-0.19 $Y=1.66 $X2=1.825 $Y2=0.74
cc_105 VPB N_TE_B_c_328_n 0.011301f $X=-0.19 $Y=1.66 $X2=1.9 $Y2=1.26
cc_106 VPB N_TE_B_c_347_n 0.0153042f $X=-0.19 $Y=1.66 $X2=2.255 $Y2=0.74
cc_107 VPB N_TE_B_c_329_n 0.00949546f $X=-0.19 $Y=1.66 $X2=2.33 $Y2=1.26
cc_108 VPB N_TE_B_c_349_n 0.0148758f $X=-0.19 $Y=1.66 $X2=2.685 $Y2=0.74
cc_109 VPB N_TE_B_c_330_n 0.011301f $X=-0.19 $Y=1.66 $X2=2.76 $Y2=1.26
cc_110 VPB N_TE_B_c_351_n 0.0153042f $X=-0.19 $Y=1.66 $X2=3.185 $Y2=0.74
cc_111 VPB N_TE_B_c_331_n 0.00949546f $X=-0.19 $Y=1.66 $X2=3.26 $Y2=1.26
cc_112 VPB N_TE_B_c_353_n 0.014896f $X=-0.19 $Y=1.66 $X2=3.615 $Y2=0.74
cc_113 VPB N_TE_B_c_332_n 0.011301f $X=-0.19 $Y=1.66 $X2=3.69 $Y2=1.26
cc_114 VPB N_TE_B_c_355_n 0.0153627f $X=-0.19 $Y=1.66 $X2=4.115 $Y2=0.74
cc_115 VPB N_TE_B_c_333_n 0.00952409f $X=-0.19 $Y=1.66 $X2=4.19 $Y2=1.26
cc_116 VPB N_TE_B_c_357_n 0.0156617f $X=-0.19 $Y=1.66 $X2=4.545 $Y2=0.74
cc_117 VPB N_TE_B_c_334_n 0.0159984f $X=-0.19 $Y=1.66 $X2=4.62 $Y2=1.26
cc_118 VPB N_TE_B_c_359_n 0.0159922f $X=-0.19 $Y=1.66 $X2=4.975 $Y2=0.74
cc_119 VPB N_TE_B_c_335_n 0.00460475f $X=-0.19 $Y=1.66 $X2=1.825 $Y2=1.26
cc_120 VPB N_TE_B_c_336_n 0.00397414f $X=-0.19 $Y=1.66 $X2=2.255 $Y2=1.26
cc_121 VPB N_TE_B_c_337_n 0.00397414f $X=-0.19 $Y=1.66 $X2=2.685 $Y2=1.26
cc_122 VPB N_TE_B_c_338_n 0.00397414f $X=-0.19 $Y=1.66 $X2=3.185 $Y2=1.26
cc_123 VPB N_TE_B_c_339_n 0.00397414f $X=-0.19 $Y=1.66 $X2=3.615 $Y2=1.26
cc_124 VPB N_TE_B_c_340_n 0.00397414f $X=-0.19 $Y=1.66 $X2=4.115 $Y2=1.26
cc_125 VPB N_TE_B_c_341_n 0.00401369f $X=-0.19 $Y=1.66 $X2=4.545 $Y2=1.26
cc_126 VPB N_A_c_503_n 0.014745f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_127 VPB N_A_c_504_n 0.0147373f $X=-0.19 $Y=1.66 $X2=2.18 $Y2=1.26
cc_128 VPB N_A_c_505_n 0.0150228f $X=-0.19 $Y=1.66 $X2=2.685 $Y2=1.185
cc_129 VPB N_A_c_506_n 0.0150478f $X=-0.19 $Y=1.66 $X2=3.185 $Y2=0.74
cc_130 VPB N_A_c_507_n 0.014664f $X=-0.19 $Y=1.66 $X2=3.69 $Y2=1.26
cc_131 VPB N_A_c_508_n 0.014664f $X=-0.19 $Y=1.66 $X2=4.545 $Y2=0.74
cc_132 VPB N_A_c_509_n 0.014664f $X=-0.19 $Y=1.66 $X2=1.19 $Y2=1.185
cc_133 VPB N_A_c_510_n 0.0186669f $X=-0.19 $Y=1.66 $X2=2.685 $Y2=1.26
cc_134 VPB A 0.0275176f $X=-0.19 $Y=1.66 $X2=1.02 $Y2=1.13
cc_135 VPB N_A_c_502_n 0.102977f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_VPWR_c_653_n 0.0121909f $X=-0.19 $Y=1.66 $X2=2.255 $Y2=0.74
cc_137 VPB N_VPWR_c_654_n 0.0589698f $X=-0.19 $Y=1.66 $X2=2.33 $Y2=1.26
cc_138 VPB N_VPWR_c_655_n 0.00572483f $X=-0.19 $Y=1.66 $X2=3.185 $Y2=1.185
cc_139 VPB N_VPWR_c_656_n 0.0175706f $X=-0.19 $Y=1.66 $X2=3.26 $Y2=1.26
cc_140 VPB N_VPWR_c_657_n 0.00511574f $X=-0.19 $Y=1.66 $X2=4.04 $Y2=1.26
cc_141 VPB N_VPWR_c_658_n 0.0175706f $X=-0.19 $Y=1.66 $X2=4.115 $Y2=0.74
cc_142 VPB N_VPWR_c_659_n 0.00521035f $X=-0.19 $Y=1.66 $X2=4.545 $Y2=0.74
cc_143 VPB N_VPWR_c_660_n 0.0186948f $X=-0.19 $Y=1.66 $X2=4.975 $Y2=1.185
cc_144 VPB N_VPWR_c_661_n 0.00858913f $X=-0.19 $Y=1.66 $X2=1.825 $Y2=1.26
cc_145 VPB N_VPWR_c_662_n 0.0328287f $X=-0.19 $Y=1.66 $X2=3.615 $Y2=1.26
cc_146 VPB N_VPWR_c_663_n 0.0992334f $X=-0.19 $Y=1.66 $X2=1.02 $Y2=0.49
cc_147 VPB N_VPWR_c_652_n 0.102005f $X=-0.19 $Y=1.66 $X2=1.19 $Y2=0.49
cc_148 VPB N_VPWR_c_665_n 0.00614127f $X=-0.19 $Y=1.66 $X2=1.19 $Y2=1.17
cc_149 VPB N_VPWR_c_666_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0.985 $Y2=1.335
cc_150 VPB N_VPWR_c_667_n 0.00614127f $X=-0.19 $Y=1.66 $X2=1.19 $Y2=1.17
cc_151 VPB N_VPWR_c_668_n 0.00631788f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_152 VPB N_A_239_368#_c_758_n 0.0124897f $X=-0.19 $Y=1.66 $X2=3.615 $Y2=0.74
cc_153 VPB N_A_239_368#_c_759_n 0.0063143f $X=-0.19 $Y=1.66 $X2=4.115 $Y2=1.185
cc_154 VPB N_A_239_368#_c_760_n 9.07775e-19 $X=-0.19 $Y=1.66 $X2=4.115 $Y2=0.74
cc_155 VPB N_A_239_368#_c_761_n 0.00216998f $X=-0.19 $Y=1.66 $X2=4.19 $Y2=1.26
cc_156 VPB N_A_239_368#_c_762_n 0.0063143f $X=-0.19 $Y=1.66 $X2=4.9 $Y2=1.26
cc_157 VPB N_A_239_368#_c_763_n 0.00216998f $X=-0.19 $Y=1.66 $X2=4.975 $Y2=0.74
cc_158 VPB N_A_239_368#_c_764_n 0.0063143f $X=-0.19 $Y=1.66 $X2=2.685 $Y2=1.26
cc_159 VPB N_A_239_368#_c_765_n 0.00257348f $X=-0.19 $Y=1.66 $X2=4.545 $Y2=1.26
cc_160 VPB N_A_239_368#_c_766_n 0.00213603f $X=-0.19 $Y=1.66 $X2=1.02 $Y2=0.49
cc_161 VPB N_A_239_368#_c_767_n 0.0021839f $X=-0.19 $Y=1.66 $X2=1.19 $Y2=0.49
cc_162 VPB N_A_239_368#_c_768_n 0.00294772f $X=-0.19 $Y=1.66 $X2=0.985 $Y2=1.17
cc_163 VPB N_A_239_368#_c_769_n 0.0030474f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_164 VPB N_A_239_368#_c_770_n 0.0124059f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_165 VPB N_A_239_368#_c_771_n 0.0354954f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_166 VPB N_A_239_368#_c_772_n 9.26938e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_167 VPB N_A_239_368#_c_773_n 0.0021839f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_168 VPB N_A_239_368#_c_774_n 0.00123754f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_169 VPB N_A_239_368#_c_775_n 0.00123754f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_170 VPB N_Z_c_938_n 0.00107462f $X=-0.19 $Y=1.66 $X2=3.26 $Y2=1.26
cc_171 VPB N_Z_c_934_n 0.00276498f $X=-0.19 $Y=1.66 $X2=1.19 $Y2=0.49
cc_172 VPB N_Z_c_940_n 0.00332871f $X=-0.19 $Y=1.66 $X2=1.19 $Y2=0.49
cc_173 N_A_126_74#_c_198_n N_TE_B_M1032_g 0.00136832f $X=1.19 $Y=0.49 $X2=0
+ $Y2=0
cc_174 N_A_126_74#_c_199_n N_TE_B_M1032_g 0.0175459f $X=1.19 $Y=0.49 $X2=0 $Y2=0
cc_175 N_A_126_74#_c_200_n N_TE_B_M1032_g 0.00683255f $X=1.19 $Y=1.17 $X2=0
+ $Y2=0
cc_176 N_A_126_74#_c_174_n N_TE_B_c_326_n 0.00105979f $X=1.355 $Y=1.26 $X2=0
+ $Y2=0
cc_177 N_A_126_74#_c_197_n N_TE_B_c_326_n 0.0341742f $X=0.78 $Y=1.985 $X2=0
+ $Y2=0
cc_178 N_A_126_74#_c_200_n N_TE_B_c_326_n 0.00141415f $X=1.19 $Y=1.17 $X2=0
+ $Y2=0
cc_179 N_A_126_74#_c_174_n N_TE_B_c_327_n 0.0138531f $X=1.355 $Y=1.26 $X2=0
+ $Y2=0
cc_180 N_A_126_74#_c_197_n N_TE_B_c_327_n 0.023773f $X=0.78 $Y=1.985 $X2=0 $Y2=0
cc_181 N_A_126_74#_c_200_n N_TE_B_c_327_n 0.00461804f $X=1.19 $Y=1.17 $X2=0
+ $Y2=0
cc_182 N_A_126_74#_c_197_n N_TE_B_c_345_n 0.00223123f $X=0.78 $Y=1.985 $X2=0
+ $Y2=0
cc_183 N_A_126_74#_c_190_n N_TE_B_c_328_n 0.0138531f $X=1.825 $Y=1.26 $X2=0
+ $Y2=0
cc_184 N_A_126_74#_c_191_n N_TE_B_c_329_n 0.0138531f $X=2.255 $Y=1.26 $X2=0
+ $Y2=0
cc_185 N_A_126_74#_c_192_n N_TE_B_c_330_n 0.0138531f $X=2.685 $Y=1.26 $X2=0
+ $Y2=0
cc_186 N_A_126_74#_c_193_n N_TE_B_c_331_n 0.0138531f $X=3.185 $Y=1.26 $X2=0
+ $Y2=0
cc_187 N_A_126_74#_c_194_n N_TE_B_c_332_n 0.0138531f $X=3.615 $Y=1.26 $X2=0
+ $Y2=0
cc_188 N_A_126_74#_c_195_n N_TE_B_c_333_n 0.0138531f $X=4.115 $Y=1.26 $X2=0
+ $Y2=0
cc_189 N_A_126_74#_c_196_n N_TE_B_c_334_n 0.0138531f $X=4.545 $Y=1.26 $X2=0
+ $Y2=0
cc_190 N_A_126_74#_c_173_n N_TE_B_c_335_n 0.0138531f $X=1.75 $Y=1.26 $X2=0 $Y2=0
cc_191 N_A_126_74#_c_176_n N_TE_B_c_336_n 0.0138531f $X=2.18 $Y=1.26 $X2=0 $Y2=0
cc_192 N_A_126_74#_c_178_n N_TE_B_c_337_n 0.0138531f $X=2.61 $Y=1.26 $X2=0 $Y2=0
cc_193 N_A_126_74#_c_180_n N_TE_B_c_338_n 0.0138531f $X=3.11 $Y=1.26 $X2=0 $Y2=0
cc_194 N_A_126_74#_c_182_n N_TE_B_c_339_n 0.0138531f $X=3.54 $Y=1.26 $X2=0 $Y2=0
cc_195 N_A_126_74#_c_184_n N_TE_B_c_340_n 0.0138531f $X=4.04 $Y=1.26 $X2=0 $Y2=0
cc_196 N_A_126_74#_c_186_n N_TE_B_c_341_n 0.0138531f $X=4.47 $Y=1.26 $X2=0 $Y2=0
cc_197 N_A_126_74#_c_200_n TE_B 0.0333272f $X=1.19 $Y=1.17 $X2=0 $Y2=0
cc_198 N_A_126_74#_c_189_n N_A_M1004_g 0.0160416f $X=4.975 $Y=1.185 $X2=0 $Y2=0
cc_199 N_A_126_74#_c_197_n N_VPWR_c_654_n 0.0451069f $X=0.78 $Y=1.985 $X2=0
+ $Y2=0
cc_200 N_A_126_74#_c_197_n N_VPWR_c_662_n 0.0145938f $X=0.78 $Y=1.985 $X2=0
+ $Y2=0
cc_201 N_A_126_74#_c_197_n N_VPWR_c_652_n 0.0120466f $X=0.78 $Y=1.985 $X2=0
+ $Y2=0
cc_202 N_A_126_74#_c_197_n N_A_239_368#_c_758_n 0.0755732f $X=0.78 $Y=1.985
+ $X2=0 $Y2=0
cc_203 N_A_126_74#_c_173_n N_A_239_368#_c_759_n 0.00107716f $X=1.75 $Y=1.26
+ $X2=0 $Y2=0
cc_204 N_A_126_74#_c_174_n N_A_239_368#_c_760_n 6.32757e-19 $X=1.355 $Y=1.26
+ $X2=0 $Y2=0
cc_205 N_A_126_74#_c_197_n N_A_239_368#_c_760_n 0.0116261f $X=0.78 $Y=1.985
+ $X2=0 $Y2=0
cc_206 N_A_126_74#_c_200_n N_A_239_368#_c_760_n 0.00886618f $X=1.19 $Y=1.17
+ $X2=0 $Y2=0
cc_207 N_A_126_74#_c_178_n N_A_239_368#_c_762_n 6.15194e-19 $X=2.61 $Y=1.26
+ $X2=0 $Y2=0
cc_208 N_A_126_74#_c_182_n N_A_239_368#_c_764_n 6.15637e-19 $X=3.54 $Y=1.26
+ $X2=0 $Y2=0
cc_209 N_A_126_74#_c_176_n N_A_239_368#_c_783_n 2.1586e-19 $X=2.18 $Y=1.26 $X2=0
+ $Y2=0
cc_210 N_A_126_74#_c_180_n N_A_239_368#_c_784_n 2.15823e-19 $X=3.11 $Y=1.26
+ $X2=0 $Y2=0
cc_211 N_A_126_74#_c_184_n N_A_239_368#_c_772_n 4.19958e-19 $X=4.04 $Y=1.26
+ $X2=0 $Y2=0
cc_212 N_A_126_74#_c_188_n N_Z_c_934_n 3.54739e-19 $X=4.9 $Y=1.26 $X2=0 $Y2=0
cc_213 N_A_126_74#_c_198_n N_VGND_c_1053_n 0.0257911f $X=1.19 $Y=0.49 $X2=0
+ $Y2=0
cc_214 N_A_126_74#_c_199_n N_VGND_c_1053_n 4.50615e-19 $X=1.19 $Y=0.49 $X2=0
+ $Y2=0
cc_215 N_A_126_74#_c_175_n N_VGND_c_1054_n 0.0148429f $X=1.825 $Y=1.185 $X2=0
+ $Y2=0
cc_216 N_A_126_74#_c_176_n N_VGND_c_1054_n 0.00230361f $X=2.18 $Y=1.26 $X2=0
+ $Y2=0
cc_217 N_A_126_74#_c_177_n N_VGND_c_1054_n 0.00198331f $X=2.255 $Y=1.185 $X2=0
+ $Y2=0
cc_218 N_A_126_74#_c_198_n N_VGND_c_1054_n 7.79228e-19 $X=1.19 $Y=0.49 $X2=0
+ $Y2=0
cc_219 N_A_126_74#_c_199_n N_VGND_c_1054_n 2.62006e-19 $X=1.19 $Y=0.49 $X2=0
+ $Y2=0
cc_220 N_A_126_74#_c_177_n N_VGND_c_1055_n 6.14817e-19 $X=2.255 $Y=1.185 $X2=0
+ $Y2=0
cc_221 N_A_126_74#_c_179_n N_VGND_c_1055_n 0.0134319f $X=2.685 $Y=1.185 $X2=0
+ $Y2=0
cc_222 N_A_126_74#_c_180_n N_VGND_c_1055_n 0.00391613f $X=3.11 $Y=1.26 $X2=0
+ $Y2=0
cc_223 N_A_126_74#_c_181_n N_VGND_c_1055_n 0.00581358f $X=3.185 $Y=1.185 $X2=0
+ $Y2=0
cc_224 N_A_126_74#_c_181_n N_VGND_c_1056_n 6.13445e-19 $X=3.185 $Y=1.185 $X2=0
+ $Y2=0
cc_225 N_A_126_74#_c_183_n N_VGND_c_1056_n 0.0134156f $X=3.615 $Y=1.185 $X2=0
+ $Y2=0
cc_226 N_A_126_74#_c_184_n N_VGND_c_1056_n 0.00391613f $X=4.04 $Y=1.26 $X2=0
+ $Y2=0
cc_227 N_A_126_74#_c_185_n N_VGND_c_1056_n 0.00581358f $X=4.115 $Y=1.185 $X2=0
+ $Y2=0
cc_228 N_A_126_74#_c_185_n N_VGND_c_1057_n 5.77505e-19 $X=4.115 $Y=1.185 $X2=0
+ $Y2=0
cc_229 N_A_126_74#_c_187_n N_VGND_c_1057_n 0.0115133f $X=4.545 $Y=1.185 $X2=0
+ $Y2=0
cc_230 N_A_126_74#_c_188_n N_VGND_c_1057_n 0.00205835f $X=4.9 $Y=1.26 $X2=0
+ $Y2=0
cc_231 N_A_126_74#_c_189_n N_VGND_c_1057_n 0.010743f $X=4.975 $Y=1.185 $X2=0
+ $Y2=0
cc_232 N_A_126_74#_c_175_n N_VGND_c_1058_n 0.00383152f $X=1.825 $Y=1.185 $X2=0
+ $Y2=0
cc_233 N_A_126_74#_c_198_n N_VGND_c_1058_n 0.0320951f $X=1.19 $Y=0.49 $X2=0
+ $Y2=0
cc_234 N_A_126_74#_c_199_n N_VGND_c_1058_n 0.00191653f $X=1.19 $Y=0.49 $X2=0
+ $Y2=0
cc_235 N_A_126_74#_c_177_n N_VGND_c_1060_n 0.00434272f $X=2.255 $Y=1.185 $X2=0
+ $Y2=0
cc_236 N_A_126_74#_c_179_n N_VGND_c_1060_n 0.00383152f $X=2.685 $Y=1.185 $X2=0
+ $Y2=0
cc_237 N_A_126_74#_c_181_n N_VGND_c_1062_n 0.00434272f $X=3.185 $Y=1.185 $X2=0
+ $Y2=0
cc_238 N_A_126_74#_c_183_n N_VGND_c_1062_n 0.00383152f $X=3.615 $Y=1.185 $X2=0
+ $Y2=0
cc_239 N_A_126_74#_c_185_n N_VGND_c_1064_n 0.00434272f $X=4.115 $Y=1.185 $X2=0
+ $Y2=0
cc_240 N_A_126_74#_c_187_n N_VGND_c_1064_n 0.00383152f $X=4.545 $Y=1.185 $X2=0
+ $Y2=0
cc_241 N_A_126_74#_c_189_n N_VGND_c_1066_n 0.00383152f $X=4.975 $Y=1.185 $X2=0
+ $Y2=0
cc_242 N_A_126_74#_c_175_n N_VGND_c_1067_n 0.00762539f $X=1.825 $Y=1.185 $X2=0
+ $Y2=0
cc_243 N_A_126_74#_c_177_n N_VGND_c_1067_n 0.00820284f $X=2.255 $Y=1.185 $X2=0
+ $Y2=0
cc_244 N_A_126_74#_c_179_n N_VGND_c_1067_n 0.0075754f $X=2.685 $Y=1.185 $X2=0
+ $Y2=0
cc_245 N_A_126_74#_c_181_n N_VGND_c_1067_n 0.00820718f $X=3.185 $Y=1.185 $X2=0
+ $Y2=0
cc_246 N_A_126_74#_c_183_n N_VGND_c_1067_n 0.0075754f $X=3.615 $Y=1.185 $X2=0
+ $Y2=0
cc_247 N_A_126_74#_c_185_n N_VGND_c_1067_n 0.00820718f $X=4.115 $Y=1.185 $X2=0
+ $Y2=0
cc_248 N_A_126_74#_c_187_n N_VGND_c_1067_n 0.0075754f $X=4.545 $Y=1.185 $X2=0
+ $Y2=0
cc_249 N_A_126_74#_c_189_n N_VGND_c_1067_n 0.00757637f $X=4.975 $Y=1.185 $X2=0
+ $Y2=0
cc_250 N_A_126_74#_c_198_n N_VGND_c_1067_n 0.0247858f $X=1.19 $Y=0.49 $X2=0
+ $Y2=0
cc_251 N_A_126_74#_c_173_n N_A_293_74#_c_1160_n 0.00966561f $X=1.75 $Y=1.26
+ $X2=0 $Y2=0
cc_252 N_A_126_74#_c_175_n N_A_293_74#_c_1160_n 0.00143488f $X=1.825 $Y=1.185
+ $X2=0 $Y2=0
cc_253 N_A_126_74#_c_198_n N_A_293_74#_c_1160_n 0.0739685f $X=1.19 $Y=0.49 $X2=0
+ $Y2=0
cc_254 N_A_126_74#_c_199_n N_A_293_74#_c_1160_n 0.00633652f $X=1.19 $Y=0.49
+ $X2=0 $Y2=0
cc_255 N_A_126_74#_c_173_n N_A_293_74#_c_1161_n 0.00283425f $X=1.75 $Y=1.26
+ $X2=0 $Y2=0
cc_256 N_A_126_74#_c_176_n N_A_293_74#_c_1161_n 0.00750207f $X=2.18 $Y=1.26
+ $X2=0 $Y2=0
cc_257 N_A_126_74#_c_190_n N_A_293_74#_c_1161_n 0.00728747f $X=1.825 $Y=1.26
+ $X2=0 $Y2=0
cc_258 N_A_126_74#_c_191_n N_A_293_74#_c_1161_n 0.00663107f $X=2.255 $Y=1.26
+ $X2=0 $Y2=0
cc_259 N_A_126_74#_c_173_n N_A_293_74#_c_1162_n 0.00209968f $X=1.75 $Y=1.26
+ $X2=0 $Y2=0
cc_260 N_A_126_74#_c_197_n N_A_293_74#_c_1162_n 0.0050605f $X=0.78 $Y=1.985
+ $X2=0 $Y2=0
cc_261 N_A_126_74#_c_200_n N_A_293_74#_c_1162_n 0.00294869f $X=1.19 $Y=1.17
+ $X2=0 $Y2=0
cc_262 N_A_126_74#_c_175_n N_A_293_74#_c_1163_n 4.44315e-19 $X=1.825 $Y=1.185
+ $X2=0 $Y2=0
cc_263 N_A_126_74#_c_177_n N_A_293_74#_c_1163_n 0.0106978f $X=2.255 $Y=1.185
+ $X2=0 $Y2=0
cc_264 N_A_126_74#_c_178_n N_A_293_74#_c_1163_n 0.0100752f $X=2.61 $Y=1.26 $X2=0
+ $Y2=0
cc_265 N_A_126_74#_c_179_n N_A_293_74#_c_1163_n 0.00195128f $X=2.685 $Y=1.185
+ $X2=0 $Y2=0
cc_266 N_A_126_74#_c_191_n N_A_293_74#_c_1163_n 0.00333129f $X=2.255 $Y=1.26
+ $X2=0 $Y2=0
cc_267 N_A_126_74#_c_178_n N_A_293_74#_c_1164_n 0.00283425f $X=2.61 $Y=1.26
+ $X2=0 $Y2=0
cc_268 N_A_126_74#_c_180_n N_A_293_74#_c_1164_n 0.00841771f $X=3.11 $Y=1.26
+ $X2=0 $Y2=0
cc_269 N_A_126_74#_c_192_n N_A_293_74#_c_1164_n 0.00728747f $X=2.685 $Y=1.26
+ $X2=0 $Y2=0
cc_270 N_A_126_74#_c_193_n N_A_293_74#_c_1164_n 0.00663107f $X=3.185 $Y=1.26
+ $X2=0 $Y2=0
cc_271 N_A_126_74#_c_179_n N_A_293_74#_c_1165_n 4.87722e-19 $X=2.685 $Y=1.185
+ $X2=0 $Y2=0
cc_272 N_A_126_74#_c_181_n N_A_293_74#_c_1165_n 0.0106102f $X=3.185 $Y=1.185
+ $X2=0 $Y2=0
cc_273 N_A_126_74#_c_182_n N_A_293_74#_c_1165_n 0.0100752f $X=3.54 $Y=1.26 $X2=0
+ $Y2=0
cc_274 N_A_126_74#_c_183_n N_A_293_74#_c_1165_n 0.00195128f $X=3.615 $Y=1.185
+ $X2=0 $Y2=0
cc_275 N_A_126_74#_c_193_n N_A_293_74#_c_1165_n 0.00552993f $X=3.185 $Y=1.26
+ $X2=0 $Y2=0
cc_276 N_A_126_74#_c_182_n N_A_293_74#_c_1166_n 0.00283425f $X=3.54 $Y=1.26
+ $X2=0 $Y2=0
cc_277 N_A_126_74#_c_184_n N_A_293_74#_c_1166_n 0.00841166f $X=4.04 $Y=1.26
+ $X2=0 $Y2=0
cc_278 N_A_126_74#_c_194_n N_A_293_74#_c_1166_n 0.00728747f $X=3.615 $Y=1.26
+ $X2=0 $Y2=0
cc_279 N_A_126_74#_c_195_n N_A_293_74#_c_1166_n 0.00663107f $X=4.115 $Y=1.26
+ $X2=0 $Y2=0
cc_280 N_A_126_74#_c_183_n N_A_293_74#_c_1167_n 4.87722e-19 $X=3.615 $Y=1.185
+ $X2=0 $Y2=0
cc_281 N_A_126_74#_c_185_n N_A_293_74#_c_1167_n 0.0106102f $X=4.115 $Y=1.185
+ $X2=0 $Y2=0
cc_282 N_A_126_74#_c_186_n N_A_293_74#_c_1167_n 0.0039817f $X=4.47 $Y=1.26 $X2=0
+ $Y2=0
cc_283 N_A_126_74#_c_187_n N_A_293_74#_c_1167_n 0.00229866f $X=4.545 $Y=1.185
+ $X2=0 $Y2=0
cc_284 N_A_126_74#_c_195_n N_A_293_74#_c_1167_n 0.0011642f $X=4.115 $Y=1.26
+ $X2=0 $Y2=0
cc_285 N_A_126_74#_c_186_n N_A_293_74#_c_1168_n 0.00314343f $X=4.47 $Y=1.26
+ $X2=0 $Y2=0
cc_286 N_A_126_74#_c_188_n N_A_293_74#_c_1168_n 0.0164668f $X=4.9 $Y=1.26 $X2=0
+ $Y2=0
cc_287 N_A_126_74#_c_196_n N_A_293_74#_c_1168_n 0.00815912f $X=4.545 $Y=1.26
+ $X2=0 $Y2=0
cc_288 N_A_126_74#_c_189_n N_A_293_74#_c_1169_n 9.48753e-19 $X=4.975 $Y=1.185
+ $X2=0 $Y2=0
cc_289 N_A_126_74#_c_189_n N_A_293_74#_c_1170_n 0.0026408f $X=4.975 $Y=1.185
+ $X2=0 $Y2=0
cc_290 N_A_126_74#_c_178_n N_A_293_74#_c_1175_n 0.00209812f $X=2.61 $Y=1.26
+ $X2=0 $Y2=0
cc_291 N_A_126_74#_c_191_n N_A_293_74#_c_1175_n 2.34165e-19 $X=2.255 $Y=1.26
+ $X2=0 $Y2=0
cc_292 N_A_126_74#_c_182_n N_A_293_74#_c_1176_n 0.00209812f $X=3.54 $Y=1.26
+ $X2=0 $Y2=0
cc_293 N_A_126_74#_c_193_n N_A_293_74#_c_1176_n 2.34165e-19 $X=3.185 $Y=1.26
+ $X2=0 $Y2=0
cc_294 N_A_126_74#_c_186_n N_A_293_74#_c_1177_n 0.00399647f $X=4.47 $Y=1.26
+ $X2=0 $Y2=0
cc_295 N_A_126_74#_c_195_n N_A_293_74#_c_1177_n 0.00511841f $X=4.115 $Y=1.26
+ $X2=0 $Y2=0
cc_296 N_TE_B_c_359_n N_A_c_503_n 0.0120492f $X=4.965 $Y=1.765 $X2=0 $Y2=0
cc_297 N_TE_B_c_334_n N_A_c_502_n 0.00905775f $X=4.875 $Y=1.65 $X2=0 $Y2=0
cc_298 N_TE_B_c_326_n N_VPWR_c_654_n 0.0366774f $X=0.555 $Y=1.765 $X2=0 $Y2=0
cc_299 TE_B N_VPWR_c_654_n 0.0253033f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_300 N_TE_B_c_345_n N_VPWR_c_655_n 0.0170945f $X=1.565 $Y=1.765 $X2=0 $Y2=0
cc_301 N_TE_B_c_328_n N_VPWR_c_655_n 0.00166497f $X=1.975 $Y=1.65 $X2=0 $Y2=0
cc_302 N_TE_B_c_347_n N_VPWR_c_655_n 0.00693368f $X=2.065 $Y=1.765 $X2=0 $Y2=0
cc_303 N_TE_B_c_347_n N_VPWR_c_656_n 0.00445602f $X=2.065 $Y=1.765 $X2=0 $Y2=0
cc_304 N_TE_B_c_349_n N_VPWR_c_656_n 0.00413917f $X=2.515 $Y=1.765 $X2=0 $Y2=0
cc_305 N_TE_B_c_347_n N_VPWR_c_657_n 6.37984e-19 $X=2.065 $Y=1.765 $X2=0 $Y2=0
cc_306 N_TE_B_c_349_n N_VPWR_c_657_n 0.0139335f $X=2.515 $Y=1.765 $X2=0 $Y2=0
cc_307 N_TE_B_c_330_n N_VPWR_c_657_n 0.00166497f $X=2.925 $Y=1.65 $X2=0 $Y2=0
cc_308 N_TE_B_c_351_n N_VPWR_c_657_n 0.00693368f $X=3.015 $Y=1.765 $X2=0 $Y2=0
cc_309 N_TE_B_c_351_n N_VPWR_c_658_n 0.00445602f $X=3.015 $Y=1.765 $X2=0 $Y2=0
cc_310 N_TE_B_c_353_n N_VPWR_c_658_n 0.00413917f $X=3.465 $Y=1.765 $X2=0 $Y2=0
cc_311 N_TE_B_c_351_n N_VPWR_c_659_n 6.37984e-19 $X=3.015 $Y=1.765 $X2=0 $Y2=0
cc_312 N_TE_B_c_353_n N_VPWR_c_659_n 0.0139335f $X=3.465 $Y=1.765 $X2=0 $Y2=0
cc_313 N_TE_B_c_332_n N_VPWR_c_659_n 0.00166497f $X=3.875 $Y=1.65 $X2=0 $Y2=0
cc_314 N_TE_B_c_355_n N_VPWR_c_659_n 0.00699801f $X=3.965 $Y=1.765 $X2=0 $Y2=0
cc_315 N_TE_B_c_355_n N_VPWR_c_660_n 0.00445602f $X=3.965 $Y=1.765 $X2=0 $Y2=0
cc_316 N_TE_B_c_357_n N_VPWR_c_660_n 0.00445602f $X=4.415 $Y=1.765 $X2=0 $Y2=0
cc_317 N_TE_B_c_357_n N_VPWR_c_661_n 0.00598632f $X=4.415 $Y=1.765 $X2=0 $Y2=0
cc_318 N_TE_B_c_359_n N_VPWR_c_661_n 0.00546951f $X=4.965 $Y=1.765 $X2=0 $Y2=0
cc_319 N_TE_B_c_326_n N_VPWR_c_662_n 0.00445602f $X=0.555 $Y=1.765 $X2=0 $Y2=0
cc_320 N_TE_B_c_345_n N_VPWR_c_662_n 0.00413917f $X=1.565 $Y=1.765 $X2=0 $Y2=0
cc_321 N_TE_B_c_359_n N_VPWR_c_663_n 0.0044313f $X=4.965 $Y=1.765 $X2=0 $Y2=0
cc_322 N_TE_B_c_326_n N_VPWR_c_652_n 0.00865368f $X=0.555 $Y=1.765 $X2=0 $Y2=0
cc_323 N_TE_B_c_345_n N_VPWR_c_652_n 0.00822528f $X=1.565 $Y=1.765 $X2=0 $Y2=0
cc_324 N_TE_B_c_347_n N_VPWR_c_652_n 0.00857378f $X=2.065 $Y=1.765 $X2=0 $Y2=0
cc_325 N_TE_B_c_349_n N_VPWR_c_652_n 0.00817726f $X=2.515 $Y=1.765 $X2=0 $Y2=0
cc_326 N_TE_B_c_351_n N_VPWR_c_652_n 0.00857378f $X=3.015 $Y=1.765 $X2=0 $Y2=0
cc_327 N_TE_B_c_353_n N_VPWR_c_652_n 0.00817726f $X=3.465 $Y=1.765 $X2=0 $Y2=0
cc_328 N_TE_B_c_355_n N_VPWR_c_652_n 0.00857378f $X=3.965 $Y=1.765 $X2=0 $Y2=0
cc_329 N_TE_B_c_357_n N_VPWR_c_652_n 0.00857797f $X=4.415 $Y=1.765 $X2=0 $Y2=0
cc_330 N_TE_B_c_359_n N_VPWR_c_652_n 0.00853652f $X=4.965 $Y=1.765 $X2=0 $Y2=0
cc_331 N_TE_B_c_326_n N_A_239_368#_c_758_n 0.0019935f $X=0.555 $Y=1.765 $X2=0
+ $Y2=0
cc_332 N_TE_B_c_345_n N_A_239_368#_c_758_n 0.00894148f $X=1.565 $Y=1.765 $X2=0
+ $Y2=0
cc_333 N_TE_B_c_327_n N_A_239_368#_c_759_n 0.0017174f $X=1.475 $Y=1.65 $X2=0
+ $Y2=0
cc_334 N_TE_B_c_345_n N_A_239_368#_c_759_n 0.00952222f $X=1.565 $Y=1.765 $X2=0
+ $Y2=0
cc_335 N_TE_B_c_328_n N_A_239_368#_c_759_n 0.00938446f $X=1.975 $Y=1.65 $X2=0
+ $Y2=0
cc_336 N_TE_B_c_347_n N_A_239_368#_c_759_n 0.00775614f $X=2.065 $Y=1.765 $X2=0
+ $Y2=0
cc_337 N_TE_B_c_335_n N_A_239_368#_c_759_n 0.00514292f $X=1.565 $Y=1.67 $X2=0
+ $Y2=0
cc_338 N_TE_B_c_336_n N_A_239_368#_c_759_n 0.00327334f $X=2.065 $Y=1.67 $X2=0
+ $Y2=0
cc_339 N_TE_B_c_326_n N_A_239_368#_c_760_n 4.62965e-19 $X=0.555 $Y=1.765 $X2=0
+ $Y2=0
cc_340 N_TE_B_c_327_n N_A_239_368#_c_760_n 0.0114653f $X=1.475 $Y=1.65 $X2=0
+ $Y2=0
cc_341 N_TE_B_c_345_n N_A_239_368#_c_761_n 7.7138e-19 $X=1.565 $Y=1.765 $X2=0
+ $Y2=0
cc_342 N_TE_B_c_347_n N_A_239_368#_c_761_n 0.0134555f $X=2.065 $Y=1.765 $X2=0
+ $Y2=0
cc_343 N_TE_B_c_349_n N_A_239_368#_c_761_n 0.00741212f $X=2.515 $Y=1.765 $X2=0
+ $Y2=0
cc_344 N_TE_B_c_329_n N_A_239_368#_c_762_n 0.00141557f $X=2.425 $Y=1.65 $X2=0
+ $Y2=0
cc_345 N_TE_B_c_349_n N_A_239_368#_c_762_n 0.00899887f $X=2.515 $Y=1.765 $X2=0
+ $Y2=0
cc_346 N_TE_B_c_330_n N_A_239_368#_c_762_n 0.00938534f $X=2.925 $Y=1.65 $X2=0
+ $Y2=0
cc_347 N_TE_B_c_351_n N_A_239_368#_c_762_n 0.00775614f $X=3.015 $Y=1.765 $X2=0
+ $Y2=0
cc_348 N_TE_B_c_337_n N_A_239_368#_c_762_n 0.00448748f $X=2.515 $Y=1.67 $X2=0
+ $Y2=0
cc_349 N_TE_B_c_338_n N_A_239_368#_c_762_n 0.00327334f $X=3.015 $Y=1.67 $X2=0
+ $Y2=0
cc_350 N_TE_B_c_349_n N_A_239_368#_c_763_n 7.7138e-19 $X=2.515 $Y=1.765 $X2=0
+ $Y2=0
cc_351 N_TE_B_c_351_n N_A_239_368#_c_763_n 0.0134555f $X=3.015 $Y=1.765 $X2=0
+ $Y2=0
cc_352 N_TE_B_c_353_n N_A_239_368#_c_763_n 0.00741212f $X=3.465 $Y=1.765 $X2=0
+ $Y2=0
cc_353 N_TE_B_c_331_n N_A_239_368#_c_764_n 0.00141557f $X=3.375 $Y=1.65 $X2=0
+ $Y2=0
cc_354 N_TE_B_c_353_n N_A_239_368#_c_764_n 0.00899887f $X=3.465 $Y=1.765 $X2=0
+ $Y2=0
cc_355 N_TE_B_c_332_n N_A_239_368#_c_764_n 0.00938534f $X=3.875 $Y=1.65 $X2=0
+ $Y2=0
cc_356 N_TE_B_c_355_n N_A_239_368#_c_764_n 0.00800872f $X=3.965 $Y=1.765 $X2=0
+ $Y2=0
cc_357 N_TE_B_c_339_n N_A_239_368#_c_764_n 0.00448793f $X=3.465 $Y=1.67 $X2=0
+ $Y2=0
cc_358 N_TE_B_c_340_n N_A_239_368#_c_764_n 0.0037082f $X=3.965 $Y=1.67 $X2=0
+ $Y2=0
cc_359 N_TE_B_c_355_n N_A_239_368#_c_765_n 0.0085677f $X=3.965 $Y=1.765 $X2=0
+ $Y2=0
cc_360 N_TE_B_c_357_n N_A_239_368#_c_765_n 0.0103138f $X=4.415 $Y=1.765 $X2=0
+ $Y2=0
cc_361 N_TE_B_c_359_n N_A_239_368#_c_765_n 6.63528e-19 $X=4.965 $Y=1.765 $X2=0
+ $Y2=0
cc_362 N_TE_B_c_334_n N_A_239_368#_c_817_n 0.00748522f $X=4.875 $Y=1.65 $X2=0
+ $Y2=0
cc_363 N_TE_B_c_359_n N_A_239_368#_c_817_n 0.0124894f $X=4.965 $Y=1.765 $X2=0
+ $Y2=0
cc_364 N_TE_B_c_359_n N_A_239_368#_c_819_n 4.20803e-19 $X=4.965 $Y=1.765 $X2=0
+ $Y2=0
cc_365 N_TE_B_c_357_n N_A_239_368#_c_820_n 6.4805e-19 $X=4.415 $Y=1.765 $X2=0
+ $Y2=0
cc_366 N_TE_B_c_359_n N_A_239_368#_c_820_n 0.00920373f $X=4.965 $Y=1.765 $X2=0
+ $Y2=0
cc_367 N_TE_B_c_359_n N_A_239_368#_c_767_n 0.00313312f $X=4.965 $Y=1.765 $X2=0
+ $Y2=0
cc_368 N_TE_B_c_347_n N_A_239_368#_c_783_n 9.70881e-19 $X=2.065 $Y=1.765 $X2=0
+ $Y2=0
cc_369 N_TE_B_c_329_n N_A_239_368#_c_783_n 0.00814436f $X=2.425 $Y=1.65 $X2=0
+ $Y2=0
cc_370 N_TE_B_c_336_n N_A_239_368#_c_783_n 0.00133274f $X=2.065 $Y=1.67 $X2=0
+ $Y2=0
cc_371 N_TE_B_c_351_n N_A_239_368#_c_784_n 9.70881e-19 $X=3.015 $Y=1.765 $X2=0
+ $Y2=0
cc_372 N_TE_B_c_331_n N_A_239_368#_c_784_n 0.00814391f $X=3.375 $Y=1.65 $X2=0
+ $Y2=0
cc_373 N_TE_B_c_338_n N_A_239_368#_c_784_n 0.00133274f $X=3.015 $Y=1.67 $X2=0
+ $Y2=0
cc_374 N_TE_B_c_353_n N_A_239_368#_c_772_n 8.00899e-19 $X=3.465 $Y=1.765 $X2=0
+ $Y2=0
cc_375 N_TE_B_c_355_n N_A_239_368#_c_772_n 0.00660358f $X=3.965 $Y=1.765 $X2=0
+ $Y2=0
cc_376 N_TE_B_c_333_n N_A_239_368#_c_772_n 0.00996496f $X=4.325 $Y=1.65 $X2=0
+ $Y2=0
cc_377 N_TE_B_c_357_n N_A_239_368#_c_772_n 0.0155478f $X=4.415 $Y=1.765 $X2=0
+ $Y2=0
cc_378 N_TE_B_c_359_n N_A_239_368#_c_772_n 0.00165413f $X=4.965 $Y=1.765 $X2=0
+ $Y2=0
cc_379 N_TE_B_c_340_n N_A_239_368#_c_772_n 0.0016238f $X=3.965 $Y=1.67 $X2=0
+ $Y2=0
cc_380 N_TE_B_c_341_n N_A_239_368#_c_772_n 0.0056829f $X=4.415 $Y=1.67 $X2=0
+ $Y2=0
cc_381 N_TE_B_c_334_n N_Z_c_934_n 0.0117352f $X=4.875 $Y=1.65 $X2=0 $Y2=0
cc_382 N_TE_B_c_359_n N_Z_c_934_n 0.00204317f $X=4.965 $Y=1.765 $X2=0 $Y2=0
cc_383 N_TE_B_M1032_g N_VGND_c_1053_n 0.0148726f $X=0.555 $Y=0.74 $X2=0 $Y2=0
cc_384 N_TE_B_c_326_n N_VGND_c_1053_n 0.00148634f $X=0.555 $Y=1.765 $X2=0 $Y2=0
cc_385 TE_B N_VGND_c_1053_n 0.0207716f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_386 N_TE_B_M1032_g N_VGND_c_1058_n 0.00383152f $X=0.555 $Y=0.74 $X2=0 $Y2=0
cc_387 N_TE_B_M1032_g N_VGND_c_1067_n 0.00762539f $X=0.555 $Y=0.74 $X2=0 $Y2=0
cc_388 N_TE_B_c_328_n N_A_293_74#_c_1161_n 0.00395446f $X=1.975 $Y=1.65 $X2=0
+ $Y2=0
cc_389 N_TE_B_c_335_n N_A_293_74#_c_1162_n 0.00139793f $X=1.565 $Y=1.67 $X2=0
+ $Y2=0
cc_390 N_TE_B_c_337_n N_A_293_74#_c_1164_n 0.00443434f $X=2.515 $Y=1.67 $X2=0
+ $Y2=0
cc_391 N_TE_B_c_339_n N_A_293_74#_c_1166_n 0.00447887f $X=3.465 $Y=1.67 $X2=0
+ $Y2=0
cc_392 N_TE_B_c_334_n N_A_293_74#_c_1168_n 3.86969e-19 $X=4.875 $Y=1.65 $X2=0
+ $Y2=0
cc_393 N_TE_B_c_341_n N_A_293_74#_c_1168_n 0.00439745f $X=4.415 $Y=1.67 $X2=0
+ $Y2=0
cc_394 N_TE_B_c_329_n N_A_293_74#_c_1175_n 0.00197752f $X=2.425 $Y=1.65 $X2=0
+ $Y2=0
cc_395 N_TE_B_c_331_n N_A_293_74#_c_1176_n 0.00194861f $X=3.375 $Y=1.65 $X2=0
+ $Y2=0
cc_396 N_TE_B_c_333_n N_A_293_74#_c_1177_n 0.00191711f $X=4.325 $Y=1.65 $X2=0
+ $Y2=0
cc_397 N_A_c_503_n N_VPWR_c_663_n 0.00278257f $X=5.415 $Y=1.765 $X2=0 $Y2=0
cc_398 N_A_c_504_n N_VPWR_c_663_n 0.00278257f $X=5.865 $Y=1.765 $X2=0 $Y2=0
cc_399 N_A_c_505_n N_VPWR_c_663_n 0.00278257f $X=6.315 $Y=1.765 $X2=0 $Y2=0
cc_400 N_A_c_506_n N_VPWR_c_663_n 0.00278271f $X=6.815 $Y=1.765 $X2=0 $Y2=0
cc_401 N_A_c_507_n N_VPWR_c_663_n 0.00278271f $X=7.265 $Y=1.765 $X2=0 $Y2=0
cc_402 N_A_c_508_n N_VPWR_c_663_n 0.00278271f $X=7.715 $Y=1.765 $X2=0 $Y2=0
cc_403 N_A_c_509_n N_VPWR_c_663_n 0.00278271f $X=8.165 $Y=1.765 $X2=0 $Y2=0
cc_404 N_A_c_510_n N_VPWR_c_663_n 0.00278271f $X=8.615 $Y=1.765 $X2=0 $Y2=0
cc_405 N_A_c_503_n N_VPWR_c_652_n 0.00353905f $X=5.415 $Y=1.765 $X2=0 $Y2=0
cc_406 N_A_c_504_n N_VPWR_c_652_n 0.00353822f $X=5.865 $Y=1.765 $X2=0 $Y2=0
cc_407 N_A_c_505_n N_VPWR_c_652_n 0.00354283f $X=6.315 $Y=1.765 $X2=0 $Y2=0
cc_408 N_A_c_506_n N_VPWR_c_652_n 0.00354284f $X=6.815 $Y=1.765 $X2=0 $Y2=0
cc_409 N_A_c_507_n N_VPWR_c_652_n 0.00353823f $X=7.265 $Y=1.765 $X2=0 $Y2=0
cc_410 N_A_c_508_n N_VPWR_c_652_n 0.00353823f $X=7.715 $Y=1.765 $X2=0 $Y2=0
cc_411 N_A_c_509_n N_VPWR_c_652_n 0.00353823f $X=8.165 $Y=1.765 $X2=0 $Y2=0
cc_412 N_A_c_510_n N_VPWR_c_652_n 0.00357317f $X=8.615 $Y=1.765 $X2=0 $Y2=0
cc_413 N_A_c_503_n N_A_239_368#_c_819_n 0.00191419f $X=5.415 $Y=1.765 $X2=0
+ $Y2=0
cc_414 N_A_c_503_n N_A_239_368#_c_820_n 0.00919154f $X=5.415 $Y=1.765 $X2=0
+ $Y2=0
cc_415 N_A_c_504_n N_A_239_368#_c_820_n 6.22492e-19 $X=5.865 $Y=1.765 $X2=0
+ $Y2=0
cc_416 N_A_c_503_n N_A_239_368#_c_766_n 0.0108414f $X=5.415 $Y=1.765 $X2=0 $Y2=0
cc_417 N_A_c_504_n N_A_239_368#_c_766_n 0.0108414f $X=5.865 $Y=1.765 $X2=0 $Y2=0
cc_418 N_A_c_503_n N_A_239_368#_c_767_n 0.00171731f $X=5.415 $Y=1.765 $X2=0
+ $Y2=0
cc_419 N_A_c_503_n N_A_239_368#_c_842_n 5.7112e-19 $X=5.415 $Y=1.765 $X2=0 $Y2=0
cc_420 N_A_c_504_n N_A_239_368#_c_842_n 0.00766499f $X=5.865 $Y=1.765 $X2=0
+ $Y2=0
cc_421 N_A_c_505_n N_A_239_368#_c_842_n 0.00756708f $X=6.315 $Y=1.765 $X2=0
+ $Y2=0
cc_422 N_A_c_506_n N_A_239_368#_c_842_n 7.75606e-19 $X=6.815 $Y=1.765 $X2=0
+ $Y2=0
cc_423 N_A_c_505_n N_A_239_368#_c_768_n 0.0111147f $X=6.315 $Y=1.765 $X2=0 $Y2=0
cc_424 N_A_c_506_n N_A_239_368#_c_768_n 0.0131082f $X=6.815 $Y=1.765 $X2=0 $Y2=0
cc_425 N_A_c_507_n N_A_239_368#_c_769_n 0.0128349f $X=7.265 $Y=1.765 $X2=0 $Y2=0
cc_426 N_A_c_508_n N_A_239_368#_c_769_n 0.0128349f $X=7.715 $Y=1.765 $X2=0 $Y2=0
cc_427 N_A_c_509_n N_A_239_368#_c_770_n 0.0128349f $X=8.165 $Y=1.765 $X2=0 $Y2=0
cc_428 N_A_c_510_n N_A_239_368#_c_770_n 0.0137046f $X=8.615 $Y=1.765 $X2=0 $Y2=0
cc_429 A N_A_239_368#_c_771_n 0.0211447f $X=8.795 $Y=1.58 $X2=0 $Y2=0
cc_430 N_A_c_504_n N_A_239_368#_c_773_n 0.00175197f $X=5.865 $Y=1.765 $X2=0
+ $Y2=0
cc_431 N_A_c_505_n N_A_239_368#_c_773_n 0.00175197f $X=6.315 $Y=1.765 $X2=0
+ $Y2=0
cc_432 N_A_M1004_g N_Z_c_944_n 0.00431189f $X=5.405 $Y=0.74 $X2=0 $Y2=0
cc_433 N_A_M1004_g N_Z_c_931_n 0.00432757f $X=5.405 $Y=0.74 $X2=0 $Y2=0
cc_434 N_A_M1007_g N_Z_c_931_n 0.00522824f $X=5.835 $Y=0.74 $X2=0 $Y2=0
cc_435 A N_Z_c_931_n 0.0107752f $X=8.795 $Y=1.58 $X2=0 $Y2=0
cc_436 N_A_c_502_n N_Z_c_931_n 0.0179489f $X=8.615 $Y=1.557 $X2=0 $Y2=0
cc_437 N_A_c_503_n N_Z_c_938_n 0.00352902f $X=5.415 $Y=1.765 $X2=0 $Y2=0
cc_438 N_A_c_504_n N_Z_c_938_n 0.00352902f $X=5.865 $Y=1.765 $X2=0 $Y2=0
cc_439 N_A_c_503_n N_Z_c_951_n 0.00279093f $X=5.415 $Y=1.765 $X2=0 $Y2=0
cc_440 N_A_c_504_n N_Z_c_951_n 0.00554349f $X=5.865 $Y=1.765 $X2=0 $Y2=0
cc_441 N_A_c_504_n N_Z_c_953_n 0.0172359f $X=5.865 $Y=1.765 $X2=0 $Y2=0
cc_442 N_A_c_505_n N_Z_c_953_n 0.0151078f $X=6.315 $Y=1.765 $X2=0 $Y2=0
cc_443 A N_Z_c_953_n 0.029833f $X=8.795 $Y=1.58 $X2=0 $Y2=0
cc_444 N_A_c_502_n N_Z_c_953_n 0.00236017f $X=8.615 $Y=1.557 $X2=0 $Y2=0
cc_445 N_A_c_506_n N_Z_c_957_n 0.00999032f $X=6.815 $Y=1.765 $X2=0 $Y2=0
cc_446 N_A_c_507_n N_Z_c_957_n 5.7112e-19 $X=7.265 $Y=1.765 $X2=0 $Y2=0
cc_447 N_A_M1013_g N_Z_c_932_n 0.00881059f $X=6.695 $Y=0.74 $X2=0 $Y2=0
cc_448 N_A_M1017_g N_Z_c_932_n 0.0125415f $X=7.195 $Y=0.74 $X2=0 $Y2=0
cc_449 N_A_c_502_n N_Z_c_932_n 0.00394597f $X=8.615 $Y=1.557 $X2=0 $Y2=0
cc_450 N_A_c_506_n N_Z_c_962_n 0.0120074f $X=6.815 $Y=1.765 $X2=0 $Y2=0
cc_451 N_A_c_507_n N_Z_c_962_n 0.0120074f $X=7.265 $Y=1.765 $X2=0 $Y2=0
cc_452 A N_Z_c_962_n 0.0393875f $X=8.795 $Y=1.58 $X2=0 $Y2=0
cc_453 N_A_c_502_n N_Z_c_962_n 0.00131036f $X=8.615 $Y=1.557 $X2=0 $Y2=0
cc_454 N_A_M1022_g N_Z_c_933_n 0.0121483f $X=7.625 $Y=0.74 $X2=0 $Y2=0
cc_455 N_A_M1024_g N_Z_c_933_n 0.0125508f $X=8.055 $Y=0.74 $X2=0 $Y2=0
cc_456 N_A_M1029_g N_Z_c_933_n 0.00249598f $X=8.625 $Y=0.74 $X2=0 $Y2=0
cc_457 A N_Z_c_933_n 0.0788927f $X=8.795 $Y=1.58 $X2=0 $Y2=0
cc_458 N_A_c_502_n N_Z_c_933_n 0.00790514f $X=8.615 $Y=1.557 $X2=0 $Y2=0
cc_459 N_A_c_508_n N_Z_c_971_n 0.0120074f $X=7.715 $Y=1.765 $X2=0 $Y2=0
cc_460 N_A_c_509_n N_Z_c_971_n 0.0119526f $X=8.165 $Y=1.765 $X2=0 $Y2=0
cc_461 A N_Z_c_971_n 0.0393875f $X=8.795 $Y=1.58 $X2=0 $Y2=0
cc_462 N_A_c_502_n N_Z_c_971_n 0.00130754f $X=8.615 $Y=1.557 $X2=0 $Y2=0
cc_463 N_A_c_503_n N_Z_c_934_n 0.00504225f $X=5.415 $Y=1.765 $X2=0 $Y2=0
cc_464 N_A_c_502_n N_Z_c_934_n 0.0113896f $X=8.615 $Y=1.557 $X2=0 $Y2=0
cc_465 N_A_c_503_n N_Z_c_940_n 0.00198966f $X=5.415 $Y=1.765 $X2=0 $Y2=0
cc_466 A N_Z_c_940_n 0.0142664f $X=8.795 $Y=1.58 $X2=0 $Y2=0
cc_467 N_A_c_502_n N_Z_c_940_n 0.0129759f $X=8.615 $Y=1.557 $X2=0 $Y2=0
cc_468 N_A_M1007_g N_Z_c_935_n 0.0187836f $X=5.835 $Y=0.74 $X2=0 $Y2=0
cc_469 N_A_M1010_g N_Z_c_935_n 0.0122111f $X=6.265 $Y=0.74 $X2=0 $Y2=0
cc_470 A N_Z_c_935_n 0.0208778f $X=8.795 $Y=1.58 $X2=0 $Y2=0
cc_471 N_A_c_502_n N_Z_c_935_n 0.00221617f $X=8.615 $Y=1.557 $X2=0 $Y2=0
cc_472 N_A_M1010_g N_Z_c_936_n 0.00330153f $X=6.265 $Y=0.74 $X2=0 $Y2=0
cc_473 N_A_M1013_g N_Z_c_936_n 0.00638767f $X=6.695 $Y=0.74 $X2=0 $Y2=0
cc_474 N_A_M1017_g N_Z_c_936_n 7.96756e-19 $X=7.195 $Y=0.74 $X2=0 $Y2=0
cc_475 A N_Z_c_936_n 0.077942f $X=8.795 $Y=1.58 $X2=0 $Y2=0
cc_476 N_A_c_502_n N_Z_c_936_n 0.00229127f $X=8.615 $Y=1.557 $X2=0 $Y2=0
cc_477 N_A_c_506_n N_Z_c_989_n 4.27055e-19 $X=6.815 $Y=1.765 $X2=0 $Y2=0
cc_478 A N_Z_c_989_n 0.025478f $X=8.795 $Y=1.58 $X2=0 $Y2=0
cc_479 N_A_c_502_n N_Z_c_989_n 0.00167458f $X=8.615 $Y=1.557 $X2=0 $Y2=0
cc_480 A N_Z_c_937_n 0.0143877f $X=8.795 $Y=1.58 $X2=0 $Y2=0
cc_481 N_A_c_502_n N_Z_c_937_n 0.00231317f $X=8.615 $Y=1.557 $X2=0 $Y2=0
cc_482 N_A_c_506_n N_Z_c_994_n 5.7112e-19 $X=6.815 $Y=1.765 $X2=0 $Y2=0
cc_483 N_A_c_507_n N_Z_c_994_n 0.0105121f $X=7.265 $Y=1.765 $X2=0 $Y2=0
cc_484 N_A_c_508_n N_Z_c_994_n 0.0105121f $X=7.715 $Y=1.765 $X2=0 $Y2=0
cc_485 N_A_c_509_n N_Z_c_994_n 5.7112e-19 $X=8.165 $Y=1.765 $X2=0 $Y2=0
cc_486 A N_Z_c_994_n 0.0237598f $X=8.795 $Y=1.58 $X2=0 $Y2=0
cc_487 N_A_c_502_n N_Z_c_994_n 0.00144162f $X=8.615 $Y=1.557 $X2=0 $Y2=0
cc_488 N_A_c_508_n N_Z_c_1000_n 5.7112e-19 $X=7.715 $Y=1.765 $X2=0 $Y2=0
cc_489 N_A_c_509_n N_Z_c_1000_n 0.0105121f $X=8.165 $Y=1.765 $X2=0 $Y2=0
cc_490 N_A_c_510_n N_Z_c_1000_n 0.011241f $X=8.615 $Y=1.765 $X2=0 $Y2=0
cc_491 A N_Z_c_1000_n 0.0237598f $X=8.795 $Y=1.58 $X2=0 $Y2=0
cc_492 N_A_c_502_n N_Z_c_1000_n 0.00144904f $X=8.615 $Y=1.557 $X2=0 $Y2=0
cc_493 N_A_M1004_g N_VGND_c_1057_n 2.43373e-19 $X=5.405 $Y=0.74 $X2=0 $Y2=0
cc_494 N_A_M1004_g N_VGND_c_1066_n 0.00278271f $X=5.405 $Y=0.74 $X2=0 $Y2=0
cc_495 N_A_M1007_g N_VGND_c_1066_n 0.00278271f $X=5.835 $Y=0.74 $X2=0 $Y2=0
cc_496 N_A_M1010_g N_VGND_c_1066_n 0.00278271f $X=6.265 $Y=0.74 $X2=0 $Y2=0
cc_497 N_A_M1013_g N_VGND_c_1066_n 0.00278271f $X=6.695 $Y=0.74 $X2=0 $Y2=0
cc_498 N_A_M1017_g N_VGND_c_1066_n 0.00279469f $X=7.195 $Y=0.74 $X2=0 $Y2=0
cc_499 N_A_M1022_g N_VGND_c_1066_n 0.00278247f $X=7.625 $Y=0.74 $X2=0 $Y2=0
cc_500 N_A_M1024_g N_VGND_c_1066_n 0.00278247f $X=8.055 $Y=0.74 $X2=0 $Y2=0
cc_501 N_A_M1029_g N_VGND_c_1066_n 0.00278247f $X=8.625 $Y=0.74 $X2=0 $Y2=0
cc_502 N_A_M1004_g N_VGND_c_1067_n 0.00353526f $X=5.405 $Y=0.74 $X2=0 $Y2=0
cc_503 N_A_M1007_g N_VGND_c_1067_n 0.00353428f $X=5.835 $Y=0.74 $X2=0 $Y2=0
cc_504 N_A_M1010_g N_VGND_c_1067_n 0.00353428f $X=6.265 $Y=0.74 $X2=0 $Y2=0
cc_505 N_A_M1013_g N_VGND_c_1067_n 0.00354087f $X=6.695 $Y=0.74 $X2=0 $Y2=0
cc_506 N_A_M1017_g N_VGND_c_1067_n 0.00353176f $X=7.195 $Y=0.74 $X2=0 $Y2=0
cc_507 N_A_M1022_g N_VGND_c_1067_n 0.00353427f $X=7.625 $Y=0.74 $X2=0 $Y2=0
cc_508 N_A_M1024_g N_VGND_c_1067_n 0.0035466f $X=8.055 $Y=0.74 $X2=0 $Y2=0
cc_509 N_A_M1029_g N_VGND_c_1067_n 0.00358318f $X=8.625 $Y=0.74 $X2=0 $Y2=0
cc_510 N_A_M1004_g N_A_293_74#_c_1168_n 0.00136516f $X=5.405 $Y=0.74 $X2=0 $Y2=0
cc_511 N_A_c_502_n N_A_293_74#_c_1168_n 9.50669e-19 $X=8.615 $Y=1.557 $X2=0
+ $Y2=0
cc_512 N_A_M1004_g N_A_293_74#_c_1170_n 9.59994e-19 $X=5.405 $Y=0.74 $X2=0 $Y2=0
cc_513 N_A_M1004_g N_A_293_74#_c_1171_n 0.0169972f $X=5.405 $Y=0.74 $X2=0 $Y2=0
cc_514 N_A_M1007_g N_A_293_74#_c_1171_n 0.013026f $X=5.835 $Y=0.74 $X2=0 $Y2=0
cc_515 N_A_M1010_g N_A_293_74#_c_1171_n 0.013026f $X=6.265 $Y=0.74 $X2=0 $Y2=0
cc_516 N_A_M1013_g N_A_293_74#_c_1171_n 0.0149406f $X=6.695 $Y=0.74 $X2=0 $Y2=0
cc_517 N_A_M1017_g N_A_293_74#_c_1172_n 0.00847867f $X=7.195 $Y=0.74 $X2=0 $Y2=0
cc_518 N_A_M1022_g N_A_293_74#_c_1172_n 0.00792642f $X=7.625 $Y=0.74 $X2=0 $Y2=0
cc_519 N_A_M1017_g N_A_293_74#_c_1243_n 5.56395e-19 $X=7.195 $Y=0.74 $X2=0 $Y2=0
cc_520 N_A_M1022_g N_A_293_74#_c_1243_n 0.00628318f $X=7.625 $Y=0.74 $X2=0 $Y2=0
cc_521 N_A_M1024_g N_A_293_74#_c_1243_n 0.00682969f $X=8.055 $Y=0.74 $X2=0 $Y2=0
cc_522 N_A_M1029_g N_A_293_74#_c_1243_n 6.35778e-19 $X=8.625 $Y=0.74 $X2=0 $Y2=0
cc_523 N_A_M1024_g N_A_293_74#_c_1173_n 0.00864553f $X=8.055 $Y=0.74 $X2=0 $Y2=0
cc_524 N_A_M1029_g N_A_293_74#_c_1173_n 0.0136117f $X=8.625 $Y=0.74 $X2=0 $Y2=0
cc_525 N_A_M1024_g N_A_293_74#_c_1174_n 7.53751e-19 $X=8.055 $Y=0.74 $X2=0 $Y2=0
cc_526 N_A_M1029_g N_A_293_74#_c_1174_n 0.0111505f $X=8.625 $Y=0.74 $X2=0 $Y2=0
cc_527 A N_A_293_74#_c_1174_n 0.023753f $X=8.795 $Y=1.58 $X2=0 $Y2=0
cc_528 N_A_M1013_g N_A_293_74#_c_1178_n 9.09403e-19 $X=6.695 $Y=0.74 $X2=0 $Y2=0
cc_529 N_A_M1017_g N_A_293_74#_c_1178_n 0.00935344f $X=7.195 $Y=0.74 $X2=0 $Y2=0
cc_530 N_A_M1022_g N_A_293_74#_c_1178_n 6.38633e-19 $X=7.625 $Y=0.74 $X2=0 $Y2=0
cc_531 N_A_M1022_g N_A_293_74#_c_1179_n 0.00254906f $X=7.625 $Y=0.74 $X2=0 $Y2=0
cc_532 N_A_M1024_g N_A_293_74#_c_1179_n 0.00254906f $X=8.055 $Y=0.74 $X2=0 $Y2=0
cc_533 N_VPWR_c_655_n N_A_239_368#_c_758_n 0.0654044f $X=1.79 $Y=2.09 $X2=0
+ $Y2=0
cc_534 N_VPWR_c_662_n N_A_239_368#_c_758_n 0.011066f $X=1.625 $Y=3.33 $X2=0
+ $Y2=0
cc_535 N_VPWR_c_652_n N_A_239_368#_c_758_n 0.00915947f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_536 N_VPWR_c_655_n N_A_239_368#_c_759_n 0.023488f $X=1.79 $Y=2.09 $X2=0 $Y2=0
cc_537 N_VPWR_c_655_n N_A_239_368#_c_761_n 0.0358509f $X=1.79 $Y=2.09 $X2=0
+ $Y2=0
cc_538 N_VPWR_c_656_n N_A_239_368#_c_761_n 0.0110241f $X=2.575 $Y=3.33 $X2=0
+ $Y2=0
cc_539 N_VPWR_c_657_n N_A_239_368#_c_761_n 0.0654044f $X=2.74 $Y=2.09 $X2=0
+ $Y2=0
cc_540 N_VPWR_c_652_n N_A_239_368#_c_761_n 0.00909194f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_541 N_VPWR_c_657_n N_A_239_368#_c_762_n 0.023488f $X=2.74 $Y=2.09 $X2=0 $Y2=0
cc_542 N_VPWR_c_657_n N_A_239_368#_c_763_n 0.0358509f $X=2.74 $Y=2.09 $X2=0
+ $Y2=0
cc_543 N_VPWR_c_658_n N_A_239_368#_c_763_n 0.0110241f $X=3.525 $Y=3.33 $X2=0
+ $Y2=0
cc_544 N_VPWR_c_659_n N_A_239_368#_c_763_n 0.0654044f $X=3.69 $Y=2.09 $X2=0
+ $Y2=0
cc_545 N_VPWR_c_652_n N_A_239_368#_c_763_n 0.00909194f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_546 N_VPWR_c_659_n N_A_239_368#_c_764_n 0.023488f $X=3.69 $Y=2.09 $X2=0 $Y2=0
cc_547 N_VPWR_c_660_n N_A_239_368#_c_765_n 0.014552f $X=4.525 $Y=3.33 $X2=0
+ $Y2=0
cc_548 N_VPWR_c_661_n N_A_239_368#_c_765_n 0.0266809f $X=4.69 $Y=2.455 $X2=0
+ $Y2=0
cc_549 N_VPWR_c_652_n N_A_239_368#_c_765_n 0.0119791f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_550 N_VPWR_M1027_d N_A_239_368#_c_817_n 0.00747406f $X=4.49 $Y=1.84 $X2=0
+ $Y2=0
cc_551 N_VPWR_c_661_n N_A_239_368#_c_817_n 0.0232685f $X=4.69 $Y=2.455 $X2=0
+ $Y2=0
cc_552 N_VPWR_c_663_n N_A_239_368#_c_766_n 0.03588f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_553 N_VPWR_c_652_n N_A_239_368#_c_766_n 0.0201952f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_554 N_VPWR_c_661_n N_A_239_368#_c_767_n 0.0119239f $X=4.69 $Y=2.455 $X2=0
+ $Y2=0
cc_555 N_VPWR_c_663_n N_A_239_368#_c_767_n 0.0235512f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_556 N_VPWR_c_652_n N_A_239_368#_c_767_n 0.0126924f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_557 N_VPWR_c_663_n N_A_239_368#_c_768_n 0.0442078f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_558 N_VPWR_c_652_n N_A_239_368#_c_768_n 0.0250141f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_559 N_VPWR_c_663_n N_A_239_368#_c_769_n 0.0460938f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_560 N_VPWR_c_652_n N_A_239_368#_c_769_n 0.0260732f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_561 N_VPWR_c_663_n N_A_239_368#_c_770_n 0.0640155f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_562 N_VPWR_c_652_n N_A_239_368#_c_770_n 0.0357926f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_563 N_VPWR_c_659_n N_A_239_368#_c_772_n 0.0375771f $X=3.69 $Y=2.09 $X2=0
+ $Y2=0
cc_564 N_VPWR_c_663_n N_A_239_368#_c_773_n 0.0235512f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_565 N_VPWR_c_652_n N_A_239_368#_c_773_n 0.0126924f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_566 N_VPWR_c_663_n N_A_239_368#_c_774_n 0.0121867f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_567 N_VPWR_c_652_n N_A_239_368#_c_774_n 0.00660921f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_568 N_VPWR_c_663_n N_A_239_368#_c_775_n 0.0121867f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_569 N_VPWR_c_652_n N_A_239_368#_c_775_n 0.00660921f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_570 N_A_239_368#_c_766_n N_Z_M1001_d 0.00247267f $X=5.925 $Y=2.99 $X2=0 $Y2=0
cc_571 N_A_239_368#_c_768_n N_Z_M1009_d 0.00250873f $X=6.955 $Y=2.99 $X2=0 $Y2=0
cc_572 N_A_239_368#_c_769_n N_Z_M1014_d 0.00197722f $X=7.855 $Y=2.99 $X2=0 $Y2=0
cc_573 N_A_239_368#_c_770_n N_Z_M1025_d 0.00197722f $X=8.755 $Y=2.99 $X2=0 $Y2=0
cc_574 N_A_239_368#_c_820_n N_Z_c_951_n 0.039994f $X=5.19 $Y=2.815 $X2=0 $Y2=0
cc_575 N_A_239_368#_c_766_n N_Z_c_951_n 0.012787f $X=5.925 $Y=2.99 $X2=0 $Y2=0
cc_576 N_A_239_368#_c_842_n N_Z_c_951_n 0.0289859f $X=6.09 $Y=2.455 $X2=0 $Y2=0
cc_577 N_A_239_368#_M1006_s N_Z_c_953_n 0.00359365f $X=5.94 $Y=1.84 $X2=0 $Y2=0
cc_578 N_A_239_368#_c_842_n N_Z_c_953_n 0.0171813f $X=6.09 $Y=2.455 $X2=0 $Y2=0
cc_579 N_A_239_368#_c_768_n N_Z_c_957_n 0.018923f $X=6.955 $Y=2.99 $X2=0 $Y2=0
cc_580 N_A_239_368#_c_902_p N_Z_c_957_n 0.0289859f $X=7.04 $Y=2.455 $X2=0 $Y2=0
cc_581 N_A_239_368#_M1011_s N_Z_c_962_n 0.00408911f $X=6.89 $Y=1.84 $X2=0 $Y2=0
cc_582 N_A_239_368#_c_902_p N_Z_c_962_n 0.0136682f $X=7.04 $Y=2.455 $X2=0 $Y2=0
cc_583 N_A_239_368#_M1021_s N_Z_c_971_n 0.00408911f $X=7.79 $Y=1.84 $X2=0 $Y2=0
cc_584 N_A_239_368#_c_906_p N_Z_c_971_n 0.0136682f $X=7.94 $Y=2.455 $X2=0 $Y2=0
cc_585 N_A_239_368#_c_817_n N_Z_c_934_n 0.00690535f $X=5.025 $Y=2.035 $X2=0
+ $Y2=0
cc_586 N_A_239_368#_c_819_n N_Z_c_934_n 0.0224729f $X=5.19 $Y=2.12 $X2=0 $Y2=0
cc_587 N_A_239_368#_c_772_n N_Z_c_934_n 0.00444027f $X=4.26 $Y=1.75 $X2=0 $Y2=0
cc_588 N_A_239_368#_c_819_n N_Z_c_1023_n 0.013092f $X=5.19 $Y=2.12 $X2=0 $Y2=0
cc_589 N_A_239_368#_c_902_p N_Z_c_994_n 0.0289859f $X=7.04 $Y=2.455 $X2=0 $Y2=0
cc_590 N_A_239_368#_c_769_n N_Z_c_994_n 0.0160777f $X=7.855 $Y=2.99 $X2=0 $Y2=0
cc_591 N_A_239_368#_c_906_p N_Z_c_994_n 0.0289859f $X=7.94 $Y=2.455 $X2=0 $Y2=0
cc_592 N_A_239_368#_c_906_p N_Z_c_1000_n 0.0289859f $X=7.94 $Y=2.455 $X2=0 $Y2=0
cc_593 N_A_239_368#_c_770_n N_Z_c_1000_n 0.0160777f $X=8.755 $Y=2.99 $X2=0 $Y2=0
cc_594 N_A_239_368#_c_771_n N_Z_c_1000_n 0.0533059f $X=8.84 $Y=2.115 $X2=0 $Y2=0
cc_595 N_A_239_368#_c_759_n N_A_293_74#_c_1161_n 0.0276514f $X=2.125 $Y=1.75
+ $X2=0 $Y2=0
cc_596 N_A_239_368#_c_783_n N_A_293_74#_c_1161_n 0.0128886f $X=2.25 $Y=1.75
+ $X2=0 $Y2=0
cc_597 N_A_239_368#_c_759_n N_A_293_74#_c_1162_n 0.0123447f $X=2.125 $Y=1.75
+ $X2=0 $Y2=0
cc_598 N_A_239_368#_c_762_n N_A_293_74#_c_1164_n 0.0334284f $X=3.075 $Y=1.75
+ $X2=0 $Y2=0
cc_599 N_A_239_368#_c_784_n N_A_293_74#_c_1164_n 0.0114485f $X=3.2 $Y=1.75 $X2=0
+ $Y2=0
cc_600 N_A_239_368#_c_764_n N_A_293_74#_c_1166_n 0.0347493f $X=4.025 $Y=1.75
+ $X2=0 $Y2=0
cc_601 N_A_239_368#_c_772_n N_A_293_74#_c_1166_n 0.00993644f $X=4.26 $Y=1.75
+ $X2=0 $Y2=0
cc_602 N_A_239_368#_c_817_n N_A_293_74#_c_1168_n 0.0115593f $X=5.025 $Y=2.035
+ $X2=0 $Y2=0
cc_603 N_A_239_368#_c_772_n N_A_293_74#_c_1168_n 0.00412109f $X=4.26 $Y=1.75
+ $X2=0 $Y2=0
cc_604 N_A_239_368#_c_762_n N_A_293_74#_c_1175_n 0.0130422f $X=3.075 $Y=1.75
+ $X2=0 $Y2=0
cc_605 N_A_239_368#_c_783_n N_A_293_74#_c_1175_n 0.00562336f $X=2.25 $Y=1.75
+ $X2=0 $Y2=0
cc_606 N_A_239_368#_c_764_n N_A_293_74#_c_1176_n 0.0115863f $X=4.025 $Y=1.75
+ $X2=0 $Y2=0
cc_607 N_A_239_368#_c_784_n N_A_293_74#_c_1176_n 0.00723003f $X=3.2 $Y=1.75
+ $X2=0 $Y2=0
cc_608 N_A_239_368#_c_772_n N_A_293_74#_c_1177_n 0.0199108f $X=4.26 $Y=1.75
+ $X2=0 $Y2=0
cc_609 N_Z_c_935_n N_A_293_74#_M1007_s 0.00177442f $X=6.315 $Y=0.975 $X2=0 $Y2=0
cc_610 N_Z_c_932_n N_A_293_74#_M1013_s 0.0025999f $X=7.325 $Y=1.095 $X2=0 $Y2=0
cc_611 N_Z_c_933_n N_A_293_74#_M1022_s 0.00182874f $X=8.175 $Y=1.095 $X2=0 $Y2=0
cc_612 N_Z_c_931_n N_A_293_74#_c_1168_n 0.01351f $X=5.59 $Y=1.55 $X2=0 $Y2=0
cc_613 N_Z_c_934_n N_A_293_74#_c_1168_n 0.0284919f $X=5.455 $Y=1.665 $X2=0 $Y2=0
cc_614 N_Z_c_944_n N_A_293_74#_c_1170_n 0.0151706f $X=5.59 $Y=1.13 $X2=0 $Y2=0
cc_615 N_Z_c_931_n N_A_293_74#_c_1170_n 0.00560041f $X=5.59 $Y=1.55 $X2=0 $Y2=0
cc_616 N_Z_M1004_d N_A_293_74#_c_1171_n 0.00180346f $X=5.48 $Y=0.37 $X2=0 $Y2=0
cc_617 N_Z_M1010_d N_A_293_74#_c_1171_n 0.00180787f $X=6.34 $Y=0.37 $X2=0 $Y2=0
cc_618 N_Z_c_944_n N_A_293_74#_c_1171_n 0.0156016f $X=5.59 $Y=1.13 $X2=0 $Y2=0
cc_619 N_Z_c_932_n N_A_293_74#_c_1171_n 0.00438759f $X=7.325 $Y=1.095 $X2=0
+ $Y2=0
cc_620 N_Z_c_935_n N_A_293_74#_c_1171_n 0.0497987f $X=6.315 $Y=0.975 $X2=0 $Y2=0
cc_621 N_Z_M1017_d N_A_293_74#_c_1172_n 0.00184993f $X=7.27 $Y=0.37 $X2=0 $Y2=0
cc_622 N_Z_c_932_n N_A_293_74#_c_1172_n 0.00305575f $X=7.325 $Y=1.095 $X2=0
+ $Y2=0
cc_623 N_Z_c_1044_p N_A_293_74#_c_1172_n 0.0113217f $X=7.41 $Y=0.78 $X2=0 $Y2=0
cc_624 N_Z_c_933_n N_A_293_74#_c_1172_n 0.00304353f $X=8.175 $Y=1.095 $X2=0
+ $Y2=0
cc_625 N_Z_c_933_n N_A_293_74#_c_1243_n 0.0157867f $X=8.175 $Y=1.095 $X2=0 $Y2=0
cc_626 N_Z_M1024_d N_A_293_74#_c_1173_n 0.00358944f $X=8.13 $Y=0.37 $X2=0 $Y2=0
cc_627 N_Z_c_933_n N_A_293_74#_c_1173_n 0.00304353f $X=8.175 $Y=1.095 $X2=0
+ $Y2=0
cc_628 N_Z_c_1049_p N_A_293_74#_c_1173_n 0.02087f $X=8.34 $Y=0.78 $X2=0 $Y2=0
cc_629 N_Z_c_933_n N_A_293_74#_c_1174_n 0.00540984f $X=8.175 $Y=1.095 $X2=0
+ $Y2=0
cc_630 N_Z_c_932_n N_A_293_74#_c_1178_n 0.0194125f $X=7.325 $Y=1.095 $X2=0 $Y2=0
cc_631 N_VGND_c_1054_n N_A_293_74#_c_1160_n 0.0281649f $X=2.04 $Y=0.515 $X2=0
+ $Y2=0
cc_632 N_VGND_c_1058_n N_A_293_74#_c_1160_n 0.00749631f $X=1.875 $Y=0 $X2=0
+ $Y2=0
cc_633 N_VGND_c_1067_n N_A_293_74#_c_1160_n 0.0062048f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_634 N_VGND_c_1054_n N_A_293_74#_c_1161_n 0.0198684f $X=2.04 $Y=0.515 $X2=0
+ $Y2=0
cc_635 N_VGND_c_1054_n N_A_293_74#_c_1163_n 0.0282477f $X=2.04 $Y=0.515 $X2=0
+ $Y2=0
cc_636 N_VGND_c_1055_n N_A_293_74#_c_1163_n 0.0294122f $X=2.9 $Y=0.515 $X2=0
+ $Y2=0
cc_637 N_VGND_c_1060_n N_A_293_74#_c_1163_n 0.0109942f $X=2.735 $Y=0 $X2=0 $Y2=0
cc_638 N_VGND_c_1067_n N_A_293_74#_c_1163_n 0.00904371f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_639 N_VGND_c_1055_n N_A_293_74#_c_1164_n 0.0263224f $X=2.9 $Y=0.515 $X2=0
+ $Y2=0
cc_640 N_VGND_c_1055_n N_A_293_74#_c_1165_n 0.0296294f $X=2.9 $Y=0.515 $X2=0
+ $Y2=0
cc_641 N_VGND_c_1056_n N_A_293_74#_c_1165_n 0.0294122f $X=3.83 $Y=0.515 $X2=0
+ $Y2=0
cc_642 N_VGND_c_1062_n N_A_293_74#_c_1165_n 0.0109942f $X=3.665 $Y=0 $X2=0 $Y2=0
cc_643 N_VGND_c_1067_n N_A_293_74#_c_1165_n 0.00904371f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_644 N_VGND_c_1056_n N_A_293_74#_c_1166_n 0.0263224f $X=3.83 $Y=0.515 $X2=0
+ $Y2=0
cc_645 N_VGND_c_1056_n N_A_293_74#_c_1167_n 0.0296294f $X=3.83 $Y=0.515 $X2=0
+ $Y2=0
cc_646 N_VGND_c_1057_n N_A_293_74#_c_1167_n 0.0254585f $X=4.76 $Y=0.515 $X2=0
+ $Y2=0
cc_647 N_VGND_c_1064_n N_A_293_74#_c_1167_n 0.0109942f $X=4.595 $Y=0 $X2=0 $Y2=0
cc_648 N_VGND_c_1067_n N_A_293_74#_c_1167_n 0.00904371f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_649 N_VGND_c_1057_n N_A_293_74#_c_1168_n 0.0204885f $X=4.76 $Y=0.515 $X2=0
+ $Y2=0
cc_650 N_VGND_c_1057_n N_A_293_74#_c_1169_n 0.0175237f $X=4.76 $Y=0.515 $X2=0
+ $Y2=0
cc_651 N_VGND_c_1066_n N_A_293_74#_c_1169_n 0.0121867f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_652 N_VGND_c_1067_n N_A_293_74#_c_1169_n 0.00660921f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_653 N_VGND_c_1066_n N_A_293_74#_c_1171_n 0.102335f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_654 N_VGND_c_1067_n N_A_293_74#_c_1171_n 0.0560806f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_655 N_VGND_c_1066_n N_A_293_74#_c_1172_n 0.0333877f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_656 N_VGND_c_1067_n N_A_293_74#_c_1172_n 0.0187857f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_657 N_VGND_c_1066_n N_A_293_74#_c_1173_n 0.0659488f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_658 N_VGND_c_1067_n N_A_293_74#_c_1173_n 0.0367612f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_659 N_VGND_c_1066_n N_A_293_74#_c_1178_n 0.0231199f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_660 N_VGND_c_1067_n N_A_293_74#_c_1178_n 0.0125837f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_661 N_VGND_c_1066_n N_A_293_74#_c_1179_n 0.0231739f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_662 N_VGND_c_1067_n N_A_293_74#_c_1179_n 0.0125425f $X=8.88 $Y=0 $X2=0 $Y2=0
