* File: sky130_fd_sc_ls__o21ai_4.pex.spice
* Created: Wed Sep  2 11:18:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__O21AI_4%A1 3 5 7 10 12 14 17 19 21 24 26 28 34 35 51
+ 54
c85 35 0 1.69044e-19 $X=1.68 $Y=1.665
c86 10 0 7.72498e-20 $X=0.925 $Y=0.74
r87 51 52 6.90365 $w=3.84e-07 $l=5.5e-08 $layer=POLY_cond $X=1.8 $Y=1.542
+ $X2=1.855 $Y2=1.542
r88 49 51 21.3385 $w=3.84e-07 $l=1.7e-07 $layer=POLY_cond $X=1.63 $Y=1.542
+ $X2=1.8 $Y2=1.542
r89 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.63
+ $Y=1.485 $X2=1.63 $Y2=1.485
r90 47 49 28.2422 $w=3.84e-07 $l=2.25e-07 $layer=POLY_cond $X=1.405 $Y=1.542
+ $X2=1.63 $Y2=1.542
r91 46 47 6.27604 $w=3.84e-07 $l=5e-08 $layer=POLY_cond $X=1.355 $Y=1.542
+ $X2=1.405 $Y2=1.542
r92 45 50 8.84058 $w=4.58e-07 $l=3.4e-07 $layer=LI1_cond $X=1.29 $Y=1.55
+ $X2=1.63 $Y2=1.55
r93 44 46 8.15885 $w=3.84e-07 $l=6.5e-08 $layer=POLY_cond $X=1.29 $Y=1.542
+ $X2=1.355 $Y2=1.542
r94 44 45 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.29
+ $Y=1.485 $X2=1.29 $Y2=1.485
r95 42 44 42.0495 $w=3.84e-07 $l=3.35e-07 $layer=POLY_cond $X=0.955 $Y=1.542
+ $X2=1.29 $Y2=1.542
r96 41 42 3.76562 $w=3.84e-07 $l=3e-08 $layer=POLY_cond $X=0.925 $Y=1.542
+ $X2=0.955 $Y2=1.542
r97 38 39 1.25521 $w=3.84e-07 $l=1e-08 $layer=POLY_cond $X=0.495 $Y=1.542
+ $X2=0.505 $Y2=1.542
r98 35 50 1.30009 $w=4.58e-07 $l=5e-08 $layer=LI1_cond $X=1.68 $Y=1.55 $X2=1.63
+ $Y2=1.55
r99 34 45 2.34015 $w=4.58e-07 $l=9e-08 $layer=LI1_cond $X=1.2 $Y=1.55 $X2=1.29
+ $Y2=1.55
r100 34 54 3.96409 $w=4.58e-07 $l=1.15e-07 $layer=LI1_cond $X=1.2 $Y=1.55
+ $X2=1.085 $Y2=1.55
r101 32 41 39.5391 $w=3.84e-07 $l=3.15e-07 $layer=POLY_cond $X=0.61 $Y=1.542
+ $X2=0.925 $Y2=1.542
r102 32 39 13.1797 $w=3.84e-07 $l=1.05e-07 $layer=POLY_cond $X=0.61 $Y=1.542
+ $X2=0.505 $Y2=1.542
r103 31 54 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=0.61 $Y=1.485
+ $X2=1.085 $Y2=1.485
r104 31 32 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.61
+ $Y=1.485 $X2=0.61 $Y2=1.485
r105 26 52 24.8669 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=1.855 $Y=1.765
+ $X2=1.855 $Y2=1.542
r106 26 28 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.855 $Y=1.765
+ $X2=1.855 $Y2=2.4
r107 22 51 24.8669 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=1.8 $Y=1.32
+ $X2=1.8 $Y2=1.542
r108 22 24 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.8 $Y=1.32 $X2=1.8
+ $Y2=0.74
r109 19 47 24.8669 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=1.405 $Y=1.765
+ $X2=1.405 $Y2=1.542
r110 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.405 $Y=1.765
+ $X2=1.405 $Y2=2.4
r111 15 46 24.8669 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=1.355 $Y=1.32
+ $X2=1.355 $Y2=1.542
r112 15 17 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.355 $Y=1.32
+ $X2=1.355 $Y2=0.74
r113 12 42 24.8669 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=0.955 $Y=1.765
+ $X2=0.955 $Y2=1.542
r114 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.955 $Y=1.765
+ $X2=0.955 $Y2=2.4
r115 8 41 24.8669 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=0.925 $Y=1.32
+ $X2=0.925 $Y2=1.542
r116 8 10 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=0.925 $Y=1.32
+ $X2=0.925 $Y2=0.74
r117 5 39 24.8669 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=1.542
r118 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.4
r119 1 38 24.8669 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=0.495 $Y=1.32
+ $X2=0.495 $Y2=1.542
r120 1 3 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=0.495 $Y=1.32
+ $X2=0.495 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__O21AI_4%B1 1 3 4 6 7 9 10 12 13 15 16 17 18 20 21 22
+ 34
c72 18 0 1.87103e-19 $X=3.52 $Y=1.185
c73 13 0 6.95413e-20 $X=3.09 $Y=1.185
c74 7 0 6.95413e-20 $X=2.66 $Y=1.185
c75 4 0 6.11875e-20 $X=2.305 $Y=1.765
c76 1 0 1.88681e-19 $X=2.23 $Y=1.185
r77 33 35 9.83673 $w=4.41e-07 $l=9e-08 $layer=POLY_cond $X=3 $Y=1.475 $X2=3.09
+ $Y2=1.475
r78 33 34 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3
+ $Y=1.385 $X2=3 $Y2=1.385
r79 31 33 26.7778 $w=4.41e-07 $l=2.45e-07 $layer=POLY_cond $X=2.755 $Y=1.475
+ $X2=3 $Y2=1.475
r80 30 31 10.3832 $w=4.41e-07 $l=9.5e-08 $layer=POLY_cond $X=2.66 $Y=1.475
+ $X2=2.755 $Y2=1.475
r81 28 30 37.161 $w=4.41e-07 $l=3.4e-07 $layer=POLY_cond $X=2.32 $Y=1.475
+ $X2=2.66 $Y2=1.475
r82 28 29 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.32
+ $Y=1.385 $X2=2.32 $Y2=1.385
r83 26 28 1.63946 $w=4.41e-07 $l=1.5e-08 $layer=POLY_cond $X=2.305 $Y=1.475
+ $X2=2.32 $Y2=1.475
r84 25 26 8.19728 $w=4.41e-07 $l=7.5e-08 $layer=POLY_cond $X=2.23 $Y=1.475
+ $X2=2.305 $Y2=1.475
r85 22 34 11.213 $w=3.68e-07 $l=3.6e-07 $layer=LI1_cond $X=2.64 $Y=1.365 $X2=3
+ $Y2=1.365
r86 22 29 9.96707 $w=3.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2.64 $Y=1.365
+ $X2=2.32 $Y2=1.365
r87 21 29 4.98354 $w=3.68e-07 $l=1.6e-07 $layer=LI1_cond $X=2.16 $Y=1.365
+ $X2=2.32 $Y2=1.365
r88 18 20 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=3.52 $Y=1.185
+ $X2=3.52 $Y2=0.74
r89 17 35 30.6324 $w=4.41e-07 $l=2.497e-07 $layer=POLY_cond $X=3.165 $Y=1.26
+ $X2=3.09 $Y2=1.475
r90 16 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.445 $Y=1.26
+ $X2=3.52 $Y2=1.185
r91 16 17 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.445 $Y=1.26
+ $X2=3.165 $Y2=1.26
r92 13 35 28.2648 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=3.09 $Y=1.185
+ $X2=3.09 $Y2=1.475
r93 13 15 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=3.09 $Y=1.185
+ $X2=3.09 $Y2=0.74
r94 10 31 28.2648 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.755 $Y=1.765
+ $X2=2.755 $Y2=1.475
r95 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.755 $Y=1.765
+ $X2=2.755 $Y2=2.4
r96 7 30 28.2648 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.66 $Y=1.185
+ $X2=2.66 $Y2=1.475
r97 7 9 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.66 $Y=1.185
+ $X2=2.66 $Y2=0.74
r98 4 26 28.2648 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.305 $Y=1.765
+ $X2=2.305 $Y2=1.475
r99 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.305 $Y=1.765
+ $X2=2.305 $Y2=2.4
r100 1 25 28.2648 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.23 $Y=1.185
+ $X2=2.23 $Y2=1.475
r101 1 3 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.23 $Y=1.185
+ $X2=2.23 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__O21AI_4%A2 1 3 6 8 10 13 15 17 20 22 24 27 29 30 31
+ 32 49
c79 8 0 6.77325e-20 $X=4.35 $Y=1.765
r80 49 50 1.93834 $w=3.73e-07 $l=1.5e-08 $layer=POLY_cond $X=5.25 $Y=1.557
+ $X2=5.265 $Y2=1.557
r81 47 49 12.9223 $w=3.73e-07 $l=1e-07 $layer=POLY_cond $X=5.15 $Y=1.557
+ $X2=5.25 $Y2=1.557
r82 47 48 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.15
+ $Y=1.515 $X2=5.15 $Y2=1.515
r83 45 47 40.7051 $w=3.73e-07 $l=3.15e-07 $layer=POLY_cond $X=4.835 $Y=1.557
+ $X2=5.15 $Y2=1.557
r84 44 45 4.52279 $w=3.73e-07 $l=3.5e-08 $layer=POLY_cond $X=4.8 $Y=1.557
+ $X2=4.835 $Y2=1.557
r85 43 44 51.0429 $w=3.73e-07 $l=3.95e-07 $layer=POLY_cond $X=4.405 $Y=1.557
+ $X2=4.8 $Y2=1.557
r86 42 43 7.10724 $w=3.73e-07 $l=5.5e-08 $layer=POLY_cond $X=4.35 $Y=1.557
+ $X2=4.405 $Y2=1.557
r87 40 42 28.429 $w=3.73e-07 $l=2.2e-07 $layer=POLY_cond $X=4.13 $Y=1.557
+ $X2=4.35 $Y2=1.557
r88 40 41 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.13
+ $Y=1.515 $X2=4.13 $Y2=1.515
r89 38 40 20.0295 $w=3.73e-07 $l=1.55e-07 $layer=POLY_cond $X=3.975 $Y=1.557
+ $X2=4.13 $Y2=1.557
r90 32 48 9.91637 $w=4.28e-07 $l=3.7e-07 $layer=LI1_cond $X=5.52 $Y=1.565
+ $X2=5.15 $Y2=1.565
r91 31 48 2.94811 $w=4.28e-07 $l=1.1e-07 $layer=LI1_cond $X=5.04 $Y=1.565
+ $X2=5.15 $Y2=1.565
r92 30 31 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=4.56 $Y=1.565
+ $X2=5.04 $Y2=1.565
r93 30 41 11.5244 $w=4.28e-07 $l=4.3e-07 $layer=LI1_cond $X=4.56 $Y=1.565
+ $X2=4.13 $Y2=1.565
r94 29 41 1.34005 $w=4.28e-07 $l=5e-08 $layer=LI1_cond $X=4.08 $Y=1.565 $X2=4.13
+ $Y2=1.565
r95 25 50 24.162 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.265 $Y=1.35
+ $X2=5.265 $Y2=1.557
r96 25 27 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.265 $Y=1.35
+ $X2=5.265 $Y2=0.74
r97 22 49 24.162 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=5.25 $Y=1.765
+ $X2=5.25 $Y2=1.557
r98 22 24 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.25 $Y=1.765
+ $X2=5.25 $Y2=2.4
r99 18 45 24.162 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.835 $Y=1.35
+ $X2=4.835 $Y2=1.557
r100 18 20 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.835 $Y=1.35
+ $X2=4.835 $Y2=0.74
r101 15 44 24.162 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=4.8 $Y=1.765
+ $X2=4.8 $Y2=1.557
r102 15 17 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.8 $Y=1.765
+ $X2=4.8 $Y2=2.4
r103 11 43 24.162 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.405 $Y=1.35
+ $X2=4.405 $Y2=1.557
r104 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.405 $Y=1.35
+ $X2=4.405 $Y2=0.74
r105 8 42 24.162 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=4.35 $Y=1.765
+ $X2=4.35 $Y2=1.557
r106 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.35 $Y=1.765
+ $X2=4.35 $Y2=2.4
r107 4 38 24.162 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.975 $Y=1.35
+ $X2=3.975 $Y2=1.557
r108 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.975 $Y=1.35
+ $X2=3.975 $Y2=0.74
r109 1 38 16.1528 $w=3.73e-07 $l=2.63181e-07 $layer=POLY_cond $X=3.85 $Y=1.765
+ $X2=3.975 $Y2=1.557
r110 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.85 $Y=1.765
+ $X2=3.85 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__O21AI_4%VPWR 1 2 3 4 13 15 21 25 29 32 33 34 40 44
+ 54 55 61 64
r70 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r71 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r72 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r73 54 55 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r74 52 55 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=5.52 $Y2=3.33
r75 52 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r76 51 54 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=3.6 $Y=3.33
+ $X2=5.52 $Y2=3.33
r77 51 52 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r78 49 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.23 $Y=3.33
+ $X2=3.065 $Y2=3.33
r79 49 51 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.23 $Y=3.33 $X2=3.6
+ $Y2=3.33
r80 48 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r81 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r82 45 61 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.245 $Y=3.33
+ $X2=2.12 $Y2=3.33
r83 45 47 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=2.245 $Y=3.33
+ $X2=2.64 $Y2=3.33
r84 44 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.9 $Y=3.33
+ $X2=3.065 $Y2=3.33
r85 44 47 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=2.9 $Y=3.33 $X2=2.64
+ $Y2=3.33
r86 43 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r87 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r88 40 61 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.995 $Y=3.33
+ $X2=2.12 $Y2=3.33
r89 40 42 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.995 $Y=3.33
+ $X2=1.68 $Y2=3.33
r90 39 43 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r91 39 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r92 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r93 36 58 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.182 $Y2=3.33
r94 36 38 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.72 $Y2=3.33
r95 34 65 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=3.12 $Y2=3.33
r96 34 48 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=2.64 $Y2=3.33
r97 32 38 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.095 $Y=3.33
+ $X2=0.72 $Y2=3.33
r98 32 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.095 $Y=3.33
+ $X2=1.18 $Y2=3.33
r99 31 42 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=1.265 $Y=3.33
+ $X2=1.68 $Y2=3.33
r100 31 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.265 $Y=3.33
+ $X2=1.18 $Y2=3.33
r101 27 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.065 $Y=3.245
+ $X2=3.065 $Y2=3.33
r102 27 29 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=3.065 $Y=3.245
+ $X2=3.065 $Y2=2.805
r103 23 61 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.12 $Y=3.245
+ $X2=2.12 $Y2=3.33
r104 23 25 20.283 $w=2.48e-07 $l=4.4e-07 $layer=LI1_cond $X=2.12 $Y=3.245
+ $X2=2.12 $Y2=2.805
r105 19 33 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.18 $Y=3.245
+ $X2=1.18 $Y2=3.33
r106 19 21 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=1.18 $Y=3.245
+ $X2=1.18 $Y2=2.455
r107 15 18 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=0.24 $Y=1.985
+ $X2=0.24 $Y2=2.815
r108 13 58 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.182 $Y2=3.33
r109 13 18 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.24 $Y2=2.815
r110 4 29 600 $w=1.7e-07 $l=1.0761e-06 $layer=licon1_PDIFF $count=1 $X=2.83
+ $Y=1.84 $X2=3.065 $Y2=2.805
r111 3 25 600 $w=1.7e-07 $l=1.03729e-06 $layer=licon1_PDIFF $count=1 $X=1.93
+ $Y=1.84 $X2=2.08 $Y2=2.805
r112 2 21 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=1.03
+ $Y=1.84 $X2=1.18 $Y2=2.455
r113 1 18 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r114 1 15 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_LS__O21AI_4%A_116_368# 1 2 3 4 5 16 18 20 22 23 26 28 30
+ 31 32 33 36 38 42 50 53
c94 30 0 6.77325e-20 $X=3.625 $Y=2.46
r95 42 45 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=5.515 $Y=2.115
+ $X2=5.515 $Y2=2.815
r96 40 45 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=5.515 $Y=2.905
+ $X2=5.515 $Y2=2.815
r97 39 53 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.66 $Y=2.99
+ $X2=4.575 $Y2=2.99
r98 38 40 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.39 $Y=2.99
+ $X2=5.515 $Y2=2.905
r99 38 39 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=5.39 $Y=2.99
+ $X2=4.66 $Y2=2.99
r100 34 53 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.575 $Y=2.905
+ $X2=4.575 $Y2=2.99
r101 34 36 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=4.575 $Y=2.905
+ $X2=4.575 $Y2=2.455
r102 32 53 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.49 $Y=2.99
+ $X2=4.575 $Y2=2.99
r103 32 33 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=4.49 $Y=2.99 $X2=3.79
+ $Y2=2.99
r104 31 33 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.625 $Y=2.905
+ $X2=3.79 $Y2=2.99
r105 30 52 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.625 $Y=2.46
+ $X2=3.625 $Y2=2.375
r106 30 31 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=3.625 $Y=2.46
+ $X2=3.625 $Y2=2.905
r107 29 50 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.795 $Y=2.375
+ $X2=1.63 $Y2=2.375
r108 28 52 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.46 $Y=2.375
+ $X2=3.625 $Y2=2.375
r109 28 29 108.626 $w=1.68e-07 $l=1.665e-06 $layer=LI1_cond $X=3.46 $Y=2.375
+ $X2=1.795 $Y2=2.375
r110 24 50 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.63 $Y=2.46
+ $X2=1.63 $Y2=2.375
r111 24 26 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=1.63 $Y=2.46
+ $X2=1.63 $Y2=2.815
r112 23 50 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.63 $Y=2.29
+ $X2=1.63 $Y2=2.375
r113 22 49 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.63 $Y=2.12 $X2=1.63
+ $Y2=2.035
r114 22 23 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=1.63 $Y=2.12
+ $X2=1.63 $Y2=2.29
r115 21 47 4.70058 $w=1.7e-07 $l=1.94808e-07 $layer=LI1_cond $X=0.895 $Y=2.035
+ $X2=0.73 $Y2=1.97
r116 20 49 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.465 $Y=2.035
+ $X2=1.63 $Y2=2.035
r117 20 21 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.465 $Y=2.035
+ $X2=0.895 $Y2=2.035
r118 16 47 3.0656 $w=3.3e-07 $l=1.5e-07 $layer=LI1_cond $X=0.73 $Y=2.12 $X2=0.73
+ $Y2=1.97
r119 16 18 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=0.73 $Y=2.12
+ $X2=0.73 $Y2=2.815
r120 5 45 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=5.325
+ $Y=1.84 $X2=5.475 $Y2=2.815
r121 5 42 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=5.325
+ $Y=1.84 $X2=5.475 $Y2=2.115
r122 4 36 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=4.425
+ $Y=1.84 $X2=4.575 $Y2=2.455
r123 3 52 300 $w=1.7e-07 $l=6.83667e-07 $layer=licon1_PDIFF $count=2 $X=3.48
+ $Y=1.84 $X2=3.625 $Y2=2.455
r124 2 49 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=1.48
+ $Y=1.84 $X2=1.63 $Y2=2.115
r125 2 26 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.48
+ $Y=1.84 $X2=1.63 $Y2=2.815
r126 1 47 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.84 $X2=0.73 $Y2=1.985
r127 1 18 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.84 $X2=0.73 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_LS__O21AI_4%Y 1 2 3 4 5 16 20 24 28 33 38 43 45 46 49
r76 51 52 1.97128 $w=3.78e-07 $l=6.5e-08 $layer=LI1_cond $X=3.525 $Y=1.97
+ $X2=3.525 $Y2=2.035
r77 46 51 9.24987 $w=3.78e-07 $l=3.05e-07 $layer=LI1_cond $X=3.525 $Y=1.665
+ $X2=3.525 $Y2=1.97
r78 46 49 7.05482 $w=3.78e-07 $l=1.15e-07 $layer=LI1_cond $X=3.525 $Y=1.665
+ $X2=3.525 $Y2=1.55
r79 41 49 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=3.42 $Y=1.01
+ $X2=3.42 $Y2=1.55
r80 33 35 5.76222 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=2.405 $Y=0.8
+ $X2=2.405 $Y2=0.925
r81 29 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.29 $Y=2.035
+ $X2=4.125 $Y2=2.035
r82 28 45 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.86 $Y=2.035
+ $X2=5.025 $Y2=2.035
r83 28 29 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=4.86 $Y=2.035
+ $X2=4.29 $Y2=2.035
r84 25 52 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.715 $Y=2.035
+ $X2=3.525 $Y2=2.035
r85 24 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.96 $Y=2.035
+ $X2=4.125 $Y2=2.035
r86 24 25 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=3.96 $Y=2.035
+ $X2=3.715 $Y2=2.035
r87 21 35 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.53 $Y=0.925
+ $X2=2.405 $Y2=0.925
r88 20 41 5.2986 $w=2.83e-07 $l=8.5e-08 $layer=LI1_cond $X=3.362 $Y=0.925
+ $X2=3.362 $Y2=1.01
r89 20 38 5.05457 $w=2.83e-07 $l=1.25e-07 $layer=LI1_cond $X=3.362 $Y=0.925
+ $X2=3.362 $Y2=0.8
r90 20 21 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.22 $Y=0.925
+ $X2=2.53 $Y2=0.925
r91 16 51 2.12414 $w=3e-07 $l=1.9e-07 $layer=LI1_cond $X=3.335 $Y=1.97 $X2=3.525
+ $Y2=1.97
r92 16 18 30.9239 $w=2.98e-07 $l=8.05e-07 $layer=LI1_cond $X=3.335 $Y=1.97
+ $X2=2.53 $Y2=1.97
r93 5 45 300 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=2 $X=4.875
+ $Y=1.84 $X2=5.025 $Y2=2.115
r94 4 43 300 $w=1.7e-07 $l=3.61421e-07 $layer=licon1_PDIFF $count=2 $X=3.925
+ $Y=1.84 $X2=4.125 $Y2=2.115
r95 3 18 600 $w=1.7e-07 $l=2.33238e-07 $layer=licon1_PDIFF $count=1 $X=2.38
+ $Y=1.84 $X2=2.53 $Y2=2.01
r96 2 38 182 $w=1.7e-07 $l=4.95076e-07 $layer=licon1_NDIFF $count=1 $X=3.165
+ $Y=0.37 $X2=3.305 $Y2=0.8
r97 1 33 182 $w=1.7e-07 $l=4.95076e-07 $layer=licon1_NDIFF $count=1 $X=2.305
+ $Y=0.37 $X2=2.445 $Y2=0.8
.ends

.subckt PM_SKY130_FD_SC_LS__O21AI_4%A_27_74# 1 2 3 4 5 6 7 24 26 27 30 32 38 39
+ 40 45 46 47 50 52 56 59 62 67
c101 59 0 7.72498e-20 $X=1.14 $Y=0.965
c102 40 0 6.95413e-20 $X=3.675 $Y=0.34
c103 38 0 6.95413e-20 $X=2.71 $Y=0.34
r104 62 65 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=2.875 $Y=0.34
+ $X2=2.875 $Y2=0.55
r105 59 60 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=1.14 $Y=0.925
+ $X2=1.14 $Y2=1.065
r106 54 56 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=5.52 $Y=1.01
+ $X2=5.52 $Y2=0.515
r107 53 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.705 $Y=1.095
+ $X2=4.62 $Y2=1.095
r108 52 54 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.395 $Y=1.095
+ $X2=5.52 $Y2=1.01
r109 52 53 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.395 $Y=1.095
+ $X2=4.705 $Y2=1.095
r110 48 67 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.62 $Y=1.01
+ $X2=4.62 $Y2=1.095
r111 48 50 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=4.62 $Y=1.01
+ $X2=4.62 $Y2=0.515
r112 46 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.535 $Y=1.095
+ $X2=4.62 $Y2=1.095
r113 46 47 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.535 $Y=1.095
+ $X2=3.845 $Y2=1.095
r114 43 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.76 $Y=1.01
+ $X2=3.845 $Y2=1.095
r115 43 45 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=3.76 $Y=1.01
+ $X2=3.76 $Y2=0.515
r116 42 45 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=3.76 $Y=0.425
+ $X2=3.76 $Y2=0.515
r117 41 62 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.04 $Y=0.34
+ $X2=2.875 $Y2=0.34
r118 40 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.675 $Y=0.34
+ $X2=3.76 $Y2=0.425
r119 40 41 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=3.675 $Y=0.34
+ $X2=3.04 $Y2=0.34
r120 38 62 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.71 $Y=0.34
+ $X2=2.875 $Y2=0.34
r121 38 39 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=2.71 $Y=0.34
+ $X2=2.1 $Y2=0.34
r122 35 37 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.015 $Y=0.84
+ $X2=2.015 $Y2=0.495
r123 34 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.015 $Y=0.425
+ $X2=2.1 $Y2=0.34
r124 34 37 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=2.015 $Y=0.425
+ $X2=2.015 $Y2=0.495
r125 33 59 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.225 $Y=0.925
+ $X2=1.14 $Y2=0.925
r126 32 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.93 $Y=0.925
+ $X2=2.015 $Y2=0.84
r127 32 33 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=1.93 $Y=0.925
+ $X2=1.225 $Y2=0.925
r128 28 59 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=0.84
+ $X2=1.14 $Y2=0.925
r129 28 30 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.14 $Y=0.84
+ $X2=1.14 $Y2=0.515
r130 26 60 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.055 $Y=1.065
+ $X2=1.14 $Y2=1.065
r131 26 27 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.055 $Y=1.065
+ $X2=0.365 $Y2=1.065
r132 22 27 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.24 $Y=0.98
+ $X2=0.365 $Y2=1.065
r133 22 24 21.4354 $w=2.48e-07 $l=4.65e-07 $layer=LI1_cond $X=0.24 $Y=0.98
+ $X2=0.24 $Y2=0.515
r134 7 56 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.34
+ $Y=0.37 $X2=5.48 $Y2=0.515
r135 6 50 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.48
+ $Y=0.37 $X2=4.62 $Y2=0.515
r136 5 45 91 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=2 $X=3.595
+ $Y=0.37 $X2=3.76 $Y2=0.515
r137 4 65 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=2.735
+ $Y=0.37 $X2=2.875 $Y2=0.55
r138 3 37 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.875
+ $Y=0.37 $X2=2.015 $Y2=0.495
r139 2 59 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=1
+ $Y=0.37 $X2=1.14 $Y2=0.965
r140 2 30 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1
+ $Y=0.37 $X2=1.14 $Y2=0.515
r141 1 24 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__O21AI_4%VGND 1 2 3 4 15 19 21 25 29 31 33 38 43 50
+ 51 54 57 60 63
c84 25 0 1.87103e-19 $X=4.19 $Y=0.595
c85 19 0 1.88681e-19 $X=1.57 $Y=0.55
r86 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r87 60 61 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r88 57 58 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r89 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r90 51 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r91 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r92 48 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.215 $Y=0 $X2=5.05
+ $Y2=0
r93 48 50 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.215 $Y=0 $X2=5.52
+ $Y2=0
r94 47 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r95 47 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r96 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r97 44 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.355 $Y=0 $X2=4.19
+ $Y2=0
r98 44 46 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=4.355 $Y=0 $X2=4.56
+ $Y2=0
r99 43 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.885 $Y=0 $X2=5.05
+ $Y2=0
r100 43 46 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=4.885 $Y=0
+ $X2=4.56 $Y2=0
r101 42 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r102 42 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r103 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r104 39 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=0.71
+ $Y2=0
r105 39 41 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=1.2
+ $Y2=0
r106 38 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.405 $Y=0 $X2=1.57
+ $Y2=0
r107 38 41 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.405 $Y=0 $X2=1.2
+ $Y2=0
r108 36 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r109 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r110 33 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.71
+ $Y2=0
r111 33 35 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0
+ $X2=0.24 $Y2=0
r112 31 61 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=2.88 $Y=0 $X2=4.08
+ $Y2=0
r113 31 58 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=2.88 $Y=0 $X2=1.68
+ $Y2=0
r114 27 63 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.05 $Y=0.085
+ $X2=5.05 $Y2=0
r115 27 29 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=5.05 $Y=0.085
+ $X2=5.05 $Y2=0.595
r116 23 60 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.19 $Y=0.085
+ $X2=4.19 $Y2=0
r117 23 25 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=4.19 $Y=0.085
+ $X2=4.19 $Y2=0.595
r118 22 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.735 $Y=0 $X2=1.57
+ $Y2=0
r119 21 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.025 $Y=0 $X2=4.19
+ $Y2=0
r120 21 22 149.401 $w=1.68e-07 $l=2.29e-06 $layer=LI1_cond $X=4.025 $Y=0
+ $X2=1.735 $Y2=0
r121 17 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.57 $Y=0.085
+ $X2=1.57 $Y2=0
r122 17 19 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=1.57 $Y=0.085
+ $X2=1.57 $Y2=0.55
r123 13 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0
r124 13 15 18.6835 $w=3.28e-07 $l=5.35e-07 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0.62
r125 4 29 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=4.91
+ $Y=0.37 $X2=5.05 $Y2=0.595
r126 3 25 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=4.05
+ $Y=0.37 $X2=4.19 $Y2=0.595
r127 2 19 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=1.43 $Y=0.37
+ $X2=1.57 $Y2=0.55
r128 1 15 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.62
.ends

