# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_ls__nor3b_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.680000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.440000 1.220000 6.595000 1.550000 ;
        RECT 6.365000 1.180000 6.595000 1.220000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.350000 1.815000 1.780000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.363000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.765000 1.180000 7.095000 1.550000 ;
    END
  END C_N
  PIN Y
    ANTENNADIFFAREA  1.985500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.615000 0.350000 0.945000 1.010000 ;
        RECT 0.615000 1.010000 5.935000 1.050000 ;
        RECT 0.615000 1.050000 3.805000 1.150000 ;
        RECT 0.615000 1.150000 2.275000 1.180000 ;
        RECT 1.615000 0.350000 1.945000 0.980000 ;
        RECT 1.615000 0.980000 5.935000 1.010000 ;
        RECT 2.045000 1.180000 2.275000 1.820000 ;
        RECT 2.045000 1.820000 3.720000 2.070000 ;
        RECT 2.625000 0.350000 2.795000 0.980000 ;
        RECT 3.475000 0.350000 3.805000 0.880000 ;
        RECT 3.475000 0.880000 5.935000 0.980000 ;
        RECT 4.475000 0.350000 4.805000 0.880000 ;
        RECT 5.605000 0.350000 5.935000 0.880000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.680000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 7.680000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.680000 0.085000 ;
      RECT 0.000000  3.245000 7.680000 3.415000 ;
      RECT 0.115000  0.085000 0.445000 1.130000 ;
      RECT 0.115000  1.950000 0.445000 2.905000 ;
      RECT 0.115000  2.905000 2.370000 3.075000 ;
      RECT 0.615000  1.950000 1.870000 2.120000 ;
      RECT 0.615000  2.120000 0.945000 2.735000 ;
      RECT 1.115000  0.085000 1.445000 0.840000 ;
      RECT 1.145000  2.290000 1.315000 2.905000 ;
      RECT 1.525000  2.120000 1.870000 2.240000 ;
      RECT 1.525000  2.240000 5.100000 2.410000 ;
      RECT 1.525000  2.410000 1.855000 2.735000 ;
      RECT 2.040000  2.580000 4.170000 2.750000 ;
      RECT 2.040000  2.750000 2.370000 2.905000 ;
      RECT 2.115000  0.085000 2.445000 0.810000 ;
      RECT 2.580000  1.320000 4.195000 1.650000 ;
      RECT 2.940000  2.750000 3.270000 2.910000 ;
      RECT 2.975000  0.085000 3.305000 0.810000 ;
      RECT 3.840000  2.750000 4.170000 2.910000 ;
      RECT 3.890000  1.650000 4.195000 1.720000 ;
      RECT 3.890000  1.720000 7.565000 1.890000 ;
      RECT 3.975000  0.085000 4.305000 0.710000 ;
      RECT 4.400000  2.580000 4.730000 3.245000 ;
      RECT 4.795000  2.060000 6.080000 2.230000 ;
      RECT 4.795000  2.230000 5.100000 2.240000 ;
      RECT 4.930000  2.410000 5.100000 2.990000 ;
      RECT 4.975000  0.085000 5.435000 0.680000 ;
      RECT 5.300000  2.400000 5.630000 3.245000 ;
      RECT 5.810000  2.230000 6.080000 2.990000 ;
      RECT 6.105000  0.085000 6.435000 1.010000 ;
      RECT 6.250000  2.060000 6.580000 3.245000 ;
      RECT 6.605000  0.350000 7.565000 1.010000 ;
      RECT 6.785000  1.890000 7.055000 2.700000 ;
      RECT 7.235000  2.060000 7.565000 3.245000 ;
      RECT 7.395000  1.010000 7.565000 1.720000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
  END
END sky130_fd_sc_ls__nor3b_4
