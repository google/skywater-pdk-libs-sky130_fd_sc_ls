* NGSPICE file created from sky130_fd_sc_ls__ebufn_2.ext - technology: sky130A

.subckt sky130_fd_sc_ls__ebufn_2 A TE_B VGND VNB VPB VPWR Z
M1000 a_84_48# A VGND VNB nshort w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=4.797e+11p ps=4.17e+06u
M1001 VPWR TE_B a_33_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=1.0815e+12p pd=6.56e+06u as=1.0528e+12p ps=8.6e+06u
M1002 a_33_368# TE_B VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPWR TE_B a_283_48# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.95e+11p ps=2.59e+06u
M1004 VGND a_283_48# a_27_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=7.289e+11p ps=6.41e+06u
M1005 a_27_74# a_283_48# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_84_48# A VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.95e+11p pd=2.59e+06u as=0p ps=0u
M1007 Z a_84_48# a_27_74# VNB nshort w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1008 a_27_74# a_84_48# Z VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND TE_B a_283_48# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1010 a_33_368# a_84_48# Z VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.92e+11p ps=2.94e+06u
M1011 Z a_84_48# a_33_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

