* NGSPICE file created from sky130_fd_sc_ls__a311o_2.ext - technology: sky130A

.subckt sky130_fd_sc_ls__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
M1000 VPWR A2 a_330_392# VPB phighvt w=1e+06u l=150000u
+  ad=1.251e+12p pd=8.85e+06u as=6.6e+11p ps=5.32e+06u
M1001 a_423_74# A2 a_351_74# VNB nshort w=740000u l=150000u
+  ad=2.886e+11p pd=2.26e+06u as=1.554e+11p ps=1.9e+06u
M1002 a_21_270# C1 a_660_392# VPB phighvt w=1e+06u l=150000u
+  ad=2.75e+11p pd=2.55e+06u as=2.7e+11p ps=2.54e+06u
M1003 VGND a_21_270# X VNB nshort w=740000u l=150000u
+  ad=7.955e+11p pd=6.59e+06u as=2.072e+11p ps=2.04e+06u
M1004 VGND B1 a_21_270# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=4.847e+11p ps=4.27e+06u
M1005 a_660_392# B1 a_330_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_351_74# A3 VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR a_21_270# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.36e+11p ps=2.84e+06u
M1008 a_21_270# C1 VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 X a_21_270# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 X a_21_270# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_330_392# A1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_21_270# A1 a_423_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_330_392# A3 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

