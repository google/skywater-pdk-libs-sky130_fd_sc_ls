* File: sky130_fd_sc_ls__sdfstp_1.pex.spice
* Created: Fri Aug 28 14:04:15 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__SDFSTP_1%SCE 2 3 5 8 10 13 14 16 19 23 24 25 28 29
+ 33 36
c88 33 0 9.32299e-20 $X=0.72 $Y=1.665
c89 28 0 1.0138e-19 $X=1.955 $Y=1.425
c90 25 0 3.03849e-20 $X=1.79 $Y=1.525
c91 3 0 1.54286e-19 $X=0.5 $Y=2.245
r92 37 42 2.62366 $w=3.72e-07 $l=8e-08 $layer=LI1_cond $X=0.63 $Y=1.445 $X2=0.63
+ $Y2=1.525
r93 36 37 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.515
+ $Y=1.445 $X2=0.515 $Y2=1.445
r94 33 42 4.5914 $w=3.72e-07 $l=1.4e-07 $layer=LI1_cond $X=0.63 $Y=1.665
+ $X2=0.63 $Y2=1.525
r95 29 39 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.955 $Y=1.425
+ $X2=1.955 $Y2=1.26
r96 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.955
+ $Y=1.425 $X2=1.955 $Y2=1.425
r97 26 42 5.3395 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=0.835 $Y=1.525
+ $X2=0.63 $Y2=1.525
r98 25 28 4.51938 $w=2.53e-07 $l=1e-07 $layer=LI1_cond $X=1.917 $Y=1.525
+ $X2=1.917 $Y2=1.425
r99 25 26 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=1.79 $Y=1.525
+ $X2=0.835 $Y2=1.525
r100 23 36 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=0.515 $Y=1.8
+ $X2=0.515 $Y2=1.445
r101 23 24 12.8678 $w=2.55e-07 $l=7.5e-08 $layer=POLY_cond $X=0.515 $Y=1.8
+ $X2=0.515 $Y2=1.875
r102 22 36 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.515 $Y=1.28
+ $X2=0.515 $Y2=1.445
r103 19 39 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.935 $Y=0.58
+ $X2=1.935 $Y2=1.26
r104 14 16 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.95 $Y=2.245
+ $X2=0.95 $Y2=2.64
r105 13 14 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.95 $Y=2.155
+ $X2=0.95 $Y2=2.245
r106 12 13 79.6855 $w=1.8e-07 $l=2.05e-07 $layer=POLY_cond $X=0.95 $Y=1.95
+ $X2=0.95 $Y2=2.155
r107 11 24 13.0648 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.68 $Y=1.875
+ $X2=0.515 $Y2=1.875
r108 10 12 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=0.86 $Y=1.875
+ $X2=0.95 $Y2=1.95
r109 10 11 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=0.86 $Y=1.875
+ $X2=0.68 $Y2=1.875
r110 8 22 358.936 $w=1.5e-07 $l=7e-07 $layer=POLY_cond $X=0.575 $Y=0.58
+ $X2=0.575 $Y2=1.28
r111 3 5 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.5 $Y=2.245 $X2=0.5
+ $Y2=2.64
r112 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.5 $Y=2.155 $X2=0.5
+ $Y2=2.245
r113 1 24 12.8678 $w=2.55e-07 $l=8.21584e-08 $layer=POLY_cond $X=0.5 $Y=1.95
+ $X2=0.515 $Y2=1.875
r114 1 2 79.6855 $w=1.8e-07 $l=2.05e-07 $layer=POLY_cond $X=0.5 $Y=1.95 $X2=0.5
+ $Y2=2.155
.ends

.subckt PM_SKY130_FD_SC_LS__SDFSTP_1%A_27_464# 1 2 9 11 13 16 19 22 24 28 31 33
+ 34 38
c83 28 0 2.18476e-19 $X=1.955 $Y=1.995
c84 22 0 1.67103e-19 $X=1.79 $Y=2.405
c85 19 0 1.54286e-19 $X=0.17 $Y=2.3
c86 9 0 9.6166e-20 $X=1.115 $Y=0.58
r87 38 41 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.055 $Y=1.105
+ $X2=1.055 $Y2=0.94
r88 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.055
+ $Y=1.105 $X2=1.055 $Y2=1.105
r89 34 37 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=1.055 $Y=1.025
+ $X2=1.055 $Y2=1.105
r90 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.955
+ $Y=1.995 $X2=1.955 $Y2=1.995
r91 26 28 14.688 $w=2.53e-07 $l=3.25e-07 $layer=LI1_cond $X=1.917 $Y=2.32
+ $X2=1.917 $Y2=1.995
r92 25 31 3.51065 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=0.525 $Y=1.025
+ $X2=0.305 $Y2=1.025
r93 24 34 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.89 $Y=1.025
+ $X2=1.055 $Y2=1.025
r94 24 25 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.89 $Y=1.025
+ $X2=0.525 $Y2=1.025
r95 23 33 2.32734 $w=1.7e-07 $l=1.42913e-07 $layer=LI1_cond $X=0.36 $Y=2.405
+ $X2=0.222 $Y2=2.395
r96 22 26 7.17723 $w=1.7e-07 $l=1.64085e-07 $layer=LI1_cond $X=1.79 $Y=2.405
+ $X2=1.917 $Y2=2.32
r97 22 23 93.2941 $w=1.68e-07 $l=1.43e-06 $layer=LI1_cond $X=1.79 $Y=2.405
+ $X2=0.36 $Y2=2.405
r98 19 33 4.10697 $w=2.22e-07 $l=1.18174e-07 $layer=LI1_cond $X=0.17 $Y=2.3
+ $X2=0.222 $Y2=2.395
r99 18 31 3.10218 $w=3.05e-07 $l=1.72337e-07 $layer=LI1_cond $X=0.17 $Y=1.11
+ $X2=0.305 $Y2=1.025
r100 18 19 77.6364 $w=1.68e-07 $l=1.19e-06 $layer=LI1_cond $X=0.17 $Y=1.11
+ $X2=0.17 $Y2=2.3
r101 14 31 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.305 $Y=0.94
+ $X2=0.305 $Y2=1.025
r102 14 16 9.42908 $w=4.38e-07 $l=3.6e-07 $layer=LI1_cond $X=0.305 $Y=0.94
+ $X2=0.305 $Y2=0.58
r103 11 29 52.2586 $w=2.99e-07 $l=2.7157e-07 $layer=POLY_cond $X=2 $Y=2.245
+ $X2=1.955 $Y2=1.995
r104 11 13 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2 $Y=2.245 $X2=2
+ $Y2=2.64
r105 9 41 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=1.115 $Y=0.58
+ $X2=1.115 $Y2=0.94
r106 2 33 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.32 $X2=0.275 $Y2=2.465
r107 1 16 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.215
+ $Y=0.37 $X2=0.36 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_LS__SDFSTP_1%D 1 3 6 8 12
c36 1 0 1.37721e-19 $X=1.37 $Y=2.245
r37 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.415
+ $Y=1.985 $X2=1.415 $Y2=1.985
r38 8 12 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=1.2 $Y=1.985
+ $X2=1.415 $Y2=1.985
r39 4 11 38.5718 $w=2.96e-07 $l=2.05122e-07 $layer=POLY_cond $X=1.505 $Y=1.82
+ $X2=1.415 $Y2=1.985
r40 4 6 635.83 $w=1.5e-07 $l=1.24e-06 $layer=POLY_cond $X=1.505 $Y=1.82
+ $X2=1.505 $Y2=0.58
r41 1 11 54.0414 $w=2.96e-07 $l=2.81603e-07 $layer=POLY_cond $X=1.37 $Y=2.245
+ $X2=1.415 $Y2=1.985
r42 1 3 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.37 $Y=2.245
+ $X2=1.37 $Y2=2.64
.ends

.subckt PM_SKY130_FD_SC_LS__SDFSTP_1%SCD 1 3 4 6 7 8 9 10 14 16
c45 16 0 2.47679e-19 $X=2.68 $Y=1.985
c46 8 0 6.18088e-20 $X=2.64 $Y=1.295
c47 4 0 2.3928e-19 $X=2.42 $Y=2.245
r48 14 19 12.0163 $w=4.85e-07 $l=1.08185e-07 $layer=POLY_cond $X=2.602 $Y=1.382
+ $X2=2.677 $Y2=1.305
r49 14 16 66.5202 $w=4.85e-07 $l=6.03e-07 $layer=POLY_cond $X=2.602 $Y=1.382
+ $X2=2.602 $Y2=1.985
r50 10 16 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.68
+ $Y=1.985 $X2=2.68 $Y2=1.985
r51 9 10 14.7513 $w=2.48e-07 $l=3.2e-07 $layer=LI1_cond $X=2.68 $Y=1.665
+ $X2=2.68 $Y2=1.985
r52 8 9 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=2.68 $Y=1.295 $X2=2.68
+ $Y2=1.665
r53 8 19 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.68
+ $Y=1.305 $X2=2.68 $Y2=1.305
r54 7 16 1.65473 $w=4.85e-07 $l=1.5e-08 $layer=POLY_cond $X=2.602 $Y=2 $X2=2.602
+ $Y2=1.985
r55 4 7 30.6727 $w=3.85e-07 $l=3.23442e-07 $layer=POLY_cond $X=2.42 $Y=2.245
+ $X2=2.602 $Y2=2
r56 4 6 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.42 $Y=2.245
+ $X2=2.42 $Y2=2.64
r57 1 19 76.956 $w=3.4e-07 $l=5.85103e-07 $layer=POLY_cond $X=2.325 $Y=0.87
+ $X2=2.677 $Y2=1.305
r58 1 3 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.325 $Y=0.87
+ $X2=2.325 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_LS__SDFSTP_1%CLK 1 3 4 6 7
c34 4 0 6.18088e-20 $X=3.515 $Y=1.765
r35 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.44
+ $Y=1.385 $X2=3.44 $Y2=1.385
r36 7 11 4.98354 $w=3.68e-07 $l=1.6e-07 $layer=LI1_cond $X=3.6 $Y=1.365 $X2=3.44
+ $Y2=1.365
r37 4 10 77.2841 $w=2.7e-07 $l=4.15812e-07 $layer=POLY_cond $X=3.515 $Y=1.765
+ $X2=3.44 $Y2=1.385
r38 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.515 $Y=1.765
+ $X2=3.515 $Y2=2.4
r39 1 10 38.9026 $w=2.7e-07 $l=2.03101e-07 $layer=POLY_cond $X=3.355 $Y=1.22
+ $X2=3.44 $Y2=1.385
r40 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.355 $Y=1.22 $X2=3.355
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__SDFSTP_1%A_800_74# 1 2 7 9 14 16 18 20 21 23 26 30
+ 32 33 34 35 38 42 44 46 47 50 51 52 54 55 56 58 59 60 63 66 69 71 77 78 83
c252 78 0 1.57372e-19 $X=5.675 $Y=1.78
c253 55 0 1.72794e-19 $X=7.775 $Y=2.055
c254 21 0 1.54803e-19 $X=8.945 $Y=1.795
r255 72 83 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=8.835 $Y=1.285
+ $X2=8.945 $Y2=1.285
r256 72 80 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=8.835 $Y=1.285
+ $X2=8.745 $Y2=1.285
r257 71 73 18.3241 $w=2.53e-07 $l=3.8e-07 $layer=LI1_cond $X=8.835 $Y=1.285
+ $X2=8.835 $Y2=1.665
r258 71 72 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.835
+ $Y=1.285 $X2=8.835 $Y2=1.285
r259 67 78 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=5.615 $Y=1.78
+ $X2=5.675 $Y2=1.78
r260 67 77 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.615 $Y=1.78
+ $X2=5.45 $Y2=1.78
r261 66 68 6.4562 $w=2.74e-07 $l=1.45e-07 $layer=LI1_cond $X=5.615 $Y=1.78
+ $X2=5.76 $Y2=1.78
r262 66 67 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.615
+ $Y=1.78 $X2=5.615 $Y2=1.78
r263 59 73 3.06467 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.67 $Y=1.665
+ $X2=8.835 $Y2=1.665
r264 59 60 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=8.67 $Y=1.665
+ $X2=7.945 $Y2=1.665
r265 57 60 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.86 $Y=1.75
+ $X2=7.945 $Y2=1.665
r266 57 58 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=7.86 $Y=1.75
+ $X2=7.86 $Y2=1.97
r267 55 58 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.775 $Y=2.055
+ $X2=7.86 $Y2=1.97
r268 55 56 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=7.775 $Y=2.055
+ $X2=7.495 $Y2=2.055
r269 53 56 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.41 $Y=2.14
+ $X2=7.495 $Y2=2.055
r270 53 54 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=7.41 $Y=2.14
+ $X2=7.41 $Y2=2.895
r271 51 54 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.325 $Y=2.98
+ $X2=7.41 $Y2=2.895
r272 51 52 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=7.325 $Y=2.98
+ $X2=6.815 $Y2=2.98
r273 50 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.73 $Y=2.895
+ $X2=6.815 $Y2=2.98
r274 49 50 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=6.73 $Y=2.515
+ $X2=6.73 $Y2=2.895
r275 48 69 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.845 $Y=2.43
+ $X2=5.76 $Y2=2.43
r276 47 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.645 $Y=2.43
+ $X2=6.73 $Y2=2.515
r277 47 48 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=6.645 $Y=2.43
+ $X2=5.845 $Y2=2.43
r278 45 69 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.76 $Y=2.515
+ $X2=5.76 $Y2=2.43
r279 45 46 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=5.76 $Y=2.515
+ $X2=5.76 $Y2=2.895
r280 44 69 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.76 $Y=2.345
+ $X2=5.76 $Y2=2.43
r281 43 68 3.52985 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.76 $Y=1.945
+ $X2=5.76 $Y2=1.78
r282 43 44 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=5.76 $Y=1.945
+ $X2=5.76 $Y2=2.345
r283 42 63 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.12 $Y=0.935
+ $X2=5.12 $Y2=1.02
r284 41 42 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=5.12 $Y=0.425
+ $X2=5.12 $Y2=0.935
r285 39 75 16.1096 $w=3.74e-07 $l=1.25e-07 $layer=POLY_cond $X=4.947 $Y=1.565
+ $X2=4.947 $Y2=1.69
r286 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.905
+ $Y=1.565 $X2=4.905 $Y2=1.565
r287 36 63 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=4.895 $Y=1.02
+ $X2=5.12 $Y2=1.02
r288 36 38 24.0965 $w=2.18e-07 $l=4.6e-07 $layer=LI1_cond $X=4.895 $Y=1.105
+ $X2=4.895 $Y2=1.565
r289 34 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.675 $Y=2.98
+ $X2=5.76 $Y2=2.895
r290 34 35 91.3369 $w=1.68e-07 $l=1.4e-06 $layer=LI1_cond $X=5.675 $Y=2.98
+ $X2=4.275 $Y2=2.98
r291 32 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.035 $Y=0.34
+ $X2=5.12 $Y2=0.425
r292 32 33 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=5.035 $Y=0.34
+ $X2=4.225 $Y2=0.34
r293 28 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.19 $Y=2.895
+ $X2=4.275 $Y2=2.98
r294 28 30 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=4.19 $Y=2.895
+ $X2=4.19 $Y2=2.78
r295 24 33 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.1 $Y=0.425
+ $X2=4.225 $Y2=0.34
r296 24 26 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=4.1 $Y=0.425 $X2=4.1
+ $Y2=0.515
r297 21 23 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=8.945 $Y=1.795
+ $X2=8.945 $Y2=2.08
r298 20 21 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=8.945 $Y=1.705
+ $X2=8.945 $Y2=1.795
r299 19 83 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=8.945 $Y=1.45
+ $X2=8.945 $Y2=1.285
r300 19 20 99.121 $w=1.8e-07 $l=2.55e-07 $layer=POLY_cond $X=8.945 $Y=1.45
+ $X2=8.945 $Y2=1.705
r301 16 80 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.745 $Y=1.12
+ $X2=8.745 $Y2=1.285
r302 16 18 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=8.745 $Y=1.12
+ $X2=8.745 $Y2=0.69
r303 12 78 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.675 $Y=1.615
+ $X2=5.675 $Y2=1.78
r304 12 14 512.766 $w=1.5e-07 $l=1e-06 $layer=POLY_cond $X=5.675 $Y=1.615
+ $X2=5.675 $Y2=0.615
r305 11 75 24.2268 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=5.155 $Y=1.69
+ $X2=4.947 $Y2=1.69
r306 11 77 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=5.155 $Y=1.69
+ $X2=5.45 $Y2=1.69
r307 7 75 84.8702 $w=3.74e-07 $l=5.75986e-07 $layer=POLY_cond $X=5.065 $Y=2.21
+ $X2=4.947 $Y2=1.69
r308 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=5.065 $Y=2.21
+ $X2=5.065 $Y2=2.495
r309 2 30 600 $w=1.7e-07 $l=1.01223e-06 $layer=licon1_PDIFF $count=1 $X=4.04
+ $Y=1.84 $X2=4.19 $Y2=2.78
r310 1 26 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4 $Y=0.37
+ $X2=4.14 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__SDFSTP_1%A_1198_55# 1 2 7 9 10 12 14 15 17 21 24 29
+ 36 42
c93 24 0 3.56679e-19 $X=6.18 $Y=1.96
c94 17 0 3.34354e-20 $X=6.675 $Y=0.945
c95 10 0 1.82591e-19 $X=6.08 $Y=2.21
r96 36 38 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=6.84 $Y=0.8
+ $X2=6.84 $Y2=0.945
r97 33 42 16.6207 $w=2.61e-07 $l=9e-08 $layer=POLY_cond $X=6.36 $Y=1.1 $X2=6.27
+ $Y2=1.1
r98 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.36
+ $Y=1.1 $X2=6.36 $Y2=1.1
r99 29 32 7.44286 $w=2.38e-07 $l=1.55e-07 $layer=LI1_cond $X=6.36 $Y=0.945
+ $X2=6.36 $Y2=1.1
r100 24 27 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=6.18 $Y=1.96
+ $X2=6.18 $Y2=2.09
r101 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.18
+ $Y=1.96 $X2=6.18 $Y2=1.96
r102 19 21 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=7.07 $Y=2.175
+ $X2=7.07 $Y2=2.495
r103 18 29 2.75731 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=6.48 $Y=0.945
+ $X2=6.36 $Y2=0.945
r104 17 38 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.675 $Y=0.945
+ $X2=6.84 $Y2=0.945
r105 17 18 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=6.675 $Y=0.945
+ $X2=6.48 $Y2=0.945
r106 16 27 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.345 $Y=2.09
+ $X2=6.18 $Y2=2.09
r107 15 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.985 $Y=2.09
+ $X2=7.07 $Y2=2.175
r108 15 16 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=6.985 $Y=2.09
+ $X2=6.345 $Y2=2.09
r109 14 25 38.5462 $w=3.19e-07 $l=2.10286e-07 $layer=POLY_cond $X=6.27 $Y=1.795
+ $X2=6.167 $Y2=1.96
r110 13 42 15.717 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.27 $Y=1.265
+ $X2=6.27 $Y2=1.1
r111 13 14 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=6.27 $Y=1.265
+ $X2=6.27 $Y2=1.795
r112 10 25 51.3895 $w=3.19e-07 $l=2.90259e-07 $layer=POLY_cond $X=6.08 $Y=2.21
+ $X2=6.167 $Y2=1.96
r113 10 12 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.08 $Y=2.21
+ $X2=6.08 $Y2=2.495
r114 7 42 37.8582 $w=2.61e-07 $l=2.75409e-07 $layer=POLY_cond $X=6.065 $Y=0.935
+ $X2=6.27 $Y2=1.1
r115 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.065 $Y=0.935
+ $X2=6.065 $Y2=0.615
r116 2 21 600 $w=1.7e-07 $l=2.86182e-07 $layer=licon1_PDIFF $count=1 $X=6.89
+ $Y=2.285 $X2=7.07 $Y2=2.495
r117 1 36 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=6.695
+ $Y=0.59 $X2=6.84 $Y2=0.8
.ends

.subckt PM_SKY130_FD_SC_LS__SDFSTP_1%A_998_81# 1 2 8 9 11 14 16 17 19 20 22 25
+ 31 33 34 35 39 41 42 48 49 51 55 60 62 64
c169 60 0 1.55656e-19 $X=6.77 $Y=1.67
c170 48 0 1.82591e-19 $X=5.34 $Y=2.495
c171 39 0 1.72794e-19 $X=7.905 $Y=1.265
c172 14 0 3.34354e-20 $X=7.055 $Y=1.09
c173 9 0 4.36509e-20 $X=6.815 $Y=2.21
r174 60 65 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.77 $Y=1.67
+ $X2=6.77 $Y2=1.835
r175 60 64 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.77 $Y=1.67
+ $X2=6.77 $Y2=1.505
r176 59 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.77
+ $Y=1.67 $X2=6.77 $Y2=1.67
r177 51 53 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=5.985 $Y=1.36
+ $X2=5.985 $Y2=1.52
r178 48 49 10.7321 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=5.34 $Y=2.495
+ $X2=5.34 $Y2=2.265
r179 42 68 11.4762 $w=3.78e-07 $l=9e-08 $layer=POLY_cond $X=8.265 $Y=1.375
+ $X2=8.355 $Y2=1.375
r180 42 66 36.9788 $w=3.78e-07 $l=2.9e-07 $layer=POLY_cond $X=8.265 $Y=1.375
+ $X2=7.975 $Y2=1.375
r181 41 42 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.265
+ $Y=1.285 $X2=8.265 $Y2=1.285
r182 39 62 6.93634 $w=2.88e-07 $l=1.45e-07 $layer=LI1_cond $X=7.905 $Y=1.265
+ $X2=7.76 $Y2=1.265
r183 39 41 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=7.905 $Y=1.265
+ $X2=8.265 $Y2=1.265
r184 38 55 3.76007 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=6.935 $Y=1.285
+ $X2=6.792 $Y2=1.285
r185 38 62 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=6.935 $Y=1.285
+ $X2=7.76 $Y2=1.285
r186 36 53 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.07 $Y=1.52
+ $X2=5.985 $Y2=1.52
r187 35 59 6.06549 $w=2.83e-07 $l=1.5e-07 $layer=LI1_cond $X=6.792 $Y=1.52
+ $X2=6.792 $Y2=1.67
r188 35 55 9.5026 $w=2.83e-07 $l=2.35e-07 $layer=LI1_cond $X=6.792 $Y=1.52
+ $X2=6.792 $Y2=1.285
r189 35 36 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=6.65 $Y=1.52
+ $X2=6.07 $Y2=1.52
r190 33 51 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.9 $Y=1.36
+ $X2=5.985 $Y2=1.36
r191 33 34 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=5.9 $Y=1.36
+ $X2=5.625 $Y2=1.36
r192 29 34 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=5.5 $Y=1.36
+ $X2=5.625 $Y2=1.36
r193 29 44 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=5.5 $Y=1.36
+ $X2=5.26 $Y2=1.36
r194 29 31 30.4245 $w=2.48e-07 $l=6.6e-07 $layer=LI1_cond $X=5.5 $Y=1.275
+ $X2=5.5 $Y2=0.615
r195 27 44 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.26 $Y=1.445
+ $X2=5.26 $Y2=1.36
r196 27 49 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=5.26 $Y=1.445
+ $X2=5.26 $Y2=2.265
r197 23 25 115.372 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=6.83 $Y=1.165
+ $X2=7.055 $Y2=1.165
r198 20 68 24.4846 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=8.355 $Y=1.12
+ $X2=8.355 $Y2=1.375
r199 20 22 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=8.355 $Y=1.12
+ $X2=8.355 $Y2=0.69
r200 17 66 24.4846 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=7.975 $Y=1.63
+ $X2=7.975 $Y2=1.375
r201 17 19 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=7.975 $Y=1.63
+ $X2=7.975 $Y2=2.205
r202 14 25 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.055 $Y=1.09
+ $X2=7.055 $Y2=1.165
r203 14 16 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=7.055 $Y=1.09
+ $X2=7.055 $Y2=0.8
r204 12 23 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.83 $Y=1.24
+ $X2=6.83 $Y2=1.165
r205 12 64 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=6.83 $Y=1.24
+ $X2=6.83 $Y2=1.505
r206 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.815 $Y=2.21
+ $X2=6.815 $Y2=2.495
r207 8 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.815 $Y=2.12 $X2=6.815
+ $Y2=2.21
r208 8 65 110.782 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=6.815 $Y=2.12
+ $X2=6.815 $Y2=1.835
r209 2 48 600 $w=1.7e-07 $l=2.93428e-07 $layer=licon1_PDIFF $count=1 $X=5.14
+ $Y=2.285 $X2=5.34 $Y2=2.495
r210 1 31 182 $w=1.7e-07 $l=5.65332e-07 $layer=licon1_NDIFF $count=1 $X=4.99
+ $Y=0.405 $X2=5.46 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_LS__SDFSTP_1%SET_B 2 3 5 8 12 15 16 18 21 22 23 24 29 32
+ 35 36 43
r139 35 38 39.5669 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=7.332 $Y=1.67
+ $X2=7.332 $Y2=1.835
r140 35 37 48.8634 $w=3.75e-07 $l=1.9e-07 $layer=POLY_cond $X=7.332 $Y=1.67
+ $X2=7.332 $Y2=1.48
r141 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.31
+ $Y=1.67 $X2=7.31 $Y2=1.67
r142 32 43 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=10.865
+ $Y=1.545 $X2=10.865 $Y2=1.545
r143 29 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=1.665
+ $X2=10.8 $Y2=1.665
r144 26 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=1.665
+ $X2=7.44 $Y2=1.665
r145 24 26 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.585 $Y=1.665
+ $X2=7.44 $Y2=1.665
r146 23 29 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=10.655 $Y=1.665
+ $X2=10.8 $Y2=1.665
r147 23 24 3.7995 $w=1.4e-07 $l=3.07e-06 $layer=MET1_cond $X=10.655 $Y=1.665
+ $X2=7.585 $Y2=1.665
r148 21 32 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=10.865 $Y=1.885
+ $X2=10.865 $Y2=1.545
r149 21 22 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.865 $Y=1.885
+ $X2=10.865 $Y2=2.05
r150 20 32 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.865 $Y=1.38
+ $X2=10.865 $Y2=1.545
r151 16 18 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=10.94 $Y=2.465
+ $X2=10.94 $Y2=2.75
r152 15 16 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=10.94 $Y=2.375
+ $X2=10.94 $Y2=2.465
r153 15 22 126.331 $w=1.8e-07 $l=3.25e-07 $layer=POLY_cond $X=10.94 $Y=2.375
+ $X2=10.94 $Y2=2.05
r154 12 20 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=10.775 $Y=0.58
+ $X2=10.775 $Y2=1.38
r155 8 37 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=7.445 $Y=0.8
+ $X2=7.445 $Y2=1.48
r156 3 5 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.295 $Y=2.21
+ $X2=7.295 $Y2=2.495
r157 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=7.295 $Y=2.12 $X2=7.295
+ $Y2=2.21
r158 2 38 110.782 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=7.295 $Y=2.12
+ $X2=7.295 $Y2=1.835
.ends

.subckt PM_SKY130_FD_SC_LS__SDFSTP_1%A_599_74# 1 2 9 11 13 15 16 17 19 20 21 22
+ 23 26 28 29 30 32 33 37 39 40 44 47 49 51 52 56 59 60 61 66 69
c190 51 0 1.92727e-19 $X=9.497 $Y=1.795
c191 30 0 1.34962e-19 $X=5.565 $Y=2.78
r192 70 71 5.58841 $w=3.45e-07 $l=4e-08 $layer=POLY_cond $X=3.925 $Y=1.557
+ $X2=3.965 $Y2=1.557
r193 67 71 11.8754 $w=3.45e-07 $l=8.5e-08 $layer=POLY_cond $X=4.05 $Y=1.557
+ $X2=3.965 $Y2=1.557
r194 66 67 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.05
+ $Y=1.515 $X2=4.05 $Y2=1.515
r195 64 66 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=4.05 $Y=1.82
+ $X2=4.05 $Y2=1.515
r196 61 63 6.68417 $w=2.48e-07 $l=1.45e-07 $layer=LI1_cond $X=3.145 $Y=1.945
+ $X2=3.29 $Y2=1.945
r197 60 64 6.98653 $w=2.5e-07 $l=2.18746e-07 $layer=LI1_cond $X=3.885 $Y=1.945
+ $X2=4.05 $Y2=1.82
r198 60 63 27.4281 $w=2.48e-07 $l=5.95e-07 $layer=LI1_cond $X=3.885 $Y=1.945
+ $X2=3.29 $Y2=1.945
r199 59 61 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.06 $Y=1.82
+ $X2=3.145 $Y2=1.945
r200 59 69 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=3.06 $Y=1.82
+ $X2=3.06 $Y2=1.01
r201 54 69 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.14 $Y=0.845
+ $X2=3.14 $Y2=1.01
r202 54 56 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=3.14 $Y=0.845
+ $X2=3.14 $Y2=0.515
r203 45 47 46.1489 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.455 $Y=2.385
+ $X2=4.545 $Y2=2.385
r204 44 51 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=9.505 $Y=2.37
+ $X2=9.505 $Y2=1.795
r205 42 52 81.8353 $w=1.8e-07 $l=2.05e-07 $layer=POLY_cond $X=9.505 $Y=2.945
+ $X2=9.505 $Y2=3.15
r206 42 44 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=9.505 $Y=2.945
+ $X2=9.505 $Y2=2.37
r207 40 51 35.2692 $w=1.95e-07 $l=9.7e-08 $layer=POLY_cond $X=9.497 $Y=1.698
+ $X2=9.497 $Y2=1.795
r208 39 50 36.6888 $w=1.95e-07 $l=9.7e-08 $layer=POLY_cond $X=9.497 $Y=1.507
+ $X2=9.497 $Y2=1.41
r209 39 40 64.9551 $w=1.95e-07 $l=1.91e-07 $layer=POLY_cond $X=9.497 $Y=1.507
+ $X2=9.497 $Y2=1.698
r210 37 50 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=9.475 $Y=0.58
+ $X2=9.475 $Y2=1.41
r211 34 49 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=5.655 $Y=3.15
+ $X2=5.565 $Y2=3.15
r212 33 52 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=9.415 $Y=3.15
+ $X2=9.505 $Y2=3.15
r213 33 34 1928 $w=1.5e-07 $l=3.76e-06 $layer=POLY_cond $X=9.415 $Y=3.15
+ $X2=5.655 $Y2=3.15
r214 30 32 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=5.565 $Y=2.78
+ $X2=5.565 $Y2=2.495
r215 29 49 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=5.565 $Y=3.075
+ $X2=5.565 $Y2=3.15
r216 28 30 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.565 $Y=2.87
+ $X2=5.565 $Y2=2.78
r217 28 29 79.6855 $w=1.8e-07 $l=2.05e-07 $layer=POLY_cond $X=5.565 $Y=2.87
+ $X2=5.565 $Y2=3.075
r218 24 26 217.926 $w=1.5e-07 $l=4.25e-07 $layer=POLY_cond $X=4.915 $Y=1.04
+ $X2=4.915 $Y2=0.615
r219 22 49 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=5.475 $Y=3.15
+ $X2=5.565 $Y2=3.15
r220 22 23 438.415 $w=1.5e-07 $l=8.55e-07 $layer=POLY_cond $X=5.475 $Y=3.15
+ $X2=4.62 $Y2=3.15
r221 20 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.84 $Y=1.115
+ $X2=4.915 $Y2=1.04
r222 20 21 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=4.84 $Y=1.115
+ $X2=4.53 $Y2=1.115
r223 19 23 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.545 $Y=3.075
+ $X2=4.62 $Y2=3.15
r224 18 47 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.545 $Y=2.46
+ $X2=4.545 $Y2=2.385
r225 18 19 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=4.545 $Y=2.46
+ $X2=4.545 $Y2=3.075
r226 17 45 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.455 $Y=2.31
+ $X2=4.455 $Y2=2.385
r227 16 67 56.5826 $w=3.45e-07 $l=4.05e-07 $layer=POLY_cond $X=4.455 $Y=1.557
+ $X2=4.05 $Y2=1.557
r228 16 17 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=4.455 $Y=1.68
+ $X2=4.455 $Y2=2.31
r229 15 16 22.2839 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.455 $Y=1.35
+ $X2=4.455 $Y2=1.557
r230 14 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.455 $Y=1.19
+ $X2=4.53 $Y2=1.115
r231 14 15 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=4.455 $Y=1.19
+ $X2=4.455 $Y2=1.35
r232 11 71 22.2839 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.965 $Y=1.765
+ $X2=3.965 $Y2=1.557
r233 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.965 $Y=1.765
+ $X2=3.965 $Y2=2.4
r234 7 70 22.2839 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.925 $Y=1.35
+ $X2=3.925 $Y2=1.557
r235 7 9 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.925 $Y=1.35
+ $X2=3.925 $Y2=0.74
r236 2 63 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=3.145
+ $Y=1.84 $X2=3.29 $Y2=1.985
r237 1 56 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=2.995
+ $Y=0.37 $X2=3.14 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__SDFSTP_1%A_1958_48# 1 2 7 9 11 12 14 15 19 23 27 32
+ 34 35 36 37 41
r96 36 37 8.63679 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=11.74 $Y=2.22
+ $X2=11.74 $Y2=2.39
r97 33 41 11.2481 $w=4.45e-07 $l=9e-08 $layer=POLY_cond $X=10.295 $Y=1.087
+ $X2=10.385 $Y2=1.087
r98 32 34 6.83261 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=10.295 $Y=1.145
+ $X2=10.46 $Y2=1.145
r99 32 33 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=10.295
+ $Y=1.145 $X2=10.295 $Y2=1.145
r100 29 35 4.47619 $w=2.72e-07 $l=5.63383e-07 $layer=LI1_cond $X=11.855 $Y=1.21
+ $X2=11.395 $Y2=0.98
r101 29 36 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=11.855 $Y=1.21
+ $X2=11.855 $Y2=2.22
r102 27 37 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=11.705 $Y=2.75
+ $X2=11.705 $Y2=2.39
r103 21 35 4.47619 $w=2.72e-07 $l=1.87e-07 $layer=LI1_cond $X=11.582 $Y=0.98
+ $X2=11.395 $Y2=0.98
r104 21 23 12.2927 $w=3.73e-07 $l=4e-07 $layer=LI1_cond $X=11.582 $Y=0.98
+ $X2=11.582 $Y2=0.58
r105 19 35 1.95968 $w=2.3e-07 $l=1.15e-07 $layer=LI1_cond $X=11.395 $Y=1.095
+ $X2=11.395 $Y2=0.98
r106 19 34 46.8493 $w=2.28e-07 $l=9.35e-07 $layer=LI1_cond $X=11.395 $Y=1.095
+ $X2=10.46 $Y2=1.095
r107 15 16 30.488 $w=1.66e-07 $l=1.05e-07 $layer=POLY_cond $X=10.385 $Y=2.377
+ $X2=10.49 $Y2=2.377
r108 12 16 5.24352 $w=1.5e-07 $l=8.8e-08 $layer=POLY_cond $X=10.49 $Y=2.465
+ $X2=10.49 $Y2=2.377
r109 12 14 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=10.49 $Y=2.465
+ $X2=10.49 $Y2=2.75
r110 11 15 5.24352 $w=1.5e-07 $l=8.7e-08 $layer=POLY_cond $X=10.385 $Y=2.29
+ $X2=10.385 $Y2=2.377
r111 10 41 28.4889 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=10.385 $Y=1.31
+ $X2=10.385 $Y2=1.087
r112 10 11 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=10.385 $Y=1.31
+ $X2=10.385 $Y2=2.29
r113 7 33 53.7407 $w=4.45e-07 $l=4.3e-07 $layer=POLY_cond $X=9.865 $Y=1.087
+ $X2=10.295 $Y2=1.087
r114 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=9.865 $Y=0.865
+ $X2=9.865 $Y2=0.58
r115 2 27 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=11.57
+ $Y=2.54 $X2=11.705 $Y2=2.75
r116 1 23 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=11.42
+ $Y=0.37 $X2=11.56 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_LS__SDFSTP_1%A_1764_74# 1 2 3 12 14 15 16 18 21 25 27 29
+ 32 33 34 36 40 43 44 47 48 49 52 56 57 60 62 65 66 67
c155 47 0 7.36644e-20 $X=10.15 $Y=2.22
c156 40 0 1.19062e-19 $X=9.275 $Y=2.015
r157 62 64 15.4168 $w=5.68e-07 $l=4.25e-07 $layer=LI1_cond $X=9.08 $Y=0.515
+ $X2=9.08 $Y2=0.94
r158 60 66 3.46198 $w=2.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=11.285 $Y=2.22
+ $X2=11.185 $Y2=2.305
r159 60 67 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=11.285 $Y=2.22
+ $X2=11.285 $Y2=2.05
r160 56 57 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=11.435
+ $Y=1.545 $X2=11.435 $Y2=1.545
r161 54 67 9.656 $w=3.98e-07 $l=2e-07 $layer=LI1_cond $X=11.4 $Y=1.85 $X2=11.4
+ $Y2=2.05
r162 54 56 8.78738 $w=3.98e-07 $l=3.05e-07 $layer=LI1_cond $X=11.4 $Y=1.85
+ $X2=11.4 $Y2=1.545
r163 50 66 3.46198 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.185 $Y=2.39
+ $X2=11.185 $Y2=2.305
r164 50 52 11.213 $w=3.68e-07 $l=3.6e-07 $layer=LI1_cond $X=11.185 $Y=2.39
+ $X2=11.185 $Y2=2.75
r165 48 66 3.05049 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=11 $Y=2.305
+ $X2=11.185 $Y2=2.305
r166 48 49 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=11 $Y=2.305
+ $X2=10.235 $Y2=2.305
r167 47 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.15 $Y=2.22
+ $X2=10.235 $Y2=2.305
r168 46 47 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=10.15 $Y=1.79
+ $X2=10.15 $Y2=2.22
r169 45 65 2.32734 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=9.365 $Y=1.705
+ $X2=9.227 $Y2=1.705
r170 44 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.065 $Y=1.705
+ $X2=10.15 $Y2=1.79
r171 44 45 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=10.065 $Y=1.705
+ $X2=9.365 $Y2=1.705
r172 43 65 4.10697 $w=2.22e-07 $l=1.08305e-07 $layer=LI1_cond $X=9.28 $Y=1.62
+ $X2=9.227 $Y2=1.705
r173 43 64 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=9.28 $Y=1.62
+ $X2=9.28 $Y2=0.94
r174 38 65 4.10697 $w=2.22e-07 $l=8.5e-08 $layer=LI1_cond $X=9.227 $Y=1.79
+ $X2=9.227 $Y2=1.705
r175 38 40 9.42908 $w=2.73e-07 $l=2.25e-07 $layer=LI1_cond $X=9.227 $Y=1.79
+ $X2=9.227 $Y2=2.015
r176 35 36 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=12.75 $Y=1.865
+ $X2=12.92 $Y2=1.865
r177 32 57 42.841 $w=3.3e-07 $l=2.45e-07 $layer=POLY_cond $X=11.435 $Y=1.79
+ $X2=11.435 $Y2=1.545
r178 31 57 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=11.435 $Y=1.38
+ $X2=11.435 $Y2=1.545
r179 27 36 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.92 $Y=1.94
+ $X2=12.92 $Y2=1.865
r180 27 29 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=12.92 $Y=1.94
+ $X2=12.92 $Y2=2.435
r181 23 35 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.75 $Y=1.79
+ $X2=12.75 $Y2=1.865
r182 23 25 489.691 $w=1.5e-07 $l=9.55e-07 $layer=POLY_cond $X=12.75 $Y=1.79
+ $X2=12.75 $Y2=0.835
r183 22 34 15.6241 $w=2.05e-07 $l=9.87421e-08 $layer=POLY_cond $X=12.02 $Y=1.865
+ $X2=11.945 $Y2=1.92
r184 21 35 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.675 $Y=1.865
+ $X2=12.75 $Y2=1.865
r185 21 22 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=12.675 $Y=1.865
+ $X2=12.02 $Y2=1.865
r186 19 34 9.82985 $w=1.5e-07 $l=1.3e-07 $layer=POLY_cond $X=11.945 $Y=2.05
+ $X2=11.945 $Y2=1.92
r187 19 33 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=11.945 $Y=2.05
+ $X2=11.945 $Y2=2.29
r188 16 33 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=11.93 $Y=2.465
+ $X2=11.93 $Y2=2.29
r189 16 18 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=11.93 $Y=2.465
+ $X2=11.93 $Y2=2.75
r190 15 32 27.4267 $w=2.6e-07 $l=2.20624e-07 $layer=POLY_cond $X=11.6 $Y=1.92
+ $X2=11.435 $Y2=1.79
r191 14 34 15.6241 $w=2.05e-07 $l=7.5e-08 $layer=POLY_cond $X=11.87 $Y=1.92
+ $X2=11.945 $Y2=1.92
r192 14 15 64.5024 $w=2.6e-07 $l=2.7e-07 $layer=POLY_cond $X=11.87 $Y=1.92
+ $X2=11.6 $Y2=1.92
r193 12 31 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=11.345 $Y=0.58
+ $X2=11.345 $Y2=1.38
r194 3 52 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=11.015
+ $Y=2.54 $X2=11.165 $Y2=2.75
r195 2 40 600 $w=1.7e-07 $l=3.19374e-07 $layer=licon1_PDIFF $count=1 $X=9.02
+ $Y=1.87 $X2=9.275 $Y2=2.015
r196 1 62 91 $w=1.7e-07 $l=3.14245e-07 $layer=licon1_NDIFF $count=2 $X=8.82
+ $Y=0.37 $X2=9.07 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__SDFSTP_1%A_2395_112# 1 2 7 9 10 12 18 23 27 32 33 35
+ 36
r62 31 33 2.05777 $w=4.63e-07 $l=8e-08 $layer=LI1_cond $X=12.535 $Y=0.772
+ $X2=12.615 $Y2=0.772
r63 31 32 5.26869 $w=4.63e-07 $l=1.65e-07 $layer=LI1_cond $X=12.535 $Y=0.772
+ $X2=12.37 $Y2=0.772
r64 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.23
+ $Y=1.385 $X2=13.23 $Y2=1.385
r65 25 35 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.7 $Y=1.385
+ $X2=12.615 $Y2=1.385
r66 25 27 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=12.7 $Y=1.385
+ $X2=13.23 $Y2=1.385
r67 23 36 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=12.695 $Y=2.16
+ $X2=12.695 $Y2=1.995
r68 19 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.615 $Y=1.55
+ $X2=12.615 $Y2=1.385
r69 19 36 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=12.615 $Y=1.55
+ $X2=12.615 $Y2=1.995
r70 18 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.615 $Y=1.22
+ $X2=12.615 $Y2=1.385
r71 17 33 6.7035 $w=1.7e-07 $l=2.33e-07 $layer=LI1_cond $X=12.615 $Y=1.005
+ $X2=12.615 $Y2=0.772
r72 17 18 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=12.615 $Y=1.005
+ $X2=12.615 $Y2=1.22
r73 15 32 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=12.12 $Y=0.705
+ $X2=12.37 $Y2=0.705
r74 10 28 68.9212 $w=3.43e-07 $l=4.4238e-07 $layer=POLY_cond $X=13.425 $Y=1.765
+ $X2=13.29 $Y2=1.385
r75 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=13.425 $Y=1.765
+ $X2=13.425 $Y2=2.4
r76 7 28 38.7084 $w=3.43e-07 $l=1.83916e-07 $layer=POLY_cond $X=13.33 $Y=1.22
+ $X2=13.29 $Y2=1.385
r77 7 9 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=13.33 $Y=1.22 $X2=13.33
+ $Y2=0.74
r78 2 23 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=12.56
+ $Y=2.015 $X2=12.695 $Y2=2.16
r79 1 31 182 $w=1.7e-07 $l=6.85857e-07 $layer=licon1_NDIFF $count=1 $X=11.975
+ $Y=0.56 $X2=12.535 $Y2=0.84
r80 1 15 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=11.975
+ $Y=0.56 $X2=12.12 $Y2=0.705
.ends

.subckt PM_SKY130_FD_SC_LS__SDFSTP_1%VPWR 1 2 3 4 5 6 7 8 27 31 33 37 41 45 49
+ 53 57 60 61 63 64 66 67 69 70 71 73 78 108 114 115 118 121 124 127
r161 127 128 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=3.33
+ $X2=13.2 $Y2=3.33
r162 124 125 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r163 122 125 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r164 121 122 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r165 118 119 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r166 115 128 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=3.33
+ $X2=13.2 $Y2=3.33
r167 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=3.33
+ $X2=13.68 $Y2=3.33
r168 112 127 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.36 $Y=3.33
+ $X2=13.195 $Y2=3.33
r169 112 114 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=13.36 $Y=3.33
+ $X2=13.68 $Y2=3.33
r170 111 128 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=13.2 $Y2=3.33
r171 110 111 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r172 108 127 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.03 $Y=3.33
+ $X2=13.195 $Y2=3.33
r173 108 110 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=13.03 $Y=3.33
+ $X2=12.72 $Y2=3.33
r174 107 111 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=12.72 $Y2=3.33
r175 106 107 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r176 104 107 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=11.76 $Y2=3.33
r177 103 106 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=10.8 $Y=3.33
+ $X2=11.76 $Y2=3.33
r178 103 104 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r179 101 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=10.8 $Y2=3.33
r180 100 101 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r181 98 101 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=10.32 $Y2=3.33
r182 97 100 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=7.92 $Y=3.33
+ $X2=10.32 $Y2=3.33
r183 97 98 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r184 95 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r185 94 95 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r186 91 94 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=6.48 $Y=3.33
+ $X2=7.44 $Y2=3.33
r187 91 92 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r188 89 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r189 88 89 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r190 86 89 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=6 $Y2=3.33
r191 86 125 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r192 85 88 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.08 $Y=3.33 $X2=6
+ $Y2=3.33
r193 85 86 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r194 83 124 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.905 $Y=3.33
+ $X2=3.74 $Y2=3.33
r195 83 85 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.905 $Y=3.33
+ $X2=4.08 $Y2=3.33
r196 82 122 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r197 82 119 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r198 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r199 79 118 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.89 $Y=3.33
+ $X2=0.725 $Y2=3.33
r200 79 81 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.89 $Y=3.33
+ $X2=1.2 $Y2=3.33
r201 78 121 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.565 $Y=3.33
+ $X2=2.73 $Y2=3.33
r202 78 81 89.0535 $w=1.68e-07 $l=1.365e-06 $layer=LI1_cond $X=2.565 $Y=3.33
+ $X2=1.2 $Y2=3.33
r203 76 119 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r204 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r205 73 118 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.56 $Y=3.33
+ $X2=0.725 $Y2=3.33
r206 73 75 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.56 $Y=3.33
+ $X2=0.24 $Y2=3.33
r207 71 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.44 $Y2=3.33
r208 71 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6.48 $Y2=3.33
r209 69 106 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=12.07 $Y=3.33
+ $X2=11.76 $Y2=3.33
r210 69 70 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.07 $Y=3.33
+ $X2=12.195 $Y2=3.33
r211 68 110 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=12.32 $Y=3.33
+ $X2=12.72 $Y2=3.33
r212 68 70 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.32 $Y=3.33
+ $X2=12.195 $Y2=3.33
r213 67 103 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.715 $Y=3.33
+ $X2=10.8 $Y2=3.33
r214 66 100 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=10.63 $Y=3.33
+ $X2=10.32 $Y2=3.33
r215 66 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.63 $Y=3.33
+ $X2=10.715 $Y2=3.33
r216 63 94 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=7.665 $Y=3.33
+ $X2=7.44 $Y2=3.33
r217 63 64 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.665 $Y=3.33
+ $X2=7.79 $Y2=3.33
r218 62 97 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=7.915 $Y=3.33
+ $X2=7.92 $Y2=3.33
r219 62 64 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.915 $Y=3.33
+ $X2=7.79 $Y2=3.33
r220 60 88 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=6.225 $Y=3.33
+ $X2=6 $Y2=3.33
r221 60 61 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.225 $Y=3.33
+ $X2=6.35 $Y2=3.33
r222 59 91 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=6.475 $Y=3.33
+ $X2=6.48 $Y2=3.33
r223 59 61 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.475 $Y=3.33
+ $X2=6.35 $Y2=3.33
r224 55 127 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.195 $Y=3.245
+ $X2=13.195 $Y2=3.33
r225 55 57 37.8909 $w=3.28e-07 $l=1.085e-06 $layer=LI1_cond $X=13.195 $Y=3.245
+ $X2=13.195 $Y2=2.16
r226 51 70 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=12.195 $Y=3.245
+ $X2=12.195 $Y2=3.33
r227 51 53 21.8964 $w=2.48e-07 $l=4.75e-07 $layer=LI1_cond $X=12.195 $Y=3.245
+ $X2=12.195 $Y2=2.77
r228 47 67 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.715 $Y=3.245
+ $X2=10.715 $Y2=3.33
r229 47 49 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=10.715 $Y=3.245
+ $X2=10.715 $Y2=2.77
r230 43 64 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.79 $Y=3.245
+ $X2=7.79 $Y2=3.33
r231 43 45 33.6513 $w=2.48e-07 $l=7.3e-07 $layer=LI1_cond $X=7.79 $Y=3.245
+ $X2=7.79 $Y2=2.515
r232 39 61 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.35 $Y=3.245
+ $X2=6.35 $Y2=3.33
r233 39 41 18.2086 $w=2.48e-07 $l=3.95e-07 $layer=LI1_cond $X=6.35 $Y=3.245
+ $X2=6.35 $Y2=2.85
r234 35 124 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.74 $Y=3.245
+ $X2=3.74 $Y2=3.33
r235 35 37 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=3.74 $Y=3.245
+ $X2=3.74 $Y2=2.78
r236 34 121 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.895 $Y=3.33
+ $X2=2.73 $Y2=3.33
r237 33 124 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.575 $Y=3.33
+ $X2=3.74 $Y2=3.33
r238 33 34 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.575 $Y=3.33
+ $X2=2.895 $Y2=3.33
r239 29 121 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.73 $Y=3.245
+ $X2=2.73 $Y2=3.33
r240 29 31 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=2.73 $Y=3.245
+ $X2=2.73 $Y2=2.995
r241 25 118 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.725 $Y=3.245
+ $X2=0.725 $Y2=3.33
r242 25 27 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=0.725 $Y=3.245
+ $X2=0.725 $Y2=2.78
r243 8 57 300 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=2 $X=12.995
+ $Y=2.015 $X2=13.195 $Y2=2.16
r244 7 53 600 $w=1.7e-07 $l=2.95635e-07 $layer=licon1_PDIFF $count=1 $X=12.005
+ $Y=2.54 $X2=12.155 $Y2=2.77
r245 6 49 600 $w=1.7e-07 $l=2.95635e-07 $layer=licon1_PDIFF $count=1 $X=10.565
+ $Y=2.54 $X2=10.715 $Y2=2.77
r246 5 45 600 $w=1.7e-07 $l=4.81456e-07 $layer=licon1_PDIFF $count=1 $X=7.37
+ $Y=2.285 $X2=7.75 $Y2=2.515
r247 4 41 600 $w=1.7e-07 $l=6.72309e-07 $layer=licon1_PDIFF $count=1 $X=6.155
+ $Y=2.285 $X2=6.39 $Y2=2.85
r248 3 37 600 $w=1.7e-07 $l=1.01223e-06 $layer=licon1_PDIFF $count=1 $X=3.59
+ $Y=1.84 $X2=3.74 $Y2=2.78
r249 2 31 600 $w=1.7e-07 $l=7.83741e-07 $layer=licon1_PDIFF $count=1 $X=2.495
+ $Y=2.32 $X2=2.73 $Y2=2.995
r250 1 27 600 $w=1.7e-07 $l=5.29717e-07 $layer=licon1_PDIFF $count=1 $X=0.575
+ $Y=2.32 $X2=0.725 $Y2=2.78
.ends

.subckt PM_SKY130_FD_SC_LS__SDFSTP_1%A_289_464# 1 2 3 4 13 19 21 22 24 25 30 31
+ 34 41 44 46
c123 46 0 1.34962e-19 $X=4.84 $Y=2.495
c124 24 0 4.44907e-20 $X=2.3 $Y=2.49
c125 22 0 9.6166e-20 $X=1.885 $Y=1.005
r126 38 41 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.53 $Y=0.68
+ $X2=4.7 $Y2=0.68
r127 34 36 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.32 $Y=2.325
+ $X2=3.32 $Y2=2.575
r128 30 46 7.64504 $w=4.83e-07 $l=3.1e-07 $layer=LI1_cond $X=4.53 $Y=2.482
+ $X2=4.84 $Y2=2.482
r129 30 44 7.45324 $w=4.83e-07 $l=8.5e-08 $layer=LI1_cond $X=4.53 $Y=2.482
+ $X2=4.445 $Y2=2.482
r130 29 38 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.53 $Y=0.765
+ $X2=4.53 $Y2=0.68
r131 29 30 96.2299 $w=1.68e-07 $l=1.475e-06 $layer=LI1_cond $X=4.53 $Y=0.765
+ $X2=4.53 $Y2=2.24
r132 28 34 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.405 $Y=2.325
+ $X2=3.32 $Y2=2.325
r133 28 44 67.8503 $w=1.68e-07 $l=1.04e-06 $layer=LI1_cond $X=3.405 $Y=2.325
+ $X2=4.445 $Y2=2.325
r134 26 31 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.385 $Y=2.575
+ $X2=2.3 $Y2=2.575
r135 25 36 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.235 $Y=2.575
+ $X2=3.32 $Y2=2.575
r136 25 26 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=3.235 $Y=2.575
+ $X2=2.385 $Y2=2.575
r137 24 31 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.3 $Y=2.49 $X2=2.3
+ $Y2=2.575
r138 23 24 91.3369 $w=1.68e-07 $l=1.4e-06 $layer=LI1_cond $X=2.3 $Y=1.09 $X2=2.3
+ $Y2=2.49
r139 21 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.215 $Y=1.005
+ $X2=2.3 $Y2=1.09
r140 21 22 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.215 $Y=1.005
+ $X2=1.885 $Y2=1.005
r141 17 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.72 $Y=0.92
+ $X2=1.885 $Y2=1.005
r142 17 19 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=1.72 $Y=0.92
+ $X2=1.72 $Y2=0.58
r143 13 31 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=2.3 $Y=2.785
+ $X2=2.3 $Y2=2.575
r144 13 15 24.4318 $w=2.48e-07 $l=5.3e-07 $layer=LI1_cond $X=2.215 $Y=2.785
+ $X2=1.685 $Y2=2.785
r145 4 46 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=4.695
+ $Y=2.285 $X2=4.84 $Y2=2.495
r146 3 15 600 $w=1.7e-07 $l=5.31625e-07 $layer=licon1_PDIFF $count=1 $X=1.445
+ $Y=2.32 $X2=1.685 $Y2=2.745
r147 2 41 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=4.555
+ $Y=0.405 $X2=4.7 $Y2=0.68
r148 1 19 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.58
+ $Y=0.37 $X2=1.72 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_LS__SDFSTP_1%A_1610_341# 1 2 9 11 12 15
r44 13 15 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=9.73 $Y=2.35
+ $X2=9.73 $Y2=2.125
r45 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.565 $Y=2.435
+ $X2=9.73 $Y2=2.35
r46 11 12 78.2888 $w=1.68e-07 $l=1.2e-06 $layer=LI1_cond $X=9.565 $Y=2.435
+ $X2=8.365 $Y2=2.435
r47 7 12 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=8.24 $Y=2.35
+ $X2=8.365 $Y2=2.435
r48 7 9 12.2159 $w=2.48e-07 $l=2.65e-07 $layer=LI1_cond $X=8.24 $Y=2.35 $X2=8.24
+ $Y2=2.085
r49 2 15 300 $w=1.7e-07 $l=3.21364e-07 $layer=licon1_PDIFF $count=2 $X=9.58
+ $Y=1.87 $X2=9.73 $Y2=2.125
r50 1 9 300 $w=1.7e-07 $l=4.48776e-07 $layer=licon1_PDIFF $count=2 $X=8.05
+ $Y=1.705 $X2=8.2 $Y2=2.085
.ends

.subckt PM_SKY130_FD_SC_LS__SDFSTP_1%A_1721_374# 1 2 7 11 14
c30 14 0 1.54803e-19 $X=8.75 $Y=2.855
r31 14 16 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=8.75 $Y=2.855
+ $X2=8.75 $Y2=2.99
r32 9 11 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=10.265 $Y=2.905
+ $X2=10.265 $Y2=2.77
r33 8 16 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.915 $Y=2.99
+ $X2=8.75 $Y2=2.99
r34 7 9 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=10.1 $Y=2.99
+ $X2=10.265 $Y2=2.905
r35 7 8 77.3102 $w=1.68e-07 $l=1.185e-06 $layer=LI1_cond $X=10.1 $Y=2.99
+ $X2=8.915 $Y2=2.99
r36 2 11 600 $w=1.7e-07 $l=2.89741e-07 $layer=licon1_PDIFF $count=1 $X=10.13
+ $Y=2.54 $X2=10.265 $Y2=2.77
r37 1 14 600 $w=1.7e-07 $l=1.05501e-06 $layer=licon1_PDIFF $count=1 $X=8.605
+ $Y=1.87 $X2=8.75 $Y2=2.855
.ends

.subckt PM_SKY130_FD_SC_LS__SDFSTP_1%Q 1 2 7 8 9 10 11 12 13 23
r17 12 13 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=13.69 $Y=2.405
+ $X2=13.69 $Y2=2.775
r18 11 12 19.361 $w=2.48e-07 $l=4.2e-07 $layer=LI1_cond $X=13.69 $Y=1.985
+ $X2=13.69 $Y2=2.405
r19 10 11 14.7513 $w=2.48e-07 $l=3.2e-07 $layer=LI1_cond $X=13.69 $Y=1.665
+ $X2=13.69 $Y2=1.985
r20 9 10 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=13.69 $Y=1.295
+ $X2=13.69 $Y2=1.665
r21 9 43 11.2939 $w=2.48e-07 $l=2.45e-07 $layer=LI1_cond $X=13.69 $Y=1.295
+ $X2=13.69 $Y2=1.05
r22 8 43 5.37855 $w=4.33e-07 $l=1.25e-07 $layer=LI1_cond $X=13.597 $Y=0.925
+ $X2=13.597 $Y2=1.05
r23 8 21 2.43735 $w=4.33e-07 $l=9.2e-08 $layer=LI1_cond $X=13.597 $Y=0.925
+ $X2=13.597 $Y2=0.833
r24 7 21 7.36504 $w=4.33e-07 $l=2.78e-07 $layer=LI1_cond $X=13.597 $Y=0.555
+ $X2=13.597 $Y2=0.833
r25 7 23 1.05972 $w=4.33e-07 $l=4e-08 $layer=LI1_cond $X=13.597 $Y=0.555
+ $X2=13.597 $Y2=0.515
r26 2 13 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=13.5
+ $Y=1.84 $X2=13.65 $Y2=2.815
r27 2 11 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=13.5
+ $Y=1.84 $X2=13.65 $Y2=1.985
r28 1 23 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=13.405
+ $Y=0.37 $X2=13.545 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__SDFSTP_1%VGND 1 2 3 4 5 6 7 26 30 34 38 42 46 50 53
+ 54 56 57 59 60 62 63 64 73 84 105 106 109 112 115
c133 26 0 3.03849e-20 $X=0.86 $Y=0.56
r134 115 116 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r135 112 113 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r136 109 110 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0
+ $X2=0.72 $Y2=0
r137 105 106 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.68 $Y=0
+ $X2=13.68 $Y2=0
r138 103 106 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=12.72 $Y=0
+ $X2=13.68 $Y2=0
r139 102 103 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r140 100 103 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=12.72 $Y2=0
r141 99 102 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=11.28 $Y=0
+ $X2=12.72 $Y2=0
r142 99 100 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r143 97 100 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=11.28 $Y2=0
r144 96 97 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=10.8 $Y=0 $X2=10.8
+ $Y2=0
r145 94 97 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=8.4 $Y=0 $X2=10.8
+ $Y2=0
r146 94 116 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=7.92
+ $Y2=0
r147 93 96 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=8.4 $Y=0 $X2=10.8
+ $Y2=0
r148 93 94 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r149 91 115 15.0812 $w=1.7e-07 $l=4.25e-07 $layer=LI1_cond $X=8.305 $Y=0
+ $X2=7.88 $Y2=0
r150 91 93 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=8.305 $Y=0 $X2=8.4
+ $Y2=0
r151 90 116 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=7.92 $Y2=0
r152 89 90 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r153 86 89 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=6.48 $Y=0 $X2=7.44
+ $Y2=0
r154 86 87 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r155 84 115 15.0812 $w=1.7e-07 $l=4.25e-07 $layer=LI1_cond $X=7.455 $Y=0
+ $X2=7.88 $Y2=0
r156 84 89 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=7.455 $Y=0 $X2=7.44
+ $Y2=0
r157 83 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r158 82 83 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6
+ $Y2=0
r159 80 83 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.08 $Y=0 $X2=6
+ $Y2=0
r160 80 113 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r161 79 82 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.08 $Y=0 $X2=6
+ $Y2=0
r162 79 80 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r163 77 112 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.805 $Y=0
+ $X2=3.64 $Y2=0
r164 77 79 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3.805 $Y=0
+ $X2=4.08 $Y2=0
r165 76 113 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r166 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r167 73 112 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.475 $Y=0
+ $X2=3.64 $Y2=0
r168 73 75 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=3.475 $Y=0
+ $X2=3.12 $Y2=0
r169 72 76 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r170 71 72 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r171 69 72 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r172 69 110 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r173 68 71 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r174 68 69 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r175 66 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.025 $Y=0
+ $X2=0.86 $Y2=0
r176 66 68 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.025 $Y=0 $X2=1.2
+ $Y2=0
r177 64 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r178 64 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=6.48
+ $Y2=0
r179 62 102 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=12.88 $Y=0
+ $X2=12.72 $Y2=0
r180 62 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.88 $Y=0
+ $X2=13.045 $Y2=0
r181 61 105 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=13.21 $Y=0
+ $X2=13.68 $Y2=0
r182 61 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.21 $Y=0
+ $X2=13.045 $Y2=0
r183 59 96 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=10.825 $Y=0
+ $X2=10.8 $Y2=0
r184 59 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.825 $Y=0
+ $X2=10.99 $Y2=0
r185 58 99 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=11.155 $Y=0
+ $X2=11.28 $Y2=0
r186 58 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.155 $Y=0
+ $X2=10.99 $Y2=0
r187 56 82 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=6.115 $Y=0 $X2=6
+ $Y2=0
r188 56 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.115 $Y=0 $X2=6.28
+ $Y2=0
r189 55 86 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=6.445 $Y=0 $X2=6.48
+ $Y2=0
r190 55 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.445 $Y=0 $X2=6.28
+ $Y2=0
r191 53 71 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.375 $Y=0
+ $X2=2.16 $Y2=0
r192 53 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.375 $Y=0 $X2=2.54
+ $Y2=0
r193 52 75 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=2.705 $Y=0
+ $X2=3.12 $Y2=0
r194 52 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.705 $Y=0 $X2=2.54
+ $Y2=0
r195 48 63 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.045 $Y=0.085
+ $X2=13.045 $Y2=0
r196 48 50 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=13.045 $Y=0.085
+ $X2=13.045 $Y2=0.515
r197 44 60 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.99 $Y=0.085
+ $X2=10.99 $Y2=0
r198 44 46 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=10.99 $Y=0.085
+ $X2=10.99 $Y2=0.58
r199 40 115 3.24638 $w=8.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.88 $Y=0.085
+ $X2=7.88 $Y2=0
r200 40 42 6.17176 $w=8.48e-07 $l=4.3e-07 $layer=LI1_cond $X=7.88 $Y=0.085
+ $X2=7.88 $Y2=0.515
r201 36 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.28 $Y=0.085
+ $X2=6.28 $Y2=0
r202 36 38 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=6.28 $Y=0.085
+ $X2=6.28 $Y2=0.575
r203 32 112 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.64 $Y=0.085
+ $X2=3.64 $Y2=0
r204 32 34 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.64 $Y=0.085
+ $X2=3.64 $Y2=0.515
r205 28 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.54 $Y=0.085
+ $X2=2.54 $Y2=0
r206 28 30 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=2.54 $Y=0.085
+ $X2=2.54 $Y2=0.55
r207 24 109 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.86 $Y=0.085
+ $X2=0.86 $Y2=0
r208 24 26 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=0.86 $Y=0.085
+ $X2=0.86 $Y2=0.56
r209 7 50 91 $w=1.7e-07 $l=2.41454e-07 $layer=licon1_NDIFF $count=2 $X=12.825
+ $Y=0.56 $X2=13.045 $Y2=0.515
r210 6 46 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=10.85
+ $Y=0.37 $X2=10.99 $Y2=0.58
r211 5 42 45.5 $w=1.7e-07 $l=6.5643e-07 $layer=licon1_NDIFF $count=4 $X=7.52
+ $Y=0.59 $X2=8.14 $Y2=0.515
r212 4 38 182 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_NDIFF $count=1 $X=6.14
+ $Y=0.405 $X2=6.28 $Y2=0.575
r213 3 34 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=3.43
+ $Y=0.37 $X2=3.64 $Y2=0.515
r214 2 30 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=2.4 $Y=0.37
+ $X2=2.54 $Y2=0.55
r215 1 26 182 $w=1.7e-07 $l=2.89828e-07 $layer=licon1_NDIFF $count=1 $X=0.65
+ $Y=0.37 $X2=0.86 $Y2=0.56
.ends

