* NGSPICE file created from sky130_fd_sc_ls__a221o_2.ext - technology: sky130A

.subckt sky130_fd_sc_ls__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
M1000 a_316_392# B1 a_515_392# VPB phighvt w=1e+06u l=150000u
+  ad=6e+11p pd=5.2e+06u as=5.75e+11p ps=5.15e+06u
M1001 VPWR A1 a_316_392# VPB phighvt w=1e+06u l=150000u
+  ad=9.81e+11p pd=8.31e+06u as=0p ps=0u
M1002 a_337_74# A2 VGND VNB nshort w=740000u l=150000u
+  ad=1.554e+11p pd=1.9e+06u as=8.362e+11p ps=6.7e+06u
M1003 a_515_392# B2 a_316_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_603_74# B1 a_89_260# VNB nshort w=740000u l=150000u
+  ad=1.554e+11p pd=1.9e+06u as=8.029e+11p ps=5.13e+06u
M1005 a_89_260# C1 a_515_392# VPB phighvt w=1e+06u l=150000u
+  ad=2.75e+11p pd=2.55e+06u as=0p ps=0u
M1006 VGND B2 a_603_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_89_260# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=0p ps=0u
M1008 VPWR a_89_260# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_89_260# C1 VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_316_392# A2 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_89_260# A1 a_337_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 X a_89_260# VGND VNB nshort w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1013 VGND a_89_260# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

