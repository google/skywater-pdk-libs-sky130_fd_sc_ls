* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__xnor3_2 A B C VGND VNB VPB VPWR X
X0 a_1027_48# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X1 a_27_373# a_83_247# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 X a_1057_74# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X3 a_83_247# B a_329_81# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X4 a_332_373# a_397_21# a_27_373# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X5 VGND a_1057_74# X VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X6 a_397_21# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X7 X a_1057_74# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X8 a_83_247# B a_332_373# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X9 a_397_21# B VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X10 a_1057_74# C a_332_373# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X11 a_1057_74# C a_329_81# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X12 a_332_373# a_1027_48# a_1057_74# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X13 a_27_373# a_83_247# VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X14 a_1027_48# C VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 a_329_81# a_397_21# a_83_247# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X16 VPWR a_1057_74# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X17 a_329_81# a_1027_48# a_1057_74# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X18 a_27_373# B a_332_373# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X19 a_27_373# B a_329_81# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X20 a_329_81# a_397_21# a_27_373# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X21 VPWR A a_83_247# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X22 VGND A a_83_247# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X23 a_332_373# a_397_21# a_83_247# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
.ends
