* File: sky130_fd_sc_ls__xor2_1.pxi.spice
* Created: Wed Sep  2 11:30:53 2020
* 
x_PM_SKY130_FD_SC_LS__XOR2_1%B N_B_c_68_n N_B_M1003_g N_B_M1000_g N_B_M1002_g
+ N_B_c_64_n N_B_M1004_g N_B_c_65_n B N_B_c_66_n N_B_c_67_n
+ PM_SKY130_FD_SC_LS__XOR2_1%B
x_PM_SKY130_FD_SC_LS__XOR2_1%A N_A_c_130_n N_A_M1006_g N_A_M1005_g N_A_c_132_n
+ N_A_c_133_n N_A_c_134_n N_A_c_135_n N_A_c_141_n N_A_M1007_g N_A_M1001_g
+ N_A_c_137_n A N_A_c_138_n PM_SKY130_FD_SC_LS__XOR2_1%A
x_PM_SKY130_FD_SC_LS__XOR2_1%A_194_125# N_A_194_125#_M1005_d
+ N_A_194_125#_M1003_d N_A_194_125#_M1009_g N_A_194_125#_c_189_n
+ N_A_194_125#_M1008_g N_A_194_125#_c_190_n N_A_194_125#_c_195_n
+ N_A_194_125#_c_227_n N_A_194_125#_c_207_n N_A_194_125#_c_196_n
+ N_A_194_125#_c_191_n N_A_194_125#_c_198_n N_A_194_125#_c_192_n
+ PM_SKY130_FD_SC_LS__XOR2_1%A_194_125#
x_PM_SKY130_FD_SC_LS__XOR2_1%VPWR N_VPWR_M1006_s N_VPWR_M1007_d N_VPWR_c_270_n
+ N_VPWR_c_271_n N_VPWR_c_272_n N_VPWR_c_273_n VPWR N_VPWR_c_274_n
+ N_VPWR_c_275_n N_VPWR_c_269_n N_VPWR_c_277_n PM_SKY130_FD_SC_LS__XOR2_1%VPWR
x_PM_SKY130_FD_SC_LS__XOR2_1%A_355_368# N_A_355_368#_M1007_s
+ N_A_355_368#_M1004_d N_A_355_368#_c_315_n N_A_355_368#_c_313_n
+ N_A_355_368#_c_314_n PM_SKY130_FD_SC_LS__XOR2_1%A_355_368#
x_PM_SKY130_FD_SC_LS__XOR2_1%X N_X_M1002_d N_X_M1008_d N_X_c_337_n N_X_c_340_n
+ N_X_c_341_n N_X_c_338_n X X N_X_c_344_n X PM_SKY130_FD_SC_LS__XOR2_1%X
x_PM_SKY130_FD_SC_LS__XOR2_1%VGND N_VGND_M1005_s N_VGND_M1000_d N_VGND_M1009_d
+ N_VGND_c_371_n N_VGND_c_372_n N_VGND_c_373_n N_VGND_c_374_n N_VGND_c_375_n
+ N_VGND_c_376_n N_VGND_c_377_n N_VGND_c_378_n N_VGND_c_379_n VGND
+ N_VGND_c_380_n PM_SKY130_FD_SC_LS__XOR2_1%VGND
cc_1 VNB N_B_M1000_g 0.0242428f $X=-0.19 $Y=-0.245 $X2=1.69 $Y2=0.9
cc_2 VNB N_B_M1002_g 0.0213738f $X=-0.19 $Y=-0.245 $X2=2.59 $Y2=0.805
cc_3 VNB N_B_c_64_n 0.0227963f $X=-0.19 $Y=-0.245 $X2=2.755 $Y2=1.765
cc_4 VNB N_B_c_65_n 0.0341405f $X=-0.19 $Y=-0.245 $X2=1.45 $Y2=1.53
cc_5 VNB N_B_c_66_n 0.00214447f $X=-0.19 $Y=-0.245 $X2=2.68 $Y2=1.515
cc_6 VNB N_B_c_67_n 0.0156482f $X=-0.19 $Y=-0.245 $X2=2.515 $Y2=1.565
cc_7 VNB N_A_c_130_n 0.034051f $X=-0.19 $Y=-0.245 $X2=1.135 $Y2=1.885
cc_8 VNB N_A_M1005_g 0.0355836f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_c_132_n 0.0949481f $X=-0.19 $Y=-0.245 $X2=2.59 $Y2=1.35
cc_10 VNB N_A_c_133_n 0.0125025f $X=-0.19 $Y=-0.245 $X2=2.59 $Y2=0.805
cc_11 VNB N_A_c_134_n 0.00594968f $X=-0.19 $Y=-0.245 $X2=2.59 $Y2=0.805
cc_12 VNB N_A_c_135_n 0.0149528f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_M1001_g 0.0165166f $X=-0.19 $Y=-0.245 $X2=1.45 $Y2=1.53
cc_14 VNB N_A_c_137_n 0.0616888f $X=-0.19 $Y=-0.245 $X2=2.555 $Y2=1.58
cc_15 VNB N_A_c_138_n 0.0280619f $X=-0.19 $Y=-0.245 $X2=2.68 $Y2=1.515
cc_16 VNB N_A_194_125#_M1009_g 0.0223322f $X=-0.19 $Y=-0.245 $X2=2.59 $Y2=0.805
cc_17 VNB N_A_194_125#_c_189_n 0.0345849f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_194_125#_c_190_n 0.00571579f $X=-0.19 $Y=-0.245 $X2=2.515 $Y2=1.53
cc_19 VNB N_A_194_125#_c_191_n 2.29747e-19 $X=-0.19 $Y=-0.245 $X2=2.68 $Y2=1.515
cc_20 VNB N_A_194_125#_c_192_n 0.00598789f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_VPWR_c_269_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_X_c_337_n 0.0123304f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_X_c_338_n 0.0241086f $X=-0.19 $Y=-0.245 $X2=1.45 $Y2=1.53
cc_24 VNB X 0.00313365f $X=-0.19 $Y=-0.245 $X2=1.45 $Y2=1.53
cc_25 VNB N_VGND_c_371_n 0.0193241f $X=-0.19 $Y=-0.245 $X2=2.59 $Y2=0.805
cc_26 VNB N_VGND_c_372_n 0.0506729f $X=-0.19 $Y=-0.245 $X2=2.755 $Y2=1.765
cc_27 VNB N_VGND_c_373_n 0.0138262f $X=-0.19 $Y=-0.245 $X2=1.45 $Y2=1.53
cc_28 VNB N_VGND_c_374_n 0.0153054f $X=-0.19 $Y=-0.245 $X2=1.135 $Y2=1.885
cc_29 VNB N_VGND_c_375_n 0.0294831f $X=-0.19 $Y=-0.245 $X2=2.68 $Y2=1.515
cc_30 VNB N_VGND_c_376_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=2.68 $Y2=1.515
cc_31 VNB N_VGND_c_377_n 0.0116899f $X=-0.19 $Y=-0.245 $X2=2.68 $Y2=1.515
cc_32 VNB N_VGND_c_378_n 0.0295747f $X=-0.19 $Y=-0.245 $X2=2.64 $Y2=1.565
cc_33 VNB N_VGND_c_379_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=2.515 $Y2=1.565
cc_34 VNB N_VGND_c_380_n 0.241744f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VPB N_B_c_68_n 0.0204565f $X=-0.19 $Y=1.66 $X2=1.135 $Y2=1.885
cc_36 VPB N_B_c_64_n 0.0273121f $X=-0.19 $Y=1.66 $X2=2.755 $Y2=1.765
cc_37 VPB N_B_c_65_n 0.041089f $X=-0.19 $Y=1.66 $X2=1.45 $Y2=1.53
cc_38 VPB N_B_c_66_n 0.00340301f $X=-0.19 $Y=1.66 $X2=2.68 $Y2=1.515
cc_39 VPB N_B_c_67_n 0.00639331f $X=-0.19 $Y=1.66 $X2=2.515 $Y2=1.565
cc_40 VPB N_A_c_130_n 0.039586f $X=-0.19 $Y=1.66 $X2=1.135 $Y2=1.885
cc_41 VPB N_A_c_135_n 6.4402e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_42 VPB N_A_c_141_n 0.0269683f $X=-0.19 $Y=1.66 $X2=2.755 $Y2=1.765
cc_43 VPB N_A_194_125#_c_189_n 0.0266887f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_44 VPB N_A_194_125#_c_190_n 0.00291248f $X=-0.19 $Y=1.66 $X2=2.515 $Y2=1.53
cc_45 VPB N_A_194_125#_c_195_n 0.0130106f $X=-0.19 $Y=1.66 $X2=1.45 $Y2=1.53
cc_46 VPB N_A_194_125#_c_196_n 0.011415f $X=-0.19 $Y=1.66 $X2=1.69 $Y2=1.625
cc_47 VPB N_A_194_125#_c_191_n 0.00132592f $X=-0.19 $Y=1.66 $X2=2.68 $Y2=1.515
cc_48 VPB N_A_194_125#_c_198_n 0.00274616f $X=-0.19 $Y=1.66 $X2=2.515 $Y2=1.565
cc_49 VPB N_VPWR_c_270_n 0.0515201f $X=-0.19 $Y=1.66 $X2=2.59 $Y2=0.805
cc_50 VPB N_VPWR_c_271_n 0.00460404f $X=-0.19 $Y=1.66 $X2=2.515 $Y2=1.53
cc_51 VPB N_VPWR_c_272_n 0.0124854f $X=-0.19 $Y=1.66 $X2=1.45 $Y2=1.53
cc_52 VPB N_VPWR_c_273_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_274_n 0.043458f $X=-0.19 $Y=1.66 $X2=2.68 $Y2=1.515
cc_54 VPB N_VPWR_c_275_n 0.0328281f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_269_n 0.0841696f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_277_n 0.00808603f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_A_355_368#_c_313_n 0.00945387f $X=-0.19 $Y=1.66 $X2=2.755 $Y2=2.4
cc_58 VPB N_A_355_368#_c_314_n 0.00289794f $X=-0.19 $Y=1.66 $X2=1.45 $Y2=1.53
cc_59 VPB N_X_c_340_n 0.0431477f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_X_c_341_n 0.0111298f $X=-0.19 $Y=1.66 $X2=1.45 $Y2=1.53
cc_61 VPB N_X_c_338_n 0.00772436f $X=-0.19 $Y=1.66 $X2=1.45 $Y2=1.53
cc_62 N_B_c_68_n N_A_c_130_n 0.0517042f $X=1.135 $Y=1.885 $X2=-0.19 $Y2=-0.245
cc_63 N_B_c_65_n N_A_c_130_n 0.0170646f $X=1.45 $Y=1.53 $X2=-0.19 $Y2=-0.245
cc_64 N_B_M1000_g N_A_M1005_g 0.00791998f $X=1.69 $Y=0.9 $X2=0 $Y2=0
cc_65 N_B_M1000_g N_A_c_132_n 0.00897099f $X=1.69 $Y=0.9 $X2=0 $Y2=0
cc_66 N_B_M1000_g N_A_c_134_n 0.00857291f $X=1.69 $Y=0.9 $X2=0 $Y2=0
cc_67 N_B_c_64_n N_A_c_135_n 0.0350595f $X=2.755 $Y=1.765 $X2=0 $Y2=0
cc_68 N_B_c_65_n N_A_c_135_n 0.00857291f $X=1.45 $Y=1.53 $X2=0 $Y2=0
cc_69 N_B_c_67_n N_A_c_135_n 0.0190794f $X=2.515 $Y=1.565 $X2=0 $Y2=0
cc_70 N_B_c_64_n N_A_c_141_n 0.0395361f $X=2.755 $Y=1.765 $X2=0 $Y2=0
cc_71 N_B_c_65_n N_A_c_141_n 0.00368422f $X=1.45 $Y=1.53 $X2=0 $Y2=0
cc_72 N_B_c_66_n N_A_c_141_n 0.00191225f $X=2.68 $Y=1.515 $X2=0 $Y2=0
cc_73 N_B_c_67_n N_A_c_141_n 0.00374038f $X=2.515 $Y=1.565 $X2=0 $Y2=0
cc_74 N_B_M1000_g N_A_M1001_g 0.0119366f $X=1.69 $Y=0.9 $X2=0 $Y2=0
cc_75 N_B_M1002_g N_A_M1001_g 0.0350595f $X=2.59 $Y=0.805 $X2=0 $Y2=0
cc_76 N_B_M1002_g N_A_194_125#_M1009_g 0.017662f $X=2.59 $Y=0.805 $X2=0 $Y2=0
cc_77 N_B_c_64_n N_A_194_125#_c_189_n 0.0515053f $X=2.755 $Y=1.765 $X2=0 $Y2=0
cc_78 N_B_c_66_n N_A_194_125#_c_189_n 4.88812e-19 $X=2.68 $Y=1.515 $X2=0 $Y2=0
cc_79 N_B_c_68_n N_A_194_125#_c_190_n 0.00309103f $X=1.135 $Y=1.885 $X2=0 $Y2=0
cc_80 N_B_M1000_g N_A_194_125#_c_190_n 0.00509445f $X=1.69 $Y=0.9 $X2=0 $Y2=0
cc_81 N_B_c_65_n N_A_194_125#_c_190_n 0.0130411f $X=1.45 $Y=1.53 $X2=0 $Y2=0
cc_82 N_B_c_67_n N_A_194_125#_c_190_n 0.0262124f $X=2.515 $Y=1.565 $X2=0 $Y2=0
cc_83 N_B_c_68_n N_A_194_125#_c_195_n 0.0192913f $X=1.135 $Y=1.885 $X2=0 $Y2=0
cc_84 N_B_M1000_g N_A_194_125#_c_207_n 0.00436246f $X=1.69 $Y=0.9 $X2=0 $Y2=0
cc_85 N_B_c_65_n N_A_194_125#_c_207_n 0.011061f $X=1.45 $Y=1.53 $X2=0 $Y2=0
cc_86 N_B_c_67_n N_A_194_125#_c_207_n 0.0152632f $X=2.515 $Y=1.565 $X2=0 $Y2=0
cc_87 N_B_c_64_n N_A_194_125#_c_196_n 0.012205f $X=2.755 $Y=1.765 $X2=0 $Y2=0
cc_88 N_B_c_65_n N_A_194_125#_c_196_n 0.00561489f $X=1.45 $Y=1.53 $X2=0 $Y2=0
cc_89 N_B_c_66_n N_A_194_125#_c_196_n 0.0226668f $X=2.68 $Y=1.515 $X2=0 $Y2=0
cc_90 N_B_c_67_n N_A_194_125#_c_196_n 0.0528266f $X=2.515 $Y=1.565 $X2=0 $Y2=0
cc_91 N_B_c_64_n N_A_194_125#_c_191_n 0.00395687f $X=2.755 $Y=1.765 $X2=0 $Y2=0
cc_92 N_B_c_66_n N_A_194_125#_c_191_n 0.00957646f $X=2.68 $Y=1.515 $X2=0 $Y2=0
cc_93 N_B_c_68_n N_A_194_125#_c_198_n 0.00808399f $X=1.135 $Y=1.885 $X2=0 $Y2=0
cc_94 N_B_c_65_n N_A_194_125#_c_198_n 0.0096596f $X=1.45 $Y=1.53 $X2=0 $Y2=0
cc_95 N_B_c_67_n N_A_194_125#_c_198_n 0.0149541f $X=2.515 $Y=1.565 $X2=0 $Y2=0
cc_96 N_B_M1002_g N_A_194_125#_c_192_n 5.92648e-19 $X=2.59 $Y=0.805 $X2=0 $Y2=0
cc_97 N_B_c_64_n N_A_194_125#_c_192_n 0.00105206f $X=2.755 $Y=1.765 $X2=0 $Y2=0
cc_98 N_B_c_66_n N_A_194_125#_c_192_n 0.0243048f $X=2.68 $Y=1.515 $X2=0 $Y2=0
cc_99 N_B_c_68_n N_VPWR_c_270_n 0.00148391f $X=1.135 $Y=1.885 $X2=0 $Y2=0
cc_100 N_B_c_64_n N_VPWR_c_271_n 0.0127571f $X=2.755 $Y=1.765 $X2=0 $Y2=0
cc_101 N_B_c_68_n N_VPWR_c_274_n 0.00291513f $X=1.135 $Y=1.885 $X2=0 $Y2=0
cc_102 N_B_c_64_n N_VPWR_c_275_n 0.00413917f $X=2.755 $Y=1.765 $X2=0 $Y2=0
cc_103 N_B_c_68_n N_VPWR_c_269_n 0.00364018f $X=1.135 $Y=1.885 $X2=0 $Y2=0
cc_104 N_B_c_64_n N_VPWR_c_269_n 0.00818241f $X=2.755 $Y=1.765 $X2=0 $Y2=0
cc_105 N_B_c_64_n N_A_355_368#_c_315_n 0.0154234f $X=2.755 $Y=1.765 $X2=0 $Y2=0
cc_106 N_B_c_68_n N_A_355_368#_c_313_n 9.28949e-19 $X=1.135 $Y=1.885 $X2=0 $Y2=0
cc_107 N_B_c_64_n N_A_355_368#_c_314_n 0.00283124f $X=2.755 $Y=1.765 $X2=0 $Y2=0
cc_108 N_B_M1002_g X 0.0144534f $X=2.59 $Y=0.805 $X2=0 $Y2=0
cc_109 N_B_M1002_g N_X_c_344_n 0.00594253f $X=2.59 $Y=0.805 $X2=0 $Y2=0
cc_110 N_B_c_64_n N_X_c_344_n 0.00454365f $X=2.755 $Y=1.765 $X2=0 $Y2=0
cc_111 N_B_c_66_n N_X_c_344_n 0.0210499f $X=2.68 $Y=1.515 $X2=0 $Y2=0
cc_112 N_B_M1000_g N_VGND_c_373_n 0.00705087f $X=1.69 $Y=0.9 $X2=0 $Y2=0
cc_113 N_B_M1002_g N_VGND_c_373_n 0.00272515f $X=2.59 $Y=0.805 $X2=0 $Y2=0
cc_114 N_B_c_67_n N_VGND_c_373_n 0.0286839f $X=2.515 $Y=1.565 $X2=0 $Y2=0
cc_115 N_B_M1002_g N_VGND_c_374_n 6.01743e-19 $X=2.59 $Y=0.805 $X2=0 $Y2=0
cc_116 N_B_M1002_g N_VGND_c_378_n 0.00395427f $X=2.59 $Y=0.805 $X2=0 $Y2=0
cc_117 N_B_M1000_g N_VGND_c_380_n 9.49986e-19 $X=1.69 $Y=0.9 $X2=0 $Y2=0
cc_118 N_B_M1002_g N_VGND_c_380_n 0.00525227f $X=2.59 $Y=0.805 $X2=0 $Y2=0
cc_119 N_A_c_130_n N_A_194_125#_c_190_n 0.0123887f $X=0.715 $Y=1.885 $X2=0 $Y2=0
cc_120 N_A_M1005_g N_A_194_125#_c_190_n 0.00959846f $X=0.895 $Y=0.9 $X2=0 $Y2=0
cc_121 N_A_c_138_n N_A_194_125#_c_190_n 0.034045f $X=0.61 $Y=1.45 $X2=0 $Y2=0
cc_122 N_A_c_130_n N_A_194_125#_c_195_n 0.00703532f $X=0.715 $Y=1.885 $X2=0
+ $Y2=0
cc_123 N_A_c_141_n N_A_194_125#_c_195_n 0.00406169f $X=2.185 $Y=1.765 $X2=0
+ $Y2=0
cc_124 N_A_M1005_g N_A_194_125#_c_227_n 0.00589874f $X=0.895 $Y=0.9 $X2=0 $Y2=0
cc_125 N_A_c_132_n N_A_194_125#_c_227_n 0.00100425f $X=2.125 $Y=0.18 $X2=0 $Y2=0
cc_126 N_A_c_132_n N_A_194_125#_c_207_n 0.00843612f $X=2.125 $Y=0.18 $X2=0 $Y2=0
cc_127 N_A_c_141_n N_A_194_125#_c_196_n 0.0136239f $X=2.185 $Y=1.765 $X2=0 $Y2=0
cc_128 N_A_c_130_n N_A_194_125#_c_198_n 0.00143427f $X=0.715 $Y=1.885 $X2=0
+ $Y2=0
cc_129 N_A_c_130_n N_VPWR_c_270_n 0.018623f $X=0.715 $Y=1.885 $X2=0 $Y2=0
cc_130 N_A_c_137_n N_VPWR_c_270_n 0.00633983f $X=0.625 $Y=1.45 $X2=0 $Y2=0
cc_131 N_A_c_138_n N_VPWR_c_270_n 0.0173129f $X=0.61 $Y=1.45 $X2=0 $Y2=0
cc_132 N_A_c_141_n N_VPWR_c_271_n 0.0146814f $X=2.185 $Y=1.765 $X2=0 $Y2=0
cc_133 N_A_c_130_n N_VPWR_c_274_n 0.00413917f $X=0.715 $Y=1.885 $X2=0 $Y2=0
cc_134 N_A_c_141_n N_VPWR_c_274_n 0.00444681f $X=2.185 $Y=1.765 $X2=0 $Y2=0
cc_135 N_A_c_130_n N_VPWR_c_269_n 0.00817532f $X=0.715 $Y=1.885 $X2=0 $Y2=0
cc_136 N_A_c_141_n N_VPWR_c_269_n 0.00882517f $X=2.185 $Y=1.765 $X2=0 $Y2=0
cc_137 N_A_c_141_n N_A_355_368#_c_315_n 0.0132362f $X=2.185 $Y=1.765 $X2=0 $Y2=0
cc_138 N_A_c_141_n N_A_355_368#_c_313_n 4.61562e-19 $X=2.185 $Y=1.765 $X2=0
+ $Y2=0
cc_139 N_A_M1001_g X 0.00192367f $X=2.2 $Y=0.805 $X2=0 $Y2=0
cc_140 N_A_M1001_g N_X_c_344_n 5.78169e-19 $X=2.2 $Y=0.805 $X2=0 $Y2=0
cc_141 N_A_c_133_n N_VGND_c_372_n 0.0232133f $X=0.97 $Y=0.18 $X2=0 $Y2=0
cc_142 N_A_c_137_n N_VGND_c_372_n 0.00360255f $X=0.625 $Y=1.45 $X2=0 $Y2=0
cc_143 N_A_c_138_n N_VGND_c_372_n 0.0484114f $X=0.61 $Y=1.45 $X2=0 $Y2=0
cc_144 N_A_c_132_n N_VGND_c_373_n 0.0226627f $X=2.125 $Y=0.18 $X2=0 $Y2=0
cc_145 N_A_c_134_n N_VGND_c_373_n 9.08308e-19 $X=2.185 $Y=1.34 $X2=0 $Y2=0
cc_146 N_A_M1001_g N_VGND_c_373_n 0.0204272f $X=2.2 $Y=0.805 $X2=0 $Y2=0
cc_147 N_A_c_133_n N_VGND_c_375_n 0.0292218f $X=0.97 $Y=0.18 $X2=0 $Y2=0
cc_148 N_A_c_132_n N_VGND_c_378_n 0.00486043f $X=2.125 $Y=0.18 $X2=0 $Y2=0
cc_149 N_A_c_132_n N_VGND_c_380_n 0.0354577f $X=2.125 $Y=0.18 $X2=0 $Y2=0
cc_150 N_A_c_133_n N_VGND_c_380_n 0.0106607f $X=0.97 $Y=0.18 $X2=0 $Y2=0
cc_151 N_A_194_125#_c_196_n N_VPWR_M1007_d 0.00728707f $X=3.025 $Y=2.035 $X2=0
+ $Y2=0
cc_152 N_A_194_125#_c_190_n N_VPWR_c_270_n 4.78333e-19 $X=1.03 $Y=1.95 $X2=0
+ $Y2=0
cc_153 N_A_194_125#_c_195_n N_VPWR_c_270_n 0.0463803f $X=1.36 $Y=2.815 $X2=0
+ $Y2=0
cc_154 N_A_194_125#_c_198_n N_VPWR_c_270_n 0.00933212f $X=1.36 $Y=2.115 $X2=0
+ $Y2=0
cc_155 N_A_194_125#_c_189_n N_VPWR_c_271_n 6.05438e-19 $X=3.255 $Y=1.765 $X2=0
+ $Y2=0
cc_156 N_A_194_125#_c_195_n N_VPWR_c_274_n 0.0253425f $X=1.36 $Y=2.815 $X2=0
+ $Y2=0
cc_157 N_A_194_125#_c_189_n N_VPWR_c_275_n 0.00445602f $X=3.255 $Y=1.765 $X2=0
+ $Y2=0
cc_158 N_A_194_125#_c_189_n N_VPWR_c_269_n 0.00862596f $X=3.255 $Y=1.765 $X2=0
+ $Y2=0
cc_159 N_A_194_125#_c_195_n N_VPWR_c_269_n 0.020624f $X=1.36 $Y=2.815 $X2=0
+ $Y2=0
cc_160 N_A_194_125#_c_195_n A_158_392# 0.00901843f $X=1.36 $Y=2.815 $X2=-0.19
+ $Y2=-0.245
cc_161 N_A_194_125#_c_198_n A_158_392# 0.00172559f $X=1.36 $Y=2.115 $X2=-0.19
+ $Y2=-0.245
cc_162 N_A_194_125#_c_196_n N_A_355_368#_M1007_s 0.00794845f $X=3.025 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_163 N_A_194_125#_c_196_n N_A_355_368#_M1004_d 0.00774505f $X=3.025 $Y=2.035
+ $X2=0 $Y2=0
cc_164 N_A_194_125#_c_191_n N_A_355_368#_M1004_d 0.00128638f $X=3.11 $Y=1.95
+ $X2=0 $Y2=0
cc_165 N_A_194_125#_c_196_n N_A_355_368#_c_315_n 0.042526f $X=3.025 $Y=2.035
+ $X2=0 $Y2=0
cc_166 N_A_194_125#_c_195_n N_A_355_368#_c_313_n 0.0492557f $X=1.36 $Y=2.815
+ $X2=0 $Y2=0
cc_167 N_A_194_125#_c_196_n N_A_355_368#_c_313_n 0.0243359f $X=3.025 $Y=2.035
+ $X2=0 $Y2=0
cc_168 N_A_194_125#_c_189_n N_A_355_368#_c_314_n 0.00762227f $X=3.255 $Y=1.765
+ $X2=0 $Y2=0
cc_169 N_A_194_125#_c_196_n N_A_355_368#_c_314_n 0.0208833f $X=3.025 $Y=2.035
+ $X2=0 $Y2=0
cc_170 N_A_194_125#_M1009_g N_X_c_337_n 0.0166901f $X=3.16 $Y=0.805 $X2=0 $Y2=0
cc_171 N_A_194_125#_c_189_n N_X_c_337_n 0.00430636f $X=3.255 $Y=1.765 $X2=0
+ $Y2=0
cc_172 N_A_194_125#_c_192_n N_X_c_337_n 0.0245397f $X=3.25 $Y=1.485 $X2=0 $Y2=0
cc_173 N_A_194_125#_c_189_n N_X_c_341_n 0.02399f $X=3.255 $Y=1.765 $X2=0 $Y2=0
cc_174 N_A_194_125#_c_191_n N_X_c_341_n 0.00518254f $X=3.11 $Y=1.95 $X2=0 $Y2=0
cc_175 N_A_194_125#_c_192_n N_X_c_341_n 0.00413233f $X=3.25 $Y=1.485 $X2=0 $Y2=0
cc_176 N_A_194_125#_M1009_g N_X_c_338_n 0.00477786f $X=3.16 $Y=0.805 $X2=0 $Y2=0
cc_177 N_A_194_125#_c_189_n N_X_c_338_n 0.00569949f $X=3.255 $Y=1.765 $X2=0
+ $Y2=0
cc_178 N_A_194_125#_c_191_n N_X_c_338_n 0.00651169f $X=3.11 $Y=1.95 $X2=0 $Y2=0
cc_179 N_A_194_125#_c_192_n N_X_c_338_n 0.0250916f $X=3.25 $Y=1.485 $X2=0 $Y2=0
cc_180 N_A_194_125#_M1009_g X 0.00974015f $X=3.16 $Y=0.805 $X2=0 $Y2=0
cc_181 N_A_194_125#_M1009_g N_VGND_c_374_n 0.00972215f $X=3.16 $Y=0.805 $X2=0
+ $Y2=0
cc_182 N_A_194_125#_c_227_n N_VGND_c_375_n 0.00228482f $X=1.115 $Y=0.875 $X2=0
+ $Y2=0
cc_183 N_A_194_125#_c_207_n N_VGND_c_375_n 0.00771542f $X=1.475 $Y=0.875 $X2=0
+ $Y2=0
cc_184 N_A_194_125#_M1009_g N_VGND_c_378_n 0.00441186f $X=3.16 $Y=0.805 $X2=0
+ $Y2=0
cc_185 N_A_194_125#_M1009_g N_VGND_c_380_n 0.0044119f $X=3.16 $Y=0.805 $X2=0
+ $Y2=0
cc_186 N_A_194_125#_c_227_n N_VGND_c_380_n 0.00415706f $X=1.115 $Y=0.875 $X2=0
+ $Y2=0
cc_187 N_A_194_125#_c_207_n N_VGND_c_380_n 0.012469f $X=1.475 $Y=0.875 $X2=0
+ $Y2=0
cc_188 N_VPWR_M1007_d N_A_355_368#_c_315_n 0.0071329f $X=2.26 $Y=1.84 $X2=0
+ $Y2=0
cc_189 N_VPWR_c_271_n N_A_355_368#_c_315_n 0.0241655f $X=2.475 $Y=2.815 $X2=0
+ $Y2=0
cc_190 N_VPWR_c_271_n N_A_355_368#_c_313_n 0.01373f $X=2.475 $Y=2.815 $X2=0
+ $Y2=0
cc_191 N_VPWR_c_274_n N_A_355_368#_c_313_n 0.0146513f $X=2.255 $Y=3.33 $X2=0
+ $Y2=0
cc_192 N_VPWR_c_269_n N_A_355_368#_c_313_n 0.0121202f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_193 N_VPWR_c_271_n N_A_355_368#_c_314_n 0.01373f $X=2.475 $Y=2.815 $X2=0
+ $Y2=0
cc_194 N_VPWR_c_275_n N_A_355_368#_c_314_n 0.0146094f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_195 N_VPWR_c_269_n N_A_355_368#_c_314_n 0.0120527f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_196 N_VPWR_c_275_n N_X_c_340_n 0.0173129f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_197 N_VPWR_c_269_n N_X_c_340_n 0.0143301f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_198 N_A_355_368#_c_314_n N_X_c_340_n 0.0202848f $X=3.03 $Y=2.455 $X2=0 $Y2=0
cc_199 N_X_c_337_n N_VGND_M1009_d 0.0136501f $X=3.585 $Y=1.065 $X2=0 $Y2=0
cc_200 N_X_c_338_n N_VGND_M1009_d 3.82603e-19 $X=3.56 $Y=1.82 $X2=0 $Y2=0
cc_201 X N_VGND_c_373_n 0.0229507f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_202 N_X_c_344_n N_VGND_c_373_n 0.00716572f $X=2.747 $Y=0.98 $X2=0 $Y2=0
cc_203 N_X_c_337_n N_VGND_c_374_n 0.0171814f $X=3.585 $Y=1.065 $X2=0 $Y2=0
cc_204 X N_VGND_c_374_n 0.0201618f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_205 X N_VGND_c_378_n 0.0152785f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_206 X N_VGND_c_380_n 0.0155747f $X=2.555 $Y=0.47 $X2=0 $Y2=0
