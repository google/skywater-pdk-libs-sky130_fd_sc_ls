* File: sky130_fd_sc_ls__ha_1.spice
* Created: Fri Aug 28 13:27:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__ha_1.pex.spice"
.subckt sky130_fd_sc_ls__ha_1  VNB VPB B A SUM VPWR COUT VGND
* 
* VGND	VGND
* COUT	COUT
* VPWR	VPWR
* SUM	SUM
* A	A
* B	B
* VPB	VPB
* VNB	VNB
MM1011 N_VGND_M1011_d N_A_83_260#_M1011_g N_SUM_M1011_s VNB NSHORT L=0.15 W=0.74
+ AD=0.19515 AS=0.2109 PD=2.05 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1007 N_A_305_130#_M1007_d N_A_239_294#_M1007_g N_A_83_260#_M1007_s VNB NSHORT
+ L=0.15 W=0.64 AD=0.0896 AS=0.1726 PD=0.92 PS=1.85 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1008 N_VGND_M1008_d N_B_M1008_g N_A_305_130#_M1007_d VNB NSHORT L=0.15 W=0.64
+ AD=0.125537 AS=0.0896 PD=1.065 PS=0.92 NRD=1.872 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1013 N_A_305_130#_M1013_d N_A_M1013_g N_VGND_M1008_d VNB NSHORT L=0.15 W=0.64
+ AD=0.1824 AS=0.125537 PD=1.85 PS=1.065 NRD=0 NRS=16.872 M=1 R=4.26667
+ SA=75001.1 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1000 A_695_119# N_B_M1000_g N_A_239_294#_M1000_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0672 AS=0.1824 PD=0.85 PS=1.85 NRD=9.372 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75001.1 A=0.096 P=1.58 MULT=1
MM1009 N_VGND_M1009_d N_A_M1009_g A_695_119# VNB NSHORT L=0.15 W=0.64
+ AD=0.115478 AS=0.0672 PD=1.01101 PS=0.85 NRD=0 NRS=9.372 M=1 R=4.26667
+ SA=75000.6 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1005 N_COUT_M1005_d N_A_239_294#_M1005_g N_VGND_M1009_d VNB NSHORT L=0.15
+ W=0.74 AD=0.2109 AS=0.133522 PD=2.05 PS=1.16899 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75000.9 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1006 N_VPWR_M1006_d N_A_83_260#_M1006_g N_SUM_M1006_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.407086 AS=0.3304 PD=2.07429 PS=2.83 NRD=35.1645 NRS=1.7533 M=1
+ R=7.46667 SA=75000.2 SB=75002.8 A=0.168 P=2.54 MULT=1
MM1002 N_A_83_260#_M1002_d N_A_239_294#_M1002_g N_VPWR_M1006_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.155491 AS=0.305314 PD=1.23717 PS=1.55571 NRD=2.3443
+ NRS=51.5943 M=1 R=5.6 SA=75001.1 SB=75002.8 A=0.126 P=1.98 MULT=1
MM1003 A_386_392# N_B_M1003_g N_A_83_260#_M1002_d VPB PHIGHVT L=0.15 W=1 AD=0.21
+ AS=0.185109 PD=1.42 PS=1.47283 NRD=30.5153 NRS=12.7853 M=1 R=6.66667
+ SA=75001.3 SB=75002.3 A=0.15 P=2.3 MULT=1
MM1012 N_VPWR_M1012_d N_A_M1012_g A_386_392# VPB PHIGHVT L=0.15 W=1 AD=0.331196
+ AS=0.21 PD=1.82065 PS=1.42 NRD=1.9503 NRS=30.5153 M=1 R=6.66667 SA=75001.9
+ SB=75001.7 A=0.15 P=2.3 MULT=1
MM1010 N_A_239_294#_M1010_d N_B_M1010_g N_VPWR_M1012_d VPB PHIGHVT L=0.15 W=0.84
+ AD=0.126 AS=0.278204 PD=1.14 PS=1.52935 NRD=2.3443 NRS=2.3443 M=1 R=5.6
+ SA=75002.7 SB=75001.2 A=0.126 P=1.98 MULT=1
MM1001 N_VPWR_M1001_d N_A_M1001_g N_A_239_294#_M1010_d VPB PHIGHVT L=0.15 W=0.84
+ AD=0.1758 AS=0.126 PD=1.30286 PS=1.14 NRD=14.0658 NRS=2.3443 M=1 R=5.6
+ SA=75003.2 SB=75000.8 A=0.126 P=1.98 MULT=1
MM1004 N_COUT_M1004_d N_A_239_294#_M1004_g N_VPWR_M1001_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.3304 AS=0.2344 PD=2.83 PS=1.73714 NRD=1.7533 NRS=10.5395 M=1
+ R=7.46667 SA=75002.8 SB=75000.2 A=0.168 P=2.54 MULT=1
DX14_noxref VNB VPB NWDIODE A=9.471 P=14.32
c_87 VPB 0 2.55746e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_ls__ha_1.pxi.spice"
*
.ends
*
*
