* NGSPICE file created from sky130_fd_sc_ls__einvn_1.ext - technology: sky130A

.subckt sky130_fd_sc_ls__einvn_1 A TE_B VGND VNB VPB VPWR Z
M1000 a_281_100# a_22_46# VGND VNB nshort w=740000u l=150000u
+  ad=1.776e+11p pd=1.96e+06u as=2.564e+11p ps=2.36e+06u
M1001 Z A a_278_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=3.024e+11p ps=2.78e+06u
M1002 Z A a_281_100# VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1003 a_278_368# TE_B VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.88e+11p ps=3.01e+06u
M1004 VGND TE_B a_22_46# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.218e+11p ps=1.42e+06u
M1005 VPWR TE_B a_22_46# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.888e+11p ps=1.87e+06u
.ends

