* NGSPICE file created from sky130_fd_sc_ls__decap_8.ext - technology: sky130A

.subckt sky130_fd_sc_ls__decap_8 VGND VNB VPB VPWR
M1000 VGND VPWR VGND VNB nshort w=420000u l=1e+06u
+  ad=6.279e+11p pd=5.51e+06u as=0p ps=0u
M1001 VGND VPWR VGND VNB nshort w=420000u l=1e+06u
+  ad=0p pd=0u as=0p ps=0u
M1002 VPWR VGND VPWR VPB phighvt w=1e+06u l=1e+06u
+  ad=1.57e+12p pd=9.14e+06u as=0p ps=0u
M1003 VPWR VGND VPWR VPB phighvt w=1e+06u l=1e+06u
+  ad=0p pd=0u as=0p ps=0u
.ends

