# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ls__o41ai_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ls__o41ai_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.240000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.350000 1.350000 6.115000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.765000 1.350000 5.155000 1.680000 ;
        RECT 4.925000 1.680000 5.155000 1.780000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005000 1.350000 3.455000 1.780000 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.405000 1.350000 2.755000 1.780000 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.280000 0.455000 1.180000 ;
        RECT 0.125000 1.180000 0.900000 1.550000 ;
        RECT 0.125000 1.550000 0.455000 1.630000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.879200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.635000 1.720000 2.235000 1.890000 ;
        RECT 0.635000 1.890000 0.805000 2.980000 ;
        RECT 1.070000 0.645000 1.400000 1.550000 ;
        RECT 1.070000 1.550000 2.235000 1.720000 ;
        RECT 2.035000 1.890000 2.235000 2.735000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 6.240000 0.085000 ;
        RECT 2.070000  0.085000 2.400000 0.795000 ;
        RECT 3.000000  0.085000 3.330000 0.795000 ;
        RECT 3.960000  0.085000 4.290000 0.795000 ;
        RECT 4.960000  0.085000 5.290000 0.795000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.240000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 6.240000 3.415000 ;
        RECT 0.105000 1.820000 0.435000 3.245000 ;
        RECT 1.005000 2.060000 1.335000 3.245000 ;
        RECT 5.435000 2.290000 5.605000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 6.240000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.640000 0.255000 1.900000 0.425000 ;
      RECT 0.640000 0.425000 0.890000 1.010000 ;
      RECT 1.535000 2.060000 1.865000 2.905000 ;
      RECT 1.535000 2.905000 2.765000 3.075000 ;
      RECT 1.570000 0.425000 1.900000 1.010000 ;
      RECT 1.570000 1.010000 5.790000 1.180000 ;
      RECT 2.435000 1.950000 3.800000 2.120000 ;
      RECT 2.435000 2.120000 2.765000 2.905000 ;
      RECT 2.580000 0.350000 2.830000 1.010000 ;
      RECT 3.020000 2.290000 3.270000 2.905000 ;
      RECT 3.020000 2.905000 4.705000 3.075000 ;
      RECT 3.470000 2.120000 3.800000 2.735000 ;
      RECT 3.510000 0.350000 3.790000 1.010000 ;
      RECT 4.005000 1.850000 4.335000 1.950000 ;
      RECT 4.005000 1.950000 6.135000 2.120000 ;
      RECT 4.005000 2.120000 4.335000 2.735000 ;
      RECT 4.460000 0.350000 4.790000 1.010000 ;
      RECT 4.535000 2.290000 4.705000 2.905000 ;
      RECT 4.905000 2.120000 5.235000 2.980000 ;
      RECT 5.460000 0.350000 5.790000 1.010000 ;
      RECT 5.805000 2.120000 6.135000 2.980000 ;
  END
END sky130_fd_sc_ls__o41ai_2
