* File: sky130_fd_sc_ls__sdlclkp_4.pex.spice
* Created: Fri Aug 28 14:06:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__SDLCLKP_4%SCE 1 3 6 8 12
r23 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.62 $X2=0.385 $Y2=1.62
r24 8 12 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=0.24 $Y=1.62
+ $X2=0.385 $Y2=1.62
r25 4 11 38.5661 $w=3.24e-07 $l=2.14173e-07 $layer=POLY_cond $X=0.52 $Y=1.455
+ $X2=0.407 $Y2=1.62
r26 4 6 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.52 $Y=1.455
+ $X2=0.52 $Y2=0.99
r27 1 11 55.6741 $w=3.24e-07 $l=3.25331e-07 $layer=POLY_cond $X=0.505 $Y=1.9
+ $X2=0.407 $Y2=1.62
r28 1 3 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.505 $Y=1.9 $X2=0.505
+ $Y2=2.395
.ends

.subckt PM_SKY130_FD_SC_LS__SDLCLKP_4%GATE 1 3 6 8
c31 8 0 1.03187e-19 $X=1.2 $Y=1.665
r32 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1 $Y=1.62
+ $X2=1 $Y2=1.62
r33 8 12 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=1.2 $Y=1.62 $X2=1
+ $Y2=1.62
r34 4 11 38.6072 $w=2.91e-07 $l=1.67481e-07 $layer=POLY_cond $X=0.995 $Y=1.455
+ $X2=1 $Y2=1.62
r35 4 6 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.995 $Y=1.455
+ $X2=0.995 $Y2=0.99
r36 1 11 57.6553 $w=2.91e-07 $l=3.15278e-07 $layer=POLY_cond $X=0.925 $Y=1.9
+ $X2=1 $Y2=1.62
r37 1 3 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.925 $Y=1.9 $X2=0.925
+ $Y2=2.395
.ends

.subckt PM_SKY130_FD_SC_LS__SDLCLKP_4%A_354_105# 1 2 7 9 10 14 18 20 21 24 26 28
+ 30
c79 28 0 3.22822e-20 $X=2.53 $Y=1.65
c80 14 0 1.62426e-20 $X=3.645 $Y=0.58
c81 7 0 1.84961e-19 $X=3.315 $Y=1.82
r82 31 35 10.378 $w=4.18e-07 $l=9e-08 $layer=POLY_cond $X=3.165 $Y=1.57
+ $X2=3.165 $Y2=1.48
r83 30 33 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=3.09 $Y=1.57 $X2=3.09
+ $Y2=1.65
r84 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.09
+ $Y=1.57 $X2=3.09 $Y2=1.57
r85 27 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.695 $Y=1.65
+ $X2=2.53 $Y2=1.65
r86 26 33 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.925 $Y=1.65
+ $X2=3.09 $Y2=1.65
r87 26 27 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=2.925 $Y=1.65
+ $X2=2.695 $Y2=1.65
r88 22 28 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.53 $Y=1.735
+ $X2=2.53 $Y2=1.65
r89 22 24 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=2.53 $Y=1.735
+ $X2=2.53 $Y2=1.975
r90 20 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.365 $Y=1.65
+ $X2=2.53 $Y2=1.65
r91 20 21 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=2.365 $Y=1.65
+ $X2=2.075 $Y2=1.65
r92 16 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.95 $Y=1.565
+ $X2=2.075 $Y2=1.65
r93 16 18 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=1.95 $Y=1.565
+ $X2=1.95 $Y2=1.12
r94 12 14 423.032 $w=1.5e-07 $l=8.25e-07 $layer=POLY_cond $X=3.645 $Y=1.405
+ $X2=3.645 $Y2=0.58
r95 11 35 26.9416 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=3.405 $Y=1.48
+ $X2=3.165 $Y2=1.48
r96 10 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.57 $Y=1.48
+ $X2=3.645 $Y2=1.405
r97 10 11 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.57 $Y=1.48
+ $X2=3.405 $Y2=1.48
r98 7 31 49.7565 $w=4.18e-07 $l=3.16228e-07 $layer=POLY_cond $X=3.315 $Y=1.82
+ $X2=3.165 $Y2=1.57
r99 7 9 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=3.315 $Y=1.82
+ $X2=3.315 $Y2=2.315
r100 2 24 600 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=1 $X=2.295
+ $Y=2.12 $X2=2.53 $Y2=1.975
r101 1 18 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=1.77
+ $Y=0.525 $X2=1.91 $Y2=1.12
.ends

.subckt PM_SKY130_FD_SC_LS__SDLCLKP_4%A_324_79# 1 2 7 9 10 11 13 14 17 18 19 20
+ 22 24 25 26 27 29 30 33 34 35 37 38 39 41 42 43 47 50 57 58 60 61
c164 58 0 1.06701e-19 $X=5.607 $Y=1.82
c165 47 0 1.46172e-19 $X=5.67 $Y=0.515
c166 42 0 9.27061e-20 $X=5.445 $Y=0.34
c167 38 0 6.61483e-20 $X=4.605 $Y=0.98
c168 33 0 1.62426e-20 $X=2.89 $Y=1.065
c169 30 0 1.84961e-19 $X=2.805 $Y=1.15
c170 11 0 1.84401e-19 $X=1.77 $Y=1.415
r171 58 60 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=5.53 $Y=1.82
+ $X2=5.53 $Y2=1.01
r172 57 58 8.46614 $w=3.33e-07 $l=1.65e-07 $layer=LI1_cond $X=5.607 $Y=1.985
+ $X2=5.607 $Y2=1.82
r173 54 61 13.7476 $w=4.45e-07 $l=1.1e-07 $layer=POLY_cond $X=2.352 $Y=1.23
+ $X2=2.352 $Y2=1.12
r174 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.41
+ $Y=1.23 $X2=2.41 $Y2=1.23
r175 50 53 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=2.41 $Y=1.15 $X2=2.41
+ $Y2=1.23
r176 45 60 9.49412 $w=3.88e-07 $l=1.95e-07 $layer=LI1_cond $X=5.64 $Y=0.815
+ $X2=5.64 $Y2=1.01
r177 45 47 8.86495 $w=3.88e-07 $l=3e-07 $layer=LI1_cond $X=5.64 $Y=0.815
+ $X2=5.64 $Y2=0.515
r178 44 47 2.65948 $w=3.88e-07 $l=9e-08 $layer=LI1_cond $X=5.64 $Y=0.425
+ $X2=5.64 $Y2=0.515
r179 42 44 8.28377 $w=1.7e-07 $l=2.33666e-07 $layer=LI1_cond $X=5.445 $Y=0.34
+ $X2=5.64 $Y2=0.425
r180 42 43 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.445 $Y=0.34
+ $X2=4.775 $Y2=0.34
r181 40 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.69 $Y=0.425
+ $X2=4.775 $Y2=0.34
r182 40 41 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=4.69 $Y=0.425
+ $X2=4.69 $Y2=0.895
r183 38 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.605 $Y=0.98
+ $X2=4.69 $Y2=0.895
r184 38 39 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.605 $Y=0.98
+ $X2=3.935 $Y2=0.98
r185 37 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.85 $Y=0.895
+ $X2=3.935 $Y2=0.98
r186 36 37 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=3.85 $Y=0.44
+ $X2=3.85 $Y2=0.895
r187 34 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.765 $Y=0.355
+ $X2=3.85 $Y2=0.44
r188 34 35 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=3.765 $Y=0.355
+ $X2=2.975 $Y2=0.355
r189 32 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.89 $Y=0.44
+ $X2=2.975 $Y2=0.355
r190 32 33 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=2.89 $Y=0.44
+ $X2=2.89 $Y2=1.065
r191 31 50 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.575 $Y=1.15
+ $X2=2.41 $Y2=1.15
r192 30 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.805 $Y=1.15
+ $X2=2.89 $Y2=1.065
r193 30 31 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=2.805 $Y=1.15
+ $X2=2.575 $Y2=1.15
r194 27 29 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.85 $Y=2.77
+ $X2=3.85 $Y2=2.485
r195 25 27 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.85 $Y=2.86 $X2=3.85
+ $Y2=2.77
r196 25 26 83.5726 $w=1.8e-07 $l=2.15e-07 $layer=POLY_cond $X=3.85 $Y=2.86
+ $X2=3.85 $Y2=3.075
r197 22 24 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=3.095 $Y=1.045
+ $X2=3.095 $Y2=0.645
r198 21 61 28.4889 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=2.575 $Y=1.12
+ $X2=2.352 $Y2=1.12
r199 20 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.02 $Y=1.12
+ $X2=3.095 $Y2=1.045
r200 20 21 228.181 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=3.02 $Y=1.12
+ $X2=2.575 $Y2=1.12
r201 18 26 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=3.76 $Y=3.15
+ $X2=3.85 $Y2=3.075
r202 18 19 743.511 $w=1.5e-07 $l=1.45e-06 $layer=POLY_cond $X=3.76 $Y=3.15
+ $X2=2.31 $Y2=3.15
r203 15 19 26.9307 $w=1.5e-07 $l=1.53542e-07 $layer=POLY_cond $X=2.22 $Y=3.035
+ $X2=2.31 $Y2=3.15
r204 15 17 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.22 $Y=3.035
+ $X2=2.22 $Y2=2.54
r205 14 17 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.22 $Y=2.045
+ $X2=2.22 $Y2=2.54
r206 13 14 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.22 $Y=1.955
+ $X2=2.22 $Y2=2.045
r207 13 65 180.75 $w=1.8e-07 $l=4.65e-07 $layer=POLY_cond $X=2.22 $Y=1.955
+ $X2=2.22 $Y2=1.49
r208 10 65 29.7069 $w=4.45e-07 $l=7.5e-08 $layer=POLY_cond $X=2.352 $Y=1.415
+ $X2=2.352 $Y2=1.49
r209 10 54 23.121 $w=4.45e-07 $l=1.85e-07 $layer=POLY_cond $X=2.352 $Y=1.415
+ $X2=2.352 $Y2=1.23
r210 10 11 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=2.13 $Y=1.415
+ $X2=1.77 $Y2=1.415
r211 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.695 $Y=1.34
+ $X2=1.77 $Y2=1.415
r212 7 9 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.695 $Y=1.34
+ $X2=1.695 $Y2=0.895
r213 2 57 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=5.46
+ $Y=1.84 $X2=5.605 $Y2=1.985
r214 1 47 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=5.525
+ $Y=0.37 $X2=5.67 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__SDLCLKP_4%A_792_48# 1 2 9 12 13 15 18 20 22 23 26 29
+ 32 33 36 37 39 43 49 50 52 58
c127 23 0 6.61483e-20 $X=4.88 $Y=1.82
c128 20 0 1.06371e-19 $X=7.015 $Y=1.765
c129 9 0 1.23505e-19 $X=4.035 $Y=0.58
r130 52 54 10.9068 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=5.11 $Y=0.83
+ $X2=5.11 $Y2=1.065
r131 44 58 25.3549 $w=3.3e-07 $l=1.45e-07 $layer=POLY_cond $X=4.125 $Y=1.74
+ $X2=4.27 $Y2=1.74
r132 44 55 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.125 $Y=1.74
+ $X2=4.035 $Y2=1.74
r133 43 46 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=4.125 $Y=1.74
+ $X2=4.125 $Y2=1.82
r134 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.125
+ $Y=1.74 $X2=4.125 $Y2=1.74
r135 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.865
+ $Y=1.465 $X2=6.865 $Y2=1.465
r136 37 39 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=6.455 $Y=1.465
+ $X2=6.865 $Y2=1.465
r137 35 37 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.37 $Y=1.63
+ $X2=6.455 $Y2=1.465
r138 35 36 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=6.37 $Y=1.63
+ $X2=6.37 $Y2=2.24
r139 34 50 4.4465 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=5.27 $Y=2.325
+ $X2=5.075 $Y2=2.325
r140 33 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.285 $Y=2.325
+ $X2=6.37 $Y2=2.24
r141 33 34 66.2193 $w=1.68e-07 $l=1.015e-06 $layer=LI1_cond $X=6.285 $Y=2.325
+ $X2=5.27 $Y2=2.325
r142 32 49 3.351 $w=2.8e-07 $l=1.46458e-07 $layer=LI1_cond $X=5.185 $Y=1.735
+ $X2=5.075 $Y2=1.82
r143 32 54 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.185 $Y=1.735
+ $X2=5.185 $Y2=1.065
r144 27 50 2.47594 $w=3.9e-07 $l=8.5e-08 $layer=LI1_cond $X=5.075 $Y=2.41
+ $X2=5.075 $Y2=2.325
r145 27 29 9.45594 $w=3.88e-07 $l=3.2e-07 $layer=LI1_cond $X=5.075 $Y=2.41
+ $X2=5.075 $Y2=2.73
r146 26 50 2.47594 $w=3.9e-07 $l=8.5e-08 $layer=LI1_cond $X=5.075 $Y=2.24
+ $X2=5.075 $Y2=2.325
r147 25 49 3.351 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=5.075 $Y=1.905
+ $X2=5.075 $Y2=1.82
r148 25 26 9.89919 $w=3.88e-07 $l=3.35e-07 $layer=LI1_cond $X=5.075 $Y=1.905
+ $X2=5.075 $Y2=2.24
r149 24 46 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.29 $Y=1.82
+ $X2=4.125 $Y2=1.82
r150 23 49 3.18746 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=4.88 $Y=1.82
+ $X2=5.075 $Y2=1.82
r151 23 24 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=4.88 $Y=1.82
+ $X2=4.29 $Y2=1.82
r152 20 40 57.8651 $w=3.39e-07 $l=3.51994e-07 $layer=POLY_cond $X=7.015 $Y=1.765
+ $X2=6.902 $Y2=1.465
r153 20 22 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.015 $Y=1.765
+ $X2=7.015 $Y2=2.4
r154 16 40 38.6704 $w=3.39e-07 $l=2.19499e-07 $layer=POLY_cond $X=6.775 $Y=1.3
+ $X2=6.902 $Y2=1.465
r155 16 18 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=6.775 $Y=1.3
+ $X2=6.775 $Y2=0.74
r156 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.27 $Y=2.2 $X2=4.27
+ $Y2=2.485
r157 12 13 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=4.27 $Y=2.11 $X2=4.27
+ $Y2=2.2
r158 11 58 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.27 $Y=1.905
+ $X2=4.27 $Y2=1.74
r159 11 12 79.6855 $w=1.8e-07 $l=2.05e-07 $layer=POLY_cond $X=4.27 $Y=1.905
+ $X2=4.27 $Y2=2.11
r160 7 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.035 $Y=1.575
+ $X2=4.035 $Y2=1.74
r161 7 9 510.202 $w=1.5e-07 $l=9.95e-07 $layer=POLY_cond $X=4.035 $Y=1.575
+ $X2=4.035 $Y2=0.58
r162 2 49 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=4.895
+ $Y=1.755 $X2=5.045 $Y2=1.9
r163 2 29 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=4.895
+ $Y=1.755 $X2=5.045 $Y2=2.73
r164 1 52 182 $w=1.7e-07 $l=5.25357e-07 $layer=licon1_NDIFF $count=1 $X=4.97
+ $Y=0.37 $X2=5.11 $Y2=0.83
.ends

.subckt PM_SKY130_FD_SC_LS__SDLCLKP_4%A_634_74# 1 2 7 9 10 12 14 17 21 26 28 29
c75 26 0 1.23505e-19 $X=3.51 $Y=0.775
r76 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.765
+ $Y=1.4 $X2=4.765 $Y2=1.4
r77 29 32 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=4.765 $Y=1.32 $X2=4.765
+ $Y2=1.4
r78 24 26 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=3.33 $Y=0.775
+ $X2=3.51 $Y2=0.775
r79 22 28 2.36881 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=3.705 $Y=1.32
+ $X2=3.565 $Y2=1.32
r80 21 29 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.6 $Y=1.32
+ $X2=4.765 $Y2=1.32
r81 21 22 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=4.6 $Y=1.32
+ $X2=3.705 $Y2=1.32
r82 17 19 21.4025 $w=2.78e-07 $l=5.2e-07 $layer=LI1_cond $X=3.565 $Y=2.07
+ $X2=3.565 $Y2=2.59
r83 15 28 4.06715 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=3.565 $Y=1.405
+ $X2=3.565 $Y2=1.32
r84 15 17 27.3705 $w=2.78e-07 $l=6.65e-07 $layer=LI1_cond $X=3.565 $Y=1.405
+ $X2=3.565 $Y2=2.07
r85 14 28 4.06715 $w=2.25e-07 $l=1.09087e-07 $layer=LI1_cond $X=3.51 $Y=1.235
+ $X2=3.565 $Y2=1.32
r86 13 26 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.51 $Y=0.94
+ $X2=3.51 $Y2=0.775
r87 13 14 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.51 $Y=0.94
+ $X2=3.51 $Y2=1.235
r88 10 33 38.5495 $w=3.2e-07 $l=2.13014e-07 $layer=POLY_cond $X=4.895 $Y=1.235
+ $X2=4.785 $Y2=1.4
r89 10 12 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=4.895 $Y=1.235
+ $X2=4.895 $Y2=0.74
r90 7 33 55.8714 $w=3.2e-07 $l=2.96985e-07 $layer=POLY_cond $X=4.82 $Y=1.68
+ $X2=4.785 $Y2=1.4
r91 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.82 $Y=1.68 $X2=4.82
+ $Y2=2.315
r92 2 19 600 $w=1.7e-07 $l=7.66339e-07 $layer=licon1_PDIFF $count=1 $X=3.39
+ $Y=1.895 $X2=3.54 $Y2=2.59
r93 2 17 600 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=1 $X=3.39
+ $Y=1.895 $X2=3.54 $Y2=2.07
r94 1 24 182 $w=1.7e-07 $l=4.78357e-07 $layer=licon1_NDIFF $count=1 $X=3.17
+ $Y=0.37 $X2=3.33 $Y2=0.775
.ends

.subckt PM_SKY130_FD_SC_LS__SDLCLKP_4%CLK 1 3 4 6 7 9 10 12 13 20
c53 13 0 1.06371e-19 $X=6 $Y=1.295
c54 10 0 2.38878e-19 $X=6.385 $Y=1.22
c55 1 0 1.06701e-19 $X=5.835 $Y=1.765
r56 20 21 1.65068 $w=4.38e-07 $l=1.5e-08 $layer=POLY_cond $X=6.37 $Y=1.492
+ $X2=6.385 $Y2=1.492
r57 18 20 46.2192 $w=4.38e-07 $l=4.2e-07 $layer=POLY_cond $X=5.95 $Y=1.492
+ $X2=6.37 $Y2=1.492
r58 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.95
+ $Y=1.385 $X2=5.95 $Y2=1.385
r59 16 18 7.15297 $w=4.38e-07 $l=6.5e-08 $layer=POLY_cond $X=5.885 $Y=1.492
+ $X2=5.95 $Y2=1.492
r60 15 16 5.50228 $w=4.38e-07 $l=5e-08 $layer=POLY_cond $X=5.835 $Y=1.492
+ $X2=5.885 $Y2=1.492
r61 13 19 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=5.95 $Y=1.295 $X2=5.95
+ $Y2=1.385
r62 10 21 28.0956 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=6.385 $Y=1.22
+ $X2=6.385 $Y2=1.492
r63 10 12 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=6.385 $Y=1.22
+ $X2=6.385 $Y2=0.74
r64 7 20 28.0956 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=6.37 $Y=1.765
+ $X2=6.37 $Y2=1.492
r65 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.37 $Y=1.765
+ $X2=6.37 $Y2=2.4
r66 4 16 28.0956 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=5.885 $Y=1.22
+ $X2=5.885 $Y2=1.492
r67 4 6 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.885 $Y=1.22 $X2=5.885
+ $Y2=0.74
r68 1 15 28.0956 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=5.835 $Y=1.765
+ $X2=5.835 $Y2=1.492
r69 1 3 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=5.835 $Y=1.765
+ $X2=5.835 $Y2=2.26
.ends

.subckt PM_SKY130_FD_SC_LS__SDLCLKP_4%A_1289_368# 1 2 7 9 12 14 16 19 21 23 26
+ 28 30 33 37 43 45 46 47 48 50 52 58 61 70
c123 33 0 1.19111e-20 $X=9.105 $Y=0.74
r124 70 71 1.87792 $w=3.85e-07 $l=1.5e-08 $layer=POLY_cond $X=9.09 $Y=1.532
+ $X2=9.105 $Y2=1.532
r125 69 70 51.9558 $w=3.85e-07 $l=4.15e-07 $layer=POLY_cond $X=8.675 $Y=1.532
+ $X2=9.09 $Y2=1.532
r126 68 69 10.0156 $w=3.85e-07 $l=8e-08 $layer=POLY_cond $X=8.595 $Y=1.532
+ $X2=8.675 $Y2=1.532
r127 65 66 18.7792 $w=3.85e-07 $l=1.5e-07 $layer=POLY_cond $X=8.095 $Y=1.532
+ $X2=8.245 $Y2=1.532
r128 64 65 41.3143 $w=3.85e-07 $l=3.3e-07 $layer=POLY_cond $X=7.765 $Y=1.532
+ $X2=8.095 $Y2=1.532
r129 59 68 40.6883 $w=3.85e-07 $l=3.25e-07 $layer=POLY_cond $X=8.27 $Y=1.532
+ $X2=8.595 $Y2=1.532
r130 59 66 3.12987 $w=3.85e-07 $l=2.5e-08 $layer=POLY_cond $X=8.27 $Y=1.532
+ $X2=8.245 $Y2=1.532
r131 58 59 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=8.27
+ $Y=1.465 $X2=8.27 $Y2=1.465
r132 56 64 21.9091 $w=3.85e-07 $l=1.75e-07 $layer=POLY_cond $X=7.59 $Y=1.532
+ $X2=7.765 $Y2=1.532
r133 56 62 9.38961 $w=3.85e-07 $l=7.5e-08 $layer=POLY_cond $X=7.59 $Y=1.532
+ $X2=7.515 $Y2=1.532
r134 55 58 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=7.59 $Y=1.465
+ $X2=8.27 $Y2=1.465
r135 55 56 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=7.59
+ $Y=1.465 $X2=7.59 $Y2=1.465
r136 53 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.535 $Y=1.465
+ $X2=7.45 $Y2=1.465
r137 53 55 1.92074 $w=3.28e-07 $l=5.5e-08 $layer=LI1_cond $X=7.535 $Y=1.465
+ $X2=7.59 $Y2=1.465
r138 51 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.45 $Y=1.63
+ $X2=7.45 $Y2=1.465
r139 51 52 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=7.45 $Y=1.63
+ $X2=7.45 $Y2=1.8
r140 50 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.45 $Y=1.3
+ $X2=7.45 $Y2=1.465
r141 49 50 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=7.45 $Y=1.13
+ $X2=7.45 $Y2=1.3
r142 47 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.365 $Y=1.045
+ $X2=7.45 $Y2=1.13
r143 47 48 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=7.365 $Y=1.045
+ $X2=7.155 $Y2=1.045
r144 45 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.365 $Y=1.885
+ $X2=7.45 $Y2=1.8
r145 45 46 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=7.365 $Y=1.885
+ $X2=6.955 $Y2=1.885
r146 41 48 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.99 $Y=0.96
+ $X2=7.155 $Y2=1.045
r147 41 43 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=6.99 $Y=0.96
+ $X2=6.99 $Y2=0.515
r148 37 39 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=6.79 $Y=1.985
+ $X2=6.79 $Y2=2.815
r149 35 46 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.79 $Y=1.97
+ $X2=6.955 $Y2=1.885
r150 35 37 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=6.79 $Y=1.97
+ $X2=6.79 $Y2=1.985
r151 31 71 24.9301 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=9.105 $Y=1.3
+ $X2=9.105 $Y2=1.532
r152 31 33 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=9.105 $Y=1.3
+ $X2=9.105 $Y2=0.74
r153 28 70 24.9301 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=9.09 $Y=1.765
+ $X2=9.09 $Y2=1.532
r154 28 30 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=9.09 $Y=1.765
+ $X2=9.09 $Y2=2.4
r155 24 69 24.9301 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=8.675 $Y=1.3
+ $X2=8.675 $Y2=1.532
r156 24 26 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=8.675 $Y=1.3
+ $X2=8.675 $Y2=0.74
r157 21 68 24.9301 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=8.595 $Y=1.765
+ $X2=8.595 $Y2=1.532
r158 21 23 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.595 $Y=1.765
+ $X2=8.595 $Y2=2.4
r159 17 66 24.9301 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=8.245 $Y=1.3
+ $X2=8.245 $Y2=1.532
r160 17 19 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=8.245 $Y=1.3
+ $X2=8.245 $Y2=0.74
r161 14 65 24.9301 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=8.095 $Y=1.765
+ $X2=8.095 $Y2=1.532
r162 14 16 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.095 $Y=1.765
+ $X2=8.095 $Y2=2.4
r163 10 64 24.9301 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=7.765 $Y=1.3
+ $X2=7.765 $Y2=1.532
r164 10 12 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=7.765 $Y=1.3
+ $X2=7.765 $Y2=0.74
r165 7 62 24.9301 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=7.515 $Y=1.765
+ $X2=7.515 $Y2=1.532
r166 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.515 $Y=1.765
+ $X2=7.515 $Y2=2.4
r167 2 39 400 $w=1.7e-07 $l=1.13446e-06 $layer=licon1_PDIFF $count=1 $X=6.445
+ $Y=1.84 $X2=6.79 $Y2=2.815
r168 2 37 400 $w=1.7e-07 $l=4.11157e-07 $layer=licon1_PDIFF $count=1 $X=6.445
+ $Y=1.84 $X2=6.79 $Y2=1.985
r169 1 43 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.85
+ $Y=0.37 $X2=6.99 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__SDLCLKP_4%VPWR 1 2 3 4 5 6 7 22 24 28 34 38 42 44 46
+ 51 52 53 55 60 68 77 81 90 97 100 103 107
r108 106 107 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r109 103 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r110 100 101 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r111 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r112 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r113 85 107 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=9.36 $Y2=3.33
r114 85 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=8.4 $Y2=3.33
r115 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r116 82 103 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.485 $Y=3.33
+ $X2=8.36 $Y2=3.33
r117 82 84 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=8.485 $Y=3.33
+ $X2=8.88 $Y2=3.33
r118 81 106 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=9.155 $Y=3.33
+ $X2=9.377 $Y2=3.33
r119 81 84 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=9.155 $Y=3.33
+ $X2=8.88 $Y2=3.33
r120 80 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r121 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r122 77 103 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.235 $Y=3.33
+ $X2=8.36 $Y2=3.33
r123 77 79 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=8.235 $Y=3.33
+ $X2=7.92 $Y2=3.33
r124 76 80 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.92 $Y2=3.33
r125 76 101 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6 $Y2=3.33
r126 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r127 73 100 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.31 $Y=3.33
+ $X2=6.145 $Y2=3.33
r128 73 75 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=6.31 $Y=3.33
+ $X2=6.96 $Y2=3.33
r129 72 101 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=6 $Y2=3.33
r130 71 72 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r131 69 97 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.68 $Y=3.33
+ $X2=4.555 $Y2=3.33
r132 69 71 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=4.68 $Y=3.33
+ $X2=5.04 $Y2=3.33
r133 68 100 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.98 $Y=3.33
+ $X2=6.145 $Y2=3.33
r134 68 71 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=5.98 $Y=3.33
+ $X2=5.04 $Y2=3.33
r135 67 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r136 66 67 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r137 64 67 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=4.08 $Y2=3.33
r138 64 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r139 63 66 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=4.08 $Y2=3.33
r140 63 64 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r141 60 97 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.43 $Y=3.33
+ $X2=4.555 $Y2=3.33
r142 60 66 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=4.43 $Y=3.33
+ $X2=4.08 $Y2=3.33
r143 59 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r144 59 88 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.24 $Y2=3.33
r145 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r146 56 87 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.222 $Y2=3.33
r147 56 58 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=1.2 $Y2=3.33
r148 55 63 8.47627 $w=1.7e-07 $l=3.08e-07 $layer=LI1_cond $X=1.852 $Y=3.33
+ $X2=2.16 $Y2=3.33
r149 55 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r150 55 90 10.7939 $w=6.13e-07 $l=5.55e-07 $layer=LI1_cond $X=1.852 $Y=3.33
+ $X2=1.852 $Y2=2.775
r151 55 58 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.545 $Y=3.33
+ $X2=1.2 $Y2=3.33
r152 53 72 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.8 $Y=3.33
+ $X2=5.04 $Y2=3.33
r153 53 98 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.8 $Y=3.33
+ $X2=4.56 $Y2=3.33
r154 51 75 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=7.125 $Y=3.33
+ $X2=6.96 $Y2=3.33
r155 51 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.125 $Y=3.33
+ $X2=7.29 $Y2=3.33
r156 50 79 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=7.455 $Y=3.33
+ $X2=7.92 $Y2=3.33
r157 50 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.455 $Y=3.33
+ $X2=7.29 $Y2=3.33
r158 46 49 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=9.32 $Y=1.985
+ $X2=9.32 $Y2=2.815
r159 44 106 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=9.32 $Y=3.245
+ $X2=9.377 $Y2=3.33
r160 44 49 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=9.32 $Y=3.245
+ $X2=9.32 $Y2=2.815
r161 40 103 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.36 $Y=3.245
+ $X2=8.36 $Y2=3.33
r162 40 42 43.3319 $w=2.48e-07 $l=9.4e-07 $layer=LI1_cond $X=8.36 $Y=3.245
+ $X2=8.36 $Y2=2.305
r163 36 52 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.29 $Y=3.245
+ $X2=7.29 $Y2=3.33
r164 36 38 32.8272 $w=3.28e-07 $l=9.4e-07 $layer=LI1_cond $X=7.29 $Y=3.245
+ $X2=7.29 $Y2=2.305
r165 32 100 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.145 $Y=3.245
+ $X2=6.145 $Y2=3.33
r166 32 34 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=6.145 $Y=3.245
+ $X2=6.145 $Y2=2.745
r167 28 31 22.5879 $w=2.48e-07 $l=4.9e-07 $layer=LI1_cond $X=4.555 $Y=2.24
+ $X2=4.555 $Y2=2.73
r168 26 97 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.555 $Y=3.245
+ $X2=4.555 $Y2=3.33
r169 26 31 23.7403 $w=2.48e-07 $l=5.15e-07 $layer=LI1_cond $X=4.555 $Y=3.245
+ $X2=4.555 $Y2=2.73
r170 22 87 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.222 $Y2=3.33
r171 22 24 39.2878 $w=3.28e-07 $l=1.125e-06 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.28 $Y2=2.12
r172 7 49 400 $w=1.7e-07 $l=1.04964e-06 $layer=licon1_PDIFF $count=1 $X=9.165
+ $Y=1.84 $X2=9.32 $Y2=2.815
r173 7 46 400 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=1 $X=9.165
+ $Y=1.84 $X2=9.32 $Y2=1.985
r174 6 42 300 $w=1.7e-07 $l=5.34766e-07 $layer=licon1_PDIFF $count=2 $X=8.17
+ $Y=1.84 $X2=8.32 $Y2=2.305
r175 5 38 300 $w=1.7e-07 $l=5.5608e-07 $layer=licon1_PDIFF $count=2 $X=7.09
+ $Y=1.84 $X2=7.29 $Y2=2.305
r176 4 34 600 $w=1.7e-07 $l=1.01573e-06 $layer=licon1_PDIFF $count=1 $X=5.91
+ $Y=1.84 $X2=6.145 $Y2=2.745
r177 3 31 600 $w=1.7e-07 $l=5.6637e-07 $layer=licon1_PDIFF $count=1 $X=4.345
+ $Y=2.275 $X2=4.595 $Y2=2.73
r178 3 28 600 $w=1.7e-07 $l=2.66927e-07 $layer=licon1_PDIFF $count=1 $X=4.345
+ $Y=2.275 $X2=4.595 $Y2=2.24
r179 2 90 600 $w=1.7e-07 $l=8.41071e-07 $layer=licon1_PDIFF $count=1 $X=1.565
+ $Y=2.12 $X2=1.99 $Y2=2.775
r180 1 24 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.975 $X2=0.28 $Y2=2.12
.ends

.subckt PM_SKY130_FD_SC_LS__SDLCLKP_4%A_119_143# 1 2 3 4 15 17 18 22 25 29 32 35
+ 36 38 39
c93 38 0 3.22822e-20 $X=2.525 $Y=0.62
c94 35 0 8.1214e-20 $X=1.655 $Y=2.217
r95 38 39 11.007 $w=5.43e-07 $l=2.2e-07 $layer=LI1_cond $X=2.525 $Y=0.622
+ $X2=2.305 $Y2=0.622
r96 27 29 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=3.09 $Y=2.31 $X2=3.09
+ $Y2=2.07
r97 25 27 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.925 $Y=2.395
+ $X2=3.09 $Y2=2.31
r98 25 35 82.8556 $w=1.68e-07 $l=1.27e-06 $layer=LI1_cond $X=2.925 $Y=2.395
+ $X2=1.655 $Y2=2.395
r99 24 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.655 $Y=0.7 $X2=1.57
+ $Y2=0.7
r100 24 39 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.655 $Y=0.7
+ $X2=2.305 $Y2=0.7
r101 22 35 7.85017 $w=5.23e-07 $l=8.5e-08 $layer=LI1_cond $X=1.57 $Y=2.217
+ $X2=1.655 $Y2=2.217
r102 22 32 9.56863 $w=5.23e-07 $l=4.2e-07 $layer=LI1_cond $X=1.57 $Y=2.217
+ $X2=1.15 $Y2=2.217
r103 21 36 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.57 $Y=0.785
+ $X2=1.57 $Y2=0.7
r104 21 22 76.3316 $w=1.68e-07 $l=1.17e-06 $layer=LI1_cond $X=1.57 $Y=0.785
+ $X2=1.57 $Y2=1.955
r105 17 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.485 $Y=0.7
+ $X2=1.57 $Y2=0.7
r106 17 18 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=1.485 $Y=0.7
+ $X2=0.945 $Y2=0.7
r107 13 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.78 $Y=0.785
+ $X2=0.945 $Y2=0.7
r108 13 15 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=0.78 $Y=0.785
+ $X2=0.78 $Y2=0.99
r109 4 29 300 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=2 $X=2.945
+ $Y=1.895 $X2=3.09 $Y2=2.07
r110 3 32 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=1
+ $Y=1.975 $X2=1.15 $Y2=2.12
r111 2 38 182 $w=1.7e-07 $l=3.3541e-07 $layer=licon1_NDIFF $count=1 $X=2.325
+ $Y=0.37 $X2=2.525 $Y2=0.62
r112 1 15 182 $w=1.7e-07 $l=3.55668e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.715 $X2=0.78 $Y2=0.99
.ends

.subckt PM_SKY130_FD_SC_LS__SDLCLKP_4%GCLK 1 2 3 4 15 21 23 24 25 26 29 35 38 39
+ 40 42
c71 25 0 1.19111e-20 $X=8.725 $Y=1.045
r72 40 45 4.56667 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=8.89 $Y=1.295
+ $X2=8.89 $Y2=1.41
r73 40 42 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=8.89 $Y=1.295
+ $X2=8.89 $Y2=1.045
r74 38 39 3.19717 $w=2.95e-07 $l=1.00995e-07 $layer=LI1_cond $X=8.855 $Y=1.8
+ $X2=8.82 $Y2=1.885
r75 38 45 17.2866 $w=2.58e-07 $l=3.9e-07 $layer=LI1_cond $X=8.855 $Y=1.8
+ $X2=8.855 $Y2=1.41
r76 33 42 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=8.89 $Y=0.96
+ $X2=8.89 $Y2=1.045
r77 33 35 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=8.89 $Y=0.96
+ $X2=8.89 $Y2=0.515
r78 29 31 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=8.82 $Y=1.985
+ $X2=8.82 $Y2=2.815
r79 27 39 3.19717 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=8.82 $Y=1.97
+ $X2=8.82 $Y2=1.885
r80 27 29 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=8.82 $Y=1.97
+ $X2=8.82 $Y2=1.985
r81 25 42 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.725 $Y=1.045
+ $X2=8.89 $Y2=1.045
r82 25 26 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=8.725 $Y=1.045
+ $X2=8.115 $Y2=1.045
r83 23 39 3.3845 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.655 $Y=1.885
+ $X2=8.82 $Y2=1.885
r84 23 24 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=8.655 $Y=1.885
+ $X2=8.035 $Y2=1.885
r85 19 26 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=7.99 $Y=0.96
+ $X2=8.115 $Y2=1.045
r86 19 21 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=7.99 $Y=0.96
+ $X2=7.99 $Y2=0.515
r87 15 17 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=7.87 $Y=1.985
+ $X2=7.87 $Y2=2.815
r88 13 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.87 $Y=1.97
+ $X2=8.035 $Y2=1.885
r89 13 15 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=7.87 $Y=1.97
+ $X2=7.87 $Y2=1.985
r90 4 31 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=8.67
+ $Y=1.84 $X2=8.82 $Y2=2.815
r91 4 29 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=8.67
+ $Y=1.84 $X2=8.82 $Y2=1.985
r92 3 17 400 $w=1.7e-07 $l=1.10618e-06 $layer=licon1_PDIFF $count=1 $X=7.59
+ $Y=1.84 $X2=7.87 $Y2=2.815
r93 3 15 400 $w=1.7e-07 $l=3.44964e-07 $layer=licon1_PDIFF $count=1 $X=7.59
+ $Y=1.84 $X2=7.87 $Y2=1.985
r94 2 35 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.75
+ $Y=0.37 $X2=8.89 $Y2=0.515
r95 1 21 91 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_NDIFF $count=2 $X=7.84
+ $Y=0.37 $X2=8.03 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__SDLCLKP_4%VGND 1 2 3 4 5 6 7 22 24 26 30 34 38 42 44
+ 46 49 50 52 53 54 69 73 78 88 94 97 101
r120 100 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r121 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r122 94 95 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r123 88 91 7.33373 $w=4.38e-07 $l=2.8e-07 $layer=LI1_cond $X=1.345 $Y=0
+ $X2=1.345 $Y2=0.28
r124 88 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r125 85 89 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r126 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r127 82 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0
+ $X2=9.36 $Y2=0
r128 82 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=8.4
+ $Y2=0
r129 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r130 79 97 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.545 $Y=0 $X2=8.42
+ $Y2=0
r131 79 81 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=8.545 $Y=0
+ $X2=8.88 $Y2=0
r132 78 100 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=9.235 $Y=0
+ $X2=9.417 $Y2=0
r133 78 81 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=9.235 $Y=0
+ $X2=8.88 $Y2=0
r134 77 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.4
+ $Y2=0
r135 77 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=7.44
+ $Y2=0
r136 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r137 74 94 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.635 $Y=0 $X2=7.51
+ $Y2=0
r138 74 76 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=7.635 $Y=0
+ $X2=7.92 $Y2=0
r139 73 97 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.295 $Y=0 $X2=8.42
+ $Y2=0
r140 73 76 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=8.295 $Y=0
+ $X2=7.92 $Y2=0
r141 72 95 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=7.44
+ $Y2=0
r142 71 72 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r143 69 94 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.385 $Y=0 $X2=7.51
+ $Y2=0
r144 69 71 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=7.385 $Y=0
+ $X2=6.48 $Y2=0
r145 68 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r146 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6 $Y2=0
r147 64 67 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=4.56 $Y=0 $X2=6
+ $Y2=0
r148 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r149 62 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r150 61 62 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r151 59 62 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=1.68 $Y=0 $X2=4.08
+ $Y2=0
r152 59 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r153 58 61 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=1.68 $Y=0 $X2=4.08
+ $Y2=0
r154 58 59 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r155 56 88 6.36164 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=1.565 $Y=0 $X2=1.345
+ $Y2=0
r156 56 58 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=1.565 $Y=0
+ $X2=1.68 $Y2=0
r157 54 68 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=4.8 $Y=0 $X2=6
+ $Y2=0
r158 54 65 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.8 $Y=0 $X2=4.56
+ $Y2=0
r159 52 67 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=6.005 $Y=0 $X2=6
+ $Y2=0
r160 52 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.005 $Y=0 $X2=6.17
+ $Y2=0
r161 51 71 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=6.335 $Y=0
+ $X2=6.48 $Y2=0
r162 51 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.335 $Y=0 $X2=6.17
+ $Y2=0
r163 49 61 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=4.105 $Y=0 $X2=4.08
+ $Y2=0
r164 49 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.105 $Y=0 $X2=4.27
+ $Y2=0
r165 48 64 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=4.435 $Y=0
+ $X2=4.56 $Y2=0
r166 48 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.435 $Y=0 $X2=4.27
+ $Y2=0
r167 44 100 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=9.36 $Y=0.085
+ $X2=9.417 $Y2=0
r168 44 46 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=9.36 $Y=0.085
+ $X2=9.36 $Y2=0.515
r169 40 97 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.42 $Y=0.085
+ $X2=8.42 $Y2=0
r170 40 42 22.3574 $w=2.48e-07 $l=4.85e-07 $layer=LI1_cond $X=8.42 $Y=0.085
+ $X2=8.42 $Y2=0.57
r171 36 94 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.51 $Y=0.085
+ $X2=7.51 $Y2=0
r172 36 38 22.3574 $w=2.48e-07 $l=4.85e-07 $layer=LI1_cond $X=7.51 $Y=0.085
+ $X2=7.51 $Y2=0.57
r173 32 53 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.17 $Y=0.085
+ $X2=6.17 $Y2=0
r174 32 34 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=6.17 $Y=0.085
+ $X2=6.17 $Y2=0.515
r175 28 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.27 $Y=0.085
+ $X2=4.27 $Y2=0
r176 28 30 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=4.27 $Y=0.085
+ $X2=4.27 $Y2=0.535
r177 27 84 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=0
+ $X2=0.222 $Y2=0
r178 26 88 6.36164 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=1.125 $Y=0 $X2=1.345
+ $Y2=0
r179 26 27 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.125 $Y=0
+ $X2=0.445 $Y2=0
r180 22 84 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.222 $Y2=0
r181 22 24 31.6049 $w=3.28e-07 $l=9.05e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.28 $Y2=0.99
r182 7 46 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.18
+ $Y=0.37 $X2=9.32 $Y2=0.515
r183 6 42 182 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=1 $X=8.32
+ $Y=0.37 $X2=8.46 $Y2=0.57
r184 5 38 182 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_NDIFF $count=1 $X=7.405
+ $Y=0.37 $X2=7.55 $Y2=0.57
r185 4 34 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=5.96
+ $Y=0.37 $X2=6.17 $Y2=0.515
r186 3 30 182 $w=1.7e-07 $l=2.31571e-07 $layer=licon1_NDIFF $count=1 $X=4.11
+ $Y=0.37 $X2=4.27 $Y2=0.535
r187 2 91 182 $w=1.7e-07 $l=5.55743e-07 $layer=licon1_NDIFF $count=1 $X=1.07
+ $Y=0.715 $X2=1.345 $Y2=0.28
r188 1 24 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.715 $X2=0.28 $Y2=0.99
.ends

