* File: sky130_fd_sc_ls__a41oi_2.pex.spice
* Created: Wed Sep  2 10:53:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__A41OI_2%B1 1 3 6 8 10 11 12 18 19
c40 19 0 6.4631e-20 $X=0.92 $Y=1.515
c41 8 0 5.79802e-20 $X=1.005 $Y=1.765
r42 18 20 10.9253 $w=3.75e-07 $l=8.5e-08 $layer=POLY_cond $X=0.92 $Y=1.557
+ $X2=1.005 $Y2=1.557
r43 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.92
+ $Y=1.515 $X2=0.92 $Y2=1.515
r44 16 18 45.6293 $w=3.75e-07 $l=3.55e-07 $layer=POLY_cond $X=0.565 $Y=1.557
+ $X2=0.92 $Y2=1.557
r45 15 16 7.712 $w=3.75e-07 $l=6e-08 $layer=POLY_cond $X=0.505 $Y=1.557
+ $X2=0.565 $Y2=1.557
r46 12 19 5.3602 $w=4.28e-07 $l=2e-07 $layer=LI1_cond $X=0.72 $Y=1.565 $X2=0.92
+ $Y2=1.565
r47 11 12 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.24 $Y=1.565
+ $X2=0.72 $Y2=1.565
r48 8 20 24.2915 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.005 $Y=1.765
+ $X2=1.005 $Y2=1.557
r49 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.005 $Y=1.765
+ $X2=1.005 $Y2=2.4
r50 4 16 24.2915 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.565 $Y=1.35
+ $X2=0.565 $Y2=1.557
r51 4 6 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.565 $Y=1.35
+ $X2=0.565 $Y2=0.79
r52 1 15 24.2915 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=1.557
r53 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__A41OI_2%A1 1 3 6 10 12 14 15 21 22
c66 21 0 5.79802e-20 $X=1.58 $Y=1.515
c67 10 0 1.05836e-19 $X=1.985 $Y=0.74
c68 1 0 6.4631e-20 $X=1.505 $Y=1.765
r69 20 22 60.4365 $w=3.23e-07 $l=4.05e-07 $layer=POLY_cond $X=1.58 $Y=1.557
+ $X2=1.985 $Y2=1.557
r70 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.58
+ $Y=1.515 $X2=1.58 $Y2=1.515
r71 18 20 3.73065 $w=3.23e-07 $l=2.5e-08 $layer=POLY_cond $X=1.555 $Y=1.557
+ $X2=1.58 $Y2=1.557
r72 17 18 7.4613 $w=3.23e-07 $l=5e-08 $layer=POLY_cond $X=1.505 $Y=1.557
+ $X2=1.555 $Y2=1.557
r73 15 21 4.54912 $w=3.78e-07 $l=1.5e-07 $layer=LI1_cond $X=1.605 $Y=1.665
+ $X2=1.605 $Y2=1.515
r74 12 22 38.7988 $w=3.23e-07 $l=3.48827e-07 $layer=POLY_cond $X=2.245 $Y=1.765
+ $X2=1.985 $Y2=1.557
r75 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.245 $Y=1.765
+ $X2=2.245 $Y2=2.4
r76 8 22 20.7134 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.985 $Y=1.35
+ $X2=1.985 $Y2=1.557
r77 8 10 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.985 $Y=1.35
+ $X2=1.985 $Y2=0.74
r78 4 18 20.7134 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.555 $Y=1.35
+ $X2=1.555 $Y2=1.557
r79 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.555 $Y=1.35
+ $X2=1.555 $Y2=0.74
r80 1 17 20.7134 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.505 $Y=1.765
+ $X2=1.505 $Y2=1.557
r81 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.505 $Y=1.765
+ $X2=1.505 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__A41OI_2%A2 1 3 4 6 7 9 10 12 15 16 23
c68 23 0 7.08412e-20 $X=3.17 $Y=1.465
c69 16 0 1.16641e-20 $X=3.6 $Y=1.665
r70 23 25 8.31034 $w=4.35e-07 $l=7.5e-08 $layer=POLY_cond $X=3.17 $Y=1.475
+ $X2=3.245 $Y2=1.475
r71 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.17
+ $Y=1.465 $X2=3.17 $Y2=1.465
r72 21 23 28.2552 $w=4.35e-07 $l=2.55e-07 $layer=POLY_cond $X=2.915 $Y=1.475
+ $X2=3.17 $Y2=1.475
r73 20 21 24.377 $w=4.35e-07 $l=2.2e-07 $layer=POLY_cond $X=2.695 $Y=1.475
+ $X2=2.915 $Y2=1.475
r74 16 24 10.7149 $w=4.78e-07 $l=4.3e-07 $layer=LI1_cond $X=3.6 $Y=1.54 $X2=3.17
+ $Y2=1.54
r75 15 24 1.24592 $w=4.78e-07 $l=5e-08 $layer=LI1_cond $X=3.12 $Y=1.54 $X2=3.17
+ $Y2=1.54
r76 10 25 27.9254 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=3.245 $Y=1.765
+ $X2=3.245 $Y2=1.475
r77 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.245 $Y=1.765
+ $X2=3.245 $Y2=2.4
r78 7 21 27.9254 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.915 $Y=1.185
+ $X2=2.915 $Y2=1.475
r79 7 9 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.915 $Y=1.185
+ $X2=2.915 $Y2=0.74
r80 4 20 27.9254 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.695 $Y=1.765
+ $X2=2.695 $Y2=1.475
r81 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.695 $Y=1.765
+ $X2=2.695 $Y2=2.4
r82 1 20 23.269 $w=4.35e-07 $l=3.80789e-07 $layer=POLY_cond $X=2.485 $Y=1.185
+ $X2=2.695 $Y2=1.475
r83 1 3 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.485 $Y=1.185
+ $X2=2.485 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__A41OI_2%A3 2 3 5 8 10 12 15 17 18 24
c60 18 0 2.26957e-19 $X=4.56 $Y=1.665
c61 10 0 1.16641e-20 $X=4.245 $Y=1.765
r62 24 26 17.9256 $w=2.42e-07 $l=9e-08 $layer=POLY_cond $X=4.245 $Y=1.5
+ $X2=4.335 $Y2=1.5
r63 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.245
+ $Y=1.515 $X2=4.245 $Y2=1.515
r64 22 24 67.719 $w=2.42e-07 $l=3.4e-07 $layer=POLY_cond $X=3.905 $Y=1.5
+ $X2=4.245 $Y2=1.5
r65 18 25 8.44232 $w=4.28e-07 $l=3.15e-07 $layer=LI1_cond $X=4.56 $Y=1.565
+ $X2=4.245 $Y2=1.565
r66 17 25 4.42216 $w=4.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.08 $Y=1.565
+ $X2=4.245 $Y2=1.565
r67 13 26 13.9682 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=4.335 $Y=1.35
+ $X2=4.335 $Y2=1.5
r68 13 15 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.335 $Y=1.35
+ $X2=4.335 $Y2=0.74
r69 10 24 13.9682 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=4.245 $Y=1.765
+ $X2=4.245 $Y2=1.5
r70 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.245 $Y=1.765
+ $X2=4.245 $Y2=2.4
r71 6 22 13.9682 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=3.905 $Y=1.35
+ $X2=3.905 $Y2=1.5
r72 6 8 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.905 $Y=1.35
+ $X2=3.905 $Y2=0.74
r73 3 5 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.695 $Y=1.765
+ $X2=3.695 $Y2=2.4
r74 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.695 $Y=1.675 $X2=3.695
+ $Y2=1.765
r75 1 22 41.8264 $w=2.42e-07 $l=2.1e-07 $layer=POLY_cond $X=3.695 $Y=1.5
+ $X2=3.905 $Y2=1.5
r76 1 2 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=3.695 $Y=1.5
+ $X2=3.695 $Y2=1.675
.ends

.subckt PM_SKY130_FD_SC_LS__A41OI_2%A4 3 5 7 8 10 13 15 16 24
c40 5 0 1.56116e-19 $X=4.78 $Y=1.765
c41 3 0 1.52326e-19 $X=4.765 $Y=0.74
r42 24 25 1.9127 $w=3.78e-07 $l=1.5e-08 $layer=POLY_cond $X=5.23 $Y=1.557
+ $X2=5.245 $Y2=1.557
r43 22 24 17.8519 $w=3.78e-07 $l=1.4e-07 $layer=POLY_cond $X=5.09 $Y=1.557
+ $X2=5.23 $Y2=1.557
r44 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.09
+ $Y=1.515 $X2=5.09 $Y2=1.515
r45 20 22 39.5291 $w=3.78e-07 $l=3.1e-07 $layer=POLY_cond $X=4.78 $Y=1.557
+ $X2=5.09 $Y2=1.557
r46 19 20 1.9127 $w=3.78e-07 $l=1.5e-08 $layer=POLY_cond $X=4.765 $Y=1.557
+ $X2=4.78 $Y2=1.557
r47 16 23 11.5244 $w=4.28e-07 $l=4.3e-07 $layer=LI1_cond $X=5.52 $Y=1.565
+ $X2=5.09 $Y2=1.565
r48 15 23 1.34005 $w=4.28e-07 $l=5e-08 $layer=LI1_cond $X=5.04 $Y=1.565 $X2=5.09
+ $Y2=1.565
r49 11 25 24.4846 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.245 $Y=1.35
+ $X2=5.245 $Y2=1.557
r50 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.245 $Y=1.35
+ $X2=5.245 $Y2=0.74
r51 8 24 24.4846 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=5.23 $Y=1.765
+ $X2=5.23 $Y2=1.557
r52 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.23 $Y=1.765
+ $X2=5.23 $Y2=2.4
r53 5 20 24.4846 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=4.78 $Y=1.765
+ $X2=4.78 $Y2=1.557
r54 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.78 $Y=1.765
+ $X2=4.78 $Y2=2.4
r55 1 19 24.4846 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.765 $Y=1.35
+ $X2=4.765 $Y2=1.557
r56 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.765 $Y=1.35
+ $X2=4.765 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__A41OI_2%A_27_368# 1 2 3 4 5 6 21 25 26 27 28 29 31
+ 32 35 37 41 43 47 49 51 53 59 61 63
r97 51 65 2.71076 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.492 $Y=2.12
+ $X2=5.492 $Y2=2.035
r98 51 53 12.0912 $w=3.03e-07 $l=3.2e-07 $layer=LI1_cond $X=5.492 $Y=2.12
+ $X2=5.492 $Y2=2.44
r99 50 63 9.23004 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=4.67 $Y=2.035
+ $X2=4.487 $Y2=2.035
r100 49 65 4.84748 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=5.34 $Y=2.035
+ $X2=5.492 $Y2=2.035
r101 49 50 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.34 $Y=2.035
+ $X2=4.67 $Y2=2.035
r102 45 63 1.2012 $w=3.65e-07 $l=8.5e-08 $layer=LI1_cond $X=4.487 $Y=2.12
+ $X2=4.487 $Y2=2.035
r103 45 47 10.1036 $w=3.63e-07 $l=3.2e-07 $layer=LI1_cond $X=4.487 $Y=2.12
+ $X2=4.487 $Y2=2.44
r104 44 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.635 $Y=2.035
+ $X2=3.47 $Y2=2.035
r105 43 63 9.23004 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=4.305 $Y=2.035
+ $X2=4.487 $Y2=2.035
r106 43 44 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.305 $Y=2.035
+ $X2=3.635 $Y2=2.035
r107 39 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.47 $Y=2.12
+ $X2=3.47 $Y2=2.035
r108 39 41 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=3.47 $Y=2.12
+ $X2=3.47 $Y2=2.815
r109 38 58 4.70058 $w=1.7e-07 $l=1.94808e-07 $layer=LI1_cond $X=2.635 $Y=2.035
+ $X2=2.47 $Y2=1.97
r110 37 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.305 $Y=2.035
+ $X2=3.47 $Y2=2.035
r111 37 38 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.305 $Y=2.035
+ $X2=2.635 $Y2=2.035
r112 33 59 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.47 $Y=2.46
+ $X2=2.47 $Y2=2.375
r113 33 35 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=2.47 $Y=2.46
+ $X2=2.47 $Y2=2.815
r114 32 59 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.47 $Y=2.29
+ $X2=2.47 $Y2=2.375
r115 31 58 3.0656 $w=3.3e-07 $l=1.5e-07 $layer=LI1_cond $X=2.47 $Y=2.12 $X2=2.47
+ $Y2=1.97
r116 31 32 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=2.47 $Y=2.12
+ $X2=2.47 $Y2=2.29
r117 30 56 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.445 $Y=2.375
+ $X2=1.28 $Y2=2.375
r118 29 59 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.305 $Y=2.375
+ $X2=2.47 $Y2=2.375
r119 29 30 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=2.305 $Y=2.375
+ $X2=1.445 $Y2=2.375
r120 27 56 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.28 $Y=2.46 $X2=1.28
+ $Y2=2.375
r121 27 28 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=1.28 $Y=2.46
+ $X2=1.28 $Y2=2.905
r122 25 28 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.115 $Y=2.99
+ $X2=1.28 $Y2=2.905
r123 25 26 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.115 $Y=2.99
+ $X2=0.445 $Y2=2.99
r124 21 24 27.0649 $w=3.28e-07 $l=7.75e-07 $layer=LI1_cond $X=0.28 $Y=2.04
+ $X2=0.28 $Y2=2.815
r125 19 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=2.905
+ $X2=0.445 $Y2=2.99
r126 19 24 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.28 $Y=2.905
+ $X2=0.28 $Y2=2.815
r127 6 65 600 $w=1.7e-07 $l=2.63106e-07 $layer=licon1_PDIFF $count=1 $X=5.305
+ $Y=1.84 $X2=5.465 $Y2=2.035
r128 6 53 300 $w=1.7e-07 $l=6.75278e-07 $layer=licon1_PDIFF $count=2 $X=5.305
+ $Y=1.84 $X2=5.465 $Y2=2.44
r129 5 63 600 $w=1.7e-07 $l=2.64953e-07 $layer=licon1_PDIFF $count=1 $X=4.32
+ $Y=1.84 $X2=4.485 $Y2=2.035
r130 5 47 300 $w=1.7e-07 $l=6.77495e-07 $layer=licon1_PDIFF $count=2 $X=4.32
+ $Y=1.84 $X2=4.485 $Y2=2.44
r131 4 61 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=3.32
+ $Y=1.84 $X2=3.47 $Y2=2.115
r132 4 41 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=3.32
+ $Y=1.84 $X2=3.47 $Y2=2.815
r133 3 58 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.32
+ $Y=1.84 $X2=2.47 $Y2=1.985
r134 3 35 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.32
+ $Y=1.84 $X2=2.47 $Y2=2.815
r135 2 56 300 $w=1.7e-07 $l=6.62495e-07 $layer=licon1_PDIFF $count=2 $X=1.08
+ $Y=1.84 $X2=1.28 $Y2=2.41
r136 1 24 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r137 1 21 400 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.04
.ends

.subckt PM_SKY130_FD_SC_LS__A41OI_2%Y 1 2 3 12 16 17 18 22 25 27 29 30 33 35
r67 33 35 1.30115 $w=3.08e-07 $l=3.5e-08 $layer=LI1_cond $X=2.12 $Y=1.26
+ $X2=2.12 $Y2=1.295
r68 30 33 2.40394 $w=2.03e-07 $l=4e-08 $layer=LI1_cond $X=2.16 $Y=1.135 $X2=2.12
+ $Y2=1.135
r69 30 35 0.92939 $w=3.08e-07 $l=2.5e-08 $layer=LI1_cond $X=2.12 $Y=1.32
+ $X2=2.12 $Y2=1.295
r70 28 30 6.50573 $w=3.08e-07 $l=1.75e-07 $layer=LI1_cond $X=2.12 $Y=1.495
+ $X2=2.12 $Y2=1.32
r71 28 29 8.09553 $w=3.08e-07 $l=1.55e-07 $layer=LI1_cond $X=2.12 $Y=1.495
+ $X2=2.12 $Y2=1.65
r72 25 29 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=2.05 $Y=1.95 $X2=2.05
+ $Y2=1.65
r73 20 33 18.6305 $w=2.03e-07 $l=3.1e-07 $layer=LI1_cond $X=1.81 $Y=1.135
+ $X2=2.12 $Y2=1.135
r74 20 22 11.5244 $w=2.48e-07 $l=2.5e-07 $layer=LI1_cond $X=1.81 $Y=1.01
+ $X2=1.81 $Y2=0.76
r75 19 27 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=2.035
+ $X2=0.78 $Y2=2.035
r76 18 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.965 $Y=2.035
+ $X2=2.05 $Y2=1.95
r77 18 19 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=1.965 $Y=2.035
+ $X2=0.945 $Y2=2.035
r78 16 20 7.87053 $w=2.03e-07 $l=1.43614e-07 $layer=LI1_cond $X=1.685 $Y=1.095
+ $X2=1.81 $Y2=1.135
r79 16 17 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=1.685 $Y=1.095
+ $X2=0.945 $Y2=1.095
r80 10 17 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.78 $Y=1.01
+ $X2=0.945 $Y2=1.095
r81 10 12 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=0.78 $Y=1.01
+ $X2=0.78 $Y2=0.565
r82 3 27 300 $w=1.7e-07 $l=3.61421e-07 $layer=licon1_PDIFF $count=2 $X=0.58
+ $Y=1.84 $X2=0.78 $Y2=2.115
r83 2 22 182 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_NDIFF $count=1 $X=1.63
+ $Y=0.37 $X2=1.77 $Y2=0.76
r84 1 12 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.64
+ $Y=0.42 $X2=0.78 $Y2=0.565
.ends

.subckt PM_SKY130_FD_SC_LS__A41OI_2%VPWR 1 2 3 4 15 19 23 27 30 31 33 34 35 37
+ 49 55 56 59 62
r74 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r75 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r76 56 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=5.04 $Y2=3.33
r77 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r78 53 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.17 $Y=3.33
+ $X2=5.005 $Y2=3.33
r79 53 55 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=5.17 $Y=3.33
+ $X2=5.52 $Y2=3.33
r80 52 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r81 51 52 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r82 49 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.84 $Y=3.33
+ $X2=5.005 $Y2=3.33
r83 49 51 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=4.84 $Y=3.33
+ $X2=4.56 $Y2=3.33
r84 48 52 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r85 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r86 45 60 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=1.68 $Y2=3.33
r87 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r88 42 59 11.5608 $w=1.7e-07 $l=2.6e-07 $layer=LI1_cond $X=2.135 $Y=3.33
+ $X2=1.875 $Y2=3.33
r89 42 44 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=2.135 $Y=3.33
+ $X2=2.64 $Y2=3.33
r90 40 60 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.68 $Y2=3.33
r91 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r92 37 59 11.5608 $w=1.7e-07 $l=2.6e-07 $layer=LI1_cond $X=1.615 $Y=3.33
+ $X2=1.875 $Y2=3.33
r93 37 39 89.7059 $w=1.68e-07 $l=1.375e-06 $layer=LI1_cond $X=1.615 $Y=3.33
+ $X2=0.24 $Y2=3.33
r94 35 48 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=3.6 $Y2=3.33
r95 35 45 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=2.64 $Y2=3.33
r96 33 47 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=3.805 $Y=3.33
+ $X2=3.6 $Y2=3.33
r97 33 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.805 $Y=3.33
+ $X2=3.97 $Y2=3.33
r98 32 51 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=4.135 $Y=3.33
+ $X2=4.56 $Y2=3.33
r99 32 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.135 $Y=3.33
+ $X2=3.97 $Y2=3.33
r100 30 44 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.805 $Y=3.33
+ $X2=2.64 $Y2=3.33
r101 30 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.805 $Y=3.33
+ $X2=2.97 $Y2=3.33
r102 29 47 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=3.135 $Y=3.33
+ $X2=3.6 $Y2=3.33
r103 29 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.135 $Y=3.33
+ $X2=2.97 $Y2=3.33
r104 25 62 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.005 $Y=3.245
+ $X2=5.005 $Y2=3.33
r105 25 27 29.1603 $w=3.28e-07 $l=8.35e-07 $layer=LI1_cond $X=5.005 $Y=3.245
+ $X2=5.005 $Y2=2.41
r106 21 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.97 $Y=3.245
+ $X2=3.97 $Y2=3.33
r107 21 23 29.1603 $w=3.28e-07 $l=8.35e-07 $layer=LI1_cond $X=3.97 $Y=3.245
+ $X2=3.97 $Y2=2.41
r108 17 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.97 $Y=3.245
+ $X2=2.97 $Y2=3.33
r109 17 19 29.1603 $w=3.28e-07 $l=8.35e-07 $layer=LI1_cond $X=2.97 $Y=3.245
+ $X2=2.97 $Y2=2.41
r110 13 59 2.17428 $w=5.2e-07 $l=8.5e-08 $layer=LI1_cond $X=1.875 $Y=3.245
+ $X2=1.875 $Y2=3.33
r111 13 15 10.6957 $w=5.18e-07 $l=4.65e-07 $layer=LI1_cond $X=1.875 $Y=3.245
+ $X2=1.875 $Y2=2.78
r112 4 27 300 $w=1.7e-07 $l=6.40625e-07 $layer=licon1_PDIFF $count=2 $X=4.855
+ $Y=1.84 $X2=5.005 $Y2=2.41
r113 3 23 300 $w=1.7e-07 $l=6.62495e-07 $layer=licon1_PDIFF $count=2 $X=3.77
+ $Y=1.84 $X2=3.97 $Y2=2.41
r114 2 19 300 $w=1.7e-07 $l=6.62495e-07 $layer=licon1_PDIFF $count=2 $X=2.77
+ $Y=1.84 $X2=2.97 $Y2=2.41
r115 1 15 600 $w=1.7e-07 $l=1.07745e-06 $layer=licon1_PDIFF $count=1 $X=1.58
+ $Y=1.84 $X2=1.875 $Y2=2.78
.ends

.subckt PM_SKY130_FD_SC_LS__A41OI_2%VGND 1 2 7 9 13 15 17 27 28 34
r53 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r54 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r55 28 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r56 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r57 25 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.145 $Y=0 $X2=4.98
+ $Y2=0
r58 25 27 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=5.145 $Y=0 $X2=5.52
+ $Y2=0
r59 24 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r60 23 24 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r61 21 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r62 20 23 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=0.72 $Y=0 $X2=4.56
+ $Y2=0
r63 20 21 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=0.72 $Y=0
+ $X2=0.72 $Y2=0
r64 18 31 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.222
+ $Y2=0
r65 18 20 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.72
+ $Y2=0
r66 17 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.815 $Y=0 $X2=4.98
+ $Y2=0
r67 17 23 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=4.815 $Y=0 $X2=4.56
+ $Y2=0
r68 15 24 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=2.88 $Y=0 $X2=4.56
+ $Y2=0
r69 15 21 0.602067 $w=4.9e-07 $l=2.16e-06 $layer=MET1_cond $X=2.88 $Y=0 $X2=0.72
+ $Y2=0
r70 11 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.98 $Y=0.085
+ $X2=4.98 $Y2=0
r71 11 13 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=4.98 $Y=0.085
+ $X2=4.98 $Y2=0.675
r72 7 31 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.222 $Y2=0
r73 7 9 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.28 $Y=0.085 $X2=0.28
+ $Y2=0.565
r74 2 13 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=4.84
+ $Y=0.37 $X2=4.98 $Y2=0.675
r75 1 9 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.42 $X2=0.28 $Y2=0.565
.ends

.subckt PM_SKY130_FD_SC_LS__A41OI_2%A_239_74# 1 2 3 12 14 15 17 20 24
r44 24 27 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=3.13 $Y=0.835 $X2=3.13
+ $Y2=0.915
r45 21 23 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.355 $Y=0.835
+ $X2=2.23 $Y2=0.835
r46 20 24 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.965 $Y=0.835
+ $X2=3.13 $Y2=0.835
r47 20 21 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=2.965 $Y=0.835
+ $X2=2.355 $Y2=0.835
r48 17 23 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.23 $Y=0.75 $X2=2.23
+ $Y2=0.835
r49 17 19 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=2.23 $Y=0.75
+ $X2=2.23 $Y2=0.495
r50 16 19 3.22684 $w=2.48e-07 $l=7e-08 $layer=LI1_cond $X=2.23 $Y=0.425 $X2=2.23
+ $Y2=0.495
r51 14 16 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.105 $Y=0.34
+ $X2=2.23 $Y2=0.425
r52 14 15 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=2.105 $Y=0.34
+ $X2=1.505 $Y2=0.34
r53 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.34 $Y=0.425
+ $X2=1.505 $Y2=0.34
r54 10 12 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=1.34 $Y=0.425
+ $X2=1.34 $Y2=0.675
r55 3 27 182 $w=1.7e-07 $l=6.11003e-07 $layer=licon1_NDIFF $count=1 $X=2.99
+ $Y=0.37 $X2=3.13 $Y2=0.915
r56 2 23 182 $w=1.7e-07 $l=5.60245e-07 $layer=licon1_NDIFF $count=1 $X=2.06
+ $Y=0.37 $X2=2.27 $Y2=0.835
r57 2 19 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=2.06
+ $Y=0.37 $X2=2.27 $Y2=0.495
r58 1 12 182 $w=1.7e-07 $l=3.70473e-07 $layer=licon1_NDIFF $count=1 $X=1.195
+ $Y=0.37 $X2=1.34 $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_LS__A41OI_2%A_512_74# 1 2 12 13
c21 13 0 1.05836e-19 $X=3.955 $Y=0.505
c22 12 0 1.52326e-19 $X=4.12 $Y=0.515
r23 12 13 6.3908 $w=3.48e-07 $l=1.65e-07 $layer=LI1_cond $X=4.12 $Y=0.505
+ $X2=3.955 $Y2=0.505
r24 9 13 57.8526 $w=2.48e-07 $l=1.255e-06 $layer=LI1_cond $X=2.7 $Y=0.455
+ $X2=3.955 $Y2=0.455
r25 2 12 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.98
+ $Y=0.37 $X2=4.12 $Y2=0.515
r26 1 9 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=2.56
+ $Y=0.37 $X2=2.7 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LS__A41OI_2%A_709_74# 1 2 3 10 16 18 22 25
r37 20 22 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=5.48 $Y=1.01
+ $X2=5.48 $Y2=0.515
r38 19 25 4.06715 $w=2.25e-07 $l=1.18427e-07 $layer=LI1_cond $X=4.635 $Y=1.095
+ $X2=4.55 $Y2=1.015
r39 18 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.315 $Y=1.095
+ $X2=5.48 $Y2=1.01
r40 18 19 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=5.315 $Y=1.095
+ $X2=4.635 $Y2=1.095
r41 14 25 2.36881 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.55 $Y=0.85
+ $X2=4.55 $Y2=1.015
r42 14 16 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=4.55 $Y=0.85
+ $X2=4.55 $Y2=0.515
r43 10 25 4.06715 $w=2.25e-07 $l=9.66954e-08 $layer=LI1_cond $X=4.465 $Y=0.99
+ $X2=4.55 $Y2=1.015
r44 10 12 31.898 $w=2.78e-07 $l=7.75e-07 $layer=LI1_cond $X=4.465 $Y=0.99
+ $X2=3.69 $Y2=0.99
r45 3 22 91 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=2 $X=5.32
+ $Y=0.37 $X2=5.48 $Y2=0.515
r46 2 25 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=4.41
+ $Y=0.37 $X2=4.55 $Y2=0.965
r47 2 16 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=4.41
+ $Y=0.37 $X2=4.55 $Y2=0.515
r48 1 12 182 $w=1.7e-07 $l=6.4846e-07 $layer=licon1_NDIFF $count=1 $X=3.545
+ $Y=0.37 $X2=3.69 $Y2=0.95
.ends

