* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__dlclkp_2 CLK GATE VGND VNB VPB VPWR GCLK
M1000 VPWR CLK a_315_48# VPB phighvt w=840000u l=150000u
+  ad=2.6426e+12p pd=1.594e+07u as=2.646e+11p ps=2.31e+06u
M1001 a_83_244# a_315_338# a_264_392# VPB phighvt w=1e+06u l=150000u
+  ad=4.267e+11p pd=3.3e+06u as=2.7e+11p ps=2.54e+06u
M1002 GCLK a_1041_387# VGND VNB nshort w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=1.45355e+12p ps=1.19e+07u
M1003 a_315_338# a_315_48# VPWR VPB phighvt w=840000u l=150000u
+  ad=2.478e+11p pd=2.27e+06u as=0p ps=0u
M1004 a_1041_387# CLK VPWR VPB phighvt w=1e+06u l=150000u
+  ad=3.25e+11p pd=2.65e+06u as=0p ps=0u
M1005 a_264_392# GATE VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_494_118# a_315_338# a_83_244# VNB nshort w=420000u l=150000u
+  ad=1.54875e+11p pd=1.7e+06u as=3.049e+11p ps=2.47e+06u
M1007 VGND a_1041_387# GCLK VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND a_27_74# a_494_118# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_315_338# a_315_48# VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1010 GCLK a_1041_387# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=0p ps=0u
M1011 VPWR a_83_244# a_27_74# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.304e+11p ps=2.83e+06u
M1012 a_267_74# GATE VGND VNB nshort w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1013 a_83_244# a_315_48# a_267_74# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND CLK a_315_48# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1015 a_1041_387# a_27_74# a_1044_119# VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=1.554e+11p ps=1.9e+06u
M1016 VPWR a_27_74# a_508_508# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1017 VPWR a_1041_387# GCLK VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND a_83_244# a_27_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1019 a_1044_119# CLK VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_508_508# a_315_48# a_83_244# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPWR a_27_74# a_1041_387# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
