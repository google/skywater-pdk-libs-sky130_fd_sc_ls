* File: sky130_fd_sc_ls__sdfxbp_2.pxi.spice
* Created: Wed Sep  2 11:28:20 2020
* 
x_PM_SKY130_FD_SC_LS__SDFXBP_2%A_36_74# N_A_36_74#_M1032_s N_A_36_74#_M1023_s
+ N_A_36_74#_M1012_g N_A_36_74#_c_273_n N_A_36_74#_M1006_g N_A_36_74#_c_269_n
+ N_A_36_74#_c_270_n N_A_36_74#_c_275_n N_A_36_74#_c_276_n N_A_36_74#_c_277_n
+ N_A_36_74#_c_278_n N_A_36_74#_c_271_n N_A_36_74#_c_272_n N_A_36_74#_c_280_n
+ PM_SKY130_FD_SC_LS__SDFXBP_2%A_36_74#
x_PM_SKY130_FD_SC_LS__SDFXBP_2%SCE N_SCE_c_352_n N_SCE_c_360_n N_SCE_c_361_n
+ N_SCE_c_353_n N_SCE_M1032_g N_SCE_c_362_n N_SCE_M1023_g N_SCE_c_363_n
+ N_SCE_c_364_n N_SCE_M1030_g N_SCE_c_354_n N_SCE_M1026_g N_SCE_c_365_n
+ N_SCE_c_355_n N_SCE_c_356_n SCE N_SCE_c_357_n N_SCE_c_358_n
+ PM_SKY130_FD_SC_LS__SDFXBP_2%SCE
x_PM_SKY130_FD_SC_LS__SDFXBP_2%D N_D_M1013_g N_D_c_430_n N_D_c_431_n N_D_M1003_g
+ D N_D_c_428_n N_D_c_429_n PM_SKY130_FD_SC_LS__SDFXBP_2%D
x_PM_SKY130_FD_SC_LS__SDFXBP_2%SCD N_SCD_c_469_n N_SCD_M1027_g N_SCD_M1024_g SCD
+ N_SCD_c_471_n PM_SKY130_FD_SC_LS__SDFXBP_2%SCD
x_PM_SKY130_FD_SC_LS__SDFXBP_2%CLK N_CLK_M1000_g N_CLK_c_504_n N_CLK_M1001_g CLK
+ N_CLK_c_503_n PM_SKY130_FD_SC_LS__SDFXBP_2%CLK
x_PM_SKY130_FD_SC_LS__SDFXBP_2%A_828_74# N_A_828_74#_M1011_d N_A_828_74#_M1031_d
+ N_A_828_74#_c_559_n N_A_828_74#_M1035_g N_A_828_74#_M1028_g
+ N_A_828_74#_c_539_n N_A_828_74#_M1033_g N_A_828_74#_c_560_n
+ N_A_828_74#_c_561_n N_A_828_74#_M1036_g N_A_828_74#_c_540_n
+ N_A_828_74#_c_563_n N_A_828_74#_c_541_n N_A_828_74#_c_542_n
+ N_A_828_74#_c_543_n N_A_828_74#_c_544_n N_A_828_74#_c_545_n
+ N_A_828_74#_c_546_n N_A_828_74#_c_547_n N_A_828_74#_c_616_p
+ N_A_828_74#_c_548_n N_A_828_74#_c_549_n N_A_828_74#_c_550_n
+ N_A_828_74#_c_565_n N_A_828_74#_c_551_n N_A_828_74#_c_552_n
+ N_A_828_74#_c_553_n N_A_828_74#_c_554_n N_A_828_74#_c_555_n
+ N_A_828_74#_c_556_n N_A_828_74#_c_557_n N_A_828_74#_c_558_n
+ PM_SKY130_FD_SC_LS__SDFXBP_2%A_828_74#
x_PM_SKY130_FD_SC_LS__SDFXBP_2%A_630_74# N_A_630_74#_M1000_d N_A_630_74#_M1001_d
+ N_A_630_74#_M1011_g N_A_630_74#_c_738_n N_A_630_74#_c_755_n
+ N_A_630_74#_M1031_g N_A_630_74#_c_739_n N_A_630_74#_M1017_g
+ N_A_630_74#_c_741_n N_A_630_74#_c_758_n N_A_630_74#_c_759_n
+ N_A_630_74#_M1015_g N_A_630_74#_c_760_n N_A_630_74#_M1016_g
+ N_A_630_74#_c_742_n N_A_630_74#_c_743_n N_A_630_74#_M1008_g
+ N_A_630_74#_c_744_n N_A_630_74#_c_745_n N_A_630_74#_c_746_n
+ N_A_630_74#_c_747_n N_A_630_74#_c_763_n N_A_630_74#_c_748_n
+ N_A_630_74#_c_749_n N_A_630_74#_c_781_n N_A_630_74#_c_764_n
+ N_A_630_74#_c_750_n N_A_630_74#_c_766_n N_A_630_74#_c_831_p
+ N_A_630_74#_c_858_p N_A_630_74#_c_767_n N_A_630_74#_c_751_n
+ N_A_630_74#_c_768_n N_A_630_74#_c_752_n N_A_630_74#_c_753_n
+ PM_SKY130_FD_SC_LS__SDFXBP_2%A_630_74#
x_PM_SKY130_FD_SC_LS__SDFXBP_2%A_1243_48# N_A_1243_48#_M1018_d
+ N_A_1243_48#_M1038_d N_A_1243_48#_M1014_g N_A_1243_48#_c_940_n
+ N_A_1243_48#_c_947_n N_A_1243_48#_M1004_g N_A_1243_48#_c_941_n
+ N_A_1243_48#_c_942_n N_A_1243_48#_c_943_n N_A_1243_48#_c_948_n
+ N_A_1243_48#_c_944_n N_A_1243_48#_c_945_n
+ PM_SKY130_FD_SC_LS__SDFXBP_2%A_1243_48#
x_PM_SKY130_FD_SC_LS__SDFXBP_2%A_1021_97# N_A_1021_97#_M1017_d
+ N_A_1021_97#_M1035_d N_A_1021_97#_M1018_g N_A_1021_97#_c_1010_n
+ N_A_1021_97#_M1038_g N_A_1021_97#_c_1011_n N_A_1021_97#_c_1012_n
+ N_A_1021_97#_c_1034_n N_A_1021_97#_c_1013_n N_A_1021_97#_c_1017_n
+ N_A_1021_97#_c_1018_n N_A_1021_97#_c_1014_n
+ PM_SKY130_FD_SC_LS__SDFXBP_2%A_1021_97#
x_PM_SKY130_FD_SC_LS__SDFXBP_2%A_1711_48# N_A_1711_48#_M1025_d
+ N_A_1711_48#_M1007_d N_A_1711_48#_c_1092_n N_A_1711_48#_M1009_g
+ N_A_1711_48#_c_1093_n N_A_1711_48#_c_1094_n N_A_1711_48#_c_1111_n
+ N_A_1711_48#_M1029_g N_A_1711_48#_c_1095_n N_A_1711_48#_c_1096_n
+ N_A_1711_48#_c_1097_n N_A_1711_48#_M1010_g N_A_1711_48#_M1022_g
+ N_A_1711_48#_c_1099_n N_A_1711_48#_c_1100_n N_A_1711_48#_c_1115_n
+ N_A_1711_48#_M1020_g N_A_1711_48#_M1037_g N_A_1711_48#_c_1102_n
+ N_A_1711_48#_c_1103_n N_A_1711_48#_c_1117_n N_A_1711_48#_M1005_g
+ N_A_1711_48#_M1021_g N_A_1711_48#_c_1105_n N_A_1711_48#_c_1106_n
+ N_A_1711_48#_c_1118_n N_A_1711_48#_c_1119_n N_A_1711_48#_c_1107_n
+ N_A_1711_48#_c_1108_n N_A_1711_48#_c_1194_p N_A_1711_48#_c_1109_n
+ N_A_1711_48#_c_1121_n N_A_1711_48#_c_1110_n
+ PM_SKY130_FD_SC_LS__SDFXBP_2%A_1711_48#
x_PM_SKY130_FD_SC_LS__SDFXBP_2%A_1511_74# N_A_1511_74#_M1033_d
+ N_A_1511_74#_M1016_d N_A_1511_74#_M1025_g N_A_1511_74#_c_1256_n
+ N_A_1511_74#_c_1266_n N_A_1511_74#_M1007_g N_A_1511_74#_c_1267_n
+ N_A_1511_74#_c_1268_n N_A_1511_74#_c_1257_n N_A_1511_74#_c_1269_n
+ N_A_1511_74#_c_1270_n N_A_1511_74#_c_1258_n N_A_1511_74#_c_1259_n
+ N_A_1511_74#_c_1260_n N_A_1511_74#_c_1272_n N_A_1511_74#_c_1261_n
+ N_A_1511_74#_c_1262_n N_A_1511_74#_c_1263_n N_A_1511_74#_c_1264_n
+ PM_SKY130_FD_SC_LS__SDFXBP_2%A_1511_74#
x_PM_SKY130_FD_SC_LS__SDFXBP_2%A_2322_368# N_A_2322_368#_M1021_s
+ N_A_2322_368#_M1005_s N_A_2322_368#_c_1372_n N_A_2322_368#_M1002_g
+ N_A_2322_368#_M1019_g N_A_2322_368#_M1039_g N_A_2322_368#_c_1373_n
+ N_A_2322_368#_M1034_g N_A_2322_368#_c_1368_n N_A_2322_368#_c_1374_n
+ N_A_2322_368#_c_1369_n N_A_2322_368#_c_1370_n N_A_2322_368#_c_1371_n
+ PM_SKY130_FD_SC_LS__SDFXBP_2%A_2322_368#
x_PM_SKY130_FD_SC_LS__SDFXBP_2%VPWR N_VPWR_M1023_d N_VPWR_M1027_d N_VPWR_M1031_s
+ N_VPWR_M1004_d N_VPWR_M1029_d N_VPWR_M1010_s N_VPWR_M1020_s N_VPWR_M1005_d
+ N_VPWR_M1034_d N_VPWR_c_1440_n N_VPWR_c_1441_n N_VPWR_c_1442_n N_VPWR_c_1443_n
+ N_VPWR_c_1444_n N_VPWR_c_1445_n N_VPWR_c_1446_n N_VPWR_c_1447_n
+ N_VPWR_c_1448_n N_VPWR_c_1449_n N_VPWR_c_1450_n N_VPWR_c_1451_n
+ N_VPWR_c_1452_n N_VPWR_c_1453_n N_VPWR_c_1454_n N_VPWR_c_1455_n
+ N_VPWR_c_1456_n N_VPWR_c_1457_n N_VPWR_c_1458_n VPWR N_VPWR_c_1459_n
+ N_VPWR_c_1460_n N_VPWR_c_1461_n N_VPWR_c_1462_n N_VPWR_c_1463_n
+ N_VPWR_c_1464_n N_VPWR_c_1465_n N_VPWR_c_1466_n N_VPWR_c_1467_n
+ N_VPWR_c_1439_n PM_SKY130_FD_SC_LS__SDFXBP_2%VPWR
x_PM_SKY130_FD_SC_LS__SDFXBP_2%A_301_74# N_A_301_74#_M1013_d N_A_301_74#_M1017_s
+ N_A_301_74#_M1003_d N_A_301_74#_M1035_s N_A_301_74#_c_1618_n
+ N_A_301_74#_c_1619_n N_A_301_74#_c_1605_n N_A_301_74#_c_1606_n
+ N_A_301_74#_c_1607_n N_A_301_74#_c_1608_n N_A_301_74#_c_1613_n
+ N_A_301_74#_c_1614_n N_A_301_74#_c_1609_n N_A_301_74#_c_1610_n
+ N_A_301_74#_c_1611_n N_A_301_74#_c_1615_n N_A_301_74#_c_1665_n
+ N_A_301_74#_c_1616_n N_A_301_74#_c_1714_n N_A_301_74#_c_1617_n
+ PM_SKY130_FD_SC_LS__SDFXBP_2%A_301_74#
x_PM_SKY130_FD_SC_LS__SDFXBP_2%Q N_Q_M1022_d N_Q_M1010_d N_Q_c_1734_n
+ N_Q_c_1731_n N_Q_c_1736_n Q Q Q PM_SKY130_FD_SC_LS__SDFXBP_2%Q
x_PM_SKY130_FD_SC_LS__SDFXBP_2%Q_N N_Q_N_M1019_d N_Q_N_M1002_s N_Q_N_c_1770_n
+ N_Q_N_c_1772_n Q_N Q_N Q_N PM_SKY130_FD_SC_LS__SDFXBP_2%Q_N
x_PM_SKY130_FD_SC_LS__SDFXBP_2%VGND N_VGND_M1032_d N_VGND_M1024_d N_VGND_M1011_s
+ N_VGND_M1014_d N_VGND_M1009_d N_VGND_M1022_s N_VGND_M1037_s N_VGND_M1021_d
+ N_VGND_M1039_s N_VGND_c_1799_n N_VGND_c_1800_n N_VGND_c_1801_n N_VGND_c_1802_n
+ N_VGND_c_1803_n N_VGND_c_1804_n N_VGND_c_1805_n N_VGND_c_1806_n
+ N_VGND_c_1807_n N_VGND_c_1808_n N_VGND_c_1809_n N_VGND_c_1810_n
+ N_VGND_c_1811_n N_VGND_c_1812_n N_VGND_c_1938_n VGND N_VGND_c_1813_n
+ N_VGND_c_1814_n N_VGND_c_1815_n N_VGND_c_1816_n N_VGND_c_1817_n
+ N_VGND_c_1818_n N_VGND_c_1819_n N_VGND_c_1820_n N_VGND_c_1821_n
+ N_VGND_c_1822_n N_VGND_c_1823_n N_VGND_c_1824_n N_VGND_c_1825_n
+ PM_SKY130_FD_SC_LS__SDFXBP_2%VGND
cc_1 VNB N_A_36_74#_M1012_g 0.0464821f $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=0.58
cc_2 VNB N_A_36_74#_c_269_n 0.0230916f $X=-0.19 $Y=-0.245 $X2=0.965 $Y2=1.635
cc_3 VNB N_A_36_74#_c_270_n 0.027073f $X=-0.19 $Y=-0.245 $X2=0.17 $Y2=1.47
cc_4 VNB N_A_36_74#_c_271_n 0.0193228f $X=-0.19 $Y=-0.245 $X2=0.325 $Y2=0.54
cc_5 VNB N_A_36_74#_c_272_n 0.0100127f $X=-0.19 $Y=-0.245 $X2=0.83 $Y2=1.635
cc_6 VNB N_SCE_c_352_n 0.0257263f $X=-0.19 $Y=-0.245 $X2=0.21 $Y2=2.265
cc_7 VNB N_SCE_c_353_n 0.0221696f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_SCE_c_354_n 0.0191896f $X=-0.19 $Y=-0.245 $X2=0.17 $Y2=1.47
cc_9 VNB N_SCE_c_355_n 0.0530904f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_SCE_c_356_n 0.0533134f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=2.055
cc_11 VNB N_SCE_c_357_n 0.0100347f $X=-0.19 $Y=-0.245 $X2=0.17 $Y2=1.635
cc_12 VNB N_SCE_c_358_n 0.0160413f $X=-0.19 $Y=-0.245 $X2=2.03 $Y2=1.89
cc_13 VNB N_D_M1013_g 0.0520573f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_D_c_428_n 0.0187805f $X=-0.19 $Y=-0.245 $X2=2.04 $Y2=2.585
cc_15 VNB N_D_c_429_n 0.00858587f $X=-0.19 $Y=-0.245 $X2=0.965 $Y2=1.635
cc_16 VNB N_SCD_M1024_g 0.0663333f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_CLK_M1000_g 0.032682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB CLK 0.00268784f $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=0.58
cc_19 VNB N_CLK_c_503_n 0.0435265f $X=-0.19 $Y=-0.245 $X2=2.04 $Y2=2.19
cc_20 VNB N_A_828_74#_M1028_g 0.0210539f $X=-0.19 $Y=-0.245 $X2=2.04 $Y2=2.585
cc_21 VNB N_A_828_74#_c_539_n 0.0177049f $X=-0.19 $Y=-0.245 $X2=0.965 $Y2=1.635
cc_22 VNB N_A_828_74#_c_540_n 0.00573146f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=2.055
cc_23 VNB N_A_828_74#_c_541_n 0.0106507f $X=-0.19 $Y=-0.245 $X2=0.325 $Y2=0.54
cc_24 VNB N_A_828_74#_c_542_n 0.0177202f $X=-0.19 $Y=-0.245 $X2=0.17 $Y2=1.635
cc_25 VNB N_A_828_74#_c_543_n 0.0036407f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_828_74#_c_544_n 0.00611811f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.635
cc_27 VNB N_A_828_74#_c_545_n 0.0175499f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.635
cc_28 VNB N_A_828_74#_c_546_n 4.98048e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_828_74#_c_547_n 0.00755014f $X=-0.19 $Y=-0.245 $X2=2.03 $Y2=1.89
cc_30 VNB N_A_828_74#_c_548_n 0.00453192f $X=-0.19 $Y=-0.245 $X2=2.03 $Y2=2.055
cc_31 VNB N_A_828_74#_c_549_n 0.00181452f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_828_74#_c_550_n 0.00996222f $X=-0.19 $Y=-0.245 $X2=2.03 $Y2=1.89
cc_33 VNB N_A_828_74#_c_551_n 0.00123754f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_828_74#_c_552_n 0.00708924f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_828_74#_c_553_n 0.0333274f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_828_74#_c_554_n 0.00690044f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_828_74#_c_555_n 0.0406871f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_828_74#_c_556_n 8.79381e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_828_74#_c_557_n 0.00265789f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_828_74#_c_558_n 0.0328554f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_630_74#_M1011_g 0.0310251f $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=0.58
cc_42 VNB N_A_630_74#_c_738_n 0.00571277f $X=-0.19 $Y=-0.245 $X2=2.04 $Y2=2.19
cc_43 VNB N_A_630_74#_c_739_n 0.011214f $X=-0.19 $Y=-0.245 $X2=0.17 $Y2=1.47
cc_44 VNB N_A_630_74#_M1017_g 0.0563562f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_630_74#_c_741_n 0.0321584f $X=-0.19 $Y=-0.245 $X2=0.83 $Y2=1.97
cc_46 VNB N_A_630_74#_c_742_n 0.0356248f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.635
cc_47 VNB N_A_630_74#_c_743_n 0.0171287f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.635
cc_48 VNB N_A_630_74#_c_744_n 0.00496867f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_630_74#_c_745_n 7.16371e-19 $X=-0.19 $Y=-0.245 $X2=2.03 $Y2=1.89
cc_50 VNB N_A_630_74#_c_746_n 0.0206099f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_630_74#_c_747_n 0.00956599f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_630_74#_c_748_n 0.0161594f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_630_74#_c_749_n 0.00283021f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_630_74#_c_750_n 0.028187f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_630_74#_c_751_n 0.0057714f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_630_74#_c_752_n 0.00255947f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_630_74#_c_753_n 0.0142198f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_1243_48#_M1014_g 0.0299074f $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=0.58
cc_59 VNB N_A_1243_48#_c_940_n 0.0200763f $X=-0.19 $Y=-0.245 $X2=2.04 $Y2=2.585
cc_60 VNB N_A_1243_48#_c_941_n 0.0105146f $X=-0.19 $Y=-0.245 $X2=0.17 $Y2=1.47
cc_61 VNB N_A_1243_48#_c_942_n 0.0348374f $X=-0.19 $Y=-0.245 $X2=0.355 $Y2=2.41
cc_62 VNB N_A_1243_48#_c_943_n 0.00303124f $X=-0.19 $Y=-0.245 $X2=1.865
+ $Y2=2.055
cc_63 VNB N_A_1243_48#_c_944_n 0.00592303f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_1243_48#_c_945_n 0.00230825f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_1021_97#_M1018_g 0.0509144f $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=0.58
cc_66 VNB N_A_1021_97#_c_1010_n 0.0108586f $X=-0.19 $Y=-0.245 $X2=2.04 $Y2=2.19
cc_67 VNB N_A_1021_97#_c_1011_n 0.0163848f $X=-0.19 $Y=-0.245 $X2=0.17 $Y2=0.73
cc_68 VNB N_A_1021_97#_c_1012_n 0.00798764f $X=-0.19 $Y=-0.245 $X2=0.302
+ $Y2=2.41
cc_69 VNB N_A_1021_97#_c_1013_n 0.00413267f $X=-0.19 $Y=-0.245 $X2=0.915
+ $Y2=2.055
cc_70 VNB N_A_1021_97#_c_1014_n 0.00234454f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_1711_48#_c_1092_n 0.0189169f $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=1.47
cc_72 VNB N_A_1711_48#_c_1093_n 0.022038f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_1711_48#_c_1094_n 0.00621707f $X=-0.19 $Y=-0.245 $X2=2.04 $Y2=2.19
cc_74 VNB N_A_1711_48#_c_1095_n 0.0334997f $X=-0.19 $Y=-0.245 $X2=0.17 $Y2=1.47
cc_75 VNB N_A_1711_48#_c_1096_n 0.0575969f $X=-0.19 $Y=-0.245 $X2=0.302 $Y2=1.8
cc_76 VNB N_A_1711_48#_c_1097_n 0.015362f $X=-0.19 $Y=-0.245 $X2=0.355 $Y2=2.41
cc_77 VNB N_A_1711_48#_M1022_g 0.0236667f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=2.055
cc_78 VNB N_A_1711_48#_c_1099_n 0.0132804f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_1711_48#_c_1100_n 0.0125197f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_1711_48#_M1037_g 0.0228514f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.635
cc_81 VNB N_A_1711_48#_c_1102_n 0.0553787f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_1711_48#_c_1103_n 0.0133157f $X=-0.19 $Y=-0.245 $X2=2.03 $Y2=1.89
cc_83 VNB N_A_1711_48#_M1021_g 0.0240308f $X=-0.19 $Y=-0.245 $X2=2.03 $Y2=1.89
cc_84 VNB N_A_1711_48#_c_1105_n 0.00294508f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_1711_48#_c_1106_n 0.0055596f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_1711_48#_c_1107_n 0.00587191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_1711_48#_c_1108_n 6.43454e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_1711_48#_c_1109_n 0.00872918f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_1711_48#_c_1110_n 0.00241988f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_1511_74#_c_1256_n 0.00692266f $X=-0.19 $Y=-0.245 $X2=2.04 $Y2=2.19
cc_91 VNB N_A_1511_74#_c_1257_n 0.0143329f $X=-0.19 $Y=-0.245 $X2=1.865
+ $Y2=2.055
cc_92 VNB N_A_1511_74#_c_1258_n 0.00316682f $X=-0.19 $Y=-0.245 $X2=0.325
+ $Y2=0.54
cc_93 VNB N_A_1511_74#_c_1259_n 0.0102043f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_1511_74#_c_1260_n 0.00591385f $X=-0.19 $Y=-0.245 $X2=0.302
+ $Y2=1.635
cc_95 VNB N_A_1511_74#_c_1261_n 0.00598581f $X=-0.19 $Y=-0.245 $X2=0.75
+ $Y2=1.635
cc_96 VNB N_A_1511_74#_c_1262_n 0.00376276f $X=-0.19 $Y=-0.245 $X2=2.03 $Y2=1.89
cc_97 VNB N_A_1511_74#_c_1263_n 0.0356373f $X=-0.19 $Y=-0.245 $X2=2.03 $Y2=2.055
cc_98 VNB N_A_1511_74#_c_1264_n 0.0204387f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_A_2322_368#_M1019_g 0.0221608f $X=-0.19 $Y=-0.245 $X2=2.04 $Y2=2.585
cc_100 VNB N_A_2322_368#_M1039_g 0.0224961f $X=-0.19 $Y=-0.245 $X2=0.17 $Y2=1.47
cc_101 VNB N_A_2322_368#_c_1368_n 0.00801417f $X=-0.19 $Y=-0.245 $X2=1.865
+ $Y2=2.055
cc_102 VNB N_A_2322_368#_c_1369_n 0.0107941f $X=-0.19 $Y=-0.245 $X2=0.75
+ $Y2=1.635
cc_103 VNB N_A_2322_368#_c_1370_n 0.0025337f $X=-0.19 $Y=-0.245 $X2=0.83
+ $Y2=1.635
cc_104 VNB N_A_2322_368#_c_1371_n 0.0471384f $X=-0.19 $Y=-0.245 $X2=2.03
+ $Y2=1.89
cc_105 VNB N_VPWR_c_1439_n 0.561729f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_A_301_74#_c_1605_n 0.00841669f $X=-0.19 $Y=-0.245 $X2=0.83 $Y2=1.97
cc_107 VNB N_A_301_74#_c_1606_n 0.0166024f $X=-0.19 $Y=-0.245 $X2=1.865
+ $Y2=2.055
cc_108 VNB N_A_301_74#_c_1607_n 0.0124226f $X=-0.19 $Y=-0.245 $X2=0.915
+ $Y2=2.055
cc_109 VNB N_A_301_74#_c_1608_n 0.00226495f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_A_301_74#_c_1609_n 0.00793804f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_A_301_74#_c_1610_n 0.00294352f $X=-0.19 $Y=-0.245 $X2=0.302
+ $Y2=1.635
cc_112 VNB N_A_301_74#_c_1611_n 0.016819f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.635
cc_113 VNB N_Q_c_1731_n 0.00247093f $X=-0.19 $Y=-0.245 $X2=0.17 $Y2=0.73
cc_114 VNB Q 0.00240191f $X=-0.19 $Y=-0.245 $X2=0.302 $Y2=1.8
cc_115 VNB Q 0.00176823f $X=-0.19 $Y=-0.245 $X2=0.302 $Y2=2.41
cc_116 VNB N_Q_N_c_1770_n 0.0148262f $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=1.47
cc_117 VNB Q_N 0.0259261f $X=-0.19 $Y=-0.245 $X2=0.17 $Y2=1.47
cc_118 VNB N_VGND_c_1799_n 0.00641221f $X=-0.19 $Y=-0.245 $X2=0.302 $Y2=1.635
cc_119 VNB N_VGND_c_1800_n 0.0143164f $X=-0.19 $Y=-0.245 $X2=0.83 $Y2=1.635
cc_120 VNB N_VGND_c_1801_n 0.0113387f $X=-0.19 $Y=-0.245 $X2=2.03 $Y2=2.055
cc_121 VNB N_VGND_c_1802_n 0.00619653f $X=-0.19 $Y=-0.245 $X2=2.03 $Y2=1.89
cc_122 VNB N_VGND_c_1803_n 0.0186543f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB N_VGND_c_1804_n 0.0237579f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_VGND_c_1805_n 0.0105835f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_1806_n 0.00274125f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_1807_n 0.0121789f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_VGND_c_1808_n 0.0240848f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_1809_n 0.0472928f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_1810_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_1811_n 0.0209223f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_1812_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_VGND_c_1813_n 0.0558968f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_VGND_c_1814_n 0.0528991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_VGND_c_1815_n 0.0201672f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_VGND_c_1816_n 0.019013f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_VGND_c_1817_n 0.0216352f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_VGND_c_1818_n 0.0172267f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB N_VGND_c_1819_n 0.0261411f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VNB N_VGND_c_1820_n 0.00613227f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_VGND_c_1821_n 0.0240346f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_141 VNB N_VGND_c_1822_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_142 VNB N_VGND_c_1823_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_143 VNB N_VGND_c_1824_n 0.00630956f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_144 VNB N_VGND_c_1825_n 0.742528f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_145 VPB N_A_36_74#_c_273_n 0.0570354f $X=-0.19 $Y=1.66 $X2=2.04 $Y2=2.19
cc_146 VPB N_A_36_74#_c_269_n 0.019329f $X=-0.19 $Y=1.66 $X2=0.965 $Y2=1.635
cc_147 VPB N_A_36_74#_c_275_n 0.0536724f $X=-0.19 $Y=1.66 $X2=0.355 $Y2=2.41
cc_148 VPB N_A_36_74#_c_276_n 0.0032166f $X=-0.19 $Y=1.66 $X2=0.83 $Y2=1.97
cc_149 VPB N_A_36_74#_c_277_n 0.0230799f $X=-0.19 $Y=1.66 $X2=1.865 $Y2=2.055
cc_150 VPB N_A_36_74#_c_278_n 5.35807e-19 $X=-0.19 $Y=1.66 $X2=0.915 $Y2=2.055
cc_151 VPB N_A_36_74#_c_272_n 0.00704567f $X=-0.19 $Y=1.66 $X2=0.83 $Y2=1.635
cc_152 VPB N_A_36_74#_c_280_n 0.00613935f $X=-0.19 $Y=1.66 $X2=2.03 $Y2=1.89
cc_153 VPB N_SCE_c_352_n 0.022762f $X=-0.19 $Y=1.66 $X2=0.21 $Y2=2.265
cc_154 VPB N_SCE_c_360_n 0.0184239f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_155 VPB N_SCE_c_361_n 0.0109496f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_156 VPB N_SCE_c_362_n 0.0176252f $X=-0.19 $Y=1.66 $X2=1.04 $Y2=0.58
cc_157 VPB N_SCE_c_363_n 0.0195802f $X=-0.19 $Y=1.66 $X2=2.04 $Y2=2.19
cc_158 VPB N_SCE_c_364_n 0.0142664f $X=-0.19 $Y=1.66 $X2=2.04 $Y2=2.585
cc_159 VPB N_SCE_c_365_n 0.00512496f $X=-0.19 $Y=1.66 $X2=0.355 $Y2=2.41
cc_160 VPB N_D_c_430_n 0.0179397f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_161 VPB N_D_c_431_n 0.0219397f $X=-0.19 $Y=1.66 $X2=1.04 $Y2=1.47
cc_162 VPB N_D_c_428_n 0.0127342f $X=-0.19 $Y=1.66 $X2=2.04 $Y2=2.585
cc_163 VPB N_D_c_429_n 0.00476594f $X=-0.19 $Y=1.66 $X2=0.965 $Y2=1.635
cc_164 VPB N_SCD_c_469_n 0.0555514f $X=-0.19 $Y=1.66 $X2=0.18 $Y2=0.37
cc_165 VPB N_SCD_M1024_g 0.00880265f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_166 VPB N_SCD_c_471_n 0.00678985f $X=-0.19 $Y=1.66 $X2=2.04 $Y2=2.585
cc_167 VPB N_CLK_c_504_n 0.021554f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_168 VPB CLK 0.0042588f $X=-0.19 $Y=1.66 $X2=1.04 $Y2=0.58
cc_169 VPB N_CLK_c_503_n 0.015843f $X=-0.19 $Y=1.66 $X2=2.04 $Y2=2.19
cc_170 VPB N_A_828_74#_c_559_n 0.0192302f $X=-0.19 $Y=1.66 $X2=1.04 $Y2=1.47
cc_171 VPB N_A_828_74#_c_560_n 0.0136492f $X=-0.19 $Y=1.66 $X2=0.302 $Y2=2.41
cc_172 VPB N_A_828_74#_c_561_n 0.0232052f $X=-0.19 $Y=1.66 $X2=0.355 $Y2=2.41
cc_173 VPB N_A_828_74#_c_540_n 0.017918f $X=-0.19 $Y=1.66 $X2=0.915 $Y2=2.055
cc_174 VPB N_A_828_74#_c_563_n 0.012659f $X=-0.19 $Y=1.66 $X2=0.17 $Y2=0.54
cc_175 VPB N_A_828_74#_c_544_n 0.0138005f $X=-0.19 $Y=1.66 $X2=0.75 $Y2=1.635
cc_176 VPB N_A_828_74#_c_565_n 0.0540189f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_177 VPB N_A_630_74#_c_738_n 0.0105095f $X=-0.19 $Y=1.66 $X2=2.04 $Y2=2.19
cc_178 VPB N_A_630_74#_c_755_n 0.022056f $X=-0.19 $Y=1.66 $X2=2.04 $Y2=2.585
cc_179 VPB N_A_630_74#_c_739_n 0.0134097f $X=-0.19 $Y=1.66 $X2=0.17 $Y2=1.47
cc_180 VPB N_A_630_74#_c_741_n 0.0258197f $X=-0.19 $Y=1.66 $X2=0.83 $Y2=1.97
cc_181 VPB N_A_630_74#_c_758_n 0.0226372f $X=-0.19 $Y=1.66 $X2=0.17 $Y2=0.54
cc_182 VPB N_A_630_74#_c_759_n 0.0424539f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_183 VPB N_A_630_74#_c_760_n 0.0186738f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_184 VPB N_A_630_74#_c_744_n 0.00167153f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_185 VPB N_A_630_74#_c_745_n 0.00464422f $X=-0.19 $Y=1.66 $X2=2.03 $Y2=1.89
cc_186 VPB N_A_630_74#_c_763_n 0.00558792f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_187 VPB N_A_630_74#_c_764_n 0.00369325f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_188 VPB N_A_630_74#_c_750_n 0.0158138f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_189 VPB N_A_630_74#_c_766_n 0.00256525f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_190 VPB N_A_630_74#_c_767_n 0.00279391f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_191 VPB N_A_630_74#_c_768_n 0.00424858f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_192 VPB N_A_630_74#_c_752_n 7.45923e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_193 VPB N_A_630_74#_c_753_n 0.0450813f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_194 VPB N_A_1243_48#_c_940_n 0.0370272f $X=-0.19 $Y=1.66 $X2=2.04 $Y2=2.585
cc_195 VPB N_A_1243_48#_c_947_n 0.0225479f $X=-0.19 $Y=1.66 $X2=2.04 $Y2=2.585
cc_196 VPB N_A_1243_48#_c_948_n 0.00333166f $X=-0.19 $Y=1.66 $X2=0.325 $Y2=0.54
cc_197 VPB N_A_1243_48#_c_944_n 0.00823746f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_198 VPB N_A_1021_97#_c_1010_n 0.0573711f $X=-0.19 $Y=1.66 $X2=2.04 $Y2=2.19
cc_199 VPB N_A_1021_97#_c_1012_n 0.0125318f $X=-0.19 $Y=1.66 $X2=0.302 $Y2=2.41
cc_200 VPB N_A_1021_97#_c_1017_n 0.00888065f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_201 VPB N_A_1021_97#_c_1018_n 0.00921162f $X=-0.19 $Y=1.66 $X2=0.325 $Y2=0.54
cc_202 VPB N_A_1021_97#_c_1014_n 0.0039159f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_203 VPB N_A_1711_48#_c_1111_n 0.0537782f $X=-0.19 $Y=1.66 $X2=2.04 $Y2=2.585
cc_204 VPB N_A_1711_48#_c_1095_n 0.0231212f $X=-0.19 $Y=1.66 $X2=0.17 $Y2=1.47
cc_205 VPB N_A_1711_48#_c_1097_n 0.024502f $X=-0.19 $Y=1.66 $X2=0.355 $Y2=2.41
cc_206 VPB N_A_1711_48#_c_1100_n 8.53067e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_207 VPB N_A_1711_48#_c_1115_n 0.0236313f $X=-0.19 $Y=1.66 $X2=0.17 $Y2=1.635
cc_208 VPB N_A_1711_48#_c_1103_n 9.71585e-19 $X=-0.19 $Y=1.66 $X2=2.03 $Y2=1.89
cc_209 VPB N_A_1711_48#_c_1117_n 0.0252442f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_210 VPB N_A_1711_48#_c_1118_n 0.0106358f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_211 VPB N_A_1711_48#_c_1119_n 0.00854044f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_212 VPB N_A_1711_48#_c_1108_n 0.00629202f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_213 VPB N_A_1711_48#_c_1121_n 0.0104973f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_214 VPB N_A_1511_74#_c_1256_n 0.00874501f $X=-0.19 $Y=1.66 $X2=2.04 $Y2=2.19
cc_215 VPB N_A_1511_74#_c_1266_n 0.0256894f $X=-0.19 $Y=1.66 $X2=2.04 $Y2=2.585
cc_216 VPB N_A_1511_74#_c_1267_n 0.00347435f $X=-0.19 $Y=1.66 $X2=0.302 $Y2=1.8
cc_217 VPB N_A_1511_74#_c_1268_n 0.00571717f $X=-0.19 $Y=1.66 $X2=0.355 $Y2=2.41
cc_218 VPB N_A_1511_74#_c_1269_n 0.015837f $X=-0.19 $Y=1.66 $X2=0.17 $Y2=0.54
cc_219 VPB N_A_1511_74#_c_1270_n 0.00199812f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_220 VPB N_A_1511_74#_c_1258_n 6.58716e-19 $X=-0.19 $Y=1.66 $X2=0.325 $Y2=0.54
cc_221 VPB N_A_1511_74#_c_1272_n 0.00387282f $X=-0.19 $Y=1.66 $X2=0.75 $Y2=1.635
cc_222 VPB N_A_2322_368#_c_1372_n 0.0163328f $X=-0.19 $Y=1.66 $X2=1.04 $Y2=1.47
cc_223 VPB N_A_2322_368#_c_1373_n 0.0171853f $X=-0.19 $Y=1.66 $X2=0.302 $Y2=2.41
cc_224 VPB N_A_2322_368#_c_1374_n 0.015347f $X=-0.19 $Y=1.66 $X2=0.325 $Y2=0.54
cc_225 VPB N_A_2322_368#_c_1371_n 0.0140201f $X=-0.19 $Y=1.66 $X2=2.03 $Y2=1.89
cc_226 VPB N_VPWR_c_1440_n 0.00817207f $X=-0.19 $Y=1.66 $X2=0.17 $Y2=1.635
cc_227 VPB N_VPWR_c_1441_n 0.0122054f $X=-0.19 $Y=1.66 $X2=0.75 $Y2=1.635
cc_228 VPB N_VPWR_c_1442_n 0.0197665f $X=-0.19 $Y=1.66 $X2=2.03 $Y2=1.89
cc_229 VPB N_VPWR_c_1443_n 0.0091289f $X=-0.19 $Y=1.66 $X2=2.03 $Y2=2.055
cc_230 VPB N_VPWR_c_1444_n 0.0204201f $X=-0.19 $Y=1.66 $X2=2.03 $Y2=1.89
cc_231 VPB N_VPWR_c_1445_n 0.00147296f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_232 VPB N_VPWR_c_1446_n 0.0157674f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_233 VPB N_VPWR_c_1447_n 0.00751242f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_234 VPB N_VPWR_c_1448_n 0.0152249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_235 VPB N_VPWR_c_1449_n 0.0116916f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_236 VPB N_VPWR_c_1450_n 0.0349184f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_237 VPB N_VPWR_c_1451_n 0.0221649f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_238 VPB N_VPWR_c_1452_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_239 VPB N_VPWR_c_1453_n 0.0490287f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_240 VPB N_VPWR_c_1454_n 0.00805426f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_241 VPB N_VPWR_c_1455_n 0.0152746f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_242 VPB N_VPWR_c_1456_n 0.0595113f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_243 VPB N_VPWR_c_1457_n 0.0198114f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_244 VPB N_VPWR_c_1458_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_245 VPB N_VPWR_c_1459_n 0.0312042f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_246 VPB N_VPWR_c_1460_n 0.0550499f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_247 VPB N_VPWR_c_1461_n 0.0185253f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_248 VPB N_VPWR_c_1462_n 0.0213015f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_249 VPB N_VPWR_c_1463_n 0.0182909f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_250 VPB N_VPWR_c_1464_n 0.00614248f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_251 VPB N_VPWR_c_1465_n 0.0107576f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_252 VPB N_VPWR_c_1466_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_253 VPB N_VPWR_c_1467_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_254 VPB N_VPWR_c_1439_n 0.186563f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_255 VPB N_A_301_74#_c_1608_n 0.00378781f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_256 VPB N_A_301_74#_c_1613_n 0.00828904f $X=-0.19 $Y=1.66 $X2=0.325 $Y2=0.54
cc_257 VPB N_A_301_74#_c_1614_n 6.88992e-19 $X=-0.19 $Y=1.66 $X2=0.17 $Y2=1.635
cc_258 VPB N_A_301_74#_c_1615_n 0.00755526f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_259 VPB N_A_301_74#_c_1616_n 0.00322246f $X=-0.19 $Y=1.66 $X2=2.03 $Y2=1.89
cc_260 VPB N_A_301_74#_c_1617_n 0.00854763f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_261 VPB N_Q_c_1734_n 0.00216998f $X=-0.19 $Y=1.66 $X2=1.04 $Y2=0.58
cc_262 VPB N_Q_c_1731_n 8.5811e-19 $X=-0.19 $Y=1.66 $X2=0.17 $Y2=0.73
cc_263 VPB N_Q_c_1736_n 0.00169544f $X=-0.19 $Y=1.66 $X2=0.17 $Y2=1.47
cc_264 VPB N_Q_N_c_1772_n 0.00243101f $X=-0.19 $Y=1.66 $X2=2.04 $Y2=2.585
cc_265 VPB Q_N 0.00860152f $X=-0.19 $Y=1.66 $X2=0.17 $Y2=1.47
cc_266 VPB Q_N 0.0172577f $X=-0.19 $Y=1.66 $X2=0.302 $Y2=2.41
cc_267 N_A_36_74#_M1012_g N_SCE_c_352_n 0.00365204f $X=1.04 $Y=0.58 $X2=0 $Y2=0
cc_268 N_A_36_74#_c_269_n N_SCE_c_352_n 0.0181416f $X=0.965 $Y=1.635 $X2=0 $Y2=0
cc_269 N_A_36_74#_c_270_n N_SCE_c_352_n 0.0150312f $X=0.17 $Y=1.47 $X2=0 $Y2=0
cc_270 N_A_36_74#_c_275_n N_SCE_c_352_n 0.0104604f $X=0.355 $Y=2.41 $X2=0 $Y2=0
cc_271 N_A_36_74#_c_276_n N_SCE_c_352_n 6.96051e-19 $X=0.83 $Y=1.97 $X2=0 $Y2=0
cc_272 N_A_36_74#_c_272_n N_SCE_c_352_n 0.0181742f $X=0.83 $Y=1.635 $X2=0 $Y2=0
cc_273 N_A_36_74#_c_269_n N_SCE_c_360_n 0.0301061f $X=0.965 $Y=1.635 $X2=0 $Y2=0
cc_274 N_A_36_74#_c_275_n N_SCE_c_360_n 0.0138037f $X=0.355 $Y=2.41 $X2=0 $Y2=0
cc_275 N_A_36_74#_c_272_n N_SCE_c_360_n 0.00411717f $X=0.83 $Y=1.635 $X2=0 $Y2=0
cc_276 N_A_36_74#_c_275_n N_SCE_c_361_n 0.00835712f $X=0.355 $Y=2.41 $X2=0 $Y2=0
cc_277 N_A_36_74#_M1012_g N_SCE_c_353_n 0.0153057f $X=1.04 $Y=0.58 $X2=0 $Y2=0
cc_278 N_A_36_74#_c_270_n N_SCE_c_353_n 0.00547775f $X=0.17 $Y=1.47 $X2=0 $Y2=0
cc_279 N_A_36_74#_c_271_n N_SCE_c_353_n 0.00485153f $X=0.325 $Y=0.54 $X2=0 $Y2=0
cc_280 N_A_36_74#_c_275_n N_SCE_c_362_n 0.0191458f $X=0.355 $Y=2.41 $X2=0 $Y2=0
cc_281 N_A_36_74#_c_277_n N_SCE_c_363_n 0.0141402f $X=1.865 $Y=2.055 $X2=0 $Y2=0
cc_282 N_A_36_74#_c_278_n N_SCE_c_363_n 0.00645861f $X=0.915 $Y=2.055 $X2=0
+ $Y2=0
cc_283 N_A_36_74#_c_273_n N_SCE_c_355_n 0.00695671f $X=2.04 $Y=2.19 $X2=0 $Y2=0
cc_284 N_A_36_74#_c_280_n N_SCE_c_355_n 0.00166786f $X=2.03 $Y=1.89 $X2=0 $Y2=0
cc_285 N_A_36_74#_M1012_g N_SCE_c_356_n 0.0214013f $X=1.04 $Y=0.58 $X2=0 $Y2=0
cc_286 N_A_36_74#_c_269_n N_SCE_c_356_n 0.00889754f $X=0.965 $Y=1.635 $X2=0
+ $Y2=0
cc_287 N_A_36_74#_c_270_n N_SCE_c_356_n 0.0127879f $X=0.17 $Y=1.47 $X2=0 $Y2=0
cc_288 N_A_36_74#_c_271_n N_SCE_c_356_n 0.00812187f $X=0.325 $Y=0.54 $X2=0 $Y2=0
cc_289 N_A_36_74#_c_272_n N_SCE_c_356_n 0.00757297f $X=0.83 $Y=1.635 $X2=0 $Y2=0
cc_290 N_A_36_74#_c_273_n N_SCE_c_357_n 2.43991e-19 $X=2.04 $Y=2.19 $X2=0 $Y2=0
cc_291 N_A_36_74#_c_280_n N_SCE_c_357_n 0.00681972f $X=2.03 $Y=1.89 $X2=0 $Y2=0
cc_292 N_A_36_74#_M1012_g N_SCE_c_358_n 0.0230183f $X=1.04 $Y=0.58 $X2=0 $Y2=0
cc_293 N_A_36_74#_c_269_n N_SCE_c_358_n 0.00597298f $X=0.965 $Y=1.635 $X2=0
+ $Y2=0
cc_294 N_A_36_74#_c_270_n N_SCE_c_358_n 0.0249855f $X=0.17 $Y=1.47 $X2=0 $Y2=0
cc_295 N_A_36_74#_c_271_n N_SCE_c_358_n 0.00335915f $X=0.325 $Y=0.54 $X2=0 $Y2=0
cc_296 N_A_36_74#_c_272_n N_SCE_c_358_n 0.0292685f $X=0.83 $Y=1.635 $X2=0 $Y2=0
cc_297 N_A_36_74#_M1012_g N_D_M1013_g 0.06651f $X=1.04 $Y=0.58 $X2=0 $Y2=0
cc_298 N_A_36_74#_c_273_n N_D_c_430_n 0.0196743f $X=2.04 $Y=2.19 $X2=0 $Y2=0
cc_299 N_A_36_74#_c_276_n N_D_c_430_n 0.0040545f $X=0.83 $Y=1.97 $X2=0 $Y2=0
cc_300 N_A_36_74#_c_277_n N_D_c_430_n 0.00819153f $X=1.865 $Y=2.055 $X2=0 $Y2=0
cc_301 N_A_36_74#_c_280_n N_D_c_430_n 0.00125029f $X=2.03 $Y=1.89 $X2=0 $Y2=0
cc_302 N_A_36_74#_c_273_n N_D_c_431_n 0.0163506f $X=2.04 $Y=2.19 $X2=0 $Y2=0
cc_303 N_A_36_74#_c_277_n N_D_c_431_n 0.00921209f $X=1.865 $Y=2.055 $X2=0 $Y2=0
cc_304 N_A_36_74#_c_273_n N_D_c_428_n 0.00472913f $X=2.04 $Y=2.19 $X2=0 $Y2=0
cc_305 N_A_36_74#_c_269_n N_D_c_428_n 0.0214888f $X=0.965 $Y=1.635 $X2=0 $Y2=0
cc_306 N_A_36_74#_c_277_n N_D_c_428_n 0.00371768f $X=1.865 $Y=2.055 $X2=0 $Y2=0
cc_307 N_A_36_74#_c_273_n N_D_c_429_n 2.57473e-19 $X=2.04 $Y=2.19 $X2=0 $Y2=0
cc_308 N_A_36_74#_c_269_n N_D_c_429_n 0.00926354f $X=0.965 $Y=1.635 $X2=0 $Y2=0
cc_309 N_A_36_74#_c_277_n N_D_c_429_n 0.0430314f $X=1.865 $Y=2.055 $X2=0 $Y2=0
cc_310 N_A_36_74#_c_272_n N_D_c_429_n 0.0273977f $X=0.83 $Y=1.635 $X2=0 $Y2=0
cc_311 N_A_36_74#_c_280_n N_D_c_429_n 0.00491403f $X=2.03 $Y=1.89 $X2=0 $Y2=0
cc_312 N_A_36_74#_c_273_n N_SCD_c_469_n 0.0544451f $X=2.04 $Y=2.19 $X2=-0.19
+ $Y2=-0.245
cc_313 N_A_36_74#_c_280_n N_SCD_c_469_n 0.00142356f $X=2.03 $Y=1.89 $X2=-0.19
+ $Y2=-0.245
cc_314 N_A_36_74#_c_273_n N_SCD_M1024_g 0.0022386f $X=2.04 $Y=2.19 $X2=0 $Y2=0
cc_315 N_A_36_74#_c_280_n N_SCD_M1024_g 3.06975e-19 $X=2.03 $Y=1.89 $X2=0 $Y2=0
cc_316 N_A_36_74#_c_273_n N_SCD_c_471_n 0.00136139f $X=2.04 $Y=2.19 $X2=0 $Y2=0
cc_317 N_A_36_74#_c_280_n N_SCD_c_471_n 0.0237414f $X=2.03 $Y=1.89 $X2=0 $Y2=0
cc_318 N_A_36_74#_c_275_n N_VPWR_c_1440_n 0.0422703f $X=0.355 $Y=2.41 $X2=0
+ $Y2=0
cc_319 N_A_36_74#_c_277_n N_VPWR_c_1440_n 0.00826449f $X=1.865 $Y=2.055 $X2=0
+ $Y2=0
cc_320 N_A_36_74#_c_278_n N_VPWR_c_1440_n 0.0118028f $X=0.915 $Y=2.055 $X2=0
+ $Y2=0
cc_321 N_A_36_74#_c_272_n N_VPWR_c_1440_n 5.44119e-19 $X=0.83 $Y=1.635 $X2=0
+ $Y2=0
cc_322 N_A_36_74#_c_275_n N_VPWR_c_1451_n 0.0158129f $X=0.355 $Y=2.41 $X2=0
+ $Y2=0
cc_323 N_A_36_74#_c_273_n N_VPWR_c_1453_n 0.00523995f $X=2.04 $Y=2.19 $X2=0
+ $Y2=0
cc_324 N_A_36_74#_c_273_n N_VPWR_c_1439_n 0.00528353f $X=2.04 $Y=2.19 $X2=0
+ $Y2=0
cc_325 N_A_36_74#_c_275_n N_VPWR_c_1439_n 0.0154507f $X=0.355 $Y=2.41 $X2=0
+ $Y2=0
cc_326 N_A_36_74#_M1012_g N_A_301_74#_c_1618_n 6.99132e-19 $X=1.04 $Y=0.58 $X2=0
+ $Y2=0
cc_327 N_A_36_74#_c_273_n N_A_301_74#_c_1619_n 0.00970262f $X=2.04 $Y=2.19 $X2=0
+ $Y2=0
cc_328 N_A_36_74#_c_280_n N_A_301_74#_c_1619_n 0.0110596f $X=2.03 $Y=1.89 $X2=0
+ $Y2=0
cc_329 N_A_36_74#_c_273_n N_A_301_74#_c_1616_n 0.00937278f $X=2.04 $Y=2.19 $X2=0
+ $Y2=0
cc_330 N_A_36_74#_c_277_n N_A_301_74#_c_1616_n 0.0168838f $X=1.865 $Y=2.055
+ $X2=0 $Y2=0
cc_331 N_A_36_74#_c_280_n N_A_301_74#_c_1616_n 0.00728111f $X=2.03 $Y=1.89 $X2=0
+ $Y2=0
cc_332 N_A_36_74#_M1012_g N_VGND_c_1799_n 0.0107959f $X=1.04 $Y=0.58 $X2=0 $Y2=0
cc_333 N_A_36_74#_c_271_n N_VGND_c_1799_n 0.0154676f $X=0.325 $Y=0.54 $X2=0
+ $Y2=0
cc_334 N_A_36_74#_M1012_g N_VGND_c_1809_n 0.00383152f $X=1.04 $Y=0.58 $X2=0
+ $Y2=0
cc_335 N_A_36_74#_c_271_n N_VGND_c_1819_n 0.0171909f $X=0.325 $Y=0.54 $X2=0
+ $Y2=0
cc_336 N_A_36_74#_M1012_g N_VGND_c_1825_n 0.0075725f $X=1.04 $Y=0.58 $X2=0 $Y2=0
cc_337 N_A_36_74#_c_271_n N_VGND_c_1825_n 0.0145444f $X=0.325 $Y=0.54 $X2=0
+ $Y2=0
cc_338 N_SCE_c_354_n N_D_M1013_g 0.0125462f $X=2.175 $Y=0.9 $X2=0 $Y2=0
cc_339 N_SCE_c_355_n N_D_M1013_g 0.0181291f $X=2.1 $Y=1.065 $X2=0 $Y2=0
cc_340 N_SCE_c_357_n N_D_M1013_g 0.00293704f $X=1.91 $Y=1.065 $X2=0 $Y2=0
cc_341 N_SCE_c_358_n N_D_M1013_g 0.020051f $X=1.565 $Y=1.02 $X2=0 $Y2=0
cc_342 N_SCE_c_363_n N_D_c_430_n 0.00884233f $X=1.04 $Y=2.115 $X2=0 $Y2=0
cc_343 N_SCE_c_364_n N_D_c_431_n 0.0378564f $X=1.115 $Y=2.19 $X2=0 $Y2=0
cc_344 N_SCE_c_358_n N_D_c_428_n 0.00437854f $X=1.565 $Y=1.02 $X2=0 $Y2=0
cc_345 N_SCE_c_363_n N_D_c_429_n 5.83509e-19 $X=1.04 $Y=2.115 $X2=0 $Y2=0
cc_346 N_SCE_c_358_n N_D_c_429_n 0.0350954f $X=1.565 $Y=1.02 $X2=0 $Y2=0
cc_347 N_SCE_c_354_n N_SCD_M1024_g 0.0494463f $X=2.175 $Y=0.9 $X2=0 $Y2=0
cc_348 N_SCE_c_362_n N_VPWR_c_1440_n 0.0135431f $X=0.665 $Y=2.19 $X2=0 $Y2=0
cc_349 N_SCE_c_363_n N_VPWR_c_1440_n 0.00254598f $X=1.04 $Y=2.115 $X2=0 $Y2=0
cc_350 N_SCE_c_364_n N_VPWR_c_1440_n 0.0149392f $X=1.115 $Y=2.19 $X2=0 $Y2=0
cc_351 N_SCE_c_362_n N_VPWR_c_1451_n 0.0048289f $X=0.665 $Y=2.19 $X2=0 $Y2=0
cc_352 N_SCE_c_364_n N_VPWR_c_1453_n 0.0048289f $X=1.115 $Y=2.19 $X2=0 $Y2=0
cc_353 N_SCE_c_362_n N_VPWR_c_1439_n 0.0047904f $X=0.665 $Y=2.19 $X2=0 $Y2=0
cc_354 N_SCE_c_364_n N_VPWR_c_1439_n 0.0047904f $X=1.115 $Y=2.19 $X2=0 $Y2=0
cc_355 N_SCE_c_354_n N_A_301_74#_c_1618_n 0.0180824f $X=2.175 $Y=0.9 $X2=0 $Y2=0
cc_356 N_SCE_c_355_n N_A_301_74#_c_1618_n 0.00183369f $X=2.1 $Y=1.065 $X2=0
+ $Y2=0
cc_357 N_SCE_c_357_n N_A_301_74#_c_1618_n 0.0391871f $X=1.91 $Y=1.065 $X2=0
+ $Y2=0
cc_358 N_SCE_c_358_n N_A_301_74#_c_1618_n 0.00322043f $X=1.565 $Y=1.02 $X2=0
+ $Y2=0
cc_359 N_SCE_c_354_n N_A_301_74#_c_1605_n 0.00915416f $X=2.175 $Y=0.9 $X2=0
+ $Y2=0
cc_360 N_SCE_c_355_n N_A_301_74#_c_1605_n 0.00685179f $X=2.1 $Y=1.065 $X2=0
+ $Y2=0
cc_361 N_SCE_c_357_n N_A_301_74#_c_1605_n 0.0320316f $X=1.91 $Y=1.065 $X2=0
+ $Y2=0
cc_362 N_SCE_c_353_n N_VGND_c_1799_n 0.00515645f $X=0.54 $Y=0.9 $X2=0 $Y2=0
cc_363 N_SCE_c_356_n N_VGND_c_1799_n 0.00215627f $X=0.59 $Y=1.065 $X2=0 $Y2=0
cc_364 N_SCE_c_358_n N_VGND_c_1799_n 0.0247894f $X=1.565 $Y=1.02 $X2=0 $Y2=0
cc_365 N_SCE_c_354_n N_VGND_c_1809_n 0.0029698f $X=2.175 $Y=0.9 $X2=0 $Y2=0
cc_366 N_SCE_c_353_n N_VGND_c_1819_n 0.00433162f $X=0.54 $Y=0.9 $X2=0 $Y2=0
cc_367 N_SCE_c_353_n N_VGND_c_1825_n 0.00820923f $X=0.54 $Y=0.9 $X2=0 $Y2=0
cc_368 N_SCE_c_354_n N_VGND_c_1825_n 0.00366067f $X=2.175 $Y=0.9 $X2=0 $Y2=0
cc_369 N_D_c_431_n N_VPWR_c_1440_n 0.00234372f $X=1.535 $Y=2.19 $X2=0 $Y2=0
cc_370 N_D_c_431_n N_VPWR_c_1453_n 0.00537957f $X=1.535 $Y=2.19 $X2=0 $Y2=0
cc_371 N_D_c_431_n N_VPWR_c_1439_n 0.00528353f $X=1.535 $Y=2.19 $X2=0 $Y2=0
cc_372 N_D_M1013_g N_A_301_74#_c_1618_n 0.00965085f $X=1.43 $Y=0.58 $X2=0 $Y2=0
cc_373 N_D_c_428_n N_A_301_74#_c_1607_n 3.1107e-19 $X=1.49 $Y=1.635 $X2=0 $Y2=0
cc_374 N_D_c_429_n N_A_301_74#_c_1607_n 0.00167835f $X=1.49 $Y=1.635 $X2=0 $Y2=0
cc_375 N_D_c_431_n N_A_301_74#_c_1616_n 0.0022363f $X=1.535 $Y=2.19 $X2=0 $Y2=0
cc_376 N_D_M1013_g N_VGND_c_1799_n 0.00191703f $X=1.43 $Y=0.58 $X2=0 $Y2=0
cc_377 N_D_M1013_g N_VGND_c_1809_n 0.00434051f $X=1.43 $Y=0.58 $X2=0 $Y2=0
cc_378 N_D_M1013_g N_VGND_c_1825_n 0.00820483f $X=1.43 $Y=0.58 $X2=0 $Y2=0
cc_379 N_SCD_M1024_g N_CLK_M1000_g 0.0258612f $X=2.565 $Y=0.58 $X2=0 $Y2=0
cc_380 N_SCD_c_469_n N_CLK_c_504_n 0.0219077f $X=2.525 $Y=2.19 $X2=0 $Y2=0
cc_381 N_SCD_M1024_g N_CLK_c_503_n 0.00425489f $X=2.565 $Y=0.58 $X2=0 $Y2=0
cc_382 N_SCD_M1024_g N_A_630_74#_c_749_n 2.6175e-19 $X=2.565 $Y=0.58 $X2=0 $Y2=0
cc_383 N_SCD_c_469_n N_VPWR_c_1441_n 0.0101015f $X=2.525 $Y=2.19 $X2=0 $Y2=0
cc_384 N_SCD_c_469_n N_VPWR_c_1453_n 0.00537957f $X=2.525 $Y=2.19 $X2=0 $Y2=0
cc_385 N_SCD_c_469_n N_VPWR_c_1439_n 0.00528353f $X=2.525 $Y=2.19 $X2=0 $Y2=0
cc_386 N_SCD_M1024_g N_A_301_74#_c_1618_n 0.00233346f $X=2.565 $Y=0.58 $X2=0
+ $Y2=0
cc_387 N_SCD_c_469_n N_A_301_74#_c_1619_n 0.0140024f $X=2.525 $Y=2.19 $X2=0
+ $Y2=0
cc_388 N_SCD_c_471_n N_A_301_74#_c_1619_n 0.0186802f $X=2.57 $Y=1.94 $X2=0 $Y2=0
cc_389 N_SCD_M1024_g N_A_301_74#_c_1605_n 0.0105762f $X=2.565 $Y=0.58 $X2=0
+ $Y2=0
cc_390 N_SCD_c_469_n N_A_301_74#_c_1606_n 0.00109452f $X=2.525 $Y=2.19 $X2=0
+ $Y2=0
cc_391 N_SCD_M1024_g N_A_301_74#_c_1606_n 0.0172141f $X=2.565 $Y=0.58 $X2=0
+ $Y2=0
cc_392 N_SCD_c_471_n N_A_301_74#_c_1606_n 0.0185388f $X=2.57 $Y=1.94 $X2=0 $Y2=0
cc_393 N_SCD_c_471_n N_A_301_74#_c_1607_n 5.67649e-19 $X=2.57 $Y=1.94 $X2=0
+ $Y2=0
cc_394 N_SCD_c_469_n N_A_301_74#_c_1608_n 0.00547308f $X=2.525 $Y=2.19 $X2=0
+ $Y2=0
cc_395 N_SCD_M1024_g N_A_301_74#_c_1608_n 0.00503488f $X=2.565 $Y=0.58 $X2=0
+ $Y2=0
cc_396 N_SCD_c_471_n N_A_301_74#_c_1608_n 0.0294561f $X=2.57 $Y=1.94 $X2=0 $Y2=0
cc_397 N_SCD_c_469_n N_A_301_74#_c_1616_n 0.00207884f $X=2.525 $Y=2.19 $X2=0
+ $Y2=0
cc_398 N_SCD_M1024_g N_VGND_c_1800_n 0.00901403f $X=2.565 $Y=0.58 $X2=0 $Y2=0
cc_399 N_SCD_M1024_g N_VGND_c_1809_n 0.00461464f $X=2.565 $Y=0.58 $X2=0 $Y2=0
cc_400 N_SCD_M1024_g N_VGND_c_1825_n 0.00908835f $X=2.565 $Y=0.58 $X2=0 $Y2=0
cc_401 N_CLK_M1000_g N_A_630_74#_c_747_n 0.00873769f $X=3.075 $Y=0.74 $X2=0
+ $Y2=0
cc_402 N_CLK_c_504_n N_A_630_74#_c_763_n 0.00298207f $X=3.235 $Y=1.765 $X2=0
+ $Y2=0
cc_403 CLK N_A_630_74#_c_763_n 0.0295753f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_404 N_CLK_c_503_n N_A_630_74#_c_763_n 0.0014347f $X=3.235 $Y=1.557 $X2=0
+ $Y2=0
cc_405 CLK N_A_630_74#_c_748_n 0.01799f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_406 N_CLK_c_503_n N_A_630_74#_c_748_n 0.00313668f $X=3.235 $Y=1.557 $X2=0
+ $Y2=0
cc_407 N_CLK_M1000_g N_A_630_74#_c_749_n 0.00517378f $X=3.075 $Y=0.74 $X2=0
+ $Y2=0
cc_408 CLK N_A_630_74#_c_749_n 0.0163194f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_409 N_CLK_c_503_n N_A_630_74#_c_749_n 0.0101557f $X=3.235 $Y=1.557 $X2=0
+ $Y2=0
cc_410 CLK N_A_630_74#_c_781_n 0.0339485f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_411 N_CLK_c_503_n N_A_630_74#_c_781_n 3.18999e-19 $X=3.235 $Y=1.557 $X2=0
+ $Y2=0
cc_412 N_CLK_c_504_n N_A_630_74#_c_764_n 0.00381308f $X=3.235 $Y=1.765 $X2=0
+ $Y2=0
cc_413 CLK N_A_630_74#_c_750_n 0.00311129f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_414 N_CLK_c_503_n N_A_630_74#_c_750_n 0.0218835f $X=3.235 $Y=1.557 $X2=0
+ $Y2=0
cc_415 N_CLK_c_504_n N_VPWR_c_1441_n 0.012405f $X=3.235 $Y=1.765 $X2=0 $Y2=0
cc_416 N_CLK_c_504_n N_VPWR_c_1459_n 0.00461464f $X=3.235 $Y=1.765 $X2=0 $Y2=0
cc_417 N_CLK_c_504_n N_VPWR_c_1439_n 0.00461447f $X=3.235 $Y=1.765 $X2=0 $Y2=0
cc_418 CLK N_A_301_74#_c_1606_n 0.0138901f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_419 N_CLK_c_503_n N_A_301_74#_c_1606_n 0.0132518f $X=3.235 $Y=1.557 $X2=0
+ $Y2=0
cc_420 N_CLK_c_504_n N_A_301_74#_c_1608_n 0.0114065f $X=3.235 $Y=1.765 $X2=0
+ $Y2=0
cc_421 CLK N_A_301_74#_c_1608_n 0.0198473f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_422 N_CLK_c_503_n N_A_301_74#_c_1608_n 0.00273453f $X=3.235 $Y=1.557 $X2=0
+ $Y2=0
cc_423 N_CLK_c_504_n N_A_301_74#_c_1613_n 0.0185105f $X=3.235 $Y=1.765 $X2=0
+ $Y2=0
cc_424 CLK N_A_301_74#_c_1613_n 7.83337e-19 $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_425 N_CLK_M1000_g N_VGND_c_1800_n 0.00355958f $X=3.075 $Y=0.74 $X2=0 $Y2=0
cc_426 N_CLK_M1000_g N_VGND_c_1801_n 0.0037599f $X=3.075 $Y=0.74 $X2=0 $Y2=0
cc_427 N_CLK_M1000_g N_VGND_c_1811_n 0.00434272f $X=3.075 $Y=0.74 $X2=0 $Y2=0
cc_428 N_CLK_M1000_g N_VGND_c_1825_n 0.00826076f $X=3.075 $Y=0.74 $X2=0 $Y2=0
cc_429 N_A_828_74#_c_541_n N_A_630_74#_M1011_g 0.00158979f $X=4.28 $Y=0.515
+ $X2=0 $Y2=0
cc_430 N_A_828_74#_c_543_n N_A_630_74#_M1011_g 0.00266901f $X=4.445 $Y=0.34
+ $X2=0 $Y2=0
cc_431 N_A_828_74#_c_541_n N_A_630_74#_c_738_n 0.00206007f $X=4.28 $Y=0.515
+ $X2=0 $Y2=0
cc_432 N_A_828_74#_c_544_n N_A_630_74#_c_755_n 0.00321054f $X=5.155 $Y=2.005
+ $X2=0 $Y2=0
cc_433 N_A_828_74#_c_565_n N_A_630_74#_c_755_n 0.0050478f $X=5.17 $Y=2.17 $X2=0
+ $Y2=0
cc_434 N_A_828_74#_c_544_n N_A_630_74#_c_739_n 0.00894894f $X=5.155 $Y=2.005
+ $X2=0 $Y2=0
cc_435 N_A_828_74#_M1028_g N_A_630_74#_M1017_g 0.00631135f $X=5.79 $Y=0.695
+ $X2=0 $Y2=0
cc_436 N_A_828_74#_c_541_n N_A_630_74#_M1017_g 0.00316746f $X=4.28 $Y=0.515
+ $X2=0 $Y2=0
cc_437 N_A_828_74#_c_542_n N_A_630_74#_M1017_g 0.00929412f $X=5.07 $Y=0.34 $X2=0
+ $Y2=0
cc_438 N_A_828_74#_c_544_n N_A_630_74#_M1017_g 0.0313046f $X=5.155 $Y=2.005
+ $X2=0 $Y2=0
cc_439 N_A_828_74#_c_551_n N_A_630_74#_M1017_g 0.00216186f $X=5.155 $Y=0.34
+ $X2=0 $Y2=0
cc_440 N_A_828_74#_c_553_n N_A_630_74#_M1017_g 0.00465058f $X=5.84 $Y=1.21 $X2=0
+ $Y2=0
cc_441 N_A_828_74#_c_544_n N_A_630_74#_c_741_n 0.00917518f $X=5.155 $Y=2.005
+ $X2=0 $Y2=0
cc_442 N_A_828_74#_c_547_n N_A_630_74#_c_741_n 2.28181e-19 $X=6.84 $Y=0.855
+ $X2=0 $Y2=0
cc_443 N_A_828_74#_c_565_n N_A_630_74#_c_741_n 0.00735373f $X=5.17 $Y=2.17 $X2=0
+ $Y2=0
cc_444 N_A_828_74#_c_552_n N_A_630_74#_c_741_n 8.19781e-19 $X=5.915 $Y=0.855
+ $X2=0 $Y2=0
cc_445 N_A_828_74#_c_553_n N_A_630_74#_c_741_n 0.0181631f $X=5.84 $Y=1.21 $X2=0
+ $Y2=0
cc_446 N_A_828_74#_c_565_n N_A_630_74#_c_758_n 0.00364152f $X=5.17 $Y=2.17 $X2=0
+ $Y2=0
cc_447 N_A_828_74#_c_559_n N_A_630_74#_c_759_n 0.011667f $X=5.475 $Y=2.42 $X2=0
+ $Y2=0
cc_448 N_A_828_74#_c_565_n N_A_630_74#_c_759_n 0.00853179f $X=5.17 $Y=2.17 $X2=0
+ $Y2=0
cc_449 N_A_828_74#_c_561_n N_A_630_74#_c_760_n 0.0123454f $X=8.38 $Y=2.465 $X2=0
+ $Y2=0
cc_450 N_A_828_74#_c_563_n N_A_630_74#_c_760_n 0.00602601f $X=8.395 $Y=2.14
+ $X2=0 $Y2=0
cc_451 N_A_828_74#_c_550_n N_A_630_74#_c_742_n 0.012422f $X=8.35 $Y=1.31 $X2=0
+ $Y2=0
cc_452 N_A_828_74#_c_554_n N_A_630_74#_c_742_n 0.00145481f $X=7.615 $Y=1.195
+ $X2=0 $Y2=0
cc_453 N_A_828_74#_c_555_n N_A_630_74#_c_742_n 0.0212282f $X=7.615 $Y=1.195
+ $X2=0 $Y2=0
cc_454 N_A_828_74#_c_557_n N_A_630_74#_c_742_n 0.00114576f $X=8.515 $Y=1.31
+ $X2=0 $Y2=0
cc_455 N_A_828_74#_c_558_n N_A_630_74#_c_742_n 0.0172616f $X=8.515 $Y=1.39 $X2=0
+ $Y2=0
cc_456 N_A_828_74#_c_539_n N_A_630_74#_c_743_n 0.00579087f $X=7.48 $Y=1.03 $X2=0
+ $Y2=0
cc_457 N_A_828_74#_c_548_n N_A_630_74#_c_743_n 0.00218367f $X=7.52 $Y=0.34 $X2=0
+ $Y2=0
cc_458 N_A_828_74#_c_556_n N_A_630_74#_c_743_n 6.68163e-19 $X=7.65 $Y=1.03 $X2=0
+ $Y2=0
cc_459 N_A_828_74#_c_544_n N_A_630_74#_c_745_n 0.00454449f $X=5.155 $Y=2.005
+ $X2=0 $Y2=0
cc_460 N_A_828_74#_c_565_n N_A_630_74#_c_745_n 0.0181742f $X=5.17 $Y=2.17 $X2=0
+ $Y2=0
cc_461 N_A_828_74#_c_539_n N_A_630_74#_c_746_n 0.00384688f $X=7.48 $Y=1.03 $X2=0
+ $Y2=0
cc_462 N_A_828_74#_c_550_n N_A_630_74#_c_746_n 0.00111322f $X=8.35 $Y=1.31 $X2=0
+ $Y2=0
cc_463 N_A_828_74#_c_556_n N_A_630_74#_c_746_n 0.00125326f $X=7.65 $Y=1.03 $X2=0
+ $Y2=0
cc_464 N_A_828_74#_c_541_n N_A_630_74#_c_748_n 0.00581604f $X=4.28 $Y=0.515
+ $X2=0 $Y2=0
cc_465 N_A_828_74#_c_540_n N_A_630_74#_c_752_n 6.22426e-19 $X=8.395 $Y=1.99
+ $X2=0 $Y2=0
cc_466 N_A_828_74#_c_550_n N_A_630_74#_c_752_n 0.00747515f $X=8.35 $Y=1.31 $X2=0
+ $Y2=0
cc_467 N_A_828_74#_c_554_n N_A_630_74#_c_752_n 0.0159884f $X=7.615 $Y=1.195
+ $X2=0 $Y2=0
cc_468 N_A_828_74#_c_555_n N_A_630_74#_c_752_n 2.52598e-19 $X=7.615 $Y=1.195
+ $X2=0 $Y2=0
cc_469 N_A_828_74#_c_540_n N_A_630_74#_c_753_n 0.0227211f $X=8.395 $Y=1.99 $X2=0
+ $Y2=0
cc_470 N_A_828_74#_c_563_n N_A_630_74#_c_753_n 0.00142452f $X=8.395 $Y=2.14
+ $X2=0 $Y2=0
cc_471 N_A_828_74#_c_550_n N_A_630_74#_c_753_n 0.00417837f $X=8.35 $Y=1.31 $X2=0
+ $Y2=0
cc_472 N_A_828_74#_c_554_n N_A_630_74#_c_753_n 8.28969e-19 $X=7.615 $Y=1.195
+ $X2=0 $Y2=0
cc_473 N_A_828_74#_c_555_n N_A_630_74#_c_753_n 0.0118401f $X=7.615 $Y=1.195
+ $X2=0 $Y2=0
cc_474 N_A_828_74#_c_548_n N_A_1243_48#_M1018_d 0.00176461f $X=7.52 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_475 N_A_828_74#_M1028_g N_A_1243_48#_M1014_g 0.0184976f $X=5.79 $Y=0.695
+ $X2=0 $Y2=0
cc_476 N_A_828_74#_c_545_n N_A_1243_48#_M1014_g 0.00288087f $X=5.91 $Y=0.34
+ $X2=0 $Y2=0
cc_477 N_A_828_74#_c_546_n N_A_1243_48#_M1014_g 0.00514734f $X=5.995 $Y=0.77
+ $X2=0 $Y2=0
cc_478 N_A_828_74#_c_547_n N_A_1243_48#_M1014_g 0.0131292f $X=6.84 $Y=0.855
+ $X2=0 $Y2=0
cc_479 N_A_828_74#_c_616_p N_A_1243_48#_M1014_g 0.00235398f $X=6.925 $Y=0.77
+ $X2=0 $Y2=0
cc_480 N_A_828_74#_c_549_n N_A_1243_48#_M1014_g 3.8049e-19 $X=7.01 $Y=0.34 $X2=0
+ $Y2=0
cc_481 N_A_828_74#_c_552_n N_A_1243_48#_M1014_g 0.0055586f $X=5.915 $Y=0.855
+ $X2=0 $Y2=0
cc_482 N_A_828_74#_c_553_n N_A_1243_48#_M1014_g 0.0205366f $X=5.84 $Y=1.21 $X2=0
+ $Y2=0
cc_483 N_A_828_74#_c_547_n N_A_1243_48#_c_941_n 0.0591813f $X=6.84 $Y=0.855
+ $X2=0 $Y2=0
cc_484 N_A_828_74#_c_552_n N_A_1243_48#_c_941_n 0.0222623f $X=5.915 $Y=0.855
+ $X2=0 $Y2=0
cc_485 N_A_828_74#_c_553_n N_A_1243_48#_c_941_n 2.65259e-19 $X=5.84 $Y=1.21
+ $X2=0 $Y2=0
cc_486 N_A_828_74#_c_547_n N_A_1243_48#_c_942_n 0.00565722f $X=6.84 $Y=0.855
+ $X2=0 $Y2=0
cc_487 N_A_828_74#_c_539_n N_A_1243_48#_c_943_n 0.00139608f $X=7.48 $Y=1.03
+ $X2=0 $Y2=0
cc_488 N_A_828_74#_c_547_n N_A_1243_48#_c_943_n 0.00787896f $X=6.84 $Y=0.855
+ $X2=0 $Y2=0
cc_489 N_A_828_74#_c_548_n N_A_1243_48#_c_943_n 0.0126348f $X=7.52 $Y=0.34 $X2=0
+ $Y2=0
cc_490 N_A_828_74#_c_556_n N_A_1243_48#_c_943_n 0.0246758f $X=7.65 $Y=1.03 $X2=0
+ $Y2=0
cc_491 N_A_828_74#_c_554_n N_A_1243_48#_c_945_n 0.0237863f $X=7.615 $Y=1.195
+ $X2=0 $Y2=0
cc_492 N_A_828_74#_c_555_n N_A_1243_48#_c_945_n 0.00226443f $X=7.615 $Y=1.195
+ $X2=0 $Y2=0
cc_493 N_A_828_74#_c_544_n N_A_1021_97#_M1017_d 0.00470085f $X=5.155 $Y=2.005
+ $X2=-0.19 $Y2=-0.245
cc_494 N_A_828_74#_c_539_n N_A_1021_97#_M1018_g 0.0317322f $X=7.48 $Y=1.03 $X2=0
+ $Y2=0
cc_495 N_A_828_74#_c_547_n N_A_1021_97#_M1018_g 0.00565986f $X=6.84 $Y=0.855
+ $X2=0 $Y2=0
cc_496 N_A_828_74#_c_616_p N_A_1021_97#_M1018_g 0.00925239f $X=6.925 $Y=0.77
+ $X2=0 $Y2=0
cc_497 N_A_828_74#_c_548_n N_A_1021_97#_M1018_g 0.00937415f $X=7.52 $Y=0.34
+ $X2=0 $Y2=0
cc_498 N_A_828_74#_c_549_n N_A_1021_97#_M1018_g 0.00288658f $X=7.01 $Y=0.34
+ $X2=0 $Y2=0
cc_499 N_A_828_74#_c_554_n N_A_1021_97#_M1018_g 3.42484e-19 $X=7.615 $Y=1.195
+ $X2=0 $Y2=0
cc_500 N_A_828_74#_c_556_n N_A_1021_97#_M1018_g 6.06864e-19 $X=7.65 $Y=1.03
+ $X2=0 $Y2=0
cc_501 N_A_828_74#_M1028_g N_A_1021_97#_c_1011_n 0.00177723f $X=5.79 $Y=0.695
+ $X2=0 $Y2=0
cc_502 N_A_828_74#_c_552_n N_A_1021_97#_c_1011_n 0.0323932f $X=5.915 $Y=0.855
+ $X2=0 $Y2=0
cc_503 N_A_828_74#_c_553_n N_A_1021_97#_c_1011_n 0.00361611f $X=5.84 $Y=1.21
+ $X2=0 $Y2=0
cc_504 N_A_828_74#_c_547_n N_A_1021_97#_c_1012_n 0.00495776f $X=6.84 $Y=0.855
+ $X2=0 $Y2=0
cc_505 N_A_828_74#_c_552_n N_A_1021_97#_c_1012_n 0.0230462f $X=5.915 $Y=0.855
+ $X2=0 $Y2=0
cc_506 N_A_828_74#_c_553_n N_A_1021_97#_c_1012_n 0.00230734f $X=5.84 $Y=1.21
+ $X2=0 $Y2=0
cc_507 N_A_828_74#_M1028_g N_A_1021_97#_c_1034_n 0.00418303f $X=5.79 $Y=0.695
+ $X2=0 $Y2=0
cc_508 N_A_828_74#_c_544_n N_A_1021_97#_c_1034_n 0.0739505f $X=5.155 $Y=2.005
+ $X2=0 $Y2=0
cc_509 N_A_828_74#_c_545_n N_A_1021_97#_c_1034_n 0.0224673f $X=5.91 $Y=0.34
+ $X2=0 $Y2=0
cc_510 N_A_828_74#_c_544_n N_A_1021_97#_c_1013_n 0.0132809f $X=5.155 $Y=2.005
+ $X2=0 $Y2=0
cc_511 N_A_828_74#_c_565_n N_A_1021_97#_c_1013_n 6.34912e-19 $X=5.17 $Y=2.17
+ $X2=0 $Y2=0
cc_512 N_A_828_74#_c_559_n N_A_1021_97#_c_1017_n 0.00757202f $X=5.475 $Y=2.42
+ $X2=0 $Y2=0
cc_513 N_A_828_74#_c_559_n N_A_1021_97#_c_1018_n 0.00270086f $X=5.475 $Y=2.42
+ $X2=0 $Y2=0
cc_514 N_A_828_74#_c_544_n N_A_1021_97#_c_1018_n 0.0386717f $X=5.155 $Y=2.005
+ $X2=0 $Y2=0
cc_515 N_A_828_74#_c_565_n N_A_1021_97#_c_1018_n 0.0105257f $X=5.17 $Y=2.17
+ $X2=0 $Y2=0
cc_516 N_A_828_74#_c_558_n N_A_1711_48#_c_1094_n 0.00814818f $X=8.515 $Y=1.39
+ $X2=0 $Y2=0
cc_517 N_A_828_74#_c_560_n N_A_1711_48#_c_1111_n 0.0169882f $X=8.38 $Y=2.375
+ $X2=0 $Y2=0
cc_518 N_A_828_74#_c_561_n N_A_1711_48#_c_1111_n 0.0283714f $X=8.38 $Y=2.465
+ $X2=0 $Y2=0
cc_519 N_A_828_74#_c_563_n N_A_1711_48#_c_1111_n 0.00555967f $X=8.395 $Y=2.14
+ $X2=0 $Y2=0
cc_520 N_A_828_74#_c_540_n N_A_1711_48#_c_1095_n 0.0146785f $X=8.395 $Y=1.99
+ $X2=0 $Y2=0
cc_521 N_A_828_74#_c_557_n N_A_1711_48#_c_1095_n 3.80732e-19 $X=8.515 $Y=1.31
+ $X2=0 $Y2=0
cc_522 N_A_828_74#_c_558_n N_A_1711_48#_c_1095_n 0.0205378f $X=8.515 $Y=1.39
+ $X2=0 $Y2=0
cc_523 N_A_828_74#_c_560_n N_A_1711_48#_c_1118_n 9.02254e-19 $X=8.38 $Y=2.375
+ $X2=0 $Y2=0
cc_524 N_A_828_74#_c_563_n N_A_1711_48#_c_1118_n 3.0415e-19 $X=8.395 $Y=2.14
+ $X2=0 $Y2=0
cc_525 N_A_828_74#_c_548_n N_A_1511_74#_M1033_d 5.36554e-19 $X=7.52 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_526 N_A_828_74#_c_556_n N_A_1511_74#_M1033_d 0.00492103f $X=7.65 $Y=1.03
+ $X2=-0.19 $Y2=-0.245
cc_527 N_A_828_74#_c_560_n N_A_1511_74#_c_1267_n 0.00282381f $X=8.38 $Y=2.375
+ $X2=0 $Y2=0
cc_528 N_A_828_74#_c_561_n N_A_1511_74#_c_1268_n 0.0128811f $X=8.38 $Y=2.465
+ $X2=0 $Y2=0
cc_529 N_A_828_74#_c_550_n N_A_1511_74#_c_1257_n 0.012009f $X=8.35 $Y=1.31 $X2=0
+ $Y2=0
cc_530 N_A_828_74#_c_557_n N_A_1511_74#_c_1257_n 0.0247442f $X=8.515 $Y=1.31
+ $X2=0 $Y2=0
cc_531 N_A_828_74#_c_558_n N_A_1511_74#_c_1257_n 0.00178652f $X=8.515 $Y=1.39
+ $X2=0 $Y2=0
cc_532 N_A_828_74#_c_540_n N_A_1511_74#_c_1269_n 0.0154537f $X=8.395 $Y=1.99
+ $X2=0 $Y2=0
cc_533 N_A_828_74#_c_563_n N_A_1511_74#_c_1269_n 0.00265181f $X=8.395 $Y=2.14
+ $X2=0 $Y2=0
cc_534 N_A_828_74#_c_550_n N_A_1511_74#_c_1269_n 0.00550527f $X=8.35 $Y=1.31
+ $X2=0 $Y2=0
cc_535 N_A_828_74#_c_557_n N_A_1511_74#_c_1269_n 0.0241867f $X=8.515 $Y=1.31
+ $X2=0 $Y2=0
cc_536 N_A_828_74#_c_558_n N_A_1511_74#_c_1269_n 0.00406216f $X=8.515 $Y=1.39
+ $X2=0 $Y2=0
cc_537 N_A_828_74#_c_550_n N_A_1511_74#_c_1270_n 0.00850562f $X=8.35 $Y=1.31
+ $X2=0 $Y2=0
cc_538 N_A_828_74#_c_540_n N_A_1511_74#_c_1258_n 0.0028736f $X=8.395 $Y=1.99
+ $X2=0 $Y2=0
cc_539 N_A_828_74#_c_557_n N_A_1511_74#_c_1258_n 0.0243882f $X=8.515 $Y=1.31
+ $X2=0 $Y2=0
cc_540 N_A_828_74#_c_558_n N_A_1511_74#_c_1258_n 0.0018137f $X=8.515 $Y=1.39
+ $X2=0 $Y2=0
cc_541 N_A_828_74#_c_539_n N_A_1511_74#_c_1260_n 0.00179f $X=7.48 $Y=1.03 $X2=0
+ $Y2=0
cc_542 N_A_828_74#_c_548_n N_A_1511_74#_c_1260_n 0.00648406f $X=7.52 $Y=0.34
+ $X2=0 $Y2=0
cc_543 N_A_828_74#_c_550_n N_A_1511_74#_c_1260_n 0.0203321f $X=8.35 $Y=1.31
+ $X2=0 $Y2=0
cc_544 N_A_828_74#_c_554_n N_A_1511_74#_c_1260_n 0.00148722f $X=7.615 $Y=1.195
+ $X2=0 $Y2=0
cc_545 N_A_828_74#_c_556_n N_A_1511_74#_c_1260_n 0.0398855f $X=7.65 $Y=1.03
+ $X2=0 $Y2=0
cc_546 N_A_828_74#_c_540_n N_A_1511_74#_c_1272_n 0.00234025f $X=8.395 $Y=1.99
+ $X2=0 $Y2=0
cc_547 N_A_828_74#_c_563_n N_A_1511_74#_c_1272_n 0.00282381f $X=8.395 $Y=2.14
+ $X2=0 $Y2=0
cc_548 N_A_828_74#_c_561_n N_VPWR_c_1443_n 0.00152232f $X=8.38 $Y=2.465 $X2=0
+ $Y2=0
cc_549 N_A_828_74#_c_559_n N_VPWR_c_1456_n 0.00500196f $X=5.475 $Y=2.42 $X2=0
+ $Y2=0
cc_550 N_A_828_74#_c_561_n N_VPWR_c_1460_n 0.00461464f $X=8.38 $Y=2.465 $X2=0
+ $Y2=0
cc_551 N_A_828_74#_c_559_n N_VPWR_c_1439_n 0.005315f $X=5.475 $Y=2.42 $X2=0
+ $Y2=0
cc_552 N_A_828_74#_c_561_n N_VPWR_c_1439_n 0.00983553f $X=8.38 $Y=2.465 $X2=0
+ $Y2=0
cc_553 N_A_828_74#_c_544_n N_A_301_74#_c_1614_n 0.0362105f $X=5.155 $Y=2.005
+ $X2=0 $Y2=0
cc_554 N_A_828_74#_c_565_n N_A_301_74#_c_1614_n 3.12271e-19 $X=5.17 $Y=2.17
+ $X2=0 $Y2=0
cc_555 N_A_828_74#_c_541_n N_A_301_74#_c_1609_n 4.37372e-19 $X=4.28 $Y=0.515
+ $X2=0 $Y2=0
cc_556 N_A_828_74#_c_544_n N_A_301_74#_c_1609_n 0.0343342f $X=5.155 $Y=2.005
+ $X2=0 $Y2=0
cc_557 N_A_828_74#_c_541_n N_A_301_74#_c_1610_n 0.00962346f $X=4.28 $Y=0.515
+ $X2=0 $Y2=0
cc_558 N_A_828_74#_c_541_n N_A_301_74#_c_1611_n 0.0374588f $X=4.28 $Y=0.515
+ $X2=0 $Y2=0
cc_559 N_A_828_74#_c_542_n N_A_301_74#_c_1611_n 0.0192119f $X=5.07 $Y=0.34 $X2=0
+ $Y2=0
cc_560 N_A_828_74#_c_544_n N_A_301_74#_c_1611_n 0.0528515f $X=5.155 $Y=2.005
+ $X2=0 $Y2=0
cc_561 N_A_828_74#_M1031_d N_A_301_74#_c_1615_n 0.00364477f $X=4.54 $Y=1.84
+ $X2=0 $Y2=0
cc_562 N_A_828_74#_c_544_n N_A_301_74#_c_1615_n 0.020128f $X=5.155 $Y=2.005
+ $X2=0 $Y2=0
cc_563 N_A_828_74#_c_565_n N_A_301_74#_c_1615_n 0.00181381f $X=5.17 $Y=2.17
+ $X2=0 $Y2=0
cc_564 N_A_828_74#_M1031_d N_A_301_74#_c_1665_n 0.00742992f $X=4.54 $Y=1.84
+ $X2=0 $Y2=0
cc_565 N_A_828_74#_c_559_n N_A_301_74#_c_1665_n 0.0018585f $X=5.475 $Y=2.42
+ $X2=0 $Y2=0
cc_566 N_A_828_74#_c_544_n N_A_301_74#_c_1665_n 0.0113655f $X=5.155 $Y=2.005
+ $X2=0 $Y2=0
cc_567 N_A_828_74#_c_565_n N_A_301_74#_c_1665_n 0.0012864f $X=5.17 $Y=2.17 $X2=0
+ $Y2=0
cc_568 N_A_828_74#_c_559_n N_A_301_74#_c_1617_n 0.0022555f $X=5.475 $Y=2.42
+ $X2=0 $Y2=0
cc_569 N_A_828_74#_c_544_n N_A_301_74#_c_1617_n 0.0205765f $X=5.155 $Y=2.005
+ $X2=0 $Y2=0
cc_570 N_A_828_74#_c_565_n N_A_301_74#_c_1617_n 0.00576151f $X=5.17 $Y=2.17
+ $X2=0 $Y2=0
cc_571 N_A_828_74#_c_547_n N_VGND_M1014_d 0.00655131f $X=6.84 $Y=0.855 $X2=0
+ $Y2=0
cc_572 N_A_828_74#_c_616_p N_VGND_M1014_d 0.004181f $X=6.925 $Y=0.77 $X2=0 $Y2=0
cc_573 N_A_828_74#_c_549_n N_VGND_M1014_d 5.37788e-19 $X=7.01 $Y=0.34 $X2=0
+ $Y2=0
cc_574 N_A_828_74#_c_543_n N_VGND_c_1801_n 0.0112234f $X=4.445 $Y=0.34 $X2=0
+ $Y2=0
cc_575 N_A_828_74#_c_545_n N_VGND_c_1802_n 0.0103385f $X=5.91 $Y=0.34 $X2=0
+ $Y2=0
cc_576 N_A_828_74#_c_546_n N_VGND_c_1802_n 0.00929617f $X=5.995 $Y=0.77 $X2=0
+ $Y2=0
cc_577 N_A_828_74#_c_547_n N_VGND_c_1802_n 0.0212699f $X=6.84 $Y=0.855 $X2=0
+ $Y2=0
cc_578 N_A_828_74#_c_616_p N_VGND_c_1802_n 0.0133374f $X=6.925 $Y=0.77 $X2=0
+ $Y2=0
cc_579 N_A_828_74#_c_549_n N_VGND_c_1802_n 0.0148563f $X=7.01 $Y=0.34 $X2=0
+ $Y2=0
cc_580 N_A_828_74#_M1028_g N_VGND_c_1813_n 7.35405e-19 $X=5.79 $Y=0.695 $X2=0
+ $Y2=0
cc_581 N_A_828_74#_c_542_n N_VGND_c_1813_n 0.0402032f $X=5.07 $Y=0.34 $X2=0
+ $Y2=0
cc_582 N_A_828_74#_c_543_n N_VGND_c_1813_n 0.0179217f $X=4.445 $Y=0.34 $X2=0
+ $Y2=0
cc_583 N_A_828_74#_c_545_n N_VGND_c_1813_n 0.0552887f $X=5.91 $Y=0.34 $X2=0
+ $Y2=0
cc_584 N_A_828_74#_c_551_n N_VGND_c_1813_n 0.0121867f $X=5.155 $Y=0.34 $X2=0
+ $Y2=0
cc_585 N_A_828_74#_c_539_n N_VGND_c_1814_n 0.00278237f $X=7.48 $Y=1.03 $X2=0
+ $Y2=0
cc_586 N_A_828_74#_c_548_n N_VGND_c_1814_n 0.0441951f $X=7.52 $Y=0.34 $X2=0
+ $Y2=0
cc_587 N_A_828_74#_c_549_n N_VGND_c_1814_n 0.0120704f $X=7.01 $Y=0.34 $X2=0
+ $Y2=0
cc_588 N_A_828_74#_c_539_n N_VGND_c_1825_n 0.00355939f $X=7.48 $Y=1.03 $X2=0
+ $Y2=0
cc_589 N_A_828_74#_c_542_n N_VGND_c_1825_n 0.0234906f $X=5.07 $Y=0.34 $X2=0
+ $Y2=0
cc_590 N_A_828_74#_c_543_n N_VGND_c_1825_n 0.00971942f $X=4.445 $Y=0.34 $X2=0
+ $Y2=0
cc_591 N_A_828_74#_c_545_n N_VGND_c_1825_n 0.0317917f $X=5.91 $Y=0.34 $X2=0
+ $Y2=0
cc_592 N_A_828_74#_c_547_n N_VGND_c_1825_n 0.0160936f $X=6.84 $Y=0.855 $X2=0
+ $Y2=0
cc_593 N_A_828_74#_c_548_n N_VGND_c_1825_n 0.0245704f $X=7.52 $Y=0.34 $X2=0
+ $Y2=0
cc_594 N_A_828_74#_c_549_n N_VGND_c_1825_n 0.00645034f $X=7.01 $Y=0.34 $X2=0
+ $Y2=0
cc_595 N_A_828_74#_c_551_n N_VGND_c_1825_n 0.00660921f $X=5.155 $Y=0.34 $X2=0
+ $Y2=0
cc_596 N_A_828_74#_c_545_n A_1173_97# 6.68967e-19 $X=5.91 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_597 N_A_828_74#_c_546_n A_1173_97# 0.00496712f $X=5.995 $Y=0.77 $X2=-0.19
+ $Y2=-0.245
cc_598 N_A_828_74#_c_547_n A_1173_97# 0.00145432f $X=6.84 $Y=0.855 $X2=-0.19
+ $Y2=-0.245
cc_599 N_A_828_74#_c_552_n A_1173_97# 5.94185e-19 $X=5.915 $Y=0.855 $X2=-0.19
+ $Y2=-0.245
cc_600 N_A_630_74#_c_831_p N_A_1243_48#_M1038_d 0.0208715f $X=7.565 $Y=2.7 $X2=0
+ $Y2=0
cc_601 N_A_630_74#_c_767_n N_A_1243_48#_M1038_d 0.00950379f $X=7.65 $Y=2.615
+ $X2=0 $Y2=0
cc_602 N_A_630_74#_c_741_n N_A_1243_48#_c_940_n 0.0394473f $X=5.8 $Y=1.69 $X2=0
+ $Y2=0
cc_603 N_A_630_74#_c_759_n N_A_1243_48#_c_940_n 0.00873558f $X=6.01 $Y=2.42
+ $X2=0 $Y2=0
cc_604 N_A_630_74#_c_766_n N_A_1243_48#_c_940_n 0.00371687f $X=6.12 $Y=2.615
+ $X2=0 $Y2=0
cc_605 N_A_630_74#_c_768_n N_A_1243_48#_c_940_n 0.00757656f $X=6.12 $Y=2.08
+ $X2=0 $Y2=0
cc_606 N_A_630_74#_c_759_n N_A_1243_48#_c_947_n 0.0288723f $X=6.01 $Y=2.42 $X2=0
+ $Y2=0
cc_607 N_A_630_74#_c_766_n N_A_1243_48#_c_947_n 0.0040898f $X=6.12 $Y=2.615
+ $X2=0 $Y2=0
cc_608 N_A_630_74#_c_831_p N_A_1243_48#_c_947_n 0.0163967f $X=7.565 $Y=2.7 $X2=0
+ $Y2=0
cc_609 N_A_630_74#_c_831_p N_A_1243_48#_c_948_n 0.0180145f $X=7.565 $Y=2.7 $X2=0
+ $Y2=0
cc_610 N_A_630_74#_c_767_n N_A_1243_48#_c_948_n 0.0249467f $X=7.65 $Y=2.615
+ $X2=0 $Y2=0
cc_611 N_A_630_74#_c_742_n N_A_1243_48#_c_944_n 0.00408593f $X=8.065 $Y=1.6
+ $X2=0 $Y2=0
cc_612 N_A_630_74#_c_752_n N_A_1243_48#_c_944_n 0.0325509f $X=7.73 $Y=1.765
+ $X2=0 $Y2=0
cc_613 N_A_630_74#_c_753_n N_A_1243_48#_c_944_n 0.00269918f $X=7.845 $Y=1.822
+ $X2=0 $Y2=0
cc_614 N_A_630_74#_c_742_n N_A_1243_48#_c_945_n 2.64577e-19 $X=8.065 $Y=1.6
+ $X2=0 $Y2=0
cc_615 N_A_630_74#_c_753_n N_A_1021_97#_M1018_g 2.97215e-19 $X=7.845 $Y=1.822
+ $X2=0 $Y2=0
cc_616 N_A_630_74#_c_760_n N_A_1021_97#_c_1010_n 0.0127665f $X=7.845 $Y=2.045
+ $X2=0 $Y2=0
cc_617 N_A_630_74#_c_831_p N_A_1021_97#_c_1010_n 0.0179214f $X=7.565 $Y=2.7
+ $X2=0 $Y2=0
cc_618 N_A_630_74#_c_767_n N_A_1021_97#_c_1010_n 0.00323365f $X=7.65 $Y=2.615
+ $X2=0 $Y2=0
cc_619 N_A_630_74#_c_753_n N_A_1021_97#_c_1010_n 0.008321f $X=7.845 $Y=1.822
+ $X2=0 $Y2=0
cc_620 N_A_630_74#_c_741_n N_A_1021_97#_c_1012_n 0.0205571f $X=5.8 $Y=1.69 $X2=0
+ $Y2=0
cc_621 N_A_630_74#_c_768_n N_A_1021_97#_c_1012_n 0.026299f $X=6.12 $Y=2.08 $X2=0
+ $Y2=0
cc_622 N_A_630_74#_M1017_g N_A_1021_97#_c_1034_n 0.00331691f $X=5.03 $Y=0.695
+ $X2=0 $Y2=0
cc_623 N_A_630_74#_M1017_g N_A_1021_97#_c_1013_n 2.27645e-19 $X=5.03 $Y=0.695
+ $X2=0 $Y2=0
cc_624 N_A_630_74#_c_741_n N_A_1021_97#_c_1013_n 0.0122841f $X=5.8 $Y=1.69 $X2=0
+ $Y2=0
cc_625 N_A_630_74#_c_759_n N_A_1021_97#_c_1017_n 0.00929725f $X=6.01 $Y=2.42
+ $X2=0 $Y2=0
cc_626 N_A_630_74#_c_766_n N_A_1021_97#_c_1017_n 0.010429f $X=6.12 $Y=2.615
+ $X2=0 $Y2=0
cc_627 N_A_630_74#_c_858_p N_A_1021_97#_c_1017_n 0.014098f $X=6.205 $Y=2.7 $X2=0
+ $Y2=0
cc_628 N_A_630_74#_c_768_n N_A_1021_97#_c_1017_n 0.00123739f $X=6.12 $Y=2.08
+ $X2=0 $Y2=0
cc_629 N_A_630_74#_c_741_n N_A_1021_97#_c_1018_n 0.00457114f $X=5.8 $Y=1.69
+ $X2=0 $Y2=0
cc_630 N_A_630_74#_c_758_n N_A_1021_97#_c_1018_n 0.0100595f $X=5.965 $Y=2.08
+ $X2=0 $Y2=0
cc_631 N_A_630_74#_c_759_n N_A_1021_97#_c_1018_n 0.00170079f $X=6.01 $Y=2.42
+ $X2=0 $Y2=0
cc_632 N_A_630_74#_c_766_n N_A_1021_97#_c_1018_n 0.00937204f $X=6.12 $Y=2.615
+ $X2=0 $Y2=0
cc_633 N_A_630_74#_c_768_n N_A_1021_97#_c_1018_n 0.0248982f $X=6.12 $Y=2.08
+ $X2=0 $Y2=0
cc_634 N_A_630_74#_c_831_p N_A_1021_97#_c_1014_n 0.00616686f $X=7.565 $Y=2.7
+ $X2=0 $Y2=0
cc_635 N_A_630_74#_c_768_n N_A_1021_97#_c_1014_n 9.7786e-19 $X=6.12 $Y=2.08
+ $X2=0 $Y2=0
cc_636 N_A_630_74#_c_743_n N_A_1711_48#_c_1092_n 0.0199822f $X=8.24 $Y=0.865
+ $X2=0 $Y2=0
cc_637 N_A_630_74#_c_746_n N_A_1711_48#_c_1094_n 0.0199822f $X=8.24 $Y=0.94
+ $X2=0 $Y2=0
cc_638 N_A_630_74#_c_760_n N_A_1511_74#_c_1267_n 0.00256776f $X=7.845 $Y=2.045
+ $X2=0 $Y2=0
cc_639 N_A_630_74#_c_767_n N_A_1511_74#_c_1267_n 0.0200013f $X=7.65 $Y=2.615
+ $X2=0 $Y2=0
cc_640 N_A_630_74#_c_753_n N_A_1511_74#_c_1267_n 0.00564347f $X=7.845 $Y=1.822
+ $X2=0 $Y2=0
cc_641 N_A_630_74#_c_760_n N_A_1511_74#_c_1268_n 0.0159121f $X=7.845 $Y=2.045
+ $X2=0 $Y2=0
cc_642 N_A_630_74#_c_746_n N_A_1511_74#_c_1257_n 0.00996416f $X=8.24 $Y=0.94
+ $X2=0 $Y2=0
cc_643 N_A_630_74#_c_752_n N_A_1511_74#_c_1270_n 0.0142007f $X=7.73 $Y=1.765
+ $X2=0 $Y2=0
cc_644 N_A_630_74#_c_753_n N_A_1511_74#_c_1270_n 0.00569571f $X=7.845 $Y=1.822
+ $X2=0 $Y2=0
cc_645 N_A_630_74#_c_742_n N_A_1511_74#_c_1260_n 0.00338372f $X=8.065 $Y=1.6
+ $X2=0 $Y2=0
cc_646 N_A_630_74#_c_743_n N_A_1511_74#_c_1260_n 0.0107359f $X=8.24 $Y=0.865
+ $X2=0 $Y2=0
cc_647 N_A_630_74#_c_746_n N_A_1511_74#_c_1260_n 0.00913705f $X=8.24 $Y=0.94
+ $X2=0 $Y2=0
cc_648 N_A_630_74#_c_760_n N_A_1511_74#_c_1272_n 4.67692e-19 $X=7.845 $Y=2.045
+ $X2=0 $Y2=0
cc_649 N_A_630_74#_c_767_n N_A_1511_74#_c_1272_n 0.00801539f $X=7.65 $Y=2.615
+ $X2=0 $Y2=0
cc_650 N_A_630_74#_c_752_n N_A_1511_74#_c_1272_n 0.00296848f $X=7.73 $Y=1.765
+ $X2=0 $Y2=0
cc_651 N_A_630_74#_c_753_n N_A_1511_74#_c_1272_n 0.00141097f $X=7.845 $Y=1.822
+ $X2=0 $Y2=0
cc_652 N_A_630_74#_c_763_n N_VPWR_M1031_s 0.00228424f $X=3.855 $Y=2.075 $X2=0
+ $Y2=0
cc_653 N_A_630_74#_c_831_p N_VPWR_M1004_d 0.0146075f $X=7.565 $Y=2.7 $X2=0 $Y2=0
cc_654 N_A_630_74#_c_755_n N_VPWR_c_1442_n 0.0191626f $X=4.465 $Y=1.765 $X2=0
+ $Y2=0
cc_655 N_A_630_74#_c_831_p N_VPWR_c_1455_n 0.0242646f $X=7.565 $Y=2.7 $X2=0
+ $Y2=0
cc_656 N_A_630_74#_c_755_n N_VPWR_c_1456_n 0.00413917f $X=4.465 $Y=1.765 $X2=0
+ $Y2=0
cc_657 N_A_630_74#_c_759_n N_VPWR_c_1456_n 0.00499599f $X=6.01 $Y=2.42 $X2=0
+ $Y2=0
cc_658 N_A_630_74#_c_831_p N_VPWR_c_1456_n 0.00675146f $X=7.565 $Y=2.7 $X2=0
+ $Y2=0
cc_659 N_A_630_74#_c_858_p N_VPWR_c_1456_n 0.00326019f $X=6.205 $Y=2.7 $X2=0
+ $Y2=0
cc_660 N_A_630_74#_c_760_n N_VPWR_c_1460_n 0.00445602f $X=7.845 $Y=2.045 $X2=0
+ $Y2=0
cc_661 N_A_630_74#_c_831_p N_VPWR_c_1460_n 0.0167786f $X=7.565 $Y=2.7 $X2=0
+ $Y2=0
cc_662 N_A_630_74#_c_755_n N_VPWR_c_1439_n 0.00407755f $X=4.465 $Y=1.765 $X2=0
+ $Y2=0
cc_663 N_A_630_74#_c_759_n N_VPWR_c_1439_n 0.005315f $X=6.01 $Y=2.42 $X2=0 $Y2=0
cc_664 N_A_630_74#_c_760_n N_VPWR_c_1439_n 0.00861536f $X=7.845 $Y=2.045 $X2=0
+ $Y2=0
cc_665 N_A_630_74#_c_831_p N_VPWR_c_1439_n 0.0379767f $X=7.565 $Y=2.7 $X2=0
+ $Y2=0
cc_666 N_A_630_74#_c_858_p N_VPWR_c_1439_n 0.00538561f $X=6.205 $Y=2.7 $X2=0
+ $Y2=0
cc_667 N_A_630_74#_c_763_n N_A_301_74#_c_1608_n 0.0171788f $X=3.855 $Y=2.075
+ $X2=0 $Y2=0
cc_668 N_A_630_74#_M1001_d N_A_301_74#_c_1613_n 0.0162485f $X=3.31 $Y=1.84 $X2=0
+ $Y2=0
cc_669 N_A_630_74#_c_763_n N_A_301_74#_c_1613_n 0.0578524f $X=3.855 $Y=2.075
+ $X2=0 $Y2=0
cc_670 N_A_630_74#_c_750_n N_A_301_74#_c_1613_n 0.00506726f $X=3.975 $Y=1.515
+ $X2=0 $Y2=0
cc_671 N_A_630_74#_c_738_n N_A_301_74#_c_1614_n 0.00583402f $X=4.39 $Y=1.69
+ $X2=0 $Y2=0
cc_672 N_A_630_74#_c_755_n N_A_301_74#_c_1614_n 0.0201f $X=4.465 $Y=1.765 $X2=0
+ $Y2=0
cc_673 N_A_630_74#_c_744_n N_A_301_74#_c_1614_n 0.00367614f $X=4.465 $Y=1.69
+ $X2=0 $Y2=0
cc_674 N_A_630_74#_c_763_n N_A_301_74#_c_1614_n 0.0203395f $X=3.855 $Y=2.075
+ $X2=0 $Y2=0
cc_675 N_A_630_74#_c_764_n N_A_301_74#_c_1614_n 0.0220906f $X=3.975 $Y=1.515
+ $X2=0 $Y2=0
cc_676 N_A_630_74#_c_739_n N_A_301_74#_c_1609_n 0.0157016f $X=4.955 $Y=1.69
+ $X2=0 $Y2=0
cc_677 N_A_630_74#_M1017_g N_A_301_74#_c_1609_n 0.00307597f $X=5.03 $Y=0.695
+ $X2=0 $Y2=0
cc_678 N_A_630_74#_c_744_n N_A_301_74#_c_1609_n 0.00670241f $X=4.465 $Y=1.69
+ $X2=0 $Y2=0
cc_679 N_A_630_74#_c_738_n N_A_301_74#_c_1610_n 0.00301454f $X=4.39 $Y=1.69
+ $X2=0 $Y2=0
cc_680 N_A_630_74#_c_744_n N_A_301_74#_c_1610_n 9.14984e-19 $X=4.465 $Y=1.69
+ $X2=0 $Y2=0
cc_681 N_A_630_74#_c_764_n N_A_301_74#_c_1610_n 0.0137931f $X=3.975 $Y=1.515
+ $X2=0 $Y2=0
cc_682 N_A_630_74#_c_750_n N_A_301_74#_c_1610_n 0.00330803f $X=3.975 $Y=1.515
+ $X2=0 $Y2=0
cc_683 N_A_630_74#_M1011_g N_A_301_74#_c_1611_n 0.00663286f $X=4.065 $Y=0.74
+ $X2=0 $Y2=0
cc_684 N_A_630_74#_M1017_g N_A_301_74#_c_1611_n 0.0127542f $X=5.03 $Y=0.695
+ $X2=0 $Y2=0
cc_685 N_A_630_74#_c_748_n N_A_301_74#_c_1611_n 0.00151783f $X=3.855 $Y=1.095
+ $X2=0 $Y2=0
cc_686 N_A_630_74#_c_781_n N_A_301_74#_c_1611_n 0.00400785f $X=3.975 $Y=1.47
+ $X2=0 $Y2=0
cc_687 N_A_630_74#_c_751_n N_A_301_74#_c_1611_n 0.00466727f $X=3.975 $Y=1.35
+ $X2=0 $Y2=0
cc_688 N_A_630_74#_c_755_n N_A_301_74#_c_1665_n 0.017739f $X=4.465 $Y=1.765
+ $X2=0 $Y2=0
cc_689 N_A_630_74#_c_755_n N_A_301_74#_c_1617_n 0.00666737f $X=4.465 $Y=1.765
+ $X2=0 $Y2=0
cc_690 N_A_630_74#_c_766_n A_1217_499# 0.0013628f $X=6.12 $Y=2.615 $X2=-0.19
+ $Y2=-0.245
cc_691 N_A_630_74#_c_831_p A_1217_499# 0.00494057f $X=7.565 $Y=2.7 $X2=-0.19
+ $Y2=-0.245
cc_692 N_A_630_74#_c_858_p A_1217_499# 0.001001f $X=6.205 $Y=2.7 $X2=-0.19
+ $Y2=-0.245
cc_693 N_A_630_74#_c_748_n N_VGND_M1011_s 0.00302243f $X=3.855 $Y=1.095 $X2=0
+ $Y2=0
cc_694 N_A_630_74#_c_747_n N_VGND_c_1800_n 0.0243474f $X=3.29 $Y=0.515 $X2=0
+ $Y2=0
cc_695 N_A_630_74#_c_749_n N_VGND_c_1800_n 0.00555794f $X=3.455 $Y=1.095 $X2=0
+ $Y2=0
cc_696 N_A_630_74#_M1011_g N_VGND_c_1801_n 0.0120174f $X=4.065 $Y=0.74 $X2=0
+ $Y2=0
cc_697 N_A_630_74#_c_747_n N_VGND_c_1801_n 0.033035f $X=3.29 $Y=0.515 $X2=0
+ $Y2=0
cc_698 N_A_630_74#_c_748_n N_VGND_c_1801_n 0.0228363f $X=3.855 $Y=1.095 $X2=0
+ $Y2=0
cc_699 N_A_630_74#_c_750_n N_VGND_c_1801_n 5.13376e-19 $X=3.975 $Y=1.515 $X2=0
+ $Y2=0
cc_700 N_A_630_74#_c_747_n N_VGND_c_1811_n 0.0145639f $X=3.29 $Y=0.515 $X2=0
+ $Y2=0
cc_701 N_A_630_74#_M1011_g N_VGND_c_1813_n 0.00383152f $X=4.065 $Y=0.74 $X2=0
+ $Y2=0
cc_702 N_A_630_74#_M1017_g N_VGND_c_1813_n 7.53287e-19 $X=5.03 $Y=0.695 $X2=0
+ $Y2=0
cc_703 N_A_630_74#_c_743_n N_VGND_c_1814_n 0.00433139f $X=8.24 $Y=0.865 $X2=0
+ $Y2=0
cc_704 N_A_630_74#_c_743_n N_VGND_c_1821_n 0.00158462f $X=8.24 $Y=0.865 $X2=0
+ $Y2=0
cc_705 N_A_630_74#_M1011_g N_VGND_c_1825_n 0.00762539f $X=4.065 $Y=0.74 $X2=0
+ $Y2=0
cc_706 N_A_630_74#_c_743_n N_VGND_c_1825_n 0.00819726f $X=8.24 $Y=0.865 $X2=0
+ $Y2=0
cc_707 N_A_630_74#_c_747_n N_VGND_c_1825_n 0.0119984f $X=3.29 $Y=0.515 $X2=0
+ $Y2=0
cc_708 N_A_1243_48#_M1014_g N_A_1021_97#_M1018_g 0.0103168f $X=6.29 $Y=0.58
+ $X2=0 $Y2=0
cc_709 N_A_1243_48#_c_940_n N_A_1021_97#_M1018_g 0.00574023f $X=6.43 $Y=2.33
+ $X2=0 $Y2=0
cc_710 N_A_1243_48#_c_941_n N_A_1021_97#_M1018_g 0.0235078f $X=7.18 $Y=1.257
+ $X2=0 $Y2=0
cc_711 N_A_1243_48#_c_942_n N_A_1021_97#_M1018_g 0.00958924f $X=6.415 $Y=1.24
+ $X2=0 $Y2=0
cc_712 N_A_1243_48#_c_943_n N_A_1021_97#_M1018_g 0.00417413f $X=7.265 $Y=0.765
+ $X2=0 $Y2=0
cc_713 N_A_1243_48#_c_944_n N_A_1021_97#_M1018_g 0.00725494f $X=7.252 $Y=2.115
+ $X2=0 $Y2=0
cc_714 N_A_1243_48#_c_940_n N_A_1021_97#_c_1010_n 0.0351265f $X=6.43 $Y=2.33
+ $X2=0 $Y2=0
cc_715 N_A_1243_48#_c_947_n N_A_1021_97#_c_1010_n 0.0165372f $X=6.43 $Y=2.42
+ $X2=0 $Y2=0
cc_716 N_A_1243_48#_c_941_n N_A_1021_97#_c_1010_n 0.00219584f $X=7.18 $Y=1.257
+ $X2=0 $Y2=0
cc_717 N_A_1243_48#_c_948_n N_A_1021_97#_c_1010_n 0.00810163f $X=7.29 $Y=2.28
+ $X2=0 $Y2=0
cc_718 N_A_1243_48#_c_944_n N_A_1021_97#_c_1010_n 0.00835127f $X=7.252 $Y=2.115
+ $X2=0 $Y2=0
cc_719 N_A_1243_48#_M1014_g N_A_1021_97#_c_1011_n 4.90972e-19 $X=6.29 $Y=0.58
+ $X2=0 $Y2=0
cc_720 N_A_1243_48#_c_941_n N_A_1021_97#_c_1011_n 8.05791e-19 $X=7.18 $Y=1.257
+ $X2=0 $Y2=0
cc_721 N_A_1243_48#_c_940_n N_A_1021_97#_c_1012_n 0.016971f $X=6.43 $Y=2.33
+ $X2=0 $Y2=0
cc_722 N_A_1243_48#_c_941_n N_A_1021_97#_c_1012_n 0.0357047f $X=7.18 $Y=1.257
+ $X2=0 $Y2=0
cc_723 N_A_1243_48#_c_942_n N_A_1021_97#_c_1012_n 0.00480266f $X=6.415 $Y=1.24
+ $X2=0 $Y2=0
cc_724 N_A_1243_48#_c_940_n N_A_1021_97#_c_1014_n 0.00141301f $X=6.43 $Y=2.33
+ $X2=0 $Y2=0
cc_725 N_A_1243_48#_c_941_n N_A_1021_97#_c_1014_n 0.0229799f $X=7.18 $Y=1.257
+ $X2=0 $Y2=0
cc_726 N_A_1243_48#_c_944_n N_A_1021_97#_c_1014_n 0.0274223f $X=7.252 $Y=2.115
+ $X2=0 $Y2=0
cc_727 N_A_1243_48#_c_947_n N_VPWR_c_1455_n 0.00259711f $X=6.43 $Y=2.42 $X2=0
+ $Y2=0
cc_728 N_A_1243_48#_c_947_n N_VPWR_c_1456_n 0.00408705f $X=6.43 $Y=2.42 $X2=0
+ $Y2=0
cc_729 N_A_1243_48#_c_947_n N_VPWR_c_1439_n 0.005315f $X=6.43 $Y=2.42 $X2=0
+ $Y2=0
cc_730 N_A_1243_48#_M1014_g N_VGND_c_1802_n 0.00774989f $X=6.29 $Y=0.58 $X2=0
+ $Y2=0
cc_731 N_A_1243_48#_M1014_g N_VGND_c_1813_n 0.00383152f $X=6.29 $Y=0.58 $X2=0
+ $Y2=0
cc_732 N_A_1243_48#_M1014_g N_VGND_c_1825_n 0.00374269f $X=6.29 $Y=0.58 $X2=0
+ $Y2=0
cc_733 N_A_1021_97#_c_1010_n N_VPWR_c_1455_n 0.0044203f $X=7.05 $Y=2.045 $X2=0
+ $Y2=0
cc_734 N_A_1021_97#_c_1017_n N_VPWR_c_1456_n 0.0132031f $X=5.7 $Y=2.705 $X2=0
+ $Y2=0
cc_735 N_A_1021_97#_c_1010_n N_VPWR_c_1460_n 0.00316125f $X=7.05 $Y=2.045 $X2=0
+ $Y2=0
cc_736 N_A_1021_97#_c_1010_n N_VPWR_c_1439_n 0.00399737f $X=7.05 $Y=2.045 $X2=0
+ $Y2=0
cc_737 N_A_1021_97#_c_1017_n N_VPWR_c_1439_n 0.0127229f $X=5.7 $Y=2.705 $X2=0
+ $Y2=0
cc_738 N_A_1021_97#_c_1017_n N_A_301_74#_c_1617_n 0.0336878f $X=5.7 $Y=2.705
+ $X2=0 $Y2=0
cc_739 N_A_1021_97#_M1018_g N_VGND_c_1802_n 0.00139143f $X=7.05 $Y=0.645 $X2=0
+ $Y2=0
cc_740 N_A_1021_97#_M1018_g N_VGND_c_1814_n 0.00278237f $X=7.05 $Y=0.645 $X2=0
+ $Y2=0
cc_741 N_A_1021_97#_M1018_g N_VGND_c_1825_n 0.00355939f $X=7.05 $Y=0.645 $X2=0
+ $Y2=0
cc_742 N_A_1711_48#_c_1095_n N_A_1511_74#_c_1256_n 0.0101627f $X=8.965 $Y=2.05
+ $X2=0 $Y2=0
cc_743 N_A_1711_48#_c_1108_n N_A_1511_74#_c_1256_n 0.00907266f $X=9.865 $Y=1.94
+ $X2=0 $Y2=0
cc_744 N_A_1711_48#_c_1111_n N_A_1511_74#_c_1266_n 0.0124837f $X=8.8 $Y=2.465
+ $X2=0 $Y2=0
cc_745 N_A_1711_48#_c_1095_n N_A_1511_74#_c_1266_n 0.0135738f $X=8.965 $Y=2.05
+ $X2=0 $Y2=0
cc_746 N_A_1711_48#_c_1118_n N_A_1511_74#_c_1266_n 0.0189022f $X=9.6 $Y=2.22
+ $X2=0 $Y2=0
cc_747 N_A_1711_48#_c_1119_n N_A_1511_74#_c_1266_n 0.0153364f $X=9.765 $Y=2.815
+ $X2=0 $Y2=0
cc_748 N_A_1711_48#_c_1108_n N_A_1511_74#_c_1266_n 0.0018588f $X=9.865 $Y=1.94
+ $X2=0 $Y2=0
cc_749 N_A_1711_48#_c_1121_n N_A_1511_74#_c_1266_n 0.00453858f $X=9.765 $Y=2.105
+ $X2=0 $Y2=0
cc_750 N_A_1711_48#_c_1093_n N_A_1511_74#_c_1257_n 0.00543249f $X=8.89 $Y=0.94
+ $X2=0 $Y2=0
cc_751 N_A_1711_48#_c_1094_n N_A_1511_74#_c_1257_n 0.00954595f $X=8.705 $Y=0.94
+ $X2=0 $Y2=0
cc_752 N_A_1711_48#_c_1095_n N_A_1511_74#_c_1257_n 3.99884e-19 $X=8.965 $Y=2.05
+ $X2=0 $Y2=0
cc_753 N_A_1711_48#_c_1111_n N_A_1511_74#_c_1269_n 0.00474408f $X=8.8 $Y=2.465
+ $X2=0 $Y2=0
cc_754 N_A_1711_48#_c_1095_n N_A_1511_74#_c_1269_n 0.00944756f $X=8.965 $Y=2.05
+ $X2=0 $Y2=0
cc_755 N_A_1711_48#_c_1118_n N_A_1511_74#_c_1269_n 0.0240911f $X=9.6 $Y=2.22
+ $X2=0 $Y2=0
cc_756 N_A_1711_48#_c_1095_n N_A_1511_74#_c_1258_n 0.0125868f $X=8.965 $Y=2.05
+ $X2=0 $Y2=0
cc_757 N_A_1711_48#_c_1095_n N_A_1511_74#_c_1259_n 0.00394677f $X=8.965 $Y=2.05
+ $X2=0 $Y2=0
cc_758 N_A_1711_48#_c_1092_n N_A_1511_74#_c_1260_n 0.00189006f $X=8.63 $Y=0.865
+ $X2=0 $Y2=0
cc_759 N_A_1711_48#_c_1118_n N_A_1511_74#_c_1272_n 0.0121329f $X=9.6 $Y=2.22
+ $X2=0 $Y2=0
cc_760 N_A_1711_48#_c_1093_n N_A_1511_74#_c_1261_n 0.0061338f $X=8.89 $Y=0.94
+ $X2=0 $Y2=0
cc_761 N_A_1711_48#_c_1095_n N_A_1511_74#_c_1261_n 0.00668193f $X=8.965 $Y=2.05
+ $X2=0 $Y2=0
cc_762 N_A_1711_48#_c_1095_n N_A_1511_74#_c_1262_n 0.00122141f $X=8.965 $Y=2.05
+ $X2=0 $Y2=0
cc_763 N_A_1711_48#_c_1096_n N_A_1511_74#_c_1262_n 2.34832e-19 $X=10.44 $Y=1.465
+ $X2=0 $Y2=0
cc_764 N_A_1711_48#_c_1118_n N_A_1511_74#_c_1262_n 0.00949851f $X=9.6 $Y=2.22
+ $X2=0 $Y2=0
cc_765 N_A_1711_48#_c_1107_n N_A_1511_74#_c_1262_n 0.0166503f $X=9.865 $Y=1.3
+ $X2=0 $Y2=0
cc_766 N_A_1711_48#_c_1109_n N_A_1511_74#_c_1262_n 0.0019473f $X=9.725 $Y=0.62
+ $X2=0 $Y2=0
cc_767 N_A_1711_48#_c_1121_n N_A_1511_74#_c_1262_n 3.79292e-19 $X=9.765 $Y=2.105
+ $X2=0 $Y2=0
cc_768 N_A_1711_48#_c_1110_n N_A_1511_74#_c_1262_n 0.0210827f $X=9.865 $Y=1.465
+ $X2=0 $Y2=0
cc_769 N_A_1711_48#_c_1095_n N_A_1511_74#_c_1263_n 0.016294f $X=8.965 $Y=2.05
+ $X2=0 $Y2=0
cc_770 N_A_1711_48#_c_1096_n N_A_1511_74#_c_1263_n 0.012283f $X=10.44 $Y=1.465
+ $X2=0 $Y2=0
cc_771 N_A_1711_48#_c_1118_n N_A_1511_74#_c_1263_n 8.42398e-19 $X=9.6 $Y=2.22
+ $X2=0 $Y2=0
cc_772 N_A_1711_48#_c_1107_n N_A_1511_74#_c_1263_n 0.00185629f $X=9.865 $Y=1.3
+ $X2=0 $Y2=0
cc_773 N_A_1711_48#_c_1110_n N_A_1511_74#_c_1263_n 0.00423969f $X=9.865 $Y=1.465
+ $X2=0 $Y2=0
cc_774 N_A_1711_48#_c_1093_n N_A_1511_74#_c_1264_n 0.011098f $X=8.89 $Y=0.94
+ $X2=0 $Y2=0
cc_775 N_A_1711_48#_c_1107_n N_A_1511_74#_c_1264_n 0.00674353f $X=9.865 $Y=1.3
+ $X2=0 $Y2=0
cc_776 N_A_1711_48#_c_1109_n N_A_1511_74#_c_1264_n 0.0145622f $X=9.725 $Y=0.62
+ $X2=0 $Y2=0
cc_777 N_A_1711_48#_c_1117_n N_A_2322_368#_c_1372_n 0.0157799f $X=11.97 $Y=1.765
+ $X2=0 $Y2=0
cc_778 N_A_1711_48#_M1021_g N_A_2322_368#_M1019_g 0.0127598f $X=11.99 $Y=0.81
+ $X2=0 $Y2=0
cc_779 N_A_1711_48#_M1037_g N_A_2322_368#_c_1368_n 0.00371293f $X=11 $Y=0.74
+ $X2=0 $Y2=0
cc_780 N_A_1711_48#_c_1102_n N_A_2322_368#_c_1368_n 0.00699854f $X=11.88
+ $Y=1.375 $X2=0 $Y2=0
cc_781 N_A_1711_48#_M1021_g N_A_2322_368#_c_1368_n 0.0129616f $X=11.99 $Y=0.81
+ $X2=0 $Y2=0
cc_782 N_A_1711_48#_c_1106_n N_A_2322_368#_c_1368_n 4.37334e-19 $X=11.972
+ $Y=1.375 $X2=0 $Y2=0
cc_783 N_A_1711_48#_c_1100_n N_A_2322_368#_c_1374_n 0.00190857f $X=10.98
+ $Y=1.675 $X2=0 $Y2=0
cc_784 N_A_1711_48#_c_1115_n N_A_2322_368#_c_1374_n 0.00266445f $X=10.98
+ $Y=1.765 $X2=0 $Y2=0
cc_785 N_A_1711_48#_c_1103_n N_A_2322_368#_c_1374_n 9.29488e-19 $X=11.97
+ $Y=1.675 $X2=0 $Y2=0
cc_786 N_A_1711_48#_c_1117_n N_A_2322_368#_c_1374_n 0.0176452f $X=11.97 $Y=1.765
+ $X2=0 $Y2=0
cc_787 N_A_1711_48#_c_1103_n N_A_2322_368#_c_1369_n 0.0105363f $X=11.97 $Y=1.675
+ $X2=0 $Y2=0
cc_788 N_A_1711_48#_c_1106_n N_A_2322_368#_c_1369_n 0.00932161f $X=11.972
+ $Y=1.375 $X2=0 $Y2=0
cc_789 N_A_1711_48#_c_1100_n N_A_2322_368#_c_1370_n 0.00351192f $X=10.98
+ $Y=1.675 $X2=0 $Y2=0
cc_790 N_A_1711_48#_c_1102_n N_A_2322_368#_c_1370_n 0.0125974f $X=11.88 $Y=1.375
+ $X2=0 $Y2=0
cc_791 N_A_1711_48#_c_1103_n N_A_2322_368#_c_1370_n 0.00668695f $X=11.97
+ $Y=1.675 $X2=0 $Y2=0
cc_792 N_A_1711_48#_c_1106_n N_A_2322_368#_c_1370_n 7.34482e-19 $X=11.972
+ $Y=1.375 $X2=0 $Y2=0
cc_793 N_A_1711_48#_c_1103_n N_A_2322_368#_c_1371_n 0.0112528f $X=11.97 $Y=1.675
+ $X2=0 $Y2=0
cc_794 N_A_1711_48#_c_1106_n N_A_2322_368#_c_1371_n 0.00462619f $X=11.972
+ $Y=1.375 $X2=0 $Y2=0
cc_795 N_A_1711_48#_c_1118_n N_VPWR_M1029_d 0.00926404f $X=9.6 $Y=2.22 $X2=0
+ $Y2=0
cc_796 N_A_1711_48#_c_1111_n N_VPWR_c_1443_n 0.0204893f $X=8.8 $Y=2.465 $X2=0
+ $Y2=0
cc_797 N_A_1711_48#_c_1118_n N_VPWR_c_1443_n 0.0309547f $X=9.6 $Y=2.22 $X2=0
+ $Y2=0
cc_798 N_A_1711_48#_c_1119_n N_VPWR_c_1443_n 0.0133529f $X=9.765 $Y=2.815 $X2=0
+ $Y2=0
cc_799 N_A_1711_48#_c_1096_n N_VPWR_c_1444_n 0.00571957f $X=10.44 $Y=1.465 $X2=0
+ $Y2=0
cc_800 N_A_1711_48#_c_1097_n N_VPWR_c_1444_n 0.008783f $X=10.53 $Y=1.765 $X2=0
+ $Y2=0
cc_801 N_A_1711_48#_c_1119_n N_VPWR_c_1444_n 0.0454184f $X=9.765 $Y=2.815 $X2=0
+ $Y2=0
cc_802 N_A_1711_48#_c_1108_n N_VPWR_c_1444_n 0.00857316f $X=9.865 $Y=1.94 $X2=0
+ $Y2=0
cc_803 N_A_1711_48#_c_1194_p N_VPWR_c_1444_n 0.0192372f $X=10.445 $Y=1.465 $X2=0
+ $Y2=0
cc_804 N_A_1711_48#_c_1121_n N_VPWR_c_1444_n 0.0347849f $X=9.765 $Y=2.105 $X2=0
+ $Y2=0
cc_805 N_A_1711_48#_c_1097_n N_VPWR_c_1445_n 2.86313e-19 $X=10.53 $Y=1.765 $X2=0
+ $Y2=0
cc_806 N_A_1711_48#_c_1115_n N_VPWR_c_1445_n 0.00286015f $X=10.98 $Y=1.765 $X2=0
+ $Y2=0
cc_807 N_A_1711_48#_c_1097_n N_VPWR_c_1446_n 3.36435e-19 $X=10.53 $Y=1.765 $X2=0
+ $Y2=0
cc_808 N_A_1711_48#_c_1115_n N_VPWR_c_1446_n 0.0123087f $X=10.98 $Y=1.765 $X2=0
+ $Y2=0
cc_809 N_A_1711_48#_c_1117_n N_VPWR_c_1446_n 0.00281486f $X=11.97 $Y=1.765 $X2=0
+ $Y2=0
cc_810 N_A_1711_48#_c_1115_n N_VPWR_c_1447_n 0.00161121f $X=10.98 $Y=1.765 $X2=0
+ $Y2=0
cc_811 N_A_1711_48#_c_1102_n N_VPWR_c_1447_n 0.00697717f $X=11.88 $Y=1.375 $X2=0
+ $Y2=0
cc_812 N_A_1711_48#_c_1117_n N_VPWR_c_1447_n 0.00174105f $X=11.97 $Y=1.765 $X2=0
+ $Y2=0
cc_813 N_A_1711_48#_c_1117_n N_VPWR_c_1448_n 0.012056f $X=11.97 $Y=1.765 $X2=0
+ $Y2=0
cc_814 N_A_1711_48#_c_1119_n N_VPWR_c_1457_n 0.0154862f $X=9.765 $Y=2.815 $X2=0
+ $Y2=0
cc_815 N_A_1711_48#_c_1111_n N_VPWR_c_1460_n 0.00413917f $X=8.8 $Y=2.465 $X2=0
+ $Y2=0
cc_816 N_A_1711_48#_c_1097_n N_VPWR_c_1461_n 0.00445602f $X=10.53 $Y=1.765 $X2=0
+ $Y2=0
cc_817 N_A_1711_48#_c_1115_n N_VPWR_c_1461_n 0.00413917f $X=10.98 $Y=1.765 $X2=0
+ $Y2=0
cc_818 N_A_1711_48#_c_1117_n N_VPWR_c_1462_n 0.00481995f $X=11.97 $Y=1.765 $X2=0
+ $Y2=0
cc_819 N_A_1711_48#_c_1111_n N_VPWR_c_1439_n 0.00852225f $X=8.8 $Y=2.465 $X2=0
+ $Y2=0
cc_820 N_A_1711_48#_c_1097_n N_VPWR_c_1439_n 0.00862391f $X=10.53 $Y=1.765 $X2=0
+ $Y2=0
cc_821 N_A_1711_48#_c_1115_n N_VPWR_c_1439_n 0.00817726f $X=10.98 $Y=1.765 $X2=0
+ $Y2=0
cc_822 N_A_1711_48#_c_1117_n N_VPWR_c_1439_n 0.00508379f $X=11.97 $Y=1.765 $X2=0
+ $Y2=0
cc_823 N_A_1711_48#_c_1119_n N_VPWR_c_1439_n 0.0127853f $X=9.765 $Y=2.815 $X2=0
+ $Y2=0
cc_824 N_A_1711_48#_c_1097_n N_Q_c_1734_n 0.0116539f $X=10.53 $Y=1.765 $X2=0
+ $Y2=0
cc_825 N_A_1711_48#_c_1115_n N_Q_c_1734_n 0.0039888f $X=10.98 $Y=1.765 $X2=0
+ $Y2=0
cc_826 N_A_1711_48#_c_1097_n N_Q_c_1731_n 0.00376613f $X=10.53 $Y=1.765 $X2=0
+ $Y2=0
cc_827 N_A_1711_48#_M1022_g N_Q_c_1731_n 0.002587f $X=10.57 $Y=0.74 $X2=0 $Y2=0
cc_828 N_A_1711_48#_c_1099_n N_Q_c_1731_n 0.00739816f $X=10.89 $Y=1.375 $X2=0
+ $Y2=0
cc_829 N_A_1711_48#_c_1100_n N_Q_c_1731_n 0.00678318f $X=10.98 $Y=1.675 $X2=0
+ $Y2=0
cc_830 N_A_1711_48#_c_1115_n N_Q_c_1731_n 0.00432314f $X=10.98 $Y=1.765 $X2=0
+ $Y2=0
cc_831 N_A_1711_48#_M1037_g N_Q_c_1731_n 0.00508906f $X=11 $Y=0.74 $X2=0 $Y2=0
cc_832 N_A_1711_48#_c_1105_n N_Q_c_1731_n 0.00502889f $X=10.982 $Y=1.375 $X2=0
+ $Y2=0
cc_833 N_A_1711_48#_c_1194_p N_Q_c_1731_n 0.0256544f $X=10.445 $Y=1.465 $X2=0
+ $Y2=0
cc_834 N_A_1711_48#_c_1097_n N_Q_c_1736_n 0.00432091f $X=10.53 $Y=1.765 $X2=0
+ $Y2=0
cc_835 N_A_1711_48#_c_1099_n N_Q_c_1736_n 0.00338114f $X=10.89 $Y=1.375 $X2=0
+ $Y2=0
cc_836 N_A_1711_48#_c_1115_n N_Q_c_1736_n 0.0049909f $X=10.98 $Y=1.765 $X2=0
+ $Y2=0
cc_837 N_A_1711_48#_c_1108_n N_Q_c_1736_n 5.50555e-19 $X=9.865 $Y=1.94 $X2=0
+ $Y2=0
cc_838 N_A_1711_48#_c_1194_p N_Q_c_1736_n 0.00153914f $X=10.445 $Y=1.465 $X2=0
+ $Y2=0
cc_839 N_A_1711_48#_M1022_g Q 0.00772833f $X=10.57 $Y=0.74 $X2=0 $Y2=0
cc_840 N_A_1711_48#_M1037_g Q 0.00788704f $X=11 $Y=0.74 $X2=0 $Y2=0
cc_841 N_A_1711_48#_M1022_g Q 0.00260726f $X=10.57 $Y=0.74 $X2=0 $Y2=0
cc_842 N_A_1711_48#_c_1099_n Q 0.00120743f $X=10.89 $Y=1.375 $X2=0 $Y2=0
cc_843 N_A_1711_48#_M1037_g Q 0.00202916f $X=11 $Y=0.74 $X2=0 $Y2=0
cc_844 N_A_1711_48#_c_1096_n N_VGND_c_1803_n 0.00763556f $X=10.44 $Y=1.465 $X2=0
+ $Y2=0
cc_845 N_A_1711_48#_M1022_g N_VGND_c_1803_n 0.0198727f $X=10.57 $Y=0.74 $X2=0
+ $Y2=0
cc_846 N_A_1711_48#_c_1194_p N_VGND_c_1803_n 0.0276236f $X=10.445 $Y=1.465 $X2=0
+ $Y2=0
cc_847 N_A_1711_48#_c_1109_n N_VGND_c_1803_n 0.0645059f $X=9.725 $Y=0.62 $X2=0
+ $Y2=0
cc_848 N_A_1711_48#_M1037_g N_VGND_c_1804_n 0.00647412f $X=11 $Y=0.74 $X2=0
+ $Y2=0
cc_849 N_A_1711_48#_c_1102_n N_VGND_c_1804_n 0.00879713f $X=11.88 $Y=1.375 $X2=0
+ $Y2=0
cc_850 N_A_1711_48#_M1021_g N_VGND_c_1804_n 0.00408841f $X=11.99 $Y=0.81 $X2=0
+ $Y2=0
cc_851 N_A_1711_48#_M1021_g N_VGND_c_1805_n 0.0053693f $X=11.99 $Y=0.81 $X2=0
+ $Y2=0
cc_852 N_A_1711_48#_c_1092_n N_VGND_c_1814_n 0.00384553f $X=8.63 $Y=0.865 $X2=0
+ $Y2=0
cc_853 N_A_1711_48#_c_1109_n N_VGND_c_1815_n 0.0170752f $X=9.725 $Y=0.62 $X2=0
+ $Y2=0
cc_854 N_A_1711_48#_M1022_g N_VGND_c_1816_n 0.00434272f $X=10.57 $Y=0.74 $X2=0
+ $Y2=0
cc_855 N_A_1711_48#_M1037_g N_VGND_c_1816_n 0.00434272f $X=11 $Y=0.74 $X2=0
+ $Y2=0
cc_856 N_A_1711_48#_M1021_g N_VGND_c_1817_n 0.0047467f $X=11.99 $Y=0.81 $X2=0
+ $Y2=0
cc_857 N_A_1711_48#_c_1092_n N_VGND_c_1821_n 0.0120622f $X=8.63 $Y=0.865 $X2=0
+ $Y2=0
cc_858 N_A_1711_48#_c_1093_n N_VGND_c_1821_n 0.00784852f $X=8.89 $Y=0.94 $X2=0
+ $Y2=0
cc_859 N_A_1711_48#_c_1109_n N_VGND_c_1821_n 0.0149377f $X=9.725 $Y=0.62 $X2=0
+ $Y2=0
cc_860 N_A_1711_48#_c_1092_n N_VGND_c_1825_n 0.0075725f $X=8.63 $Y=0.865 $X2=0
+ $Y2=0
cc_861 N_A_1711_48#_M1022_g N_VGND_c_1825_n 0.00825059f $X=10.57 $Y=0.74 $X2=0
+ $Y2=0
cc_862 N_A_1711_48#_M1037_g N_VGND_c_1825_n 0.00825283f $X=11 $Y=0.74 $X2=0
+ $Y2=0
cc_863 N_A_1711_48#_M1021_g N_VGND_c_1825_n 0.00508379f $X=11.99 $Y=0.81 $X2=0
+ $Y2=0
cc_864 N_A_1711_48#_c_1109_n N_VGND_c_1825_n 0.0141497f $X=9.725 $Y=0.62 $X2=0
+ $Y2=0
cc_865 N_A_1511_74#_c_1266_n N_VPWR_c_1443_n 0.0065215f $X=9.54 $Y=1.885 $X2=0
+ $Y2=0
cc_866 N_A_1511_74#_c_1268_n N_VPWR_c_1443_n 0.00953279f $X=8.07 $Y=2.815 $X2=0
+ $Y2=0
cc_867 N_A_1511_74#_c_1266_n N_VPWR_c_1444_n 0.00419871f $X=9.54 $Y=1.885 $X2=0
+ $Y2=0
cc_868 N_A_1511_74#_c_1266_n N_VPWR_c_1457_n 0.00445602f $X=9.54 $Y=1.885 $X2=0
+ $Y2=0
cc_869 N_A_1511_74#_c_1268_n N_VPWR_c_1460_n 0.0145938f $X=8.07 $Y=2.815 $X2=0
+ $Y2=0
cc_870 N_A_1511_74#_c_1266_n N_VPWR_c_1439_n 0.00863833f $X=9.54 $Y=1.885 $X2=0
+ $Y2=0
cc_871 N_A_1511_74#_c_1268_n N_VPWR_c_1439_n 0.0120466f $X=8.07 $Y=2.815 $X2=0
+ $Y2=0
cc_872 N_A_1511_74#_c_1259_n N_VGND_M1009_d 0.00152837f $X=9.28 $Y=1.14 $X2=0
+ $Y2=0
cc_873 N_A_1511_74#_c_1262_n N_VGND_M1009_d 0.00160992f $X=9.445 $Y=1.14 $X2=0
+ $Y2=0
cc_874 N_A_1511_74#_c_1264_n N_VGND_c_1803_n 0.00375193f $X=9.455 $Y=1.22 $X2=0
+ $Y2=0
cc_875 N_A_1511_74#_c_1260_n N_VGND_c_1814_n 0.0144717f $X=8.025 $Y=0.58 $X2=0
+ $Y2=0
cc_876 N_A_1511_74#_c_1264_n N_VGND_c_1815_n 0.00434272f $X=9.455 $Y=1.22 $X2=0
+ $Y2=0
cc_877 N_A_1511_74#_c_1257_n N_VGND_c_1821_n 0.0106389f $X=8.85 $Y=0.97 $X2=0
+ $Y2=0
cc_878 N_A_1511_74#_c_1259_n N_VGND_c_1821_n 0.0128493f $X=9.28 $Y=1.14 $X2=0
+ $Y2=0
cc_879 N_A_1511_74#_c_1260_n N_VGND_c_1821_n 0.0123089f $X=8.025 $Y=0.58 $X2=0
+ $Y2=0
cc_880 N_A_1511_74#_c_1261_n N_VGND_c_1821_n 0.0146416f $X=8.935 $Y=0.97 $X2=0
+ $Y2=0
cc_881 N_A_1511_74#_c_1262_n N_VGND_c_1821_n 0.00511089f $X=9.445 $Y=1.14 $X2=0
+ $Y2=0
cc_882 N_A_1511_74#_c_1263_n N_VGND_c_1821_n 5.45988e-19 $X=9.445 $Y=1.385 $X2=0
+ $Y2=0
cc_883 N_A_1511_74#_c_1264_n N_VGND_c_1821_n 0.00557841f $X=9.455 $Y=1.22 $X2=0
+ $Y2=0
cc_884 N_A_1511_74#_c_1260_n N_VGND_c_1825_n 0.0119991f $X=8.025 $Y=0.58 $X2=0
+ $Y2=0
cc_885 N_A_1511_74#_c_1264_n N_VGND_c_1825_n 0.00830058f $X=9.455 $Y=1.22 $X2=0
+ $Y2=0
cc_886 N_A_2322_368#_c_1374_n N_VPWR_c_1447_n 0.0741374f $X=11.745 $Y=1.985
+ $X2=0 $Y2=0
cc_887 N_A_2322_368#_c_1372_n N_VPWR_c_1448_n 0.00772238f $X=12.495 $Y=1.765
+ $X2=0 $Y2=0
cc_888 N_A_2322_368#_c_1374_n N_VPWR_c_1448_n 0.0711612f $X=11.745 $Y=1.985
+ $X2=0 $Y2=0
cc_889 N_A_2322_368#_c_1369_n N_VPWR_c_1448_n 0.0219385f $X=12.57 $Y=1.485 $X2=0
+ $Y2=0
cc_890 N_A_2322_368#_c_1372_n N_VPWR_c_1450_n 5.28947e-19 $X=12.495 $Y=1.765
+ $X2=0 $Y2=0
cc_891 N_A_2322_368#_c_1373_n N_VPWR_c_1450_n 0.0117933f $X=12.945 $Y=1.765
+ $X2=0 $Y2=0
cc_892 N_A_2322_368#_c_1374_n N_VPWR_c_1462_n 0.0097982f $X=11.745 $Y=1.985
+ $X2=0 $Y2=0
cc_893 N_A_2322_368#_c_1372_n N_VPWR_c_1463_n 0.00445602f $X=12.495 $Y=1.765
+ $X2=0 $Y2=0
cc_894 N_A_2322_368#_c_1373_n N_VPWR_c_1463_n 0.00413917f $X=12.945 $Y=1.765
+ $X2=0 $Y2=0
cc_895 N_A_2322_368#_c_1372_n N_VPWR_c_1439_n 0.00862391f $X=12.495 $Y=1.765
+ $X2=0 $Y2=0
cc_896 N_A_2322_368#_c_1373_n N_VPWR_c_1439_n 0.00817726f $X=12.945 $Y=1.765
+ $X2=0 $Y2=0
cc_897 N_A_2322_368#_c_1374_n N_VPWR_c_1439_n 0.0111907f $X=11.745 $Y=1.985
+ $X2=0 $Y2=0
cc_898 N_A_2322_368#_c_1368_n N_Q_c_1731_n 0.00539511f $X=11.775 $Y=0.665 $X2=0
+ $Y2=0
cc_899 N_A_2322_368#_c_1374_n N_Q_c_1731_n 0.00488341f $X=11.745 $Y=1.985 $X2=0
+ $Y2=0
cc_900 N_A_2322_368#_c_1370_n N_Q_c_1731_n 0.00932649f $X=11.76 $Y=1.485 $X2=0
+ $Y2=0
cc_901 N_A_2322_368#_M1019_g N_Q_N_c_1770_n 0.00419288f $X=12.5 $Y=0.76 $X2=0
+ $Y2=0
cc_902 N_A_2322_368#_M1039_g N_Q_N_c_1770_n 0.0188457f $X=12.945 $Y=0.76 $X2=0
+ $Y2=0
cc_903 N_A_2322_368#_c_1369_n N_Q_N_c_1770_n 0.0142268f $X=12.57 $Y=1.485 $X2=0
+ $Y2=0
cc_904 N_A_2322_368#_c_1371_n N_Q_N_c_1770_n 0.0032855f $X=12.945 $Y=1.542 $X2=0
+ $Y2=0
cc_905 N_A_2322_368#_c_1372_n N_Q_N_c_1772_n 0.00943074f $X=12.495 $Y=1.765
+ $X2=0 $Y2=0
cc_906 N_A_2322_368#_c_1373_n N_Q_N_c_1772_n 3.88029e-19 $X=12.945 $Y=1.765
+ $X2=0 $Y2=0
cc_907 N_A_2322_368#_M1039_g Q_N 0.0068339f $X=12.945 $Y=0.76 $X2=0 $Y2=0
cc_908 N_A_2322_368#_c_1373_n Q_N 0.0022049f $X=12.945 $Y=1.765 $X2=0 $Y2=0
cc_909 N_A_2322_368#_c_1369_n Q_N 0.0159506f $X=12.57 $Y=1.485 $X2=0 $Y2=0
cc_910 N_A_2322_368#_c_1371_n Q_N 0.0156589f $X=12.945 $Y=1.542 $X2=0 $Y2=0
cc_911 N_A_2322_368#_c_1372_n Q_N 0.00386859f $X=12.495 $Y=1.765 $X2=0 $Y2=0
cc_912 N_A_2322_368#_c_1373_n Q_N 0.0223155f $X=12.945 $Y=1.765 $X2=0 $Y2=0
cc_913 N_A_2322_368#_c_1369_n Q_N 0.0141835f $X=12.57 $Y=1.485 $X2=0 $Y2=0
cc_914 N_A_2322_368#_c_1371_n Q_N 0.00899713f $X=12.945 $Y=1.542 $X2=0 $Y2=0
cc_915 N_A_2322_368#_c_1368_n N_VGND_c_1804_n 0.0417545f $X=11.775 $Y=0.665
+ $X2=0 $Y2=0
cc_916 N_A_2322_368#_M1019_g N_VGND_c_1805_n 0.00828604f $X=12.5 $Y=0.76 $X2=0
+ $Y2=0
cc_917 N_A_2322_368#_M1039_g N_VGND_c_1805_n 0.00139894f $X=12.945 $Y=0.76 $X2=0
+ $Y2=0
cc_918 N_A_2322_368#_M1019_g N_VGND_c_1806_n 4.25008e-19 $X=12.5 $Y=0.76 $X2=0
+ $Y2=0
cc_919 N_A_2322_368#_c_1368_n N_VGND_c_1806_n 0.0221622f $X=11.775 $Y=0.665
+ $X2=0 $Y2=0
cc_920 N_A_2322_368#_c_1369_n N_VGND_c_1806_n 0.0228231f $X=12.57 $Y=1.485 $X2=0
+ $Y2=0
cc_921 N_A_2322_368#_M1019_g N_VGND_c_1808_n 0.00139971f $X=12.5 $Y=0.76 $X2=0
+ $Y2=0
cc_922 N_A_2322_368#_M1039_g N_VGND_c_1808_n 0.0118008f $X=12.945 $Y=0.76 $X2=0
+ $Y2=0
cc_923 N_A_2322_368#_M1019_g N_VGND_c_1938_n 0.00359505f $X=12.5 $Y=0.76 $X2=0
+ $Y2=0
cc_924 N_A_2322_368#_c_1369_n N_VGND_c_1938_n 0.00137637f $X=12.57 $Y=1.485
+ $X2=0 $Y2=0
cc_925 N_A_2322_368#_c_1368_n N_VGND_c_1817_n 0.00757218f $X=11.775 $Y=0.665
+ $X2=0 $Y2=0
cc_926 N_A_2322_368#_M1019_g N_VGND_c_1818_n 0.00468165f $X=12.5 $Y=0.76 $X2=0
+ $Y2=0
cc_927 N_A_2322_368#_M1039_g N_VGND_c_1818_n 0.00468165f $X=12.945 $Y=0.76 $X2=0
+ $Y2=0
cc_928 N_A_2322_368#_M1019_g N_VGND_c_1825_n 0.00453141f $X=12.5 $Y=0.76 $X2=0
+ $Y2=0
cc_929 N_A_2322_368#_M1039_g N_VGND_c_1825_n 0.00453141f $X=12.945 $Y=0.76 $X2=0
+ $Y2=0
cc_930 N_A_2322_368#_c_1368_n N_VGND_c_1825_n 0.0114347f $X=11.775 $Y=0.665
+ $X2=0 $Y2=0
cc_931 N_VPWR_M1027_d N_A_301_74#_c_1619_n 0.0117101f $X=2.6 $Y=2.265 $X2=0
+ $Y2=0
cc_932 N_VPWR_c_1441_n N_A_301_74#_c_1619_n 0.020145f $X=2.88 $Y=2.875 $X2=0
+ $Y2=0
cc_933 N_VPWR_c_1439_n N_A_301_74#_c_1619_n 0.024843f $X=13.2 $Y=3.33 $X2=0
+ $Y2=0
cc_934 N_VPWR_M1027_d N_A_301_74#_c_1608_n 0.0144814f $X=2.6 $Y=2.265 $X2=0
+ $Y2=0
cc_935 N_VPWR_M1027_d N_A_301_74#_c_1613_n 4.01762e-19 $X=2.6 $Y=2.265 $X2=0
+ $Y2=0
cc_936 N_VPWR_M1031_s N_A_301_74#_c_1613_n 0.0056789f $X=4.095 $Y=1.84 $X2=0
+ $Y2=0
cc_937 N_VPWR_c_1442_n N_A_301_74#_c_1613_n 0.0150387f $X=4.24 $Y=2.805 $X2=0
+ $Y2=0
cc_938 N_VPWR_c_1439_n N_A_301_74#_c_1613_n 0.0349768f $X=13.2 $Y=3.33 $X2=0
+ $Y2=0
cc_939 N_VPWR_M1031_s N_A_301_74#_c_1614_n 0.010278f $X=4.095 $Y=1.84 $X2=0
+ $Y2=0
cc_940 N_VPWR_c_1456_n N_A_301_74#_c_1615_n 0.00574705f $X=6.575 $Y=3.33 $X2=0
+ $Y2=0
cc_941 N_VPWR_c_1439_n N_A_301_74#_c_1615_n 0.00948569f $X=13.2 $Y=3.33 $X2=0
+ $Y2=0
cc_942 N_VPWR_M1031_s N_A_301_74#_c_1665_n 7.28257e-19 $X=4.095 $Y=1.84 $X2=0
+ $Y2=0
cc_943 N_VPWR_c_1442_n N_A_301_74#_c_1665_n 0.00703764f $X=4.24 $Y=2.805 $X2=0
+ $Y2=0
cc_944 N_VPWR_c_1456_n N_A_301_74#_c_1665_n 0.00272086f $X=6.575 $Y=3.33 $X2=0
+ $Y2=0
cc_945 N_VPWR_c_1439_n N_A_301_74#_c_1665_n 0.0107375f $X=13.2 $Y=3.33 $X2=0
+ $Y2=0
cc_946 N_VPWR_c_1440_n N_A_301_74#_c_1616_n 0.00545176f $X=0.89 $Y=2.41 $X2=0
+ $Y2=0
cc_947 N_VPWR_c_1453_n N_A_301_74#_c_1616_n 0.0118538f $X=2.67 $Y=3.33 $X2=0
+ $Y2=0
cc_948 N_VPWR_c_1439_n N_A_301_74#_c_1616_n 0.0116474f $X=13.2 $Y=3.33 $X2=0
+ $Y2=0
cc_949 N_VPWR_M1027_d N_A_301_74#_c_1714_n 0.00240288f $X=2.6 $Y=2.265 $X2=0
+ $Y2=0
cc_950 N_VPWR_c_1441_n N_A_301_74#_c_1714_n 0.0143529f $X=2.88 $Y=2.875 $X2=0
+ $Y2=0
cc_951 N_VPWR_c_1439_n N_A_301_74#_c_1714_n 8.67729e-19 $X=13.2 $Y=3.33 $X2=0
+ $Y2=0
cc_952 N_VPWR_c_1456_n N_A_301_74#_c_1617_n 0.00908144f $X=6.575 $Y=3.33 $X2=0
+ $Y2=0
cc_953 N_VPWR_c_1439_n N_A_301_74#_c_1617_n 0.00876884f $X=13.2 $Y=3.33 $X2=0
+ $Y2=0
cc_954 N_VPWR_c_1445_n N_Q_c_1734_n 0.0563195f $X=11.205 $Y=2.305 $X2=0 $Y2=0
cc_955 N_VPWR_c_1447_n N_Q_c_1734_n 0.00900415f $X=11.205 $Y=1.985 $X2=0 $Y2=0
cc_956 N_VPWR_c_1461_n N_Q_c_1734_n 0.0110241f $X=11.04 $Y=3.33 $X2=0 $Y2=0
cc_957 N_VPWR_c_1439_n N_Q_c_1734_n 0.00909194f $X=13.2 $Y=3.33 $X2=0 $Y2=0
cc_958 N_VPWR_c_1444_n N_Q_c_1736_n 0.076487f $X=10.305 $Y=1.985 $X2=0 $Y2=0
cc_959 N_VPWR_c_1447_n N_Q_c_1736_n 0.0115032f $X=11.205 $Y=1.985 $X2=0 $Y2=0
cc_960 N_VPWR_c_1448_n N_Q_N_c_1772_n 0.0550023f $X=12.27 $Y=1.985 $X2=0 $Y2=0
cc_961 N_VPWR_c_1450_n N_Q_N_c_1772_n 0.0255358f $X=13.17 $Y=2.405 $X2=0 $Y2=0
cc_962 N_VPWR_c_1463_n N_Q_N_c_1772_n 0.0123628f $X=13.005 $Y=3.33 $X2=0 $Y2=0
cc_963 N_VPWR_c_1439_n N_Q_N_c_1772_n 0.0101999f $X=13.2 $Y=3.33 $X2=0 $Y2=0
cc_964 N_VPWR_M1034_d Q_N 0.00426951f $X=13.02 $Y=1.84 $X2=0 $Y2=0
cc_965 N_VPWR_c_1448_n Q_N 0.0233786f $X=12.27 $Y=1.985 $X2=0 $Y2=0
cc_966 N_VPWR_c_1450_n Q_N 0.0213356f $X=13.17 $Y=2.405 $X2=0 $Y2=0
cc_967 N_A_301_74#_c_1619_n A_423_453# 0.012064f $X=2.925 $Y=2.455 $X2=-0.19
+ $Y2=-0.245
cc_968 N_A_301_74#_c_1618_n N_VGND_c_1799_n 0.00833256f $X=2.245 $Y=0.515 $X2=0
+ $Y2=0
cc_969 N_A_301_74#_c_1605_n N_VGND_c_1800_n 0.0223267f $X=2.33 $Y=1.35 $X2=0
+ $Y2=0
cc_970 N_A_301_74#_c_1606_n N_VGND_c_1800_n 0.0175851f $X=2.925 $Y=1.435 $X2=0
+ $Y2=0
cc_971 N_A_301_74#_c_1618_n N_VGND_c_1809_n 0.029956f $X=2.245 $Y=0.515 $X2=0
+ $Y2=0
cc_972 N_A_301_74#_c_1618_n N_VGND_c_1825_n 0.0318853f $X=2.245 $Y=0.515 $X2=0
+ $Y2=0
cc_973 N_A_301_74#_c_1618_n A_450_74# 0.00397798f $X=2.245 $Y=0.515 $X2=-0.19
+ $Y2=-0.245
cc_974 N_A_301_74#_c_1605_n A_450_74# 0.00148509f $X=2.33 $Y=1.35 $X2=-0.19
+ $Y2=-0.245
cc_975 Q N_VGND_c_1803_n 0.0308109f $X=10.715 $Y=0.47 $X2=0 $Y2=0
cc_976 Q N_VGND_c_1804_n 0.0293763f $X=10.715 $Y=0.47 $X2=0 $Y2=0
cc_977 Q N_VGND_c_1816_n 0.0144922f $X=10.715 $Y=0.47 $X2=0 $Y2=0
cc_978 Q N_VGND_c_1825_n 0.0118826f $X=10.715 $Y=0.47 $X2=0 $Y2=0
cc_979 N_Q_N_c_1770_n N_VGND_M1039_s 0.00302692f $X=13.075 $Y=1.025 $X2=0 $Y2=0
cc_980 N_Q_N_c_1770_n N_VGND_c_1806_n 0.0111722f $X=13.075 $Y=1.025 $X2=0 $Y2=0
cc_981 N_Q_N_c_1770_n N_VGND_c_1808_n 0.0234536f $X=13.075 $Y=1.025 $X2=0 $Y2=0
