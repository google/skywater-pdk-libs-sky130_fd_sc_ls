* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__fa_2 A B CIN VGND VNB VPB VPWR COUT SUM
X0 VPWR A a_683_347# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 VGND a_992_347# SUM VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X2 a_1205_79# A VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X3 SUM a_992_347# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X4 VPWR CIN a_683_347# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 VGND a_336_347# COUT VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X6 a_701_79# a_336_347# a_992_347# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X7 COUT a_336_347# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X8 a_27_378# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 a_683_347# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 VPWR B a_27_378# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 a_27_79# A VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X12 a_27_79# CIN a_336_347# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X13 VPWR a_992_347# SUM VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X14 a_992_347# CIN a_1119_79# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X15 a_1119_79# B a_1205_79# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X16 a_1202_368# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X17 a_683_347# a_336_347# a_992_347# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X18 VGND B a_27_79# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X19 a_992_347# CIN a_1094_347# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X20 a_484_347# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X21 a_487_79# A VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X22 a_1094_347# B a_1202_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X23 COUT a_336_347# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X24 VGND CIN a_701_79# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X25 a_27_378# CIN a_336_347# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X26 a_336_347# B a_484_347# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X27 SUM a_992_347# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X28 VGND A a_701_79# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X29 VPWR a_336_347# COUT VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X30 a_336_347# B a_487_79# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X31 a_701_79# B VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
.ends
