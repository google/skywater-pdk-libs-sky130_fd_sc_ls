* File: sky130_fd_sc_ls__dlrtn_1.pxi.spice
* Created: Wed Sep  2 11:03:38 2020
* 
x_PM_SKY130_FD_SC_LS__DLRTN_1%D N_D_M1012_g N_D_c_126_n N_D_M1000_g D
+ PM_SKY130_FD_SC_LS__DLRTN_1%D
x_PM_SKY130_FD_SC_LS__DLRTN_1%GATE_N N_GATE_N_M1001_g N_GATE_N_c_152_n
+ N_GATE_N_M1019_g GATE_N PM_SKY130_FD_SC_LS__DLRTN_1%GATE_N
x_PM_SKY130_FD_SC_LS__DLRTN_1%A_232_98# N_A_232_98#_M1001_d N_A_232_98#_M1019_d
+ N_A_232_98#_c_185_n N_A_232_98#_M1009_g N_A_232_98#_M1015_g
+ N_A_232_98#_M1017_g N_A_232_98#_c_193_n N_A_232_98#_c_194_n
+ N_A_232_98#_M1003_g N_A_232_98#_c_188_n N_A_232_98#_c_196_n
+ N_A_232_98#_c_189_n N_A_232_98#_c_197_n N_A_232_98#_c_190_n
+ N_A_232_98#_c_199_n N_A_232_98#_c_200_n N_A_232_98#_c_201_n
+ N_A_232_98#_c_202_n N_A_232_98#_c_203_n PM_SKY130_FD_SC_LS__DLRTN_1%A_232_98#
x_PM_SKY130_FD_SC_LS__DLRTN_1%A_27_136# N_A_27_136#_M1012_s N_A_27_136#_M1000_s
+ N_A_27_136#_c_308_n N_A_27_136#_c_309_n N_A_27_136#_c_319_n
+ N_A_27_136#_M1005_g N_A_27_136#_c_310_n N_A_27_136#_c_311_n
+ N_A_27_136#_M1011_g N_A_27_136#_c_312_n N_A_27_136#_c_313_n
+ N_A_27_136#_c_314_n N_A_27_136#_c_315_n N_A_27_136#_c_316_n
+ N_A_27_136#_c_320_n N_A_27_136#_c_317_n PM_SKY130_FD_SC_LS__DLRTN_1%A_27_136#
x_PM_SKY130_FD_SC_LS__DLRTN_1%A_357_392# N_A_357_392#_M1015_s
+ N_A_357_392#_M1009_s N_A_357_392#_c_389_n N_A_357_392#_M1002_g
+ N_A_357_392#_M1007_g N_A_357_392#_c_391_n N_A_357_392#_c_397_n
+ N_A_357_392#_c_398_n N_A_357_392#_c_392_n N_A_357_392#_c_393_n
+ N_A_357_392#_c_394_n N_A_357_392#_c_395_n N_A_357_392#_c_399_n
+ PM_SKY130_FD_SC_LS__DLRTN_1%A_357_392#
x_PM_SKY130_FD_SC_LS__DLRTN_1%A_897_406# N_A_897_406#_M1013_s
+ N_A_897_406#_M1010_d N_A_897_406#_c_492_n N_A_897_406#_M1018_g
+ N_A_897_406#_M1004_g N_A_897_406#_c_484_n N_A_897_406#_M1014_g
+ N_A_897_406#_c_486_n N_A_897_406#_M1006_g N_A_897_406#_c_487_n
+ N_A_897_406#_c_495_n N_A_897_406#_c_488_n N_A_897_406#_c_496_n
+ N_A_897_406#_c_489_n N_A_897_406#_c_497_n N_A_897_406#_c_490_n
+ N_A_897_406#_c_499_n N_A_897_406#_c_491_n
+ PM_SKY130_FD_SC_LS__DLRTN_1%A_897_406#
x_PM_SKY130_FD_SC_LS__DLRTN_1%A_654_392# N_A_654_392#_M1017_d
+ N_A_654_392#_M1002_d N_A_654_392#_c_595_n N_A_654_392#_c_596_n
+ N_A_654_392#_c_605_n N_A_654_392#_M1010_g N_A_654_392#_c_597_n
+ N_A_654_392#_M1013_g N_A_654_392#_c_598_n N_A_654_392#_c_607_n
+ N_A_654_392#_c_608_n N_A_654_392#_c_609_n N_A_654_392#_c_610_n
+ N_A_654_392#_c_599_n N_A_654_392#_c_600_n N_A_654_392#_c_601_n
+ N_A_654_392#_c_602_n N_A_654_392#_c_603_n N_A_654_392#_c_604_n
+ PM_SKY130_FD_SC_LS__DLRTN_1%A_654_392#
x_PM_SKY130_FD_SC_LS__DLRTN_1%RESET_B N_RESET_B_c_702_n N_RESET_B_M1008_g
+ N_RESET_B_c_703_n N_RESET_B_M1016_g RESET_B
+ PM_SKY130_FD_SC_LS__DLRTN_1%RESET_B
x_PM_SKY130_FD_SC_LS__DLRTN_1%VPWR N_VPWR_M1000_d N_VPWR_M1009_d N_VPWR_M1018_d
+ N_VPWR_M1016_d N_VPWR_c_737_n N_VPWR_c_738_n N_VPWR_c_739_n N_VPWR_c_740_n
+ N_VPWR_c_741_n VPWR N_VPWR_c_742_n N_VPWR_c_743_n N_VPWR_c_744_n
+ N_VPWR_c_736_n N_VPWR_c_746_n N_VPWR_c_747_n N_VPWR_c_748_n
+ PM_SKY130_FD_SC_LS__DLRTN_1%VPWR
x_PM_SKY130_FD_SC_LS__DLRTN_1%Q N_Q_M1014_d N_Q_M1006_d N_Q_c_810_n N_Q_c_811_n
+ Q Q Q Q N_Q_c_812_n PM_SKY130_FD_SC_LS__DLRTN_1%Q
x_PM_SKY130_FD_SC_LS__DLRTN_1%VGND N_VGND_M1012_d N_VGND_M1015_d N_VGND_M1004_d
+ N_VGND_M1008_d N_VGND_c_832_n N_VGND_c_833_n N_VGND_c_834_n N_VGND_c_835_n
+ N_VGND_c_836_n N_VGND_c_837_n VGND N_VGND_c_838_n N_VGND_c_839_n
+ N_VGND_c_840_n N_VGND_c_841_n N_VGND_c_842_n N_VGND_c_843_n
+ PM_SKY130_FD_SC_LS__DLRTN_1%VGND
cc_1 VNB N_D_M1012_g 0.028833f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.955
cc_2 VNB N_D_c_126_n 0.0252084f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.895
cc_3 VNB D 0.00388042f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_4 VNB N_GATE_N_M1001_g 0.0314648f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.955
cc_5 VNB N_GATE_N_c_152_n 0.0197831f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.895
cc_6 VNB GATE_N 0.0017082f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_7 VNB N_A_232_98#_c_185_n 0.0174347f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.39
cc_8 VNB N_A_232_98#_M1015_g 0.027213f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.615
cc_9 VNB N_A_232_98#_M1017_g 0.049147f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_232_98#_c_188_n 0.0342904f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_232_98#_c_189_n 0.00893275f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_232_98#_c_190_n 0.0134414f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_136#_c_308_n 0.0447037f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.39
cc_14 VNB N_A_27_136#_c_309_n 0.00414301f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_15 VNB N_A_27_136#_c_310_n 0.033783f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.615
cc_16 VNB N_A_27_136#_c_311_n 0.0166671f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_27_136#_c_312_n 0.0125907f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_27_136#_c_313_n 0.0131232f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_27_136#_c_314_n 0.0115633f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_27_136#_c_315_n 0.00337621f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_27_136#_c_316_n 0.0132007f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_27_136#_c_317_n 0.0193493f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_357_392#_c_389_n 0.0173696f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.39
cc_24 VNB N_A_357_392#_M1007_g 0.0319639f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.615
cc_25 VNB N_A_357_392#_c_391_n 0.00242021f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.615
cc_26 VNB N_A_357_392#_c_392_n 0.00190671f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_357_392#_c_393_n 0.0194901f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_357_392#_c_394_n 0.0312515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_357_392#_c_395_n 0.0043822f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_897_406#_M1004_g 0.0440734f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.615
cc_31 VNB N_A_897_406#_c_484_n 0.0127126f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.615
cc_32 VNB N_A_897_406#_M1014_g 0.0298216f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_897_406#_c_486_n 0.0339664f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_897_406#_c_487_n 0.00957668f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_897_406#_c_488_n 0.00892155f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_897_406#_c_489_n 0.0037106f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_897_406#_c_490_n 0.00551864f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_897_406#_c_491_n 0.00881731f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_654_392#_c_595_n 0.0220846f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.39
cc_40 VNB N_A_654_392#_c_596_n 0.020671f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_41 VNB N_A_654_392#_c_597_n 0.0176306f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.615
cc_42 VNB N_A_654_392#_c_598_n 0.0121055f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_654_392#_c_599_n 0.0028741f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_654_392#_c_600_n 0.0176552f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_654_392#_c_601_n 0.00257655f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_654_392#_c_602_n 0.00398174f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_654_392#_c_603_n 0.00400951f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_654_392#_c_604_n 0.0123765f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_RESET_B_c_702_n 0.0183781f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.45
cc_50 VNB N_RESET_B_c_703_n 0.0405077f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB RESET_B 0.0101043f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.39
cc_52 VNB N_VPWR_c_736_n 0.302998f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_Q_c_810_n 0.0275421f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_Q_c_811_n 0.0151501f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.615
cc_55 VNB N_Q_c_812_n 0.0251008f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_832_n 0.00999694f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.615
cc_57 VNB N_VGND_c_833_n 0.00984624f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_834_n 0.0439944f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_835_n 0.00635026f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_836_n 0.0328251f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_837_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_838_n 0.0194325f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_839_n 0.0223814f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_840_n 0.416002f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_841_n 0.023189f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_842_n 0.0375862f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_843_n 0.0279221f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VPB N_D_c_126_n 0.0442086f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.895
cc_69 VPB D 0.00137322f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_70 VPB N_GATE_N_c_152_n 0.0425388f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.895
cc_71 VPB GATE_N 0.00232335f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_72 VPB N_A_232_98#_c_185_n 0.0361213f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=2.39
cc_73 VPB N_A_232_98#_M1017_g 0.00462336f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_A_232_98#_c_193_n 0.0105215f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_A_232_98#_c_194_n 0.0710897f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_A_232_98#_c_188_n 0.0139115f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_A_232_98#_c_196_n 0.0198893f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_A_232_98#_c_197_n 0.00545165f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 VPB N_A_232_98#_c_190_n 0.0069577f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 VPB N_A_232_98#_c_199_n 0.00837753f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_A_232_98#_c_200_n 0.00911126f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 VPB N_A_232_98#_c_201_n 0.00402733f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 VPB N_A_232_98#_c_202_n 0.0110241f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_84 VPB N_A_232_98#_c_203_n 0.00530584f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_A_27_136#_c_309_n 0.00806868f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_86 VPB N_A_27_136#_c_319_n 0.0217632f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_A_27_136#_c_320_n 0.0448422f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_A_27_136#_c_317_n 0.0137996f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_A_357_392#_c_389_n 0.0350524f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=2.39
cc_90 VPB N_A_357_392#_c_397_n 0.0138632f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB N_A_357_392#_c_398_n 0.00108801f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_92 VPB N_A_357_392#_c_399_n 0.00288783f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_A_897_406#_c_492_n 0.0623617f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=2.39
cc_94 VPB N_A_897_406#_c_484_n 0.0258438f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.615
cc_95 VPB N_A_897_406#_c_486_n 0.029474f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB N_A_897_406#_c_495_n 0.010104f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_A_897_406#_c_496_n 0.00698864f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_A_897_406#_c_497_n 0.00968685f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB N_A_897_406#_c_490_n 6.80603e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 VPB N_A_897_406#_c_499_n 0.00393712f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB N_A_897_406#_c_491_n 0.00211738f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_102 VPB N_A_654_392#_c_605_n 0.0180852f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 VPB N_A_654_392#_c_598_n 0.0214382f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB N_A_654_392#_c_607_n 0.00358759f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_105 VPB N_A_654_392#_c_608_n 0.00569705f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_A_654_392#_c_609_n 0.0233987f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB N_A_654_392#_c_610_n 0.00173401f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_A_654_392#_c_603_n 0.00311577f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_109 VPB N_RESET_B_c_703_n 0.0239354f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_110 VPB N_VPWR_c_737_n 0.0303098f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_VPWR_c_738_n 0.0140923f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_739_n 0.0142191f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_VPWR_c_740_n 0.0362164f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_VPWR_c_741_n 0.00631473f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_VPWR_c_742_n 0.0565095f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_VPWR_c_743_n 0.0241717f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_744_n 0.0189171f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_736_n 0.11316f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_746_n 0.0272551f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_747_n 0.0344519f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_748_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB Q 0.0138432f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB Q 0.041687f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_Q_c_812_n 0.0075608f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 N_D_M1012_g N_GATE_N_M1001_g 0.0243459f $X=0.495 $Y=0.955 $X2=0 $Y2=0
cc_126 N_D_c_126_n N_GATE_N_c_152_n 0.0388821f $X=0.51 $Y=1.895 $X2=0 $Y2=0
cc_127 D N_GATE_N_c_152_n 0.00201746f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_128 N_D_c_126_n GATE_N 3.62002e-19 $X=0.51 $Y=1.895 $X2=0 $Y2=0
cc_129 D GATE_N 0.0264884f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_130 N_D_M1012_g N_A_232_98#_c_189_n 0.00114236f $X=0.495 $Y=0.955 $X2=0 $Y2=0
cc_131 N_D_M1012_g N_A_27_136#_c_312_n 0.00672937f $X=0.495 $Y=0.955 $X2=0 $Y2=0
cc_132 N_D_M1012_g N_A_27_136#_c_313_n 0.0118249f $X=0.495 $Y=0.955 $X2=0 $Y2=0
cc_133 N_D_M1012_g N_A_27_136#_c_314_n 0.00420241f $X=0.495 $Y=0.955 $X2=0 $Y2=0
cc_134 N_D_M1012_g N_A_27_136#_c_316_n 0.00637197f $X=0.495 $Y=0.955 $X2=0 $Y2=0
cc_135 D N_A_27_136#_c_316_n 6.29576e-19 $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_136 N_D_c_126_n N_A_27_136#_c_320_n 0.0145926f $X=0.51 $Y=1.895 $X2=0 $Y2=0
cc_137 D N_A_27_136#_c_320_n 0.00111755f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_138 N_D_M1012_g N_A_27_136#_c_317_n 0.0169137f $X=0.495 $Y=0.955 $X2=0 $Y2=0
cc_139 D N_A_27_136#_c_317_n 0.0251401f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_140 N_D_c_126_n N_VPWR_c_737_n 0.0145591f $X=0.51 $Y=1.895 $X2=0 $Y2=0
cc_141 D N_VPWR_c_737_n 0.0153846f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_142 N_D_c_126_n N_VPWR_c_736_n 0.00499434f $X=0.51 $Y=1.895 $X2=0 $Y2=0
cc_143 N_D_c_126_n N_VPWR_c_746_n 0.00463894f $X=0.51 $Y=1.895 $X2=0 $Y2=0
cc_144 N_D_M1012_g N_VGND_c_838_n 0.00297615f $X=0.495 $Y=0.955 $X2=0 $Y2=0
cc_145 N_D_M1012_g N_VGND_c_840_n 0.00454494f $X=0.495 $Y=0.955 $X2=0 $Y2=0
cc_146 N_GATE_N_M1001_g N_A_232_98#_c_188_n 0.00268628f $X=1.085 $Y=0.86 $X2=0
+ $Y2=0
cc_147 N_GATE_N_c_152_n N_A_232_98#_c_188_n 0.0116346f $X=1.13 $Y=1.895 $X2=0
+ $Y2=0
cc_148 GATE_N N_A_232_98#_c_188_n 2.4045e-19 $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_149 N_GATE_N_M1001_g N_A_232_98#_c_189_n 0.0111812f $X=1.085 $Y=0.86 $X2=0
+ $Y2=0
cc_150 N_GATE_N_c_152_n N_A_232_98#_c_189_n 0.00124885f $X=1.13 $Y=1.895 $X2=0
+ $Y2=0
cc_151 GATE_N N_A_232_98#_c_189_n 0.0185311f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_152 N_GATE_N_c_152_n N_A_232_98#_c_197_n 0.00700717f $X=1.13 $Y=1.895 $X2=0
+ $Y2=0
cc_153 N_GATE_N_M1001_g N_A_232_98#_c_190_n 0.00486829f $X=1.085 $Y=0.86 $X2=0
+ $Y2=0
cc_154 N_GATE_N_c_152_n N_A_232_98#_c_190_n 0.00135318f $X=1.13 $Y=1.895 $X2=0
+ $Y2=0
cc_155 GATE_N N_A_232_98#_c_190_n 0.0177666f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_156 N_GATE_N_c_152_n N_A_232_98#_c_200_n 0.00390615f $X=1.13 $Y=1.895 $X2=0
+ $Y2=0
cc_157 N_GATE_N_c_152_n N_A_232_98#_c_202_n 0.00450473f $X=1.13 $Y=1.895 $X2=0
+ $Y2=0
cc_158 GATE_N N_A_232_98#_c_202_n 0.0120553f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_159 N_GATE_N_c_152_n N_A_232_98#_c_203_n 0.00762749f $X=1.13 $Y=1.895 $X2=0
+ $Y2=0
cc_160 GATE_N N_A_232_98#_c_203_n 0.0082296f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_161 N_GATE_N_M1001_g N_A_27_136#_c_312_n 0.00178342f $X=1.085 $Y=0.86 $X2=0
+ $Y2=0
cc_162 N_GATE_N_M1001_g N_A_27_136#_c_313_n 0.0155433f $X=1.085 $Y=0.86 $X2=0
+ $Y2=0
cc_163 N_GATE_N_c_152_n N_A_357_392#_c_399_n 5.76387e-19 $X=1.13 $Y=1.895 $X2=0
+ $Y2=0
cc_164 N_GATE_N_c_152_n N_VPWR_c_737_n 0.0120148f $X=1.13 $Y=1.895 $X2=0 $Y2=0
cc_165 N_GATE_N_c_152_n N_VPWR_c_740_n 0.00463088f $X=1.13 $Y=1.895 $X2=0 $Y2=0
cc_166 N_GATE_N_c_152_n N_VPWR_c_736_n 0.00499434f $X=1.13 $Y=1.895 $X2=0 $Y2=0
cc_167 N_GATE_N_M1001_g N_VGND_c_840_n 0.00508379f $X=1.085 $Y=0.86 $X2=0 $Y2=0
cc_168 N_GATE_N_M1001_g N_VGND_c_841_n 0.00210264f $X=1.085 $Y=0.86 $X2=0 $Y2=0
cc_169 N_GATE_N_M1001_g N_VGND_c_842_n 0.00374721f $X=1.085 $Y=0.86 $X2=0 $Y2=0
cc_170 N_A_232_98#_c_185_n N_A_27_136#_c_308_n 0.00433445f $X=2.155 $Y=1.885
+ $X2=0 $Y2=0
cc_171 N_A_232_98#_M1015_g N_A_27_136#_c_308_n 0.0167468f $X=2.225 $Y=0.78 $X2=0
+ $Y2=0
cc_172 N_A_232_98#_c_185_n N_A_27_136#_c_309_n 0.00851977f $X=2.155 $Y=1.885
+ $X2=0 $Y2=0
cc_173 N_A_232_98#_c_185_n N_A_27_136#_c_319_n 0.0252751f $X=2.155 $Y=1.885
+ $X2=0 $Y2=0
cc_174 N_A_232_98#_c_199_n N_A_27_136#_c_319_n 0.0141293f $X=3.915 $Y=2.605
+ $X2=0 $Y2=0
cc_175 N_A_232_98#_M1017_g N_A_27_136#_c_311_n 0.0550157f $X=3.72 $Y=0.69 $X2=0
+ $Y2=0
cc_176 N_A_232_98#_c_189_n N_A_27_136#_c_312_n 0.00886663f $X=1.505 $Y=1.085
+ $X2=0 $Y2=0
cc_177 N_A_232_98#_M1001_d N_A_27_136#_c_313_n 0.00639363f $X=1.16 $Y=0.49 $X2=0
+ $Y2=0
cc_178 N_A_232_98#_M1015_g N_A_27_136#_c_313_n 0.0168663f $X=2.225 $Y=0.78 $X2=0
+ $Y2=0
cc_179 N_A_232_98#_c_188_n N_A_27_136#_c_313_n 0.00122731f $X=2.065 $Y=1.505
+ $X2=0 $Y2=0
cc_180 N_A_232_98#_c_189_n N_A_27_136#_c_313_n 0.0289436f $X=1.505 $Y=1.085
+ $X2=0 $Y2=0
cc_181 N_A_232_98#_c_190_n N_A_27_136#_c_313_n 0.0193437f $X=1.59 $Y=1.67 $X2=0
+ $Y2=0
cc_182 N_A_232_98#_c_185_n N_A_27_136#_c_315_n 4.50657e-19 $X=2.155 $Y=1.885
+ $X2=0 $Y2=0
cc_183 N_A_232_98#_M1015_g N_A_27_136#_c_315_n 0.0113783f $X=2.225 $Y=0.78 $X2=0
+ $Y2=0
cc_184 N_A_232_98#_c_199_n N_A_357_392#_M1009_s 0.00942365f $X=3.915 $Y=2.605
+ $X2=0 $Y2=0
cc_185 N_A_232_98#_M1017_g N_A_357_392#_c_389_n 0.0180503f $X=3.72 $Y=0.69 $X2=0
+ $Y2=0
cc_186 N_A_232_98#_c_193_n N_A_357_392#_c_389_n 0.00673467f $X=3.875 $Y=2.03
+ $X2=0 $Y2=0
cc_187 N_A_232_98#_c_194_n N_A_357_392#_c_389_n 0.0150798f $X=3.89 $Y=2.465
+ $X2=0 $Y2=0
cc_188 N_A_232_98#_c_196_n N_A_357_392#_c_389_n 0.00339685f $X=3.875 $Y=1.805
+ $X2=0 $Y2=0
cc_189 N_A_232_98#_c_199_n N_A_357_392#_c_389_n 0.0142012f $X=3.915 $Y=2.605
+ $X2=0 $Y2=0
cc_190 N_A_232_98#_c_201_n N_A_357_392#_c_389_n 4.59072e-19 $X=4.08 $Y=2.195
+ $X2=0 $Y2=0
cc_191 N_A_232_98#_M1017_g N_A_357_392#_M1007_g 0.0215197f $X=3.72 $Y=0.69 $X2=0
+ $Y2=0
cc_192 N_A_232_98#_c_185_n N_A_357_392#_c_391_n 0.0217374f $X=2.155 $Y=1.885
+ $X2=0 $Y2=0
cc_193 N_A_232_98#_M1015_g N_A_357_392#_c_391_n 0.00592463f $X=2.225 $Y=0.78
+ $X2=0 $Y2=0
cc_194 N_A_232_98#_c_190_n N_A_357_392#_c_391_n 0.0315194f $X=1.59 $Y=1.67 $X2=0
+ $Y2=0
cc_195 N_A_232_98#_c_203_n N_A_357_392#_c_391_n 0.00641126f $X=1.432 $Y=1.95
+ $X2=0 $Y2=0
cc_196 N_A_232_98#_c_185_n N_A_357_392#_c_397_n 0.00187077f $X=2.155 $Y=1.885
+ $X2=0 $Y2=0
cc_197 N_A_232_98#_c_199_n N_A_357_392#_c_397_n 0.0247998f $X=3.915 $Y=2.605
+ $X2=0 $Y2=0
cc_198 N_A_232_98#_M1017_g N_A_357_392#_c_398_n 0.00119138f $X=3.72 $Y=0.69
+ $X2=0 $Y2=0
cc_199 N_A_232_98#_c_196_n N_A_357_392#_c_398_n 2.01574e-19 $X=3.875 $Y=1.805
+ $X2=0 $Y2=0
cc_200 N_A_232_98#_M1017_g N_A_357_392#_c_393_n 0.0228752f $X=3.72 $Y=0.69 $X2=0
+ $Y2=0
cc_201 N_A_232_98#_c_196_n N_A_357_392#_c_393_n 0.00101863f $X=3.875 $Y=1.805
+ $X2=0 $Y2=0
cc_202 N_A_232_98#_M1017_g N_A_357_392#_c_394_n 0.021337f $X=3.72 $Y=0.69 $X2=0
+ $Y2=0
cc_203 N_A_232_98#_c_194_n N_A_357_392#_c_394_n 0.00434555f $X=3.89 $Y=2.465
+ $X2=0 $Y2=0
cc_204 N_A_232_98#_c_185_n N_A_357_392#_c_395_n 3.54466e-19 $X=2.155 $Y=1.885
+ $X2=0 $Y2=0
cc_205 N_A_232_98#_M1015_g N_A_357_392#_c_395_n 0.00649689f $X=2.225 $Y=0.78
+ $X2=0 $Y2=0
cc_206 N_A_232_98#_c_188_n N_A_357_392#_c_395_n 0.00523096f $X=2.065 $Y=1.505
+ $X2=0 $Y2=0
cc_207 N_A_232_98#_c_190_n N_A_357_392#_c_395_n 0.026826f $X=1.59 $Y=1.67 $X2=0
+ $Y2=0
cc_208 N_A_232_98#_c_185_n N_A_357_392#_c_399_n 0.0184871f $X=2.155 $Y=1.885
+ $X2=0 $Y2=0
cc_209 N_A_232_98#_c_188_n N_A_357_392#_c_399_n 0.00514254f $X=2.065 $Y=1.505
+ $X2=0 $Y2=0
cc_210 N_A_232_98#_c_190_n N_A_357_392#_c_399_n 0.00494207f $X=1.59 $Y=1.67
+ $X2=0 $Y2=0
cc_211 N_A_232_98#_c_199_n N_A_357_392#_c_399_n 0.025181f $X=3.915 $Y=2.605
+ $X2=0 $Y2=0
cc_212 N_A_232_98#_c_203_n N_A_357_392#_c_399_n 0.0435783f $X=1.432 $Y=1.95
+ $X2=0 $Y2=0
cc_213 N_A_232_98#_c_194_n N_A_897_406#_c_492_n 0.0327659f $X=3.89 $Y=2.465
+ $X2=0 $Y2=0
cc_214 N_A_232_98#_c_199_n N_A_897_406#_c_492_n 0.00194059f $X=3.915 $Y=2.605
+ $X2=0 $Y2=0
cc_215 N_A_232_98#_c_201_n N_A_897_406#_c_492_n 0.00418318f $X=4.08 $Y=2.195
+ $X2=0 $Y2=0
cc_216 N_A_232_98#_c_196_n N_A_897_406#_c_484_n 0.00574774f $X=3.875 $Y=1.805
+ $X2=0 $Y2=0
cc_217 N_A_232_98#_c_194_n N_A_897_406#_c_495_n 0.00127573f $X=3.89 $Y=2.465
+ $X2=0 $Y2=0
cc_218 N_A_232_98#_c_201_n N_A_897_406#_c_495_n 0.0198487f $X=4.08 $Y=2.195
+ $X2=0 $Y2=0
cc_219 N_A_232_98#_c_199_n N_A_654_392#_M1002_d 0.0117896f $X=3.915 $Y=2.605
+ $X2=0 $Y2=0
cc_220 N_A_232_98#_c_194_n N_A_654_392#_c_607_n 0.00216866f $X=3.89 $Y=2.465
+ $X2=0 $Y2=0
cc_221 N_A_232_98#_c_199_n N_A_654_392#_c_607_n 0.0332943f $X=3.915 $Y=2.605
+ $X2=0 $Y2=0
cc_222 N_A_232_98#_c_201_n N_A_654_392#_c_607_n 0.013958f $X=4.08 $Y=2.195 $X2=0
+ $Y2=0
cc_223 N_A_232_98#_c_193_n N_A_654_392#_c_608_n 0.0058042f $X=3.875 $Y=2.03
+ $X2=0 $Y2=0
cc_224 N_A_232_98#_c_196_n N_A_654_392#_c_608_n 0.00325234f $X=3.875 $Y=1.805
+ $X2=0 $Y2=0
cc_225 N_A_232_98#_c_201_n N_A_654_392#_c_608_n 0.0112343f $X=4.08 $Y=2.195
+ $X2=0 $Y2=0
cc_226 N_A_232_98#_M1017_g N_A_654_392#_c_609_n 0.00176148f $X=3.72 $Y=0.69
+ $X2=0 $Y2=0
cc_227 N_A_232_98#_c_194_n N_A_654_392#_c_609_n 0.00129168f $X=3.89 $Y=2.465
+ $X2=0 $Y2=0
cc_228 N_A_232_98#_c_196_n N_A_654_392#_c_609_n 0.0119896f $X=3.875 $Y=1.805
+ $X2=0 $Y2=0
cc_229 N_A_232_98#_c_199_n N_A_654_392#_c_609_n 0.00394489f $X=3.915 $Y=2.605
+ $X2=0 $Y2=0
cc_230 N_A_232_98#_c_201_n N_A_654_392#_c_609_n 0.0260226f $X=4.08 $Y=2.195
+ $X2=0 $Y2=0
cc_231 N_A_232_98#_M1017_g N_A_654_392#_c_610_n 0.00198035f $X=3.72 $Y=0.69
+ $X2=0 $Y2=0
cc_232 N_A_232_98#_c_196_n N_A_654_392#_c_610_n 0.00200433f $X=3.875 $Y=1.805
+ $X2=0 $Y2=0
cc_233 N_A_232_98#_M1017_g N_A_654_392#_c_599_n 7.62689e-19 $X=3.72 $Y=0.69
+ $X2=0 $Y2=0
cc_234 N_A_232_98#_M1017_g N_A_654_392#_c_601_n 0.00113438f $X=3.72 $Y=0.69
+ $X2=0 $Y2=0
cc_235 N_A_232_98#_c_199_n N_VPWR_M1009_d 0.0113312f $X=3.915 $Y=2.605 $X2=0
+ $Y2=0
cc_236 N_A_232_98#_c_200_n N_VPWR_c_737_n 0.0218701f $X=1.675 $Y=2.605 $X2=0
+ $Y2=0
cc_237 N_A_232_98#_c_202_n N_VPWR_c_737_n 0.0393897f $X=1.355 $Y=2.115 $X2=0
+ $Y2=0
cc_238 N_A_232_98#_c_185_n N_VPWR_c_738_n 0.00201997f $X=2.155 $Y=1.885 $X2=0
+ $Y2=0
cc_239 N_A_232_98#_c_199_n N_VPWR_c_738_n 0.0250768f $X=3.915 $Y=2.605 $X2=0
+ $Y2=0
cc_240 N_A_232_98#_c_185_n N_VPWR_c_740_n 0.00361055f $X=2.155 $Y=1.885 $X2=0
+ $Y2=0
cc_241 N_A_232_98#_c_199_n N_VPWR_c_740_n 0.00982449f $X=3.915 $Y=2.605 $X2=0
+ $Y2=0
cc_242 N_A_232_98#_c_200_n N_VPWR_c_740_n 0.0133755f $X=1.675 $Y=2.605 $X2=0
+ $Y2=0
cc_243 N_A_232_98#_c_194_n N_VPWR_c_742_n 0.00326703f $X=3.89 $Y=2.465 $X2=0
+ $Y2=0
cc_244 N_A_232_98#_c_199_n N_VPWR_c_742_n 0.0252287f $X=3.915 $Y=2.605 $X2=0
+ $Y2=0
cc_245 N_A_232_98#_c_185_n N_VPWR_c_736_n 0.0049649f $X=2.155 $Y=1.885 $X2=0
+ $Y2=0
cc_246 N_A_232_98#_c_194_n N_VPWR_c_736_n 0.00418893f $X=3.89 $Y=2.465 $X2=0
+ $Y2=0
cc_247 N_A_232_98#_c_199_n N_VPWR_c_736_n 0.0634281f $X=3.915 $Y=2.605 $X2=0
+ $Y2=0
cc_248 N_A_232_98#_c_200_n N_VPWR_c_736_n 0.0162101f $X=1.675 $Y=2.605 $X2=0
+ $Y2=0
cc_249 N_A_232_98#_c_194_n N_VPWR_c_747_n 0.001799f $X=3.89 $Y=2.465 $X2=0 $Y2=0
cc_250 N_A_232_98#_c_199_n N_VPWR_c_747_n 0.00735006f $X=3.915 $Y=2.605 $X2=0
+ $Y2=0
cc_251 N_A_232_98#_c_199_n A_570_392# 0.00557976f $X=3.915 $Y=2.605 $X2=-0.19
+ $Y2=-0.245
cc_252 N_A_232_98#_c_199_n A_793_508# 0.0067331f $X=3.915 $Y=2.605 $X2=-0.19
+ $Y2=-0.245
cc_253 N_A_232_98#_M1017_g N_VGND_c_834_n 0.00461464f $X=3.72 $Y=0.69 $X2=0
+ $Y2=0
cc_254 N_A_232_98#_M1015_g N_VGND_c_840_n 0.00533081f $X=2.225 $Y=0.78 $X2=0
+ $Y2=0
cc_255 N_A_232_98#_M1017_g N_VGND_c_840_n 0.00909529f $X=3.72 $Y=0.69 $X2=0
+ $Y2=0
cc_256 N_A_232_98#_M1015_g N_VGND_c_842_n 0.00414982f $X=2.225 $Y=0.78 $X2=0
+ $Y2=0
cc_257 N_A_232_98#_M1015_g N_VGND_c_843_n 0.0060117f $X=2.225 $Y=0.78 $X2=0
+ $Y2=0
cc_258 N_A_27_136#_c_313_n N_A_357_392#_M1015_s 0.00690466f $X=2.535 $Y=0.665
+ $X2=-0.19 $Y2=-0.245
cc_259 N_A_27_136#_c_308_n N_A_357_392#_c_389_n 0.0209724f $X=2.775 $Y=1.59
+ $X2=0 $Y2=0
cc_260 N_A_27_136#_c_309_n N_A_357_392#_c_389_n 0.00573481f $X=2.775 $Y=1.795
+ $X2=0 $Y2=0
cc_261 N_A_27_136#_c_319_n N_A_357_392#_c_389_n 0.0598349f $X=2.775 $Y=1.885
+ $X2=0 $Y2=0
cc_262 N_A_27_136#_c_310_n N_A_357_392#_c_389_n 0.0214145f $X=3.255 $Y=1.16
+ $X2=0 $Y2=0
cc_263 N_A_27_136#_c_315_n N_A_357_392#_c_389_n 3.38535e-19 $X=2.7 $Y=1.425
+ $X2=0 $Y2=0
cc_264 N_A_27_136#_c_308_n N_A_357_392#_c_391_n 0.00125202f $X=2.775 $Y=1.59
+ $X2=0 $Y2=0
cc_265 N_A_27_136#_c_309_n N_A_357_392#_c_391_n 0.0014328f $X=2.775 $Y=1.795
+ $X2=0 $Y2=0
cc_266 N_A_27_136#_c_315_n N_A_357_392#_c_391_n 0.0199283f $X=2.7 $Y=1.425 $X2=0
+ $Y2=0
cc_267 N_A_27_136#_c_308_n N_A_357_392#_c_397_n 9.68515e-19 $X=2.775 $Y=1.59
+ $X2=0 $Y2=0
cc_268 N_A_27_136#_c_319_n N_A_357_392#_c_397_n 0.0143888f $X=2.775 $Y=1.885
+ $X2=0 $Y2=0
cc_269 N_A_27_136#_c_310_n N_A_357_392#_c_397_n 0.00455655f $X=3.255 $Y=1.16
+ $X2=0 $Y2=0
cc_270 N_A_27_136#_c_315_n N_A_357_392#_c_397_n 0.0189066f $X=2.7 $Y=1.425 $X2=0
+ $Y2=0
cc_271 N_A_27_136#_c_308_n N_A_357_392#_c_398_n 0.00149274f $X=2.775 $Y=1.59
+ $X2=0 $Y2=0
cc_272 N_A_27_136#_c_309_n N_A_357_392#_c_398_n 0.00141758f $X=2.775 $Y=1.795
+ $X2=0 $Y2=0
cc_273 N_A_27_136#_c_315_n N_A_357_392#_c_398_n 0.00440446f $X=2.7 $Y=1.425
+ $X2=0 $Y2=0
cc_274 N_A_27_136#_c_308_n N_A_357_392#_c_392_n 0.00497266f $X=2.775 $Y=1.59
+ $X2=0 $Y2=0
cc_275 N_A_27_136#_c_310_n N_A_357_392#_c_392_n 0.021332f $X=3.255 $Y=1.16 $X2=0
+ $Y2=0
cc_276 N_A_27_136#_c_315_n N_A_357_392#_c_392_n 0.0231983f $X=2.7 $Y=1.425 $X2=0
+ $Y2=0
cc_277 N_A_27_136#_c_313_n N_A_357_392#_c_395_n 0.025204f $X=2.535 $Y=0.665
+ $X2=0 $Y2=0
cc_278 N_A_27_136#_c_315_n N_A_357_392#_c_395_n 0.0130374f $X=2.7 $Y=1.425 $X2=0
+ $Y2=0
cc_279 N_A_27_136#_c_319_n N_A_654_392#_c_607_n 8.04279e-19 $X=2.775 $Y=1.885
+ $X2=0 $Y2=0
cc_280 N_A_27_136#_c_320_n N_VPWR_c_737_n 0.0594947f $X=0.285 $Y=2.115 $X2=0
+ $Y2=0
cc_281 N_A_27_136#_c_319_n N_VPWR_c_738_n 0.00860015f $X=2.775 $Y=1.885 $X2=0
+ $Y2=0
cc_282 N_A_27_136#_c_319_n N_VPWR_c_742_n 0.00326738f $X=2.775 $Y=1.885 $X2=0
+ $Y2=0
cc_283 N_A_27_136#_c_319_n N_VPWR_c_736_n 0.0041926f $X=2.775 $Y=1.885 $X2=0
+ $Y2=0
cc_284 N_A_27_136#_c_320_n N_VPWR_c_736_n 0.011795f $X=0.285 $Y=2.115 $X2=0
+ $Y2=0
cc_285 N_A_27_136#_c_320_n N_VPWR_c_746_n 0.00972743f $X=0.285 $Y=2.115 $X2=0
+ $Y2=0
cc_286 N_A_27_136#_c_313_n N_VGND_M1012_d 0.0162931f $X=2.535 $Y=0.665 $X2=-0.19
+ $Y2=-0.245
cc_287 N_A_27_136#_c_313_n N_VGND_M1015_d 0.0184311f $X=2.535 $Y=0.665 $X2=0
+ $Y2=0
cc_288 N_A_27_136#_c_315_n N_VGND_M1015_d 0.011441f $X=2.7 $Y=1.425 $X2=0 $Y2=0
cc_289 N_A_27_136#_c_311_n N_VGND_c_834_n 0.00461464f $X=3.33 $Y=1.085 $X2=0
+ $Y2=0
cc_290 N_A_27_136#_c_313_n N_VGND_c_838_n 0.00345394f $X=2.535 $Y=0.665 $X2=0
+ $Y2=0
cc_291 N_A_27_136#_c_314_n N_VGND_c_838_n 0.00791634f $X=0.445 $Y=0.665 $X2=0
+ $Y2=0
cc_292 N_A_27_136#_c_311_n N_VGND_c_840_n 0.00913019f $X=3.33 $Y=1.085 $X2=0
+ $Y2=0
cc_293 N_A_27_136#_c_313_n N_VGND_c_840_n 0.0511453f $X=2.535 $Y=0.665 $X2=0
+ $Y2=0
cc_294 N_A_27_136#_c_314_n N_VGND_c_840_n 0.011025f $X=0.445 $Y=0.665 $X2=0
+ $Y2=0
cc_295 N_A_27_136#_c_313_n N_VGND_c_841_n 0.0246008f $X=2.535 $Y=0.665 $X2=0
+ $Y2=0
cc_296 N_A_27_136#_c_313_n N_VGND_c_842_n 0.0258079f $X=2.535 $Y=0.665 $X2=0
+ $Y2=0
cc_297 N_A_27_136#_c_308_n N_VGND_c_843_n 0.00817797f $X=2.775 $Y=1.59 $X2=0
+ $Y2=0
cc_298 N_A_27_136#_c_311_n N_VGND_c_843_n 0.00642663f $X=3.33 $Y=1.085 $X2=0
+ $Y2=0
cc_299 N_A_27_136#_c_313_n N_VGND_c_843_n 0.0404537f $X=2.535 $Y=0.665 $X2=0
+ $Y2=0
cc_300 N_A_357_392#_M1007_g N_A_897_406#_M1004_g 0.0427152f $X=4.195 $Y=0.58
+ $X2=0 $Y2=0
cc_301 N_A_357_392#_c_393_n N_A_897_406#_M1004_g 0.00116465f $X=4.17 $Y=1.355
+ $X2=0 $Y2=0
cc_302 N_A_357_392#_c_394_n N_A_897_406#_M1004_g 0.0179408f $X=4.17 $Y=1.355
+ $X2=0 $Y2=0
cc_303 N_A_357_392#_c_394_n N_A_897_406#_c_484_n 0.00150268f $X=4.17 $Y=1.355
+ $X2=0 $Y2=0
cc_304 N_A_357_392#_c_397_n N_A_654_392#_M1002_d 0.00134049f $X=3.075 $Y=1.925
+ $X2=0 $Y2=0
cc_305 N_A_357_392#_c_389_n N_A_654_392#_c_607_n 0.00387534f $X=3.195 $Y=1.885
+ $X2=0 $Y2=0
cc_306 N_A_357_392#_c_397_n N_A_654_392#_c_607_n 0.00745454f $X=3.075 $Y=1.925
+ $X2=0 $Y2=0
cc_307 N_A_357_392#_c_393_n N_A_654_392#_c_607_n 0.00494788f $X=4.17 $Y=1.355
+ $X2=0 $Y2=0
cc_308 N_A_357_392#_c_389_n N_A_654_392#_c_608_n 0.00321088f $X=3.195 $Y=1.885
+ $X2=0 $Y2=0
cc_309 N_A_357_392#_c_397_n N_A_654_392#_c_608_n 0.0125414f $X=3.075 $Y=1.925
+ $X2=0 $Y2=0
cc_310 N_A_357_392#_c_393_n N_A_654_392#_c_609_n 0.0449862f $X=4.17 $Y=1.355
+ $X2=0 $Y2=0
cc_311 N_A_357_392#_c_394_n N_A_654_392#_c_609_n 0.00440959f $X=4.17 $Y=1.355
+ $X2=0 $Y2=0
cc_312 N_A_357_392#_c_389_n N_A_654_392#_c_610_n 8.30345e-19 $X=3.195 $Y=1.885
+ $X2=0 $Y2=0
cc_313 N_A_357_392#_c_397_n N_A_654_392#_c_610_n 0.00187356f $X=3.075 $Y=1.925
+ $X2=0 $Y2=0
cc_314 N_A_357_392#_c_398_n N_A_654_392#_c_610_n 0.0128753f $X=3.24 $Y=1.61
+ $X2=0 $Y2=0
cc_315 N_A_357_392#_c_393_n N_A_654_392#_c_610_n 0.0141411f $X=4.17 $Y=1.355
+ $X2=0 $Y2=0
cc_316 N_A_357_392#_M1007_g N_A_654_392#_c_599_n 0.0102957f $X=4.195 $Y=0.58
+ $X2=0 $Y2=0
cc_317 N_A_357_392#_M1007_g N_A_654_392#_c_600_n 0.00848162f $X=4.195 $Y=0.58
+ $X2=0 $Y2=0
cc_318 N_A_357_392#_c_393_n N_A_654_392#_c_600_n 0.0137779f $X=4.17 $Y=1.355
+ $X2=0 $Y2=0
cc_319 N_A_357_392#_c_394_n N_A_654_392#_c_600_n 0.00145734f $X=4.17 $Y=1.355
+ $X2=0 $Y2=0
cc_320 N_A_357_392#_M1007_g N_A_654_392#_c_601_n 0.00270231f $X=4.195 $Y=0.58
+ $X2=0 $Y2=0
cc_321 N_A_357_392#_c_393_n N_A_654_392#_c_601_n 0.0284678f $X=4.17 $Y=1.355
+ $X2=0 $Y2=0
cc_322 N_A_357_392#_c_394_n N_A_654_392#_c_601_n 0.00267329f $X=4.17 $Y=1.355
+ $X2=0 $Y2=0
cc_323 N_A_357_392#_c_393_n N_A_654_392#_c_602_n 0.00345296f $X=4.17 $Y=1.355
+ $X2=0 $Y2=0
cc_324 N_A_357_392#_c_393_n N_A_654_392#_c_603_n 0.00746488f $X=4.17 $Y=1.355
+ $X2=0 $Y2=0
cc_325 N_A_357_392#_c_397_n N_VPWR_M1009_d 0.00671554f $X=3.075 $Y=1.925 $X2=0
+ $Y2=0
cc_326 N_A_357_392#_c_389_n N_VPWR_c_742_n 0.00326738f $X=3.195 $Y=1.885 $X2=0
+ $Y2=0
cc_327 N_A_357_392#_c_389_n N_VPWR_c_736_n 0.00416973f $X=3.195 $Y=1.885 $X2=0
+ $Y2=0
cc_328 N_A_357_392#_c_397_n A_570_392# 0.00284769f $X=3.075 $Y=1.925 $X2=-0.19
+ $Y2=-0.245
cc_329 N_A_357_392#_M1007_g N_VGND_c_832_n 0.00151896f $X=4.195 $Y=0.58 $X2=0
+ $Y2=0
cc_330 N_A_357_392#_M1007_g N_VGND_c_834_n 0.00434272f $X=4.195 $Y=0.58 $X2=0
+ $Y2=0
cc_331 N_A_357_392#_M1007_g N_VGND_c_840_n 0.00448673f $X=4.195 $Y=0.58 $X2=0
+ $Y2=0
cc_332 N_A_897_406#_c_497_n N_A_654_392#_c_595_n 0.0023113f $X=5.715 $Y=1.805
+ $X2=0 $Y2=0
cc_333 N_A_897_406#_c_490_n N_A_654_392#_c_595_n 0.010923f $X=5.715 $Y=1.72
+ $X2=0 $Y2=0
cc_334 N_A_897_406#_M1004_g N_A_654_392#_c_596_n 0.00666444f $X=4.62 $Y=0.58
+ $X2=0 $Y2=0
cc_335 N_A_897_406#_c_489_n N_A_654_392#_c_596_n 0.00949746f $X=5.437 $Y=1.13
+ $X2=0 $Y2=0
cc_336 N_A_897_406#_c_492_n N_A_654_392#_c_605_n 0.00451717f $X=4.575 $Y=2.465
+ $X2=0 $Y2=0
cc_337 N_A_897_406#_c_484_n N_A_654_392#_c_605_n 0.00467639f $X=4.65 $Y=2.03
+ $X2=0 $Y2=0
cc_338 N_A_897_406#_c_495_n N_A_654_392#_c_605_n 0.0118431f $X=5.465 $Y=2.195
+ $X2=0 $Y2=0
cc_339 N_A_897_406#_c_497_n N_A_654_392#_c_605_n 0.0290042f $X=5.715 $Y=1.805
+ $X2=0 $Y2=0
cc_340 N_A_897_406#_c_499_n N_A_654_392#_c_605_n 0.00820023f $X=5.8 $Y=2.34
+ $X2=0 $Y2=0
cc_341 N_A_897_406#_c_488_n N_A_654_392#_c_597_n 0.0147933f $X=5.405 $Y=0.515
+ $X2=0 $Y2=0
cc_342 N_A_897_406#_c_489_n N_A_654_392#_c_597_n 0.00476794f $X=5.437 $Y=1.13
+ $X2=0 $Y2=0
cc_343 N_A_897_406#_c_490_n N_A_654_392#_c_597_n 0.00192894f $X=5.715 $Y=1.72
+ $X2=0 $Y2=0
cc_344 N_A_897_406#_c_484_n N_A_654_392#_c_598_n 0.0101642f $X=4.65 $Y=2.03
+ $X2=0 $Y2=0
cc_345 N_A_897_406#_c_495_n N_A_654_392#_c_598_n 0.00855638f $X=5.465 $Y=2.195
+ $X2=0 $Y2=0
cc_346 N_A_897_406#_c_497_n N_A_654_392#_c_598_n 0.00204104f $X=5.715 $Y=1.805
+ $X2=0 $Y2=0
cc_347 N_A_897_406#_c_490_n N_A_654_392#_c_598_n 0.00655086f $X=5.715 $Y=1.72
+ $X2=0 $Y2=0
cc_348 N_A_897_406#_c_492_n N_A_654_392#_c_609_n 0.0038768f $X=4.575 $Y=2.465
+ $X2=0 $Y2=0
cc_349 N_A_897_406#_c_484_n N_A_654_392#_c_609_n 0.0147233f $X=4.65 $Y=2.03
+ $X2=0 $Y2=0
cc_350 N_A_897_406#_c_487_n N_A_654_392#_c_609_n 4.39555e-19 $X=4.635 $Y=1.49
+ $X2=0 $Y2=0
cc_351 N_A_897_406#_c_495_n N_A_654_392#_c_609_n 0.0309417f $X=5.465 $Y=2.195
+ $X2=0 $Y2=0
cc_352 N_A_897_406#_M1004_g N_A_654_392#_c_599_n 0.00179535f $X=4.62 $Y=0.58
+ $X2=0 $Y2=0
cc_353 N_A_897_406#_M1004_g N_A_654_392#_c_600_n 0.0153082f $X=4.62 $Y=0.58
+ $X2=0 $Y2=0
cc_354 N_A_897_406#_c_487_n N_A_654_392#_c_600_n 7.81529e-19 $X=4.635 $Y=1.49
+ $X2=0 $Y2=0
cc_355 N_A_897_406#_c_488_n N_A_654_392#_c_600_n 0.0151911f $X=5.405 $Y=0.515
+ $X2=0 $Y2=0
cc_356 N_A_897_406#_M1004_g N_A_654_392#_c_602_n 0.00650161f $X=4.62 $Y=0.58
+ $X2=0 $Y2=0
cc_357 N_A_897_406#_c_489_n N_A_654_392#_c_602_n 0.00880982f $X=5.437 $Y=1.13
+ $X2=0 $Y2=0
cc_358 N_A_897_406#_c_490_n N_A_654_392#_c_602_n 0.00622767f $X=5.715 $Y=1.72
+ $X2=0 $Y2=0
cc_359 N_A_897_406#_M1004_g N_A_654_392#_c_603_n 4.02061e-19 $X=4.62 $Y=0.58
+ $X2=0 $Y2=0
cc_360 N_A_897_406#_c_487_n N_A_654_392#_c_603_n 0.00573586f $X=4.635 $Y=1.49
+ $X2=0 $Y2=0
cc_361 N_A_897_406#_c_495_n N_A_654_392#_c_603_n 0.0242337f $X=5.465 $Y=2.195
+ $X2=0 $Y2=0
cc_362 N_A_897_406#_c_489_n N_A_654_392#_c_603_n 0.00457555f $X=5.437 $Y=1.13
+ $X2=0 $Y2=0
cc_363 N_A_897_406#_c_490_n N_A_654_392#_c_603_n 0.034501f $X=5.715 $Y=1.72
+ $X2=0 $Y2=0
cc_364 N_A_897_406#_c_487_n N_A_654_392#_c_604_n 0.00974488f $X=4.635 $Y=1.49
+ $X2=0 $Y2=0
cc_365 N_A_897_406#_c_490_n N_A_654_392#_c_604_n 2.42207e-19 $X=5.715 $Y=1.72
+ $X2=0 $Y2=0
cc_366 N_A_897_406#_M1014_g N_RESET_B_c_702_n 0.0197034f $X=6.6 $Y=0.74
+ $X2=-0.19 $Y2=-0.245
cc_367 N_A_897_406#_c_488_n N_RESET_B_c_702_n 0.00312003f $X=5.405 $Y=0.515
+ $X2=-0.19 $Y2=-0.245
cc_368 N_A_897_406#_M1014_g N_RESET_B_c_703_n 0.00457497f $X=6.6 $Y=0.74 $X2=0
+ $Y2=0
cc_369 N_A_897_406#_c_486_n N_RESET_B_c_703_n 0.0451007f $X=6.695 $Y=1.765 $X2=0
+ $Y2=0
cc_370 N_A_897_406#_c_496_n N_RESET_B_c_703_n 0.0166029f $X=6.415 $Y=1.805 $X2=0
+ $Y2=0
cc_371 N_A_897_406#_c_497_n N_RESET_B_c_703_n 0.015505f $X=5.715 $Y=1.805 $X2=0
+ $Y2=0
cc_372 N_A_897_406#_c_490_n N_RESET_B_c_703_n 0.00451451f $X=5.715 $Y=1.72 $X2=0
+ $Y2=0
cc_373 N_A_897_406#_c_491_n N_RESET_B_c_703_n 0.00503565f $X=6.61 $Y=1.485 $X2=0
+ $Y2=0
cc_374 N_A_897_406#_M1014_g RESET_B 0.00149724f $X=6.6 $Y=0.74 $X2=0 $Y2=0
cc_375 N_A_897_406#_c_486_n RESET_B 2.70907e-19 $X=6.695 $Y=1.765 $X2=0 $Y2=0
cc_376 N_A_897_406#_c_496_n RESET_B 0.0198218f $X=6.415 $Y=1.805 $X2=0 $Y2=0
cc_377 N_A_897_406#_c_497_n RESET_B 0.00674165f $X=5.715 $Y=1.805 $X2=0 $Y2=0
cc_378 N_A_897_406#_c_490_n RESET_B 0.0218949f $X=5.715 $Y=1.72 $X2=0 $Y2=0
cc_379 N_A_897_406#_c_491_n RESET_B 0.0177152f $X=6.61 $Y=1.485 $X2=0 $Y2=0
cc_380 N_A_897_406#_c_495_n N_VPWR_M1018_d 0.00655572f $X=5.465 $Y=2.195 $X2=0
+ $Y2=0
cc_381 N_A_897_406#_c_496_n N_VPWR_M1016_d 0.00230596f $X=6.415 $Y=1.805 $X2=0
+ $Y2=0
cc_382 N_A_897_406#_c_491_n N_VPWR_M1016_d 0.00203861f $X=6.61 $Y=1.485 $X2=0
+ $Y2=0
cc_383 N_A_897_406#_c_486_n N_VPWR_c_739_n 0.0113564f $X=6.695 $Y=1.765 $X2=0
+ $Y2=0
cc_384 N_A_897_406#_c_496_n N_VPWR_c_739_n 0.0128995f $X=6.415 $Y=1.805 $X2=0
+ $Y2=0
cc_385 N_A_897_406#_c_497_n N_VPWR_c_739_n 0.0438551f $X=5.715 $Y=1.805 $X2=0
+ $Y2=0
cc_386 N_A_897_406#_c_491_n N_VPWR_c_739_n 0.0131716f $X=6.61 $Y=1.485 $X2=0
+ $Y2=0
cc_387 N_A_897_406#_c_492_n N_VPWR_c_742_n 0.00415318f $X=4.575 $Y=2.465 $X2=0
+ $Y2=0
cc_388 N_A_897_406#_c_499_n N_VPWR_c_743_n 0.00983421f $X=5.8 $Y=2.34 $X2=0
+ $Y2=0
cc_389 N_A_897_406#_c_486_n N_VPWR_c_744_n 0.00445602f $X=6.695 $Y=1.765 $X2=0
+ $Y2=0
cc_390 N_A_897_406#_c_492_n N_VPWR_c_736_n 0.00854473f $X=4.575 $Y=2.465 $X2=0
+ $Y2=0
cc_391 N_A_897_406#_c_486_n N_VPWR_c_736_n 0.00865213f $X=6.695 $Y=1.765 $X2=0
+ $Y2=0
cc_392 N_A_897_406#_c_499_n N_VPWR_c_736_n 0.011205f $X=5.8 $Y=2.34 $X2=0 $Y2=0
cc_393 N_A_897_406#_c_492_n N_VPWR_c_747_n 0.0213766f $X=4.575 $Y=2.465 $X2=0
+ $Y2=0
cc_394 N_A_897_406#_c_495_n N_VPWR_c_747_n 0.0634565f $X=5.465 $Y=2.195 $X2=0
+ $Y2=0
cc_395 N_A_897_406#_c_499_n N_VPWR_c_747_n 0.0234615f $X=5.8 $Y=2.34 $X2=0 $Y2=0
cc_396 N_A_897_406#_M1014_g N_Q_c_810_n 0.015485f $X=6.6 $Y=0.74 $X2=0 $Y2=0
cc_397 N_A_897_406#_c_486_n N_Q_c_811_n 7.88609e-19 $X=6.695 $Y=1.765 $X2=0
+ $Y2=0
cc_398 N_A_897_406#_c_491_n N_Q_c_811_n 0.00342799f $X=6.61 $Y=1.485 $X2=0 $Y2=0
cc_399 N_A_897_406#_c_486_n Q 0.00413071f $X=6.695 $Y=1.765 $X2=0 $Y2=0
cc_400 N_A_897_406#_c_491_n Q 0.00509501f $X=6.61 $Y=1.485 $X2=0 $Y2=0
cc_401 N_A_897_406#_c_486_n Q 0.0116369f $X=6.695 $Y=1.765 $X2=0 $Y2=0
cc_402 N_A_897_406#_M1014_g N_Q_c_812_n 0.00429103f $X=6.6 $Y=0.74 $X2=0 $Y2=0
cc_403 N_A_897_406#_c_486_n N_Q_c_812_n 0.0101667f $X=6.695 $Y=1.765 $X2=0 $Y2=0
cc_404 N_A_897_406#_c_491_n N_Q_c_812_n 0.0307041f $X=6.61 $Y=1.485 $X2=0 $Y2=0
cc_405 N_A_897_406#_M1004_g N_VGND_c_832_n 0.0112076f $X=4.62 $Y=0.58 $X2=0
+ $Y2=0
cc_406 N_A_897_406#_c_488_n N_VGND_c_832_n 0.022605f $X=5.405 $Y=0.515 $X2=0
+ $Y2=0
cc_407 N_A_897_406#_M1014_g N_VGND_c_833_n 0.00734264f $X=6.6 $Y=0.74 $X2=0
+ $Y2=0
cc_408 N_A_897_406#_c_488_n N_VGND_c_833_n 0.0108156f $X=5.405 $Y=0.515 $X2=0
+ $Y2=0
cc_409 N_A_897_406#_c_491_n N_VGND_c_833_n 0.00303799f $X=6.61 $Y=1.485 $X2=0
+ $Y2=0
cc_410 N_A_897_406#_M1004_g N_VGND_c_834_n 0.00383152f $X=4.62 $Y=0.58 $X2=0
+ $Y2=0
cc_411 N_A_897_406#_c_488_n N_VGND_c_836_n 0.01727f $X=5.405 $Y=0.515 $X2=0
+ $Y2=0
cc_412 N_A_897_406#_M1014_g N_VGND_c_839_n 0.00461464f $X=6.6 $Y=0.74 $X2=0
+ $Y2=0
cc_413 N_A_897_406#_M1004_g N_VGND_c_840_n 0.00386109f $X=4.62 $Y=0.58 $X2=0
+ $Y2=0
cc_414 N_A_897_406#_M1014_g N_VGND_c_840_n 0.00913693f $X=6.6 $Y=0.74 $X2=0
+ $Y2=0
cc_415 N_A_897_406#_c_488_n N_VGND_c_840_n 0.0140855f $X=5.405 $Y=0.515 $X2=0
+ $Y2=0
cc_416 N_A_654_392#_c_597_n N_RESET_B_c_702_n 0.0491811f $X=5.62 $Y=1.185
+ $X2=-0.19 $Y2=-0.245
cc_417 N_A_654_392#_c_595_n N_RESET_B_c_703_n 0.00764716f $X=5.545 $Y=1.26 $X2=0
+ $Y2=0
cc_418 N_A_654_392#_c_605_n N_RESET_B_c_703_n 0.0218678f $X=5.49 $Y=1.765 $X2=0
+ $Y2=0
cc_419 N_A_654_392#_c_598_n N_RESET_B_c_703_n 0.00442103f $X=5.13 $Y=1.575 $X2=0
+ $Y2=0
cc_420 N_A_654_392#_c_604_n N_RESET_B_c_703_n 7.92081e-19 $X=5.13 $Y=1.465 $X2=0
+ $Y2=0
cc_421 N_A_654_392#_c_597_n RESET_B 0.0011065f $X=5.62 $Y=1.185 $X2=0 $Y2=0
cc_422 N_A_654_392#_c_605_n N_VPWR_c_743_n 0.00444645f $X=5.49 $Y=1.765 $X2=0
+ $Y2=0
cc_423 N_A_654_392#_c_605_n N_VPWR_c_736_n 0.00460931f $X=5.49 $Y=1.765 $X2=0
+ $Y2=0
cc_424 N_A_654_392#_c_605_n N_VPWR_c_747_n 0.00952195f $X=5.49 $Y=1.765 $X2=0
+ $Y2=0
cc_425 N_A_654_392#_c_597_n N_VGND_c_832_n 0.0033649f $X=5.62 $Y=1.185 $X2=0
+ $Y2=0
cc_426 N_A_654_392#_c_599_n N_VGND_c_832_n 0.00986285f $X=3.98 $Y=0.58 $X2=0
+ $Y2=0
cc_427 N_A_654_392#_c_600_n N_VGND_c_832_n 0.0255573f $X=4.9 $Y=0.935 $X2=0
+ $Y2=0
cc_428 N_A_654_392#_c_599_n N_VGND_c_834_n 0.0145482f $X=3.98 $Y=0.58 $X2=0
+ $Y2=0
cc_429 N_A_654_392#_c_597_n N_VGND_c_836_n 0.00360627f $X=5.62 $Y=1.185 $X2=0
+ $Y2=0
cc_430 N_A_654_392#_c_597_n N_VGND_c_840_n 0.00587514f $X=5.62 $Y=1.185 $X2=0
+ $Y2=0
cc_431 N_A_654_392#_c_599_n N_VGND_c_840_n 0.0119922f $X=3.98 $Y=0.58 $X2=0
+ $Y2=0
cc_432 N_A_654_392#_c_600_n N_VGND_c_840_n 0.0197026f $X=4.9 $Y=0.935 $X2=0
+ $Y2=0
cc_433 N_A_654_392#_c_599_n N_VGND_c_843_n 6.72815e-19 $X=3.98 $Y=0.58 $X2=0
+ $Y2=0
cc_434 N_RESET_B_c_703_n N_VPWR_c_739_n 0.0119374f $X=6.11 $Y=1.765 $X2=0 $Y2=0
cc_435 N_RESET_B_c_703_n N_VPWR_c_743_n 0.0049405f $X=6.11 $Y=1.765 $X2=0 $Y2=0
cc_436 N_RESET_B_c_703_n N_VPWR_c_736_n 0.00508379f $X=6.11 $Y=1.765 $X2=0 $Y2=0
cc_437 N_RESET_B_c_703_n N_VPWR_c_747_n 5.43541e-19 $X=6.11 $Y=1.765 $X2=0 $Y2=0
cc_438 N_RESET_B_c_703_n Q 9.71254e-19 $X=6.11 $Y=1.765 $X2=0 $Y2=0
cc_439 N_RESET_B_c_702_n N_VGND_c_833_n 0.00740995f $X=6.01 $Y=1.22 $X2=0 $Y2=0
cc_440 N_RESET_B_c_703_n N_VGND_c_833_n 6.53093e-19 $X=6.11 $Y=1.765 $X2=0 $Y2=0
cc_441 RESET_B N_VGND_c_833_n 0.00812328f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_442 N_RESET_B_c_702_n N_VGND_c_836_n 0.00461464f $X=6.01 $Y=1.22 $X2=0 $Y2=0
cc_443 N_RESET_B_c_702_n N_VGND_c_840_n 0.00909437f $X=6.01 $Y=1.22 $X2=0 $Y2=0
cc_444 N_VPWR_c_739_n Q 0.0357739f $X=6.42 $Y=2.145 $X2=0 $Y2=0
cc_445 N_VPWR_c_744_n Q 0.0159324f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_446 N_VPWR_c_736_n Q 0.0131546f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_447 N_Q_c_810_n N_VGND_c_833_n 0.00118878f $X=6.895 $Y=0.515 $X2=0 $Y2=0
cc_448 N_Q_c_810_n N_VGND_c_839_n 0.0170898f $X=6.895 $Y=0.515 $X2=0 $Y2=0
cc_449 N_Q_c_810_n N_VGND_c_840_n 0.0141455f $X=6.895 $Y=0.515 $X2=0 $Y2=0
