* File: sky130_fd_sc_ls__nand2b_2.pxi.spice
* Created: Fri Aug 28 13:32:47 2020
* 
x_PM_SKY130_FD_SC_LS__NAND2B_2%A_N N_A_N_M1008_g N_A_N_c_72_n N_A_N_M1006_g A_N
+ N_A_N_c_73_n PM_SKY130_FD_SC_LS__NAND2B_2%A_N
x_PM_SKY130_FD_SC_LS__NAND2B_2%A_27_74# N_A_27_74#_M1008_s N_A_27_74#_M1006_s
+ N_A_27_74#_c_99_n N_A_27_74#_c_100_n N_A_27_74#_c_114_n N_A_27_74#_M1000_g
+ N_A_27_74#_M1004_g N_A_27_74#_c_102_n N_A_27_74#_c_103_n N_A_27_74#_c_116_n
+ N_A_27_74#_M1007_g N_A_27_74#_M1009_g N_A_27_74#_c_105_n N_A_27_74#_c_106_n
+ N_A_27_74#_c_107_n N_A_27_74#_c_108_n N_A_27_74#_c_109_n N_A_27_74#_c_126_n
+ N_A_27_74#_c_110_n N_A_27_74#_c_111_n N_A_27_74#_c_118_n N_A_27_74#_c_112_n
+ PM_SKY130_FD_SC_LS__NAND2B_2%A_27_74#
x_PM_SKY130_FD_SC_LS__NAND2B_2%B N_B_c_202_n N_B_M1001_g N_B_M1002_g N_B_c_203_n
+ N_B_M1003_g N_B_M1005_g B N_B_c_200_n N_B_c_201_n
+ PM_SKY130_FD_SC_LS__NAND2B_2%B
x_PM_SKY130_FD_SC_LS__NAND2B_2%VPWR N_VPWR_M1006_d N_VPWR_M1007_d N_VPWR_M1003_s
+ N_VPWR_c_249_n N_VPWR_c_250_n N_VPWR_c_251_n N_VPWR_c_252_n N_VPWR_c_253_n
+ N_VPWR_c_254_n VPWR N_VPWR_c_255_n N_VPWR_c_256_n N_VPWR_c_257_n
+ N_VPWR_c_248_n PM_SKY130_FD_SC_LS__NAND2B_2%VPWR
x_PM_SKY130_FD_SC_LS__NAND2B_2%Y N_Y_M1004_d N_Y_M1000_s N_Y_M1001_d N_Y_c_299_n
+ N_Y_c_295_n N_Y_c_296_n N_Y_c_297_n N_Y_c_316_n Y Y
+ PM_SKY130_FD_SC_LS__NAND2B_2%Y
x_PM_SKY130_FD_SC_LS__NAND2B_2%VGND N_VGND_M1008_d N_VGND_M1002_d N_VGND_c_338_n
+ N_VGND_c_339_n VGND N_VGND_c_340_n N_VGND_c_341_n N_VGND_c_342_n
+ N_VGND_c_343_n N_VGND_c_344_n N_VGND_c_345_n PM_SKY130_FD_SC_LS__NAND2B_2%VGND
x_PM_SKY130_FD_SC_LS__NAND2B_2%A_242_74# N_A_242_74#_M1004_s N_A_242_74#_M1009_s
+ N_A_242_74#_M1005_s N_A_242_74#_c_378_n N_A_242_74#_c_379_n
+ N_A_242_74#_c_387_n N_A_242_74#_c_405_n N_A_242_74#_c_380_n
+ N_A_242_74#_c_381_n N_A_242_74#_c_409_n N_A_242_74#_c_382_n
+ N_A_242_74#_c_383_n N_A_242_74#_c_384_n N_A_242_74#_c_385_n
+ PM_SKY130_FD_SC_LS__NAND2B_2%A_242_74#
cc_1 VNB N_A_N_M1008_g 0.0408957f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.69
cc_2 VNB N_A_N_c_72_n 0.0308261f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_3 VNB N_A_N_c_73_n 0.0158471f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.515
cc_4 VNB N_A_27_74#_c_99_n 0.0240853f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.34
cc_5 VNB N_A_27_74#_c_100_n 0.0122346f $X=-0.19 $Y=-0.245 $X2=0.41 $Y2=1.515
cc_6 VNB N_A_27_74#_M1004_g 0.0237949f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.565
cc_7 VNB N_A_27_74#_c_102_n 0.00882279f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_27_74#_c_103_n 0.0103245f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_27_74#_M1009_g 0.0206469f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_27_74#_c_105_n 0.00593864f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_27_74#_c_106_n 0.00594687f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_74#_c_107_n 0.0277086f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_74#_c_108_n 0.0111309f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_74#_c_109_n 0.0102604f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_74#_c_110_n 0.0216805f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_27_74#_c_111_n 0.00301676f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_27_74#_c_112_n 0.0370399f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_B_M1002_g 0.02374f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.34
cc_19 VNB N_B_M1005_g 0.0284162f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.565
cc_20 VNB N_B_c_200_n 0.00107131f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_B_c_201_n 0.0386336f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VPWR_c_248_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_Y_c_295_n 0.00171224f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.565
cc_24 VNB N_Y_c_296_n 0.00541157f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_Y_c_297_n 6.45006e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB Y 0.00338874f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_338_n 0.0145875f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_339_n 0.00945073f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.565
cc_29 VNB N_VGND_c_340_n 0.0191515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_341_n 0.0419632f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_342_n 0.0196288f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_343_n 0.21982f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_344_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_345_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_242_74#_c_378_n 0.00386622f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.565
cc_36 VNB N_A_242_74#_c_379_n 0.00500698f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_242_74#_c_380_n 0.00403194f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_242_74#_c_381_n 0.00442536f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_242_74#_c_382_n 0.0259999f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_242_74#_c_383_n 0.0254393f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_242_74#_c_384_n 0.00270215f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_242_74#_c_385_n 0.0116965f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VPB N_A_N_c_72_n 0.0346343f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_44 VPB N_A_N_c_73_n 0.00796889f $X=-0.19 $Y=1.66 $X2=0.405 $Y2=1.515
cc_45 VPB N_A_27_74#_c_100_n 9.06264e-19 $X=-0.19 $Y=1.66 $X2=0.41 $Y2=1.515
cc_46 VPB N_A_27_74#_c_114_n 0.0241891f $X=-0.19 $Y=1.66 $X2=0.405 $Y2=1.515
cc_47 VPB N_A_27_74#_c_103_n 7.64781e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 VPB N_A_27_74#_c_116_n 0.0206347f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 VPB N_A_27_74#_c_111_n 0.00412606f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_A_27_74#_c_118_n 0.0389799f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_51 VPB N_B_c_202_n 0.0151507f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.35
cc_52 VPB N_B_c_203_n 0.0172531f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_53 VPB N_B_c_200_n 0.00284491f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_B_c_201_n 0.0205815f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_249_n 0.0155479f $X=-0.19 $Y=1.66 $X2=0.405 $Y2=1.515
cc_56 VPB N_VPWR_c_250_n 0.00329129f $X=-0.19 $Y=1.66 $X2=0.405 $Y2=1.565
cc_57 VPB N_VPWR_c_251_n 0.0120118f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_252_n 0.0190928f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_253_n 0.0231902f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_254_n 0.00709097f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_255_n 0.0290546f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_256_n 0.0177589f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_257_n 0.00601765f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_248_n 0.074124f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_Y_c_299_n 0.00365845f $X=-0.19 $Y=1.66 $X2=0.41 $Y2=1.515
cc_66 VPB Y 0.00271805f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_A_242_74#_c_379_n 0.00214346f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_A_242_74#_c_387_n 0.00721688f $X=-0.19 $Y=1.66 $X2=0.405 $Y2=1.565
cc_69 VPB N_A_242_74#_c_383_n 0.0272713f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 N_A_N_M1008_g N_A_27_74#_c_107_n 0.0131663f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_71 N_A_N_M1008_g N_A_27_74#_c_108_n 0.0123128f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_72 N_A_N_c_72_n N_A_27_74#_c_108_n 2.84881e-19 $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_73 N_A_N_c_73_n N_A_27_74#_c_108_n 0.00908651f $X=0.405 $Y=1.515 $X2=0 $Y2=0
cc_74 N_A_N_M1008_g N_A_27_74#_c_109_n 0.00417698f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_75 N_A_N_c_72_n N_A_27_74#_c_109_n 0.00419865f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_76 N_A_N_c_73_n N_A_27_74#_c_109_n 0.0278644f $X=0.405 $Y=1.515 $X2=0 $Y2=0
cc_77 N_A_N_c_72_n N_A_27_74#_c_126_n 0.0137387f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_78 N_A_N_c_73_n N_A_27_74#_c_126_n 0.00908651f $X=0.405 $Y=1.515 $X2=0 $Y2=0
cc_79 N_A_N_M1008_g N_A_27_74#_c_110_n 0.00111356f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_80 N_A_N_c_73_n N_A_27_74#_c_110_n 0.00710963f $X=0.405 $Y=1.515 $X2=0 $Y2=0
cc_81 N_A_N_c_72_n N_A_27_74#_c_111_n 0.00836613f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_82 N_A_N_c_73_n N_A_27_74#_c_111_n 0.01865f $X=0.405 $Y=1.515 $X2=0 $Y2=0
cc_83 N_A_N_c_72_n N_A_27_74#_c_118_n 0.0203471f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_84 N_A_N_c_73_n N_A_27_74#_c_118_n 0.0255992f $X=0.405 $Y=1.515 $X2=0 $Y2=0
cc_85 N_A_N_M1008_g N_A_27_74#_c_112_n 0.0178386f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_86 N_A_N_c_72_n N_VPWR_c_249_n 0.0166183f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_87 N_A_N_c_72_n N_VPWR_c_253_n 0.00481995f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_88 N_A_N_c_72_n N_VPWR_c_248_n 0.00508379f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_89 N_A_N_M1008_g N_VGND_c_338_n 0.00708561f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_90 N_A_N_M1008_g N_VGND_c_340_n 0.00434272f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_91 N_A_N_M1008_g N_VGND_c_343_n 0.00828717f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_92 N_A_N_M1008_g N_A_242_74#_c_378_n 0.00353982f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_93 N_A_27_74#_c_116_n N_B_c_202_n 0.04059f $X=1.955 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_94 N_A_27_74#_M1009_g N_B_M1002_g 0.0187832f $X=2 $Y=0.74 $X2=0 $Y2=0
cc_95 N_A_27_74#_c_103_n N_B_c_201_n 0.0119172f $X=1.955 $Y=1.675 $X2=0 $Y2=0
cc_96 N_A_27_74#_c_106_n N_B_c_201_n 0.00655909f $X=1.97 $Y=1.395 $X2=0 $Y2=0
cc_97 N_A_27_74#_c_126_n N_VPWR_M1006_d 0.016662f $X=0.805 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_98 N_A_27_74#_c_111_n N_VPWR_M1006_d 0.00367869f $X=0.89 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_99 N_A_27_74#_c_114_n N_VPWR_c_249_n 0.0187016f $X=1.505 $Y=1.765 $X2=0 $Y2=0
cc_100 N_A_27_74#_c_126_n N_VPWR_c_249_n 0.0216282f $X=0.805 $Y=2.035 $X2=0
+ $Y2=0
cc_101 N_A_27_74#_c_118_n N_VPWR_c_249_n 0.0304896f $X=0.28 $Y=2.115 $X2=0 $Y2=0
cc_102 N_A_27_74#_c_114_n N_VPWR_c_250_n 0.00181708f $X=1.505 $Y=1.765 $X2=0
+ $Y2=0
cc_103 N_A_27_74#_c_116_n N_VPWR_c_250_n 0.00886652f $X=1.955 $Y=1.765 $X2=0
+ $Y2=0
cc_104 N_A_27_74#_c_118_n N_VPWR_c_253_n 0.0097982f $X=0.28 $Y=2.115 $X2=0 $Y2=0
cc_105 N_A_27_74#_c_114_n N_VPWR_c_255_n 0.00461464f $X=1.505 $Y=1.765 $X2=0
+ $Y2=0
cc_106 N_A_27_74#_c_116_n N_VPWR_c_255_n 0.00413917f $X=1.955 $Y=1.765 $X2=0
+ $Y2=0
cc_107 N_A_27_74#_c_114_n N_VPWR_c_248_n 0.0045722f $X=1.505 $Y=1.765 $X2=0
+ $Y2=0
cc_108 N_A_27_74#_c_116_n N_VPWR_c_248_n 0.00403181f $X=1.955 $Y=1.765 $X2=0
+ $Y2=0
cc_109 N_A_27_74#_c_118_n N_VPWR_c_248_n 0.0111907f $X=0.28 $Y=2.115 $X2=0 $Y2=0
cc_110 N_A_27_74#_c_114_n N_Y_c_299_n 0.00149728f $X=1.505 $Y=1.765 $X2=0 $Y2=0
cc_111 N_A_27_74#_c_102_n N_Y_c_299_n 0.00213792f $X=1.865 $Y=1.395 $X2=0 $Y2=0
cc_112 N_A_27_74#_c_116_n N_Y_c_299_n 0.0162581f $X=1.955 $Y=1.765 $X2=0 $Y2=0
cc_113 N_A_27_74#_M1004_g N_Y_c_295_n 0.00122852f $X=1.57 $Y=0.74 $X2=0 $Y2=0
cc_114 N_A_27_74#_M1009_g N_Y_c_295_n 0.00296465f $X=2 $Y=0.74 $X2=0 $Y2=0
cc_115 N_A_27_74#_M1009_g N_Y_c_296_n 0.00903645f $X=2 $Y=0.74 $X2=0 $Y2=0
cc_116 N_A_27_74#_c_106_n N_Y_c_296_n 0.00560489f $X=1.97 $Y=1.395 $X2=0 $Y2=0
cc_117 N_A_27_74#_M1004_g N_Y_c_297_n 8.9081e-19 $X=1.57 $Y=0.74 $X2=0 $Y2=0
cc_118 N_A_27_74#_c_102_n N_Y_c_297_n 0.00760002f $X=1.865 $Y=1.395 $X2=0 $Y2=0
cc_119 N_A_27_74#_c_103_n Y 0.00415246f $X=1.955 $Y=1.675 $X2=0 $Y2=0
cc_120 N_A_27_74#_c_116_n Y 7.5187e-19 $X=1.955 $Y=1.765 $X2=0 $Y2=0
cc_121 N_A_27_74#_c_106_n Y 0.00367039f $X=1.97 $Y=1.395 $X2=0 $Y2=0
cc_122 N_A_27_74#_M1004_g N_VGND_c_338_n 0.00162304f $X=1.57 $Y=0.74 $X2=0 $Y2=0
cc_123 N_A_27_74#_c_107_n N_VGND_c_338_n 0.0191484f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_124 N_A_27_74#_c_108_n N_VGND_c_338_n 0.0150968f $X=0.805 $Y=1.095 $X2=0
+ $Y2=0
cc_125 N_A_27_74#_c_110_n N_VGND_c_338_n 0.00641171f $X=0.89 $Y=1.47 $X2=0 $Y2=0
cc_126 N_A_27_74#_c_112_n N_VGND_c_338_n 3.97306e-19 $X=0.97 $Y=1.305 $X2=0
+ $Y2=0
cc_127 N_A_27_74#_c_107_n N_VGND_c_340_n 0.0145639f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_128 N_A_27_74#_M1004_g N_VGND_c_341_n 0.00278247f $X=1.57 $Y=0.74 $X2=0 $Y2=0
cc_129 N_A_27_74#_M1009_g N_VGND_c_341_n 0.00278247f $X=2 $Y=0.74 $X2=0 $Y2=0
cc_130 N_A_27_74#_M1004_g N_VGND_c_343_n 0.00358425f $X=1.57 $Y=0.74 $X2=0 $Y2=0
cc_131 N_A_27_74#_M1009_g N_VGND_c_343_n 0.00353524f $X=2 $Y=0.74 $X2=0 $Y2=0
cc_132 N_A_27_74#_c_107_n N_VGND_c_343_n 0.0119984f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_133 N_A_27_74#_M1004_g N_A_242_74#_c_378_n 0.0053576f $X=1.57 $Y=0.74 $X2=0
+ $Y2=0
cc_134 N_A_27_74#_M1009_g N_A_242_74#_c_378_n 7.03865e-19 $X=2 $Y=0.74 $X2=0
+ $Y2=0
cc_135 N_A_27_74#_c_99_n N_A_242_74#_c_379_n 0.00877596f $X=1.415 $Y=1.395 $X2=0
+ $Y2=0
cc_136 N_A_27_74#_c_100_n N_A_242_74#_c_379_n 0.00766209f $X=1.505 $Y=1.675
+ $X2=0 $Y2=0
cc_137 N_A_27_74#_c_114_n N_A_242_74#_c_379_n 0.0225541f $X=1.505 $Y=1.765 $X2=0
+ $Y2=0
cc_138 N_A_27_74#_M1004_g N_A_242_74#_c_379_n 0.00360253f $X=1.57 $Y=0.74 $X2=0
+ $Y2=0
cc_139 N_A_27_74#_c_103_n N_A_242_74#_c_379_n 9.1341e-19 $X=1.955 $Y=1.675 $X2=0
+ $Y2=0
cc_140 N_A_27_74#_c_116_n N_A_242_74#_c_379_n 0.00114138f $X=1.955 $Y=1.765
+ $X2=0 $Y2=0
cc_141 N_A_27_74#_c_105_n N_A_242_74#_c_379_n 0.0055455f $X=1.53 $Y=1.395 $X2=0
+ $Y2=0
cc_142 N_A_27_74#_c_126_n N_A_242_74#_c_379_n 0.00847604f $X=0.805 $Y=2.035
+ $X2=0 $Y2=0
cc_143 N_A_27_74#_c_110_n N_A_242_74#_c_379_n 0.0313128f $X=0.89 $Y=1.47 $X2=0
+ $Y2=0
cc_144 N_A_27_74#_c_111_n N_A_242_74#_c_379_n 0.0224633f $X=0.89 $Y=1.95 $X2=0
+ $Y2=0
cc_145 N_A_27_74#_c_112_n N_A_242_74#_c_379_n 6.08793e-19 $X=0.97 $Y=1.305 $X2=0
+ $Y2=0
cc_146 N_A_27_74#_c_114_n N_A_242_74#_c_387_n 0.0106545f $X=1.505 $Y=1.765 $X2=0
+ $Y2=0
cc_147 N_A_27_74#_c_116_n N_A_242_74#_c_387_n 0.0117527f $X=1.955 $Y=1.765 $X2=0
+ $Y2=0
cc_148 N_A_27_74#_c_114_n N_A_242_74#_c_405_n 0.00470556f $X=1.505 $Y=1.765
+ $X2=0 $Y2=0
cc_149 N_A_27_74#_M1004_g N_A_242_74#_c_380_n 0.0100711f $X=1.57 $Y=0.74 $X2=0
+ $Y2=0
cc_150 N_A_27_74#_M1009_g N_A_242_74#_c_380_n 0.0119194f $X=2 $Y=0.74 $X2=0
+ $Y2=0
cc_151 N_A_27_74#_M1004_g N_A_242_74#_c_381_n 0.00281658f $X=1.57 $Y=0.74 $X2=0
+ $Y2=0
cc_152 N_A_27_74#_M1004_g N_A_242_74#_c_409_n 7.28037e-19 $X=1.57 $Y=0.74 $X2=0
+ $Y2=0
cc_153 N_A_27_74#_M1009_g N_A_242_74#_c_409_n 0.00893796f $X=2 $Y=0.74 $X2=0
+ $Y2=0
cc_154 N_A_27_74#_c_99_n N_A_242_74#_c_384_n 0.00386604f $X=1.415 $Y=1.395 $X2=0
+ $Y2=0
cc_155 N_A_27_74#_M1004_g N_A_242_74#_c_384_n 0.00290614f $X=1.57 $Y=0.74 $X2=0
+ $Y2=0
cc_156 N_B_c_202_n N_VPWR_c_250_n 0.00871578f $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_157 N_B_c_203_n N_VPWR_c_250_n 0.00112373f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_158 N_B_c_202_n N_VPWR_c_252_n 0.00112373f $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_159 N_B_c_203_n N_VPWR_c_252_n 0.00974588f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_160 N_B_c_202_n N_VPWR_c_256_n 0.00413917f $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_161 N_B_c_203_n N_VPWR_c_256_n 0.00413917f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_162 N_B_c_202_n N_VPWR_c_248_n 0.00403181f $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_163 N_B_c_203_n N_VPWR_c_248_n 0.00403181f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_164 N_B_M1002_g N_Y_c_296_n 0.0038121f $X=2.43 $Y=0.74 $X2=0 $Y2=0
cc_165 N_B_c_200_n N_Y_c_296_n 0.00332636f $X=2.61 $Y=1.515 $X2=0 $Y2=0
cc_166 N_B_c_201_n N_Y_c_296_n 3.62014e-19 $X=2.855 $Y=1.557 $X2=0 $Y2=0
cc_167 N_B_c_202_n N_Y_c_316_n 0.0143919f $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_168 N_B_c_203_n N_Y_c_316_n 0.00403377f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_169 N_B_c_200_n N_Y_c_316_n 0.0225186f $X=2.61 $Y=1.515 $X2=0 $Y2=0
cc_170 N_B_c_201_n N_Y_c_316_n 0.00133815f $X=2.855 $Y=1.557 $X2=0 $Y2=0
cc_171 N_B_c_202_n Y 0.00110805f $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_172 N_B_c_200_n Y 0.0299194f $X=2.61 $Y=1.515 $X2=0 $Y2=0
cc_173 N_B_c_201_n Y 0.00316826f $X=2.855 $Y=1.557 $X2=0 $Y2=0
cc_174 N_B_c_202_n Y 0.00108874f $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_175 N_B_M1002_g N_VGND_c_339_n 0.00188034f $X=2.43 $Y=0.74 $X2=0 $Y2=0
cc_176 N_B_M1005_g N_VGND_c_339_n 0.00533745f $X=2.865 $Y=0.74 $X2=0 $Y2=0
cc_177 N_B_c_200_n N_VGND_c_339_n 0.0119403f $X=2.61 $Y=1.515 $X2=0 $Y2=0
cc_178 N_B_c_201_n N_VGND_c_339_n 8.04984e-19 $X=2.855 $Y=1.557 $X2=0 $Y2=0
cc_179 N_B_M1002_g N_VGND_c_341_n 0.00430908f $X=2.43 $Y=0.74 $X2=0 $Y2=0
cc_180 N_B_M1005_g N_VGND_c_342_n 0.00434272f $X=2.865 $Y=0.74 $X2=0 $Y2=0
cc_181 N_B_M1002_g N_VGND_c_343_n 0.0081583f $X=2.43 $Y=0.74 $X2=0 $Y2=0
cc_182 N_B_M1005_g N_VGND_c_343_n 0.00824104f $X=2.865 $Y=0.74 $X2=0 $Y2=0
cc_183 N_B_c_202_n N_A_242_74#_c_387_n 0.0118038f $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_184 N_B_c_203_n N_A_242_74#_c_387_n 0.0172709f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_185 N_B_M1002_g N_A_242_74#_c_380_n 0.00323029f $X=2.43 $Y=0.74 $X2=0 $Y2=0
cc_186 N_B_M1002_g N_A_242_74#_c_409_n 0.00835413f $X=2.43 $Y=0.74 $X2=0 $Y2=0
cc_187 N_B_M1005_g N_A_242_74#_c_382_n 0.00826065f $X=2.865 $Y=0.74 $X2=0 $Y2=0
cc_188 N_B_c_203_n N_A_242_74#_c_383_n 0.0175143f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_189 N_B_M1005_g N_A_242_74#_c_383_n 0.00778767f $X=2.865 $Y=0.74 $X2=0 $Y2=0
cc_190 N_B_c_200_n N_A_242_74#_c_383_n 0.021203f $X=2.61 $Y=1.515 $X2=0 $Y2=0
cc_191 N_B_c_201_n N_A_242_74#_c_383_n 0.0112879f $X=2.855 $Y=1.557 $X2=0 $Y2=0
cc_192 N_B_M1005_g N_A_242_74#_c_385_n 0.00333567f $X=2.865 $Y=0.74 $X2=0 $Y2=0
cc_193 N_B_c_201_n N_A_242_74#_c_385_n 2.15716e-19 $X=2.855 $Y=1.557 $X2=0 $Y2=0
cc_194 N_VPWR_M1007_d Y 0.00206339f $X=2.03 $Y=1.84 $X2=0 $Y2=0
cc_195 N_VPWR_M1006_d N_A_242_74#_c_379_n 0.0114702f $X=0.58 $Y=1.84 $X2=0 $Y2=0
cc_196 N_VPWR_c_249_n N_A_242_74#_c_379_n 0.00524486f $X=0.915 $Y=2.405 $X2=0
+ $Y2=0
cc_197 N_VPWR_M1007_d N_A_242_74#_c_387_n 0.00391935f $X=2.03 $Y=1.84 $X2=0
+ $Y2=0
cc_198 N_VPWR_M1003_s N_A_242_74#_c_387_n 0.00692961f $X=2.93 $Y=1.84 $X2=0
+ $Y2=0
cc_199 N_VPWR_c_250_n N_A_242_74#_c_387_n 0.0167754f $X=2.18 $Y=2.805 $X2=0
+ $Y2=0
cc_200 N_VPWR_c_252_n N_A_242_74#_c_387_n 0.0228134f $X=3.08 $Y=2.805 $X2=0
+ $Y2=0
cc_201 N_VPWR_c_248_n N_A_242_74#_c_387_n 0.0387921f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_202 N_VPWR_M1006_d N_A_242_74#_c_405_n 0.00359043f $X=0.58 $Y=1.84 $X2=0
+ $Y2=0
cc_203 N_VPWR_c_249_n N_A_242_74#_c_405_n 0.0124718f $X=0.915 $Y=2.405 $X2=0
+ $Y2=0
cc_204 N_VPWR_c_248_n N_A_242_74#_c_405_n 0.00661702f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_205 N_VPWR_M1003_s N_A_242_74#_c_383_n 0.00974914f $X=2.93 $Y=1.84 $X2=0
+ $Y2=0
cc_206 N_Y_c_299_n N_A_242_74#_c_379_n 0.0298028f $X=2.045 $Y=2.01 $X2=0 $Y2=0
cc_207 N_Y_c_295_n N_A_242_74#_c_379_n 0.0067072f $X=1.785 $Y=0.825 $X2=0 $Y2=0
cc_208 N_Y_c_297_n N_A_242_74#_c_379_n 0.0110286f $X=1.87 $Y=1.305 $X2=0 $Y2=0
cc_209 Y N_A_242_74#_c_379_n 0.0122293f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_210 N_Y_M1000_s N_A_242_74#_c_387_n 0.00578049f $X=1.58 $Y=1.84 $X2=0 $Y2=0
cc_211 N_Y_M1001_d N_A_242_74#_c_387_n 0.00542821f $X=2.48 $Y=1.84 $X2=0 $Y2=0
cc_212 N_Y_c_299_n N_A_242_74#_c_387_n 0.0245513f $X=2.045 $Y=2.01 $X2=0 $Y2=0
cc_213 N_Y_c_316_n N_A_242_74#_c_387_n 0.0253647f $X=2.63 $Y=2.115 $X2=0 $Y2=0
cc_214 Y N_A_242_74#_c_387_n 0.0151327f $X=2.075 $Y=1.95 $X2=0 $Y2=0
cc_215 N_Y_M1004_d N_A_242_74#_c_380_n 0.00191292f $X=1.645 $Y=0.37 $X2=0 $Y2=0
cc_216 N_Y_c_295_n N_A_242_74#_c_380_n 0.0107548f $X=1.785 $Y=0.825 $X2=0 $Y2=0
cc_217 N_Y_c_296_n N_A_242_74#_c_409_n 0.0178056f $X=2.045 $Y=1.305 $X2=0 $Y2=0
cc_218 N_Y_c_316_n N_A_242_74#_c_383_n 0.0132513f $X=2.63 $Y=2.115 $X2=0 $Y2=0
cc_219 N_VGND_c_338_n N_A_242_74#_c_378_n 0.0220879f $X=0.71 $Y=0.675 $X2=0
+ $Y2=0
cc_220 N_VGND_c_339_n N_A_242_74#_c_380_n 0.010974f $X=2.645 $Y=0.515 $X2=0
+ $Y2=0
cc_221 N_VGND_c_341_n N_A_242_74#_c_380_n 0.0568424f $X=2.56 $Y=0 $X2=0 $Y2=0
cc_222 N_VGND_c_343_n N_A_242_74#_c_380_n 0.0313831f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_223 N_VGND_c_338_n N_A_242_74#_c_381_n 0.00962616f $X=0.71 $Y=0.675 $X2=0
+ $Y2=0
cc_224 N_VGND_c_341_n N_A_242_74#_c_381_n 0.0236115f $X=2.56 $Y=0 $X2=0 $Y2=0
cc_225 N_VGND_c_343_n N_A_242_74#_c_381_n 0.0127234f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_226 N_VGND_c_339_n N_A_242_74#_c_382_n 0.053968f $X=2.645 $Y=0.515 $X2=0
+ $Y2=0
cc_227 N_VGND_c_342_n N_A_242_74#_c_382_n 0.0145639f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_228 N_VGND_c_343_n N_A_242_74#_c_382_n 0.0119984f $X=3.12 $Y=0 $X2=0 $Y2=0
