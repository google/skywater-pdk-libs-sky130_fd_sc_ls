* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__nor3b_4 A B C_N VGND VNB VPB VPWR Y
X0 VGND C_N a_468_264# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X1 a_27_368# B a_126_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X2 VGND B Y VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X3 a_27_368# a_468_264# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X4 VPWR A a_126_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X5 Y B VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X7 a_126_368# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X8 a_27_368# B a_126_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X9 a_27_368# a_468_264# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X10 a_126_368# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X11 a_468_264# C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X12 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X13 VGND a_468_264# Y VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X14 a_126_368# B a_27_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X15 Y a_468_264# a_27_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X16 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X17 Y a_468_264# a_27_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X18 a_126_368# B a_27_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X19 VPWR A a_126_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X20 Y B VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X21 Y a_468_264# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X22 VPWR C_N a_468_264# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X23 VGND a_468_264# Y VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X24 Y a_468_264# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X25 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X26 VGND B Y VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
.ends
