* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
X0 a_602_392# B1 a_517_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 VPWR A2 a_517_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 VGND C1 a_105_280# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X3 VGND a_105_280# X VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X4 X a_105_280# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X5 a_105_280# C1 VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X6 a_105_280# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X7 VGND a_105_280# X VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X8 X a_105_280# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X9 a_105_280# C1 a_602_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 X a_105_280# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X11 a_1064_123# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X12 X a_105_280# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X13 VPWR a_105_280# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X14 VGND A2 a_1064_123# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X15 a_105_280# A1 a_1064_123# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X16 a_517_392# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X17 a_517_392# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X18 a_517_392# B1 a_602_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 VPWR A1 a_517_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X20 a_1064_123# A1 a_105_280# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X21 VGND B1 a_105_280# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X22 VPWR a_105_280# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X23 a_602_392# C1 a_105_280# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends
