* File: sky130_fd_sc_ls__a222o_1.pxi.spice
* Created: Wed Sep  2 10:49:46 2020
* 
x_PM_SKY130_FD_SC_LS__A222O_1%C1 N_C1_c_85_n N_C1_c_90_n N_C1_M1009_g
+ N_C1_M1006_g C1 C1 N_C1_c_86_n N_C1_c_87_n N_C1_c_88_n
+ PM_SKY130_FD_SC_LS__A222O_1%C1
x_PM_SKY130_FD_SC_LS__A222O_1%C2 N_C2_c_115_n N_C2_M1013_g N_C2_c_116_n
+ N_C2_c_120_n N_C2_M1011_g C2 N_C2_c_118_n PM_SKY130_FD_SC_LS__A222O_1%C2
x_PM_SKY130_FD_SC_LS__A222O_1%B2 N_B2_c_162_n N_B2_M1012_g N_B2_c_158_n
+ N_B2_M1007_g N_B2_c_164_n B2 N_B2_c_161_n PM_SKY130_FD_SC_LS__A222O_1%B2
x_PM_SKY130_FD_SC_LS__A222O_1%B1 N_B1_M1002_g N_B1_M1008_g N_B1_c_207_n
+ N_B1_c_212_n B1 B1 N_B1_c_208_n N_B1_c_209_n N_B1_c_210_n
+ PM_SKY130_FD_SC_LS__A222O_1%B1
x_PM_SKY130_FD_SC_LS__A222O_1%A1 N_A1_M1004_g N_A1_c_249_n N_A1_c_254_n
+ N_A1_M1003_g N_A1_c_255_n A1 N_A1_c_251_n N_A1_c_252_n
+ PM_SKY130_FD_SC_LS__A222O_1%A1
x_PM_SKY130_FD_SC_LS__A222O_1%A2 N_A2_M1001_g N_A2_c_287_n N_A2_c_292_n
+ N_A2_M1010_g A2 N_A2_c_289_n N_A2_c_290_n PM_SKY130_FD_SC_LS__A222O_1%A2
x_PM_SKY130_FD_SC_LS__A222O_1%A_32_74# N_A_32_74#_M1006_s N_A_32_74#_M1008_d
+ N_A_32_74#_M1009_d N_A_32_74#_c_328_n N_A_32_74#_M1005_g N_A_32_74#_M1000_g
+ N_A_32_74#_c_330_n N_A_32_74#_c_340_n N_A_32_74#_c_331_n N_A_32_74#_c_337_n
+ N_A_32_74#_c_367_n N_A_32_74#_c_332_n N_A_32_74#_c_351_n N_A_32_74#_c_333_n
+ N_A_32_74#_c_356_n N_A_32_74#_c_334_n N_A_32_74#_c_335_n
+ PM_SKY130_FD_SC_LS__A222O_1%A_32_74#
x_PM_SKY130_FD_SC_LS__A222O_1%A_27_390# N_A_27_390#_M1009_s N_A_27_390#_M1011_d
+ N_A_27_390#_M1002_d N_A_27_390#_c_431_n N_A_27_390#_c_432_n
+ N_A_27_390#_c_433_n N_A_27_390#_c_434_n N_A_27_390#_c_435_n
+ N_A_27_390#_c_436_n N_A_27_390#_c_437_n PM_SKY130_FD_SC_LS__A222O_1%A_27_390#
x_PM_SKY130_FD_SC_LS__A222O_1%A_337_390# N_A_337_390#_M1012_d
+ N_A_337_390#_M1003_d N_A_337_390#_c_476_n N_A_337_390#_c_477_n
+ N_A_337_390#_c_478_n N_A_337_390#_c_479_n
+ PM_SKY130_FD_SC_LS__A222O_1%A_337_390#
x_PM_SKY130_FD_SC_LS__A222O_1%VPWR N_VPWR_M1003_s N_VPWR_M1010_d N_VPWR_c_513_n
+ N_VPWR_c_514_n N_VPWR_c_515_n N_VPWR_c_516_n VPWR N_VPWR_c_517_n
+ N_VPWR_c_518_n N_VPWR_c_512_n N_VPWR_c_520_n PM_SKY130_FD_SC_LS__A222O_1%VPWR
x_PM_SKY130_FD_SC_LS__A222O_1%X N_X_M1000_d N_X_M1005_d N_X_c_560_n N_X_c_561_n
+ X X X X N_X_c_562_n PM_SKY130_FD_SC_LS__A222O_1%X
x_PM_SKY130_FD_SC_LS__A222O_1%VGND N_VGND_M1013_d N_VGND_M1001_d VGND
+ N_VGND_c_588_n N_VGND_c_589_n N_VGND_c_590_n N_VGND_c_591_n N_VGND_c_592_n
+ PM_SKY130_FD_SC_LS__A222O_1%VGND
cc_1 VNB N_C1_c_85_n 0.014917f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.785
cc_2 VNB N_C1_c_86_n 0.0415775f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.285
cc_3 VNB N_C1_c_87_n 0.0243057f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.285
cc_4 VNB N_C1_c_88_n 0.0238394f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.12
cc_5 VNB N_C2_c_115_n 0.0211034f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.45
cc_6 VNB N_C2_c_116_n 0.0126102f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.45
cc_7 VNB C2 0.00372322f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_8 VNB N_C2_c_118_n 0.0473823f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_B2_c_158_n 0.00756866f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.45
cc_10 VNB N_B2_M1007_g 0.0250785f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.69
cc_11 VNB B2 0.00699165f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_B2_c_161_n 0.0286499f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.285
cc_13 VNB N_B1_c_207_n 0.0136647f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_14 VNB N_B1_c_208_n 0.0401895f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.12
cc_15 VNB N_B1_c_209_n 0.00896147f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.45
cc_16 VNB N_B1_c_210_n 0.0235135f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.285
cc_17 VNB N_A1_c_249_n 0.0130874f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.45
cc_18 VNB A1 0.00802928f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.285
cc_19 VNB N_A1_c_251_n 0.0303908f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.12
cc_20 VNB N_A1_c_252_n 0.0235136f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.285
cc_21 VNB N_A2_c_287_n 0.0114015f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.45
cc_22 VNB A2 0.00857517f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_23 VNB N_A2_c_289_n 0.0290381f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A2_c_290_n 0.0188217f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.285
cc_25 VNB N_A_32_74#_c_328_n 0.0370482f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_26 VNB N_A_32_74#_M1000_g 0.0292321f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.285
cc_27 VNB N_A_32_74#_c_330_n 0.0189692f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_32_74#_c_331_n 0.00721971f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.665
cc_29 VNB N_A_32_74#_c_332_n 0.00282281f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_32_74#_c_333_n 0.00768644f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_32_74#_c_334_n 0.00712101f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_32_74#_c_335_n 0.00281093f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VPWR_c_512_n 0.203486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_X_c_560_n 0.0265168f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_35 VNB N_X_c_561_n 0.0133911f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.285
cc_36 VNB N_X_c_562_n 0.0247034f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_588_n 0.0703162f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.285
cc_38 VNB N_VGND_c_589_n 0.0189863f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_590_n 0.271043f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_591_n 0.0299712f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_592_n 0.0244424f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VPB N_C1_c_85_n 0.00885027f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.785
cc_43 VPB N_C1_c_90_n 0.0279981f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.875
cc_44 VPB N_C1_c_87_n 0.00822918f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.285
cc_45 VPB N_C2_c_116_n 0.00737721f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.45
cc_46 VPB N_C2_c_120_n 0.021942f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.12
cc_47 VPB C2 0.00305182f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_48 VPB N_B2_c_162_n 0.0149731f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.45
cc_49 VPB N_B2_c_158_n 0.0014731f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.45
cc_50 VPB N_B2_c_164_n 0.0184489f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_51 VPB B2 0.00262299f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_B1_c_207_n 0.0086808f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_53 VPB N_B1_c_212_n 0.0273095f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_54 VPB N_B1_c_209_n 0.00739206f $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.45
cc_55 VPB N_A1_c_249_n 0.0018398f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.45
cc_56 VPB N_A1_c_254_n 0.0172824f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.12
cc_57 VPB N_A1_c_255_n 0.0193789f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_A2_c_287_n 0.00559538f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.45
cc_59 VPB N_A2_c_292_n 0.0227094f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.12
cc_60 VPB N_A_32_74#_c_328_n 0.0297366f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_61 VPB N_A_32_74#_c_337_n 0.00272263f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_A_32_74#_c_333_n 0.00558651f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_A_27_390#_c_431_n 0.0363365f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_A_27_390#_c_432_n 0.00391743f $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.12
cc_65 VPB N_A_27_390#_c_433_n 0.0098742f $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.45
cc_66 VPB N_A_27_390#_c_434_n 0.00684298f $X=-0.19 $Y=1.66 $X2=0.337 $Y2=1.295
cc_67 VPB N_A_27_390#_c_435_n 0.00794963f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_A_27_390#_c_436_n 0.00565834f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_A_27_390#_c_437_n 0.0022931f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_A_337_390#_c_476_n 0.0146376f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_71 VPB N_A_337_390#_c_477_n 0.00705207f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_A_337_390#_c_478_n 0.00277636f $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.285
cc_73 VPB N_A_337_390#_c_479_n 0.0067323f $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.12
cc_74 VPB N_VPWR_c_513_n 0.017915f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_75 VPB N_VPWR_c_514_n 0.015585f $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.285
cc_76 VPB N_VPWR_c_515_n 0.0679823f $X=-0.19 $Y=1.66 $X2=0.337 $Y2=1.285
cc_77 VPB N_VPWR_c_516_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_517_n 0.0200251f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_518_n 0.0189562f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_512_n 0.0912132f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_520_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 VPB X 0.0135031f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.285
cc_83 VPB X 0.0415177f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_84 VPB N_X_c_562_n 0.00775552f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 N_C1_c_88_n N_C2_c_115_n 0.0266007f $X=0.407 $Y=1.12 $X2=-0.19 $Y2=-0.245
cc_86 N_C1_c_85_n N_C2_c_116_n 0.00407741f $X=0.505 $Y=1.785 $X2=0 $Y2=0
cc_87 N_C1_c_90_n N_C2_c_120_n 0.0207527f $X=0.505 $Y=1.875 $X2=0 $Y2=0
cc_88 N_C1_c_86_n N_C2_c_118_n 0.0306781f $X=0.385 $Y=1.285 $X2=0 $Y2=0
cc_89 N_C1_c_88_n N_A_32_74#_c_330_n 0.00793201f $X=0.407 $Y=1.12 $X2=0 $Y2=0
cc_90 N_C1_c_87_n N_A_32_74#_c_340_n 0.0059763f $X=0.385 $Y=1.285 $X2=0 $Y2=0
cc_91 N_C1_c_88_n N_A_32_74#_c_340_n 0.00946381f $X=0.407 $Y=1.12 $X2=0 $Y2=0
cc_92 N_C1_c_86_n N_A_32_74#_c_331_n 0.00158451f $X=0.385 $Y=1.285 $X2=0 $Y2=0
cc_93 N_C1_c_87_n N_A_32_74#_c_331_n 0.026304f $X=0.385 $Y=1.285 $X2=0 $Y2=0
cc_94 N_C1_c_88_n N_A_32_74#_c_331_n 7.14797e-19 $X=0.407 $Y=1.12 $X2=0 $Y2=0
cc_95 N_C1_c_90_n N_A_32_74#_c_333_n 0.00946312f $X=0.505 $Y=1.875 $X2=0 $Y2=0
cc_96 N_C1_c_87_n N_A_32_74#_c_333_n 0.0512661f $X=0.385 $Y=1.285 $X2=0 $Y2=0
cc_97 N_C1_c_88_n N_A_32_74#_c_333_n 0.0108286f $X=0.407 $Y=1.12 $X2=0 $Y2=0
cc_98 N_C1_c_90_n N_A_27_390#_c_431_n 0.0130457f $X=0.505 $Y=1.875 $X2=0 $Y2=0
cc_99 N_C1_c_86_n N_A_27_390#_c_431_n 6.85165e-19 $X=0.385 $Y=1.285 $X2=0 $Y2=0
cc_100 N_C1_c_87_n N_A_27_390#_c_431_n 0.026435f $X=0.385 $Y=1.285 $X2=0 $Y2=0
cc_101 N_C1_c_90_n N_A_27_390#_c_432_n 0.0114648f $X=0.505 $Y=1.875 $X2=0 $Y2=0
cc_102 N_C1_c_90_n N_A_27_390#_c_433_n 0.00282905f $X=0.505 $Y=1.875 $X2=0 $Y2=0
cc_103 N_C1_c_90_n N_VPWR_c_515_n 0.00390694f $X=0.505 $Y=1.875 $X2=0 $Y2=0
cc_104 N_C1_c_90_n N_VPWR_c_512_n 0.00542671f $X=0.505 $Y=1.875 $X2=0 $Y2=0
cc_105 N_C1_c_88_n N_VGND_c_590_n 0.00437003f $X=0.407 $Y=1.12 $X2=0 $Y2=0
cc_106 N_C1_c_88_n N_VGND_c_591_n 0.00434272f $X=0.407 $Y=1.12 $X2=0 $Y2=0
cc_107 N_C1_c_88_n N_VGND_c_592_n 0.00126064f $X=0.407 $Y=1.12 $X2=0 $Y2=0
cc_108 N_C2_c_120_n N_B2_c_162_n 0.0197621f $X=1.11 $Y=1.875 $X2=-0.19
+ $Y2=-0.245
cc_109 C2 N_B2_M1007_g 3.3883e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_110 N_C2_c_118_n N_B2_M1007_g 0.0016358f $X=1.11 $Y=1.285 $X2=0 $Y2=0
cc_111 N_C2_c_116_n N_B2_c_164_n 0.00734891f $X=1.11 $Y=1.785 $X2=0 $Y2=0
cc_112 C2 N_B2_c_164_n 5.04794e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_113 N_C2_c_116_n B2 6.69477e-19 $X=1.11 $Y=1.785 $X2=0 $Y2=0
cc_114 C2 B2 0.0465362f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_115 N_C2_c_118_n B2 9.0494e-19 $X=1.11 $Y=1.285 $X2=0 $Y2=0
cc_116 N_C2_c_116_n N_B2_c_161_n 0.0066094f $X=1.11 $Y=1.785 $X2=0 $Y2=0
cc_117 C2 N_B2_c_161_n 0.00116331f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_118 N_C2_c_118_n N_B2_c_161_n 0.0175466f $X=1.11 $Y=1.285 $X2=0 $Y2=0
cc_119 N_C2_c_115_n N_A_32_74#_c_330_n 0.00159871f $X=0.91 $Y=1.12 $X2=0 $Y2=0
cc_120 N_C2_c_120_n N_A_32_74#_c_337_n 0.0108705f $X=1.11 $Y=1.875 $X2=0 $Y2=0
cc_121 N_C2_c_118_n N_A_32_74#_c_337_n 0.00364036f $X=1.11 $Y=1.285 $X2=0 $Y2=0
cc_122 N_C2_c_115_n N_A_32_74#_c_351_n 0.0040045f $X=0.91 $Y=1.12 $X2=0 $Y2=0
cc_123 N_C2_c_115_n N_A_32_74#_c_333_n 0.00811889f $X=0.91 $Y=1.12 $X2=0 $Y2=0
cc_124 N_C2_c_120_n N_A_32_74#_c_333_n 0.00124989f $X=1.11 $Y=1.875 $X2=0 $Y2=0
cc_125 C2 N_A_32_74#_c_333_n 0.0475893f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_126 N_C2_c_118_n N_A_32_74#_c_333_n 0.0116709f $X=1.11 $Y=1.285 $X2=0 $Y2=0
cc_127 N_C2_c_115_n N_A_32_74#_c_356_n 0.0111662f $X=0.91 $Y=1.12 $X2=0 $Y2=0
cc_128 C2 N_A_32_74#_c_356_n 0.0256857f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_129 N_C2_c_118_n N_A_32_74#_c_356_n 0.00982054f $X=1.11 $Y=1.285 $X2=0 $Y2=0
cc_130 N_C2_c_120_n N_A_27_390#_c_431_n 9.29186e-19 $X=1.11 $Y=1.875 $X2=0 $Y2=0
cc_131 N_C2_c_120_n N_A_27_390#_c_432_n 0.0144113f $X=1.11 $Y=1.875 $X2=0 $Y2=0
cc_132 N_C2_c_120_n N_A_27_390#_c_434_n 0.00525241f $X=1.11 $Y=1.875 $X2=0 $Y2=0
cc_133 C2 N_A_27_390#_c_434_n 0.0156932f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_134 N_C2_c_118_n N_A_27_390#_c_434_n 6.89403e-19 $X=1.11 $Y=1.285 $X2=0 $Y2=0
cc_135 N_C2_c_120_n N_VPWR_c_515_n 0.00390708f $X=1.11 $Y=1.875 $X2=0 $Y2=0
cc_136 N_C2_c_120_n N_VPWR_c_512_n 0.00542671f $X=1.11 $Y=1.875 $X2=0 $Y2=0
cc_137 N_C2_c_115_n N_VGND_c_590_n 0.00369441f $X=0.91 $Y=1.12 $X2=0 $Y2=0
cc_138 N_C2_c_115_n N_VGND_c_591_n 0.00383152f $X=0.91 $Y=1.12 $X2=0 $Y2=0
cc_139 N_C2_c_115_n N_VGND_c_592_n 0.0102512f $X=0.91 $Y=1.12 $X2=0 $Y2=0
cc_140 N_B2_c_158_n N_B1_c_207_n 0.00738059f $X=1.675 $Y=1.69 $X2=0 $Y2=0
cc_141 B2 N_B1_c_207_n 0.00200975f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_142 N_B2_c_161_n N_B1_c_207_n 0.012376f $X=1.765 $Y=1.345 $X2=0 $Y2=0
cc_143 N_B2_c_162_n N_B1_c_212_n 0.0248509f $X=1.61 $Y=1.875 $X2=0 $Y2=0
cc_144 N_B2_c_164_n N_B1_c_212_n 0.00327331f $X=1.61 $Y=1.782 $X2=0 $Y2=0
cc_145 N_B2_M1007_g N_B1_c_208_n 0.012376f $X=1.855 $Y=0.69 $X2=0 $Y2=0
cc_146 B2 N_B1_c_208_n 0.00122615f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_147 N_B2_c_158_n N_B1_c_209_n 2.23407e-19 $X=1.675 $Y=1.69 $X2=0 $Y2=0
cc_148 N_B2_M1007_g N_B1_c_209_n 3.3231e-19 $X=1.855 $Y=0.69 $X2=0 $Y2=0
cc_149 B2 N_B1_c_209_n 0.0307418f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_150 N_B2_c_161_n N_B1_c_209_n 3.65571e-19 $X=1.765 $Y=1.345 $X2=0 $Y2=0
cc_151 N_B2_M1007_g N_B1_c_210_n 0.0467273f $X=1.855 $Y=0.69 $X2=0 $Y2=0
cc_152 N_B2_M1007_g N_A_32_74#_c_356_n 0.0136055f $X=1.855 $Y=0.69 $X2=0 $Y2=0
cc_153 B2 N_A_32_74#_c_356_n 0.0204678f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_154 N_B2_c_161_n N_A_32_74#_c_356_n 0.00425903f $X=1.765 $Y=1.345 $X2=0 $Y2=0
cc_155 N_B2_M1007_g N_A_32_74#_c_334_n 0.0016437f $X=1.855 $Y=0.69 $X2=0 $Y2=0
cc_156 N_B2_c_162_n N_A_27_390#_c_434_n 0.0120044f $X=1.61 $Y=1.875 $X2=0 $Y2=0
cc_157 N_B2_c_164_n N_A_27_390#_c_434_n 7.1313e-19 $X=1.61 $Y=1.782 $X2=0 $Y2=0
cc_158 N_B2_c_162_n N_A_27_390#_c_435_n 0.0114074f $X=1.61 $Y=1.875 $X2=0 $Y2=0
cc_159 N_B2_c_162_n N_A_27_390#_c_436_n 8.51498e-19 $X=1.61 $Y=1.875 $X2=0 $Y2=0
cc_160 N_B2_c_162_n N_A_27_390#_c_437_n 0.00203163f $X=1.61 $Y=1.875 $X2=0 $Y2=0
cc_161 N_B2_c_162_n N_A_337_390#_c_479_n 0.00135425f $X=1.61 $Y=1.875 $X2=0
+ $Y2=0
cc_162 N_B2_c_164_n N_A_337_390#_c_479_n 8.838e-19 $X=1.61 $Y=1.782 $X2=0 $Y2=0
cc_163 B2 N_A_337_390#_c_479_n 0.0192235f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_164 N_B2_c_161_n N_A_337_390#_c_479_n 8.10809e-19 $X=1.765 $Y=1.345 $X2=0
+ $Y2=0
cc_165 N_B2_c_162_n N_VPWR_c_515_n 0.00390694f $X=1.61 $Y=1.875 $X2=0 $Y2=0
cc_166 N_B2_c_162_n N_VPWR_c_512_n 0.00542671f $X=1.61 $Y=1.875 $X2=0 $Y2=0
cc_167 N_B2_M1007_g N_VGND_c_588_n 0.00383152f $X=1.855 $Y=0.69 $X2=0 $Y2=0
cc_168 N_B2_M1007_g N_VGND_c_590_n 0.00369533f $X=1.855 $Y=0.69 $X2=0 $Y2=0
cc_169 N_B2_M1007_g N_VGND_c_592_n 0.0101986f $X=1.855 $Y=0.69 $X2=0 $Y2=0
cc_170 N_B1_c_209_n N_A1_c_249_n 0.00933156f $X=2.385 $Y=1.285 $X2=0 $Y2=0
cc_171 N_B1_c_207_n A1 2.03024e-19 $X=2.207 $Y=1.79 $X2=0 $Y2=0
cc_172 N_B1_c_208_n A1 3.06869e-19 $X=2.385 $Y=1.285 $X2=0 $Y2=0
cc_173 N_B1_c_209_n A1 0.0331959f $X=2.385 $Y=1.285 $X2=0 $Y2=0
cc_174 N_B1_c_208_n N_A1_c_251_n 0.0101376f $X=2.385 $Y=1.285 $X2=0 $Y2=0
cc_175 N_B1_c_209_n N_A1_c_251_n 0.00134319f $X=2.385 $Y=1.285 $X2=0 $Y2=0
cc_176 N_B1_c_209_n N_A_32_74#_c_356_n 0.0434877f $X=2.385 $Y=1.285 $X2=0 $Y2=0
cc_177 N_B1_c_210_n N_A_32_74#_c_356_n 0.00961672f $X=2.345 $Y=1.12 $X2=0 $Y2=0
cc_178 N_B1_c_208_n N_A_32_74#_c_334_n 0.00162761f $X=2.385 $Y=1.285 $X2=0 $Y2=0
cc_179 N_B1_c_210_n N_A_32_74#_c_334_n 0.00978938f $X=2.345 $Y=1.12 $X2=0 $Y2=0
cc_180 N_B1_c_212_n N_A_27_390#_c_434_n 9.82651e-19 $X=2.207 $Y=1.875 $X2=0
+ $Y2=0
cc_181 N_B1_c_212_n N_A_27_390#_c_435_n 0.0142364f $X=2.207 $Y=1.875 $X2=0 $Y2=0
cc_182 N_B1_c_212_n N_A_27_390#_c_436_n 0.0081748f $X=2.207 $Y=1.875 $X2=0 $Y2=0
cc_183 N_B1_c_212_n N_A_337_390#_c_476_n 0.0200545f $X=2.207 $Y=1.875 $X2=0
+ $Y2=0
cc_184 N_B1_c_208_n N_A_337_390#_c_476_n 8.35191e-19 $X=2.385 $Y=1.285 $X2=0
+ $Y2=0
cc_185 N_B1_c_209_n N_A_337_390#_c_476_n 0.0419755f $X=2.385 $Y=1.285 $X2=0
+ $Y2=0
cc_186 N_B1_c_212_n N_A_337_390#_c_479_n 0.00986926f $X=2.207 $Y=1.875 $X2=0
+ $Y2=0
cc_187 N_B1_c_212_n N_VPWR_c_513_n 0.00171611f $X=2.207 $Y=1.875 $X2=0 $Y2=0
cc_188 N_B1_c_212_n N_VPWR_c_515_n 0.00390694f $X=2.207 $Y=1.875 $X2=0 $Y2=0
cc_189 N_B1_c_212_n N_VPWR_c_512_n 0.00542671f $X=2.207 $Y=1.875 $X2=0 $Y2=0
cc_190 N_B1_c_210_n N_VGND_c_588_n 0.00432706f $X=2.345 $Y=1.12 $X2=0 $Y2=0
cc_191 N_B1_c_210_n N_VGND_c_590_n 0.00438903f $X=2.345 $Y=1.12 $X2=0 $Y2=0
cc_192 N_B1_c_210_n N_VGND_c_592_n 0.00122056f $X=2.345 $Y=1.12 $X2=0 $Y2=0
cc_193 N_A1_c_249_n N_A2_c_287_n 0.00876246f $X=3.18 $Y=1.69 $X2=0 $Y2=0
cc_194 N_A1_c_255_n N_A2_c_287_n 0.00826139f $X=3.26 $Y=1.765 $X2=0 $Y2=0
cc_195 N_A1_c_254_n N_A2_c_292_n 0.00847822f $X=3.26 $Y=1.84 $X2=0 $Y2=0
cc_196 N_A1_c_249_n A2 5.72071e-19 $X=3.18 $Y=1.69 $X2=0 $Y2=0
cc_197 A1 A2 0.0253547f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_198 N_A1_c_251_n A2 0.00148118f $X=3.09 $Y=1.285 $X2=0 $Y2=0
cc_199 A1 N_A2_c_289_n 4.13361e-19 $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_200 N_A1_c_251_n N_A2_c_289_n 0.0324045f $X=3.09 $Y=1.285 $X2=0 $Y2=0
cc_201 N_A1_c_252_n N_A2_c_290_n 0.0324045f $X=3.09 $Y=1.12 $X2=0 $Y2=0
cc_202 N_A1_c_252_n N_A_32_74#_c_367_n 0.00806212f $X=3.09 $Y=1.12 $X2=0 $Y2=0
cc_203 A1 N_A_32_74#_c_334_n 0.023365f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_204 N_A1_c_251_n N_A_32_74#_c_334_n 0.00400401f $X=3.09 $Y=1.285 $X2=0 $Y2=0
cc_205 N_A1_c_252_n N_A_32_74#_c_334_n 0.00976723f $X=3.09 $Y=1.12 $X2=0 $Y2=0
cc_206 N_A1_c_254_n N_A_337_390#_c_476_n 0.0162531f $X=3.26 $Y=1.84 $X2=0 $Y2=0
cc_207 N_A1_c_255_n N_A_337_390#_c_476_n 0.00217f $X=3.26 $Y=1.765 $X2=0 $Y2=0
cc_208 A1 N_A_337_390#_c_476_n 0.0114382f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_209 N_A1_c_251_n N_A_337_390#_c_476_n 9.0515e-19 $X=3.09 $Y=1.285 $X2=0 $Y2=0
cc_210 N_A1_c_254_n N_A_337_390#_c_477_n 0.0039201f $X=3.26 $Y=1.84 $X2=0 $Y2=0
cc_211 N_A1_c_255_n N_A_337_390#_c_477_n 6.99035e-19 $X=3.26 $Y=1.765 $X2=0
+ $Y2=0
cc_212 N_A1_c_254_n N_A_337_390#_c_478_n 0.0139037f $X=3.26 $Y=1.84 $X2=0 $Y2=0
cc_213 N_A1_c_254_n N_VPWR_c_513_n 0.0172277f $X=3.26 $Y=1.84 $X2=0 $Y2=0
cc_214 N_A1_c_254_n N_VPWR_c_517_n 0.00530811f $X=3.26 $Y=1.84 $X2=0 $Y2=0
cc_215 N_A1_c_254_n N_VPWR_c_512_n 0.005315f $X=3.26 $Y=1.84 $X2=0 $Y2=0
cc_216 N_A1_c_252_n N_VGND_c_588_n 0.00557855f $X=3.09 $Y=1.12 $X2=0 $Y2=0
cc_217 N_A1_c_252_n N_VGND_c_590_n 0.00438903f $X=3.09 $Y=1.12 $X2=0 $Y2=0
cc_218 N_A2_c_287_n N_A_32_74#_c_328_n 0.0145442f $X=3.71 $Y=1.75 $X2=0 $Y2=0
cc_219 N_A2_c_292_n N_A_32_74#_c_328_n 0.0248102f $X=3.71 $Y=1.84 $X2=0 $Y2=0
cc_220 A2 N_A_32_74#_c_328_n 4.88188e-19 $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_221 N_A2_c_289_n N_A_32_74#_c_328_n 0.00945972f $X=3.66 $Y=1.285 $X2=0 $Y2=0
cc_222 N_A2_c_289_n N_A_32_74#_M1000_g 0.00426644f $X=3.66 $Y=1.285 $X2=0 $Y2=0
cc_223 N_A2_c_290_n N_A_32_74#_M1000_g 0.0133207f $X=3.66 $Y=1.12 $X2=0 $Y2=0
cc_224 A2 N_A_32_74#_c_367_n 0.0228539f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_225 N_A2_c_289_n N_A_32_74#_c_367_n 0.00452134f $X=3.66 $Y=1.285 $X2=0 $Y2=0
cc_226 N_A2_c_290_n N_A_32_74#_c_367_n 0.012296f $X=3.66 $Y=1.12 $X2=0 $Y2=0
cc_227 A2 N_A_32_74#_c_332_n 0.0124561f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_228 N_A2_c_289_n N_A_32_74#_c_332_n 6.3503e-19 $X=3.66 $Y=1.285 $X2=0 $Y2=0
cc_229 N_A2_c_290_n N_A_32_74#_c_332_n 0.00310754f $X=3.66 $Y=1.12 $X2=0 $Y2=0
cc_230 N_A2_c_290_n N_A_32_74#_c_334_n 0.00162108f $X=3.66 $Y=1.12 $X2=0 $Y2=0
cc_231 N_A2_c_287_n N_A_32_74#_c_335_n 0.00221602f $X=3.71 $Y=1.75 $X2=0 $Y2=0
cc_232 A2 N_A_32_74#_c_335_n 0.0183844f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_233 N_A2_c_289_n N_A_32_74#_c_335_n 5.13863e-19 $X=3.66 $Y=1.285 $X2=0 $Y2=0
cc_234 N_A2_c_292_n N_A_337_390#_c_477_n 0.00355712f $X=3.71 $Y=1.84 $X2=0 $Y2=0
cc_235 A2 N_A_337_390#_c_477_n 0.00879649f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_236 N_A2_c_289_n N_A_337_390#_c_477_n 7.51809e-19 $X=3.66 $Y=1.285 $X2=0
+ $Y2=0
cc_237 N_A2_c_292_n N_A_337_390#_c_478_n 0.00882327f $X=3.71 $Y=1.84 $X2=0 $Y2=0
cc_238 N_A2_c_292_n N_VPWR_c_514_n 0.0131787f $X=3.71 $Y=1.84 $X2=0 $Y2=0
cc_239 N_A2_c_292_n N_VPWR_c_517_n 0.00530811f $X=3.71 $Y=1.84 $X2=0 $Y2=0
cc_240 N_A2_c_292_n N_VPWR_c_512_n 0.005315f $X=3.71 $Y=1.84 $X2=0 $Y2=0
cc_241 N_A2_c_292_n X 5.37073e-19 $X=3.71 $Y=1.84 $X2=0 $Y2=0
cc_242 N_A2_c_290_n N_VGND_c_588_n 0.0178758f $X=3.66 $Y=1.12 $X2=0 $Y2=0
cc_243 N_A2_c_290_n N_VGND_c_590_n 0.00371083f $X=3.66 $Y=1.12 $X2=0 $Y2=0
cc_244 N_A_32_74#_c_337_n N_A_27_390#_c_431_n 0.0415813f $X=0.885 $Y=2.095 $X2=0
+ $Y2=0
cc_245 N_A_32_74#_M1009_d N_A_27_390#_c_432_n 0.00616839f $X=0.58 $Y=1.95 $X2=0
+ $Y2=0
cc_246 N_A_32_74#_c_337_n N_A_27_390#_c_432_n 0.0205214f $X=0.885 $Y=2.095 $X2=0
+ $Y2=0
cc_247 N_A_32_74#_c_337_n N_A_27_390#_c_434_n 0.0309585f $X=0.885 $Y=2.095 $X2=0
+ $Y2=0
cc_248 N_A_32_74#_c_328_n N_VPWR_c_514_n 0.0139217f $X=4.295 $Y=1.765 $X2=0
+ $Y2=0
cc_249 N_A_32_74#_c_335_n N_VPWR_c_514_n 0.0093499f $X=4.205 $Y=1.465 $X2=0
+ $Y2=0
cc_250 N_A_32_74#_c_328_n N_VPWR_c_518_n 0.00445602f $X=4.295 $Y=1.765 $X2=0
+ $Y2=0
cc_251 N_A_32_74#_c_328_n N_VPWR_c_512_n 0.00865213f $X=4.295 $Y=1.765 $X2=0
+ $Y2=0
cc_252 N_A_32_74#_M1000_g N_X_c_560_n 0.0138767f $X=4.305 $Y=0.74 $X2=0 $Y2=0
cc_253 N_A_32_74#_c_332_n N_X_c_560_n 0.00750685f $X=4.1 $Y=1.3 $X2=0 $Y2=0
cc_254 N_A_32_74#_c_328_n N_X_c_561_n 2.30445e-19 $X=4.295 $Y=1.765 $X2=0 $Y2=0
cc_255 N_A_32_74#_M1000_g N_X_c_561_n 0.00297544f $X=4.305 $Y=0.74 $X2=0 $Y2=0
cc_256 N_A_32_74#_c_335_n N_X_c_561_n 0.00111755f $X=4.205 $Y=1.465 $X2=0 $Y2=0
cc_257 N_A_32_74#_c_328_n X 0.00390015f $X=4.295 $Y=1.765 $X2=0 $Y2=0
cc_258 N_A_32_74#_c_335_n X 0.00102175f $X=4.205 $Y=1.465 $X2=0 $Y2=0
cc_259 N_A_32_74#_c_328_n X 0.0110443f $X=4.295 $Y=1.765 $X2=0 $Y2=0
cc_260 N_A_32_74#_c_328_n N_X_c_562_n 0.0125762f $X=4.295 $Y=1.765 $X2=0 $Y2=0
cc_261 N_A_32_74#_M1000_g N_X_c_562_n 0.00255192f $X=4.305 $Y=0.74 $X2=0 $Y2=0
cc_262 N_A_32_74#_c_332_n N_X_c_562_n 0.00541114f $X=4.1 $Y=1.3 $X2=0 $Y2=0
cc_263 N_A_32_74#_c_335_n N_X_c_562_n 0.0249107f $X=4.205 $Y=1.465 $X2=0 $Y2=0
cc_264 N_A_32_74#_c_340_n A_119_74# 0.00383368f $X=0.72 $Y=0.865 $X2=-0.19
+ $Y2=-0.245
cc_265 N_A_32_74#_c_351_n A_119_74# 0.00130602f $X=0.805 $Y=0.865 $X2=-0.19
+ $Y2=-0.245
cc_266 N_A_32_74#_c_333_n A_119_74# 6.66187e-19 $X=0.885 $Y=1.93 $X2=-0.19
+ $Y2=-0.245
cc_267 N_A_32_74#_c_356_n N_VGND_M1013_d 0.0224135f $X=2.295 $Y=0.64 $X2=-0.19
+ $Y2=-0.245
cc_268 N_A_32_74#_c_367_n N_VGND_M1001_d 0.0163508f $X=4.015 $Y=0.865 $X2=0
+ $Y2=0
cc_269 N_A_32_74#_c_332_n N_VGND_M1001_d 0.00355979f $X=4.1 $Y=1.3 $X2=0 $Y2=0
cc_270 N_A_32_74#_c_328_n N_VGND_c_588_n 4.00439e-19 $X=4.295 $Y=1.765 $X2=0
+ $Y2=0
cc_271 N_A_32_74#_M1000_g N_VGND_c_588_n 0.00583725f $X=4.305 $Y=0.74 $X2=0
+ $Y2=0
cc_272 N_A_32_74#_c_367_n N_VGND_c_588_n 0.0401368f $X=4.015 $Y=0.865 $X2=0
+ $Y2=0
cc_273 N_A_32_74#_c_334_n N_VGND_c_588_n 0.0496465f $X=3.13 $Y=0.64 $X2=0 $Y2=0
cc_274 N_A_32_74#_M1000_g N_VGND_c_589_n 0.00434272f $X=4.305 $Y=0.74 $X2=0
+ $Y2=0
cc_275 N_A_32_74#_M1000_g N_VGND_c_590_n 0.00826002f $X=4.305 $Y=0.74 $X2=0
+ $Y2=0
cc_276 N_A_32_74#_c_330_n N_VGND_c_590_n 0.0119472f $X=0.305 $Y=0.515 $X2=0
+ $Y2=0
cc_277 N_A_32_74#_c_340_n N_VGND_c_590_n 0.0081717f $X=0.72 $Y=0.865 $X2=0 $Y2=0
cc_278 N_A_32_74#_c_367_n N_VGND_c_590_n 0.0180838f $X=4.015 $Y=0.865 $X2=0
+ $Y2=0
cc_279 N_A_32_74#_c_351_n N_VGND_c_590_n 0.00663982f $X=0.805 $Y=0.865 $X2=0
+ $Y2=0
cc_280 N_A_32_74#_c_356_n N_VGND_c_590_n 0.0210815f $X=2.295 $Y=0.64 $X2=0 $Y2=0
cc_281 N_A_32_74#_c_334_n N_VGND_c_590_n 0.0308511f $X=3.13 $Y=0.64 $X2=0 $Y2=0
cc_282 N_A_32_74#_c_330_n N_VGND_c_591_n 0.0144324f $X=0.305 $Y=0.515 $X2=0
+ $Y2=0
cc_283 N_A_32_74#_c_330_n N_VGND_c_592_n 0.00836615f $X=0.305 $Y=0.515 $X2=0
+ $Y2=0
cc_284 N_A_32_74#_c_356_n N_VGND_c_592_n 0.0545917f $X=2.295 $Y=0.64 $X2=0 $Y2=0
cc_285 N_A_32_74#_c_334_n N_VGND_c_592_n 0.00952048f $X=3.13 $Y=0.64 $X2=0 $Y2=0
cc_286 N_A_32_74#_c_356_n A_386_74# 0.0072096f $X=2.295 $Y=0.64 $X2=-0.19
+ $Y2=-0.245
cc_287 N_A_32_74#_c_367_n A_651_74# 0.0072096f $X=4.015 $Y=0.865 $X2=-0.19
+ $Y2=-0.245
cc_288 N_A_27_390#_c_435_n N_A_337_390#_M1012_d 0.0041451f $X=2.26 $Y=2.99
+ $X2=-0.19 $Y2=1.66
cc_289 N_A_27_390#_M1002_d N_A_337_390#_c_476_n 0.00587162f $X=2.275 $Y=1.95
+ $X2=0 $Y2=0
cc_290 N_A_27_390#_c_436_n N_A_337_390#_c_476_n 0.0219924f $X=2.425 $Y=2.465
+ $X2=0 $Y2=0
cc_291 N_A_27_390#_c_434_n N_A_337_390#_c_479_n 0.00833463f $X=1.385 $Y=2.095
+ $X2=0 $Y2=0
cc_292 N_A_27_390#_c_435_n N_A_337_390#_c_479_n 0.0233667f $X=2.26 $Y=2.99 $X2=0
+ $Y2=0
cc_293 N_A_27_390#_c_436_n N_A_337_390#_c_479_n 0.0287017f $X=2.425 $Y=2.465
+ $X2=0 $Y2=0
cc_294 N_A_27_390#_c_435_n N_VPWR_c_513_n 0.0121618f $X=2.26 $Y=2.99 $X2=0 $Y2=0
cc_295 N_A_27_390#_c_436_n N_VPWR_c_513_n 0.0407548f $X=2.425 $Y=2.465 $X2=0
+ $Y2=0
cc_296 N_A_27_390#_c_432_n N_VPWR_c_515_n 0.0490392f $X=1.22 $Y=2.99 $X2=0 $Y2=0
cc_297 N_A_27_390#_c_433_n N_VPWR_c_515_n 0.0236039f $X=0.445 $Y=2.99 $X2=0
+ $Y2=0
cc_298 N_A_27_390#_c_435_n N_VPWR_c_515_n 0.0685025f $X=2.26 $Y=2.99 $X2=0 $Y2=0
cc_299 N_A_27_390#_c_437_n N_VPWR_c_515_n 0.0236039f $X=1.385 $Y=2.99 $X2=0
+ $Y2=0
cc_300 N_A_27_390#_c_432_n N_VPWR_c_512_n 0.0289696f $X=1.22 $Y=2.99 $X2=0 $Y2=0
cc_301 N_A_27_390#_c_433_n N_VPWR_c_512_n 0.0128208f $X=0.445 $Y=2.99 $X2=0
+ $Y2=0
cc_302 N_A_27_390#_c_435_n N_VPWR_c_512_n 0.0393555f $X=2.26 $Y=2.99 $X2=0 $Y2=0
cc_303 N_A_27_390#_c_437_n N_VPWR_c_512_n 0.0128208f $X=1.385 $Y=2.99 $X2=0
+ $Y2=0
cc_304 N_A_337_390#_c_476_n N_VPWR_M1003_s 0.010717f $X=3.32 $Y=2.045 $X2=-0.19
+ $Y2=1.66
cc_305 N_A_337_390#_c_476_n N_VPWR_c_513_n 0.025036f $X=3.32 $Y=2.045 $X2=0
+ $Y2=0
cc_306 N_A_337_390#_c_478_n N_VPWR_c_513_n 0.0246172f $X=3.485 $Y=2.77 $X2=0
+ $Y2=0
cc_307 N_A_337_390#_c_477_n N_VPWR_c_514_n 0.0165339f $X=3.485 $Y=2.13 $X2=0
+ $Y2=0
cc_308 N_A_337_390#_c_478_n N_VPWR_c_514_n 0.0541034f $X=3.485 $Y=2.77 $X2=0
+ $Y2=0
cc_309 N_A_337_390#_c_478_n N_VPWR_c_517_n 0.0123111f $X=3.485 $Y=2.77 $X2=0
+ $Y2=0
cc_310 N_A_337_390#_c_478_n N_VPWR_c_512_n 0.0117546f $X=3.485 $Y=2.77 $X2=0
+ $Y2=0
cc_311 N_VPWR_c_514_n X 0.0419219f $X=4.02 $Y=2.06 $X2=0 $Y2=0
cc_312 N_VPWR_c_518_n X 0.0157093f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_313 N_VPWR_c_512_n X 0.0129699f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_314 N_X_c_560_n N_VGND_c_588_n 0.0107229f $X=4.52 $Y=0.515 $X2=0 $Y2=0
cc_315 N_X_c_560_n N_VGND_c_589_n 0.0156794f $X=4.52 $Y=0.515 $X2=0 $Y2=0
cc_316 N_X_c_560_n N_VGND_c_590_n 0.0129217f $X=4.52 $Y=0.515 $X2=0 $Y2=0
